* NGSPICE file created from opamp114.ext - technology: sky130A

.subckt opamp114 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 a_n2140_13878.t20 a_n2318_13878.t24 a_n2318_13878.t25 vdd.t228 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X1 CSoutput.t111 a_n7636_8799.t32 vdd.t240 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X2 a_n2140_13878.t4 a_n2318_13878.t48 vdd.t239 vdd.t238 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 vdd.t179 a_n7636_8799.t33 CSoutput.t110 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X4 gnd.t238 gnd.t235 gnd.t237 gnd.t236 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X5 commonsourceibias.t47 commonsourceibias.t46 gnd.t82 gnd.t78 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X6 gnd.t257 commonsourceibias.t48 CSoutput.t136 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 gnd.t234 gnd.t232 gnd.t233 gnd.t220 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X8 a_n7636_8799.t5 plus.t5 a_n2903_n3924.t35 gnd.t109 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X9 output.t19 outputibias.t8 gnd.t261 gnd.t260 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X10 output.t15 CSoutput.t144 vdd.t117 gnd.t25 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X11 CSoutput.t109 a_n7636_8799.t34 vdd.t94 vdd.t93 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X12 gnd.t58 commonsourceibias.t49 CSoutput.t14 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X13 minus.t4 gnd.t229 gnd.t231 gnd.t230 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X14 gnd.t114 commonsourceibias.t44 commonsourceibias.t45 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X15 vdd.t92 vdd.t90 vdd.t91 vdd.t51 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X16 a_n2318_8322.t27 a_n2318_13878.t49 a_n7636_8799.t12 vdd.t237 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X17 gnd.t77 commonsourceibias.t50 CSoutput.t116 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X18 outputibias.t7 outputibias.t6 gnd.t56 gnd.t55 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X19 output.t14 CSoutput.t145 vdd.t118 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X20 CSoutput.t108 a_n7636_8799.t35 vdd.t154 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X21 vdd.t159 a_n7636_8799.t36 CSoutput.t107 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X22 a_n7636_8799.t17 a_n2318_13878.t50 a_n2318_8322.t26 vdd.t226 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X23 a_n2318_13878.t46 minus.t5 a_n2903_n3924.t18 gnd.t106 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X24 a_n7636_8799.t22 plus.t6 a_n2903_n3924.t34 gnd.t125 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X25 gnd.t7 commonsourceibias.t42 commonsourceibias.t43 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X26 CSoutput.t106 a_n7636_8799.t37 vdd.t107 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X27 vdd.t263 a_n7636_8799.t38 CSoutput.t105 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X28 a_n2318_13878.t47 minus.t6 a_n2903_n3924.t19 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X29 vdd.t104 a_n7636_8799.t39 CSoutput.t104 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X30 a_n7636_8799.t8 a_n2318_13878.t51 a_n2318_8322.t25 vdd.t193 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X31 CSoutput.t118 commonsourceibias.t51 gnd.t81 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 CSoutput.t146 a_n2318_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X33 gnd.t86 commonsourceibias.t40 commonsourceibias.t41 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X34 vdd.t89 vdd.t87 vdd.t88 vdd.t18 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X35 CSoutput.t103 a_n7636_8799.t40 vdd.t181 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X36 a_n2903_n3924.t33 plus.t7 a_n7636_8799.t2 gnd.t105 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X37 vdd.t174 CSoutput.t147 output.t13 gnd.t23 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X38 vdd.t175 CSoutput.t148 output.t12 gnd.t22 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X39 CSoutput.t102 a_n7636_8799.t41 vdd.t170 vdd.t169 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X40 a_n2903_n3924.t17 minus.t7 a_n2318_13878.t45 gnd.t250 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X41 CSoutput.t126 commonsourceibias.t52 gnd.t123 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X42 a_n2903_n3924.t3 diffpairibias.t16 gnd.t120 gnd.t119 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X43 CSoutput.t101 a_n7636_8799.t42 vdd.t262 vdd.t93 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X44 CSoutput.t131 commonsourceibias.t53 gnd.t130 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X45 a_n2140_13878.t19 a_n2318_13878.t10 a_n2318_13878.t11 vdd.t201 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X46 a_n2318_13878.t31 a_n2318_13878.t30 a_n2140_13878.t18 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X47 vdd.t86 vdd.t84 vdd.t85 vdd.t51 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X48 CSoutput.t132 commonsourceibias.t54 gnd.t240 gnd.t78 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X49 CSoutput.t100 a_n7636_8799.t43 vdd.t116 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X50 gnd.t228 gnd.t226 plus.t4 gnd.t227 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X51 vdd.t83 vdd.t81 vdd.t82 vdd.t64 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X52 vdd.t180 a_n7636_8799.t44 CSoutput.t99 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X53 a_n2903_n3924.t32 plus.t8 a_n7636_8799.t24 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X54 diffpairibias.t15 diffpairibias.t14 gnd.t65 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X55 gnd.t225 gnd.t223 gnd.t224 gnd.t220 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X56 a_n7636_8799.t10 a_n2318_13878.t52 a_n2318_8322.t24 vdd.t219 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X57 vdd.t1 a_n7636_8799.t45 CSoutput.t98 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X58 vdd.t264 a_n7636_8799.t46 CSoutput.t97 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X59 CSoutput.t96 a_n7636_8799.t47 vdd.t5 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X60 gnd.t129 commonsourceibias.t55 CSoutput.t130 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X61 gnd.t3 commonsourceibias.t56 CSoutput.t1 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X62 diffpairibias.t13 diffpairibias.t12 gnd.t99 gnd.t98 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X63 CSoutput.t95 a_n7636_8799.t48 vdd.t106 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X64 output.t11 CSoutput.t149 vdd.t176 gnd.t21 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X65 gnd.t128 commonsourceibias.t57 CSoutput.t129 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X66 commonsourceibias.t39 commonsourceibias.t38 gnd.t85 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X67 vdd.t144 CSoutput.t150 output.t10 gnd.t20 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X68 CSoutput.t94 a_n7636_8799.t49 vdd.t156 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X69 vdd.t261 a_n7636_8799.t50 CSoutput.t93 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X70 CSoutput.t92 a_n7636_8799.t51 vdd.t244 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X71 CSoutput.t91 a_n7636_8799.t52 vdd.t3 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X72 CSoutput.t90 a_n7636_8799.t53 vdd.t243 vdd.t169 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X73 a_n2903_n3924.t16 minus.t8 a_n2318_13878.t44 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X74 a_n2903_n3924.t31 plus.t9 a_n7636_8799.t23 gnd.t239 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X75 gnd.t243 commonsourceibias.t58 CSoutput.t134 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X76 commonsourceibias.t37 commonsourceibias.t36 gnd.t111 gnd.t72 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X77 vdd.t10 a_n7636_8799.t54 CSoutput.t89 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X78 a_n2903_n3924.t39 diffpairibias.t17 gnd.t277 gnd.t276 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X79 gnd.t68 commonsourceibias.t34 commonsourceibias.t35 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 vdd.t16 a_n7636_8799.t55 CSoutput.t88 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X81 vdd.t257 a_n7636_8799.t56 CSoutput.t87 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X82 a_n7636_8799.t19 a_n2318_13878.t53 a_n2318_8322.t23 vdd.t227 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X83 a_n2318_13878.t3 a_n2318_13878.t2 a_n2140_13878.t17 vdd.t237 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X84 a_n2903_n3924.t30 plus.t10 a_n7636_8799.t4 gnd.t108 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X85 a_n2318_13878.t17 a_n2318_13878.t16 a_n2140_13878.t16 vdd.t196 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X86 gnd.t281 commonsourceibias.t32 commonsourceibias.t33 gnd.t93 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X87 commonsourceibias.t31 commonsourceibias.t30 gnd.t127 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 outputibias.t5 outputibias.t4 gnd.t50 gnd.t49 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X89 CSoutput.t86 a_n7636_8799.t57 vdd.t256 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X90 vdd.t266 a_n7636_8799.t58 CSoutput.t85 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X91 CSoutput.t12 commonsourceibias.t59 gnd.t48 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X92 vdd.t145 CSoutput.t151 output.t9 gnd.t19 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X93 vdd.t80 vdd.t78 vdd.t79 vdd.t30 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X94 CSoutput.t84 a_n7636_8799.t59 vdd.t265 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X95 vdd.t77 vdd.t75 vdd.t76 vdd.t68 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X96 CSoutput.t6 commonsourceibias.t60 gnd.t33 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X97 vdd.t74 vdd.t71 vdd.t73 vdd.t72 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X98 gnd.t258 commonsourceibias.t61 CSoutput.t137 gnd.t93 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X99 gnd.t222 gnd.t219 gnd.t221 gnd.t220 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X100 commonsourceibias.t29 commonsourceibias.t28 gnd.t110 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X101 CSoutput.t117 commonsourceibias.t62 gnd.t79 gnd.t78 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X102 CSoutput.t152 a_n2318_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X103 outputibias.t3 outputibias.t2 gnd.t256 gnd.t255 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X104 a_n2318_8322.t11 a_n2318_13878.t54 vdd.t236 vdd.t235 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X105 vdd.t234 a_n2318_13878.t55 a_n2318_8322.t10 vdd.t233 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X106 a_n2318_13878.t7 a_n2318_13878.t6 a_n2140_13878.t15 vdd.t203 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X107 gnd.t218 gnd.t216 minus.t3 gnd.t217 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X108 CSoutput.t83 a_n7636_8799.t60 vdd.t191 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X109 CSoutput.t82 a_n7636_8799.t61 vdd.t182 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X110 a_n2903_n3924.t2 diffpairibias.t18 gnd.t102 gnd.t101 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X111 gnd.t215 gnd.t213 gnd.t214 gnd.t161 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X112 commonsourceibias.t27 commonsourceibias.t26 gnd.t40 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X113 vdd.t232 a_n2318_13878.t56 a_n2140_13878.t0 vdd.t231 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X114 vdd.t70 vdd.t67 vdd.t69 vdd.t68 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X115 vdd.t241 a_n7636_8799.t62 CSoutput.t81 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X116 gnd.t268 commonsourceibias.t24 commonsourceibias.t25 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X117 gnd.t75 commonsourceibias.t63 CSoutput.t115 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X118 a_n7636_8799.t18 a_n2318_13878.t57 a_n2318_8322.t22 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X119 a_n2318_8322.t9 a_n2318_13878.t58 vdd.t230 vdd.t229 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X120 vdd.t66 vdd.t63 vdd.t65 vdd.t64 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X121 gnd.t52 commonsourceibias.t64 CSoutput.t13 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X122 a_n7636_8799.t25 plus.t11 a_n2903_n3924.t29 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X123 gnd.t61 commonsourceibias.t65 CSoutput.t15 gnd.t60 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X124 vdd.t245 a_n7636_8799.t63 CSoutput.t80 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X125 vdd.t95 a_n7636_8799.t64 CSoutput.t79 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X126 a_n2318_13878.t23 a_n2318_13878.t22 a_n2140_13878.t14 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X127 CSoutput.t78 a_n7636_8799.t65 vdd.t157 vdd.t123 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X128 a_n7636_8799.t30 plus.t12 a_n2903_n3924.t28 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X129 diffpairibias.t11 diffpairibias.t10 gnd.t104 gnd.t103 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X130 CSoutput.t77 a_n7636_8799.t66 vdd.t177 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X131 a_n7636_8799.t20 a_n2318_13878.t59 a_n2318_8322.t21 vdd.t228 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X132 gnd.t89 commonsourceibias.t66 CSoutput.t120 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X133 a_n2140_13878.t13 a_n2318_13878.t12 a_n2318_13878.t13 vdd.t227 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X134 gnd.t212 gnd.t210 gnd.t211 gnd.t139 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X135 outputibias.t1 outputibias.t0 gnd.t54 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X136 vdd.t62 vdd.t60 vdd.t61 vdd.t30 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X137 gnd.t74 commonsourceibias.t67 CSoutput.t114 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X138 CSoutput.t153 a_n2318_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X139 a_n2140_13878.t12 a_n2318_13878.t18 a_n2318_13878.t19 vdd.t226 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X140 CSoutput.t76 a_n7636_8799.t67 vdd.t267 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X141 vdd.t225 a_n2318_13878.t60 a_n2318_8322.t8 vdd.t224 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X142 CSoutput.t139 commonsourceibias.t68 gnd.t266 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X143 CSoutput.t154 a_n2318_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X144 a_n2318_13878.t21 a_n2318_13878.t20 a_n2140_13878.t11 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X145 vdd.t190 a_n7636_8799.t68 CSoutput.t75 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X146 a_n2903_n3924.t27 plus.t13 a_n7636_8799.t1 gnd.t76 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X147 a_n2318_13878.t43 minus.t9 a_n2903_n3924.t15 gnd.t109 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X148 plus.t3 gnd.t207 gnd.t209 gnd.t208 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X149 vdd.t158 a_n7636_8799.t69 CSoutput.t74 vdd.t133 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X150 gnd.t206 gnd.t204 minus.t2 gnd.t205 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X151 gnd.t203 gnd.t200 gnd.t202 gnd.t201 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X152 a_n2903_n3924.t0 diffpairibias.t19 gnd.t91 gnd.t90 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X153 CSoutput.t135 commonsourceibias.t69 gnd.t244 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X154 a_n7636_8799.t27 plus.t14 a_n2903_n3924.t26 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X155 CSoutput.t112 commonsourceibias.t70 gnd.t70 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X156 a_n2903_n3924.t36 diffpairibias.t20 gnd.t265 gnd.t264 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X157 vdd.t122 CSoutput.t155 output.t8 gnd.t18 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X158 vdd.t167 a_n7636_8799.t70 CSoutput.t73 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X159 vdd.t168 a_n7636_8799.t71 CSoutput.t72 vdd.t161 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X160 gnd.t94 commonsourceibias.t71 CSoutput.t122 gnd.t93 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X161 CSoutput.t9 commonsourceibias.t72 gnd.t39 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X162 a_n7636_8799.t26 plus.t15 a_n2903_n3924.t25 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X163 CSoutput.t71 a_n7636_8799.t72 vdd.t120 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X164 CSoutput.t70 a_n7636_8799.t73 vdd.t121 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X165 CSoutput.t69 a_n7636_8799.t74 vdd.t147 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X166 a_n2140_13878.t22 a_n2318_13878.t61 vdd.t223 vdd.t222 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X167 gnd.t199 gnd.t197 gnd.t198 gnd.t157 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X168 diffpairibias.t9 diffpairibias.t8 gnd.t63 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X169 vdd.t59 vdd.t57 vdd.t58 vdd.t47 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X170 vdd.t221 a_n2318_13878.t62 a_n2140_13878.t21 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X171 a_n2318_13878.t36 minus.t10 a_n2903_n3924.t8 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X172 vdd.t149 a_n7636_8799.t75 CSoutput.t68 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X173 CSoutput.t67 a_n7636_8799.t76 vdd.t165 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X174 a_n2903_n3924.t24 plus.t16 a_n7636_8799.t31 gnd.t250 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X175 vdd.t56 vdd.t54 vdd.t55 vdd.t47 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X176 CSoutput.t138 commonsourceibias.t73 gnd.t263 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X177 gnd.t282 commonsourceibias.t74 CSoutput.t143 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X178 a_n2140_13878.t10 a_n2318_13878.t0 a_n2318_13878.t1 vdd.t219 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X179 gnd.t87 commonsourceibias.t22 commonsourceibias.t23 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X180 gnd.t95 commonsourceibias.t75 CSoutput.t123 gnd.t60 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X181 vdd.t166 a_n7636_8799.t77 CSoutput.t66 vdd.t133 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X182 a_n2318_8322.t20 a_n2318_13878.t63 a_n7636_8799.t6 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X183 gnd.t92 commonsourceibias.t76 CSoutput.t121 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X184 a_n2903_n3924.t7 minus.t11 a_n2318_13878.t35 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X185 vdd.t141 a_n7636_8799.t78 CSoutput.t65 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X186 CSoutput.t64 a_n7636_8799.t79 vdd.t142 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X187 diffpairibias.t7 diffpairibias.t6 gnd.t279 gnd.t278 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X188 vdd.t160 a_n7636_8799.t80 CSoutput.t63 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X189 vdd.t162 a_n7636_8799.t81 CSoutput.t62 vdd.t161 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X190 vdd.t218 a_n2318_13878.t64 a_n2318_8322.t7 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X191 gnd.t267 commonsourceibias.t20 commonsourceibias.t21 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X192 gnd.t196 gnd.t194 minus.t1 gnd.t195 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X193 plus.t2 gnd.t191 gnd.t193 gnd.t192 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X194 CSoutput.t142 commonsourceibias.t77 gnd.t273 gnd.t72 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X195 gnd.t190 gnd.t188 gnd.t189 gnd.t157 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X196 gnd.t187 gnd.t185 gnd.t186 gnd.t143 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X197 CSoutput.t141 commonsourceibias.t78 gnd.t272 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X198 a_n2140_13878.t3 a_n2318_13878.t65 vdd.t216 vdd.t215 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X199 vdd.t114 a_n7636_8799.t82 CSoutput.t61 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X200 CSoutput.t60 a_n7636_8799.t83 vdd.t115 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X201 CSoutput.t59 a_n7636_8799.t84 vdd.t7 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X202 gnd.t26 commonsourceibias.t18 commonsourceibias.t19 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X203 vdd.t53 vdd.t50 vdd.t52 vdd.t51 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X204 gnd.t184 gnd.t181 gnd.t183 gnd.t182 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X205 a_n2318_8322.t19 a_n2318_13878.t66 a_n7636_8799.t15 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X206 vdd.t213 a_n2318_13878.t67 a_n2318_8322.t6 vdd.t212 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X207 vdd.t49 vdd.t46 vdd.t48 vdd.t47 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X208 CSoutput.t58 a_n7636_8799.t85 vdd.t8 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X209 CSoutput.t119 commonsourceibias.t79 gnd.t84 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X210 a_n2903_n3924.t37 diffpairibias.t21 gnd.t270 gnd.t269 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X211 output.t7 CSoutput.t156 vdd.t253 gnd.t17 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X212 CSoutput.t57 a_n7636_8799.t86 vdd.t135 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X213 vdd.t137 a_n7636_8799.t87 CSoutput.t56 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X214 a_n7636_8799.t3 plus.t17 a_n2903_n3924.t23 gnd.t106 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X215 a_n2318_13878.t42 minus.t12 a_n2903_n3924.t14 gnd.t125 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X216 CSoutput.t125 commonsourceibias.t80 gnd.t107 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X217 vdd.t112 a_n7636_8799.t88 CSoutput.t55 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X218 vdd.t113 a_n7636_8799.t89 CSoutput.t54 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X219 a_n2903_n3924.t13 minus.t13 a_n2318_13878.t41 gnd.t239 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X220 CSoutput.t157 a_n2318_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X221 CSoutput.t128 commonsourceibias.t81 gnd.t126 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X222 vdd.t45 vdd.t43 vdd.t44 vdd.t26 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X223 gnd.t1 commonsourceibias.t82 CSoutput.t0 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X224 output.t18 outputibias.t9 gnd.t252 gnd.t251 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X225 output.t6 CSoutput.t158 vdd.t254 gnd.t16 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X226 vdd.t42 vdd.t39 vdd.t41 vdd.t40 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X227 vdd.t129 a_n7636_8799.t90 CSoutput.t53 vdd.t108 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X228 a_n2903_n3924.t12 minus.t14 a_n2318_13878.t40 gnd.t108 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X229 gnd.t180 gnd.t178 gnd.t179 gnd.t150 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X230 CSoutput.t52 a_n7636_8799.t91 vdd.t131 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X231 CSoutput.t51 a_n7636_8799.t92 vdd.t151 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X232 a_n2140_13878.t9 a_n2318_13878.t28 a_n2318_13878.t29 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X233 a_n2903_n3924.t11 minus.t15 a_n2318_13878.t39 gnd.t105 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X234 a_n2318_8322.t18 a_n2318_13878.t68 a_n7636_8799.t16 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X235 gnd.t177 gnd.t175 gnd.t176 gnd.t150 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X236 output.t17 outputibias.t10 gnd.t116 gnd.t115 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X237 diffpairibias.t5 diffpairibias.t4 gnd.t122 gnd.t121 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X238 CSoutput.t50 a_n7636_8799.t93 vdd.t153 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X239 CSoutput.t49 a_n7636_8799.t94 vdd.t124 vdd.t123 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X240 vdd.t125 a_n7636_8799.t95 CSoutput.t48 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X241 gnd.t124 commonsourceibias.t83 CSoutput.t127 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X242 CSoutput.t11 commonsourceibias.t84 gnd.t46 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X243 vdd.t101 a_n7636_8799.t96 CSoutput.t47 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X244 CSoutput.t46 a_n7636_8799.t97 vdd.t103 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X245 a_n2318_8322.t5 a_n2318_13878.t69 vdd.t210 vdd.t209 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X246 gnd.t44 commonsourceibias.t85 CSoutput.t10 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X247 gnd.t71 commonsourceibias.t16 commonsourceibias.t17 gnd.t60 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X248 output.t5 CSoutput.t159 vdd.t247 gnd.t15 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X249 vdd.t38 vdd.t36 vdd.t37 vdd.t22 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X250 a_n2903_n3924.t10 minus.t16 a_n2318_13878.t38 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X251 gnd.t174 gnd.t171 gnd.t173 gnd.t172 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X252 vdd.t208 a_n2318_13878.t70 a_n2140_13878.t1 vdd.t207 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X253 gnd.t170 gnd.t167 gnd.t169 gnd.t168 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X254 CSoutput.t45 a_n7636_8799.t98 vdd.t97 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X255 CSoutput.t44 a_n7636_8799.t99 vdd.t99 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X256 vdd.t12 a_n7636_8799.t100 CSoutput.t43 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X257 vdd.t14 a_n7636_8799.t101 CSoutput.t42 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X258 gnd.t166 gnd.t164 gnd.t165 gnd.t143 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X259 CSoutput.t113 commonsourceibias.t86 gnd.t73 gnd.t72 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X260 gnd.t163 gnd.t160 gnd.t162 gnd.t161 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X261 CSoutput.t4 commonsourceibias.t87 gnd.t30 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X262 gnd.t159 gnd.t156 gnd.t158 gnd.t157 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X263 vdd.t248 CSoutput.t160 output.t4 gnd.t14 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X264 vdd.t35 vdd.t33 vdd.t34 vdd.t26 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X265 gnd.t155 gnd.t153 plus.t1 gnd.t154 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X266 a_n7636_8799.t11 a_n2318_13878.t71 a_n2318_8322.t17 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X267 a_n2318_8322.t16 a_n2318_13878.t72 a_n7636_8799.t9 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X268 CSoutput.t41 a_n7636_8799.t102 vdd.t186 vdd.t169 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X269 a_n2140_13878.t2 a_n2318_13878.t73 vdd.t205 vdd.t204 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X270 vdd.t187 a_n7636_8799.t103 CSoutput.t40 vdd.t161 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X271 vdd.t184 a_n7636_8799.t104 CSoutput.t39 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X272 CSoutput.t38 a_n7636_8799.t105 vdd.t185 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 a_n2903_n3924.t22 plus.t18 a_n7636_8799.t29 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X274 output.t16 outputibias.t11 gnd.t118 gnd.t117 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X275 a_n2318_8322.t15 a_n2318_13878.t74 a_n7636_8799.t7 vdd.t203 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X276 a_n2318_13878.t37 minus.t17 a_n2903_n3924.t9 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X277 CSoutput.t140 commonsourceibias.t88 gnd.t271 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 CSoutput.t37 a_n7636_8799.t106 vdd.t132 vdd.t123 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X279 vdd.t134 a_n7636_8799.t107 CSoutput.t36 vdd.t133 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X280 vdd.t249 CSoutput.t161 output.t3 gnd.t13 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X281 CSoutput.t35 a_n7636_8799.t108 vdd.t127 vdd.t126 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X282 CSoutput.t34 a_n7636_8799.t109 vdd.t128 vdd.t126 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X283 a_n2140_13878.t8 a_n2318_13878.t26 a_n2318_13878.t27 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X284 commonsourceibias.t15 commonsourceibias.t14 gnd.t59 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X285 output.t2 CSoutput.t162 vdd.t250 gnd.t12 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X286 vdd.t258 a_n7636_8799.t110 CSoutput.t33 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X287 vdd.t32 vdd.t29 vdd.t31 vdd.t30 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X288 gnd.t35 commonsourceibias.t89 CSoutput.t7 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X289 vdd.t28 vdd.t25 vdd.t27 vdd.t26 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X290 gnd.t100 commonsourceibias.t90 CSoutput.t124 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X291 output.t1 CSoutput.t163 vdd.t251 gnd.t11 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X292 vdd.t259 a_n7636_8799.t111 CSoutput.t32 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X293 vdd.t109 a_n7636_8799.t112 CSoutput.t31 vdd.t108 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X294 gnd.t152 gnd.t149 gnd.t151 gnd.t150 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X295 a_n2903_n3924.t5 minus.t18 a_n2318_13878.t33 gnd.t76 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X296 a_n2903_n3924.t38 diffpairibias.t22 gnd.t275 gnd.t274 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X297 CSoutput.t30 a_n7636_8799.t113 vdd.t111 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X298 a_n7636_8799.t21 a_n2318_13878.t75 a_n2318_8322.t14 vdd.t201 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X299 a_n2318_13878.t5 a_n2318_13878.t4 a_n2140_13878.t7 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X300 gnd.t5 commonsourceibias.t91 CSoutput.t2 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X301 commonsourceibias.t13 commonsourceibias.t12 gnd.t80 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X302 CSoutput.t29 a_n7636_8799.t114 vdd.t260 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X303 vdd.t139 a_n7636_8799.t115 CSoutput.t28 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X304 vdd.t163 a_n7636_8799.t116 CSoutput.t27 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X305 CSoutput.t26 a_n7636_8799.t117 vdd.t171 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X306 vdd.t173 a_n7636_8799.t118 CSoutput.t25 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X307 minus.t0 gnd.t146 gnd.t148 gnd.t147 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X308 gnd.t137 gnd.t135 plus.t0 gnd.t136 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X309 diffpairibias.t3 diffpairibias.t2 gnd.t113 gnd.t112 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X310 a_n2318_8322.t13 a_n2318_13878.t76 a_n7636_8799.t14 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X311 a_n2318_13878.t32 minus.t19 a_n2903_n3924.t4 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X312 vdd.t255 a_n7636_8799.t119 CSoutput.t24 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X313 commonsourceibias.t11 commonsourceibias.t10 gnd.t28 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X314 gnd.t241 commonsourceibias.t92 CSoutput.t133 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X315 CSoutput.t164 a_n2318_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X316 diffpairibias.t1 diffpairibias.t0 gnd.t42 gnd.t41 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X317 CSoutput.t3 commonsourceibias.t93 gnd.t9 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X318 vdd.t252 CSoutput.t165 output.t0 gnd.t10 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X319 CSoutput.t23 a_n7636_8799.t120 vdd.t242 vdd.t126 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X320 vdd.t198 a_n2318_13878.t77 a_n2140_13878.t23 vdd.t197 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X321 vdd.t24 vdd.t21 vdd.t23 vdd.t22 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X322 vdd.t20 vdd.t17 vdd.t19 vdd.t18 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X323 vdd.t246 a_n7636_8799.t121 CSoutput.t22 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X324 gnd.t145 gnd.t142 gnd.t144 gnd.t143 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X325 CSoutput.t5 commonsourceibias.t94 gnd.t31 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X326 vdd.t178 a_n7636_8799.t122 CSoutput.t21 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X327 CSoutput.t20 a_n7636_8799.t123 vdd.t143 vdd.t93 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X328 commonsourceibias.t9 commonsourceibias.t8 gnd.t259 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X329 a_n7636_8799.t28 plus.t19 a_n2903_n3924.t21 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X330 a_n2318_8322.t12 a_n2318_13878.t78 a_n7636_8799.t13 vdd.t196 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X331 CSoutput.t8 commonsourceibias.t95 gnd.t37 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X332 a_n2318_13878.t34 minus.t20 a_n2903_n3924.t6 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X333 vdd.t189 a_n7636_8799.t124 CSoutput.t19 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X334 CSoutput.t18 a_n7636_8799.t125 vdd.t119 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X335 vdd.t155 a_n7636_8799.t126 CSoutput.t17 vdd.t108 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X336 gnd.t283 commonsourceibias.t6 commonsourceibias.t7 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X337 commonsourceibias.t5 commonsourceibias.t4 gnd.t254 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X338 a_n2318_8322.t4 a_n2318_13878.t79 vdd.t195 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X339 a_n2140_13878.t6 a_n2318_13878.t14 a_n2318_13878.t15 vdd.t193 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X340 gnd.t141 gnd.t138 gnd.t140 gnd.t139 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X341 vdd.t164 a_n7636_8799.t127 CSoutput.t16 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X342 a_n2903_n3924.t20 plus.t20 a_n7636_8799.t0 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X343 commonsourceibias.t3 commonsourceibias.t2 gnd.t262 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X344 a_n2318_13878.t9 a_n2318_13878.t8 a_n2140_13878.t5 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X345 gnd.t280 commonsourceibias.t0 commonsourceibias.t1 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X346 a_n2903_n3924.t1 diffpairibias.t23 gnd.t97 gnd.t96 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X347 gnd.t134 gnd.t131 gnd.t133 gnd.t132 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
R0 a_n2318_13878.n57 a_n2318_13878.t6 533.335
R1 a_n2318_13878.n112 a_n2318_13878.t0 512.366
R2 a_n2318_13878.n64 a_n2318_13878.t4 512.366
R3 a_n2318_13878.n111 a_n2318_13878.t28 512.366
R4 a_n2318_13878.n110 a_n2318_13878.t2 512.366
R5 a_n2318_13878.n65 a_n2318_13878.t26 512.366
R6 a_n2318_13878.n109 a_n2318_13878.t22 512.366
R7 a_n2318_13878.n51 a_n2318_13878.t78 533.335
R8 a_n2318_13878.n108 a_n2318_13878.t59 512.366
R9 a_n2318_13878.n74 a_n2318_13878.t63 512.366
R10 a_n2318_13878.n107 a_n2318_13878.t53 512.366
R11 a_n2318_13878.n106 a_n2318_13878.t68 512.366
R12 a_n2318_13878.n75 a_n2318_13878.t75 512.366
R13 a_n2318_13878.n105 a_n2318_13878.t76 512.366
R14 a_n2318_13878.n36 a_n2318_13878.t16 533.335
R15 a_n2318_13878.n86 a_n2318_13878.t24 512.366
R16 a_n2318_13878.n87 a_n2318_13878.t8 512.366
R17 a_n2318_13878.n88 a_n2318_13878.t12 512.366
R18 a_n2318_13878.n89 a_n2318_13878.t30 512.366
R19 a_n2318_13878.n79 a_n2318_13878.t10 512.366
R20 a_n2318_13878.n90 a_n2318_13878.t20 512.366
R21 a_n2318_13878.n29 a_n2318_13878.t74 533.335
R22 a_n2318_13878.n81 a_n2318_13878.t52 512.366
R23 a_n2318_13878.n82 a_n2318_13878.t72 512.366
R24 a_n2318_13878.n83 a_n2318_13878.t71 512.366
R25 a_n2318_13878.n84 a_n2318_13878.t49 512.366
R26 a_n2318_13878.n80 a_n2318_13878.t57 512.366
R27 a_n2318_13878.n85 a_n2318_13878.t66 512.366
R28 a_n2318_13878.n102 a_n2318_13878.t65 512.366
R29 a_n2318_13878.n92 a_n2318_13878.t56 512.366
R30 a_n2318_13878.n103 a_n2318_13878.t48 512.366
R31 a_n2318_13878.n100 a_n2318_13878.t73 512.366
R32 a_n2318_13878.n93 a_n2318_13878.t62 512.366
R33 a_n2318_13878.n101 a_n2318_13878.t61 512.366
R34 a_n2318_13878.n98 a_n2318_13878.t69 512.366
R35 a_n2318_13878.n94 a_n2318_13878.t55 512.366
R36 a_n2318_13878.n99 a_n2318_13878.t54 512.366
R37 a_n2318_13878.n96 a_n2318_13878.t58 512.366
R38 a_n2318_13878.n95 a_n2318_13878.t67 512.366
R39 a_n2318_13878.n97 a_n2318_13878.t79 512.366
R40 a_n2318_13878.n63 a_n2318_13878.n28 70.1674
R41 a_n2318_13878.n56 a_n2318_13878.n6 70.1674
R42 a_n2318_13878.n18 a_n2318_13878.n42 70.1674
R43 a_n2318_13878.n21 a_n2318_13878.n35 70.1674
R44 a_n2318_13878.n85 a_n2318_13878.n35 20.9683
R45 a_n2318_13878.n34 a_n2318_13878.n22 72.3034
R46 a_n2318_13878.n34 a_n2318_13878.n80 16.6962
R47 a_n2318_13878.n22 a_n2318_13878.n33 77.6622
R48 a_n2318_13878.n84 a_n2318_13878.n33 5.97853
R49 a_n2318_13878.n32 a_n2318_13878.n23 77.6622
R50 a_n2318_13878.n23 a_n2318_13878.n31 72.3034
R51 a_n2318_13878.n81 a_n2318_13878.n29 20.9683
R52 a_n2318_13878.n30 a_n2318_13878.n29 70.1674
R53 a_n2318_13878.n90 a_n2318_13878.n42 20.9683
R54 a_n2318_13878.n41 a_n2318_13878.n19 72.3034
R55 a_n2318_13878.n41 a_n2318_13878.n79 16.6962
R56 a_n2318_13878.n19 a_n2318_13878.n40 77.6622
R57 a_n2318_13878.n89 a_n2318_13878.n40 5.97853
R58 a_n2318_13878.n39 a_n2318_13878.n20 77.6622
R59 a_n2318_13878.n20 a_n2318_13878.n38 72.3034
R60 a_n2318_13878.n86 a_n2318_13878.n36 20.9683
R61 a_n2318_13878.n37 a_n2318_13878.n36 70.1674
R62 a_n2318_13878.n9 a_n2318_13878.n50 70.1674
R63 a_n2318_13878.n11 a_n2318_13878.n48 70.1674
R64 a_n2318_13878.n13 a_n2318_13878.n46 70.1674
R65 a_n2318_13878.n16 a_n2318_13878.n44 70.1674
R66 a_n2318_13878.n97 a_n2318_13878.n44 20.9683
R67 a_n2318_13878.n43 a_n2318_13878.n17 75.0448
R68 a_n2318_13878.n43 a_n2318_13878.n95 11.2134
R69 a_n2318_13878.n17 a_n2318_13878.n96 161.3
R70 a_n2318_13878.n99 a_n2318_13878.n46 20.9683
R71 a_n2318_13878.n45 a_n2318_13878.n14 75.0448
R72 a_n2318_13878.n45 a_n2318_13878.n94 11.2134
R73 a_n2318_13878.n14 a_n2318_13878.n98 161.3
R74 a_n2318_13878.n101 a_n2318_13878.n48 20.9683
R75 a_n2318_13878.n47 a_n2318_13878.n12 75.0448
R76 a_n2318_13878.n47 a_n2318_13878.n93 11.2134
R77 a_n2318_13878.n12 a_n2318_13878.n100 161.3
R78 a_n2318_13878.n103 a_n2318_13878.n50 20.9683
R79 a_n2318_13878.n49 a_n2318_13878.n10 75.0448
R80 a_n2318_13878.n49 a_n2318_13878.n92 11.2134
R81 a_n2318_13878.n10 a_n2318_13878.n102 161.3
R82 a_n2318_13878.n105 a_n2318_13878.n56 20.9683
R83 a_n2318_13878.n7 a_n2318_13878.n55 72.3034
R84 a_n2318_13878.n55 a_n2318_13878.n75 16.6962
R85 a_n2318_13878.n54 a_n2318_13878.n7 77.6622
R86 a_n2318_13878.n106 a_n2318_13878.n54 5.97853
R87 a_n2318_13878.n53 a_n2318_13878.n5 77.6622
R88 a_n2318_13878.n5 a_n2318_13878.n52 72.3034
R89 a_n2318_13878.n108 a_n2318_13878.n51 20.9683
R90 a_n2318_13878.n8 a_n2318_13878.n51 70.1674
R91 a_n2318_13878.n109 a_n2318_13878.n63 20.9683
R92 a_n2318_13878.n28 a_n2318_13878.n62 72.3034
R93 a_n2318_13878.n62 a_n2318_13878.n65 16.6962
R94 a_n2318_13878.n61 a_n2318_13878.n60 77.6622
R95 a_n2318_13878.n110 a_n2318_13878.n61 5.97853
R96 a_n2318_13878.n59 a_n2318_13878.n4 77.6622
R97 a_n2318_13878.n4 a_n2318_13878.n58 72.3034
R98 a_n2318_13878.n112 a_n2318_13878.n57 20.9683
R99 a_n2318_13878.n3 a_n2318_13878.n57 70.1674
R100 a_n2318_13878.n1 a_n2318_13878.n72 81.4626
R101 a_n2318_13878.n2 a_n2318_13878.n68 81.4626
R102 a_n2318_13878.n2 a_n2318_13878.n66 81.4626
R103 a_n2318_13878.n1 a_n2318_13878.n73 80.9324
R104 a_n2318_13878.n1 a_n2318_13878.n71 80.9324
R105 a_n2318_13878.n0 a_n2318_13878.n70 80.9324
R106 a_n2318_13878.n2 a_n2318_13878.n69 80.9324
R107 a_n2318_13878.n2 a_n2318_13878.n67 80.9324
R108 a_n2318_13878.n26 a_n2318_13878.t15 74.6477
R109 a_n2318_13878.n24 a_n2318_13878.t17 74.6477
R110 a_n2318_13878.n27 a_n2318_13878.t7 74.2899
R111 a_n2318_13878.n25 a_n2318_13878.t19 74.2897
R112 a_n2318_13878.n26 a_n2318_13878.n114 70.6783
R113 a_n2318_13878.n26 a_n2318_13878.n115 70.6783
R114 a_n2318_13878.n25 a_n2318_13878.n78 70.6783
R115 a_n2318_13878.n24 a_n2318_13878.n77 70.6783
R116 a_n2318_13878.n24 a_n2318_13878.n76 70.6783
R117 a_n2318_13878.n116 a_n2318_13878.n27 70.6782
R118 a_n2318_13878.n111 a_n2318_13878.n110 48.2005
R119 a_n2318_13878.n63 a_n2318_13878.t14 533.335
R120 a_n2318_13878.n107 a_n2318_13878.n106 48.2005
R121 a_n2318_13878.n56 a_n2318_13878.t50 533.335
R122 a_n2318_13878.n89 a_n2318_13878.n88 48.2005
R123 a_n2318_13878.t18 a_n2318_13878.n42 533.335
R124 a_n2318_13878.n84 a_n2318_13878.n83 48.2005
R125 a_n2318_13878.t51 a_n2318_13878.n35 533.335
R126 a_n2318_13878.n102 a_n2318_13878.n92 48.2005
R127 a_n2318_13878.t70 a_n2318_13878.n50 533.335
R128 a_n2318_13878.n100 a_n2318_13878.n93 48.2005
R129 a_n2318_13878.t77 a_n2318_13878.n48 533.335
R130 a_n2318_13878.n98 a_n2318_13878.n94 48.2005
R131 a_n2318_13878.t64 a_n2318_13878.n46 533.335
R132 a_n2318_13878.n96 a_n2318_13878.n95 48.2005
R133 a_n2318_13878.t60 a_n2318_13878.n44 533.335
R134 a_n2318_13878.n58 a_n2318_13878.n64 16.6962
R135 a_n2318_13878.n109 a_n2318_13878.n62 27.6507
R136 a_n2318_13878.n52 a_n2318_13878.n74 16.6962
R137 a_n2318_13878.n105 a_n2318_13878.n55 27.6507
R138 a_n2318_13878.n87 a_n2318_13878.n38 16.6962
R139 a_n2318_13878.n90 a_n2318_13878.n41 27.6507
R140 a_n2318_13878.n82 a_n2318_13878.n31 16.6962
R141 a_n2318_13878.n85 a_n2318_13878.n34 27.6507
R142 a_n2318_13878.n59 a_n2318_13878.n64 41.7634
R143 a_n2318_13878.n53 a_n2318_13878.n74 41.7634
R144 a_n2318_13878.n87 a_n2318_13878.n39 41.7634
R145 a_n2318_13878.n82 a_n2318_13878.n32 41.7634
R146 a_n2318_13878.n103 a_n2318_13878.n49 35.3134
R147 a_n2318_13878.n101 a_n2318_13878.n47 35.3134
R148 a_n2318_13878.n99 a_n2318_13878.n45 35.3134
R149 a_n2318_13878.n97 a_n2318_13878.n43 35.3134
R150 a_n2318_13878.n28 a_n2318_13878.n1 23.891
R151 a_n2318_13878.n30 a_n2318_13878.n15 12.705
R152 a_n2318_13878.n6 a_n2318_13878.n104 12.5005
R153 a_n2318_13878.n59 a_n2318_13878.n111 5.97853
R154 a_n2318_13878.n61 a_n2318_13878.n65 41.7634
R155 a_n2318_13878.n53 a_n2318_13878.n107 5.97853
R156 a_n2318_13878.n54 a_n2318_13878.n75 41.7634
R157 a_n2318_13878.n88 a_n2318_13878.n39 5.97853
R158 a_n2318_13878.n79 a_n2318_13878.n40 41.7634
R159 a_n2318_13878.n83 a_n2318_13878.n32 5.97853
R160 a_n2318_13878.n80 a_n2318_13878.n33 41.7634
R161 a_n2318_13878.n0 a_n2318_13878.n2 32.5247
R162 a_n2318_13878.n113 a_n2318_13878.n3 11.1956
R163 a_n2318_13878.n112 a_n2318_13878.n58 27.6507
R164 a_n2318_13878.n108 a_n2318_13878.n52 27.6507
R165 a_n2318_13878.n38 a_n2318_13878.n86 27.6507
R166 a_n2318_13878.n31 a_n2318_13878.n81 27.6507
R167 a_n2318_13878.n91 a_n2318_13878.n25 9.85898
R168 a_n2318_13878.n17 a_n2318_13878.n15 8.73345
R169 a_n2318_13878.n104 a_n2318_13878.n9 8.73345
R170 a_n2318_13878.n91 a_n2318_13878.n18 7.36035
R171 a_n2318_13878.n27 a_n2318_13878.n113 6.01559
R172 a_n2318_13878.n104 a_n2318_13878.n91 5.3452
R173 a_n2318_13878.n37 a_n2318_13878.n21 4.01186
R174 a_n2318_13878.n28 a_n2318_13878.n8 4.0079
R175 a_n2318_13878.n114 a_n2318_13878.t27 3.61217
R176 a_n2318_13878.n114 a_n2318_13878.t23 3.61217
R177 a_n2318_13878.n115 a_n2318_13878.t29 3.61217
R178 a_n2318_13878.n115 a_n2318_13878.t3 3.61217
R179 a_n2318_13878.n78 a_n2318_13878.t11 3.61217
R180 a_n2318_13878.n78 a_n2318_13878.t21 3.61217
R181 a_n2318_13878.n77 a_n2318_13878.t13 3.61217
R182 a_n2318_13878.n77 a_n2318_13878.t31 3.61217
R183 a_n2318_13878.n76 a_n2318_13878.t25 3.61217
R184 a_n2318_13878.n76 a_n2318_13878.t9 3.61217
R185 a_n2318_13878.t1 a_n2318_13878.n116 3.61217
R186 a_n2318_13878.n116 a_n2318_13878.t5 3.61217
R187 a_n2318_13878.n72 a_n2318_13878.t38 2.82907
R188 a_n2318_13878.n72 a_n2318_13878.t34 2.82907
R189 a_n2318_13878.n73 a_n2318_13878.t35 2.82907
R190 a_n2318_13878.n73 a_n2318_13878.t36 2.82907
R191 a_n2318_13878.n71 a_n2318_13878.t45 2.82907
R192 a_n2318_13878.n71 a_n2318_13878.t47 2.82907
R193 a_n2318_13878.n70 a_n2318_13878.t39 2.82907
R194 a_n2318_13878.n70 a_n2318_13878.t42 2.82907
R195 a_n2318_13878.n68 a_n2318_13878.t40 2.82907
R196 a_n2318_13878.n68 a_n2318_13878.t37 2.82907
R197 a_n2318_13878.n69 a_n2318_13878.t33 2.82907
R198 a_n2318_13878.n69 a_n2318_13878.t32 2.82907
R199 a_n2318_13878.n67 a_n2318_13878.t44 2.82907
R200 a_n2318_13878.n67 a_n2318_13878.t46 2.82907
R201 a_n2318_13878.n66 a_n2318_13878.t41 2.82907
R202 a_n2318_13878.n66 a_n2318_13878.t43 2.82907
R203 a_n2318_13878.n113 a_n2318_13878.n15 1.30542
R204 a_n2318_13878.n27 a_n2318_13878.n26 1.07378
R205 a_n2318_13878.n25 a_n2318_13878.n24 1.07378
R206 a_n2318_13878.n1 a_n2318_13878.n0 1.06084
R207 a_n2318_13878.n12 a_n2318_13878.n13 1.04595
R208 a_n2318_13878.n23 a_n2318_13878.n22 0.758076
R209 a_n2318_13878.n22 a_n2318_13878.n21 0.758076
R210 a_n2318_13878.n20 a_n2318_13878.n19 0.758076
R211 a_n2318_13878.n19 a_n2318_13878.n18 0.758076
R212 a_n2318_13878.n17 a_n2318_13878.n16 0.758076
R213 a_n2318_13878.n14 a_n2318_13878.n13 0.758076
R214 a_n2318_13878.n12 a_n2318_13878.n11 0.758076
R215 a_n2318_13878.n10 a_n2318_13878.n9 0.758076
R216 a_n2318_13878.n7 a_n2318_13878.n5 0.758076
R217 a_n2318_13878.n7 a_n2318_13878.n6 0.758076
R218 a_n2318_13878.n60 a_n2318_13878.n4 0.758076
R219 a_n2318_13878.n60 a_n2318_13878.n28 0.724161
R220 a_n2318_13878.n14 a_n2318_13878.n16 0.67853
R221 a_n2318_13878.n10 a_n2318_13878.n11 0.67853
R222 a_n2318_13878.n4 a_n2318_13878.n3 0.568682
R223 a_n2318_13878.n5 a_n2318_13878.n8 0.568682
R224 a_n2318_13878.n37 a_n2318_13878.n20 0.568682
R225 a_n2318_13878.n30 a_n2318_13878.n23 0.568682
R226 a_n2140_13878.n21 a_n2140_13878.n20 98.9632
R227 a_n2140_13878.n2 a_n2140_13878.n0 98.7517
R228 a_n2140_13878.n18 a_n2140_13878.n17 98.6055
R229 a_n2140_13878.n20 a_n2140_13878.n19 98.6055
R230 a_n2140_13878.n6 a_n2140_13878.n5 98.6055
R231 a_n2140_13878.n4 a_n2140_13878.n3 98.6055
R232 a_n2140_13878.n2 a_n2140_13878.n1 98.6055
R233 a_n2140_13878.n16 a_n2140_13878.n15 98.6054
R234 a_n2140_13878.n8 a_n2140_13878.t2 74.6477
R235 a_n2140_13878.n13 a_n2140_13878.t1 74.2899
R236 a_n2140_13878.n10 a_n2140_13878.t3 74.2899
R237 a_n2140_13878.n9 a_n2140_13878.t23 74.2899
R238 a_n2140_13878.n12 a_n2140_13878.n11 70.6783
R239 a_n2140_13878.n8 a_n2140_13878.n7 70.6783
R240 a_n2140_13878.n14 a_n2140_13878.n6 14.2849
R241 a_n2140_13878.n16 a_n2140_13878.n14 11.9339
R242 a_n2140_13878.n14 a_n2140_13878.n13 6.95632
R243 a_n2140_13878.n15 a_n2140_13878.t11 3.61217
R244 a_n2140_13878.n15 a_n2140_13878.t12 3.61217
R245 a_n2140_13878.n17 a_n2140_13878.t18 3.61217
R246 a_n2140_13878.n17 a_n2140_13878.t19 3.61217
R247 a_n2140_13878.n19 a_n2140_13878.t5 3.61217
R248 a_n2140_13878.n19 a_n2140_13878.t13 3.61217
R249 a_n2140_13878.n11 a_n2140_13878.t0 3.61217
R250 a_n2140_13878.n11 a_n2140_13878.t4 3.61217
R251 a_n2140_13878.n7 a_n2140_13878.t21 3.61217
R252 a_n2140_13878.n7 a_n2140_13878.t22 3.61217
R253 a_n2140_13878.n5 a_n2140_13878.t14 3.61217
R254 a_n2140_13878.n5 a_n2140_13878.t6 3.61217
R255 a_n2140_13878.n3 a_n2140_13878.t17 3.61217
R256 a_n2140_13878.n3 a_n2140_13878.t8 3.61217
R257 a_n2140_13878.n1 a_n2140_13878.t7 3.61217
R258 a_n2140_13878.n1 a_n2140_13878.t9 3.61217
R259 a_n2140_13878.n0 a_n2140_13878.t15 3.61217
R260 a_n2140_13878.n0 a_n2140_13878.t10 3.61217
R261 a_n2140_13878.n21 a_n2140_13878.t16 3.61217
R262 a_n2140_13878.t20 a_n2140_13878.n21 3.61217
R263 a_n2140_13878.n9 a_n2140_13878.n8 0.358259
R264 a_n2140_13878.n12 a_n2140_13878.n10 0.358259
R265 a_n2140_13878.n13 a_n2140_13878.n12 0.358259
R266 a_n2140_13878.n20 a_n2140_13878.n18 0.358259
R267 a_n2140_13878.n18 a_n2140_13878.n16 0.358259
R268 a_n2140_13878.n4 a_n2140_13878.n2 0.146627
R269 a_n2140_13878.n6 a_n2140_13878.n4 0.146627
R270 a_n2140_13878.n10 a_n2140_13878.n9 0.101793
R271 vdd.n315 vdd.n279 756.745
R272 vdd.n260 vdd.n224 756.745
R273 vdd.n217 vdd.n181 756.745
R274 vdd.n162 vdd.n126 756.745
R275 vdd.n120 vdd.n84 756.745
R276 vdd.n65 vdd.n29 756.745
R277 vdd.n2046 vdd.n2010 756.745
R278 vdd.n2101 vdd.n2065 756.745
R279 vdd.n1948 vdd.n1912 756.745
R280 vdd.n2003 vdd.n1967 756.745
R281 vdd.n1851 vdd.n1815 756.745
R282 vdd.n1906 vdd.n1870 756.745
R283 vdd.n1224 vdd.t21 640.208
R284 vdd.n952 vdd.t63 640.208
R285 vdd.n1244 vdd.t36 640.208
R286 vdd.n943 vdd.t81 640.208
R287 vdd.n843 vdd.t39 640.208
R288 vdd.n2621 vdd.t75 640.208
R289 vdd.n804 vdd.t87 640.208
R290 vdd.n2618 vdd.t67 640.208
R291 vdd.n768 vdd.t17 640.208
R292 vdd.n1014 vdd.t71 640.208
R293 vdd.n1510 vdd.t54 592.009
R294 vdd.n1666 vdd.t46 592.009
R295 vdd.n1702 vdd.t57 592.009
R296 vdd.n2186 vdd.t29 592.009
R297 vdd.n1161 vdd.t60 592.009
R298 vdd.n1121 vdd.t78 592.009
R299 vdd.n405 vdd.t50 592.009
R300 vdd.n419 vdd.t84 592.009
R301 vdd.n431 vdd.t90 592.009
R302 vdd.n723 vdd.t33 592.009
R303 vdd.n686 vdd.t43 592.009
R304 vdd.n3105 vdd.t25 592.009
R305 vdd.n316 vdd.n315 585
R306 vdd.n314 vdd.n281 585
R307 vdd.n313 vdd.n312 585
R308 vdd.n284 vdd.n282 585
R309 vdd.n307 vdd.n306 585
R310 vdd.n305 vdd.n304 585
R311 vdd.n288 vdd.n287 585
R312 vdd.n299 vdd.n298 585
R313 vdd.n297 vdd.n296 585
R314 vdd.n292 vdd.n291 585
R315 vdd.n261 vdd.n260 585
R316 vdd.n259 vdd.n226 585
R317 vdd.n258 vdd.n257 585
R318 vdd.n229 vdd.n227 585
R319 vdd.n252 vdd.n251 585
R320 vdd.n250 vdd.n249 585
R321 vdd.n233 vdd.n232 585
R322 vdd.n244 vdd.n243 585
R323 vdd.n242 vdd.n241 585
R324 vdd.n237 vdd.n236 585
R325 vdd.n218 vdd.n217 585
R326 vdd.n216 vdd.n183 585
R327 vdd.n215 vdd.n214 585
R328 vdd.n186 vdd.n184 585
R329 vdd.n209 vdd.n208 585
R330 vdd.n207 vdd.n206 585
R331 vdd.n190 vdd.n189 585
R332 vdd.n201 vdd.n200 585
R333 vdd.n199 vdd.n198 585
R334 vdd.n194 vdd.n193 585
R335 vdd.n163 vdd.n162 585
R336 vdd.n161 vdd.n128 585
R337 vdd.n160 vdd.n159 585
R338 vdd.n131 vdd.n129 585
R339 vdd.n154 vdd.n153 585
R340 vdd.n152 vdd.n151 585
R341 vdd.n135 vdd.n134 585
R342 vdd.n146 vdd.n145 585
R343 vdd.n144 vdd.n143 585
R344 vdd.n139 vdd.n138 585
R345 vdd.n121 vdd.n120 585
R346 vdd.n119 vdd.n86 585
R347 vdd.n118 vdd.n117 585
R348 vdd.n89 vdd.n87 585
R349 vdd.n112 vdd.n111 585
R350 vdd.n110 vdd.n109 585
R351 vdd.n93 vdd.n92 585
R352 vdd.n104 vdd.n103 585
R353 vdd.n102 vdd.n101 585
R354 vdd.n97 vdd.n96 585
R355 vdd.n66 vdd.n65 585
R356 vdd.n64 vdd.n31 585
R357 vdd.n63 vdd.n62 585
R358 vdd.n34 vdd.n32 585
R359 vdd.n57 vdd.n56 585
R360 vdd.n55 vdd.n54 585
R361 vdd.n38 vdd.n37 585
R362 vdd.n49 vdd.n48 585
R363 vdd.n47 vdd.n46 585
R364 vdd.n42 vdd.n41 585
R365 vdd.n2047 vdd.n2046 585
R366 vdd.n2045 vdd.n2012 585
R367 vdd.n2044 vdd.n2043 585
R368 vdd.n2015 vdd.n2013 585
R369 vdd.n2038 vdd.n2037 585
R370 vdd.n2036 vdd.n2035 585
R371 vdd.n2019 vdd.n2018 585
R372 vdd.n2030 vdd.n2029 585
R373 vdd.n2028 vdd.n2027 585
R374 vdd.n2023 vdd.n2022 585
R375 vdd.n2102 vdd.n2101 585
R376 vdd.n2100 vdd.n2067 585
R377 vdd.n2099 vdd.n2098 585
R378 vdd.n2070 vdd.n2068 585
R379 vdd.n2093 vdd.n2092 585
R380 vdd.n2091 vdd.n2090 585
R381 vdd.n2074 vdd.n2073 585
R382 vdd.n2085 vdd.n2084 585
R383 vdd.n2083 vdd.n2082 585
R384 vdd.n2078 vdd.n2077 585
R385 vdd.n1949 vdd.n1948 585
R386 vdd.n1947 vdd.n1914 585
R387 vdd.n1946 vdd.n1945 585
R388 vdd.n1917 vdd.n1915 585
R389 vdd.n1940 vdd.n1939 585
R390 vdd.n1938 vdd.n1937 585
R391 vdd.n1921 vdd.n1920 585
R392 vdd.n1932 vdd.n1931 585
R393 vdd.n1930 vdd.n1929 585
R394 vdd.n1925 vdd.n1924 585
R395 vdd.n2004 vdd.n2003 585
R396 vdd.n2002 vdd.n1969 585
R397 vdd.n2001 vdd.n2000 585
R398 vdd.n1972 vdd.n1970 585
R399 vdd.n1995 vdd.n1994 585
R400 vdd.n1993 vdd.n1992 585
R401 vdd.n1976 vdd.n1975 585
R402 vdd.n1987 vdd.n1986 585
R403 vdd.n1985 vdd.n1984 585
R404 vdd.n1980 vdd.n1979 585
R405 vdd.n1852 vdd.n1851 585
R406 vdd.n1850 vdd.n1817 585
R407 vdd.n1849 vdd.n1848 585
R408 vdd.n1820 vdd.n1818 585
R409 vdd.n1843 vdd.n1842 585
R410 vdd.n1841 vdd.n1840 585
R411 vdd.n1824 vdd.n1823 585
R412 vdd.n1835 vdd.n1834 585
R413 vdd.n1833 vdd.n1832 585
R414 vdd.n1828 vdd.n1827 585
R415 vdd.n1907 vdd.n1906 585
R416 vdd.n1905 vdd.n1872 585
R417 vdd.n1904 vdd.n1903 585
R418 vdd.n1875 vdd.n1873 585
R419 vdd.n1898 vdd.n1897 585
R420 vdd.n1896 vdd.n1895 585
R421 vdd.n1879 vdd.n1878 585
R422 vdd.n1890 vdd.n1889 585
R423 vdd.n1888 vdd.n1887 585
R424 vdd.n1883 vdd.n1882 585
R425 vdd.n445 vdd.n370 462.44
R426 vdd.n3343 vdd.n372 462.44
R427 vdd.n3238 vdd.n657 462.44
R428 vdd.n3236 vdd.n660 462.44
R429 vdd.n2181 vdd.n1409 462.44
R430 vdd.n2184 vdd.n2183 462.44
R431 vdd.n1737 vdd.n1507 462.44
R432 vdd.n1734 vdd.n1505 462.44
R433 vdd.n293 vdd.t244 329.043
R434 vdd.n238 vdd.t168 329.043
R435 vdd.n195 vdd.t191 329.043
R436 vdd.n140 vdd.t162 329.043
R437 vdd.n98 vdd.t151 329.043
R438 vdd.n43 vdd.t187 329.043
R439 vdd.n2024 vdd.t170 329.043
R440 vdd.n2079 vdd.t109 329.043
R441 vdd.n1926 vdd.t243 329.043
R442 vdd.n1981 vdd.t155 329.043
R443 vdd.n1829 vdd.t186 329.043
R444 vdd.n1884 vdd.t129 329.043
R445 vdd.n1510 vdd.t56 319.788
R446 vdd.n1666 vdd.t49 319.788
R447 vdd.n1702 vdd.t59 319.788
R448 vdd.n2186 vdd.t31 319.788
R449 vdd.n1161 vdd.t61 319.788
R450 vdd.n1121 vdd.t79 319.788
R451 vdd.n405 vdd.t52 319.788
R452 vdd.n419 vdd.t85 319.788
R453 vdd.n431 vdd.t91 319.788
R454 vdd.n723 vdd.t35 319.788
R455 vdd.n686 vdd.t45 319.788
R456 vdd.n3105 vdd.t28 319.788
R457 vdd.n1511 vdd.t55 303.69
R458 vdd.n1667 vdd.t48 303.69
R459 vdd.n1703 vdd.t58 303.69
R460 vdd.n2187 vdd.t32 303.69
R461 vdd.n1162 vdd.t62 303.69
R462 vdd.n1122 vdd.t80 303.69
R463 vdd.n406 vdd.t53 303.69
R464 vdd.n420 vdd.t86 303.69
R465 vdd.n432 vdd.t92 303.69
R466 vdd.n724 vdd.t34 303.69
R467 vdd.n687 vdd.t44 303.69
R468 vdd.n3106 vdd.t27 303.69
R469 vdd.n2853 vdd.n898 291.221
R470 vdd.n3067 vdd.n778 291.221
R471 vdd.n3004 vdd.n775 291.221
R472 vdd.n2785 vdd.n2784 291.221
R473 vdd.n2581 vdd.n940 291.221
R474 vdd.n2512 vdd.n2511 291.221
R475 vdd.n1280 vdd.n1279 291.221
R476 vdd.n2332 vdd.n1046 291.221
R477 vdd.n2983 vdd.n776 291.221
R478 vdd.n3070 vdd.n3069 291.221
R479 vdd.n2689 vdd.n2615 291.221
R480 vdd.n2857 vdd.n902 291.221
R481 vdd.n2509 vdd.n950 291.221
R482 vdd.n948 vdd.n922 291.221
R483 vdd.n1358 vdd.n1087 291.221
R484 vdd.n2336 vdd.n1051 291.221
R485 vdd.n2985 vdd.n776 185
R486 vdd.n3068 vdd.n776 185
R487 vdd.n2987 vdd.n2986 185
R488 vdd.n2986 vdd.n774 185
R489 vdd.n2988 vdd.n810 185
R490 vdd.n2998 vdd.n810 185
R491 vdd.n2989 vdd.n819 185
R492 vdd.n819 vdd.n817 185
R493 vdd.n2991 vdd.n2990 185
R494 vdd.n2992 vdd.n2991 185
R495 vdd.n2944 vdd.n818 185
R496 vdd.n818 vdd.n814 185
R497 vdd.n2943 vdd.n2942 185
R498 vdd.n2942 vdd.n2941 185
R499 vdd.n821 vdd.n820 185
R500 vdd.n822 vdd.n821 185
R501 vdd.n2934 vdd.n2933 185
R502 vdd.n2935 vdd.n2934 185
R503 vdd.n2932 vdd.n831 185
R504 vdd.n831 vdd.n828 185
R505 vdd.n2931 vdd.n2930 185
R506 vdd.n2930 vdd.n2929 185
R507 vdd.n833 vdd.n832 185
R508 vdd.n841 vdd.n833 185
R509 vdd.n2922 vdd.n2921 185
R510 vdd.n2923 vdd.n2922 185
R511 vdd.n2919 vdd.n842 185
R512 vdd.n849 vdd.n842 185
R513 vdd.n2918 vdd.n2917 185
R514 vdd.n2917 vdd.n2916 185
R515 vdd.n845 vdd.n844 185
R516 vdd.n846 vdd.n845 185
R517 vdd.n2909 vdd.n2908 185
R518 vdd.n2910 vdd.n2909 185
R519 vdd.n2907 vdd.n856 185
R520 vdd.n856 vdd.n853 185
R521 vdd.n2906 vdd.n2905 185
R522 vdd.n2905 vdd.n2904 185
R523 vdd.n858 vdd.n857 185
R524 vdd.n866 vdd.n858 185
R525 vdd.n2897 vdd.n2896 185
R526 vdd.n2898 vdd.n2897 185
R527 vdd.n2895 vdd.n867 185
R528 vdd.n872 vdd.n867 185
R529 vdd.n2894 vdd.n2893 185
R530 vdd.n2893 vdd.n2892 185
R531 vdd.n869 vdd.n868 185
R532 vdd.n2764 vdd.n869 185
R533 vdd.n2885 vdd.n2884 185
R534 vdd.n2886 vdd.n2885 185
R535 vdd.n2883 vdd.n879 185
R536 vdd.n879 vdd.n876 185
R537 vdd.n2882 vdd.n2881 185
R538 vdd.n2881 vdd.n2880 185
R539 vdd.n881 vdd.n880 185
R540 vdd.n882 vdd.n881 185
R541 vdd.n2873 vdd.n2872 185
R542 vdd.n2874 vdd.n2873 185
R543 vdd.n2871 vdd.n891 185
R544 vdd.n891 vdd.n888 185
R545 vdd.n2870 vdd.n2869 185
R546 vdd.n2869 vdd.n2868 185
R547 vdd.n893 vdd.n892 185
R548 vdd.n2779 vdd.n893 185
R549 vdd.n2861 vdd.n2860 185
R550 vdd.n2862 vdd.n2861 185
R551 vdd.n2859 vdd.n902 185
R552 vdd.n902 vdd.n899 185
R553 vdd.n2858 vdd.n2857 185
R554 vdd.n904 vdd.n903 185
R555 vdd.n2625 vdd.n2624 185
R556 vdd.n2627 vdd.n2626 185
R557 vdd.n2629 vdd.n2628 185
R558 vdd.n2631 vdd.n2630 185
R559 vdd.n2633 vdd.n2632 185
R560 vdd.n2635 vdd.n2634 185
R561 vdd.n2637 vdd.n2636 185
R562 vdd.n2639 vdd.n2638 185
R563 vdd.n2641 vdd.n2640 185
R564 vdd.n2643 vdd.n2642 185
R565 vdd.n2645 vdd.n2644 185
R566 vdd.n2647 vdd.n2646 185
R567 vdd.n2649 vdd.n2648 185
R568 vdd.n2651 vdd.n2650 185
R569 vdd.n2653 vdd.n2652 185
R570 vdd.n2655 vdd.n2654 185
R571 vdd.n2657 vdd.n2656 185
R572 vdd.n2659 vdd.n2658 185
R573 vdd.n2661 vdd.n2660 185
R574 vdd.n2663 vdd.n2662 185
R575 vdd.n2665 vdd.n2664 185
R576 vdd.n2667 vdd.n2666 185
R577 vdd.n2669 vdd.n2668 185
R578 vdd.n2671 vdd.n2670 185
R579 vdd.n2673 vdd.n2672 185
R580 vdd.n2675 vdd.n2674 185
R581 vdd.n2677 vdd.n2676 185
R582 vdd.n2679 vdd.n2678 185
R583 vdd.n2681 vdd.n2680 185
R584 vdd.n2683 vdd.n2682 185
R585 vdd.n2685 vdd.n2684 185
R586 vdd.n2687 vdd.n2686 185
R587 vdd.n2688 vdd.n2615 185
R588 vdd.n2855 vdd.n2615 185
R589 vdd.n3071 vdd.n3070 185
R590 vdd.n3072 vdd.n767 185
R591 vdd.n3074 vdd.n3073 185
R592 vdd.n3076 vdd.n765 185
R593 vdd.n3078 vdd.n3077 185
R594 vdd.n3079 vdd.n764 185
R595 vdd.n3081 vdd.n3080 185
R596 vdd.n3083 vdd.n762 185
R597 vdd.n3085 vdd.n3084 185
R598 vdd.n3086 vdd.n761 185
R599 vdd.n3088 vdd.n3087 185
R600 vdd.n3090 vdd.n759 185
R601 vdd.n3092 vdd.n3091 185
R602 vdd.n3093 vdd.n758 185
R603 vdd.n3095 vdd.n3094 185
R604 vdd.n3097 vdd.n757 185
R605 vdd.n3098 vdd.n754 185
R606 vdd.n3101 vdd.n3100 185
R607 vdd.n755 vdd.n753 185
R608 vdd.n2957 vdd.n2956 185
R609 vdd.n2959 vdd.n2958 185
R610 vdd.n2961 vdd.n2953 185
R611 vdd.n2963 vdd.n2962 185
R612 vdd.n2964 vdd.n2952 185
R613 vdd.n2966 vdd.n2965 185
R614 vdd.n2968 vdd.n2950 185
R615 vdd.n2970 vdd.n2969 185
R616 vdd.n2971 vdd.n2949 185
R617 vdd.n2973 vdd.n2972 185
R618 vdd.n2975 vdd.n2947 185
R619 vdd.n2977 vdd.n2976 185
R620 vdd.n2978 vdd.n2946 185
R621 vdd.n2980 vdd.n2979 185
R622 vdd.n2982 vdd.n2945 185
R623 vdd.n2984 vdd.n2983 185
R624 vdd.n2983 vdd.n756 185
R625 vdd.n3069 vdd.n771 185
R626 vdd.n3069 vdd.n3068 185
R627 vdd.n2692 vdd.n773 185
R628 vdd.n774 vdd.n773 185
R629 vdd.n2693 vdd.n809 185
R630 vdd.n2998 vdd.n809 185
R631 vdd.n2695 vdd.n2694 185
R632 vdd.n2694 vdd.n817 185
R633 vdd.n2696 vdd.n816 185
R634 vdd.n2992 vdd.n816 185
R635 vdd.n2698 vdd.n2697 185
R636 vdd.n2697 vdd.n814 185
R637 vdd.n2699 vdd.n824 185
R638 vdd.n2941 vdd.n824 185
R639 vdd.n2701 vdd.n2700 185
R640 vdd.n2700 vdd.n822 185
R641 vdd.n2702 vdd.n830 185
R642 vdd.n2935 vdd.n830 185
R643 vdd.n2704 vdd.n2703 185
R644 vdd.n2703 vdd.n828 185
R645 vdd.n2705 vdd.n835 185
R646 vdd.n2929 vdd.n835 185
R647 vdd.n2707 vdd.n2706 185
R648 vdd.n2706 vdd.n841 185
R649 vdd.n2708 vdd.n840 185
R650 vdd.n2923 vdd.n840 185
R651 vdd.n2710 vdd.n2709 185
R652 vdd.n2709 vdd.n849 185
R653 vdd.n2711 vdd.n848 185
R654 vdd.n2916 vdd.n848 185
R655 vdd.n2713 vdd.n2712 185
R656 vdd.n2712 vdd.n846 185
R657 vdd.n2714 vdd.n855 185
R658 vdd.n2910 vdd.n855 185
R659 vdd.n2716 vdd.n2715 185
R660 vdd.n2715 vdd.n853 185
R661 vdd.n2717 vdd.n860 185
R662 vdd.n2904 vdd.n860 185
R663 vdd.n2719 vdd.n2718 185
R664 vdd.n2718 vdd.n866 185
R665 vdd.n2720 vdd.n865 185
R666 vdd.n2898 vdd.n865 185
R667 vdd.n2722 vdd.n2721 185
R668 vdd.n2721 vdd.n872 185
R669 vdd.n2723 vdd.n871 185
R670 vdd.n2892 vdd.n871 185
R671 vdd.n2766 vdd.n2765 185
R672 vdd.n2765 vdd.n2764 185
R673 vdd.n2767 vdd.n878 185
R674 vdd.n2886 vdd.n878 185
R675 vdd.n2769 vdd.n2768 185
R676 vdd.n2768 vdd.n876 185
R677 vdd.n2770 vdd.n884 185
R678 vdd.n2880 vdd.n884 185
R679 vdd.n2772 vdd.n2771 185
R680 vdd.n2771 vdd.n882 185
R681 vdd.n2773 vdd.n890 185
R682 vdd.n2874 vdd.n890 185
R683 vdd.n2775 vdd.n2774 185
R684 vdd.n2774 vdd.n888 185
R685 vdd.n2776 vdd.n895 185
R686 vdd.n2868 vdd.n895 185
R687 vdd.n2778 vdd.n2777 185
R688 vdd.n2779 vdd.n2778 185
R689 vdd.n2691 vdd.n901 185
R690 vdd.n2862 vdd.n901 185
R691 vdd.n2690 vdd.n2689 185
R692 vdd.n2689 vdd.n899 185
R693 vdd.n2181 vdd.n2180 185
R694 vdd.n2182 vdd.n2181 185
R695 vdd.n1410 vdd.n1408 185
R696 vdd.n1408 vdd.n1407 185
R697 vdd.n2176 vdd.n2175 185
R698 vdd.n2175 vdd.n2174 185
R699 vdd.n1413 vdd.n1412 185
R700 vdd.n1414 vdd.n1413 185
R701 vdd.n2163 vdd.n2162 185
R702 vdd.n2164 vdd.n2163 185
R703 vdd.n1422 vdd.n1421 185
R704 vdd.n2155 vdd.n1421 185
R705 vdd.n2158 vdd.n2157 185
R706 vdd.n2157 vdd.n2156 185
R707 vdd.n1425 vdd.n1424 185
R708 vdd.n1431 vdd.n1425 185
R709 vdd.n2146 vdd.n2145 185
R710 vdd.n2147 vdd.n2146 185
R711 vdd.n1433 vdd.n1432 185
R712 vdd.n2138 vdd.n1432 185
R713 vdd.n2141 vdd.n2140 185
R714 vdd.n2140 vdd.n2139 185
R715 vdd.n1436 vdd.n1435 185
R716 vdd.n1437 vdd.n1436 185
R717 vdd.n2129 vdd.n2128 185
R718 vdd.n2130 vdd.n2129 185
R719 vdd.n1445 vdd.n1444 185
R720 vdd.n1444 vdd.n1443 185
R721 vdd.n2124 vdd.n2123 185
R722 vdd.n2123 vdd.n2122 185
R723 vdd.n1448 vdd.n1447 185
R724 vdd.n1454 vdd.n1448 185
R725 vdd.n2113 vdd.n2112 185
R726 vdd.n2114 vdd.n2113 185
R727 vdd.n1456 vdd.n1455 185
R728 vdd.n1810 vdd.n1455 185
R729 vdd.n1813 vdd.n1812 185
R730 vdd.n1812 vdd.n1811 185
R731 vdd.n1459 vdd.n1458 185
R732 vdd.n1466 vdd.n1459 185
R733 vdd.n1801 vdd.n1800 185
R734 vdd.n1802 vdd.n1801 185
R735 vdd.n1468 vdd.n1467 185
R736 vdd.n1467 vdd.n1465 185
R737 vdd.n1796 vdd.n1795 185
R738 vdd.n1795 vdd.n1794 185
R739 vdd.n1471 vdd.n1470 185
R740 vdd.n1472 vdd.n1471 185
R741 vdd.n1785 vdd.n1784 185
R742 vdd.n1786 vdd.n1785 185
R743 vdd.n1479 vdd.n1478 185
R744 vdd.n1777 vdd.n1478 185
R745 vdd.n1780 vdd.n1779 185
R746 vdd.n1779 vdd.n1778 185
R747 vdd.n1482 vdd.n1481 185
R748 vdd.n1488 vdd.n1482 185
R749 vdd.n1768 vdd.n1767 185
R750 vdd.n1769 vdd.n1768 185
R751 vdd.n1490 vdd.n1489 185
R752 vdd.n1760 vdd.n1489 185
R753 vdd.n1763 vdd.n1762 185
R754 vdd.n1762 vdd.n1761 185
R755 vdd.n1493 vdd.n1492 185
R756 vdd.n1494 vdd.n1493 185
R757 vdd.n1751 vdd.n1750 185
R758 vdd.n1752 vdd.n1751 185
R759 vdd.n1502 vdd.n1501 185
R760 vdd.n1501 vdd.n1500 185
R761 vdd.n1746 vdd.n1745 185
R762 vdd.n1745 vdd.n1744 185
R763 vdd.n1505 vdd.n1504 185
R764 vdd.n1506 vdd.n1505 185
R765 vdd.n1734 vdd.n1733 185
R766 vdd.n1732 vdd.n1545 185
R767 vdd.n1547 vdd.n1544 185
R768 vdd.n1736 vdd.n1544 185
R769 vdd.n1728 vdd.n1549 185
R770 vdd.n1727 vdd.n1550 185
R771 vdd.n1726 vdd.n1551 185
R772 vdd.n1554 vdd.n1552 185
R773 vdd.n1722 vdd.n1555 185
R774 vdd.n1721 vdd.n1556 185
R775 vdd.n1720 vdd.n1557 185
R776 vdd.n1560 vdd.n1558 185
R777 vdd.n1716 vdd.n1561 185
R778 vdd.n1715 vdd.n1562 185
R779 vdd.n1714 vdd.n1563 185
R780 vdd.n1566 vdd.n1564 185
R781 vdd.n1710 vdd.n1567 185
R782 vdd.n1709 vdd.n1568 185
R783 vdd.n1708 vdd.n1569 185
R784 vdd.n1700 vdd.n1570 185
R785 vdd.n1704 vdd.n1701 185
R786 vdd.n1699 vdd.n1572 185
R787 vdd.n1698 vdd.n1573 185
R788 vdd.n1576 vdd.n1574 185
R789 vdd.n1694 vdd.n1577 185
R790 vdd.n1693 vdd.n1578 185
R791 vdd.n1692 vdd.n1579 185
R792 vdd.n1582 vdd.n1580 185
R793 vdd.n1688 vdd.n1583 185
R794 vdd.n1687 vdd.n1584 185
R795 vdd.n1686 vdd.n1585 185
R796 vdd.n1588 vdd.n1586 185
R797 vdd.n1682 vdd.n1589 185
R798 vdd.n1681 vdd.n1590 185
R799 vdd.n1680 vdd.n1591 185
R800 vdd.n1594 vdd.n1592 185
R801 vdd.n1676 vdd.n1595 185
R802 vdd.n1675 vdd.n1596 185
R803 vdd.n1674 vdd.n1597 185
R804 vdd.n1600 vdd.n1598 185
R805 vdd.n1670 vdd.n1601 185
R806 vdd.n1669 vdd.n1602 185
R807 vdd.n1668 vdd.n1665 185
R808 vdd.n1605 vdd.n1603 185
R809 vdd.n1661 vdd.n1606 185
R810 vdd.n1660 vdd.n1607 185
R811 vdd.n1659 vdd.n1608 185
R812 vdd.n1611 vdd.n1609 185
R813 vdd.n1655 vdd.n1612 185
R814 vdd.n1654 vdd.n1613 185
R815 vdd.n1653 vdd.n1614 185
R816 vdd.n1617 vdd.n1615 185
R817 vdd.n1649 vdd.n1618 185
R818 vdd.n1648 vdd.n1619 185
R819 vdd.n1647 vdd.n1620 185
R820 vdd.n1623 vdd.n1621 185
R821 vdd.n1643 vdd.n1624 185
R822 vdd.n1642 vdd.n1625 185
R823 vdd.n1641 vdd.n1626 185
R824 vdd.n1629 vdd.n1627 185
R825 vdd.n1637 vdd.n1630 185
R826 vdd.n1636 vdd.n1631 185
R827 vdd.n1635 vdd.n1632 185
R828 vdd.n1633 vdd.n1513 185
R829 vdd.n1738 vdd.n1737 185
R830 vdd.n1737 vdd.n1736 185
R831 vdd.n2185 vdd.n2184 185
R832 vdd.n2189 vdd.n1403 185
R833 vdd.n1402 vdd.n1396 185
R834 vdd.n1400 vdd.n1399 185
R835 vdd.n1398 vdd.n1192 185
R836 vdd.n2193 vdd.n1189 185
R837 vdd.n2195 vdd.n2194 185
R838 vdd.n2197 vdd.n1187 185
R839 vdd.n2199 vdd.n2198 185
R840 vdd.n2200 vdd.n1182 185
R841 vdd.n2202 vdd.n2201 185
R842 vdd.n2204 vdd.n1180 185
R843 vdd.n2206 vdd.n2205 185
R844 vdd.n2207 vdd.n1175 185
R845 vdd.n2209 vdd.n2208 185
R846 vdd.n2211 vdd.n1173 185
R847 vdd.n2213 vdd.n2212 185
R848 vdd.n2214 vdd.n1169 185
R849 vdd.n2216 vdd.n2215 185
R850 vdd.n2218 vdd.n1166 185
R851 vdd.n2220 vdd.n2219 185
R852 vdd.n1167 vdd.n1160 185
R853 vdd.n2224 vdd.n1164 185
R854 vdd.n2225 vdd.n1156 185
R855 vdd.n2227 vdd.n2226 185
R856 vdd.n2229 vdd.n1154 185
R857 vdd.n2231 vdd.n2230 185
R858 vdd.n2232 vdd.n1149 185
R859 vdd.n2234 vdd.n2233 185
R860 vdd.n2236 vdd.n1147 185
R861 vdd.n2238 vdd.n2237 185
R862 vdd.n2239 vdd.n1142 185
R863 vdd.n2241 vdd.n2240 185
R864 vdd.n2243 vdd.n1140 185
R865 vdd.n2245 vdd.n2244 185
R866 vdd.n2246 vdd.n1135 185
R867 vdd.n2248 vdd.n2247 185
R868 vdd.n2250 vdd.n1133 185
R869 vdd.n2252 vdd.n2251 185
R870 vdd.n2253 vdd.n1129 185
R871 vdd.n2255 vdd.n2254 185
R872 vdd.n2257 vdd.n1126 185
R873 vdd.n2259 vdd.n2258 185
R874 vdd.n1127 vdd.n1120 185
R875 vdd.n2263 vdd.n1124 185
R876 vdd.n2264 vdd.n1116 185
R877 vdd.n2266 vdd.n2265 185
R878 vdd.n2268 vdd.n1114 185
R879 vdd.n2270 vdd.n2269 185
R880 vdd.n2271 vdd.n1109 185
R881 vdd.n2273 vdd.n2272 185
R882 vdd.n2275 vdd.n1107 185
R883 vdd.n2277 vdd.n2276 185
R884 vdd.n2278 vdd.n1102 185
R885 vdd.n2280 vdd.n2279 185
R886 vdd.n2282 vdd.n1100 185
R887 vdd.n2284 vdd.n2283 185
R888 vdd.n2285 vdd.n1098 185
R889 vdd.n2287 vdd.n2286 185
R890 vdd.n2290 vdd.n2289 185
R891 vdd.n2292 vdd.n2291 185
R892 vdd.n2294 vdd.n1096 185
R893 vdd.n2296 vdd.n2295 185
R894 vdd.n1409 vdd.n1095 185
R895 vdd.n2183 vdd.n1406 185
R896 vdd.n2183 vdd.n2182 185
R897 vdd.n1417 vdd.n1405 185
R898 vdd.n1407 vdd.n1405 185
R899 vdd.n2173 vdd.n2172 185
R900 vdd.n2174 vdd.n2173 185
R901 vdd.n1416 vdd.n1415 185
R902 vdd.n1415 vdd.n1414 185
R903 vdd.n2166 vdd.n2165 185
R904 vdd.n2165 vdd.n2164 185
R905 vdd.n1420 vdd.n1419 185
R906 vdd.n2155 vdd.n1420 185
R907 vdd.n2154 vdd.n2153 185
R908 vdd.n2156 vdd.n2154 185
R909 vdd.n1427 vdd.n1426 185
R910 vdd.n1431 vdd.n1426 185
R911 vdd.n2149 vdd.n2148 185
R912 vdd.n2148 vdd.n2147 185
R913 vdd.n1430 vdd.n1429 185
R914 vdd.n2138 vdd.n1430 185
R915 vdd.n2137 vdd.n2136 185
R916 vdd.n2139 vdd.n2137 185
R917 vdd.n1439 vdd.n1438 185
R918 vdd.n1438 vdd.n1437 185
R919 vdd.n2132 vdd.n2131 185
R920 vdd.n2131 vdd.n2130 185
R921 vdd.n1442 vdd.n1441 185
R922 vdd.n1443 vdd.n1442 185
R923 vdd.n2121 vdd.n2120 185
R924 vdd.n2122 vdd.n2121 185
R925 vdd.n1450 vdd.n1449 185
R926 vdd.n1454 vdd.n1449 185
R927 vdd.n2116 vdd.n2115 185
R928 vdd.n2115 vdd.n2114 185
R929 vdd.n1453 vdd.n1452 185
R930 vdd.n1810 vdd.n1453 185
R931 vdd.n1809 vdd.n1808 185
R932 vdd.n1811 vdd.n1809 185
R933 vdd.n1461 vdd.n1460 185
R934 vdd.n1466 vdd.n1460 185
R935 vdd.n1804 vdd.n1803 185
R936 vdd.n1803 vdd.n1802 185
R937 vdd.n1464 vdd.n1463 185
R938 vdd.n1465 vdd.n1464 185
R939 vdd.n1793 vdd.n1792 185
R940 vdd.n1794 vdd.n1793 185
R941 vdd.n1474 vdd.n1473 185
R942 vdd.n1473 vdd.n1472 185
R943 vdd.n1788 vdd.n1787 185
R944 vdd.n1787 vdd.n1786 185
R945 vdd.n1477 vdd.n1476 185
R946 vdd.n1777 vdd.n1477 185
R947 vdd.n1776 vdd.n1775 185
R948 vdd.n1778 vdd.n1776 185
R949 vdd.n1484 vdd.n1483 185
R950 vdd.n1488 vdd.n1483 185
R951 vdd.n1771 vdd.n1770 185
R952 vdd.n1770 vdd.n1769 185
R953 vdd.n1487 vdd.n1486 185
R954 vdd.n1760 vdd.n1487 185
R955 vdd.n1759 vdd.n1758 185
R956 vdd.n1761 vdd.n1759 185
R957 vdd.n1496 vdd.n1495 185
R958 vdd.n1495 vdd.n1494 185
R959 vdd.n1754 vdd.n1753 185
R960 vdd.n1753 vdd.n1752 185
R961 vdd.n1499 vdd.n1498 185
R962 vdd.n1500 vdd.n1499 185
R963 vdd.n1743 vdd.n1742 185
R964 vdd.n1744 vdd.n1743 185
R965 vdd.n1508 vdd.n1507 185
R966 vdd.n1507 vdd.n1506 185
R967 vdd.n942 vdd.n940 185
R968 vdd.n2510 vdd.n940 185
R969 vdd.n2432 vdd.n960 185
R970 vdd.n960 vdd.n947 185
R971 vdd.n2434 vdd.n2433 185
R972 vdd.n2435 vdd.n2434 185
R973 vdd.n2431 vdd.n959 185
R974 vdd.n1309 vdd.n959 185
R975 vdd.n2430 vdd.n2429 185
R976 vdd.n2429 vdd.n2428 185
R977 vdd.n962 vdd.n961 185
R978 vdd.n963 vdd.n962 185
R979 vdd.n2419 vdd.n2418 185
R980 vdd.n2420 vdd.n2419 185
R981 vdd.n2417 vdd.n973 185
R982 vdd.n973 vdd.n970 185
R983 vdd.n2416 vdd.n2415 185
R984 vdd.n2415 vdd.n2414 185
R985 vdd.n975 vdd.n974 185
R986 vdd.n976 vdd.n975 185
R987 vdd.n2407 vdd.n2406 185
R988 vdd.n2408 vdd.n2407 185
R989 vdd.n2405 vdd.n984 185
R990 vdd.n989 vdd.n984 185
R991 vdd.n2404 vdd.n2403 185
R992 vdd.n2403 vdd.n2402 185
R993 vdd.n986 vdd.n985 185
R994 vdd.n995 vdd.n986 185
R995 vdd.n2395 vdd.n2394 185
R996 vdd.n2396 vdd.n2395 185
R997 vdd.n2393 vdd.n996 185
R998 vdd.n1330 vdd.n996 185
R999 vdd.n2392 vdd.n2391 185
R1000 vdd.n2391 vdd.n2390 185
R1001 vdd.n998 vdd.n997 185
R1002 vdd.n999 vdd.n998 185
R1003 vdd.n2383 vdd.n2382 185
R1004 vdd.n2384 vdd.n2383 185
R1005 vdd.n2381 vdd.n1008 185
R1006 vdd.n1008 vdd.n1005 185
R1007 vdd.n2380 vdd.n2379 185
R1008 vdd.n2379 vdd.n2378 185
R1009 vdd.n1010 vdd.n1009 185
R1010 vdd.n1019 vdd.n1010 185
R1011 vdd.n2370 vdd.n2369 185
R1012 vdd.n2371 vdd.n2370 185
R1013 vdd.n2368 vdd.n1020 185
R1014 vdd.n1026 vdd.n1020 185
R1015 vdd.n2367 vdd.n2366 185
R1016 vdd.n2366 vdd.n2365 185
R1017 vdd.n1022 vdd.n1021 185
R1018 vdd.n1023 vdd.n1022 185
R1019 vdd.n2358 vdd.n2357 185
R1020 vdd.n2359 vdd.n2358 185
R1021 vdd.n2356 vdd.n1033 185
R1022 vdd.n1033 vdd.n1030 185
R1023 vdd.n2355 vdd.n2354 185
R1024 vdd.n2354 vdd.n2353 185
R1025 vdd.n1035 vdd.n1034 185
R1026 vdd.n1036 vdd.n1035 185
R1027 vdd.n2346 vdd.n2345 185
R1028 vdd.n2347 vdd.n2346 185
R1029 vdd.n2344 vdd.n1044 185
R1030 vdd.n1050 vdd.n1044 185
R1031 vdd.n2343 vdd.n2342 185
R1032 vdd.n2342 vdd.n2341 185
R1033 vdd.n1046 vdd.n1045 185
R1034 vdd.n1047 vdd.n1046 185
R1035 vdd.n2332 vdd.n2331 185
R1036 vdd.n2330 vdd.n1089 185
R1037 vdd.n2329 vdd.n1088 185
R1038 vdd.n2334 vdd.n1088 185
R1039 vdd.n2328 vdd.n2327 185
R1040 vdd.n2326 vdd.n2325 185
R1041 vdd.n2324 vdd.n2323 185
R1042 vdd.n2322 vdd.n2321 185
R1043 vdd.n2320 vdd.n2319 185
R1044 vdd.n2318 vdd.n2317 185
R1045 vdd.n2316 vdd.n2315 185
R1046 vdd.n2314 vdd.n2313 185
R1047 vdd.n2312 vdd.n2311 185
R1048 vdd.n2310 vdd.n2309 185
R1049 vdd.n2308 vdd.n2307 185
R1050 vdd.n2306 vdd.n2305 185
R1051 vdd.n2304 vdd.n2303 185
R1052 vdd.n2302 vdd.n2301 185
R1053 vdd.n2300 vdd.n2299 185
R1054 vdd.n1246 vdd.n1090 185
R1055 vdd.n1248 vdd.n1247 185
R1056 vdd.n1250 vdd.n1249 185
R1057 vdd.n1252 vdd.n1251 185
R1058 vdd.n1254 vdd.n1253 185
R1059 vdd.n1256 vdd.n1255 185
R1060 vdd.n1258 vdd.n1257 185
R1061 vdd.n1260 vdd.n1259 185
R1062 vdd.n1262 vdd.n1261 185
R1063 vdd.n1264 vdd.n1263 185
R1064 vdd.n1266 vdd.n1265 185
R1065 vdd.n1268 vdd.n1267 185
R1066 vdd.n1270 vdd.n1269 185
R1067 vdd.n1272 vdd.n1271 185
R1068 vdd.n1275 vdd.n1274 185
R1069 vdd.n1277 vdd.n1276 185
R1070 vdd.n1279 vdd.n1278 185
R1071 vdd.n2513 vdd.n2512 185
R1072 vdd.n2515 vdd.n2514 185
R1073 vdd.n2517 vdd.n2516 185
R1074 vdd.n2520 vdd.n2519 185
R1075 vdd.n2522 vdd.n2521 185
R1076 vdd.n2524 vdd.n2523 185
R1077 vdd.n2526 vdd.n2525 185
R1078 vdd.n2528 vdd.n2527 185
R1079 vdd.n2530 vdd.n2529 185
R1080 vdd.n2532 vdd.n2531 185
R1081 vdd.n2534 vdd.n2533 185
R1082 vdd.n2536 vdd.n2535 185
R1083 vdd.n2538 vdd.n2537 185
R1084 vdd.n2540 vdd.n2539 185
R1085 vdd.n2542 vdd.n2541 185
R1086 vdd.n2544 vdd.n2543 185
R1087 vdd.n2546 vdd.n2545 185
R1088 vdd.n2548 vdd.n2547 185
R1089 vdd.n2550 vdd.n2549 185
R1090 vdd.n2552 vdd.n2551 185
R1091 vdd.n2554 vdd.n2553 185
R1092 vdd.n2556 vdd.n2555 185
R1093 vdd.n2558 vdd.n2557 185
R1094 vdd.n2560 vdd.n2559 185
R1095 vdd.n2562 vdd.n2561 185
R1096 vdd.n2564 vdd.n2563 185
R1097 vdd.n2566 vdd.n2565 185
R1098 vdd.n2568 vdd.n2567 185
R1099 vdd.n2570 vdd.n2569 185
R1100 vdd.n2572 vdd.n2571 185
R1101 vdd.n2574 vdd.n2573 185
R1102 vdd.n2576 vdd.n2575 185
R1103 vdd.n2578 vdd.n2577 185
R1104 vdd.n2579 vdd.n941 185
R1105 vdd.n2581 vdd.n2580 185
R1106 vdd.n2582 vdd.n2581 185
R1107 vdd.n2511 vdd.n945 185
R1108 vdd.n2511 vdd.n2510 185
R1109 vdd.n1307 vdd.n946 185
R1110 vdd.n947 vdd.n946 185
R1111 vdd.n1308 vdd.n957 185
R1112 vdd.n2435 vdd.n957 185
R1113 vdd.n1311 vdd.n1310 185
R1114 vdd.n1310 vdd.n1309 185
R1115 vdd.n1312 vdd.n964 185
R1116 vdd.n2428 vdd.n964 185
R1117 vdd.n1314 vdd.n1313 185
R1118 vdd.n1313 vdd.n963 185
R1119 vdd.n1315 vdd.n971 185
R1120 vdd.n2420 vdd.n971 185
R1121 vdd.n1317 vdd.n1316 185
R1122 vdd.n1316 vdd.n970 185
R1123 vdd.n1318 vdd.n977 185
R1124 vdd.n2414 vdd.n977 185
R1125 vdd.n1320 vdd.n1319 185
R1126 vdd.n1319 vdd.n976 185
R1127 vdd.n1321 vdd.n982 185
R1128 vdd.n2408 vdd.n982 185
R1129 vdd.n1323 vdd.n1322 185
R1130 vdd.n1322 vdd.n989 185
R1131 vdd.n1324 vdd.n987 185
R1132 vdd.n2402 vdd.n987 185
R1133 vdd.n1326 vdd.n1325 185
R1134 vdd.n1325 vdd.n995 185
R1135 vdd.n1327 vdd.n993 185
R1136 vdd.n2396 vdd.n993 185
R1137 vdd.n1329 vdd.n1328 185
R1138 vdd.n1330 vdd.n1329 185
R1139 vdd.n1306 vdd.n1000 185
R1140 vdd.n2390 vdd.n1000 185
R1141 vdd.n1305 vdd.n1304 185
R1142 vdd.n1304 vdd.n999 185
R1143 vdd.n1303 vdd.n1006 185
R1144 vdd.n2384 vdd.n1006 185
R1145 vdd.n1302 vdd.n1301 185
R1146 vdd.n1301 vdd.n1005 185
R1147 vdd.n1300 vdd.n1011 185
R1148 vdd.n2378 vdd.n1011 185
R1149 vdd.n1299 vdd.n1298 185
R1150 vdd.n1298 vdd.n1019 185
R1151 vdd.n1297 vdd.n1017 185
R1152 vdd.n2371 vdd.n1017 185
R1153 vdd.n1296 vdd.n1295 185
R1154 vdd.n1295 vdd.n1026 185
R1155 vdd.n1294 vdd.n1024 185
R1156 vdd.n2365 vdd.n1024 185
R1157 vdd.n1293 vdd.n1292 185
R1158 vdd.n1292 vdd.n1023 185
R1159 vdd.n1291 vdd.n1031 185
R1160 vdd.n2359 vdd.n1031 185
R1161 vdd.n1290 vdd.n1289 185
R1162 vdd.n1289 vdd.n1030 185
R1163 vdd.n1288 vdd.n1037 185
R1164 vdd.n2353 vdd.n1037 185
R1165 vdd.n1287 vdd.n1286 185
R1166 vdd.n1286 vdd.n1036 185
R1167 vdd.n1285 vdd.n1042 185
R1168 vdd.n2347 vdd.n1042 185
R1169 vdd.n1284 vdd.n1283 185
R1170 vdd.n1283 vdd.n1050 185
R1171 vdd.n1282 vdd.n1048 185
R1172 vdd.n2341 vdd.n1048 185
R1173 vdd.n1281 vdd.n1280 185
R1174 vdd.n1280 vdd.n1047 185
R1175 vdd.n370 vdd.n369 185
R1176 vdd.n3346 vdd.n370 185
R1177 vdd.n3349 vdd.n3348 185
R1178 vdd.n3348 vdd.n3347 185
R1179 vdd.n3350 vdd.n364 185
R1180 vdd.n364 vdd.n363 185
R1181 vdd.n3352 vdd.n3351 185
R1182 vdd.n3353 vdd.n3352 185
R1183 vdd.n359 vdd.n358 185
R1184 vdd.n3354 vdd.n359 185
R1185 vdd.n3357 vdd.n3356 185
R1186 vdd.n3356 vdd.n3355 185
R1187 vdd.n3358 vdd.n353 185
R1188 vdd.n3328 vdd.n353 185
R1189 vdd.n3360 vdd.n3359 185
R1190 vdd.n3361 vdd.n3360 185
R1191 vdd.n348 vdd.n347 185
R1192 vdd.n3362 vdd.n348 185
R1193 vdd.n3365 vdd.n3364 185
R1194 vdd.n3364 vdd.n3363 185
R1195 vdd.n3366 vdd.n342 185
R1196 vdd.n349 vdd.n342 185
R1197 vdd.n3368 vdd.n3367 185
R1198 vdd.n3369 vdd.n3368 185
R1199 vdd.n338 vdd.n337 185
R1200 vdd.n3370 vdd.n338 185
R1201 vdd.n3373 vdd.n3372 185
R1202 vdd.n3372 vdd.n3371 185
R1203 vdd.n3374 vdd.n333 185
R1204 vdd.n333 vdd.n332 185
R1205 vdd.n3376 vdd.n3375 185
R1206 vdd.n3377 vdd.n3376 185
R1207 vdd.n327 vdd.n325 185
R1208 vdd.n3378 vdd.n327 185
R1209 vdd.n3381 vdd.n3380 185
R1210 vdd.n3380 vdd.n3379 185
R1211 vdd.n326 vdd.n324 185
R1212 vdd.n328 vdd.n326 185
R1213 vdd.n3304 vdd.n3303 185
R1214 vdd.n3305 vdd.n3304 185
R1215 vdd.n615 vdd.n614 185
R1216 vdd.n614 vdd.n613 185
R1217 vdd.n3299 vdd.n3298 185
R1218 vdd.n3298 vdd.n3297 185
R1219 vdd.n618 vdd.n617 185
R1220 vdd.n624 vdd.n618 185
R1221 vdd.n3285 vdd.n3284 185
R1222 vdd.n3286 vdd.n3285 185
R1223 vdd.n626 vdd.n625 185
R1224 vdd.n3277 vdd.n625 185
R1225 vdd.n3280 vdd.n3279 185
R1226 vdd.n3279 vdd.n3278 185
R1227 vdd.n629 vdd.n628 185
R1228 vdd.n636 vdd.n629 185
R1229 vdd.n3268 vdd.n3267 185
R1230 vdd.n3269 vdd.n3268 185
R1231 vdd.n638 vdd.n637 185
R1232 vdd.n637 vdd.n635 185
R1233 vdd.n3263 vdd.n3262 185
R1234 vdd.n3262 vdd.n3261 185
R1235 vdd.n641 vdd.n640 185
R1236 vdd.n642 vdd.n641 185
R1237 vdd.n3252 vdd.n3251 185
R1238 vdd.n3253 vdd.n3252 185
R1239 vdd.n650 vdd.n649 185
R1240 vdd.n649 vdd.n648 185
R1241 vdd.n3247 vdd.n3246 185
R1242 vdd.n3246 vdd.n3245 185
R1243 vdd.n653 vdd.n652 185
R1244 vdd.n659 vdd.n653 185
R1245 vdd.n3236 vdd.n3235 185
R1246 vdd.n3237 vdd.n3236 185
R1247 vdd.n3232 vdd.n660 185
R1248 vdd.n3231 vdd.n3230 185
R1249 vdd.n3228 vdd.n662 185
R1250 vdd.n3228 vdd.n658 185
R1251 vdd.n3227 vdd.n3226 185
R1252 vdd.n3225 vdd.n3224 185
R1253 vdd.n3223 vdd.n3222 185
R1254 vdd.n3221 vdd.n3220 185
R1255 vdd.n3219 vdd.n668 185
R1256 vdd.n3217 vdd.n3216 185
R1257 vdd.n3215 vdd.n669 185
R1258 vdd.n3214 vdd.n3213 185
R1259 vdd.n3211 vdd.n674 185
R1260 vdd.n3209 vdd.n3208 185
R1261 vdd.n3207 vdd.n675 185
R1262 vdd.n3206 vdd.n3205 185
R1263 vdd.n3203 vdd.n680 185
R1264 vdd.n3201 vdd.n3200 185
R1265 vdd.n3199 vdd.n681 185
R1266 vdd.n3198 vdd.n3197 185
R1267 vdd.n3195 vdd.n688 185
R1268 vdd.n3193 vdd.n3192 185
R1269 vdd.n3191 vdd.n689 185
R1270 vdd.n3190 vdd.n3189 185
R1271 vdd.n3187 vdd.n694 185
R1272 vdd.n3185 vdd.n3184 185
R1273 vdd.n3183 vdd.n695 185
R1274 vdd.n3182 vdd.n3181 185
R1275 vdd.n3179 vdd.n700 185
R1276 vdd.n3177 vdd.n3176 185
R1277 vdd.n3175 vdd.n701 185
R1278 vdd.n3174 vdd.n3173 185
R1279 vdd.n3171 vdd.n706 185
R1280 vdd.n3169 vdd.n3168 185
R1281 vdd.n3167 vdd.n707 185
R1282 vdd.n3166 vdd.n3165 185
R1283 vdd.n3163 vdd.n712 185
R1284 vdd.n3161 vdd.n3160 185
R1285 vdd.n3159 vdd.n713 185
R1286 vdd.n3158 vdd.n3157 185
R1287 vdd.n3155 vdd.n718 185
R1288 vdd.n3153 vdd.n3152 185
R1289 vdd.n3151 vdd.n719 185
R1290 vdd.n728 vdd.n722 185
R1291 vdd.n3147 vdd.n3146 185
R1292 vdd.n3144 vdd.n726 185
R1293 vdd.n3143 vdd.n3142 185
R1294 vdd.n3141 vdd.n3140 185
R1295 vdd.n3139 vdd.n732 185
R1296 vdd.n3137 vdd.n3136 185
R1297 vdd.n3135 vdd.n733 185
R1298 vdd.n3134 vdd.n3133 185
R1299 vdd.n3131 vdd.n738 185
R1300 vdd.n3129 vdd.n3128 185
R1301 vdd.n3127 vdd.n739 185
R1302 vdd.n3126 vdd.n3125 185
R1303 vdd.n3123 vdd.n744 185
R1304 vdd.n3121 vdd.n3120 185
R1305 vdd.n3119 vdd.n745 185
R1306 vdd.n3118 vdd.n3117 185
R1307 vdd.n3115 vdd.n3114 185
R1308 vdd.n3113 vdd.n3112 185
R1309 vdd.n3111 vdd.n3110 185
R1310 vdd.n3109 vdd.n3108 185
R1311 vdd.n3104 vdd.n657 185
R1312 vdd.n658 vdd.n657 185
R1313 vdd.n3343 vdd.n3342 185
R1314 vdd.n599 vdd.n404 185
R1315 vdd.n598 vdd.n597 185
R1316 vdd.n596 vdd.n595 185
R1317 vdd.n594 vdd.n409 185
R1318 vdd.n590 vdd.n589 185
R1319 vdd.n588 vdd.n587 185
R1320 vdd.n586 vdd.n585 185
R1321 vdd.n584 vdd.n411 185
R1322 vdd.n580 vdd.n579 185
R1323 vdd.n578 vdd.n577 185
R1324 vdd.n576 vdd.n575 185
R1325 vdd.n574 vdd.n413 185
R1326 vdd.n570 vdd.n569 185
R1327 vdd.n568 vdd.n567 185
R1328 vdd.n566 vdd.n565 185
R1329 vdd.n564 vdd.n415 185
R1330 vdd.n560 vdd.n559 185
R1331 vdd.n558 vdd.n557 185
R1332 vdd.n556 vdd.n555 185
R1333 vdd.n554 vdd.n417 185
R1334 vdd.n550 vdd.n549 185
R1335 vdd.n548 vdd.n547 185
R1336 vdd.n546 vdd.n545 185
R1337 vdd.n544 vdd.n421 185
R1338 vdd.n540 vdd.n539 185
R1339 vdd.n538 vdd.n537 185
R1340 vdd.n536 vdd.n535 185
R1341 vdd.n534 vdd.n423 185
R1342 vdd.n530 vdd.n529 185
R1343 vdd.n528 vdd.n527 185
R1344 vdd.n526 vdd.n525 185
R1345 vdd.n524 vdd.n425 185
R1346 vdd.n520 vdd.n519 185
R1347 vdd.n518 vdd.n517 185
R1348 vdd.n516 vdd.n515 185
R1349 vdd.n514 vdd.n427 185
R1350 vdd.n510 vdd.n509 185
R1351 vdd.n508 vdd.n507 185
R1352 vdd.n506 vdd.n505 185
R1353 vdd.n504 vdd.n429 185
R1354 vdd.n500 vdd.n499 185
R1355 vdd.n498 vdd.n497 185
R1356 vdd.n496 vdd.n495 185
R1357 vdd.n494 vdd.n433 185
R1358 vdd.n490 vdd.n489 185
R1359 vdd.n488 vdd.n487 185
R1360 vdd.n486 vdd.n485 185
R1361 vdd.n484 vdd.n435 185
R1362 vdd.n480 vdd.n479 185
R1363 vdd.n478 vdd.n477 185
R1364 vdd.n476 vdd.n475 185
R1365 vdd.n474 vdd.n437 185
R1366 vdd.n470 vdd.n469 185
R1367 vdd.n468 vdd.n467 185
R1368 vdd.n466 vdd.n465 185
R1369 vdd.n464 vdd.n439 185
R1370 vdd.n460 vdd.n459 185
R1371 vdd.n458 vdd.n457 185
R1372 vdd.n456 vdd.n455 185
R1373 vdd.n454 vdd.n441 185
R1374 vdd.n450 vdd.n449 185
R1375 vdd.n448 vdd.n447 185
R1376 vdd.n446 vdd.n445 185
R1377 vdd.n3339 vdd.n372 185
R1378 vdd.n3346 vdd.n372 185
R1379 vdd.n3338 vdd.n371 185
R1380 vdd.n3347 vdd.n371 185
R1381 vdd.n3337 vdd.n3336 185
R1382 vdd.n3336 vdd.n363 185
R1383 vdd.n602 vdd.n362 185
R1384 vdd.n3353 vdd.n362 185
R1385 vdd.n3332 vdd.n361 185
R1386 vdd.n3354 vdd.n361 185
R1387 vdd.n3331 vdd.n360 185
R1388 vdd.n3355 vdd.n360 185
R1389 vdd.n3330 vdd.n3329 185
R1390 vdd.n3329 vdd.n3328 185
R1391 vdd.n604 vdd.n352 185
R1392 vdd.n3361 vdd.n352 185
R1393 vdd.n3324 vdd.n351 185
R1394 vdd.n3362 vdd.n351 185
R1395 vdd.n3323 vdd.n350 185
R1396 vdd.n3363 vdd.n350 185
R1397 vdd.n3322 vdd.n3321 185
R1398 vdd.n3321 vdd.n349 185
R1399 vdd.n606 vdd.n341 185
R1400 vdd.n3369 vdd.n341 185
R1401 vdd.n3317 vdd.n340 185
R1402 vdd.n3370 vdd.n340 185
R1403 vdd.n3316 vdd.n339 185
R1404 vdd.n3371 vdd.n339 185
R1405 vdd.n3315 vdd.n3314 185
R1406 vdd.n3314 vdd.n332 185
R1407 vdd.n608 vdd.n331 185
R1408 vdd.n3377 vdd.n331 185
R1409 vdd.n3310 vdd.n330 185
R1410 vdd.n3378 vdd.n330 185
R1411 vdd.n3309 vdd.n329 185
R1412 vdd.n3379 vdd.n329 185
R1413 vdd.n3308 vdd.n3307 185
R1414 vdd.n3307 vdd.n328 185
R1415 vdd.n3306 vdd.n610 185
R1416 vdd.n3306 vdd.n3305 185
R1417 vdd.n3294 vdd.n612 185
R1418 vdd.n613 vdd.n612 185
R1419 vdd.n3296 vdd.n3295 185
R1420 vdd.n3297 vdd.n3296 185
R1421 vdd.n620 vdd.n619 185
R1422 vdd.n624 vdd.n619 185
R1423 vdd.n3288 vdd.n3287 185
R1424 vdd.n3287 vdd.n3286 185
R1425 vdd.n623 vdd.n622 185
R1426 vdd.n3277 vdd.n623 185
R1427 vdd.n3276 vdd.n3275 185
R1428 vdd.n3278 vdd.n3276 185
R1429 vdd.n631 vdd.n630 185
R1430 vdd.n636 vdd.n630 185
R1431 vdd.n3271 vdd.n3270 185
R1432 vdd.n3270 vdd.n3269 185
R1433 vdd.n634 vdd.n633 185
R1434 vdd.n635 vdd.n634 185
R1435 vdd.n3260 vdd.n3259 185
R1436 vdd.n3261 vdd.n3260 185
R1437 vdd.n644 vdd.n643 185
R1438 vdd.n643 vdd.n642 185
R1439 vdd.n3255 vdd.n3254 185
R1440 vdd.n3254 vdd.n3253 185
R1441 vdd.n647 vdd.n646 185
R1442 vdd.n648 vdd.n647 185
R1443 vdd.n3244 vdd.n3243 185
R1444 vdd.n3245 vdd.n3244 185
R1445 vdd.n655 vdd.n654 185
R1446 vdd.n659 vdd.n654 185
R1447 vdd.n3239 vdd.n3238 185
R1448 vdd.n3238 vdd.n3237 185
R1449 vdd.n2853 vdd.n2852 185
R1450 vdd.n2851 vdd.n2617 185
R1451 vdd.n2850 vdd.n2616 185
R1452 vdd.n2855 vdd.n2616 185
R1453 vdd.n2849 vdd.n2848 185
R1454 vdd.n2847 vdd.n2846 185
R1455 vdd.n2845 vdd.n2844 185
R1456 vdd.n2843 vdd.n2842 185
R1457 vdd.n2841 vdd.n2840 185
R1458 vdd.n2839 vdd.n2838 185
R1459 vdd.n2837 vdd.n2836 185
R1460 vdd.n2835 vdd.n2834 185
R1461 vdd.n2833 vdd.n2832 185
R1462 vdd.n2831 vdd.n2830 185
R1463 vdd.n2829 vdd.n2828 185
R1464 vdd.n2827 vdd.n2826 185
R1465 vdd.n2825 vdd.n2824 185
R1466 vdd.n2823 vdd.n2822 185
R1467 vdd.n2821 vdd.n2820 185
R1468 vdd.n2819 vdd.n2818 185
R1469 vdd.n2817 vdd.n2816 185
R1470 vdd.n2815 vdd.n2814 185
R1471 vdd.n2813 vdd.n2812 185
R1472 vdd.n2811 vdd.n2810 185
R1473 vdd.n2809 vdd.n2808 185
R1474 vdd.n2807 vdd.n2806 185
R1475 vdd.n2805 vdd.n2804 185
R1476 vdd.n2803 vdd.n2802 185
R1477 vdd.n2801 vdd.n2800 185
R1478 vdd.n2799 vdd.n2798 185
R1479 vdd.n2797 vdd.n2796 185
R1480 vdd.n2795 vdd.n2794 185
R1481 vdd.n2793 vdd.n2792 185
R1482 vdd.n2790 vdd.n2789 185
R1483 vdd.n2788 vdd.n2787 185
R1484 vdd.n2786 vdd.n2785 185
R1485 vdd.n3005 vdd.n3004 185
R1486 vdd.n3006 vdd.n803 185
R1487 vdd.n3008 vdd.n3007 185
R1488 vdd.n3010 vdd.n801 185
R1489 vdd.n3012 vdd.n3011 185
R1490 vdd.n3013 vdd.n800 185
R1491 vdd.n3015 vdd.n3014 185
R1492 vdd.n3017 vdd.n798 185
R1493 vdd.n3019 vdd.n3018 185
R1494 vdd.n3020 vdd.n797 185
R1495 vdd.n3022 vdd.n3021 185
R1496 vdd.n3024 vdd.n795 185
R1497 vdd.n3026 vdd.n3025 185
R1498 vdd.n3027 vdd.n794 185
R1499 vdd.n3029 vdd.n3028 185
R1500 vdd.n3031 vdd.n792 185
R1501 vdd.n3033 vdd.n3032 185
R1502 vdd.n3035 vdd.n791 185
R1503 vdd.n3037 vdd.n3036 185
R1504 vdd.n3039 vdd.n789 185
R1505 vdd.n3041 vdd.n3040 185
R1506 vdd.n3042 vdd.n788 185
R1507 vdd.n3044 vdd.n3043 185
R1508 vdd.n3046 vdd.n786 185
R1509 vdd.n3048 vdd.n3047 185
R1510 vdd.n3049 vdd.n785 185
R1511 vdd.n3051 vdd.n3050 185
R1512 vdd.n3053 vdd.n783 185
R1513 vdd.n3055 vdd.n3054 185
R1514 vdd.n3056 vdd.n782 185
R1515 vdd.n3058 vdd.n3057 185
R1516 vdd.n3060 vdd.n781 185
R1517 vdd.n3061 vdd.n780 185
R1518 vdd.n3064 vdd.n3063 185
R1519 vdd.n3065 vdd.n778 185
R1520 vdd.n778 vdd.n756 185
R1521 vdd.n3002 vdd.n775 185
R1522 vdd.n3068 vdd.n775 185
R1523 vdd.n3001 vdd.n3000 185
R1524 vdd.n3000 vdd.n774 185
R1525 vdd.n2999 vdd.n807 185
R1526 vdd.n2999 vdd.n2998 185
R1527 vdd.n2733 vdd.n808 185
R1528 vdd.n817 vdd.n808 185
R1529 vdd.n2734 vdd.n815 185
R1530 vdd.n2992 vdd.n815 185
R1531 vdd.n2736 vdd.n2735 185
R1532 vdd.n2735 vdd.n814 185
R1533 vdd.n2737 vdd.n823 185
R1534 vdd.n2941 vdd.n823 185
R1535 vdd.n2739 vdd.n2738 185
R1536 vdd.n2738 vdd.n822 185
R1537 vdd.n2740 vdd.n829 185
R1538 vdd.n2935 vdd.n829 185
R1539 vdd.n2742 vdd.n2741 185
R1540 vdd.n2741 vdd.n828 185
R1541 vdd.n2743 vdd.n834 185
R1542 vdd.n2929 vdd.n834 185
R1543 vdd.n2745 vdd.n2744 185
R1544 vdd.n2744 vdd.n841 185
R1545 vdd.n2746 vdd.n839 185
R1546 vdd.n2923 vdd.n839 185
R1547 vdd.n2748 vdd.n2747 185
R1548 vdd.n2747 vdd.n849 185
R1549 vdd.n2749 vdd.n847 185
R1550 vdd.n2916 vdd.n847 185
R1551 vdd.n2751 vdd.n2750 185
R1552 vdd.n2750 vdd.n846 185
R1553 vdd.n2752 vdd.n854 185
R1554 vdd.n2910 vdd.n854 185
R1555 vdd.n2754 vdd.n2753 185
R1556 vdd.n2753 vdd.n853 185
R1557 vdd.n2755 vdd.n859 185
R1558 vdd.n2904 vdd.n859 185
R1559 vdd.n2757 vdd.n2756 185
R1560 vdd.n2756 vdd.n866 185
R1561 vdd.n2758 vdd.n864 185
R1562 vdd.n2898 vdd.n864 185
R1563 vdd.n2760 vdd.n2759 185
R1564 vdd.n2759 vdd.n872 185
R1565 vdd.n2761 vdd.n870 185
R1566 vdd.n2892 vdd.n870 185
R1567 vdd.n2763 vdd.n2762 185
R1568 vdd.n2764 vdd.n2763 185
R1569 vdd.n2732 vdd.n877 185
R1570 vdd.n2886 vdd.n877 185
R1571 vdd.n2731 vdd.n2730 185
R1572 vdd.n2730 vdd.n876 185
R1573 vdd.n2729 vdd.n883 185
R1574 vdd.n2880 vdd.n883 185
R1575 vdd.n2728 vdd.n2727 185
R1576 vdd.n2727 vdd.n882 185
R1577 vdd.n2726 vdd.n889 185
R1578 vdd.n2874 vdd.n889 185
R1579 vdd.n2725 vdd.n2724 185
R1580 vdd.n2724 vdd.n888 185
R1581 vdd.n2620 vdd.n894 185
R1582 vdd.n2868 vdd.n894 185
R1583 vdd.n2781 vdd.n2780 185
R1584 vdd.n2780 vdd.n2779 185
R1585 vdd.n2782 vdd.n900 185
R1586 vdd.n2862 vdd.n900 185
R1587 vdd.n2784 vdd.n2783 185
R1588 vdd.n2784 vdd.n899 185
R1589 vdd.n898 vdd.n897 185
R1590 vdd.n899 vdd.n898 185
R1591 vdd.n2864 vdd.n2863 185
R1592 vdd.n2863 vdd.n2862 185
R1593 vdd.n2865 vdd.n896 185
R1594 vdd.n2779 vdd.n896 185
R1595 vdd.n2867 vdd.n2866 185
R1596 vdd.n2868 vdd.n2867 185
R1597 vdd.n887 vdd.n886 185
R1598 vdd.n888 vdd.n887 185
R1599 vdd.n2876 vdd.n2875 185
R1600 vdd.n2875 vdd.n2874 185
R1601 vdd.n2877 vdd.n885 185
R1602 vdd.n885 vdd.n882 185
R1603 vdd.n2879 vdd.n2878 185
R1604 vdd.n2880 vdd.n2879 185
R1605 vdd.n875 vdd.n874 185
R1606 vdd.n876 vdd.n875 185
R1607 vdd.n2888 vdd.n2887 185
R1608 vdd.n2887 vdd.n2886 185
R1609 vdd.n2889 vdd.n873 185
R1610 vdd.n2764 vdd.n873 185
R1611 vdd.n2891 vdd.n2890 185
R1612 vdd.n2892 vdd.n2891 185
R1613 vdd.n863 vdd.n862 185
R1614 vdd.n872 vdd.n863 185
R1615 vdd.n2900 vdd.n2899 185
R1616 vdd.n2899 vdd.n2898 185
R1617 vdd.n2901 vdd.n861 185
R1618 vdd.n866 vdd.n861 185
R1619 vdd.n2903 vdd.n2902 185
R1620 vdd.n2904 vdd.n2903 185
R1621 vdd.n852 vdd.n851 185
R1622 vdd.n853 vdd.n852 185
R1623 vdd.n2912 vdd.n2911 185
R1624 vdd.n2911 vdd.n2910 185
R1625 vdd.n2913 vdd.n850 185
R1626 vdd.n850 vdd.n846 185
R1627 vdd.n2915 vdd.n2914 185
R1628 vdd.n2916 vdd.n2915 185
R1629 vdd.n838 vdd.n837 185
R1630 vdd.n849 vdd.n838 185
R1631 vdd.n2925 vdd.n2924 185
R1632 vdd.n2924 vdd.n2923 185
R1633 vdd.n2926 vdd.n836 185
R1634 vdd.n841 vdd.n836 185
R1635 vdd.n2928 vdd.n2927 185
R1636 vdd.n2929 vdd.n2928 185
R1637 vdd.n827 vdd.n826 185
R1638 vdd.n828 vdd.n827 185
R1639 vdd.n2937 vdd.n2936 185
R1640 vdd.n2936 vdd.n2935 185
R1641 vdd.n2938 vdd.n825 185
R1642 vdd.n825 vdd.n822 185
R1643 vdd.n2940 vdd.n2939 185
R1644 vdd.n2941 vdd.n2940 185
R1645 vdd.n813 vdd.n812 185
R1646 vdd.n814 vdd.n813 185
R1647 vdd.n2994 vdd.n2993 185
R1648 vdd.n2993 vdd.n2992 185
R1649 vdd.n2995 vdd.n811 185
R1650 vdd.n817 vdd.n811 185
R1651 vdd.n2997 vdd.n2996 185
R1652 vdd.n2998 vdd.n2997 185
R1653 vdd.n779 vdd.n777 185
R1654 vdd.n777 vdd.n774 185
R1655 vdd.n3067 vdd.n3066 185
R1656 vdd.n3068 vdd.n3067 185
R1657 vdd.n2509 vdd.n2508 185
R1658 vdd.n2510 vdd.n2509 185
R1659 vdd.n951 vdd.n949 185
R1660 vdd.n949 vdd.n947 185
R1661 vdd.n2424 vdd.n958 185
R1662 vdd.n2435 vdd.n958 185
R1663 vdd.n2425 vdd.n967 185
R1664 vdd.n1309 vdd.n967 185
R1665 vdd.n2427 vdd.n2426 185
R1666 vdd.n2428 vdd.n2427 185
R1667 vdd.n2423 vdd.n966 185
R1668 vdd.n966 vdd.n963 185
R1669 vdd.n2422 vdd.n2421 185
R1670 vdd.n2421 vdd.n2420 185
R1671 vdd.n969 vdd.n968 185
R1672 vdd.n970 vdd.n969 185
R1673 vdd.n2413 vdd.n2412 185
R1674 vdd.n2414 vdd.n2413 185
R1675 vdd.n2411 vdd.n979 185
R1676 vdd.n979 vdd.n976 185
R1677 vdd.n2410 vdd.n2409 185
R1678 vdd.n2409 vdd.n2408 185
R1679 vdd.n981 vdd.n980 185
R1680 vdd.n989 vdd.n981 185
R1681 vdd.n2401 vdd.n2400 185
R1682 vdd.n2402 vdd.n2401 185
R1683 vdd.n2399 vdd.n990 185
R1684 vdd.n995 vdd.n990 185
R1685 vdd.n2398 vdd.n2397 185
R1686 vdd.n2397 vdd.n2396 185
R1687 vdd.n992 vdd.n991 185
R1688 vdd.n1330 vdd.n992 185
R1689 vdd.n2389 vdd.n2388 185
R1690 vdd.n2390 vdd.n2389 185
R1691 vdd.n2387 vdd.n1002 185
R1692 vdd.n1002 vdd.n999 185
R1693 vdd.n2386 vdd.n2385 185
R1694 vdd.n2385 vdd.n2384 185
R1695 vdd.n1004 vdd.n1003 185
R1696 vdd.n1005 vdd.n1004 185
R1697 vdd.n2377 vdd.n2376 185
R1698 vdd.n2378 vdd.n2377 185
R1699 vdd.n2374 vdd.n1013 185
R1700 vdd.n1019 vdd.n1013 185
R1701 vdd.n2373 vdd.n2372 185
R1702 vdd.n2372 vdd.n2371 185
R1703 vdd.n1016 vdd.n1015 185
R1704 vdd.n1026 vdd.n1016 185
R1705 vdd.n2364 vdd.n2363 185
R1706 vdd.n2365 vdd.n2364 185
R1707 vdd.n2362 vdd.n1027 185
R1708 vdd.n1027 vdd.n1023 185
R1709 vdd.n2361 vdd.n2360 185
R1710 vdd.n2360 vdd.n2359 185
R1711 vdd.n1029 vdd.n1028 185
R1712 vdd.n1030 vdd.n1029 185
R1713 vdd.n2352 vdd.n2351 185
R1714 vdd.n2353 vdd.n2352 185
R1715 vdd.n2350 vdd.n1039 185
R1716 vdd.n1039 vdd.n1036 185
R1717 vdd.n2349 vdd.n2348 185
R1718 vdd.n2348 vdd.n2347 185
R1719 vdd.n1041 vdd.n1040 185
R1720 vdd.n1050 vdd.n1041 185
R1721 vdd.n2340 vdd.n2339 185
R1722 vdd.n2341 vdd.n2340 185
R1723 vdd.n2338 vdd.n1051 185
R1724 vdd.n1051 vdd.n1047 185
R1725 vdd.n2440 vdd.n922 185
R1726 vdd.n2582 vdd.n922 185
R1727 vdd.n2442 vdd.n2441 185
R1728 vdd.n2444 vdd.n2443 185
R1729 vdd.n2446 vdd.n2445 185
R1730 vdd.n2448 vdd.n2447 185
R1731 vdd.n2450 vdd.n2449 185
R1732 vdd.n2452 vdd.n2451 185
R1733 vdd.n2454 vdd.n2453 185
R1734 vdd.n2456 vdd.n2455 185
R1735 vdd.n2458 vdd.n2457 185
R1736 vdd.n2460 vdd.n2459 185
R1737 vdd.n2462 vdd.n2461 185
R1738 vdd.n2464 vdd.n2463 185
R1739 vdd.n2466 vdd.n2465 185
R1740 vdd.n2468 vdd.n2467 185
R1741 vdd.n2470 vdd.n2469 185
R1742 vdd.n2472 vdd.n2471 185
R1743 vdd.n2474 vdd.n2473 185
R1744 vdd.n2476 vdd.n2475 185
R1745 vdd.n2478 vdd.n2477 185
R1746 vdd.n2480 vdd.n2479 185
R1747 vdd.n2482 vdd.n2481 185
R1748 vdd.n2484 vdd.n2483 185
R1749 vdd.n2486 vdd.n2485 185
R1750 vdd.n2488 vdd.n2487 185
R1751 vdd.n2490 vdd.n2489 185
R1752 vdd.n2492 vdd.n2491 185
R1753 vdd.n2494 vdd.n2493 185
R1754 vdd.n2496 vdd.n2495 185
R1755 vdd.n2498 vdd.n2497 185
R1756 vdd.n2500 vdd.n2499 185
R1757 vdd.n2502 vdd.n2501 185
R1758 vdd.n2504 vdd.n2503 185
R1759 vdd.n2506 vdd.n2505 185
R1760 vdd.n2507 vdd.n950 185
R1761 vdd.n2439 vdd.n948 185
R1762 vdd.n2510 vdd.n948 185
R1763 vdd.n2438 vdd.n2437 185
R1764 vdd.n2437 vdd.n947 185
R1765 vdd.n2436 vdd.n955 185
R1766 vdd.n2436 vdd.n2435 185
R1767 vdd.n1227 vdd.n956 185
R1768 vdd.n1309 vdd.n956 185
R1769 vdd.n1228 vdd.n965 185
R1770 vdd.n2428 vdd.n965 185
R1771 vdd.n1230 vdd.n1229 185
R1772 vdd.n1229 vdd.n963 185
R1773 vdd.n1231 vdd.n972 185
R1774 vdd.n2420 vdd.n972 185
R1775 vdd.n1233 vdd.n1232 185
R1776 vdd.n1232 vdd.n970 185
R1777 vdd.n1234 vdd.n978 185
R1778 vdd.n2414 vdd.n978 185
R1779 vdd.n1236 vdd.n1235 185
R1780 vdd.n1235 vdd.n976 185
R1781 vdd.n1237 vdd.n983 185
R1782 vdd.n2408 vdd.n983 185
R1783 vdd.n1239 vdd.n1238 185
R1784 vdd.n1238 vdd.n989 185
R1785 vdd.n1240 vdd.n988 185
R1786 vdd.n2402 vdd.n988 185
R1787 vdd.n1242 vdd.n1241 185
R1788 vdd.n1241 vdd.n995 185
R1789 vdd.n1243 vdd.n994 185
R1790 vdd.n2396 vdd.n994 185
R1791 vdd.n1332 vdd.n1331 185
R1792 vdd.n1331 vdd.n1330 185
R1793 vdd.n1333 vdd.n1001 185
R1794 vdd.n2390 vdd.n1001 185
R1795 vdd.n1335 vdd.n1334 185
R1796 vdd.n1334 vdd.n999 185
R1797 vdd.n1336 vdd.n1007 185
R1798 vdd.n2384 vdd.n1007 185
R1799 vdd.n1338 vdd.n1337 185
R1800 vdd.n1337 vdd.n1005 185
R1801 vdd.n1339 vdd.n1012 185
R1802 vdd.n2378 vdd.n1012 185
R1803 vdd.n1341 vdd.n1340 185
R1804 vdd.n1340 vdd.n1019 185
R1805 vdd.n1342 vdd.n1018 185
R1806 vdd.n2371 vdd.n1018 185
R1807 vdd.n1344 vdd.n1343 185
R1808 vdd.n1343 vdd.n1026 185
R1809 vdd.n1345 vdd.n1025 185
R1810 vdd.n2365 vdd.n1025 185
R1811 vdd.n1347 vdd.n1346 185
R1812 vdd.n1346 vdd.n1023 185
R1813 vdd.n1348 vdd.n1032 185
R1814 vdd.n2359 vdd.n1032 185
R1815 vdd.n1350 vdd.n1349 185
R1816 vdd.n1349 vdd.n1030 185
R1817 vdd.n1351 vdd.n1038 185
R1818 vdd.n2353 vdd.n1038 185
R1819 vdd.n1353 vdd.n1352 185
R1820 vdd.n1352 vdd.n1036 185
R1821 vdd.n1354 vdd.n1043 185
R1822 vdd.n2347 vdd.n1043 185
R1823 vdd.n1356 vdd.n1355 185
R1824 vdd.n1355 vdd.n1050 185
R1825 vdd.n1357 vdd.n1049 185
R1826 vdd.n2341 vdd.n1049 185
R1827 vdd.n1359 vdd.n1358 185
R1828 vdd.n1358 vdd.n1047 185
R1829 vdd.n2337 vdd.n2336 185
R1830 vdd.n1053 vdd.n1052 185
R1831 vdd.n1194 vdd.n1193 185
R1832 vdd.n1196 vdd.n1195 185
R1833 vdd.n1198 vdd.n1197 185
R1834 vdd.n1200 vdd.n1199 185
R1835 vdd.n1202 vdd.n1201 185
R1836 vdd.n1204 vdd.n1203 185
R1837 vdd.n1206 vdd.n1205 185
R1838 vdd.n1208 vdd.n1207 185
R1839 vdd.n1210 vdd.n1209 185
R1840 vdd.n1212 vdd.n1211 185
R1841 vdd.n1214 vdd.n1213 185
R1842 vdd.n1216 vdd.n1215 185
R1843 vdd.n1218 vdd.n1217 185
R1844 vdd.n1220 vdd.n1219 185
R1845 vdd.n1222 vdd.n1221 185
R1846 vdd.n1393 vdd.n1223 185
R1847 vdd.n1392 vdd.n1391 185
R1848 vdd.n1390 vdd.n1389 185
R1849 vdd.n1388 vdd.n1387 185
R1850 vdd.n1386 vdd.n1385 185
R1851 vdd.n1384 vdd.n1383 185
R1852 vdd.n1382 vdd.n1381 185
R1853 vdd.n1380 vdd.n1379 185
R1854 vdd.n1378 vdd.n1377 185
R1855 vdd.n1376 vdd.n1375 185
R1856 vdd.n1374 vdd.n1373 185
R1857 vdd.n1372 vdd.n1371 185
R1858 vdd.n1370 vdd.n1369 185
R1859 vdd.n1368 vdd.n1367 185
R1860 vdd.n1366 vdd.n1365 185
R1861 vdd.n1364 vdd.n1363 185
R1862 vdd.n1362 vdd.n1361 185
R1863 vdd.n1360 vdd.n1087 185
R1864 vdd.n2334 vdd.n1087 185
R1865 vdd.n2334 vdd.n1054 179.345
R1866 vdd.n756 vdd.n658 179.345
R1867 vdd.n315 vdd.n314 171.744
R1868 vdd.n314 vdd.n313 171.744
R1869 vdd.n313 vdd.n282 171.744
R1870 vdd.n306 vdd.n282 171.744
R1871 vdd.n306 vdd.n305 171.744
R1872 vdd.n305 vdd.n287 171.744
R1873 vdd.n298 vdd.n287 171.744
R1874 vdd.n298 vdd.n297 171.744
R1875 vdd.n297 vdd.n291 171.744
R1876 vdd.n260 vdd.n259 171.744
R1877 vdd.n259 vdd.n258 171.744
R1878 vdd.n258 vdd.n227 171.744
R1879 vdd.n251 vdd.n227 171.744
R1880 vdd.n251 vdd.n250 171.744
R1881 vdd.n250 vdd.n232 171.744
R1882 vdd.n243 vdd.n232 171.744
R1883 vdd.n243 vdd.n242 171.744
R1884 vdd.n242 vdd.n236 171.744
R1885 vdd.n217 vdd.n216 171.744
R1886 vdd.n216 vdd.n215 171.744
R1887 vdd.n215 vdd.n184 171.744
R1888 vdd.n208 vdd.n184 171.744
R1889 vdd.n208 vdd.n207 171.744
R1890 vdd.n207 vdd.n189 171.744
R1891 vdd.n200 vdd.n189 171.744
R1892 vdd.n200 vdd.n199 171.744
R1893 vdd.n199 vdd.n193 171.744
R1894 vdd.n162 vdd.n161 171.744
R1895 vdd.n161 vdd.n160 171.744
R1896 vdd.n160 vdd.n129 171.744
R1897 vdd.n153 vdd.n129 171.744
R1898 vdd.n153 vdd.n152 171.744
R1899 vdd.n152 vdd.n134 171.744
R1900 vdd.n145 vdd.n134 171.744
R1901 vdd.n145 vdd.n144 171.744
R1902 vdd.n144 vdd.n138 171.744
R1903 vdd.n120 vdd.n119 171.744
R1904 vdd.n119 vdd.n118 171.744
R1905 vdd.n118 vdd.n87 171.744
R1906 vdd.n111 vdd.n87 171.744
R1907 vdd.n111 vdd.n110 171.744
R1908 vdd.n110 vdd.n92 171.744
R1909 vdd.n103 vdd.n92 171.744
R1910 vdd.n103 vdd.n102 171.744
R1911 vdd.n102 vdd.n96 171.744
R1912 vdd.n65 vdd.n64 171.744
R1913 vdd.n64 vdd.n63 171.744
R1914 vdd.n63 vdd.n32 171.744
R1915 vdd.n56 vdd.n32 171.744
R1916 vdd.n56 vdd.n55 171.744
R1917 vdd.n55 vdd.n37 171.744
R1918 vdd.n48 vdd.n37 171.744
R1919 vdd.n48 vdd.n47 171.744
R1920 vdd.n47 vdd.n41 171.744
R1921 vdd.n2046 vdd.n2045 171.744
R1922 vdd.n2045 vdd.n2044 171.744
R1923 vdd.n2044 vdd.n2013 171.744
R1924 vdd.n2037 vdd.n2013 171.744
R1925 vdd.n2037 vdd.n2036 171.744
R1926 vdd.n2036 vdd.n2018 171.744
R1927 vdd.n2029 vdd.n2018 171.744
R1928 vdd.n2029 vdd.n2028 171.744
R1929 vdd.n2028 vdd.n2022 171.744
R1930 vdd.n2101 vdd.n2100 171.744
R1931 vdd.n2100 vdd.n2099 171.744
R1932 vdd.n2099 vdd.n2068 171.744
R1933 vdd.n2092 vdd.n2068 171.744
R1934 vdd.n2092 vdd.n2091 171.744
R1935 vdd.n2091 vdd.n2073 171.744
R1936 vdd.n2084 vdd.n2073 171.744
R1937 vdd.n2084 vdd.n2083 171.744
R1938 vdd.n2083 vdd.n2077 171.744
R1939 vdd.n1948 vdd.n1947 171.744
R1940 vdd.n1947 vdd.n1946 171.744
R1941 vdd.n1946 vdd.n1915 171.744
R1942 vdd.n1939 vdd.n1915 171.744
R1943 vdd.n1939 vdd.n1938 171.744
R1944 vdd.n1938 vdd.n1920 171.744
R1945 vdd.n1931 vdd.n1920 171.744
R1946 vdd.n1931 vdd.n1930 171.744
R1947 vdd.n1930 vdd.n1924 171.744
R1948 vdd.n2003 vdd.n2002 171.744
R1949 vdd.n2002 vdd.n2001 171.744
R1950 vdd.n2001 vdd.n1970 171.744
R1951 vdd.n1994 vdd.n1970 171.744
R1952 vdd.n1994 vdd.n1993 171.744
R1953 vdd.n1993 vdd.n1975 171.744
R1954 vdd.n1986 vdd.n1975 171.744
R1955 vdd.n1986 vdd.n1985 171.744
R1956 vdd.n1985 vdd.n1979 171.744
R1957 vdd.n1851 vdd.n1850 171.744
R1958 vdd.n1850 vdd.n1849 171.744
R1959 vdd.n1849 vdd.n1818 171.744
R1960 vdd.n1842 vdd.n1818 171.744
R1961 vdd.n1842 vdd.n1841 171.744
R1962 vdd.n1841 vdd.n1823 171.744
R1963 vdd.n1834 vdd.n1823 171.744
R1964 vdd.n1834 vdd.n1833 171.744
R1965 vdd.n1833 vdd.n1827 171.744
R1966 vdd.n1906 vdd.n1905 171.744
R1967 vdd.n1905 vdd.n1904 171.744
R1968 vdd.n1904 vdd.n1873 171.744
R1969 vdd.n1897 vdd.n1873 171.744
R1970 vdd.n1897 vdd.n1896 171.744
R1971 vdd.n1896 vdd.n1878 171.744
R1972 vdd.n1889 vdd.n1878 171.744
R1973 vdd.n1889 vdd.n1888 171.744
R1974 vdd.n1888 vdd.n1882 171.744
R1975 vdd.n449 vdd.n448 146.341
R1976 vdd.n455 vdd.n454 146.341
R1977 vdd.n459 vdd.n458 146.341
R1978 vdd.n465 vdd.n464 146.341
R1979 vdd.n469 vdd.n468 146.341
R1980 vdd.n475 vdd.n474 146.341
R1981 vdd.n479 vdd.n478 146.341
R1982 vdd.n485 vdd.n484 146.341
R1983 vdd.n489 vdd.n488 146.341
R1984 vdd.n495 vdd.n494 146.341
R1985 vdd.n499 vdd.n498 146.341
R1986 vdd.n505 vdd.n504 146.341
R1987 vdd.n509 vdd.n508 146.341
R1988 vdd.n515 vdd.n514 146.341
R1989 vdd.n519 vdd.n518 146.341
R1990 vdd.n525 vdd.n524 146.341
R1991 vdd.n529 vdd.n528 146.341
R1992 vdd.n535 vdd.n534 146.341
R1993 vdd.n539 vdd.n538 146.341
R1994 vdd.n545 vdd.n544 146.341
R1995 vdd.n549 vdd.n548 146.341
R1996 vdd.n555 vdd.n554 146.341
R1997 vdd.n559 vdd.n558 146.341
R1998 vdd.n565 vdd.n564 146.341
R1999 vdd.n569 vdd.n568 146.341
R2000 vdd.n575 vdd.n574 146.341
R2001 vdd.n579 vdd.n578 146.341
R2002 vdd.n585 vdd.n584 146.341
R2003 vdd.n589 vdd.n588 146.341
R2004 vdd.n595 vdd.n594 146.341
R2005 vdd.n597 vdd.n404 146.341
R2006 vdd.n3238 vdd.n654 146.341
R2007 vdd.n3244 vdd.n654 146.341
R2008 vdd.n3244 vdd.n647 146.341
R2009 vdd.n3254 vdd.n647 146.341
R2010 vdd.n3254 vdd.n643 146.341
R2011 vdd.n3260 vdd.n643 146.341
R2012 vdd.n3260 vdd.n634 146.341
R2013 vdd.n3270 vdd.n634 146.341
R2014 vdd.n3270 vdd.n630 146.341
R2015 vdd.n3276 vdd.n630 146.341
R2016 vdd.n3276 vdd.n623 146.341
R2017 vdd.n3287 vdd.n623 146.341
R2018 vdd.n3287 vdd.n619 146.341
R2019 vdd.n3296 vdd.n619 146.341
R2020 vdd.n3296 vdd.n612 146.341
R2021 vdd.n3306 vdd.n612 146.341
R2022 vdd.n3307 vdd.n3306 146.341
R2023 vdd.n3307 vdd.n329 146.341
R2024 vdd.n330 vdd.n329 146.341
R2025 vdd.n331 vdd.n330 146.341
R2026 vdd.n3314 vdd.n331 146.341
R2027 vdd.n3314 vdd.n339 146.341
R2028 vdd.n340 vdd.n339 146.341
R2029 vdd.n341 vdd.n340 146.341
R2030 vdd.n3321 vdd.n341 146.341
R2031 vdd.n3321 vdd.n350 146.341
R2032 vdd.n351 vdd.n350 146.341
R2033 vdd.n352 vdd.n351 146.341
R2034 vdd.n3329 vdd.n352 146.341
R2035 vdd.n3329 vdd.n360 146.341
R2036 vdd.n361 vdd.n360 146.341
R2037 vdd.n362 vdd.n361 146.341
R2038 vdd.n3336 vdd.n362 146.341
R2039 vdd.n3336 vdd.n371 146.341
R2040 vdd.n372 vdd.n371 146.341
R2041 vdd.n3230 vdd.n3228 146.341
R2042 vdd.n3228 vdd.n3227 146.341
R2043 vdd.n3224 vdd.n3223 146.341
R2044 vdd.n3220 vdd.n3219 146.341
R2045 vdd.n3217 vdd.n669 146.341
R2046 vdd.n3213 vdd.n3211 146.341
R2047 vdd.n3209 vdd.n675 146.341
R2048 vdd.n3205 vdd.n3203 146.341
R2049 vdd.n3201 vdd.n681 146.341
R2050 vdd.n3197 vdd.n3195 146.341
R2051 vdd.n3193 vdd.n689 146.341
R2052 vdd.n3189 vdd.n3187 146.341
R2053 vdd.n3185 vdd.n695 146.341
R2054 vdd.n3181 vdd.n3179 146.341
R2055 vdd.n3177 vdd.n701 146.341
R2056 vdd.n3173 vdd.n3171 146.341
R2057 vdd.n3169 vdd.n707 146.341
R2058 vdd.n3165 vdd.n3163 146.341
R2059 vdd.n3161 vdd.n713 146.341
R2060 vdd.n3157 vdd.n3155 146.341
R2061 vdd.n3153 vdd.n719 146.341
R2062 vdd.n3146 vdd.n728 146.341
R2063 vdd.n3144 vdd.n3143 146.341
R2064 vdd.n3140 vdd.n3139 146.341
R2065 vdd.n3137 vdd.n733 146.341
R2066 vdd.n3133 vdd.n3131 146.341
R2067 vdd.n3129 vdd.n739 146.341
R2068 vdd.n3125 vdd.n3123 146.341
R2069 vdd.n3121 vdd.n745 146.341
R2070 vdd.n3117 vdd.n3115 146.341
R2071 vdd.n3112 vdd.n3111 146.341
R2072 vdd.n3108 vdd.n657 146.341
R2073 vdd.n3236 vdd.n653 146.341
R2074 vdd.n3246 vdd.n653 146.341
R2075 vdd.n3246 vdd.n649 146.341
R2076 vdd.n3252 vdd.n649 146.341
R2077 vdd.n3252 vdd.n641 146.341
R2078 vdd.n3262 vdd.n641 146.341
R2079 vdd.n3262 vdd.n637 146.341
R2080 vdd.n3268 vdd.n637 146.341
R2081 vdd.n3268 vdd.n629 146.341
R2082 vdd.n3279 vdd.n629 146.341
R2083 vdd.n3279 vdd.n625 146.341
R2084 vdd.n3285 vdd.n625 146.341
R2085 vdd.n3285 vdd.n618 146.341
R2086 vdd.n3298 vdd.n618 146.341
R2087 vdd.n3298 vdd.n614 146.341
R2088 vdd.n3304 vdd.n614 146.341
R2089 vdd.n3304 vdd.n326 146.341
R2090 vdd.n3380 vdd.n326 146.341
R2091 vdd.n3380 vdd.n327 146.341
R2092 vdd.n3376 vdd.n327 146.341
R2093 vdd.n3376 vdd.n333 146.341
R2094 vdd.n3372 vdd.n333 146.341
R2095 vdd.n3372 vdd.n338 146.341
R2096 vdd.n3368 vdd.n338 146.341
R2097 vdd.n3368 vdd.n342 146.341
R2098 vdd.n3364 vdd.n342 146.341
R2099 vdd.n3364 vdd.n348 146.341
R2100 vdd.n3360 vdd.n348 146.341
R2101 vdd.n3360 vdd.n353 146.341
R2102 vdd.n3356 vdd.n353 146.341
R2103 vdd.n3356 vdd.n359 146.341
R2104 vdd.n3352 vdd.n359 146.341
R2105 vdd.n3352 vdd.n364 146.341
R2106 vdd.n3348 vdd.n364 146.341
R2107 vdd.n3348 vdd.n370 146.341
R2108 vdd.n2295 vdd.n2294 146.341
R2109 vdd.n2292 vdd.n2289 146.341
R2110 vdd.n2287 vdd.n1098 146.341
R2111 vdd.n2283 vdd.n2282 146.341
R2112 vdd.n2280 vdd.n1102 146.341
R2113 vdd.n2276 vdd.n2275 146.341
R2114 vdd.n2273 vdd.n1109 146.341
R2115 vdd.n2269 vdd.n2268 146.341
R2116 vdd.n2266 vdd.n1116 146.341
R2117 vdd.n1127 vdd.n1124 146.341
R2118 vdd.n2258 vdd.n2257 146.341
R2119 vdd.n2255 vdd.n1129 146.341
R2120 vdd.n2251 vdd.n2250 146.341
R2121 vdd.n2248 vdd.n1135 146.341
R2122 vdd.n2244 vdd.n2243 146.341
R2123 vdd.n2241 vdd.n1142 146.341
R2124 vdd.n2237 vdd.n2236 146.341
R2125 vdd.n2234 vdd.n1149 146.341
R2126 vdd.n2230 vdd.n2229 146.341
R2127 vdd.n2227 vdd.n1156 146.341
R2128 vdd.n1167 vdd.n1164 146.341
R2129 vdd.n2219 vdd.n2218 146.341
R2130 vdd.n2216 vdd.n1169 146.341
R2131 vdd.n2212 vdd.n2211 146.341
R2132 vdd.n2209 vdd.n1175 146.341
R2133 vdd.n2205 vdd.n2204 146.341
R2134 vdd.n2202 vdd.n1182 146.341
R2135 vdd.n2198 vdd.n2197 146.341
R2136 vdd.n2195 vdd.n1189 146.341
R2137 vdd.n1400 vdd.n1398 146.341
R2138 vdd.n1403 vdd.n1402 146.341
R2139 vdd.n1743 vdd.n1507 146.341
R2140 vdd.n1743 vdd.n1499 146.341
R2141 vdd.n1753 vdd.n1499 146.341
R2142 vdd.n1753 vdd.n1495 146.341
R2143 vdd.n1759 vdd.n1495 146.341
R2144 vdd.n1759 vdd.n1487 146.341
R2145 vdd.n1770 vdd.n1487 146.341
R2146 vdd.n1770 vdd.n1483 146.341
R2147 vdd.n1776 vdd.n1483 146.341
R2148 vdd.n1776 vdd.n1477 146.341
R2149 vdd.n1787 vdd.n1477 146.341
R2150 vdd.n1787 vdd.n1473 146.341
R2151 vdd.n1793 vdd.n1473 146.341
R2152 vdd.n1793 vdd.n1464 146.341
R2153 vdd.n1803 vdd.n1464 146.341
R2154 vdd.n1803 vdd.n1460 146.341
R2155 vdd.n1809 vdd.n1460 146.341
R2156 vdd.n1809 vdd.n1453 146.341
R2157 vdd.n2115 vdd.n1453 146.341
R2158 vdd.n2115 vdd.n1449 146.341
R2159 vdd.n2121 vdd.n1449 146.341
R2160 vdd.n2121 vdd.n1442 146.341
R2161 vdd.n2131 vdd.n1442 146.341
R2162 vdd.n2131 vdd.n1438 146.341
R2163 vdd.n2137 vdd.n1438 146.341
R2164 vdd.n2137 vdd.n1430 146.341
R2165 vdd.n2148 vdd.n1430 146.341
R2166 vdd.n2148 vdd.n1426 146.341
R2167 vdd.n2154 vdd.n1426 146.341
R2168 vdd.n2154 vdd.n1420 146.341
R2169 vdd.n2165 vdd.n1420 146.341
R2170 vdd.n2165 vdd.n1415 146.341
R2171 vdd.n2173 vdd.n1415 146.341
R2172 vdd.n2173 vdd.n1405 146.341
R2173 vdd.n2183 vdd.n1405 146.341
R2174 vdd.n1545 vdd.n1544 146.341
R2175 vdd.n1549 vdd.n1544 146.341
R2176 vdd.n1551 vdd.n1550 146.341
R2177 vdd.n1555 vdd.n1554 146.341
R2178 vdd.n1557 vdd.n1556 146.341
R2179 vdd.n1561 vdd.n1560 146.341
R2180 vdd.n1563 vdd.n1562 146.341
R2181 vdd.n1567 vdd.n1566 146.341
R2182 vdd.n1569 vdd.n1568 146.341
R2183 vdd.n1701 vdd.n1700 146.341
R2184 vdd.n1573 vdd.n1572 146.341
R2185 vdd.n1577 vdd.n1576 146.341
R2186 vdd.n1579 vdd.n1578 146.341
R2187 vdd.n1583 vdd.n1582 146.341
R2188 vdd.n1585 vdd.n1584 146.341
R2189 vdd.n1589 vdd.n1588 146.341
R2190 vdd.n1591 vdd.n1590 146.341
R2191 vdd.n1595 vdd.n1594 146.341
R2192 vdd.n1597 vdd.n1596 146.341
R2193 vdd.n1601 vdd.n1600 146.341
R2194 vdd.n1665 vdd.n1602 146.341
R2195 vdd.n1606 vdd.n1605 146.341
R2196 vdd.n1608 vdd.n1607 146.341
R2197 vdd.n1612 vdd.n1611 146.341
R2198 vdd.n1614 vdd.n1613 146.341
R2199 vdd.n1618 vdd.n1617 146.341
R2200 vdd.n1620 vdd.n1619 146.341
R2201 vdd.n1624 vdd.n1623 146.341
R2202 vdd.n1626 vdd.n1625 146.341
R2203 vdd.n1630 vdd.n1629 146.341
R2204 vdd.n1632 vdd.n1631 146.341
R2205 vdd.n1737 vdd.n1513 146.341
R2206 vdd.n1745 vdd.n1505 146.341
R2207 vdd.n1745 vdd.n1501 146.341
R2208 vdd.n1751 vdd.n1501 146.341
R2209 vdd.n1751 vdd.n1493 146.341
R2210 vdd.n1762 vdd.n1493 146.341
R2211 vdd.n1762 vdd.n1489 146.341
R2212 vdd.n1768 vdd.n1489 146.341
R2213 vdd.n1768 vdd.n1482 146.341
R2214 vdd.n1779 vdd.n1482 146.341
R2215 vdd.n1779 vdd.n1478 146.341
R2216 vdd.n1785 vdd.n1478 146.341
R2217 vdd.n1785 vdd.n1471 146.341
R2218 vdd.n1795 vdd.n1471 146.341
R2219 vdd.n1795 vdd.n1467 146.341
R2220 vdd.n1801 vdd.n1467 146.341
R2221 vdd.n1801 vdd.n1459 146.341
R2222 vdd.n1812 vdd.n1459 146.341
R2223 vdd.n1812 vdd.n1455 146.341
R2224 vdd.n2113 vdd.n1455 146.341
R2225 vdd.n2113 vdd.n1448 146.341
R2226 vdd.n2123 vdd.n1448 146.341
R2227 vdd.n2123 vdd.n1444 146.341
R2228 vdd.n2129 vdd.n1444 146.341
R2229 vdd.n2129 vdd.n1436 146.341
R2230 vdd.n2140 vdd.n1436 146.341
R2231 vdd.n2140 vdd.n1432 146.341
R2232 vdd.n2146 vdd.n1432 146.341
R2233 vdd.n2146 vdd.n1425 146.341
R2234 vdd.n2157 vdd.n1425 146.341
R2235 vdd.n2157 vdd.n1421 146.341
R2236 vdd.n2163 vdd.n1421 146.341
R2237 vdd.n2163 vdd.n1413 146.341
R2238 vdd.n2175 vdd.n1413 146.341
R2239 vdd.n2175 vdd.n1408 146.341
R2240 vdd.n2181 vdd.n1408 146.341
R2241 vdd.n1224 vdd.t24 127.284
R2242 vdd.n952 vdd.t65 127.284
R2243 vdd.n1244 vdd.t38 127.284
R2244 vdd.n943 vdd.t82 127.284
R2245 vdd.n843 vdd.t41 127.284
R2246 vdd.n843 vdd.t42 127.284
R2247 vdd.n2621 vdd.t77 127.284
R2248 vdd.n804 vdd.t88 127.284
R2249 vdd.n2618 vdd.t70 127.284
R2250 vdd.n768 vdd.t19 127.284
R2251 vdd.n1014 vdd.t73 127.284
R2252 vdd.n1014 vdd.t74 127.284
R2253 vdd.n22 vdd.n20 117.314
R2254 vdd.n17 vdd.n15 117.314
R2255 vdd.n27 vdd.n26 116.927
R2256 vdd.n24 vdd.n23 116.927
R2257 vdd.n22 vdd.n21 116.927
R2258 vdd.n17 vdd.n16 116.927
R2259 vdd.n19 vdd.n18 116.927
R2260 vdd.n27 vdd.n25 116.927
R2261 vdd.n1225 vdd.t23 111.188
R2262 vdd.n953 vdd.t66 111.188
R2263 vdd.n1245 vdd.t37 111.188
R2264 vdd.n944 vdd.t83 111.188
R2265 vdd.n2622 vdd.t76 111.188
R2266 vdd.n805 vdd.t89 111.188
R2267 vdd.n2619 vdd.t69 111.188
R2268 vdd.n769 vdd.t20 111.188
R2269 vdd.n2863 vdd.n898 99.5127
R2270 vdd.n2863 vdd.n896 99.5127
R2271 vdd.n2867 vdd.n896 99.5127
R2272 vdd.n2867 vdd.n887 99.5127
R2273 vdd.n2875 vdd.n887 99.5127
R2274 vdd.n2875 vdd.n885 99.5127
R2275 vdd.n2879 vdd.n885 99.5127
R2276 vdd.n2879 vdd.n875 99.5127
R2277 vdd.n2887 vdd.n875 99.5127
R2278 vdd.n2887 vdd.n873 99.5127
R2279 vdd.n2891 vdd.n873 99.5127
R2280 vdd.n2891 vdd.n863 99.5127
R2281 vdd.n2899 vdd.n863 99.5127
R2282 vdd.n2899 vdd.n861 99.5127
R2283 vdd.n2903 vdd.n861 99.5127
R2284 vdd.n2903 vdd.n852 99.5127
R2285 vdd.n2911 vdd.n852 99.5127
R2286 vdd.n2911 vdd.n850 99.5127
R2287 vdd.n2915 vdd.n850 99.5127
R2288 vdd.n2915 vdd.n838 99.5127
R2289 vdd.n2924 vdd.n838 99.5127
R2290 vdd.n2924 vdd.n836 99.5127
R2291 vdd.n2928 vdd.n836 99.5127
R2292 vdd.n2928 vdd.n827 99.5127
R2293 vdd.n2936 vdd.n827 99.5127
R2294 vdd.n2936 vdd.n825 99.5127
R2295 vdd.n2940 vdd.n825 99.5127
R2296 vdd.n2940 vdd.n813 99.5127
R2297 vdd.n2993 vdd.n813 99.5127
R2298 vdd.n2993 vdd.n811 99.5127
R2299 vdd.n2997 vdd.n811 99.5127
R2300 vdd.n2997 vdd.n777 99.5127
R2301 vdd.n3067 vdd.n777 99.5127
R2302 vdd.n3063 vdd.n778 99.5127
R2303 vdd.n3061 vdd.n3060 99.5127
R2304 vdd.n3058 vdd.n782 99.5127
R2305 vdd.n3054 vdd.n3053 99.5127
R2306 vdd.n3051 vdd.n785 99.5127
R2307 vdd.n3047 vdd.n3046 99.5127
R2308 vdd.n3044 vdd.n788 99.5127
R2309 vdd.n3040 vdd.n3039 99.5127
R2310 vdd.n3037 vdd.n791 99.5127
R2311 vdd.n3032 vdd.n3031 99.5127
R2312 vdd.n3029 vdd.n794 99.5127
R2313 vdd.n3025 vdd.n3024 99.5127
R2314 vdd.n3022 vdd.n797 99.5127
R2315 vdd.n3018 vdd.n3017 99.5127
R2316 vdd.n3015 vdd.n800 99.5127
R2317 vdd.n3011 vdd.n3010 99.5127
R2318 vdd.n3008 vdd.n803 99.5127
R2319 vdd.n2784 vdd.n900 99.5127
R2320 vdd.n2780 vdd.n900 99.5127
R2321 vdd.n2780 vdd.n894 99.5127
R2322 vdd.n2724 vdd.n894 99.5127
R2323 vdd.n2724 vdd.n889 99.5127
R2324 vdd.n2727 vdd.n889 99.5127
R2325 vdd.n2727 vdd.n883 99.5127
R2326 vdd.n2730 vdd.n883 99.5127
R2327 vdd.n2730 vdd.n877 99.5127
R2328 vdd.n2763 vdd.n877 99.5127
R2329 vdd.n2763 vdd.n870 99.5127
R2330 vdd.n2759 vdd.n870 99.5127
R2331 vdd.n2759 vdd.n864 99.5127
R2332 vdd.n2756 vdd.n864 99.5127
R2333 vdd.n2756 vdd.n859 99.5127
R2334 vdd.n2753 vdd.n859 99.5127
R2335 vdd.n2753 vdd.n854 99.5127
R2336 vdd.n2750 vdd.n854 99.5127
R2337 vdd.n2750 vdd.n847 99.5127
R2338 vdd.n2747 vdd.n847 99.5127
R2339 vdd.n2747 vdd.n839 99.5127
R2340 vdd.n2744 vdd.n839 99.5127
R2341 vdd.n2744 vdd.n834 99.5127
R2342 vdd.n2741 vdd.n834 99.5127
R2343 vdd.n2741 vdd.n829 99.5127
R2344 vdd.n2738 vdd.n829 99.5127
R2345 vdd.n2738 vdd.n823 99.5127
R2346 vdd.n2735 vdd.n823 99.5127
R2347 vdd.n2735 vdd.n815 99.5127
R2348 vdd.n815 vdd.n808 99.5127
R2349 vdd.n2999 vdd.n808 99.5127
R2350 vdd.n3000 vdd.n2999 99.5127
R2351 vdd.n3000 vdd.n775 99.5127
R2352 vdd.n2617 vdd.n2616 99.5127
R2353 vdd.n2848 vdd.n2616 99.5127
R2354 vdd.n2846 vdd.n2845 99.5127
R2355 vdd.n2842 vdd.n2841 99.5127
R2356 vdd.n2838 vdd.n2837 99.5127
R2357 vdd.n2834 vdd.n2833 99.5127
R2358 vdd.n2830 vdd.n2829 99.5127
R2359 vdd.n2826 vdd.n2825 99.5127
R2360 vdd.n2822 vdd.n2821 99.5127
R2361 vdd.n2818 vdd.n2817 99.5127
R2362 vdd.n2814 vdd.n2813 99.5127
R2363 vdd.n2810 vdd.n2809 99.5127
R2364 vdd.n2806 vdd.n2805 99.5127
R2365 vdd.n2802 vdd.n2801 99.5127
R2366 vdd.n2798 vdd.n2797 99.5127
R2367 vdd.n2794 vdd.n2793 99.5127
R2368 vdd.n2789 vdd.n2788 99.5127
R2369 vdd.n2581 vdd.n941 99.5127
R2370 vdd.n2577 vdd.n2576 99.5127
R2371 vdd.n2573 vdd.n2572 99.5127
R2372 vdd.n2569 vdd.n2568 99.5127
R2373 vdd.n2565 vdd.n2564 99.5127
R2374 vdd.n2561 vdd.n2560 99.5127
R2375 vdd.n2557 vdd.n2556 99.5127
R2376 vdd.n2553 vdd.n2552 99.5127
R2377 vdd.n2549 vdd.n2548 99.5127
R2378 vdd.n2545 vdd.n2544 99.5127
R2379 vdd.n2541 vdd.n2540 99.5127
R2380 vdd.n2537 vdd.n2536 99.5127
R2381 vdd.n2533 vdd.n2532 99.5127
R2382 vdd.n2529 vdd.n2528 99.5127
R2383 vdd.n2525 vdd.n2524 99.5127
R2384 vdd.n2521 vdd.n2520 99.5127
R2385 vdd.n2516 vdd.n2515 99.5127
R2386 vdd.n1280 vdd.n1048 99.5127
R2387 vdd.n1283 vdd.n1048 99.5127
R2388 vdd.n1283 vdd.n1042 99.5127
R2389 vdd.n1286 vdd.n1042 99.5127
R2390 vdd.n1286 vdd.n1037 99.5127
R2391 vdd.n1289 vdd.n1037 99.5127
R2392 vdd.n1289 vdd.n1031 99.5127
R2393 vdd.n1292 vdd.n1031 99.5127
R2394 vdd.n1292 vdd.n1024 99.5127
R2395 vdd.n1295 vdd.n1024 99.5127
R2396 vdd.n1295 vdd.n1017 99.5127
R2397 vdd.n1298 vdd.n1017 99.5127
R2398 vdd.n1298 vdd.n1011 99.5127
R2399 vdd.n1301 vdd.n1011 99.5127
R2400 vdd.n1301 vdd.n1006 99.5127
R2401 vdd.n1304 vdd.n1006 99.5127
R2402 vdd.n1304 vdd.n1000 99.5127
R2403 vdd.n1329 vdd.n1000 99.5127
R2404 vdd.n1329 vdd.n993 99.5127
R2405 vdd.n1325 vdd.n993 99.5127
R2406 vdd.n1325 vdd.n987 99.5127
R2407 vdd.n1322 vdd.n987 99.5127
R2408 vdd.n1322 vdd.n982 99.5127
R2409 vdd.n1319 vdd.n982 99.5127
R2410 vdd.n1319 vdd.n977 99.5127
R2411 vdd.n1316 vdd.n977 99.5127
R2412 vdd.n1316 vdd.n971 99.5127
R2413 vdd.n1313 vdd.n971 99.5127
R2414 vdd.n1313 vdd.n964 99.5127
R2415 vdd.n1310 vdd.n964 99.5127
R2416 vdd.n1310 vdd.n957 99.5127
R2417 vdd.n957 vdd.n946 99.5127
R2418 vdd.n2511 vdd.n946 99.5127
R2419 vdd.n1089 vdd.n1088 99.5127
R2420 vdd.n2327 vdd.n1088 99.5127
R2421 vdd.n2325 vdd.n2324 99.5127
R2422 vdd.n2321 vdd.n2320 99.5127
R2423 vdd.n2317 vdd.n2316 99.5127
R2424 vdd.n2313 vdd.n2312 99.5127
R2425 vdd.n2309 vdd.n2308 99.5127
R2426 vdd.n2305 vdd.n2304 99.5127
R2427 vdd.n2301 vdd.n2300 99.5127
R2428 vdd.n1247 vdd.n1246 99.5127
R2429 vdd.n1251 vdd.n1250 99.5127
R2430 vdd.n1255 vdd.n1254 99.5127
R2431 vdd.n1259 vdd.n1258 99.5127
R2432 vdd.n1263 vdd.n1262 99.5127
R2433 vdd.n1267 vdd.n1266 99.5127
R2434 vdd.n1271 vdd.n1270 99.5127
R2435 vdd.n1276 vdd.n1275 99.5127
R2436 vdd.n2342 vdd.n1046 99.5127
R2437 vdd.n2342 vdd.n1044 99.5127
R2438 vdd.n2346 vdd.n1044 99.5127
R2439 vdd.n2346 vdd.n1035 99.5127
R2440 vdd.n2354 vdd.n1035 99.5127
R2441 vdd.n2354 vdd.n1033 99.5127
R2442 vdd.n2358 vdd.n1033 99.5127
R2443 vdd.n2358 vdd.n1022 99.5127
R2444 vdd.n2366 vdd.n1022 99.5127
R2445 vdd.n2366 vdd.n1020 99.5127
R2446 vdd.n2370 vdd.n1020 99.5127
R2447 vdd.n2370 vdd.n1010 99.5127
R2448 vdd.n2379 vdd.n1010 99.5127
R2449 vdd.n2379 vdd.n1008 99.5127
R2450 vdd.n2383 vdd.n1008 99.5127
R2451 vdd.n2383 vdd.n998 99.5127
R2452 vdd.n2391 vdd.n998 99.5127
R2453 vdd.n2391 vdd.n996 99.5127
R2454 vdd.n2395 vdd.n996 99.5127
R2455 vdd.n2395 vdd.n986 99.5127
R2456 vdd.n2403 vdd.n986 99.5127
R2457 vdd.n2403 vdd.n984 99.5127
R2458 vdd.n2407 vdd.n984 99.5127
R2459 vdd.n2407 vdd.n975 99.5127
R2460 vdd.n2415 vdd.n975 99.5127
R2461 vdd.n2415 vdd.n973 99.5127
R2462 vdd.n2419 vdd.n973 99.5127
R2463 vdd.n2419 vdd.n962 99.5127
R2464 vdd.n2429 vdd.n962 99.5127
R2465 vdd.n2429 vdd.n959 99.5127
R2466 vdd.n2434 vdd.n959 99.5127
R2467 vdd.n2434 vdd.n960 99.5127
R2468 vdd.n960 vdd.n940 99.5127
R2469 vdd.n2983 vdd.n2982 99.5127
R2470 vdd.n2980 vdd.n2946 99.5127
R2471 vdd.n2976 vdd.n2975 99.5127
R2472 vdd.n2973 vdd.n2949 99.5127
R2473 vdd.n2969 vdd.n2968 99.5127
R2474 vdd.n2966 vdd.n2952 99.5127
R2475 vdd.n2962 vdd.n2961 99.5127
R2476 vdd.n2959 vdd.n2956 99.5127
R2477 vdd.n3100 vdd.n755 99.5127
R2478 vdd.n3098 vdd.n3097 99.5127
R2479 vdd.n3095 vdd.n758 99.5127
R2480 vdd.n3091 vdd.n3090 99.5127
R2481 vdd.n3088 vdd.n761 99.5127
R2482 vdd.n3084 vdd.n3083 99.5127
R2483 vdd.n3081 vdd.n764 99.5127
R2484 vdd.n3077 vdd.n3076 99.5127
R2485 vdd.n3074 vdd.n767 99.5127
R2486 vdd.n2689 vdd.n901 99.5127
R2487 vdd.n2778 vdd.n901 99.5127
R2488 vdd.n2778 vdd.n895 99.5127
R2489 vdd.n2774 vdd.n895 99.5127
R2490 vdd.n2774 vdd.n890 99.5127
R2491 vdd.n2771 vdd.n890 99.5127
R2492 vdd.n2771 vdd.n884 99.5127
R2493 vdd.n2768 vdd.n884 99.5127
R2494 vdd.n2768 vdd.n878 99.5127
R2495 vdd.n2765 vdd.n878 99.5127
R2496 vdd.n2765 vdd.n871 99.5127
R2497 vdd.n2721 vdd.n871 99.5127
R2498 vdd.n2721 vdd.n865 99.5127
R2499 vdd.n2718 vdd.n865 99.5127
R2500 vdd.n2718 vdd.n860 99.5127
R2501 vdd.n2715 vdd.n860 99.5127
R2502 vdd.n2715 vdd.n855 99.5127
R2503 vdd.n2712 vdd.n855 99.5127
R2504 vdd.n2712 vdd.n848 99.5127
R2505 vdd.n2709 vdd.n848 99.5127
R2506 vdd.n2709 vdd.n840 99.5127
R2507 vdd.n2706 vdd.n840 99.5127
R2508 vdd.n2706 vdd.n835 99.5127
R2509 vdd.n2703 vdd.n835 99.5127
R2510 vdd.n2703 vdd.n830 99.5127
R2511 vdd.n2700 vdd.n830 99.5127
R2512 vdd.n2700 vdd.n824 99.5127
R2513 vdd.n2697 vdd.n824 99.5127
R2514 vdd.n2697 vdd.n816 99.5127
R2515 vdd.n2694 vdd.n816 99.5127
R2516 vdd.n2694 vdd.n809 99.5127
R2517 vdd.n809 vdd.n773 99.5127
R2518 vdd.n3069 vdd.n773 99.5127
R2519 vdd.n2624 vdd.n904 99.5127
R2520 vdd.n2628 vdd.n2627 99.5127
R2521 vdd.n2632 vdd.n2631 99.5127
R2522 vdd.n2636 vdd.n2635 99.5127
R2523 vdd.n2640 vdd.n2639 99.5127
R2524 vdd.n2644 vdd.n2643 99.5127
R2525 vdd.n2648 vdd.n2647 99.5127
R2526 vdd.n2652 vdd.n2651 99.5127
R2527 vdd.n2656 vdd.n2655 99.5127
R2528 vdd.n2660 vdd.n2659 99.5127
R2529 vdd.n2664 vdd.n2663 99.5127
R2530 vdd.n2668 vdd.n2667 99.5127
R2531 vdd.n2672 vdd.n2671 99.5127
R2532 vdd.n2676 vdd.n2675 99.5127
R2533 vdd.n2680 vdd.n2679 99.5127
R2534 vdd.n2684 vdd.n2683 99.5127
R2535 vdd.n2686 vdd.n2615 99.5127
R2536 vdd.n2861 vdd.n902 99.5127
R2537 vdd.n2861 vdd.n893 99.5127
R2538 vdd.n2869 vdd.n893 99.5127
R2539 vdd.n2869 vdd.n891 99.5127
R2540 vdd.n2873 vdd.n891 99.5127
R2541 vdd.n2873 vdd.n881 99.5127
R2542 vdd.n2881 vdd.n881 99.5127
R2543 vdd.n2881 vdd.n879 99.5127
R2544 vdd.n2885 vdd.n879 99.5127
R2545 vdd.n2885 vdd.n869 99.5127
R2546 vdd.n2893 vdd.n869 99.5127
R2547 vdd.n2893 vdd.n867 99.5127
R2548 vdd.n2897 vdd.n867 99.5127
R2549 vdd.n2897 vdd.n858 99.5127
R2550 vdd.n2905 vdd.n858 99.5127
R2551 vdd.n2905 vdd.n856 99.5127
R2552 vdd.n2909 vdd.n856 99.5127
R2553 vdd.n2909 vdd.n845 99.5127
R2554 vdd.n2917 vdd.n845 99.5127
R2555 vdd.n2917 vdd.n842 99.5127
R2556 vdd.n2922 vdd.n842 99.5127
R2557 vdd.n2922 vdd.n833 99.5127
R2558 vdd.n2930 vdd.n833 99.5127
R2559 vdd.n2930 vdd.n831 99.5127
R2560 vdd.n2934 vdd.n831 99.5127
R2561 vdd.n2934 vdd.n821 99.5127
R2562 vdd.n2942 vdd.n821 99.5127
R2563 vdd.n2942 vdd.n818 99.5127
R2564 vdd.n2991 vdd.n818 99.5127
R2565 vdd.n2991 vdd.n819 99.5127
R2566 vdd.n819 vdd.n810 99.5127
R2567 vdd.n2986 vdd.n810 99.5127
R2568 vdd.n2986 vdd.n776 99.5127
R2569 vdd.n2505 vdd.n2504 99.5127
R2570 vdd.n2501 vdd.n2500 99.5127
R2571 vdd.n2497 vdd.n2496 99.5127
R2572 vdd.n2493 vdd.n2492 99.5127
R2573 vdd.n2489 vdd.n2488 99.5127
R2574 vdd.n2485 vdd.n2484 99.5127
R2575 vdd.n2481 vdd.n2480 99.5127
R2576 vdd.n2477 vdd.n2476 99.5127
R2577 vdd.n2473 vdd.n2472 99.5127
R2578 vdd.n2469 vdd.n2468 99.5127
R2579 vdd.n2465 vdd.n2464 99.5127
R2580 vdd.n2461 vdd.n2460 99.5127
R2581 vdd.n2457 vdd.n2456 99.5127
R2582 vdd.n2453 vdd.n2452 99.5127
R2583 vdd.n2449 vdd.n2448 99.5127
R2584 vdd.n2445 vdd.n2444 99.5127
R2585 vdd.n2441 vdd.n922 99.5127
R2586 vdd.n1358 vdd.n1049 99.5127
R2587 vdd.n1355 vdd.n1049 99.5127
R2588 vdd.n1355 vdd.n1043 99.5127
R2589 vdd.n1352 vdd.n1043 99.5127
R2590 vdd.n1352 vdd.n1038 99.5127
R2591 vdd.n1349 vdd.n1038 99.5127
R2592 vdd.n1349 vdd.n1032 99.5127
R2593 vdd.n1346 vdd.n1032 99.5127
R2594 vdd.n1346 vdd.n1025 99.5127
R2595 vdd.n1343 vdd.n1025 99.5127
R2596 vdd.n1343 vdd.n1018 99.5127
R2597 vdd.n1340 vdd.n1018 99.5127
R2598 vdd.n1340 vdd.n1012 99.5127
R2599 vdd.n1337 vdd.n1012 99.5127
R2600 vdd.n1337 vdd.n1007 99.5127
R2601 vdd.n1334 vdd.n1007 99.5127
R2602 vdd.n1334 vdd.n1001 99.5127
R2603 vdd.n1331 vdd.n1001 99.5127
R2604 vdd.n1331 vdd.n994 99.5127
R2605 vdd.n1241 vdd.n994 99.5127
R2606 vdd.n1241 vdd.n988 99.5127
R2607 vdd.n1238 vdd.n988 99.5127
R2608 vdd.n1238 vdd.n983 99.5127
R2609 vdd.n1235 vdd.n983 99.5127
R2610 vdd.n1235 vdd.n978 99.5127
R2611 vdd.n1232 vdd.n978 99.5127
R2612 vdd.n1232 vdd.n972 99.5127
R2613 vdd.n1229 vdd.n972 99.5127
R2614 vdd.n1229 vdd.n965 99.5127
R2615 vdd.n965 vdd.n956 99.5127
R2616 vdd.n2436 vdd.n956 99.5127
R2617 vdd.n2437 vdd.n2436 99.5127
R2618 vdd.n2437 vdd.n948 99.5127
R2619 vdd.n1193 vdd.n1053 99.5127
R2620 vdd.n1197 vdd.n1196 99.5127
R2621 vdd.n1201 vdd.n1200 99.5127
R2622 vdd.n1205 vdd.n1204 99.5127
R2623 vdd.n1209 vdd.n1208 99.5127
R2624 vdd.n1213 vdd.n1212 99.5127
R2625 vdd.n1217 vdd.n1216 99.5127
R2626 vdd.n1221 vdd.n1220 99.5127
R2627 vdd.n1391 vdd.n1223 99.5127
R2628 vdd.n1389 vdd.n1388 99.5127
R2629 vdd.n1385 vdd.n1384 99.5127
R2630 vdd.n1381 vdd.n1380 99.5127
R2631 vdd.n1377 vdd.n1376 99.5127
R2632 vdd.n1373 vdd.n1372 99.5127
R2633 vdd.n1369 vdd.n1368 99.5127
R2634 vdd.n1365 vdd.n1364 99.5127
R2635 vdd.n1361 vdd.n1087 99.5127
R2636 vdd.n2340 vdd.n1051 99.5127
R2637 vdd.n2340 vdd.n1041 99.5127
R2638 vdd.n2348 vdd.n1041 99.5127
R2639 vdd.n2348 vdd.n1039 99.5127
R2640 vdd.n2352 vdd.n1039 99.5127
R2641 vdd.n2352 vdd.n1029 99.5127
R2642 vdd.n2360 vdd.n1029 99.5127
R2643 vdd.n2360 vdd.n1027 99.5127
R2644 vdd.n2364 vdd.n1027 99.5127
R2645 vdd.n2364 vdd.n1016 99.5127
R2646 vdd.n2372 vdd.n1016 99.5127
R2647 vdd.n2372 vdd.n1013 99.5127
R2648 vdd.n2377 vdd.n1013 99.5127
R2649 vdd.n2377 vdd.n1004 99.5127
R2650 vdd.n2385 vdd.n1004 99.5127
R2651 vdd.n2385 vdd.n1002 99.5127
R2652 vdd.n2389 vdd.n1002 99.5127
R2653 vdd.n2389 vdd.n992 99.5127
R2654 vdd.n2397 vdd.n992 99.5127
R2655 vdd.n2397 vdd.n990 99.5127
R2656 vdd.n2401 vdd.n990 99.5127
R2657 vdd.n2401 vdd.n981 99.5127
R2658 vdd.n2409 vdd.n981 99.5127
R2659 vdd.n2409 vdd.n979 99.5127
R2660 vdd.n2413 vdd.n979 99.5127
R2661 vdd.n2413 vdd.n969 99.5127
R2662 vdd.n2421 vdd.n969 99.5127
R2663 vdd.n2421 vdd.n966 99.5127
R2664 vdd.n2427 vdd.n966 99.5127
R2665 vdd.n2427 vdd.n967 99.5127
R2666 vdd.n967 vdd.n958 99.5127
R2667 vdd.n958 vdd.n949 99.5127
R2668 vdd.n2509 vdd.n949 99.5127
R2669 vdd.n9 vdd.n7 98.9633
R2670 vdd.n2 vdd.n0 98.9633
R2671 vdd.n9 vdd.n8 98.6055
R2672 vdd.n11 vdd.n10 98.6055
R2673 vdd.n13 vdd.n12 98.6055
R2674 vdd.n6 vdd.n5 98.6055
R2675 vdd.n4 vdd.n3 98.6055
R2676 vdd.n2 vdd.n1 98.6055
R2677 vdd.t244 vdd.n291 85.8723
R2678 vdd.t168 vdd.n236 85.8723
R2679 vdd.t191 vdd.n193 85.8723
R2680 vdd.t162 vdd.n138 85.8723
R2681 vdd.t151 vdd.n96 85.8723
R2682 vdd.t187 vdd.n41 85.8723
R2683 vdd.t170 vdd.n2022 85.8723
R2684 vdd.t109 vdd.n2077 85.8723
R2685 vdd.t243 vdd.n1924 85.8723
R2686 vdd.t155 vdd.n1979 85.8723
R2687 vdd.t186 vdd.n1827 85.8723
R2688 vdd.t129 vdd.n1882 85.8723
R2689 vdd.n2920 vdd.n843 78.546
R2690 vdd.n2375 vdd.n1014 78.546
R2691 vdd.n278 vdd.n277 75.1835
R2692 vdd.n276 vdd.n275 75.1835
R2693 vdd.n274 vdd.n273 75.1835
R2694 vdd.n272 vdd.n271 75.1835
R2695 vdd.n270 vdd.n269 75.1835
R2696 vdd.n268 vdd.n267 75.1835
R2697 vdd.n266 vdd.n265 75.1835
R2698 vdd.n180 vdd.n179 75.1835
R2699 vdd.n178 vdd.n177 75.1835
R2700 vdd.n176 vdd.n175 75.1835
R2701 vdd.n174 vdd.n173 75.1835
R2702 vdd.n172 vdd.n171 75.1835
R2703 vdd.n170 vdd.n169 75.1835
R2704 vdd.n168 vdd.n167 75.1835
R2705 vdd.n83 vdd.n82 75.1835
R2706 vdd.n81 vdd.n80 75.1835
R2707 vdd.n79 vdd.n78 75.1835
R2708 vdd.n77 vdd.n76 75.1835
R2709 vdd.n75 vdd.n74 75.1835
R2710 vdd.n73 vdd.n72 75.1835
R2711 vdd.n71 vdd.n70 75.1835
R2712 vdd.n2052 vdd.n2051 75.1835
R2713 vdd.n2054 vdd.n2053 75.1835
R2714 vdd.n2056 vdd.n2055 75.1835
R2715 vdd.n2058 vdd.n2057 75.1835
R2716 vdd.n2060 vdd.n2059 75.1835
R2717 vdd.n2062 vdd.n2061 75.1835
R2718 vdd.n2064 vdd.n2063 75.1835
R2719 vdd.n1954 vdd.n1953 75.1835
R2720 vdd.n1956 vdd.n1955 75.1835
R2721 vdd.n1958 vdd.n1957 75.1835
R2722 vdd.n1960 vdd.n1959 75.1835
R2723 vdd.n1962 vdd.n1961 75.1835
R2724 vdd.n1964 vdd.n1963 75.1835
R2725 vdd.n1966 vdd.n1965 75.1835
R2726 vdd.n1857 vdd.n1856 75.1835
R2727 vdd.n1859 vdd.n1858 75.1835
R2728 vdd.n1861 vdd.n1860 75.1835
R2729 vdd.n1863 vdd.n1862 75.1835
R2730 vdd.n1865 vdd.n1864 75.1835
R2731 vdd.n1867 vdd.n1866 75.1835
R2732 vdd.n1869 vdd.n1868 75.1835
R2733 vdd.n2856 vdd.n2855 72.8958
R2734 vdd.n2855 vdd.n2599 72.8958
R2735 vdd.n2855 vdd.n2600 72.8958
R2736 vdd.n2855 vdd.n2601 72.8958
R2737 vdd.n2855 vdd.n2602 72.8958
R2738 vdd.n2855 vdd.n2603 72.8958
R2739 vdd.n2855 vdd.n2604 72.8958
R2740 vdd.n2855 vdd.n2605 72.8958
R2741 vdd.n2855 vdd.n2606 72.8958
R2742 vdd.n2855 vdd.n2607 72.8958
R2743 vdd.n2855 vdd.n2608 72.8958
R2744 vdd.n2855 vdd.n2609 72.8958
R2745 vdd.n2855 vdd.n2610 72.8958
R2746 vdd.n2855 vdd.n2611 72.8958
R2747 vdd.n2855 vdd.n2612 72.8958
R2748 vdd.n2855 vdd.n2613 72.8958
R2749 vdd.n2855 vdd.n2614 72.8958
R2750 vdd.n772 vdd.n756 72.8958
R2751 vdd.n3075 vdd.n756 72.8958
R2752 vdd.n766 vdd.n756 72.8958
R2753 vdd.n3082 vdd.n756 72.8958
R2754 vdd.n763 vdd.n756 72.8958
R2755 vdd.n3089 vdd.n756 72.8958
R2756 vdd.n760 vdd.n756 72.8958
R2757 vdd.n3096 vdd.n756 72.8958
R2758 vdd.n3099 vdd.n756 72.8958
R2759 vdd.n2955 vdd.n756 72.8958
R2760 vdd.n2960 vdd.n756 72.8958
R2761 vdd.n2954 vdd.n756 72.8958
R2762 vdd.n2967 vdd.n756 72.8958
R2763 vdd.n2951 vdd.n756 72.8958
R2764 vdd.n2974 vdd.n756 72.8958
R2765 vdd.n2948 vdd.n756 72.8958
R2766 vdd.n2981 vdd.n756 72.8958
R2767 vdd.n2334 vdd.n2333 72.8958
R2768 vdd.n2334 vdd.n1055 72.8958
R2769 vdd.n2334 vdd.n1056 72.8958
R2770 vdd.n2334 vdd.n1057 72.8958
R2771 vdd.n2334 vdd.n1058 72.8958
R2772 vdd.n2334 vdd.n1059 72.8958
R2773 vdd.n2334 vdd.n1060 72.8958
R2774 vdd.n2334 vdd.n1061 72.8958
R2775 vdd.n2334 vdd.n1062 72.8958
R2776 vdd.n2334 vdd.n1063 72.8958
R2777 vdd.n2334 vdd.n1064 72.8958
R2778 vdd.n2334 vdd.n1065 72.8958
R2779 vdd.n2334 vdd.n1066 72.8958
R2780 vdd.n2334 vdd.n1067 72.8958
R2781 vdd.n2334 vdd.n1068 72.8958
R2782 vdd.n2334 vdd.n1069 72.8958
R2783 vdd.n2334 vdd.n1070 72.8958
R2784 vdd.n2582 vdd.n923 72.8958
R2785 vdd.n2582 vdd.n924 72.8958
R2786 vdd.n2582 vdd.n925 72.8958
R2787 vdd.n2582 vdd.n926 72.8958
R2788 vdd.n2582 vdd.n927 72.8958
R2789 vdd.n2582 vdd.n928 72.8958
R2790 vdd.n2582 vdd.n929 72.8958
R2791 vdd.n2582 vdd.n930 72.8958
R2792 vdd.n2582 vdd.n931 72.8958
R2793 vdd.n2582 vdd.n932 72.8958
R2794 vdd.n2582 vdd.n933 72.8958
R2795 vdd.n2582 vdd.n934 72.8958
R2796 vdd.n2582 vdd.n935 72.8958
R2797 vdd.n2582 vdd.n936 72.8958
R2798 vdd.n2582 vdd.n937 72.8958
R2799 vdd.n2582 vdd.n938 72.8958
R2800 vdd.n2582 vdd.n939 72.8958
R2801 vdd.n2855 vdd.n2854 72.8958
R2802 vdd.n2855 vdd.n2583 72.8958
R2803 vdd.n2855 vdd.n2584 72.8958
R2804 vdd.n2855 vdd.n2585 72.8958
R2805 vdd.n2855 vdd.n2586 72.8958
R2806 vdd.n2855 vdd.n2587 72.8958
R2807 vdd.n2855 vdd.n2588 72.8958
R2808 vdd.n2855 vdd.n2589 72.8958
R2809 vdd.n2855 vdd.n2590 72.8958
R2810 vdd.n2855 vdd.n2591 72.8958
R2811 vdd.n2855 vdd.n2592 72.8958
R2812 vdd.n2855 vdd.n2593 72.8958
R2813 vdd.n2855 vdd.n2594 72.8958
R2814 vdd.n2855 vdd.n2595 72.8958
R2815 vdd.n2855 vdd.n2596 72.8958
R2816 vdd.n2855 vdd.n2597 72.8958
R2817 vdd.n2855 vdd.n2598 72.8958
R2818 vdd.n3003 vdd.n756 72.8958
R2819 vdd.n3009 vdd.n756 72.8958
R2820 vdd.n802 vdd.n756 72.8958
R2821 vdd.n3016 vdd.n756 72.8958
R2822 vdd.n799 vdd.n756 72.8958
R2823 vdd.n3023 vdd.n756 72.8958
R2824 vdd.n796 vdd.n756 72.8958
R2825 vdd.n3030 vdd.n756 72.8958
R2826 vdd.n793 vdd.n756 72.8958
R2827 vdd.n3038 vdd.n756 72.8958
R2828 vdd.n790 vdd.n756 72.8958
R2829 vdd.n3045 vdd.n756 72.8958
R2830 vdd.n787 vdd.n756 72.8958
R2831 vdd.n3052 vdd.n756 72.8958
R2832 vdd.n784 vdd.n756 72.8958
R2833 vdd.n3059 vdd.n756 72.8958
R2834 vdd.n3062 vdd.n756 72.8958
R2835 vdd.n2582 vdd.n921 72.8958
R2836 vdd.n2582 vdd.n920 72.8958
R2837 vdd.n2582 vdd.n919 72.8958
R2838 vdd.n2582 vdd.n918 72.8958
R2839 vdd.n2582 vdd.n917 72.8958
R2840 vdd.n2582 vdd.n916 72.8958
R2841 vdd.n2582 vdd.n915 72.8958
R2842 vdd.n2582 vdd.n914 72.8958
R2843 vdd.n2582 vdd.n913 72.8958
R2844 vdd.n2582 vdd.n912 72.8958
R2845 vdd.n2582 vdd.n911 72.8958
R2846 vdd.n2582 vdd.n910 72.8958
R2847 vdd.n2582 vdd.n909 72.8958
R2848 vdd.n2582 vdd.n908 72.8958
R2849 vdd.n2582 vdd.n907 72.8958
R2850 vdd.n2582 vdd.n906 72.8958
R2851 vdd.n2582 vdd.n905 72.8958
R2852 vdd.n2335 vdd.n2334 72.8958
R2853 vdd.n2334 vdd.n1071 72.8958
R2854 vdd.n2334 vdd.n1072 72.8958
R2855 vdd.n2334 vdd.n1073 72.8958
R2856 vdd.n2334 vdd.n1074 72.8958
R2857 vdd.n2334 vdd.n1075 72.8958
R2858 vdd.n2334 vdd.n1076 72.8958
R2859 vdd.n2334 vdd.n1077 72.8958
R2860 vdd.n2334 vdd.n1078 72.8958
R2861 vdd.n2334 vdd.n1079 72.8958
R2862 vdd.n2334 vdd.n1080 72.8958
R2863 vdd.n2334 vdd.n1081 72.8958
R2864 vdd.n2334 vdd.n1082 72.8958
R2865 vdd.n2334 vdd.n1083 72.8958
R2866 vdd.n2334 vdd.n1084 72.8958
R2867 vdd.n2334 vdd.n1085 72.8958
R2868 vdd.n2334 vdd.n1086 72.8958
R2869 vdd.n1736 vdd.n1735 66.2847
R2870 vdd.n1736 vdd.n1514 66.2847
R2871 vdd.n1736 vdd.n1515 66.2847
R2872 vdd.n1736 vdd.n1516 66.2847
R2873 vdd.n1736 vdd.n1517 66.2847
R2874 vdd.n1736 vdd.n1518 66.2847
R2875 vdd.n1736 vdd.n1519 66.2847
R2876 vdd.n1736 vdd.n1520 66.2847
R2877 vdd.n1736 vdd.n1521 66.2847
R2878 vdd.n1736 vdd.n1522 66.2847
R2879 vdd.n1736 vdd.n1523 66.2847
R2880 vdd.n1736 vdd.n1524 66.2847
R2881 vdd.n1736 vdd.n1525 66.2847
R2882 vdd.n1736 vdd.n1526 66.2847
R2883 vdd.n1736 vdd.n1527 66.2847
R2884 vdd.n1736 vdd.n1528 66.2847
R2885 vdd.n1736 vdd.n1529 66.2847
R2886 vdd.n1736 vdd.n1530 66.2847
R2887 vdd.n1736 vdd.n1531 66.2847
R2888 vdd.n1736 vdd.n1532 66.2847
R2889 vdd.n1736 vdd.n1533 66.2847
R2890 vdd.n1736 vdd.n1534 66.2847
R2891 vdd.n1736 vdd.n1535 66.2847
R2892 vdd.n1736 vdd.n1536 66.2847
R2893 vdd.n1736 vdd.n1537 66.2847
R2894 vdd.n1736 vdd.n1538 66.2847
R2895 vdd.n1736 vdd.n1539 66.2847
R2896 vdd.n1736 vdd.n1540 66.2847
R2897 vdd.n1736 vdd.n1541 66.2847
R2898 vdd.n1736 vdd.n1542 66.2847
R2899 vdd.n1736 vdd.n1543 66.2847
R2900 vdd.n1404 vdd.n1054 66.2847
R2901 vdd.n1401 vdd.n1054 66.2847
R2902 vdd.n1397 vdd.n1054 66.2847
R2903 vdd.n2196 vdd.n1054 66.2847
R2904 vdd.n1188 vdd.n1054 66.2847
R2905 vdd.n2203 vdd.n1054 66.2847
R2906 vdd.n1181 vdd.n1054 66.2847
R2907 vdd.n2210 vdd.n1054 66.2847
R2908 vdd.n1174 vdd.n1054 66.2847
R2909 vdd.n2217 vdd.n1054 66.2847
R2910 vdd.n1168 vdd.n1054 66.2847
R2911 vdd.n1163 vdd.n1054 66.2847
R2912 vdd.n2228 vdd.n1054 66.2847
R2913 vdd.n1155 vdd.n1054 66.2847
R2914 vdd.n2235 vdd.n1054 66.2847
R2915 vdd.n1148 vdd.n1054 66.2847
R2916 vdd.n2242 vdd.n1054 66.2847
R2917 vdd.n1141 vdd.n1054 66.2847
R2918 vdd.n2249 vdd.n1054 66.2847
R2919 vdd.n1134 vdd.n1054 66.2847
R2920 vdd.n2256 vdd.n1054 66.2847
R2921 vdd.n1128 vdd.n1054 66.2847
R2922 vdd.n1123 vdd.n1054 66.2847
R2923 vdd.n2267 vdd.n1054 66.2847
R2924 vdd.n1115 vdd.n1054 66.2847
R2925 vdd.n2274 vdd.n1054 66.2847
R2926 vdd.n1108 vdd.n1054 66.2847
R2927 vdd.n2281 vdd.n1054 66.2847
R2928 vdd.n1101 vdd.n1054 66.2847
R2929 vdd.n2288 vdd.n1054 66.2847
R2930 vdd.n2293 vdd.n1054 66.2847
R2931 vdd.n1097 vdd.n1054 66.2847
R2932 vdd.n3229 vdd.n658 66.2847
R2933 vdd.n663 vdd.n658 66.2847
R2934 vdd.n666 vdd.n658 66.2847
R2935 vdd.n3218 vdd.n658 66.2847
R2936 vdd.n3212 vdd.n658 66.2847
R2937 vdd.n3210 vdd.n658 66.2847
R2938 vdd.n3204 vdd.n658 66.2847
R2939 vdd.n3202 vdd.n658 66.2847
R2940 vdd.n3196 vdd.n658 66.2847
R2941 vdd.n3194 vdd.n658 66.2847
R2942 vdd.n3188 vdd.n658 66.2847
R2943 vdd.n3186 vdd.n658 66.2847
R2944 vdd.n3180 vdd.n658 66.2847
R2945 vdd.n3178 vdd.n658 66.2847
R2946 vdd.n3172 vdd.n658 66.2847
R2947 vdd.n3170 vdd.n658 66.2847
R2948 vdd.n3164 vdd.n658 66.2847
R2949 vdd.n3162 vdd.n658 66.2847
R2950 vdd.n3156 vdd.n658 66.2847
R2951 vdd.n3154 vdd.n658 66.2847
R2952 vdd.n727 vdd.n658 66.2847
R2953 vdd.n3145 vdd.n658 66.2847
R2954 vdd.n729 vdd.n658 66.2847
R2955 vdd.n3138 vdd.n658 66.2847
R2956 vdd.n3132 vdd.n658 66.2847
R2957 vdd.n3130 vdd.n658 66.2847
R2958 vdd.n3124 vdd.n658 66.2847
R2959 vdd.n3122 vdd.n658 66.2847
R2960 vdd.n3116 vdd.n658 66.2847
R2961 vdd.n750 vdd.n658 66.2847
R2962 vdd.n752 vdd.n658 66.2847
R2963 vdd.n3345 vdd.n3344 66.2847
R2964 vdd.n3345 vdd.n403 66.2847
R2965 vdd.n3345 vdd.n402 66.2847
R2966 vdd.n3345 vdd.n401 66.2847
R2967 vdd.n3345 vdd.n400 66.2847
R2968 vdd.n3345 vdd.n399 66.2847
R2969 vdd.n3345 vdd.n398 66.2847
R2970 vdd.n3345 vdd.n397 66.2847
R2971 vdd.n3345 vdd.n396 66.2847
R2972 vdd.n3345 vdd.n395 66.2847
R2973 vdd.n3345 vdd.n394 66.2847
R2974 vdd.n3345 vdd.n393 66.2847
R2975 vdd.n3345 vdd.n392 66.2847
R2976 vdd.n3345 vdd.n391 66.2847
R2977 vdd.n3345 vdd.n390 66.2847
R2978 vdd.n3345 vdd.n389 66.2847
R2979 vdd.n3345 vdd.n388 66.2847
R2980 vdd.n3345 vdd.n387 66.2847
R2981 vdd.n3345 vdd.n386 66.2847
R2982 vdd.n3345 vdd.n385 66.2847
R2983 vdd.n3345 vdd.n384 66.2847
R2984 vdd.n3345 vdd.n383 66.2847
R2985 vdd.n3345 vdd.n382 66.2847
R2986 vdd.n3345 vdd.n381 66.2847
R2987 vdd.n3345 vdd.n380 66.2847
R2988 vdd.n3345 vdd.n379 66.2847
R2989 vdd.n3345 vdd.n378 66.2847
R2990 vdd.n3345 vdd.n377 66.2847
R2991 vdd.n3345 vdd.n376 66.2847
R2992 vdd.n3345 vdd.n375 66.2847
R2993 vdd.n3345 vdd.n374 66.2847
R2994 vdd.n3345 vdd.n373 66.2847
R2995 vdd.n448 vdd.n373 52.4337
R2996 vdd.n454 vdd.n374 52.4337
R2997 vdd.n458 vdd.n375 52.4337
R2998 vdd.n464 vdd.n376 52.4337
R2999 vdd.n468 vdd.n377 52.4337
R3000 vdd.n474 vdd.n378 52.4337
R3001 vdd.n478 vdd.n379 52.4337
R3002 vdd.n484 vdd.n380 52.4337
R3003 vdd.n488 vdd.n381 52.4337
R3004 vdd.n494 vdd.n382 52.4337
R3005 vdd.n498 vdd.n383 52.4337
R3006 vdd.n504 vdd.n384 52.4337
R3007 vdd.n508 vdd.n385 52.4337
R3008 vdd.n514 vdd.n386 52.4337
R3009 vdd.n518 vdd.n387 52.4337
R3010 vdd.n524 vdd.n388 52.4337
R3011 vdd.n528 vdd.n389 52.4337
R3012 vdd.n534 vdd.n390 52.4337
R3013 vdd.n538 vdd.n391 52.4337
R3014 vdd.n544 vdd.n392 52.4337
R3015 vdd.n548 vdd.n393 52.4337
R3016 vdd.n554 vdd.n394 52.4337
R3017 vdd.n558 vdd.n395 52.4337
R3018 vdd.n564 vdd.n396 52.4337
R3019 vdd.n568 vdd.n397 52.4337
R3020 vdd.n574 vdd.n398 52.4337
R3021 vdd.n578 vdd.n399 52.4337
R3022 vdd.n584 vdd.n400 52.4337
R3023 vdd.n588 vdd.n401 52.4337
R3024 vdd.n594 vdd.n402 52.4337
R3025 vdd.n597 vdd.n403 52.4337
R3026 vdd.n3344 vdd.n3343 52.4337
R3027 vdd.n3229 vdd.n660 52.4337
R3028 vdd.n3227 vdd.n663 52.4337
R3029 vdd.n3223 vdd.n666 52.4337
R3030 vdd.n3219 vdd.n3218 52.4337
R3031 vdd.n3212 vdd.n669 52.4337
R3032 vdd.n3211 vdd.n3210 52.4337
R3033 vdd.n3204 vdd.n675 52.4337
R3034 vdd.n3203 vdd.n3202 52.4337
R3035 vdd.n3196 vdd.n681 52.4337
R3036 vdd.n3195 vdd.n3194 52.4337
R3037 vdd.n3188 vdd.n689 52.4337
R3038 vdd.n3187 vdd.n3186 52.4337
R3039 vdd.n3180 vdd.n695 52.4337
R3040 vdd.n3179 vdd.n3178 52.4337
R3041 vdd.n3172 vdd.n701 52.4337
R3042 vdd.n3171 vdd.n3170 52.4337
R3043 vdd.n3164 vdd.n707 52.4337
R3044 vdd.n3163 vdd.n3162 52.4337
R3045 vdd.n3156 vdd.n713 52.4337
R3046 vdd.n3155 vdd.n3154 52.4337
R3047 vdd.n727 vdd.n719 52.4337
R3048 vdd.n3146 vdd.n3145 52.4337
R3049 vdd.n3143 vdd.n729 52.4337
R3050 vdd.n3139 vdd.n3138 52.4337
R3051 vdd.n3132 vdd.n733 52.4337
R3052 vdd.n3131 vdd.n3130 52.4337
R3053 vdd.n3124 vdd.n739 52.4337
R3054 vdd.n3123 vdd.n3122 52.4337
R3055 vdd.n3116 vdd.n745 52.4337
R3056 vdd.n3115 vdd.n750 52.4337
R3057 vdd.n3111 vdd.n752 52.4337
R3058 vdd.n2295 vdd.n1097 52.4337
R3059 vdd.n2293 vdd.n2292 52.4337
R3060 vdd.n2288 vdd.n2287 52.4337
R3061 vdd.n2283 vdd.n1101 52.4337
R3062 vdd.n2281 vdd.n2280 52.4337
R3063 vdd.n2276 vdd.n1108 52.4337
R3064 vdd.n2274 vdd.n2273 52.4337
R3065 vdd.n2269 vdd.n1115 52.4337
R3066 vdd.n2267 vdd.n2266 52.4337
R3067 vdd.n1124 vdd.n1123 52.4337
R3068 vdd.n2258 vdd.n1128 52.4337
R3069 vdd.n2256 vdd.n2255 52.4337
R3070 vdd.n2251 vdd.n1134 52.4337
R3071 vdd.n2249 vdd.n2248 52.4337
R3072 vdd.n2244 vdd.n1141 52.4337
R3073 vdd.n2242 vdd.n2241 52.4337
R3074 vdd.n2237 vdd.n1148 52.4337
R3075 vdd.n2235 vdd.n2234 52.4337
R3076 vdd.n2230 vdd.n1155 52.4337
R3077 vdd.n2228 vdd.n2227 52.4337
R3078 vdd.n1164 vdd.n1163 52.4337
R3079 vdd.n2219 vdd.n1168 52.4337
R3080 vdd.n2217 vdd.n2216 52.4337
R3081 vdd.n2212 vdd.n1174 52.4337
R3082 vdd.n2210 vdd.n2209 52.4337
R3083 vdd.n2205 vdd.n1181 52.4337
R3084 vdd.n2203 vdd.n2202 52.4337
R3085 vdd.n2198 vdd.n1188 52.4337
R3086 vdd.n2196 vdd.n2195 52.4337
R3087 vdd.n1398 vdd.n1397 52.4337
R3088 vdd.n1402 vdd.n1401 52.4337
R3089 vdd.n2184 vdd.n1404 52.4337
R3090 vdd.n1735 vdd.n1734 52.4337
R3091 vdd.n1549 vdd.n1514 52.4337
R3092 vdd.n1551 vdd.n1515 52.4337
R3093 vdd.n1555 vdd.n1516 52.4337
R3094 vdd.n1557 vdd.n1517 52.4337
R3095 vdd.n1561 vdd.n1518 52.4337
R3096 vdd.n1563 vdd.n1519 52.4337
R3097 vdd.n1567 vdd.n1520 52.4337
R3098 vdd.n1569 vdd.n1521 52.4337
R3099 vdd.n1701 vdd.n1522 52.4337
R3100 vdd.n1573 vdd.n1523 52.4337
R3101 vdd.n1577 vdd.n1524 52.4337
R3102 vdd.n1579 vdd.n1525 52.4337
R3103 vdd.n1583 vdd.n1526 52.4337
R3104 vdd.n1585 vdd.n1527 52.4337
R3105 vdd.n1589 vdd.n1528 52.4337
R3106 vdd.n1591 vdd.n1529 52.4337
R3107 vdd.n1595 vdd.n1530 52.4337
R3108 vdd.n1597 vdd.n1531 52.4337
R3109 vdd.n1601 vdd.n1532 52.4337
R3110 vdd.n1665 vdd.n1533 52.4337
R3111 vdd.n1606 vdd.n1534 52.4337
R3112 vdd.n1608 vdd.n1535 52.4337
R3113 vdd.n1612 vdd.n1536 52.4337
R3114 vdd.n1614 vdd.n1537 52.4337
R3115 vdd.n1618 vdd.n1538 52.4337
R3116 vdd.n1620 vdd.n1539 52.4337
R3117 vdd.n1624 vdd.n1540 52.4337
R3118 vdd.n1626 vdd.n1541 52.4337
R3119 vdd.n1630 vdd.n1542 52.4337
R3120 vdd.n1632 vdd.n1543 52.4337
R3121 vdd.n1735 vdd.n1545 52.4337
R3122 vdd.n1550 vdd.n1514 52.4337
R3123 vdd.n1554 vdd.n1515 52.4337
R3124 vdd.n1556 vdd.n1516 52.4337
R3125 vdd.n1560 vdd.n1517 52.4337
R3126 vdd.n1562 vdd.n1518 52.4337
R3127 vdd.n1566 vdd.n1519 52.4337
R3128 vdd.n1568 vdd.n1520 52.4337
R3129 vdd.n1700 vdd.n1521 52.4337
R3130 vdd.n1572 vdd.n1522 52.4337
R3131 vdd.n1576 vdd.n1523 52.4337
R3132 vdd.n1578 vdd.n1524 52.4337
R3133 vdd.n1582 vdd.n1525 52.4337
R3134 vdd.n1584 vdd.n1526 52.4337
R3135 vdd.n1588 vdd.n1527 52.4337
R3136 vdd.n1590 vdd.n1528 52.4337
R3137 vdd.n1594 vdd.n1529 52.4337
R3138 vdd.n1596 vdd.n1530 52.4337
R3139 vdd.n1600 vdd.n1531 52.4337
R3140 vdd.n1602 vdd.n1532 52.4337
R3141 vdd.n1605 vdd.n1533 52.4337
R3142 vdd.n1607 vdd.n1534 52.4337
R3143 vdd.n1611 vdd.n1535 52.4337
R3144 vdd.n1613 vdd.n1536 52.4337
R3145 vdd.n1617 vdd.n1537 52.4337
R3146 vdd.n1619 vdd.n1538 52.4337
R3147 vdd.n1623 vdd.n1539 52.4337
R3148 vdd.n1625 vdd.n1540 52.4337
R3149 vdd.n1629 vdd.n1541 52.4337
R3150 vdd.n1631 vdd.n1542 52.4337
R3151 vdd.n1543 vdd.n1513 52.4337
R3152 vdd.n1404 vdd.n1403 52.4337
R3153 vdd.n1401 vdd.n1400 52.4337
R3154 vdd.n1397 vdd.n1189 52.4337
R3155 vdd.n2197 vdd.n2196 52.4337
R3156 vdd.n1188 vdd.n1182 52.4337
R3157 vdd.n2204 vdd.n2203 52.4337
R3158 vdd.n1181 vdd.n1175 52.4337
R3159 vdd.n2211 vdd.n2210 52.4337
R3160 vdd.n1174 vdd.n1169 52.4337
R3161 vdd.n2218 vdd.n2217 52.4337
R3162 vdd.n1168 vdd.n1167 52.4337
R3163 vdd.n1163 vdd.n1156 52.4337
R3164 vdd.n2229 vdd.n2228 52.4337
R3165 vdd.n1155 vdd.n1149 52.4337
R3166 vdd.n2236 vdd.n2235 52.4337
R3167 vdd.n1148 vdd.n1142 52.4337
R3168 vdd.n2243 vdd.n2242 52.4337
R3169 vdd.n1141 vdd.n1135 52.4337
R3170 vdd.n2250 vdd.n2249 52.4337
R3171 vdd.n1134 vdd.n1129 52.4337
R3172 vdd.n2257 vdd.n2256 52.4337
R3173 vdd.n1128 vdd.n1127 52.4337
R3174 vdd.n1123 vdd.n1116 52.4337
R3175 vdd.n2268 vdd.n2267 52.4337
R3176 vdd.n1115 vdd.n1109 52.4337
R3177 vdd.n2275 vdd.n2274 52.4337
R3178 vdd.n1108 vdd.n1102 52.4337
R3179 vdd.n2282 vdd.n2281 52.4337
R3180 vdd.n1101 vdd.n1098 52.4337
R3181 vdd.n2289 vdd.n2288 52.4337
R3182 vdd.n2294 vdd.n2293 52.4337
R3183 vdd.n1409 vdd.n1097 52.4337
R3184 vdd.n3230 vdd.n3229 52.4337
R3185 vdd.n3224 vdd.n663 52.4337
R3186 vdd.n3220 vdd.n666 52.4337
R3187 vdd.n3218 vdd.n3217 52.4337
R3188 vdd.n3213 vdd.n3212 52.4337
R3189 vdd.n3210 vdd.n3209 52.4337
R3190 vdd.n3205 vdd.n3204 52.4337
R3191 vdd.n3202 vdd.n3201 52.4337
R3192 vdd.n3197 vdd.n3196 52.4337
R3193 vdd.n3194 vdd.n3193 52.4337
R3194 vdd.n3189 vdd.n3188 52.4337
R3195 vdd.n3186 vdd.n3185 52.4337
R3196 vdd.n3181 vdd.n3180 52.4337
R3197 vdd.n3178 vdd.n3177 52.4337
R3198 vdd.n3173 vdd.n3172 52.4337
R3199 vdd.n3170 vdd.n3169 52.4337
R3200 vdd.n3165 vdd.n3164 52.4337
R3201 vdd.n3162 vdd.n3161 52.4337
R3202 vdd.n3157 vdd.n3156 52.4337
R3203 vdd.n3154 vdd.n3153 52.4337
R3204 vdd.n728 vdd.n727 52.4337
R3205 vdd.n3145 vdd.n3144 52.4337
R3206 vdd.n3140 vdd.n729 52.4337
R3207 vdd.n3138 vdd.n3137 52.4337
R3208 vdd.n3133 vdd.n3132 52.4337
R3209 vdd.n3130 vdd.n3129 52.4337
R3210 vdd.n3125 vdd.n3124 52.4337
R3211 vdd.n3122 vdd.n3121 52.4337
R3212 vdd.n3117 vdd.n3116 52.4337
R3213 vdd.n3112 vdd.n750 52.4337
R3214 vdd.n3108 vdd.n752 52.4337
R3215 vdd.n3344 vdd.n404 52.4337
R3216 vdd.n595 vdd.n403 52.4337
R3217 vdd.n589 vdd.n402 52.4337
R3218 vdd.n585 vdd.n401 52.4337
R3219 vdd.n579 vdd.n400 52.4337
R3220 vdd.n575 vdd.n399 52.4337
R3221 vdd.n569 vdd.n398 52.4337
R3222 vdd.n565 vdd.n397 52.4337
R3223 vdd.n559 vdd.n396 52.4337
R3224 vdd.n555 vdd.n395 52.4337
R3225 vdd.n549 vdd.n394 52.4337
R3226 vdd.n545 vdd.n393 52.4337
R3227 vdd.n539 vdd.n392 52.4337
R3228 vdd.n535 vdd.n391 52.4337
R3229 vdd.n529 vdd.n390 52.4337
R3230 vdd.n525 vdd.n389 52.4337
R3231 vdd.n519 vdd.n388 52.4337
R3232 vdd.n515 vdd.n387 52.4337
R3233 vdd.n509 vdd.n386 52.4337
R3234 vdd.n505 vdd.n385 52.4337
R3235 vdd.n499 vdd.n384 52.4337
R3236 vdd.n495 vdd.n383 52.4337
R3237 vdd.n489 vdd.n382 52.4337
R3238 vdd.n485 vdd.n381 52.4337
R3239 vdd.n479 vdd.n380 52.4337
R3240 vdd.n475 vdd.n379 52.4337
R3241 vdd.n469 vdd.n378 52.4337
R3242 vdd.n465 vdd.n377 52.4337
R3243 vdd.n459 vdd.n376 52.4337
R3244 vdd.n455 vdd.n375 52.4337
R3245 vdd.n449 vdd.n374 52.4337
R3246 vdd.n445 vdd.n373 52.4337
R3247 vdd.t204 vdd.t217 51.4683
R3248 vdd.n266 vdd.n264 42.0461
R3249 vdd.n168 vdd.n166 42.0461
R3250 vdd.n71 vdd.n69 42.0461
R3251 vdd.n2052 vdd.n2050 42.0461
R3252 vdd.n1954 vdd.n1952 42.0461
R3253 vdd.n1857 vdd.n1855 42.0461
R3254 vdd.n320 vdd.n319 41.6884
R3255 vdd.n222 vdd.n221 41.6884
R3256 vdd.n125 vdd.n124 41.6884
R3257 vdd.n2106 vdd.n2105 41.6884
R3258 vdd.n2008 vdd.n2007 41.6884
R3259 vdd.n1911 vdd.n1910 41.6884
R3260 vdd.n1512 vdd.n1511 41.1157
R3261 vdd.n1668 vdd.n1667 41.1157
R3262 vdd.n1704 vdd.n1703 41.1157
R3263 vdd.n407 vdd.n406 41.1157
R3264 vdd.n547 vdd.n420 41.1157
R3265 vdd.n433 vdd.n432 41.1157
R3266 vdd.n3062 vdd.n3061 39.2114
R3267 vdd.n3059 vdd.n3058 39.2114
R3268 vdd.n3054 vdd.n784 39.2114
R3269 vdd.n3052 vdd.n3051 39.2114
R3270 vdd.n3047 vdd.n787 39.2114
R3271 vdd.n3045 vdd.n3044 39.2114
R3272 vdd.n3040 vdd.n790 39.2114
R3273 vdd.n3038 vdd.n3037 39.2114
R3274 vdd.n3032 vdd.n793 39.2114
R3275 vdd.n3030 vdd.n3029 39.2114
R3276 vdd.n3025 vdd.n796 39.2114
R3277 vdd.n3023 vdd.n3022 39.2114
R3278 vdd.n3018 vdd.n799 39.2114
R3279 vdd.n3016 vdd.n3015 39.2114
R3280 vdd.n3011 vdd.n802 39.2114
R3281 vdd.n3009 vdd.n3008 39.2114
R3282 vdd.n3004 vdd.n3003 39.2114
R3283 vdd.n2854 vdd.n2853 39.2114
R3284 vdd.n2848 vdd.n2583 39.2114
R3285 vdd.n2845 vdd.n2584 39.2114
R3286 vdd.n2841 vdd.n2585 39.2114
R3287 vdd.n2837 vdd.n2586 39.2114
R3288 vdd.n2833 vdd.n2587 39.2114
R3289 vdd.n2829 vdd.n2588 39.2114
R3290 vdd.n2825 vdd.n2589 39.2114
R3291 vdd.n2821 vdd.n2590 39.2114
R3292 vdd.n2817 vdd.n2591 39.2114
R3293 vdd.n2813 vdd.n2592 39.2114
R3294 vdd.n2809 vdd.n2593 39.2114
R3295 vdd.n2805 vdd.n2594 39.2114
R3296 vdd.n2801 vdd.n2595 39.2114
R3297 vdd.n2797 vdd.n2596 39.2114
R3298 vdd.n2793 vdd.n2597 39.2114
R3299 vdd.n2788 vdd.n2598 39.2114
R3300 vdd.n2577 vdd.n939 39.2114
R3301 vdd.n2573 vdd.n938 39.2114
R3302 vdd.n2569 vdd.n937 39.2114
R3303 vdd.n2565 vdd.n936 39.2114
R3304 vdd.n2561 vdd.n935 39.2114
R3305 vdd.n2557 vdd.n934 39.2114
R3306 vdd.n2553 vdd.n933 39.2114
R3307 vdd.n2549 vdd.n932 39.2114
R3308 vdd.n2545 vdd.n931 39.2114
R3309 vdd.n2541 vdd.n930 39.2114
R3310 vdd.n2537 vdd.n929 39.2114
R3311 vdd.n2533 vdd.n928 39.2114
R3312 vdd.n2529 vdd.n927 39.2114
R3313 vdd.n2525 vdd.n926 39.2114
R3314 vdd.n2521 vdd.n925 39.2114
R3315 vdd.n2516 vdd.n924 39.2114
R3316 vdd.n2512 vdd.n923 39.2114
R3317 vdd.n2333 vdd.n2332 39.2114
R3318 vdd.n2327 vdd.n1055 39.2114
R3319 vdd.n2324 vdd.n1056 39.2114
R3320 vdd.n2320 vdd.n1057 39.2114
R3321 vdd.n2316 vdd.n1058 39.2114
R3322 vdd.n2312 vdd.n1059 39.2114
R3323 vdd.n2308 vdd.n1060 39.2114
R3324 vdd.n2304 vdd.n1061 39.2114
R3325 vdd.n2300 vdd.n1062 39.2114
R3326 vdd.n1247 vdd.n1063 39.2114
R3327 vdd.n1251 vdd.n1064 39.2114
R3328 vdd.n1255 vdd.n1065 39.2114
R3329 vdd.n1259 vdd.n1066 39.2114
R3330 vdd.n1263 vdd.n1067 39.2114
R3331 vdd.n1267 vdd.n1068 39.2114
R3332 vdd.n1271 vdd.n1069 39.2114
R3333 vdd.n1276 vdd.n1070 39.2114
R3334 vdd.n2981 vdd.n2980 39.2114
R3335 vdd.n2976 vdd.n2948 39.2114
R3336 vdd.n2974 vdd.n2973 39.2114
R3337 vdd.n2969 vdd.n2951 39.2114
R3338 vdd.n2967 vdd.n2966 39.2114
R3339 vdd.n2962 vdd.n2954 39.2114
R3340 vdd.n2960 vdd.n2959 39.2114
R3341 vdd.n2955 vdd.n755 39.2114
R3342 vdd.n3099 vdd.n3098 39.2114
R3343 vdd.n3096 vdd.n3095 39.2114
R3344 vdd.n3091 vdd.n760 39.2114
R3345 vdd.n3089 vdd.n3088 39.2114
R3346 vdd.n3084 vdd.n763 39.2114
R3347 vdd.n3082 vdd.n3081 39.2114
R3348 vdd.n3077 vdd.n766 39.2114
R3349 vdd.n3075 vdd.n3074 39.2114
R3350 vdd.n3070 vdd.n772 39.2114
R3351 vdd.n2857 vdd.n2856 39.2114
R3352 vdd.n2624 vdd.n2599 39.2114
R3353 vdd.n2628 vdd.n2600 39.2114
R3354 vdd.n2632 vdd.n2601 39.2114
R3355 vdd.n2636 vdd.n2602 39.2114
R3356 vdd.n2640 vdd.n2603 39.2114
R3357 vdd.n2644 vdd.n2604 39.2114
R3358 vdd.n2648 vdd.n2605 39.2114
R3359 vdd.n2652 vdd.n2606 39.2114
R3360 vdd.n2656 vdd.n2607 39.2114
R3361 vdd.n2660 vdd.n2608 39.2114
R3362 vdd.n2664 vdd.n2609 39.2114
R3363 vdd.n2668 vdd.n2610 39.2114
R3364 vdd.n2672 vdd.n2611 39.2114
R3365 vdd.n2676 vdd.n2612 39.2114
R3366 vdd.n2680 vdd.n2613 39.2114
R3367 vdd.n2684 vdd.n2614 39.2114
R3368 vdd.n2856 vdd.n904 39.2114
R3369 vdd.n2627 vdd.n2599 39.2114
R3370 vdd.n2631 vdd.n2600 39.2114
R3371 vdd.n2635 vdd.n2601 39.2114
R3372 vdd.n2639 vdd.n2602 39.2114
R3373 vdd.n2643 vdd.n2603 39.2114
R3374 vdd.n2647 vdd.n2604 39.2114
R3375 vdd.n2651 vdd.n2605 39.2114
R3376 vdd.n2655 vdd.n2606 39.2114
R3377 vdd.n2659 vdd.n2607 39.2114
R3378 vdd.n2663 vdd.n2608 39.2114
R3379 vdd.n2667 vdd.n2609 39.2114
R3380 vdd.n2671 vdd.n2610 39.2114
R3381 vdd.n2675 vdd.n2611 39.2114
R3382 vdd.n2679 vdd.n2612 39.2114
R3383 vdd.n2683 vdd.n2613 39.2114
R3384 vdd.n2686 vdd.n2614 39.2114
R3385 vdd.n772 vdd.n767 39.2114
R3386 vdd.n3076 vdd.n3075 39.2114
R3387 vdd.n766 vdd.n764 39.2114
R3388 vdd.n3083 vdd.n3082 39.2114
R3389 vdd.n763 vdd.n761 39.2114
R3390 vdd.n3090 vdd.n3089 39.2114
R3391 vdd.n760 vdd.n758 39.2114
R3392 vdd.n3097 vdd.n3096 39.2114
R3393 vdd.n3100 vdd.n3099 39.2114
R3394 vdd.n2956 vdd.n2955 39.2114
R3395 vdd.n2961 vdd.n2960 39.2114
R3396 vdd.n2954 vdd.n2952 39.2114
R3397 vdd.n2968 vdd.n2967 39.2114
R3398 vdd.n2951 vdd.n2949 39.2114
R3399 vdd.n2975 vdd.n2974 39.2114
R3400 vdd.n2948 vdd.n2946 39.2114
R3401 vdd.n2982 vdd.n2981 39.2114
R3402 vdd.n2333 vdd.n1089 39.2114
R3403 vdd.n2325 vdd.n1055 39.2114
R3404 vdd.n2321 vdd.n1056 39.2114
R3405 vdd.n2317 vdd.n1057 39.2114
R3406 vdd.n2313 vdd.n1058 39.2114
R3407 vdd.n2309 vdd.n1059 39.2114
R3408 vdd.n2305 vdd.n1060 39.2114
R3409 vdd.n2301 vdd.n1061 39.2114
R3410 vdd.n1246 vdd.n1062 39.2114
R3411 vdd.n1250 vdd.n1063 39.2114
R3412 vdd.n1254 vdd.n1064 39.2114
R3413 vdd.n1258 vdd.n1065 39.2114
R3414 vdd.n1262 vdd.n1066 39.2114
R3415 vdd.n1266 vdd.n1067 39.2114
R3416 vdd.n1270 vdd.n1068 39.2114
R3417 vdd.n1275 vdd.n1069 39.2114
R3418 vdd.n1279 vdd.n1070 39.2114
R3419 vdd.n2515 vdd.n923 39.2114
R3420 vdd.n2520 vdd.n924 39.2114
R3421 vdd.n2524 vdd.n925 39.2114
R3422 vdd.n2528 vdd.n926 39.2114
R3423 vdd.n2532 vdd.n927 39.2114
R3424 vdd.n2536 vdd.n928 39.2114
R3425 vdd.n2540 vdd.n929 39.2114
R3426 vdd.n2544 vdd.n930 39.2114
R3427 vdd.n2548 vdd.n931 39.2114
R3428 vdd.n2552 vdd.n932 39.2114
R3429 vdd.n2556 vdd.n933 39.2114
R3430 vdd.n2560 vdd.n934 39.2114
R3431 vdd.n2564 vdd.n935 39.2114
R3432 vdd.n2568 vdd.n936 39.2114
R3433 vdd.n2572 vdd.n937 39.2114
R3434 vdd.n2576 vdd.n938 39.2114
R3435 vdd.n941 vdd.n939 39.2114
R3436 vdd.n2854 vdd.n2617 39.2114
R3437 vdd.n2846 vdd.n2583 39.2114
R3438 vdd.n2842 vdd.n2584 39.2114
R3439 vdd.n2838 vdd.n2585 39.2114
R3440 vdd.n2834 vdd.n2586 39.2114
R3441 vdd.n2830 vdd.n2587 39.2114
R3442 vdd.n2826 vdd.n2588 39.2114
R3443 vdd.n2822 vdd.n2589 39.2114
R3444 vdd.n2818 vdd.n2590 39.2114
R3445 vdd.n2814 vdd.n2591 39.2114
R3446 vdd.n2810 vdd.n2592 39.2114
R3447 vdd.n2806 vdd.n2593 39.2114
R3448 vdd.n2802 vdd.n2594 39.2114
R3449 vdd.n2798 vdd.n2595 39.2114
R3450 vdd.n2794 vdd.n2596 39.2114
R3451 vdd.n2789 vdd.n2597 39.2114
R3452 vdd.n2785 vdd.n2598 39.2114
R3453 vdd.n3003 vdd.n803 39.2114
R3454 vdd.n3010 vdd.n3009 39.2114
R3455 vdd.n802 vdd.n800 39.2114
R3456 vdd.n3017 vdd.n3016 39.2114
R3457 vdd.n799 vdd.n797 39.2114
R3458 vdd.n3024 vdd.n3023 39.2114
R3459 vdd.n796 vdd.n794 39.2114
R3460 vdd.n3031 vdd.n3030 39.2114
R3461 vdd.n793 vdd.n791 39.2114
R3462 vdd.n3039 vdd.n3038 39.2114
R3463 vdd.n790 vdd.n788 39.2114
R3464 vdd.n3046 vdd.n3045 39.2114
R3465 vdd.n787 vdd.n785 39.2114
R3466 vdd.n3053 vdd.n3052 39.2114
R3467 vdd.n784 vdd.n782 39.2114
R3468 vdd.n3060 vdd.n3059 39.2114
R3469 vdd.n3063 vdd.n3062 39.2114
R3470 vdd.n950 vdd.n905 39.2114
R3471 vdd.n2504 vdd.n906 39.2114
R3472 vdd.n2500 vdd.n907 39.2114
R3473 vdd.n2496 vdd.n908 39.2114
R3474 vdd.n2492 vdd.n909 39.2114
R3475 vdd.n2488 vdd.n910 39.2114
R3476 vdd.n2484 vdd.n911 39.2114
R3477 vdd.n2480 vdd.n912 39.2114
R3478 vdd.n2476 vdd.n913 39.2114
R3479 vdd.n2472 vdd.n914 39.2114
R3480 vdd.n2468 vdd.n915 39.2114
R3481 vdd.n2464 vdd.n916 39.2114
R3482 vdd.n2460 vdd.n917 39.2114
R3483 vdd.n2456 vdd.n918 39.2114
R3484 vdd.n2452 vdd.n919 39.2114
R3485 vdd.n2448 vdd.n920 39.2114
R3486 vdd.n2444 vdd.n921 39.2114
R3487 vdd.n2336 vdd.n2335 39.2114
R3488 vdd.n1193 vdd.n1071 39.2114
R3489 vdd.n1197 vdd.n1072 39.2114
R3490 vdd.n1201 vdd.n1073 39.2114
R3491 vdd.n1205 vdd.n1074 39.2114
R3492 vdd.n1209 vdd.n1075 39.2114
R3493 vdd.n1213 vdd.n1076 39.2114
R3494 vdd.n1217 vdd.n1077 39.2114
R3495 vdd.n1221 vdd.n1078 39.2114
R3496 vdd.n1391 vdd.n1079 39.2114
R3497 vdd.n1388 vdd.n1080 39.2114
R3498 vdd.n1384 vdd.n1081 39.2114
R3499 vdd.n1380 vdd.n1082 39.2114
R3500 vdd.n1376 vdd.n1083 39.2114
R3501 vdd.n1372 vdd.n1084 39.2114
R3502 vdd.n1368 vdd.n1085 39.2114
R3503 vdd.n1364 vdd.n1086 39.2114
R3504 vdd.n2441 vdd.n921 39.2114
R3505 vdd.n2445 vdd.n920 39.2114
R3506 vdd.n2449 vdd.n919 39.2114
R3507 vdd.n2453 vdd.n918 39.2114
R3508 vdd.n2457 vdd.n917 39.2114
R3509 vdd.n2461 vdd.n916 39.2114
R3510 vdd.n2465 vdd.n915 39.2114
R3511 vdd.n2469 vdd.n914 39.2114
R3512 vdd.n2473 vdd.n913 39.2114
R3513 vdd.n2477 vdd.n912 39.2114
R3514 vdd.n2481 vdd.n911 39.2114
R3515 vdd.n2485 vdd.n910 39.2114
R3516 vdd.n2489 vdd.n909 39.2114
R3517 vdd.n2493 vdd.n908 39.2114
R3518 vdd.n2497 vdd.n907 39.2114
R3519 vdd.n2501 vdd.n906 39.2114
R3520 vdd.n2505 vdd.n905 39.2114
R3521 vdd.n2335 vdd.n1053 39.2114
R3522 vdd.n1196 vdd.n1071 39.2114
R3523 vdd.n1200 vdd.n1072 39.2114
R3524 vdd.n1204 vdd.n1073 39.2114
R3525 vdd.n1208 vdd.n1074 39.2114
R3526 vdd.n1212 vdd.n1075 39.2114
R3527 vdd.n1216 vdd.n1076 39.2114
R3528 vdd.n1220 vdd.n1077 39.2114
R3529 vdd.n1223 vdd.n1078 39.2114
R3530 vdd.n1389 vdd.n1079 39.2114
R3531 vdd.n1385 vdd.n1080 39.2114
R3532 vdd.n1381 vdd.n1081 39.2114
R3533 vdd.n1377 vdd.n1082 39.2114
R3534 vdd.n1373 vdd.n1083 39.2114
R3535 vdd.n1369 vdd.n1084 39.2114
R3536 vdd.n1365 vdd.n1085 39.2114
R3537 vdd.n1361 vdd.n1086 39.2114
R3538 vdd.n2188 vdd.n2187 37.2369
R3539 vdd.n2224 vdd.n1162 37.2369
R3540 vdd.n2263 vdd.n1122 37.2369
R3541 vdd.n3151 vdd.n724 37.2369
R3542 vdd.n688 vdd.n687 37.2369
R3543 vdd.n3107 vdd.n3106 37.2369
R3544 vdd.n2331 vdd.n1045 31.0639
R3545 vdd.n2580 vdd.n942 31.0639
R3546 vdd.n2513 vdd.n945 31.0639
R3547 vdd.n1281 vdd.n1278 31.0639
R3548 vdd.n2786 vdd.n2783 31.0639
R3549 vdd.n3005 vdd.n3002 31.0639
R3550 vdd.n2852 vdd.n897 31.0639
R3551 vdd.n3066 vdd.n3065 31.0639
R3552 vdd.n2985 vdd.n2984 31.0639
R3553 vdd.n3071 vdd.n771 31.0639
R3554 vdd.n2690 vdd.n2688 31.0639
R3555 vdd.n2859 vdd.n2858 31.0639
R3556 vdd.n2338 vdd.n2337 31.0639
R3557 vdd.n2508 vdd.n2507 31.0639
R3558 vdd.n2440 vdd.n2439 31.0639
R3559 vdd.n1360 vdd.n1359 31.0639
R3560 vdd.n1226 vdd.n1225 30.449
R3561 vdd.n954 vdd.n953 30.449
R3562 vdd.n1273 vdd.n1245 30.449
R3563 vdd.n2518 vdd.n944 30.449
R3564 vdd.n2623 vdd.n2622 30.449
R3565 vdd.n806 vdd.n805 30.449
R3566 vdd.n2791 vdd.n2619 30.449
R3567 vdd.n770 vdd.n769 30.449
R3568 vdd.n1742 vdd.n1508 19.3944
R3569 vdd.n1742 vdd.n1498 19.3944
R3570 vdd.n1754 vdd.n1498 19.3944
R3571 vdd.n1754 vdd.n1496 19.3944
R3572 vdd.n1758 vdd.n1496 19.3944
R3573 vdd.n1758 vdd.n1486 19.3944
R3574 vdd.n1771 vdd.n1486 19.3944
R3575 vdd.n1771 vdd.n1484 19.3944
R3576 vdd.n1775 vdd.n1484 19.3944
R3577 vdd.n1775 vdd.n1476 19.3944
R3578 vdd.n1788 vdd.n1476 19.3944
R3579 vdd.n1788 vdd.n1474 19.3944
R3580 vdd.n1792 vdd.n1474 19.3944
R3581 vdd.n1792 vdd.n1463 19.3944
R3582 vdd.n1804 vdd.n1463 19.3944
R3583 vdd.n1804 vdd.n1461 19.3944
R3584 vdd.n1808 vdd.n1461 19.3944
R3585 vdd.n1808 vdd.n1452 19.3944
R3586 vdd.n2116 vdd.n1452 19.3944
R3587 vdd.n2116 vdd.n1450 19.3944
R3588 vdd.n2120 vdd.n1450 19.3944
R3589 vdd.n2120 vdd.n1441 19.3944
R3590 vdd.n2132 vdd.n1441 19.3944
R3591 vdd.n2132 vdd.n1439 19.3944
R3592 vdd.n2136 vdd.n1439 19.3944
R3593 vdd.n2136 vdd.n1429 19.3944
R3594 vdd.n2149 vdd.n1429 19.3944
R3595 vdd.n2149 vdd.n1427 19.3944
R3596 vdd.n2153 vdd.n1427 19.3944
R3597 vdd.n2153 vdd.n1419 19.3944
R3598 vdd.n2166 vdd.n1419 19.3944
R3599 vdd.n2166 vdd.n1416 19.3944
R3600 vdd.n2172 vdd.n1416 19.3944
R3601 vdd.n2172 vdd.n1417 19.3944
R3602 vdd.n1417 vdd.n1406 19.3944
R3603 vdd.n1661 vdd.n1603 19.3944
R3604 vdd.n1661 vdd.n1660 19.3944
R3605 vdd.n1660 vdd.n1659 19.3944
R3606 vdd.n1659 vdd.n1609 19.3944
R3607 vdd.n1655 vdd.n1609 19.3944
R3608 vdd.n1655 vdd.n1654 19.3944
R3609 vdd.n1654 vdd.n1653 19.3944
R3610 vdd.n1653 vdd.n1615 19.3944
R3611 vdd.n1649 vdd.n1615 19.3944
R3612 vdd.n1649 vdd.n1648 19.3944
R3613 vdd.n1648 vdd.n1647 19.3944
R3614 vdd.n1647 vdd.n1621 19.3944
R3615 vdd.n1643 vdd.n1621 19.3944
R3616 vdd.n1643 vdd.n1642 19.3944
R3617 vdd.n1642 vdd.n1641 19.3944
R3618 vdd.n1641 vdd.n1627 19.3944
R3619 vdd.n1637 vdd.n1627 19.3944
R3620 vdd.n1637 vdd.n1636 19.3944
R3621 vdd.n1636 vdd.n1635 19.3944
R3622 vdd.n1635 vdd.n1633 19.3944
R3623 vdd.n1699 vdd.n1698 19.3944
R3624 vdd.n1698 vdd.n1574 19.3944
R3625 vdd.n1694 vdd.n1574 19.3944
R3626 vdd.n1694 vdd.n1693 19.3944
R3627 vdd.n1693 vdd.n1692 19.3944
R3628 vdd.n1692 vdd.n1580 19.3944
R3629 vdd.n1688 vdd.n1580 19.3944
R3630 vdd.n1688 vdd.n1687 19.3944
R3631 vdd.n1687 vdd.n1686 19.3944
R3632 vdd.n1686 vdd.n1586 19.3944
R3633 vdd.n1682 vdd.n1586 19.3944
R3634 vdd.n1682 vdd.n1681 19.3944
R3635 vdd.n1681 vdd.n1680 19.3944
R3636 vdd.n1680 vdd.n1592 19.3944
R3637 vdd.n1676 vdd.n1592 19.3944
R3638 vdd.n1676 vdd.n1675 19.3944
R3639 vdd.n1675 vdd.n1674 19.3944
R3640 vdd.n1674 vdd.n1598 19.3944
R3641 vdd.n1670 vdd.n1598 19.3944
R3642 vdd.n1670 vdd.n1669 19.3944
R3643 vdd.n1733 vdd.n1732 19.3944
R3644 vdd.n1732 vdd.n1547 19.3944
R3645 vdd.n1728 vdd.n1547 19.3944
R3646 vdd.n1728 vdd.n1727 19.3944
R3647 vdd.n1727 vdd.n1726 19.3944
R3648 vdd.n1726 vdd.n1552 19.3944
R3649 vdd.n1722 vdd.n1552 19.3944
R3650 vdd.n1722 vdd.n1721 19.3944
R3651 vdd.n1721 vdd.n1720 19.3944
R3652 vdd.n1720 vdd.n1558 19.3944
R3653 vdd.n1716 vdd.n1558 19.3944
R3654 vdd.n1716 vdd.n1715 19.3944
R3655 vdd.n1715 vdd.n1714 19.3944
R3656 vdd.n1714 vdd.n1564 19.3944
R3657 vdd.n1710 vdd.n1564 19.3944
R3658 vdd.n1710 vdd.n1709 19.3944
R3659 vdd.n1709 vdd.n1708 19.3944
R3660 vdd.n1708 vdd.n1570 19.3944
R3661 vdd.n2220 vdd.n1160 19.3944
R3662 vdd.n2220 vdd.n1166 19.3944
R3663 vdd.n2215 vdd.n1166 19.3944
R3664 vdd.n2215 vdd.n2214 19.3944
R3665 vdd.n2214 vdd.n2213 19.3944
R3666 vdd.n2213 vdd.n1173 19.3944
R3667 vdd.n2208 vdd.n1173 19.3944
R3668 vdd.n2208 vdd.n2207 19.3944
R3669 vdd.n2207 vdd.n2206 19.3944
R3670 vdd.n2206 vdd.n1180 19.3944
R3671 vdd.n2201 vdd.n1180 19.3944
R3672 vdd.n2201 vdd.n2200 19.3944
R3673 vdd.n2200 vdd.n2199 19.3944
R3674 vdd.n2199 vdd.n1187 19.3944
R3675 vdd.n2194 vdd.n1187 19.3944
R3676 vdd.n2194 vdd.n2193 19.3944
R3677 vdd.n1399 vdd.n1192 19.3944
R3678 vdd.n2189 vdd.n1396 19.3944
R3679 vdd.n2259 vdd.n1120 19.3944
R3680 vdd.n2259 vdd.n1126 19.3944
R3681 vdd.n2254 vdd.n1126 19.3944
R3682 vdd.n2254 vdd.n2253 19.3944
R3683 vdd.n2253 vdd.n2252 19.3944
R3684 vdd.n2252 vdd.n1133 19.3944
R3685 vdd.n2247 vdd.n1133 19.3944
R3686 vdd.n2247 vdd.n2246 19.3944
R3687 vdd.n2246 vdd.n2245 19.3944
R3688 vdd.n2245 vdd.n1140 19.3944
R3689 vdd.n2240 vdd.n1140 19.3944
R3690 vdd.n2240 vdd.n2239 19.3944
R3691 vdd.n2239 vdd.n2238 19.3944
R3692 vdd.n2238 vdd.n1147 19.3944
R3693 vdd.n2233 vdd.n1147 19.3944
R3694 vdd.n2233 vdd.n2232 19.3944
R3695 vdd.n2232 vdd.n2231 19.3944
R3696 vdd.n2231 vdd.n1154 19.3944
R3697 vdd.n2226 vdd.n1154 19.3944
R3698 vdd.n2226 vdd.n2225 19.3944
R3699 vdd.n2296 vdd.n1095 19.3944
R3700 vdd.n2296 vdd.n1096 19.3944
R3701 vdd.n2291 vdd.n2290 19.3944
R3702 vdd.n2286 vdd.n2285 19.3944
R3703 vdd.n2285 vdd.n2284 19.3944
R3704 vdd.n2284 vdd.n1100 19.3944
R3705 vdd.n2279 vdd.n1100 19.3944
R3706 vdd.n2279 vdd.n2278 19.3944
R3707 vdd.n2278 vdd.n2277 19.3944
R3708 vdd.n2277 vdd.n1107 19.3944
R3709 vdd.n2272 vdd.n1107 19.3944
R3710 vdd.n2272 vdd.n2271 19.3944
R3711 vdd.n2271 vdd.n2270 19.3944
R3712 vdd.n2270 vdd.n1114 19.3944
R3713 vdd.n2265 vdd.n1114 19.3944
R3714 vdd.n2265 vdd.n2264 19.3944
R3715 vdd.n1746 vdd.n1504 19.3944
R3716 vdd.n1746 vdd.n1502 19.3944
R3717 vdd.n1750 vdd.n1502 19.3944
R3718 vdd.n1750 vdd.n1492 19.3944
R3719 vdd.n1763 vdd.n1492 19.3944
R3720 vdd.n1763 vdd.n1490 19.3944
R3721 vdd.n1767 vdd.n1490 19.3944
R3722 vdd.n1767 vdd.n1481 19.3944
R3723 vdd.n1780 vdd.n1481 19.3944
R3724 vdd.n1780 vdd.n1479 19.3944
R3725 vdd.n1784 vdd.n1479 19.3944
R3726 vdd.n1784 vdd.n1470 19.3944
R3727 vdd.n1796 vdd.n1470 19.3944
R3728 vdd.n1796 vdd.n1468 19.3944
R3729 vdd.n1800 vdd.n1468 19.3944
R3730 vdd.n1800 vdd.n1458 19.3944
R3731 vdd.n1813 vdd.n1458 19.3944
R3732 vdd.n1813 vdd.n1456 19.3944
R3733 vdd.n2112 vdd.n1456 19.3944
R3734 vdd.n2112 vdd.n1447 19.3944
R3735 vdd.n2124 vdd.n1447 19.3944
R3736 vdd.n2124 vdd.n1445 19.3944
R3737 vdd.n2128 vdd.n1445 19.3944
R3738 vdd.n2128 vdd.n1435 19.3944
R3739 vdd.n2141 vdd.n1435 19.3944
R3740 vdd.n2141 vdd.n1433 19.3944
R3741 vdd.n2145 vdd.n1433 19.3944
R3742 vdd.n2145 vdd.n1424 19.3944
R3743 vdd.n2158 vdd.n1424 19.3944
R3744 vdd.n2158 vdd.n1422 19.3944
R3745 vdd.n2162 vdd.n1422 19.3944
R3746 vdd.n2162 vdd.n1412 19.3944
R3747 vdd.n2176 vdd.n1412 19.3944
R3748 vdd.n2176 vdd.n1410 19.3944
R3749 vdd.n2180 vdd.n1410 19.3944
R3750 vdd.n3239 vdd.n655 19.3944
R3751 vdd.n3243 vdd.n655 19.3944
R3752 vdd.n3243 vdd.n646 19.3944
R3753 vdd.n3255 vdd.n646 19.3944
R3754 vdd.n3255 vdd.n644 19.3944
R3755 vdd.n3259 vdd.n644 19.3944
R3756 vdd.n3259 vdd.n633 19.3944
R3757 vdd.n3271 vdd.n633 19.3944
R3758 vdd.n3271 vdd.n631 19.3944
R3759 vdd.n3275 vdd.n631 19.3944
R3760 vdd.n3275 vdd.n622 19.3944
R3761 vdd.n3288 vdd.n622 19.3944
R3762 vdd.n3288 vdd.n620 19.3944
R3763 vdd.n3295 vdd.n620 19.3944
R3764 vdd.n3295 vdd.n3294 19.3944
R3765 vdd.n3294 vdd.n610 19.3944
R3766 vdd.n3308 vdd.n610 19.3944
R3767 vdd.n3309 vdd.n3308 19.3944
R3768 vdd.n3310 vdd.n3309 19.3944
R3769 vdd.n3310 vdd.n608 19.3944
R3770 vdd.n3315 vdd.n608 19.3944
R3771 vdd.n3316 vdd.n3315 19.3944
R3772 vdd.n3317 vdd.n3316 19.3944
R3773 vdd.n3317 vdd.n606 19.3944
R3774 vdd.n3322 vdd.n606 19.3944
R3775 vdd.n3323 vdd.n3322 19.3944
R3776 vdd.n3324 vdd.n3323 19.3944
R3777 vdd.n3324 vdd.n604 19.3944
R3778 vdd.n3330 vdd.n604 19.3944
R3779 vdd.n3331 vdd.n3330 19.3944
R3780 vdd.n3332 vdd.n3331 19.3944
R3781 vdd.n3332 vdd.n602 19.3944
R3782 vdd.n3337 vdd.n602 19.3944
R3783 vdd.n3338 vdd.n3337 19.3944
R3784 vdd.n3339 vdd.n3338 19.3944
R3785 vdd.n550 vdd.n417 19.3944
R3786 vdd.n556 vdd.n417 19.3944
R3787 vdd.n557 vdd.n556 19.3944
R3788 vdd.n560 vdd.n557 19.3944
R3789 vdd.n560 vdd.n415 19.3944
R3790 vdd.n566 vdd.n415 19.3944
R3791 vdd.n567 vdd.n566 19.3944
R3792 vdd.n570 vdd.n567 19.3944
R3793 vdd.n570 vdd.n413 19.3944
R3794 vdd.n576 vdd.n413 19.3944
R3795 vdd.n577 vdd.n576 19.3944
R3796 vdd.n580 vdd.n577 19.3944
R3797 vdd.n580 vdd.n411 19.3944
R3798 vdd.n586 vdd.n411 19.3944
R3799 vdd.n587 vdd.n586 19.3944
R3800 vdd.n590 vdd.n587 19.3944
R3801 vdd.n590 vdd.n409 19.3944
R3802 vdd.n596 vdd.n409 19.3944
R3803 vdd.n598 vdd.n596 19.3944
R3804 vdd.n599 vdd.n598 19.3944
R3805 vdd.n497 vdd.n496 19.3944
R3806 vdd.n500 vdd.n497 19.3944
R3807 vdd.n500 vdd.n429 19.3944
R3808 vdd.n506 vdd.n429 19.3944
R3809 vdd.n507 vdd.n506 19.3944
R3810 vdd.n510 vdd.n507 19.3944
R3811 vdd.n510 vdd.n427 19.3944
R3812 vdd.n516 vdd.n427 19.3944
R3813 vdd.n517 vdd.n516 19.3944
R3814 vdd.n520 vdd.n517 19.3944
R3815 vdd.n520 vdd.n425 19.3944
R3816 vdd.n526 vdd.n425 19.3944
R3817 vdd.n527 vdd.n526 19.3944
R3818 vdd.n530 vdd.n527 19.3944
R3819 vdd.n530 vdd.n423 19.3944
R3820 vdd.n536 vdd.n423 19.3944
R3821 vdd.n537 vdd.n536 19.3944
R3822 vdd.n540 vdd.n537 19.3944
R3823 vdd.n540 vdd.n421 19.3944
R3824 vdd.n546 vdd.n421 19.3944
R3825 vdd.n447 vdd.n446 19.3944
R3826 vdd.n450 vdd.n447 19.3944
R3827 vdd.n450 vdd.n441 19.3944
R3828 vdd.n456 vdd.n441 19.3944
R3829 vdd.n457 vdd.n456 19.3944
R3830 vdd.n460 vdd.n457 19.3944
R3831 vdd.n460 vdd.n439 19.3944
R3832 vdd.n466 vdd.n439 19.3944
R3833 vdd.n467 vdd.n466 19.3944
R3834 vdd.n470 vdd.n467 19.3944
R3835 vdd.n470 vdd.n437 19.3944
R3836 vdd.n476 vdd.n437 19.3944
R3837 vdd.n477 vdd.n476 19.3944
R3838 vdd.n480 vdd.n477 19.3944
R3839 vdd.n480 vdd.n435 19.3944
R3840 vdd.n486 vdd.n435 19.3944
R3841 vdd.n487 vdd.n486 19.3944
R3842 vdd.n490 vdd.n487 19.3944
R3843 vdd.n3235 vdd.n652 19.3944
R3844 vdd.n3247 vdd.n652 19.3944
R3845 vdd.n3247 vdd.n650 19.3944
R3846 vdd.n3251 vdd.n650 19.3944
R3847 vdd.n3251 vdd.n640 19.3944
R3848 vdd.n3263 vdd.n640 19.3944
R3849 vdd.n3263 vdd.n638 19.3944
R3850 vdd.n3267 vdd.n638 19.3944
R3851 vdd.n3267 vdd.n628 19.3944
R3852 vdd.n3280 vdd.n628 19.3944
R3853 vdd.n3280 vdd.n626 19.3944
R3854 vdd.n3284 vdd.n626 19.3944
R3855 vdd.n3284 vdd.n617 19.3944
R3856 vdd.n3299 vdd.n617 19.3944
R3857 vdd.n3299 vdd.n615 19.3944
R3858 vdd.n3303 vdd.n615 19.3944
R3859 vdd.n3303 vdd.n324 19.3944
R3860 vdd.n3381 vdd.n324 19.3944
R3861 vdd.n3381 vdd.n325 19.3944
R3862 vdd.n3375 vdd.n325 19.3944
R3863 vdd.n3375 vdd.n3374 19.3944
R3864 vdd.n3374 vdd.n3373 19.3944
R3865 vdd.n3373 vdd.n337 19.3944
R3866 vdd.n3367 vdd.n337 19.3944
R3867 vdd.n3367 vdd.n3366 19.3944
R3868 vdd.n3366 vdd.n3365 19.3944
R3869 vdd.n3365 vdd.n347 19.3944
R3870 vdd.n3359 vdd.n347 19.3944
R3871 vdd.n3359 vdd.n3358 19.3944
R3872 vdd.n3358 vdd.n3357 19.3944
R3873 vdd.n3357 vdd.n358 19.3944
R3874 vdd.n3351 vdd.n358 19.3944
R3875 vdd.n3351 vdd.n3350 19.3944
R3876 vdd.n3350 vdd.n3349 19.3944
R3877 vdd.n3349 vdd.n369 19.3944
R3878 vdd.n3192 vdd.n3191 19.3944
R3879 vdd.n3191 vdd.n3190 19.3944
R3880 vdd.n3190 vdd.n694 19.3944
R3881 vdd.n3184 vdd.n694 19.3944
R3882 vdd.n3184 vdd.n3183 19.3944
R3883 vdd.n3183 vdd.n3182 19.3944
R3884 vdd.n3182 vdd.n700 19.3944
R3885 vdd.n3176 vdd.n700 19.3944
R3886 vdd.n3176 vdd.n3175 19.3944
R3887 vdd.n3175 vdd.n3174 19.3944
R3888 vdd.n3174 vdd.n706 19.3944
R3889 vdd.n3168 vdd.n706 19.3944
R3890 vdd.n3168 vdd.n3167 19.3944
R3891 vdd.n3167 vdd.n3166 19.3944
R3892 vdd.n3166 vdd.n712 19.3944
R3893 vdd.n3160 vdd.n712 19.3944
R3894 vdd.n3160 vdd.n3159 19.3944
R3895 vdd.n3159 vdd.n3158 19.3944
R3896 vdd.n3158 vdd.n718 19.3944
R3897 vdd.n3152 vdd.n718 19.3944
R3898 vdd.n3232 vdd.n3231 19.3944
R3899 vdd.n3231 vdd.n662 19.3944
R3900 vdd.n3226 vdd.n3225 19.3944
R3901 vdd.n3222 vdd.n3221 19.3944
R3902 vdd.n3221 vdd.n668 19.3944
R3903 vdd.n3216 vdd.n668 19.3944
R3904 vdd.n3216 vdd.n3215 19.3944
R3905 vdd.n3215 vdd.n3214 19.3944
R3906 vdd.n3214 vdd.n674 19.3944
R3907 vdd.n3208 vdd.n674 19.3944
R3908 vdd.n3208 vdd.n3207 19.3944
R3909 vdd.n3207 vdd.n3206 19.3944
R3910 vdd.n3206 vdd.n680 19.3944
R3911 vdd.n3200 vdd.n680 19.3944
R3912 vdd.n3200 vdd.n3199 19.3944
R3913 vdd.n3199 vdd.n3198 19.3944
R3914 vdd.n3147 vdd.n722 19.3944
R3915 vdd.n3147 vdd.n726 19.3944
R3916 vdd.n3142 vdd.n726 19.3944
R3917 vdd.n3142 vdd.n3141 19.3944
R3918 vdd.n3141 vdd.n732 19.3944
R3919 vdd.n3136 vdd.n732 19.3944
R3920 vdd.n3136 vdd.n3135 19.3944
R3921 vdd.n3135 vdd.n3134 19.3944
R3922 vdd.n3134 vdd.n738 19.3944
R3923 vdd.n3128 vdd.n738 19.3944
R3924 vdd.n3128 vdd.n3127 19.3944
R3925 vdd.n3127 vdd.n3126 19.3944
R3926 vdd.n3126 vdd.n744 19.3944
R3927 vdd.n3120 vdd.n744 19.3944
R3928 vdd.n3120 vdd.n3119 19.3944
R3929 vdd.n3119 vdd.n3118 19.3944
R3930 vdd.n3114 vdd.n3113 19.3944
R3931 vdd.n3110 vdd.n3109 19.3944
R3932 vdd.n1668 vdd.n1603 19.0066
R3933 vdd.n2224 vdd.n1160 19.0066
R3934 vdd.n550 vdd.n547 19.0066
R3935 vdd.n3151 vdd.n722 19.0066
R3936 vdd.n1736 vdd.n1506 18.5924
R3937 vdd.n2182 vdd.n1054 18.5924
R3938 vdd.n3237 vdd.n658 18.5924
R3939 vdd.n3346 vdd.n3345 18.5924
R3940 vdd.n1225 vdd.n1224 16.0975
R3941 vdd.n953 vdd.n952 16.0975
R3942 vdd.n1511 vdd.n1510 16.0975
R3943 vdd.n1667 vdd.n1666 16.0975
R3944 vdd.n1703 vdd.n1702 16.0975
R3945 vdd.n2187 vdd.n2186 16.0975
R3946 vdd.n1162 vdd.n1161 16.0975
R3947 vdd.n1122 vdd.n1121 16.0975
R3948 vdd.n1245 vdd.n1244 16.0975
R3949 vdd.n944 vdd.n943 16.0975
R3950 vdd.n2622 vdd.n2621 16.0975
R3951 vdd.n406 vdd.n405 16.0975
R3952 vdd.n420 vdd.n419 16.0975
R3953 vdd.n432 vdd.n431 16.0975
R3954 vdd.n724 vdd.n723 16.0975
R3955 vdd.n687 vdd.n686 16.0975
R3956 vdd.n805 vdd.n804 16.0975
R3957 vdd.n2619 vdd.n2618 16.0975
R3958 vdd.n3106 vdd.n3105 16.0975
R3959 vdd.n769 vdd.n768 16.0975
R3960 vdd.t217 vdd.n2582 15.4182
R3961 vdd.n2855 vdd.t204 15.4182
R3962 vdd.n28 vdd.n27 14.5238
R3963 vdd.n2334 vdd.n1047 14.0578
R3964 vdd.n3068 vdd.n756 14.0578
R3965 vdd.n316 vdd.n281 13.1884
R3966 vdd.n261 vdd.n226 13.1884
R3967 vdd.n218 vdd.n183 13.1884
R3968 vdd.n163 vdd.n128 13.1884
R3969 vdd.n121 vdd.n86 13.1884
R3970 vdd.n66 vdd.n31 13.1884
R3971 vdd.n2047 vdd.n2012 13.1884
R3972 vdd.n2102 vdd.n2067 13.1884
R3973 vdd.n1949 vdd.n1914 13.1884
R3974 vdd.n2004 vdd.n1969 13.1884
R3975 vdd.n1852 vdd.n1817 13.1884
R3976 vdd.n1907 vdd.n1872 13.1884
R3977 vdd.n1704 vdd.n1699 12.9944
R3978 vdd.n1704 vdd.n1570 12.9944
R3979 vdd.n2263 vdd.n1120 12.9944
R3980 vdd.n2264 vdd.n2263 12.9944
R3981 vdd.n496 vdd.n433 12.9944
R3982 vdd.n490 vdd.n433 12.9944
R3983 vdd.n3192 vdd.n688 12.9944
R3984 vdd.n3198 vdd.n688 12.9944
R3985 vdd.n317 vdd.n279 12.8005
R3986 vdd.n312 vdd.n283 12.8005
R3987 vdd.n262 vdd.n224 12.8005
R3988 vdd.n257 vdd.n228 12.8005
R3989 vdd.n219 vdd.n181 12.8005
R3990 vdd.n214 vdd.n185 12.8005
R3991 vdd.n164 vdd.n126 12.8005
R3992 vdd.n159 vdd.n130 12.8005
R3993 vdd.n122 vdd.n84 12.8005
R3994 vdd.n117 vdd.n88 12.8005
R3995 vdd.n67 vdd.n29 12.8005
R3996 vdd.n62 vdd.n33 12.8005
R3997 vdd.n2048 vdd.n2010 12.8005
R3998 vdd.n2043 vdd.n2014 12.8005
R3999 vdd.n2103 vdd.n2065 12.8005
R4000 vdd.n2098 vdd.n2069 12.8005
R4001 vdd.n1950 vdd.n1912 12.8005
R4002 vdd.n1945 vdd.n1916 12.8005
R4003 vdd.n2005 vdd.n1967 12.8005
R4004 vdd.n2000 vdd.n1971 12.8005
R4005 vdd.n1853 vdd.n1815 12.8005
R4006 vdd.n1848 vdd.n1819 12.8005
R4007 vdd.n1908 vdd.n1870 12.8005
R4008 vdd.n1903 vdd.n1874 12.8005
R4009 vdd.n311 vdd.n284 12.0247
R4010 vdd.n256 vdd.n229 12.0247
R4011 vdd.n213 vdd.n186 12.0247
R4012 vdd.n158 vdd.n131 12.0247
R4013 vdd.n116 vdd.n89 12.0247
R4014 vdd.n61 vdd.n34 12.0247
R4015 vdd.n2042 vdd.n2015 12.0247
R4016 vdd.n2097 vdd.n2070 12.0247
R4017 vdd.n1944 vdd.n1917 12.0247
R4018 vdd.n1999 vdd.n1972 12.0247
R4019 vdd.n1847 vdd.n1820 12.0247
R4020 vdd.n1902 vdd.n1875 12.0247
R4021 vdd.n1744 vdd.n1506 11.337
R4022 vdd.n1752 vdd.n1500 11.337
R4023 vdd.n1752 vdd.n1494 11.337
R4024 vdd.n1761 vdd.n1494 11.337
R4025 vdd.n1769 vdd.n1488 11.337
R4026 vdd.n1778 vdd.n1777 11.337
R4027 vdd.n1794 vdd.n1472 11.337
R4028 vdd.n1802 vdd.n1465 11.337
R4029 vdd.n1811 vdd.n1810 11.337
R4030 vdd.n2114 vdd.n1454 11.337
R4031 vdd.n2130 vdd.n1443 11.337
R4032 vdd.n2139 vdd.n1437 11.337
R4033 vdd.n2147 vdd.n1431 11.337
R4034 vdd.n2156 vdd.n2155 11.337
R4035 vdd.n2164 vdd.n1414 11.337
R4036 vdd.n2174 vdd.n1414 11.337
R4037 vdd.n2182 vdd.n1407 11.337
R4038 vdd.n3237 vdd.n659 11.337
R4039 vdd.n3245 vdd.n648 11.337
R4040 vdd.n3253 vdd.n648 11.337
R4041 vdd.n3261 vdd.n642 11.337
R4042 vdd.n3269 vdd.n635 11.337
R4043 vdd.n3278 vdd.n3277 11.337
R4044 vdd.n3286 vdd.n624 11.337
R4045 vdd.n3305 vdd.n613 11.337
R4046 vdd.n3379 vdd.n328 11.337
R4047 vdd.n3377 vdd.n332 11.337
R4048 vdd.n3371 vdd.n3370 11.337
R4049 vdd.n3363 vdd.n349 11.337
R4050 vdd.n3362 vdd.n3361 11.337
R4051 vdd.n3355 vdd.n3354 11.337
R4052 vdd.n3354 vdd.n3353 11.337
R4053 vdd.n3353 vdd.n363 11.337
R4054 vdd.n3347 vdd.n3346 11.337
R4055 vdd.n308 vdd.n307 11.249
R4056 vdd.n253 vdd.n252 11.249
R4057 vdd.n210 vdd.n209 11.249
R4058 vdd.n155 vdd.n154 11.249
R4059 vdd.n113 vdd.n112 11.249
R4060 vdd.n58 vdd.n57 11.249
R4061 vdd.n2039 vdd.n2038 11.249
R4062 vdd.n2094 vdd.n2093 11.249
R4063 vdd.n1941 vdd.n1940 11.249
R4064 vdd.n1996 vdd.n1995 11.249
R4065 vdd.n1844 vdd.n1843 11.249
R4066 vdd.n1899 vdd.n1898 11.249
R4067 vdd.n2164 vdd.t169 10.7702
R4068 vdd.n3253 vdd.t161 10.7702
R4069 vdd.n293 vdd.n292 10.7238
R4070 vdd.n238 vdd.n237 10.7238
R4071 vdd.n195 vdd.n194 10.7238
R4072 vdd.n140 vdd.n139 10.7238
R4073 vdd.n98 vdd.n97 10.7238
R4074 vdd.n43 vdd.n42 10.7238
R4075 vdd.n2024 vdd.n2023 10.7238
R4076 vdd.n2079 vdd.n2078 10.7238
R4077 vdd.n1926 vdd.n1925 10.7238
R4078 vdd.n1981 vdd.n1980 10.7238
R4079 vdd.n1829 vdd.n1828 10.7238
R4080 vdd.n1884 vdd.n1883 10.7238
R4081 vdd.n2510 vdd.t235 10.6568
R4082 vdd.t220 vdd.n899 10.6568
R4083 vdd.n2343 vdd.n1045 10.6151
R4084 vdd.n2344 vdd.n2343 10.6151
R4085 vdd.n2345 vdd.n2344 10.6151
R4086 vdd.n2345 vdd.n1034 10.6151
R4087 vdd.n2355 vdd.n1034 10.6151
R4088 vdd.n2356 vdd.n2355 10.6151
R4089 vdd.n2357 vdd.n2356 10.6151
R4090 vdd.n2357 vdd.n1021 10.6151
R4091 vdd.n2367 vdd.n1021 10.6151
R4092 vdd.n2368 vdd.n2367 10.6151
R4093 vdd.n2369 vdd.n2368 10.6151
R4094 vdd.n2369 vdd.n1009 10.6151
R4095 vdd.n2380 vdd.n1009 10.6151
R4096 vdd.n2381 vdd.n2380 10.6151
R4097 vdd.n2382 vdd.n2381 10.6151
R4098 vdd.n2382 vdd.n997 10.6151
R4099 vdd.n2392 vdd.n997 10.6151
R4100 vdd.n2393 vdd.n2392 10.6151
R4101 vdd.n2394 vdd.n2393 10.6151
R4102 vdd.n2394 vdd.n985 10.6151
R4103 vdd.n2404 vdd.n985 10.6151
R4104 vdd.n2405 vdd.n2404 10.6151
R4105 vdd.n2406 vdd.n2405 10.6151
R4106 vdd.n2406 vdd.n974 10.6151
R4107 vdd.n2416 vdd.n974 10.6151
R4108 vdd.n2417 vdd.n2416 10.6151
R4109 vdd.n2418 vdd.n2417 10.6151
R4110 vdd.n2418 vdd.n961 10.6151
R4111 vdd.n2430 vdd.n961 10.6151
R4112 vdd.n2431 vdd.n2430 10.6151
R4113 vdd.n2433 vdd.n2431 10.6151
R4114 vdd.n2433 vdd.n2432 10.6151
R4115 vdd.n2432 vdd.n942 10.6151
R4116 vdd.n2580 vdd.n2579 10.6151
R4117 vdd.n2579 vdd.n2578 10.6151
R4118 vdd.n2578 vdd.n2575 10.6151
R4119 vdd.n2575 vdd.n2574 10.6151
R4120 vdd.n2574 vdd.n2571 10.6151
R4121 vdd.n2571 vdd.n2570 10.6151
R4122 vdd.n2570 vdd.n2567 10.6151
R4123 vdd.n2567 vdd.n2566 10.6151
R4124 vdd.n2566 vdd.n2563 10.6151
R4125 vdd.n2563 vdd.n2562 10.6151
R4126 vdd.n2562 vdd.n2559 10.6151
R4127 vdd.n2559 vdd.n2558 10.6151
R4128 vdd.n2558 vdd.n2555 10.6151
R4129 vdd.n2555 vdd.n2554 10.6151
R4130 vdd.n2554 vdd.n2551 10.6151
R4131 vdd.n2551 vdd.n2550 10.6151
R4132 vdd.n2550 vdd.n2547 10.6151
R4133 vdd.n2547 vdd.n2546 10.6151
R4134 vdd.n2546 vdd.n2543 10.6151
R4135 vdd.n2543 vdd.n2542 10.6151
R4136 vdd.n2542 vdd.n2539 10.6151
R4137 vdd.n2539 vdd.n2538 10.6151
R4138 vdd.n2538 vdd.n2535 10.6151
R4139 vdd.n2535 vdd.n2534 10.6151
R4140 vdd.n2534 vdd.n2531 10.6151
R4141 vdd.n2531 vdd.n2530 10.6151
R4142 vdd.n2530 vdd.n2527 10.6151
R4143 vdd.n2527 vdd.n2526 10.6151
R4144 vdd.n2526 vdd.n2523 10.6151
R4145 vdd.n2523 vdd.n2522 10.6151
R4146 vdd.n2522 vdd.n2519 10.6151
R4147 vdd.n2517 vdd.n2514 10.6151
R4148 vdd.n2514 vdd.n2513 10.6151
R4149 vdd.n1282 vdd.n1281 10.6151
R4150 vdd.n1284 vdd.n1282 10.6151
R4151 vdd.n1285 vdd.n1284 10.6151
R4152 vdd.n1287 vdd.n1285 10.6151
R4153 vdd.n1288 vdd.n1287 10.6151
R4154 vdd.n1290 vdd.n1288 10.6151
R4155 vdd.n1291 vdd.n1290 10.6151
R4156 vdd.n1293 vdd.n1291 10.6151
R4157 vdd.n1294 vdd.n1293 10.6151
R4158 vdd.n1296 vdd.n1294 10.6151
R4159 vdd.n1297 vdd.n1296 10.6151
R4160 vdd.n1299 vdd.n1297 10.6151
R4161 vdd.n1300 vdd.n1299 10.6151
R4162 vdd.n1302 vdd.n1300 10.6151
R4163 vdd.n1303 vdd.n1302 10.6151
R4164 vdd.n1305 vdd.n1303 10.6151
R4165 vdd.n1306 vdd.n1305 10.6151
R4166 vdd.n1328 vdd.n1306 10.6151
R4167 vdd.n1328 vdd.n1327 10.6151
R4168 vdd.n1327 vdd.n1326 10.6151
R4169 vdd.n1326 vdd.n1324 10.6151
R4170 vdd.n1324 vdd.n1323 10.6151
R4171 vdd.n1323 vdd.n1321 10.6151
R4172 vdd.n1321 vdd.n1320 10.6151
R4173 vdd.n1320 vdd.n1318 10.6151
R4174 vdd.n1318 vdd.n1317 10.6151
R4175 vdd.n1317 vdd.n1315 10.6151
R4176 vdd.n1315 vdd.n1314 10.6151
R4177 vdd.n1314 vdd.n1312 10.6151
R4178 vdd.n1312 vdd.n1311 10.6151
R4179 vdd.n1311 vdd.n1308 10.6151
R4180 vdd.n1308 vdd.n1307 10.6151
R4181 vdd.n1307 vdd.n945 10.6151
R4182 vdd.n2331 vdd.n2330 10.6151
R4183 vdd.n2330 vdd.n2329 10.6151
R4184 vdd.n2329 vdd.n2328 10.6151
R4185 vdd.n2328 vdd.n2326 10.6151
R4186 vdd.n2326 vdd.n2323 10.6151
R4187 vdd.n2323 vdd.n2322 10.6151
R4188 vdd.n2322 vdd.n2319 10.6151
R4189 vdd.n2319 vdd.n2318 10.6151
R4190 vdd.n2318 vdd.n2315 10.6151
R4191 vdd.n2315 vdd.n2314 10.6151
R4192 vdd.n2314 vdd.n2311 10.6151
R4193 vdd.n2311 vdd.n2310 10.6151
R4194 vdd.n2310 vdd.n2307 10.6151
R4195 vdd.n2307 vdd.n2306 10.6151
R4196 vdd.n2306 vdd.n2303 10.6151
R4197 vdd.n2303 vdd.n2302 10.6151
R4198 vdd.n2302 vdd.n2299 10.6151
R4199 vdd.n2299 vdd.n1090 10.6151
R4200 vdd.n1248 vdd.n1090 10.6151
R4201 vdd.n1249 vdd.n1248 10.6151
R4202 vdd.n1252 vdd.n1249 10.6151
R4203 vdd.n1253 vdd.n1252 10.6151
R4204 vdd.n1256 vdd.n1253 10.6151
R4205 vdd.n1257 vdd.n1256 10.6151
R4206 vdd.n1260 vdd.n1257 10.6151
R4207 vdd.n1261 vdd.n1260 10.6151
R4208 vdd.n1264 vdd.n1261 10.6151
R4209 vdd.n1265 vdd.n1264 10.6151
R4210 vdd.n1268 vdd.n1265 10.6151
R4211 vdd.n1269 vdd.n1268 10.6151
R4212 vdd.n1272 vdd.n1269 10.6151
R4213 vdd.n1277 vdd.n1274 10.6151
R4214 vdd.n1278 vdd.n1277 10.6151
R4215 vdd.n2783 vdd.n2782 10.6151
R4216 vdd.n2782 vdd.n2781 10.6151
R4217 vdd.n2781 vdd.n2620 10.6151
R4218 vdd.n2725 vdd.n2620 10.6151
R4219 vdd.n2726 vdd.n2725 10.6151
R4220 vdd.n2728 vdd.n2726 10.6151
R4221 vdd.n2729 vdd.n2728 10.6151
R4222 vdd.n2731 vdd.n2729 10.6151
R4223 vdd.n2732 vdd.n2731 10.6151
R4224 vdd.n2762 vdd.n2732 10.6151
R4225 vdd.n2762 vdd.n2761 10.6151
R4226 vdd.n2761 vdd.n2760 10.6151
R4227 vdd.n2760 vdd.n2758 10.6151
R4228 vdd.n2758 vdd.n2757 10.6151
R4229 vdd.n2757 vdd.n2755 10.6151
R4230 vdd.n2755 vdd.n2754 10.6151
R4231 vdd.n2754 vdd.n2752 10.6151
R4232 vdd.n2752 vdd.n2751 10.6151
R4233 vdd.n2751 vdd.n2749 10.6151
R4234 vdd.n2749 vdd.n2748 10.6151
R4235 vdd.n2748 vdd.n2746 10.6151
R4236 vdd.n2746 vdd.n2745 10.6151
R4237 vdd.n2745 vdd.n2743 10.6151
R4238 vdd.n2743 vdd.n2742 10.6151
R4239 vdd.n2742 vdd.n2740 10.6151
R4240 vdd.n2740 vdd.n2739 10.6151
R4241 vdd.n2739 vdd.n2737 10.6151
R4242 vdd.n2737 vdd.n2736 10.6151
R4243 vdd.n2736 vdd.n2734 10.6151
R4244 vdd.n2734 vdd.n2733 10.6151
R4245 vdd.n2733 vdd.n807 10.6151
R4246 vdd.n3001 vdd.n807 10.6151
R4247 vdd.n3002 vdd.n3001 10.6151
R4248 vdd.n2852 vdd.n2851 10.6151
R4249 vdd.n2851 vdd.n2850 10.6151
R4250 vdd.n2850 vdd.n2849 10.6151
R4251 vdd.n2849 vdd.n2847 10.6151
R4252 vdd.n2847 vdd.n2844 10.6151
R4253 vdd.n2844 vdd.n2843 10.6151
R4254 vdd.n2843 vdd.n2840 10.6151
R4255 vdd.n2840 vdd.n2839 10.6151
R4256 vdd.n2839 vdd.n2836 10.6151
R4257 vdd.n2836 vdd.n2835 10.6151
R4258 vdd.n2835 vdd.n2832 10.6151
R4259 vdd.n2832 vdd.n2831 10.6151
R4260 vdd.n2831 vdd.n2828 10.6151
R4261 vdd.n2828 vdd.n2827 10.6151
R4262 vdd.n2827 vdd.n2824 10.6151
R4263 vdd.n2824 vdd.n2823 10.6151
R4264 vdd.n2823 vdd.n2820 10.6151
R4265 vdd.n2820 vdd.n2819 10.6151
R4266 vdd.n2819 vdd.n2816 10.6151
R4267 vdd.n2816 vdd.n2815 10.6151
R4268 vdd.n2815 vdd.n2812 10.6151
R4269 vdd.n2812 vdd.n2811 10.6151
R4270 vdd.n2811 vdd.n2808 10.6151
R4271 vdd.n2808 vdd.n2807 10.6151
R4272 vdd.n2807 vdd.n2804 10.6151
R4273 vdd.n2804 vdd.n2803 10.6151
R4274 vdd.n2803 vdd.n2800 10.6151
R4275 vdd.n2800 vdd.n2799 10.6151
R4276 vdd.n2799 vdd.n2796 10.6151
R4277 vdd.n2796 vdd.n2795 10.6151
R4278 vdd.n2795 vdd.n2792 10.6151
R4279 vdd.n2790 vdd.n2787 10.6151
R4280 vdd.n2787 vdd.n2786 10.6151
R4281 vdd.n2864 vdd.n897 10.6151
R4282 vdd.n2865 vdd.n2864 10.6151
R4283 vdd.n2866 vdd.n2865 10.6151
R4284 vdd.n2866 vdd.n886 10.6151
R4285 vdd.n2876 vdd.n886 10.6151
R4286 vdd.n2877 vdd.n2876 10.6151
R4287 vdd.n2878 vdd.n2877 10.6151
R4288 vdd.n2878 vdd.n874 10.6151
R4289 vdd.n2888 vdd.n874 10.6151
R4290 vdd.n2889 vdd.n2888 10.6151
R4291 vdd.n2890 vdd.n2889 10.6151
R4292 vdd.n2890 vdd.n862 10.6151
R4293 vdd.n2900 vdd.n862 10.6151
R4294 vdd.n2901 vdd.n2900 10.6151
R4295 vdd.n2902 vdd.n2901 10.6151
R4296 vdd.n2902 vdd.n851 10.6151
R4297 vdd.n2912 vdd.n851 10.6151
R4298 vdd.n2913 vdd.n2912 10.6151
R4299 vdd.n2914 vdd.n2913 10.6151
R4300 vdd.n2914 vdd.n837 10.6151
R4301 vdd.n2925 vdd.n837 10.6151
R4302 vdd.n2926 vdd.n2925 10.6151
R4303 vdd.n2927 vdd.n2926 10.6151
R4304 vdd.n2927 vdd.n826 10.6151
R4305 vdd.n2937 vdd.n826 10.6151
R4306 vdd.n2938 vdd.n2937 10.6151
R4307 vdd.n2939 vdd.n2938 10.6151
R4308 vdd.n2939 vdd.n812 10.6151
R4309 vdd.n2994 vdd.n812 10.6151
R4310 vdd.n2995 vdd.n2994 10.6151
R4311 vdd.n2996 vdd.n2995 10.6151
R4312 vdd.n2996 vdd.n779 10.6151
R4313 vdd.n3066 vdd.n779 10.6151
R4314 vdd.n3065 vdd.n3064 10.6151
R4315 vdd.n3064 vdd.n780 10.6151
R4316 vdd.n781 vdd.n780 10.6151
R4317 vdd.n3057 vdd.n781 10.6151
R4318 vdd.n3057 vdd.n3056 10.6151
R4319 vdd.n3056 vdd.n3055 10.6151
R4320 vdd.n3055 vdd.n783 10.6151
R4321 vdd.n3050 vdd.n783 10.6151
R4322 vdd.n3050 vdd.n3049 10.6151
R4323 vdd.n3049 vdd.n3048 10.6151
R4324 vdd.n3048 vdd.n786 10.6151
R4325 vdd.n3043 vdd.n786 10.6151
R4326 vdd.n3043 vdd.n3042 10.6151
R4327 vdd.n3042 vdd.n3041 10.6151
R4328 vdd.n3041 vdd.n789 10.6151
R4329 vdd.n3036 vdd.n789 10.6151
R4330 vdd.n3036 vdd.n3035 10.6151
R4331 vdd.n3035 vdd.n3033 10.6151
R4332 vdd.n3033 vdd.n792 10.6151
R4333 vdd.n3028 vdd.n792 10.6151
R4334 vdd.n3028 vdd.n3027 10.6151
R4335 vdd.n3027 vdd.n3026 10.6151
R4336 vdd.n3026 vdd.n795 10.6151
R4337 vdd.n3021 vdd.n795 10.6151
R4338 vdd.n3021 vdd.n3020 10.6151
R4339 vdd.n3020 vdd.n3019 10.6151
R4340 vdd.n3019 vdd.n798 10.6151
R4341 vdd.n3014 vdd.n798 10.6151
R4342 vdd.n3014 vdd.n3013 10.6151
R4343 vdd.n3013 vdd.n3012 10.6151
R4344 vdd.n3012 vdd.n801 10.6151
R4345 vdd.n3007 vdd.n3006 10.6151
R4346 vdd.n3006 vdd.n3005 10.6151
R4347 vdd.n2984 vdd.n2945 10.6151
R4348 vdd.n2979 vdd.n2945 10.6151
R4349 vdd.n2979 vdd.n2978 10.6151
R4350 vdd.n2978 vdd.n2977 10.6151
R4351 vdd.n2977 vdd.n2947 10.6151
R4352 vdd.n2972 vdd.n2947 10.6151
R4353 vdd.n2972 vdd.n2971 10.6151
R4354 vdd.n2971 vdd.n2970 10.6151
R4355 vdd.n2970 vdd.n2950 10.6151
R4356 vdd.n2965 vdd.n2950 10.6151
R4357 vdd.n2965 vdd.n2964 10.6151
R4358 vdd.n2964 vdd.n2963 10.6151
R4359 vdd.n2963 vdd.n2953 10.6151
R4360 vdd.n2958 vdd.n2953 10.6151
R4361 vdd.n2958 vdd.n2957 10.6151
R4362 vdd.n2957 vdd.n753 10.6151
R4363 vdd.n3101 vdd.n753 10.6151
R4364 vdd.n3101 vdd.n754 10.6151
R4365 vdd.n757 vdd.n754 10.6151
R4366 vdd.n3094 vdd.n757 10.6151
R4367 vdd.n3094 vdd.n3093 10.6151
R4368 vdd.n3093 vdd.n3092 10.6151
R4369 vdd.n3092 vdd.n759 10.6151
R4370 vdd.n3087 vdd.n759 10.6151
R4371 vdd.n3087 vdd.n3086 10.6151
R4372 vdd.n3086 vdd.n3085 10.6151
R4373 vdd.n3085 vdd.n762 10.6151
R4374 vdd.n3080 vdd.n762 10.6151
R4375 vdd.n3080 vdd.n3079 10.6151
R4376 vdd.n3079 vdd.n3078 10.6151
R4377 vdd.n3078 vdd.n765 10.6151
R4378 vdd.n3073 vdd.n3072 10.6151
R4379 vdd.n3072 vdd.n3071 10.6151
R4380 vdd.n2691 vdd.n2690 10.6151
R4381 vdd.n2777 vdd.n2691 10.6151
R4382 vdd.n2777 vdd.n2776 10.6151
R4383 vdd.n2776 vdd.n2775 10.6151
R4384 vdd.n2775 vdd.n2773 10.6151
R4385 vdd.n2773 vdd.n2772 10.6151
R4386 vdd.n2772 vdd.n2770 10.6151
R4387 vdd.n2770 vdd.n2769 10.6151
R4388 vdd.n2769 vdd.n2767 10.6151
R4389 vdd.n2767 vdd.n2766 10.6151
R4390 vdd.n2766 vdd.n2723 10.6151
R4391 vdd.n2723 vdd.n2722 10.6151
R4392 vdd.n2722 vdd.n2720 10.6151
R4393 vdd.n2720 vdd.n2719 10.6151
R4394 vdd.n2719 vdd.n2717 10.6151
R4395 vdd.n2717 vdd.n2716 10.6151
R4396 vdd.n2716 vdd.n2714 10.6151
R4397 vdd.n2714 vdd.n2713 10.6151
R4398 vdd.n2713 vdd.n2711 10.6151
R4399 vdd.n2711 vdd.n2710 10.6151
R4400 vdd.n2710 vdd.n2708 10.6151
R4401 vdd.n2708 vdd.n2707 10.6151
R4402 vdd.n2707 vdd.n2705 10.6151
R4403 vdd.n2705 vdd.n2704 10.6151
R4404 vdd.n2704 vdd.n2702 10.6151
R4405 vdd.n2702 vdd.n2701 10.6151
R4406 vdd.n2701 vdd.n2699 10.6151
R4407 vdd.n2699 vdd.n2698 10.6151
R4408 vdd.n2698 vdd.n2696 10.6151
R4409 vdd.n2696 vdd.n2695 10.6151
R4410 vdd.n2695 vdd.n2693 10.6151
R4411 vdd.n2693 vdd.n2692 10.6151
R4412 vdd.n2692 vdd.n771 10.6151
R4413 vdd.n2858 vdd.n903 10.6151
R4414 vdd.n2625 vdd.n903 10.6151
R4415 vdd.n2626 vdd.n2625 10.6151
R4416 vdd.n2629 vdd.n2626 10.6151
R4417 vdd.n2630 vdd.n2629 10.6151
R4418 vdd.n2633 vdd.n2630 10.6151
R4419 vdd.n2634 vdd.n2633 10.6151
R4420 vdd.n2637 vdd.n2634 10.6151
R4421 vdd.n2638 vdd.n2637 10.6151
R4422 vdd.n2641 vdd.n2638 10.6151
R4423 vdd.n2642 vdd.n2641 10.6151
R4424 vdd.n2645 vdd.n2642 10.6151
R4425 vdd.n2646 vdd.n2645 10.6151
R4426 vdd.n2649 vdd.n2646 10.6151
R4427 vdd.n2650 vdd.n2649 10.6151
R4428 vdd.n2653 vdd.n2650 10.6151
R4429 vdd.n2654 vdd.n2653 10.6151
R4430 vdd.n2657 vdd.n2654 10.6151
R4431 vdd.n2658 vdd.n2657 10.6151
R4432 vdd.n2661 vdd.n2658 10.6151
R4433 vdd.n2662 vdd.n2661 10.6151
R4434 vdd.n2665 vdd.n2662 10.6151
R4435 vdd.n2666 vdd.n2665 10.6151
R4436 vdd.n2669 vdd.n2666 10.6151
R4437 vdd.n2670 vdd.n2669 10.6151
R4438 vdd.n2673 vdd.n2670 10.6151
R4439 vdd.n2674 vdd.n2673 10.6151
R4440 vdd.n2677 vdd.n2674 10.6151
R4441 vdd.n2678 vdd.n2677 10.6151
R4442 vdd.n2681 vdd.n2678 10.6151
R4443 vdd.n2682 vdd.n2681 10.6151
R4444 vdd.n2687 vdd.n2685 10.6151
R4445 vdd.n2688 vdd.n2687 10.6151
R4446 vdd.n2860 vdd.n2859 10.6151
R4447 vdd.n2860 vdd.n892 10.6151
R4448 vdd.n2870 vdd.n892 10.6151
R4449 vdd.n2871 vdd.n2870 10.6151
R4450 vdd.n2872 vdd.n2871 10.6151
R4451 vdd.n2872 vdd.n880 10.6151
R4452 vdd.n2882 vdd.n880 10.6151
R4453 vdd.n2883 vdd.n2882 10.6151
R4454 vdd.n2884 vdd.n2883 10.6151
R4455 vdd.n2884 vdd.n868 10.6151
R4456 vdd.n2894 vdd.n868 10.6151
R4457 vdd.n2895 vdd.n2894 10.6151
R4458 vdd.n2896 vdd.n2895 10.6151
R4459 vdd.n2896 vdd.n857 10.6151
R4460 vdd.n2906 vdd.n857 10.6151
R4461 vdd.n2907 vdd.n2906 10.6151
R4462 vdd.n2908 vdd.n2907 10.6151
R4463 vdd.n2908 vdd.n844 10.6151
R4464 vdd.n2918 vdd.n844 10.6151
R4465 vdd.n2919 vdd.n2918 10.6151
R4466 vdd.n2921 vdd.n832 10.6151
R4467 vdd.n2931 vdd.n832 10.6151
R4468 vdd.n2932 vdd.n2931 10.6151
R4469 vdd.n2933 vdd.n2932 10.6151
R4470 vdd.n2933 vdd.n820 10.6151
R4471 vdd.n2943 vdd.n820 10.6151
R4472 vdd.n2944 vdd.n2943 10.6151
R4473 vdd.n2990 vdd.n2944 10.6151
R4474 vdd.n2990 vdd.n2989 10.6151
R4475 vdd.n2989 vdd.n2988 10.6151
R4476 vdd.n2988 vdd.n2987 10.6151
R4477 vdd.n2987 vdd.n2985 10.6151
R4478 vdd.n2339 vdd.n2338 10.6151
R4479 vdd.n2339 vdd.n1040 10.6151
R4480 vdd.n2349 vdd.n1040 10.6151
R4481 vdd.n2350 vdd.n2349 10.6151
R4482 vdd.n2351 vdd.n2350 10.6151
R4483 vdd.n2351 vdd.n1028 10.6151
R4484 vdd.n2361 vdd.n1028 10.6151
R4485 vdd.n2362 vdd.n2361 10.6151
R4486 vdd.n2363 vdd.n2362 10.6151
R4487 vdd.n2363 vdd.n1015 10.6151
R4488 vdd.n2373 vdd.n1015 10.6151
R4489 vdd.n2374 vdd.n2373 10.6151
R4490 vdd.n2376 vdd.n1003 10.6151
R4491 vdd.n2386 vdd.n1003 10.6151
R4492 vdd.n2387 vdd.n2386 10.6151
R4493 vdd.n2388 vdd.n2387 10.6151
R4494 vdd.n2388 vdd.n991 10.6151
R4495 vdd.n2398 vdd.n991 10.6151
R4496 vdd.n2399 vdd.n2398 10.6151
R4497 vdd.n2400 vdd.n2399 10.6151
R4498 vdd.n2400 vdd.n980 10.6151
R4499 vdd.n2410 vdd.n980 10.6151
R4500 vdd.n2411 vdd.n2410 10.6151
R4501 vdd.n2412 vdd.n2411 10.6151
R4502 vdd.n2412 vdd.n968 10.6151
R4503 vdd.n2422 vdd.n968 10.6151
R4504 vdd.n2423 vdd.n2422 10.6151
R4505 vdd.n2426 vdd.n2423 10.6151
R4506 vdd.n2426 vdd.n2425 10.6151
R4507 vdd.n2425 vdd.n2424 10.6151
R4508 vdd.n2424 vdd.n951 10.6151
R4509 vdd.n2508 vdd.n951 10.6151
R4510 vdd.n2507 vdd.n2506 10.6151
R4511 vdd.n2506 vdd.n2503 10.6151
R4512 vdd.n2503 vdd.n2502 10.6151
R4513 vdd.n2502 vdd.n2499 10.6151
R4514 vdd.n2499 vdd.n2498 10.6151
R4515 vdd.n2498 vdd.n2495 10.6151
R4516 vdd.n2495 vdd.n2494 10.6151
R4517 vdd.n2494 vdd.n2491 10.6151
R4518 vdd.n2491 vdd.n2490 10.6151
R4519 vdd.n2490 vdd.n2487 10.6151
R4520 vdd.n2487 vdd.n2486 10.6151
R4521 vdd.n2486 vdd.n2483 10.6151
R4522 vdd.n2483 vdd.n2482 10.6151
R4523 vdd.n2482 vdd.n2479 10.6151
R4524 vdd.n2479 vdd.n2478 10.6151
R4525 vdd.n2478 vdd.n2475 10.6151
R4526 vdd.n2475 vdd.n2474 10.6151
R4527 vdd.n2474 vdd.n2471 10.6151
R4528 vdd.n2471 vdd.n2470 10.6151
R4529 vdd.n2470 vdd.n2467 10.6151
R4530 vdd.n2467 vdd.n2466 10.6151
R4531 vdd.n2466 vdd.n2463 10.6151
R4532 vdd.n2463 vdd.n2462 10.6151
R4533 vdd.n2462 vdd.n2459 10.6151
R4534 vdd.n2459 vdd.n2458 10.6151
R4535 vdd.n2458 vdd.n2455 10.6151
R4536 vdd.n2455 vdd.n2454 10.6151
R4537 vdd.n2454 vdd.n2451 10.6151
R4538 vdd.n2451 vdd.n2450 10.6151
R4539 vdd.n2450 vdd.n2447 10.6151
R4540 vdd.n2447 vdd.n2446 10.6151
R4541 vdd.n2443 vdd.n2442 10.6151
R4542 vdd.n2442 vdd.n2440 10.6151
R4543 vdd.n1359 vdd.n1357 10.6151
R4544 vdd.n1357 vdd.n1356 10.6151
R4545 vdd.n1356 vdd.n1354 10.6151
R4546 vdd.n1354 vdd.n1353 10.6151
R4547 vdd.n1353 vdd.n1351 10.6151
R4548 vdd.n1351 vdd.n1350 10.6151
R4549 vdd.n1350 vdd.n1348 10.6151
R4550 vdd.n1348 vdd.n1347 10.6151
R4551 vdd.n1347 vdd.n1345 10.6151
R4552 vdd.n1345 vdd.n1344 10.6151
R4553 vdd.n1344 vdd.n1342 10.6151
R4554 vdd.n1342 vdd.n1341 10.6151
R4555 vdd.n1341 vdd.n1339 10.6151
R4556 vdd.n1339 vdd.n1338 10.6151
R4557 vdd.n1338 vdd.n1336 10.6151
R4558 vdd.n1336 vdd.n1335 10.6151
R4559 vdd.n1335 vdd.n1333 10.6151
R4560 vdd.n1333 vdd.n1332 10.6151
R4561 vdd.n1332 vdd.n1243 10.6151
R4562 vdd.n1243 vdd.n1242 10.6151
R4563 vdd.n1242 vdd.n1240 10.6151
R4564 vdd.n1240 vdd.n1239 10.6151
R4565 vdd.n1239 vdd.n1237 10.6151
R4566 vdd.n1237 vdd.n1236 10.6151
R4567 vdd.n1236 vdd.n1234 10.6151
R4568 vdd.n1234 vdd.n1233 10.6151
R4569 vdd.n1233 vdd.n1231 10.6151
R4570 vdd.n1231 vdd.n1230 10.6151
R4571 vdd.n1230 vdd.n1228 10.6151
R4572 vdd.n1228 vdd.n1227 10.6151
R4573 vdd.n1227 vdd.n955 10.6151
R4574 vdd.n2438 vdd.n955 10.6151
R4575 vdd.n2439 vdd.n2438 10.6151
R4576 vdd.n2337 vdd.n1052 10.6151
R4577 vdd.n1194 vdd.n1052 10.6151
R4578 vdd.n1195 vdd.n1194 10.6151
R4579 vdd.n1198 vdd.n1195 10.6151
R4580 vdd.n1199 vdd.n1198 10.6151
R4581 vdd.n1202 vdd.n1199 10.6151
R4582 vdd.n1203 vdd.n1202 10.6151
R4583 vdd.n1206 vdd.n1203 10.6151
R4584 vdd.n1207 vdd.n1206 10.6151
R4585 vdd.n1210 vdd.n1207 10.6151
R4586 vdd.n1211 vdd.n1210 10.6151
R4587 vdd.n1214 vdd.n1211 10.6151
R4588 vdd.n1215 vdd.n1214 10.6151
R4589 vdd.n1218 vdd.n1215 10.6151
R4590 vdd.n1219 vdd.n1218 10.6151
R4591 vdd.n1222 vdd.n1219 10.6151
R4592 vdd.n1393 vdd.n1222 10.6151
R4593 vdd.n1393 vdd.n1392 10.6151
R4594 vdd.n1392 vdd.n1390 10.6151
R4595 vdd.n1390 vdd.n1387 10.6151
R4596 vdd.n1387 vdd.n1386 10.6151
R4597 vdd.n1386 vdd.n1383 10.6151
R4598 vdd.n1383 vdd.n1382 10.6151
R4599 vdd.n1382 vdd.n1379 10.6151
R4600 vdd.n1379 vdd.n1378 10.6151
R4601 vdd.n1378 vdd.n1375 10.6151
R4602 vdd.n1375 vdd.n1374 10.6151
R4603 vdd.n1374 vdd.n1371 10.6151
R4604 vdd.n1371 vdd.n1370 10.6151
R4605 vdd.n1370 vdd.n1367 10.6151
R4606 vdd.n1367 vdd.n1366 10.6151
R4607 vdd.n1363 vdd.n1362 10.6151
R4608 vdd.n1362 vdd.n1360 10.6151
R4609 vdd.t15 vdd.n2138 10.5435
R4610 vdd.n636 vdd.t102 10.5435
R4611 vdd.n304 vdd.n286 10.4732
R4612 vdd.n249 vdd.n231 10.4732
R4613 vdd.n206 vdd.n188 10.4732
R4614 vdd.n151 vdd.n133 10.4732
R4615 vdd.n109 vdd.n91 10.4732
R4616 vdd.n54 vdd.n36 10.4732
R4617 vdd.n2035 vdd.n2017 10.4732
R4618 vdd.n2090 vdd.n2072 10.4732
R4619 vdd.n1937 vdd.n1919 10.4732
R4620 vdd.n1992 vdd.n1974 10.4732
R4621 vdd.n1840 vdd.n1822 10.4732
R4622 vdd.n1895 vdd.n1877 10.4732
R4623 vdd.n2122 vdd.t152 10.3167
R4624 vdd.n3297 vdd.t11 10.3167
R4625 vdd.t148 vdd.n1466 10.09
R4626 vdd.n2174 vdd.t30 10.09
R4627 vdd.n3245 vdd.t26 10.09
R4628 vdd.n3378 vdd.t98 10.09
R4629 vdd.n1786 vdd.t123 9.86327
R4630 vdd.n3369 vdd.t0 9.86327
R4631 vdd.n2299 vdd.n2298 9.78206
R4632 vdd.n3035 vdd.n3034 9.78206
R4633 vdd.n3102 vdd.n3101 9.78206
R4634 vdd.n2191 vdd.n1393 9.78206
R4635 vdd.n303 vdd.n288 9.69747
R4636 vdd.n248 vdd.n233 9.69747
R4637 vdd.n205 vdd.n190 9.69747
R4638 vdd.n150 vdd.n135 9.69747
R4639 vdd.n108 vdd.n93 9.69747
R4640 vdd.n53 vdd.n38 9.69747
R4641 vdd.n2034 vdd.n2019 9.69747
R4642 vdd.n2089 vdd.n2074 9.69747
R4643 vdd.n1936 vdd.n1921 9.69747
R4644 vdd.n1991 vdd.n1976 9.69747
R4645 vdd.n1839 vdd.n1824 9.69747
R4646 vdd.n1894 vdd.n1879 9.69747
R4647 vdd.t108 vdd.n1760 9.63654
R4648 vdd.n3328 vdd.t150 9.63654
R4649 vdd.n319 vdd.n318 9.45567
R4650 vdd.n264 vdd.n263 9.45567
R4651 vdd.n221 vdd.n220 9.45567
R4652 vdd.n166 vdd.n165 9.45567
R4653 vdd.n124 vdd.n123 9.45567
R4654 vdd.n69 vdd.n68 9.45567
R4655 vdd.n2050 vdd.n2049 9.45567
R4656 vdd.n2105 vdd.n2104 9.45567
R4657 vdd.n1952 vdd.n1951 9.45567
R4658 vdd.n2007 vdd.n2006 9.45567
R4659 vdd.n1855 vdd.n1854 9.45567
R4660 vdd.n1910 vdd.n1909 9.45567
R4661 vdd.n2261 vdd.n1120 9.3005
R4662 vdd.n2260 vdd.n2259 9.3005
R4663 vdd.n1126 vdd.n1125 9.3005
R4664 vdd.n2254 vdd.n1130 9.3005
R4665 vdd.n2253 vdd.n1131 9.3005
R4666 vdd.n2252 vdd.n1132 9.3005
R4667 vdd.n1136 vdd.n1133 9.3005
R4668 vdd.n2247 vdd.n1137 9.3005
R4669 vdd.n2246 vdd.n1138 9.3005
R4670 vdd.n2245 vdd.n1139 9.3005
R4671 vdd.n1143 vdd.n1140 9.3005
R4672 vdd.n2240 vdd.n1144 9.3005
R4673 vdd.n2239 vdd.n1145 9.3005
R4674 vdd.n2238 vdd.n1146 9.3005
R4675 vdd.n1150 vdd.n1147 9.3005
R4676 vdd.n2233 vdd.n1151 9.3005
R4677 vdd.n2232 vdd.n1152 9.3005
R4678 vdd.n2231 vdd.n1153 9.3005
R4679 vdd.n1157 vdd.n1154 9.3005
R4680 vdd.n2226 vdd.n1158 9.3005
R4681 vdd.n2225 vdd.n1159 9.3005
R4682 vdd.n2224 vdd.n2223 9.3005
R4683 vdd.n2222 vdd.n1160 9.3005
R4684 vdd.n2221 vdd.n2220 9.3005
R4685 vdd.n1166 vdd.n1165 9.3005
R4686 vdd.n2215 vdd.n1170 9.3005
R4687 vdd.n2214 vdd.n1171 9.3005
R4688 vdd.n2213 vdd.n1172 9.3005
R4689 vdd.n1176 vdd.n1173 9.3005
R4690 vdd.n2208 vdd.n1177 9.3005
R4691 vdd.n2207 vdd.n1178 9.3005
R4692 vdd.n2206 vdd.n1179 9.3005
R4693 vdd.n1183 vdd.n1180 9.3005
R4694 vdd.n2201 vdd.n1184 9.3005
R4695 vdd.n2200 vdd.n1185 9.3005
R4696 vdd.n2199 vdd.n1186 9.3005
R4697 vdd.n1190 vdd.n1187 9.3005
R4698 vdd.n2194 vdd.n1191 9.3005
R4699 vdd.n2263 vdd.n2262 9.3005
R4700 vdd.n2285 vdd.n1091 9.3005
R4701 vdd.n2284 vdd.n1099 9.3005
R4702 vdd.n1103 vdd.n1100 9.3005
R4703 vdd.n2279 vdd.n1104 9.3005
R4704 vdd.n2278 vdd.n1105 9.3005
R4705 vdd.n2277 vdd.n1106 9.3005
R4706 vdd.n1110 vdd.n1107 9.3005
R4707 vdd.n2272 vdd.n1111 9.3005
R4708 vdd.n2271 vdd.n1112 9.3005
R4709 vdd.n2270 vdd.n1113 9.3005
R4710 vdd.n1117 vdd.n1114 9.3005
R4711 vdd.n2265 vdd.n1118 9.3005
R4712 vdd.n2264 vdd.n1119 9.3005
R4713 vdd.n2297 vdd.n2296 9.3005
R4714 vdd.n1095 vdd.n1094 9.3005
R4715 vdd.n2110 vdd.n1456 9.3005
R4716 vdd.n2112 vdd.n2111 9.3005
R4717 vdd.n1447 vdd.n1446 9.3005
R4718 vdd.n2125 vdd.n2124 9.3005
R4719 vdd.n2126 vdd.n1445 9.3005
R4720 vdd.n2128 vdd.n2127 9.3005
R4721 vdd.n1435 vdd.n1434 9.3005
R4722 vdd.n2142 vdd.n2141 9.3005
R4723 vdd.n2143 vdd.n1433 9.3005
R4724 vdd.n2145 vdd.n2144 9.3005
R4725 vdd.n1424 vdd.n1423 9.3005
R4726 vdd.n2159 vdd.n2158 9.3005
R4727 vdd.n2160 vdd.n1422 9.3005
R4728 vdd.n2162 vdd.n2161 9.3005
R4729 vdd.n1412 vdd.n1411 9.3005
R4730 vdd.n2177 vdd.n2176 9.3005
R4731 vdd.n2178 vdd.n1410 9.3005
R4732 vdd.n2180 vdd.n2179 9.3005
R4733 vdd.n295 vdd.n294 9.3005
R4734 vdd.n290 vdd.n289 9.3005
R4735 vdd.n301 vdd.n300 9.3005
R4736 vdd.n303 vdd.n302 9.3005
R4737 vdd.n286 vdd.n285 9.3005
R4738 vdd.n309 vdd.n308 9.3005
R4739 vdd.n311 vdd.n310 9.3005
R4740 vdd.n283 vdd.n280 9.3005
R4741 vdd.n318 vdd.n317 9.3005
R4742 vdd.n240 vdd.n239 9.3005
R4743 vdd.n235 vdd.n234 9.3005
R4744 vdd.n246 vdd.n245 9.3005
R4745 vdd.n248 vdd.n247 9.3005
R4746 vdd.n231 vdd.n230 9.3005
R4747 vdd.n254 vdd.n253 9.3005
R4748 vdd.n256 vdd.n255 9.3005
R4749 vdd.n228 vdd.n225 9.3005
R4750 vdd.n263 vdd.n262 9.3005
R4751 vdd.n197 vdd.n196 9.3005
R4752 vdd.n192 vdd.n191 9.3005
R4753 vdd.n203 vdd.n202 9.3005
R4754 vdd.n205 vdd.n204 9.3005
R4755 vdd.n188 vdd.n187 9.3005
R4756 vdd.n211 vdd.n210 9.3005
R4757 vdd.n213 vdd.n212 9.3005
R4758 vdd.n185 vdd.n182 9.3005
R4759 vdd.n220 vdd.n219 9.3005
R4760 vdd.n142 vdd.n141 9.3005
R4761 vdd.n137 vdd.n136 9.3005
R4762 vdd.n148 vdd.n147 9.3005
R4763 vdd.n150 vdd.n149 9.3005
R4764 vdd.n133 vdd.n132 9.3005
R4765 vdd.n156 vdd.n155 9.3005
R4766 vdd.n158 vdd.n157 9.3005
R4767 vdd.n130 vdd.n127 9.3005
R4768 vdd.n165 vdd.n164 9.3005
R4769 vdd.n100 vdd.n99 9.3005
R4770 vdd.n95 vdd.n94 9.3005
R4771 vdd.n106 vdd.n105 9.3005
R4772 vdd.n108 vdd.n107 9.3005
R4773 vdd.n91 vdd.n90 9.3005
R4774 vdd.n114 vdd.n113 9.3005
R4775 vdd.n116 vdd.n115 9.3005
R4776 vdd.n88 vdd.n85 9.3005
R4777 vdd.n123 vdd.n122 9.3005
R4778 vdd.n45 vdd.n44 9.3005
R4779 vdd.n40 vdd.n39 9.3005
R4780 vdd.n51 vdd.n50 9.3005
R4781 vdd.n53 vdd.n52 9.3005
R4782 vdd.n36 vdd.n35 9.3005
R4783 vdd.n59 vdd.n58 9.3005
R4784 vdd.n61 vdd.n60 9.3005
R4785 vdd.n33 vdd.n30 9.3005
R4786 vdd.n68 vdd.n67 9.3005
R4787 vdd.n3151 vdd.n3150 9.3005
R4788 vdd.n3152 vdd.n721 9.3005
R4789 vdd.n720 vdd.n718 9.3005
R4790 vdd.n3158 vdd.n717 9.3005
R4791 vdd.n3159 vdd.n716 9.3005
R4792 vdd.n3160 vdd.n715 9.3005
R4793 vdd.n714 vdd.n712 9.3005
R4794 vdd.n3166 vdd.n711 9.3005
R4795 vdd.n3167 vdd.n710 9.3005
R4796 vdd.n3168 vdd.n709 9.3005
R4797 vdd.n708 vdd.n706 9.3005
R4798 vdd.n3174 vdd.n705 9.3005
R4799 vdd.n3175 vdd.n704 9.3005
R4800 vdd.n3176 vdd.n703 9.3005
R4801 vdd.n702 vdd.n700 9.3005
R4802 vdd.n3182 vdd.n699 9.3005
R4803 vdd.n3183 vdd.n698 9.3005
R4804 vdd.n3184 vdd.n697 9.3005
R4805 vdd.n696 vdd.n694 9.3005
R4806 vdd.n3190 vdd.n693 9.3005
R4807 vdd.n3191 vdd.n692 9.3005
R4808 vdd.n3192 vdd.n691 9.3005
R4809 vdd.n690 vdd.n688 9.3005
R4810 vdd.n3198 vdd.n685 9.3005
R4811 vdd.n3199 vdd.n684 9.3005
R4812 vdd.n3200 vdd.n683 9.3005
R4813 vdd.n682 vdd.n680 9.3005
R4814 vdd.n3206 vdd.n679 9.3005
R4815 vdd.n3207 vdd.n678 9.3005
R4816 vdd.n3208 vdd.n677 9.3005
R4817 vdd.n676 vdd.n674 9.3005
R4818 vdd.n3214 vdd.n673 9.3005
R4819 vdd.n3215 vdd.n672 9.3005
R4820 vdd.n3216 vdd.n671 9.3005
R4821 vdd.n670 vdd.n668 9.3005
R4822 vdd.n3221 vdd.n667 9.3005
R4823 vdd.n3231 vdd.n661 9.3005
R4824 vdd.n3233 vdd.n3232 9.3005
R4825 vdd.n652 vdd.n651 9.3005
R4826 vdd.n3248 vdd.n3247 9.3005
R4827 vdd.n3249 vdd.n650 9.3005
R4828 vdd.n3251 vdd.n3250 9.3005
R4829 vdd.n640 vdd.n639 9.3005
R4830 vdd.n3264 vdd.n3263 9.3005
R4831 vdd.n3265 vdd.n638 9.3005
R4832 vdd.n3267 vdd.n3266 9.3005
R4833 vdd.n628 vdd.n627 9.3005
R4834 vdd.n3281 vdd.n3280 9.3005
R4835 vdd.n3282 vdd.n626 9.3005
R4836 vdd.n3284 vdd.n3283 9.3005
R4837 vdd.n617 vdd.n616 9.3005
R4838 vdd.n3300 vdd.n3299 9.3005
R4839 vdd.n3301 vdd.n615 9.3005
R4840 vdd.n3303 vdd.n3302 9.3005
R4841 vdd.n324 vdd.n322 9.3005
R4842 vdd.n3235 vdd.n3234 9.3005
R4843 vdd.n3382 vdd.n3381 9.3005
R4844 vdd.n325 vdd.n323 9.3005
R4845 vdd.n3375 vdd.n334 9.3005
R4846 vdd.n3374 vdd.n335 9.3005
R4847 vdd.n3373 vdd.n336 9.3005
R4848 vdd.n343 vdd.n337 9.3005
R4849 vdd.n3367 vdd.n344 9.3005
R4850 vdd.n3366 vdd.n345 9.3005
R4851 vdd.n3365 vdd.n346 9.3005
R4852 vdd.n354 vdd.n347 9.3005
R4853 vdd.n3359 vdd.n355 9.3005
R4854 vdd.n3358 vdd.n356 9.3005
R4855 vdd.n3357 vdd.n357 9.3005
R4856 vdd.n365 vdd.n358 9.3005
R4857 vdd.n3351 vdd.n366 9.3005
R4858 vdd.n3350 vdd.n367 9.3005
R4859 vdd.n3349 vdd.n368 9.3005
R4860 vdd.n443 vdd.n369 9.3005
R4861 vdd.n447 vdd.n442 9.3005
R4862 vdd.n451 vdd.n450 9.3005
R4863 vdd.n452 vdd.n441 9.3005
R4864 vdd.n456 vdd.n453 9.3005
R4865 vdd.n457 vdd.n440 9.3005
R4866 vdd.n461 vdd.n460 9.3005
R4867 vdd.n462 vdd.n439 9.3005
R4868 vdd.n466 vdd.n463 9.3005
R4869 vdd.n467 vdd.n438 9.3005
R4870 vdd.n471 vdd.n470 9.3005
R4871 vdd.n472 vdd.n437 9.3005
R4872 vdd.n476 vdd.n473 9.3005
R4873 vdd.n477 vdd.n436 9.3005
R4874 vdd.n481 vdd.n480 9.3005
R4875 vdd.n482 vdd.n435 9.3005
R4876 vdd.n486 vdd.n483 9.3005
R4877 vdd.n487 vdd.n434 9.3005
R4878 vdd.n491 vdd.n490 9.3005
R4879 vdd.n492 vdd.n433 9.3005
R4880 vdd.n496 vdd.n493 9.3005
R4881 vdd.n497 vdd.n430 9.3005
R4882 vdd.n501 vdd.n500 9.3005
R4883 vdd.n502 vdd.n429 9.3005
R4884 vdd.n506 vdd.n503 9.3005
R4885 vdd.n507 vdd.n428 9.3005
R4886 vdd.n511 vdd.n510 9.3005
R4887 vdd.n512 vdd.n427 9.3005
R4888 vdd.n516 vdd.n513 9.3005
R4889 vdd.n517 vdd.n426 9.3005
R4890 vdd.n521 vdd.n520 9.3005
R4891 vdd.n522 vdd.n425 9.3005
R4892 vdd.n526 vdd.n523 9.3005
R4893 vdd.n527 vdd.n424 9.3005
R4894 vdd.n531 vdd.n530 9.3005
R4895 vdd.n532 vdd.n423 9.3005
R4896 vdd.n536 vdd.n533 9.3005
R4897 vdd.n537 vdd.n422 9.3005
R4898 vdd.n541 vdd.n540 9.3005
R4899 vdd.n542 vdd.n421 9.3005
R4900 vdd.n546 vdd.n543 9.3005
R4901 vdd.n547 vdd.n418 9.3005
R4902 vdd.n551 vdd.n550 9.3005
R4903 vdd.n552 vdd.n417 9.3005
R4904 vdd.n556 vdd.n553 9.3005
R4905 vdd.n557 vdd.n416 9.3005
R4906 vdd.n561 vdd.n560 9.3005
R4907 vdd.n562 vdd.n415 9.3005
R4908 vdd.n566 vdd.n563 9.3005
R4909 vdd.n567 vdd.n414 9.3005
R4910 vdd.n571 vdd.n570 9.3005
R4911 vdd.n572 vdd.n413 9.3005
R4912 vdd.n576 vdd.n573 9.3005
R4913 vdd.n577 vdd.n412 9.3005
R4914 vdd.n581 vdd.n580 9.3005
R4915 vdd.n582 vdd.n411 9.3005
R4916 vdd.n586 vdd.n583 9.3005
R4917 vdd.n587 vdd.n410 9.3005
R4918 vdd.n591 vdd.n590 9.3005
R4919 vdd.n592 vdd.n409 9.3005
R4920 vdd.n596 vdd.n593 9.3005
R4921 vdd.n598 vdd.n408 9.3005
R4922 vdd.n600 vdd.n599 9.3005
R4923 vdd.n3342 vdd.n3341 9.3005
R4924 vdd.n446 vdd.n444 9.3005
R4925 vdd.n3241 vdd.n655 9.3005
R4926 vdd.n3243 vdd.n3242 9.3005
R4927 vdd.n646 vdd.n645 9.3005
R4928 vdd.n3256 vdd.n3255 9.3005
R4929 vdd.n3257 vdd.n644 9.3005
R4930 vdd.n3259 vdd.n3258 9.3005
R4931 vdd.n633 vdd.n632 9.3005
R4932 vdd.n3272 vdd.n3271 9.3005
R4933 vdd.n3273 vdd.n631 9.3005
R4934 vdd.n3275 vdd.n3274 9.3005
R4935 vdd.n622 vdd.n621 9.3005
R4936 vdd.n3289 vdd.n3288 9.3005
R4937 vdd.n3290 vdd.n620 9.3005
R4938 vdd.n3295 vdd.n3291 9.3005
R4939 vdd.n3294 vdd.n3293 9.3005
R4940 vdd.n3292 vdd.n610 9.3005
R4941 vdd.n3308 vdd.n611 9.3005
R4942 vdd.n3309 vdd.n609 9.3005
R4943 vdd.n3311 vdd.n3310 9.3005
R4944 vdd.n3312 vdd.n608 9.3005
R4945 vdd.n3315 vdd.n3313 9.3005
R4946 vdd.n3316 vdd.n607 9.3005
R4947 vdd.n3318 vdd.n3317 9.3005
R4948 vdd.n3319 vdd.n606 9.3005
R4949 vdd.n3322 vdd.n3320 9.3005
R4950 vdd.n3323 vdd.n605 9.3005
R4951 vdd.n3325 vdd.n3324 9.3005
R4952 vdd.n3326 vdd.n604 9.3005
R4953 vdd.n3330 vdd.n3327 9.3005
R4954 vdd.n3331 vdd.n603 9.3005
R4955 vdd.n3333 vdd.n3332 9.3005
R4956 vdd.n3334 vdd.n602 9.3005
R4957 vdd.n3337 vdd.n3335 9.3005
R4958 vdd.n3338 vdd.n601 9.3005
R4959 vdd.n3340 vdd.n3339 9.3005
R4960 vdd.n3240 vdd.n3239 9.3005
R4961 vdd.n3104 vdd.n656 9.3005
R4962 vdd.n3109 vdd.n3103 9.3005
R4963 vdd.n3119 vdd.n748 9.3005
R4964 vdd.n3120 vdd.n747 9.3005
R4965 vdd.n746 vdd.n744 9.3005
R4966 vdd.n3126 vdd.n743 9.3005
R4967 vdd.n3127 vdd.n742 9.3005
R4968 vdd.n3128 vdd.n741 9.3005
R4969 vdd.n740 vdd.n738 9.3005
R4970 vdd.n3134 vdd.n737 9.3005
R4971 vdd.n3135 vdd.n736 9.3005
R4972 vdd.n3136 vdd.n735 9.3005
R4973 vdd.n734 vdd.n732 9.3005
R4974 vdd.n3141 vdd.n731 9.3005
R4975 vdd.n3142 vdd.n730 9.3005
R4976 vdd.n726 vdd.n725 9.3005
R4977 vdd.n3148 vdd.n3147 9.3005
R4978 vdd.n3149 vdd.n722 9.3005
R4979 vdd.n2190 vdd.n2189 9.3005
R4980 vdd.n2185 vdd.n1395 9.3005
R4981 vdd.n1742 vdd.n1741 9.3005
R4982 vdd.n1498 vdd.n1497 9.3005
R4983 vdd.n1755 vdd.n1754 9.3005
R4984 vdd.n1756 vdd.n1496 9.3005
R4985 vdd.n1758 vdd.n1757 9.3005
R4986 vdd.n1486 vdd.n1485 9.3005
R4987 vdd.n1772 vdd.n1771 9.3005
R4988 vdd.n1773 vdd.n1484 9.3005
R4989 vdd.n1775 vdd.n1774 9.3005
R4990 vdd.n1476 vdd.n1475 9.3005
R4991 vdd.n1789 vdd.n1788 9.3005
R4992 vdd.n1790 vdd.n1474 9.3005
R4993 vdd.n1792 vdd.n1791 9.3005
R4994 vdd.n1463 vdd.n1462 9.3005
R4995 vdd.n1805 vdd.n1804 9.3005
R4996 vdd.n1806 vdd.n1461 9.3005
R4997 vdd.n1808 vdd.n1807 9.3005
R4998 vdd.n1452 vdd.n1451 9.3005
R4999 vdd.n2117 vdd.n2116 9.3005
R5000 vdd.n2118 vdd.n1450 9.3005
R5001 vdd.n2120 vdd.n2119 9.3005
R5002 vdd.n1441 vdd.n1440 9.3005
R5003 vdd.n2133 vdd.n2132 9.3005
R5004 vdd.n2134 vdd.n1439 9.3005
R5005 vdd.n2136 vdd.n2135 9.3005
R5006 vdd.n1429 vdd.n1428 9.3005
R5007 vdd.n2150 vdd.n2149 9.3005
R5008 vdd.n2151 vdd.n1427 9.3005
R5009 vdd.n2153 vdd.n2152 9.3005
R5010 vdd.n1419 vdd.n1418 9.3005
R5011 vdd.n2167 vdd.n2166 9.3005
R5012 vdd.n2168 vdd.n1416 9.3005
R5013 vdd.n2172 vdd.n2171 9.3005
R5014 vdd.n2170 vdd.n1417 9.3005
R5015 vdd.n2169 vdd.n1406 9.3005
R5016 vdd.n1740 vdd.n1508 9.3005
R5017 vdd.n1633 vdd.n1509 9.3005
R5018 vdd.n1635 vdd.n1634 9.3005
R5019 vdd.n1636 vdd.n1628 9.3005
R5020 vdd.n1638 vdd.n1637 9.3005
R5021 vdd.n1639 vdd.n1627 9.3005
R5022 vdd.n1641 vdd.n1640 9.3005
R5023 vdd.n1642 vdd.n1622 9.3005
R5024 vdd.n1644 vdd.n1643 9.3005
R5025 vdd.n1645 vdd.n1621 9.3005
R5026 vdd.n1647 vdd.n1646 9.3005
R5027 vdd.n1648 vdd.n1616 9.3005
R5028 vdd.n1650 vdd.n1649 9.3005
R5029 vdd.n1651 vdd.n1615 9.3005
R5030 vdd.n1653 vdd.n1652 9.3005
R5031 vdd.n1654 vdd.n1610 9.3005
R5032 vdd.n1656 vdd.n1655 9.3005
R5033 vdd.n1657 vdd.n1609 9.3005
R5034 vdd.n1659 vdd.n1658 9.3005
R5035 vdd.n1660 vdd.n1604 9.3005
R5036 vdd.n1662 vdd.n1661 9.3005
R5037 vdd.n1663 vdd.n1603 9.3005
R5038 vdd.n1668 vdd.n1664 9.3005
R5039 vdd.n1669 vdd.n1599 9.3005
R5040 vdd.n1671 vdd.n1670 9.3005
R5041 vdd.n1672 vdd.n1598 9.3005
R5042 vdd.n1674 vdd.n1673 9.3005
R5043 vdd.n1675 vdd.n1593 9.3005
R5044 vdd.n1677 vdd.n1676 9.3005
R5045 vdd.n1678 vdd.n1592 9.3005
R5046 vdd.n1680 vdd.n1679 9.3005
R5047 vdd.n1681 vdd.n1587 9.3005
R5048 vdd.n1683 vdd.n1682 9.3005
R5049 vdd.n1684 vdd.n1586 9.3005
R5050 vdd.n1686 vdd.n1685 9.3005
R5051 vdd.n1687 vdd.n1581 9.3005
R5052 vdd.n1689 vdd.n1688 9.3005
R5053 vdd.n1690 vdd.n1580 9.3005
R5054 vdd.n1692 vdd.n1691 9.3005
R5055 vdd.n1693 vdd.n1575 9.3005
R5056 vdd.n1695 vdd.n1694 9.3005
R5057 vdd.n1696 vdd.n1574 9.3005
R5058 vdd.n1698 vdd.n1697 9.3005
R5059 vdd.n1699 vdd.n1571 9.3005
R5060 vdd.n1705 vdd.n1704 9.3005
R5061 vdd.n1706 vdd.n1570 9.3005
R5062 vdd.n1708 vdd.n1707 9.3005
R5063 vdd.n1709 vdd.n1565 9.3005
R5064 vdd.n1711 vdd.n1710 9.3005
R5065 vdd.n1712 vdd.n1564 9.3005
R5066 vdd.n1714 vdd.n1713 9.3005
R5067 vdd.n1715 vdd.n1559 9.3005
R5068 vdd.n1717 vdd.n1716 9.3005
R5069 vdd.n1718 vdd.n1558 9.3005
R5070 vdd.n1720 vdd.n1719 9.3005
R5071 vdd.n1721 vdd.n1553 9.3005
R5072 vdd.n1723 vdd.n1722 9.3005
R5073 vdd.n1724 vdd.n1552 9.3005
R5074 vdd.n1726 vdd.n1725 9.3005
R5075 vdd.n1727 vdd.n1548 9.3005
R5076 vdd.n1729 vdd.n1728 9.3005
R5077 vdd.n1730 vdd.n1547 9.3005
R5078 vdd.n1732 vdd.n1731 9.3005
R5079 vdd.n1733 vdd.n1546 9.3005
R5080 vdd.n1739 vdd.n1738 9.3005
R5081 vdd.n1747 vdd.n1746 9.3005
R5082 vdd.n1748 vdd.n1502 9.3005
R5083 vdd.n1750 vdd.n1749 9.3005
R5084 vdd.n1492 vdd.n1491 9.3005
R5085 vdd.n1764 vdd.n1763 9.3005
R5086 vdd.n1765 vdd.n1490 9.3005
R5087 vdd.n1767 vdd.n1766 9.3005
R5088 vdd.n1481 vdd.n1480 9.3005
R5089 vdd.n1781 vdd.n1780 9.3005
R5090 vdd.n1782 vdd.n1479 9.3005
R5091 vdd.n1784 vdd.n1783 9.3005
R5092 vdd.n1470 vdd.n1469 9.3005
R5093 vdd.n1797 vdd.n1796 9.3005
R5094 vdd.n1798 vdd.n1468 9.3005
R5095 vdd.n1800 vdd.n1799 9.3005
R5096 vdd.n1458 vdd.n1457 9.3005
R5097 vdd.n1814 vdd.n1813 9.3005
R5098 vdd.n1504 vdd.n1503 9.3005
R5099 vdd.n2026 vdd.n2025 9.3005
R5100 vdd.n2021 vdd.n2020 9.3005
R5101 vdd.n2032 vdd.n2031 9.3005
R5102 vdd.n2034 vdd.n2033 9.3005
R5103 vdd.n2017 vdd.n2016 9.3005
R5104 vdd.n2040 vdd.n2039 9.3005
R5105 vdd.n2042 vdd.n2041 9.3005
R5106 vdd.n2014 vdd.n2011 9.3005
R5107 vdd.n2049 vdd.n2048 9.3005
R5108 vdd.n2081 vdd.n2080 9.3005
R5109 vdd.n2076 vdd.n2075 9.3005
R5110 vdd.n2087 vdd.n2086 9.3005
R5111 vdd.n2089 vdd.n2088 9.3005
R5112 vdd.n2072 vdd.n2071 9.3005
R5113 vdd.n2095 vdd.n2094 9.3005
R5114 vdd.n2097 vdd.n2096 9.3005
R5115 vdd.n2069 vdd.n2066 9.3005
R5116 vdd.n2104 vdd.n2103 9.3005
R5117 vdd.n1928 vdd.n1927 9.3005
R5118 vdd.n1923 vdd.n1922 9.3005
R5119 vdd.n1934 vdd.n1933 9.3005
R5120 vdd.n1936 vdd.n1935 9.3005
R5121 vdd.n1919 vdd.n1918 9.3005
R5122 vdd.n1942 vdd.n1941 9.3005
R5123 vdd.n1944 vdd.n1943 9.3005
R5124 vdd.n1916 vdd.n1913 9.3005
R5125 vdd.n1951 vdd.n1950 9.3005
R5126 vdd.n1983 vdd.n1982 9.3005
R5127 vdd.n1978 vdd.n1977 9.3005
R5128 vdd.n1989 vdd.n1988 9.3005
R5129 vdd.n1991 vdd.n1990 9.3005
R5130 vdd.n1974 vdd.n1973 9.3005
R5131 vdd.n1997 vdd.n1996 9.3005
R5132 vdd.n1999 vdd.n1998 9.3005
R5133 vdd.n1971 vdd.n1968 9.3005
R5134 vdd.n2006 vdd.n2005 9.3005
R5135 vdd.n1831 vdd.n1830 9.3005
R5136 vdd.n1826 vdd.n1825 9.3005
R5137 vdd.n1837 vdd.n1836 9.3005
R5138 vdd.n1839 vdd.n1838 9.3005
R5139 vdd.n1822 vdd.n1821 9.3005
R5140 vdd.n1845 vdd.n1844 9.3005
R5141 vdd.n1847 vdd.n1846 9.3005
R5142 vdd.n1819 vdd.n1816 9.3005
R5143 vdd.n1854 vdd.n1853 9.3005
R5144 vdd.n1886 vdd.n1885 9.3005
R5145 vdd.n1881 vdd.n1880 9.3005
R5146 vdd.n1892 vdd.n1891 9.3005
R5147 vdd.n1894 vdd.n1893 9.3005
R5148 vdd.n1877 vdd.n1876 9.3005
R5149 vdd.n1900 vdd.n1899 9.3005
R5150 vdd.n1902 vdd.n1901 9.3005
R5151 vdd.n1874 vdd.n1871 9.3005
R5152 vdd.n1909 vdd.n1908 9.3005
R5153 vdd.n1760 vdd.t110 9.18308
R5154 vdd.n3328 vdd.t9 9.18308
R5155 vdd.n1786 vdd.t138 8.95635
R5156 vdd.t105 vdd.n3369 8.95635
R5157 vdd.n300 vdd.n299 8.92171
R5158 vdd.n245 vdd.n244 8.92171
R5159 vdd.n202 vdd.n201 8.92171
R5160 vdd.n147 vdd.n146 8.92171
R5161 vdd.n105 vdd.n104 8.92171
R5162 vdd.n50 vdd.n49 8.92171
R5163 vdd.n2031 vdd.n2030 8.92171
R5164 vdd.n2086 vdd.n2085 8.92171
R5165 vdd.n1933 vdd.n1932 8.92171
R5166 vdd.n1988 vdd.n1987 8.92171
R5167 vdd.n1836 vdd.n1835 8.92171
R5168 vdd.n1891 vdd.n1890 8.92171
R5169 vdd.n223 vdd.n125 8.81535
R5170 vdd.n2009 vdd.n1911 8.81535
R5171 vdd.n1466 vdd.t130 8.72962
R5172 vdd.t140 vdd.n3378 8.72962
R5173 vdd.n2122 vdd.t13 8.50289
R5174 vdd.n3297 vdd.t93 8.50289
R5175 vdd.n28 vdd.n14 8.42249
R5176 vdd.n2138 vdd.t6 8.27616
R5177 vdd.t136 vdd.n636 8.27616
R5178 vdd.n3384 vdd.n3383 8.16225
R5179 vdd.n2109 vdd.n2108 8.16225
R5180 vdd.n296 vdd.n290 8.14595
R5181 vdd.n241 vdd.n235 8.14595
R5182 vdd.n198 vdd.n192 8.14595
R5183 vdd.n143 vdd.n137 8.14595
R5184 vdd.n101 vdd.n95 8.14595
R5185 vdd.n46 vdd.n40 8.14595
R5186 vdd.n2027 vdd.n2021 8.14595
R5187 vdd.n2082 vdd.n2076 8.14595
R5188 vdd.n1929 vdd.n1923 8.14595
R5189 vdd.n1984 vdd.n1978 8.14595
R5190 vdd.n1832 vdd.n1826 8.14595
R5191 vdd.n1887 vdd.n1881 8.14595
R5192 vdd.t47 vdd.n1500 7.8227
R5193 vdd.t51 vdd.n363 7.8227
R5194 vdd.n2341 vdd.n1047 7.70933
R5195 vdd.n2341 vdd.n1050 7.70933
R5196 vdd.n2347 vdd.n1036 7.70933
R5197 vdd.n2353 vdd.n1036 7.70933
R5198 vdd.n2353 vdd.n1030 7.70933
R5199 vdd.n2359 vdd.n1030 7.70933
R5200 vdd.n2365 vdd.n1023 7.70933
R5201 vdd.n2365 vdd.n1026 7.70933
R5202 vdd.n2371 vdd.n1019 7.70933
R5203 vdd.n2378 vdd.n1005 7.70933
R5204 vdd.n2384 vdd.n1005 7.70933
R5205 vdd.n2390 vdd.n999 7.70933
R5206 vdd.n2396 vdd.n995 7.70933
R5207 vdd.n2402 vdd.n989 7.70933
R5208 vdd.n2414 vdd.n976 7.70933
R5209 vdd.n2420 vdd.n970 7.70933
R5210 vdd.n2420 vdd.n963 7.70933
R5211 vdd.n2428 vdd.n963 7.70933
R5212 vdd.n2510 vdd.n947 7.70933
R5213 vdd.n2862 vdd.n899 7.70933
R5214 vdd.n2874 vdd.n888 7.70933
R5215 vdd.n2874 vdd.n882 7.70933
R5216 vdd.n2880 vdd.n882 7.70933
R5217 vdd.n2886 vdd.n876 7.70933
R5218 vdd.n2892 vdd.n872 7.70933
R5219 vdd.n2898 vdd.n866 7.70933
R5220 vdd.n2910 vdd.n853 7.70933
R5221 vdd.n2916 vdd.n846 7.70933
R5222 vdd.n2916 vdd.n849 7.70933
R5223 vdd.n2923 vdd.n841 7.70933
R5224 vdd.n2929 vdd.n828 7.70933
R5225 vdd.n2935 vdd.n828 7.70933
R5226 vdd.n2941 vdd.n822 7.70933
R5227 vdd.n2941 vdd.n814 7.70933
R5228 vdd.n2992 vdd.n814 7.70933
R5229 vdd.n2992 vdd.n817 7.70933
R5230 vdd.n2998 vdd.n774 7.70933
R5231 vdd.n3068 vdd.n774 7.70933
R5232 vdd.n2921 vdd.n2920 7.49318
R5233 vdd.n2375 vdd.n2374 7.49318
R5234 vdd.n295 vdd.n292 7.3702
R5235 vdd.n240 vdd.n237 7.3702
R5236 vdd.n197 vdd.n194 7.3702
R5237 vdd.n142 vdd.n139 7.3702
R5238 vdd.n100 vdd.n97 7.3702
R5239 vdd.n45 vdd.n42 7.3702
R5240 vdd.n2026 vdd.n2023 7.3702
R5241 vdd.n2081 vdd.n2078 7.3702
R5242 vdd.n1928 vdd.n1925 7.3702
R5243 vdd.n1983 vdd.n1980 7.3702
R5244 vdd.n1831 vdd.n1828 7.3702
R5245 vdd.n1886 vdd.n1883 7.3702
R5246 vdd.n2359 vdd.t203 7.36923
R5247 vdd.t226 vdd.n822 7.36923
R5248 vdd.n2435 vdd.t233 7.25587
R5249 vdd.n2779 vdd.t222 7.25587
R5250 vdd.n1669 vdd.n1668 6.98232
R5251 vdd.n2225 vdd.n2224 6.98232
R5252 vdd.n547 vdd.n546 6.98232
R5253 vdd.n3152 vdd.n3151 6.98232
R5254 vdd.n2156 vdd.t188 6.91577
R5255 vdd.n3261 vdd.t2 6.91577
R5256 vdd.t146 vdd.n1437 6.68904
R5257 vdd.n3277 vdd.t100 6.68904
R5258 vdd.n2114 vdd.t172 6.46231
R5259 vdd.n3305 vdd.t96 6.46231
R5260 vdd.n3384 vdd.n321 6.32949
R5261 vdd.n2108 vdd.n2107 6.32949
R5262 vdd.t4 vdd.n1465 6.23558
R5263 vdd.t183 vdd.n332 6.23558
R5264 vdd.n1778 vdd.t133 6.00885
R5265 vdd.n3363 vdd.t126 6.00885
R5266 vdd.t194 vdd.n976 5.89549
R5267 vdd.n2886 vdd.t231 5.89549
R5268 vdd.n296 vdd.n295 5.81868
R5269 vdd.n241 vdd.n240 5.81868
R5270 vdd.n198 vdd.n197 5.81868
R5271 vdd.n143 vdd.n142 5.81868
R5272 vdd.n101 vdd.n100 5.81868
R5273 vdd.n46 vdd.n45 5.81868
R5274 vdd.n2027 vdd.n2026 5.81868
R5275 vdd.n2082 vdd.n2081 5.81868
R5276 vdd.n1929 vdd.n1928 5.81868
R5277 vdd.n1984 vdd.n1983 5.81868
R5278 vdd.n1832 vdd.n1831 5.81868
R5279 vdd.n1887 vdd.n1886 5.81868
R5280 vdd.n2518 vdd.n2517 5.77611
R5281 vdd.n1274 vdd.n1273 5.77611
R5282 vdd.n2791 vdd.n2790 5.77611
R5283 vdd.n3007 vdd.n806 5.77611
R5284 vdd.n3073 vdd.n770 5.77611
R5285 vdd.n2685 vdd.n2623 5.77611
R5286 vdd.n2443 vdd.n954 5.77611
R5287 vdd.n1363 vdd.n1226 5.77611
R5288 vdd.n1738 vdd.n1512 5.62474
R5289 vdd.n2188 vdd.n2185 5.62474
R5290 vdd.n3342 vdd.n407 5.62474
R5291 vdd.n3107 vdd.n3104 5.62474
R5292 vdd.t206 vdd.n999 5.55539
R5293 vdd.n2390 vdd.t237 5.55539
R5294 vdd.t227 vdd.n853 5.55539
R5295 vdd.n2910 vdd.t211 5.55539
R5296 vdd.n1019 vdd.t72 5.44203
R5297 vdd.n2923 vdd.t40 5.44203
R5298 vdd.n1488 vdd.t133 5.32866
R5299 vdd.n2347 vdd.t22 5.32866
R5300 vdd.n1309 vdd.t64 5.32866
R5301 vdd.n2868 vdd.t68 5.32866
R5302 vdd.n817 vdd.t18 5.32866
R5303 vdd.t126 vdd.n3362 5.32866
R5304 vdd.n1794 vdd.t4 5.10193
R5305 vdd.n3371 vdd.t183 5.10193
R5306 vdd.n299 vdd.n290 5.04292
R5307 vdd.n244 vdd.n235 5.04292
R5308 vdd.n201 vdd.n192 5.04292
R5309 vdd.n146 vdd.n137 5.04292
R5310 vdd.n104 vdd.n95 5.04292
R5311 vdd.n49 vdd.n40 5.04292
R5312 vdd.n2030 vdd.n2021 5.04292
R5313 vdd.n2085 vdd.n2076 5.04292
R5314 vdd.n1932 vdd.n1923 5.04292
R5315 vdd.n1987 vdd.n1978 5.04292
R5316 vdd.n1835 vdd.n1826 5.04292
R5317 vdd.n1890 vdd.n1881 5.04292
R5318 vdd.n2396 vdd.t229 4.98857
R5319 vdd.n866 vdd.t207 4.98857
R5320 vdd.n1810 vdd.t172 4.8752
R5321 vdd.t202 vdd.t212 4.8752
R5322 vdd.t193 vdd.t224 4.8752
R5323 vdd.t215 vdd.t196 4.8752
R5324 vdd.t238 vdd.t192 4.8752
R5325 vdd.t96 vdd.n328 4.8752
R5326 vdd.n2519 vdd.n2518 4.83952
R5327 vdd.n1273 vdd.n1272 4.83952
R5328 vdd.n2792 vdd.n2791 4.83952
R5329 vdd.n806 vdd.n801 4.83952
R5330 vdd.n770 vdd.n765 4.83952
R5331 vdd.n2682 vdd.n2623 4.83952
R5332 vdd.n2446 vdd.n954 4.83952
R5333 vdd.n1366 vdd.n1226 4.83952
R5334 vdd.n2193 vdd.n2192 4.74817
R5335 vdd.n1399 vdd.n1394 4.74817
R5336 vdd.n1096 vdd.n1093 4.74817
R5337 vdd.n2286 vdd.n1092 4.74817
R5338 vdd.n2291 vdd.n1093 4.74817
R5339 vdd.n2290 vdd.n1092 4.74817
R5340 vdd.n664 vdd.n662 4.74817
R5341 vdd.n3222 vdd.n665 4.74817
R5342 vdd.n3225 vdd.n665 4.74817
R5343 vdd.n3226 vdd.n664 4.74817
R5344 vdd.n3114 vdd.n749 4.74817
R5345 vdd.n3110 vdd.n751 4.74817
R5346 vdd.n3113 vdd.n751 4.74817
R5347 vdd.n3118 vdd.n749 4.74817
R5348 vdd.n2192 vdd.n1192 4.74817
R5349 vdd.n1396 vdd.n1394 4.74817
R5350 vdd.n321 vdd.n320 4.7074
R5351 vdd.n223 vdd.n222 4.7074
R5352 vdd.n2107 vdd.n2106 4.7074
R5353 vdd.n2009 vdd.n2008 4.7074
R5354 vdd.n2130 vdd.t146 4.64847
R5355 vdd.n2371 vdd.t219 4.64847
R5356 vdd.n989 vdd.t214 4.64847
R5357 vdd.n2892 vdd.t228 4.64847
R5358 vdd.n841 vdd.t199 4.64847
R5359 vdd.n3286 vdd.t100 4.64847
R5360 vdd.n1431 vdd.t188 4.42174
R5361 vdd.t2 vdd.n635 4.42174
R5362 vdd.n300 vdd.n288 4.26717
R5363 vdd.n245 vdd.n233 4.26717
R5364 vdd.n202 vdd.n190 4.26717
R5365 vdd.n147 vdd.n135 4.26717
R5366 vdd.n105 vdd.n93 4.26717
R5367 vdd.n50 vdd.n38 4.26717
R5368 vdd.n2031 vdd.n2019 4.26717
R5369 vdd.n2086 vdd.n2074 4.26717
R5370 vdd.n1933 vdd.n1921 4.26717
R5371 vdd.n1988 vdd.n1976 4.26717
R5372 vdd.n1836 vdd.n1824 4.26717
R5373 vdd.n1891 vdd.n1879 4.26717
R5374 vdd.n321 vdd.n223 4.10845
R5375 vdd.n2107 vdd.n2009 4.10845
R5376 vdd.n277 vdd.t127 4.06363
R5377 vdd.n277 vdd.t167 4.06363
R5378 vdd.n275 vdd.t106 4.06363
R5379 vdd.n275 vdd.t104 4.06363
R5380 vdd.n273 vdd.t154 4.06363
R5381 vdd.n273 vdd.t184 4.06363
R5382 vdd.n271 vdd.t135 4.06363
R5383 vdd.n271 vdd.t159 4.06363
R5384 vdd.n269 vdd.t94 4.06363
R5385 vdd.n269 vdd.t112 4.06363
R5386 vdd.n267 vdd.t115 4.06363
R5387 vdd.n267 vdd.t114 4.06363
R5388 vdd.n265 vdd.t3 4.06363
R5389 vdd.n265 vdd.t163 4.06363
R5390 vdd.n179 vdd.t242 4.06363
R5391 vdd.n179 vdd.t160 4.06363
R5392 vdd.n177 vdd.t265 4.06363
R5393 vdd.n177 vdd.t1 4.06363
R5394 vdd.n175 vdd.t116 4.06363
R5395 vdd.n175 vdd.t255 4.06363
R5396 vdd.n173 vdd.t97 4.06363
R5397 vdd.n173 vdd.t180 4.06363
R5398 vdd.n171 vdd.t262 4.06363
R5399 vdd.n171 vdd.t12 4.06363
R5400 vdd.n169 vdd.t103 4.06363
R5401 vdd.n169 vdd.t101 4.06363
R5402 vdd.n167 vdd.t182 4.06363
R5403 vdd.n167 vdd.t164 4.06363
R5404 vdd.n82 vdd.t128 4.06363
R5405 vdd.n82 vdd.t10 4.06363
R5406 vdd.n80 vdd.t260 4.06363
R5407 vdd.n80 vdd.t95 4.06363
R5408 vdd.n78 vdd.t99 4.06363
R5409 vdd.n78 vdd.t264 4.06363
R5410 vdd.n76 vdd.t171 4.06363
R5411 vdd.n76 vdd.t141 4.06363
R5412 vdd.n74 vdd.t143 4.06363
R5413 vdd.n74 vdd.t125 4.06363
R5414 vdd.n72 vdd.t107 4.06363
R5415 vdd.n72 vdd.t257 4.06363
R5416 vdd.n70 vdd.t156 4.06363
R5417 vdd.n70 vdd.t137 4.06363
R5418 vdd.n2051 vdd.t121 4.06363
R5419 vdd.n2051 vdd.t259 4.06363
R5420 vdd.n2053 vdd.t240 4.06363
R5421 vdd.n2053 vdd.t16 4.06363
R5422 vdd.n2055 vdd.t256 4.06363
R5423 vdd.n2055 vdd.t113 4.06363
R5424 vdd.n2057 vdd.t131 4.06363
R5425 vdd.n2057 vdd.t266 4.06363
R5426 vdd.n2059 vdd.t267 4.06363
R5427 vdd.n2059 vdd.t190 4.06363
R5428 vdd.n2061 vdd.t124 4.06363
R5429 vdd.n2061 vdd.t258 4.06363
R5430 vdd.n2063 vdd.t111 4.06363
R5431 vdd.n2063 vdd.t158 4.06363
R5432 vdd.n1953 vdd.t7 4.06363
R5433 vdd.n1953 vdd.t189 4.06363
R5434 vdd.n1955 vdd.t181 4.06363
R5435 vdd.n1955 vdd.t241 4.06363
R5436 vdd.n1957 vdd.t177 4.06363
R5437 vdd.n1957 vdd.t14 4.06363
R5438 vdd.n1959 vdd.t185 4.06363
R5439 vdd.n1959 vdd.t245 4.06363
R5440 vdd.n1961 vdd.t165 4.06363
R5441 vdd.n1961 vdd.t149 4.06363
R5442 vdd.n1963 vdd.t132 4.06363
R5443 vdd.n1963 vdd.t178 4.06363
R5444 vdd.n1965 vdd.t119 4.06363
R5445 vdd.n1965 vdd.t166 4.06363
R5446 vdd.n1856 vdd.t8 4.06363
R5447 vdd.n1856 vdd.t261 4.06363
R5448 vdd.n1858 vdd.t147 4.06363
R5449 vdd.n1858 vdd.t263 4.06363
R5450 vdd.n1860 vdd.t153 4.06363
R5451 vdd.n1860 vdd.t246 4.06363
R5452 vdd.n1862 vdd.t142 4.06363
R5453 vdd.n1862 vdd.t173 4.06363
R5454 vdd.n1864 vdd.t5 4.06363
R5455 vdd.n1864 vdd.t179 4.06363
R5456 vdd.n1866 vdd.t157 4.06363
R5457 vdd.n1866 vdd.t139 4.06363
R5458 vdd.n1868 vdd.t120 4.06363
R5459 vdd.n1868 vdd.t134 4.06363
R5460 vdd.n26 vdd.t251 3.9605
R5461 vdd.n26 vdd.t252 3.9605
R5462 vdd.n23 vdd.t176 3.9605
R5463 vdd.n23 vdd.t248 3.9605
R5464 vdd.n21 vdd.t254 3.9605
R5465 vdd.n21 vdd.t122 3.9605
R5466 vdd.n20 vdd.t118 3.9605
R5467 vdd.n20 vdd.t174 3.9605
R5468 vdd.n15 vdd.t253 3.9605
R5469 vdd.n15 vdd.t175 3.9605
R5470 vdd.n16 vdd.t117 3.9605
R5471 vdd.n16 vdd.t249 3.9605
R5472 vdd.n18 vdd.t247 3.9605
R5473 vdd.n18 vdd.t144 3.9605
R5474 vdd.n25 vdd.t250 3.9605
R5475 vdd.n25 vdd.t145 3.9605
R5476 vdd.n2428 vdd.t209 3.85492
R5477 vdd.n1309 vdd.t209 3.85492
R5478 vdd.n2868 vdd.t197 3.85492
R5479 vdd.t197 vdd.n888 3.85492
R5480 vdd.n7 vdd.t239 3.61217
R5481 vdd.n7 vdd.t208 3.61217
R5482 vdd.n8 vdd.t216 3.61217
R5483 vdd.n8 vdd.t232 3.61217
R5484 vdd.n10 vdd.t223 3.61217
R5485 vdd.n10 vdd.t198 3.61217
R5486 vdd.n12 vdd.t205 3.61217
R5487 vdd.n12 vdd.t221 3.61217
R5488 vdd.n5 vdd.t236 3.61217
R5489 vdd.n5 vdd.t218 3.61217
R5490 vdd.n3 vdd.t210 3.61217
R5491 vdd.n3 vdd.t234 3.61217
R5492 vdd.n1 vdd.t195 3.61217
R5493 vdd.n1 vdd.t225 3.61217
R5494 vdd.n0 vdd.t230 3.61217
R5495 vdd.n0 vdd.t213 3.61217
R5496 vdd.n1744 vdd.t47 3.51482
R5497 vdd.n3347 vdd.t51 3.51482
R5498 vdd.n304 vdd.n303 3.49141
R5499 vdd.n249 vdd.n248 3.49141
R5500 vdd.n206 vdd.n205 3.49141
R5501 vdd.n151 vdd.n150 3.49141
R5502 vdd.n109 vdd.n108 3.49141
R5503 vdd.n54 vdd.n53 3.49141
R5504 vdd.n2035 vdd.n2034 3.49141
R5505 vdd.n2090 vdd.n2089 3.49141
R5506 vdd.n1937 vdd.n1936 3.49141
R5507 vdd.n1992 vdd.n1991 3.49141
R5508 vdd.n1840 vdd.n1839 3.49141
R5509 vdd.n1895 vdd.n1894 3.49141
R5510 vdd.n2582 vdd.t235 3.40145
R5511 vdd.n2855 vdd.t220 3.40145
R5512 vdd.n2920 vdd.n2919 3.12245
R5513 vdd.n2376 vdd.n2375 3.12245
R5514 vdd.n2147 vdd.t6 3.06136
R5515 vdd.n1026 vdd.t219 3.06136
R5516 vdd.n2408 vdd.t214 3.06136
R5517 vdd.n2764 vdd.t228 3.06136
R5518 vdd.n2929 vdd.t199 3.06136
R5519 vdd.n3269 vdd.t136 3.06136
R5520 vdd.t13 vdd.n1443 2.83463
R5521 vdd.n624 vdd.t93 2.83463
R5522 vdd.n1330 vdd.t229 2.72126
R5523 vdd.n2904 vdd.t207 2.72126
R5524 vdd.n307 vdd.n286 2.71565
R5525 vdd.n252 vdd.n231 2.71565
R5526 vdd.n209 vdd.n188 2.71565
R5527 vdd.n154 vdd.n133 2.71565
R5528 vdd.n112 vdd.n91 2.71565
R5529 vdd.n57 vdd.n36 2.71565
R5530 vdd.n2038 vdd.n2017 2.71565
R5531 vdd.n2093 vdd.n2072 2.71565
R5532 vdd.n1940 vdd.n1919 2.71565
R5533 vdd.n1995 vdd.n1974 2.71565
R5534 vdd.n1843 vdd.n1822 2.71565
R5535 vdd.n1898 vdd.n1877 2.71565
R5536 vdd.n1811 vdd.t130 2.6079
R5537 vdd.n3379 vdd.t140 2.6079
R5538 vdd.t224 vdd.n970 2.49453
R5539 vdd.n2880 vdd.t215 2.49453
R5540 vdd.n294 vdd.n293 2.4129
R5541 vdd.n239 vdd.n238 2.4129
R5542 vdd.n196 vdd.n195 2.4129
R5543 vdd.n141 vdd.n140 2.4129
R5544 vdd.n99 vdd.n98 2.4129
R5545 vdd.n44 vdd.n43 2.4129
R5546 vdd.n2025 vdd.n2024 2.4129
R5547 vdd.n2080 vdd.n2079 2.4129
R5548 vdd.n1927 vdd.n1926 2.4129
R5549 vdd.n1982 vdd.n1981 2.4129
R5550 vdd.n1830 vdd.n1829 2.4129
R5551 vdd.n1885 vdd.n1884 2.4129
R5552 vdd.t138 vdd.n1472 2.38117
R5553 vdd.n1050 vdd.t22 2.38117
R5554 vdd.n2435 vdd.t64 2.38117
R5555 vdd.n2779 vdd.t68 2.38117
R5556 vdd.n2998 vdd.t18 2.38117
R5557 vdd.n3370 vdd.t105 2.38117
R5558 vdd.n2298 vdd.n1093 2.27742
R5559 vdd.n2298 vdd.n1092 2.27742
R5560 vdd.n3034 vdd.n665 2.27742
R5561 vdd.n3034 vdd.n664 2.27742
R5562 vdd.n3102 vdd.n751 2.27742
R5563 vdd.n3102 vdd.n749 2.27742
R5564 vdd.n2192 vdd.n2191 2.27742
R5565 vdd.n2191 vdd.n1394 2.27742
R5566 vdd.n1769 vdd.t110 2.15444
R5567 vdd.n2384 vdd.t206 2.15444
R5568 vdd.n1330 vdd.t237 2.15444
R5569 vdd.n2904 vdd.t227 2.15444
R5570 vdd.t211 vdd.n846 2.15444
R5571 vdd.n3361 vdd.t9 2.15444
R5572 vdd.n308 vdd.n284 1.93989
R5573 vdd.n253 vdd.n229 1.93989
R5574 vdd.n210 vdd.n186 1.93989
R5575 vdd.n155 vdd.n131 1.93989
R5576 vdd.n113 vdd.n89 1.93989
R5577 vdd.n58 vdd.n34 1.93989
R5578 vdd.n2039 vdd.n2015 1.93989
R5579 vdd.n2094 vdd.n2070 1.93989
R5580 vdd.n1941 vdd.n1917 1.93989
R5581 vdd.n1996 vdd.n1972 1.93989
R5582 vdd.n1844 vdd.n1820 1.93989
R5583 vdd.n1899 vdd.n1875 1.93989
R5584 vdd.n2408 vdd.t194 1.81434
R5585 vdd.n2764 vdd.t231 1.81434
R5586 vdd.n1761 vdd.t108 1.70098
R5587 vdd.n3355 vdd.t150 1.70098
R5588 vdd.n2402 vdd.t212 1.58761
R5589 vdd.n872 vdd.t238 1.58761
R5590 vdd.n1777 vdd.t123 1.47425
R5591 vdd.n349 vdd.t0 1.47425
R5592 vdd.n1802 vdd.t148 1.24752
R5593 vdd.t30 vdd.n1407 1.24752
R5594 vdd.n2378 vdd.t200 1.24752
R5595 vdd.n995 vdd.t202 1.24752
R5596 vdd.n2898 vdd.t192 1.24752
R5597 vdd.n849 vdd.t201 1.24752
R5598 vdd.n659 vdd.t26 1.24752
R5599 vdd.t98 vdd.n3377 1.24752
R5600 vdd.n319 vdd.n279 1.16414
R5601 vdd.n312 vdd.n311 1.16414
R5602 vdd.n264 vdd.n224 1.16414
R5603 vdd.n257 vdd.n256 1.16414
R5604 vdd.n221 vdd.n181 1.16414
R5605 vdd.n214 vdd.n213 1.16414
R5606 vdd.n166 vdd.n126 1.16414
R5607 vdd.n159 vdd.n158 1.16414
R5608 vdd.n124 vdd.n84 1.16414
R5609 vdd.n117 vdd.n116 1.16414
R5610 vdd.n69 vdd.n29 1.16414
R5611 vdd.n62 vdd.n61 1.16414
R5612 vdd.n2050 vdd.n2010 1.16414
R5613 vdd.n2043 vdd.n2042 1.16414
R5614 vdd.n2105 vdd.n2065 1.16414
R5615 vdd.n2098 vdd.n2097 1.16414
R5616 vdd.n1952 vdd.n1912 1.16414
R5617 vdd.n1945 vdd.n1944 1.16414
R5618 vdd.n2007 vdd.n1967 1.16414
R5619 vdd.n2000 vdd.n1999 1.16414
R5620 vdd.n1855 vdd.n1815 1.16414
R5621 vdd.n1848 vdd.n1847 1.16414
R5622 vdd.n1910 vdd.n1870 1.16414
R5623 vdd.n1903 vdd.n1902 1.16414
R5624 vdd.n1454 vdd.t152 1.02079
R5625 vdd.t72 vdd.t200 1.02079
R5626 vdd.t201 vdd.t40 1.02079
R5627 vdd.t11 vdd.n613 1.02079
R5628 vdd.n1633 vdd.n1512 0.970197
R5629 vdd.n2189 vdd.n2188 0.970197
R5630 vdd.n599 vdd.n407 0.970197
R5631 vdd.n3109 vdd.n3107 0.970197
R5632 vdd.n2108 vdd.n28 0.956323
R5633 vdd vdd.n3384 0.94849
R5634 vdd.n2139 vdd.t15 0.794056
R5635 vdd.n3278 vdd.t102 0.794056
R5636 vdd.n2155 vdd.t169 0.567326
R5637 vdd.t161 vdd.n642 0.567326
R5638 vdd.n2179 vdd.n1094 0.482207
R5639 vdd.n3234 vdd.n3233 0.482207
R5640 vdd.n444 vdd.n443 0.482207
R5641 vdd.n3341 vdd.n3340 0.482207
R5642 vdd.n3240 vdd.n656 0.482207
R5643 vdd.n2169 vdd.n1395 0.482207
R5644 vdd.n1740 vdd.n1739 0.482207
R5645 vdd.n1546 vdd.n1503 0.482207
R5646 vdd.n4 vdd.n2 0.459552
R5647 vdd.n11 vdd.n9 0.459552
R5648 vdd.t233 vdd.n947 0.453961
R5649 vdd.n2862 vdd.t222 0.453961
R5650 vdd.n317 vdd.n316 0.388379
R5651 vdd.n283 vdd.n281 0.388379
R5652 vdd.n262 vdd.n261 0.388379
R5653 vdd.n228 vdd.n226 0.388379
R5654 vdd.n219 vdd.n218 0.388379
R5655 vdd.n185 vdd.n183 0.388379
R5656 vdd.n164 vdd.n163 0.388379
R5657 vdd.n130 vdd.n128 0.388379
R5658 vdd.n122 vdd.n121 0.388379
R5659 vdd.n88 vdd.n86 0.388379
R5660 vdd.n67 vdd.n66 0.388379
R5661 vdd.n33 vdd.n31 0.388379
R5662 vdd.n2048 vdd.n2047 0.388379
R5663 vdd.n2014 vdd.n2012 0.388379
R5664 vdd.n2103 vdd.n2102 0.388379
R5665 vdd.n2069 vdd.n2067 0.388379
R5666 vdd.n1950 vdd.n1949 0.388379
R5667 vdd.n1916 vdd.n1914 0.388379
R5668 vdd.n2005 vdd.n2004 0.388379
R5669 vdd.n1971 vdd.n1969 0.388379
R5670 vdd.n1853 vdd.n1852 0.388379
R5671 vdd.n1819 vdd.n1817 0.388379
R5672 vdd.n1908 vdd.n1907 0.388379
R5673 vdd.n1874 vdd.n1872 0.388379
R5674 vdd.n19 vdd.n17 0.387128
R5675 vdd.n24 vdd.n22 0.387128
R5676 vdd.n6 vdd.n4 0.358259
R5677 vdd.n13 vdd.n11 0.358259
R5678 vdd.n268 vdd.n266 0.358259
R5679 vdd.n270 vdd.n268 0.358259
R5680 vdd.n272 vdd.n270 0.358259
R5681 vdd.n274 vdd.n272 0.358259
R5682 vdd.n276 vdd.n274 0.358259
R5683 vdd.n278 vdd.n276 0.358259
R5684 vdd.n320 vdd.n278 0.358259
R5685 vdd.n170 vdd.n168 0.358259
R5686 vdd.n172 vdd.n170 0.358259
R5687 vdd.n174 vdd.n172 0.358259
R5688 vdd.n176 vdd.n174 0.358259
R5689 vdd.n178 vdd.n176 0.358259
R5690 vdd.n180 vdd.n178 0.358259
R5691 vdd.n222 vdd.n180 0.358259
R5692 vdd.n73 vdd.n71 0.358259
R5693 vdd.n75 vdd.n73 0.358259
R5694 vdd.n77 vdd.n75 0.358259
R5695 vdd.n79 vdd.n77 0.358259
R5696 vdd.n81 vdd.n79 0.358259
R5697 vdd.n83 vdd.n81 0.358259
R5698 vdd.n125 vdd.n83 0.358259
R5699 vdd.n2106 vdd.n2064 0.358259
R5700 vdd.n2064 vdd.n2062 0.358259
R5701 vdd.n2062 vdd.n2060 0.358259
R5702 vdd.n2060 vdd.n2058 0.358259
R5703 vdd.n2058 vdd.n2056 0.358259
R5704 vdd.n2056 vdd.n2054 0.358259
R5705 vdd.n2054 vdd.n2052 0.358259
R5706 vdd.n2008 vdd.n1966 0.358259
R5707 vdd.n1966 vdd.n1964 0.358259
R5708 vdd.n1964 vdd.n1962 0.358259
R5709 vdd.n1962 vdd.n1960 0.358259
R5710 vdd.n1960 vdd.n1958 0.358259
R5711 vdd.n1958 vdd.n1956 0.358259
R5712 vdd.n1956 vdd.n1954 0.358259
R5713 vdd.n1911 vdd.n1869 0.358259
R5714 vdd.n1869 vdd.n1867 0.358259
R5715 vdd.n1867 vdd.n1865 0.358259
R5716 vdd.n1865 vdd.n1863 0.358259
R5717 vdd.n1863 vdd.n1861 0.358259
R5718 vdd.n1861 vdd.n1859 0.358259
R5719 vdd.n1859 vdd.n1857 0.358259
R5720 vdd.t203 vdd.n1023 0.340595
R5721 vdd.n2414 vdd.t193 0.340595
R5722 vdd.t196 vdd.n876 0.340595
R5723 vdd.n2935 vdd.t226 0.340595
R5724 vdd.n14 vdd.n6 0.334552
R5725 vdd.n14 vdd.n13 0.334552
R5726 vdd.n27 vdd.n19 0.21707
R5727 vdd.n27 vdd.n24 0.21707
R5728 vdd.n318 vdd.n280 0.155672
R5729 vdd.n310 vdd.n280 0.155672
R5730 vdd.n310 vdd.n309 0.155672
R5731 vdd.n309 vdd.n285 0.155672
R5732 vdd.n302 vdd.n285 0.155672
R5733 vdd.n302 vdd.n301 0.155672
R5734 vdd.n301 vdd.n289 0.155672
R5735 vdd.n294 vdd.n289 0.155672
R5736 vdd.n263 vdd.n225 0.155672
R5737 vdd.n255 vdd.n225 0.155672
R5738 vdd.n255 vdd.n254 0.155672
R5739 vdd.n254 vdd.n230 0.155672
R5740 vdd.n247 vdd.n230 0.155672
R5741 vdd.n247 vdd.n246 0.155672
R5742 vdd.n246 vdd.n234 0.155672
R5743 vdd.n239 vdd.n234 0.155672
R5744 vdd.n220 vdd.n182 0.155672
R5745 vdd.n212 vdd.n182 0.155672
R5746 vdd.n212 vdd.n211 0.155672
R5747 vdd.n211 vdd.n187 0.155672
R5748 vdd.n204 vdd.n187 0.155672
R5749 vdd.n204 vdd.n203 0.155672
R5750 vdd.n203 vdd.n191 0.155672
R5751 vdd.n196 vdd.n191 0.155672
R5752 vdd.n165 vdd.n127 0.155672
R5753 vdd.n157 vdd.n127 0.155672
R5754 vdd.n157 vdd.n156 0.155672
R5755 vdd.n156 vdd.n132 0.155672
R5756 vdd.n149 vdd.n132 0.155672
R5757 vdd.n149 vdd.n148 0.155672
R5758 vdd.n148 vdd.n136 0.155672
R5759 vdd.n141 vdd.n136 0.155672
R5760 vdd.n123 vdd.n85 0.155672
R5761 vdd.n115 vdd.n85 0.155672
R5762 vdd.n115 vdd.n114 0.155672
R5763 vdd.n114 vdd.n90 0.155672
R5764 vdd.n107 vdd.n90 0.155672
R5765 vdd.n107 vdd.n106 0.155672
R5766 vdd.n106 vdd.n94 0.155672
R5767 vdd.n99 vdd.n94 0.155672
R5768 vdd.n68 vdd.n30 0.155672
R5769 vdd.n60 vdd.n30 0.155672
R5770 vdd.n60 vdd.n59 0.155672
R5771 vdd.n59 vdd.n35 0.155672
R5772 vdd.n52 vdd.n35 0.155672
R5773 vdd.n52 vdd.n51 0.155672
R5774 vdd.n51 vdd.n39 0.155672
R5775 vdd.n44 vdd.n39 0.155672
R5776 vdd.n2049 vdd.n2011 0.155672
R5777 vdd.n2041 vdd.n2011 0.155672
R5778 vdd.n2041 vdd.n2040 0.155672
R5779 vdd.n2040 vdd.n2016 0.155672
R5780 vdd.n2033 vdd.n2016 0.155672
R5781 vdd.n2033 vdd.n2032 0.155672
R5782 vdd.n2032 vdd.n2020 0.155672
R5783 vdd.n2025 vdd.n2020 0.155672
R5784 vdd.n2104 vdd.n2066 0.155672
R5785 vdd.n2096 vdd.n2066 0.155672
R5786 vdd.n2096 vdd.n2095 0.155672
R5787 vdd.n2095 vdd.n2071 0.155672
R5788 vdd.n2088 vdd.n2071 0.155672
R5789 vdd.n2088 vdd.n2087 0.155672
R5790 vdd.n2087 vdd.n2075 0.155672
R5791 vdd.n2080 vdd.n2075 0.155672
R5792 vdd.n1951 vdd.n1913 0.155672
R5793 vdd.n1943 vdd.n1913 0.155672
R5794 vdd.n1943 vdd.n1942 0.155672
R5795 vdd.n1942 vdd.n1918 0.155672
R5796 vdd.n1935 vdd.n1918 0.155672
R5797 vdd.n1935 vdd.n1934 0.155672
R5798 vdd.n1934 vdd.n1922 0.155672
R5799 vdd.n1927 vdd.n1922 0.155672
R5800 vdd.n2006 vdd.n1968 0.155672
R5801 vdd.n1998 vdd.n1968 0.155672
R5802 vdd.n1998 vdd.n1997 0.155672
R5803 vdd.n1997 vdd.n1973 0.155672
R5804 vdd.n1990 vdd.n1973 0.155672
R5805 vdd.n1990 vdd.n1989 0.155672
R5806 vdd.n1989 vdd.n1977 0.155672
R5807 vdd.n1982 vdd.n1977 0.155672
R5808 vdd.n1854 vdd.n1816 0.155672
R5809 vdd.n1846 vdd.n1816 0.155672
R5810 vdd.n1846 vdd.n1845 0.155672
R5811 vdd.n1845 vdd.n1821 0.155672
R5812 vdd.n1838 vdd.n1821 0.155672
R5813 vdd.n1838 vdd.n1837 0.155672
R5814 vdd.n1837 vdd.n1825 0.155672
R5815 vdd.n1830 vdd.n1825 0.155672
R5816 vdd.n1909 vdd.n1871 0.155672
R5817 vdd.n1901 vdd.n1871 0.155672
R5818 vdd.n1901 vdd.n1900 0.155672
R5819 vdd.n1900 vdd.n1876 0.155672
R5820 vdd.n1893 vdd.n1876 0.155672
R5821 vdd.n1893 vdd.n1892 0.155672
R5822 vdd.n1892 vdd.n1880 0.155672
R5823 vdd.n1885 vdd.n1880 0.155672
R5824 vdd.n1099 vdd.n1091 0.152939
R5825 vdd.n1103 vdd.n1099 0.152939
R5826 vdd.n1104 vdd.n1103 0.152939
R5827 vdd.n1105 vdd.n1104 0.152939
R5828 vdd.n1106 vdd.n1105 0.152939
R5829 vdd.n1110 vdd.n1106 0.152939
R5830 vdd.n1111 vdd.n1110 0.152939
R5831 vdd.n1112 vdd.n1111 0.152939
R5832 vdd.n1113 vdd.n1112 0.152939
R5833 vdd.n1117 vdd.n1113 0.152939
R5834 vdd.n1118 vdd.n1117 0.152939
R5835 vdd.n1119 vdd.n1118 0.152939
R5836 vdd.n2262 vdd.n1119 0.152939
R5837 vdd.n2262 vdd.n2261 0.152939
R5838 vdd.n2261 vdd.n2260 0.152939
R5839 vdd.n2260 vdd.n1125 0.152939
R5840 vdd.n1130 vdd.n1125 0.152939
R5841 vdd.n1131 vdd.n1130 0.152939
R5842 vdd.n1132 vdd.n1131 0.152939
R5843 vdd.n1136 vdd.n1132 0.152939
R5844 vdd.n1137 vdd.n1136 0.152939
R5845 vdd.n1138 vdd.n1137 0.152939
R5846 vdd.n1139 vdd.n1138 0.152939
R5847 vdd.n1143 vdd.n1139 0.152939
R5848 vdd.n1144 vdd.n1143 0.152939
R5849 vdd.n1145 vdd.n1144 0.152939
R5850 vdd.n1146 vdd.n1145 0.152939
R5851 vdd.n1150 vdd.n1146 0.152939
R5852 vdd.n1151 vdd.n1150 0.152939
R5853 vdd.n1152 vdd.n1151 0.152939
R5854 vdd.n1153 vdd.n1152 0.152939
R5855 vdd.n1157 vdd.n1153 0.152939
R5856 vdd.n1158 vdd.n1157 0.152939
R5857 vdd.n1159 vdd.n1158 0.152939
R5858 vdd.n2223 vdd.n1159 0.152939
R5859 vdd.n2223 vdd.n2222 0.152939
R5860 vdd.n2222 vdd.n2221 0.152939
R5861 vdd.n2221 vdd.n1165 0.152939
R5862 vdd.n1170 vdd.n1165 0.152939
R5863 vdd.n1171 vdd.n1170 0.152939
R5864 vdd.n1172 vdd.n1171 0.152939
R5865 vdd.n1176 vdd.n1172 0.152939
R5866 vdd.n1177 vdd.n1176 0.152939
R5867 vdd.n1178 vdd.n1177 0.152939
R5868 vdd.n1179 vdd.n1178 0.152939
R5869 vdd.n1183 vdd.n1179 0.152939
R5870 vdd.n1184 vdd.n1183 0.152939
R5871 vdd.n1185 vdd.n1184 0.152939
R5872 vdd.n1186 vdd.n1185 0.152939
R5873 vdd.n1190 vdd.n1186 0.152939
R5874 vdd.n1191 vdd.n1190 0.152939
R5875 vdd.n2297 vdd.n1094 0.152939
R5876 vdd.n2111 vdd.n2110 0.152939
R5877 vdd.n2111 vdd.n1446 0.152939
R5878 vdd.n2125 vdd.n1446 0.152939
R5879 vdd.n2126 vdd.n2125 0.152939
R5880 vdd.n2127 vdd.n2126 0.152939
R5881 vdd.n2127 vdd.n1434 0.152939
R5882 vdd.n2142 vdd.n1434 0.152939
R5883 vdd.n2143 vdd.n2142 0.152939
R5884 vdd.n2144 vdd.n2143 0.152939
R5885 vdd.n2144 vdd.n1423 0.152939
R5886 vdd.n2159 vdd.n1423 0.152939
R5887 vdd.n2160 vdd.n2159 0.152939
R5888 vdd.n2161 vdd.n2160 0.152939
R5889 vdd.n2161 vdd.n1411 0.152939
R5890 vdd.n2177 vdd.n1411 0.152939
R5891 vdd.n2178 vdd.n2177 0.152939
R5892 vdd.n2179 vdd.n2178 0.152939
R5893 vdd.n670 vdd.n667 0.152939
R5894 vdd.n671 vdd.n670 0.152939
R5895 vdd.n672 vdd.n671 0.152939
R5896 vdd.n673 vdd.n672 0.152939
R5897 vdd.n676 vdd.n673 0.152939
R5898 vdd.n677 vdd.n676 0.152939
R5899 vdd.n678 vdd.n677 0.152939
R5900 vdd.n679 vdd.n678 0.152939
R5901 vdd.n682 vdd.n679 0.152939
R5902 vdd.n683 vdd.n682 0.152939
R5903 vdd.n684 vdd.n683 0.152939
R5904 vdd.n685 vdd.n684 0.152939
R5905 vdd.n690 vdd.n685 0.152939
R5906 vdd.n691 vdd.n690 0.152939
R5907 vdd.n692 vdd.n691 0.152939
R5908 vdd.n693 vdd.n692 0.152939
R5909 vdd.n696 vdd.n693 0.152939
R5910 vdd.n697 vdd.n696 0.152939
R5911 vdd.n698 vdd.n697 0.152939
R5912 vdd.n699 vdd.n698 0.152939
R5913 vdd.n702 vdd.n699 0.152939
R5914 vdd.n703 vdd.n702 0.152939
R5915 vdd.n704 vdd.n703 0.152939
R5916 vdd.n705 vdd.n704 0.152939
R5917 vdd.n708 vdd.n705 0.152939
R5918 vdd.n709 vdd.n708 0.152939
R5919 vdd.n710 vdd.n709 0.152939
R5920 vdd.n711 vdd.n710 0.152939
R5921 vdd.n714 vdd.n711 0.152939
R5922 vdd.n715 vdd.n714 0.152939
R5923 vdd.n716 vdd.n715 0.152939
R5924 vdd.n717 vdd.n716 0.152939
R5925 vdd.n720 vdd.n717 0.152939
R5926 vdd.n721 vdd.n720 0.152939
R5927 vdd.n3150 vdd.n721 0.152939
R5928 vdd.n3150 vdd.n3149 0.152939
R5929 vdd.n3149 vdd.n3148 0.152939
R5930 vdd.n3148 vdd.n725 0.152939
R5931 vdd.n730 vdd.n725 0.152939
R5932 vdd.n731 vdd.n730 0.152939
R5933 vdd.n734 vdd.n731 0.152939
R5934 vdd.n735 vdd.n734 0.152939
R5935 vdd.n736 vdd.n735 0.152939
R5936 vdd.n737 vdd.n736 0.152939
R5937 vdd.n740 vdd.n737 0.152939
R5938 vdd.n741 vdd.n740 0.152939
R5939 vdd.n742 vdd.n741 0.152939
R5940 vdd.n743 vdd.n742 0.152939
R5941 vdd.n746 vdd.n743 0.152939
R5942 vdd.n747 vdd.n746 0.152939
R5943 vdd.n748 vdd.n747 0.152939
R5944 vdd.n3233 vdd.n661 0.152939
R5945 vdd.n3234 vdd.n651 0.152939
R5946 vdd.n3248 vdd.n651 0.152939
R5947 vdd.n3249 vdd.n3248 0.152939
R5948 vdd.n3250 vdd.n3249 0.152939
R5949 vdd.n3250 vdd.n639 0.152939
R5950 vdd.n3264 vdd.n639 0.152939
R5951 vdd.n3265 vdd.n3264 0.152939
R5952 vdd.n3266 vdd.n3265 0.152939
R5953 vdd.n3266 vdd.n627 0.152939
R5954 vdd.n3281 vdd.n627 0.152939
R5955 vdd.n3282 vdd.n3281 0.152939
R5956 vdd.n3283 vdd.n3282 0.152939
R5957 vdd.n3283 vdd.n616 0.152939
R5958 vdd.n3300 vdd.n616 0.152939
R5959 vdd.n3301 vdd.n3300 0.152939
R5960 vdd.n3302 vdd.n3301 0.152939
R5961 vdd.n3302 vdd.n322 0.152939
R5962 vdd.n3382 vdd.n323 0.152939
R5963 vdd.n334 vdd.n323 0.152939
R5964 vdd.n335 vdd.n334 0.152939
R5965 vdd.n336 vdd.n335 0.152939
R5966 vdd.n343 vdd.n336 0.152939
R5967 vdd.n344 vdd.n343 0.152939
R5968 vdd.n345 vdd.n344 0.152939
R5969 vdd.n346 vdd.n345 0.152939
R5970 vdd.n354 vdd.n346 0.152939
R5971 vdd.n355 vdd.n354 0.152939
R5972 vdd.n356 vdd.n355 0.152939
R5973 vdd.n357 vdd.n356 0.152939
R5974 vdd.n365 vdd.n357 0.152939
R5975 vdd.n366 vdd.n365 0.152939
R5976 vdd.n367 vdd.n366 0.152939
R5977 vdd.n368 vdd.n367 0.152939
R5978 vdd.n443 vdd.n368 0.152939
R5979 vdd.n444 vdd.n442 0.152939
R5980 vdd.n451 vdd.n442 0.152939
R5981 vdd.n452 vdd.n451 0.152939
R5982 vdd.n453 vdd.n452 0.152939
R5983 vdd.n453 vdd.n440 0.152939
R5984 vdd.n461 vdd.n440 0.152939
R5985 vdd.n462 vdd.n461 0.152939
R5986 vdd.n463 vdd.n462 0.152939
R5987 vdd.n463 vdd.n438 0.152939
R5988 vdd.n471 vdd.n438 0.152939
R5989 vdd.n472 vdd.n471 0.152939
R5990 vdd.n473 vdd.n472 0.152939
R5991 vdd.n473 vdd.n436 0.152939
R5992 vdd.n481 vdd.n436 0.152939
R5993 vdd.n482 vdd.n481 0.152939
R5994 vdd.n483 vdd.n482 0.152939
R5995 vdd.n483 vdd.n434 0.152939
R5996 vdd.n491 vdd.n434 0.152939
R5997 vdd.n492 vdd.n491 0.152939
R5998 vdd.n493 vdd.n492 0.152939
R5999 vdd.n493 vdd.n430 0.152939
R6000 vdd.n501 vdd.n430 0.152939
R6001 vdd.n502 vdd.n501 0.152939
R6002 vdd.n503 vdd.n502 0.152939
R6003 vdd.n503 vdd.n428 0.152939
R6004 vdd.n511 vdd.n428 0.152939
R6005 vdd.n512 vdd.n511 0.152939
R6006 vdd.n513 vdd.n512 0.152939
R6007 vdd.n513 vdd.n426 0.152939
R6008 vdd.n521 vdd.n426 0.152939
R6009 vdd.n522 vdd.n521 0.152939
R6010 vdd.n523 vdd.n522 0.152939
R6011 vdd.n523 vdd.n424 0.152939
R6012 vdd.n531 vdd.n424 0.152939
R6013 vdd.n532 vdd.n531 0.152939
R6014 vdd.n533 vdd.n532 0.152939
R6015 vdd.n533 vdd.n422 0.152939
R6016 vdd.n541 vdd.n422 0.152939
R6017 vdd.n542 vdd.n541 0.152939
R6018 vdd.n543 vdd.n542 0.152939
R6019 vdd.n543 vdd.n418 0.152939
R6020 vdd.n551 vdd.n418 0.152939
R6021 vdd.n552 vdd.n551 0.152939
R6022 vdd.n553 vdd.n552 0.152939
R6023 vdd.n553 vdd.n416 0.152939
R6024 vdd.n561 vdd.n416 0.152939
R6025 vdd.n562 vdd.n561 0.152939
R6026 vdd.n563 vdd.n562 0.152939
R6027 vdd.n563 vdd.n414 0.152939
R6028 vdd.n571 vdd.n414 0.152939
R6029 vdd.n572 vdd.n571 0.152939
R6030 vdd.n573 vdd.n572 0.152939
R6031 vdd.n573 vdd.n412 0.152939
R6032 vdd.n581 vdd.n412 0.152939
R6033 vdd.n582 vdd.n581 0.152939
R6034 vdd.n583 vdd.n582 0.152939
R6035 vdd.n583 vdd.n410 0.152939
R6036 vdd.n591 vdd.n410 0.152939
R6037 vdd.n592 vdd.n591 0.152939
R6038 vdd.n593 vdd.n592 0.152939
R6039 vdd.n593 vdd.n408 0.152939
R6040 vdd.n600 vdd.n408 0.152939
R6041 vdd.n3341 vdd.n600 0.152939
R6042 vdd.n3241 vdd.n3240 0.152939
R6043 vdd.n3242 vdd.n3241 0.152939
R6044 vdd.n3242 vdd.n645 0.152939
R6045 vdd.n3256 vdd.n645 0.152939
R6046 vdd.n3257 vdd.n3256 0.152939
R6047 vdd.n3258 vdd.n3257 0.152939
R6048 vdd.n3258 vdd.n632 0.152939
R6049 vdd.n3272 vdd.n632 0.152939
R6050 vdd.n3273 vdd.n3272 0.152939
R6051 vdd.n3274 vdd.n3273 0.152939
R6052 vdd.n3274 vdd.n621 0.152939
R6053 vdd.n3289 vdd.n621 0.152939
R6054 vdd.n3290 vdd.n3289 0.152939
R6055 vdd.n3291 vdd.n3290 0.152939
R6056 vdd.n3293 vdd.n3291 0.152939
R6057 vdd.n3293 vdd.n3292 0.152939
R6058 vdd.n3292 vdd.n611 0.152939
R6059 vdd.n611 vdd.n609 0.152939
R6060 vdd.n3311 vdd.n609 0.152939
R6061 vdd.n3312 vdd.n3311 0.152939
R6062 vdd.n3313 vdd.n3312 0.152939
R6063 vdd.n3313 vdd.n607 0.152939
R6064 vdd.n3318 vdd.n607 0.152939
R6065 vdd.n3319 vdd.n3318 0.152939
R6066 vdd.n3320 vdd.n3319 0.152939
R6067 vdd.n3320 vdd.n605 0.152939
R6068 vdd.n3325 vdd.n605 0.152939
R6069 vdd.n3326 vdd.n3325 0.152939
R6070 vdd.n3327 vdd.n3326 0.152939
R6071 vdd.n3327 vdd.n603 0.152939
R6072 vdd.n3333 vdd.n603 0.152939
R6073 vdd.n3334 vdd.n3333 0.152939
R6074 vdd.n3335 vdd.n3334 0.152939
R6075 vdd.n3335 vdd.n601 0.152939
R6076 vdd.n3340 vdd.n601 0.152939
R6077 vdd.n3103 vdd.n656 0.152939
R6078 vdd.n2190 vdd.n1395 0.152939
R6079 vdd.n1741 vdd.n1740 0.152939
R6080 vdd.n1741 vdd.n1497 0.152939
R6081 vdd.n1755 vdd.n1497 0.152939
R6082 vdd.n1756 vdd.n1755 0.152939
R6083 vdd.n1757 vdd.n1756 0.152939
R6084 vdd.n1757 vdd.n1485 0.152939
R6085 vdd.n1772 vdd.n1485 0.152939
R6086 vdd.n1773 vdd.n1772 0.152939
R6087 vdd.n1774 vdd.n1773 0.152939
R6088 vdd.n1774 vdd.n1475 0.152939
R6089 vdd.n1789 vdd.n1475 0.152939
R6090 vdd.n1790 vdd.n1789 0.152939
R6091 vdd.n1791 vdd.n1790 0.152939
R6092 vdd.n1791 vdd.n1462 0.152939
R6093 vdd.n1805 vdd.n1462 0.152939
R6094 vdd.n1806 vdd.n1805 0.152939
R6095 vdd.n1807 vdd.n1806 0.152939
R6096 vdd.n1807 vdd.n1451 0.152939
R6097 vdd.n2117 vdd.n1451 0.152939
R6098 vdd.n2118 vdd.n2117 0.152939
R6099 vdd.n2119 vdd.n2118 0.152939
R6100 vdd.n2119 vdd.n1440 0.152939
R6101 vdd.n2133 vdd.n1440 0.152939
R6102 vdd.n2134 vdd.n2133 0.152939
R6103 vdd.n2135 vdd.n2134 0.152939
R6104 vdd.n2135 vdd.n1428 0.152939
R6105 vdd.n2150 vdd.n1428 0.152939
R6106 vdd.n2151 vdd.n2150 0.152939
R6107 vdd.n2152 vdd.n2151 0.152939
R6108 vdd.n2152 vdd.n1418 0.152939
R6109 vdd.n2167 vdd.n1418 0.152939
R6110 vdd.n2168 vdd.n2167 0.152939
R6111 vdd.n2171 vdd.n2168 0.152939
R6112 vdd.n2171 vdd.n2170 0.152939
R6113 vdd.n2170 vdd.n2169 0.152939
R6114 vdd.n1731 vdd.n1546 0.152939
R6115 vdd.n1731 vdd.n1730 0.152939
R6116 vdd.n1730 vdd.n1729 0.152939
R6117 vdd.n1729 vdd.n1548 0.152939
R6118 vdd.n1725 vdd.n1548 0.152939
R6119 vdd.n1725 vdd.n1724 0.152939
R6120 vdd.n1724 vdd.n1723 0.152939
R6121 vdd.n1723 vdd.n1553 0.152939
R6122 vdd.n1719 vdd.n1553 0.152939
R6123 vdd.n1719 vdd.n1718 0.152939
R6124 vdd.n1718 vdd.n1717 0.152939
R6125 vdd.n1717 vdd.n1559 0.152939
R6126 vdd.n1713 vdd.n1559 0.152939
R6127 vdd.n1713 vdd.n1712 0.152939
R6128 vdd.n1712 vdd.n1711 0.152939
R6129 vdd.n1711 vdd.n1565 0.152939
R6130 vdd.n1707 vdd.n1565 0.152939
R6131 vdd.n1707 vdd.n1706 0.152939
R6132 vdd.n1706 vdd.n1705 0.152939
R6133 vdd.n1705 vdd.n1571 0.152939
R6134 vdd.n1697 vdd.n1571 0.152939
R6135 vdd.n1697 vdd.n1696 0.152939
R6136 vdd.n1696 vdd.n1695 0.152939
R6137 vdd.n1695 vdd.n1575 0.152939
R6138 vdd.n1691 vdd.n1575 0.152939
R6139 vdd.n1691 vdd.n1690 0.152939
R6140 vdd.n1690 vdd.n1689 0.152939
R6141 vdd.n1689 vdd.n1581 0.152939
R6142 vdd.n1685 vdd.n1581 0.152939
R6143 vdd.n1685 vdd.n1684 0.152939
R6144 vdd.n1684 vdd.n1683 0.152939
R6145 vdd.n1683 vdd.n1587 0.152939
R6146 vdd.n1679 vdd.n1587 0.152939
R6147 vdd.n1679 vdd.n1678 0.152939
R6148 vdd.n1678 vdd.n1677 0.152939
R6149 vdd.n1677 vdd.n1593 0.152939
R6150 vdd.n1673 vdd.n1593 0.152939
R6151 vdd.n1673 vdd.n1672 0.152939
R6152 vdd.n1672 vdd.n1671 0.152939
R6153 vdd.n1671 vdd.n1599 0.152939
R6154 vdd.n1664 vdd.n1599 0.152939
R6155 vdd.n1664 vdd.n1663 0.152939
R6156 vdd.n1663 vdd.n1662 0.152939
R6157 vdd.n1662 vdd.n1604 0.152939
R6158 vdd.n1658 vdd.n1604 0.152939
R6159 vdd.n1658 vdd.n1657 0.152939
R6160 vdd.n1657 vdd.n1656 0.152939
R6161 vdd.n1656 vdd.n1610 0.152939
R6162 vdd.n1652 vdd.n1610 0.152939
R6163 vdd.n1652 vdd.n1651 0.152939
R6164 vdd.n1651 vdd.n1650 0.152939
R6165 vdd.n1650 vdd.n1616 0.152939
R6166 vdd.n1646 vdd.n1616 0.152939
R6167 vdd.n1646 vdd.n1645 0.152939
R6168 vdd.n1645 vdd.n1644 0.152939
R6169 vdd.n1644 vdd.n1622 0.152939
R6170 vdd.n1640 vdd.n1622 0.152939
R6171 vdd.n1640 vdd.n1639 0.152939
R6172 vdd.n1639 vdd.n1638 0.152939
R6173 vdd.n1638 vdd.n1628 0.152939
R6174 vdd.n1634 vdd.n1628 0.152939
R6175 vdd.n1634 vdd.n1509 0.152939
R6176 vdd.n1739 vdd.n1509 0.152939
R6177 vdd.n1747 vdd.n1503 0.152939
R6178 vdd.n1748 vdd.n1747 0.152939
R6179 vdd.n1749 vdd.n1748 0.152939
R6180 vdd.n1749 vdd.n1491 0.152939
R6181 vdd.n1764 vdd.n1491 0.152939
R6182 vdd.n1765 vdd.n1764 0.152939
R6183 vdd.n1766 vdd.n1765 0.152939
R6184 vdd.n1766 vdd.n1480 0.152939
R6185 vdd.n1781 vdd.n1480 0.152939
R6186 vdd.n1782 vdd.n1781 0.152939
R6187 vdd.n1783 vdd.n1782 0.152939
R6188 vdd.n1783 vdd.n1469 0.152939
R6189 vdd.n1797 vdd.n1469 0.152939
R6190 vdd.n1798 vdd.n1797 0.152939
R6191 vdd.n1799 vdd.n1798 0.152939
R6192 vdd.n1799 vdd.n1457 0.152939
R6193 vdd.n1814 vdd.n1457 0.152939
R6194 vdd.n2298 vdd.n2297 0.110256
R6195 vdd.n3034 vdd.n661 0.110256
R6196 vdd.n3103 vdd.n3102 0.110256
R6197 vdd.n2191 vdd.n2190 0.110256
R6198 vdd.n2110 vdd.n2109 0.0695946
R6199 vdd.n3383 vdd.n322 0.0695946
R6200 vdd.n3383 vdd.n3382 0.0695946
R6201 vdd.n2109 vdd.n1814 0.0695946
R6202 vdd.n2298 vdd.n1091 0.0431829
R6203 vdd.n2191 vdd.n1191 0.0431829
R6204 vdd.n3034 vdd.n667 0.0431829
R6205 vdd.n3102 vdd.n748 0.0431829
R6206 vdd vdd.n28 0.00833333
R6207 a_n7636_8799.n176 a_n7636_8799.t51 485.149
R6208 a_n7636_8799.n192 a_n7636_8799.t60 485.149
R6209 a_n7636_8799.n209 a_n7636_8799.t92 485.149
R6210 a_n7636_8799.n125 a_n7636_8799.t112 485.149
R6211 a_n7636_8799.n141 a_n7636_8799.t126 485.149
R6212 a_n7636_8799.n158 a_n7636_8799.t90 485.149
R6213 a_n7636_8799.n186 a_n7636_8799.t71 464.166
R6214 a_n7636_8799.n185 a_n7636_8799.t52 464.166
R6215 a_n7636_8799.n171 a_n7636_8799.t116 464.166
R6216 a_n7636_8799.n184 a_n7636_8799.t83 464.166
R6217 a_n7636_8799.n183 a_n7636_8799.t82 464.166
R6218 a_n7636_8799.n172 a_n7636_8799.t34 464.166
R6219 a_n7636_8799.n182 a_n7636_8799.t88 464.166
R6220 a_n7636_8799.n181 a_n7636_8799.t86 464.166
R6221 a_n7636_8799.n173 a_n7636_8799.t36 464.166
R6222 a_n7636_8799.n180 a_n7636_8799.t35 464.166
R6223 a_n7636_8799.n179 a_n7636_8799.t104 464.166
R6224 a_n7636_8799.n174 a_n7636_8799.t48 464.166
R6225 a_n7636_8799.n178 a_n7636_8799.t39 464.166
R6226 a_n7636_8799.n177 a_n7636_8799.t108 464.166
R6227 a_n7636_8799.n175 a_n7636_8799.t70 464.166
R6228 a_n7636_8799.n202 a_n7636_8799.t81 464.166
R6229 a_n7636_8799.n201 a_n7636_8799.t61 464.166
R6230 a_n7636_8799.n187 a_n7636_8799.t127 464.166
R6231 a_n7636_8799.n200 a_n7636_8799.t97 464.166
R6232 a_n7636_8799.n199 a_n7636_8799.t96 464.166
R6233 a_n7636_8799.n188 a_n7636_8799.t42 464.166
R6234 a_n7636_8799.n198 a_n7636_8799.t100 464.166
R6235 a_n7636_8799.n197 a_n7636_8799.t98 464.166
R6236 a_n7636_8799.n189 a_n7636_8799.t44 464.166
R6237 a_n7636_8799.n196 a_n7636_8799.t43 464.166
R6238 a_n7636_8799.n195 a_n7636_8799.t119 464.166
R6239 a_n7636_8799.n190 a_n7636_8799.t59 464.166
R6240 a_n7636_8799.n194 a_n7636_8799.t45 464.166
R6241 a_n7636_8799.n193 a_n7636_8799.t120 464.166
R6242 a_n7636_8799.n191 a_n7636_8799.t80 464.166
R6243 a_n7636_8799.n219 a_n7636_8799.t103 464.166
R6244 a_n7636_8799.n218 a_n7636_8799.t49 464.166
R6245 a_n7636_8799.n204 a_n7636_8799.t87 464.166
R6246 a_n7636_8799.n217 a_n7636_8799.t37 464.166
R6247 a_n7636_8799.n216 a_n7636_8799.t56 464.166
R6248 a_n7636_8799.n205 a_n7636_8799.t123 464.166
R6249 a_n7636_8799.n215 a_n7636_8799.t95 464.166
R6250 a_n7636_8799.n214 a_n7636_8799.t117 464.166
R6251 a_n7636_8799.n206 a_n7636_8799.t78 464.166
R6252 a_n7636_8799.n213 a_n7636_8799.t99 464.166
R6253 a_n7636_8799.n212 a_n7636_8799.t46 464.166
R6254 a_n7636_8799.n207 a_n7636_8799.t114 464.166
R6255 a_n7636_8799.n211 a_n7636_8799.t64 464.166
R6256 a_n7636_8799.n210 a_n7636_8799.t109 464.166
R6257 a_n7636_8799.n208 a_n7636_8799.t54 464.166
R6258 a_n7636_8799.n124 a_n7636_8799.t113 464.166
R6259 a_n7636_8799.n127 a_n7636_8799.t69 464.166
R6260 a_n7636_8799.n123 a_n7636_8799.t94 464.166
R6261 a_n7636_8799.n128 a_n7636_8799.t110 464.166
R6262 a_n7636_8799.n129 a_n7636_8799.t67 464.166
R6263 a_n7636_8799.n130 a_n7636_8799.t68 464.166
R6264 a_n7636_8799.n131 a_n7636_8799.t91 464.166
R6265 a_n7636_8799.n122 a_n7636_8799.t58 464.166
R6266 a_n7636_8799.n132 a_n7636_8799.t57 464.166
R6267 a_n7636_8799.n133 a_n7636_8799.t89 464.166
R6268 a_n7636_8799.n134 a_n7636_8799.t32 464.166
R6269 a_n7636_8799.n135 a_n7636_8799.t55 464.166
R6270 a_n7636_8799.n121 a_n7636_8799.t73 464.166
R6271 a_n7636_8799.n136 a_n7636_8799.t111 464.166
R6272 a_n7636_8799.n140 a_n7636_8799.t125 464.166
R6273 a_n7636_8799.n143 a_n7636_8799.t77 464.166
R6274 a_n7636_8799.n139 a_n7636_8799.t106 464.166
R6275 a_n7636_8799.n144 a_n7636_8799.t122 464.166
R6276 a_n7636_8799.n145 a_n7636_8799.t76 464.166
R6277 a_n7636_8799.n146 a_n7636_8799.t75 464.166
R6278 a_n7636_8799.n147 a_n7636_8799.t105 464.166
R6279 a_n7636_8799.n138 a_n7636_8799.t63 464.166
R6280 a_n7636_8799.n148 a_n7636_8799.t66 464.166
R6281 a_n7636_8799.n149 a_n7636_8799.t101 464.166
R6282 a_n7636_8799.n150 a_n7636_8799.t40 464.166
R6283 a_n7636_8799.n151 a_n7636_8799.t62 464.166
R6284 a_n7636_8799.n137 a_n7636_8799.t84 464.166
R6285 a_n7636_8799.n152 a_n7636_8799.t124 464.166
R6286 a_n7636_8799.n157 a_n7636_8799.t72 464.166
R6287 a_n7636_8799.n160 a_n7636_8799.t107 464.166
R6288 a_n7636_8799.n156 a_n7636_8799.t65 464.166
R6289 a_n7636_8799.n161 a_n7636_8799.t115 464.166
R6290 a_n7636_8799.n162 a_n7636_8799.t47 464.166
R6291 a_n7636_8799.n163 a_n7636_8799.t33 464.166
R6292 a_n7636_8799.n164 a_n7636_8799.t79 464.166
R6293 a_n7636_8799.n155 a_n7636_8799.t118 464.166
R6294 a_n7636_8799.n165 a_n7636_8799.t93 464.166
R6295 a_n7636_8799.n166 a_n7636_8799.t121 464.166
R6296 a_n7636_8799.n167 a_n7636_8799.t74 464.166
R6297 a_n7636_8799.n168 a_n7636_8799.t38 464.166
R6298 a_n7636_8799.n154 a_n7636_8799.t85 464.166
R6299 a_n7636_8799.n169 a_n7636_8799.t50 464.166
R6300 a_n7636_8799.n51 a_n7636_8799.n33 74.4178
R6301 a_n7636_8799.n177 a_n7636_8799.n51 12.4674
R6302 a_n7636_8799.n50 a_n7636_8799.n33 80.107
R6303 a_n7636_8799.n50 a_n7636_8799.n178 1.08907
R6304 a_n7636_8799.n34 a_n7636_8799.n49 75.3623
R6305 a_n7636_8799.n48 a_n7636_8799.n34 70.3058
R6306 a_n7636_8799.n36 a_n7636_8799.n47 70.1674
R6307 a_n7636_8799.n47 a_n7636_8799.n173 20.9683
R6308 a_n7636_8799.n46 a_n7636_8799.n36 75.0448
R6309 a_n7636_8799.n181 a_n7636_8799.n46 11.2134
R6310 a_n7636_8799.n45 a_n7636_8799.n35 80.4688
R6311 a_n7636_8799.n35 a_n7636_8799.n44 74.73
R6312 a_n7636_8799.n43 a_n7636_8799.n37 70.1674
R6313 a_n7636_8799.n184 a_n7636_8799.n43 20.9683
R6314 a_n7636_8799.n37 a_n7636_8799.n42 70.5844
R6315 a_n7636_8799.n42 a_n7636_8799.n171 20.1342
R6316 a_n7636_8799.n41 a_n7636_8799.n38 75.6825
R6317 a_n7636_8799.n185 a_n7636_8799.n41 9.93802
R6318 a_n7636_8799.n38 a_n7636_8799.n186 161.3
R6319 a_n7636_8799.n62 a_n7636_8799.n27 74.4178
R6320 a_n7636_8799.n193 a_n7636_8799.n62 12.4674
R6321 a_n7636_8799.n61 a_n7636_8799.n27 80.107
R6322 a_n7636_8799.n61 a_n7636_8799.n194 1.08907
R6323 a_n7636_8799.n28 a_n7636_8799.n60 75.3623
R6324 a_n7636_8799.n59 a_n7636_8799.n28 70.3058
R6325 a_n7636_8799.n30 a_n7636_8799.n58 70.1674
R6326 a_n7636_8799.n58 a_n7636_8799.n189 20.9683
R6327 a_n7636_8799.n57 a_n7636_8799.n30 75.0448
R6328 a_n7636_8799.n197 a_n7636_8799.n57 11.2134
R6329 a_n7636_8799.n56 a_n7636_8799.n29 80.4688
R6330 a_n7636_8799.n29 a_n7636_8799.n55 74.73
R6331 a_n7636_8799.n54 a_n7636_8799.n31 70.1674
R6332 a_n7636_8799.n200 a_n7636_8799.n54 20.9683
R6333 a_n7636_8799.n31 a_n7636_8799.n53 70.5844
R6334 a_n7636_8799.n53 a_n7636_8799.n187 20.1342
R6335 a_n7636_8799.n52 a_n7636_8799.n32 75.6825
R6336 a_n7636_8799.n201 a_n7636_8799.n52 9.93802
R6337 a_n7636_8799.n32 a_n7636_8799.n202 161.3
R6338 a_n7636_8799.n73 a_n7636_8799.n21 74.4178
R6339 a_n7636_8799.n210 a_n7636_8799.n73 12.4674
R6340 a_n7636_8799.n72 a_n7636_8799.n21 80.107
R6341 a_n7636_8799.n72 a_n7636_8799.n211 1.08907
R6342 a_n7636_8799.n22 a_n7636_8799.n71 75.3623
R6343 a_n7636_8799.n70 a_n7636_8799.n22 70.3058
R6344 a_n7636_8799.n24 a_n7636_8799.n69 70.1674
R6345 a_n7636_8799.n69 a_n7636_8799.n206 20.9683
R6346 a_n7636_8799.n68 a_n7636_8799.n24 75.0448
R6347 a_n7636_8799.n214 a_n7636_8799.n68 11.2134
R6348 a_n7636_8799.n67 a_n7636_8799.n23 80.4688
R6349 a_n7636_8799.n23 a_n7636_8799.n66 74.73
R6350 a_n7636_8799.n65 a_n7636_8799.n25 70.1674
R6351 a_n7636_8799.n217 a_n7636_8799.n65 20.9683
R6352 a_n7636_8799.n25 a_n7636_8799.n64 70.5844
R6353 a_n7636_8799.n64 a_n7636_8799.n204 20.1342
R6354 a_n7636_8799.n63 a_n7636_8799.n26 75.6825
R6355 a_n7636_8799.n218 a_n7636_8799.n63 9.93802
R6356 a_n7636_8799.n26 a_n7636_8799.n219 161.3
R6357 a_n7636_8799.n16 a_n7636_8799.n84 70.1674
R6358 a_n7636_8799.n136 a_n7636_8799.n84 20.9683
R6359 a_n7636_8799.n83 a_n7636_8799.n16 74.4178
R6360 a_n7636_8799.n83 a_n7636_8799.n121 12.4674
R6361 a_n7636_8799.n15 a_n7636_8799.n82 80.107
R6362 a_n7636_8799.n135 a_n7636_8799.n82 1.08907
R6363 a_n7636_8799.n81 a_n7636_8799.n15 75.3623
R6364 a_n7636_8799.n17 a_n7636_8799.n80 70.3058
R6365 a_n7636_8799.n79 a_n7636_8799.n17 70.1674
R6366 a_n7636_8799.n79 a_n7636_8799.n122 20.9683
R6367 a_n7636_8799.n18 a_n7636_8799.n78 75.0448
R6368 a_n7636_8799.n131 a_n7636_8799.n78 11.2134
R6369 a_n7636_8799.n77 a_n7636_8799.n18 80.4688
R6370 a_n7636_8799.n19 a_n7636_8799.n76 74.73
R6371 a_n7636_8799.n75 a_n7636_8799.n19 70.1674
R6372 a_n7636_8799.n75 a_n7636_8799.n123 20.9683
R6373 a_n7636_8799.n20 a_n7636_8799.n74 70.5844
R6374 a_n7636_8799.n127 a_n7636_8799.n74 20.1342
R6375 a_n7636_8799.n126 a_n7636_8799.n20 161.3
R6376 a_n7636_8799.n10 a_n7636_8799.n95 70.1674
R6377 a_n7636_8799.n152 a_n7636_8799.n95 20.9683
R6378 a_n7636_8799.n94 a_n7636_8799.n10 74.4178
R6379 a_n7636_8799.n94 a_n7636_8799.n137 12.4674
R6380 a_n7636_8799.n9 a_n7636_8799.n93 80.107
R6381 a_n7636_8799.n151 a_n7636_8799.n93 1.08907
R6382 a_n7636_8799.n92 a_n7636_8799.n9 75.3623
R6383 a_n7636_8799.n11 a_n7636_8799.n91 70.3058
R6384 a_n7636_8799.n90 a_n7636_8799.n11 70.1674
R6385 a_n7636_8799.n90 a_n7636_8799.n138 20.9683
R6386 a_n7636_8799.n12 a_n7636_8799.n89 75.0448
R6387 a_n7636_8799.n147 a_n7636_8799.n89 11.2134
R6388 a_n7636_8799.n88 a_n7636_8799.n12 80.4688
R6389 a_n7636_8799.n13 a_n7636_8799.n87 74.73
R6390 a_n7636_8799.n86 a_n7636_8799.n13 70.1674
R6391 a_n7636_8799.n86 a_n7636_8799.n139 20.9683
R6392 a_n7636_8799.n14 a_n7636_8799.n85 70.5844
R6393 a_n7636_8799.n143 a_n7636_8799.n85 20.1342
R6394 a_n7636_8799.n142 a_n7636_8799.n14 161.3
R6395 a_n7636_8799.n4 a_n7636_8799.n106 70.1674
R6396 a_n7636_8799.n169 a_n7636_8799.n106 20.9683
R6397 a_n7636_8799.n105 a_n7636_8799.n4 74.4178
R6398 a_n7636_8799.n105 a_n7636_8799.n154 12.4674
R6399 a_n7636_8799.n3 a_n7636_8799.n104 80.107
R6400 a_n7636_8799.n168 a_n7636_8799.n104 1.08907
R6401 a_n7636_8799.n103 a_n7636_8799.n3 75.3623
R6402 a_n7636_8799.n5 a_n7636_8799.n102 70.3058
R6403 a_n7636_8799.n101 a_n7636_8799.n5 70.1674
R6404 a_n7636_8799.n101 a_n7636_8799.n155 20.9683
R6405 a_n7636_8799.n6 a_n7636_8799.n100 75.0448
R6406 a_n7636_8799.n164 a_n7636_8799.n100 11.2134
R6407 a_n7636_8799.n99 a_n7636_8799.n6 80.4688
R6408 a_n7636_8799.n7 a_n7636_8799.n98 74.73
R6409 a_n7636_8799.n97 a_n7636_8799.n7 70.1674
R6410 a_n7636_8799.n97 a_n7636_8799.n156 20.9683
R6411 a_n7636_8799.n8 a_n7636_8799.n96 70.5844
R6412 a_n7636_8799.n160 a_n7636_8799.n96 20.1342
R6413 a_n7636_8799.n159 a_n7636_8799.n8 161.3
R6414 a_n7636_8799.n226 a_n7636_8799.n107 98.9633
R6415 a_n7636_8799.n39 a_n7636_8799.n108 98.9631
R6416 a_n7636_8799.n40 a_n7636_8799.n224 98.6055
R6417 a_n7636_8799.n40 a_n7636_8799.n225 98.6055
R6418 a_n7636_8799.n39 a_n7636_8799.n109 98.6055
R6419 a_n7636_8799.n39 a_n7636_8799.n110 98.6055
R6420 a_n7636_8799.n112 a_n7636_8799.n111 98.6055
R6421 a_n7636_8799.n227 a_n7636_8799.n226 98.6054
R6422 a_n7636_8799.n1 a_n7636_8799.n113 81.4626
R6423 a_n7636_8799.n2 a_n7636_8799.n117 81.4626
R6424 a_n7636_8799.n2 a_n7636_8799.n115 81.4626
R6425 a_n7636_8799.n0 a_n7636_8799.n119 80.9324
R6426 a_n7636_8799.n1 a_n7636_8799.n120 80.9324
R6427 a_n7636_8799.n1 a_n7636_8799.n114 80.9324
R6428 a_n7636_8799.n2 a_n7636_8799.n118 80.9324
R6429 a_n7636_8799.n2 a_n7636_8799.n116 80.9324
R6430 a_n7636_8799.n33 a_n7636_8799.n176 70.4033
R6431 a_n7636_8799.n27 a_n7636_8799.n192 70.4033
R6432 a_n7636_8799.n21 a_n7636_8799.n209 70.4033
R6433 a_n7636_8799.n20 a_n7636_8799.n125 70.4033
R6434 a_n7636_8799.n14 a_n7636_8799.n141 70.4033
R6435 a_n7636_8799.n8 a_n7636_8799.n158 70.4033
R6436 a_n7636_8799.n186 a_n7636_8799.n185 48.2005
R6437 a_n7636_8799.n43 a_n7636_8799.n183 20.9683
R6438 a_n7636_8799.n182 a_n7636_8799.n181 48.2005
R6439 a_n7636_8799.n180 a_n7636_8799.n47 20.9683
R6440 a_n7636_8799.n178 a_n7636_8799.n174 48.2005
R6441 a_n7636_8799.n202 a_n7636_8799.n201 48.2005
R6442 a_n7636_8799.n54 a_n7636_8799.n199 20.9683
R6443 a_n7636_8799.n198 a_n7636_8799.n197 48.2005
R6444 a_n7636_8799.n196 a_n7636_8799.n58 20.9683
R6445 a_n7636_8799.n194 a_n7636_8799.n190 48.2005
R6446 a_n7636_8799.n219 a_n7636_8799.n218 48.2005
R6447 a_n7636_8799.n65 a_n7636_8799.n216 20.9683
R6448 a_n7636_8799.n215 a_n7636_8799.n214 48.2005
R6449 a_n7636_8799.n213 a_n7636_8799.n69 20.9683
R6450 a_n7636_8799.n211 a_n7636_8799.n207 48.2005
R6451 a_n7636_8799.n128 a_n7636_8799.n75 20.9683
R6452 a_n7636_8799.n131 a_n7636_8799.n130 48.2005
R6453 a_n7636_8799.n132 a_n7636_8799.n79 20.9683
R6454 a_n7636_8799.n135 a_n7636_8799.n134 48.2005
R6455 a_n7636_8799.t41 a_n7636_8799.n84 485.135
R6456 a_n7636_8799.n144 a_n7636_8799.n86 20.9683
R6457 a_n7636_8799.n147 a_n7636_8799.n146 48.2005
R6458 a_n7636_8799.n148 a_n7636_8799.n90 20.9683
R6459 a_n7636_8799.n151 a_n7636_8799.n150 48.2005
R6460 a_n7636_8799.t53 a_n7636_8799.n95 485.135
R6461 a_n7636_8799.n161 a_n7636_8799.n97 20.9683
R6462 a_n7636_8799.n164 a_n7636_8799.n163 48.2005
R6463 a_n7636_8799.n165 a_n7636_8799.n101 20.9683
R6464 a_n7636_8799.n168 a_n7636_8799.n167 48.2005
R6465 a_n7636_8799.t102 a_n7636_8799.n106 485.135
R6466 a_n7636_8799.n45 a_n7636_8799.n172 47.835
R6467 a_n7636_8799.n48 a_n7636_8799.n179 20.6913
R6468 a_n7636_8799.n56 a_n7636_8799.n188 47.835
R6469 a_n7636_8799.n59 a_n7636_8799.n195 20.6913
R6470 a_n7636_8799.n67 a_n7636_8799.n205 47.835
R6471 a_n7636_8799.n70 a_n7636_8799.n212 20.6913
R6472 a_n7636_8799.n129 a_n7636_8799.n77 47.835
R6473 a_n7636_8799.n133 a_n7636_8799.n80 20.6913
R6474 a_n7636_8799.n145 a_n7636_8799.n88 47.835
R6475 a_n7636_8799.n149 a_n7636_8799.n91 20.6913
R6476 a_n7636_8799.n162 a_n7636_8799.n99 47.835
R6477 a_n7636_8799.n166 a_n7636_8799.n102 20.6913
R6478 a_n7636_8799.n184 a_n7636_8799.n42 22.3251
R6479 a_n7636_8799.n200 a_n7636_8799.n53 22.3251
R6480 a_n7636_8799.n217 a_n7636_8799.n64 22.3251
R6481 a_n7636_8799.n123 a_n7636_8799.n74 22.3251
R6482 a_n7636_8799.n139 a_n7636_8799.n85 22.3251
R6483 a_n7636_8799.n156 a_n7636_8799.n96 22.3251
R6484 a_n7636_8799.n223 a_n7636_8799.n112 31.7372
R6485 a_n7636_8799.n51 a_n7636_8799.n175 33.6462
R6486 a_n7636_8799.n62 a_n7636_8799.n191 33.6462
R6487 a_n7636_8799.n73 a_n7636_8799.n208 33.6462
R6488 a_n7636_8799.n127 a_n7636_8799.n126 27.0217
R6489 a_n7636_8799.n136 a_n7636_8799.n83 33.6462
R6490 a_n7636_8799.n143 a_n7636_8799.n142 27.0217
R6491 a_n7636_8799.n152 a_n7636_8799.n94 33.6462
R6492 a_n7636_8799.n160 a_n7636_8799.n159 27.0217
R6493 a_n7636_8799.n169 a_n7636_8799.n105 33.6462
R6494 a_n7636_8799.n44 a_n7636_8799.n172 11.843
R6495 a_n7636_8799.n179 a_n7636_8799.n49 36.139
R6496 a_n7636_8799.n55 a_n7636_8799.n188 11.843
R6497 a_n7636_8799.n195 a_n7636_8799.n60 36.139
R6498 a_n7636_8799.n66 a_n7636_8799.n205 11.843
R6499 a_n7636_8799.n212 a_n7636_8799.n71 36.139
R6500 a_n7636_8799.n129 a_n7636_8799.n76 11.843
R6501 a_n7636_8799.n133 a_n7636_8799.n81 36.139
R6502 a_n7636_8799.n145 a_n7636_8799.n87 11.843
R6503 a_n7636_8799.n149 a_n7636_8799.n92 36.139
R6504 a_n7636_8799.n162 a_n7636_8799.n98 11.843
R6505 a_n7636_8799.n166 a_n7636_8799.n103 36.139
R6506 a_n7636_8799.n46 a_n7636_8799.n173 35.3134
R6507 a_n7636_8799.n57 a_n7636_8799.n189 35.3134
R6508 a_n7636_8799.n68 a_n7636_8799.n206 35.3134
R6509 a_n7636_8799.n122 a_n7636_8799.n78 35.3134
R6510 a_n7636_8799.n138 a_n7636_8799.n89 35.3134
R6511 a_n7636_8799.n155 a_n7636_8799.n100 35.3134
R6512 a_n7636_8799.n183 a_n7636_8799.n44 34.4824
R6513 a_n7636_8799.n49 a_n7636_8799.n174 10.5784
R6514 a_n7636_8799.n199 a_n7636_8799.n55 34.4824
R6515 a_n7636_8799.n60 a_n7636_8799.n190 10.5784
R6516 a_n7636_8799.n216 a_n7636_8799.n66 34.4824
R6517 a_n7636_8799.n71 a_n7636_8799.n207 10.5784
R6518 a_n7636_8799.n76 a_n7636_8799.n128 34.4824
R6519 a_n7636_8799.n134 a_n7636_8799.n81 10.5784
R6520 a_n7636_8799.n87 a_n7636_8799.n144 34.4824
R6521 a_n7636_8799.n150 a_n7636_8799.n92 10.5784
R6522 a_n7636_8799.n98 a_n7636_8799.n161 34.4824
R6523 a_n7636_8799.n167 a_n7636_8799.n103 10.5784
R6524 a_n7636_8799.n41 a_n7636_8799.n171 36.9592
R6525 a_n7636_8799.n52 a_n7636_8799.n187 36.9592
R6526 a_n7636_8799.n63 a_n7636_8799.n204 36.9592
R6527 a_n7636_8799.n126 a_n7636_8799.n124 21.1793
R6528 a_n7636_8799.n142 a_n7636_8799.n140 21.1793
R6529 a_n7636_8799.n159 a_n7636_8799.n157 21.1793
R6530 a_n7636_8799.n176 a_n7636_8799.n175 20.9576
R6531 a_n7636_8799.n192 a_n7636_8799.n191 20.9576
R6532 a_n7636_8799.n209 a_n7636_8799.n208 20.9576
R6533 a_n7636_8799.n125 a_n7636_8799.n124 20.9576
R6534 a_n7636_8799.n141 a_n7636_8799.n140 20.9576
R6535 a_n7636_8799.n158 a_n7636_8799.n157 20.9576
R6536 a_n7636_8799.n40 a_n7636_8799.n223 18.8589
R6537 a_n7636_8799.n222 a_n7636_8799.n1 12.3339
R6538 a_n7636_8799.n223 a_n7636_8799.n222 11.4887
R6539 a_n7636_8799.n203 a_n7636_8799.n38 9.07815
R6540 a_n7636_8799.n153 a_n7636_8799.n16 9.07815
R6541 a_n7636_8799.n221 a_n7636_8799.n170 6.96667
R6542 a_n7636_8799.n221 a_n7636_8799.n220 6.62419
R6543 a_n7636_8799.n203 a_n7636_8799.n32 4.9702
R6544 a_n7636_8799.n220 a_n7636_8799.n26 4.9702
R6545 a_n7636_8799.n153 a_n7636_8799.n10 4.9702
R6546 a_n7636_8799.n170 a_n7636_8799.n4 4.9702
R6547 a_n7636_8799.n220 a_n7636_8799.n203 4.10845
R6548 a_n7636_8799.n170 a_n7636_8799.n153 4.10845
R6549 a_n7636_8799.n224 a_n7636_8799.t14 3.61217
R6550 a_n7636_8799.n224 a_n7636_8799.t17 3.61217
R6551 a_n7636_8799.n225 a_n7636_8799.t16 3.61217
R6552 a_n7636_8799.n225 a_n7636_8799.t21 3.61217
R6553 a_n7636_8799.n107 a_n7636_8799.t13 3.61217
R6554 a_n7636_8799.n107 a_n7636_8799.t20 3.61217
R6555 a_n7636_8799.n108 a_n7636_8799.t15 3.61217
R6556 a_n7636_8799.n108 a_n7636_8799.t8 3.61217
R6557 a_n7636_8799.n109 a_n7636_8799.t12 3.61217
R6558 a_n7636_8799.n109 a_n7636_8799.t18 3.61217
R6559 a_n7636_8799.n110 a_n7636_8799.t9 3.61217
R6560 a_n7636_8799.n110 a_n7636_8799.t11 3.61217
R6561 a_n7636_8799.n111 a_n7636_8799.t7 3.61217
R6562 a_n7636_8799.n111 a_n7636_8799.t10 3.61217
R6563 a_n7636_8799.t6 a_n7636_8799.n227 3.61217
R6564 a_n7636_8799.n227 a_n7636_8799.t19 3.61217
R6565 a_n7636_8799.n222 a_n7636_8799.n221 3.4105
R6566 a_n7636_8799.n119 a_n7636_8799.t4 2.82907
R6567 a_n7636_8799.n119 a_n7636_8799.t30 2.82907
R6568 a_n7636_8799.n120 a_n7636_8799.t1 2.82907
R6569 a_n7636_8799.n120 a_n7636_8799.t27 2.82907
R6570 a_n7636_8799.n114 a_n7636_8799.t29 2.82907
R6571 a_n7636_8799.n114 a_n7636_8799.t3 2.82907
R6572 a_n7636_8799.n113 a_n7636_8799.t23 2.82907
R6573 a_n7636_8799.n113 a_n7636_8799.t5 2.82907
R6574 a_n7636_8799.n117 a_n7636_8799.t24 2.82907
R6575 a_n7636_8799.n117 a_n7636_8799.t25 2.82907
R6576 a_n7636_8799.n118 a_n7636_8799.t0 2.82907
R6577 a_n7636_8799.n118 a_n7636_8799.t28 2.82907
R6578 a_n7636_8799.n116 a_n7636_8799.t31 2.82907
R6579 a_n7636_8799.n116 a_n7636_8799.t26 2.82907
R6580 a_n7636_8799.n115 a_n7636_8799.t2 2.82907
R6581 a_n7636_8799.n115 a_n7636_8799.t22 2.82907
R6582 a_n7636_8799.n50 a_n7636_8799.n177 47.0982
R6583 a_n7636_8799.n61 a_n7636_8799.n193 47.0982
R6584 a_n7636_8799.n72 a_n7636_8799.n210 47.0982
R6585 a_n7636_8799.n121 a_n7636_8799.n82 47.0982
R6586 a_n7636_8799.n137 a_n7636_8799.n93 47.0982
R6587 a_n7636_8799.n154 a_n7636_8799.n104 47.0982
R6588 a_n7636_8799.n0 a_n7636_8799.n2 33.2634
R6589 a_n7636_8799.n45 a_n7636_8799.n182 0.365327
R6590 a_n7636_8799.n180 a_n7636_8799.n48 21.4216
R6591 a_n7636_8799.n56 a_n7636_8799.n198 0.365327
R6592 a_n7636_8799.n196 a_n7636_8799.n59 21.4216
R6593 a_n7636_8799.n67 a_n7636_8799.n215 0.365327
R6594 a_n7636_8799.n213 a_n7636_8799.n70 21.4216
R6595 a_n7636_8799.n130 a_n7636_8799.n77 0.365327
R6596 a_n7636_8799.n80 a_n7636_8799.n132 21.4216
R6597 a_n7636_8799.n146 a_n7636_8799.n88 0.365327
R6598 a_n7636_8799.n91 a_n7636_8799.n148 21.4216
R6599 a_n7636_8799.n163 a_n7636_8799.n99 0.365327
R6600 a_n7636_8799.n102 a_n7636_8799.n165 21.4216
R6601 a_n7636_8799.n34 a_n7636_8799.n33 1.13686
R6602 a_n7636_8799.n28 a_n7636_8799.n27 1.13686
R6603 a_n7636_8799.n22 a_n7636_8799.n21 1.13686
R6604 a_n7636_8799.n16 a_n7636_8799.n15 1.13686
R6605 a_n7636_8799.n10 a_n7636_8799.n9 1.13686
R6606 a_n7636_8799.n4 a_n7636_8799.n3 1.13686
R6607 a_n7636_8799.n1 a_n7636_8799.n0 1.06084
R6608 a_n7636_8799.n38 a_n7636_8799.n37 0.758076
R6609 a_n7636_8799.n35 a_n7636_8799.n37 0.758076
R6610 a_n7636_8799.n36 a_n7636_8799.n35 0.758076
R6611 a_n7636_8799.n36 a_n7636_8799.n34 0.758076
R6612 a_n7636_8799.n32 a_n7636_8799.n31 0.758076
R6613 a_n7636_8799.n29 a_n7636_8799.n31 0.758076
R6614 a_n7636_8799.n30 a_n7636_8799.n29 0.758076
R6615 a_n7636_8799.n30 a_n7636_8799.n28 0.758076
R6616 a_n7636_8799.n26 a_n7636_8799.n25 0.758076
R6617 a_n7636_8799.n23 a_n7636_8799.n25 0.758076
R6618 a_n7636_8799.n24 a_n7636_8799.n23 0.758076
R6619 a_n7636_8799.n24 a_n7636_8799.n22 0.758076
R6620 a_n7636_8799.n19 a_n7636_8799.n20 0.758076
R6621 a_n7636_8799.n18 a_n7636_8799.n19 0.758076
R6622 a_n7636_8799.n17 a_n7636_8799.n18 0.758076
R6623 a_n7636_8799.n15 a_n7636_8799.n17 0.758076
R6624 a_n7636_8799.n13 a_n7636_8799.n14 0.758076
R6625 a_n7636_8799.n12 a_n7636_8799.n13 0.758076
R6626 a_n7636_8799.n11 a_n7636_8799.n12 0.758076
R6627 a_n7636_8799.n9 a_n7636_8799.n11 0.758076
R6628 a_n7636_8799.n7 a_n7636_8799.n8 0.758076
R6629 a_n7636_8799.n6 a_n7636_8799.n7 0.758076
R6630 a_n7636_8799.n5 a_n7636_8799.n6 0.758076
R6631 a_n7636_8799.n3 a_n7636_8799.n5 0.758076
R6632 a_n7636_8799.n226 a_n7636_8799.n40 0.716017
R6633 a_n7636_8799.n112 a_n7636_8799.n39 0.716017
R6634 CSoutput.n19 CSoutput.t145 184.661
R6635 CSoutput.n78 CSoutput.n77 165.8
R6636 CSoutput.n76 CSoutput.n0 165.8
R6637 CSoutput.n75 CSoutput.n74 165.8
R6638 CSoutput.n73 CSoutput.n72 165.8
R6639 CSoutput.n71 CSoutput.n2 165.8
R6640 CSoutput.n69 CSoutput.n68 165.8
R6641 CSoutput.n67 CSoutput.n3 165.8
R6642 CSoutput.n66 CSoutput.n65 165.8
R6643 CSoutput.n63 CSoutput.n4 165.8
R6644 CSoutput.n61 CSoutput.n60 165.8
R6645 CSoutput.n59 CSoutput.n5 165.8
R6646 CSoutput.n58 CSoutput.n57 165.8
R6647 CSoutput.n55 CSoutput.n6 165.8
R6648 CSoutput.n54 CSoutput.n53 165.8
R6649 CSoutput.n52 CSoutput.n51 165.8
R6650 CSoutput.n50 CSoutput.n8 165.8
R6651 CSoutput.n48 CSoutput.n47 165.8
R6652 CSoutput.n46 CSoutput.n9 165.8
R6653 CSoutput.n45 CSoutput.n44 165.8
R6654 CSoutput.n42 CSoutput.n10 165.8
R6655 CSoutput.n41 CSoutput.n40 165.8
R6656 CSoutput.n39 CSoutput.n38 165.8
R6657 CSoutput.n37 CSoutput.n12 165.8
R6658 CSoutput.n35 CSoutput.n34 165.8
R6659 CSoutput.n33 CSoutput.n13 165.8
R6660 CSoutput.n32 CSoutput.n31 165.8
R6661 CSoutput.n29 CSoutput.n14 165.8
R6662 CSoutput.n28 CSoutput.n27 165.8
R6663 CSoutput.n26 CSoutput.n25 165.8
R6664 CSoutput.n24 CSoutput.n16 165.8
R6665 CSoutput.n22 CSoutput.n21 165.8
R6666 CSoutput.n20 CSoutput.n17 165.8
R6667 CSoutput.n77 CSoutput.t148 162.194
R6668 CSoutput.n18 CSoutput.t147 120.501
R6669 CSoutput.n23 CSoutput.t158 120.501
R6670 CSoutput.n15 CSoutput.t155 120.501
R6671 CSoutput.n30 CSoutput.t149 120.501
R6672 CSoutput.n36 CSoutput.t160 120.501
R6673 CSoutput.n11 CSoutput.t162 120.501
R6674 CSoutput.n43 CSoutput.t151 120.501
R6675 CSoutput.n49 CSoutput.t163 120.501
R6676 CSoutput.n7 CSoutput.t165 120.501
R6677 CSoutput.n56 CSoutput.t159 120.501
R6678 CSoutput.n62 CSoutput.t150 120.501
R6679 CSoutput.n64 CSoutput.t144 120.501
R6680 CSoutput.n70 CSoutput.t161 120.501
R6681 CSoutput.n1 CSoutput.t156 120.501
R6682 CSoutput.n310 CSoutput.n308 103.469
R6683 CSoutput.n294 CSoutput.n292 103.469
R6684 CSoutput.n279 CSoutput.n277 103.469
R6685 CSoutput.n112 CSoutput.n110 103.469
R6686 CSoutput.n96 CSoutput.n94 103.469
R6687 CSoutput.n81 CSoutput.n79 103.469
R6688 CSoutput.n320 CSoutput.n319 103.111
R6689 CSoutput.n318 CSoutput.n317 103.111
R6690 CSoutput.n316 CSoutput.n315 103.111
R6691 CSoutput.n314 CSoutput.n313 103.111
R6692 CSoutput.n312 CSoutput.n311 103.111
R6693 CSoutput.n310 CSoutput.n309 103.111
R6694 CSoutput.n306 CSoutput.n305 103.111
R6695 CSoutput.n304 CSoutput.n303 103.111
R6696 CSoutput.n302 CSoutput.n301 103.111
R6697 CSoutput.n300 CSoutput.n299 103.111
R6698 CSoutput.n298 CSoutput.n297 103.111
R6699 CSoutput.n296 CSoutput.n295 103.111
R6700 CSoutput.n294 CSoutput.n293 103.111
R6701 CSoutput.n291 CSoutput.n290 103.111
R6702 CSoutput.n289 CSoutput.n288 103.111
R6703 CSoutput.n287 CSoutput.n286 103.111
R6704 CSoutput.n285 CSoutput.n284 103.111
R6705 CSoutput.n283 CSoutput.n282 103.111
R6706 CSoutput.n281 CSoutput.n280 103.111
R6707 CSoutput.n279 CSoutput.n278 103.111
R6708 CSoutput.n112 CSoutput.n111 103.111
R6709 CSoutput.n114 CSoutput.n113 103.111
R6710 CSoutput.n116 CSoutput.n115 103.111
R6711 CSoutput.n118 CSoutput.n117 103.111
R6712 CSoutput.n120 CSoutput.n119 103.111
R6713 CSoutput.n122 CSoutput.n121 103.111
R6714 CSoutput.n124 CSoutput.n123 103.111
R6715 CSoutput.n96 CSoutput.n95 103.111
R6716 CSoutput.n98 CSoutput.n97 103.111
R6717 CSoutput.n100 CSoutput.n99 103.111
R6718 CSoutput.n102 CSoutput.n101 103.111
R6719 CSoutput.n104 CSoutput.n103 103.111
R6720 CSoutput.n106 CSoutput.n105 103.111
R6721 CSoutput.n108 CSoutput.n107 103.111
R6722 CSoutput.n81 CSoutput.n80 103.111
R6723 CSoutput.n83 CSoutput.n82 103.111
R6724 CSoutput.n85 CSoutput.n84 103.111
R6725 CSoutput.n87 CSoutput.n86 103.111
R6726 CSoutput.n89 CSoutput.n88 103.111
R6727 CSoutput.n91 CSoutput.n90 103.111
R6728 CSoutput.n93 CSoutput.n92 103.111
R6729 CSoutput.n322 CSoutput.n321 103.111
R6730 CSoutput.n338 CSoutput.n336 81.5057
R6731 CSoutput.n327 CSoutput.n325 81.5057
R6732 CSoutput.n362 CSoutput.n360 81.5057
R6733 CSoutput.n351 CSoutput.n349 81.5057
R6734 CSoutput.n346 CSoutput.n345 80.9324
R6735 CSoutput.n344 CSoutput.n343 80.9324
R6736 CSoutput.n342 CSoutput.n341 80.9324
R6737 CSoutput.n340 CSoutput.n339 80.9324
R6738 CSoutput.n338 CSoutput.n337 80.9324
R6739 CSoutput.n335 CSoutput.n334 80.9324
R6740 CSoutput.n333 CSoutput.n332 80.9324
R6741 CSoutput.n331 CSoutput.n330 80.9324
R6742 CSoutput.n329 CSoutput.n328 80.9324
R6743 CSoutput.n327 CSoutput.n326 80.9324
R6744 CSoutput.n362 CSoutput.n361 80.9324
R6745 CSoutput.n364 CSoutput.n363 80.9324
R6746 CSoutput.n366 CSoutput.n365 80.9324
R6747 CSoutput.n368 CSoutput.n367 80.9324
R6748 CSoutput.n370 CSoutput.n369 80.9324
R6749 CSoutput.n351 CSoutput.n350 80.9324
R6750 CSoutput.n353 CSoutput.n352 80.9324
R6751 CSoutput.n355 CSoutput.n354 80.9324
R6752 CSoutput.n357 CSoutput.n356 80.9324
R6753 CSoutput.n359 CSoutput.n358 80.9324
R6754 CSoutput.n25 CSoutput.n24 48.1486
R6755 CSoutput.n69 CSoutput.n3 48.1486
R6756 CSoutput.n38 CSoutput.n37 48.1486
R6757 CSoutput.n42 CSoutput.n41 48.1486
R6758 CSoutput.n51 CSoutput.n50 48.1486
R6759 CSoutput.n55 CSoutput.n54 48.1486
R6760 CSoutput.n22 CSoutput.n17 46.462
R6761 CSoutput.n72 CSoutput.n71 46.462
R6762 CSoutput.n20 CSoutput.n19 44.9055
R6763 CSoutput.n29 CSoutput.n28 43.7635
R6764 CSoutput.n65 CSoutput.n63 43.7635
R6765 CSoutput.n35 CSoutput.n13 41.7396
R6766 CSoutput.n57 CSoutput.n5 41.7396
R6767 CSoutput.n44 CSoutput.n9 37.0171
R6768 CSoutput.n48 CSoutput.n9 37.0171
R6769 CSoutput.n76 CSoutput.n75 34.9932
R6770 CSoutput.n31 CSoutput.n13 32.2947
R6771 CSoutput.n61 CSoutput.n5 32.2947
R6772 CSoutput.n30 CSoutput.n29 29.6014
R6773 CSoutput.n63 CSoutput.n62 29.6014
R6774 CSoutput.n19 CSoutput.n18 28.4085
R6775 CSoutput.n18 CSoutput.n17 25.1176
R6776 CSoutput.n72 CSoutput.n1 25.1176
R6777 CSoutput.n43 CSoutput.n42 22.0922
R6778 CSoutput.n50 CSoutput.n49 22.0922
R6779 CSoutput.n77 CSoutput.n76 21.8586
R6780 CSoutput.n37 CSoutput.n36 18.9681
R6781 CSoutput.n56 CSoutput.n55 18.9681
R6782 CSoutput.n25 CSoutput.n15 17.6292
R6783 CSoutput.n64 CSoutput.n3 17.6292
R6784 CSoutput.n24 CSoutput.n23 15.844
R6785 CSoutput.n70 CSoutput.n69 15.844
R6786 CSoutput.n38 CSoutput.n11 14.5051
R6787 CSoutput.n54 CSoutput.n7 14.5051
R6788 CSoutput.n373 CSoutput.n78 11.6139
R6789 CSoutput.n41 CSoutput.n11 11.3811
R6790 CSoutput.n51 CSoutput.n7 11.3811
R6791 CSoutput.n23 CSoutput.n22 10.0422
R6792 CSoutput.n71 CSoutput.n70 10.0422
R6793 CSoutput.n307 CSoutput.n291 9.25285
R6794 CSoutput.n109 CSoutput.n93 9.25285
R6795 CSoutput.n347 CSoutput.n335 8.97993
R6796 CSoutput.n371 CSoutput.n359 8.97993
R6797 CSoutput.n348 CSoutput.n324 8.61621
R6798 CSoutput.n28 CSoutput.n15 8.25698
R6799 CSoutput.n65 CSoutput.n64 8.25698
R6800 CSoutput.n348 CSoutput.n347 7.89345
R6801 CSoutput.n372 CSoutput.n371 7.89345
R6802 CSoutput.n324 CSoutput.n323 7.12641
R6803 CSoutput.n126 CSoutput.n125 7.12641
R6804 CSoutput.n36 CSoutput.n35 6.91809
R6805 CSoutput.n57 CSoutput.n56 6.91809
R6806 CSoutput.n347 CSoutput.n346 5.25266
R6807 CSoutput.n371 CSoutput.n370 5.25266
R6808 CSoutput.n323 CSoutput.n322 5.1449
R6809 CSoutput.n307 CSoutput.n306 5.1449
R6810 CSoutput.n125 CSoutput.n124 5.1449
R6811 CSoutput.n109 CSoutput.n108 5.1449
R6812 CSoutput.n373 CSoutput.n126 5.02377
R6813 CSoutput.n217 CSoutput.n170 4.5005
R6814 CSoutput.n186 CSoutput.n170 4.5005
R6815 CSoutput.n181 CSoutput.n165 4.5005
R6816 CSoutput.n181 CSoutput.n167 4.5005
R6817 CSoutput.n181 CSoutput.n164 4.5005
R6818 CSoutput.n181 CSoutput.n168 4.5005
R6819 CSoutput.n181 CSoutput.n163 4.5005
R6820 CSoutput.n181 CSoutput.t152 4.5005
R6821 CSoutput.n181 CSoutput.n162 4.5005
R6822 CSoutput.n181 CSoutput.n169 4.5005
R6823 CSoutput.n181 CSoutput.n170 4.5005
R6824 CSoutput.n179 CSoutput.n165 4.5005
R6825 CSoutput.n179 CSoutput.n167 4.5005
R6826 CSoutput.n179 CSoutput.n164 4.5005
R6827 CSoutput.n179 CSoutput.n168 4.5005
R6828 CSoutput.n179 CSoutput.n163 4.5005
R6829 CSoutput.n179 CSoutput.t152 4.5005
R6830 CSoutput.n179 CSoutput.n162 4.5005
R6831 CSoutput.n179 CSoutput.n169 4.5005
R6832 CSoutput.n179 CSoutput.n170 4.5005
R6833 CSoutput.n178 CSoutput.n165 4.5005
R6834 CSoutput.n178 CSoutput.n167 4.5005
R6835 CSoutput.n178 CSoutput.n164 4.5005
R6836 CSoutput.n178 CSoutput.n168 4.5005
R6837 CSoutput.n178 CSoutput.n163 4.5005
R6838 CSoutput.n178 CSoutput.t152 4.5005
R6839 CSoutput.n178 CSoutput.n162 4.5005
R6840 CSoutput.n178 CSoutput.n169 4.5005
R6841 CSoutput.n178 CSoutput.n170 4.5005
R6842 CSoutput.n263 CSoutput.n165 4.5005
R6843 CSoutput.n263 CSoutput.n167 4.5005
R6844 CSoutput.n263 CSoutput.n164 4.5005
R6845 CSoutput.n263 CSoutput.n168 4.5005
R6846 CSoutput.n263 CSoutput.n163 4.5005
R6847 CSoutput.n263 CSoutput.t152 4.5005
R6848 CSoutput.n263 CSoutput.n162 4.5005
R6849 CSoutput.n263 CSoutput.n169 4.5005
R6850 CSoutput.n263 CSoutput.n170 4.5005
R6851 CSoutput.n261 CSoutput.n165 4.5005
R6852 CSoutput.n261 CSoutput.n167 4.5005
R6853 CSoutput.n261 CSoutput.n164 4.5005
R6854 CSoutput.n261 CSoutput.n168 4.5005
R6855 CSoutput.n261 CSoutput.n163 4.5005
R6856 CSoutput.n261 CSoutput.t152 4.5005
R6857 CSoutput.n261 CSoutput.n162 4.5005
R6858 CSoutput.n261 CSoutput.n169 4.5005
R6859 CSoutput.n259 CSoutput.n165 4.5005
R6860 CSoutput.n259 CSoutput.n167 4.5005
R6861 CSoutput.n259 CSoutput.n164 4.5005
R6862 CSoutput.n259 CSoutput.n168 4.5005
R6863 CSoutput.n259 CSoutput.n163 4.5005
R6864 CSoutput.n259 CSoutput.t152 4.5005
R6865 CSoutput.n259 CSoutput.n162 4.5005
R6866 CSoutput.n259 CSoutput.n169 4.5005
R6867 CSoutput.n189 CSoutput.n165 4.5005
R6868 CSoutput.n189 CSoutput.n167 4.5005
R6869 CSoutput.n189 CSoutput.n164 4.5005
R6870 CSoutput.n189 CSoutput.n168 4.5005
R6871 CSoutput.n189 CSoutput.n163 4.5005
R6872 CSoutput.n189 CSoutput.t152 4.5005
R6873 CSoutput.n189 CSoutput.n162 4.5005
R6874 CSoutput.n189 CSoutput.n169 4.5005
R6875 CSoutput.n189 CSoutput.n170 4.5005
R6876 CSoutput.n188 CSoutput.n165 4.5005
R6877 CSoutput.n188 CSoutput.n167 4.5005
R6878 CSoutput.n188 CSoutput.n164 4.5005
R6879 CSoutput.n188 CSoutput.n168 4.5005
R6880 CSoutput.n188 CSoutput.n163 4.5005
R6881 CSoutput.n188 CSoutput.t152 4.5005
R6882 CSoutput.n188 CSoutput.n162 4.5005
R6883 CSoutput.n188 CSoutput.n169 4.5005
R6884 CSoutput.n188 CSoutput.n170 4.5005
R6885 CSoutput.n192 CSoutput.n165 4.5005
R6886 CSoutput.n192 CSoutput.n167 4.5005
R6887 CSoutput.n192 CSoutput.n164 4.5005
R6888 CSoutput.n192 CSoutput.n168 4.5005
R6889 CSoutput.n192 CSoutput.n163 4.5005
R6890 CSoutput.n192 CSoutput.t152 4.5005
R6891 CSoutput.n192 CSoutput.n162 4.5005
R6892 CSoutput.n192 CSoutput.n169 4.5005
R6893 CSoutput.n192 CSoutput.n170 4.5005
R6894 CSoutput.n191 CSoutput.n165 4.5005
R6895 CSoutput.n191 CSoutput.n167 4.5005
R6896 CSoutput.n191 CSoutput.n164 4.5005
R6897 CSoutput.n191 CSoutput.n168 4.5005
R6898 CSoutput.n191 CSoutput.n163 4.5005
R6899 CSoutput.n191 CSoutput.t152 4.5005
R6900 CSoutput.n191 CSoutput.n162 4.5005
R6901 CSoutput.n191 CSoutput.n169 4.5005
R6902 CSoutput.n191 CSoutput.n170 4.5005
R6903 CSoutput.n174 CSoutput.n165 4.5005
R6904 CSoutput.n174 CSoutput.n167 4.5005
R6905 CSoutput.n174 CSoutput.n164 4.5005
R6906 CSoutput.n174 CSoutput.n168 4.5005
R6907 CSoutput.n174 CSoutput.n163 4.5005
R6908 CSoutput.n174 CSoutput.t152 4.5005
R6909 CSoutput.n174 CSoutput.n162 4.5005
R6910 CSoutput.n174 CSoutput.n169 4.5005
R6911 CSoutput.n174 CSoutput.n170 4.5005
R6912 CSoutput.n266 CSoutput.n165 4.5005
R6913 CSoutput.n266 CSoutput.n167 4.5005
R6914 CSoutput.n266 CSoutput.n164 4.5005
R6915 CSoutput.n266 CSoutput.n168 4.5005
R6916 CSoutput.n266 CSoutput.n163 4.5005
R6917 CSoutput.n266 CSoutput.t152 4.5005
R6918 CSoutput.n266 CSoutput.n162 4.5005
R6919 CSoutput.n266 CSoutput.n169 4.5005
R6920 CSoutput.n266 CSoutput.n170 4.5005
R6921 CSoutput.n253 CSoutput.n224 4.5005
R6922 CSoutput.n253 CSoutput.n230 4.5005
R6923 CSoutput.n211 CSoutput.n200 4.5005
R6924 CSoutput.n211 CSoutput.n202 4.5005
R6925 CSoutput.n211 CSoutput.n199 4.5005
R6926 CSoutput.n211 CSoutput.n203 4.5005
R6927 CSoutput.n211 CSoutput.n198 4.5005
R6928 CSoutput.n211 CSoutput.t146 4.5005
R6929 CSoutput.n211 CSoutput.n197 4.5005
R6930 CSoutput.n211 CSoutput.n204 4.5005
R6931 CSoutput.n253 CSoutput.n211 4.5005
R6932 CSoutput.n232 CSoutput.n200 4.5005
R6933 CSoutput.n232 CSoutput.n202 4.5005
R6934 CSoutput.n232 CSoutput.n199 4.5005
R6935 CSoutput.n232 CSoutput.n203 4.5005
R6936 CSoutput.n232 CSoutput.n198 4.5005
R6937 CSoutput.n232 CSoutput.t146 4.5005
R6938 CSoutput.n232 CSoutput.n197 4.5005
R6939 CSoutput.n232 CSoutput.n204 4.5005
R6940 CSoutput.n253 CSoutput.n232 4.5005
R6941 CSoutput.n210 CSoutput.n200 4.5005
R6942 CSoutput.n210 CSoutput.n202 4.5005
R6943 CSoutput.n210 CSoutput.n199 4.5005
R6944 CSoutput.n210 CSoutput.n203 4.5005
R6945 CSoutput.n210 CSoutput.n198 4.5005
R6946 CSoutput.n210 CSoutput.t146 4.5005
R6947 CSoutput.n210 CSoutput.n197 4.5005
R6948 CSoutput.n210 CSoutput.n204 4.5005
R6949 CSoutput.n253 CSoutput.n210 4.5005
R6950 CSoutput.n234 CSoutput.n200 4.5005
R6951 CSoutput.n234 CSoutput.n202 4.5005
R6952 CSoutput.n234 CSoutput.n199 4.5005
R6953 CSoutput.n234 CSoutput.n203 4.5005
R6954 CSoutput.n234 CSoutput.n198 4.5005
R6955 CSoutput.n234 CSoutput.t146 4.5005
R6956 CSoutput.n234 CSoutput.n197 4.5005
R6957 CSoutput.n234 CSoutput.n204 4.5005
R6958 CSoutput.n253 CSoutput.n234 4.5005
R6959 CSoutput.n200 CSoutput.n195 4.5005
R6960 CSoutput.n202 CSoutput.n195 4.5005
R6961 CSoutput.n199 CSoutput.n195 4.5005
R6962 CSoutput.n203 CSoutput.n195 4.5005
R6963 CSoutput.n198 CSoutput.n195 4.5005
R6964 CSoutput.t146 CSoutput.n195 4.5005
R6965 CSoutput.n197 CSoutput.n195 4.5005
R6966 CSoutput.n204 CSoutput.n195 4.5005
R6967 CSoutput.n256 CSoutput.n200 4.5005
R6968 CSoutput.n256 CSoutput.n202 4.5005
R6969 CSoutput.n256 CSoutput.n199 4.5005
R6970 CSoutput.n256 CSoutput.n203 4.5005
R6971 CSoutput.n256 CSoutput.n198 4.5005
R6972 CSoutput.n256 CSoutput.t146 4.5005
R6973 CSoutput.n256 CSoutput.n197 4.5005
R6974 CSoutput.n256 CSoutput.n204 4.5005
R6975 CSoutput.n254 CSoutput.n200 4.5005
R6976 CSoutput.n254 CSoutput.n202 4.5005
R6977 CSoutput.n254 CSoutput.n199 4.5005
R6978 CSoutput.n254 CSoutput.n203 4.5005
R6979 CSoutput.n254 CSoutput.n198 4.5005
R6980 CSoutput.n254 CSoutput.t146 4.5005
R6981 CSoutput.n254 CSoutput.n197 4.5005
R6982 CSoutput.n254 CSoutput.n204 4.5005
R6983 CSoutput.n254 CSoutput.n253 4.5005
R6984 CSoutput.n236 CSoutput.n200 4.5005
R6985 CSoutput.n236 CSoutput.n202 4.5005
R6986 CSoutput.n236 CSoutput.n199 4.5005
R6987 CSoutput.n236 CSoutput.n203 4.5005
R6988 CSoutput.n236 CSoutput.n198 4.5005
R6989 CSoutput.n236 CSoutput.t146 4.5005
R6990 CSoutput.n236 CSoutput.n197 4.5005
R6991 CSoutput.n236 CSoutput.n204 4.5005
R6992 CSoutput.n253 CSoutput.n236 4.5005
R6993 CSoutput.n208 CSoutput.n200 4.5005
R6994 CSoutput.n208 CSoutput.n202 4.5005
R6995 CSoutput.n208 CSoutput.n199 4.5005
R6996 CSoutput.n208 CSoutput.n203 4.5005
R6997 CSoutput.n208 CSoutput.n198 4.5005
R6998 CSoutput.n208 CSoutput.t146 4.5005
R6999 CSoutput.n208 CSoutput.n197 4.5005
R7000 CSoutput.n208 CSoutput.n204 4.5005
R7001 CSoutput.n253 CSoutput.n208 4.5005
R7002 CSoutput.n238 CSoutput.n200 4.5005
R7003 CSoutput.n238 CSoutput.n202 4.5005
R7004 CSoutput.n238 CSoutput.n199 4.5005
R7005 CSoutput.n238 CSoutput.n203 4.5005
R7006 CSoutput.n238 CSoutput.n198 4.5005
R7007 CSoutput.n238 CSoutput.t146 4.5005
R7008 CSoutput.n238 CSoutput.n197 4.5005
R7009 CSoutput.n238 CSoutput.n204 4.5005
R7010 CSoutput.n253 CSoutput.n238 4.5005
R7011 CSoutput.n207 CSoutput.n200 4.5005
R7012 CSoutput.n207 CSoutput.n202 4.5005
R7013 CSoutput.n207 CSoutput.n199 4.5005
R7014 CSoutput.n207 CSoutput.n203 4.5005
R7015 CSoutput.n207 CSoutput.n198 4.5005
R7016 CSoutput.n207 CSoutput.t146 4.5005
R7017 CSoutput.n207 CSoutput.n197 4.5005
R7018 CSoutput.n207 CSoutput.n204 4.5005
R7019 CSoutput.n253 CSoutput.n207 4.5005
R7020 CSoutput.n252 CSoutput.n200 4.5005
R7021 CSoutput.n252 CSoutput.n202 4.5005
R7022 CSoutput.n252 CSoutput.n199 4.5005
R7023 CSoutput.n252 CSoutput.n203 4.5005
R7024 CSoutput.n252 CSoutput.n198 4.5005
R7025 CSoutput.n252 CSoutput.t146 4.5005
R7026 CSoutput.n252 CSoutput.n197 4.5005
R7027 CSoutput.n252 CSoutput.n204 4.5005
R7028 CSoutput.n253 CSoutput.n252 4.5005
R7029 CSoutput.n251 CSoutput.n136 4.5005
R7030 CSoutput.n152 CSoutput.n136 4.5005
R7031 CSoutput.n147 CSoutput.n131 4.5005
R7032 CSoutput.n147 CSoutput.n133 4.5005
R7033 CSoutput.n147 CSoutput.n130 4.5005
R7034 CSoutput.n147 CSoutput.n134 4.5005
R7035 CSoutput.n147 CSoutput.n129 4.5005
R7036 CSoutput.n147 CSoutput.t164 4.5005
R7037 CSoutput.n147 CSoutput.n128 4.5005
R7038 CSoutput.n147 CSoutput.n135 4.5005
R7039 CSoutput.n147 CSoutput.n136 4.5005
R7040 CSoutput.n145 CSoutput.n131 4.5005
R7041 CSoutput.n145 CSoutput.n133 4.5005
R7042 CSoutput.n145 CSoutput.n130 4.5005
R7043 CSoutput.n145 CSoutput.n134 4.5005
R7044 CSoutput.n145 CSoutput.n129 4.5005
R7045 CSoutput.n145 CSoutput.t164 4.5005
R7046 CSoutput.n145 CSoutput.n128 4.5005
R7047 CSoutput.n145 CSoutput.n135 4.5005
R7048 CSoutput.n145 CSoutput.n136 4.5005
R7049 CSoutput.n144 CSoutput.n131 4.5005
R7050 CSoutput.n144 CSoutput.n133 4.5005
R7051 CSoutput.n144 CSoutput.n130 4.5005
R7052 CSoutput.n144 CSoutput.n134 4.5005
R7053 CSoutput.n144 CSoutput.n129 4.5005
R7054 CSoutput.n144 CSoutput.t164 4.5005
R7055 CSoutput.n144 CSoutput.n128 4.5005
R7056 CSoutput.n144 CSoutput.n135 4.5005
R7057 CSoutput.n144 CSoutput.n136 4.5005
R7058 CSoutput.n273 CSoutput.n131 4.5005
R7059 CSoutput.n273 CSoutput.n133 4.5005
R7060 CSoutput.n273 CSoutput.n130 4.5005
R7061 CSoutput.n273 CSoutput.n134 4.5005
R7062 CSoutput.n273 CSoutput.n129 4.5005
R7063 CSoutput.n273 CSoutput.t164 4.5005
R7064 CSoutput.n273 CSoutput.n128 4.5005
R7065 CSoutput.n273 CSoutput.n135 4.5005
R7066 CSoutput.n273 CSoutput.n136 4.5005
R7067 CSoutput.n271 CSoutput.n131 4.5005
R7068 CSoutput.n271 CSoutput.n133 4.5005
R7069 CSoutput.n271 CSoutput.n130 4.5005
R7070 CSoutput.n271 CSoutput.n134 4.5005
R7071 CSoutput.n271 CSoutput.n129 4.5005
R7072 CSoutput.n271 CSoutput.t164 4.5005
R7073 CSoutput.n271 CSoutput.n128 4.5005
R7074 CSoutput.n271 CSoutput.n135 4.5005
R7075 CSoutput.n269 CSoutput.n131 4.5005
R7076 CSoutput.n269 CSoutput.n133 4.5005
R7077 CSoutput.n269 CSoutput.n130 4.5005
R7078 CSoutput.n269 CSoutput.n134 4.5005
R7079 CSoutput.n269 CSoutput.n129 4.5005
R7080 CSoutput.n269 CSoutput.t164 4.5005
R7081 CSoutput.n269 CSoutput.n128 4.5005
R7082 CSoutput.n269 CSoutput.n135 4.5005
R7083 CSoutput.n155 CSoutput.n131 4.5005
R7084 CSoutput.n155 CSoutput.n133 4.5005
R7085 CSoutput.n155 CSoutput.n130 4.5005
R7086 CSoutput.n155 CSoutput.n134 4.5005
R7087 CSoutput.n155 CSoutput.n129 4.5005
R7088 CSoutput.n155 CSoutput.t164 4.5005
R7089 CSoutput.n155 CSoutput.n128 4.5005
R7090 CSoutput.n155 CSoutput.n135 4.5005
R7091 CSoutput.n155 CSoutput.n136 4.5005
R7092 CSoutput.n154 CSoutput.n131 4.5005
R7093 CSoutput.n154 CSoutput.n133 4.5005
R7094 CSoutput.n154 CSoutput.n130 4.5005
R7095 CSoutput.n154 CSoutput.n134 4.5005
R7096 CSoutput.n154 CSoutput.n129 4.5005
R7097 CSoutput.n154 CSoutput.t164 4.5005
R7098 CSoutput.n154 CSoutput.n128 4.5005
R7099 CSoutput.n154 CSoutput.n135 4.5005
R7100 CSoutput.n154 CSoutput.n136 4.5005
R7101 CSoutput.n158 CSoutput.n131 4.5005
R7102 CSoutput.n158 CSoutput.n133 4.5005
R7103 CSoutput.n158 CSoutput.n130 4.5005
R7104 CSoutput.n158 CSoutput.n134 4.5005
R7105 CSoutput.n158 CSoutput.n129 4.5005
R7106 CSoutput.n158 CSoutput.t164 4.5005
R7107 CSoutput.n158 CSoutput.n128 4.5005
R7108 CSoutput.n158 CSoutput.n135 4.5005
R7109 CSoutput.n158 CSoutput.n136 4.5005
R7110 CSoutput.n157 CSoutput.n131 4.5005
R7111 CSoutput.n157 CSoutput.n133 4.5005
R7112 CSoutput.n157 CSoutput.n130 4.5005
R7113 CSoutput.n157 CSoutput.n134 4.5005
R7114 CSoutput.n157 CSoutput.n129 4.5005
R7115 CSoutput.n157 CSoutput.t164 4.5005
R7116 CSoutput.n157 CSoutput.n128 4.5005
R7117 CSoutput.n157 CSoutput.n135 4.5005
R7118 CSoutput.n157 CSoutput.n136 4.5005
R7119 CSoutput.n140 CSoutput.n131 4.5005
R7120 CSoutput.n140 CSoutput.n133 4.5005
R7121 CSoutput.n140 CSoutput.n130 4.5005
R7122 CSoutput.n140 CSoutput.n134 4.5005
R7123 CSoutput.n140 CSoutput.n129 4.5005
R7124 CSoutput.n140 CSoutput.t164 4.5005
R7125 CSoutput.n140 CSoutput.n128 4.5005
R7126 CSoutput.n140 CSoutput.n135 4.5005
R7127 CSoutput.n140 CSoutput.n136 4.5005
R7128 CSoutput.n276 CSoutput.n131 4.5005
R7129 CSoutput.n276 CSoutput.n133 4.5005
R7130 CSoutput.n276 CSoutput.n130 4.5005
R7131 CSoutput.n276 CSoutput.n134 4.5005
R7132 CSoutput.n276 CSoutput.n129 4.5005
R7133 CSoutput.n276 CSoutput.t164 4.5005
R7134 CSoutput.n276 CSoutput.n128 4.5005
R7135 CSoutput.n276 CSoutput.n135 4.5005
R7136 CSoutput.n276 CSoutput.n136 4.5005
R7137 CSoutput.n323 CSoutput.n307 4.10845
R7138 CSoutput.n125 CSoutput.n109 4.10845
R7139 CSoutput.n321 CSoutput.t73 4.06363
R7140 CSoutput.n321 CSoutput.t92 4.06363
R7141 CSoutput.n319 CSoutput.t104 4.06363
R7142 CSoutput.n319 CSoutput.t35 4.06363
R7143 CSoutput.n317 CSoutput.t39 4.06363
R7144 CSoutput.n317 CSoutput.t95 4.06363
R7145 CSoutput.n315 CSoutput.t107 4.06363
R7146 CSoutput.n315 CSoutput.t108 4.06363
R7147 CSoutput.n313 CSoutput.t55 4.06363
R7148 CSoutput.n313 CSoutput.t57 4.06363
R7149 CSoutput.n311 CSoutput.t61 4.06363
R7150 CSoutput.n311 CSoutput.t109 4.06363
R7151 CSoutput.n309 CSoutput.t27 4.06363
R7152 CSoutput.n309 CSoutput.t60 4.06363
R7153 CSoutput.n308 CSoutput.t72 4.06363
R7154 CSoutput.n308 CSoutput.t91 4.06363
R7155 CSoutput.n305 CSoutput.t63 4.06363
R7156 CSoutput.n305 CSoutput.t83 4.06363
R7157 CSoutput.n303 CSoutput.t98 4.06363
R7158 CSoutput.n303 CSoutput.t23 4.06363
R7159 CSoutput.n301 CSoutput.t24 4.06363
R7160 CSoutput.n301 CSoutput.t84 4.06363
R7161 CSoutput.n299 CSoutput.t99 4.06363
R7162 CSoutput.n299 CSoutput.t100 4.06363
R7163 CSoutput.n297 CSoutput.t43 4.06363
R7164 CSoutput.n297 CSoutput.t45 4.06363
R7165 CSoutput.n295 CSoutput.t47 4.06363
R7166 CSoutput.n295 CSoutput.t101 4.06363
R7167 CSoutput.n293 CSoutput.t16 4.06363
R7168 CSoutput.n293 CSoutput.t46 4.06363
R7169 CSoutput.n292 CSoutput.t62 4.06363
R7170 CSoutput.n292 CSoutput.t82 4.06363
R7171 CSoutput.n290 CSoutput.t89 4.06363
R7172 CSoutput.n290 CSoutput.t51 4.06363
R7173 CSoutput.n288 CSoutput.t79 4.06363
R7174 CSoutput.n288 CSoutput.t34 4.06363
R7175 CSoutput.n286 CSoutput.t97 4.06363
R7176 CSoutput.n286 CSoutput.t29 4.06363
R7177 CSoutput.n284 CSoutput.t65 4.06363
R7178 CSoutput.n284 CSoutput.t44 4.06363
R7179 CSoutput.n282 CSoutput.t48 4.06363
R7180 CSoutput.n282 CSoutput.t26 4.06363
R7181 CSoutput.n280 CSoutput.t87 4.06363
R7182 CSoutput.n280 CSoutput.t20 4.06363
R7183 CSoutput.n278 CSoutput.t56 4.06363
R7184 CSoutput.n278 CSoutput.t106 4.06363
R7185 CSoutput.n277 CSoutput.t40 4.06363
R7186 CSoutput.n277 CSoutput.t94 4.06363
R7187 CSoutput.n110 CSoutput.t32 4.06363
R7188 CSoutput.n110 CSoutput.t102 4.06363
R7189 CSoutput.n111 CSoutput.t88 4.06363
R7190 CSoutput.n111 CSoutput.t70 4.06363
R7191 CSoutput.n113 CSoutput.t54 4.06363
R7192 CSoutput.n113 CSoutput.t111 4.06363
R7193 CSoutput.n115 CSoutput.t85 4.06363
R7194 CSoutput.n115 CSoutput.t86 4.06363
R7195 CSoutput.n117 CSoutput.t75 4.06363
R7196 CSoutput.n117 CSoutput.t52 4.06363
R7197 CSoutput.n119 CSoutput.t33 4.06363
R7198 CSoutput.n119 CSoutput.t76 4.06363
R7199 CSoutput.n121 CSoutput.t74 4.06363
R7200 CSoutput.n121 CSoutput.t49 4.06363
R7201 CSoutput.n123 CSoutput.t31 4.06363
R7202 CSoutput.n123 CSoutput.t30 4.06363
R7203 CSoutput.n94 CSoutput.t19 4.06363
R7204 CSoutput.n94 CSoutput.t90 4.06363
R7205 CSoutput.n95 CSoutput.t81 4.06363
R7206 CSoutput.n95 CSoutput.t59 4.06363
R7207 CSoutput.n97 CSoutput.t42 4.06363
R7208 CSoutput.n97 CSoutput.t103 4.06363
R7209 CSoutput.n99 CSoutput.t80 4.06363
R7210 CSoutput.n99 CSoutput.t77 4.06363
R7211 CSoutput.n101 CSoutput.t68 4.06363
R7212 CSoutput.n101 CSoutput.t38 4.06363
R7213 CSoutput.n103 CSoutput.t21 4.06363
R7214 CSoutput.n103 CSoutput.t67 4.06363
R7215 CSoutput.n105 CSoutput.t66 4.06363
R7216 CSoutput.n105 CSoutput.t37 4.06363
R7217 CSoutput.n107 CSoutput.t17 4.06363
R7218 CSoutput.n107 CSoutput.t18 4.06363
R7219 CSoutput.n79 CSoutput.t93 4.06363
R7220 CSoutput.n79 CSoutput.t41 4.06363
R7221 CSoutput.n80 CSoutput.t105 4.06363
R7222 CSoutput.n80 CSoutput.t58 4.06363
R7223 CSoutput.n82 CSoutput.t22 4.06363
R7224 CSoutput.n82 CSoutput.t69 4.06363
R7225 CSoutput.n84 CSoutput.t25 4.06363
R7226 CSoutput.n84 CSoutput.t50 4.06363
R7227 CSoutput.n86 CSoutput.t110 4.06363
R7228 CSoutput.n86 CSoutput.t64 4.06363
R7229 CSoutput.n88 CSoutput.t28 4.06363
R7230 CSoutput.n88 CSoutput.t96 4.06363
R7231 CSoutput.n90 CSoutput.t36 4.06363
R7232 CSoutput.n90 CSoutput.t78 4.06363
R7233 CSoutput.n92 CSoutput.t53 4.06363
R7234 CSoutput.n92 CSoutput.t71 4.06363
R7235 CSoutput.n44 CSoutput.n43 3.79402
R7236 CSoutput.n49 CSoutput.n48 3.79402
R7237 CSoutput.n373 CSoutput.n372 3.57343
R7238 CSoutput.n345 CSoutput.t129 2.82907
R7239 CSoutput.n345 CSoutput.t132 2.82907
R7240 CSoutput.n343 CSoutput.t134 2.82907
R7241 CSoutput.n343 CSoutput.t139 2.82907
R7242 CSoutput.n341 CSoutput.t2 2.82907
R7243 CSoutput.n341 CSoutput.t6 2.82907
R7244 CSoutput.n339 CSoutput.t120 2.82907
R7245 CSoutput.n339 CSoutput.t142 2.82907
R7246 CSoutput.n337 CSoutput.t14 2.82907
R7247 CSoutput.n337 CSoutput.t8 2.82907
R7248 CSoutput.n336 CSoutput.t137 2.82907
R7249 CSoutput.n336 CSoutput.t9 2.82907
R7250 CSoutput.n334 CSoutput.t13 2.82907
R7251 CSoutput.n334 CSoutput.t117 2.82907
R7252 CSoutput.n332 CSoutput.t114 2.82907
R7253 CSoutput.n332 CSoutput.t141 2.82907
R7254 CSoutput.n330 CSoutput.t116 2.82907
R7255 CSoutput.n330 CSoutput.t135 2.82907
R7256 CSoutput.n328 CSoutput.t121 2.82907
R7257 CSoutput.n328 CSoutput.t113 2.82907
R7258 CSoutput.n326 CSoutput.t130 2.82907
R7259 CSoutput.n326 CSoutput.t131 2.82907
R7260 CSoutput.n325 CSoutput.t122 2.82907
R7261 CSoutput.n325 CSoutput.t128 2.82907
R7262 CSoutput.n360 CSoutput.t10 2.82907
R7263 CSoutput.n360 CSoutput.t138 2.82907
R7264 CSoutput.n361 CSoutput.t1 2.82907
R7265 CSoutput.n361 CSoutput.t3 2.82907
R7266 CSoutput.n363 CSoutput.t7 2.82907
R7267 CSoutput.n363 CSoutput.t119 2.82907
R7268 CSoutput.n365 CSoutput.t143 2.82907
R7269 CSoutput.n365 CSoutput.t4 2.82907
R7270 CSoutput.n367 CSoutput.t0 2.82907
R7271 CSoutput.n367 CSoutput.t112 2.82907
R7272 CSoutput.n369 CSoutput.t15 2.82907
R7273 CSoutput.n369 CSoutput.t126 2.82907
R7274 CSoutput.n349 CSoutput.t133 2.82907
R7275 CSoutput.n349 CSoutput.t11 2.82907
R7276 CSoutput.n350 CSoutput.t115 2.82907
R7277 CSoutput.n350 CSoutput.t118 2.82907
R7278 CSoutput.n352 CSoutput.t136 2.82907
R7279 CSoutput.n352 CSoutput.t140 2.82907
R7280 CSoutput.n354 CSoutput.t127 2.82907
R7281 CSoutput.n354 CSoutput.t5 2.82907
R7282 CSoutput.n356 CSoutput.t124 2.82907
R7283 CSoutput.n356 CSoutput.t125 2.82907
R7284 CSoutput.n358 CSoutput.t123 2.82907
R7285 CSoutput.n358 CSoutput.t12 2.82907
R7286 CSoutput.n372 CSoutput.n348 2.75627
R7287 CSoutput.n324 CSoutput.n126 2.57547
R7288 CSoutput.n75 CSoutput.n1 2.45513
R7289 CSoutput.n217 CSoutput.n215 2.251
R7290 CSoutput.n217 CSoutput.n214 2.251
R7291 CSoutput.n217 CSoutput.n213 2.251
R7292 CSoutput.n217 CSoutput.n212 2.251
R7293 CSoutput.n186 CSoutput.n185 2.251
R7294 CSoutput.n186 CSoutput.n184 2.251
R7295 CSoutput.n186 CSoutput.n183 2.251
R7296 CSoutput.n186 CSoutput.n182 2.251
R7297 CSoutput.n259 CSoutput.n258 2.251
R7298 CSoutput.n224 CSoutput.n222 2.251
R7299 CSoutput.n224 CSoutput.n221 2.251
R7300 CSoutput.n224 CSoutput.n220 2.251
R7301 CSoutput.n242 CSoutput.n224 2.251
R7302 CSoutput.n230 CSoutput.n229 2.251
R7303 CSoutput.n230 CSoutput.n228 2.251
R7304 CSoutput.n230 CSoutput.n227 2.251
R7305 CSoutput.n230 CSoutput.n226 2.251
R7306 CSoutput.n256 CSoutput.n196 2.251
R7307 CSoutput.n251 CSoutput.n249 2.251
R7308 CSoutput.n251 CSoutput.n248 2.251
R7309 CSoutput.n251 CSoutput.n247 2.251
R7310 CSoutput.n251 CSoutput.n246 2.251
R7311 CSoutput.n152 CSoutput.n151 2.251
R7312 CSoutput.n152 CSoutput.n150 2.251
R7313 CSoutput.n152 CSoutput.n149 2.251
R7314 CSoutput.n152 CSoutput.n148 2.251
R7315 CSoutput.n269 CSoutput.n268 2.251
R7316 CSoutput.n186 CSoutput.n166 2.2505
R7317 CSoutput.n181 CSoutput.n166 2.2505
R7318 CSoutput.n179 CSoutput.n166 2.2505
R7319 CSoutput.n178 CSoutput.n166 2.2505
R7320 CSoutput.n263 CSoutput.n166 2.2505
R7321 CSoutput.n261 CSoutput.n166 2.2505
R7322 CSoutput.n259 CSoutput.n166 2.2505
R7323 CSoutput.n189 CSoutput.n166 2.2505
R7324 CSoutput.n188 CSoutput.n166 2.2505
R7325 CSoutput.n192 CSoutput.n166 2.2505
R7326 CSoutput.n191 CSoutput.n166 2.2505
R7327 CSoutput.n174 CSoutput.n166 2.2505
R7328 CSoutput.n266 CSoutput.n166 2.2505
R7329 CSoutput.n266 CSoutput.n265 2.2505
R7330 CSoutput.n230 CSoutput.n201 2.2505
R7331 CSoutput.n211 CSoutput.n201 2.2505
R7332 CSoutput.n232 CSoutput.n201 2.2505
R7333 CSoutput.n210 CSoutput.n201 2.2505
R7334 CSoutput.n234 CSoutput.n201 2.2505
R7335 CSoutput.n201 CSoutput.n195 2.2505
R7336 CSoutput.n256 CSoutput.n201 2.2505
R7337 CSoutput.n254 CSoutput.n201 2.2505
R7338 CSoutput.n236 CSoutput.n201 2.2505
R7339 CSoutput.n208 CSoutput.n201 2.2505
R7340 CSoutput.n238 CSoutput.n201 2.2505
R7341 CSoutput.n207 CSoutput.n201 2.2505
R7342 CSoutput.n252 CSoutput.n201 2.2505
R7343 CSoutput.n252 CSoutput.n205 2.2505
R7344 CSoutput.n152 CSoutput.n132 2.2505
R7345 CSoutput.n147 CSoutput.n132 2.2505
R7346 CSoutput.n145 CSoutput.n132 2.2505
R7347 CSoutput.n144 CSoutput.n132 2.2505
R7348 CSoutput.n273 CSoutput.n132 2.2505
R7349 CSoutput.n271 CSoutput.n132 2.2505
R7350 CSoutput.n269 CSoutput.n132 2.2505
R7351 CSoutput.n155 CSoutput.n132 2.2505
R7352 CSoutput.n154 CSoutput.n132 2.2505
R7353 CSoutput.n158 CSoutput.n132 2.2505
R7354 CSoutput.n157 CSoutput.n132 2.2505
R7355 CSoutput.n140 CSoutput.n132 2.2505
R7356 CSoutput.n276 CSoutput.n132 2.2505
R7357 CSoutput.n276 CSoutput.n275 2.2505
R7358 CSoutput.n194 CSoutput.n187 2.25024
R7359 CSoutput.n194 CSoutput.n180 2.25024
R7360 CSoutput.n262 CSoutput.n194 2.25024
R7361 CSoutput.n194 CSoutput.n190 2.25024
R7362 CSoutput.n194 CSoutput.n193 2.25024
R7363 CSoutput.n194 CSoutput.n161 2.25024
R7364 CSoutput.n244 CSoutput.n241 2.25024
R7365 CSoutput.n244 CSoutput.n240 2.25024
R7366 CSoutput.n244 CSoutput.n239 2.25024
R7367 CSoutput.n244 CSoutput.n206 2.25024
R7368 CSoutput.n244 CSoutput.n243 2.25024
R7369 CSoutput.n245 CSoutput.n244 2.25024
R7370 CSoutput.n160 CSoutput.n153 2.25024
R7371 CSoutput.n160 CSoutput.n146 2.25024
R7372 CSoutput.n272 CSoutput.n160 2.25024
R7373 CSoutput.n160 CSoutput.n156 2.25024
R7374 CSoutput.n160 CSoutput.n159 2.25024
R7375 CSoutput.n160 CSoutput.n127 2.25024
R7376 CSoutput.n261 CSoutput.n171 1.50111
R7377 CSoutput.n209 CSoutput.n195 1.50111
R7378 CSoutput.n271 CSoutput.n137 1.50111
R7379 CSoutput.n217 CSoutput.n216 1.501
R7380 CSoutput.n224 CSoutput.n223 1.501
R7381 CSoutput.n251 CSoutput.n250 1.501
R7382 CSoutput.n265 CSoutput.n176 1.12536
R7383 CSoutput.n265 CSoutput.n177 1.12536
R7384 CSoutput.n265 CSoutput.n264 1.12536
R7385 CSoutput.n225 CSoutput.n205 1.12536
R7386 CSoutput.n231 CSoutput.n205 1.12536
R7387 CSoutput.n233 CSoutput.n205 1.12536
R7388 CSoutput.n275 CSoutput.n142 1.12536
R7389 CSoutput.n275 CSoutput.n143 1.12536
R7390 CSoutput.n275 CSoutput.n274 1.12536
R7391 CSoutput.n265 CSoutput.n172 1.12536
R7392 CSoutput.n265 CSoutput.n173 1.12536
R7393 CSoutput.n265 CSoutput.n175 1.12536
R7394 CSoutput.n255 CSoutput.n205 1.12536
R7395 CSoutput.n235 CSoutput.n205 1.12536
R7396 CSoutput.n237 CSoutput.n205 1.12536
R7397 CSoutput.n275 CSoutput.n138 1.12536
R7398 CSoutput.n275 CSoutput.n139 1.12536
R7399 CSoutput.n275 CSoutput.n141 1.12536
R7400 CSoutput.n31 CSoutput.n30 0.669944
R7401 CSoutput.n62 CSoutput.n61 0.669944
R7402 CSoutput.n340 CSoutput.n338 0.573776
R7403 CSoutput.n342 CSoutput.n340 0.573776
R7404 CSoutput.n344 CSoutput.n342 0.573776
R7405 CSoutput.n346 CSoutput.n344 0.573776
R7406 CSoutput.n329 CSoutput.n327 0.573776
R7407 CSoutput.n331 CSoutput.n329 0.573776
R7408 CSoutput.n333 CSoutput.n331 0.573776
R7409 CSoutput.n335 CSoutput.n333 0.573776
R7410 CSoutput.n370 CSoutput.n368 0.573776
R7411 CSoutput.n368 CSoutput.n366 0.573776
R7412 CSoutput.n366 CSoutput.n364 0.573776
R7413 CSoutput.n364 CSoutput.n362 0.573776
R7414 CSoutput.n359 CSoutput.n357 0.573776
R7415 CSoutput.n357 CSoutput.n355 0.573776
R7416 CSoutput.n355 CSoutput.n353 0.573776
R7417 CSoutput.n353 CSoutput.n351 0.573776
R7418 CSoutput.n373 CSoutput.n276 0.53442
R7419 CSoutput.n312 CSoutput.n310 0.358259
R7420 CSoutput.n314 CSoutput.n312 0.358259
R7421 CSoutput.n316 CSoutput.n314 0.358259
R7422 CSoutput.n318 CSoutput.n316 0.358259
R7423 CSoutput.n320 CSoutput.n318 0.358259
R7424 CSoutput.n322 CSoutput.n320 0.358259
R7425 CSoutput.n296 CSoutput.n294 0.358259
R7426 CSoutput.n298 CSoutput.n296 0.358259
R7427 CSoutput.n300 CSoutput.n298 0.358259
R7428 CSoutput.n302 CSoutput.n300 0.358259
R7429 CSoutput.n304 CSoutput.n302 0.358259
R7430 CSoutput.n306 CSoutput.n304 0.358259
R7431 CSoutput.n281 CSoutput.n279 0.358259
R7432 CSoutput.n283 CSoutput.n281 0.358259
R7433 CSoutput.n285 CSoutput.n283 0.358259
R7434 CSoutput.n287 CSoutput.n285 0.358259
R7435 CSoutput.n289 CSoutput.n287 0.358259
R7436 CSoutput.n291 CSoutput.n289 0.358259
R7437 CSoutput.n124 CSoutput.n122 0.358259
R7438 CSoutput.n122 CSoutput.n120 0.358259
R7439 CSoutput.n120 CSoutput.n118 0.358259
R7440 CSoutput.n118 CSoutput.n116 0.358259
R7441 CSoutput.n116 CSoutput.n114 0.358259
R7442 CSoutput.n114 CSoutput.n112 0.358259
R7443 CSoutput.n108 CSoutput.n106 0.358259
R7444 CSoutput.n106 CSoutput.n104 0.358259
R7445 CSoutput.n104 CSoutput.n102 0.358259
R7446 CSoutput.n102 CSoutput.n100 0.358259
R7447 CSoutput.n100 CSoutput.n98 0.358259
R7448 CSoutput.n98 CSoutput.n96 0.358259
R7449 CSoutput.n93 CSoutput.n91 0.358259
R7450 CSoutput.n91 CSoutput.n89 0.358259
R7451 CSoutput.n89 CSoutput.n87 0.358259
R7452 CSoutput.n87 CSoutput.n85 0.358259
R7453 CSoutput.n85 CSoutput.n83 0.358259
R7454 CSoutput.n83 CSoutput.n81 0.358259
R7455 CSoutput.n21 CSoutput.n20 0.169105
R7456 CSoutput.n21 CSoutput.n16 0.169105
R7457 CSoutput.n26 CSoutput.n16 0.169105
R7458 CSoutput.n27 CSoutput.n26 0.169105
R7459 CSoutput.n27 CSoutput.n14 0.169105
R7460 CSoutput.n32 CSoutput.n14 0.169105
R7461 CSoutput.n33 CSoutput.n32 0.169105
R7462 CSoutput.n34 CSoutput.n33 0.169105
R7463 CSoutput.n34 CSoutput.n12 0.169105
R7464 CSoutput.n39 CSoutput.n12 0.169105
R7465 CSoutput.n40 CSoutput.n39 0.169105
R7466 CSoutput.n40 CSoutput.n10 0.169105
R7467 CSoutput.n45 CSoutput.n10 0.169105
R7468 CSoutput.n46 CSoutput.n45 0.169105
R7469 CSoutput.n47 CSoutput.n46 0.169105
R7470 CSoutput.n47 CSoutput.n8 0.169105
R7471 CSoutput.n52 CSoutput.n8 0.169105
R7472 CSoutput.n53 CSoutput.n52 0.169105
R7473 CSoutput.n53 CSoutput.n6 0.169105
R7474 CSoutput.n58 CSoutput.n6 0.169105
R7475 CSoutput.n59 CSoutput.n58 0.169105
R7476 CSoutput.n60 CSoutput.n59 0.169105
R7477 CSoutput.n60 CSoutput.n4 0.169105
R7478 CSoutput.n66 CSoutput.n4 0.169105
R7479 CSoutput.n67 CSoutput.n66 0.169105
R7480 CSoutput.n68 CSoutput.n67 0.169105
R7481 CSoutput.n68 CSoutput.n2 0.169105
R7482 CSoutput.n73 CSoutput.n2 0.169105
R7483 CSoutput.n74 CSoutput.n73 0.169105
R7484 CSoutput.n74 CSoutput.n0 0.169105
R7485 CSoutput.n78 CSoutput.n0 0.169105
R7486 CSoutput.n219 CSoutput.n218 0.0910737
R7487 CSoutput.n270 CSoutput.n267 0.0723685
R7488 CSoutput.n224 CSoutput.n219 0.0522944
R7489 CSoutput.n267 CSoutput.n266 0.0499135
R7490 CSoutput.n218 CSoutput.n217 0.0499135
R7491 CSoutput.n252 CSoutput.n251 0.0464294
R7492 CSoutput.n260 CSoutput.n257 0.0391444
R7493 CSoutput.n219 CSoutput.t154 0.023435
R7494 CSoutput.n267 CSoutput.t153 0.02262
R7495 CSoutput.n218 CSoutput.t157 0.02262
R7496 CSoutput CSoutput.n373 0.0052
R7497 CSoutput.n189 CSoutput.n172 0.00365111
R7498 CSoutput.n192 CSoutput.n173 0.00365111
R7499 CSoutput.n175 CSoutput.n174 0.00365111
R7500 CSoutput.n217 CSoutput.n176 0.00365111
R7501 CSoutput.n181 CSoutput.n177 0.00365111
R7502 CSoutput.n264 CSoutput.n178 0.00365111
R7503 CSoutput.n255 CSoutput.n254 0.00365111
R7504 CSoutput.n235 CSoutput.n208 0.00365111
R7505 CSoutput.n237 CSoutput.n207 0.00365111
R7506 CSoutput.n225 CSoutput.n224 0.00365111
R7507 CSoutput.n231 CSoutput.n211 0.00365111
R7508 CSoutput.n233 CSoutput.n210 0.00365111
R7509 CSoutput.n155 CSoutput.n138 0.00365111
R7510 CSoutput.n158 CSoutput.n139 0.00365111
R7511 CSoutput.n141 CSoutput.n140 0.00365111
R7512 CSoutput.n251 CSoutput.n142 0.00365111
R7513 CSoutput.n147 CSoutput.n143 0.00365111
R7514 CSoutput.n274 CSoutput.n144 0.00365111
R7515 CSoutput.n186 CSoutput.n176 0.00340054
R7516 CSoutput.n179 CSoutput.n177 0.00340054
R7517 CSoutput.n264 CSoutput.n263 0.00340054
R7518 CSoutput.n259 CSoutput.n172 0.00340054
R7519 CSoutput.n188 CSoutput.n173 0.00340054
R7520 CSoutput.n191 CSoutput.n175 0.00340054
R7521 CSoutput.n230 CSoutput.n225 0.00340054
R7522 CSoutput.n232 CSoutput.n231 0.00340054
R7523 CSoutput.n234 CSoutput.n233 0.00340054
R7524 CSoutput.n256 CSoutput.n255 0.00340054
R7525 CSoutput.n236 CSoutput.n235 0.00340054
R7526 CSoutput.n238 CSoutput.n237 0.00340054
R7527 CSoutput.n152 CSoutput.n142 0.00340054
R7528 CSoutput.n145 CSoutput.n143 0.00340054
R7529 CSoutput.n274 CSoutput.n273 0.00340054
R7530 CSoutput.n269 CSoutput.n138 0.00340054
R7531 CSoutput.n154 CSoutput.n139 0.00340054
R7532 CSoutput.n157 CSoutput.n141 0.00340054
R7533 CSoutput.n187 CSoutput.n181 0.00252698
R7534 CSoutput.n180 CSoutput.n178 0.00252698
R7535 CSoutput.n262 CSoutput.n261 0.00252698
R7536 CSoutput.n190 CSoutput.n188 0.00252698
R7537 CSoutput.n193 CSoutput.n191 0.00252698
R7538 CSoutput.n266 CSoutput.n161 0.00252698
R7539 CSoutput.n187 CSoutput.n186 0.00252698
R7540 CSoutput.n180 CSoutput.n179 0.00252698
R7541 CSoutput.n263 CSoutput.n262 0.00252698
R7542 CSoutput.n190 CSoutput.n189 0.00252698
R7543 CSoutput.n193 CSoutput.n192 0.00252698
R7544 CSoutput.n174 CSoutput.n161 0.00252698
R7545 CSoutput.n241 CSoutput.n211 0.00252698
R7546 CSoutput.n240 CSoutput.n210 0.00252698
R7547 CSoutput.n239 CSoutput.n195 0.00252698
R7548 CSoutput.n236 CSoutput.n206 0.00252698
R7549 CSoutput.n243 CSoutput.n238 0.00252698
R7550 CSoutput.n252 CSoutput.n245 0.00252698
R7551 CSoutput.n241 CSoutput.n230 0.00252698
R7552 CSoutput.n240 CSoutput.n232 0.00252698
R7553 CSoutput.n239 CSoutput.n234 0.00252698
R7554 CSoutput.n254 CSoutput.n206 0.00252698
R7555 CSoutput.n243 CSoutput.n208 0.00252698
R7556 CSoutput.n245 CSoutput.n207 0.00252698
R7557 CSoutput.n153 CSoutput.n147 0.00252698
R7558 CSoutput.n146 CSoutput.n144 0.00252698
R7559 CSoutput.n272 CSoutput.n271 0.00252698
R7560 CSoutput.n156 CSoutput.n154 0.00252698
R7561 CSoutput.n159 CSoutput.n157 0.00252698
R7562 CSoutput.n276 CSoutput.n127 0.00252698
R7563 CSoutput.n153 CSoutput.n152 0.00252698
R7564 CSoutput.n146 CSoutput.n145 0.00252698
R7565 CSoutput.n273 CSoutput.n272 0.00252698
R7566 CSoutput.n156 CSoutput.n155 0.00252698
R7567 CSoutput.n159 CSoutput.n158 0.00252698
R7568 CSoutput.n140 CSoutput.n127 0.00252698
R7569 CSoutput.n261 CSoutput.n260 0.0020275
R7570 CSoutput.n260 CSoutput.n259 0.0020275
R7571 CSoutput.n257 CSoutput.n195 0.0020275
R7572 CSoutput.n257 CSoutput.n256 0.0020275
R7573 CSoutput.n271 CSoutput.n270 0.0020275
R7574 CSoutput.n270 CSoutput.n269 0.0020275
R7575 CSoutput.n171 CSoutput.n170 0.00166668
R7576 CSoutput.n253 CSoutput.n209 0.00166668
R7577 CSoutput.n137 CSoutput.n136 0.00166668
R7578 CSoutput.n275 CSoutput.n137 0.00133328
R7579 CSoutput.n209 CSoutput.n205 0.00133328
R7580 CSoutput.n265 CSoutput.n171 0.00133328
R7581 CSoutput.n268 CSoutput.n160 0.001
R7582 CSoutput.n246 CSoutput.n160 0.001
R7583 CSoutput.n148 CSoutput.n128 0.001
R7584 CSoutput.n247 CSoutput.n128 0.001
R7585 CSoutput.n149 CSoutput.n129 0.001
R7586 CSoutput.n248 CSoutput.n129 0.001
R7587 CSoutput.n150 CSoutput.n130 0.001
R7588 CSoutput.n249 CSoutput.n130 0.001
R7589 CSoutput.n151 CSoutput.n131 0.001
R7590 CSoutput.n250 CSoutput.n131 0.001
R7591 CSoutput.n244 CSoutput.n196 0.001
R7592 CSoutput.n244 CSoutput.n242 0.001
R7593 CSoutput.n226 CSoutput.n197 0.001
R7594 CSoutput.n220 CSoutput.n197 0.001
R7595 CSoutput.n227 CSoutput.n198 0.001
R7596 CSoutput.n221 CSoutput.n198 0.001
R7597 CSoutput.n228 CSoutput.n199 0.001
R7598 CSoutput.n222 CSoutput.n199 0.001
R7599 CSoutput.n229 CSoutput.n200 0.001
R7600 CSoutput.n223 CSoutput.n200 0.001
R7601 CSoutput.n258 CSoutput.n194 0.001
R7602 CSoutput.n212 CSoutput.n194 0.001
R7603 CSoutput.n182 CSoutput.n162 0.001
R7604 CSoutput.n213 CSoutput.n162 0.001
R7605 CSoutput.n183 CSoutput.n163 0.001
R7606 CSoutput.n214 CSoutput.n163 0.001
R7607 CSoutput.n184 CSoutput.n164 0.001
R7608 CSoutput.n215 CSoutput.n164 0.001
R7609 CSoutput.n185 CSoutput.n165 0.001
R7610 CSoutput.n216 CSoutput.n165 0.001
R7611 CSoutput.n216 CSoutput.n166 0.001
R7612 CSoutput.n215 CSoutput.n167 0.001
R7613 CSoutput.n214 CSoutput.n168 0.001
R7614 CSoutput.n213 CSoutput.t152 0.001
R7615 CSoutput.n212 CSoutput.n169 0.001
R7616 CSoutput.n185 CSoutput.n167 0.001
R7617 CSoutput.n184 CSoutput.n168 0.001
R7618 CSoutput.n183 CSoutput.t152 0.001
R7619 CSoutput.n182 CSoutput.n169 0.001
R7620 CSoutput.n258 CSoutput.n170 0.001
R7621 CSoutput.n223 CSoutput.n201 0.001
R7622 CSoutput.n222 CSoutput.n202 0.001
R7623 CSoutput.n221 CSoutput.n203 0.001
R7624 CSoutput.n220 CSoutput.t146 0.001
R7625 CSoutput.n242 CSoutput.n204 0.001
R7626 CSoutput.n229 CSoutput.n202 0.001
R7627 CSoutput.n228 CSoutput.n203 0.001
R7628 CSoutput.n227 CSoutput.t146 0.001
R7629 CSoutput.n226 CSoutput.n204 0.001
R7630 CSoutput.n253 CSoutput.n196 0.001
R7631 CSoutput.n250 CSoutput.n132 0.001
R7632 CSoutput.n249 CSoutput.n133 0.001
R7633 CSoutput.n248 CSoutput.n134 0.001
R7634 CSoutput.n247 CSoutput.t164 0.001
R7635 CSoutput.n246 CSoutput.n135 0.001
R7636 CSoutput.n151 CSoutput.n133 0.001
R7637 CSoutput.n150 CSoutput.n134 0.001
R7638 CSoutput.n149 CSoutput.t164 0.001
R7639 CSoutput.n148 CSoutput.n135 0.001
R7640 CSoutput.n268 CSoutput.n136 0.001
R7641 gnd.n6535 gnd.n403 2174.34
R7642 gnd.n3785 gnd.n3555 939.716
R7643 gnd.n6844 gnd.n84 838.452
R7644 gnd.n7007 gnd.n80 838.452
R7645 gnd.n5111 gnd.n1128 838.452
R7646 gnd.n5030 gnd.n1130 838.452
R7647 gnd.n5853 gnd.n997 838.452
R7648 gnd.n4141 gnd.n995 838.452
R7649 gnd.n3642 gnd.n3583 838.452
R7650 gnd.n3787 gnd.n2098 838.452
R7651 gnd.n7005 gnd.n86 819.232
R7652 gnd.n154 gnd.n82 819.232
R7653 gnd.n5461 gnd.n1127 819.232
R7654 gnd.n5706 gnd.n1131 819.232
R7655 gnd.n5855 gnd.n992 819.232
R7656 gnd.n4308 gnd.n994 819.232
R7657 gnd.n3707 gnd.n3706 819.232
R7658 gnd.n3783 gnd.n2094 819.232
R7659 gnd.n4187 gnd.n1002 771.183
R7660 gnd.n5724 gnd.n1105 771.183
R7661 gnd.n4070 gnd.n1928 771.183
R7662 gnd.n5144 gnd.n1107 771.183
R7663 gnd.n3463 gnd.n2106 766.379
R7664 gnd.n3466 gnd.n3465 766.379
R7665 gnd.n2704 gnd.n2607 766.379
R7666 gnd.n2700 gnd.n2605 766.379
R7667 gnd.n3554 gnd.n2128 756.769
R7668 gnd.n3457 gnd.n3456 756.769
R7669 gnd.n2797 gnd.n2514 756.769
R7670 gnd.n2795 gnd.n2517 756.769
R7671 gnd.n6116 gnd.n656 756.769
R7672 gnd.n6536 gnd.n404 756.769
R7673 gnd.n6749 gnd.n277 756.769
R7674 gnd.n5948 gnd.n826 756.769
R7675 gnd.n6117 gnd.n6116 585
R7676 gnd.n6116 gnd.n6115 585
R7677 gnd.n660 gnd.n659 585
R7678 gnd.n6114 gnd.n660 585
R7679 gnd.n6112 gnd.n6111 585
R7680 gnd.n6113 gnd.n6112 585
R7681 gnd.n6110 gnd.n662 585
R7682 gnd.n662 gnd.n661 585
R7683 gnd.n6109 gnd.n6108 585
R7684 gnd.n6108 gnd.n6107 585
R7685 gnd.n667 gnd.n666 585
R7686 gnd.n6106 gnd.n667 585
R7687 gnd.n6104 gnd.n6103 585
R7688 gnd.n6105 gnd.n6104 585
R7689 gnd.n6102 gnd.n669 585
R7690 gnd.n669 gnd.n668 585
R7691 gnd.n6101 gnd.n6100 585
R7692 gnd.n6100 gnd.n6099 585
R7693 gnd.n675 gnd.n674 585
R7694 gnd.n6098 gnd.n675 585
R7695 gnd.n6096 gnd.n6095 585
R7696 gnd.n6097 gnd.n6096 585
R7697 gnd.n6094 gnd.n677 585
R7698 gnd.n677 gnd.n676 585
R7699 gnd.n6093 gnd.n6092 585
R7700 gnd.n6092 gnd.n6091 585
R7701 gnd.n683 gnd.n682 585
R7702 gnd.n6090 gnd.n683 585
R7703 gnd.n6088 gnd.n6087 585
R7704 gnd.n6089 gnd.n6088 585
R7705 gnd.n6086 gnd.n685 585
R7706 gnd.n685 gnd.n684 585
R7707 gnd.n6085 gnd.n6084 585
R7708 gnd.n6084 gnd.n6083 585
R7709 gnd.n691 gnd.n690 585
R7710 gnd.n6082 gnd.n691 585
R7711 gnd.n6080 gnd.n6079 585
R7712 gnd.n6081 gnd.n6080 585
R7713 gnd.n6078 gnd.n693 585
R7714 gnd.n693 gnd.n692 585
R7715 gnd.n6077 gnd.n6076 585
R7716 gnd.n6076 gnd.n6075 585
R7717 gnd.n699 gnd.n698 585
R7718 gnd.n6074 gnd.n699 585
R7719 gnd.n6072 gnd.n6071 585
R7720 gnd.n6073 gnd.n6072 585
R7721 gnd.n6070 gnd.n701 585
R7722 gnd.n701 gnd.n700 585
R7723 gnd.n6069 gnd.n6068 585
R7724 gnd.n6068 gnd.n6067 585
R7725 gnd.n707 gnd.n706 585
R7726 gnd.n6066 gnd.n707 585
R7727 gnd.n6064 gnd.n6063 585
R7728 gnd.n6065 gnd.n6064 585
R7729 gnd.n6062 gnd.n709 585
R7730 gnd.n709 gnd.n708 585
R7731 gnd.n6061 gnd.n6060 585
R7732 gnd.n6060 gnd.n6059 585
R7733 gnd.n715 gnd.n714 585
R7734 gnd.n6058 gnd.n715 585
R7735 gnd.n6056 gnd.n6055 585
R7736 gnd.n6057 gnd.n6056 585
R7737 gnd.n6054 gnd.n717 585
R7738 gnd.n717 gnd.n716 585
R7739 gnd.n6053 gnd.n6052 585
R7740 gnd.n6052 gnd.n6051 585
R7741 gnd.n723 gnd.n722 585
R7742 gnd.n6050 gnd.n723 585
R7743 gnd.n6048 gnd.n6047 585
R7744 gnd.n6049 gnd.n6048 585
R7745 gnd.n6046 gnd.n725 585
R7746 gnd.n725 gnd.n724 585
R7747 gnd.n6045 gnd.n6044 585
R7748 gnd.n6044 gnd.n6043 585
R7749 gnd.n731 gnd.n730 585
R7750 gnd.n6042 gnd.n731 585
R7751 gnd.n6040 gnd.n6039 585
R7752 gnd.n6041 gnd.n6040 585
R7753 gnd.n6038 gnd.n733 585
R7754 gnd.n733 gnd.n732 585
R7755 gnd.n6037 gnd.n6036 585
R7756 gnd.n6036 gnd.n6035 585
R7757 gnd.n739 gnd.n738 585
R7758 gnd.n6034 gnd.n739 585
R7759 gnd.n6032 gnd.n6031 585
R7760 gnd.n6033 gnd.n6032 585
R7761 gnd.n6030 gnd.n741 585
R7762 gnd.n741 gnd.n740 585
R7763 gnd.n6029 gnd.n6028 585
R7764 gnd.n6028 gnd.n6027 585
R7765 gnd.n747 gnd.n746 585
R7766 gnd.n6026 gnd.n747 585
R7767 gnd.n6024 gnd.n6023 585
R7768 gnd.n6025 gnd.n6024 585
R7769 gnd.n6022 gnd.n749 585
R7770 gnd.n749 gnd.n748 585
R7771 gnd.n6021 gnd.n6020 585
R7772 gnd.n6020 gnd.n6019 585
R7773 gnd.n755 gnd.n754 585
R7774 gnd.n6018 gnd.n755 585
R7775 gnd.n6016 gnd.n6015 585
R7776 gnd.n6017 gnd.n6016 585
R7777 gnd.n6014 gnd.n757 585
R7778 gnd.n757 gnd.n756 585
R7779 gnd.n6013 gnd.n6012 585
R7780 gnd.n6012 gnd.n6011 585
R7781 gnd.n763 gnd.n762 585
R7782 gnd.n6010 gnd.n763 585
R7783 gnd.n6008 gnd.n6007 585
R7784 gnd.n6009 gnd.n6008 585
R7785 gnd.n6006 gnd.n765 585
R7786 gnd.n765 gnd.n764 585
R7787 gnd.n6005 gnd.n6004 585
R7788 gnd.n6004 gnd.n6003 585
R7789 gnd.n771 gnd.n770 585
R7790 gnd.n6002 gnd.n771 585
R7791 gnd.n6000 gnd.n5999 585
R7792 gnd.n6001 gnd.n6000 585
R7793 gnd.n5998 gnd.n773 585
R7794 gnd.n773 gnd.n772 585
R7795 gnd.n5997 gnd.n5996 585
R7796 gnd.n5996 gnd.n5995 585
R7797 gnd.n779 gnd.n778 585
R7798 gnd.n5994 gnd.n779 585
R7799 gnd.n5992 gnd.n5991 585
R7800 gnd.n5993 gnd.n5992 585
R7801 gnd.n5990 gnd.n781 585
R7802 gnd.n781 gnd.n780 585
R7803 gnd.n5989 gnd.n5988 585
R7804 gnd.n5988 gnd.n5987 585
R7805 gnd.n787 gnd.n786 585
R7806 gnd.n5986 gnd.n787 585
R7807 gnd.n5984 gnd.n5983 585
R7808 gnd.n5985 gnd.n5984 585
R7809 gnd.n5982 gnd.n789 585
R7810 gnd.n789 gnd.n788 585
R7811 gnd.n5981 gnd.n5980 585
R7812 gnd.n5980 gnd.n5979 585
R7813 gnd.n795 gnd.n794 585
R7814 gnd.n5978 gnd.n795 585
R7815 gnd.n5976 gnd.n5975 585
R7816 gnd.n5977 gnd.n5976 585
R7817 gnd.n5974 gnd.n797 585
R7818 gnd.n797 gnd.n796 585
R7819 gnd.n5973 gnd.n5972 585
R7820 gnd.n5972 gnd.n5971 585
R7821 gnd.n803 gnd.n802 585
R7822 gnd.n5970 gnd.n803 585
R7823 gnd.n5968 gnd.n5967 585
R7824 gnd.n5969 gnd.n5968 585
R7825 gnd.n5966 gnd.n805 585
R7826 gnd.n805 gnd.n804 585
R7827 gnd.n5965 gnd.n5964 585
R7828 gnd.n5964 gnd.n5963 585
R7829 gnd.n811 gnd.n810 585
R7830 gnd.n5962 gnd.n811 585
R7831 gnd.n5960 gnd.n5959 585
R7832 gnd.n5961 gnd.n5960 585
R7833 gnd.n5958 gnd.n813 585
R7834 gnd.n813 gnd.n812 585
R7835 gnd.n5957 gnd.n5956 585
R7836 gnd.n5956 gnd.n5955 585
R7837 gnd.n819 gnd.n818 585
R7838 gnd.n5954 gnd.n819 585
R7839 gnd.n5952 gnd.n5951 585
R7840 gnd.n5953 gnd.n5952 585
R7841 gnd.n5950 gnd.n821 585
R7842 gnd.n821 gnd.n820 585
R7843 gnd.n657 gnd.n656 585
R7844 gnd.n656 gnd.n655 585
R7845 gnd.n6122 gnd.n6121 585
R7846 gnd.n6123 gnd.n6122 585
R7847 gnd.n654 gnd.n653 585
R7848 gnd.n6124 gnd.n654 585
R7849 gnd.n6127 gnd.n6126 585
R7850 gnd.n6126 gnd.n6125 585
R7851 gnd.n651 gnd.n650 585
R7852 gnd.n650 gnd.n649 585
R7853 gnd.n6132 gnd.n6131 585
R7854 gnd.n6133 gnd.n6132 585
R7855 gnd.n648 gnd.n647 585
R7856 gnd.n6134 gnd.n648 585
R7857 gnd.n6137 gnd.n6136 585
R7858 gnd.n6136 gnd.n6135 585
R7859 gnd.n645 gnd.n644 585
R7860 gnd.n644 gnd.n643 585
R7861 gnd.n6142 gnd.n6141 585
R7862 gnd.n6143 gnd.n6142 585
R7863 gnd.n642 gnd.n641 585
R7864 gnd.n6144 gnd.n642 585
R7865 gnd.n6147 gnd.n6146 585
R7866 gnd.n6146 gnd.n6145 585
R7867 gnd.n639 gnd.n638 585
R7868 gnd.n638 gnd.n637 585
R7869 gnd.n6152 gnd.n6151 585
R7870 gnd.n6153 gnd.n6152 585
R7871 gnd.n636 gnd.n635 585
R7872 gnd.n6154 gnd.n636 585
R7873 gnd.n6157 gnd.n6156 585
R7874 gnd.n6156 gnd.n6155 585
R7875 gnd.n633 gnd.n632 585
R7876 gnd.n632 gnd.n631 585
R7877 gnd.n6162 gnd.n6161 585
R7878 gnd.n6163 gnd.n6162 585
R7879 gnd.n630 gnd.n629 585
R7880 gnd.n6164 gnd.n630 585
R7881 gnd.n6167 gnd.n6166 585
R7882 gnd.n6166 gnd.n6165 585
R7883 gnd.n627 gnd.n626 585
R7884 gnd.n626 gnd.n625 585
R7885 gnd.n6172 gnd.n6171 585
R7886 gnd.n6173 gnd.n6172 585
R7887 gnd.n624 gnd.n623 585
R7888 gnd.n6174 gnd.n624 585
R7889 gnd.n6177 gnd.n6176 585
R7890 gnd.n6176 gnd.n6175 585
R7891 gnd.n621 gnd.n620 585
R7892 gnd.n620 gnd.n619 585
R7893 gnd.n6182 gnd.n6181 585
R7894 gnd.n6183 gnd.n6182 585
R7895 gnd.n618 gnd.n617 585
R7896 gnd.n6184 gnd.n618 585
R7897 gnd.n6187 gnd.n6186 585
R7898 gnd.n6186 gnd.n6185 585
R7899 gnd.n615 gnd.n614 585
R7900 gnd.n614 gnd.n613 585
R7901 gnd.n6192 gnd.n6191 585
R7902 gnd.n6193 gnd.n6192 585
R7903 gnd.n612 gnd.n611 585
R7904 gnd.n6194 gnd.n612 585
R7905 gnd.n6197 gnd.n6196 585
R7906 gnd.n6196 gnd.n6195 585
R7907 gnd.n609 gnd.n608 585
R7908 gnd.n608 gnd.n607 585
R7909 gnd.n6202 gnd.n6201 585
R7910 gnd.n6203 gnd.n6202 585
R7911 gnd.n606 gnd.n605 585
R7912 gnd.n6204 gnd.n606 585
R7913 gnd.n6207 gnd.n6206 585
R7914 gnd.n6206 gnd.n6205 585
R7915 gnd.n603 gnd.n602 585
R7916 gnd.n602 gnd.n601 585
R7917 gnd.n6212 gnd.n6211 585
R7918 gnd.n6213 gnd.n6212 585
R7919 gnd.n600 gnd.n599 585
R7920 gnd.n6214 gnd.n600 585
R7921 gnd.n6217 gnd.n6216 585
R7922 gnd.n6216 gnd.n6215 585
R7923 gnd.n597 gnd.n596 585
R7924 gnd.n596 gnd.n595 585
R7925 gnd.n6222 gnd.n6221 585
R7926 gnd.n6223 gnd.n6222 585
R7927 gnd.n594 gnd.n593 585
R7928 gnd.n6224 gnd.n594 585
R7929 gnd.n6227 gnd.n6226 585
R7930 gnd.n6226 gnd.n6225 585
R7931 gnd.n591 gnd.n590 585
R7932 gnd.n590 gnd.n589 585
R7933 gnd.n6232 gnd.n6231 585
R7934 gnd.n6233 gnd.n6232 585
R7935 gnd.n588 gnd.n587 585
R7936 gnd.n6234 gnd.n588 585
R7937 gnd.n6237 gnd.n6236 585
R7938 gnd.n6236 gnd.n6235 585
R7939 gnd.n585 gnd.n584 585
R7940 gnd.n584 gnd.n583 585
R7941 gnd.n6242 gnd.n6241 585
R7942 gnd.n6243 gnd.n6242 585
R7943 gnd.n582 gnd.n581 585
R7944 gnd.n6244 gnd.n582 585
R7945 gnd.n6247 gnd.n6246 585
R7946 gnd.n6246 gnd.n6245 585
R7947 gnd.n579 gnd.n578 585
R7948 gnd.n578 gnd.n577 585
R7949 gnd.n6252 gnd.n6251 585
R7950 gnd.n6253 gnd.n6252 585
R7951 gnd.n576 gnd.n575 585
R7952 gnd.n6254 gnd.n576 585
R7953 gnd.n6257 gnd.n6256 585
R7954 gnd.n6256 gnd.n6255 585
R7955 gnd.n573 gnd.n572 585
R7956 gnd.n572 gnd.n571 585
R7957 gnd.n6262 gnd.n6261 585
R7958 gnd.n6263 gnd.n6262 585
R7959 gnd.n570 gnd.n569 585
R7960 gnd.n6264 gnd.n570 585
R7961 gnd.n6267 gnd.n6266 585
R7962 gnd.n6266 gnd.n6265 585
R7963 gnd.n567 gnd.n566 585
R7964 gnd.n566 gnd.n565 585
R7965 gnd.n6272 gnd.n6271 585
R7966 gnd.n6273 gnd.n6272 585
R7967 gnd.n564 gnd.n563 585
R7968 gnd.n6274 gnd.n564 585
R7969 gnd.n6277 gnd.n6276 585
R7970 gnd.n6276 gnd.n6275 585
R7971 gnd.n561 gnd.n560 585
R7972 gnd.n560 gnd.n559 585
R7973 gnd.n6282 gnd.n6281 585
R7974 gnd.n6283 gnd.n6282 585
R7975 gnd.n558 gnd.n557 585
R7976 gnd.n6284 gnd.n558 585
R7977 gnd.n6287 gnd.n6286 585
R7978 gnd.n6286 gnd.n6285 585
R7979 gnd.n555 gnd.n554 585
R7980 gnd.n554 gnd.n553 585
R7981 gnd.n6292 gnd.n6291 585
R7982 gnd.n6293 gnd.n6292 585
R7983 gnd.n552 gnd.n551 585
R7984 gnd.n6294 gnd.n552 585
R7985 gnd.n6297 gnd.n6296 585
R7986 gnd.n6296 gnd.n6295 585
R7987 gnd.n549 gnd.n548 585
R7988 gnd.n548 gnd.n547 585
R7989 gnd.n6302 gnd.n6301 585
R7990 gnd.n6303 gnd.n6302 585
R7991 gnd.n546 gnd.n545 585
R7992 gnd.n6304 gnd.n546 585
R7993 gnd.n6307 gnd.n6306 585
R7994 gnd.n6306 gnd.n6305 585
R7995 gnd.n543 gnd.n542 585
R7996 gnd.n542 gnd.n541 585
R7997 gnd.n6312 gnd.n6311 585
R7998 gnd.n6313 gnd.n6312 585
R7999 gnd.n540 gnd.n539 585
R8000 gnd.n6314 gnd.n540 585
R8001 gnd.n6317 gnd.n6316 585
R8002 gnd.n6316 gnd.n6315 585
R8003 gnd.n537 gnd.n536 585
R8004 gnd.n536 gnd.n535 585
R8005 gnd.n6322 gnd.n6321 585
R8006 gnd.n6323 gnd.n6322 585
R8007 gnd.n534 gnd.n533 585
R8008 gnd.n6324 gnd.n534 585
R8009 gnd.n6327 gnd.n6326 585
R8010 gnd.n6326 gnd.n6325 585
R8011 gnd.n531 gnd.n530 585
R8012 gnd.n530 gnd.n529 585
R8013 gnd.n6332 gnd.n6331 585
R8014 gnd.n6333 gnd.n6332 585
R8015 gnd.n528 gnd.n527 585
R8016 gnd.n6334 gnd.n528 585
R8017 gnd.n6337 gnd.n6336 585
R8018 gnd.n6336 gnd.n6335 585
R8019 gnd.n525 gnd.n524 585
R8020 gnd.n524 gnd.n523 585
R8021 gnd.n6342 gnd.n6341 585
R8022 gnd.n6343 gnd.n6342 585
R8023 gnd.n522 gnd.n521 585
R8024 gnd.n6344 gnd.n522 585
R8025 gnd.n6347 gnd.n6346 585
R8026 gnd.n6346 gnd.n6345 585
R8027 gnd.n519 gnd.n518 585
R8028 gnd.n518 gnd.n517 585
R8029 gnd.n6352 gnd.n6351 585
R8030 gnd.n6353 gnd.n6352 585
R8031 gnd.n516 gnd.n515 585
R8032 gnd.n6354 gnd.n516 585
R8033 gnd.n6357 gnd.n6356 585
R8034 gnd.n6356 gnd.n6355 585
R8035 gnd.n513 gnd.n512 585
R8036 gnd.n512 gnd.n511 585
R8037 gnd.n6362 gnd.n6361 585
R8038 gnd.n6363 gnd.n6362 585
R8039 gnd.n510 gnd.n509 585
R8040 gnd.n6364 gnd.n510 585
R8041 gnd.n6367 gnd.n6366 585
R8042 gnd.n6366 gnd.n6365 585
R8043 gnd.n507 gnd.n506 585
R8044 gnd.n506 gnd.n505 585
R8045 gnd.n6372 gnd.n6371 585
R8046 gnd.n6373 gnd.n6372 585
R8047 gnd.n504 gnd.n503 585
R8048 gnd.n6374 gnd.n504 585
R8049 gnd.n6377 gnd.n6376 585
R8050 gnd.n6376 gnd.n6375 585
R8051 gnd.n501 gnd.n500 585
R8052 gnd.n500 gnd.n499 585
R8053 gnd.n6382 gnd.n6381 585
R8054 gnd.n6383 gnd.n6382 585
R8055 gnd.n498 gnd.n497 585
R8056 gnd.n6384 gnd.n498 585
R8057 gnd.n6387 gnd.n6386 585
R8058 gnd.n6386 gnd.n6385 585
R8059 gnd.n495 gnd.n494 585
R8060 gnd.n494 gnd.n493 585
R8061 gnd.n6392 gnd.n6391 585
R8062 gnd.n6393 gnd.n6392 585
R8063 gnd.n492 gnd.n491 585
R8064 gnd.n6394 gnd.n492 585
R8065 gnd.n6397 gnd.n6396 585
R8066 gnd.n6396 gnd.n6395 585
R8067 gnd.n489 gnd.n488 585
R8068 gnd.n488 gnd.n487 585
R8069 gnd.n6402 gnd.n6401 585
R8070 gnd.n6403 gnd.n6402 585
R8071 gnd.n486 gnd.n485 585
R8072 gnd.n6404 gnd.n486 585
R8073 gnd.n6407 gnd.n6406 585
R8074 gnd.n6406 gnd.n6405 585
R8075 gnd.n483 gnd.n482 585
R8076 gnd.n482 gnd.n481 585
R8077 gnd.n6412 gnd.n6411 585
R8078 gnd.n6413 gnd.n6412 585
R8079 gnd.n480 gnd.n479 585
R8080 gnd.n6414 gnd.n480 585
R8081 gnd.n6417 gnd.n6416 585
R8082 gnd.n6416 gnd.n6415 585
R8083 gnd.n477 gnd.n476 585
R8084 gnd.n476 gnd.n475 585
R8085 gnd.n6422 gnd.n6421 585
R8086 gnd.n6423 gnd.n6422 585
R8087 gnd.n474 gnd.n473 585
R8088 gnd.n6424 gnd.n474 585
R8089 gnd.n6427 gnd.n6426 585
R8090 gnd.n6426 gnd.n6425 585
R8091 gnd.n471 gnd.n470 585
R8092 gnd.n470 gnd.n469 585
R8093 gnd.n6432 gnd.n6431 585
R8094 gnd.n6433 gnd.n6432 585
R8095 gnd.n468 gnd.n467 585
R8096 gnd.n6434 gnd.n468 585
R8097 gnd.n6437 gnd.n6436 585
R8098 gnd.n6436 gnd.n6435 585
R8099 gnd.n465 gnd.n464 585
R8100 gnd.n464 gnd.n463 585
R8101 gnd.n6442 gnd.n6441 585
R8102 gnd.n6443 gnd.n6442 585
R8103 gnd.n462 gnd.n461 585
R8104 gnd.n6444 gnd.n462 585
R8105 gnd.n6447 gnd.n6446 585
R8106 gnd.n6446 gnd.n6445 585
R8107 gnd.n459 gnd.n458 585
R8108 gnd.n458 gnd.n457 585
R8109 gnd.n6452 gnd.n6451 585
R8110 gnd.n6453 gnd.n6452 585
R8111 gnd.n456 gnd.n455 585
R8112 gnd.n6454 gnd.n456 585
R8113 gnd.n6457 gnd.n6456 585
R8114 gnd.n6456 gnd.n6455 585
R8115 gnd.n453 gnd.n452 585
R8116 gnd.n452 gnd.n451 585
R8117 gnd.n6462 gnd.n6461 585
R8118 gnd.n6463 gnd.n6462 585
R8119 gnd.n450 gnd.n449 585
R8120 gnd.n6464 gnd.n450 585
R8121 gnd.n6467 gnd.n6466 585
R8122 gnd.n6466 gnd.n6465 585
R8123 gnd.n447 gnd.n446 585
R8124 gnd.n446 gnd.n445 585
R8125 gnd.n6472 gnd.n6471 585
R8126 gnd.n6473 gnd.n6472 585
R8127 gnd.n444 gnd.n443 585
R8128 gnd.n6474 gnd.n444 585
R8129 gnd.n6477 gnd.n6476 585
R8130 gnd.n6476 gnd.n6475 585
R8131 gnd.n441 gnd.n440 585
R8132 gnd.n440 gnd.n439 585
R8133 gnd.n6482 gnd.n6481 585
R8134 gnd.n6483 gnd.n6482 585
R8135 gnd.n438 gnd.n437 585
R8136 gnd.n6484 gnd.n438 585
R8137 gnd.n6487 gnd.n6486 585
R8138 gnd.n6486 gnd.n6485 585
R8139 gnd.n435 gnd.n434 585
R8140 gnd.n434 gnd.n433 585
R8141 gnd.n6492 gnd.n6491 585
R8142 gnd.n6493 gnd.n6492 585
R8143 gnd.n432 gnd.n431 585
R8144 gnd.n6494 gnd.n432 585
R8145 gnd.n6497 gnd.n6496 585
R8146 gnd.n6496 gnd.n6495 585
R8147 gnd.n429 gnd.n428 585
R8148 gnd.n428 gnd.n427 585
R8149 gnd.n6502 gnd.n6501 585
R8150 gnd.n6503 gnd.n6502 585
R8151 gnd.n426 gnd.n425 585
R8152 gnd.n6504 gnd.n426 585
R8153 gnd.n6507 gnd.n6506 585
R8154 gnd.n6506 gnd.n6505 585
R8155 gnd.n423 gnd.n422 585
R8156 gnd.n422 gnd.n421 585
R8157 gnd.n6512 gnd.n6511 585
R8158 gnd.n6513 gnd.n6512 585
R8159 gnd.n420 gnd.n419 585
R8160 gnd.n6514 gnd.n420 585
R8161 gnd.n6517 gnd.n6516 585
R8162 gnd.n6516 gnd.n6515 585
R8163 gnd.n417 gnd.n416 585
R8164 gnd.n416 gnd.n415 585
R8165 gnd.n6522 gnd.n6521 585
R8166 gnd.n6523 gnd.n6522 585
R8167 gnd.n414 gnd.n413 585
R8168 gnd.n6524 gnd.n414 585
R8169 gnd.n6527 gnd.n6526 585
R8170 gnd.n6526 gnd.n6525 585
R8171 gnd.n411 gnd.n410 585
R8172 gnd.n410 gnd.n409 585
R8173 gnd.n6532 gnd.n6531 585
R8174 gnd.n6533 gnd.n6532 585
R8175 gnd.n408 gnd.n407 585
R8176 gnd.n6534 gnd.n408 585
R8177 gnd.n6537 gnd.n6536 585
R8178 gnd.n6536 gnd.n6535 585
R8179 gnd.n6748 gnd.n281 585
R8180 gnd.n6748 gnd.n6747 585
R8181 gnd.n6742 gnd.n282 585
R8182 gnd.n6746 gnd.n282 585
R8183 gnd.n6744 gnd.n6743 585
R8184 gnd.n6745 gnd.n6744 585
R8185 gnd.n285 gnd.n284 585
R8186 gnd.n284 gnd.n283 585
R8187 gnd.n6737 gnd.n6736 585
R8188 gnd.n6736 gnd.n6735 585
R8189 gnd.n288 gnd.n287 585
R8190 gnd.n6734 gnd.n288 585
R8191 gnd.n6732 gnd.n6731 585
R8192 gnd.n6733 gnd.n6732 585
R8193 gnd.n291 gnd.n290 585
R8194 gnd.n290 gnd.n289 585
R8195 gnd.n6727 gnd.n6726 585
R8196 gnd.n6726 gnd.n6725 585
R8197 gnd.n294 gnd.n293 585
R8198 gnd.n6724 gnd.n294 585
R8199 gnd.n6722 gnd.n6721 585
R8200 gnd.n6723 gnd.n6722 585
R8201 gnd.n297 gnd.n296 585
R8202 gnd.n296 gnd.n295 585
R8203 gnd.n6717 gnd.n6716 585
R8204 gnd.n6716 gnd.n6715 585
R8205 gnd.n300 gnd.n299 585
R8206 gnd.n6714 gnd.n300 585
R8207 gnd.n6712 gnd.n6711 585
R8208 gnd.n6713 gnd.n6712 585
R8209 gnd.n303 gnd.n302 585
R8210 gnd.n302 gnd.n301 585
R8211 gnd.n6707 gnd.n6706 585
R8212 gnd.n6706 gnd.n6705 585
R8213 gnd.n306 gnd.n305 585
R8214 gnd.n6704 gnd.n306 585
R8215 gnd.n6702 gnd.n6701 585
R8216 gnd.n6703 gnd.n6702 585
R8217 gnd.n309 gnd.n308 585
R8218 gnd.n308 gnd.n307 585
R8219 gnd.n6697 gnd.n6696 585
R8220 gnd.n6696 gnd.n6695 585
R8221 gnd.n312 gnd.n311 585
R8222 gnd.n6694 gnd.n312 585
R8223 gnd.n6692 gnd.n6691 585
R8224 gnd.n6693 gnd.n6692 585
R8225 gnd.n315 gnd.n314 585
R8226 gnd.n314 gnd.n313 585
R8227 gnd.n6687 gnd.n6686 585
R8228 gnd.n6686 gnd.n6685 585
R8229 gnd.n318 gnd.n317 585
R8230 gnd.n6684 gnd.n318 585
R8231 gnd.n6682 gnd.n6681 585
R8232 gnd.n6683 gnd.n6682 585
R8233 gnd.n321 gnd.n320 585
R8234 gnd.n320 gnd.n319 585
R8235 gnd.n6677 gnd.n6676 585
R8236 gnd.n6676 gnd.n6675 585
R8237 gnd.n324 gnd.n323 585
R8238 gnd.n6674 gnd.n324 585
R8239 gnd.n6672 gnd.n6671 585
R8240 gnd.n6673 gnd.n6672 585
R8241 gnd.n327 gnd.n326 585
R8242 gnd.n326 gnd.n325 585
R8243 gnd.n6667 gnd.n6666 585
R8244 gnd.n6666 gnd.n6665 585
R8245 gnd.n330 gnd.n329 585
R8246 gnd.n6664 gnd.n330 585
R8247 gnd.n6662 gnd.n6661 585
R8248 gnd.n6663 gnd.n6662 585
R8249 gnd.n333 gnd.n332 585
R8250 gnd.n332 gnd.n331 585
R8251 gnd.n6657 gnd.n6656 585
R8252 gnd.n6656 gnd.n6655 585
R8253 gnd.n336 gnd.n335 585
R8254 gnd.n6654 gnd.n336 585
R8255 gnd.n6652 gnd.n6651 585
R8256 gnd.n6653 gnd.n6652 585
R8257 gnd.n339 gnd.n338 585
R8258 gnd.n338 gnd.n337 585
R8259 gnd.n6647 gnd.n6646 585
R8260 gnd.n6646 gnd.n6645 585
R8261 gnd.n342 gnd.n341 585
R8262 gnd.n6644 gnd.n342 585
R8263 gnd.n6642 gnd.n6641 585
R8264 gnd.n6643 gnd.n6642 585
R8265 gnd.n345 gnd.n344 585
R8266 gnd.n344 gnd.n343 585
R8267 gnd.n6637 gnd.n6636 585
R8268 gnd.n6636 gnd.n6635 585
R8269 gnd.n348 gnd.n347 585
R8270 gnd.n6634 gnd.n348 585
R8271 gnd.n6632 gnd.n6631 585
R8272 gnd.n6633 gnd.n6632 585
R8273 gnd.n351 gnd.n350 585
R8274 gnd.n350 gnd.n349 585
R8275 gnd.n6627 gnd.n6626 585
R8276 gnd.n6626 gnd.n6625 585
R8277 gnd.n354 gnd.n353 585
R8278 gnd.n6624 gnd.n354 585
R8279 gnd.n6622 gnd.n6621 585
R8280 gnd.n6623 gnd.n6622 585
R8281 gnd.n357 gnd.n356 585
R8282 gnd.n356 gnd.n355 585
R8283 gnd.n6617 gnd.n6616 585
R8284 gnd.n6616 gnd.n6615 585
R8285 gnd.n360 gnd.n359 585
R8286 gnd.n6614 gnd.n360 585
R8287 gnd.n6612 gnd.n6611 585
R8288 gnd.n6613 gnd.n6612 585
R8289 gnd.n363 gnd.n362 585
R8290 gnd.n362 gnd.n361 585
R8291 gnd.n6607 gnd.n6606 585
R8292 gnd.n6606 gnd.n6605 585
R8293 gnd.n366 gnd.n365 585
R8294 gnd.n6604 gnd.n366 585
R8295 gnd.n6602 gnd.n6601 585
R8296 gnd.n6603 gnd.n6602 585
R8297 gnd.n369 gnd.n368 585
R8298 gnd.n368 gnd.n367 585
R8299 gnd.n6597 gnd.n6596 585
R8300 gnd.n6596 gnd.n6595 585
R8301 gnd.n372 gnd.n371 585
R8302 gnd.n6594 gnd.n372 585
R8303 gnd.n6592 gnd.n6591 585
R8304 gnd.n6593 gnd.n6592 585
R8305 gnd.n375 gnd.n374 585
R8306 gnd.n374 gnd.n373 585
R8307 gnd.n6587 gnd.n6586 585
R8308 gnd.n6586 gnd.n6585 585
R8309 gnd.n378 gnd.n377 585
R8310 gnd.n6584 gnd.n378 585
R8311 gnd.n6582 gnd.n6581 585
R8312 gnd.n6583 gnd.n6582 585
R8313 gnd.n381 gnd.n380 585
R8314 gnd.n380 gnd.n379 585
R8315 gnd.n6577 gnd.n6576 585
R8316 gnd.n6576 gnd.n6575 585
R8317 gnd.n384 gnd.n383 585
R8318 gnd.n6574 gnd.n384 585
R8319 gnd.n6572 gnd.n6571 585
R8320 gnd.n6573 gnd.n6572 585
R8321 gnd.n387 gnd.n386 585
R8322 gnd.n386 gnd.n385 585
R8323 gnd.n6567 gnd.n6566 585
R8324 gnd.n6566 gnd.n6565 585
R8325 gnd.n390 gnd.n389 585
R8326 gnd.n6564 gnd.n390 585
R8327 gnd.n6562 gnd.n6561 585
R8328 gnd.n6563 gnd.n6562 585
R8329 gnd.n393 gnd.n392 585
R8330 gnd.n392 gnd.n391 585
R8331 gnd.n6557 gnd.n6556 585
R8332 gnd.n6556 gnd.n6555 585
R8333 gnd.n396 gnd.n395 585
R8334 gnd.n6554 gnd.n396 585
R8335 gnd.n6552 gnd.n6551 585
R8336 gnd.n6553 gnd.n6552 585
R8337 gnd.n399 gnd.n398 585
R8338 gnd.n398 gnd.n397 585
R8339 gnd.n6547 gnd.n6546 585
R8340 gnd.n6546 gnd.n6545 585
R8341 gnd.n402 gnd.n401 585
R8342 gnd.n6544 gnd.n402 585
R8343 gnd.n6542 gnd.n6541 585
R8344 gnd.n6543 gnd.n6542 585
R8345 gnd.n405 gnd.n404 585
R8346 gnd.n404 gnd.n403 585
R8347 gnd.n5853 gnd.n5852 585
R8348 gnd.n5854 gnd.n5853 585
R8349 gnd.n982 gnd.n981 585
R8350 gnd.n4301 gnd.n982 585
R8351 gnd.n5862 gnd.n5861 585
R8352 gnd.n5861 gnd.n5860 585
R8353 gnd.n5863 gnd.n976 585
R8354 gnd.n4005 gnd.n976 585
R8355 gnd.n5865 gnd.n5864 585
R8356 gnd.n5866 gnd.n5865 585
R8357 gnd.n961 gnd.n960 585
R8358 gnd.n3996 gnd.n961 585
R8359 gnd.n5874 gnd.n5873 585
R8360 gnd.n5873 gnd.n5872 585
R8361 gnd.n5875 gnd.n955 585
R8362 gnd.n3992 gnd.n955 585
R8363 gnd.n5877 gnd.n5876 585
R8364 gnd.n5878 gnd.n5877 585
R8365 gnd.n939 gnd.n938 585
R8366 gnd.n3985 gnd.n939 585
R8367 gnd.n5886 gnd.n5885 585
R8368 gnd.n5885 gnd.n5884 585
R8369 gnd.n5887 gnd.n933 585
R8370 gnd.n4022 gnd.n933 585
R8371 gnd.n5889 gnd.n5888 585
R8372 gnd.n5890 gnd.n5889 585
R8373 gnd.n920 gnd.n919 585
R8374 gnd.n3977 gnd.n920 585
R8375 gnd.n5898 gnd.n5897 585
R8376 gnd.n5897 gnd.n5896 585
R8377 gnd.n5899 gnd.n914 585
R8378 gnd.n3969 gnd.n914 585
R8379 gnd.n5901 gnd.n5900 585
R8380 gnd.n5902 gnd.n5901 585
R8381 gnd.n915 gnd.n913 585
R8382 gnd.n3956 gnd.n913 585
R8383 gnd.n3938 gnd.n3937 585
R8384 gnd.n3937 gnd.n2014 585
R8385 gnd.n3939 gnd.n2024 585
R8386 gnd.n3948 gnd.n2024 585
R8387 gnd.n3941 gnd.n3940 585
R8388 gnd.n3942 gnd.n3941 585
R8389 gnd.n2031 gnd.n2030 585
R8390 gnd.n3928 gnd.n2030 585
R8391 gnd.n3916 gnd.n3915 585
R8392 gnd.n3917 gnd.n3916 585
R8393 gnd.n3914 gnd.n3910 585
R8394 gnd.n3920 gnd.n3910 585
R8395 gnd.n893 gnd.n892 585
R8396 gnd.n3893 gnd.n893 585
R8397 gnd.n5912 gnd.n5911 585
R8398 gnd.n5911 gnd.n5910 585
R8399 gnd.n5913 gnd.n887 585
R8400 gnd.n3883 gnd.n887 585
R8401 gnd.n5915 gnd.n5914 585
R8402 gnd.n5916 gnd.n5915 585
R8403 gnd.n872 gnd.n871 585
R8404 gnd.n3873 gnd.n872 585
R8405 gnd.n5924 gnd.n5923 585
R8406 gnd.n5923 gnd.n5922 585
R8407 gnd.n5925 gnd.n866 585
R8408 gnd.n3839 gnd.n866 585
R8409 gnd.n5927 gnd.n5926 585
R8410 gnd.n5928 gnd.n5927 585
R8411 gnd.n851 gnd.n850 585
R8412 gnd.n3845 gnd.n851 585
R8413 gnd.n5936 gnd.n5935 585
R8414 gnd.n5935 gnd.n5934 585
R8415 gnd.n5937 gnd.n845 585
R8416 gnd.n3825 gnd.n845 585
R8417 gnd.n5939 gnd.n5938 585
R8418 gnd.n5940 gnd.n5939 585
R8419 gnd.n846 gnd.n844 585
R8420 gnd.n844 gnd.n830 585
R8421 gnd.n3794 gnd.n831 585
R8422 gnd.n5946 gnd.n831 585
R8423 gnd.n3796 gnd.n3795 585
R8424 gnd.n3795 gnd.n827 585
R8425 gnd.n3797 gnd.n2089 585
R8426 gnd.n3812 gnd.n2089 585
R8427 gnd.n2101 gnd.n2099 585
R8428 gnd.n2099 gnd.n2087 585
R8429 gnd.n3802 gnd.n3801 585
R8430 gnd.n3803 gnd.n3802 585
R8431 gnd.n2100 gnd.n2098 585
R8432 gnd.n2098 gnd.n2095 585
R8433 gnd.n3788 gnd.n3787 585
R8434 gnd.n2104 gnd.n2103 585
R8435 gnd.n3596 gnd.n3595 585
R8436 gnd.n3598 gnd.n3597 585
R8437 gnd.n3600 gnd.n3599 585
R8438 gnd.n3604 gnd.n3592 585
R8439 gnd.n3606 gnd.n3605 585
R8440 gnd.n3608 gnd.n3607 585
R8441 gnd.n3610 gnd.n3609 585
R8442 gnd.n3614 gnd.n3590 585
R8443 gnd.n3616 gnd.n3615 585
R8444 gnd.n3618 gnd.n3617 585
R8445 gnd.n3620 gnd.n3619 585
R8446 gnd.n3624 gnd.n3588 585
R8447 gnd.n3626 gnd.n3625 585
R8448 gnd.n3628 gnd.n3627 585
R8449 gnd.n3630 gnd.n3629 585
R8450 gnd.n3586 gnd.n3582 585
R8451 gnd.n3642 gnd.n3641 585
R8452 gnd.n3785 gnd.n3642 585
R8453 gnd.n4142 gnd.n4141 585
R8454 gnd.n4139 gnd.n4133 585
R8455 gnd.n4149 gnd.n4130 585
R8456 gnd.n4150 gnd.n4128 585
R8457 gnd.n4127 gnd.n4120 585
R8458 gnd.n4157 gnd.n4119 585
R8459 gnd.n4158 gnd.n4118 585
R8460 gnd.n4116 gnd.n4108 585
R8461 gnd.n4165 gnd.n4107 585
R8462 gnd.n4166 gnd.n4105 585
R8463 gnd.n4104 gnd.n4097 585
R8464 gnd.n4173 gnd.n4096 585
R8465 gnd.n4174 gnd.n4095 585
R8466 gnd.n4093 gnd.n4086 585
R8467 gnd.n4181 gnd.n4085 585
R8468 gnd.n4182 gnd.n4083 585
R8469 gnd.n4082 gnd.n4078 585
R8470 gnd.n4080 gnd.n4079 585
R8471 gnd.n999 gnd.n997 585
R8472 gnd.n1870 gnd.n997 585
R8473 gnd.n1906 gnd.n995 585
R8474 gnd.n5854 gnd.n995 585
R8475 gnd.n4300 gnd.n4299 585
R8476 gnd.n4301 gnd.n4300 585
R8477 gnd.n1905 gnd.n985 585
R8478 gnd.n5860 gnd.n985 585
R8479 gnd.n4008 gnd.n4006 585
R8480 gnd.n4006 gnd.n4005 585
R8481 gnd.n4009 gnd.n974 585
R8482 gnd.n5866 gnd.n974 585
R8483 gnd.n4010 gnd.n1997 585
R8484 gnd.n3996 gnd.n1997 585
R8485 gnd.n1995 gnd.n963 585
R8486 gnd.n5872 gnd.n963 585
R8487 gnd.n4014 gnd.n1994 585
R8488 gnd.n3992 gnd.n1994 585
R8489 gnd.n4015 gnd.n953 585
R8490 gnd.n5878 gnd.n953 585
R8491 gnd.n4016 gnd.n1993 585
R8492 gnd.n3985 gnd.n1993 585
R8493 gnd.n1990 gnd.n942 585
R8494 gnd.n5884 gnd.n942 585
R8495 gnd.n4021 gnd.n4020 585
R8496 gnd.n4022 gnd.n4021 585
R8497 gnd.n1989 gnd.n932 585
R8498 gnd.n5890 gnd.n932 585
R8499 gnd.n3976 gnd.n3975 585
R8500 gnd.n3977 gnd.n3976 585
R8501 gnd.n2005 gnd.n922 585
R8502 gnd.n5896 gnd.n922 585
R8503 gnd.n3971 gnd.n3970 585
R8504 gnd.n3970 gnd.n3969 585
R8505 gnd.n2007 gnd.n911 585
R8506 gnd.n5902 gnd.n911 585
R8507 gnd.n3955 gnd.n3954 585
R8508 gnd.n3956 gnd.n3955 585
R8509 gnd.n2017 gnd.n2016 585
R8510 gnd.n2016 gnd.n2014 585
R8511 gnd.n3950 gnd.n3949 585
R8512 gnd.n3949 gnd.n3948 585
R8513 gnd.n2020 gnd.n2019 585
R8514 gnd.n3942 gnd.n2020 585
R8515 gnd.n3927 gnd.n3926 585
R8516 gnd.n3928 gnd.n3927 585
R8517 gnd.n2051 gnd.n2050 585
R8518 gnd.n3917 gnd.n2050 585
R8519 gnd.n3922 gnd.n3921 585
R8520 gnd.n3921 gnd.n3920 585
R8521 gnd.n2054 gnd.n2053 585
R8522 gnd.n3893 gnd.n2054 585
R8523 gnd.n3880 gnd.n896 585
R8524 gnd.n5910 gnd.n896 585
R8525 gnd.n3882 gnd.n3881 585
R8526 gnd.n3883 gnd.n3882 585
R8527 gnd.n2064 gnd.n885 585
R8528 gnd.n5916 gnd.n885 585
R8529 gnd.n3875 gnd.n3874 585
R8530 gnd.n3874 gnd.n3873 585
R8531 gnd.n2066 gnd.n875 585
R8532 gnd.n5922 gnd.n875 585
R8533 gnd.n3841 gnd.n3840 585
R8534 gnd.n3840 gnd.n3839 585
R8535 gnd.n3842 gnd.n864 585
R8536 gnd.n5928 gnd.n864 585
R8537 gnd.n3844 gnd.n3843 585
R8538 gnd.n3845 gnd.n3844 585
R8539 gnd.n2074 gnd.n854 585
R8540 gnd.n5934 gnd.n854 585
R8541 gnd.n3824 gnd.n3823 585
R8542 gnd.n3825 gnd.n3824 585
R8543 gnd.n2082 gnd.n842 585
R8544 gnd.n5940 gnd.n842 585
R8545 gnd.n3818 gnd.n3817 585
R8546 gnd.n3817 gnd.n830 585
R8547 gnd.n3816 gnd.n829 585
R8548 gnd.n5946 gnd.n829 585
R8549 gnd.n3815 gnd.n3814 585
R8550 gnd.n3814 gnd.n827 585
R8551 gnd.n3813 gnd.n2084 585
R8552 gnd.n3813 gnd.n3812 585
R8553 gnd.n3636 gnd.n2086 585
R8554 gnd.n2087 gnd.n2086 585
R8555 gnd.n3637 gnd.n2097 585
R8556 gnd.n3803 gnd.n2097 585
R8557 gnd.n3638 gnd.n3583 585
R8558 gnd.n3583 gnd.n2095 585
R8559 gnd.n6910 gnd.n84 585
R8560 gnd.n7006 gnd.n84 585
R8561 gnd.n6911 gnd.n6842 585
R8562 gnd.n6842 gnd.n81 585
R8563 gnd.n6912 gnd.n162 585
R8564 gnd.n6926 gnd.n162 585
R8565 gnd.n173 gnd.n171 585
R8566 gnd.n171 gnd.n161 585
R8567 gnd.n6917 gnd.n6916 585
R8568 gnd.n6918 gnd.n6917 585
R8569 gnd.n172 gnd.n170 585
R8570 gnd.n180 gnd.n170 585
R8571 gnd.n6838 gnd.n6837 585
R8572 gnd.n6837 gnd.n6836 585
R8573 gnd.n176 gnd.n175 585
R8574 gnd.n261 gnd.n176 585
R8575 gnd.n6827 gnd.n6826 585
R8576 gnd.n6828 gnd.n6827 585
R8577 gnd.n190 gnd.n189 585
R8578 gnd.n266 gnd.n189 585
R8579 gnd.n6822 gnd.n6821 585
R8580 gnd.n6821 gnd.n6820 585
R8581 gnd.n193 gnd.n192 585
R8582 gnd.n6763 gnd.n193 585
R8583 gnd.n6811 gnd.n6810 585
R8584 gnd.n6812 gnd.n6811 585
R8585 gnd.n205 gnd.n204 585
R8586 gnd.n6768 gnd.n204 585
R8587 gnd.n6806 gnd.n6805 585
R8588 gnd.n6805 gnd.n6804 585
R8589 gnd.n208 gnd.n207 585
R8590 gnd.n6772 gnd.n208 585
R8591 gnd.n6795 gnd.n6794 585
R8592 gnd.n6796 gnd.n6795 585
R8593 gnd.n227 gnd.n226 585
R8594 gnd.n6777 gnd.n226 585
R8595 gnd.n6790 gnd.n6789 585
R8596 gnd.n6789 gnd.n6788 585
R8597 gnd.n230 gnd.n229 585
R8598 gnd.n6783 gnd.n230 585
R8599 gnd.n5669 gnd.n5667 585
R8600 gnd.n5667 gnd.n5666 585
R8601 gnd.n5670 gnd.n1169 585
R8602 gnd.n1170 gnd.n1169 585
R8603 gnd.n5671 gnd.n1168 585
R8604 gnd.n5638 gnd.n1168 585
R8605 gnd.n1175 gnd.n1166 585
R8606 gnd.n1176 gnd.n1175 585
R8607 gnd.n5675 gnd.n1165 585
R8608 gnd.n5629 gnd.n1165 585
R8609 gnd.n5676 gnd.n1164 585
R8610 gnd.n5506 gnd.n1164 585
R8611 gnd.n5677 gnd.n1163 585
R8612 gnd.n5619 gnd.n1163 585
R8613 gnd.n1204 gnd.n1161 585
R8614 gnd.n1205 gnd.n1204 585
R8615 gnd.n5681 gnd.n1160 585
R8616 gnd.n5613 gnd.n1160 585
R8617 gnd.n5682 gnd.n1159 585
R8618 gnd.n5595 gnd.n1159 585
R8619 gnd.n5683 gnd.n1158 585
R8620 gnd.n1212 gnd.n1158 585
R8621 gnd.n1223 gnd.n1156 585
R8622 gnd.n5586 gnd.n1223 585
R8623 gnd.n5687 gnd.n1155 585
R8624 gnd.n1233 gnd.n1155 585
R8625 gnd.n5688 gnd.n1154 585
R8626 gnd.n5575 gnd.n1154 585
R8627 gnd.n5689 gnd.n1153 585
R8628 gnd.n5563 gnd.n1153 585
R8629 gnd.n1240 gnd.n1151 585
R8630 gnd.n1241 gnd.n1240 585
R8631 gnd.n5693 gnd.n1150 585
R8632 gnd.n5554 gnd.n1150 585
R8633 gnd.n5694 gnd.n1149 585
R8634 gnd.n5526 gnd.n1149 585
R8635 gnd.n5695 gnd.n1148 585
R8636 gnd.n5544 gnd.n1148 585
R8637 gnd.n1145 gnd.n1143 585
R8638 gnd.n5477 gnd.n1143 585
R8639 gnd.n5700 gnd.n5699 585
R8640 gnd.n5701 gnd.n5700 585
R8641 gnd.n1144 gnd.n1142 585
R8642 gnd.n5468 gnd.n1142 585
R8643 gnd.n5026 gnd.n1130 585
R8644 gnd.n5707 gnd.n1130 585
R8645 gnd.n5030 gnd.n5029 585
R8646 gnd.n5032 gnd.n5023 585
R8647 gnd.n5035 gnd.n5034 585
R8648 gnd.n5016 gnd.n5015 585
R8649 gnd.n5049 gnd.n5048 585
R8650 gnd.n5051 gnd.n5014 585
R8651 gnd.n5054 gnd.n5053 585
R8652 gnd.n5007 gnd.n5006 585
R8653 gnd.n5068 gnd.n5067 585
R8654 gnd.n5070 gnd.n5005 585
R8655 gnd.n5073 gnd.n5072 585
R8656 gnd.n4998 gnd.n4997 585
R8657 gnd.n5087 gnd.n5086 585
R8658 gnd.n5089 gnd.n4996 585
R8659 gnd.n5092 gnd.n5091 585
R8660 gnd.n4989 gnd.n4988 585
R8661 gnd.n5108 gnd.n5107 585
R8662 gnd.n5110 gnd.n4987 585
R8663 gnd.n5112 gnd.n5111 585
R8664 gnd.n5111 gnd.n1118 585
R8665 gnd.n6881 gnd.n80 585
R8666 gnd.n6882 gnd.n6880 585
R8667 gnd.n6883 gnd.n6876 585
R8668 gnd.n6874 gnd.n6872 585
R8669 gnd.n6887 gnd.n6871 585
R8670 gnd.n6888 gnd.n6869 585
R8671 gnd.n6889 gnd.n6868 585
R8672 gnd.n6866 gnd.n6864 585
R8673 gnd.n6893 gnd.n6863 585
R8674 gnd.n6894 gnd.n6861 585
R8675 gnd.n6895 gnd.n6860 585
R8676 gnd.n6858 gnd.n6856 585
R8677 gnd.n6899 gnd.n6855 585
R8678 gnd.n6900 gnd.n6853 585
R8679 gnd.n6901 gnd.n6852 585
R8680 gnd.n6850 gnd.n6848 585
R8681 gnd.n6905 gnd.n6847 585
R8682 gnd.n6906 gnd.n6845 585
R8683 gnd.n6907 gnd.n6844 585
R8684 gnd.n6844 gnd.n83 585
R8685 gnd.n7008 gnd.n7007 585
R8686 gnd.n7007 gnd.n7006 585
R8687 gnd.n79 gnd.n77 585
R8688 gnd.n81 gnd.n79 585
R8689 gnd.n7012 gnd.n76 585
R8690 gnd.n6926 gnd.n76 585
R8691 gnd.n7013 gnd.n75 585
R8692 gnd.n161 gnd.n75 585
R8693 gnd.n7014 gnd.n74 585
R8694 gnd.n6918 gnd.n74 585
R8695 gnd.n179 gnd.n72 585
R8696 gnd.n180 gnd.n179 585
R8697 gnd.n7018 gnd.n71 585
R8698 gnd.n6836 gnd.n71 585
R8699 gnd.n7019 gnd.n70 585
R8700 gnd.n261 gnd.n70 585
R8701 gnd.n7020 gnd.n69 585
R8702 gnd.n6828 gnd.n69 585
R8703 gnd.n265 gnd.n67 585
R8704 gnd.n266 gnd.n265 585
R8705 gnd.n7024 gnd.n66 585
R8706 gnd.n6820 gnd.n66 585
R8707 gnd.n7025 gnd.n65 585
R8708 gnd.n6763 gnd.n65 585
R8709 gnd.n7026 gnd.n64 585
R8710 gnd.n6812 gnd.n64 585
R8711 gnd.n6767 gnd.n62 585
R8712 gnd.n6768 gnd.n6767 585
R8713 gnd.n7030 gnd.n61 585
R8714 gnd.n6804 gnd.n61 585
R8715 gnd.n7031 gnd.n60 585
R8716 gnd.n6772 gnd.n60 585
R8717 gnd.n7032 gnd.n59 585
R8718 gnd.n6796 gnd.n59 585
R8719 gnd.n6776 gnd.n57 585
R8720 gnd.n6777 gnd.n6776 585
R8721 gnd.n7036 gnd.n56 585
R8722 gnd.n6788 gnd.n56 585
R8723 gnd.n7037 gnd.n55 585
R8724 gnd.n6783 gnd.n55 585
R8725 gnd.n7038 gnd.n54 585
R8726 gnd.n5666 gnd.n54 585
R8727 gnd.n1178 gnd.n52 585
R8728 gnd.n1178 gnd.n1170 585
R8729 gnd.n1189 gnd.n1179 585
R8730 gnd.n5638 gnd.n1179 585
R8731 gnd.n1190 gnd.n1187 585
R8732 gnd.n1187 gnd.n1176 585
R8733 gnd.n5627 gnd.n5626 585
R8734 gnd.n5629 gnd.n5627 585
R8735 gnd.n1188 gnd.n1186 585
R8736 gnd.n5506 gnd.n1186 585
R8737 gnd.n5621 gnd.n5620 585
R8738 gnd.n5620 gnd.n5619 585
R8739 gnd.n1193 gnd.n1192 585
R8740 gnd.n1205 gnd.n1193 585
R8741 gnd.n1216 gnd.n1203 585
R8742 gnd.n5613 gnd.n1203 585
R8743 gnd.n5594 gnd.n5593 585
R8744 gnd.n5595 gnd.n5594 585
R8745 gnd.n1215 gnd.n1214 585
R8746 gnd.n1214 gnd.n1212 585
R8747 gnd.n5588 gnd.n5587 585
R8748 gnd.n5587 gnd.n5586 585
R8749 gnd.n1219 gnd.n1218 585
R8750 gnd.n1233 gnd.n1219 585
R8751 gnd.n1245 gnd.n1232 585
R8752 gnd.n5575 gnd.n1232 585
R8753 gnd.n5562 gnd.n5561 585
R8754 gnd.n5563 gnd.n5562 585
R8755 gnd.n1244 gnd.n1243 585
R8756 gnd.n1243 gnd.n1241 585
R8757 gnd.n5556 gnd.n5555 585
R8758 gnd.n5555 gnd.n5554 585
R8759 gnd.n1248 gnd.n1247 585
R8760 gnd.n5526 gnd.n1248 585
R8761 gnd.n1263 gnd.n1258 585
R8762 gnd.n5544 gnd.n1258 585
R8763 gnd.n5476 gnd.n5475 585
R8764 gnd.n5477 gnd.n5476 585
R8765 gnd.n1262 gnd.n1140 585
R8766 gnd.n5701 gnd.n1140 585
R8767 gnd.n5470 gnd.n5469 585
R8768 gnd.n5469 gnd.n5468 585
R8769 gnd.n1265 gnd.n1128 585
R8770 gnd.n5707 gnd.n1128 585
R8771 gnd.n3463 gnd.n3462 585
R8772 gnd.n3464 gnd.n3463 585
R8773 gnd.n2181 gnd.n2180 585
R8774 gnd.n2187 gnd.n2180 585
R8775 gnd.n3438 gnd.n2199 585
R8776 gnd.n2199 gnd.n2186 585
R8777 gnd.n3440 gnd.n3439 585
R8778 gnd.n3441 gnd.n3440 585
R8779 gnd.n2200 gnd.n2198 585
R8780 gnd.n2198 gnd.n2194 585
R8781 gnd.n3172 gnd.n3171 585
R8782 gnd.n3171 gnd.n3170 585
R8783 gnd.n2205 gnd.n2204 585
R8784 gnd.n3141 gnd.n2205 585
R8785 gnd.n3161 gnd.n3160 585
R8786 gnd.n3160 gnd.n3159 585
R8787 gnd.n2212 gnd.n2211 585
R8788 gnd.n3147 gnd.n2212 585
R8789 gnd.n3117 gnd.n2232 585
R8790 gnd.n2232 gnd.n2231 585
R8791 gnd.n3119 gnd.n3118 585
R8792 gnd.n3120 gnd.n3119 585
R8793 gnd.n2233 gnd.n2230 585
R8794 gnd.n2241 gnd.n2230 585
R8795 gnd.n3095 gnd.n2253 585
R8796 gnd.n2253 gnd.n2240 585
R8797 gnd.n3097 gnd.n3096 585
R8798 gnd.n3098 gnd.n3097 585
R8799 gnd.n2254 gnd.n2252 585
R8800 gnd.n2252 gnd.n2248 585
R8801 gnd.n3083 gnd.n3082 585
R8802 gnd.n3082 gnd.n3081 585
R8803 gnd.n2259 gnd.n2258 585
R8804 gnd.n2269 gnd.n2259 585
R8805 gnd.n3071 gnd.n3070 585
R8806 gnd.n3070 gnd.n3069 585
R8807 gnd.n2266 gnd.n2265 585
R8808 gnd.n3057 gnd.n2266 585
R8809 gnd.n3031 gnd.n2287 585
R8810 gnd.n2287 gnd.n2276 585
R8811 gnd.n3033 gnd.n3032 585
R8812 gnd.n3034 gnd.n3033 585
R8813 gnd.n2288 gnd.n2286 585
R8814 gnd.n2296 gnd.n2286 585
R8815 gnd.n3009 gnd.n2308 585
R8816 gnd.n2308 gnd.n2295 585
R8817 gnd.n3011 gnd.n3010 585
R8818 gnd.n3012 gnd.n3011 585
R8819 gnd.n2309 gnd.n2307 585
R8820 gnd.n2307 gnd.n2303 585
R8821 gnd.n2997 gnd.n2996 585
R8822 gnd.n2996 gnd.n2995 585
R8823 gnd.n2314 gnd.n2313 585
R8824 gnd.n2323 gnd.n2314 585
R8825 gnd.n2986 gnd.n2985 585
R8826 gnd.n2985 gnd.n2984 585
R8827 gnd.n2321 gnd.n2320 585
R8828 gnd.n2972 gnd.n2321 585
R8829 gnd.n2410 gnd.n2409 585
R8830 gnd.n2410 gnd.n2330 585
R8831 gnd.n2929 gnd.n2928 585
R8832 gnd.n2928 gnd.n2927 585
R8833 gnd.n2930 gnd.n2404 585
R8834 gnd.n2415 gnd.n2404 585
R8835 gnd.n2932 gnd.n2931 585
R8836 gnd.n2933 gnd.n2932 585
R8837 gnd.n2405 gnd.n2403 585
R8838 gnd.n2428 gnd.n2403 585
R8839 gnd.n2388 gnd.n2387 585
R8840 gnd.n2391 gnd.n2388 585
R8841 gnd.n2943 gnd.n2942 585
R8842 gnd.n2942 gnd.n2941 585
R8843 gnd.n2944 gnd.n2382 585
R8844 gnd.n2903 gnd.n2382 585
R8845 gnd.n2946 gnd.n2945 585
R8846 gnd.n2947 gnd.n2946 585
R8847 gnd.n2383 gnd.n2381 585
R8848 gnd.n2442 gnd.n2381 585
R8849 gnd.n2895 gnd.n2894 585
R8850 gnd.n2894 gnd.n2893 585
R8851 gnd.n2439 gnd.n2438 585
R8852 gnd.n2877 gnd.n2439 585
R8853 gnd.n2864 gnd.n2458 585
R8854 gnd.n2458 gnd.n2457 585
R8855 gnd.n2866 gnd.n2865 585
R8856 gnd.n2867 gnd.n2866 585
R8857 gnd.n2459 gnd.n2456 585
R8858 gnd.n2465 gnd.n2456 585
R8859 gnd.n2845 gnd.n2844 585
R8860 gnd.n2846 gnd.n2845 585
R8861 gnd.n2476 gnd.n2475 585
R8862 gnd.n2475 gnd.n2471 585
R8863 gnd.n2835 gnd.n2834 585
R8864 gnd.n2836 gnd.n2835 585
R8865 gnd.n2486 gnd.n2485 585
R8866 gnd.n2491 gnd.n2485 585
R8867 gnd.n2813 gnd.n2504 585
R8868 gnd.n2504 gnd.n2490 585
R8869 gnd.n2815 gnd.n2814 585
R8870 gnd.n2816 gnd.n2815 585
R8871 gnd.n2505 gnd.n2503 585
R8872 gnd.n2503 gnd.n2499 585
R8873 gnd.n2804 gnd.n2803 585
R8874 gnd.n2805 gnd.n2804 585
R8875 gnd.n2512 gnd.n2511 585
R8876 gnd.n2516 gnd.n2511 585
R8877 gnd.n2781 gnd.n2533 585
R8878 gnd.n2533 gnd.n2515 585
R8879 gnd.n2783 gnd.n2782 585
R8880 gnd.n2784 gnd.n2783 585
R8881 gnd.n2534 gnd.n2532 585
R8882 gnd.n2532 gnd.n2523 585
R8883 gnd.n2776 gnd.n2775 585
R8884 gnd.n2775 gnd.n2774 585
R8885 gnd.n2581 gnd.n2580 585
R8886 gnd.n2582 gnd.n2581 585
R8887 gnd.n2735 gnd.n2734 585
R8888 gnd.n2736 gnd.n2735 585
R8889 gnd.n2591 gnd.n2590 585
R8890 gnd.n2590 gnd.n2589 585
R8891 gnd.n2730 gnd.n2729 585
R8892 gnd.n2729 gnd.n2728 585
R8893 gnd.n2594 gnd.n2593 585
R8894 gnd.n2595 gnd.n2594 585
R8895 gnd.n2719 gnd.n2718 585
R8896 gnd.n2720 gnd.n2719 585
R8897 gnd.n2602 gnd.n2601 585
R8898 gnd.n2711 gnd.n2601 585
R8899 gnd.n2714 gnd.n2713 585
R8900 gnd.n2713 gnd.n2712 585
R8901 gnd.n2605 gnd.n2604 585
R8902 gnd.n2606 gnd.n2605 585
R8903 gnd.n2700 gnd.n2699 585
R8904 gnd.n2698 gnd.n2624 585
R8905 gnd.n2697 gnd.n2623 585
R8906 gnd.n2702 gnd.n2623 585
R8907 gnd.n2696 gnd.n2695 585
R8908 gnd.n2694 gnd.n2693 585
R8909 gnd.n2692 gnd.n2691 585
R8910 gnd.n2690 gnd.n2689 585
R8911 gnd.n2688 gnd.n2687 585
R8912 gnd.n2686 gnd.n2685 585
R8913 gnd.n2684 gnd.n2683 585
R8914 gnd.n2682 gnd.n2681 585
R8915 gnd.n2680 gnd.n2679 585
R8916 gnd.n2678 gnd.n2677 585
R8917 gnd.n2676 gnd.n2675 585
R8918 gnd.n2674 gnd.n2673 585
R8919 gnd.n2672 gnd.n2671 585
R8920 gnd.n2670 gnd.n2669 585
R8921 gnd.n2668 gnd.n2667 585
R8922 gnd.n2666 gnd.n2665 585
R8923 gnd.n2664 gnd.n2663 585
R8924 gnd.n2662 gnd.n2661 585
R8925 gnd.n2660 gnd.n2659 585
R8926 gnd.n2658 gnd.n2657 585
R8927 gnd.n2656 gnd.n2655 585
R8928 gnd.n2654 gnd.n2653 585
R8929 gnd.n2611 gnd.n2610 585
R8930 gnd.n2705 gnd.n2704 585
R8931 gnd.n3467 gnd.n3466 585
R8932 gnd.n3469 gnd.n3468 585
R8933 gnd.n3471 gnd.n3470 585
R8934 gnd.n3473 gnd.n3472 585
R8935 gnd.n3475 gnd.n3474 585
R8936 gnd.n3477 gnd.n3476 585
R8937 gnd.n3479 gnd.n3478 585
R8938 gnd.n3481 gnd.n3480 585
R8939 gnd.n3483 gnd.n3482 585
R8940 gnd.n3485 gnd.n3484 585
R8941 gnd.n3487 gnd.n3486 585
R8942 gnd.n3489 gnd.n3488 585
R8943 gnd.n3491 gnd.n3490 585
R8944 gnd.n3493 gnd.n3492 585
R8945 gnd.n3495 gnd.n3494 585
R8946 gnd.n3497 gnd.n3496 585
R8947 gnd.n3499 gnd.n3498 585
R8948 gnd.n3501 gnd.n3500 585
R8949 gnd.n3503 gnd.n3502 585
R8950 gnd.n3505 gnd.n3504 585
R8951 gnd.n3507 gnd.n3506 585
R8952 gnd.n3509 gnd.n3508 585
R8953 gnd.n3511 gnd.n3510 585
R8954 gnd.n3513 gnd.n3512 585
R8955 gnd.n3515 gnd.n3514 585
R8956 gnd.n3516 gnd.n2148 585
R8957 gnd.n3517 gnd.n2106 585
R8958 gnd.n3555 gnd.n2106 585
R8959 gnd.n3465 gnd.n2178 585
R8960 gnd.n3465 gnd.n3464 585
R8961 gnd.n3134 gnd.n2177 585
R8962 gnd.n2187 gnd.n2177 585
R8963 gnd.n3136 gnd.n3135 585
R8964 gnd.n3135 gnd.n2186 585
R8965 gnd.n3137 gnd.n2196 585
R8966 gnd.n3441 gnd.n2196 585
R8967 gnd.n3139 gnd.n3138 585
R8968 gnd.n3138 gnd.n2194 585
R8969 gnd.n3140 gnd.n2207 585
R8970 gnd.n3170 gnd.n2207 585
R8971 gnd.n3143 gnd.n3142 585
R8972 gnd.n3142 gnd.n3141 585
R8973 gnd.n3144 gnd.n2214 585
R8974 gnd.n3159 gnd.n2214 585
R8975 gnd.n3146 gnd.n3145 585
R8976 gnd.n3147 gnd.n3146 585
R8977 gnd.n2224 gnd.n2223 585
R8978 gnd.n2231 gnd.n2223 585
R8979 gnd.n3122 gnd.n3121 585
R8980 gnd.n3121 gnd.n3120 585
R8981 gnd.n2227 gnd.n2226 585
R8982 gnd.n2241 gnd.n2227 585
R8983 gnd.n3047 gnd.n3046 585
R8984 gnd.n3046 gnd.n2240 585
R8985 gnd.n3048 gnd.n2250 585
R8986 gnd.n3098 gnd.n2250 585
R8987 gnd.n3050 gnd.n3049 585
R8988 gnd.n3049 gnd.n2248 585
R8989 gnd.n3051 gnd.n2261 585
R8990 gnd.n3081 gnd.n2261 585
R8991 gnd.n3053 gnd.n3052 585
R8992 gnd.n3052 gnd.n2269 585
R8993 gnd.n3054 gnd.n2268 585
R8994 gnd.n3069 gnd.n2268 585
R8995 gnd.n3056 gnd.n3055 585
R8996 gnd.n3057 gnd.n3056 585
R8997 gnd.n2280 gnd.n2279 585
R8998 gnd.n2279 gnd.n2276 585
R8999 gnd.n3036 gnd.n3035 585
R9000 gnd.n3035 gnd.n3034 585
R9001 gnd.n2283 gnd.n2282 585
R9002 gnd.n2296 gnd.n2283 585
R9003 gnd.n2960 gnd.n2959 585
R9004 gnd.n2959 gnd.n2295 585
R9005 gnd.n2961 gnd.n2305 585
R9006 gnd.n3012 gnd.n2305 585
R9007 gnd.n2963 gnd.n2962 585
R9008 gnd.n2962 gnd.n2303 585
R9009 gnd.n2964 gnd.n2316 585
R9010 gnd.n2995 gnd.n2316 585
R9011 gnd.n2966 gnd.n2965 585
R9012 gnd.n2965 gnd.n2323 585
R9013 gnd.n2967 gnd.n2322 585
R9014 gnd.n2984 gnd.n2322 585
R9015 gnd.n2969 gnd.n2968 585
R9016 gnd.n2972 gnd.n2969 585
R9017 gnd.n2333 gnd.n2332 585
R9018 gnd.n2332 gnd.n2330 585
R9019 gnd.n2412 gnd.n2411 585
R9020 gnd.n2927 gnd.n2411 585
R9021 gnd.n2414 gnd.n2413 585
R9022 gnd.n2415 gnd.n2414 585
R9023 gnd.n2425 gnd.n2401 585
R9024 gnd.n2933 gnd.n2401 585
R9025 gnd.n2427 gnd.n2426 585
R9026 gnd.n2428 gnd.n2427 585
R9027 gnd.n2424 gnd.n2423 585
R9028 gnd.n2424 gnd.n2391 585
R9029 gnd.n2422 gnd.n2389 585
R9030 gnd.n2941 gnd.n2389 585
R9031 gnd.n2378 gnd.n2376 585
R9032 gnd.n2903 gnd.n2378 585
R9033 gnd.n2949 gnd.n2948 585
R9034 gnd.n2948 gnd.n2947 585
R9035 gnd.n2377 gnd.n2375 585
R9036 gnd.n2442 gnd.n2377 585
R9037 gnd.n2874 gnd.n2441 585
R9038 gnd.n2893 gnd.n2441 585
R9039 gnd.n2876 gnd.n2875 585
R9040 gnd.n2877 gnd.n2876 585
R9041 gnd.n2451 gnd.n2450 585
R9042 gnd.n2457 gnd.n2450 585
R9043 gnd.n2869 gnd.n2868 585
R9044 gnd.n2868 gnd.n2867 585
R9045 gnd.n2454 gnd.n2453 585
R9046 gnd.n2465 gnd.n2454 585
R9047 gnd.n2754 gnd.n2473 585
R9048 gnd.n2846 gnd.n2473 585
R9049 gnd.n2756 gnd.n2755 585
R9050 gnd.n2755 gnd.n2471 585
R9051 gnd.n2757 gnd.n2484 585
R9052 gnd.n2836 gnd.n2484 585
R9053 gnd.n2759 gnd.n2758 585
R9054 gnd.n2759 gnd.n2491 585
R9055 gnd.n2761 gnd.n2760 585
R9056 gnd.n2760 gnd.n2490 585
R9057 gnd.n2762 gnd.n2501 585
R9058 gnd.n2816 gnd.n2501 585
R9059 gnd.n2764 gnd.n2763 585
R9060 gnd.n2763 gnd.n2499 585
R9061 gnd.n2765 gnd.n2510 585
R9062 gnd.n2805 gnd.n2510 585
R9063 gnd.n2767 gnd.n2766 585
R9064 gnd.n2767 gnd.n2516 585
R9065 gnd.n2769 gnd.n2768 585
R9066 gnd.n2768 gnd.n2515 585
R9067 gnd.n2770 gnd.n2531 585
R9068 gnd.n2784 gnd.n2531 585
R9069 gnd.n2771 gnd.n2584 585
R9070 gnd.n2584 gnd.n2523 585
R9071 gnd.n2773 gnd.n2772 585
R9072 gnd.n2774 gnd.n2773 585
R9073 gnd.n2585 gnd.n2583 585
R9074 gnd.n2583 gnd.n2582 585
R9075 gnd.n2738 gnd.n2737 585
R9076 gnd.n2737 gnd.n2736 585
R9077 gnd.n2588 gnd.n2587 585
R9078 gnd.n2589 gnd.n2588 585
R9079 gnd.n2727 gnd.n2726 585
R9080 gnd.n2728 gnd.n2727 585
R9081 gnd.n2597 gnd.n2596 585
R9082 gnd.n2596 gnd.n2595 585
R9083 gnd.n2722 gnd.n2721 585
R9084 gnd.n2721 gnd.n2720 585
R9085 gnd.n2600 gnd.n2599 585
R9086 gnd.n2711 gnd.n2600 585
R9087 gnd.n2710 gnd.n2709 585
R9088 gnd.n2712 gnd.n2710 585
R9089 gnd.n2608 gnd.n2607 585
R9090 gnd.n2607 gnd.n2606 585
R9091 gnd.n3450 gnd.n2128 585
R9092 gnd.n2128 gnd.n2105 585
R9093 gnd.n3451 gnd.n2189 585
R9094 gnd.n2189 gnd.n2179 585
R9095 gnd.n3453 gnd.n3452 585
R9096 gnd.n3454 gnd.n3453 585
R9097 gnd.n2190 gnd.n2188 585
R9098 gnd.n2197 gnd.n2188 585
R9099 gnd.n3444 gnd.n3443 585
R9100 gnd.n3443 gnd.n3442 585
R9101 gnd.n2193 gnd.n2192 585
R9102 gnd.n3169 gnd.n2193 585
R9103 gnd.n3155 gnd.n2216 585
R9104 gnd.n2216 gnd.n2206 585
R9105 gnd.n3157 gnd.n3156 585
R9106 gnd.n3158 gnd.n3157 585
R9107 gnd.n2217 gnd.n2215 585
R9108 gnd.n2215 gnd.n2213 585
R9109 gnd.n3150 gnd.n3149 585
R9110 gnd.n3149 gnd.n3148 585
R9111 gnd.n2220 gnd.n2219 585
R9112 gnd.n2229 gnd.n2220 585
R9113 gnd.n3106 gnd.n2243 585
R9114 gnd.n2243 gnd.n2228 585
R9115 gnd.n3108 gnd.n3107 585
R9116 gnd.n3109 gnd.n3108 585
R9117 gnd.n2244 gnd.n2242 585
R9118 gnd.n2251 gnd.n2242 585
R9119 gnd.n3101 gnd.n3100 585
R9120 gnd.n3100 gnd.n3099 585
R9121 gnd.n2247 gnd.n2246 585
R9122 gnd.n3080 gnd.n2247 585
R9123 gnd.n3065 gnd.n2271 585
R9124 gnd.n2271 gnd.n2260 585
R9125 gnd.n3067 gnd.n3066 585
R9126 gnd.n3068 gnd.n3067 585
R9127 gnd.n2272 gnd.n2270 585
R9128 gnd.n2270 gnd.n2267 585
R9129 gnd.n3060 gnd.n3059 585
R9130 gnd.n3059 gnd.n3058 585
R9131 gnd.n2275 gnd.n2274 585
R9132 gnd.n2285 gnd.n2275 585
R9133 gnd.n3020 gnd.n2298 585
R9134 gnd.n2298 gnd.n2284 585
R9135 gnd.n3022 gnd.n3021 585
R9136 gnd.n3023 gnd.n3022 585
R9137 gnd.n2299 gnd.n2297 585
R9138 gnd.n2306 gnd.n2297 585
R9139 gnd.n3015 gnd.n3014 585
R9140 gnd.n3014 gnd.n3013 585
R9141 gnd.n2302 gnd.n2301 585
R9142 gnd.n2994 gnd.n2302 585
R9143 gnd.n2980 gnd.n2325 585
R9144 gnd.n2325 gnd.n2315 585
R9145 gnd.n2982 gnd.n2981 585
R9146 gnd.n2983 gnd.n2982 585
R9147 gnd.n2326 gnd.n2324 585
R9148 gnd.n2971 gnd.n2324 585
R9149 gnd.n2975 gnd.n2974 585
R9150 gnd.n2974 gnd.n2973 585
R9151 gnd.n2329 gnd.n2328 585
R9152 gnd.n2926 gnd.n2329 585
R9153 gnd.n2419 gnd.n2418 585
R9154 gnd.n2420 gnd.n2419 585
R9155 gnd.n2399 gnd.n2398 585
R9156 gnd.n2402 gnd.n2399 585
R9157 gnd.n2936 gnd.n2935 585
R9158 gnd.n2935 gnd.n2934 585
R9159 gnd.n2937 gnd.n2393 585
R9160 gnd.n2429 gnd.n2393 585
R9161 gnd.n2939 gnd.n2938 585
R9162 gnd.n2940 gnd.n2939 585
R9163 gnd.n2394 gnd.n2392 585
R9164 gnd.n2904 gnd.n2392 585
R9165 gnd.n2888 gnd.n2887 585
R9166 gnd.n2887 gnd.n2380 585
R9167 gnd.n2889 gnd.n2444 585
R9168 gnd.n2444 gnd.n2379 585
R9169 gnd.n2891 gnd.n2890 585
R9170 gnd.n2892 gnd.n2891 585
R9171 gnd.n2445 gnd.n2443 585
R9172 gnd.n2443 gnd.n2440 585
R9173 gnd.n2880 gnd.n2879 585
R9174 gnd.n2879 gnd.n2878 585
R9175 gnd.n2448 gnd.n2447 585
R9176 gnd.n2455 gnd.n2448 585
R9177 gnd.n2854 gnd.n2853 585
R9178 gnd.n2855 gnd.n2854 585
R9179 gnd.n2467 gnd.n2466 585
R9180 gnd.n2474 gnd.n2466 585
R9181 gnd.n2849 gnd.n2848 585
R9182 gnd.n2848 gnd.n2847 585
R9183 gnd.n2470 gnd.n2469 585
R9184 gnd.n2837 gnd.n2470 585
R9185 gnd.n2824 gnd.n2494 585
R9186 gnd.n2494 gnd.n2493 585
R9187 gnd.n2826 gnd.n2825 585
R9188 gnd.n2827 gnd.n2826 585
R9189 gnd.n2495 gnd.n2492 585
R9190 gnd.n2502 gnd.n2492 585
R9191 gnd.n2819 gnd.n2818 585
R9192 gnd.n2818 gnd.n2817 585
R9193 gnd.n2498 gnd.n2497 585
R9194 gnd.n2806 gnd.n2498 585
R9195 gnd.n2793 gnd.n2519 585
R9196 gnd.n2519 gnd.n2518 585
R9197 gnd.n2795 gnd.n2794 585
R9198 gnd.n2796 gnd.n2795 585
R9199 gnd.n2789 gnd.n2517 585
R9200 gnd.n2788 gnd.n2787 585
R9201 gnd.n2522 gnd.n2521 585
R9202 gnd.n2785 gnd.n2522 585
R9203 gnd.n2544 gnd.n2543 585
R9204 gnd.n2547 gnd.n2546 585
R9205 gnd.n2545 gnd.n2540 585
R9206 gnd.n2552 gnd.n2551 585
R9207 gnd.n2554 gnd.n2553 585
R9208 gnd.n2557 gnd.n2556 585
R9209 gnd.n2555 gnd.n2538 585
R9210 gnd.n2562 gnd.n2561 585
R9211 gnd.n2564 gnd.n2563 585
R9212 gnd.n2567 gnd.n2566 585
R9213 gnd.n2565 gnd.n2536 585
R9214 gnd.n2572 gnd.n2571 585
R9215 gnd.n2576 gnd.n2573 585
R9216 gnd.n2577 gnd.n2514 585
R9217 gnd.n3456 gnd.n2143 585
R9218 gnd.n3523 gnd.n3522 585
R9219 gnd.n3525 gnd.n3524 585
R9220 gnd.n3527 gnd.n3526 585
R9221 gnd.n3529 gnd.n3528 585
R9222 gnd.n3531 gnd.n3530 585
R9223 gnd.n3533 gnd.n3532 585
R9224 gnd.n3535 gnd.n3534 585
R9225 gnd.n3537 gnd.n3536 585
R9226 gnd.n3539 gnd.n3538 585
R9227 gnd.n3541 gnd.n3540 585
R9228 gnd.n3543 gnd.n3542 585
R9229 gnd.n3545 gnd.n3544 585
R9230 gnd.n3548 gnd.n3547 585
R9231 gnd.n3546 gnd.n2131 585
R9232 gnd.n3552 gnd.n2129 585
R9233 gnd.n3554 gnd.n3553 585
R9234 gnd.n3555 gnd.n3554 585
R9235 gnd.n3457 gnd.n2184 585
R9236 gnd.n3457 gnd.n2105 585
R9237 gnd.n3459 gnd.n3458 585
R9238 gnd.n3458 gnd.n2179 585
R9239 gnd.n3455 gnd.n2183 585
R9240 gnd.n3455 gnd.n3454 585
R9241 gnd.n3434 gnd.n2185 585
R9242 gnd.n2197 gnd.n2185 585
R9243 gnd.n3433 gnd.n2195 585
R9244 gnd.n3442 gnd.n2195 585
R9245 gnd.n3168 gnd.n2202 585
R9246 gnd.n3169 gnd.n3168 585
R9247 gnd.n3167 gnd.n3166 585
R9248 gnd.n3167 gnd.n2206 585
R9249 gnd.n3165 gnd.n2208 585
R9250 gnd.n3158 gnd.n2208 585
R9251 gnd.n2221 gnd.n2209 585
R9252 gnd.n2221 gnd.n2213 585
R9253 gnd.n3114 gnd.n2222 585
R9254 gnd.n3148 gnd.n2222 585
R9255 gnd.n3113 gnd.n3112 585
R9256 gnd.n3112 gnd.n2229 585
R9257 gnd.n3111 gnd.n2237 585
R9258 gnd.n3111 gnd.n2228 585
R9259 gnd.n3110 gnd.n2239 585
R9260 gnd.n3110 gnd.n3109 585
R9261 gnd.n3089 gnd.n2238 585
R9262 gnd.n2251 gnd.n2238 585
R9263 gnd.n3088 gnd.n2249 585
R9264 gnd.n3099 gnd.n2249 585
R9265 gnd.n3078 gnd.n2256 585
R9266 gnd.n3080 gnd.n3078 585
R9267 gnd.n3077 gnd.n3076 585
R9268 gnd.n3077 gnd.n2260 585
R9269 gnd.n3075 gnd.n2262 585
R9270 gnd.n3068 gnd.n2262 585
R9271 gnd.n2277 gnd.n2263 585
R9272 gnd.n2277 gnd.n2267 585
R9273 gnd.n3028 gnd.n2278 585
R9274 gnd.n3058 gnd.n2278 585
R9275 gnd.n3027 gnd.n3026 585
R9276 gnd.n3026 gnd.n2285 585
R9277 gnd.n3025 gnd.n2292 585
R9278 gnd.n3025 gnd.n2284 585
R9279 gnd.n3024 gnd.n2294 585
R9280 gnd.n3024 gnd.n3023 585
R9281 gnd.n3003 gnd.n2293 585
R9282 gnd.n2306 gnd.n2293 585
R9283 gnd.n3002 gnd.n2304 585
R9284 gnd.n3013 gnd.n2304 585
R9285 gnd.n2993 gnd.n2311 585
R9286 gnd.n2994 gnd.n2993 585
R9287 gnd.n2992 gnd.n2991 585
R9288 gnd.n2992 gnd.n2315 585
R9289 gnd.n2990 gnd.n2317 585
R9290 gnd.n2983 gnd.n2317 585
R9291 gnd.n2970 gnd.n2318 585
R9292 gnd.n2971 gnd.n2970 585
R9293 gnd.n2923 gnd.n2331 585
R9294 gnd.n2973 gnd.n2331 585
R9295 gnd.n2925 gnd.n2924 585
R9296 gnd.n2926 gnd.n2925 585
R9297 gnd.n2918 gnd.n2421 585
R9298 gnd.n2421 gnd.n2420 585
R9299 gnd.n2916 gnd.n2915 585
R9300 gnd.n2915 gnd.n2402 585
R9301 gnd.n2913 gnd.n2400 585
R9302 gnd.n2934 gnd.n2400 585
R9303 gnd.n2431 gnd.n2430 585
R9304 gnd.n2430 gnd.n2429 585
R9305 gnd.n2907 gnd.n2390 585
R9306 gnd.n2940 gnd.n2390 585
R9307 gnd.n2906 gnd.n2905 585
R9308 gnd.n2905 gnd.n2904 585
R9309 gnd.n2902 gnd.n2433 585
R9310 gnd.n2902 gnd.n2380 585
R9311 gnd.n2901 gnd.n2900 585
R9312 gnd.n2901 gnd.n2379 585
R9313 gnd.n2436 gnd.n2435 585
R9314 gnd.n2892 gnd.n2435 585
R9315 gnd.n2860 gnd.n2859 585
R9316 gnd.n2859 gnd.n2440 585
R9317 gnd.n2861 gnd.n2449 585
R9318 gnd.n2878 gnd.n2449 585
R9319 gnd.n2858 gnd.n2857 585
R9320 gnd.n2857 gnd.n2455 585
R9321 gnd.n2856 gnd.n2463 585
R9322 gnd.n2856 gnd.n2855 585
R9323 gnd.n2841 gnd.n2464 585
R9324 gnd.n2474 gnd.n2464 585
R9325 gnd.n2840 gnd.n2472 585
R9326 gnd.n2847 gnd.n2472 585
R9327 gnd.n2839 gnd.n2838 585
R9328 gnd.n2838 gnd.n2837 585
R9329 gnd.n2483 gnd.n2480 585
R9330 gnd.n2493 gnd.n2483 585
R9331 gnd.n2829 gnd.n2828 585
R9332 gnd.n2828 gnd.n2827 585
R9333 gnd.n2489 gnd.n2488 585
R9334 gnd.n2502 gnd.n2489 585
R9335 gnd.n2809 gnd.n2500 585
R9336 gnd.n2817 gnd.n2500 585
R9337 gnd.n2808 gnd.n2807 585
R9338 gnd.n2807 gnd.n2806 585
R9339 gnd.n2509 gnd.n2507 585
R9340 gnd.n2518 gnd.n2509 585
R9341 gnd.n2798 gnd.n2797 585
R9342 gnd.n2797 gnd.n2796 585
R9343 gnd.n5856 gnd.n5855 585
R9344 gnd.n5855 gnd.n5854 585
R9345 gnd.n5857 gnd.n987 585
R9346 gnd.n4301 gnd.n987 585
R9347 gnd.n5859 gnd.n5858 585
R9348 gnd.n5860 gnd.n5859 585
R9349 gnd.n971 gnd.n970 585
R9350 gnd.n4005 gnd.n971 585
R9351 gnd.n5868 gnd.n5867 585
R9352 gnd.n5867 gnd.n5866 585
R9353 gnd.n5869 gnd.n965 585
R9354 gnd.n3996 gnd.n965 585
R9355 gnd.n5871 gnd.n5870 585
R9356 gnd.n5872 gnd.n5871 585
R9357 gnd.n950 gnd.n949 585
R9358 gnd.n3992 gnd.n950 585
R9359 gnd.n5880 gnd.n5879 585
R9360 gnd.n5879 gnd.n5878 585
R9361 gnd.n5881 gnd.n944 585
R9362 gnd.n3985 gnd.n944 585
R9363 gnd.n5883 gnd.n5882 585
R9364 gnd.n5884 gnd.n5883 585
R9365 gnd.n929 gnd.n928 585
R9366 gnd.n4022 gnd.n929 585
R9367 gnd.n5892 gnd.n5891 585
R9368 gnd.n5891 gnd.n5890 585
R9369 gnd.n5893 gnd.n924 585
R9370 gnd.n3977 gnd.n924 585
R9371 gnd.n5895 gnd.n5894 585
R9372 gnd.n5896 gnd.n5895 585
R9373 gnd.n908 gnd.n906 585
R9374 gnd.n3969 gnd.n908 585
R9375 gnd.n5904 gnd.n5903 585
R9376 gnd.n5903 gnd.n5902 585
R9377 gnd.n907 gnd.n905 585
R9378 gnd.n3956 gnd.n907 585
R9379 gnd.n3945 gnd.n3944 585
R9380 gnd.n3944 gnd.n2014 585
R9381 gnd.n3947 gnd.n3946 585
R9382 gnd.n3948 gnd.n3947 585
R9383 gnd.n3943 gnd.n2027 585
R9384 gnd.n3943 gnd.n3942 585
R9385 gnd.n2026 gnd.n2025 585
R9386 gnd.n3928 gnd.n2025 585
R9387 gnd.n3918 gnd.n3911 585
R9388 gnd.n3918 gnd.n3917 585
R9389 gnd.n3919 gnd.n899 585
R9390 gnd.n3920 gnd.n3919 585
R9391 gnd.n5907 gnd.n897 585
R9392 gnd.n3893 gnd.n897 585
R9393 gnd.n5909 gnd.n5908 585
R9394 gnd.n5910 gnd.n5909 585
R9395 gnd.n883 gnd.n882 585
R9396 gnd.n3883 gnd.n883 585
R9397 gnd.n5918 gnd.n5917 585
R9398 gnd.n5917 gnd.n5916 585
R9399 gnd.n5919 gnd.n877 585
R9400 gnd.n3873 gnd.n877 585
R9401 gnd.n5921 gnd.n5920 585
R9402 gnd.n5922 gnd.n5921 585
R9403 gnd.n861 gnd.n860 585
R9404 gnd.n3839 gnd.n861 585
R9405 gnd.n5930 gnd.n5929 585
R9406 gnd.n5929 gnd.n5928 585
R9407 gnd.n5931 gnd.n855 585
R9408 gnd.n3845 gnd.n855 585
R9409 gnd.n5933 gnd.n5932 585
R9410 gnd.n5934 gnd.n5933 585
R9411 gnd.n839 gnd.n838 585
R9412 gnd.n3825 gnd.n839 585
R9413 gnd.n5942 gnd.n5941 585
R9414 gnd.n5941 gnd.n5940 585
R9415 gnd.n5943 gnd.n833 585
R9416 gnd.n833 gnd.n830 585
R9417 gnd.n5945 gnd.n5944 585
R9418 gnd.n5946 gnd.n5945 585
R9419 gnd.n834 gnd.n832 585
R9420 gnd.n832 gnd.n827 585
R9421 gnd.n3811 gnd.n3810 585
R9422 gnd.n3812 gnd.n3811 585
R9423 gnd.n2091 gnd.n2090 585
R9424 gnd.n2090 gnd.n2087 585
R9425 gnd.n3805 gnd.n3804 585
R9426 gnd.n3804 gnd.n3803 585
R9427 gnd.n2094 gnd.n2093 585
R9428 gnd.n2095 gnd.n2094 585
R9429 gnd.n3783 gnd.n3782 585
R9430 gnd.n3781 gnd.n3644 585
R9431 gnd.n3780 gnd.n3643 585
R9432 gnd.n3785 gnd.n3643 585
R9433 gnd.n3779 gnd.n3778 585
R9434 gnd.n3777 gnd.n3776 585
R9435 gnd.n3775 gnd.n3774 585
R9436 gnd.n3773 gnd.n3772 585
R9437 gnd.n3771 gnd.n3770 585
R9438 gnd.n3769 gnd.n3768 585
R9439 gnd.n3767 gnd.n3766 585
R9440 gnd.n3765 gnd.n3764 585
R9441 gnd.n3763 gnd.n3762 585
R9442 gnd.n3761 gnd.n3760 585
R9443 gnd.n3759 gnd.n3758 585
R9444 gnd.n3757 gnd.n3756 585
R9445 gnd.n3755 gnd.n3754 585
R9446 gnd.n3753 gnd.n3752 585
R9447 gnd.n3751 gnd.n3750 585
R9448 gnd.n3748 gnd.n3747 585
R9449 gnd.n3746 gnd.n3745 585
R9450 gnd.n3744 gnd.n3743 585
R9451 gnd.n3742 gnd.n3741 585
R9452 gnd.n3740 gnd.n3739 585
R9453 gnd.n3738 gnd.n3737 585
R9454 gnd.n3736 gnd.n3735 585
R9455 gnd.n3734 gnd.n3733 585
R9456 gnd.n3732 gnd.n3731 585
R9457 gnd.n3730 gnd.n3729 585
R9458 gnd.n3728 gnd.n3727 585
R9459 gnd.n3726 gnd.n3725 585
R9460 gnd.n3724 gnd.n3723 585
R9461 gnd.n3722 gnd.n3721 585
R9462 gnd.n3720 gnd.n3719 585
R9463 gnd.n3718 gnd.n3717 585
R9464 gnd.n3716 gnd.n3715 585
R9465 gnd.n3714 gnd.n3713 585
R9466 gnd.n3712 gnd.n3683 585
R9467 gnd.n3687 gnd.n3684 585
R9468 gnd.n3708 gnd.n3707 585
R9469 gnd.n4308 gnd.n4307 585
R9470 gnd.n4310 gnd.n1900 585
R9471 gnd.n4312 gnd.n4311 585
R9472 gnd.n4313 gnd.n1893 585
R9473 gnd.n4315 gnd.n4314 585
R9474 gnd.n4317 gnd.n1891 585
R9475 gnd.n4319 gnd.n4318 585
R9476 gnd.n4320 gnd.n1886 585
R9477 gnd.n4322 gnd.n4321 585
R9478 gnd.n4324 gnd.n1884 585
R9479 gnd.n4326 gnd.n4325 585
R9480 gnd.n4327 gnd.n1879 585
R9481 gnd.n4329 gnd.n4328 585
R9482 gnd.n4331 gnd.n1877 585
R9483 gnd.n4333 gnd.n4332 585
R9484 gnd.n4334 gnd.n1872 585
R9485 gnd.n4336 gnd.n4335 585
R9486 gnd.n4338 gnd.n1871 585
R9487 gnd.n4339 gnd.n1814 585
R9488 gnd.n4342 gnd.n4341 585
R9489 gnd.n1815 gnd.n1807 585
R9490 gnd.n1843 gnd.n1808 585
R9491 gnd.n1845 gnd.n1844 585
R9492 gnd.n1847 gnd.n1846 585
R9493 gnd.n1849 gnd.n1848 585
R9494 gnd.n1851 gnd.n1850 585
R9495 gnd.n1853 gnd.n1852 585
R9496 gnd.n1855 gnd.n1854 585
R9497 gnd.n1857 gnd.n1856 585
R9498 gnd.n1859 gnd.n1858 585
R9499 gnd.n1861 gnd.n1860 585
R9500 gnd.n1863 gnd.n1862 585
R9501 gnd.n1865 gnd.n1864 585
R9502 gnd.n1866 gnd.n1825 585
R9503 gnd.n1868 gnd.n1867 585
R9504 gnd.n1826 gnd.n1824 585
R9505 gnd.n1827 gnd.n992 585
R9506 gnd.n1870 gnd.n992 585
R9507 gnd.n4304 gnd.n994 585
R9508 gnd.n5854 gnd.n994 585
R9509 gnd.n4303 gnd.n4302 585
R9510 gnd.n4302 gnd.n4301 585
R9511 gnd.n1904 gnd.n984 585
R9512 gnd.n5860 gnd.n984 585
R9513 gnd.n4004 gnd.n4003 585
R9514 gnd.n4005 gnd.n4004 585
R9515 gnd.n1998 gnd.n973 585
R9516 gnd.n5866 gnd.n973 585
R9517 gnd.n3998 gnd.n3997 585
R9518 gnd.n3997 gnd.n3996 585
R9519 gnd.n3995 gnd.n962 585
R9520 gnd.n5872 gnd.n962 585
R9521 gnd.n3994 gnd.n3993 585
R9522 gnd.n3993 gnd.n3992 585
R9523 gnd.n2000 gnd.n952 585
R9524 gnd.n5878 gnd.n952 585
R9525 gnd.n3987 gnd.n3986 585
R9526 gnd.n3986 gnd.n3985 585
R9527 gnd.n3984 gnd.n941 585
R9528 gnd.n5884 gnd.n941 585
R9529 gnd.n3983 gnd.n1988 585
R9530 gnd.n4022 gnd.n1988 585
R9531 gnd.n2002 gnd.n931 585
R9532 gnd.n5890 gnd.n931 585
R9533 gnd.n3979 gnd.n3978 585
R9534 gnd.n3978 gnd.n3977 585
R9535 gnd.n2004 gnd.n921 585
R9536 gnd.n5896 gnd.n921 585
R9537 gnd.n2041 gnd.n2008 585
R9538 gnd.n3969 gnd.n2008 585
R9539 gnd.n2042 gnd.n910 585
R9540 gnd.n5902 gnd.n910 585
R9541 gnd.n2043 gnd.n2015 585
R9542 gnd.n3956 gnd.n2015 585
R9543 gnd.n2045 gnd.n2044 585
R9544 gnd.n2044 gnd.n2014 585
R9545 gnd.n2046 gnd.n2022 585
R9546 gnd.n3948 gnd.n2022 585
R9547 gnd.n2047 gnd.n2029 585
R9548 gnd.n3942 gnd.n2029 585
R9549 gnd.n3930 gnd.n3929 585
R9550 gnd.n3929 gnd.n3928 585
R9551 gnd.n2048 gnd.n2035 585
R9552 gnd.n3917 gnd.n2048 585
R9553 gnd.n3890 gnd.n2056 585
R9554 gnd.n3920 gnd.n2056 585
R9555 gnd.n3892 gnd.n3891 585
R9556 gnd.n3893 gnd.n3892 585
R9557 gnd.n2061 gnd.n895 585
R9558 gnd.n5910 gnd.n895 585
R9559 gnd.n3885 gnd.n3884 585
R9560 gnd.n3884 gnd.n3883 585
R9561 gnd.n2063 gnd.n884 585
R9562 gnd.n5916 gnd.n884 585
R9563 gnd.n3835 gnd.n2067 585
R9564 gnd.n3873 gnd.n2067 585
R9565 gnd.n3836 gnd.n874 585
R9566 gnd.n5922 gnd.n874 585
R9567 gnd.n3838 gnd.n3837 585
R9568 gnd.n3839 gnd.n3838 585
R9569 gnd.n2078 gnd.n863 585
R9570 gnd.n5928 gnd.n863 585
R9571 gnd.n3829 gnd.n2073 585
R9572 gnd.n3845 gnd.n2073 585
R9573 gnd.n3828 gnd.n853 585
R9574 gnd.n5934 gnd.n853 585
R9575 gnd.n3827 gnd.n3826 585
R9576 gnd.n3826 gnd.n3825 585
R9577 gnd.n2080 gnd.n841 585
R9578 gnd.n5940 gnd.n841 585
R9579 gnd.n3696 gnd.n3695 585
R9580 gnd.n3695 gnd.n830 585
R9581 gnd.n3697 gnd.n828 585
R9582 gnd.n5946 gnd.n828 585
R9583 gnd.n3699 gnd.n3698 585
R9584 gnd.n3698 gnd.n827 585
R9585 gnd.n3700 gnd.n2088 585
R9586 gnd.n3812 gnd.n2088 585
R9587 gnd.n3690 gnd.n3689 585
R9588 gnd.n3689 gnd.n2087 585
R9589 gnd.n3704 gnd.n2096 585
R9590 gnd.n3803 gnd.n2096 585
R9591 gnd.n3706 gnd.n3705 585
R9592 gnd.n3706 gnd.n2095 585
R9593 gnd.n7005 gnd.n7004 585
R9594 gnd.n7006 gnd.n7005 585
R9595 gnd.n87 gnd.n85 585
R9596 gnd.n85 gnd.n81 585
R9597 gnd.n6925 gnd.n6924 585
R9598 gnd.n6926 gnd.n6925 585
R9599 gnd.n164 gnd.n163 585
R9600 gnd.n163 gnd.n161 585
R9601 gnd.n6920 gnd.n6919 585
R9602 gnd.n6919 gnd.n6918 585
R9603 gnd.n167 gnd.n166 585
R9604 gnd.n180 gnd.n167 585
R9605 gnd.n6835 gnd.n6834 585
R9606 gnd.n6836 gnd.n6835 585
R9607 gnd.n182 gnd.n181 585
R9608 gnd.n261 gnd.n181 585
R9609 gnd.n6830 gnd.n6829 585
R9610 gnd.n6829 gnd.n6828 585
R9611 gnd.n185 gnd.n184 585
R9612 gnd.n266 gnd.n185 585
R9613 gnd.n6819 gnd.n6818 585
R9614 gnd.n6820 gnd.n6819 585
R9615 gnd.n198 gnd.n197 585
R9616 gnd.n6763 gnd.n197 585
R9617 gnd.n6814 gnd.n6813 585
R9618 gnd.n6813 gnd.n6812 585
R9619 gnd.n201 gnd.n200 585
R9620 gnd.n6768 gnd.n201 585
R9621 gnd.n6803 gnd.n6802 585
R9622 gnd.n6804 gnd.n6803 585
R9623 gnd.n213 gnd.n212 585
R9624 gnd.n6772 gnd.n212 585
R9625 gnd.n6798 gnd.n6797 585
R9626 gnd.n6797 gnd.n6796 585
R9627 gnd.n222 gnd.n221 585
R9628 gnd.n6777 gnd.n222 585
R9629 gnd.n6787 gnd.n6786 585
R9630 gnd.n6788 gnd.n6787 585
R9631 gnd.n6785 gnd.n6784 585
R9632 gnd.n6784 gnd.n6783 585
R9633 gnd.n5632 gnd.n234 585
R9634 gnd.n5666 gnd.n234 585
R9635 gnd.n5634 gnd.n5633 585
R9636 gnd.n5634 gnd.n1170 585
R9637 gnd.n5637 gnd.n5636 585
R9638 gnd.n5638 gnd.n5637 585
R9639 gnd.n5635 gnd.n5631 585
R9640 gnd.n5631 gnd.n1176 585
R9641 gnd.n5630 gnd.n1183 585
R9642 gnd.n5630 gnd.n5629 585
R9643 gnd.n1182 gnd.n1181 585
R9644 gnd.n5506 gnd.n1181 585
R9645 gnd.n5618 gnd.n5617 585
R9646 gnd.n5619 gnd.n5618 585
R9647 gnd.n5616 gnd.n1197 585
R9648 gnd.n1205 gnd.n1197 585
R9649 gnd.n5615 gnd.n5614 585
R9650 gnd.n5614 gnd.n5613 585
R9651 gnd.n1200 gnd.n1198 585
R9652 gnd.n5595 gnd.n1200 585
R9653 gnd.n5583 gnd.n1225 585
R9654 gnd.n1225 gnd.n1212 585
R9655 gnd.n5585 gnd.n5584 585
R9656 gnd.n5586 gnd.n5585 585
R9657 gnd.n1226 gnd.n1224 585
R9658 gnd.n1233 gnd.n1224 585
R9659 gnd.n5577 gnd.n5576 585
R9660 gnd.n5576 gnd.n5575 585
R9661 gnd.n1229 gnd.n1228 585
R9662 gnd.n5563 gnd.n1229 585
R9663 gnd.n5551 gnd.n1253 585
R9664 gnd.n1253 gnd.n1241 585
R9665 gnd.n5553 gnd.n5552 585
R9666 gnd.n5554 gnd.n5553 585
R9667 gnd.n1254 gnd.n1252 585
R9668 gnd.n5526 gnd.n1252 585
R9669 gnd.n5546 gnd.n5545 585
R9670 gnd.n5545 gnd.n5544 585
R9671 gnd.n1137 gnd.n1136 585
R9672 gnd.n5477 gnd.n1137 585
R9673 gnd.n5703 gnd.n5702 585
R9674 gnd.n5702 gnd.n5701 585
R9675 gnd.n5704 gnd.n1132 585
R9676 gnd.n5468 gnd.n1132 585
R9677 gnd.n5706 gnd.n5705 585
R9678 gnd.n5707 gnd.n5706 585
R9679 gnd.n5367 gnd.n1131 585
R9680 gnd.n5372 gnd.n5370 585
R9681 gnd.n5373 gnd.n5366 585
R9682 gnd.n5373 gnd.n1118 585
R9683 gnd.n5376 gnd.n5375 585
R9684 gnd.n5364 gnd.n5363 585
R9685 gnd.n5381 gnd.n5380 585
R9686 gnd.n5383 gnd.n5362 585
R9687 gnd.n5386 gnd.n5385 585
R9688 gnd.n5360 gnd.n5359 585
R9689 gnd.n5391 gnd.n5390 585
R9690 gnd.n5393 gnd.n5358 585
R9691 gnd.n5396 gnd.n5395 585
R9692 gnd.n5356 gnd.n5355 585
R9693 gnd.n5402 gnd.n5401 585
R9694 gnd.n5404 gnd.n5354 585
R9695 gnd.n5405 gnd.n1291 585
R9696 gnd.n1289 gnd.n1288 585
R9697 gnd.n5415 gnd.n5414 585
R9698 gnd.n5417 gnd.n1287 585
R9699 gnd.n5420 gnd.n5419 585
R9700 gnd.n1285 gnd.n1284 585
R9701 gnd.n5425 gnd.n5424 585
R9702 gnd.n5427 gnd.n1283 585
R9703 gnd.n5430 gnd.n5429 585
R9704 gnd.n1281 gnd.n1280 585
R9705 gnd.n5435 gnd.n5434 585
R9706 gnd.n5437 gnd.n1279 585
R9707 gnd.n5440 gnd.n5439 585
R9708 gnd.n1277 gnd.n1276 585
R9709 gnd.n5445 gnd.n5444 585
R9710 gnd.n5447 gnd.n1275 585
R9711 gnd.n5450 gnd.n5449 585
R9712 gnd.n1273 gnd.n1272 585
R9713 gnd.n5456 gnd.n5455 585
R9714 gnd.n5458 gnd.n1271 585
R9715 gnd.n5459 gnd.n1270 585
R9716 gnd.n5462 gnd.n5461 585
R9717 gnd.n155 gnd.n154 585
R9718 gnd.n6934 gnd.n150 585
R9719 gnd.n6936 gnd.n6935 585
R9720 gnd.n6938 gnd.n148 585
R9721 gnd.n6940 gnd.n6939 585
R9722 gnd.n6941 gnd.n143 585
R9723 gnd.n6943 gnd.n6942 585
R9724 gnd.n6945 gnd.n141 585
R9725 gnd.n6947 gnd.n6946 585
R9726 gnd.n6948 gnd.n136 585
R9727 gnd.n6950 gnd.n6949 585
R9728 gnd.n6952 gnd.n134 585
R9729 gnd.n6954 gnd.n6953 585
R9730 gnd.n6955 gnd.n129 585
R9731 gnd.n6957 gnd.n6956 585
R9732 gnd.n6959 gnd.n127 585
R9733 gnd.n6961 gnd.n6960 585
R9734 gnd.n6962 gnd.n122 585
R9735 gnd.n6964 gnd.n6963 585
R9736 gnd.n6966 gnd.n120 585
R9737 gnd.n6968 gnd.n6967 585
R9738 gnd.n6972 gnd.n115 585
R9739 gnd.n6974 gnd.n6973 585
R9740 gnd.n6976 gnd.n113 585
R9741 gnd.n6978 gnd.n6977 585
R9742 gnd.n6979 gnd.n108 585
R9743 gnd.n6981 gnd.n6980 585
R9744 gnd.n6983 gnd.n106 585
R9745 gnd.n6985 gnd.n6984 585
R9746 gnd.n6986 gnd.n101 585
R9747 gnd.n6988 gnd.n6987 585
R9748 gnd.n6990 gnd.n99 585
R9749 gnd.n6992 gnd.n6991 585
R9750 gnd.n6993 gnd.n94 585
R9751 gnd.n6995 gnd.n6994 585
R9752 gnd.n6997 gnd.n92 585
R9753 gnd.n6999 gnd.n6998 585
R9754 gnd.n7000 gnd.n90 585
R9755 gnd.n7001 gnd.n86 585
R9756 gnd.n86 gnd.n83 585
R9757 gnd.n6930 gnd.n82 585
R9758 gnd.n7006 gnd.n82 585
R9759 gnd.n6929 gnd.n6928 585
R9760 gnd.n6928 gnd.n81 585
R9761 gnd.n6927 gnd.n159 585
R9762 gnd.n6927 gnd.n6926 585
R9763 gnd.n256 gnd.n160 585
R9764 gnd.n161 gnd.n160 585
R9765 gnd.n257 gnd.n169 585
R9766 gnd.n6918 gnd.n169 585
R9767 gnd.n259 gnd.n258 585
R9768 gnd.n258 gnd.n180 585
R9769 gnd.n260 gnd.n178 585
R9770 gnd.n6836 gnd.n178 585
R9771 gnd.n263 gnd.n262 585
R9772 gnd.n262 gnd.n261 585
R9773 gnd.n264 gnd.n187 585
R9774 gnd.n6828 gnd.n187 585
R9775 gnd.n268 gnd.n267 585
R9776 gnd.n267 gnd.n266 585
R9777 gnd.n269 gnd.n195 585
R9778 gnd.n6820 gnd.n195 585
R9779 gnd.n6765 gnd.n6764 585
R9780 gnd.n6764 gnd.n6763 585
R9781 gnd.n6766 gnd.n203 585
R9782 gnd.n6812 gnd.n203 585
R9783 gnd.n6770 gnd.n6769 585
R9784 gnd.n6769 gnd.n6768 585
R9785 gnd.n6771 gnd.n210 585
R9786 gnd.n6804 gnd.n210 585
R9787 gnd.n6774 gnd.n6773 585
R9788 gnd.n6773 gnd.n6772 585
R9789 gnd.n6775 gnd.n224 585
R9790 gnd.n6796 gnd.n224 585
R9791 gnd.n6779 gnd.n6778 585
R9792 gnd.n6778 gnd.n6777 585
R9793 gnd.n6780 gnd.n232 585
R9794 gnd.n6788 gnd.n232 585
R9795 gnd.n6782 gnd.n6781 585
R9796 gnd.n6783 gnd.n6782 585
R9797 gnd.n237 gnd.n236 585
R9798 gnd.n5666 gnd.n236 585
R9799 gnd.n5501 gnd.n5500 585
R9800 gnd.n5500 gnd.n1170 585
R9801 gnd.n5502 gnd.n1177 585
R9802 gnd.n5638 gnd.n1177 585
R9803 gnd.n5504 gnd.n5503 585
R9804 gnd.n5503 gnd.n1176 585
R9805 gnd.n5505 gnd.n1185 585
R9806 gnd.n5629 gnd.n1185 585
R9807 gnd.n5508 gnd.n5507 585
R9808 gnd.n5507 gnd.n5506 585
R9809 gnd.n5509 gnd.n1195 585
R9810 gnd.n5619 gnd.n1195 585
R9811 gnd.n5511 gnd.n5510 585
R9812 gnd.n5510 gnd.n1205 585
R9813 gnd.n5512 gnd.n1202 585
R9814 gnd.n5613 gnd.n1202 585
R9815 gnd.n5513 gnd.n1213 585
R9816 gnd.n5595 gnd.n1213 585
R9817 gnd.n5515 gnd.n5514 585
R9818 gnd.n5514 gnd.n1212 585
R9819 gnd.n5516 gnd.n1221 585
R9820 gnd.n5586 gnd.n1221 585
R9821 gnd.n5518 gnd.n5517 585
R9822 gnd.n5517 gnd.n1233 585
R9823 gnd.n5519 gnd.n1231 585
R9824 gnd.n5575 gnd.n1231 585
R9825 gnd.n5520 gnd.n1242 585
R9826 gnd.n5563 gnd.n1242 585
R9827 gnd.n5522 gnd.n5521 585
R9828 gnd.n5521 gnd.n1241 585
R9829 gnd.n5523 gnd.n1250 585
R9830 gnd.n5554 gnd.n1250 585
R9831 gnd.n5525 gnd.n5524 585
R9832 gnd.n5526 gnd.n5525 585
R9833 gnd.n1259 gnd.n1257 585
R9834 gnd.n5544 gnd.n1257 585
R9835 gnd.n5479 gnd.n5478 585
R9836 gnd.n5478 gnd.n5477 585
R9837 gnd.n1261 gnd.n1139 585
R9838 gnd.n5701 gnd.n1139 585
R9839 gnd.n5467 gnd.n5466 585
R9840 gnd.n5468 gnd.n5467 585
R9841 gnd.n1266 gnd.n1127 585
R9842 gnd.n5707 gnd.n1127 585
R9843 gnd.n5281 gnd.n5280 585
R9844 gnd.n5282 gnd.n5281 585
R9845 gnd.n5195 gnd.n1336 585
R9846 gnd.n1343 gnd.n1336 585
R9847 gnd.n5194 gnd.n5193 585
R9848 gnd.n5193 gnd.n5192 585
R9849 gnd.n1339 gnd.n1338 585
R9850 gnd.n4939 gnd.n1339 585
R9851 gnd.n4928 gnd.n1398 585
R9852 gnd.n1398 gnd.n1393 585
R9853 gnd.n4930 gnd.n4929 585
R9854 gnd.n4931 gnd.n4930 585
R9855 gnd.n4927 gnd.n1397 585
R9856 gnd.n4922 gnd.n1397 585
R9857 gnd.n4926 gnd.n4925 585
R9858 gnd.n4925 gnd.n4924 585
R9859 gnd.n1400 gnd.n1399 585
R9860 gnd.n4907 gnd.n1400 585
R9861 gnd.n4897 gnd.n1419 585
R9862 gnd.n1419 gnd.n1412 585
R9863 gnd.n4899 gnd.n4898 585
R9864 gnd.n4900 gnd.n4899 585
R9865 gnd.n4896 gnd.n1418 585
R9866 gnd.n4856 gnd.n1418 585
R9867 gnd.n4895 gnd.n4894 585
R9868 gnd.n4894 gnd.n4893 585
R9869 gnd.n1421 gnd.n1420 585
R9870 gnd.n4772 gnd.n1421 585
R9871 gnd.n4880 gnd.n4879 585
R9872 gnd.n4881 gnd.n4880 585
R9873 gnd.n4878 gnd.n1433 585
R9874 gnd.n1433 gnd.n1429 585
R9875 gnd.n4877 gnd.n4876 585
R9876 gnd.n4876 gnd.n4875 585
R9877 gnd.n1435 gnd.n1434 585
R9878 gnd.n4780 gnd.n1435 585
R9879 gnd.n4847 gnd.n4846 585
R9880 gnd.n4848 gnd.n4847 585
R9881 gnd.n4845 gnd.n1446 585
R9882 gnd.n1446 gnd.t242 585
R9883 gnd.n4844 gnd.n4843 585
R9884 gnd.n4843 gnd.n4842 585
R9885 gnd.n1448 gnd.n1447 585
R9886 gnd.n4787 gnd.n1448 585
R9887 gnd.n4827 gnd.n4826 585
R9888 gnd.n4828 gnd.n4827 585
R9889 gnd.n4825 gnd.n1459 585
R9890 gnd.n4820 gnd.n1459 585
R9891 gnd.n4824 gnd.n4823 585
R9892 gnd.n4823 gnd.n4822 585
R9893 gnd.n1461 gnd.n1460 585
R9894 gnd.n1473 gnd.n1461 585
R9895 gnd.n4758 gnd.n4757 585
R9896 gnd.n4758 gnd.n1472 585
R9897 gnd.n4762 gnd.n4761 585
R9898 gnd.n4761 gnd.n4760 585
R9899 gnd.n4763 gnd.n1480 585
R9900 gnd.n4800 gnd.n1480 585
R9901 gnd.n4764 gnd.n1490 585
R9902 gnd.n1490 gnd.n1489 585
R9903 gnd.n4766 gnd.n4765 585
R9904 gnd.n4767 gnd.n4766 585
R9905 gnd.n4756 gnd.n1487 585
R9906 gnd.n4750 gnd.n1487 585
R9907 gnd.n4755 gnd.n4754 585
R9908 gnd.n4754 gnd.n4753 585
R9909 gnd.n1492 gnd.n1491 585
R9910 gnd.n4739 gnd.n1492 585
R9911 gnd.n4729 gnd.n1509 585
R9912 gnd.n1509 gnd.n1501 585
R9913 gnd.n4731 gnd.n4730 585
R9914 gnd.n4732 gnd.n4731 585
R9915 gnd.n4728 gnd.n1508 585
R9916 gnd.n1513 gnd.n1508 585
R9917 gnd.n4727 gnd.n4726 585
R9918 gnd.n4726 gnd.n4725 585
R9919 gnd.n1511 gnd.n1510 585
R9920 gnd.n4682 gnd.n1511 585
R9921 gnd.n4713 gnd.n4712 585
R9922 gnd.n4714 gnd.n4713 585
R9923 gnd.n4711 gnd.n1524 585
R9924 gnd.n1524 gnd.n1520 585
R9925 gnd.n4710 gnd.n4709 585
R9926 gnd.n4709 gnd.n4708 585
R9927 gnd.n1526 gnd.n1525 585
R9928 gnd.n4672 gnd.n1526 585
R9929 gnd.n4657 gnd.n4656 585
R9930 gnd.n4656 gnd.n1536 585
R9931 gnd.n4658 gnd.n1546 585
R9932 gnd.n4641 gnd.n1546 585
R9933 gnd.n4660 gnd.n4659 585
R9934 gnd.n4661 gnd.n4660 585
R9935 gnd.n4655 gnd.n1545 585
R9936 gnd.n1545 gnd.n1542 585
R9937 gnd.n4654 gnd.n4653 585
R9938 gnd.n4653 gnd.n4652 585
R9939 gnd.n1548 gnd.n1547 585
R9940 gnd.n4632 gnd.n1548 585
R9941 gnd.n4617 gnd.n4616 585
R9942 gnd.n4616 gnd.n1559 585
R9943 gnd.n4618 gnd.n1569 585
R9944 gnd.n4605 gnd.n1569 585
R9945 gnd.n4620 gnd.n4619 585
R9946 gnd.n4621 gnd.n4620 585
R9947 gnd.n4615 gnd.n1568 585
R9948 gnd.n1568 gnd.n1565 585
R9949 gnd.n4614 gnd.n4613 585
R9950 gnd.n4613 gnd.n4612 585
R9951 gnd.n1571 gnd.n1570 585
R9952 gnd.n4548 gnd.n1571 585
R9953 gnd.n4590 gnd.n4589 585
R9954 gnd.n4591 gnd.n4590 585
R9955 gnd.n4588 gnd.n1586 585
R9956 gnd.n4583 gnd.n1586 585
R9957 gnd.n4587 gnd.n4586 585
R9958 gnd.n4586 gnd.n4585 585
R9959 gnd.n1588 gnd.n1587 585
R9960 gnd.n4576 gnd.n1588 585
R9961 gnd.n4559 gnd.n4558 585
R9962 gnd.n4558 gnd.n4557 585
R9963 gnd.n4560 gnd.n1603 585
R9964 gnd.n4435 gnd.n1603 585
R9965 gnd.n4562 gnd.n4561 585
R9966 gnd.n4563 gnd.n4562 585
R9967 gnd.n1604 gnd.n1602 585
R9968 gnd.t250 gnd.n1602 585
R9969 gnd.n4535 gnd.n4534 585
R9970 gnd.n4536 gnd.n4535 585
R9971 gnd.n4533 gnd.n1615 585
R9972 gnd.n1615 gnd.n1612 585
R9973 gnd.n4532 gnd.n4531 585
R9974 gnd.n4531 gnd.n4530 585
R9975 gnd.n1617 gnd.n1616 585
R9976 gnd.n1626 gnd.n1617 585
R9977 gnd.n4503 gnd.n4502 585
R9978 gnd.n4502 gnd.n1625 585
R9979 gnd.n4504 gnd.n1635 585
R9980 gnd.n4449 gnd.n1635 585
R9981 gnd.n4506 gnd.n4505 585
R9982 gnd.n4507 gnd.n4506 585
R9983 gnd.n4501 gnd.n1634 585
R9984 gnd.n4496 gnd.n1634 585
R9985 gnd.n4500 gnd.n4499 585
R9986 gnd.n4499 gnd.n4498 585
R9987 gnd.n1637 gnd.n1636 585
R9988 gnd.n1647 gnd.n1637 585
R9989 gnd.n4472 gnd.n4471 585
R9990 gnd.n4471 gnd.n1645 585
R9991 gnd.n4473 gnd.n1657 585
R9992 gnd.n4459 gnd.n1657 585
R9993 gnd.n4475 gnd.n4474 585
R9994 gnd.n4476 gnd.n4475 585
R9995 gnd.n4470 gnd.n1656 585
R9996 gnd.n4465 gnd.n1656 585
R9997 gnd.n4469 gnd.n4468 585
R9998 gnd.n4468 gnd.n4467 585
R9999 gnd.n1659 gnd.n1658 585
R10000 gnd.n4429 gnd.n1659 585
R10001 gnd.n4416 gnd.n1677 585
R10002 gnd.n1677 gnd.n1676 585
R10003 gnd.n4418 gnd.n4417 585
R10004 gnd.n4419 gnd.n4418 585
R10005 gnd.n4415 gnd.n1675 585
R10006 gnd.n1675 gnd.n1671 585
R10007 gnd.n4413 gnd.n4412 585
R10008 gnd.n1699 gnd.n1698 585
R10009 gnd.n4409 gnd.n4408 585
R10010 gnd.n4410 gnd.n4409 585
R10011 gnd.n4407 gnd.n1734 585
R10012 gnd.n4406 gnd.n4405 585
R10013 gnd.n4404 gnd.n4403 585
R10014 gnd.n4402 gnd.n4401 585
R10015 gnd.n4400 gnd.n4399 585
R10016 gnd.n4398 gnd.n4397 585
R10017 gnd.n4396 gnd.n4395 585
R10018 gnd.n4394 gnd.n4393 585
R10019 gnd.n4392 gnd.n4391 585
R10020 gnd.n4390 gnd.n4389 585
R10021 gnd.n4388 gnd.n4387 585
R10022 gnd.n4386 gnd.n4385 585
R10023 gnd.n4384 gnd.n4383 585
R10024 gnd.n4382 gnd.n4381 585
R10025 gnd.n4380 gnd.n4379 585
R10026 gnd.n4378 gnd.n4377 585
R10027 gnd.n4376 gnd.n4375 585
R10028 gnd.n4374 gnd.n4373 585
R10029 gnd.n4372 gnd.n4371 585
R10030 gnd.n4370 gnd.n4369 585
R10031 gnd.n4368 gnd.n4367 585
R10032 gnd.n4366 gnd.n4365 585
R10033 gnd.n4364 gnd.n4363 585
R10034 gnd.n4362 gnd.n4361 585
R10035 gnd.n4360 gnd.n4359 585
R10036 gnd.n4358 gnd.n4357 585
R10037 gnd.n4356 gnd.n4355 585
R10038 gnd.n4354 gnd.n4353 585
R10039 gnd.n4352 gnd.n4351 585
R10040 gnd.n4350 gnd.n4349 585
R10041 gnd.n4348 gnd.n1806 585
R10042 gnd.n1805 gnd.n1804 585
R10043 gnd.n1803 gnd.n1802 585
R10044 gnd.n1800 gnd.n1799 585
R10045 gnd.n1798 gnd.n1797 585
R10046 gnd.n1796 gnd.n1795 585
R10047 gnd.n1794 gnd.n1793 585
R10048 gnd.n1792 gnd.n1791 585
R10049 gnd.n1790 gnd.n1789 585
R10050 gnd.n1788 gnd.n1787 585
R10051 gnd.n1786 gnd.n1785 585
R10052 gnd.n1784 gnd.n1783 585
R10053 gnd.n1782 gnd.n1781 585
R10054 gnd.n1780 gnd.n1779 585
R10055 gnd.n1778 gnd.n1777 585
R10056 gnd.n1776 gnd.n1775 585
R10057 gnd.n1774 gnd.n1773 585
R10058 gnd.n1772 gnd.n1771 585
R10059 gnd.n1770 gnd.n1769 585
R10060 gnd.n1768 gnd.n1767 585
R10061 gnd.n1766 gnd.n1765 585
R10062 gnd.n1764 gnd.n1763 585
R10063 gnd.n1762 gnd.n1761 585
R10064 gnd.n1760 gnd.n1759 585
R10065 gnd.n1758 gnd.n1757 585
R10066 gnd.n1756 gnd.n1755 585
R10067 gnd.n1754 gnd.n1753 585
R10068 gnd.n1752 gnd.n1751 585
R10069 gnd.n1750 gnd.n1749 585
R10070 gnd.n1748 gnd.n1747 585
R10071 gnd.n1746 gnd.n1745 585
R10072 gnd.n1744 gnd.n1743 585
R10073 gnd.n5285 gnd.n5284 585
R10074 gnd.n5287 gnd.n5286 585
R10075 gnd.n5289 gnd.n5288 585
R10076 gnd.n5291 gnd.n5290 585
R10077 gnd.n5293 gnd.n5292 585
R10078 gnd.n5295 gnd.n5294 585
R10079 gnd.n5297 gnd.n5296 585
R10080 gnd.n5299 gnd.n5298 585
R10081 gnd.n5301 gnd.n5300 585
R10082 gnd.n5303 gnd.n5302 585
R10083 gnd.n5305 gnd.n5304 585
R10084 gnd.n5307 gnd.n5306 585
R10085 gnd.n5309 gnd.n5308 585
R10086 gnd.n5311 gnd.n5310 585
R10087 gnd.n5313 gnd.n5312 585
R10088 gnd.n5315 gnd.n5314 585
R10089 gnd.n5317 gnd.n5316 585
R10090 gnd.n5319 gnd.n5318 585
R10091 gnd.n5321 gnd.n5320 585
R10092 gnd.n5323 gnd.n5322 585
R10093 gnd.n5325 gnd.n5324 585
R10094 gnd.n5327 gnd.n5326 585
R10095 gnd.n5329 gnd.n5328 585
R10096 gnd.n5331 gnd.n5330 585
R10097 gnd.n5333 gnd.n5332 585
R10098 gnd.n5335 gnd.n5334 585
R10099 gnd.n5337 gnd.n5336 585
R10100 gnd.n5339 gnd.n5338 585
R10101 gnd.n5341 gnd.n5340 585
R10102 gnd.n5343 gnd.n1329 585
R10103 gnd.n5345 gnd.n5344 585
R10104 gnd.n5347 gnd.n1292 585
R10105 gnd.n5349 gnd.n5348 585
R10106 gnd.n5352 gnd.n5351 585
R10107 gnd.n1295 gnd.n1293 585
R10108 gnd.n5218 gnd.n5217 585
R10109 gnd.n5220 gnd.n5219 585
R10110 gnd.n5223 gnd.n5222 585
R10111 gnd.n5225 gnd.n5224 585
R10112 gnd.n5227 gnd.n5226 585
R10113 gnd.n5229 gnd.n5228 585
R10114 gnd.n5231 gnd.n5230 585
R10115 gnd.n5233 gnd.n5232 585
R10116 gnd.n5235 gnd.n5234 585
R10117 gnd.n5237 gnd.n5236 585
R10118 gnd.n5239 gnd.n5238 585
R10119 gnd.n5241 gnd.n5240 585
R10120 gnd.n5243 gnd.n5242 585
R10121 gnd.n5245 gnd.n5244 585
R10122 gnd.n5247 gnd.n5246 585
R10123 gnd.n5249 gnd.n5248 585
R10124 gnd.n5251 gnd.n5250 585
R10125 gnd.n5253 gnd.n5252 585
R10126 gnd.n5255 gnd.n5254 585
R10127 gnd.n5257 gnd.n5256 585
R10128 gnd.n5259 gnd.n5258 585
R10129 gnd.n5261 gnd.n5260 585
R10130 gnd.n5263 gnd.n5262 585
R10131 gnd.n5265 gnd.n5264 585
R10132 gnd.n5267 gnd.n5266 585
R10133 gnd.n5269 gnd.n5268 585
R10134 gnd.n5271 gnd.n5270 585
R10135 gnd.n5273 gnd.n5272 585
R10136 gnd.n5275 gnd.n5274 585
R10137 gnd.n5277 gnd.n5276 585
R10138 gnd.n5278 gnd.n1337 585
R10139 gnd.n5283 gnd.n1332 585
R10140 gnd.n5283 gnd.n5282 585
R10141 gnd.n4935 gnd.n1333 585
R10142 gnd.n1343 gnd.n1333 585
R10143 gnd.n4936 gnd.n1342 585
R10144 gnd.n5192 gnd.n1342 585
R10145 gnd.n4938 gnd.n4937 585
R10146 gnd.n4939 gnd.n4938 585
R10147 gnd.n4934 gnd.n1394 585
R10148 gnd.n1394 gnd.n1393 585
R10149 gnd.n4933 gnd.n4932 585
R10150 gnd.n4932 gnd.n4931 585
R10151 gnd.n1396 gnd.n1395 585
R10152 gnd.n4922 gnd.n1396 585
R10153 gnd.n4904 gnd.n1402 585
R10154 gnd.n4924 gnd.n1402 585
R10155 gnd.n4906 gnd.n4905 585
R10156 gnd.n4907 gnd.n4906 585
R10157 gnd.n4903 gnd.n1414 585
R10158 gnd.n1414 gnd.n1412 585
R10159 gnd.n4902 gnd.n4901 585
R10160 gnd.n4901 gnd.n4900 585
R10161 gnd.n1416 gnd.n1415 585
R10162 gnd.n4856 gnd.n1416 585
R10163 gnd.n4771 gnd.n1423 585
R10164 gnd.n4893 gnd.n1423 585
R10165 gnd.n4774 gnd.n4773 585
R10166 gnd.n4773 gnd.n4772 585
R10167 gnd.n4775 gnd.n1431 585
R10168 gnd.n4881 gnd.n1431 585
R10169 gnd.n4777 gnd.n4776 585
R10170 gnd.n4776 gnd.n1429 585
R10171 gnd.n4778 gnd.n1437 585
R10172 gnd.n4875 gnd.n1437 585
R10173 gnd.n4782 gnd.n4781 585
R10174 gnd.n4781 gnd.n4780 585
R10175 gnd.n4783 gnd.n1444 585
R10176 gnd.n4848 gnd.n1444 585
R10177 gnd.n4785 gnd.n4784 585
R10178 gnd.n4784 gnd.t242 585
R10179 gnd.n4786 gnd.n1450 585
R10180 gnd.n4842 gnd.n1450 585
R10181 gnd.n4789 gnd.n4788 585
R10182 gnd.n4788 gnd.n4787 585
R10183 gnd.n4790 gnd.n1457 585
R10184 gnd.n4828 gnd.n1457 585
R10185 gnd.n4791 gnd.n1464 585
R10186 gnd.n4820 gnd.n1464 585
R10187 gnd.n4792 gnd.n1463 585
R10188 gnd.n4822 gnd.n1463 585
R10189 gnd.n4794 gnd.n4793 585
R10190 gnd.n4794 gnd.n1473 585
R10191 gnd.n4796 gnd.n4795 585
R10192 gnd.n4795 gnd.n1472 585
R10193 gnd.n4797 gnd.n1483 585
R10194 gnd.n4760 gnd.n1483 585
R10195 gnd.n4799 gnd.n4798 585
R10196 gnd.n4800 gnd.n4799 585
R10197 gnd.n4770 gnd.n1482 585
R10198 gnd.n1489 gnd.n1482 585
R10199 gnd.n4769 gnd.n4768 585
R10200 gnd.n4768 gnd.n4767 585
R10201 gnd.n1485 gnd.n1484 585
R10202 gnd.n4750 gnd.n1485 585
R10203 gnd.n4736 gnd.n1494 585
R10204 gnd.n4753 gnd.n1494 585
R10205 gnd.n4738 gnd.n4737 585
R10206 gnd.n4739 gnd.n4738 585
R10207 gnd.n4735 gnd.n1503 585
R10208 gnd.n1503 gnd.n1501 585
R10209 gnd.n4734 gnd.n4733 585
R10210 gnd.n4733 gnd.n4732 585
R10211 gnd.n1505 gnd.n1504 585
R10212 gnd.n1513 gnd.n1505 585
R10213 gnd.n4679 gnd.n1512 585
R10214 gnd.n4725 gnd.n1512 585
R10215 gnd.n4681 gnd.n4680 585
R10216 gnd.n4682 gnd.n4681 585
R10217 gnd.n4678 gnd.n1522 585
R10218 gnd.n4714 gnd.n1522 585
R10219 gnd.n4677 gnd.n4676 585
R10220 gnd.n4676 gnd.n1520 585
R10221 gnd.n4675 gnd.n1528 585
R10222 gnd.n4708 gnd.n1528 585
R10223 gnd.n4674 gnd.n4673 585
R10224 gnd.n4673 gnd.n4672 585
R10225 gnd.n1535 gnd.n1534 585
R10226 gnd.n1536 gnd.n1535 585
R10227 gnd.n4640 gnd.n4639 585
R10228 gnd.n4641 gnd.n4640 585
R10229 gnd.n4638 gnd.n1543 585
R10230 gnd.n4661 gnd.n1543 585
R10231 gnd.n4637 gnd.n4636 585
R10232 gnd.n4636 gnd.n1542 585
R10233 gnd.n4635 gnd.n1550 585
R10234 gnd.n4652 gnd.n1550 585
R10235 gnd.n4634 gnd.n4633 585
R10236 gnd.n4633 gnd.n4632 585
R10237 gnd.n1558 gnd.n1557 585
R10238 gnd.n1559 gnd.n1558 585
R10239 gnd.n4607 gnd.n4606 585
R10240 gnd.n4606 gnd.n4605 585
R10241 gnd.n4608 gnd.n1566 585
R10242 gnd.n4621 gnd.n1566 585
R10243 gnd.n4609 gnd.n1575 585
R10244 gnd.n1575 gnd.n1565 585
R10245 gnd.n4611 gnd.n4610 585
R10246 gnd.n4612 gnd.n4611 585
R10247 gnd.n1576 gnd.n1574 585
R10248 gnd.n4548 gnd.n1574 585
R10249 gnd.n4580 gnd.n1585 585
R10250 gnd.n4591 gnd.n1585 585
R10251 gnd.n4582 gnd.n4581 585
R10252 gnd.n4583 gnd.n4582 585
R10253 gnd.n4579 gnd.n1590 585
R10254 gnd.n4585 gnd.n1590 585
R10255 gnd.n4578 gnd.n4577 585
R10256 gnd.n4577 gnd.n4576 585
R10257 gnd.n1592 gnd.n1591 585
R10258 gnd.n4557 gnd.n1592 585
R10259 gnd.n4437 gnd.n4436 585
R10260 gnd.n4436 gnd.n4435 585
R10261 gnd.n4438 gnd.n1600 585
R10262 gnd.n4563 gnd.n1600 585
R10263 gnd.n4440 gnd.n4439 585
R10264 gnd.n4439 gnd.t250 585
R10265 gnd.n4441 gnd.n1613 585
R10266 gnd.n4536 gnd.n1613 585
R10267 gnd.n4443 gnd.n4442 585
R10268 gnd.n4442 gnd.n1612 585
R10269 gnd.n4444 gnd.n1619 585
R10270 gnd.n4530 gnd.n1619 585
R10271 gnd.n4446 gnd.n4445 585
R10272 gnd.n4446 gnd.n1626 585
R10273 gnd.n4447 gnd.n4434 585
R10274 gnd.n4447 gnd.n1625 585
R10275 gnd.n4451 gnd.n4450 585
R10276 gnd.n4450 gnd.n4449 585
R10277 gnd.n4452 gnd.n1632 585
R10278 gnd.n4507 gnd.n1632 585
R10279 gnd.n4453 gnd.n1639 585
R10280 gnd.n4496 gnd.n1639 585
R10281 gnd.n4454 gnd.n1638 585
R10282 gnd.n4498 gnd.n1638 585
R10283 gnd.n4456 gnd.n4455 585
R10284 gnd.n4456 gnd.n1647 585
R10285 gnd.n4457 gnd.n4433 585
R10286 gnd.n4457 gnd.n1645 585
R10287 gnd.n4461 gnd.n4460 585
R10288 gnd.n4460 gnd.n4459 585
R10289 gnd.n4462 gnd.n1654 585
R10290 gnd.n4476 gnd.n1654 585
R10291 gnd.n4464 gnd.n4463 585
R10292 gnd.n4465 gnd.n4464 585
R10293 gnd.n4432 gnd.n1661 585
R10294 gnd.n4467 gnd.n1661 585
R10295 gnd.n4431 gnd.n4430 585
R10296 gnd.n4430 gnd.n4429 585
R10297 gnd.n1663 gnd.n1662 585
R10298 gnd.n1676 gnd.n1663 585
R10299 gnd.n1740 gnd.n1673 585
R10300 gnd.n4419 gnd.n1673 585
R10301 gnd.n1742 gnd.n1741 585
R10302 gnd.n1742 gnd.n1671 585
R10303 gnd.n5949 gnd.n5948 585
R10304 gnd.n5948 gnd.n5947 585
R10305 gnd.n6750 gnd.n6749 585
R10306 gnd.n6749 gnd.n168 585
R10307 gnd.n6753 gnd.n277 585
R10308 gnd.n277 gnd.n177 585
R10309 gnd.n6755 gnd.n6754 585
R10310 gnd.n6755 gnd.n188 585
R10311 gnd.n6756 gnd.n276 585
R10312 gnd.n6756 gnd.n186 585
R10313 gnd.n6758 gnd.n6757 585
R10314 gnd.n6757 gnd.n196 585
R10315 gnd.n6759 gnd.n271 585
R10316 gnd.n271 gnd.n194 585
R10317 gnd.n6761 gnd.n6760 585
R10318 gnd.n6762 gnd.n6761 585
R10319 gnd.n272 gnd.n270 585
R10320 gnd.n270 gnd.n202 585
R10321 gnd.n5652 gnd.n5651 585
R10322 gnd.n5652 gnd.n211 585
R10323 gnd.n5654 gnd.n5653 585
R10324 gnd.n5653 gnd.n209 585
R10325 gnd.n5655 gnd.n5645 585
R10326 gnd.n5645 gnd.n225 585
R10327 gnd.n5657 gnd.n5656 585
R10328 gnd.n5657 gnd.n223 585
R10329 gnd.n5658 gnd.n5644 585
R10330 gnd.n5658 gnd.n233 585
R10331 gnd.n5660 gnd.n5659 585
R10332 gnd.n5659 gnd.n231 585
R10333 gnd.n5662 gnd.n1172 585
R10334 gnd.n1172 gnd.n235 585
R10335 gnd.n5664 gnd.n5663 585
R10336 gnd.n5665 gnd.n5664 585
R10337 gnd.n5642 gnd.n1171 585
R10338 gnd.n1180 gnd.n1171 585
R10339 gnd.n5641 gnd.n5640 585
R10340 gnd.n5640 gnd.n5639 585
R10341 gnd.n5604 gnd.n1174 585
R10342 gnd.n5628 gnd.n1174 585
R10343 gnd.n5606 gnd.n5605 585
R10344 gnd.n5606 gnd.n1184 585
R10345 gnd.n5608 gnd.n5607 585
R10346 gnd.n5607 gnd.n1196 585
R10347 gnd.n5609 gnd.n1207 585
R10348 gnd.n1207 gnd.n1194 585
R10349 gnd.n5611 gnd.n5610 585
R10350 gnd.n5612 gnd.n5611 585
R10351 gnd.n1208 gnd.n1206 585
R10352 gnd.n1206 gnd.n1201 585
R10353 gnd.n5598 gnd.n5597 585
R10354 gnd.n5597 gnd.n5596 585
R10355 gnd.n1211 gnd.n1210 585
R10356 gnd.n1222 gnd.n1211 585
R10357 gnd.n5571 gnd.n1235 585
R10358 gnd.n1235 gnd.n1220 585
R10359 gnd.n5573 gnd.n5572 585
R10360 gnd.n5574 gnd.n5573 585
R10361 gnd.n1236 gnd.n1234 585
R10362 gnd.n1234 gnd.n1230 585
R10363 gnd.n5566 gnd.n5565 585
R10364 gnd.n5565 gnd.n5564 585
R10365 gnd.n1239 gnd.n1238 585
R10366 gnd.n1251 gnd.n1239 585
R10367 gnd.n5540 gnd.n5528 585
R10368 gnd.n5528 gnd.n1249 585
R10369 gnd.n5542 gnd.n5541 585
R10370 gnd.n5543 gnd.n5542 585
R10371 gnd.n5529 gnd.n5527 585
R10372 gnd.n5527 gnd.n1256 585
R10373 gnd.n5535 gnd.n5534 585
R10374 gnd.n5534 gnd.n1141 585
R10375 gnd.n5533 gnd.n5532 585
R10376 gnd.n5533 gnd.n1138 585
R10377 gnd.n1125 gnd.n1124 585
R10378 gnd.n1129 gnd.n1125 585
R10379 gnd.n5710 gnd.n5709 585
R10380 gnd.n5709 gnd.n5708 585
R10381 gnd.n5711 gnd.n1119 585
R10382 gnd.n1126 gnd.n1119 585
R10383 gnd.n5713 gnd.n5712 585
R10384 gnd.n5714 gnd.n5713 585
R10385 gnd.n1116 gnd.n1115 585
R10386 gnd.n5715 gnd.n1116 585
R10387 gnd.n5718 gnd.n5717 585
R10388 gnd.n5717 gnd.n5716 585
R10389 gnd.n5719 gnd.n1110 585
R10390 gnd.n1110 gnd.n1108 585
R10391 gnd.n5721 gnd.n5720 585
R10392 gnd.n5722 gnd.n5721 585
R10393 gnd.n1111 gnd.n1109 585
R10394 gnd.n1109 gnd.n1106 585
R10395 gnd.n5156 gnd.n5155 585
R10396 gnd.n5157 gnd.n5156 585
R10397 gnd.n1375 gnd.n1374 585
R10398 gnd.n5159 gnd.n1375 585
R10399 gnd.n5164 gnd.n5163 585
R10400 gnd.n5163 gnd.n5162 585
R10401 gnd.n5165 gnd.n1369 585
R10402 gnd.n1376 gnd.n1369 585
R10403 gnd.n5167 gnd.n5166 585
R10404 gnd.n5168 gnd.n5167 585
R10405 gnd.n1363 gnd.n1362 585
R10406 gnd.n5170 gnd.n1363 585
R10407 gnd.n5175 gnd.n5174 585
R10408 gnd.n5174 gnd.n5173 585
R10409 gnd.n5176 gnd.n1355 585
R10410 gnd.n1364 gnd.n1355 585
R10411 gnd.n5178 gnd.n5177 585
R10412 gnd.n5179 gnd.n5178 585
R10413 gnd.n1356 gnd.n1351 585
R10414 gnd.n5181 gnd.n1351 585
R10415 gnd.n5185 gnd.n1350 585
R10416 gnd.n5185 gnd.n5184 585
R10417 gnd.n5187 gnd.n5186 585
R10418 gnd.n5186 gnd.n1296 585
R10419 gnd.n5188 gnd.n1345 585
R10420 gnd.n1345 gnd.n1334 585
R10421 gnd.n5190 gnd.n5189 585
R10422 gnd.n5191 gnd.n5190 585
R10423 gnd.n1346 gnd.n1344 585
R10424 gnd.n4939 gnd.n1344 585
R10425 gnd.n4918 gnd.n1407 585
R10426 gnd.n1407 gnd.n1406 585
R10427 gnd.n4920 gnd.n4919 585
R10428 gnd.n4921 gnd.n4920 585
R10429 gnd.n1408 gnd.n1405 585
R10430 gnd.n1405 gnd.n1401 585
R10431 gnd.n4912 gnd.n4911 585
R10432 gnd.n4911 gnd.n4910 585
R10433 gnd.n1411 gnd.n1410 585
R10434 gnd.n1417 gnd.n1411 585
R10435 gnd.n4891 gnd.n4890 585
R10436 gnd.n4892 gnd.n4891 585
R10437 gnd.n1425 gnd.n1424 585
R10438 gnd.n1432 gnd.n1424 585
R10439 gnd.n4886 gnd.n4885 585
R10440 gnd.n4885 gnd.n4884 585
R10441 gnd.n1428 gnd.n1427 585
R10442 gnd.n1436 gnd.n1428 585
R10443 gnd.n4836 gnd.n1452 585
R10444 gnd.n1452 gnd.n1445 585
R10445 gnd.n4838 gnd.n4837 585
R10446 gnd.n4839 gnd.n4838 585
R10447 gnd.n1453 gnd.n1451 585
R10448 gnd.n1451 gnd.n1449 585
R10449 gnd.n4831 gnd.n4830 585
R10450 gnd.n4830 gnd.n4829 585
R10451 gnd.n1456 gnd.n1455 585
R10452 gnd.n4821 gnd.n1456 585
R10453 gnd.n4807 gnd.n4806 585
R10454 gnd.n4808 gnd.n4807 585
R10455 gnd.n1475 gnd.n1474 585
R10456 gnd.n4759 gnd.n1474 585
R10457 gnd.n4802 gnd.n4801 585
R10458 gnd.n4801 gnd.n4800 585
R10459 gnd.n1478 gnd.n1477 585
R10460 gnd.n1488 gnd.n1478 585
R10461 gnd.n4748 gnd.n4747 585
R10462 gnd.n4749 gnd.n4748 585
R10463 gnd.n1497 gnd.n1496 585
R10464 gnd.n1496 gnd.n1493 585
R10465 gnd.n4743 gnd.n4742 585
R10466 gnd.n4742 gnd.n4741 585
R10467 gnd.n1500 gnd.n1499 585
R10468 gnd.n1506 gnd.n1500 585
R10469 gnd.n4723 gnd.n4722 585
R10470 gnd.n4724 gnd.n4723 585
R10471 gnd.n1516 gnd.n1515 585
R10472 gnd.n1523 gnd.n1515 585
R10473 gnd.n4718 gnd.n4717 585
R10474 gnd.n4717 gnd.n4716 585
R10475 gnd.n1519 gnd.n1518 585
R10476 gnd.n1527 gnd.n1519 585
R10477 gnd.n4669 gnd.n4668 585
R10478 gnd.n4670 gnd.n4669 585
R10479 gnd.n1538 gnd.n1537 585
R10480 gnd.n1556 gnd.n1537 585
R10481 gnd.n4664 gnd.n4663 585
R10482 gnd.n4663 gnd.n4662 585
R10483 gnd.n1541 gnd.n1540 585
R10484 gnd.n1549 gnd.n1541 585
R10485 gnd.n4629 gnd.n4628 585
R10486 gnd.n4630 gnd.n4629 585
R10487 gnd.n1561 gnd.n1560 585
R10488 gnd.n1577 gnd.n1560 585
R10489 gnd.n4624 gnd.n4623 585
R10490 gnd.n4623 gnd.n4622 585
R10491 gnd.n1564 gnd.n1563 585
R10492 gnd.n4612 gnd.n1564 585
R10493 gnd.n4550 gnd.n4547 585
R10494 gnd.n4550 gnd.n4549 585
R10495 gnd.n4552 gnd.n4551 585
R10496 gnd.n4551 gnd.n1584 585
R10497 gnd.n4553 gnd.n1607 585
R10498 gnd.n1607 gnd.n1589 585
R10499 gnd.n4555 gnd.n4554 585
R10500 gnd.n4556 gnd.n4555 585
R10501 gnd.n1608 gnd.n1606 585
R10502 gnd.n1606 gnd.n1601 585
R10503 gnd.n4540 gnd.n4539 585
R10504 gnd.n4539 gnd.n1599 585
R10505 gnd.n4538 gnd.n1610 585
R10506 gnd.n4538 gnd.n4537 585
R10507 gnd.n4515 gnd.n1611 585
R10508 gnd.n4529 gnd.n1611 585
R10509 gnd.n4517 gnd.n4516 585
R10510 gnd.n4518 gnd.n4517 585
R10511 gnd.n1628 gnd.n1627 585
R10512 gnd.n4448 gnd.n1627 585
R10513 gnd.n4510 gnd.n4509 585
R10514 gnd.n4509 gnd.n4508 585
R10515 gnd.n1631 gnd.n1630 585
R10516 gnd.n4497 gnd.n1631 585
R10517 gnd.n4484 gnd.n4483 585
R10518 gnd.n4485 gnd.n4484 585
R10519 gnd.n1649 gnd.n1648 585
R10520 gnd.n4458 gnd.n1648 585
R10521 gnd.n4479 gnd.n4478 585
R10522 gnd.n4478 gnd.n4477 585
R10523 gnd.n1652 gnd.n1651 585
R10524 gnd.n4466 gnd.n1652 585
R10525 gnd.n4428 gnd.n4427 585
R10526 gnd.n4429 gnd.n4428 585
R10527 gnd.n1667 gnd.n1666 585
R10528 gnd.n1674 gnd.n1666 585
R10529 gnd.n4423 gnd.n4422 585
R10530 gnd.n4422 gnd.n4421 585
R10531 gnd.n1670 gnd.n1669 585
R10532 gnd.n1733 gnd.n1670 585
R10533 gnd.n4239 gnd.n4238 585
R10534 gnd.n4240 gnd.n4239 585
R10535 gnd.n1944 gnd.n1943 585
R10536 gnd.n4230 gnd.n1943 585
R10537 gnd.n4234 gnd.n4233 585
R10538 gnd.n4233 gnd.n4232 585
R10539 gnd.n1947 gnd.n1946 585
R10540 gnd.n4228 gnd.n1947 585
R10541 gnd.n4225 gnd.n4224 585
R10542 gnd.n4226 gnd.n4225 585
R10543 gnd.n1952 gnd.n1951 585
R10544 gnd.n4216 gnd.n1951 585
R10545 gnd.n4220 gnd.n4219 585
R10546 gnd.n4219 gnd.n4218 585
R10547 gnd.n1955 gnd.n1954 585
R10548 gnd.n4214 gnd.n1955 585
R10549 gnd.n4211 gnd.n4210 585
R10550 gnd.n4212 gnd.n4211 585
R10551 gnd.n1960 gnd.n1959 585
R10552 gnd.n4202 gnd.n1959 585
R10553 gnd.n4206 gnd.n4205 585
R10554 gnd.n4205 gnd.n4204 585
R10555 gnd.n1963 gnd.n1962 585
R10556 gnd.n4200 gnd.n1963 585
R10557 gnd.n4197 gnd.n4196 585
R10558 gnd.n4198 gnd.n4197 585
R10559 gnd.n1966 gnd.n1965 585
R10560 gnd.n1965 gnd.n1964 585
R10561 gnd.n4192 gnd.n4191 585
R10562 gnd.n4191 gnd.n4190 585
R10563 gnd.n1969 gnd.n1968 585
R10564 gnd.n4056 gnd.n1969 585
R10565 gnd.n4054 gnd.n4053 585
R10566 gnd.n4055 gnd.n4054 585
R10567 gnd.n1972 gnd.n1971 585
R10568 gnd.n1971 gnd.n1970 585
R10569 gnd.n4049 gnd.n4048 585
R10570 gnd.n4048 gnd.n996 585
R10571 gnd.n4047 gnd.n1974 585
R10572 gnd.n4047 gnd.n993 585
R10573 gnd.n4046 gnd.n4045 585
R10574 gnd.n4046 gnd.n986 585
R10575 gnd.n1976 gnd.n1975 585
R10576 gnd.n1975 gnd.n983 585
R10577 gnd.n4041 gnd.n4040 585
R10578 gnd.n4040 gnd.n975 585
R10579 gnd.n4039 gnd.n1978 585
R10580 gnd.n4039 gnd.n972 585
R10581 gnd.n4038 gnd.n4037 585
R10582 gnd.n4038 gnd.n964 585
R10583 gnd.n1980 gnd.n1979 585
R10584 gnd.n3991 gnd.n1979 585
R10585 gnd.n4033 gnd.n4032 585
R10586 gnd.n4032 gnd.n954 585
R10587 gnd.n4031 gnd.n1982 585
R10588 gnd.n4031 gnd.n951 585
R10589 gnd.n4030 gnd.n4029 585
R10590 gnd.n4030 gnd.n943 585
R10591 gnd.n1984 gnd.n1983 585
R10592 gnd.n1983 gnd.n940 585
R10593 gnd.n4025 gnd.n4024 585
R10594 gnd.n4024 gnd.n4023 585
R10595 gnd.n1987 gnd.n1986 585
R10596 gnd.n1987 gnd.n930 585
R10597 gnd.n3965 gnd.n2010 585
R10598 gnd.n2010 gnd.n923 585
R10599 gnd.n3967 gnd.n3966 585
R10600 gnd.n3968 gnd.n3967 585
R10601 gnd.n3961 gnd.n2009 585
R10602 gnd.n2009 gnd.n912 585
R10603 gnd.n3960 gnd.n3959 585
R10604 gnd.n3959 gnd.n909 585
R10605 gnd.n3958 gnd.n2013 585
R10606 gnd.n3958 gnd.n3957 585
R10607 gnd.n3899 gnd.n2012 585
R10608 gnd.n2023 gnd.n2012 585
R10609 gnd.n3902 gnd.n3901 585
R10610 gnd.n3902 gnd.n2021 585
R10611 gnd.n3904 gnd.n3903 585
R10612 gnd.n3903 gnd.n2028 585
R10613 gnd.n3906 gnd.n2058 585
R10614 gnd.n2058 gnd.n2049 585
R10615 gnd.n3908 gnd.n3907 585
R10616 gnd.n3909 gnd.n3908 585
R10617 gnd.n3897 gnd.n2057 585
R10618 gnd.n2057 gnd.n2055 585
R10619 gnd.n3896 gnd.n3895 585
R10620 gnd.n3895 gnd.n3894 585
R10621 gnd.n3868 gnd.n2060 585
R10622 gnd.n2060 gnd.n894 585
R10623 gnd.n3869 gnd.n2069 585
R10624 gnd.n2069 gnd.n886 585
R10625 gnd.n3871 gnd.n3870 585
R10626 gnd.n3872 gnd.n3871 585
R10627 gnd.n2070 gnd.n2068 585
R10628 gnd.n2068 gnd.n876 585
R10629 gnd.n3863 gnd.n3862 585
R10630 gnd.n3862 gnd.n873 585
R10631 gnd.n3861 gnd.n2072 585
R10632 gnd.n3861 gnd.n865 585
R10633 gnd.n3860 gnd.n3859 585
R10634 gnd.n3860 gnd.n862 585
R10635 gnd.n3848 gnd.n3847 585
R10636 gnd.n3847 gnd.n3846 585
R10637 gnd.n3855 gnd.n3854 585
R10638 gnd.n3854 gnd.n852 585
R10639 gnd.n3853 gnd.n3852 585
R10640 gnd.n3853 gnd.n843 585
R10641 gnd.n3851 gnd.n826 585
R10642 gnd.n840 gnd.n826 585
R10643 gnd.n5725 gnd.n5724 585
R10644 gnd.n5724 gnd.n5723 585
R10645 gnd.n5726 gnd.n1103 585
R10646 gnd.n5151 gnd.n1103 585
R10647 gnd.n5727 gnd.n1102 585
R10648 gnd.n5158 gnd.n1102 585
R10649 gnd.n5160 gnd.n1100 585
R10650 gnd.n5161 gnd.n5160 585
R10651 gnd.n5731 gnd.n1099 585
R10652 gnd.n1377 gnd.n1099 585
R10653 gnd.n5732 gnd.n1098 585
R10654 gnd.n1368 gnd.n1098 585
R10655 gnd.n5733 gnd.n1097 585
R10656 gnd.n5169 gnd.n1097 585
R10657 gnd.n5171 gnd.n1095 585
R10658 gnd.n5172 gnd.n5171 585
R10659 gnd.n5737 gnd.n1094 585
R10660 gnd.n1365 gnd.n1094 585
R10661 gnd.n5738 gnd.n1093 585
R10662 gnd.n1354 gnd.n1093 585
R10663 gnd.n5739 gnd.n1092 585
R10664 gnd.n5180 gnd.n1092 585
R10665 gnd.n5182 gnd.n1090 585
R10666 gnd.n5183 gnd.n5182 585
R10667 gnd.n5743 gnd.n1089 585
R10668 gnd.n1313 gnd.n1089 585
R10669 gnd.n5744 gnd.n1088 585
R10670 gnd.n1335 gnd.n1088 585
R10671 gnd.n5745 gnd.n1087 585
R10672 gnd.n4948 gnd.n1087 585
R10673 gnd.n1340 gnd.n1085 585
R10674 gnd.n1341 gnd.n1340 585
R10675 gnd.n5749 gnd.n1084 585
R10676 gnd.n4940 gnd.n1084 585
R10677 gnd.n5750 gnd.n1083 585
R10678 gnd.n1404 gnd.n1083 585
R10679 gnd.n5751 gnd.n1082 585
R10680 gnd.n4923 gnd.n1082 585
R10681 gnd.n4908 gnd.n1080 585
R10682 gnd.n4909 gnd.n4908 585
R10683 gnd.n5755 gnd.n1079 585
R10684 gnd.n4859 gnd.n1079 585
R10685 gnd.n5756 gnd.n1078 585
R10686 gnd.n4857 gnd.n1078 585
R10687 gnd.n5757 gnd.n1077 585
R10688 gnd.n1422 gnd.n1077 585
R10689 gnd.n4882 gnd.n1075 585
R10690 gnd.n4883 gnd.n4882 585
R10691 gnd.n5761 gnd.n1074 585
R10692 gnd.n4874 gnd.n1074 585
R10693 gnd.n5762 gnd.n1073 585
R10694 gnd.n4779 gnd.n1073 585
R10695 gnd.n5763 gnd.n1072 585
R10696 gnd.n4849 gnd.n1072 585
R10697 gnd.n4840 gnd.n1070 585
R10698 gnd.n4841 gnd.n4840 585
R10699 gnd.n5767 gnd.n1069 585
R10700 gnd.n1458 gnd.n1069 585
R10701 gnd.n5768 gnd.n1068 585
R10702 gnd.n4819 gnd.n1068 585
R10703 gnd.n5769 gnd.n1067 585
R10704 gnd.n1462 gnd.n1067 585
R10705 gnd.n4809 gnd.n1065 585
R10706 gnd.n4810 gnd.n4809 585
R10707 gnd.n5773 gnd.n1064 585
R10708 gnd.n1481 gnd.n1064 585
R10709 gnd.n5774 gnd.n1063 585
R10710 gnd.n1479 gnd.n1063 585
R10711 gnd.n5775 gnd.n1062 585
R10712 gnd.n1486 gnd.n1062 585
R10713 gnd.n4751 gnd.n1060 585
R10714 gnd.n4752 gnd.n4751 585
R10715 gnd.n5779 gnd.n1059 585
R10716 gnd.n4740 gnd.n1059 585
R10717 gnd.n5780 gnd.n1058 585
R10718 gnd.n1507 gnd.n1058 585
R10719 gnd.n5781 gnd.n1057 585
R10720 gnd.n1514 gnd.n1057 585
R10721 gnd.n4683 gnd.n1055 585
R10722 gnd.n4684 gnd.n4683 585
R10723 gnd.n5785 gnd.n1054 585
R10724 gnd.n4715 gnd.n1054 585
R10725 gnd.n5786 gnd.n1053 585
R10726 gnd.n4707 gnd.n1053 585
R10727 gnd.n5787 gnd.n1052 585
R10728 gnd.n4671 gnd.n1052 585
R10729 gnd.n4642 gnd.n1050 585
R10730 gnd.n4643 gnd.n4642 585
R10731 gnd.n5791 gnd.n1049 585
R10732 gnd.n1544 gnd.n1049 585
R10733 gnd.n5792 gnd.n1048 585
R10734 gnd.n4651 gnd.n1048 585
R10735 gnd.n5793 gnd.n1047 585
R10736 gnd.n4631 gnd.n1047 585
R10737 gnd.n4603 gnd.n1045 585
R10738 gnd.n4604 gnd.n4603 585
R10739 gnd.n5797 gnd.n1044 585
R10740 gnd.n1567 gnd.n1044 585
R10741 gnd.n5798 gnd.n1043 585
R10742 gnd.n1573 gnd.n1043 585
R10743 gnd.n5799 gnd.n1042 585
R10744 gnd.n1572 gnd.n1042 585
R10745 gnd.n4592 gnd.n1040 585
R10746 gnd.n4593 gnd.n4592 585
R10747 gnd.n5803 gnd.n1039 585
R10748 gnd.n4584 gnd.n1039 585
R10749 gnd.n5804 gnd.n1038 585
R10750 gnd.n4575 gnd.n1038 585
R10751 gnd.n5805 gnd.n1037 585
R10752 gnd.n1605 gnd.n1037 585
R10753 gnd.n4564 gnd.n1035 585
R10754 gnd.n4565 gnd.n4564 585
R10755 gnd.n5809 gnd.n1034 585
R10756 gnd.n1614 gnd.n1034 585
R10757 gnd.n5810 gnd.n1033 585
R10758 gnd.n4528 gnd.n1033 585
R10759 gnd.n5811 gnd.n1032 585
R10760 gnd.n1618 gnd.n1032 585
R10761 gnd.n4519 gnd.n1030 585
R10762 gnd.n4520 gnd.n4519 585
R10763 gnd.n5815 gnd.n1029 585
R10764 gnd.n1633 gnd.n1029 585
R10765 gnd.n5816 gnd.n1028 585
R10766 gnd.n4495 gnd.n1028 585
R10767 gnd.n5817 gnd.n1027 585
R10768 gnd.n1646 gnd.n1027 585
R10769 gnd.n4486 gnd.n1025 585
R10770 gnd.n4487 gnd.n4486 585
R10771 gnd.n5821 gnd.n1024 585
R10772 gnd.n1655 gnd.n1024 585
R10773 gnd.n5822 gnd.n1023 585
R10774 gnd.n1653 gnd.n1023 585
R10775 gnd.n5823 gnd.n1022 585
R10776 gnd.n1660 gnd.n1022 585
R10777 gnd.n1664 gnd.n1020 585
R10778 gnd.n1665 gnd.n1664 585
R10779 gnd.n5827 gnd.n1019 585
R10780 gnd.n4420 gnd.n1019 585
R10781 gnd.n5828 gnd.n1018 585
R10782 gnd.n4245 gnd.n1018 585
R10783 gnd.n5829 gnd.n1017 585
R10784 gnd.n1700 gnd.n1017 585
R10785 gnd.n4241 gnd.n1015 585
R10786 gnd.n4242 gnd.n4241 585
R10787 gnd.n5833 gnd.n1014 585
R10788 gnd.n4231 gnd.n1014 585
R10789 gnd.n5834 gnd.n1013 585
R10790 gnd.n4229 gnd.n1013 585
R10791 gnd.n5835 gnd.n1012 585
R10792 gnd.n4227 gnd.n1012 585
R10793 gnd.n1949 gnd.n1010 585
R10794 gnd.n1950 gnd.n1949 585
R10795 gnd.n5839 gnd.n1009 585
R10796 gnd.n4217 gnd.n1009 585
R10797 gnd.n5840 gnd.n1008 585
R10798 gnd.n4215 gnd.n1008 585
R10799 gnd.n5841 gnd.n1007 585
R10800 gnd.n4213 gnd.n1007 585
R10801 gnd.n1957 gnd.n1005 585
R10802 gnd.n1958 gnd.n1957 585
R10803 gnd.n5845 gnd.n1004 585
R10804 gnd.n4203 gnd.n1004 585
R10805 gnd.n5846 gnd.n1003 585
R10806 gnd.n4201 gnd.n1003 585
R10807 gnd.n5847 gnd.n1002 585
R10808 gnd.n4199 gnd.n1002 585
R10809 gnd.n4187 gnd.n4186 585
R10810 gnd.n4185 gnd.n4073 585
R10811 gnd.n4075 gnd.n4072 585
R10812 gnd.n4189 gnd.n4072 585
R10813 gnd.n4178 gnd.n4088 585
R10814 gnd.n4177 gnd.n4089 585
R10815 gnd.n4091 gnd.n4090 585
R10816 gnd.n4170 gnd.n4099 585
R10817 gnd.n4169 gnd.n4100 585
R10818 gnd.n4110 gnd.n4101 585
R10819 gnd.n4162 gnd.n4111 585
R10820 gnd.n4161 gnd.n4112 585
R10821 gnd.n4114 gnd.n4113 585
R10822 gnd.n4154 gnd.n4122 585
R10823 gnd.n4153 gnd.n4123 585
R10824 gnd.n4135 gnd.n4124 585
R10825 gnd.n4146 gnd.n4136 585
R10826 gnd.n4145 gnd.n4138 585
R10827 gnd.n4137 gnd.n1910 585
R10828 gnd.n4294 gnd.n1911 585
R10829 gnd.n4293 gnd.n1912 585
R10830 gnd.n4292 gnd.n1913 585
R10831 gnd.n4066 gnd.n1914 585
R10832 gnd.n4288 gnd.n1916 585
R10833 gnd.n4287 gnd.n1917 585
R10834 gnd.n4286 gnd.n1918 585
R10835 gnd.n4283 gnd.n1923 585
R10836 gnd.n4282 gnd.n1924 585
R10837 gnd.n4281 gnd.n1925 585
R10838 gnd.n4070 gnd.n1926 585
R10839 gnd.n1381 gnd.n1107 585
R10840 gnd.n5723 gnd.n1107 585
R10841 gnd.n5150 gnd.n5149 585
R10842 gnd.n5151 gnd.n5150 585
R10843 gnd.n1380 gnd.n1379 585
R10844 gnd.n5158 gnd.n1379 585
R10845 gnd.n4969 gnd.n1378 585
R10846 gnd.n5161 gnd.n1378 585
R10847 gnd.n4968 gnd.n4967 585
R10848 gnd.n4967 gnd.n1377 585
R10849 gnd.n4966 gnd.n4965 585
R10850 gnd.n4966 gnd.n1368 585
R10851 gnd.n1383 gnd.n1367 585
R10852 gnd.n5169 gnd.n1367 585
R10853 gnd.n4961 gnd.n1366 585
R10854 gnd.n5172 gnd.n1366 585
R10855 gnd.n4960 gnd.n4959 585
R10856 gnd.n4959 gnd.n1365 585
R10857 gnd.n4958 gnd.n4957 585
R10858 gnd.n4958 gnd.n1354 585
R10859 gnd.n1385 gnd.n1353 585
R10860 gnd.n5180 gnd.n1353 585
R10861 gnd.n4953 gnd.n1352 585
R10862 gnd.n5183 gnd.n1352 585
R10863 gnd.n4952 gnd.n4951 585
R10864 gnd.n4951 gnd.n1313 585
R10865 gnd.n4950 gnd.n1387 585
R10866 gnd.n4950 gnd.n1335 585
R10867 gnd.n4949 gnd.n4947 585
R10868 gnd.n4949 gnd.n4948 585
R10869 gnd.n1389 gnd.n1388 585
R10870 gnd.n1388 gnd.n1341 585
R10871 gnd.n4942 gnd.n4941 585
R10872 gnd.n4941 gnd.n4940 585
R10873 gnd.n1392 gnd.n1391 585
R10874 gnd.n1404 gnd.n1392 585
R10875 gnd.n4862 gnd.n1403 585
R10876 gnd.n4923 gnd.n1403 585
R10877 gnd.n4861 gnd.n1413 585
R10878 gnd.n4909 gnd.n1413 585
R10879 gnd.n4866 gnd.n4860 585
R10880 gnd.n4860 gnd.n4859 585
R10881 gnd.n4867 gnd.n4858 585
R10882 gnd.n4858 gnd.n4857 585
R10883 gnd.n4868 gnd.n4855 585
R10884 gnd.n4855 gnd.n1422 585
R10885 gnd.n1440 gnd.n1430 585
R10886 gnd.n4883 gnd.n1430 585
R10887 gnd.n4873 gnd.n4872 585
R10888 gnd.n4874 gnd.n4873 585
R10889 gnd.n1439 gnd.n1438 585
R10890 gnd.n4779 gnd.n1438 585
R10891 gnd.n4851 gnd.n4850 585
R10892 gnd.n4850 gnd.n4849 585
R10893 gnd.n1443 gnd.n1442 585
R10894 gnd.n4841 gnd.n1443 585
R10895 gnd.n1468 gnd.n1466 585
R10896 gnd.n1466 gnd.n1458 585
R10897 gnd.n4818 gnd.n4817 585
R10898 gnd.n4819 gnd.n4818 585
R10899 gnd.n1467 gnd.n1465 585
R10900 gnd.n1465 gnd.n1462 585
R10901 gnd.n4812 gnd.n4811 585
R10902 gnd.n4811 gnd.n4810 585
R10903 gnd.n1471 gnd.n1470 585
R10904 gnd.n1481 gnd.n1471 585
R10905 gnd.n4693 gnd.n4691 585
R10906 gnd.n4691 gnd.n1479 585
R10907 gnd.n4694 gnd.n4690 585
R10908 gnd.n4690 gnd.n1486 585
R10909 gnd.n4695 gnd.n1495 585
R10910 gnd.n4752 gnd.n1495 585
R10911 gnd.n4688 gnd.n1502 585
R10912 gnd.n4740 gnd.n1502 585
R10913 gnd.n4699 gnd.n4687 585
R10914 gnd.n4687 gnd.n1507 585
R10915 gnd.n4700 gnd.n4686 585
R10916 gnd.n4686 gnd.n1514 585
R10917 gnd.n4701 gnd.n4685 585
R10918 gnd.n4685 gnd.n4684 585
R10919 gnd.n1531 gnd.n1521 585
R10920 gnd.n4715 gnd.n1521 585
R10921 gnd.n4706 gnd.n4705 585
R10922 gnd.n4707 gnd.n4706 585
R10923 gnd.n1530 gnd.n1529 585
R10924 gnd.n4671 gnd.n1529 585
R10925 gnd.n4645 gnd.n4644 585
R10926 gnd.n4644 gnd.n4643 585
R10927 gnd.n1554 gnd.n1552 585
R10928 gnd.n1552 gnd.n1544 585
R10929 gnd.n4650 gnd.n4649 585
R10930 gnd.n4651 gnd.n4650 585
R10931 gnd.n1553 gnd.n1551 585
R10932 gnd.n4631 gnd.n1551 585
R10933 gnd.n4602 gnd.n4601 585
R10934 gnd.n4604 gnd.n4602 585
R10935 gnd.n1579 gnd.n1578 585
R10936 gnd.n1578 gnd.n1567 585
R10937 gnd.n4597 gnd.n4596 585
R10938 gnd.n4596 gnd.n1573 585
R10939 gnd.n4595 gnd.n1581 585
R10940 gnd.n4595 gnd.n1572 585
R10941 gnd.n4594 gnd.n1583 585
R10942 gnd.n4594 gnd.n4593 585
R10943 gnd.n1595 gnd.n1582 585
R10944 gnd.n4584 gnd.n1582 585
R10945 gnd.n4574 gnd.n4573 585
R10946 gnd.n4575 gnd.n4574 585
R10947 gnd.n1594 gnd.n1593 585
R10948 gnd.n1605 gnd.n1593 585
R10949 gnd.n4567 gnd.n4566 585
R10950 gnd.n4566 gnd.n4565 585
R10951 gnd.n1598 gnd.n1597 585
R10952 gnd.n1614 gnd.n1598 585
R10953 gnd.n4527 gnd.n4526 585
R10954 gnd.n4528 gnd.n4527 585
R10955 gnd.n1621 gnd.n1620 585
R10956 gnd.n1620 gnd.n1618 585
R10957 gnd.n4522 gnd.n4521 585
R10958 gnd.n4521 gnd.n4520 585
R10959 gnd.n1624 gnd.n1623 585
R10960 gnd.n1633 gnd.n1624 585
R10961 gnd.n4494 gnd.n4493 585
R10962 gnd.n4495 gnd.n4494 585
R10963 gnd.n1641 gnd.n1640 585
R10964 gnd.n1646 gnd.n1640 585
R10965 gnd.n4489 gnd.n4488 585
R10966 gnd.n4488 gnd.n4487 585
R10967 gnd.n1644 gnd.n1643 585
R10968 gnd.n1655 gnd.n1644 585
R10969 gnd.n4252 gnd.n4251 585
R10970 gnd.n4251 gnd.n1653 585
R10971 gnd.n4253 gnd.n4250 585
R10972 gnd.n4250 gnd.n1660 585
R10973 gnd.n4249 gnd.n4247 585
R10974 gnd.n4249 gnd.n1665 585
R10975 gnd.n4257 gnd.n1672 585
R10976 gnd.n4420 gnd.n1672 585
R10977 gnd.n4258 gnd.n4246 585
R10978 gnd.n4246 gnd.n4245 585
R10979 gnd.n4259 gnd.n4244 585
R10980 gnd.n4244 gnd.n1700 585
R10981 gnd.n4243 gnd.n1941 585
R10982 gnd.n4243 gnd.n4242 585
R10983 gnd.n4263 gnd.n1940 585
R10984 gnd.n4231 gnd.n1940 585
R10985 gnd.n4264 gnd.n1939 585
R10986 gnd.n4229 gnd.n1939 585
R10987 gnd.n4265 gnd.n1938 585
R10988 gnd.n4227 gnd.n1938 585
R10989 gnd.n1948 gnd.n1936 585
R10990 gnd.n1950 gnd.n1948 585
R10991 gnd.n4269 gnd.n1935 585
R10992 gnd.n4217 gnd.n1935 585
R10993 gnd.n4270 gnd.n1934 585
R10994 gnd.n4215 gnd.n1934 585
R10995 gnd.n4271 gnd.n1933 585
R10996 gnd.n4213 gnd.n1933 585
R10997 gnd.n1956 gnd.n1931 585
R10998 gnd.n1958 gnd.n1956 585
R10999 gnd.n4275 gnd.n1930 585
R11000 gnd.n4203 gnd.n1930 585
R11001 gnd.n4276 gnd.n1929 585
R11002 gnd.n4201 gnd.n1929 585
R11003 gnd.n4277 gnd.n1928 585
R11004 gnd.n4199 gnd.n1928 585
R11005 gnd.n5145 gnd.n5144 585
R11006 gnd.n5144 gnd.n1117 585
R11007 gnd.n5143 gnd.n4973 585
R11008 gnd.n5141 gnd.n5140 585
R11009 gnd.n4975 gnd.n4974 585
R11010 gnd.n5136 gnd.n5132 585
R11011 gnd.n5130 gnd.n4977 585
R11012 gnd.n5128 gnd.n5127 585
R11013 gnd.n4979 gnd.n4978 585
R11014 gnd.n5123 gnd.n5122 585
R11015 gnd.n5120 gnd.n4981 585
R11016 gnd.n5118 gnd.n5117 585
R11017 gnd.n4983 gnd.n4982 585
R11018 gnd.n5103 gnd.n5102 585
R11019 gnd.n5104 gnd.n5100 585
R11020 gnd.n5098 gnd.n4992 585
R11021 gnd.n5097 gnd.n5096 585
R11022 gnd.n5081 gnd.n4994 585
R11023 gnd.n5083 gnd.n5082 585
R11024 gnd.n5079 gnd.n5001 585
R11025 gnd.n5078 gnd.n5077 585
R11026 gnd.n5062 gnd.n5003 585
R11027 gnd.n5064 gnd.n5063 585
R11028 gnd.n5060 gnd.n5010 585
R11029 gnd.n5059 gnd.n5058 585
R11030 gnd.n5043 gnd.n5012 585
R11031 gnd.n5045 gnd.n5044 585
R11032 gnd.n5041 gnd.n5019 585
R11033 gnd.n5040 gnd.n5039 585
R11034 gnd.n5021 gnd.n1105 585
R11035 gnd.n6115 gnd.n655 530.795
R11036 gnd.n5281 gnd.n1337 511.721
R11037 gnd.n5284 gnd.n5283 511.721
R11038 gnd.n1743 gnd.n1742 511.721
R11039 gnd.n4412 gnd.n1675 511.721
R11040 gnd.n1738 gnd.t210 389.64
R11041 gnd.n1330 gnd.t160 389.64
R11042 gnd.n1735 gnd.t138 389.64
R11043 gnd.n5215 gnd.t213 389.64
R11044 gnd.n1919 gnd.t200 371.625
R11045 gnd.n6877 gnd.t185 371.625
R11046 gnd.n4985 gnd.t178 371.625
R11047 gnd.n4131 gnd.t197 371.625
R11048 gnd.n5408 gnd.t175 371.625
R11049 gnd.n1268 gnd.t149 371.625
R11050 gnd.n156 gnd.t142 371.625
R11051 gnd.n6969 gnd.t164 371.625
R11052 gnd.n3663 gnd.t232 371.625
R11053 gnd.n3685 gnd.t223 371.625
R11054 gnd.n3584 gnd.t219 371.625
R11055 gnd.n1898 gnd.t156 371.625
R11056 gnd.n1809 gnd.t188 371.625
R11057 gnd.n5133 gnd.t181 371.625
R11058 gnd.n2574 gnd.t131 323.425
R11059 gnd.n2144 gnd.t167 323.425
R11060 gnd.n3423 gnd.n3397 289.615
R11061 gnd.n3391 gnd.n3365 289.615
R11062 gnd.n3359 gnd.n3333 289.615
R11063 gnd.n3328 gnd.n3302 289.615
R11064 gnd.n3296 gnd.n3270 289.615
R11065 gnd.n3264 gnd.n3238 289.615
R11066 gnd.n3232 gnd.n3206 289.615
R11067 gnd.n3201 gnd.n3175 289.615
R11068 gnd.n2648 gnd.t235 279.217
R11069 gnd.n2170 gnd.t171 279.217
R11070 gnd.n1684 gnd.t137 260.649
R11071 gnd.n5207 gnd.t196 260.649
R11072 gnd.n4411 gnd.n4410 256.663
R11073 gnd.n4410 gnd.n1701 256.663
R11074 gnd.n4410 gnd.n1702 256.663
R11075 gnd.n4410 gnd.n1703 256.663
R11076 gnd.n4410 gnd.n1704 256.663
R11077 gnd.n4410 gnd.n1705 256.663
R11078 gnd.n4410 gnd.n1706 256.663
R11079 gnd.n4410 gnd.n1707 256.663
R11080 gnd.n4410 gnd.n1708 256.663
R11081 gnd.n4410 gnd.n1709 256.663
R11082 gnd.n4410 gnd.n1710 256.663
R11083 gnd.n4410 gnd.n1711 256.663
R11084 gnd.n4410 gnd.n1712 256.663
R11085 gnd.n4410 gnd.n1713 256.663
R11086 gnd.n4410 gnd.n1714 256.663
R11087 gnd.n4410 gnd.n1715 256.663
R11088 gnd.n4350 gnd.n4347 256.663
R11089 gnd.n4410 gnd.n1716 256.663
R11090 gnd.n4410 gnd.n1717 256.663
R11091 gnd.n4410 gnd.n1718 256.663
R11092 gnd.n4410 gnd.n1719 256.663
R11093 gnd.n4410 gnd.n1720 256.663
R11094 gnd.n4410 gnd.n1721 256.663
R11095 gnd.n4410 gnd.n1722 256.663
R11096 gnd.n4410 gnd.n1723 256.663
R11097 gnd.n4410 gnd.n1724 256.663
R11098 gnd.n4410 gnd.n1725 256.663
R11099 gnd.n4410 gnd.n1726 256.663
R11100 gnd.n4410 gnd.n1727 256.663
R11101 gnd.n4410 gnd.n1728 256.663
R11102 gnd.n4410 gnd.n1729 256.663
R11103 gnd.n4410 gnd.n1730 256.663
R11104 gnd.n4410 gnd.n1731 256.663
R11105 gnd.n4410 gnd.n1732 256.663
R11106 gnd.n5349 gnd.n1314 256.663
R11107 gnd.n5349 gnd.n1315 256.663
R11108 gnd.n5349 gnd.n1316 256.663
R11109 gnd.n5349 gnd.n1317 256.663
R11110 gnd.n5349 gnd.n1318 256.663
R11111 gnd.n5349 gnd.n1319 256.663
R11112 gnd.n5349 gnd.n1320 256.663
R11113 gnd.n5349 gnd.n1321 256.663
R11114 gnd.n5349 gnd.n1322 256.663
R11115 gnd.n5349 gnd.n1323 256.663
R11116 gnd.n5349 gnd.n1324 256.663
R11117 gnd.n5349 gnd.n1325 256.663
R11118 gnd.n5349 gnd.n1326 256.663
R11119 gnd.n5349 gnd.n1327 256.663
R11120 gnd.n5349 gnd.n1328 256.663
R11121 gnd.n5349 gnd.n5346 256.663
R11122 gnd.n5352 gnd.n1294 256.663
R11123 gnd.n5350 gnd.n5349 256.663
R11124 gnd.n5349 gnd.n1312 256.663
R11125 gnd.n5349 gnd.n1311 256.663
R11126 gnd.n5349 gnd.n1310 256.663
R11127 gnd.n5349 gnd.n1309 256.663
R11128 gnd.n5349 gnd.n1308 256.663
R11129 gnd.n5349 gnd.n1307 256.663
R11130 gnd.n5349 gnd.n1306 256.663
R11131 gnd.n5349 gnd.n1305 256.663
R11132 gnd.n5349 gnd.n1304 256.663
R11133 gnd.n5349 gnd.n1303 256.663
R11134 gnd.n5349 gnd.n1302 256.663
R11135 gnd.n5349 gnd.n1301 256.663
R11136 gnd.n5349 gnd.n1300 256.663
R11137 gnd.n5349 gnd.n1299 256.663
R11138 gnd.n5349 gnd.n1298 256.663
R11139 gnd.n5349 gnd.n1297 256.663
R11140 gnd.n3786 gnd.n3785 242.672
R11141 gnd.n3785 gnd.n3574 242.672
R11142 gnd.n3785 gnd.n3575 242.672
R11143 gnd.n3785 gnd.n3576 242.672
R11144 gnd.n3785 gnd.n3577 242.672
R11145 gnd.n3785 gnd.n3578 242.672
R11146 gnd.n3785 gnd.n3579 242.672
R11147 gnd.n3785 gnd.n3580 242.672
R11148 gnd.n3785 gnd.n3581 242.672
R11149 gnd.n4140 gnd.n1870 242.672
R11150 gnd.n4129 gnd.n1870 242.672
R11151 gnd.n4126 gnd.n1870 242.672
R11152 gnd.n4117 gnd.n1870 242.672
R11153 gnd.n4106 gnd.n1870 242.672
R11154 gnd.n4103 gnd.n1870 242.672
R11155 gnd.n4094 gnd.n1870 242.672
R11156 gnd.n4084 gnd.n1870 242.672
R11157 gnd.n4081 gnd.n1870 242.672
R11158 gnd.n5031 gnd.n1118 242.672
R11159 gnd.n5033 gnd.n1118 242.672
R11160 gnd.n5050 gnd.n1118 242.672
R11161 gnd.n5052 gnd.n1118 242.672
R11162 gnd.n5069 gnd.n1118 242.672
R11163 gnd.n5071 gnd.n1118 242.672
R11164 gnd.n5088 gnd.n1118 242.672
R11165 gnd.n5090 gnd.n1118 242.672
R11166 gnd.n5109 gnd.n1118 242.672
R11167 gnd.n6879 gnd.n83 242.672
R11168 gnd.n6875 gnd.n83 242.672
R11169 gnd.n6870 gnd.n83 242.672
R11170 gnd.n6867 gnd.n83 242.672
R11171 gnd.n6862 gnd.n83 242.672
R11172 gnd.n6859 gnd.n83 242.672
R11173 gnd.n6854 gnd.n83 242.672
R11174 gnd.n6851 gnd.n83 242.672
R11175 gnd.n6846 gnd.n83 242.672
R11176 gnd.n2702 gnd.n2701 242.672
R11177 gnd.n2702 gnd.n2612 242.672
R11178 gnd.n2702 gnd.n2613 242.672
R11179 gnd.n2702 gnd.n2614 242.672
R11180 gnd.n2702 gnd.n2615 242.672
R11181 gnd.n2702 gnd.n2616 242.672
R11182 gnd.n2702 gnd.n2617 242.672
R11183 gnd.n2702 gnd.n2618 242.672
R11184 gnd.n2702 gnd.n2619 242.672
R11185 gnd.n2702 gnd.n2620 242.672
R11186 gnd.n2702 gnd.n2621 242.672
R11187 gnd.n2702 gnd.n2622 242.672
R11188 gnd.n2703 gnd.n2702 242.672
R11189 gnd.n3555 gnd.n2119 242.672
R11190 gnd.n3555 gnd.n2118 242.672
R11191 gnd.n3555 gnd.n2117 242.672
R11192 gnd.n3555 gnd.n2116 242.672
R11193 gnd.n3555 gnd.n2115 242.672
R11194 gnd.n3555 gnd.n2114 242.672
R11195 gnd.n3555 gnd.n2113 242.672
R11196 gnd.n3555 gnd.n2112 242.672
R11197 gnd.n3555 gnd.n2111 242.672
R11198 gnd.n3555 gnd.n2110 242.672
R11199 gnd.n3555 gnd.n2109 242.672
R11200 gnd.n3555 gnd.n2108 242.672
R11201 gnd.n3555 gnd.n2107 242.672
R11202 gnd.n2786 gnd.n2785 242.672
R11203 gnd.n2785 gnd.n2524 242.672
R11204 gnd.n2785 gnd.n2525 242.672
R11205 gnd.n2785 gnd.n2526 242.672
R11206 gnd.n2785 gnd.n2527 242.672
R11207 gnd.n2785 gnd.n2528 242.672
R11208 gnd.n2785 gnd.n2529 242.672
R11209 gnd.n2785 gnd.n2530 242.672
R11210 gnd.n3555 gnd.n2120 242.672
R11211 gnd.n3555 gnd.n2121 242.672
R11212 gnd.n3555 gnd.n2122 242.672
R11213 gnd.n3555 gnd.n2123 242.672
R11214 gnd.n3555 gnd.n2124 242.672
R11215 gnd.n3555 gnd.n2125 242.672
R11216 gnd.n3555 gnd.n2126 242.672
R11217 gnd.n3555 gnd.n2127 242.672
R11218 gnd.n3785 gnd.n3784 242.672
R11219 gnd.n3785 gnd.n3556 242.672
R11220 gnd.n3785 gnd.n3557 242.672
R11221 gnd.n3785 gnd.n3558 242.672
R11222 gnd.n3785 gnd.n3559 242.672
R11223 gnd.n3785 gnd.n3560 242.672
R11224 gnd.n3785 gnd.n3561 242.672
R11225 gnd.n3785 gnd.n3562 242.672
R11226 gnd.n3785 gnd.n3563 242.672
R11227 gnd.n3785 gnd.n3564 242.672
R11228 gnd.n3785 gnd.n3565 242.672
R11229 gnd.n3785 gnd.n3566 242.672
R11230 gnd.n3785 gnd.n3567 242.672
R11231 gnd.n3785 gnd.n3568 242.672
R11232 gnd.n3785 gnd.n3569 242.672
R11233 gnd.n3785 gnd.n3570 242.672
R11234 gnd.n3785 gnd.n3571 242.672
R11235 gnd.n3785 gnd.n3572 242.672
R11236 gnd.n3785 gnd.n3573 242.672
R11237 gnd.n4309 gnd.n1870 242.672
R11238 gnd.n1901 gnd.n1870 242.672
R11239 gnd.n4316 gnd.n1870 242.672
R11240 gnd.n1892 gnd.n1870 242.672
R11241 gnd.n4323 gnd.n1870 242.672
R11242 gnd.n1885 gnd.n1870 242.672
R11243 gnd.n4330 gnd.n1870 242.672
R11244 gnd.n1878 gnd.n1870 242.672
R11245 gnd.n4337 gnd.n1870 242.672
R11246 gnd.n4340 gnd.n1870 242.672
R11247 gnd.n1870 gnd.n1816 242.672
R11248 gnd.n4346 gnd.n1811 242.672
R11249 gnd.n1870 gnd.n1817 242.672
R11250 gnd.n1870 gnd.n1818 242.672
R11251 gnd.n1870 gnd.n1819 242.672
R11252 gnd.n1870 gnd.n1820 242.672
R11253 gnd.n1870 gnd.n1821 242.672
R11254 gnd.n1870 gnd.n1822 242.672
R11255 gnd.n1870 gnd.n1823 242.672
R11256 gnd.n1870 gnd.n1869 242.672
R11257 gnd.n5371 gnd.n1118 242.672
R11258 gnd.n5374 gnd.n1118 242.672
R11259 gnd.n5382 gnd.n1118 242.672
R11260 gnd.n5384 gnd.n1118 242.672
R11261 gnd.n5392 gnd.n1118 242.672
R11262 gnd.n5394 gnd.n1118 242.672
R11263 gnd.n5403 gnd.n1118 242.672
R11264 gnd.n5406 gnd.n1118 242.672
R11265 gnd.n5410 gnd.n5407 242.672
R11266 gnd.n5353 gnd.n1118 242.672
R11267 gnd.n5416 gnd.n1118 242.672
R11268 gnd.n5418 gnd.n1118 242.672
R11269 gnd.n5426 gnd.n1118 242.672
R11270 gnd.n5428 gnd.n1118 242.672
R11271 gnd.n5436 gnd.n1118 242.672
R11272 gnd.n5438 gnd.n1118 242.672
R11273 gnd.n5446 gnd.n1118 242.672
R11274 gnd.n5448 gnd.n1118 242.672
R11275 gnd.n5457 gnd.n1118 242.672
R11276 gnd.n5460 gnd.n1118 242.672
R11277 gnd.n153 gnd.n83 242.672
R11278 gnd.n6937 gnd.n83 242.672
R11279 gnd.n149 gnd.n83 242.672
R11280 gnd.n6944 gnd.n83 242.672
R11281 gnd.n142 gnd.n83 242.672
R11282 gnd.n6951 gnd.n83 242.672
R11283 gnd.n135 gnd.n83 242.672
R11284 gnd.n6958 gnd.n83 242.672
R11285 gnd.n128 gnd.n83 242.672
R11286 gnd.n6965 gnd.n83 242.672
R11287 gnd.n121 gnd.n83 242.672
R11288 gnd.n6975 gnd.n83 242.672
R11289 gnd.n114 gnd.n83 242.672
R11290 gnd.n6982 gnd.n83 242.672
R11291 gnd.n107 gnd.n83 242.672
R11292 gnd.n6989 gnd.n83 242.672
R11293 gnd.n100 gnd.n83 242.672
R11294 gnd.n6996 gnd.n83 242.672
R11295 gnd.n93 gnd.n83 242.672
R11296 gnd.n4189 gnd.n4188 242.672
R11297 gnd.n4189 gnd.n4057 242.672
R11298 gnd.n4189 gnd.n4058 242.672
R11299 gnd.n4189 gnd.n4059 242.672
R11300 gnd.n4189 gnd.n4060 242.672
R11301 gnd.n4189 gnd.n4061 242.672
R11302 gnd.n4189 gnd.n4062 242.672
R11303 gnd.n4189 gnd.n4063 242.672
R11304 gnd.n4189 gnd.n4064 242.672
R11305 gnd.n4189 gnd.n4065 242.672
R11306 gnd.n4189 gnd.n4067 242.672
R11307 gnd.n4189 gnd.n4068 242.672
R11308 gnd.n4189 gnd.n4069 242.672
R11309 gnd.n4189 gnd.n4071 242.672
R11310 gnd.n5142 gnd.n1117 242.672
R11311 gnd.n5131 gnd.n1117 242.672
R11312 gnd.n5129 gnd.n1117 242.672
R11313 gnd.n5121 gnd.n1117 242.672
R11314 gnd.n5119 gnd.n1117 242.672
R11315 gnd.n5101 gnd.n1117 242.672
R11316 gnd.n5099 gnd.n1117 242.672
R11317 gnd.n4993 gnd.n1117 242.672
R11318 gnd.n5080 gnd.n1117 242.672
R11319 gnd.n5002 gnd.n1117 242.672
R11320 gnd.n5061 gnd.n1117 242.672
R11321 gnd.n5011 gnd.n1117 242.672
R11322 gnd.n5042 gnd.n1117 242.672
R11323 gnd.n5020 gnd.n1117 242.672
R11324 gnd.n90 gnd.n86 240.244
R11325 gnd.n6998 gnd.n6997 240.244
R11326 gnd.n6995 gnd.n94 240.244
R11327 gnd.n6991 gnd.n6990 240.244
R11328 gnd.n6988 gnd.n101 240.244
R11329 gnd.n6984 gnd.n6983 240.244
R11330 gnd.n6981 gnd.n108 240.244
R11331 gnd.n6977 gnd.n6976 240.244
R11332 gnd.n6974 gnd.n115 240.244
R11333 gnd.n6967 gnd.n6966 240.244
R11334 gnd.n6964 gnd.n122 240.244
R11335 gnd.n6960 gnd.n6959 240.244
R11336 gnd.n6957 gnd.n129 240.244
R11337 gnd.n6953 gnd.n6952 240.244
R11338 gnd.n6950 gnd.n136 240.244
R11339 gnd.n6946 gnd.n6945 240.244
R11340 gnd.n6943 gnd.n143 240.244
R11341 gnd.n6939 gnd.n6938 240.244
R11342 gnd.n6936 gnd.n150 240.244
R11343 gnd.n5467 gnd.n1127 240.244
R11344 gnd.n5467 gnd.n1139 240.244
R11345 gnd.n5478 gnd.n1139 240.244
R11346 gnd.n5478 gnd.n1257 240.244
R11347 gnd.n5525 gnd.n1257 240.244
R11348 gnd.n5525 gnd.n1250 240.244
R11349 gnd.n5521 gnd.n1250 240.244
R11350 gnd.n5521 gnd.n1242 240.244
R11351 gnd.n1242 gnd.n1231 240.244
R11352 gnd.n5517 gnd.n1231 240.244
R11353 gnd.n5517 gnd.n1221 240.244
R11354 gnd.n5514 gnd.n1221 240.244
R11355 gnd.n5514 gnd.n1213 240.244
R11356 gnd.n1213 gnd.n1202 240.244
R11357 gnd.n5510 gnd.n1202 240.244
R11358 gnd.n5510 gnd.n1195 240.244
R11359 gnd.n5507 gnd.n1195 240.244
R11360 gnd.n5507 gnd.n1185 240.244
R11361 gnd.n5503 gnd.n1185 240.244
R11362 gnd.n5503 gnd.n1177 240.244
R11363 gnd.n5500 gnd.n1177 240.244
R11364 gnd.n5500 gnd.n236 240.244
R11365 gnd.n6782 gnd.n236 240.244
R11366 gnd.n6782 gnd.n232 240.244
R11367 gnd.n6778 gnd.n232 240.244
R11368 gnd.n6778 gnd.n224 240.244
R11369 gnd.n6773 gnd.n224 240.244
R11370 gnd.n6773 gnd.n210 240.244
R11371 gnd.n6769 gnd.n210 240.244
R11372 gnd.n6769 gnd.n203 240.244
R11373 gnd.n6764 gnd.n203 240.244
R11374 gnd.n6764 gnd.n195 240.244
R11375 gnd.n267 gnd.n195 240.244
R11376 gnd.n267 gnd.n187 240.244
R11377 gnd.n262 gnd.n187 240.244
R11378 gnd.n262 gnd.n178 240.244
R11379 gnd.n258 gnd.n178 240.244
R11380 gnd.n258 gnd.n169 240.244
R11381 gnd.n169 gnd.n160 240.244
R11382 gnd.n6927 gnd.n160 240.244
R11383 gnd.n6928 gnd.n6927 240.244
R11384 gnd.n6928 gnd.n82 240.244
R11385 gnd.n5373 gnd.n5372 240.244
R11386 gnd.n5375 gnd.n5373 240.244
R11387 gnd.n5381 gnd.n5363 240.244
R11388 gnd.n5385 gnd.n5383 240.244
R11389 gnd.n5391 gnd.n5359 240.244
R11390 gnd.n5395 gnd.n5393 240.244
R11391 gnd.n5402 gnd.n5355 240.244
R11392 gnd.n5405 gnd.n5404 240.244
R11393 gnd.n5415 gnd.n1288 240.244
R11394 gnd.n5419 gnd.n5417 240.244
R11395 gnd.n5425 gnd.n1284 240.244
R11396 gnd.n5429 gnd.n5427 240.244
R11397 gnd.n5435 gnd.n1280 240.244
R11398 gnd.n5439 gnd.n5437 240.244
R11399 gnd.n5445 gnd.n1276 240.244
R11400 gnd.n5449 gnd.n5447 240.244
R11401 gnd.n5456 gnd.n1272 240.244
R11402 gnd.n5459 gnd.n5458 240.244
R11403 gnd.n5706 gnd.n1132 240.244
R11404 gnd.n5702 gnd.n1132 240.244
R11405 gnd.n5702 gnd.n1137 240.244
R11406 gnd.n5545 gnd.n1137 240.244
R11407 gnd.n5545 gnd.n1252 240.244
R11408 gnd.n5553 gnd.n1252 240.244
R11409 gnd.n5553 gnd.n1253 240.244
R11410 gnd.n1253 gnd.n1229 240.244
R11411 gnd.n5576 gnd.n1229 240.244
R11412 gnd.n5576 gnd.n1224 240.244
R11413 gnd.n5585 gnd.n1224 240.244
R11414 gnd.n5585 gnd.n1225 240.244
R11415 gnd.n1225 gnd.n1200 240.244
R11416 gnd.n5614 gnd.n1200 240.244
R11417 gnd.n5614 gnd.n1197 240.244
R11418 gnd.n5618 gnd.n1197 240.244
R11419 gnd.n5618 gnd.n1181 240.244
R11420 gnd.n5630 gnd.n1181 240.244
R11421 gnd.n5631 gnd.n5630 240.244
R11422 gnd.n5637 gnd.n5631 240.244
R11423 gnd.n5637 gnd.n5634 240.244
R11424 gnd.n5634 gnd.n234 240.244
R11425 gnd.n6784 gnd.n234 240.244
R11426 gnd.n6787 gnd.n6784 240.244
R11427 gnd.n6787 gnd.n222 240.244
R11428 gnd.n6797 gnd.n222 240.244
R11429 gnd.n6797 gnd.n212 240.244
R11430 gnd.n6803 gnd.n212 240.244
R11431 gnd.n6803 gnd.n201 240.244
R11432 gnd.n6813 gnd.n201 240.244
R11433 gnd.n6813 gnd.n197 240.244
R11434 gnd.n6819 gnd.n197 240.244
R11435 gnd.n6819 gnd.n185 240.244
R11436 gnd.n6829 gnd.n185 240.244
R11437 gnd.n6829 gnd.n181 240.244
R11438 gnd.n6835 gnd.n181 240.244
R11439 gnd.n6835 gnd.n167 240.244
R11440 gnd.n6919 gnd.n167 240.244
R11441 gnd.n6919 gnd.n163 240.244
R11442 gnd.n6925 gnd.n163 240.244
R11443 gnd.n6925 gnd.n85 240.244
R11444 gnd.n7005 gnd.n85 240.244
R11445 gnd.n1824 gnd.n992 240.244
R11446 gnd.n1868 gnd.n1825 240.244
R11447 gnd.n1864 gnd.n1863 240.244
R11448 gnd.n1860 gnd.n1859 240.244
R11449 gnd.n1856 gnd.n1855 240.244
R11450 gnd.n1852 gnd.n1851 240.244
R11451 gnd.n1848 gnd.n1847 240.244
R11452 gnd.n1844 gnd.n1843 240.244
R11453 gnd.n4341 gnd.n1815 240.244
R11454 gnd.n4339 gnd.n4338 240.244
R11455 gnd.n4336 gnd.n1872 240.244
R11456 gnd.n4332 gnd.n4331 240.244
R11457 gnd.n4329 gnd.n1879 240.244
R11458 gnd.n4325 gnd.n4324 240.244
R11459 gnd.n4322 gnd.n1886 240.244
R11460 gnd.n4318 gnd.n4317 240.244
R11461 gnd.n4315 gnd.n1893 240.244
R11462 gnd.n4311 gnd.n4310 240.244
R11463 gnd.n3706 gnd.n2096 240.244
R11464 gnd.n3689 gnd.n2096 240.244
R11465 gnd.n3689 gnd.n2088 240.244
R11466 gnd.n3698 gnd.n2088 240.244
R11467 gnd.n3698 gnd.n828 240.244
R11468 gnd.n3695 gnd.n828 240.244
R11469 gnd.n3695 gnd.n841 240.244
R11470 gnd.n3826 gnd.n841 240.244
R11471 gnd.n3826 gnd.n853 240.244
R11472 gnd.n2073 gnd.n853 240.244
R11473 gnd.n2073 gnd.n863 240.244
R11474 gnd.n3838 gnd.n863 240.244
R11475 gnd.n3838 gnd.n874 240.244
R11476 gnd.n2067 gnd.n874 240.244
R11477 gnd.n2067 gnd.n884 240.244
R11478 gnd.n3884 gnd.n884 240.244
R11479 gnd.n3884 gnd.n895 240.244
R11480 gnd.n3892 gnd.n895 240.244
R11481 gnd.n3892 gnd.n2056 240.244
R11482 gnd.n2056 gnd.n2048 240.244
R11483 gnd.n3929 gnd.n2048 240.244
R11484 gnd.n3929 gnd.n2029 240.244
R11485 gnd.n2029 gnd.n2022 240.244
R11486 gnd.n2044 gnd.n2022 240.244
R11487 gnd.n2044 gnd.n2015 240.244
R11488 gnd.n2015 gnd.n910 240.244
R11489 gnd.n2008 gnd.n910 240.244
R11490 gnd.n2008 gnd.n921 240.244
R11491 gnd.n3978 gnd.n921 240.244
R11492 gnd.n3978 gnd.n931 240.244
R11493 gnd.n1988 gnd.n931 240.244
R11494 gnd.n1988 gnd.n941 240.244
R11495 gnd.n3986 gnd.n941 240.244
R11496 gnd.n3986 gnd.n952 240.244
R11497 gnd.n3993 gnd.n952 240.244
R11498 gnd.n3993 gnd.n962 240.244
R11499 gnd.n3997 gnd.n962 240.244
R11500 gnd.n3997 gnd.n973 240.244
R11501 gnd.n4004 gnd.n973 240.244
R11502 gnd.n4004 gnd.n984 240.244
R11503 gnd.n4302 gnd.n984 240.244
R11504 gnd.n4302 gnd.n994 240.244
R11505 gnd.n3644 gnd.n3643 240.244
R11506 gnd.n3778 gnd.n3643 240.244
R11507 gnd.n3776 gnd.n3775 240.244
R11508 gnd.n3772 gnd.n3771 240.244
R11509 gnd.n3768 gnd.n3767 240.244
R11510 gnd.n3764 gnd.n3763 240.244
R11511 gnd.n3760 gnd.n3759 240.244
R11512 gnd.n3756 gnd.n3755 240.244
R11513 gnd.n3752 gnd.n3751 240.244
R11514 gnd.n3747 gnd.n3746 240.244
R11515 gnd.n3743 gnd.n3742 240.244
R11516 gnd.n3739 gnd.n3738 240.244
R11517 gnd.n3735 gnd.n3734 240.244
R11518 gnd.n3731 gnd.n3730 240.244
R11519 gnd.n3727 gnd.n3726 240.244
R11520 gnd.n3723 gnd.n3722 240.244
R11521 gnd.n3719 gnd.n3718 240.244
R11522 gnd.n3715 gnd.n3714 240.244
R11523 gnd.n3684 gnd.n3683 240.244
R11524 gnd.n3804 gnd.n2094 240.244
R11525 gnd.n3804 gnd.n2090 240.244
R11526 gnd.n3811 gnd.n2090 240.244
R11527 gnd.n3811 gnd.n832 240.244
R11528 gnd.n5945 gnd.n832 240.244
R11529 gnd.n5945 gnd.n833 240.244
R11530 gnd.n5941 gnd.n833 240.244
R11531 gnd.n5941 gnd.n839 240.244
R11532 gnd.n5933 gnd.n839 240.244
R11533 gnd.n5933 gnd.n855 240.244
R11534 gnd.n5929 gnd.n855 240.244
R11535 gnd.n5929 gnd.n861 240.244
R11536 gnd.n5921 gnd.n861 240.244
R11537 gnd.n5921 gnd.n877 240.244
R11538 gnd.n5917 gnd.n877 240.244
R11539 gnd.n5917 gnd.n883 240.244
R11540 gnd.n5909 gnd.n883 240.244
R11541 gnd.n5909 gnd.n897 240.244
R11542 gnd.n3919 gnd.n897 240.244
R11543 gnd.n3919 gnd.n3918 240.244
R11544 gnd.n3918 gnd.n2025 240.244
R11545 gnd.n3943 gnd.n2025 240.244
R11546 gnd.n3947 gnd.n3943 240.244
R11547 gnd.n3947 gnd.n3944 240.244
R11548 gnd.n3944 gnd.n907 240.244
R11549 gnd.n5903 gnd.n907 240.244
R11550 gnd.n5903 gnd.n908 240.244
R11551 gnd.n5895 gnd.n908 240.244
R11552 gnd.n5895 gnd.n924 240.244
R11553 gnd.n5891 gnd.n924 240.244
R11554 gnd.n5891 gnd.n929 240.244
R11555 gnd.n5883 gnd.n929 240.244
R11556 gnd.n5883 gnd.n944 240.244
R11557 gnd.n5879 gnd.n944 240.244
R11558 gnd.n5879 gnd.n950 240.244
R11559 gnd.n5871 gnd.n950 240.244
R11560 gnd.n5871 gnd.n965 240.244
R11561 gnd.n5867 gnd.n965 240.244
R11562 gnd.n5867 gnd.n971 240.244
R11563 gnd.n5859 gnd.n971 240.244
R11564 gnd.n5859 gnd.n987 240.244
R11565 gnd.n5855 gnd.n987 240.244
R11566 gnd.n3554 gnd.n2129 240.244
R11567 gnd.n3547 gnd.n3546 240.244
R11568 gnd.n3544 gnd.n3543 240.244
R11569 gnd.n3540 gnd.n3539 240.244
R11570 gnd.n3536 gnd.n3535 240.244
R11571 gnd.n3532 gnd.n3531 240.244
R11572 gnd.n3528 gnd.n3527 240.244
R11573 gnd.n3524 gnd.n3523 240.244
R11574 gnd.n2797 gnd.n2509 240.244
R11575 gnd.n2807 gnd.n2509 240.244
R11576 gnd.n2807 gnd.n2500 240.244
R11577 gnd.n2500 gnd.n2489 240.244
R11578 gnd.n2828 gnd.n2489 240.244
R11579 gnd.n2828 gnd.n2483 240.244
R11580 gnd.n2838 gnd.n2483 240.244
R11581 gnd.n2838 gnd.n2472 240.244
R11582 gnd.n2472 gnd.n2464 240.244
R11583 gnd.n2856 gnd.n2464 240.244
R11584 gnd.n2857 gnd.n2856 240.244
R11585 gnd.n2857 gnd.n2449 240.244
R11586 gnd.n2859 gnd.n2449 240.244
R11587 gnd.n2859 gnd.n2435 240.244
R11588 gnd.n2901 gnd.n2435 240.244
R11589 gnd.n2902 gnd.n2901 240.244
R11590 gnd.n2905 gnd.n2902 240.244
R11591 gnd.n2905 gnd.n2390 240.244
R11592 gnd.n2430 gnd.n2390 240.244
R11593 gnd.n2430 gnd.n2400 240.244
R11594 gnd.n2915 gnd.n2400 240.244
R11595 gnd.n2915 gnd.n2421 240.244
R11596 gnd.n2925 gnd.n2421 240.244
R11597 gnd.n2925 gnd.n2331 240.244
R11598 gnd.n2970 gnd.n2331 240.244
R11599 gnd.n2970 gnd.n2317 240.244
R11600 gnd.n2992 gnd.n2317 240.244
R11601 gnd.n2993 gnd.n2992 240.244
R11602 gnd.n2993 gnd.n2304 240.244
R11603 gnd.n2304 gnd.n2293 240.244
R11604 gnd.n3024 gnd.n2293 240.244
R11605 gnd.n3025 gnd.n3024 240.244
R11606 gnd.n3026 gnd.n3025 240.244
R11607 gnd.n3026 gnd.n2278 240.244
R11608 gnd.n2278 gnd.n2277 240.244
R11609 gnd.n2277 gnd.n2262 240.244
R11610 gnd.n3077 gnd.n2262 240.244
R11611 gnd.n3078 gnd.n3077 240.244
R11612 gnd.n3078 gnd.n2249 240.244
R11613 gnd.n2249 gnd.n2238 240.244
R11614 gnd.n3110 gnd.n2238 240.244
R11615 gnd.n3111 gnd.n3110 240.244
R11616 gnd.n3112 gnd.n3111 240.244
R11617 gnd.n3112 gnd.n2222 240.244
R11618 gnd.n2222 gnd.n2221 240.244
R11619 gnd.n2221 gnd.n2208 240.244
R11620 gnd.n3167 gnd.n2208 240.244
R11621 gnd.n3168 gnd.n3167 240.244
R11622 gnd.n3168 gnd.n2195 240.244
R11623 gnd.n2195 gnd.n2185 240.244
R11624 gnd.n3455 gnd.n2185 240.244
R11625 gnd.n3458 gnd.n3455 240.244
R11626 gnd.n3458 gnd.n3457 240.244
R11627 gnd.n2787 gnd.n2522 240.244
R11628 gnd.n2543 gnd.n2522 240.244
R11629 gnd.n2546 gnd.n2545 240.244
R11630 gnd.n2553 gnd.n2552 240.244
R11631 gnd.n2556 gnd.n2555 240.244
R11632 gnd.n2563 gnd.n2562 240.244
R11633 gnd.n2566 gnd.n2565 240.244
R11634 gnd.n2573 gnd.n2572 240.244
R11635 gnd.n2795 gnd.n2519 240.244
R11636 gnd.n2519 gnd.n2498 240.244
R11637 gnd.n2818 gnd.n2498 240.244
R11638 gnd.n2818 gnd.n2492 240.244
R11639 gnd.n2826 gnd.n2492 240.244
R11640 gnd.n2826 gnd.n2494 240.244
R11641 gnd.n2494 gnd.n2470 240.244
R11642 gnd.n2848 gnd.n2470 240.244
R11643 gnd.n2848 gnd.n2466 240.244
R11644 gnd.n2854 gnd.n2466 240.244
R11645 gnd.n2854 gnd.n2448 240.244
R11646 gnd.n2879 gnd.n2448 240.244
R11647 gnd.n2879 gnd.n2443 240.244
R11648 gnd.n2891 gnd.n2443 240.244
R11649 gnd.n2891 gnd.n2444 240.244
R11650 gnd.n2887 gnd.n2444 240.244
R11651 gnd.n2887 gnd.n2392 240.244
R11652 gnd.n2939 gnd.n2392 240.244
R11653 gnd.n2939 gnd.n2393 240.244
R11654 gnd.n2935 gnd.n2393 240.244
R11655 gnd.n2935 gnd.n2399 240.244
R11656 gnd.n2419 gnd.n2399 240.244
R11657 gnd.n2419 gnd.n2329 240.244
R11658 gnd.n2974 gnd.n2329 240.244
R11659 gnd.n2974 gnd.n2324 240.244
R11660 gnd.n2982 gnd.n2324 240.244
R11661 gnd.n2982 gnd.n2325 240.244
R11662 gnd.n2325 gnd.n2302 240.244
R11663 gnd.n3014 gnd.n2302 240.244
R11664 gnd.n3014 gnd.n2297 240.244
R11665 gnd.n3022 gnd.n2297 240.244
R11666 gnd.n3022 gnd.n2298 240.244
R11667 gnd.n2298 gnd.n2275 240.244
R11668 gnd.n3059 gnd.n2275 240.244
R11669 gnd.n3059 gnd.n2270 240.244
R11670 gnd.n3067 gnd.n2270 240.244
R11671 gnd.n3067 gnd.n2271 240.244
R11672 gnd.n2271 gnd.n2247 240.244
R11673 gnd.n3100 gnd.n2247 240.244
R11674 gnd.n3100 gnd.n2242 240.244
R11675 gnd.n3108 gnd.n2242 240.244
R11676 gnd.n3108 gnd.n2243 240.244
R11677 gnd.n2243 gnd.n2220 240.244
R11678 gnd.n3149 gnd.n2220 240.244
R11679 gnd.n3149 gnd.n2215 240.244
R11680 gnd.n3157 gnd.n2215 240.244
R11681 gnd.n3157 gnd.n2216 240.244
R11682 gnd.n2216 gnd.n2193 240.244
R11683 gnd.n3443 gnd.n2193 240.244
R11684 gnd.n3443 gnd.n2188 240.244
R11685 gnd.n3453 gnd.n2188 240.244
R11686 gnd.n3453 gnd.n2189 240.244
R11687 gnd.n2189 gnd.n2128 240.244
R11688 gnd.n2148 gnd.n2106 240.244
R11689 gnd.n3514 gnd.n3513 240.244
R11690 gnd.n3510 gnd.n3509 240.244
R11691 gnd.n3506 gnd.n3505 240.244
R11692 gnd.n3502 gnd.n3501 240.244
R11693 gnd.n3498 gnd.n3497 240.244
R11694 gnd.n3494 gnd.n3493 240.244
R11695 gnd.n3490 gnd.n3489 240.244
R11696 gnd.n3486 gnd.n3485 240.244
R11697 gnd.n3482 gnd.n3481 240.244
R11698 gnd.n3478 gnd.n3477 240.244
R11699 gnd.n3474 gnd.n3473 240.244
R11700 gnd.n3470 gnd.n3469 240.244
R11701 gnd.n2710 gnd.n2607 240.244
R11702 gnd.n2710 gnd.n2600 240.244
R11703 gnd.n2721 gnd.n2600 240.244
R11704 gnd.n2721 gnd.n2596 240.244
R11705 gnd.n2727 gnd.n2596 240.244
R11706 gnd.n2727 gnd.n2588 240.244
R11707 gnd.n2737 gnd.n2588 240.244
R11708 gnd.n2737 gnd.n2583 240.244
R11709 gnd.n2773 gnd.n2583 240.244
R11710 gnd.n2773 gnd.n2584 240.244
R11711 gnd.n2584 gnd.n2531 240.244
R11712 gnd.n2768 gnd.n2531 240.244
R11713 gnd.n2768 gnd.n2767 240.244
R11714 gnd.n2767 gnd.n2510 240.244
R11715 gnd.n2763 gnd.n2510 240.244
R11716 gnd.n2763 gnd.n2501 240.244
R11717 gnd.n2760 gnd.n2501 240.244
R11718 gnd.n2760 gnd.n2759 240.244
R11719 gnd.n2759 gnd.n2484 240.244
R11720 gnd.n2755 gnd.n2484 240.244
R11721 gnd.n2755 gnd.n2473 240.244
R11722 gnd.n2473 gnd.n2454 240.244
R11723 gnd.n2868 gnd.n2454 240.244
R11724 gnd.n2868 gnd.n2450 240.244
R11725 gnd.n2876 gnd.n2450 240.244
R11726 gnd.n2876 gnd.n2441 240.244
R11727 gnd.n2441 gnd.n2377 240.244
R11728 gnd.n2948 gnd.n2377 240.244
R11729 gnd.n2948 gnd.n2378 240.244
R11730 gnd.n2389 gnd.n2378 240.244
R11731 gnd.n2424 gnd.n2389 240.244
R11732 gnd.n2427 gnd.n2424 240.244
R11733 gnd.n2427 gnd.n2401 240.244
R11734 gnd.n2414 gnd.n2401 240.244
R11735 gnd.n2414 gnd.n2411 240.244
R11736 gnd.n2411 gnd.n2332 240.244
R11737 gnd.n2969 gnd.n2332 240.244
R11738 gnd.n2969 gnd.n2322 240.244
R11739 gnd.n2965 gnd.n2322 240.244
R11740 gnd.n2965 gnd.n2316 240.244
R11741 gnd.n2962 gnd.n2316 240.244
R11742 gnd.n2962 gnd.n2305 240.244
R11743 gnd.n2959 gnd.n2305 240.244
R11744 gnd.n2959 gnd.n2283 240.244
R11745 gnd.n3035 gnd.n2283 240.244
R11746 gnd.n3035 gnd.n2279 240.244
R11747 gnd.n3056 gnd.n2279 240.244
R11748 gnd.n3056 gnd.n2268 240.244
R11749 gnd.n3052 gnd.n2268 240.244
R11750 gnd.n3052 gnd.n2261 240.244
R11751 gnd.n3049 gnd.n2261 240.244
R11752 gnd.n3049 gnd.n2250 240.244
R11753 gnd.n3046 gnd.n2250 240.244
R11754 gnd.n3046 gnd.n2227 240.244
R11755 gnd.n3121 gnd.n2227 240.244
R11756 gnd.n3121 gnd.n2223 240.244
R11757 gnd.n3146 gnd.n2223 240.244
R11758 gnd.n3146 gnd.n2214 240.244
R11759 gnd.n3142 gnd.n2214 240.244
R11760 gnd.n3142 gnd.n2207 240.244
R11761 gnd.n3138 gnd.n2207 240.244
R11762 gnd.n3138 gnd.n2196 240.244
R11763 gnd.n3135 gnd.n2196 240.244
R11764 gnd.n3135 gnd.n2177 240.244
R11765 gnd.n3465 gnd.n2177 240.244
R11766 gnd.n2624 gnd.n2623 240.244
R11767 gnd.n2695 gnd.n2623 240.244
R11768 gnd.n2693 gnd.n2692 240.244
R11769 gnd.n2689 gnd.n2688 240.244
R11770 gnd.n2685 gnd.n2684 240.244
R11771 gnd.n2681 gnd.n2680 240.244
R11772 gnd.n2677 gnd.n2676 240.244
R11773 gnd.n2673 gnd.n2672 240.244
R11774 gnd.n2669 gnd.n2668 240.244
R11775 gnd.n2665 gnd.n2664 240.244
R11776 gnd.n2661 gnd.n2660 240.244
R11777 gnd.n2657 gnd.n2656 240.244
R11778 gnd.n2653 gnd.n2611 240.244
R11779 gnd.n2713 gnd.n2605 240.244
R11780 gnd.n2713 gnd.n2601 240.244
R11781 gnd.n2719 gnd.n2601 240.244
R11782 gnd.n2719 gnd.n2594 240.244
R11783 gnd.n2729 gnd.n2594 240.244
R11784 gnd.n2729 gnd.n2590 240.244
R11785 gnd.n2735 gnd.n2590 240.244
R11786 gnd.n2735 gnd.n2581 240.244
R11787 gnd.n2775 gnd.n2581 240.244
R11788 gnd.n2775 gnd.n2532 240.244
R11789 gnd.n2783 gnd.n2532 240.244
R11790 gnd.n2783 gnd.n2533 240.244
R11791 gnd.n2533 gnd.n2511 240.244
R11792 gnd.n2804 gnd.n2511 240.244
R11793 gnd.n2804 gnd.n2503 240.244
R11794 gnd.n2815 gnd.n2503 240.244
R11795 gnd.n2815 gnd.n2504 240.244
R11796 gnd.n2504 gnd.n2485 240.244
R11797 gnd.n2835 gnd.n2485 240.244
R11798 gnd.n2835 gnd.n2475 240.244
R11799 gnd.n2845 gnd.n2475 240.244
R11800 gnd.n2845 gnd.n2456 240.244
R11801 gnd.n2866 gnd.n2456 240.244
R11802 gnd.n2866 gnd.n2458 240.244
R11803 gnd.n2458 gnd.n2439 240.244
R11804 gnd.n2894 gnd.n2439 240.244
R11805 gnd.n2894 gnd.n2381 240.244
R11806 gnd.n2946 gnd.n2381 240.244
R11807 gnd.n2946 gnd.n2382 240.244
R11808 gnd.n2942 gnd.n2382 240.244
R11809 gnd.n2942 gnd.n2388 240.244
R11810 gnd.n2403 gnd.n2388 240.244
R11811 gnd.n2932 gnd.n2403 240.244
R11812 gnd.n2932 gnd.n2404 240.244
R11813 gnd.n2928 gnd.n2404 240.244
R11814 gnd.n2928 gnd.n2410 240.244
R11815 gnd.n2410 gnd.n2321 240.244
R11816 gnd.n2985 gnd.n2321 240.244
R11817 gnd.n2985 gnd.n2314 240.244
R11818 gnd.n2996 gnd.n2314 240.244
R11819 gnd.n2996 gnd.n2307 240.244
R11820 gnd.n3011 gnd.n2307 240.244
R11821 gnd.n3011 gnd.n2308 240.244
R11822 gnd.n2308 gnd.n2286 240.244
R11823 gnd.n3033 gnd.n2286 240.244
R11824 gnd.n3033 gnd.n2287 240.244
R11825 gnd.n2287 gnd.n2266 240.244
R11826 gnd.n3070 gnd.n2266 240.244
R11827 gnd.n3070 gnd.n2259 240.244
R11828 gnd.n3082 gnd.n2259 240.244
R11829 gnd.n3082 gnd.n2252 240.244
R11830 gnd.n3097 gnd.n2252 240.244
R11831 gnd.n3097 gnd.n2253 240.244
R11832 gnd.n2253 gnd.n2230 240.244
R11833 gnd.n3119 gnd.n2230 240.244
R11834 gnd.n3119 gnd.n2232 240.244
R11835 gnd.n2232 gnd.n2212 240.244
R11836 gnd.n3160 gnd.n2212 240.244
R11837 gnd.n3160 gnd.n2205 240.244
R11838 gnd.n3171 gnd.n2205 240.244
R11839 gnd.n3171 gnd.n2198 240.244
R11840 gnd.n3440 gnd.n2198 240.244
R11841 gnd.n3440 gnd.n2199 240.244
R11842 gnd.n2199 gnd.n2180 240.244
R11843 gnd.n3463 gnd.n2180 240.244
R11844 gnd.n6845 gnd.n6844 240.244
R11845 gnd.n6850 gnd.n6847 240.244
R11846 gnd.n6853 gnd.n6852 240.244
R11847 gnd.n6858 gnd.n6855 240.244
R11848 gnd.n6861 gnd.n6860 240.244
R11849 gnd.n6866 gnd.n6863 240.244
R11850 gnd.n6869 gnd.n6868 240.244
R11851 gnd.n6874 gnd.n6871 240.244
R11852 gnd.n6880 gnd.n6876 240.244
R11853 gnd.n5469 gnd.n1128 240.244
R11854 gnd.n5469 gnd.n1140 240.244
R11855 gnd.n5476 gnd.n1140 240.244
R11856 gnd.n5476 gnd.n1258 240.244
R11857 gnd.n1258 gnd.n1248 240.244
R11858 gnd.n5555 gnd.n1248 240.244
R11859 gnd.n5555 gnd.n1243 240.244
R11860 gnd.n5562 gnd.n1243 240.244
R11861 gnd.n5562 gnd.n1232 240.244
R11862 gnd.n1232 gnd.n1219 240.244
R11863 gnd.n5587 gnd.n1219 240.244
R11864 gnd.n5587 gnd.n1214 240.244
R11865 gnd.n5594 gnd.n1214 240.244
R11866 gnd.n5594 gnd.n1203 240.244
R11867 gnd.n1203 gnd.n1193 240.244
R11868 gnd.n5620 gnd.n1193 240.244
R11869 gnd.n5620 gnd.n1186 240.244
R11870 gnd.n5627 gnd.n1186 240.244
R11871 gnd.n5627 gnd.n1187 240.244
R11872 gnd.n1187 gnd.n1179 240.244
R11873 gnd.n1179 gnd.n1178 240.244
R11874 gnd.n1178 gnd.n54 240.244
R11875 gnd.n55 gnd.n54 240.244
R11876 gnd.n56 gnd.n55 240.244
R11877 gnd.n6776 gnd.n56 240.244
R11878 gnd.n6776 gnd.n59 240.244
R11879 gnd.n60 gnd.n59 240.244
R11880 gnd.n61 gnd.n60 240.244
R11881 gnd.n6767 gnd.n61 240.244
R11882 gnd.n6767 gnd.n64 240.244
R11883 gnd.n65 gnd.n64 240.244
R11884 gnd.n66 gnd.n65 240.244
R11885 gnd.n265 gnd.n66 240.244
R11886 gnd.n265 gnd.n69 240.244
R11887 gnd.n70 gnd.n69 240.244
R11888 gnd.n71 gnd.n70 240.244
R11889 gnd.n179 gnd.n71 240.244
R11890 gnd.n179 gnd.n74 240.244
R11891 gnd.n75 gnd.n74 240.244
R11892 gnd.n76 gnd.n75 240.244
R11893 gnd.n79 gnd.n76 240.244
R11894 gnd.n7007 gnd.n79 240.244
R11895 gnd.n5034 gnd.n5032 240.244
R11896 gnd.n5049 gnd.n5015 240.244
R11897 gnd.n5053 gnd.n5051 240.244
R11898 gnd.n5068 gnd.n5006 240.244
R11899 gnd.n5072 gnd.n5070 240.244
R11900 gnd.n5087 gnd.n4997 240.244
R11901 gnd.n5091 gnd.n5089 240.244
R11902 gnd.n5108 gnd.n4988 240.244
R11903 gnd.n5111 gnd.n5110 240.244
R11904 gnd.n1142 gnd.n1130 240.244
R11905 gnd.n5700 gnd.n1142 240.244
R11906 gnd.n5700 gnd.n1143 240.244
R11907 gnd.n1148 gnd.n1143 240.244
R11908 gnd.n1149 gnd.n1148 240.244
R11909 gnd.n1150 gnd.n1149 240.244
R11910 gnd.n1240 gnd.n1150 240.244
R11911 gnd.n1240 gnd.n1153 240.244
R11912 gnd.n1154 gnd.n1153 240.244
R11913 gnd.n1155 gnd.n1154 240.244
R11914 gnd.n1223 gnd.n1155 240.244
R11915 gnd.n1223 gnd.n1158 240.244
R11916 gnd.n1159 gnd.n1158 240.244
R11917 gnd.n1160 gnd.n1159 240.244
R11918 gnd.n1204 gnd.n1160 240.244
R11919 gnd.n1204 gnd.n1163 240.244
R11920 gnd.n1164 gnd.n1163 240.244
R11921 gnd.n1165 gnd.n1164 240.244
R11922 gnd.n1175 gnd.n1165 240.244
R11923 gnd.n1175 gnd.n1168 240.244
R11924 gnd.n1169 gnd.n1168 240.244
R11925 gnd.n5667 gnd.n1169 240.244
R11926 gnd.n5667 gnd.n230 240.244
R11927 gnd.n6789 gnd.n230 240.244
R11928 gnd.n6789 gnd.n226 240.244
R11929 gnd.n6795 gnd.n226 240.244
R11930 gnd.n6795 gnd.n208 240.244
R11931 gnd.n6805 gnd.n208 240.244
R11932 gnd.n6805 gnd.n204 240.244
R11933 gnd.n6811 gnd.n204 240.244
R11934 gnd.n6811 gnd.n193 240.244
R11935 gnd.n6821 gnd.n193 240.244
R11936 gnd.n6821 gnd.n189 240.244
R11937 gnd.n6827 gnd.n189 240.244
R11938 gnd.n6827 gnd.n176 240.244
R11939 gnd.n6837 gnd.n176 240.244
R11940 gnd.n6837 gnd.n170 240.244
R11941 gnd.n6917 gnd.n170 240.244
R11942 gnd.n6917 gnd.n171 240.244
R11943 gnd.n171 gnd.n162 240.244
R11944 gnd.n6842 gnd.n162 240.244
R11945 gnd.n6842 gnd.n84 240.244
R11946 gnd.n4080 gnd.n997 240.244
R11947 gnd.n4083 gnd.n4082 240.244
R11948 gnd.n4093 gnd.n4085 240.244
R11949 gnd.n4096 gnd.n4095 240.244
R11950 gnd.n4105 gnd.n4104 240.244
R11951 gnd.n4116 gnd.n4107 240.244
R11952 gnd.n4119 gnd.n4118 240.244
R11953 gnd.n4128 gnd.n4127 240.244
R11954 gnd.n4139 gnd.n4130 240.244
R11955 gnd.n3583 gnd.n2097 240.244
R11956 gnd.n2097 gnd.n2086 240.244
R11957 gnd.n3813 gnd.n2086 240.244
R11958 gnd.n3814 gnd.n3813 240.244
R11959 gnd.n3814 gnd.n829 240.244
R11960 gnd.n3817 gnd.n829 240.244
R11961 gnd.n3817 gnd.n842 240.244
R11962 gnd.n3824 gnd.n842 240.244
R11963 gnd.n3824 gnd.n854 240.244
R11964 gnd.n3844 gnd.n854 240.244
R11965 gnd.n3844 gnd.n864 240.244
R11966 gnd.n3840 gnd.n864 240.244
R11967 gnd.n3840 gnd.n875 240.244
R11968 gnd.n3874 gnd.n875 240.244
R11969 gnd.n3874 gnd.n885 240.244
R11970 gnd.n3882 gnd.n885 240.244
R11971 gnd.n3882 gnd.n896 240.244
R11972 gnd.n2054 gnd.n896 240.244
R11973 gnd.n3921 gnd.n2054 240.244
R11974 gnd.n3921 gnd.n2050 240.244
R11975 gnd.n3927 gnd.n2050 240.244
R11976 gnd.n3927 gnd.n2020 240.244
R11977 gnd.n3949 gnd.n2020 240.244
R11978 gnd.n3949 gnd.n2016 240.244
R11979 gnd.n3955 gnd.n2016 240.244
R11980 gnd.n3955 gnd.n911 240.244
R11981 gnd.n3970 gnd.n911 240.244
R11982 gnd.n3970 gnd.n922 240.244
R11983 gnd.n3976 gnd.n922 240.244
R11984 gnd.n3976 gnd.n932 240.244
R11985 gnd.n4021 gnd.n932 240.244
R11986 gnd.n4021 gnd.n942 240.244
R11987 gnd.n1993 gnd.n942 240.244
R11988 gnd.n1993 gnd.n953 240.244
R11989 gnd.n1994 gnd.n953 240.244
R11990 gnd.n1994 gnd.n963 240.244
R11991 gnd.n1997 gnd.n963 240.244
R11992 gnd.n1997 gnd.n974 240.244
R11993 gnd.n4006 gnd.n974 240.244
R11994 gnd.n4006 gnd.n985 240.244
R11995 gnd.n4300 gnd.n985 240.244
R11996 gnd.n4300 gnd.n995 240.244
R11997 gnd.n3595 gnd.n2104 240.244
R11998 gnd.n3599 gnd.n3598 240.244
R11999 gnd.n3605 gnd.n3604 240.244
R12000 gnd.n3609 gnd.n3608 240.244
R12001 gnd.n3615 gnd.n3614 240.244
R12002 gnd.n3619 gnd.n3618 240.244
R12003 gnd.n3625 gnd.n3624 240.244
R12004 gnd.n3629 gnd.n3628 240.244
R12005 gnd.n3642 gnd.n3582 240.244
R12006 gnd.n3802 gnd.n2098 240.244
R12007 gnd.n3802 gnd.n2099 240.244
R12008 gnd.n2099 gnd.n2089 240.244
R12009 gnd.n3795 gnd.n2089 240.244
R12010 gnd.n3795 gnd.n831 240.244
R12011 gnd.n844 gnd.n831 240.244
R12012 gnd.n5939 gnd.n844 240.244
R12013 gnd.n5939 gnd.n845 240.244
R12014 gnd.n5935 gnd.n845 240.244
R12015 gnd.n5935 gnd.n851 240.244
R12016 gnd.n5927 gnd.n851 240.244
R12017 gnd.n5927 gnd.n866 240.244
R12018 gnd.n5923 gnd.n866 240.244
R12019 gnd.n5923 gnd.n872 240.244
R12020 gnd.n5915 gnd.n872 240.244
R12021 gnd.n5915 gnd.n887 240.244
R12022 gnd.n5911 gnd.n887 240.244
R12023 gnd.n5911 gnd.n893 240.244
R12024 gnd.n3910 gnd.n893 240.244
R12025 gnd.n3916 gnd.n3910 240.244
R12026 gnd.n3916 gnd.n2030 240.244
R12027 gnd.n3941 gnd.n2030 240.244
R12028 gnd.n3941 gnd.n2024 240.244
R12029 gnd.n3937 gnd.n2024 240.244
R12030 gnd.n3937 gnd.n913 240.244
R12031 gnd.n5901 gnd.n913 240.244
R12032 gnd.n5901 gnd.n914 240.244
R12033 gnd.n5897 gnd.n914 240.244
R12034 gnd.n5897 gnd.n920 240.244
R12035 gnd.n5889 gnd.n920 240.244
R12036 gnd.n5889 gnd.n933 240.244
R12037 gnd.n5885 gnd.n933 240.244
R12038 gnd.n5885 gnd.n939 240.244
R12039 gnd.n5877 gnd.n939 240.244
R12040 gnd.n5877 gnd.n955 240.244
R12041 gnd.n5873 gnd.n955 240.244
R12042 gnd.n5873 gnd.n961 240.244
R12043 gnd.n5865 gnd.n961 240.244
R12044 gnd.n5865 gnd.n976 240.244
R12045 gnd.n5861 gnd.n976 240.244
R12046 gnd.n5861 gnd.n982 240.244
R12047 gnd.n5853 gnd.n982 240.244
R12048 gnd.n6122 gnd.n656 240.244
R12049 gnd.n6122 gnd.n654 240.244
R12050 gnd.n6126 gnd.n654 240.244
R12051 gnd.n6126 gnd.n650 240.244
R12052 gnd.n6132 gnd.n650 240.244
R12053 gnd.n6132 gnd.n648 240.244
R12054 gnd.n6136 gnd.n648 240.244
R12055 gnd.n6136 gnd.n644 240.244
R12056 gnd.n6142 gnd.n644 240.244
R12057 gnd.n6142 gnd.n642 240.244
R12058 gnd.n6146 gnd.n642 240.244
R12059 gnd.n6146 gnd.n638 240.244
R12060 gnd.n6152 gnd.n638 240.244
R12061 gnd.n6152 gnd.n636 240.244
R12062 gnd.n6156 gnd.n636 240.244
R12063 gnd.n6156 gnd.n632 240.244
R12064 gnd.n6162 gnd.n632 240.244
R12065 gnd.n6162 gnd.n630 240.244
R12066 gnd.n6166 gnd.n630 240.244
R12067 gnd.n6166 gnd.n626 240.244
R12068 gnd.n6172 gnd.n626 240.244
R12069 gnd.n6172 gnd.n624 240.244
R12070 gnd.n6176 gnd.n624 240.244
R12071 gnd.n6176 gnd.n620 240.244
R12072 gnd.n6182 gnd.n620 240.244
R12073 gnd.n6182 gnd.n618 240.244
R12074 gnd.n6186 gnd.n618 240.244
R12075 gnd.n6186 gnd.n614 240.244
R12076 gnd.n6192 gnd.n614 240.244
R12077 gnd.n6192 gnd.n612 240.244
R12078 gnd.n6196 gnd.n612 240.244
R12079 gnd.n6196 gnd.n608 240.244
R12080 gnd.n6202 gnd.n608 240.244
R12081 gnd.n6202 gnd.n606 240.244
R12082 gnd.n6206 gnd.n606 240.244
R12083 gnd.n6206 gnd.n602 240.244
R12084 gnd.n6212 gnd.n602 240.244
R12085 gnd.n6212 gnd.n600 240.244
R12086 gnd.n6216 gnd.n600 240.244
R12087 gnd.n6216 gnd.n596 240.244
R12088 gnd.n6222 gnd.n596 240.244
R12089 gnd.n6222 gnd.n594 240.244
R12090 gnd.n6226 gnd.n594 240.244
R12091 gnd.n6226 gnd.n590 240.244
R12092 gnd.n6232 gnd.n590 240.244
R12093 gnd.n6232 gnd.n588 240.244
R12094 gnd.n6236 gnd.n588 240.244
R12095 gnd.n6236 gnd.n584 240.244
R12096 gnd.n6242 gnd.n584 240.244
R12097 gnd.n6242 gnd.n582 240.244
R12098 gnd.n6246 gnd.n582 240.244
R12099 gnd.n6246 gnd.n578 240.244
R12100 gnd.n6252 gnd.n578 240.244
R12101 gnd.n6252 gnd.n576 240.244
R12102 gnd.n6256 gnd.n576 240.244
R12103 gnd.n6256 gnd.n572 240.244
R12104 gnd.n6262 gnd.n572 240.244
R12105 gnd.n6262 gnd.n570 240.244
R12106 gnd.n6266 gnd.n570 240.244
R12107 gnd.n6266 gnd.n566 240.244
R12108 gnd.n6272 gnd.n566 240.244
R12109 gnd.n6272 gnd.n564 240.244
R12110 gnd.n6276 gnd.n564 240.244
R12111 gnd.n6276 gnd.n560 240.244
R12112 gnd.n6282 gnd.n560 240.244
R12113 gnd.n6282 gnd.n558 240.244
R12114 gnd.n6286 gnd.n558 240.244
R12115 gnd.n6286 gnd.n554 240.244
R12116 gnd.n6292 gnd.n554 240.244
R12117 gnd.n6292 gnd.n552 240.244
R12118 gnd.n6296 gnd.n552 240.244
R12119 gnd.n6296 gnd.n548 240.244
R12120 gnd.n6302 gnd.n548 240.244
R12121 gnd.n6302 gnd.n546 240.244
R12122 gnd.n6306 gnd.n546 240.244
R12123 gnd.n6306 gnd.n542 240.244
R12124 gnd.n6312 gnd.n542 240.244
R12125 gnd.n6312 gnd.n540 240.244
R12126 gnd.n6316 gnd.n540 240.244
R12127 gnd.n6316 gnd.n536 240.244
R12128 gnd.n6322 gnd.n536 240.244
R12129 gnd.n6322 gnd.n534 240.244
R12130 gnd.n6326 gnd.n534 240.244
R12131 gnd.n6326 gnd.n530 240.244
R12132 gnd.n6332 gnd.n530 240.244
R12133 gnd.n6332 gnd.n528 240.244
R12134 gnd.n6336 gnd.n528 240.244
R12135 gnd.n6336 gnd.n524 240.244
R12136 gnd.n6342 gnd.n524 240.244
R12137 gnd.n6342 gnd.n522 240.244
R12138 gnd.n6346 gnd.n522 240.244
R12139 gnd.n6346 gnd.n518 240.244
R12140 gnd.n6352 gnd.n518 240.244
R12141 gnd.n6352 gnd.n516 240.244
R12142 gnd.n6356 gnd.n516 240.244
R12143 gnd.n6356 gnd.n512 240.244
R12144 gnd.n6362 gnd.n512 240.244
R12145 gnd.n6362 gnd.n510 240.244
R12146 gnd.n6366 gnd.n510 240.244
R12147 gnd.n6366 gnd.n506 240.244
R12148 gnd.n6372 gnd.n506 240.244
R12149 gnd.n6372 gnd.n504 240.244
R12150 gnd.n6376 gnd.n504 240.244
R12151 gnd.n6376 gnd.n500 240.244
R12152 gnd.n6382 gnd.n500 240.244
R12153 gnd.n6382 gnd.n498 240.244
R12154 gnd.n6386 gnd.n498 240.244
R12155 gnd.n6386 gnd.n494 240.244
R12156 gnd.n6392 gnd.n494 240.244
R12157 gnd.n6392 gnd.n492 240.244
R12158 gnd.n6396 gnd.n492 240.244
R12159 gnd.n6396 gnd.n488 240.244
R12160 gnd.n6402 gnd.n488 240.244
R12161 gnd.n6402 gnd.n486 240.244
R12162 gnd.n6406 gnd.n486 240.244
R12163 gnd.n6406 gnd.n482 240.244
R12164 gnd.n6412 gnd.n482 240.244
R12165 gnd.n6412 gnd.n480 240.244
R12166 gnd.n6416 gnd.n480 240.244
R12167 gnd.n6416 gnd.n476 240.244
R12168 gnd.n6422 gnd.n476 240.244
R12169 gnd.n6422 gnd.n474 240.244
R12170 gnd.n6426 gnd.n474 240.244
R12171 gnd.n6426 gnd.n470 240.244
R12172 gnd.n6432 gnd.n470 240.244
R12173 gnd.n6432 gnd.n468 240.244
R12174 gnd.n6436 gnd.n468 240.244
R12175 gnd.n6436 gnd.n464 240.244
R12176 gnd.n6442 gnd.n464 240.244
R12177 gnd.n6442 gnd.n462 240.244
R12178 gnd.n6446 gnd.n462 240.244
R12179 gnd.n6446 gnd.n458 240.244
R12180 gnd.n6452 gnd.n458 240.244
R12181 gnd.n6452 gnd.n456 240.244
R12182 gnd.n6456 gnd.n456 240.244
R12183 gnd.n6456 gnd.n452 240.244
R12184 gnd.n6462 gnd.n452 240.244
R12185 gnd.n6462 gnd.n450 240.244
R12186 gnd.n6466 gnd.n450 240.244
R12187 gnd.n6466 gnd.n446 240.244
R12188 gnd.n6472 gnd.n446 240.244
R12189 gnd.n6472 gnd.n444 240.244
R12190 gnd.n6476 gnd.n444 240.244
R12191 gnd.n6476 gnd.n440 240.244
R12192 gnd.n6482 gnd.n440 240.244
R12193 gnd.n6482 gnd.n438 240.244
R12194 gnd.n6486 gnd.n438 240.244
R12195 gnd.n6486 gnd.n434 240.244
R12196 gnd.n6492 gnd.n434 240.244
R12197 gnd.n6492 gnd.n432 240.244
R12198 gnd.n6496 gnd.n432 240.244
R12199 gnd.n6496 gnd.n428 240.244
R12200 gnd.n6502 gnd.n428 240.244
R12201 gnd.n6502 gnd.n426 240.244
R12202 gnd.n6506 gnd.n426 240.244
R12203 gnd.n6506 gnd.n422 240.244
R12204 gnd.n6512 gnd.n422 240.244
R12205 gnd.n6512 gnd.n420 240.244
R12206 gnd.n6516 gnd.n420 240.244
R12207 gnd.n6516 gnd.n416 240.244
R12208 gnd.n6522 gnd.n416 240.244
R12209 gnd.n6522 gnd.n414 240.244
R12210 gnd.n6526 gnd.n414 240.244
R12211 gnd.n6526 gnd.n410 240.244
R12212 gnd.n6532 gnd.n410 240.244
R12213 gnd.n6532 gnd.n408 240.244
R12214 gnd.n6536 gnd.n408 240.244
R12215 gnd.n6542 gnd.n404 240.244
R12216 gnd.n6542 gnd.n402 240.244
R12217 gnd.n6546 gnd.n402 240.244
R12218 gnd.n6546 gnd.n398 240.244
R12219 gnd.n6552 gnd.n398 240.244
R12220 gnd.n6552 gnd.n396 240.244
R12221 gnd.n6556 gnd.n396 240.244
R12222 gnd.n6556 gnd.n392 240.244
R12223 gnd.n6562 gnd.n392 240.244
R12224 gnd.n6562 gnd.n390 240.244
R12225 gnd.n6566 gnd.n390 240.244
R12226 gnd.n6566 gnd.n386 240.244
R12227 gnd.n6572 gnd.n386 240.244
R12228 gnd.n6572 gnd.n384 240.244
R12229 gnd.n6576 gnd.n384 240.244
R12230 gnd.n6576 gnd.n380 240.244
R12231 gnd.n6582 gnd.n380 240.244
R12232 gnd.n6582 gnd.n378 240.244
R12233 gnd.n6586 gnd.n378 240.244
R12234 gnd.n6586 gnd.n374 240.244
R12235 gnd.n6592 gnd.n374 240.244
R12236 gnd.n6592 gnd.n372 240.244
R12237 gnd.n6596 gnd.n372 240.244
R12238 gnd.n6596 gnd.n368 240.244
R12239 gnd.n6602 gnd.n368 240.244
R12240 gnd.n6602 gnd.n366 240.244
R12241 gnd.n6606 gnd.n366 240.244
R12242 gnd.n6606 gnd.n362 240.244
R12243 gnd.n6612 gnd.n362 240.244
R12244 gnd.n6612 gnd.n360 240.244
R12245 gnd.n6616 gnd.n360 240.244
R12246 gnd.n6616 gnd.n356 240.244
R12247 gnd.n6622 gnd.n356 240.244
R12248 gnd.n6622 gnd.n354 240.244
R12249 gnd.n6626 gnd.n354 240.244
R12250 gnd.n6626 gnd.n350 240.244
R12251 gnd.n6632 gnd.n350 240.244
R12252 gnd.n6632 gnd.n348 240.244
R12253 gnd.n6636 gnd.n348 240.244
R12254 gnd.n6636 gnd.n344 240.244
R12255 gnd.n6642 gnd.n344 240.244
R12256 gnd.n6642 gnd.n342 240.244
R12257 gnd.n6646 gnd.n342 240.244
R12258 gnd.n6646 gnd.n338 240.244
R12259 gnd.n6652 gnd.n338 240.244
R12260 gnd.n6652 gnd.n336 240.244
R12261 gnd.n6656 gnd.n336 240.244
R12262 gnd.n6656 gnd.n332 240.244
R12263 gnd.n6662 gnd.n332 240.244
R12264 gnd.n6662 gnd.n330 240.244
R12265 gnd.n6666 gnd.n330 240.244
R12266 gnd.n6666 gnd.n326 240.244
R12267 gnd.n6672 gnd.n326 240.244
R12268 gnd.n6672 gnd.n324 240.244
R12269 gnd.n6676 gnd.n324 240.244
R12270 gnd.n6676 gnd.n320 240.244
R12271 gnd.n6682 gnd.n320 240.244
R12272 gnd.n6682 gnd.n318 240.244
R12273 gnd.n6686 gnd.n318 240.244
R12274 gnd.n6686 gnd.n314 240.244
R12275 gnd.n6692 gnd.n314 240.244
R12276 gnd.n6692 gnd.n312 240.244
R12277 gnd.n6696 gnd.n312 240.244
R12278 gnd.n6696 gnd.n308 240.244
R12279 gnd.n6702 gnd.n308 240.244
R12280 gnd.n6702 gnd.n306 240.244
R12281 gnd.n6706 gnd.n306 240.244
R12282 gnd.n6706 gnd.n302 240.244
R12283 gnd.n6712 gnd.n302 240.244
R12284 gnd.n6712 gnd.n300 240.244
R12285 gnd.n6716 gnd.n300 240.244
R12286 gnd.n6716 gnd.n296 240.244
R12287 gnd.n6722 gnd.n296 240.244
R12288 gnd.n6722 gnd.n294 240.244
R12289 gnd.n6726 gnd.n294 240.244
R12290 gnd.n6726 gnd.n290 240.244
R12291 gnd.n6732 gnd.n290 240.244
R12292 gnd.n6732 gnd.n288 240.244
R12293 gnd.n6736 gnd.n288 240.244
R12294 gnd.n6736 gnd.n284 240.244
R12295 gnd.n6744 gnd.n284 240.244
R12296 gnd.n6744 gnd.n282 240.244
R12297 gnd.n6748 gnd.n282 240.244
R12298 gnd.n6749 gnd.n6748 240.244
R12299 gnd.n3853 gnd.n826 240.244
R12300 gnd.n3854 gnd.n3853 240.244
R12301 gnd.n3854 gnd.n3847 240.244
R12302 gnd.n3860 gnd.n3847 240.244
R12303 gnd.n3861 gnd.n3860 240.244
R12304 gnd.n3862 gnd.n3861 240.244
R12305 gnd.n3862 gnd.n2068 240.244
R12306 gnd.n3871 gnd.n2068 240.244
R12307 gnd.n3871 gnd.n2069 240.244
R12308 gnd.n2069 gnd.n2060 240.244
R12309 gnd.n3895 gnd.n2060 240.244
R12310 gnd.n3895 gnd.n2057 240.244
R12311 gnd.n3908 gnd.n2057 240.244
R12312 gnd.n3908 gnd.n2058 240.244
R12313 gnd.n3903 gnd.n2058 240.244
R12314 gnd.n3903 gnd.n3902 240.244
R12315 gnd.n3902 gnd.n2012 240.244
R12316 gnd.n3958 gnd.n2012 240.244
R12317 gnd.n3959 gnd.n3958 240.244
R12318 gnd.n3959 gnd.n2009 240.244
R12319 gnd.n3967 gnd.n2009 240.244
R12320 gnd.n3967 gnd.n2010 240.244
R12321 gnd.n2010 gnd.n1987 240.244
R12322 gnd.n4024 gnd.n1987 240.244
R12323 gnd.n4024 gnd.n1983 240.244
R12324 gnd.n4030 gnd.n1983 240.244
R12325 gnd.n4031 gnd.n4030 240.244
R12326 gnd.n4032 gnd.n4031 240.244
R12327 gnd.n4032 gnd.n1979 240.244
R12328 gnd.n4038 gnd.n1979 240.244
R12329 gnd.n4039 gnd.n4038 240.244
R12330 gnd.n4040 gnd.n4039 240.244
R12331 gnd.n4040 gnd.n1975 240.244
R12332 gnd.n4046 gnd.n1975 240.244
R12333 gnd.n4047 gnd.n4046 240.244
R12334 gnd.n4048 gnd.n4047 240.244
R12335 gnd.n4048 gnd.n1971 240.244
R12336 gnd.n4054 gnd.n1971 240.244
R12337 gnd.n4054 gnd.n1969 240.244
R12338 gnd.n4191 gnd.n1969 240.244
R12339 gnd.n4191 gnd.n1965 240.244
R12340 gnd.n4197 gnd.n1965 240.244
R12341 gnd.n4197 gnd.n1963 240.244
R12342 gnd.n4205 gnd.n1963 240.244
R12343 gnd.n4205 gnd.n1959 240.244
R12344 gnd.n4211 gnd.n1959 240.244
R12345 gnd.n4211 gnd.n1955 240.244
R12346 gnd.n4219 gnd.n1955 240.244
R12347 gnd.n4219 gnd.n1951 240.244
R12348 gnd.n4225 gnd.n1951 240.244
R12349 gnd.n4225 gnd.n1947 240.244
R12350 gnd.n4233 gnd.n1947 240.244
R12351 gnd.n4233 gnd.n1943 240.244
R12352 gnd.n4239 gnd.n1943 240.244
R12353 gnd.n4239 gnd.n1670 240.244
R12354 gnd.n4422 gnd.n1670 240.244
R12355 gnd.n4422 gnd.n1666 240.244
R12356 gnd.n4428 gnd.n1666 240.244
R12357 gnd.n4428 gnd.n1652 240.244
R12358 gnd.n4478 gnd.n1652 240.244
R12359 gnd.n4478 gnd.n1648 240.244
R12360 gnd.n4484 gnd.n1648 240.244
R12361 gnd.n4484 gnd.n1631 240.244
R12362 gnd.n4509 gnd.n1631 240.244
R12363 gnd.n4509 gnd.n1627 240.244
R12364 gnd.n4517 gnd.n1627 240.244
R12365 gnd.n4517 gnd.n1611 240.244
R12366 gnd.n4538 gnd.n1611 240.244
R12367 gnd.n4539 gnd.n4538 240.244
R12368 gnd.n4539 gnd.n1606 240.244
R12369 gnd.n4555 gnd.n1606 240.244
R12370 gnd.n4555 gnd.n1607 240.244
R12371 gnd.n4551 gnd.n1607 240.244
R12372 gnd.n4551 gnd.n4550 240.244
R12373 gnd.n4550 gnd.n1564 240.244
R12374 gnd.n4623 gnd.n1564 240.244
R12375 gnd.n4623 gnd.n1560 240.244
R12376 gnd.n4629 gnd.n1560 240.244
R12377 gnd.n4629 gnd.n1541 240.244
R12378 gnd.n4663 gnd.n1541 240.244
R12379 gnd.n4663 gnd.n1537 240.244
R12380 gnd.n4669 gnd.n1537 240.244
R12381 gnd.n4669 gnd.n1519 240.244
R12382 gnd.n4717 gnd.n1519 240.244
R12383 gnd.n4717 gnd.n1515 240.244
R12384 gnd.n4723 gnd.n1515 240.244
R12385 gnd.n4723 gnd.n1500 240.244
R12386 gnd.n4742 gnd.n1500 240.244
R12387 gnd.n4742 gnd.n1496 240.244
R12388 gnd.n4748 gnd.n1496 240.244
R12389 gnd.n4748 gnd.n1478 240.244
R12390 gnd.n4801 gnd.n1478 240.244
R12391 gnd.n4801 gnd.n1474 240.244
R12392 gnd.n4807 gnd.n1474 240.244
R12393 gnd.n4807 gnd.n1456 240.244
R12394 gnd.n4830 gnd.n1456 240.244
R12395 gnd.n4830 gnd.n1451 240.244
R12396 gnd.n4838 gnd.n1451 240.244
R12397 gnd.n4838 gnd.n1452 240.244
R12398 gnd.n1452 gnd.n1428 240.244
R12399 gnd.n4885 gnd.n1428 240.244
R12400 gnd.n4885 gnd.n1424 240.244
R12401 gnd.n4891 gnd.n1424 240.244
R12402 gnd.n4891 gnd.n1411 240.244
R12403 gnd.n4911 gnd.n1411 240.244
R12404 gnd.n4911 gnd.n1405 240.244
R12405 gnd.n4920 gnd.n1405 240.244
R12406 gnd.n4920 gnd.n1407 240.244
R12407 gnd.n1407 gnd.n1344 240.244
R12408 gnd.n5190 gnd.n1344 240.244
R12409 gnd.n5190 gnd.n1345 240.244
R12410 gnd.n5186 gnd.n1345 240.244
R12411 gnd.n5186 gnd.n5185 240.244
R12412 gnd.n5185 gnd.n1351 240.244
R12413 gnd.n5178 gnd.n1351 240.244
R12414 gnd.n5178 gnd.n1355 240.244
R12415 gnd.n5174 gnd.n1355 240.244
R12416 gnd.n5174 gnd.n1363 240.244
R12417 gnd.n5167 gnd.n1363 240.244
R12418 gnd.n5167 gnd.n1369 240.244
R12419 gnd.n5163 gnd.n1369 240.244
R12420 gnd.n5163 gnd.n1375 240.244
R12421 gnd.n5156 gnd.n1375 240.244
R12422 gnd.n5156 gnd.n1109 240.244
R12423 gnd.n5721 gnd.n1109 240.244
R12424 gnd.n5721 gnd.n1110 240.244
R12425 gnd.n5717 gnd.n1110 240.244
R12426 gnd.n5717 gnd.n1116 240.244
R12427 gnd.n5713 gnd.n1116 240.244
R12428 gnd.n5713 gnd.n1119 240.244
R12429 gnd.n5709 gnd.n1119 240.244
R12430 gnd.n5709 gnd.n1125 240.244
R12431 gnd.n5533 gnd.n1125 240.244
R12432 gnd.n5534 gnd.n5533 240.244
R12433 gnd.n5534 gnd.n5527 240.244
R12434 gnd.n5542 gnd.n5527 240.244
R12435 gnd.n5542 gnd.n5528 240.244
R12436 gnd.n5528 gnd.n1239 240.244
R12437 gnd.n5565 gnd.n1239 240.244
R12438 gnd.n5565 gnd.n1234 240.244
R12439 gnd.n5573 gnd.n1234 240.244
R12440 gnd.n5573 gnd.n1235 240.244
R12441 gnd.n1235 gnd.n1211 240.244
R12442 gnd.n5597 gnd.n1211 240.244
R12443 gnd.n5597 gnd.n1206 240.244
R12444 gnd.n5611 gnd.n1206 240.244
R12445 gnd.n5611 gnd.n1207 240.244
R12446 gnd.n5607 gnd.n1207 240.244
R12447 gnd.n5607 gnd.n5606 240.244
R12448 gnd.n5606 gnd.n1174 240.244
R12449 gnd.n5640 gnd.n1174 240.244
R12450 gnd.n5640 gnd.n1171 240.244
R12451 gnd.n5664 gnd.n1171 240.244
R12452 gnd.n5664 gnd.n1172 240.244
R12453 gnd.n5659 gnd.n1172 240.244
R12454 gnd.n5659 gnd.n5658 240.244
R12455 gnd.n5658 gnd.n5657 240.244
R12456 gnd.n5657 gnd.n5645 240.244
R12457 gnd.n5653 gnd.n5645 240.244
R12458 gnd.n5653 gnd.n5652 240.244
R12459 gnd.n5652 gnd.n270 240.244
R12460 gnd.n6761 gnd.n270 240.244
R12461 gnd.n6761 gnd.n271 240.244
R12462 gnd.n6757 gnd.n271 240.244
R12463 gnd.n6757 gnd.n6756 240.244
R12464 gnd.n6756 gnd.n6755 240.244
R12465 gnd.n6755 gnd.n277 240.244
R12466 gnd.n6116 gnd.n660 240.244
R12467 gnd.n6112 gnd.n660 240.244
R12468 gnd.n6112 gnd.n662 240.244
R12469 gnd.n6108 gnd.n662 240.244
R12470 gnd.n6108 gnd.n667 240.244
R12471 gnd.n6104 gnd.n667 240.244
R12472 gnd.n6104 gnd.n669 240.244
R12473 gnd.n6100 gnd.n669 240.244
R12474 gnd.n6100 gnd.n675 240.244
R12475 gnd.n6096 gnd.n675 240.244
R12476 gnd.n6096 gnd.n677 240.244
R12477 gnd.n6092 gnd.n677 240.244
R12478 gnd.n6092 gnd.n683 240.244
R12479 gnd.n6088 gnd.n683 240.244
R12480 gnd.n6088 gnd.n685 240.244
R12481 gnd.n6084 gnd.n685 240.244
R12482 gnd.n6084 gnd.n691 240.244
R12483 gnd.n6080 gnd.n691 240.244
R12484 gnd.n6080 gnd.n693 240.244
R12485 gnd.n6076 gnd.n693 240.244
R12486 gnd.n6076 gnd.n699 240.244
R12487 gnd.n6072 gnd.n699 240.244
R12488 gnd.n6072 gnd.n701 240.244
R12489 gnd.n6068 gnd.n701 240.244
R12490 gnd.n6068 gnd.n707 240.244
R12491 gnd.n6064 gnd.n707 240.244
R12492 gnd.n6064 gnd.n709 240.244
R12493 gnd.n6060 gnd.n709 240.244
R12494 gnd.n6060 gnd.n715 240.244
R12495 gnd.n6056 gnd.n715 240.244
R12496 gnd.n6056 gnd.n717 240.244
R12497 gnd.n6052 gnd.n717 240.244
R12498 gnd.n6052 gnd.n723 240.244
R12499 gnd.n6048 gnd.n723 240.244
R12500 gnd.n6048 gnd.n725 240.244
R12501 gnd.n6044 gnd.n725 240.244
R12502 gnd.n6044 gnd.n731 240.244
R12503 gnd.n6040 gnd.n731 240.244
R12504 gnd.n6040 gnd.n733 240.244
R12505 gnd.n6036 gnd.n733 240.244
R12506 gnd.n6036 gnd.n739 240.244
R12507 gnd.n6032 gnd.n739 240.244
R12508 gnd.n6032 gnd.n741 240.244
R12509 gnd.n6028 gnd.n741 240.244
R12510 gnd.n6028 gnd.n747 240.244
R12511 gnd.n6024 gnd.n747 240.244
R12512 gnd.n6024 gnd.n749 240.244
R12513 gnd.n6020 gnd.n749 240.244
R12514 gnd.n6020 gnd.n755 240.244
R12515 gnd.n6016 gnd.n755 240.244
R12516 gnd.n6016 gnd.n757 240.244
R12517 gnd.n6012 gnd.n757 240.244
R12518 gnd.n6012 gnd.n763 240.244
R12519 gnd.n6008 gnd.n763 240.244
R12520 gnd.n6008 gnd.n765 240.244
R12521 gnd.n6004 gnd.n765 240.244
R12522 gnd.n6004 gnd.n771 240.244
R12523 gnd.n6000 gnd.n771 240.244
R12524 gnd.n6000 gnd.n773 240.244
R12525 gnd.n5996 gnd.n773 240.244
R12526 gnd.n5996 gnd.n779 240.244
R12527 gnd.n5992 gnd.n779 240.244
R12528 gnd.n5992 gnd.n781 240.244
R12529 gnd.n5988 gnd.n781 240.244
R12530 gnd.n5988 gnd.n787 240.244
R12531 gnd.n5984 gnd.n787 240.244
R12532 gnd.n5984 gnd.n789 240.244
R12533 gnd.n5980 gnd.n789 240.244
R12534 gnd.n5980 gnd.n795 240.244
R12535 gnd.n5976 gnd.n795 240.244
R12536 gnd.n5976 gnd.n797 240.244
R12537 gnd.n5972 gnd.n797 240.244
R12538 gnd.n5972 gnd.n803 240.244
R12539 gnd.n5968 gnd.n803 240.244
R12540 gnd.n5968 gnd.n805 240.244
R12541 gnd.n5964 gnd.n805 240.244
R12542 gnd.n5964 gnd.n811 240.244
R12543 gnd.n5960 gnd.n811 240.244
R12544 gnd.n5960 gnd.n813 240.244
R12545 gnd.n5956 gnd.n813 240.244
R12546 gnd.n5956 gnd.n819 240.244
R12547 gnd.n5952 gnd.n819 240.244
R12548 gnd.n5952 gnd.n821 240.244
R12549 gnd.n5948 gnd.n821 240.244
R12550 gnd.n1003 gnd.n1002 240.244
R12551 gnd.n1004 gnd.n1003 240.244
R12552 gnd.n1957 gnd.n1004 240.244
R12553 gnd.n1957 gnd.n1007 240.244
R12554 gnd.n1008 gnd.n1007 240.244
R12555 gnd.n1009 gnd.n1008 240.244
R12556 gnd.n1949 gnd.n1009 240.244
R12557 gnd.n1949 gnd.n1012 240.244
R12558 gnd.n1013 gnd.n1012 240.244
R12559 gnd.n1014 gnd.n1013 240.244
R12560 gnd.n4241 gnd.n1014 240.244
R12561 gnd.n4241 gnd.n1017 240.244
R12562 gnd.n1018 gnd.n1017 240.244
R12563 gnd.n1019 gnd.n1018 240.244
R12564 gnd.n1664 gnd.n1019 240.244
R12565 gnd.n1664 gnd.n1022 240.244
R12566 gnd.n1023 gnd.n1022 240.244
R12567 gnd.n1024 gnd.n1023 240.244
R12568 gnd.n4486 gnd.n1024 240.244
R12569 gnd.n4486 gnd.n1027 240.244
R12570 gnd.n1028 gnd.n1027 240.244
R12571 gnd.n1029 gnd.n1028 240.244
R12572 gnd.n4519 gnd.n1029 240.244
R12573 gnd.n4519 gnd.n1032 240.244
R12574 gnd.n1033 gnd.n1032 240.244
R12575 gnd.n1034 gnd.n1033 240.244
R12576 gnd.n4564 gnd.n1034 240.244
R12577 gnd.n4564 gnd.n1037 240.244
R12578 gnd.n1038 gnd.n1037 240.244
R12579 gnd.n1039 gnd.n1038 240.244
R12580 gnd.n4592 gnd.n1039 240.244
R12581 gnd.n4592 gnd.n1042 240.244
R12582 gnd.n1043 gnd.n1042 240.244
R12583 gnd.n1044 gnd.n1043 240.244
R12584 gnd.n4603 gnd.n1044 240.244
R12585 gnd.n4603 gnd.n1047 240.244
R12586 gnd.n1048 gnd.n1047 240.244
R12587 gnd.n1049 gnd.n1048 240.244
R12588 gnd.n4642 gnd.n1049 240.244
R12589 gnd.n4642 gnd.n1052 240.244
R12590 gnd.n1053 gnd.n1052 240.244
R12591 gnd.n1054 gnd.n1053 240.244
R12592 gnd.n4683 gnd.n1054 240.244
R12593 gnd.n4683 gnd.n1057 240.244
R12594 gnd.n1058 gnd.n1057 240.244
R12595 gnd.n1059 gnd.n1058 240.244
R12596 gnd.n4751 gnd.n1059 240.244
R12597 gnd.n4751 gnd.n1062 240.244
R12598 gnd.n1063 gnd.n1062 240.244
R12599 gnd.n1064 gnd.n1063 240.244
R12600 gnd.n4809 gnd.n1064 240.244
R12601 gnd.n4809 gnd.n1067 240.244
R12602 gnd.n1068 gnd.n1067 240.244
R12603 gnd.n1069 gnd.n1068 240.244
R12604 gnd.n4840 gnd.n1069 240.244
R12605 gnd.n4840 gnd.n1072 240.244
R12606 gnd.n1073 gnd.n1072 240.244
R12607 gnd.n1074 gnd.n1073 240.244
R12608 gnd.n4882 gnd.n1074 240.244
R12609 gnd.n4882 gnd.n1077 240.244
R12610 gnd.n1078 gnd.n1077 240.244
R12611 gnd.n1079 gnd.n1078 240.244
R12612 gnd.n4908 gnd.n1079 240.244
R12613 gnd.n4908 gnd.n1082 240.244
R12614 gnd.n1083 gnd.n1082 240.244
R12615 gnd.n1084 gnd.n1083 240.244
R12616 gnd.n1340 gnd.n1084 240.244
R12617 gnd.n1340 gnd.n1087 240.244
R12618 gnd.n1088 gnd.n1087 240.244
R12619 gnd.n1089 gnd.n1088 240.244
R12620 gnd.n5182 gnd.n1089 240.244
R12621 gnd.n5182 gnd.n1092 240.244
R12622 gnd.n1093 gnd.n1092 240.244
R12623 gnd.n1094 gnd.n1093 240.244
R12624 gnd.n5171 gnd.n1094 240.244
R12625 gnd.n5171 gnd.n1097 240.244
R12626 gnd.n1098 gnd.n1097 240.244
R12627 gnd.n1099 gnd.n1098 240.244
R12628 gnd.n5160 gnd.n1099 240.244
R12629 gnd.n5160 gnd.n1102 240.244
R12630 gnd.n1103 gnd.n1102 240.244
R12631 gnd.n5724 gnd.n1103 240.244
R12632 gnd.n4073 gnd.n4072 240.244
R12633 gnd.n4088 gnd.n4072 240.244
R12634 gnd.n4090 gnd.n4089 240.244
R12635 gnd.n4100 gnd.n4099 240.244
R12636 gnd.n4111 gnd.n4110 240.244
R12637 gnd.n4113 gnd.n4112 240.244
R12638 gnd.n4123 gnd.n4122 240.244
R12639 gnd.n4136 gnd.n4135 240.244
R12640 gnd.n4138 gnd.n4137 240.244
R12641 gnd.n1912 gnd.n1911 240.244
R12642 gnd.n4066 gnd.n1913 240.244
R12643 gnd.n1917 gnd.n1916 240.244
R12644 gnd.n1923 gnd.n1918 240.244
R12645 gnd.n1925 gnd.n1924 240.244
R12646 gnd.n1929 gnd.n1928 240.244
R12647 gnd.n1930 gnd.n1929 240.244
R12648 gnd.n1956 gnd.n1930 240.244
R12649 gnd.n1956 gnd.n1933 240.244
R12650 gnd.n1934 gnd.n1933 240.244
R12651 gnd.n1935 gnd.n1934 240.244
R12652 gnd.n1948 gnd.n1935 240.244
R12653 gnd.n1948 gnd.n1938 240.244
R12654 gnd.n1939 gnd.n1938 240.244
R12655 gnd.n1940 gnd.n1939 240.244
R12656 gnd.n4243 gnd.n1940 240.244
R12657 gnd.n4244 gnd.n4243 240.244
R12658 gnd.n4246 gnd.n4244 240.244
R12659 gnd.n4246 gnd.n1672 240.244
R12660 gnd.n4249 gnd.n1672 240.244
R12661 gnd.n4250 gnd.n4249 240.244
R12662 gnd.n4251 gnd.n4250 240.244
R12663 gnd.n4251 gnd.n1644 240.244
R12664 gnd.n4488 gnd.n1644 240.244
R12665 gnd.n4488 gnd.n1640 240.244
R12666 gnd.n4494 gnd.n1640 240.244
R12667 gnd.n4494 gnd.n1624 240.244
R12668 gnd.n4521 gnd.n1624 240.244
R12669 gnd.n4521 gnd.n1620 240.244
R12670 gnd.n4527 gnd.n1620 240.244
R12671 gnd.n4527 gnd.n1598 240.244
R12672 gnd.n4566 gnd.n1598 240.244
R12673 gnd.n4566 gnd.n1593 240.244
R12674 gnd.n4574 gnd.n1593 240.244
R12675 gnd.n4574 gnd.n1582 240.244
R12676 gnd.n4594 gnd.n1582 240.244
R12677 gnd.n4595 gnd.n4594 240.244
R12678 gnd.n4596 gnd.n4595 240.244
R12679 gnd.n4596 gnd.n1578 240.244
R12680 gnd.n4602 gnd.n1578 240.244
R12681 gnd.n4602 gnd.n1551 240.244
R12682 gnd.n4650 gnd.n1551 240.244
R12683 gnd.n4650 gnd.n1552 240.244
R12684 gnd.n4644 gnd.n1552 240.244
R12685 gnd.n4644 gnd.n1529 240.244
R12686 gnd.n4706 gnd.n1529 240.244
R12687 gnd.n4706 gnd.n1521 240.244
R12688 gnd.n4685 gnd.n1521 240.244
R12689 gnd.n4686 gnd.n4685 240.244
R12690 gnd.n4687 gnd.n4686 240.244
R12691 gnd.n4687 gnd.n1502 240.244
R12692 gnd.n1502 gnd.n1495 240.244
R12693 gnd.n4690 gnd.n1495 240.244
R12694 gnd.n4691 gnd.n4690 240.244
R12695 gnd.n4691 gnd.n1471 240.244
R12696 gnd.n4811 gnd.n1471 240.244
R12697 gnd.n4811 gnd.n1465 240.244
R12698 gnd.n4818 gnd.n1465 240.244
R12699 gnd.n4818 gnd.n1466 240.244
R12700 gnd.n1466 gnd.n1443 240.244
R12701 gnd.n4850 gnd.n1443 240.244
R12702 gnd.n4850 gnd.n1438 240.244
R12703 gnd.n4873 gnd.n1438 240.244
R12704 gnd.n4873 gnd.n1430 240.244
R12705 gnd.n4855 gnd.n1430 240.244
R12706 gnd.n4858 gnd.n4855 240.244
R12707 gnd.n4860 gnd.n4858 240.244
R12708 gnd.n4860 gnd.n1413 240.244
R12709 gnd.n1413 gnd.n1403 240.244
R12710 gnd.n1403 gnd.n1392 240.244
R12711 gnd.n4941 gnd.n1392 240.244
R12712 gnd.n4941 gnd.n1388 240.244
R12713 gnd.n4949 gnd.n1388 240.244
R12714 gnd.n4950 gnd.n4949 240.244
R12715 gnd.n4951 gnd.n4950 240.244
R12716 gnd.n4951 gnd.n1352 240.244
R12717 gnd.n1353 gnd.n1352 240.244
R12718 gnd.n4958 gnd.n1353 240.244
R12719 gnd.n4959 gnd.n4958 240.244
R12720 gnd.n4959 gnd.n1366 240.244
R12721 gnd.n1367 gnd.n1366 240.244
R12722 gnd.n4966 gnd.n1367 240.244
R12723 gnd.n4967 gnd.n4966 240.244
R12724 gnd.n4967 gnd.n1378 240.244
R12725 gnd.n1379 gnd.n1378 240.244
R12726 gnd.n5150 gnd.n1379 240.244
R12727 gnd.n5150 gnd.n1107 240.244
R12728 gnd.n5041 gnd.n5040 240.244
R12729 gnd.n5044 gnd.n5043 240.244
R12730 gnd.n5060 gnd.n5059 240.244
R12731 gnd.n5063 gnd.n5062 240.244
R12732 gnd.n5079 gnd.n5078 240.244
R12733 gnd.n5082 gnd.n5081 240.244
R12734 gnd.n5098 gnd.n5097 240.244
R12735 gnd.n5102 gnd.n5100 240.244
R12736 gnd.n5118 gnd.n4982 240.244
R12737 gnd.n5122 gnd.n5120 240.244
R12738 gnd.n5128 gnd.n4978 240.244
R12739 gnd.n5132 gnd.n5130 240.244
R12740 gnd.n5141 gnd.n4974 240.244
R12741 gnd.n5144 gnd.n5143 240.244
R12742 gnd.n1684 gnd.n1683 240.132
R12743 gnd.n5207 gnd.n5206 240.132
R12744 gnd.n6123 gnd.n655 225.874
R12745 gnd.n6124 gnd.n6123 225.874
R12746 gnd.n6125 gnd.n6124 225.874
R12747 gnd.n6125 gnd.n649 225.874
R12748 gnd.n6133 gnd.n649 225.874
R12749 gnd.n6134 gnd.n6133 225.874
R12750 gnd.n6135 gnd.n6134 225.874
R12751 gnd.n6135 gnd.n643 225.874
R12752 gnd.n6143 gnd.n643 225.874
R12753 gnd.n6144 gnd.n6143 225.874
R12754 gnd.n6145 gnd.n6144 225.874
R12755 gnd.n6145 gnd.n637 225.874
R12756 gnd.n6153 gnd.n637 225.874
R12757 gnd.n6154 gnd.n6153 225.874
R12758 gnd.n6155 gnd.n6154 225.874
R12759 gnd.n6155 gnd.n631 225.874
R12760 gnd.n6163 gnd.n631 225.874
R12761 gnd.n6164 gnd.n6163 225.874
R12762 gnd.n6165 gnd.n6164 225.874
R12763 gnd.n6165 gnd.n625 225.874
R12764 gnd.n6173 gnd.n625 225.874
R12765 gnd.n6174 gnd.n6173 225.874
R12766 gnd.n6175 gnd.n6174 225.874
R12767 gnd.n6175 gnd.n619 225.874
R12768 gnd.n6183 gnd.n619 225.874
R12769 gnd.n6184 gnd.n6183 225.874
R12770 gnd.n6185 gnd.n6184 225.874
R12771 gnd.n6185 gnd.n613 225.874
R12772 gnd.n6193 gnd.n613 225.874
R12773 gnd.n6194 gnd.n6193 225.874
R12774 gnd.n6195 gnd.n6194 225.874
R12775 gnd.n6195 gnd.n607 225.874
R12776 gnd.n6203 gnd.n607 225.874
R12777 gnd.n6204 gnd.n6203 225.874
R12778 gnd.n6205 gnd.n6204 225.874
R12779 gnd.n6205 gnd.n601 225.874
R12780 gnd.n6213 gnd.n601 225.874
R12781 gnd.n6214 gnd.n6213 225.874
R12782 gnd.n6215 gnd.n6214 225.874
R12783 gnd.n6215 gnd.n595 225.874
R12784 gnd.n6223 gnd.n595 225.874
R12785 gnd.n6224 gnd.n6223 225.874
R12786 gnd.n6225 gnd.n6224 225.874
R12787 gnd.n6225 gnd.n589 225.874
R12788 gnd.n6233 gnd.n589 225.874
R12789 gnd.n6234 gnd.n6233 225.874
R12790 gnd.n6235 gnd.n6234 225.874
R12791 gnd.n6235 gnd.n583 225.874
R12792 gnd.n6243 gnd.n583 225.874
R12793 gnd.n6244 gnd.n6243 225.874
R12794 gnd.n6245 gnd.n6244 225.874
R12795 gnd.n6245 gnd.n577 225.874
R12796 gnd.n6253 gnd.n577 225.874
R12797 gnd.n6254 gnd.n6253 225.874
R12798 gnd.n6255 gnd.n6254 225.874
R12799 gnd.n6255 gnd.n571 225.874
R12800 gnd.n6263 gnd.n571 225.874
R12801 gnd.n6264 gnd.n6263 225.874
R12802 gnd.n6265 gnd.n6264 225.874
R12803 gnd.n6265 gnd.n565 225.874
R12804 gnd.n6273 gnd.n565 225.874
R12805 gnd.n6274 gnd.n6273 225.874
R12806 gnd.n6275 gnd.n6274 225.874
R12807 gnd.n6275 gnd.n559 225.874
R12808 gnd.n6283 gnd.n559 225.874
R12809 gnd.n6284 gnd.n6283 225.874
R12810 gnd.n6285 gnd.n6284 225.874
R12811 gnd.n6285 gnd.n553 225.874
R12812 gnd.n6293 gnd.n553 225.874
R12813 gnd.n6294 gnd.n6293 225.874
R12814 gnd.n6295 gnd.n6294 225.874
R12815 gnd.n6295 gnd.n547 225.874
R12816 gnd.n6303 gnd.n547 225.874
R12817 gnd.n6304 gnd.n6303 225.874
R12818 gnd.n6305 gnd.n6304 225.874
R12819 gnd.n6305 gnd.n541 225.874
R12820 gnd.n6313 gnd.n541 225.874
R12821 gnd.n6314 gnd.n6313 225.874
R12822 gnd.n6315 gnd.n6314 225.874
R12823 gnd.n6315 gnd.n535 225.874
R12824 gnd.n6323 gnd.n535 225.874
R12825 gnd.n6324 gnd.n6323 225.874
R12826 gnd.n6325 gnd.n6324 225.874
R12827 gnd.n6325 gnd.n529 225.874
R12828 gnd.n6333 gnd.n529 225.874
R12829 gnd.n6334 gnd.n6333 225.874
R12830 gnd.n6335 gnd.n6334 225.874
R12831 gnd.n6335 gnd.n523 225.874
R12832 gnd.n6343 gnd.n523 225.874
R12833 gnd.n6344 gnd.n6343 225.874
R12834 gnd.n6345 gnd.n6344 225.874
R12835 gnd.n6345 gnd.n517 225.874
R12836 gnd.n6353 gnd.n517 225.874
R12837 gnd.n6354 gnd.n6353 225.874
R12838 gnd.n6355 gnd.n6354 225.874
R12839 gnd.n6355 gnd.n511 225.874
R12840 gnd.n6363 gnd.n511 225.874
R12841 gnd.n6364 gnd.n6363 225.874
R12842 gnd.n6365 gnd.n6364 225.874
R12843 gnd.n6365 gnd.n505 225.874
R12844 gnd.n6373 gnd.n505 225.874
R12845 gnd.n6374 gnd.n6373 225.874
R12846 gnd.n6375 gnd.n6374 225.874
R12847 gnd.n6375 gnd.n499 225.874
R12848 gnd.n6383 gnd.n499 225.874
R12849 gnd.n6384 gnd.n6383 225.874
R12850 gnd.n6385 gnd.n6384 225.874
R12851 gnd.n6385 gnd.n493 225.874
R12852 gnd.n6393 gnd.n493 225.874
R12853 gnd.n6394 gnd.n6393 225.874
R12854 gnd.n6395 gnd.n6394 225.874
R12855 gnd.n6395 gnd.n487 225.874
R12856 gnd.n6403 gnd.n487 225.874
R12857 gnd.n6404 gnd.n6403 225.874
R12858 gnd.n6405 gnd.n6404 225.874
R12859 gnd.n6405 gnd.n481 225.874
R12860 gnd.n6413 gnd.n481 225.874
R12861 gnd.n6414 gnd.n6413 225.874
R12862 gnd.n6415 gnd.n6414 225.874
R12863 gnd.n6415 gnd.n475 225.874
R12864 gnd.n6423 gnd.n475 225.874
R12865 gnd.n6424 gnd.n6423 225.874
R12866 gnd.n6425 gnd.n6424 225.874
R12867 gnd.n6425 gnd.n469 225.874
R12868 gnd.n6433 gnd.n469 225.874
R12869 gnd.n6434 gnd.n6433 225.874
R12870 gnd.n6435 gnd.n6434 225.874
R12871 gnd.n6435 gnd.n463 225.874
R12872 gnd.n6443 gnd.n463 225.874
R12873 gnd.n6444 gnd.n6443 225.874
R12874 gnd.n6445 gnd.n6444 225.874
R12875 gnd.n6445 gnd.n457 225.874
R12876 gnd.n6453 gnd.n457 225.874
R12877 gnd.n6454 gnd.n6453 225.874
R12878 gnd.n6455 gnd.n6454 225.874
R12879 gnd.n6455 gnd.n451 225.874
R12880 gnd.n6463 gnd.n451 225.874
R12881 gnd.n6464 gnd.n6463 225.874
R12882 gnd.n6465 gnd.n6464 225.874
R12883 gnd.n6465 gnd.n445 225.874
R12884 gnd.n6473 gnd.n445 225.874
R12885 gnd.n6474 gnd.n6473 225.874
R12886 gnd.n6475 gnd.n6474 225.874
R12887 gnd.n6475 gnd.n439 225.874
R12888 gnd.n6483 gnd.n439 225.874
R12889 gnd.n6484 gnd.n6483 225.874
R12890 gnd.n6485 gnd.n6484 225.874
R12891 gnd.n6485 gnd.n433 225.874
R12892 gnd.n6493 gnd.n433 225.874
R12893 gnd.n6494 gnd.n6493 225.874
R12894 gnd.n6495 gnd.n6494 225.874
R12895 gnd.n6495 gnd.n427 225.874
R12896 gnd.n6503 gnd.n427 225.874
R12897 gnd.n6504 gnd.n6503 225.874
R12898 gnd.n6505 gnd.n6504 225.874
R12899 gnd.n6505 gnd.n421 225.874
R12900 gnd.n6513 gnd.n421 225.874
R12901 gnd.n6514 gnd.n6513 225.874
R12902 gnd.n6515 gnd.n6514 225.874
R12903 gnd.n6515 gnd.n415 225.874
R12904 gnd.n6523 gnd.n415 225.874
R12905 gnd.n6524 gnd.n6523 225.874
R12906 gnd.n6525 gnd.n6524 225.874
R12907 gnd.n6525 gnd.n409 225.874
R12908 gnd.n6533 gnd.n409 225.874
R12909 gnd.n6534 gnd.n6533 225.874
R12910 gnd.n6535 gnd.n6534 225.874
R12911 gnd.n2648 gnd.t238 224.174
R12912 gnd.n2170 gnd.t173 224.174
R12913 gnd.n6747 gnd.n83 215.659
R12914 gnd.n6543 gnd.n403 206.476
R12915 gnd.n6544 gnd.n6543 206.476
R12916 gnd.n6545 gnd.n6544 206.476
R12917 gnd.n6545 gnd.n397 206.476
R12918 gnd.n6553 gnd.n397 206.476
R12919 gnd.n6554 gnd.n6553 206.476
R12920 gnd.n6555 gnd.n6554 206.476
R12921 gnd.n6555 gnd.n391 206.476
R12922 gnd.n6563 gnd.n391 206.476
R12923 gnd.n6564 gnd.n6563 206.476
R12924 gnd.n6565 gnd.n6564 206.476
R12925 gnd.n6565 gnd.n385 206.476
R12926 gnd.n6573 gnd.n385 206.476
R12927 gnd.n6574 gnd.n6573 206.476
R12928 gnd.n6575 gnd.n6574 206.476
R12929 gnd.n6575 gnd.n379 206.476
R12930 gnd.n6583 gnd.n379 206.476
R12931 gnd.n6584 gnd.n6583 206.476
R12932 gnd.n6585 gnd.n6584 206.476
R12933 gnd.n6585 gnd.n373 206.476
R12934 gnd.n6593 gnd.n373 206.476
R12935 gnd.n6594 gnd.n6593 206.476
R12936 gnd.n6595 gnd.n6594 206.476
R12937 gnd.n6595 gnd.n367 206.476
R12938 gnd.n6603 gnd.n367 206.476
R12939 gnd.n6604 gnd.n6603 206.476
R12940 gnd.n6605 gnd.n6604 206.476
R12941 gnd.n6605 gnd.n361 206.476
R12942 gnd.n6613 gnd.n361 206.476
R12943 gnd.n6614 gnd.n6613 206.476
R12944 gnd.n6615 gnd.n6614 206.476
R12945 gnd.n6615 gnd.n355 206.476
R12946 gnd.n6623 gnd.n355 206.476
R12947 gnd.n6624 gnd.n6623 206.476
R12948 gnd.n6625 gnd.n6624 206.476
R12949 gnd.n6625 gnd.n349 206.476
R12950 gnd.n6633 gnd.n349 206.476
R12951 gnd.n6634 gnd.n6633 206.476
R12952 gnd.n6635 gnd.n6634 206.476
R12953 gnd.n6635 gnd.n343 206.476
R12954 gnd.n6643 gnd.n343 206.476
R12955 gnd.n6644 gnd.n6643 206.476
R12956 gnd.n6645 gnd.n6644 206.476
R12957 gnd.n6645 gnd.n337 206.476
R12958 gnd.n6653 gnd.n337 206.476
R12959 gnd.n6654 gnd.n6653 206.476
R12960 gnd.n6655 gnd.n6654 206.476
R12961 gnd.n6655 gnd.n331 206.476
R12962 gnd.n6663 gnd.n331 206.476
R12963 gnd.n6664 gnd.n6663 206.476
R12964 gnd.n6665 gnd.n6664 206.476
R12965 gnd.n6665 gnd.n325 206.476
R12966 gnd.n6673 gnd.n325 206.476
R12967 gnd.n6674 gnd.n6673 206.476
R12968 gnd.n6675 gnd.n6674 206.476
R12969 gnd.n6675 gnd.n319 206.476
R12970 gnd.n6683 gnd.n319 206.476
R12971 gnd.n6684 gnd.n6683 206.476
R12972 gnd.n6685 gnd.n6684 206.476
R12973 gnd.n6685 gnd.n313 206.476
R12974 gnd.n6693 gnd.n313 206.476
R12975 gnd.n6694 gnd.n6693 206.476
R12976 gnd.n6695 gnd.n6694 206.476
R12977 gnd.n6695 gnd.n307 206.476
R12978 gnd.n6703 gnd.n307 206.476
R12979 gnd.n6704 gnd.n6703 206.476
R12980 gnd.n6705 gnd.n6704 206.476
R12981 gnd.n6705 gnd.n301 206.476
R12982 gnd.n6713 gnd.n301 206.476
R12983 gnd.n6714 gnd.n6713 206.476
R12984 gnd.n6715 gnd.n6714 206.476
R12985 gnd.n6715 gnd.n295 206.476
R12986 gnd.n6723 gnd.n295 206.476
R12987 gnd.n6724 gnd.n6723 206.476
R12988 gnd.n6725 gnd.n6724 206.476
R12989 gnd.n6725 gnd.n289 206.476
R12990 gnd.n6733 gnd.n289 206.476
R12991 gnd.n6734 gnd.n6733 206.476
R12992 gnd.n6735 gnd.n6734 206.476
R12993 gnd.n6735 gnd.n283 206.476
R12994 gnd.n6745 gnd.n283 206.476
R12995 gnd.n6746 gnd.n6745 206.476
R12996 gnd.n6747 gnd.n6746 206.476
R12997 gnd.n5407 gnd.n5406 199.319
R12998 gnd.n5407 gnd.n5353 199.319
R12999 gnd.n1817 gnd.n1811 199.319
R13000 gnd.n1816 gnd.n1811 199.319
R13001 gnd.n1685 gnd.n1682 186.49
R13002 gnd.n5208 gnd.n5205 186.49
R13003 gnd.n3424 gnd.n3423 185
R13004 gnd.n3422 gnd.n3421 185
R13005 gnd.n3401 gnd.n3400 185
R13006 gnd.n3416 gnd.n3415 185
R13007 gnd.n3414 gnd.n3413 185
R13008 gnd.n3405 gnd.n3404 185
R13009 gnd.n3408 gnd.n3407 185
R13010 gnd.n3392 gnd.n3391 185
R13011 gnd.n3390 gnd.n3389 185
R13012 gnd.n3369 gnd.n3368 185
R13013 gnd.n3384 gnd.n3383 185
R13014 gnd.n3382 gnd.n3381 185
R13015 gnd.n3373 gnd.n3372 185
R13016 gnd.n3376 gnd.n3375 185
R13017 gnd.n3360 gnd.n3359 185
R13018 gnd.n3358 gnd.n3357 185
R13019 gnd.n3337 gnd.n3336 185
R13020 gnd.n3352 gnd.n3351 185
R13021 gnd.n3350 gnd.n3349 185
R13022 gnd.n3341 gnd.n3340 185
R13023 gnd.n3344 gnd.n3343 185
R13024 gnd.n3329 gnd.n3328 185
R13025 gnd.n3327 gnd.n3326 185
R13026 gnd.n3306 gnd.n3305 185
R13027 gnd.n3321 gnd.n3320 185
R13028 gnd.n3319 gnd.n3318 185
R13029 gnd.n3310 gnd.n3309 185
R13030 gnd.n3313 gnd.n3312 185
R13031 gnd.n3297 gnd.n3296 185
R13032 gnd.n3295 gnd.n3294 185
R13033 gnd.n3274 gnd.n3273 185
R13034 gnd.n3289 gnd.n3288 185
R13035 gnd.n3287 gnd.n3286 185
R13036 gnd.n3278 gnd.n3277 185
R13037 gnd.n3281 gnd.n3280 185
R13038 gnd.n3265 gnd.n3264 185
R13039 gnd.n3263 gnd.n3262 185
R13040 gnd.n3242 gnd.n3241 185
R13041 gnd.n3257 gnd.n3256 185
R13042 gnd.n3255 gnd.n3254 185
R13043 gnd.n3246 gnd.n3245 185
R13044 gnd.n3249 gnd.n3248 185
R13045 gnd.n3233 gnd.n3232 185
R13046 gnd.n3231 gnd.n3230 185
R13047 gnd.n3210 gnd.n3209 185
R13048 gnd.n3225 gnd.n3224 185
R13049 gnd.n3223 gnd.n3222 185
R13050 gnd.n3214 gnd.n3213 185
R13051 gnd.n3217 gnd.n3216 185
R13052 gnd.n3202 gnd.n3201 185
R13053 gnd.n3200 gnd.n3199 185
R13054 gnd.n3179 gnd.n3178 185
R13055 gnd.n3194 gnd.n3193 185
R13056 gnd.n3192 gnd.n3191 185
R13057 gnd.n3183 gnd.n3182 185
R13058 gnd.n3186 gnd.n3185 185
R13059 gnd.n2649 gnd.t237 178.987
R13060 gnd.n2171 gnd.t174 178.987
R13061 gnd.n1 gnd.t270 170.774
R13062 gnd.n7 gnd.t102 170.103
R13063 gnd.n6 gnd.t275 170.103
R13064 gnd.n5 gnd.t265 170.103
R13065 gnd.n4 gnd.t97 170.103
R13066 gnd.n3 gnd.t91 170.103
R13067 gnd.n2 gnd.t120 170.103
R13068 gnd.n1 gnd.t277 170.103
R13069 gnd.n5276 gnd.n5275 163.367
R13070 gnd.n5272 gnd.n5271 163.367
R13071 gnd.n5268 gnd.n5267 163.367
R13072 gnd.n5264 gnd.n5263 163.367
R13073 gnd.n5260 gnd.n5259 163.367
R13074 gnd.n5256 gnd.n5255 163.367
R13075 gnd.n5252 gnd.n5251 163.367
R13076 gnd.n5248 gnd.n5247 163.367
R13077 gnd.n5244 gnd.n5243 163.367
R13078 gnd.n5240 gnd.n5239 163.367
R13079 gnd.n5236 gnd.n5235 163.367
R13080 gnd.n5232 gnd.n5231 163.367
R13081 gnd.n5228 gnd.n5227 163.367
R13082 gnd.n5224 gnd.n5223 163.367
R13083 gnd.n5219 gnd.n5218 163.367
R13084 gnd.n5351 gnd.n1295 163.367
R13085 gnd.n5348 gnd.n5347 163.367
R13086 gnd.n5345 gnd.n1329 163.367
R13087 gnd.n5340 gnd.n5339 163.367
R13088 gnd.n5336 gnd.n5335 163.367
R13089 gnd.n5332 gnd.n5331 163.367
R13090 gnd.n5328 gnd.n5327 163.367
R13091 gnd.n5324 gnd.n5323 163.367
R13092 gnd.n5320 gnd.n5319 163.367
R13093 gnd.n5316 gnd.n5315 163.367
R13094 gnd.n5312 gnd.n5311 163.367
R13095 gnd.n5308 gnd.n5307 163.367
R13096 gnd.n5304 gnd.n5303 163.367
R13097 gnd.n5300 gnd.n5299 163.367
R13098 gnd.n5296 gnd.n5295 163.367
R13099 gnd.n5292 gnd.n5291 163.367
R13100 gnd.n5288 gnd.n5287 163.367
R13101 gnd.n1742 gnd.n1673 163.367
R13102 gnd.n1673 gnd.n1663 163.367
R13103 gnd.n4430 gnd.n1663 163.367
R13104 gnd.n4430 gnd.n1661 163.367
R13105 gnd.n4464 gnd.n1661 163.367
R13106 gnd.n4464 gnd.n1654 163.367
R13107 gnd.n4460 gnd.n1654 163.367
R13108 gnd.n4460 gnd.n4457 163.367
R13109 gnd.n4457 gnd.n4456 163.367
R13110 gnd.n4456 gnd.n1638 163.367
R13111 gnd.n1639 gnd.n1638 163.367
R13112 gnd.n1639 gnd.n1632 163.367
R13113 gnd.n4450 gnd.n1632 163.367
R13114 gnd.n4450 gnd.n4447 163.367
R13115 gnd.n4447 gnd.n4446 163.367
R13116 gnd.n4446 gnd.n1619 163.367
R13117 gnd.n4442 gnd.n1619 163.367
R13118 gnd.n4442 gnd.n1613 163.367
R13119 gnd.n4439 gnd.n1613 163.367
R13120 gnd.n4439 gnd.n1600 163.367
R13121 gnd.n4436 gnd.n1600 163.367
R13122 gnd.n4436 gnd.n1592 163.367
R13123 gnd.n4577 gnd.n1592 163.367
R13124 gnd.n4577 gnd.n1590 163.367
R13125 gnd.n4582 gnd.n1590 163.367
R13126 gnd.n4582 gnd.n1585 163.367
R13127 gnd.n1585 gnd.n1574 163.367
R13128 gnd.n4611 gnd.n1574 163.367
R13129 gnd.n4611 gnd.n1575 163.367
R13130 gnd.n1575 gnd.n1566 163.367
R13131 gnd.n4606 gnd.n1566 163.367
R13132 gnd.n4606 gnd.n1558 163.367
R13133 gnd.n4633 gnd.n1558 163.367
R13134 gnd.n4633 gnd.n1550 163.367
R13135 gnd.n4636 gnd.n1550 163.367
R13136 gnd.n4636 gnd.n1543 163.367
R13137 gnd.n4640 gnd.n1543 163.367
R13138 gnd.n4640 gnd.n1535 163.367
R13139 gnd.n4673 gnd.n1535 163.367
R13140 gnd.n4673 gnd.n1528 163.367
R13141 gnd.n4676 gnd.n1528 163.367
R13142 gnd.n4676 gnd.n1522 163.367
R13143 gnd.n4681 gnd.n1522 163.367
R13144 gnd.n4681 gnd.n1512 163.367
R13145 gnd.n1512 gnd.n1505 163.367
R13146 gnd.n4733 gnd.n1505 163.367
R13147 gnd.n4733 gnd.n1503 163.367
R13148 gnd.n4738 gnd.n1503 163.367
R13149 gnd.n4738 gnd.n1494 163.367
R13150 gnd.n1494 gnd.n1485 163.367
R13151 gnd.n4768 gnd.n1485 163.367
R13152 gnd.n4768 gnd.n1482 163.367
R13153 gnd.n4799 gnd.n1482 163.367
R13154 gnd.n4799 gnd.n1483 163.367
R13155 gnd.n4795 gnd.n1483 163.367
R13156 gnd.n4795 gnd.n4794 163.367
R13157 gnd.n4794 gnd.n1463 163.367
R13158 gnd.n1464 gnd.n1463 163.367
R13159 gnd.n1464 gnd.n1457 163.367
R13160 gnd.n4788 gnd.n1457 163.367
R13161 gnd.n4788 gnd.n1450 163.367
R13162 gnd.n4784 gnd.n1450 163.367
R13163 gnd.n4784 gnd.n1444 163.367
R13164 gnd.n4781 gnd.n1444 163.367
R13165 gnd.n4781 gnd.n1437 163.367
R13166 gnd.n4776 gnd.n1437 163.367
R13167 gnd.n4776 gnd.n1431 163.367
R13168 gnd.n4773 gnd.n1431 163.367
R13169 gnd.n4773 gnd.n1423 163.367
R13170 gnd.n1423 gnd.n1416 163.367
R13171 gnd.n4901 gnd.n1416 163.367
R13172 gnd.n4901 gnd.n1414 163.367
R13173 gnd.n4906 gnd.n1414 163.367
R13174 gnd.n4906 gnd.n1402 163.367
R13175 gnd.n1402 gnd.n1396 163.367
R13176 gnd.n4932 gnd.n1396 163.367
R13177 gnd.n4932 gnd.n1394 163.367
R13178 gnd.n4938 gnd.n1394 163.367
R13179 gnd.n4938 gnd.n1342 163.367
R13180 gnd.n1342 gnd.n1333 163.367
R13181 gnd.n5283 gnd.n1333 163.367
R13182 gnd.n4409 gnd.n1699 163.367
R13183 gnd.n4409 gnd.n1734 163.367
R13184 gnd.n4405 gnd.n4404 163.367
R13185 gnd.n4401 gnd.n4400 163.367
R13186 gnd.n4397 gnd.n4396 163.367
R13187 gnd.n4393 gnd.n4392 163.367
R13188 gnd.n4389 gnd.n4388 163.367
R13189 gnd.n4385 gnd.n4384 163.367
R13190 gnd.n4381 gnd.n4380 163.367
R13191 gnd.n4377 gnd.n4376 163.367
R13192 gnd.n4373 gnd.n4372 163.367
R13193 gnd.n4369 gnd.n4368 163.367
R13194 gnd.n4365 gnd.n4364 163.367
R13195 gnd.n4361 gnd.n4360 163.367
R13196 gnd.n4357 gnd.n4356 163.367
R13197 gnd.n4353 gnd.n4352 163.367
R13198 gnd.n4349 gnd.n4348 163.367
R13199 gnd.n1804 gnd.n1803 163.367
R13200 gnd.n1799 gnd.n1798 163.367
R13201 gnd.n1795 gnd.n1794 163.367
R13202 gnd.n1791 gnd.n1790 163.367
R13203 gnd.n1787 gnd.n1786 163.367
R13204 gnd.n1783 gnd.n1782 163.367
R13205 gnd.n1779 gnd.n1778 163.367
R13206 gnd.n1775 gnd.n1774 163.367
R13207 gnd.n1771 gnd.n1770 163.367
R13208 gnd.n1767 gnd.n1766 163.367
R13209 gnd.n1763 gnd.n1762 163.367
R13210 gnd.n1759 gnd.n1758 163.367
R13211 gnd.n1755 gnd.n1754 163.367
R13212 gnd.n1751 gnd.n1750 163.367
R13213 gnd.n1747 gnd.n1746 163.367
R13214 gnd.n4418 gnd.n1675 163.367
R13215 gnd.n4418 gnd.n1677 163.367
R13216 gnd.n1677 gnd.n1659 163.367
R13217 gnd.n4468 gnd.n1659 163.367
R13218 gnd.n4468 gnd.n1656 163.367
R13219 gnd.n4475 gnd.n1656 163.367
R13220 gnd.n4475 gnd.n1657 163.367
R13221 gnd.n4471 gnd.n1657 163.367
R13222 gnd.n4471 gnd.n1637 163.367
R13223 gnd.n4499 gnd.n1637 163.367
R13224 gnd.n4499 gnd.n1634 163.367
R13225 gnd.n4506 gnd.n1634 163.367
R13226 gnd.n4506 gnd.n1635 163.367
R13227 gnd.n4502 gnd.n1635 163.367
R13228 gnd.n4502 gnd.n1617 163.367
R13229 gnd.n4531 gnd.n1617 163.367
R13230 gnd.n4531 gnd.n1615 163.367
R13231 gnd.n4535 gnd.n1615 163.367
R13232 gnd.n4535 gnd.n1602 163.367
R13233 gnd.n4562 gnd.n1602 163.367
R13234 gnd.n4562 gnd.n1603 163.367
R13235 gnd.n4558 gnd.n1603 163.367
R13236 gnd.n4558 gnd.n1588 163.367
R13237 gnd.n4586 gnd.n1588 163.367
R13238 gnd.n4586 gnd.n1586 163.367
R13239 gnd.n4590 gnd.n1586 163.367
R13240 gnd.n4590 gnd.n1571 163.367
R13241 gnd.n4613 gnd.n1571 163.367
R13242 gnd.n4613 gnd.n1568 163.367
R13243 gnd.n4620 gnd.n1568 163.367
R13244 gnd.n4620 gnd.n1569 163.367
R13245 gnd.n4616 gnd.n1569 163.367
R13246 gnd.n4616 gnd.n1548 163.367
R13247 gnd.n4653 gnd.n1548 163.367
R13248 gnd.n4653 gnd.n1545 163.367
R13249 gnd.n4660 gnd.n1545 163.367
R13250 gnd.n4660 gnd.n1546 163.367
R13251 gnd.n4656 gnd.n1546 163.367
R13252 gnd.n4656 gnd.n1526 163.367
R13253 gnd.n4709 gnd.n1526 163.367
R13254 gnd.n4709 gnd.n1524 163.367
R13255 gnd.n4713 gnd.n1524 163.367
R13256 gnd.n4713 gnd.n1511 163.367
R13257 gnd.n4726 gnd.n1511 163.367
R13258 gnd.n4726 gnd.n1508 163.367
R13259 gnd.n4731 gnd.n1508 163.367
R13260 gnd.n4731 gnd.n1509 163.367
R13261 gnd.n1509 gnd.n1492 163.367
R13262 gnd.n4754 gnd.n1492 163.367
R13263 gnd.n4754 gnd.n1487 163.367
R13264 gnd.n4766 gnd.n1487 163.367
R13265 gnd.n4766 gnd.n1490 163.367
R13266 gnd.n1490 gnd.n1480 163.367
R13267 gnd.n4761 gnd.n1480 163.367
R13268 gnd.n4761 gnd.n4758 163.367
R13269 gnd.n4758 gnd.n1461 163.367
R13270 gnd.n4823 gnd.n1461 163.367
R13271 gnd.n4823 gnd.n1459 163.367
R13272 gnd.n4827 gnd.n1459 163.367
R13273 gnd.n4827 gnd.n1448 163.367
R13274 gnd.n4843 gnd.n1448 163.367
R13275 gnd.n4843 gnd.n1446 163.367
R13276 gnd.n4847 gnd.n1446 163.367
R13277 gnd.n4847 gnd.n1435 163.367
R13278 gnd.n4876 gnd.n1435 163.367
R13279 gnd.n4876 gnd.n1433 163.367
R13280 gnd.n4880 gnd.n1433 163.367
R13281 gnd.n4880 gnd.n1421 163.367
R13282 gnd.n4894 gnd.n1421 163.367
R13283 gnd.n4894 gnd.n1418 163.367
R13284 gnd.n4899 gnd.n1418 163.367
R13285 gnd.n4899 gnd.n1419 163.367
R13286 gnd.n1419 gnd.n1400 163.367
R13287 gnd.n4925 gnd.n1400 163.367
R13288 gnd.n4925 gnd.n1397 163.367
R13289 gnd.n4930 gnd.n1397 163.367
R13290 gnd.n4930 gnd.n1398 163.367
R13291 gnd.n1398 gnd.n1339 163.367
R13292 gnd.n5193 gnd.n1339 163.367
R13293 gnd.n5193 gnd.n1336 163.367
R13294 gnd.n5281 gnd.n1336 163.367
R13295 gnd.n5214 gnd.n5213 156.462
R13296 gnd.n3364 gnd.n3332 153.042
R13297 gnd.n3428 gnd.n3427 152.079
R13298 gnd.n3396 gnd.n3395 152.079
R13299 gnd.n3364 gnd.n3363 152.079
R13300 gnd.n1690 gnd.n1689 152
R13301 gnd.n1691 gnd.n1680 152
R13302 gnd.n1693 gnd.n1692 152
R13303 gnd.n1695 gnd.n1678 152
R13304 gnd.n1697 gnd.n1696 152
R13305 gnd.n5212 gnd.n5196 152
R13306 gnd.n5204 gnd.n5197 152
R13307 gnd.n5203 gnd.n5202 152
R13308 gnd.n5201 gnd.n5198 152
R13309 gnd.n5199 gnd.t194 150.546
R13310 gnd.t261 gnd.n3406 147.661
R13311 gnd.t252 gnd.n3374 147.661
R13312 gnd.t116 gnd.n3342 147.661
R13313 gnd.t118 gnd.n3311 147.661
R13314 gnd.t50 gnd.n3279 147.661
R13315 gnd.t56 gnd.n3247 147.661
R13316 gnd.t54 gnd.n3215 147.661
R13317 gnd.t256 gnd.n3184 147.661
R13318 gnd.n5350 gnd.n1294 143.351
R13319 gnd.n4347 gnd.n1715 143.351
R13320 gnd.n4347 gnd.n1716 143.351
R13321 gnd.n1687 gnd.t226 130.484
R13322 gnd.n1696 gnd.t135 126.766
R13323 gnd.n1694 gnd.t207 126.766
R13324 gnd.n1680 gnd.t153 126.766
R13325 gnd.n1688 gnd.t191 126.766
R13326 gnd.n5200 gnd.t229 126.766
R13327 gnd.n5202 gnd.t204 126.766
R13328 gnd.n5211 gnd.t146 126.766
R13329 gnd.n5213 gnd.t216 126.766
R13330 gnd.n5410 gnd.n5352 108.609
R13331 gnd.n4350 gnd.n4346 108.609
R13332 gnd.n3423 gnd.n3422 104.615
R13333 gnd.n3422 gnd.n3400 104.615
R13334 gnd.n3415 gnd.n3400 104.615
R13335 gnd.n3415 gnd.n3414 104.615
R13336 gnd.n3414 gnd.n3404 104.615
R13337 gnd.n3407 gnd.n3404 104.615
R13338 gnd.n3391 gnd.n3390 104.615
R13339 gnd.n3390 gnd.n3368 104.615
R13340 gnd.n3383 gnd.n3368 104.615
R13341 gnd.n3383 gnd.n3382 104.615
R13342 gnd.n3382 gnd.n3372 104.615
R13343 gnd.n3375 gnd.n3372 104.615
R13344 gnd.n3359 gnd.n3358 104.615
R13345 gnd.n3358 gnd.n3336 104.615
R13346 gnd.n3351 gnd.n3336 104.615
R13347 gnd.n3351 gnd.n3350 104.615
R13348 gnd.n3350 gnd.n3340 104.615
R13349 gnd.n3343 gnd.n3340 104.615
R13350 gnd.n3328 gnd.n3327 104.615
R13351 gnd.n3327 gnd.n3305 104.615
R13352 gnd.n3320 gnd.n3305 104.615
R13353 gnd.n3320 gnd.n3319 104.615
R13354 gnd.n3319 gnd.n3309 104.615
R13355 gnd.n3312 gnd.n3309 104.615
R13356 gnd.n3296 gnd.n3295 104.615
R13357 gnd.n3295 gnd.n3273 104.615
R13358 gnd.n3288 gnd.n3273 104.615
R13359 gnd.n3288 gnd.n3287 104.615
R13360 gnd.n3287 gnd.n3277 104.615
R13361 gnd.n3280 gnd.n3277 104.615
R13362 gnd.n3264 gnd.n3263 104.615
R13363 gnd.n3263 gnd.n3241 104.615
R13364 gnd.n3256 gnd.n3241 104.615
R13365 gnd.n3256 gnd.n3255 104.615
R13366 gnd.n3255 gnd.n3245 104.615
R13367 gnd.n3248 gnd.n3245 104.615
R13368 gnd.n3232 gnd.n3231 104.615
R13369 gnd.n3231 gnd.n3209 104.615
R13370 gnd.n3224 gnd.n3209 104.615
R13371 gnd.n3224 gnd.n3223 104.615
R13372 gnd.n3223 gnd.n3213 104.615
R13373 gnd.n3216 gnd.n3213 104.615
R13374 gnd.n3201 gnd.n3200 104.615
R13375 gnd.n3200 gnd.n3178 104.615
R13376 gnd.n3193 gnd.n3178 104.615
R13377 gnd.n3193 gnd.n3192 104.615
R13378 gnd.n3192 gnd.n3182 104.615
R13379 gnd.n3185 gnd.n3182 104.615
R13380 gnd.n2574 gnd.t134 100.632
R13381 gnd.n2144 gnd.t169 100.632
R13382 gnd.n6998 gnd.n93 99.6594
R13383 gnd.n6996 gnd.n6995 99.6594
R13384 gnd.n6991 gnd.n100 99.6594
R13385 gnd.n6989 gnd.n6988 99.6594
R13386 gnd.n6984 gnd.n107 99.6594
R13387 gnd.n6982 gnd.n6981 99.6594
R13388 gnd.n6977 gnd.n114 99.6594
R13389 gnd.n6975 gnd.n6974 99.6594
R13390 gnd.n6967 gnd.n121 99.6594
R13391 gnd.n6965 gnd.n6964 99.6594
R13392 gnd.n6960 gnd.n128 99.6594
R13393 gnd.n6958 gnd.n6957 99.6594
R13394 gnd.n6953 gnd.n135 99.6594
R13395 gnd.n6951 gnd.n6950 99.6594
R13396 gnd.n6946 gnd.n142 99.6594
R13397 gnd.n6944 gnd.n6943 99.6594
R13398 gnd.n6939 gnd.n149 99.6594
R13399 gnd.n6937 gnd.n6936 99.6594
R13400 gnd.n154 gnd.n153 99.6594
R13401 gnd.n5371 gnd.n1131 99.6594
R13402 gnd.n5375 gnd.n5374 99.6594
R13403 gnd.n5382 gnd.n5381 99.6594
R13404 gnd.n5385 gnd.n5384 99.6594
R13405 gnd.n5392 gnd.n5391 99.6594
R13406 gnd.n5395 gnd.n5394 99.6594
R13407 gnd.n5403 gnd.n5402 99.6594
R13408 gnd.n5406 gnd.n5405 99.6594
R13409 gnd.n5416 gnd.n5415 99.6594
R13410 gnd.n5419 gnd.n5418 99.6594
R13411 gnd.n5426 gnd.n5425 99.6594
R13412 gnd.n5429 gnd.n5428 99.6594
R13413 gnd.n5436 gnd.n5435 99.6594
R13414 gnd.n5439 gnd.n5438 99.6594
R13415 gnd.n5446 gnd.n5445 99.6594
R13416 gnd.n5449 gnd.n5448 99.6594
R13417 gnd.n5457 gnd.n5456 99.6594
R13418 gnd.n5460 gnd.n5459 99.6594
R13419 gnd.n1869 gnd.n1868 99.6594
R13420 gnd.n1864 gnd.n1823 99.6594
R13421 gnd.n1860 gnd.n1822 99.6594
R13422 gnd.n1856 gnd.n1821 99.6594
R13423 gnd.n1852 gnd.n1820 99.6594
R13424 gnd.n1848 gnd.n1819 99.6594
R13425 gnd.n1844 gnd.n1818 99.6594
R13426 gnd.n1816 gnd.n1815 99.6594
R13427 gnd.n4340 gnd.n4339 99.6594
R13428 gnd.n4337 gnd.n4336 99.6594
R13429 gnd.n4332 gnd.n1878 99.6594
R13430 gnd.n4330 gnd.n4329 99.6594
R13431 gnd.n4325 gnd.n1885 99.6594
R13432 gnd.n4323 gnd.n4322 99.6594
R13433 gnd.n4318 gnd.n1892 99.6594
R13434 gnd.n4316 gnd.n4315 99.6594
R13435 gnd.n4311 gnd.n1901 99.6594
R13436 gnd.n4309 gnd.n4308 99.6594
R13437 gnd.n3784 gnd.n3783 99.6594
R13438 gnd.n3778 gnd.n3556 99.6594
R13439 gnd.n3775 gnd.n3557 99.6594
R13440 gnd.n3771 gnd.n3558 99.6594
R13441 gnd.n3767 gnd.n3559 99.6594
R13442 gnd.n3763 gnd.n3560 99.6594
R13443 gnd.n3759 gnd.n3561 99.6594
R13444 gnd.n3755 gnd.n3562 99.6594
R13445 gnd.n3751 gnd.n3563 99.6594
R13446 gnd.n3746 gnd.n3564 99.6594
R13447 gnd.n3742 gnd.n3565 99.6594
R13448 gnd.n3738 gnd.n3566 99.6594
R13449 gnd.n3734 gnd.n3567 99.6594
R13450 gnd.n3730 gnd.n3568 99.6594
R13451 gnd.n3726 gnd.n3569 99.6594
R13452 gnd.n3722 gnd.n3570 99.6594
R13453 gnd.n3718 gnd.n3571 99.6594
R13454 gnd.n3714 gnd.n3572 99.6594
R13455 gnd.n3684 gnd.n3573 99.6594
R13456 gnd.n3546 gnd.n2127 99.6594
R13457 gnd.n3544 gnd.n2126 99.6594
R13458 gnd.n3540 gnd.n2125 99.6594
R13459 gnd.n3536 gnd.n2124 99.6594
R13460 gnd.n3532 gnd.n2123 99.6594
R13461 gnd.n3528 gnd.n2122 99.6594
R13462 gnd.n3524 gnd.n2121 99.6594
R13463 gnd.n3456 gnd.n2120 99.6594
R13464 gnd.n2786 gnd.n2517 99.6594
R13465 gnd.n2543 gnd.n2524 99.6594
R13466 gnd.n2545 gnd.n2525 99.6594
R13467 gnd.n2553 gnd.n2526 99.6594
R13468 gnd.n2555 gnd.n2527 99.6594
R13469 gnd.n2563 gnd.n2528 99.6594
R13470 gnd.n2565 gnd.n2529 99.6594
R13471 gnd.n2573 gnd.n2530 99.6594
R13472 gnd.n3514 gnd.n2107 99.6594
R13473 gnd.n3510 gnd.n2108 99.6594
R13474 gnd.n3506 gnd.n2109 99.6594
R13475 gnd.n3502 gnd.n2110 99.6594
R13476 gnd.n3498 gnd.n2111 99.6594
R13477 gnd.n3494 gnd.n2112 99.6594
R13478 gnd.n3490 gnd.n2113 99.6594
R13479 gnd.n3486 gnd.n2114 99.6594
R13480 gnd.n3482 gnd.n2115 99.6594
R13481 gnd.n3478 gnd.n2116 99.6594
R13482 gnd.n3474 gnd.n2117 99.6594
R13483 gnd.n3470 gnd.n2118 99.6594
R13484 gnd.n3466 gnd.n2119 99.6594
R13485 gnd.n2701 gnd.n2700 99.6594
R13486 gnd.n2695 gnd.n2612 99.6594
R13487 gnd.n2692 gnd.n2613 99.6594
R13488 gnd.n2688 gnd.n2614 99.6594
R13489 gnd.n2684 gnd.n2615 99.6594
R13490 gnd.n2680 gnd.n2616 99.6594
R13491 gnd.n2676 gnd.n2617 99.6594
R13492 gnd.n2672 gnd.n2618 99.6594
R13493 gnd.n2668 gnd.n2619 99.6594
R13494 gnd.n2664 gnd.n2620 99.6594
R13495 gnd.n2660 gnd.n2621 99.6594
R13496 gnd.n2656 gnd.n2622 99.6594
R13497 gnd.n2703 gnd.n2611 99.6594
R13498 gnd.n6847 gnd.n6846 99.6594
R13499 gnd.n6852 gnd.n6851 99.6594
R13500 gnd.n6855 gnd.n6854 99.6594
R13501 gnd.n6860 gnd.n6859 99.6594
R13502 gnd.n6863 gnd.n6862 99.6594
R13503 gnd.n6868 gnd.n6867 99.6594
R13504 gnd.n6871 gnd.n6870 99.6594
R13505 gnd.n6876 gnd.n6875 99.6594
R13506 gnd.n6879 gnd.n80 99.6594
R13507 gnd.n5031 gnd.n5030 99.6594
R13508 gnd.n5034 gnd.n5033 99.6594
R13509 gnd.n5050 gnd.n5049 99.6594
R13510 gnd.n5053 gnd.n5052 99.6594
R13511 gnd.n5069 gnd.n5068 99.6594
R13512 gnd.n5072 gnd.n5071 99.6594
R13513 gnd.n5088 gnd.n5087 99.6594
R13514 gnd.n5091 gnd.n5090 99.6594
R13515 gnd.n5109 gnd.n5108 99.6594
R13516 gnd.n4082 gnd.n4081 99.6594
R13517 gnd.n4085 gnd.n4084 99.6594
R13518 gnd.n4095 gnd.n4094 99.6594
R13519 gnd.n4104 gnd.n4103 99.6594
R13520 gnd.n4107 gnd.n4106 99.6594
R13521 gnd.n4118 gnd.n4117 99.6594
R13522 gnd.n4127 gnd.n4126 99.6594
R13523 gnd.n4130 gnd.n4129 99.6594
R13524 gnd.n4141 gnd.n4140 99.6594
R13525 gnd.n3787 gnd.n3786 99.6594
R13526 gnd.n3595 gnd.n3574 99.6594
R13527 gnd.n3599 gnd.n3575 99.6594
R13528 gnd.n3605 gnd.n3576 99.6594
R13529 gnd.n3609 gnd.n3577 99.6594
R13530 gnd.n3615 gnd.n3578 99.6594
R13531 gnd.n3619 gnd.n3579 99.6594
R13532 gnd.n3625 gnd.n3580 99.6594
R13533 gnd.n3629 gnd.n3581 99.6594
R13534 gnd.n3786 gnd.n2104 99.6594
R13535 gnd.n3598 gnd.n3574 99.6594
R13536 gnd.n3604 gnd.n3575 99.6594
R13537 gnd.n3608 gnd.n3576 99.6594
R13538 gnd.n3614 gnd.n3577 99.6594
R13539 gnd.n3618 gnd.n3578 99.6594
R13540 gnd.n3624 gnd.n3579 99.6594
R13541 gnd.n3628 gnd.n3580 99.6594
R13542 gnd.n3582 gnd.n3581 99.6594
R13543 gnd.n4140 gnd.n4139 99.6594
R13544 gnd.n4129 gnd.n4128 99.6594
R13545 gnd.n4126 gnd.n4119 99.6594
R13546 gnd.n4117 gnd.n4116 99.6594
R13547 gnd.n4106 gnd.n4105 99.6594
R13548 gnd.n4103 gnd.n4096 99.6594
R13549 gnd.n4094 gnd.n4093 99.6594
R13550 gnd.n4084 gnd.n4083 99.6594
R13551 gnd.n4081 gnd.n4080 99.6594
R13552 gnd.n5032 gnd.n5031 99.6594
R13553 gnd.n5033 gnd.n5015 99.6594
R13554 gnd.n5051 gnd.n5050 99.6594
R13555 gnd.n5052 gnd.n5006 99.6594
R13556 gnd.n5070 gnd.n5069 99.6594
R13557 gnd.n5071 gnd.n4997 99.6594
R13558 gnd.n5089 gnd.n5088 99.6594
R13559 gnd.n5090 gnd.n4988 99.6594
R13560 gnd.n5110 gnd.n5109 99.6594
R13561 gnd.n6880 gnd.n6879 99.6594
R13562 gnd.n6875 gnd.n6874 99.6594
R13563 gnd.n6870 gnd.n6869 99.6594
R13564 gnd.n6867 gnd.n6866 99.6594
R13565 gnd.n6862 gnd.n6861 99.6594
R13566 gnd.n6859 gnd.n6858 99.6594
R13567 gnd.n6854 gnd.n6853 99.6594
R13568 gnd.n6851 gnd.n6850 99.6594
R13569 gnd.n6846 gnd.n6845 99.6594
R13570 gnd.n2701 gnd.n2624 99.6594
R13571 gnd.n2693 gnd.n2612 99.6594
R13572 gnd.n2689 gnd.n2613 99.6594
R13573 gnd.n2685 gnd.n2614 99.6594
R13574 gnd.n2681 gnd.n2615 99.6594
R13575 gnd.n2677 gnd.n2616 99.6594
R13576 gnd.n2673 gnd.n2617 99.6594
R13577 gnd.n2669 gnd.n2618 99.6594
R13578 gnd.n2665 gnd.n2619 99.6594
R13579 gnd.n2661 gnd.n2620 99.6594
R13580 gnd.n2657 gnd.n2621 99.6594
R13581 gnd.n2653 gnd.n2622 99.6594
R13582 gnd.n2704 gnd.n2703 99.6594
R13583 gnd.n3469 gnd.n2119 99.6594
R13584 gnd.n3473 gnd.n2118 99.6594
R13585 gnd.n3477 gnd.n2117 99.6594
R13586 gnd.n3481 gnd.n2116 99.6594
R13587 gnd.n3485 gnd.n2115 99.6594
R13588 gnd.n3489 gnd.n2114 99.6594
R13589 gnd.n3493 gnd.n2113 99.6594
R13590 gnd.n3497 gnd.n2112 99.6594
R13591 gnd.n3501 gnd.n2111 99.6594
R13592 gnd.n3505 gnd.n2110 99.6594
R13593 gnd.n3509 gnd.n2109 99.6594
R13594 gnd.n3513 gnd.n2108 99.6594
R13595 gnd.n2148 gnd.n2107 99.6594
R13596 gnd.n2787 gnd.n2786 99.6594
R13597 gnd.n2546 gnd.n2524 99.6594
R13598 gnd.n2552 gnd.n2525 99.6594
R13599 gnd.n2556 gnd.n2526 99.6594
R13600 gnd.n2562 gnd.n2527 99.6594
R13601 gnd.n2566 gnd.n2528 99.6594
R13602 gnd.n2572 gnd.n2529 99.6594
R13603 gnd.n2530 gnd.n2514 99.6594
R13604 gnd.n3523 gnd.n2120 99.6594
R13605 gnd.n3527 gnd.n2121 99.6594
R13606 gnd.n3531 gnd.n2122 99.6594
R13607 gnd.n3535 gnd.n2123 99.6594
R13608 gnd.n3539 gnd.n2124 99.6594
R13609 gnd.n3543 gnd.n2125 99.6594
R13610 gnd.n3547 gnd.n2126 99.6594
R13611 gnd.n2129 gnd.n2127 99.6594
R13612 gnd.n3784 gnd.n3644 99.6594
R13613 gnd.n3776 gnd.n3556 99.6594
R13614 gnd.n3772 gnd.n3557 99.6594
R13615 gnd.n3768 gnd.n3558 99.6594
R13616 gnd.n3764 gnd.n3559 99.6594
R13617 gnd.n3760 gnd.n3560 99.6594
R13618 gnd.n3756 gnd.n3561 99.6594
R13619 gnd.n3752 gnd.n3562 99.6594
R13620 gnd.n3747 gnd.n3563 99.6594
R13621 gnd.n3743 gnd.n3564 99.6594
R13622 gnd.n3739 gnd.n3565 99.6594
R13623 gnd.n3735 gnd.n3566 99.6594
R13624 gnd.n3731 gnd.n3567 99.6594
R13625 gnd.n3727 gnd.n3568 99.6594
R13626 gnd.n3723 gnd.n3569 99.6594
R13627 gnd.n3719 gnd.n3570 99.6594
R13628 gnd.n3715 gnd.n3571 99.6594
R13629 gnd.n3683 gnd.n3572 99.6594
R13630 gnd.n3707 gnd.n3573 99.6594
R13631 gnd.n4310 gnd.n4309 99.6594
R13632 gnd.n1901 gnd.n1893 99.6594
R13633 gnd.n4317 gnd.n4316 99.6594
R13634 gnd.n1892 gnd.n1886 99.6594
R13635 gnd.n4324 gnd.n4323 99.6594
R13636 gnd.n1885 gnd.n1879 99.6594
R13637 gnd.n4331 gnd.n4330 99.6594
R13638 gnd.n1878 gnd.n1872 99.6594
R13639 gnd.n4338 gnd.n4337 99.6594
R13640 gnd.n4341 gnd.n4340 99.6594
R13641 gnd.n1843 gnd.n1817 99.6594
R13642 gnd.n1847 gnd.n1818 99.6594
R13643 gnd.n1851 gnd.n1819 99.6594
R13644 gnd.n1855 gnd.n1820 99.6594
R13645 gnd.n1859 gnd.n1821 99.6594
R13646 gnd.n1863 gnd.n1822 99.6594
R13647 gnd.n1825 gnd.n1823 99.6594
R13648 gnd.n1869 gnd.n1824 99.6594
R13649 gnd.n5372 gnd.n5371 99.6594
R13650 gnd.n5374 gnd.n5363 99.6594
R13651 gnd.n5383 gnd.n5382 99.6594
R13652 gnd.n5384 gnd.n5359 99.6594
R13653 gnd.n5393 gnd.n5392 99.6594
R13654 gnd.n5394 gnd.n5355 99.6594
R13655 gnd.n5404 gnd.n5403 99.6594
R13656 gnd.n5353 gnd.n1288 99.6594
R13657 gnd.n5417 gnd.n5416 99.6594
R13658 gnd.n5418 gnd.n1284 99.6594
R13659 gnd.n5427 gnd.n5426 99.6594
R13660 gnd.n5428 gnd.n1280 99.6594
R13661 gnd.n5437 gnd.n5436 99.6594
R13662 gnd.n5438 gnd.n1276 99.6594
R13663 gnd.n5447 gnd.n5446 99.6594
R13664 gnd.n5448 gnd.n1272 99.6594
R13665 gnd.n5458 gnd.n5457 99.6594
R13666 gnd.n5461 gnd.n5460 99.6594
R13667 gnd.n153 gnd.n150 99.6594
R13668 gnd.n6938 gnd.n6937 99.6594
R13669 gnd.n149 gnd.n143 99.6594
R13670 gnd.n6945 gnd.n6944 99.6594
R13671 gnd.n142 gnd.n136 99.6594
R13672 gnd.n6952 gnd.n6951 99.6594
R13673 gnd.n135 gnd.n129 99.6594
R13674 gnd.n6959 gnd.n6958 99.6594
R13675 gnd.n128 gnd.n122 99.6594
R13676 gnd.n6966 gnd.n6965 99.6594
R13677 gnd.n121 gnd.n115 99.6594
R13678 gnd.n6976 gnd.n6975 99.6594
R13679 gnd.n114 gnd.n108 99.6594
R13680 gnd.n6983 gnd.n6982 99.6594
R13681 gnd.n107 gnd.n101 99.6594
R13682 gnd.n6990 gnd.n6989 99.6594
R13683 gnd.n100 gnd.n94 99.6594
R13684 gnd.n6997 gnd.n6996 99.6594
R13685 gnd.n93 gnd.n90 99.6594
R13686 gnd.n4188 gnd.n4187 99.6594
R13687 gnd.n4088 gnd.n4057 99.6594
R13688 gnd.n4090 gnd.n4058 99.6594
R13689 gnd.n4100 gnd.n4059 99.6594
R13690 gnd.n4111 gnd.n4060 99.6594
R13691 gnd.n4113 gnd.n4061 99.6594
R13692 gnd.n4123 gnd.n4062 99.6594
R13693 gnd.n4136 gnd.n4063 99.6594
R13694 gnd.n4137 gnd.n4064 99.6594
R13695 gnd.n4065 gnd.n1912 99.6594
R13696 gnd.n4067 gnd.n4066 99.6594
R13697 gnd.n4068 gnd.n1917 99.6594
R13698 gnd.n4069 gnd.n1923 99.6594
R13699 gnd.n4071 gnd.n1925 99.6594
R13700 gnd.n4188 gnd.n4073 99.6594
R13701 gnd.n4089 gnd.n4057 99.6594
R13702 gnd.n4099 gnd.n4058 99.6594
R13703 gnd.n4110 gnd.n4059 99.6594
R13704 gnd.n4112 gnd.n4060 99.6594
R13705 gnd.n4122 gnd.n4061 99.6594
R13706 gnd.n4135 gnd.n4062 99.6594
R13707 gnd.n4138 gnd.n4063 99.6594
R13708 gnd.n4064 gnd.n1911 99.6594
R13709 gnd.n4065 gnd.n1913 99.6594
R13710 gnd.n4067 gnd.n1916 99.6594
R13711 gnd.n4068 gnd.n1918 99.6594
R13712 gnd.n4069 gnd.n1924 99.6594
R13713 gnd.n4071 gnd.n4070 99.6594
R13714 gnd.n5040 gnd.n5020 99.6594
R13715 gnd.n5044 gnd.n5042 99.6594
R13716 gnd.n5059 gnd.n5011 99.6594
R13717 gnd.n5063 gnd.n5061 99.6594
R13718 gnd.n5078 gnd.n5002 99.6594
R13719 gnd.n5082 gnd.n5080 99.6594
R13720 gnd.n5097 gnd.n4993 99.6594
R13721 gnd.n5100 gnd.n5099 99.6594
R13722 gnd.n5101 gnd.n4982 99.6594
R13723 gnd.n5120 gnd.n5119 99.6594
R13724 gnd.n5121 gnd.n4978 99.6594
R13725 gnd.n5130 gnd.n5129 99.6594
R13726 gnd.n5131 gnd.n4974 99.6594
R13727 gnd.n5143 gnd.n5142 99.6594
R13728 gnd.n5142 gnd.n5141 99.6594
R13729 gnd.n5132 gnd.n5131 99.6594
R13730 gnd.n5129 gnd.n5128 99.6594
R13731 gnd.n5122 gnd.n5121 99.6594
R13732 gnd.n5119 gnd.n5118 99.6594
R13733 gnd.n5102 gnd.n5101 99.6594
R13734 gnd.n5099 gnd.n5098 99.6594
R13735 gnd.n5081 gnd.n4993 99.6594
R13736 gnd.n5080 gnd.n5079 99.6594
R13737 gnd.n5062 gnd.n5002 99.6594
R13738 gnd.n5061 gnd.n5060 99.6594
R13739 gnd.n5043 gnd.n5011 99.6594
R13740 gnd.n5042 gnd.n5041 99.6594
R13741 gnd.n5020 gnd.n1105 99.6594
R13742 gnd.n1919 gnd.t203 98.63
R13743 gnd.n6877 gnd.t186 98.63
R13744 gnd.n4985 gnd.t180 98.63
R13745 gnd.n4131 gnd.t198 98.63
R13746 gnd.n5408 gnd.t177 98.63
R13747 gnd.n1268 gnd.t152 98.63
R13748 gnd.n156 gnd.t144 98.63
R13749 gnd.n6969 gnd.t165 98.63
R13750 gnd.n3663 gnd.t234 98.63
R13751 gnd.n3685 gnd.t225 98.63
R13752 gnd.n3584 gnd.t222 98.63
R13753 gnd.n1898 gnd.t158 98.63
R13754 gnd.n1809 gnd.t189 98.63
R13755 gnd.n5133 gnd.t183 98.63
R13756 gnd.n1738 gnd.t212 96.6984
R13757 gnd.n1330 gnd.t162 96.6984
R13758 gnd.n1735 gnd.t141 96.6906
R13759 gnd.n5215 gnd.t214 96.6906
R13760 gnd.n1687 gnd.n1686 81.8399
R13761 gnd.n2575 gnd.t133 74.8376
R13762 gnd.n2145 gnd.t170 74.8376
R13763 gnd.n1739 gnd.t211 72.8438
R13764 gnd.n1331 gnd.t163 72.8438
R13765 gnd.n1688 gnd.n1681 72.8411
R13766 gnd.n1694 gnd.n1679 72.8411
R13767 gnd.n5211 gnd.n5210 72.8411
R13768 gnd.n1920 gnd.t202 72.836
R13769 gnd.n1736 gnd.t140 72.836
R13770 gnd.n5216 gnd.t215 72.836
R13771 gnd.n6878 gnd.t187 72.836
R13772 gnd.n4986 gnd.t179 72.836
R13773 gnd.n4132 gnd.t199 72.836
R13774 gnd.n5409 gnd.t176 72.836
R13775 gnd.n1269 gnd.t151 72.836
R13776 gnd.n157 gnd.t145 72.836
R13777 gnd.n6970 gnd.t166 72.836
R13778 gnd.n3664 gnd.t233 72.836
R13779 gnd.n3686 gnd.t224 72.836
R13780 gnd.n3585 gnd.t221 72.836
R13781 gnd.n1899 gnd.t159 72.836
R13782 gnd.n1810 gnd.t190 72.836
R13783 gnd.n5134 gnd.t184 72.836
R13784 gnd.n5276 gnd.n1297 71.676
R13785 gnd.n5272 gnd.n1298 71.676
R13786 gnd.n5268 gnd.n1299 71.676
R13787 gnd.n5264 gnd.n1300 71.676
R13788 gnd.n5260 gnd.n1301 71.676
R13789 gnd.n5256 gnd.n1302 71.676
R13790 gnd.n5252 gnd.n1303 71.676
R13791 gnd.n5248 gnd.n1304 71.676
R13792 gnd.n5244 gnd.n1305 71.676
R13793 gnd.n5240 gnd.n1306 71.676
R13794 gnd.n5236 gnd.n1307 71.676
R13795 gnd.n5232 gnd.n1308 71.676
R13796 gnd.n5228 gnd.n1309 71.676
R13797 gnd.n5224 gnd.n1310 71.676
R13798 gnd.n5219 gnd.n1311 71.676
R13799 gnd.n1312 gnd.n1295 71.676
R13800 gnd.n5348 gnd.n1294 71.676
R13801 gnd.n5346 gnd.n5345 71.676
R13802 gnd.n5340 gnd.n1328 71.676
R13803 gnd.n5336 gnd.n1327 71.676
R13804 gnd.n5332 gnd.n1326 71.676
R13805 gnd.n5328 gnd.n1325 71.676
R13806 gnd.n5324 gnd.n1324 71.676
R13807 gnd.n5320 gnd.n1323 71.676
R13808 gnd.n5316 gnd.n1322 71.676
R13809 gnd.n5312 gnd.n1321 71.676
R13810 gnd.n5308 gnd.n1320 71.676
R13811 gnd.n5304 gnd.n1319 71.676
R13812 gnd.n5300 gnd.n1318 71.676
R13813 gnd.n5296 gnd.n1317 71.676
R13814 gnd.n5292 gnd.n1316 71.676
R13815 gnd.n5288 gnd.n1315 71.676
R13816 gnd.n5284 gnd.n1314 71.676
R13817 gnd.n4412 gnd.n4411 71.676
R13818 gnd.n1734 gnd.n1701 71.676
R13819 gnd.n4404 gnd.n1702 71.676
R13820 gnd.n4400 gnd.n1703 71.676
R13821 gnd.n4396 gnd.n1704 71.676
R13822 gnd.n4392 gnd.n1705 71.676
R13823 gnd.n4388 gnd.n1706 71.676
R13824 gnd.n4384 gnd.n1707 71.676
R13825 gnd.n4380 gnd.n1708 71.676
R13826 gnd.n4376 gnd.n1709 71.676
R13827 gnd.n4372 gnd.n1710 71.676
R13828 gnd.n4368 gnd.n1711 71.676
R13829 gnd.n4364 gnd.n1712 71.676
R13830 gnd.n4360 gnd.n1713 71.676
R13831 gnd.n4356 gnd.n1714 71.676
R13832 gnd.n4352 gnd.n1715 71.676
R13833 gnd.n4348 gnd.n1717 71.676
R13834 gnd.n1803 gnd.n1718 71.676
R13835 gnd.n1798 gnd.n1719 71.676
R13836 gnd.n1794 gnd.n1720 71.676
R13837 gnd.n1790 gnd.n1721 71.676
R13838 gnd.n1786 gnd.n1722 71.676
R13839 gnd.n1782 gnd.n1723 71.676
R13840 gnd.n1778 gnd.n1724 71.676
R13841 gnd.n1774 gnd.n1725 71.676
R13842 gnd.n1770 gnd.n1726 71.676
R13843 gnd.n1766 gnd.n1727 71.676
R13844 gnd.n1762 gnd.n1728 71.676
R13845 gnd.n1758 gnd.n1729 71.676
R13846 gnd.n1754 gnd.n1730 71.676
R13847 gnd.n1750 gnd.n1731 71.676
R13848 gnd.n1746 gnd.n1732 71.676
R13849 gnd.n4411 gnd.n1699 71.676
R13850 gnd.n4405 gnd.n1701 71.676
R13851 gnd.n4401 gnd.n1702 71.676
R13852 gnd.n4397 gnd.n1703 71.676
R13853 gnd.n4393 gnd.n1704 71.676
R13854 gnd.n4389 gnd.n1705 71.676
R13855 gnd.n4385 gnd.n1706 71.676
R13856 gnd.n4381 gnd.n1707 71.676
R13857 gnd.n4377 gnd.n1708 71.676
R13858 gnd.n4373 gnd.n1709 71.676
R13859 gnd.n4369 gnd.n1710 71.676
R13860 gnd.n4365 gnd.n1711 71.676
R13861 gnd.n4361 gnd.n1712 71.676
R13862 gnd.n4357 gnd.n1713 71.676
R13863 gnd.n4353 gnd.n1714 71.676
R13864 gnd.n4349 gnd.n1716 71.676
R13865 gnd.n1804 gnd.n1717 71.676
R13866 gnd.n1799 gnd.n1718 71.676
R13867 gnd.n1795 gnd.n1719 71.676
R13868 gnd.n1791 gnd.n1720 71.676
R13869 gnd.n1787 gnd.n1721 71.676
R13870 gnd.n1783 gnd.n1722 71.676
R13871 gnd.n1779 gnd.n1723 71.676
R13872 gnd.n1775 gnd.n1724 71.676
R13873 gnd.n1771 gnd.n1725 71.676
R13874 gnd.n1767 gnd.n1726 71.676
R13875 gnd.n1763 gnd.n1727 71.676
R13876 gnd.n1759 gnd.n1728 71.676
R13877 gnd.n1755 gnd.n1729 71.676
R13878 gnd.n1751 gnd.n1730 71.676
R13879 gnd.n1747 gnd.n1731 71.676
R13880 gnd.n1743 gnd.n1732 71.676
R13881 gnd.n5287 gnd.n1314 71.676
R13882 gnd.n5291 gnd.n1315 71.676
R13883 gnd.n5295 gnd.n1316 71.676
R13884 gnd.n5299 gnd.n1317 71.676
R13885 gnd.n5303 gnd.n1318 71.676
R13886 gnd.n5307 gnd.n1319 71.676
R13887 gnd.n5311 gnd.n1320 71.676
R13888 gnd.n5315 gnd.n1321 71.676
R13889 gnd.n5319 gnd.n1322 71.676
R13890 gnd.n5323 gnd.n1323 71.676
R13891 gnd.n5327 gnd.n1324 71.676
R13892 gnd.n5331 gnd.n1325 71.676
R13893 gnd.n5335 gnd.n1326 71.676
R13894 gnd.n5339 gnd.n1327 71.676
R13895 gnd.n1329 gnd.n1328 71.676
R13896 gnd.n5347 gnd.n5346 71.676
R13897 gnd.n5351 gnd.n5350 71.676
R13898 gnd.n5218 gnd.n1312 71.676
R13899 gnd.n5223 gnd.n1311 71.676
R13900 gnd.n5227 gnd.n1310 71.676
R13901 gnd.n5231 gnd.n1309 71.676
R13902 gnd.n5235 gnd.n1308 71.676
R13903 gnd.n5239 gnd.n1307 71.676
R13904 gnd.n5243 gnd.n1306 71.676
R13905 gnd.n5247 gnd.n1305 71.676
R13906 gnd.n5251 gnd.n1304 71.676
R13907 gnd.n5255 gnd.n1303 71.676
R13908 gnd.n5259 gnd.n1302 71.676
R13909 gnd.n5263 gnd.n1301 71.676
R13910 gnd.n5267 gnd.n1300 71.676
R13911 gnd.n5271 gnd.n1299 71.676
R13912 gnd.n5275 gnd.n1298 71.676
R13913 gnd.n1337 gnd.n1297 71.676
R13914 gnd.n8 gnd.t65 69.1507
R13915 gnd.n14 gnd.t42 68.4792
R13916 gnd.n13 gnd.t63 68.4792
R13917 gnd.n12 gnd.t104 68.4792
R13918 gnd.n11 gnd.t279 68.4792
R13919 gnd.n10 gnd.t113 68.4792
R13920 gnd.n9 gnd.t99 68.4792
R13921 gnd.n8 gnd.t122 68.4792
R13922 gnd.n2702 gnd.n2606 64.369
R13923 gnd.n3785 gnd.n2095 63.0944
R13924 gnd.n7006 gnd.n83 63.0944
R13925 gnd.n1801 gnd.n1739 59.5399
R13926 gnd.n5342 gnd.n1331 59.5399
R13927 gnd.n1737 gnd.n1736 59.5399
R13928 gnd.n5221 gnd.n5216 59.5399
R13929 gnd.n4414 gnd.n1697 59.1804
R13930 gnd.n3555 gnd.n2105 57.3586
R13931 gnd.n2361 gnd.t262 56.607
R13932 gnd.n40 gnd.t281 56.607
R13933 gnd.n2338 gnd.t263 56.407
R13934 gnd.n2349 gnd.t46 56.407
R13935 gnd.n17 gnd.t258 56.407
R13936 gnd.n28 gnd.t94 56.407
R13937 gnd.n2370 gnd.t71 55.8337
R13938 gnd.n2347 gnd.t61 55.8337
R13939 gnd.n2358 gnd.t95 55.8337
R13940 gnd.n49 gnd.t82 55.8337
R13941 gnd.n26 gnd.t240 55.8337
R13942 gnd.n37 gnd.t79 55.8337
R13943 gnd.n1685 gnd.n1684 54.358
R13944 gnd.n5208 gnd.n5207 54.358
R13945 gnd.n2361 gnd.n2360 53.0052
R13946 gnd.n2363 gnd.n2362 53.0052
R13947 gnd.n2365 gnd.n2364 53.0052
R13948 gnd.n2367 gnd.n2366 53.0052
R13949 gnd.n2369 gnd.n2368 53.0052
R13950 gnd.n2338 gnd.n2337 53.0052
R13951 gnd.n2340 gnd.n2339 53.0052
R13952 gnd.n2342 gnd.n2341 53.0052
R13953 gnd.n2344 gnd.n2343 53.0052
R13954 gnd.n2346 gnd.n2345 53.0052
R13955 gnd.n2349 gnd.n2348 53.0052
R13956 gnd.n2351 gnd.n2350 53.0052
R13957 gnd.n2353 gnd.n2352 53.0052
R13958 gnd.n2355 gnd.n2354 53.0052
R13959 gnd.n2357 gnd.n2356 53.0052
R13960 gnd.n48 gnd.n47 53.0052
R13961 gnd.n46 gnd.n45 53.0052
R13962 gnd.n44 gnd.n43 53.0052
R13963 gnd.n42 gnd.n41 53.0052
R13964 gnd.n40 gnd.n39 53.0052
R13965 gnd.n25 gnd.n24 53.0052
R13966 gnd.n23 gnd.n22 53.0052
R13967 gnd.n21 gnd.n20 53.0052
R13968 gnd.n19 gnd.n18 53.0052
R13969 gnd.n17 gnd.n16 53.0052
R13970 gnd.n36 gnd.n35 53.0052
R13971 gnd.n34 gnd.n33 53.0052
R13972 gnd.n32 gnd.n31 53.0052
R13973 gnd.n30 gnd.n29 53.0052
R13974 gnd.n28 gnd.n27 53.0052
R13975 gnd.n5199 gnd.n5198 52.4801
R13976 gnd.n3407 gnd.t261 52.3082
R13977 gnd.n3375 gnd.t252 52.3082
R13978 gnd.n3343 gnd.t116 52.3082
R13979 gnd.n3312 gnd.t118 52.3082
R13980 gnd.n3280 gnd.t50 52.3082
R13981 gnd.n3248 gnd.t56 52.3082
R13982 gnd.n3216 gnd.t54 52.3082
R13983 gnd.n3185 gnd.t256 52.3082
R13984 gnd.n3237 gnd.n3205 51.4173
R13985 gnd.n3301 gnd.n3300 50.455
R13986 gnd.n3269 gnd.n3268 50.455
R13987 gnd.n3237 gnd.n3236 50.455
R13988 gnd.n2649 gnd.n2648 45.1884
R13989 gnd.n2171 gnd.n2170 45.1884
R13990 gnd.n5279 gnd.n5214 44.3322
R13991 gnd.n1688 gnd.n1687 44.3189
R13992 gnd.n1921 gnd.n1920 42.2793
R13993 gnd.n2650 gnd.n2649 42.2793
R13994 gnd.n2172 gnd.n2171 42.2793
R13995 gnd.n2576 gnd.n2575 42.2793
R13996 gnd.n3522 gnd.n2145 42.2793
R13997 gnd.n6882 gnd.n6878 42.2793
R13998 gnd.n4987 gnd.n4986 42.2793
R13999 gnd.n4133 gnd.n4132 42.2793
R14000 gnd.n1270 gnd.n1269 42.2793
R14001 gnd.n6934 gnd.n157 42.2793
R14002 gnd.n6971 gnd.n6970 42.2793
R14003 gnd.n3749 gnd.n3664 42.2793
R14004 gnd.n3687 gnd.n3686 42.2793
R14005 gnd.n3586 gnd.n3585 42.2793
R14006 gnd.n1900 gnd.n1899 42.2793
R14007 gnd.n5135 gnd.n5134 42.2793
R14008 gnd.n1686 gnd.n1685 41.6274
R14009 gnd.n5209 gnd.n5208 41.6274
R14010 gnd.n6115 gnd.n6114 41.1297
R14011 gnd.n6114 gnd.n6113 41.1297
R14012 gnd.n6113 gnd.n661 41.1297
R14013 gnd.n6107 gnd.n661 41.1297
R14014 gnd.n6107 gnd.n6106 41.1297
R14015 gnd.n6106 gnd.n6105 41.1297
R14016 gnd.n6105 gnd.n668 41.1297
R14017 gnd.n6099 gnd.n668 41.1297
R14018 gnd.n6099 gnd.n6098 41.1297
R14019 gnd.n6098 gnd.n6097 41.1297
R14020 gnd.n6097 gnd.n676 41.1297
R14021 gnd.n6091 gnd.n676 41.1297
R14022 gnd.n6091 gnd.n6090 41.1297
R14023 gnd.n6090 gnd.n6089 41.1297
R14024 gnd.n6089 gnd.n684 41.1297
R14025 gnd.n6083 gnd.n684 41.1297
R14026 gnd.n6083 gnd.n6082 41.1297
R14027 gnd.n6082 gnd.n6081 41.1297
R14028 gnd.n6081 gnd.n692 41.1297
R14029 gnd.n6075 gnd.n692 41.1297
R14030 gnd.n6075 gnd.n6074 41.1297
R14031 gnd.n6074 gnd.n6073 41.1297
R14032 gnd.n6073 gnd.n700 41.1297
R14033 gnd.n6067 gnd.n700 41.1297
R14034 gnd.n6067 gnd.n6066 41.1297
R14035 gnd.n6066 gnd.n6065 41.1297
R14036 gnd.n6065 gnd.n708 41.1297
R14037 gnd.n6059 gnd.n708 41.1297
R14038 gnd.n6059 gnd.n6058 41.1297
R14039 gnd.n6058 gnd.n6057 41.1297
R14040 gnd.n6057 gnd.n716 41.1297
R14041 gnd.n6051 gnd.n716 41.1297
R14042 gnd.n6051 gnd.n6050 41.1297
R14043 gnd.n6050 gnd.n6049 41.1297
R14044 gnd.n6049 gnd.n724 41.1297
R14045 gnd.n6043 gnd.n724 41.1297
R14046 gnd.n6043 gnd.n6042 41.1297
R14047 gnd.n6042 gnd.n6041 41.1297
R14048 gnd.n6041 gnd.n732 41.1297
R14049 gnd.n6035 gnd.n732 41.1297
R14050 gnd.n6035 gnd.n6034 41.1297
R14051 gnd.n6034 gnd.n6033 41.1297
R14052 gnd.n6033 gnd.n740 41.1297
R14053 gnd.n6027 gnd.n740 41.1297
R14054 gnd.n6027 gnd.n6026 41.1297
R14055 gnd.n6026 gnd.n6025 41.1297
R14056 gnd.n6025 gnd.n748 41.1297
R14057 gnd.n6019 gnd.n748 41.1297
R14058 gnd.n6019 gnd.n6018 41.1297
R14059 gnd.n6018 gnd.n6017 41.1297
R14060 gnd.n6017 gnd.n756 41.1297
R14061 gnd.n6011 gnd.n756 41.1297
R14062 gnd.n6011 gnd.n6010 41.1297
R14063 gnd.n6010 gnd.n6009 41.1297
R14064 gnd.n6009 gnd.n764 41.1297
R14065 gnd.n6003 gnd.n764 41.1297
R14066 gnd.n6003 gnd.n6002 41.1297
R14067 gnd.n6002 gnd.n6001 41.1297
R14068 gnd.n6001 gnd.n772 41.1297
R14069 gnd.n5995 gnd.n772 41.1297
R14070 gnd.n5995 gnd.n5994 41.1297
R14071 gnd.n5994 gnd.n5993 41.1297
R14072 gnd.n5993 gnd.n780 41.1297
R14073 gnd.n5987 gnd.n780 41.1297
R14074 gnd.n5987 gnd.n5986 41.1297
R14075 gnd.n5986 gnd.n5985 41.1297
R14076 gnd.n5985 gnd.n788 41.1297
R14077 gnd.n5979 gnd.n788 41.1297
R14078 gnd.n5979 gnd.n5978 41.1297
R14079 gnd.n5978 gnd.n5977 41.1297
R14080 gnd.n5977 gnd.n796 41.1297
R14081 gnd.n5971 gnd.n796 41.1297
R14082 gnd.n5971 gnd.n5970 41.1297
R14083 gnd.n5970 gnd.n5969 41.1297
R14084 gnd.n5969 gnd.n804 41.1297
R14085 gnd.n5963 gnd.n804 41.1297
R14086 gnd.n5963 gnd.n5962 41.1297
R14087 gnd.n5962 gnd.n5961 41.1297
R14088 gnd.n5961 gnd.n812 41.1297
R14089 gnd.n5955 gnd.n812 41.1297
R14090 gnd.n5955 gnd.n5954 41.1297
R14091 gnd.n5954 gnd.n5953 41.1297
R14092 gnd.n5953 gnd.n820 41.1297
R14093 gnd.n1695 gnd.n1694 40.8975
R14094 gnd.n5212 gnd.n5211 40.8975
R14095 gnd.n5410 gnd.n5409 36.9518
R14096 gnd.n4346 gnd.n1810 36.9518
R14097 gnd.n1694 gnd.n1693 35.055
R14098 gnd.n1689 gnd.n1688 35.055
R14099 gnd.n5201 gnd.n5200 35.055
R14100 gnd.n5211 gnd.n5197 35.055
R14101 gnd.n5285 gnd.n1332 33.2493
R14102 gnd.n1744 gnd.n1741 33.2493
R14103 gnd.n2712 gnd.n2606 31.8661
R14104 gnd.n2712 gnd.n2711 31.8661
R14105 gnd.n2720 gnd.n2595 31.8661
R14106 gnd.n2728 gnd.n2595 31.8661
R14107 gnd.n2728 gnd.n2589 31.8661
R14108 gnd.n2736 gnd.n2589 31.8661
R14109 gnd.n2736 gnd.n2582 31.8661
R14110 gnd.n2774 gnd.n2582 31.8661
R14111 gnd.n2784 gnd.n2515 31.8661
R14112 gnd.n3803 gnd.n2095 31.8661
R14113 gnd.n3812 gnd.n2087 31.8661
R14114 gnd.n3812 gnd.n827 31.8661
R14115 gnd.n5946 gnd.n830 31.8661
R14116 gnd.n1970 gnd.n996 31.8661
R14117 gnd.n4056 gnd.n4055 31.8661
R14118 gnd.n4190 gnd.n4056 31.8661
R14119 gnd.n4198 gnd.n1964 31.8661
R14120 gnd.n5722 gnd.n1108 31.8661
R14121 gnd.n5716 gnd.n5715 31.8661
R14122 gnd.n5715 gnd.n5714 31.8661
R14123 gnd.n5708 gnd.n1126 31.8661
R14124 gnd.n6836 gnd.n180 31.8661
R14125 gnd.n6918 gnd.n161 31.8661
R14126 gnd.n6926 gnd.n161 31.8661
R14127 gnd.n7006 gnd.n81 31.8661
R14128 gnd.n1920 gnd.n1919 25.7944
R14129 gnd.n2575 gnd.n2574 25.7944
R14130 gnd.n2145 gnd.n2144 25.7944
R14131 gnd.n6878 gnd.n6877 25.7944
R14132 gnd.n4986 gnd.n4985 25.7944
R14133 gnd.n4132 gnd.n4131 25.7944
R14134 gnd.n5409 gnd.n5408 25.7944
R14135 gnd.n1269 gnd.n1268 25.7944
R14136 gnd.n157 gnd.n156 25.7944
R14137 gnd.n6970 gnd.n6969 25.7944
R14138 gnd.n3664 gnd.n3663 25.7944
R14139 gnd.n3686 gnd.n3685 25.7944
R14140 gnd.n3585 gnd.n3584 25.7944
R14141 gnd.n1899 gnd.n1898 25.7944
R14142 gnd.n1810 gnd.n1809 25.7944
R14143 gnd.n5134 gnd.n5133 25.7944
R14144 gnd.n2796 gnd.n2516 24.8557
R14145 gnd.n2806 gnd.n2499 24.8557
R14146 gnd.n2502 gnd.n2490 24.8557
R14147 gnd.n2827 gnd.n2491 24.8557
R14148 gnd.n2837 gnd.n2471 24.8557
R14149 gnd.n2847 gnd.n2846 24.8557
R14150 gnd.n2457 gnd.n2455 24.8557
R14151 gnd.n2878 gnd.n2877 24.8557
R14152 gnd.n2893 gnd.n2440 24.8557
R14153 gnd.n2947 gnd.n2379 24.8557
R14154 gnd.n2903 gnd.n2380 24.8557
R14155 gnd.n2940 gnd.n2391 24.8557
R14156 gnd.n2429 gnd.n2428 24.8557
R14157 gnd.n2934 gnd.n2933 24.8557
R14158 gnd.n2415 gnd.n2402 24.8557
R14159 gnd.n2973 gnd.n2972 24.8557
R14160 gnd.n2983 gnd.n2323 24.8557
R14161 gnd.n2995 gnd.n2315 24.8557
R14162 gnd.n2994 gnd.n2303 24.8557
R14163 gnd.n3013 gnd.n3012 24.8557
R14164 gnd.n3023 gnd.n2296 24.8557
R14165 gnd.n3034 gnd.n2284 24.8557
R14166 gnd.n3058 gnd.n3057 24.8557
R14167 gnd.n3069 gnd.n2267 24.8557
R14168 gnd.n3068 gnd.n2269 24.8557
R14169 gnd.n3081 gnd.n2260 24.8557
R14170 gnd.n3099 gnd.n3098 24.8557
R14171 gnd.n2251 gnd.n2240 24.8557
R14172 gnd.n3120 gnd.n2228 24.8557
R14173 gnd.n3148 gnd.n3147 24.8557
R14174 gnd.n3159 gnd.n2213 24.8557
R14175 gnd.n3170 gnd.n2206 24.8557
R14176 gnd.n3169 gnd.n2194 24.8557
R14177 gnd.n3442 gnd.n3441 24.8557
R14178 gnd.n3464 gnd.n2179 24.8557
R14179 gnd.n3079 gnd.n820 24.678
R14180 gnd.n1739 gnd.n1738 23.855
R14181 gnd.n1331 gnd.n1330 23.855
R14182 gnd.n1736 gnd.n1735 23.855
R14183 gnd.n5216 gnd.n5215 23.855
R14184 gnd.n2817 gnd.t255 23.2624
R14185 gnd.n2518 gnd.t132 22.6251
R14186 gnd.t117 gnd.n2523 21.3504
R14187 gnd.n4415 gnd.n4414 21.0737
R14188 gnd.n5280 gnd.n5279 21.0737
R14189 gnd.n3825 gnd.n843 21.0318
R14190 gnd.n5934 gnd.n852 21.0318
R14191 gnd.n3846 gnd.n3845 21.0318
R14192 gnd.n5928 gnd.n862 21.0318
R14193 gnd.n5922 gnd.n873 21.0318
R14194 gnd.n3873 gnd.n876 21.0318
R14195 gnd.n3883 gnd.n886 21.0318
R14196 gnd.n5910 gnd.n894 21.0318
R14197 gnd.n3894 gnd.n3893 21.0318
R14198 gnd.n3920 gnd.n2055 21.0318
R14199 gnd.n3928 gnd.n2049 21.0318
R14200 gnd.n3942 gnd.n2028 21.0318
R14201 gnd.n3948 gnd.n2021 21.0318
R14202 gnd.n2023 gnd.n2014 21.0318
R14203 gnd.n5902 gnd.n909 21.0318
R14204 gnd.n3969 gnd.n912 21.0318
R14205 gnd.n3977 gnd.n923 21.0318
R14206 gnd.n5890 gnd.n930 21.0318
R14207 gnd.n4023 gnd.n4022 21.0318
R14208 gnd.n5884 gnd.n940 21.0318
R14209 gnd.n5878 gnd.n951 21.0318
R14210 gnd.n3992 gnd.n954 21.0318
R14211 gnd.n3996 gnd.n964 21.0318
R14212 gnd.n5866 gnd.n972 21.0318
R14213 gnd.n4005 gnd.n975 21.0318
R14214 gnd.n5860 gnd.n983 21.0318
R14215 gnd.n5854 gnd.n993 21.0318
R14216 gnd.n5707 gnd.n1129 21.0318
R14217 gnd.n5701 gnd.n1141 21.0318
R14218 gnd.n5477 gnd.n1256 21.0318
R14219 gnd.n5544 gnd.n5543 21.0318
R14220 gnd.n5526 gnd.n1249 21.0318
R14221 gnd.n5564 gnd.n1241 21.0318
R14222 gnd.n5563 gnd.n1230 21.0318
R14223 gnd.n1233 gnd.n1220 21.0318
R14224 gnd.n5586 gnd.n1222 21.0318
R14225 gnd.n5596 gnd.n1212 21.0318
R14226 gnd.n5595 gnd.n1201 21.0318
R14227 gnd.n1205 gnd.n1194 21.0318
R14228 gnd.n5619 gnd.n1196 21.0318
R14229 gnd.n5629 gnd.n5628 21.0318
R14230 gnd.n5639 gnd.n1176 21.0318
R14231 gnd.n5638 gnd.n1180 21.0318
R14232 gnd.n5665 gnd.n1170 21.0318
R14233 gnd.n6783 gnd.n231 21.0318
R14234 gnd.n6788 gnd.n233 21.0318
R14235 gnd.n6777 gnd.n223 21.0318
R14236 gnd.n6796 gnd.n225 21.0318
R14237 gnd.n6804 gnd.n211 21.0318
R14238 gnd.n6768 gnd.n202 21.0318
R14239 gnd.n6763 gnd.n194 21.0318
R14240 gnd.n6820 gnd.n196 21.0318
R14241 gnd.n266 gnd.n186 21.0318
R14242 gnd.n6828 gnd.n188 21.0318
R14243 gnd.t13 gnd.n2241 20.7131
R14244 gnd.n5916 gnd.t69 20.7131
R14245 gnd.n3957 gnd.t83 20.7131
R14246 gnd.t88 gnd.n1184 20.7131
R14247 gnd.n6772 gnd.t67 20.7131
R14248 gnd.n1970 gnd.n1870 20.3945
R14249 gnd.n1126 gnd.n1118 20.3945
R14250 gnd.t15 gnd.n2276 20.0758
R14251 gnd.n5940 gnd.t60 20.0758
R14252 gnd.t43 gnd.n943 20.0758
R14253 gnd.t38 gnd.n5574 20.0758
R14254 gnd.n261 gnd.t78 20.0758
R14255 gnd.n1682 gnd.t193 19.8005
R14256 gnd.n1682 gnd.t228 19.8005
R14257 gnd.n1683 gnd.t209 19.8005
R14258 gnd.n1683 gnd.t155 19.8005
R14259 gnd.n5205 gnd.t148 19.8005
R14260 gnd.n5205 gnd.t218 19.8005
R14261 gnd.n5206 gnd.t231 19.8005
R14262 gnd.n5206 gnd.t206 19.8005
R14263 gnd.n1679 gnd.n1678 19.5087
R14264 gnd.n1692 gnd.n1679 19.5087
R14265 gnd.n1690 gnd.n1681 19.5087
R14266 gnd.n5210 gnd.n5204 19.5087
R14267 gnd.n2984 gnd.t19 19.4385
R14268 gnd.n5947 gnd.n5946 19.4385
R14269 gnd.n180 gnd.n168 19.4385
R14270 gnd.n4277 gnd.n4276 19.3944
R14271 gnd.n4276 gnd.n4275 19.3944
R14272 gnd.n4275 gnd.n1931 19.3944
R14273 gnd.n4271 gnd.n1931 19.3944
R14274 gnd.n4271 gnd.n4270 19.3944
R14275 gnd.n4270 gnd.n4269 19.3944
R14276 gnd.n4269 gnd.n1936 19.3944
R14277 gnd.n4265 gnd.n1936 19.3944
R14278 gnd.n4265 gnd.n4264 19.3944
R14279 gnd.n4264 gnd.n4263 19.3944
R14280 gnd.n4263 gnd.n1941 19.3944
R14281 gnd.n4259 gnd.n1941 19.3944
R14282 gnd.n4259 gnd.n4258 19.3944
R14283 gnd.n4258 gnd.n4257 19.3944
R14284 gnd.n4257 gnd.n4247 19.3944
R14285 gnd.n4253 gnd.n4247 19.3944
R14286 gnd.n4253 gnd.n4252 19.3944
R14287 gnd.n4252 gnd.n1643 19.3944
R14288 gnd.n4489 gnd.n1643 19.3944
R14289 gnd.n4489 gnd.n1641 19.3944
R14290 gnd.n4493 gnd.n1641 19.3944
R14291 gnd.n4493 gnd.n1623 19.3944
R14292 gnd.n4522 gnd.n1623 19.3944
R14293 gnd.n4522 gnd.n1621 19.3944
R14294 gnd.n4526 gnd.n1621 19.3944
R14295 gnd.n4526 gnd.n1597 19.3944
R14296 gnd.n4567 gnd.n1597 19.3944
R14297 gnd.n4567 gnd.n1594 19.3944
R14298 gnd.n4573 gnd.n1594 19.3944
R14299 gnd.n4573 gnd.n1595 19.3944
R14300 gnd.n1595 gnd.n1583 19.3944
R14301 gnd.n1583 gnd.n1581 19.3944
R14302 gnd.n4597 gnd.n1581 19.3944
R14303 gnd.n4597 gnd.n1579 19.3944
R14304 gnd.n4601 gnd.n1579 19.3944
R14305 gnd.n4601 gnd.n1553 19.3944
R14306 gnd.n4649 gnd.n1553 19.3944
R14307 gnd.n4649 gnd.n1554 19.3944
R14308 gnd.n4645 gnd.n1554 19.3944
R14309 gnd.n4645 gnd.n1530 19.3944
R14310 gnd.n4705 gnd.n1530 19.3944
R14311 gnd.n4705 gnd.n1531 19.3944
R14312 gnd.n4701 gnd.n1531 19.3944
R14313 gnd.n4701 gnd.n4700 19.3944
R14314 gnd.n4700 gnd.n4699 19.3944
R14315 gnd.n4699 gnd.n4688 19.3944
R14316 gnd.n4695 gnd.n4688 19.3944
R14317 gnd.n4695 gnd.n4694 19.3944
R14318 gnd.n4694 gnd.n4693 19.3944
R14319 gnd.n4693 gnd.n1470 19.3944
R14320 gnd.n4812 gnd.n1470 19.3944
R14321 gnd.n4812 gnd.n1467 19.3944
R14322 gnd.n4817 gnd.n1467 19.3944
R14323 gnd.n4817 gnd.n1468 19.3944
R14324 gnd.n1468 gnd.n1442 19.3944
R14325 gnd.n4851 gnd.n1442 19.3944
R14326 gnd.n4851 gnd.n1439 19.3944
R14327 gnd.n4872 gnd.n1439 19.3944
R14328 gnd.n4872 gnd.n1440 19.3944
R14329 gnd.n4868 gnd.n1440 19.3944
R14330 gnd.n4868 gnd.n4867 19.3944
R14331 gnd.n4867 gnd.n4866 19.3944
R14332 gnd.n4866 gnd.n4861 19.3944
R14333 gnd.n4862 gnd.n4861 19.3944
R14334 gnd.n4862 gnd.n1391 19.3944
R14335 gnd.n4942 gnd.n1391 19.3944
R14336 gnd.n4942 gnd.n1389 19.3944
R14337 gnd.n4947 gnd.n1389 19.3944
R14338 gnd.n4947 gnd.n1387 19.3944
R14339 gnd.n4952 gnd.n1387 19.3944
R14340 gnd.n4953 gnd.n4952 19.3944
R14341 gnd.n4953 gnd.n1385 19.3944
R14342 gnd.n4957 gnd.n1385 19.3944
R14343 gnd.n4960 gnd.n4957 19.3944
R14344 gnd.n4961 gnd.n4960 19.3944
R14345 gnd.n4961 gnd.n1383 19.3944
R14346 gnd.n4965 gnd.n1383 19.3944
R14347 gnd.n4968 gnd.n4965 19.3944
R14348 gnd.n4969 gnd.n4968 19.3944
R14349 gnd.n4969 gnd.n1380 19.3944
R14350 gnd.n5149 gnd.n1380 19.3944
R14351 gnd.n5149 gnd.n1381 19.3944
R14352 gnd.n4283 gnd.n4282 19.3944
R14353 gnd.n4282 gnd.n4281 19.3944
R14354 gnd.n4281 gnd.n1926 19.3944
R14355 gnd.n4186 gnd.n4185 19.3944
R14356 gnd.n4185 gnd.n4075 19.3944
R14357 gnd.n4178 gnd.n4075 19.3944
R14358 gnd.n4178 gnd.n4177 19.3944
R14359 gnd.n4177 gnd.n4091 19.3944
R14360 gnd.n4170 gnd.n4091 19.3944
R14361 gnd.n4170 gnd.n4169 19.3944
R14362 gnd.n4169 gnd.n4101 19.3944
R14363 gnd.n4162 gnd.n4101 19.3944
R14364 gnd.n4162 gnd.n4161 19.3944
R14365 gnd.n4161 gnd.n4114 19.3944
R14366 gnd.n4154 gnd.n4114 19.3944
R14367 gnd.n4154 gnd.n4153 19.3944
R14368 gnd.n4153 gnd.n4124 19.3944
R14369 gnd.n4146 gnd.n4124 19.3944
R14370 gnd.n4146 gnd.n4145 19.3944
R14371 gnd.n4145 gnd.n1910 19.3944
R14372 gnd.n4294 gnd.n1910 19.3944
R14373 gnd.n4294 gnd.n4293 19.3944
R14374 gnd.n4293 gnd.n4292 19.3944
R14375 gnd.n4292 gnd.n1914 19.3944
R14376 gnd.n4288 gnd.n1914 19.3944
R14377 gnd.n4288 gnd.n4287 19.3944
R14378 gnd.n4287 gnd.n4286 19.3944
R14379 gnd.n2699 gnd.n2698 19.3944
R14380 gnd.n2698 gnd.n2697 19.3944
R14381 gnd.n2697 gnd.n2696 19.3944
R14382 gnd.n2696 gnd.n2694 19.3944
R14383 gnd.n2694 gnd.n2691 19.3944
R14384 gnd.n2691 gnd.n2690 19.3944
R14385 gnd.n2690 gnd.n2687 19.3944
R14386 gnd.n2687 gnd.n2686 19.3944
R14387 gnd.n2686 gnd.n2683 19.3944
R14388 gnd.n2683 gnd.n2682 19.3944
R14389 gnd.n2682 gnd.n2679 19.3944
R14390 gnd.n2679 gnd.n2678 19.3944
R14391 gnd.n2678 gnd.n2675 19.3944
R14392 gnd.n2675 gnd.n2674 19.3944
R14393 gnd.n2674 gnd.n2671 19.3944
R14394 gnd.n2671 gnd.n2670 19.3944
R14395 gnd.n2670 gnd.n2667 19.3944
R14396 gnd.n2667 gnd.n2666 19.3944
R14397 gnd.n2666 gnd.n2663 19.3944
R14398 gnd.n2663 gnd.n2662 19.3944
R14399 gnd.n2662 gnd.n2659 19.3944
R14400 gnd.n2659 gnd.n2658 19.3944
R14401 gnd.n2655 gnd.n2654 19.3944
R14402 gnd.n2654 gnd.n2610 19.3944
R14403 gnd.n2705 gnd.n2610 19.3944
R14404 gnd.n3472 gnd.n3471 19.3944
R14405 gnd.n3471 gnd.n3468 19.3944
R14406 gnd.n3468 gnd.n3467 19.3944
R14407 gnd.n3517 gnd.n3516 19.3944
R14408 gnd.n3516 gnd.n3515 19.3944
R14409 gnd.n3515 gnd.n3512 19.3944
R14410 gnd.n3512 gnd.n3511 19.3944
R14411 gnd.n3511 gnd.n3508 19.3944
R14412 gnd.n3508 gnd.n3507 19.3944
R14413 gnd.n3507 gnd.n3504 19.3944
R14414 gnd.n3504 gnd.n3503 19.3944
R14415 gnd.n3503 gnd.n3500 19.3944
R14416 gnd.n3500 gnd.n3499 19.3944
R14417 gnd.n3499 gnd.n3496 19.3944
R14418 gnd.n3496 gnd.n3495 19.3944
R14419 gnd.n3495 gnd.n3492 19.3944
R14420 gnd.n3492 gnd.n3491 19.3944
R14421 gnd.n3491 gnd.n3488 19.3944
R14422 gnd.n3488 gnd.n3487 19.3944
R14423 gnd.n3487 gnd.n3484 19.3944
R14424 gnd.n3484 gnd.n3483 19.3944
R14425 gnd.n3483 gnd.n3480 19.3944
R14426 gnd.n3480 gnd.n3479 19.3944
R14427 gnd.n3479 gnd.n3476 19.3944
R14428 gnd.n3476 gnd.n3475 19.3944
R14429 gnd.n2798 gnd.n2507 19.3944
R14430 gnd.n2808 gnd.n2507 19.3944
R14431 gnd.n2809 gnd.n2808 19.3944
R14432 gnd.n2809 gnd.n2488 19.3944
R14433 gnd.n2829 gnd.n2488 19.3944
R14434 gnd.n2829 gnd.n2480 19.3944
R14435 gnd.n2839 gnd.n2480 19.3944
R14436 gnd.n2840 gnd.n2839 19.3944
R14437 gnd.n2841 gnd.n2840 19.3944
R14438 gnd.n2841 gnd.n2463 19.3944
R14439 gnd.n2858 gnd.n2463 19.3944
R14440 gnd.n2861 gnd.n2858 19.3944
R14441 gnd.n2861 gnd.n2860 19.3944
R14442 gnd.n2860 gnd.n2436 19.3944
R14443 gnd.n2900 gnd.n2436 19.3944
R14444 gnd.n2900 gnd.n2433 19.3944
R14445 gnd.n2906 gnd.n2433 19.3944
R14446 gnd.n2907 gnd.n2906 19.3944
R14447 gnd.n2907 gnd.n2431 19.3944
R14448 gnd.n2913 gnd.n2431 19.3944
R14449 gnd.n2916 gnd.n2913 19.3944
R14450 gnd.n2918 gnd.n2916 19.3944
R14451 gnd.n2924 gnd.n2918 19.3944
R14452 gnd.n2924 gnd.n2923 19.3944
R14453 gnd.n2923 gnd.n2318 19.3944
R14454 gnd.n2990 gnd.n2318 19.3944
R14455 gnd.n2991 gnd.n2990 19.3944
R14456 gnd.n2991 gnd.n2311 19.3944
R14457 gnd.n3002 gnd.n2311 19.3944
R14458 gnd.n3003 gnd.n3002 19.3944
R14459 gnd.n3003 gnd.n2294 19.3944
R14460 gnd.n2294 gnd.n2292 19.3944
R14461 gnd.n3027 gnd.n2292 19.3944
R14462 gnd.n3028 gnd.n3027 19.3944
R14463 gnd.n3028 gnd.n2263 19.3944
R14464 gnd.n3075 gnd.n2263 19.3944
R14465 gnd.n3076 gnd.n3075 19.3944
R14466 gnd.n3076 gnd.n2256 19.3944
R14467 gnd.n3088 gnd.n2256 19.3944
R14468 gnd.n3089 gnd.n3088 19.3944
R14469 gnd.n3089 gnd.n2239 19.3944
R14470 gnd.n2239 gnd.n2237 19.3944
R14471 gnd.n3113 gnd.n2237 19.3944
R14472 gnd.n3114 gnd.n3113 19.3944
R14473 gnd.n3114 gnd.n2209 19.3944
R14474 gnd.n3165 gnd.n2209 19.3944
R14475 gnd.n3166 gnd.n3165 19.3944
R14476 gnd.n3166 gnd.n2202 19.3944
R14477 gnd.n3433 gnd.n2202 19.3944
R14478 gnd.n3434 gnd.n3433 19.3944
R14479 gnd.n3434 gnd.n2183 19.3944
R14480 gnd.n3459 gnd.n2183 19.3944
R14481 gnd.n3459 gnd.n2184 19.3944
R14482 gnd.n2789 gnd.n2788 19.3944
R14483 gnd.n2788 gnd.n2521 19.3944
R14484 gnd.n2544 gnd.n2521 19.3944
R14485 gnd.n2547 gnd.n2544 19.3944
R14486 gnd.n2547 gnd.n2540 19.3944
R14487 gnd.n2551 gnd.n2540 19.3944
R14488 gnd.n2554 gnd.n2551 19.3944
R14489 gnd.n2557 gnd.n2554 19.3944
R14490 gnd.n2557 gnd.n2538 19.3944
R14491 gnd.n2561 gnd.n2538 19.3944
R14492 gnd.n2564 gnd.n2561 19.3944
R14493 gnd.n2567 gnd.n2564 19.3944
R14494 gnd.n2567 gnd.n2536 19.3944
R14495 gnd.n2571 gnd.n2536 19.3944
R14496 gnd.n2794 gnd.n2793 19.3944
R14497 gnd.n2793 gnd.n2497 19.3944
R14498 gnd.n2819 gnd.n2497 19.3944
R14499 gnd.n2819 gnd.n2495 19.3944
R14500 gnd.n2825 gnd.n2495 19.3944
R14501 gnd.n2825 gnd.n2824 19.3944
R14502 gnd.n2824 gnd.n2469 19.3944
R14503 gnd.n2849 gnd.n2469 19.3944
R14504 gnd.n2849 gnd.n2467 19.3944
R14505 gnd.n2853 gnd.n2467 19.3944
R14506 gnd.n2853 gnd.n2447 19.3944
R14507 gnd.n2880 gnd.n2447 19.3944
R14508 gnd.n2880 gnd.n2445 19.3944
R14509 gnd.n2890 gnd.n2445 19.3944
R14510 gnd.n2890 gnd.n2889 19.3944
R14511 gnd.n2889 gnd.n2888 19.3944
R14512 gnd.n2888 gnd.n2394 19.3944
R14513 gnd.n2938 gnd.n2394 19.3944
R14514 gnd.n2938 gnd.n2937 19.3944
R14515 gnd.n2937 gnd.n2936 19.3944
R14516 gnd.n2936 gnd.n2398 19.3944
R14517 gnd.n2418 gnd.n2398 19.3944
R14518 gnd.n2418 gnd.n2328 19.3944
R14519 gnd.n2975 gnd.n2328 19.3944
R14520 gnd.n2975 gnd.n2326 19.3944
R14521 gnd.n2981 gnd.n2326 19.3944
R14522 gnd.n2981 gnd.n2980 19.3944
R14523 gnd.n2980 gnd.n2301 19.3944
R14524 gnd.n3015 gnd.n2301 19.3944
R14525 gnd.n3015 gnd.n2299 19.3944
R14526 gnd.n3021 gnd.n2299 19.3944
R14527 gnd.n3021 gnd.n3020 19.3944
R14528 gnd.n3020 gnd.n2274 19.3944
R14529 gnd.n3060 gnd.n2274 19.3944
R14530 gnd.n3060 gnd.n2272 19.3944
R14531 gnd.n3066 gnd.n2272 19.3944
R14532 gnd.n3066 gnd.n3065 19.3944
R14533 gnd.n3065 gnd.n2246 19.3944
R14534 gnd.n3101 gnd.n2246 19.3944
R14535 gnd.n3101 gnd.n2244 19.3944
R14536 gnd.n3107 gnd.n2244 19.3944
R14537 gnd.n3107 gnd.n3106 19.3944
R14538 gnd.n3106 gnd.n2219 19.3944
R14539 gnd.n3150 gnd.n2219 19.3944
R14540 gnd.n3150 gnd.n2217 19.3944
R14541 gnd.n3156 gnd.n2217 19.3944
R14542 gnd.n3156 gnd.n3155 19.3944
R14543 gnd.n3155 gnd.n2192 19.3944
R14544 gnd.n3444 gnd.n2192 19.3944
R14545 gnd.n3444 gnd.n2190 19.3944
R14546 gnd.n3452 gnd.n2190 19.3944
R14547 gnd.n3452 gnd.n3451 19.3944
R14548 gnd.n3451 gnd.n3450 19.3944
R14549 gnd.n3553 gnd.n3552 19.3944
R14550 gnd.n3552 gnd.n2131 19.3944
R14551 gnd.n3548 gnd.n2131 19.3944
R14552 gnd.n3548 gnd.n3545 19.3944
R14553 gnd.n3545 gnd.n3542 19.3944
R14554 gnd.n3542 gnd.n3541 19.3944
R14555 gnd.n3541 gnd.n3538 19.3944
R14556 gnd.n3538 gnd.n3537 19.3944
R14557 gnd.n3537 gnd.n3534 19.3944
R14558 gnd.n3534 gnd.n3533 19.3944
R14559 gnd.n3533 gnd.n3530 19.3944
R14560 gnd.n3530 gnd.n3529 19.3944
R14561 gnd.n3529 gnd.n3526 19.3944
R14562 gnd.n3526 gnd.n3525 19.3944
R14563 gnd.n2709 gnd.n2608 19.3944
R14564 gnd.n2709 gnd.n2599 19.3944
R14565 gnd.n2722 gnd.n2599 19.3944
R14566 gnd.n2722 gnd.n2597 19.3944
R14567 gnd.n2726 gnd.n2597 19.3944
R14568 gnd.n2726 gnd.n2587 19.3944
R14569 gnd.n2738 gnd.n2587 19.3944
R14570 gnd.n2738 gnd.n2585 19.3944
R14571 gnd.n2772 gnd.n2585 19.3944
R14572 gnd.n2772 gnd.n2771 19.3944
R14573 gnd.n2771 gnd.n2770 19.3944
R14574 gnd.n2770 gnd.n2769 19.3944
R14575 gnd.n2769 gnd.n2766 19.3944
R14576 gnd.n2766 gnd.n2765 19.3944
R14577 gnd.n2765 gnd.n2764 19.3944
R14578 gnd.n2764 gnd.n2762 19.3944
R14579 gnd.n2762 gnd.n2761 19.3944
R14580 gnd.n2761 gnd.n2758 19.3944
R14581 gnd.n2758 gnd.n2757 19.3944
R14582 gnd.n2757 gnd.n2756 19.3944
R14583 gnd.n2756 gnd.n2754 19.3944
R14584 gnd.n2754 gnd.n2453 19.3944
R14585 gnd.n2869 gnd.n2453 19.3944
R14586 gnd.n2869 gnd.n2451 19.3944
R14587 gnd.n2875 gnd.n2451 19.3944
R14588 gnd.n2875 gnd.n2874 19.3944
R14589 gnd.n2874 gnd.n2375 19.3944
R14590 gnd.n2949 gnd.n2375 19.3944
R14591 gnd.n2949 gnd.n2376 19.3944
R14592 gnd.n2423 gnd.n2422 19.3944
R14593 gnd.n2426 gnd.n2425 19.3944
R14594 gnd.n2413 gnd.n2412 19.3944
R14595 gnd.n2968 gnd.n2333 19.3944
R14596 gnd.n2968 gnd.n2967 19.3944
R14597 gnd.n2967 gnd.n2966 19.3944
R14598 gnd.n2966 gnd.n2964 19.3944
R14599 gnd.n2964 gnd.n2963 19.3944
R14600 gnd.n2963 gnd.n2961 19.3944
R14601 gnd.n2961 gnd.n2960 19.3944
R14602 gnd.n2960 gnd.n2282 19.3944
R14603 gnd.n3036 gnd.n2282 19.3944
R14604 gnd.n3036 gnd.n2280 19.3944
R14605 gnd.n3055 gnd.n2280 19.3944
R14606 gnd.n3055 gnd.n3054 19.3944
R14607 gnd.n3054 gnd.n3053 19.3944
R14608 gnd.n3053 gnd.n3051 19.3944
R14609 gnd.n3051 gnd.n3050 19.3944
R14610 gnd.n3050 gnd.n3048 19.3944
R14611 gnd.n3048 gnd.n3047 19.3944
R14612 gnd.n3047 gnd.n2226 19.3944
R14613 gnd.n3122 gnd.n2226 19.3944
R14614 gnd.n3122 gnd.n2224 19.3944
R14615 gnd.n3145 gnd.n2224 19.3944
R14616 gnd.n3145 gnd.n3144 19.3944
R14617 gnd.n3144 gnd.n3143 19.3944
R14618 gnd.n3143 gnd.n3140 19.3944
R14619 gnd.n3140 gnd.n3139 19.3944
R14620 gnd.n3139 gnd.n3137 19.3944
R14621 gnd.n3137 gnd.n3136 19.3944
R14622 gnd.n3136 gnd.n3134 19.3944
R14623 gnd.n3134 gnd.n2178 19.3944
R14624 gnd.n2714 gnd.n2604 19.3944
R14625 gnd.n2714 gnd.n2602 19.3944
R14626 gnd.n2718 gnd.n2602 19.3944
R14627 gnd.n2718 gnd.n2593 19.3944
R14628 gnd.n2730 gnd.n2593 19.3944
R14629 gnd.n2730 gnd.n2591 19.3944
R14630 gnd.n2734 gnd.n2591 19.3944
R14631 gnd.n2734 gnd.n2580 19.3944
R14632 gnd.n2776 gnd.n2580 19.3944
R14633 gnd.n2776 gnd.n2534 19.3944
R14634 gnd.n2782 gnd.n2534 19.3944
R14635 gnd.n2782 gnd.n2781 19.3944
R14636 gnd.n2781 gnd.n2512 19.3944
R14637 gnd.n2803 gnd.n2512 19.3944
R14638 gnd.n2803 gnd.n2505 19.3944
R14639 gnd.n2814 gnd.n2505 19.3944
R14640 gnd.n2814 gnd.n2813 19.3944
R14641 gnd.n2813 gnd.n2486 19.3944
R14642 gnd.n2834 gnd.n2486 19.3944
R14643 gnd.n2834 gnd.n2476 19.3944
R14644 gnd.n2844 gnd.n2476 19.3944
R14645 gnd.n2844 gnd.n2459 19.3944
R14646 gnd.n2865 gnd.n2459 19.3944
R14647 gnd.n2865 gnd.n2864 19.3944
R14648 gnd.n2864 gnd.n2438 19.3944
R14649 gnd.n2895 gnd.n2438 19.3944
R14650 gnd.n2895 gnd.n2383 19.3944
R14651 gnd.n2945 gnd.n2383 19.3944
R14652 gnd.n2945 gnd.n2944 19.3944
R14653 gnd.n2944 gnd.n2943 19.3944
R14654 gnd.n2943 gnd.n2387 19.3944
R14655 gnd.n2405 gnd.n2387 19.3944
R14656 gnd.n2931 gnd.n2405 19.3944
R14657 gnd.n2931 gnd.n2930 19.3944
R14658 gnd.n2930 gnd.n2929 19.3944
R14659 gnd.n2929 gnd.n2409 19.3944
R14660 gnd.n2409 gnd.n2320 19.3944
R14661 gnd.n2986 gnd.n2320 19.3944
R14662 gnd.n2986 gnd.n2313 19.3944
R14663 gnd.n2997 gnd.n2313 19.3944
R14664 gnd.n2997 gnd.n2309 19.3944
R14665 gnd.n3010 gnd.n2309 19.3944
R14666 gnd.n3010 gnd.n3009 19.3944
R14667 gnd.n3009 gnd.n2288 19.3944
R14668 gnd.n3032 gnd.n2288 19.3944
R14669 gnd.n3032 gnd.n3031 19.3944
R14670 gnd.n3031 gnd.n2265 19.3944
R14671 gnd.n3071 gnd.n2265 19.3944
R14672 gnd.n3071 gnd.n2258 19.3944
R14673 gnd.n3083 gnd.n2258 19.3944
R14674 gnd.n3083 gnd.n2254 19.3944
R14675 gnd.n3096 gnd.n2254 19.3944
R14676 gnd.n3096 gnd.n3095 19.3944
R14677 gnd.n3095 gnd.n2233 19.3944
R14678 gnd.n3118 gnd.n2233 19.3944
R14679 gnd.n3118 gnd.n3117 19.3944
R14680 gnd.n3117 gnd.n2211 19.3944
R14681 gnd.n3161 gnd.n2211 19.3944
R14682 gnd.n3161 gnd.n2204 19.3944
R14683 gnd.n3172 gnd.n2204 19.3944
R14684 gnd.n3172 gnd.n2200 19.3944
R14685 gnd.n3439 gnd.n2200 19.3944
R14686 gnd.n3439 gnd.n3438 19.3944
R14687 gnd.n3438 gnd.n2181 19.3944
R14688 gnd.n3462 gnd.n2181 19.3944
R14689 gnd.n5470 gnd.n1265 19.3944
R14690 gnd.n5470 gnd.n1262 19.3944
R14691 gnd.n5475 gnd.n1262 19.3944
R14692 gnd.n5475 gnd.n1263 19.3944
R14693 gnd.n1263 gnd.n1247 19.3944
R14694 gnd.n5556 gnd.n1247 19.3944
R14695 gnd.n5556 gnd.n1244 19.3944
R14696 gnd.n5561 gnd.n1244 19.3944
R14697 gnd.n5561 gnd.n1245 19.3944
R14698 gnd.n1245 gnd.n1218 19.3944
R14699 gnd.n5588 gnd.n1218 19.3944
R14700 gnd.n5588 gnd.n1215 19.3944
R14701 gnd.n5593 gnd.n1215 19.3944
R14702 gnd.n5593 gnd.n1216 19.3944
R14703 gnd.n1216 gnd.n1192 19.3944
R14704 gnd.n5621 gnd.n1192 19.3944
R14705 gnd.n5621 gnd.n1188 19.3944
R14706 gnd.n5626 gnd.n1188 19.3944
R14707 gnd.n5626 gnd.n1190 19.3944
R14708 gnd.n1190 gnd.n1189 19.3944
R14709 gnd.n1189 gnd.n52 19.3944
R14710 gnd.n7038 gnd.n52 19.3944
R14711 gnd.n7038 gnd.n7037 19.3944
R14712 gnd.n7037 gnd.n7036 19.3944
R14713 gnd.n7036 gnd.n57 19.3944
R14714 gnd.n7032 gnd.n57 19.3944
R14715 gnd.n7032 gnd.n7031 19.3944
R14716 gnd.n7031 gnd.n7030 19.3944
R14717 gnd.n7030 gnd.n62 19.3944
R14718 gnd.n7026 gnd.n62 19.3944
R14719 gnd.n7026 gnd.n7025 19.3944
R14720 gnd.n7025 gnd.n7024 19.3944
R14721 gnd.n7024 gnd.n67 19.3944
R14722 gnd.n7020 gnd.n67 19.3944
R14723 gnd.n7020 gnd.n7019 19.3944
R14724 gnd.n7019 gnd.n7018 19.3944
R14725 gnd.n7018 gnd.n72 19.3944
R14726 gnd.n7014 gnd.n72 19.3944
R14727 gnd.n7014 gnd.n7013 19.3944
R14728 gnd.n7013 gnd.n7012 19.3944
R14729 gnd.n7012 gnd.n77 19.3944
R14730 gnd.n7008 gnd.n77 19.3944
R14731 gnd.n6907 gnd.n6906 19.3944
R14732 gnd.n6906 gnd.n6905 19.3944
R14733 gnd.n6905 gnd.n6848 19.3944
R14734 gnd.n6901 gnd.n6848 19.3944
R14735 gnd.n6901 gnd.n6900 19.3944
R14736 gnd.n6900 gnd.n6899 19.3944
R14737 gnd.n6899 gnd.n6856 19.3944
R14738 gnd.n6895 gnd.n6856 19.3944
R14739 gnd.n6895 gnd.n6894 19.3944
R14740 gnd.n6894 gnd.n6893 19.3944
R14741 gnd.n6893 gnd.n6864 19.3944
R14742 gnd.n6889 gnd.n6864 19.3944
R14743 gnd.n6889 gnd.n6888 19.3944
R14744 gnd.n6888 gnd.n6887 19.3944
R14745 gnd.n6887 gnd.n6872 19.3944
R14746 gnd.n6883 gnd.n6872 19.3944
R14747 gnd.n5029 gnd.n5023 19.3944
R14748 gnd.n5035 gnd.n5023 19.3944
R14749 gnd.n5035 gnd.n5016 19.3944
R14750 gnd.n5048 gnd.n5016 19.3944
R14751 gnd.n5048 gnd.n5014 19.3944
R14752 gnd.n5054 gnd.n5014 19.3944
R14753 gnd.n5054 gnd.n5007 19.3944
R14754 gnd.n5067 gnd.n5007 19.3944
R14755 gnd.n5067 gnd.n5005 19.3944
R14756 gnd.n5073 gnd.n5005 19.3944
R14757 gnd.n5073 gnd.n4998 19.3944
R14758 gnd.n5086 gnd.n4998 19.3944
R14759 gnd.n5086 gnd.n4996 19.3944
R14760 gnd.n5092 gnd.n4996 19.3944
R14761 gnd.n5092 gnd.n4989 19.3944
R14762 gnd.n5107 gnd.n4989 19.3944
R14763 gnd.n5026 gnd.n1144 19.3944
R14764 gnd.n5699 gnd.n1144 19.3944
R14765 gnd.n5699 gnd.n1145 19.3944
R14766 gnd.n5695 gnd.n1145 19.3944
R14767 gnd.n5695 gnd.n5694 19.3944
R14768 gnd.n5694 gnd.n5693 19.3944
R14769 gnd.n5693 gnd.n1151 19.3944
R14770 gnd.n5689 gnd.n1151 19.3944
R14771 gnd.n5689 gnd.n5688 19.3944
R14772 gnd.n5688 gnd.n5687 19.3944
R14773 gnd.n5687 gnd.n1156 19.3944
R14774 gnd.n5683 gnd.n1156 19.3944
R14775 gnd.n5683 gnd.n5682 19.3944
R14776 gnd.n5682 gnd.n5681 19.3944
R14777 gnd.n5681 gnd.n1161 19.3944
R14778 gnd.n5677 gnd.n1161 19.3944
R14779 gnd.n5677 gnd.n5676 19.3944
R14780 gnd.n5676 gnd.n5675 19.3944
R14781 gnd.n5675 gnd.n1166 19.3944
R14782 gnd.n5671 gnd.n1166 19.3944
R14783 gnd.n5671 gnd.n5670 19.3944
R14784 gnd.n5670 gnd.n5669 19.3944
R14785 gnd.n5669 gnd.n229 19.3944
R14786 gnd.n6790 gnd.n229 19.3944
R14787 gnd.n6790 gnd.n227 19.3944
R14788 gnd.n6794 gnd.n227 19.3944
R14789 gnd.n6794 gnd.n207 19.3944
R14790 gnd.n6806 gnd.n207 19.3944
R14791 gnd.n6806 gnd.n205 19.3944
R14792 gnd.n6810 gnd.n205 19.3944
R14793 gnd.n6810 gnd.n192 19.3944
R14794 gnd.n6822 gnd.n192 19.3944
R14795 gnd.n6822 gnd.n190 19.3944
R14796 gnd.n6826 gnd.n190 19.3944
R14797 gnd.n6826 gnd.n175 19.3944
R14798 gnd.n6838 gnd.n175 19.3944
R14799 gnd.n6838 gnd.n172 19.3944
R14800 gnd.n6916 gnd.n172 19.3944
R14801 gnd.n6916 gnd.n173 19.3944
R14802 gnd.n6912 gnd.n173 19.3944
R14803 gnd.n6912 gnd.n6911 19.3944
R14804 gnd.n6911 gnd.n6910 19.3944
R14805 gnd.n4079 gnd.n999 19.3944
R14806 gnd.n4079 gnd.n4078 19.3944
R14807 gnd.n4182 gnd.n4078 19.3944
R14808 gnd.n4182 gnd.n4181 19.3944
R14809 gnd.n4181 gnd.n4086 19.3944
R14810 gnd.n4174 gnd.n4086 19.3944
R14811 gnd.n4174 gnd.n4173 19.3944
R14812 gnd.n4173 gnd.n4097 19.3944
R14813 gnd.n4166 gnd.n4097 19.3944
R14814 gnd.n4166 gnd.n4165 19.3944
R14815 gnd.n4165 gnd.n4108 19.3944
R14816 gnd.n4158 gnd.n4108 19.3944
R14817 gnd.n4158 gnd.n4157 19.3944
R14818 gnd.n4157 gnd.n4120 19.3944
R14819 gnd.n4150 gnd.n4120 19.3944
R14820 gnd.n4150 gnd.n4149 19.3944
R14821 gnd.n6541 gnd.n405 19.3944
R14822 gnd.n6541 gnd.n401 19.3944
R14823 gnd.n6547 gnd.n401 19.3944
R14824 gnd.n6547 gnd.n399 19.3944
R14825 gnd.n6551 gnd.n399 19.3944
R14826 gnd.n6551 gnd.n395 19.3944
R14827 gnd.n6557 gnd.n395 19.3944
R14828 gnd.n6557 gnd.n393 19.3944
R14829 gnd.n6561 gnd.n393 19.3944
R14830 gnd.n6561 gnd.n389 19.3944
R14831 gnd.n6567 gnd.n389 19.3944
R14832 gnd.n6567 gnd.n387 19.3944
R14833 gnd.n6571 gnd.n387 19.3944
R14834 gnd.n6571 gnd.n383 19.3944
R14835 gnd.n6577 gnd.n383 19.3944
R14836 gnd.n6577 gnd.n381 19.3944
R14837 gnd.n6581 gnd.n381 19.3944
R14838 gnd.n6581 gnd.n377 19.3944
R14839 gnd.n6587 gnd.n377 19.3944
R14840 gnd.n6587 gnd.n375 19.3944
R14841 gnd.n6591 gnd.n375 19.3944
R14842 gnd.n6591 gnd.n371 19.3944
R14843 gnd.n6597 gnd.n371 19.3944
R14844 gnd.n6597 gnd.n369 19.3944
R14845 gnd.n6601 gnd.n369 19.3944
R14846 gnd.n6601 gnd.n365 19.3944
R14847 gnd.n6607 gnd.n365 19.3944
R14848 gnd.n6607 gnd.n363 19.3944
R14849 gnd.n6611 gnd.n363 19.3944
R14850 gnd.n6611 gnd.n359 19.3944
R14851 gnd.n6617 gnd.n359 19.3944
R14852 gnd.n6617 gnd.n357 19.3944
R14853 gnd.n6621 gnd.n357 19.3944
R14854 gnd.n6621 gnd.n353 19.3944
R14855 gnd.n6627 gnd.n353 19.3944
R14856 gnd.n6627 gnd.n351 19.3944
R14857 gnd.n6631 gnd.n351 19.3944
R14858 gnd.n6631 gnd.n347 19.3944
R14859 gnd.n6637 gnd.n347 19.3944
R14860 gnd.n6637 gnd.n345 19.3944
R14861 gnd.n6641 gnd.n345 19.3944
R14862 gnd.n6641 gnd.n341 19.3944
R14863 gnd.n6647 gnd.n341 19.3944
R14864 gnd.n6647 gnd.n339 19.3944
R14865 gnd.n6651 gnd.n339 19.3944
R14866 gnd.n6651 gnd.n335 19.3944
R14867 gnd.n6657 gnd.n335 19.3944
R14868 gnd.n6657 gnd.n333 19.3944
R14869 gnd.n6661 gnd.n333 19.3944
R14870 gnd.n6661 gnd.n329 19.3944
R14871 gnd.n6667 gnd.n329 19.3944
R14872 gnd.n6667 gnd.n327 19.3944
R14873 gnd.n6671 gnd.n327 19.3944
R14874 gnd.n6671 gnd.n323 19.3944
R14875 gnd.n6677 gnd.n323 19.3944
R14876 gnd.n6677 gnd.n321 19.3944
R14877 gnd.n6681 gnd.n321 19.3944
R14878 gnd.n6681 gnd.n317 19.3944
R14879 gnd.n6687 gnd.n317 19.3944
R14880 gnd.n6687 gnd.n315 19.3944
R14881 gnd.n6691 gnd.n315 19.3944
R14882 gnd.n6691 gnd.n311 19.3944
R14883 gnd.n6697 gnd.n311 19.3944
R14884 gnd.n6697 gnd.n309 19.3944
R14885 gnd.n6701 gnd.n309 19.3944
R14886 gnd.n6701 gnd.n305 19.3944
R14887 gnd.n6707 gnd.n305 19.3944
R14888 gnd.n6707 gnd.n303 19.3944
R14889 gnd.n6711 gnd.n303 19.3944
R14890 gnd.n6711 gnd.n299 19.3944
R14891 gnd.n6717 gnd.n299 19.3944
R14892 gnd.n6717 gnd.n297 19.3944
R14893 gnd.n6721 gnd.n297 19.3944
R14894 gnd.n6721 gnd.n293 19.3944
R14895 gnd.n6727 gnd.n293 19.3944
R14896 gnd.n6727 gnd.n291 19.3944
R14897 gnd.n6731 gnd.n291 19.3944
R14898 gnd.n6731 gnd.n287 19.3944
R14899 gnd.n6737 gnd.n287 19.3944
R14900 gnd.n6737 gnd.n285 19.3944
R14901 gnd.n6743 gnd.n285 19.3944
R14902 gnd.n6743 gnd.n6742 19.3944
R14903 gnd.n6742 gnd.n281 19.3944
R14904 gnd.n6750 gnd.n281 19.3944
R14905 gnd.n6121 gnd.n657 19.3944
R14906 gnd.n6121 gnd.n653 19.3944
R14907 gnd.n6127 gnd.n653 19.3944
R14908 gnd.n6127 gnd.n651 19.3944
R14909 gnd.n6131 gnd.n651 19.3944
R14910 gnd.n6131 gnd.n647 19.3944
R14911 gnd.n6137 gnd.n647 19.3944
R14912 gnd.n6137 gnd.n645 19.3944
R14913 gnd.n6141 gnd.n645 19.3944
R14914 gnd.n6141 gnd.n641 19.3944
R14915 gnd.n6147 gnd.n641 19.3944
R14916 gnd.n6147 gnd.n639 19.3944
R14917 gnd.n6151 gnd.n639 19.3944
R14918 gnd.n6151 gnd.n635 19.3944
R14919 gnd.n6157 gnd.n635 19.3944
R14920 gnd.n6157 gnd.n633 19.3944
R14921 gnd.n6161 gnd.n633 19.3944
R14922 gnd.n6161 gnd.n629 19.3944
R14923 gnd.n6167 gnd.n629 19.3944
R14924 gnd.n6167 gnd.n627 19.3944
R14925 gnd.n6171 gnd.n627 19.3944
R14926 gnd.n6171 gnd.n623 19.3944
R14927 gnd.n6177 gnd.n623 19.3944
R14928 gnd.n6177 gnd.n621 19.3944
R14929 gnd.n6181 gnd.n621 19.3944
R14930 gnd.n6181 gnd.n617 19.3944
R14931 gnd.n6187 gnd.n617 19.3944
R14932 gnd.n6187 gnd.n615 19.3944
R14933 gnd.n6191 gnd.n615 19.3944
R14934 gnd.n6191 gnd.n611 19.3944
R14935 gnd.n6197 gnd.n611 19.3944
R14936 gnd.n6197 gnd.n609 19.3944
R14937 gnd.n6201 gnd.n609 19.3944
R14938 gnd.n6201 gnd.n605 19.3944
R14939 gnd.n6207 gnd.n605 19.3944
R14940 gnd.n6207 gnd.n603 19.3944
R14941 gnd.n6211 gnd.n603 19.3944
R14942 gnd.n6211 gnd.n599 19.3944
R14943 gnd.n6217 gnd.n599 19.3944
R14944 gnd.n6217 gnd.n597 19.3944
R14945 gnd.n6221 gnd.n597 19.3944
R14946 gnd.n6221 gnd.n593 19.3944
R14947 gnd.n6227 gnd.n593 19.3944
R14948 gnd.n6227 gnd.n591 19.3944
R14949 gnd.n6231 gnd.n591 19.3944
R14950 gnd.n6231 gnd.n587 19.3944
R14951 gnd.n6237 gnd.n587 19.3944
R14952 gnd.n6237 gnd.n585 19.3944
R14953 gnd.n6241 gnd.n585 19.3944
R14954 gnd.n6241 gnd.n581 19.3944
R14955 gnd.n6247 gnd.n581 19.3944
R14956 gnd.n6247 gnd.n579 19.3944
R14957 gnd.n6251 gnd.n579 19.3944
R14958 gnd.n6251 gnd.n575 19.3944
R14959 gnd.n6257 gnd.n575 19.3944
R14960 gnd.n6257 gnd.n573 19.3944
R14961 gnd.n6261 gnd.n573 19.3944
R14962 gnd.n6261 gnd.n569 19.3944
R14963 gnd.n6267 gnd.n569 19.3944
R14964 gnd.n6267 gnd.n567 19.3944
R14965 gnd.n6271 gnd.n567 19.3944
R14966 gnd.n6271 gnd.n563 19.3944
R14967 gnd.n6277 gnd.n563 19.3944
R14968 gnd.n6277 gnd.n561 19.3944
R14969 gnd.n6281 gnd.n561 19.3944
R14970 gnd.n6281 gnd.n557 19.3944
R14971 gnd.n6287 gnd.n557 19.3944
R14972 gnd.n6287 gnd.n555 19.3944
R14973 gnd.n6291 gnd.n555 19.3944
R14974 gnd.n6291 gnd.n551 19.3944
R14975 gnd.n6297 gnd.n551 19.3944
R14976 gnd.n6297 gnd.n549 19.3944
R14977 gnd.n6301 gnd.n549 19.3944
R14978 gnd.n6301 gnd.n545 19.3944
R14979 gnd.n6307 gnd.n545 19.3944
R14980 gnd.n6307 gnd.n543 19.3944
R14981 gnd.n6311 gnd.n543 19.3944
R14982 gnd.n6311 gnd.n539 19.3944
R14983 gnd.n6317 gnd.n539 19.3944
R14984 gnd.n6317 gnd.n537 19.3944
R14985 gnd.n6321 gnd.n537 19.3944
R14986 gnd.n6321 gnd.n533 19.3944
R14987 gnd.n6327 gnd.n533 19.3944
R14988 gnd.n6327 gnd.n531 19.3944
R14989 gnd.n6331 gnd.n531 19.3944
R14990 gnd.n6331 gnd.n527 19.3944
R14991 gnd.n6337 gnd.n527 19.3944
R14992 gnd.n6337 gnd.n525 19.3944
R14993 gnd.n6341 gnd.n525 19.3944
R14994 gnd.n6341 gnd.n521 19.3944
R14995 gnd.n6347 gnd.n521 19.3944
R14996 gnd.n6347 gnd.n519 19.3944
R14997 gnd.n6351 gnd.n519 19.3944
R14998 gnd.n6351 gnd.n515 19.3944
R14999 gnd.n6357 gnd.n515 19.3944
R15000 gnd.n6357 gnd.n513 19.3944
R15001 gnd.n6361 gnd.n513 19.3944
R15002 gnd.n6361 gnd.n509 19.3944
R15003 gnd.n6367 gnd.n509 19.3944
R15004 gnd.n6367 gnd.n507 19.3944
R15005 gnd.n6371 gnd.n507 19.3944
R15006 gnd.n6371 gnd.n503 19.3944
R15007 gnd.n6377 gnd.n503 19.3944
R15008 gnd.n6377 gnd.n501 19.3944
R15009 gnd.n6381 gnd.n501 19.3944
R15010 gnd.n6381 gnd.n497 19.3944
R15011 gnd.n6387 gnd.n497 19.3944
R15012 gnd.n6387 gnd.n495 19.3944
R15013 gnd.n6391 gnd.n495 19.3944
R15014 gnd.n6391 gnd.n491 19.3944
R15015 gnd.n6397 gnd.n491 19.3944
R15016 gnd.n6397 gnd.n489 19.3944
R15017 gnd.n6401 gnd.n489 19.3944
R15018 gnd.n6401 gnd.n485 19.3944
R15019 gnd.n6407 gnd.n485 19.3944
R15020 gnd.n6407 gnd.n483 19.3944
R15021 gnd.n6411 gnd.n483 19.3944
R15022 gnd.n6411 gnd.n479 19.3944
R15023 gnd.n6417 gnd.n479 19.3944
R15024 gnd.n6417 gnd.n477 19.3944
R15025 gnd.n6421 gnd.n477 19.3944
R15026 gnd.n6421 gnd.n473 19.3944
R15027 gnd.n6427 gnd.n473 19.3944
R15028 gnd.n6427 gnd.n471 19.3944
R15029 gnd.n6431 gnd.n471 19.3944
R15030 gnd.n6431 gnd.n467 19.3944
R15031 gnd.n6437 gnd.n467 19.3944
R15032 gnd.n6437 gnd.n465 19.3944
R15033 gnd.n6441 gnd.n465 19.3944
R15034 gnd.n6441 gnd.n461 19.3944
R15035 gnd.n6447 gnd.n461 19.3944
R15036 gnd.n6447 gnd.n459 19.3944
R15037 gnd.n6451 gnd.n459 19.3944
R15038 gnd.n6451 gnd.n455 19.3944
R15039 gnd.n6457 gnd.n455 19.3944
R15040 gnd.n6457 gnd.n453 19.3944
R15041 gnd.n6461 gnd.n453 19.3944
R15042 gnd.n6461 gnd.n449 19.3944
R15043 gnd.n6467 gnd.n449 19.3944
R15044 gnd.n6467 gnd.n447 19.3944
R15045 gnd.n6471 gnd.n447 19.3944
R15046 gnd.n6471 gnd.n443 19.3944
R15047 gnd.n6477 gnd.n443 19.3944
R15048 gnd.n6477 gnd.n441 19.3944
R15049 gnd.n6481 gnd.n441 19.3944
R15050 gnd.n6481 gnd.n437 19.3944
R15051 gnd.n6487 gnd.n437 19.3944
R15052 gnd.n6487 gnd.n435 19.3944
R15053 gnd.n6491 gnd.n435 19.3944
R15054 gnd.n6491 gnd.n431 19.3944
R15055 gnd.n6497 gnd.n431 19.3944
R15056 gnd.n6497 gnd.n429 19.3944
R15057 gnd.n6501 gnd.n429 19.3944
R15058 gnd.n6501 gnd.n425 19.3944
R15059 gnd.n6507 gnd.n425 19.3944
R15060 gnd.n6507 gnd.n423 19.3944
R15061 gnd.n6511 gnd.n423 19.3944
R15062 gnd.n6511 gnd.n419 19.3944
R15063 gnd.n6517 gnd.n419 19.3944
R15064 gnd.n6517 gnd.n417 19.3944
R15065 gnd.n6521 gnd.n417 19.3944
R15066 gnd.n6521 gnd.n413 19.3944
R15067 gnd.n6527 gnd.n413 19.3944
R15068 gnd.n6527 gnd.n411 19.3944
R15069 gnd.n6531 gnd.n411 19.3944
R15070 gnd.n6531 gnd.n407 19.3944
R15071 gnd.n6537 gnd.n407 19.3944
R15072 gnd.n5370 gnd.n5367 19.3944
R15073 gnd.n5370 gnd.n5366 19.3944
R15074 gnd.n5376 gnd.n5366 19.3944
R15075 gnd.n5376 gnd.n5364 19.3944
R15076 gnd.n5380 gnd.n5364 19.3944
R15077 gnd.n5380 gnd.n5362 19.3944
R15078 gnd.n5386 gnd.n5362 19.3944
R15079 gnd.n5386 gnd.n5360 19.3944
R15080 gnd.n5390 gnd.n5360 19.3944
R15081 gnd.n5390 gnd.n5358 19.3944
R15082 gnd.n5396 gnd.n5358 19.3944
R15083 gnd.n5396 gnd.n5356 19.3944
R15084 gnd.n5401 gnd.n5356 19.3944
R15085 gnd.n5401 gnd.n5354 19.3944
R15086 gnd.n5354 gnd.n1291 19.3944
R15087 gnd.n5414 gnd.n1289 19.3944
R15088 gnd.n5414 gnd.n1287 19.3944
R15089 gnd.n5420 gnd.n1287 19.3944
R15090 gnd.n5420 gnd.n1285 19.3944
R15091 gnd.n5424 gnd.n1285 19.3944
R15092 gnd.n5424 gnd.n1283 19.3944
R15093 gnd.n5430 gnd.n1283 19.3944
R15094 gnd.n5430 gnd.n1281 19.3944
R15095 gnd.n5434 gnd.n1281 19.3944
R15096 gnd.n5434 gnd.n1279 19.3944
R15097 gnd.n5440 gnd.n1279 19.3944
R15098 gnd.n5440 gnd.n1277 19.3944
R15099 gnd.n5444 gnd.n1277 19.3944
R15100 gnd.n5444 gnd.n1275 19.3944
R15101 gnd.n5450 gnd.n1275 19.3944
R15102 gnd.n5450 gnd.n1273 19.3944
R15103 gnd.n5455 gnd.n1273 19.3944
R15104 gnd.n5455 gnd.n1271 19.3944
R15105 gnd.n5466 gnd.n1266 19.3944
R15106 gnd.n5466 gnd.n1261 19.3944
R15107 gnd.n5479 gnd.n1261 19.3944
R15108 gnd.n5479 gnd.n1259 19.3944
R15109 gnd.n5524 gnd.n1259 19.3944
R15110 gnd.n5524 gnd.n5523 19.3944
R15111 gnd.n5523 gnd.n5522 19.3944
R15112 gnd.n5522 gnd.n5520 19.3944
R15113 gnd.n5520 gnd.n5519 19.3944
R15114 gnd.n5519 gnd.n5518 19.3944
R15115 gnd.n5518 gnd.n5516 19.3944
R15116 gnd.n5516 gnd.n5515 19.3944
R15117 gnd.n5515 gnd.n5513 19.3944
R15118 gnd.n5513 gnd.n5512 19.3944
R15119 gnd.n5512 gnd.n5511 19.3944
R15120 gnd.n5511 gnd.n5509 19.3944
R15121 gnd.n5509 gnd.n5508 19.3944
R15122 gnd.n5508 gnd.n5505 19.3944
R15123 gnd.n5505 gnd.n5504 19.3944
R15124 gnd.n5504 gnd.n5502 19.3944
R15125 gnd.n5502 gnd.n5501 19.3944
R15126 gnd.n5501 gnd.n237 19.3944
R15127 gnd.n6781 gnd.n237 19.3944
R15128 gnd.n6781 gnd.n6780 19.3944
R15129 gnd.n6780 gnd.n6779 19.3944
R15130 gnd.n6779 gnd.n6775 19.3944
R15131 gnd.n6775 gnd.n6774 19.3944
R15132 gnd.n6774 gnd.n6771 19.3944
R15133 gnd.n6771 gnd.n6770 19.3944
R15134 gnd.n6770 gnd.n6766 19.3944
R15135 gnd.n6766 gnd.n6765 19.3944
R15136 gnd.n6765 gnd.n269 19.3944
R15137 gnd.n269 gnd.n268 19.3944
R15138 gnd.n268 gnd.n264 19.3944
R15139 gnd.n264 gnd.n263 19.3944
R15140 gnd.n263 gnd.n260 19.3944
R15141 gnd.n260 gnd.n259 19.3944
R15142 gnd.n259 gnd.n257 19.3944
R15143 gnd.n257 gnd.n256 19.3944
R15144 gnd.n256 gnd.n159 19.3944
R15145 gnd.n6929 gnd.n159 19.3944
R15146 gnd.n6930 gnd.n6929 19.3944
R15147 gnd.n6968 gnd.n120 19.3944
R15148 gnd.n6963 gnd.n120 19.3944
R15149 gnd.n6963 gnd.n6962 19.3944
R15150 gnd.n6962 gnd.n6961 19.3944
R15151 gnd.n6961 gnd.n127 19.3944
R15152 gnd.n6956 gnd.n127 19.3944
R15153 gnd.n6956 gnd.n6955 19.3944
R15154 gnd.n6955 gnd.n6954 19.3944
R15155 gnd.n6954 gnd.n134 19.3944
R15156 gnd.n6949 gnd.n134 19.3944
R15157 gnd.n6949 gnd.n6948 19.3944
R15158 gnd.n6948 gnd.n6947 19.3944
R15159 gnd.n6947 gnd.n141 19.3944
R15160 gnd.n6942 gnd.n141 19.3944
R15161 gnd.n6942 gnd.n6941 19.3944
R15162 gnd.n6941 gnd.n6940 19.3944
R15163 gnd.n6940 gnd.n148 19.3944
R15164 gnd.n6935 gnd.n148 19.3944
R15165 gnd.n7001 gnd.n7000 19.3944
R15166 gnd.n7000 gnd.n6999 19.3944
R15167 gnd.n6999 gnd.n92 19.3944
R15168 gnd.n6994 gnd.n92 19.3944
R15169 gnd.n6994 gnd.n6993 19.3944
R15170 gnd.n6993 gnd.n6992 19.3944
R15171 gnd.n6992 gnd.n99 19.3944
R15172 gnd.n6987 gnd.n99 19.3944
R15173 gnd.n6987 gnd.n6986 19.3944
R15174 gnd.n6986 gnd.n6985 19.3944
R15175 gnd.n6985 gnd.n106 19.3944
R15176 gnd.n6980 gnd.n106 19.3944
R15177 gnd.n6980 gnd.n6979 19.3944
R15178 gnd.n6979 gnd.n6978 19.3944
R15179 gnd.n6978 gnd.n113 19.3944
R15180 gnd.n6973 gnd.n113 19.3944
R15181 gnd.n6973 gnd.n6972 19.3944
R15182 gnd.n5705 gnd.n5704 19.3944
R15183 gnd.n5704 gnd.n5703 19.3944
R15184 gnd.n5703 gnd.n1136 19.3944
R15185 gnd.n5546 gnd.n1136 19.3944
R15186 gnd.n5546 gnd.n1254 19.3944
R15187 gnd.n5552 gnd.n1254 19.3944
R15188 gnd.n5552 gnd.n5551 19.3944
R15189 gnd.n5551 gnd.n1228 19.3944
R15190 gnd.n5577 gnd.n1228 19.3944
R15191 gnd.n5577 gnd.n1226 19.3944
R15192 gnd.n5584 gnd.n1226 19.3944
R15193 gnd.n5584 gnd.n5583 19.3944
R15194 gnd.n5583 gnd.n1198 19.3944
R15195 gnd.n5615 gnd.n1198 19.3944
R15196 gnd.n5616 gnd.n5615 19.3944
R15197 gnd.n5617 gnd.n5616 19.3944
R15198 gnd.n1183 gnd.n1182 19.3944
R15199 gnd.n5636 gnd.n5635 19.3944
R15200 gnd.n5633 gnd.n5632 19.3944
R15201 gnd.n6786 gnd.n6785 19.3944
R15202 gnd.n6798 gnd.n221 19.3944
R15203 gnd.n6798 gnd.n213 19.3944
R15204 gnd.n6802 gnd.n213 19.3944
R15205 gnd.n6802 gnd.n200 19.3944
R15206 gnd.n6814 gnd.n200 19.3944
R15207 gnd.n6814 gnd.n198 19.3944
R15208 gnd.n6818 gnd.n198 19.3944
R15209 gnd.n6818 gnd.n184 19.3944
R15210 gnd.n6830 gnd.n184 19.3944
R15211 gnd.n6830 gnd.n182 19.3944
R15212 gnd.n6834 gnd.n182 19.3944
R15213 gnd.n6834 gnd.n166 19.3944
R15214 gnd.n6920 gnd.n166 19.3944
R15215 gnd.n6920 gnd.n164 19.3944
R15216 gnd.n6924 gnd.n164 19.3944
R15217 gnd.n6924 gnd.n87 19.3944
R15218 gnd.n7004 gnd.n87 19.3944
R15219 gnd.n3852 gnd.n3851 19.3944
R15220 gnd.n3855 gnd.n3852 19.3944
R15221 gnd.n3855 gnd.n3848 19.3944
R15222 gnd.n3859 gnd.n3848 19.3944
R15223 gnd.n3859 gnd.n2072 19.3944
R15224 gnd.n3863 gnd.n2072 19.3944
R15225 gnd.n3863 gnd.n2070 19.3944
R15226 gnd.n3870 gnd.n2070 19.3944
R15227 gnd.n3870 gnd.n3869 19.3944
R15228 gnd.n3869 gnd.n3868 19.3944
R15229 gnd.n3897 gnd.n3896 19.3944
R15230 gnd.n3907 gnd.n3906 19.3944
R15231 gnd.n3904 gnd.n3901 19.3944
R15232 gnd.n3899 gnd.n2013 19.3944
R15233 gnd.n3961 gnd.n3960 19.3944
R15234 gnd.n3966 gnd.n3961 19.3944
R15235 gnd.n3966 gnd.n3965 19.3944
R15236 gnd.n3965 gnd.n1986 19.3944
R15237 gnd.n4025 gnd.n1986 19.3944
R15238 gnd.n4025 gnd.n1984 19.3944
R15239 gnd.n4029 gnd.n1984 19.3944
R15240 gnd.n4029 gnd.n1982 19.3944
R15241 gnd.n4033 gnd.n1982 19.3944
R15242 gnd.n4033 gnd.n1980 19.3944
R15243 gnd.n4037 gnd.n1980 19.3944
R15244 gnd.n4037 gnd.n1978 19.3944
R15245 gnd.n4041 gnd.n1978 19.3944
R15246 gnd.n4041 gnd.n1976 19.3944
R15247 gnd.n4045 gnd.n1976 19.3944
R15248 gnd.n4045 gnd.n1974 19.3944
R15249 gnd.n4049 gnd.n1974 19.3944
R15250 gnd.n4049 gnd.n1972 19.3944
R15251 gnd.n4053 gnd.n1972 19.3944
R15252 gnd.n4053 gnd.n1968 19.3944
R15253 gnd.n4192 gnd.n1968 19.3944
R15254 gnd.n4192 gnd.n1966 19.3944
R15255 gnd.n4196 gnd.n1966 19.3944
R15256 gnd.n4196 gnd.n1962 19.3944
R15257 gnd.n4206 gnd.n1962 19.3944
R15258 gnd.n4206 gnd.n1960 19.3944
R15259 gnd.n4210 gnd.n1960 19.3944
R15260 gnd.n4210 gnd.n1954 19.3944
R15261 gnd.n4220 gnd.n1954 19.3944
R15262 gnd.n4220 gnd.n1952 19.3944
R15263 gnd.n4224 gnd.n1952 19.3944
R15264 gnd.n4224 gnd.n1946 19.3944
R15265 gnd.n4234 gnd.n1946 19.3944
R15266 gnd.n4234 gnd.n1944 19.3944
R15267 gnd.n4238 gnd.n1944 19.3944
R15268 gnd.n4238 gnd.n1669 19.3944
R15269 gnd.n4423 gnd.n1669 19.3944
R15270 gnd.n4423 gnd.n1667 19.3944
R15271 gnd.n4427 gnd.n1667 19.3944
R15272 gnd.n4427 gnd.n1651 19.3944
R15273 gnd.n4479 gnd.n1651 19.3944
R15274 gnd.n4479 gnd.n1649 19.3944
R15275 gnd.n4483 gnd.n1649 19.3944
R15276 gnd.n4483 gnd.n1630 19.3944
R15277 gnd.n4510 gnd.n1630 19.3944
R15278 gnd.n4510 gnd.n1628 19.3944
R15279 gnd.n4516 gnd.n1628 19.3944
R15280 gnd.n4516 gnd.n4515 19.3944
R15281 gnd.n4515 gnd.n1610 19.3944
R15282 gnd.n4540 gnd.n1610 19.3944
R15283 gnd.n4540 gnd.n1608 19.3944
R15284 gnd.n4554 gnd.n1608 19.3944
R15285 gnd.n4554 gnd.n4553 19.3944
R15286 gnd.n4553 gnd.n4552 19.3944
R15287 gnd.n4552 gnd.n4547 19.3944
R15288 gnd.n4547 gnd.n1563 19.3944
R15289 gnd.n4624 gnd.n1563 19.3944
R15290 gnd.n4624 gnd.n1561 19.3944
R15291 gnd.n4628 gnd.n1561 19.3944
R15292 gnd.n4628 gnd.n1540 19.3944
R15293 gnd.n4664 gnd.n1540 19.3944
R15294 gnd.n4664 gnd.n1538 19.3944
R15295 gnd.n4668 gnd.n1538 19.3944
R15296 gnd.n4668 gnd.n1518 19.3944
R15297 gnd.n4718 gnd.n1518 19.3944
R15298 gnd.n4718 gnd.n1516 19.3944
R15299 gnd.n4722 gnd.n1516 19.3944
R15300 gnd.n4722 gnd.n1499 19.3944
R15301 gnd.n4743 gnd.n1499 19.3944
R15302 gnd.n4743 gnd.n1497 19.3944
R15303 gnd.n4747 gnd.n1497 19.3944
R15304 gnd.n4747 gnd.n1477 19.3944
R15305 gnd.n4802 gnd.n1477 19.3944
R15306 gnd.n4802 gnd.n1475 19.3944
R15307 gnd.n4806 gnd.n1475 19.3944
R15308 gnd.n4806 gnd.n1455 19.3944
R15309 gnd.n4831 gnd.n1455 19.3944
R15310 gnd.n4831 gnd.n1453 19.3944
R15311 gnd.n4837 gnd.n1453 19.3944
R15312 gnd.n4837 gnd.n4836 19.3944
R15313 gnd.n4836 gnd.n1427 19.3944
R15314 gnd.n4886 gnd.n1427 19.3944
R15315 gnd.n4886 gnd.n1425 19.3944
R15316 gnd.n4890 gnd.n1425 19.3944
R15317 gnd.n4890 gnd.n1410 19.3944
R15318 gnd.n4912 gnd.n1410 19.3944
R15319 gnd.n4912 gnd.n1408 19.3944
R15320 gnd.n4919 gnd.n1408 19.3944
R15321 gnd.n4919 gnd.n4918 19.3944
R15322 gnd.n4918 gnd.n1346 19.3944
R15323 gnd.n5189 gnd.n1346 19.3944
R15324 gnd.n5189 gnd.n5188 19.3944
R15325 gnd.n5188 gnd.n5187 19.3944
R15326 gnd.n5187 gnd.n1350 19.3944
R15327 gnd.n1356 gnd.n1350 19.3944
R15328 gnd.n5177 gnd.n1356 19.3944
R15329 gnd.n5177 gnd.n5176 19.3944
R15330 gnd.n5176 gnd.n5175 19.3944
R15331 gnd.n5175 gnd.n1362 19.3944
R15332 gnd.n5166 gnd.n1362 19.3944
R15333 gnd.n5166 gnd.n5165 19.3944
R15334 gnd.n5165 gnd.n5164 19.3944
R15335 gnd.n5164 gnd.n1374 19.3944
R15336 gnd.n5155 gnd.n1374 19.3944
R15337 gnd.n5155 gnd.n1111 19.3944
R15338 gnd.n5720 gnd.n1111 19.3944
R15339 gnd.n5720 gnd.n5719 19.3944
R15340 gnd.n5719 gnd.n5718 19.3944
R15341 gnd.n5718 gnd.n1115 19.3944
R15342 gnd.n5712 gnd.n1115 19.3944
R15343 gnd.n5712 gnd.n5711 19.3944
R15344 gnd.n5711 gnd.n5710 19.3944
R15345 gnd.n5710 gnd.n1124 19.3944
R15346 gnd.n5532 gnd.n1124 19.3944
R15347 gnd.n5535 gnd.n5532 19.3944
R15348 gnd.n5535 gnd.n5529 19.3944
R15349 gnd.n5541 gnd.n5529 19.3944
R15350 gnd.n5541 gnd.n5540 19.3944
R15351 gnd.n5540 gnd.n1238 19.3944
R15352 gnd.n5566 gnd.n1238 19.3944
R15353 gnd.n5566 gnd.n1236 19.3944
R15354 gnd.n5572 gnd.n1236 19.3944
R15355 gnd.n5572 gnd.n5571 19.3944
R15356 gnd.n5571 gnd.n1210 19.3944
R15357 gnd.n5598 gnd.n1210 19.3944
R15358 gnd.n5598 gnd.n1208 19.3944
R15359 gnd.n5610 gnd.n1208 19.3944
R15360 gnd.n5610 gnd.n5609 19.3944
R15361 gnd.n5609 gnd.n5608 19.3944
R15362 gnd.n5605 gnd.n5604 19.3944
R15363 gnd.n5642 gnd.n5641 19.3944
R15364 gnd.n5663 gnd.n5662 19.3944
R15365 gnd.n5660 gnd.n5644 19.3944
R15366 gnd.n5656 gnd.n5655 19.3944
R15367 gnd.n5655 gnd.n5654 19.3944
R15368 gnd.n5654 gnd.n5651 19.3944
R15369 gnd.n5651 gnd.n272 19.3944
R15370 gnd.n6760 gnd.n272 19.3944
R15371 gnd.n6760 gnd.n6759 19.3944
R15372 gnd.n6759 gnd.n6758 19.3944
R15373 gnd.n6758 gnd.n276 19.3944
R15374 gnd.n6754 gnd.n276 19.3944
R15375 gnd.n6754 gnd.n6753 19.3944
R15376 gnd.n3782 gnd.n3781 19.3944
R15377 gnd.n3781 gnd.n3780 19.3944
R15378 gnd.n3780 gnd.n3779 19.3944
R15379 gnd.n3779 gnd.n3777 19.3944
R15380 gnd.n3777 gnd.n3774 19.3944
R15381 gnd.n3774 gnd.n3773 19.3944
R15382 gnd.n3773 gnd.n3770 19.3944
R15383 gnd.n3770 gnd.n3769 19.3944
R15384 gnd.n3769 gnd.n3766 19.3944
R15385 gnd.n3766 gnd.n3765 19.3944
R15386 gnd.n3765 gnd.n3762 19.3944
R15387 gnd.n3762 gnd.n3761 19.3944
R15388 gnd.n3761 gnd.n3758 19.3944
R15389 gnd.n3758 gnd.n3757 19.3944
R15390 gnd.n3757 gnd.n3754 19.3944
R15391 gnd.n3754 gnd.n3753 19.3944
R15392 gnd.n3753 gnd.n3750 19.3944
R15393 gnd.n3748 gnd.n3745 19.3944
R15394 gnd.n3745 gnd.n3744 19.3944
R15395 gnd.n3744 gnd.n3741 19.3944
R15396 gnd.n3741 gnd.n3740 19.3944
R15397 gnd.n3740 gnd.n3737 19.3944
R15398 gnd.n3737 gnd.n3736 19.3944
R15399 gnd.n3736 gnd.n3733 19.3944
R15400 gnd.n3733 gnd.n3732 19.3944
R15401 gnd.n3732 gnd.n3729 19.3944
R15402 gnd.n3729 gnd.n3728 19.3944
R15403 gnd.n3728 gnd.n3725 19.3944
R15404 gnd.n3725 gnd.n3724 19.3944
R15405 gnd.n3724 gnd.n3721 19.3944
R15406 gnd.n3721 gnd.n3720 19.3944
R15407 gnd.n3720 gnd.n3717 19.3944
R15408 gnd.n3717 gnd.n3716 19.3944
R15409 gnd.n3716 gnd.n3713 19.3944
R15410 gnd.n3713 gnd.n3712 19.3944
R15411 gnd.n3801 gnd.n2100 19.3944
R15412 gnd.n3801 gnd.n2101 19.3944
R15413 gnd.n3797 gnd.n2101 19.3944
R15414 gnd.n3797 gnd.n3796 19.3944
R15415 gnd.n3796 gnd.n3794 19.3944
R15416 gnd.n3794 gnd.n846 19.3944
R15417 gnd.n5938 gnd.n846 19.3944
R15418 gnd.n5938 gnd.n5937 19.3944
R15419 gnd.n5937 gnd.n5936 19.3944
R15420 gnd.n5936 gnd.n850 19.3944
R15421 gnd.n5926 gnd.n850 19.3944
R15422 gnd.n5926 gnd.n5925 19.3944
R15423 gnd.n5925 gnd.n5924 19.3944
R15424 gnd.n5924 gnd.n871 19.3944
R15425 gnd.n5914 gnd.n871 19.3944
R15426 gnd.n5914 gnd.n5913 19.3944
R15427 gnd.n5913 gnd.n5912 19.3944
R15428 gnd.n5912 gnd.n892 19.3944
R15429 gnd.n3914 gnd.n892 19.3944
R15430 gnd.n3915 gnd.n3914 19.3944
R15431 gnd.n3915 gnd.n2031 19.3944
R15432 gnd.n3940 gnd.n2031 19.3944
R15433 gnd.n3940 gnd.n3939 19.3944
R15434 gnd.n3939 gnd.n3938 19.3944
R15435 gnd.n3938 gnd.n915 19.3944
R15436 gnd.n5900 gnd.n915 19.3944
R15437 gnd.n5900 gnd.n5899 19.3944
R15438 gnd.n5899 gnd.n5898 19.3944
R15439 gnd.n5898 gnd.n919 19.3944
R15440 gnd.n5888 gnd.n919 19.3944
R15441 gnd.n5888 gnd.n5887 19.3944
R15442 gnd.n5887 gnd.n5886 19.3944
R15443 gnd.n5886 gnd.n938 19.3944
R15444 gnd.n5876 gnd.n938 19.3944
R15445 gnd.n5876 gnd.n5875 19.3944
R15446 gnd.n5875 gnd.n5874 19.3944
R15447 gnd.n5874 gnd.n960 19.3944
R15448 gnd.n5864 gnd.n960 19.3944
R15449 gnd.n5864 gnd.n5863 19.3944
R15450 gnd.n5863 gnd.n5862 19.3944
R15451 gnd.n5862 gnd.n981 19.3944
R15452 gnd.n5852 gnd.n981 19.3944
R15453 gnd.n3788 gnd.n2103 19.3944
R15454 gnd.n3596 gnd.n2103 19.3944
R15455 gnd.n3597 gnd.n3596 19.3944
R15456 gnd.n3600 gnd.n3597 19.3944
R15457 gnd.n3600 gnd.n3592 19.3944
R15458 gnd.n3606 gnd.n3592 19.3944
R15459 gnd.n3607 gnd.n3606 19.3944
R15460 gnd.n3610 gnd.n3607 19.3944
R15461 gnd.n3610 gnd.n3590 19.3944
R15462 gnd.n3616 gnd.n3590 19.3944
R15463 gnd.n3617 gnd.n3616 19.3944
R15464 gnd.n3620 gnd.n3617 19.3944
R15465 gnd.n3620 gnd.n3588 19.3944
R15466 gnd.n3626 gnd.n3588 19.3944
R15467 gnd.n3627 gnd.n3626 19.3944
R15468 gnd.n3630 gnd.n3627 19.3944
R15469 gnd.n3638 gnd.n3637 19.3944
R15470 gnd.n3637 gnd.n3636 19.3944
R15471 gnd.n3636 gnd.n2084 19.3944
R15472 gnd.n3815 gnd.n2084 19.3944
R15473 gnd.n3816 gnd.n3815 19.3944
R15474 gnd.n3818 gnd.n3816 19.3944
R15475 gnd.n3818 gnd.n2082 19.3944
R15476 gnd.n3823 gnd.n2082 19.3944
R15477 gnd.n3823 gnd.n2074 19.3944
R15478 gnd.n3843 gnd.n2074 19.3944
R15479 gnd.n3843 gnd.n3842 19.3944
R15480 gnd.n3842 gnd.n3841 19.3944
R15481 gnd.n3841 gnd.n2066 19.3944
R15482 gnd.n3875 gnd.n2066 19.3944
R15483 gnd.n3875 gnd.n2064 19.3944
R15484 gnd.n3881 gnd.n2064 19.3944
R15485 gnd.n3881 gnd.n3880 19.3944
R15486 gnd.n3880 gnd.n2053 19.3944
R15487 gnd.n3922 gnd.n2053 19.3944
R15488 gnd.n3922 gnd.n2051 19.3944
R15489 gnd.n3926 gnd.n2051 19.3944
R15490 gnd.n3926 gnd.n2019 19.3944
R15491 gnd.n3950 gnd.n2019 19.3944
R15492 gnd.n3950 gnd.n2017 19.3944
R15493 gnd.n3954 gnd.n2017 19.3944
R15494 gnd.n3954 gnd.n2007 19.3944
R15495 gnd.n3971 gnd.n2007 19.3944
R15496 gnd.n3971 gnd.n2005 19.3944
R15497 gnd.n3975 gnd.n2005 19.3944
R15498 gnd.n3975 gnd.n1989 19.3944
R15499 gnd.n4020 gnd.n1989 19.3944
R15500 gnd.n4020 gnd.n1990 19.3944
R15501 gnd.n4016 gnd.n1990 19.3944
R15502 gnd.n4016 gnd.n4015 19.3944
R15503 gnd.n4015 gnd.n4014 19.3944
R15504 gnd.n4014 gnd.n1995 19.3944
R15505 gnd.n4010 gnd.n1995 19.3944
R15506 gnd.n4010 gnd.n4009 19.3944
R15507 gnd.n4009 gnd.n4008 19.3944
R15508 gnd.n4008 gnd.n1905 19.3944
R15509 gnd.n4299 gnd.n1905 19.3944
R15510 gnd.n4299 gnd.n1906 19.3944
R15511 gnd.n3705 gnd.n3704 19.3944
R15512 gnd.n3704 gnd.n3690 19.3944
R15513 gnd.n3700 gnd.n3690 19.3944
R15514 gnd.n3700 gnd.n3699 19.3944
R15515 gnd.n3699 gnd.n3697 19.3944
R15516 gnd.n3697 gnd.n3696 19.3944
R15517 gnd.n3696 gnd.n2080 19.3944
R15518 gnd.n3827 gnd.n2080 19.3944
R15519 gnd.n3828 gnd.n3827 19.3944
R15520 gnd.n3829 gnd.n3828 19.3944
R15521 gnd.n3829 gnd.n2078 19.3944
R15522 gnd.n3837 gnd.n2078 19.3944
R15523 gnd.n3837 gnd.n3836 19.3944
R15524 gnd.n3836 gnd.n3835 19.3944
R15525 gnd.n3835 gnd.n2063 19.3944
R15526 gnd.n3885 gnd.n2063 19.3944
R15527 gnd.n3885 gnd.n2061 19.3944
R15528 gnd.n3891 gnd.n2061 19.3944
R15529 gnd.n3891 gnd.n3890 19.3944
R15530 gnd.n3890 gnd.n2035 19.3944
R15531 gnd.n3930 gnd.n2035 19.3944
R15532 gnd.n3930 gnd.n2047 19.3944
R15533 gnd.n2047 gnd.n2046 19.3944
R15534 gnd.n2046 gnd.n2045 19.3944
R15535 gnd.n2045 gnd.n2043 19.3944
R15536 gnd.n2043 gnd.n2042 19.3944
R15537 gnd.n2042 gnd.n2041 19.3944
R15538 gnd.n2041 gnd.n2004 19.3944
R15539 gnd.n3979 gnd.n2004 19.3944
R15540 gnd.n3979 gnd.n2002 19.3944
R15541 gnd.n3983 gnd.n2002 19.3944
R15542 gnd.n3984 gnd.n3983 19.3944
R15543 gnd.n3987 gnd.n3984 19.3944
R15544 gnd.n3987 gnd.n2000 19.3944
R15545 gnd.n3994 gnd.n2000 19.3944
R15546 gnd.n3995 gnd.n3994 19.3944
R15547 gnd.n3998 gnd.n3995 19.3944
R15548 gnd.n3998 gnd.n1998 19.3944
R15549 gnd.n4003 gnd.n1998 19.3944
R15550 gnd.n4003 gnd.n1904 19.3944
R15551 gnd.n4303 gnd.n1904 19.3944
R15552 gnd.n4304 gnd.n4303 19.3944
R15553 gnd.n4342 gnd.n1807 19.3944
R15554 gnd.n4342 gnd.n1814 19.3944
R15555 gnd.n1871 gnd.n1814 19.3944
R15556 gnd.n4335 gnd.n1871 19.3944
R15557 gnd.n4335 gnd.n4334 19.3944
R15558 gnd.n4334 gnd.n4333 19.3944
R15559 gnd.n4333 gnd.n1877 19.3944
R15560 gnd.n4328 gnd.n1877 19.3944
R15561 gnd.n4328 gnd.n4327 19.3944
R15562 gnd.n4327 gnd.n4326 19.3944
R15563 gnd.n4326 gnd.n1884 19.3944
R15564 gnd.n4321 gnd.n1884 19.3944
R15565 gnd.n4321 gnd.n4320 19.3944
R15566 gnd.n4320 gnd.n4319 19.3944
R15567 gnd.n4319 gnd.n1891 19.3944
R15568 gnd.n4314 gnd.n1891 19.3944
R15569 gnd.n4314 gnd.n4313 19.3944
R15570 gnd.n4313 gnd.n4312 19.3944
R15571 gnd.n1827 gnd.n1826 19.3944
R15572 gnd.n1867 gnd.n1826 19.3944
R15573 gnd.n1867 gnd.n1866 19.3944
R15574 gnd.n1866 gnd.n1865 19.3944
R15575 gnd.n1865 gnd.n1862 19.3944
R15576 gnd.n1862 gnd.n1861 19.3944
R15577 gnd.n1861 gnd.n1858 19.3944
R15578 gnd.n1858 gnd.n1857 19.3944
R15579 gnd.n1857 gnd.n1854 19.3944
R15580 gnd.n1854 gnd.n1853 19.3944
R15581 gnd.n1853 gnd.n1850 19.3944
R15582 gnd.n1850 gnd.n1849 19.3944
R15583 gnd.n1849 gnd.n1846 19.3944
R15584 gnd.n1846 gnd.n1845 19.3944
R15585 gnd.n1845 gnd.n1808 19.3944
R15586 gnd.n3805 gnd.n2093 19.3944
R15587 gnd.n3805 gnd.n2091 19.3944
R15588 gnd.n3810 gnd.n2091 19.3944
R15589 gnd.n3810 gnd.n834 19.3944
R15590 gnd.n5944 gnd.n834 19.3944
R15591 gnd.n5944 gnd.n5943 19.3944
R15592 gnd.n5943 gnd.n5942 19.3944
R15593 gnd.n5942 gnd.n838 19.3944
R15594 gnd.n5932 gnd.n838 19.3944
R15595 gnd.n5932 gnd.n5931 19.3944
R15596 gnd.n5931 gnd.n5930 19.3944
R15597 gnd.n5930 gnd.n860 19.3944
R15598 gnd.n5920 gnd.n860 19.3944
R15599 gnd.n5920 gnd.n5919 19.3944
R15600 gnd.n5919 gnd.n5918 19.3944
R15601 gnd.n5918 gnd.n882 19.3944
R15602 gnd.n5908 gnd.n5907 19.3944
R15603 gnd.n3911 gnd.n899 19.3944
R15604 gnd.n2027 gnd.n2026 19.3944
R15605 gnd.n3946 gnd.n3945 19.3944
R15606 gnd.n5904 gnd.n905 19.3944
R15607 gnd.n5904 gnd.n906 19.3944
R15608 gnd.n5894 gnd.n906 19.3944
R15609 gnd.n5894 gnd.n5893 19.3944
R15610 gnd.n5893 gnd.n5892 19.3944
R15611 gnd.n5892 gnd.n928 19.3944
R15612 gnd.n5882 gnd.n928 19.3944
R15613 gnd.n5882 gnd.n5881 19.3944
R15614 gnd.n5881 gnd.n5880 19.3944
R15615 gnd.n5880 gnd.n949 19.3944
R15616 gnd.n5870 gnd.n949 19.3944
R15617 gnd.n5870 gnd.n5869 19.3944
R15618 gnd.n5869 gnd.n5868 19.3944
R15619 gnd.n5868 gnd.n970 19.3944
R15620 gnd.n5858 gnd.n970 19.3944
R15621 gnd.n5858 gnd.n5857 19.3944
R15622 gnd.n5857 gnd.n5856 19.3944
R15623 gnd.n6117 gnd.n659 19.3944
R15624 gnd.n6111 gnd.n659 19.3944
R15625 gnd.n6111 gnd.n6110 19.3944
R15626 gnd.n6110 gnd.n6109 19.3944
R15627 gnd.n6109 gnd.n666 19.3944
R15628 gnd.n6103 gnd.n666 19.3944
R15629 gnd.n6103 gnd.n6102 19.3944
R15630 gnd.n6102 gnd.n6101 19.3944
R15631 gnd.n6101 gnd.n674 19.3944
R15632 gnd.n6095 gnd.n674 19.3944
R15633 gnd.n6095 gnd.n6094 19.3944
R15634 gnd.n6094 gnd.n6093 19.3944
R15635 gnd.n6093 gnd.n682 19.3944
R15636 gnd.n6087 gnd.n682 19.3944
R15637 gnd.n6087 gnd.n6086 19.3944
R15638 gnd.n6086 gnd.n6085 19.3944
R15639 gnd.n6085 gnd.n690 19.3944
R15640 gnd.n6079 gnd.n690 19.3944
R15641 gnd.n6079 gnd.n6078 19.3944
R15642 gnd.n6078 gnd.n6077 19.3944
R15643 gnd.n6077 gnd.n698 19.3944
R15644 gnd.n6071 gnd.n698 19.3944
R15645 gnd.n6071 gnd.n6070 19.3944
R15646 gnd.n6070 gnd.n6069 19.3944
R15647 gnd.n6069 gnd.n706 19.3944
R15648 gnd.n6063 gnd.n706 19.3944
R15649 gnd.n6063 gnd.n6062 19.3944
R15650 gnd.n6062 gnd.n6061 19.3944
R15651 gnd.n6061 gnd.n714 19.3944
R15652 gnd.n6055 gnd.n714 19.3944
R15653 gnd.n6055 gnd.n6054 19.3944
R15654 gnd.n6054 gnd.n6053 19.3944
R15655 gnd.n6053 gnd.n722 19.3944
R15656 gnd.n6047 gnd.n722 19.3944
R15657 gnd.n6047 gnd.n6046 19.3944
R15658 gnd.n6046 gnd.n6045 19.3944
R15659 gnd.n6045 gnd.n730 19.3944
R15660 gnd.n6039 gnd.n730 19.3944
R15661 gnd.n6039 gnd.n6038 19.3944
R15662 gnd.n6038 gnd.n6037 19.3944
R15663 gnd.n6037 gnd.n738 19.3944
R15664 gnd.n6031 gnd.n738 19.3944
R15665 gnd.n6031 gnd.n6030 19.3944
R15666 gnd.n6030 gnd.n6029 19.3944
R15667 gnd.n6029 gnd.n746 19.3944
R15668 gnd.n6023 gnd.n746 19.3944
R15669 gnd.n6023 gnd.n6022 19.3944
R15670 gnd.n6022 gnd.n6021 19.3944
R15671 gnd.n6021 gnd.n754 19.3944
R15672 gnd.n6015 gnd.n754 19.3944
R15673 gnd.n6015 gnd.n6014 19.3944
R15674 gnd.n6014 gnd.n6013 19.3944
R15675 gnd.n6013 gnd.n762 19.3944
R15676 gnd.n6007 gnd.n762 19.3944
R15677 gnd.n6007 gnd.n6006 19.3944
R15678 gnd.n6006 gnd.n6005 19.3944
R15679 gnd.n6005 gnd.n770 19.3944
R15680 gnd.n5999 gnd.n770 19.3944
R15681 gnd.n5999 gnd.n5998 19.3944
R15682 gnd.n5998 gnd.n5997 19.3944
R15683 gnd.n5997 gnd.n778 19.3944
R15684 gnd.n5991 gnd.n778 19.3944
R15685 gnd.n5991 gnd.n5990 19.3944
R15686 gnd.n5990 gnd.n5989 19.3944
R15687 gnd.n5989 gnd.n786 19.3944
R15688 gnd.n5983 gnd.n786 19.3944
R15689 gnd.n5983 gnd.n5982 19.3944
R15690 gnd.n5982 gnd.n5981 19.3944
R15691 gnd.n5981 gnd.n794 19.3944
R15692 gnd.n5975 gnd.n794 19.3944
R15693 gnd.n5975 gnd.n5974 19.3944
R15694 gnd.n5974 gnd.n5973 19.3944
R15695 gnd.n5973 gnd.n802 19.3944
R15696 gnd.n5967 gnd.n802 19.3944
R15697 gnd.n5967 gnd.n5966 19.3944
R15698 gnd.n5966 gnd.n5965 19.3944
R15699 gnd.n5965 gnd.n810 19.3944
R15700 gnd.n5959 gnd.n810 19.3944
R15701 gnd.n5959 gnd.n5958 19.3944
R15702 gnd.n5958 gnd.n5957 19.3944
R15703 gnd.n5957 gnd.n818 19.3944
R15704 gnd.n5951 gnd.n818 19.3944
R15705 gnd.n5951 gnd.n5950 19.3944
R15706 gnd.n5950 gnd.n5949 19.3944
R15707 gnd.n5847 gnd.n5846 19.3944
R15708 gnd.n5846 gnd.n5845 19.3944
R15709 gnd.n5845 gnd.n1005 19.3944
R15710 gnd.n5841 gnd.n1005 19.3944
R15711 gnd.n5841 gnd.n5840 19.3944
R15712 gnd.n5840 gnd.n5839 19.3944
R15713 gnd.n5839 gnd.n1010 19.3944
R15714 gnd.n5835 gnd.n1010 19.3944
R15715 gnd.n5835 gnd.n5834 19.3944
R15716 gnd.n5834 gnd.n5833 19.3944
R15717 gnd.n5833 gnd.n1015 19.3944
R15718 gnd.n5829 gnd.n1015 19.3944
R15719 gnd.n5829 gnd.n5828 19.3944
R15720 gnd.n5828 gnd.n5827 19.3944
R15721 gnd.n5827 gnd.n1020 19.3944
R15722 gnd.n5823 gnd.n1020 19.3944
R15723 gnd.n5823 gnd.n5822 19.3944
R15724 gnd.n5822 gnd.n5821 19.3944
R15725 gnd.n5821 gnd.n1025 19.3944
R15726 gnd.n5817 gnd.n1025 19.3944
R15727 gnd.n5817 gnd.n5816 19.3944
R15728 gnd.n5816 gnd.n5815 19.3944
R15729 gnd.n5815 gnd.n1030 19.3944
R15730 gnd.n5811 gnd.n1030 19.3944
R15731 gnd.n5811 gnd.n5810 19.3944
R15732 gnd.n5810 gnd.n5809 19.3944
R15733 gnd.n5809 gnd.n1035 19.3944
R15734 gnd.n5805 gnd.n1035 19.3944
R15735 gnd.n5805 gnd.n5804 19.3944
R15736 gnd.n5804 gnd.n5803 19.3944
R15737 gnd.n5803 gnd.n1040 19.3944
R15738 gnd.n5799 gnd.n1040 19.3944
R15739 gnd.n5799 gnd.n5798 19.3944
R15740 gnd.n5798 gnd.n5797 19.3944
R15741 gnd.n5797 gnd.n1045 19.3944
R15742 gnd.n5793 gnd.n1045 19.3944
R15743 gnd.n5793 gnd.n5792 19.3944
R15744 gnd.n5792 gnd.n5791 19.3944
R15745 gnd.n5791 gnd.n1050 19.3944
R15746 gnd.n5787 gnd.n1050 19.3944
R15747 gnd.n5787 gnd.n5786 19.3944
R15748 gnd.n5786 gnd.n5785 19.3944
R15749 gnd.n5785 gnd.n1055 19.3944
R15750 gnd.n5781 gnd.n1055 19.3944
R15751 gnd.n5781 gnd.n5780 19.3944
R15752 gnd.n5780 gnd.n5779 19.3944
R15753 gnd.n5779 gnd.n1060 19.3944
R15754 gnd.n5775 gnd.n1060 19.3944
R15755 gnd.n5775 gnd.n5774 19.3944
R15756 gnd.n5774 gnd.n5773 19.3944
R15757 gnd.n5773 gnd.n1065 19.3944
R15758 gnd.n5769 gnd.n1065 19.3944
R15759 gnd.n5769 gnd.n5768 19.3944
R15760 gnd.n5768 gnd.n5767 19.3944
R15761 gnd.n5767 gnd.n1070 19.3944
R15762 gnd.n5763 gnd.n1070 19.3944
R15763 gnd.n5763 gnd.n5762 19.3944
R15764 gnd.n5762 gnd.n5761 19.3944
R15765 gnd.n5761 gnd.n1075 19.3944
R15766 gnd.n5757 gnd.n1075 19.3944
R15767 gnd.n5757 gnd.n5756 19.3944
R15768 gnd.n5756 gnd.n5755 19.3944
R15769 gnd.n5755 gnd.n1080 19.3944
R15770 gnd.n5751 gnd.n1080 19.3944
R15771 gnd.n5751 gnd.n5750 19.3944
R15772 gnd.n5750 gnd.n5749 19.3944
R15773 gnd.n5749 gnd.n1085 19.3944
R15774 gnd.n5745 gnd.n1085 19.3944
R15775 gnd.n5745 gnd.n5744 19.3944
R15776 gnd.n5744 gnd.n5743 19.3944
R15777 gnd.n5743 gnd.n1090 19.3944
R15778 gnd.n5739 gnd.n1090 19.3944
R15779 gnd.n5739 gnd.n5738 19.3944
R15780 gnd.n5738 gnd.n5737 19.3944
R15781 gnd.n5737 gnd.n1095 19.3944
R15782 gnd.n5733 gnd.n1095 19.3944
R15783 gnd.n5733 gnd.n5732 19.3944
R15784 gnd.n5732 gnd.n5731 19.3944
R15785 gnd.n5731 gnd.n1100 19.3944
R15786 gnd.n5727 gnd.n1100 19.3944
R15787 gnd.n5727 gnd.n5726 19.3944
R15788 gnd.n5726 gnd.n5725 19.3944
R15789 gnd.n5140 gnd.n4975 19.3944
R15790 gnd.n5140 gnd.n4973 19.3944
R15791 gnd.n5145 gnd.n4973 19.3944
R15792 gnd.n5039 gnd.n5021 19.3944
R15793 gnd.n5039 gnd.n5019 19.3944
R15794 gnd.n5045 gnd.n5019 19.3944
R15795 gnd.n5045 gnd.n5012 19.3944
R15796 gnd.n5058 gnd.n5012 19.3944
R15797 gnd.n5058 gnd.n5010 19.3944
R15798 gnd.n5064 gnd.n5010 19.3944
R15799 gnd.n5064 gnd.n5003 19.3944
R15800 gnd.n5077 gnd.n5003 19.3944
R15801 gnd.n5077 gnd.n5001 19.3944
R15802 gnd.n5083 gnd.n5001 19.3944
R15803 gnd.n5083 gnd.n4994 19.3944
R15804 gnd.n5096 gnd.n4994 19.3944
R15805 gnd.n5096 gnd.n4992 19.3944
R15806 gnd.n5104 gnd.n4992 19.3944
R15807 gnd.n5104 gnd.n5103 19.3944
R15808 gnd.n5103 gnd.n4983 19.3944
R15809 gnd.n5117 gnd.n4983 19.3944
R15810 gnd.n5117 gnd.n4981 19.3944
R15811 gnd.n5123 gnd.n4981 19.3944
R15812 gnd.n5123 gnd.n4979 19.3944
R15813 gnd.n5127 gnd.n4979 19.3944
R15814 gnd.n5127 gnd.n4977 19.3944
R15815 gnd.n5136 gnd.n4977 19.3944
R15816 gnd.n2941 gnd.t21 18.8012
R15817 gnd.n2926 gnd.t251 18.8012
R15818 gnd.n2785 gnd.n2784 18.4825
R15819 gnd.n5410 gnd.n1291 18.4247
R15820 gnd.n4346 gnd.n1808 18.4247
R15821 gnd.n6883 gnd.n6882 18.2308
R15822 gnd.n5107 gnd.n4987 18.2308
R15823 gnd.n4149 gnd.n4133 18.2308
R15824 gnd.n3630 gnd.n3586 18.2308
R15825 gnd.t23 gnd.n2465 18.1639
R15826 gnd.n2493 gnd.t24 17.5266
R15827 gnd.n2892 gnd.t18 16.8893
R15828 gnd.n3803 gnd.t220 16.8893
R15829 gnd.n4301 gnd.t157 16.8893
R15830 gnd.n5468 gnd.t150 16.8893
R15831 gnd.t143 gnd.n81 16.8893
R15832 gnd.n2720 gnd.t236 16.2519
R15833 gnd.n2420 gnd.t12 16.2519
R15834 gnd.n4190 gnd.n4189 15.9333
R15835 gnd.n4189 gnd.n1964 15.9333
R15836 gnd.n4199 gnd.n4198 15.9333
R15837 gnd.n4200 gnd.n4199 15.9333
R15838 gnd.n4201 gnd.n4200 15.9333
R15839 gnd.n4204 gnd.n4201 15.9333
R15840 gnd.n4203 gnd.n4202 15.9333
R15841 gnd.n4202 gnd.n1958 15.9333
R15842 gnd.n4212 gnd.n1958 15.9333
R15843 gnd.n4213 gnd.n4212 15.9333
R15844 gnd.n4214 gnd.n4213 15.9333
R15845 gnd.n4215 gnd.n4214 15.9333
R15846 gnd.n4218 gnd.n4215 15.9333
R15847 gnd.n4218 gnd.n4217 15.9333
R15848 gnd.n4216 gnd.n1950 15.9333
R15849 gnd.n4226 gnd.n1950 15.9333
R15850 gnd.n4227 gnd.n4226 15.9333
R15851 gnd.n4228 gnd.n4227 15.9333
R15852 gnd.n4229 gnd.n4228 15.9333
R15853 gnd.n4232 gnd.n4229 15.9333
R15854 gnd.n4232 gnd.n4231 15.9333
R15855 gnd.n4231 gnd.n4230 15.9333
R15856 gnd.n4242 gnd.n4240 15.9333
R15857 gnd.n4240 gnd.n1700 15.9333
R15858 gnd.n4245 gnd.n1733 15.9333
R15859 gnd.n4421 gnd.n4420 15.9333
R15860 gnd.n4429 gnd.n1665 15.9333
R15861 gnd.n4477 gnd.n1653 15.9333
R15862 gnd.n4487 gnd.n4485 15.9333
R15863 gnd.n4520 gnd.n4518 15.9333
R15864 gnd.n4565 gnd.n1599 15.9333
R15865 gnd.n4593 gnd.n1584 15.9333
R15866 gnd.n4612 gnd.n1572 15.9333
R15867 gnd.n4612 gnd.n1573 15.9333
R15868 gnd.n1556 gnd.n1544 15.9333
R15869 gnd.n4671 gnd.n1527 15.9333
R15870 gnd.n4716 gnd.n4715 15.9333
R15871 gnd.n4724 gnd.n1514 15.9333
R15872 gnd.n4800 gnd.n1479 15.9333
R15873 gnd.n4800 gnd.n1481 15.9333
R15874 gnd.n4810 gnd.n4808 15.9333
R15875 gnd.n4841 gnd.n4839 15.9333
R15876 gnd.n4884 gnd.n4883 15.9333
R15877 gnd.n4910 gnd.n4909 15.9333
R15878 gnd.n4921 gnd.n1404 15.9333
R15879 gnd.n1335 gnd.n1296 15.9333
R15880 gnd.n5184 gnd.n5183 15.9333
R15881 gnd.n5181 gnd.n5180 15.9333
R15882 gnd.n5180 gnd.n5179 15.9333
R15883 gnd.n5179 gnd.n1354 15.9333
R15884 gnd.n1364 gnd.n1354 15.9333
R15885 gnd.n1365 gnd.n1364 15.9333
R15886 gnd.n5173 gnd.n1365 15.9333
R15887 gnd.n5173 gnd.n5172 15.9333
R15888 gnd.n5172 gnd.n5170 15.9333
R15889 gnd.n5169 gnd.n5168 15.9333
R15890 gnd.n5168 gnd.n1368 15.9333
R15891 gnd.n1376 gnd.n1368 15.9333
R15892 gnd.n1377 gnd.n1376 15.9333
R15893 gnd.n5162 gnd.n1377 15.9333
R15894 gnd.n5162 gnd.n5161 15.9333
R15895 gnd.n5161 gnd.n5159 15.9333
R15896 gnd.n5159 gnd.n5158 15.9333
R15897 gnd.n5157 gnd.n5151 15.9333
R15898 gnd.n5151 gnd.n1106 15.9333
R15899 gnd.n5723 gnd.n1106 15.9333
R15900 gnd.n5723 gnd.n5722 15.9333
R15901 gnd.n1117 gnd.n1108 15.9333
R15902 gnd.n5716 gnd.n1117 15.9333
R15903 gnd.n3408 gnd.n3406 15.6674
R15904 gnd.n3376 gnd.n3374 15.6674
R15905 gnd.n3344 gnd.n3342 15.6674
R15906 gnd.n3313 gnd.n3311 15.6674
R15907 gnd.n3281 gnd.n3279 15.6674
R15908 gnd.n3249 gnd.n3247 15.6674
R15909 gnd.n3217 gnd.n3215 15.6674
R15910 gnd.n3186 gnd.n3184 15.6674
R15911 gnd.n2711 gnd.t236 15.6146
R15912 gnd.t172 gnd.n2186 15.6146
R15913 gnd.t168 gnd.n2187 15.6146
R15914 gnd.t201 gnd.n4203 15.6146
R15915 gnd.n5158 gnd.t182 15.6146
R15916 gnd.n4448 gnd.n1625 15.296
R15917 gnd.n4537 gnd.n1612 15.296
R15918 gnd.n4672 gnd.n4670 15.296
R15919 gnd.n4714 gnd.n1523 15.296
R15920 gnd.n4780 gnd.n1445 15.296
R15921 gnd.n4881 gnd.n1432 15.296
R15922 gnd.n5200 gnd.n5199 15.0827
R15923 gnd.n1686 gnd.n1681 15.0481
R15924 gnd.n5210 gnd.n5209 15.0481
R15925 gnd.n3080 gnd.t25 14.9773
R15926 gnd.t220 gnd.n2087 14.9773
R15927 gnd.n4230 gnd.t64 14.9773
R15928 gnd.t101 gnd.n5181 14.9773
R15929 gnd.n6926 gnd.t143 14.9773
R15930 gnd.n4476 gnd.n1655 14.6587
R15931 gnd.n4495 gnd.t105 14.6587
R15932 gnd.n4584 gnd.n4583 14.6587
R15933 gnd.n4605 gnd.n4604 14.6587
R15934 gnd.n4752 gnd.n4750 14.6587
R15935 gnd.n1473 gnd.n1462 14.6587
R15936 gnd.n4857 gnd.t247 14.6587
R15937 gnd.n4923 gnd.n4922 14.6587
R15938 gnd.n5282 gnd.n1335 14.6587
R15939 gnd.n5184 gnd.t217 14.6587
R15940 gnd.t49 gnd.n2229 14.34
R15941 gnd.n3158 gnd.t22 14.34
R15942 gnd.n4497 gnd.n4496 14.0214
R15943 gnd.n4563 gnd.n1601 14.0214
R15944 gnd.n4662 gnd.n4661 14.0214
R15945 gnd.n1513 gnd.n1506 14.0214
R15946 gnd.n4842 gnd.n1449 14.0214
R15947 gnd.n4856 gnd.n1417 14.0214
R15948 gnd.n2867 gnd.t115 13.7027
R15949 gnd.n1577 gnd.t90 13.7027
R15950 gnd.n4749 gnd.t278 13.7027
R15951 gnd.n2577 gnd.n2576 13.5763
R15952 gnd.n3522 gnd.n2143 13.5763
R15953 gnd.n1271 gnd.n1270 13.5763
R15954 gnd.n6935 gnd.n6934 13.5763
R15955 gnd.n3712 gnd.n3687 13.5763
R15956 gnd.n4312 gnd.n1900 13.5763
R15957 gnd.n2785 gnd.n2523 13.384
R15958 gnd.n4557 gnd.n1605 13.384
R15959 gnd.n4652 gnd.n4651 13.384
R15960 gnd.n1507 gnd.n1501 13.384
R15961 gnd.n4828 gnd.n1458 13.384
R15962 gnd.n4859 gnd.n1412 13.384
R15963 gnd.n1697 gnd.n1678 13.1884
R15964 gnd.n1692 gnd.n1691 13.1884
R15965 gnd.n1691 gnd.n1690 13.1884
R15966 gnd.n5203 gnd.n5198 13.1884
R15967 gnd.n5204 gnd.n5203 13.1884
R15968 gnd.n1693 gnd.n1680 13.146
R15969 gnd.n1689 gnd.n1680 13.146
R15970 gnd.n5202 gnd.n5201 13.146
R15971 gnd.n5202 gnd.n5197 13.146
R15972 gnd.t276 gnd.n1660 13.0654
R15973 gnd.n4940 gnd.t62 13.0654
R15974 gnd.n3409 gnd.n3405 12.8005
R15975 gnd.n3377 gnd.n3373 12.8005
R15976 gnd.n3345 gnd.n3341 12.8005
R15977 gnd.n3314 gnd.n3310 12.8005
R15978 gnd.n3282 gnd.n3278 12.8005
R15979 gnd.n3250 gnd.n3246 12.8005
R15980 gnd.n3218 gnd.n3214 12.8005
R15981 gnd.n3187 gnd.n3183 12.8005
R15982 gnd.n4458 gnd.n1645 12.7467
R15983 gnd.n4632 gnd.n4630 12.7467
R15984 gnd.n4739 gnd.n1493 12.7467
R15985 gnd.n5947 gnd.n827 12.4281
R15986 gnd.n4410 gnd.n1733 12.4281
R15987 gnd.n5349 gnd.n1296 12.4281
R15988 gnd.n6918 gnd.n168 12.4281
R15989 gnd.n2576 gnd.n2571 12.4126
R15990 gnd.n3525 gnd.n3522 12.4126
R15991 gnd.n5462 gnd.n1270 12.4126
R15992 gnd.n6934 gnd.n155 12.4126
R15993 gnd.n3708 gnd.n3687 12.4126
R15994 gnd.n4307 gnd.n1900 12.4126
R15995 gnd.n4414 gnd.n4413 12.1761
R15996 gnd.n5279 gnd.n5278 12.1761
R15997 gnd.n4507 gnd.n1633 12.1094
R15998 gnd.t250 gnd.n1614 12.1094
R15999 gnd.n4849 gnd.t242 12.1094
R16000 gnd.n4893 gnd.n1422 12.1094
R16001 gnd.n4948 gnd.t147 12.1094
R16002 gnd.n3413 gnd.n3412 12.0247
R16003 gnd.n3381 gnd.n3380 12.0247
R16004 gnd.n3349 gnd.n3348 12.0247
R16005 gnd.n3318 gnd.n3317 12.0247
R16006 gnd.n3286 gnd.n3285 12.0247
R16007 gnd.n3254 gnd.n3253 12.0247
R16008 gnd.n3222 gnd.n3221 12.0247
R16009 gnd.n3191 gnd.n3190 12.0247
R16010 gnd.n5872 gnd.t45 11.7908
R16011 gnd.n5554 gnd.t93 11.7908
R16012 gnd.n4055 gnd.n1870 11.4721
R16013 gnd.t136 gnd.n1671 11.4721
R16014 gnd.n4419 gnd.n1674 11.4721
R16015 gnd.n5191 gnd.n1343 11.4721
R16016 gnd.n5714 gnd.n1118 11.4721
R16017 gnd.n3416 gnd.n3403 11.249
R16018 gnd.n3384 gnd.n3371 11.249
R16019 gnd.n3352 gnd.n3339 11.249
R16020 gnd.n3321 gnd.n3308 11.249
R16021 gnd.n3289 gnd.n3276 11.249
R16022 gnd.n3257 gnd.n3244 11.249
R16023 gnd.n3225 gnd.n3212 11.249
R16024 gnd.n3194 gnd.n3181 11.249
R16025 gnd.n2855 gnd.t115 11.1535
R16026 gnd.t0 gnd.n865 11.1535
R16027 gnd.n5896 gnd.t2 11.1535
R16028 gnd.n4217 gnd.t269 11.1535
R16029 gnd.n4576 gnd.t98 11.1535
R16030 gnd.t264 gnd.n4820 11.1535
R16031 gnd.t41 gnd.n5169 11.1535
R16032 gnd.n5613 gnd.t36 11.1535
R16033 gnd.n6762 gnd.t27 11.1535
R16034 gnd.n840 gnd.n830 10.8348
R16035 gnd.n5940 gnd.n843 10.8348
R16036 gnd.n3825 gnd.n852 10.8348
R16037 gnd.n3845 gnd.n862 10.8348
R16038 gnd.n5928 gnd.n865 10.8348
R16039 gnd.n3839 gnd.n873 10.8348
R16040 gnd.n5922 gnd.n876 10.8348
R16041 gnd.n3873 gnd.n3872 10.8348
R16042 gnd.n5916 gnd.n886 10.8348
R16043 gnd.n3883 gnd.n894 10.8348
R16044 gnd.n3893 gnd.n2055 10.8348
R16045 gnd.n3920 gnd.n3909 10.8348
R16046 gnd.n3917 gnd.n2049 10.8348
R16047 gnd.n3928 gnd.n2028 10.8348
R16048 gnd.n3948 gnd.n2023 10.8348
R16049 gnd.n3957 gnd.n2014 10.8348
R16050 gnd.n3956 gnd.n909 10.8348
R16051 gnd.n5902 gnd.n912 10.8348
R16052 gnd.n3969 gnd.n3968 10.8348
R16053 gnd.n5896 gnd.n923 10.8348
R16054 gnd.n3977 gnd.n930 10.8348
R16055 gnd.n4022 gnd.n940 10.8348
R16056 gnd.n5884 gnd.n943 10.8348
R16057 gnd.n3985 gnd.n951 10.8348
R16058 gnd.n5878 gnd.n954 10.8348
R16059 gnd.n3992 gnd.n3991 10.8348
R16060 gnd.n5872 gnd.n964 10.8348
R16061 gnd.n3996 gnd.n972 10.8348
R16062 gnd.n5866 gnd.n975 10.8348
R16063 gnd.n4005 gnd.n983 10.8348
R16064 gnd.n5860 gnd.n986 10.8348
R16065 gnd.n4301 gnd.n993 10.8348
R16066 gnd.n5854 gnd.n996 10.8348
R16067 gnd.n4530 gnd.n1618 10.8348
R16068 gnd.n4556 gnd.t253 10.8348
R16069 gnd.n4708 gnd.n4707 10.8348
R16070 gnd.n4707 gnd.n1520 10.8348
R16071 gnd.n4829 gnd.t76 10.8348
R16072 gnd.n4875 gnd.n4874 10.8348
R16073 gnd.n5708 gnd.n5707 10.8348
R16074 gnd.n5468 gnd.n1129 10.8348
R16075 gnd.n5701 gnd.n1138 10.8348
R16076 gnd.n5477 gnd.n1141 10.8348
R16077 gnd.n5544 gnd.n1256 10.8348
R16078 gnd.n5543 gnd.n5526 10.8348
R16079 gnd.n5554 gnd.n1249 10.8348
R16080 gnd.n1251 gnd.n1241 10.8348
R16081 gnd.n5564 gnd.n5563 10.8348
R16082 gnd.n5575 gnd.n1230 10.8348
R16083 gnd.n5574 gnd.n1233 10.8348
R16084 gnd.n5586 gnd.n1220 10.8348
R16085 gnd.n5596 gnd.n5595 10.8348
R16086 gnd.n5613 gnd.n1201 10.8348
R16087 gnd.n5612 gnd.n1205 10.8348
R16088 gnd.n5619 gnd.n1194 10.8348
R16089 gnd.n5506 gnd.n1196 10.8348
R16090 gnd.n5629 gnd.n1184 10.8348
R16091 gnd.n5628 gnd.n1176 10.8348
R16092 gnd.n1180 gnd.n1170 10.8348
R16093 gnd.n5666 gnd.n5665 10.8348
R16094 gnd.n6783 gnd.n235 10.8348
R16095 gnd.n6788 gnd.n231 10.8348
R16096 gnd.n6796 gnd.n223 10.8348
R16097 gnd.n6772 gnd.n225 10.8348
R16098 gnd.n6804 gnd.n209 10.8348
R16099 gnd.n6768 gnd.n211 10.8348
R16100 gnd.n6812 gnd.n202 10.8348
R16101 gnd.n6763 gnd.n6762 10.8348
R16102 gnd.n6820 gnd.n194 10.8348
R16103 gnd.n6828 gnd.n186 10.8348
R16104 gnd.n261 gnd.n188 10.8348
R16105 gnd.n6836 gnd.n177 10.8348
R16106 gnd.n5344 gnd.n1292 10.6151
R16107 gnd.n5344 gnd.n5343 10.6151
R16108 gnd.n5341 gnd.n5338 10.6151
R16109 gnd.n5338 gnd.n5337 10.6151
R16110 gnd.n5337 gnd.n5334 10.6151
R16111 gnd.n5334 gnd.n5333 10.6151
R16112 gnd.n5333 gnd.n5330 10.6151
R16113 gnd.n5330 gnd.n5329 10.6151
R16114 gnd.n5329 gnd.n5326 10.6151
R16115 gnd.n5326 gnd.n5325 10.6151
R16116 gnd.n5325 gnd.n5322 10.6151
R16117 gnd.n5322 gnd.n5321 10.6151
R16118 gnd.n5321 gnd.n5318 10.6151
R16119 gnd.n5318 gnd.n5317 10.6151
R16120 gnd.n5317 gnd.n5314 10.6151
R16121 gnd.n5314 gnd.n5313 10.6151
R16122 gnd.n5313 gnd.n5310 10.6151
R16123 gnd.n5310 gnd.n5309 10.6151
R16124 gnd.n5309 gnd.n5306 10.6151
R16125 gnd.n5306 gnd.n5305 10.6151
R16126 gnd.n5305 gnd.n5302 10.6151
R16127 gnd.n5302 gnd.n5301 10.6151
R16128 gnd.n5301 gnd.n5298 10.6151
R16129 gnd.n5298 gnd.n5297 10.6151
R16130 gnd.n5297 gnd.n5294 10.6151
R16131 gnd.n5294 gnd.n5293 10.6151
R16132 gnd.n5293 gnd.n5290 10.6151
R16133 gnd.n5290 gnd.n5289 10.6151
R16134 gnd.n5289 gnd.n5286 10.6151
R16135 gnd.n5286 gnd.n5285 10.6151
R16136 gnd.n1741 gnd.n1740 10.6151
R16137 gnd.n1740 gnd.n1662 10.6151
R16138 gnd.n4431 gnd.n1662 10.6151
R16139 gnd.n4432 gnd.n4431 10.6151
R16140 gnd.n4463 gnd.n4432 10.6151
R16141 gnd.n4463 gnd.n4462 10.6151
R16142 gnd.n4462 gnd.n4461 10.6151
R16143 gnd.n4461 gnd.n4433 10.6151
R16144 gnd.n4455 gnd.n4433 10.6151
R16145 gnd.n4455 gnd.n4454 10.6151
R16146 gnd.n4454 gnd.n4453 10.6151
R16147 gnd.n4453 gnd.n4452 10.6151
R16148 gnd.n4452 gnd.n4451 10.6151
R16149 gnd.n4451 gnd.n4434 10.6151
R16150 gnd.n4445 gnd.n4434 10.6151
R16151 gnd.n4445 gnd.n4444 10.6151
R16152 gnd.n4444 gnd.n4443 10.6151
R16153 gnd.n4443 gnd.n4441 10.6151
R16154 gnd.n4441 gnd.n4440 10.6151
R16155 gnd.n4440 gnd.n4438 10.6151
R16156 gnd.n4438 gnd.n4437 10.6151
R16157 gnd.n4437 gnd.n1591 10.6151
R16158 gnd.n4578 gnd.n1591 10.6151
R16159 gnd.n4579 gnd.n4578 10.6151
R16160 gnd.n4581 gnd.n4579 10.6151
R16161 gnd.n4581 gnd.n4580 10.6151
R16162 gnd.n4580 gnd.n1576 10.6151
R16163 gnd.n4610 gnd.n1576 10.6151
R16164 gnd.n4610 gnd.n4609 10.6151
R16165 gnd.n4609 gnd.n4608 10.6151
R16166 gnd.n4608 gnd.n4607 10.6151
R16167 gnd.n4607 gnd.n1557 10.6151
R16168 gnd.n4634 gnd.n1557 10.6151
R16169 gnd.n4635 gnd.n4634 10.6151
R16170 gnd.n4637 gnd.n4635 10.6151
R16171 gnd.n4638 gnd.n4637 10.6151
R16172 gnd.n4639 gnd.n4638 10.6151
R16173 gnd.n4639 gnd.n1534 10.6151
R16174 gnd.n4674 gnd.n1534 10.6151
R16175 gnd.n4675 gnd.n4674 10.6151
R16176 gnd.n4677 gnd.n4675 10.6151
R16177 gnd.n4678 gnd.n4677 10.6151
R16178 gnd.n4680 gnd.n4678 10.6151
R16179 gnd.n4680 gnd.n4679 10.6151
R16180 gnd.n4679 gnd.n1504 10.6151
R16181 gnd.n4734 gnd.n1504 10.6151
R16182 gnd.n4735 gnd.n4734 10.6151
R16183 gnd.n4737 gnd.n4735 10.6151
R16184 gnd.n4737 gnd.n4736 10.6151
R16185 gnd.n4736 gnd.n1484 10.6151
R16186 gnd.n4769 gnd.n1484 10.6151
R16187 gnd.n4770 gnd.n4769 10.6151
R16188 gnd.n4798 gnd.n4770 10.6151
R16189 gnd.n4798 gnd.n4797 10.6151
R16190 gnd.n4797 gnd.n4796 10.6151
R16191 gnd.n4796 gnd.n4793 10.6151
R16192 gnd.n4793 gnd.n4792 10.6151
R16193 gnd.n4792 gnd.n4791 10.6151
R16194 gnd.n4791 gnd.n4790 10.6151
R16195 gnd.n4790 gnd.n4789 10.6151
R16196 gnd.n4789 gnd.n4786 10.6151
R16197 gnd.n4786 gnd.n4785 10.6151
R16198 gnd.n4785 gnd.n4783 10.6151
R16199 gnd.n4783 gnd.n4782 10.6151
R16200 gnd.n4782 gnd.n4778 10.6151
R16201 gnd.n4778 gnd.n4777 10.6151
R16202 gnd.n4777 gnd.n4775 10.6151
R16203 gnd.n4775 gnd.n4774 10.6151
R16204 gnd.n4774 gnd.n4771 10.6151
R16205 gnd.n4771 gnd.n1415 10.6151
R16206 gnd.n4902 gnd.n1415 10.6151
R16207 gnd.n4903 gnd.n4902 10.6151
R16208 gnd.n4905 gnd.n4903 10.6151
R16209 gnd.n4905 gnd.n4904 10.6151
R16210 gnd.n4904 gnd.n1395 10.6151
R16211 gnd.n4933 gnd.n1395 10.6151
R16212 gnd.n4934 gnd.n4933 10.6151
R16213 gnd.n4937 gnd.n4934 10.6151
R16214 gnd.n4937 gnd.n4936 10.6151
R16215 gnd.n4936 gnd.n4935 10.6151
R16216 gnd.n4935 gnd.n1332 10.6151
R16217 gnd.n1806 gnd.n1805 10.6151
R16218 gnd.n1805 gnd.n1802 10.6151
R16219 gnd.n1800 gnd.n1797 10.6151
R16220 gnd.n1797 gnd.n1796 10.6151
R16221 gnd.n1796 gnd.n1793 10.6151
R16222 gnd.n1793 gnd.n1792 10.6151
R16223 gnd.n1792 gnd.n1789 10.6151
R16224 gnd.n1789 gnd.n1788 10.6151
R16225 gnd.n1788 gnd.n1785 10.6151
R16226 gnd.n1785 gnd.n1784 10.6151
R16227 gnd.n1784 gnd.n1781 10.6151
R16228 gnd.n1781 gnd.n1780 10.6151
R16229 gnd.n1780 gnd.n1777 10.6151
R16230 gnd.n1777 gnd.n1776 10.6151
R16231 gnd.n1776 gnd.n1773 10.6151
R16232 gnd.n1773 gnd.n1772 10.6151
R16233 gnd.n1772 gnd.n1769 10.6151
R16234 gnd.n1769 gnd.n1768 10.6151
R16235 gnd.n1768 gnd.n1765 10.6151
R16236 gnd.n1765 gnd.n1764 10.6151
R16237 gnd.n1764 gnd.n1761 10.6151
R16238 gnd.n1761 gnd.n1760 10.6151
R16239 gnd.n1760 gnd.n1757 10.6151
R16240 gnd.n1757 gnd.n1756 10.6151
R16241 gnd.n1756 gnd.n1753 10.6151
R16242 gnd.n1753 gnd.n1752 10.6151
R16243 gnd.n1752 gnd.n1749 10.6151
R16244 gnd.n1749 gnd.n1748 10.6151
R16245 gnd.n1748 gnd.n1745 10.6151
R16246 gnd.n1745 gnd.n1744 10.6151
R16247 gnd.n4413 gnd.n1698 10.6151
R16248 gnd.n4408 gnd.n1698 10.6151
R16249 gnd.n4408 gnd.n4407 10.6151
R16250 gnd.n4407 gnd.n4406 10.6151
R16251 gnd.n4406 gnd.n4403 10.6151
R16252 gnd.n4403 gnd.n4402 10.6151
R16253 gnd.n4402 gnd.n4399 10.6151
R16254 gnd.n4399 gnd.n4398 10.6151
R16255 gnd.n4398 gnd.n4395 10.6151
R16256 gnd.n4395 gnd.n4394 10.6151
R16257 gnd.n4394 gnd.n4391 10.6151
R16258 gnd.n4391 gnd.n4390 10.6151
R16259 gnd.n4390 gnd.n4387 10.6151
R16260 gnd.n4387 gnd.n4386 10.6151
R16261 gnd.n4386 gnd.n4383 10.6151
R16262 gnd.n4383 gnd.n4382 10.6151
R16263 gnd.n4382 gnd.n4379 10.6151
R16264 gnd.n4379 gnd.n4378 10.6151
R16265 gnd.n4378 gnd.n4375 10.6151
R16266 gnd.n4375 gnd.n4374 10.6151
R16267 gnd.n4374 gnd.n4371 10.6151
R16268 gnd.n4371 gnd.n4370 10.6151
R16269 gnd.n4370 gnd.n4367 10.6151
R16270 gnd.n4367 gnd.n4366 10.6151
R16271 gnd.n4366 gnd.n4363 10.6151
R16272 gnd.n4363 gnd.n4362 10.6151
R16273 gnd.n4362 gnd.n4359 10.6151
R16274 gnd.n4359 gnd.n4358 10.6151
R16275 gnd.n4355 gnd.n4354 10.6151
R16276 gnd.n4354 gnd.n4351 10.6151
R16277 gnd.n5278 gnd.n5277 10.6151
R16278 gnd.n5277 gnd.n5274 10.6151
R16279 gnd.n5274 gnd.n5273 10.6151
R16280 gnd.n5273 gnd.n5270 10.6151
R16281 gnd.n5270 gnd.n5269 10.6151
R16282 gnd.n5269 gnd.n5266 10.6151
R16283 gnd.n5266 gnd.n5265 10.6151
R16284 gnd.n5265 gnd.n5262 10.6151
R16285 gnd.n5262 gnd.n5261 10.6151
R16286 gnd.n5261 gnd.n5258 10.6151
R16287 gnd.n5258 gnd.n5257 10.6151
R16288 gnd.n5257 gnd.n5254 10.6151
R16289 gnd.n5254 gnd.n5253 10.6151
R16290 gnd.n5253 gnd.n5250 10.6151
R16291 gnd.n5250 gnd.n5249 10.6151
R16292 gnd.n5249 gnd.n5246 10.6151
R16293 gnd.n5246 gnd.n5245 10.6151
R16294 gnd.n5245 gnd.n5242 10.6151
R16295 gnd.n5242 gnd.n5241 10.6151
R16296 gnd.n5241 gnd.n5238 10.6151
R16297 gnd.n5238 gnd.n5237 10.6151
R16298 gnd.n5237 gnd.n5234 10.6151
R16299 gnd.n5234 gnd.n5233 10.6151
R16300 gnd.n5233 gnd.n5230 10.6151
R16301 gnd.n5230 gnd.n5229 10.6151
R16302 gnd.n5229 gnd.n5226 10.6151
R16303 gnd.n5226 gnd.n5225 10.6151
R16304 gnd.n5225 gnd.n5222 10.6151
R16305 gnd.n5220 gnd.n5217 10.6151
R16306 gnd.n5217 gnd.n1293 10.6151
R16307 gnd.n4417 gnd.n4415 10.6151
R16308 gnd.n4417 gnd.n4416 10.6151
R16309 gnd.n4416 gnd.n1658 10.6151
R16310 gnd.n4469 gnd.n1658 10.6151
R16311 gnd.n4470 gnd.n4469 10.6151
R16312 gnd.n4474 gnd.n4470 10.6151
R16313 gnd.n4474 gnd.n4473 10.6151
R16314 gnd.n4473 gnd.n4472 10.6151
R16315 gnd.n4472 gnd.n1636 10.6151
R16316 gnd.n4500 gnd.n1636 10.6151
R16317 gnd.n4501 gnd.n4500 10.6151
R16318 gnd.n4505 gnd.n4501 10.6151
R16319 gnd.n4505 gnd.n4504 10.6151
R16320 gnd.n4504 gnd.n4503 10.6151
R16321 gnd.n4503 gnd.n1616 10.6151
R16322 gnd.n4532 gnd.n1616 10.6151
R16323 gnd.n4533 gnd.n4532 10.6151
R16324 gnd.n4534 gnd.n4533 10.6151
R16325 gnd.n4534 gnd.n1604 10.6151
R16326 gnd.n4561 gnd.n1604 10.6151
R16327 gnd.n4561 gnd.n4560 10.6151
R16328 gnd.n4560 gnd.n4559 10.6151
R16329 gnd.n4559 gnd.n1587 10.6151
R16330 gnd.n4587 gnd.n1587 10.6151
R16331 gnd.n4588 gnd.n4587 10.6151
R16332 gnd.n4589 gnd.n4588 10.6151
R16333 gnd.n4589 gnd.n1570 10.6151
R16334 gnd.n4614 gnd.n1570 10.6151
R16335 gnd.n4615 gnd.n4614 10.6151
R16336 gnd.n4619 gnd.n4615 10.6151
R16337 gnd.n4619 gnd.n4618 10.6151
R16338 gnd.n4618 gnd.n4617 10.6151
R16339 gnd.n4617 gnd.n1547 10.6151
R16340 gnd.n4654 gnd.n1547 10.6151
R16341 gnd.n4655 gnd.n4654 10.6151
R16342 gnd.n4659 gnd.n4655 10.6151
R16343 gnd.n4659 gnd.n4658 10.6151
R16344 gnd.n4658 gnd.n4657 10.6151
R16345 gnd.n4657 gnd.n1525 10.6151
R16346 gnd.n4710 gnd.n1525 10.6151
R16347 gnd.n4711 gnd.n4710 10.6151
R16348 gnd.n4712 gnd.n4711 10.6151
R16349 gnd.n4712 gnd.n1510 10.6151
R16350 gnd.n4727 gnd.n1510 10.6151
R16351 gnd.n4728 gnd.n4727 10.6151
R16352 gnd.n4730 gnd.n4728 10.6151
R16353 gnd.n4730 gnd.n4729 10.6151
R16354 gnd.n4729 gnd.n1491 10.6151
R16355 gnd.n4755 gnd.n1491 10.6151
R16356 gnd.n4756 gnd.n4755 10.6151
R16357 gnd.n4765 gnd.n4756 10.6151
R16358 gnd.n4765 gnd.n4764 10.6151
R16359 gnd.n4764 gnd.n4763 10.6151
R16360 gnd.n4763 gnd.n4762 10.6151
R16361 gnd.n4762 gnd.n4757 10.6151
R16362 gnd.n4757 gnd.n1460 10.6151
R16363 gnd.n4824 gnd.n1460 10.6151
R16364 gnd.n4825 gnd.n4824 10.6151
R16365 gnd.n4826 gnd.n4825 10.6151
R16366 gnd.n4826 gnd.n1447 10.6151
R16367 gnd.n4844 gnd.n1447 10.6151
R16368 gnd.n4845 gnd.n4844 10.6151
R16369 gnd.n4846 gnd.n4845 10.6151
R16370 gnd.n4846 gnd.n1434 10.6151
R16371 gnd.n4877 gnd.n1434 10.6151
R16372 gnd.n4878 gnd.n4877 10.6151
R16373 gnd.n4879 gnd.n4878 10.6151
R16374 gnd.n4879 gnd.n1420 10.6151
R16375 gnd.n4895 gnd.n1420 10.6151
R16376 gnd.n4896 gnd.n4895 10.6151
R16377 gnd.n4898 gnd.n4896 10.6151
R16378 gnd.n4898 gnd.n4897 10.6151
R16379 gnd.n4897 gnd.n1399 10.6151
R16380 gnd.n4926 gnd.n1399 10.6151
R16381 gnd.n4927 gnd.n4926 10.6151
R16382 gnd.n4929 gnd.n4927 10.6151
R16383 gnd.n4929 gnd.n4928 10.6151
R16384 gnd.n4928 gnd.n1338 10.6151
R16385 gnd.n5194 gnd.n1338 10.6151
R16386 gnd.n5195 gnd.n5194 10.6151
R16387 gnd.n5280 gnd.n5195 10.6151
R16388 gnd.n2774 gnd.t117 10.5161
R16389 gnd.n2231 gnd.t49 10.5161
R16390 gnd.n3141 gnd.t22 10.5161
R16391 gnd.n3894 gnd.t6 10.5161
R16392 gnd.t29 gnd.n3909 10.5161
R16393 gnd.n3917 gnd.t29 10.5161
R16394 gnd.n3942 gnd.t34 10.5161
R16395 gnd.n4529 gnd.t119 10.5161
R16396 gnd.t103 gnd.n1436 10.5161
R16397 gnd.t72 gnd.n5638 10.5161
R16398 gnd.n5666 gnd.t4 10.5161
R16399 gnd.t4 gnd.n235 10.5161
R16400 gnd.t32 gnd.n233 10.5161
R16401 gnd.n3417 gnd.n3401 10.4732
R16402 gnd.n3385 gnd.n3369 10.4732
R16403 gnd.n3353 gnd.n3337 10.4732
R16404 gnd.n3322 gnd.n3306 10.4732
R16405 gnd.n3290 gnd.n3274 10.4732
R16406 gnd.n3258 gnd.n3242 10.4732
R16407 gnd.n3226 gnd.n3210 10.4732
R16408 gnd.n3195 gnd.n3179 10.4732
R16409 gnd.n4466 gnd.t139 10.1975
R16410 gnd.n4549 gnd.n4548 10.1975
R16411 gnd.n4622 gnd.n1565 10.1975
R16412 gnd.n1489 gnd.n1488 10.1975
R16413 gnd.n4760 gnd.n4759 10.1975
R16414 gnd.n1406 gnd.t161 10.1975
R16415 gnd.n1406 gnd.n1393 10.1975
R16416 gnd.n5192 gnd.n5191 10.1975
R16417 gnd.n3846 gnd.t47 9.87883
R16418 gnd.n3839 gnd.t0 9.87883
R16419 gnd.n3968 gnd.t2 9.87883
R16420 gnd.n5890 gnd.t8 9.87883
R16421 gnd.n4643 gnd.t112 9.87883
R16422 gnd.n4684 gnd.t96 9.87883
R16423 gnd.t57 gnd.n1212 9.87883
R16424 gnd.t36 gnd.n5612 9.87883
R16425 gnd.n6812 gnd.t27 9.87883
R16426 gnd.t51 gnd.n196 9.87883
R16427 gnd.n3421 gnd.n3420 9.69747
R16428 gnd.n3389 gnd.n3388 9.69747
R16429 gnd.n3357 gnd.n3356 9.69747
R16430 gnd.n3326 gnd.n3325 9.69747
R16431 gnd.n3294 gnd.n3293 9.69747
R16432 gnd.n3262 gnd.n3261 9.69747
R16433 gnd.n3230 gnd.n3229 9.69747
R16434 gnd.n3199 gnd.n3198 9.69747
R16435 gnd.n7041 gnd.n50 9.6512
R16436 gnd.n4449 gnd.n1633 9.56018
R16437 gnd.n4536 gnd.n1614 9.56018
R16438 gnd.n4643 gnd.n1536 9.56018
R16439 gnd.n4684 gnd.n4682 9.56018
R16440 gnd.n4849 gnd.n4848 9.56018
R16441 gnd.n4772 gnd.n1422 9.56018
R16442 gnd.n4907 gnd.t195 9.56018
R16443 gnd.n5850 gnd.n999 9.45599
R16444 gnd.n5029 gnd.n5028 9.45599
R16445 gnd.n3427 gnd.n3426 9.45567
R16446 gnd.n3395 gnd.n3394 9.45567
R16447 gnd.n3363 gnd.n3362 9.45567
R16448 gnd.n3332 gnd.n3331 9.45567
R16449 gnd.n3300 gnd.n3299 9.45567
R16450 gnd.n3268 gnd.n3267 9.45567
R16451 gnd.n3236 gnd.n3235 9.45567
R16452 gnd.n3205 gnd.n3204 9.45567
R16453 gnd.n2372 gnd.n2371 9.39724
R16454 gnd.n3426 gnd.n3425 9.3005
R16455 gnd.n3399 gnd.n3398 9.3005
R16456 gnd.n3420 gnd.n3419 9.3005
R16457 gnd.n3418 gnd.n3417 9.3005
R16458 gnd.n3403 gnd.n3402 9.3005
R16459 gnd.n3412 gnd.n3411 9.3005
R16460 gnd.n3410 gnd.n3409 9.3005
R16461 gnd.n3394 gnd.n3393 9.3005
R16462 gnd.n3367 gnd.n3366 9.3005
R16463 gnd.n3388 gnd.n3387 9.3005
R16464 gnd.n3386 gnd.n3385 9.3005
R16465 gnd.n3371 gnd.n3370 9.3005
R16466 gnd.n3380 gnd.n3379 9.3005
R16467 gnd.n3378 gnd.n3377 9.3005
R16468 gnd.n3362 gnd.n3361 9.3005
R16469 gnd.n3335 gnd.n3334 9.3005
R16470 gnd.n3356 gnd.n3355 9.3005
R16471 gnd.n3354 gnd.n3353 9.3005
R16472 gnd.n3339 gnd.n3338 9.3005
R16473 gnd.n3348 gnd.n3347 9.3005
R16474 gnd.n3346 gnd.n3345 9.3005
R16475 gnd.n3331 gnd.n3330 9.3005
R16476 gnd.n3304 gnd.n3303 9.3005
R16477 gnd.n3325 gnd.n3324 9.3005
R16478 gnd.n3323 gnd.n3322 9.3005
R16479 gnd.n3308 gnd.n3307 9.3005
R16480 gnd.n3317 gnd.n3316 9.3005
R16481 gnd.n3315 gnd.n3314 9.3005
R16482 gnd.n3299 gnd.n3298 9.3005
R16483 gnd.n3272 gnd.n3271 9.3005
R16484 gnd.n3293 gnd.n3292 9.3005
R16485 gnd.n3291 gnd.n3290 9.3005
R16486 gnd.n3276 gnd.n3275 9.3005
R16487 gnd.n3285 gnd.n3284 9.3005
R16488 gnd.n3283 gnd.n3282 9.3005
R16489 gnd.n3267 gnd.n3266 9.3005
R16490 gnd.n3240 gnd.n3239 9.3005
R16491 gnd.n3261 gnd.n3260 9.3005
R16492 gnd.n3259 gnd.n3258 9.3005
R16493 gnd.n3244 gnd.n3243 9.3005
R16494 gnd.n3253 gnd.n3252 9.3005
R16495 gnd.n3251 gnd.n3250 9.3005
R16496 gnd.n3235 gnd.n3234 9.3005
R16497 gnd.n3208 gnd.n3207 9.3005
R16498 gnd.n3229 gnd.n3228 9.3005
R16499 gnd.n3227 gnd.n3226 9.3005
R16500 gnd.n3212 gnd.n3211 9.3005
R16501 gnd.n3221 gnd.n3220 9.3005
R16502 gnd.n3219 gnd.n3218 9.3005
R16503 gnd.n3204 gnd.n3203 9.3005
R16504 gnd.n3177 gnd.n3176 9.3005
R16505 gnd.n3198 gnd.n3197 9.3005
R16506 gnd.n3196 gnd.n3195 9.3005
R16507 gnd.n3181 gnd.n3180 9.3005
R16508 gnd.n3190 gnd.n3189 9.3005
R16509 gnd.n3188 gnd.n3187 9.3005
R16510 gnd.n3552 gnd.n3551 9.3005
R16511 gnd.n3550 gnd.n2131 9.3005
R16512 gnd.n3549 gnd.n3548 9.3005
R16513 gnd.n3545 gnd.n2132 9.3005
R16514 gnd.n3542 gnd.n2133 9.3005
R16515 gnd.n3541 gnd.n2134 9.3005
R16516 gnd.n3538 gnd.n2135 9.3005
R16517 gnd.n3537 gnd.n2136 9.3005
R16518 gnd.n3534 gnd.n2137 9.3005
R16519 gnd.n3533 gnd.n2138 9.3005
R16520 gnd.n3530 gnd.n2139 9.3005
R16521 gnd.n3529 gnd.n2140 9.3005
R16522 gnd.n3526 gnd.n2141 9.3005
R16523 gnd.n3525 gnd.n2142 9.3005
R16524 gnd.n3522 gnd.n3521 9.3005
R16525 gnd.n3520 gnd.n2143 9.3005
R16526 gnd.n3553 gnd.n2130 9.3005
R16527 gnd.n2793 gnd.n2792 9.3005
R16528 gnd.n2497 gnd.n2496 9.3005
R16529 gnd.n2820 gnd.n2819 9.3005
R16530 gnd.n2821 gnd.n2495 9.3005
R16531 gnd.n2825 gnd.n2822 9.3005
R16532 gnd.n2824 gnd.n2823 9.3005
R16533 gnd.n2469 gnd.n2468 9.3005
R16534 gnd.n2850 gnd.n2849 9.3005
R16535 gnd.n2851 gnd.n2467 9.3005
R16536 gnd.n2853 gnd.n2852 9.3005
R16537 gnd.n2447 gnd.n2446 9.3005
R16538 gnd.n2881 gnd.n2880 9.3005
R16539 gnd.n2882 gnd.n2445 9.3005
R16540 gnd.n2890 gnd.n2883 9.3005
R16541 gnd.n2889 gnd.n2884 9.3005
R16542 gnd.n2888 gnd.n2886 9.3005
R16543 gnd.n2885 gnd.n2394 9.3005
R16544 gnd.n2938 gnd.n2395 9.3005
R16545 gnd.n2937 gnd.n2396 9.3005
R16546 gnd.n2936 gnd.n2397 9.3005
R16547 gnd.n2416 gnd.n2398 9.3005
R16548 gnd.n2418 gnd.n2417 9.3005
R16549 gnd.n2328 gnd.n2327 9.3005
R16550 gnd.n2976 gnd.n2975 9.3005
R16551 gnd.n2977 gnd.n2326 9.3005
R16552 gnd.n2981 gnd.n2978 9.3005
R16553 gnd.n2980 gnd.n2979 9.3005
R16554 gnd.n2301 gnd.n2300 9.3005
R16555 gnd.n3016 gnd.n3015 9.3005
R16556 gnd.n3017 gnd.n2299 9.3005
R16557 gnd.n3021 gnd.n3018 9.3005
R16558 gnd.n3020 gnd.n3019 9.3005
R16559 gnd.n2274 gnd.n2273 9.3005
R16560 gnd.n3061 gnd.n3060 9.3005
R16561 gnd.n3062 gnd.n2272 9.3005
R16562 gnd.n3066 gnd.n3063 9.3005
R16563 gnd.n3065 gnd.n3064 9.3005
R16564 gnd.n2246 gnd.n2245 9.3005
R16565 gnd.n3102 gnd.n3101 9.3005
R16566 gnd.n3103 gnd.n2244 9.3005
R16567 gnd.n3107 gnd.n3104 9.3005
R16568 gnd.n3106 gnd.n3105 9.3005
R16569 gnd.n2219 gnd.n2218 9.3005
R16570 gnd.n3151 gnd.n3150 9.3005
R16571 gnd.n3152 gnd.n2217 9.3005
R16572 gnd.n3156 gnd.n3153 9.3005
R16573 gnd.n3155 gnd.n3154 9.3005
R16574 gnd.n2192 gnd.n2191 9.3005
R16575 gnd.n3445 gnd.n3444 9.3005
R16576 gnd.n3446 gnd.n2190 9.3005
R16577 gnd.n3452 gnd.n3447 9.3005
R16578 gnd.n3451 gnd.n3448 9.3005
R16579 gnd.n3450 gnd.n3449 9.3005
R16580 gnd.n2794 gnd.n2791 9.3005
R16581 gnd.n2576 gnd.n2535 9.3005
R16582 gnd.n2571 gnd.n2570 9.3005
R16583 gnd.n2569 gnd.n2536 9.3005
R16584 gnd.n2568 gnd.n2567 9.3005
R16585 gnd.n2564 gnd.n2537 9.3005
R16586 gnd.n2561 gnd.n2560 9.3005
R16587 gnd.n2559 gnd.n2538 9.3005
R16588 gnd.n2558 gnd.n2557 9.3005
R16589 gnd.n2554 gnd.n2539 9.3005
R16590 gnd.n2551 gnd.n2550 9.3005
R16591 gnd.n2549 gnd.n2540 9.3005
R16592 gnd.n2548 gnd.n2547 9.3005
R16593 gnd.n2544 gnd.n2542 9.3005
R16594 gnd.n2541 gnd.n2521 9.3005
R16595 gnd.n2788 gnd.n2520 9.3005
R16596 gnd.n2790 gnd.n2789 9.3005
R16597 gnd.n2578 gnd.n2577 9.3005
R16598 gnd.n2801 gnd.n2507 9.3005
R16599 gnd.n2808 gnd.n2508 9.3005
R16600 gnd.n2810 gnd.n2809 9.3005
R16601 gnd.n2811 gnd.n2488 9.3005
R16602 gnd.n2830 gnd.n2829 9.3005
R16603 gnd.n2832 gnd.n2480 9.3005
R16604 gnd.n2839 gnd.n2482 9.3005
R16605 gnd.n2840 gnd.n2477 9.3005
R16606 gnd.n2842 gnd.n2841 9.3005
R16607 gnd.n2478 gnd.n2463 9.3005
R16608 gnd.n2858 gnd.n2461 9.3005
R16609 gnd.n2862 gnd.n2861 9.3005
R16610 gnd.n2860 gnd.n2437 9.3005
R16611 gnd.n2897 gnd.n2436 9.3005
R16612 gnd.n2900 gnd.n2899 9.3005
R16613 gnd.n2433 gnd.n2432 9.3005
R16614 gnd.n2906 gnd.n2434 9.3005
R16615 gnd.n2908 gnd.n2907 9.3005
R16616 gnd.n2910 gnd.n2431 9.3005
R16617 gnd.n2913 gnd.n2912 9.3005
R16618 gnd.n2916 gnd.n2914 9.3005
R16619 gnd.n2918 gnd.n2917 9.3005
R16620 gnd.n2924 gnd.n2919 9.3005
R16621 gnd.n2923 gnd.n2922 9.3005
R16622 gnd.n2319 gnd.n2318 9.3005
R16623 gnd.n2990 gnd.n2989 9.3005
R16624 gnd.n2991 gnd.n2312 9.3005
R16625 gnd.n2999 gnd.n2311 9.3005
R16626 gnd.n3002 gnd.n3001 9.3005
R16627 gnd.n3004 gnd.n3003 9.3005
R16628 gnd.n3007 gnd.n2294 9.3005
R16629 gnd.n3005 gnd.n2292 9.3005
R16630 gnd.n3027 gnd.n2290 9.3005
R16631 gnd.n3029 gnd.n3028 9.3005
R16632 gnd.n2264 gnd.n2263 9.3005
R16633 gnd.n3075 gnd.n3074 9.3005
R16634 gnd.n3076 gnd.n2257 9.3005
R16635 gnd.n3085 gnd.n2256 9.3005
R16636 gnd.n3088 gnd.n3087 9.3005
R16637 gnd.n3090 gnd.n3089 9.3005
R16638 gnd.n3093 gnd.n2239 9.3005
R16639 gnd.n3091 gnd.n2237 9.3005
R16640 gnd.n3113 gnd.n2235 9.3005
R16641 gnd.n3115 gnd.n3114 9.3005
R16642 gnd.n2210 gnd.n2209 9.3005
R16643 gnd.n3165 gnd.n3164 9.3005
R16644 gnd.n3166 gnd.n2203 9.3005
R16645 gnd.n3174 gnd.n2202 9.3005
R16646 gnd.n3433 gnd.n3432 9.3005
R16647 gnd.n3435 gnd.n3434 9.3005
R16648 gnd.n3436 gnd.n2183 9.3005
R16649 gnd.n3460 gnd.n3459 9.3005
R16650 gnd.n2184 gnd.n2146 9.3005
R16651 gnd.n2799 gnd.n2798 9.3005
R16652 gnd.n3516 gnd.n2147 9.3005
R16653 gnd.n3515 gnd.n2149 9.3005
R16654 gnd.n3512 gnd.n2150 9.3005
R16655 gnd.n3511 gnd.n2151 9.3005
R16656 gnd.n3508 gnd.n2152 9.3005
R16657 gnd.n3507 gnd.n2153 9.3005
R16658 gnd.n3504 gnd.n2154 9.3005
R16659 gnd.n3503 gnd.n2155 9.3005
R16660 gnd.n3500 gnd.n2156 9.3005
R16661 gnd.n3499 gnd.n2157 9.3005
R16662 gnd.n3496 gnd.n2158 9.3005
R16663 gnd.n3495 gnd.n2159 9.3005
R16664 gnd.n3492 gnd.n2160 9.3005
R16665 gnd.n3491 gnd.n2161 9.3005
R16666 gnd.n3488 gnd.n2162 9.3005
R16667 gnd.n3487 gnd.n2163 9.3005
R16668 gnd.n3484 gnd.n2164 9.3005
R16669 gnd.n3483 gnd.n2165 9.3005
R16670 gnd.n3480 gnd.n2166 9.3005
R16671 gnd.n3479 gnd.n2167 9.3005
R16672 gnd.n3476 gnd.n2168 9.3005
R16673 gnd.n3475 gnd.n2169 9.3005
R16674 gnd.n3472 gnd.n2173 9.3005
R16675 gnd.n3471 gnd.n2174 9.3005
R16676 gnd.n3468 gnd.n2175 9.3005
R16677 gnd.n3467 gnd.n2176 9.3005
R16678 gnd.n3518 gnd.n3517 9.3005
R16679 gnd.n2968 gnd.n2952 9.3005
R16680 gnd.n2967 gnd.n2953 9.3005
R16681 gnd.n2966 gnd.n2954 9.3005
R16682 gnd.n2964 gnd.n2955 9.3005
R16683 gnd.n2963 gnd.n2956 9.3005
R16684 gnd.n2961 gnd.n2957 9.3005
R16685 gnd.n2960 gnd.n2958 9.3005
R16686 gnd.n2282 gnd.n2281 9.3005
R16687 gnd.n3037 gnd.n3036 9.3005
R16688 gnd.n3038 gnd.n2280 9.3005
R16689 gnd.n3055 gnd.n3039 9.3005
R16690 gnd.n3054 gnd.n3040 9.3005
R16691 gnd.n3053 gnd.n3041 9.3005
R16692 gnd.n3051 gnd.n3042 9.3005
R16693 gnd.n3050 gnd.n3043 9.3005
R16694 gnd.n3048 gnd.n3044 9.3005
R16695 gnd.n3047 gnd.n3045 9.3005
R16696 gnd.n2226 gnd.n2225 9.3005
R16697 gnd.n3123 gnd.n3122 9.3005
R16698 gnd.n3124 gnd.n2224 9.3005
R16699 gnd.n3145 gnd.n3125 9.3005
R16700 gnd.n3144 gnd.n3126 9.3005
R16701 gnd.n3143 gnd.n3127 9.3005
R16702 gnd.n3140 gnd.n3128 9.3005
R16703 gnd.n3139 gnd.n3129 9.3005
R16704 gnd.n3137 gnd.n3130 9.3005
R16705 gnd.n3136 gnd.n3131 9.3005
R16706 gnd.n3134 gnd.n3133 9.3005
R16707 gnd.n3132 gnd.n2178 9.3005
R16708 gnd.n2709 gnd.n2708 9.3005
R16709 gnd.n2599 gnd.n2598 9.3005
R16710 gnd.n2723 gnd.n2722 9.3005
R16711 gnd.n2724 gnd.n2597 9.3005
R16712 gnd.n2726 gnd.n2725 9.3005
R16713 gnd.n2587 gnd.n2586 9.3005
R16714 gnd.n2739 gnd.n2738 9.3005
R16715 gnd.n2740 gnd.n2585 9.3005
R16716 gnd.n2772 gnd.n2741 9.3005
R16717 gnd.n2771 gnd.n2742 9.3005
R16718 gnd.n2770 gnd.n2743 9.3005
R16719 gnd.n2769 gnd.n2744 9.3005
R16720 gnd.n2766 gnd.n2745 9.3005
R16721 gnd.n2765 gnd.n2746 9.3005
R16722 gnd.n2764 gnd.n2747 9.3005
R16723 gnd.n2762 gnd.n2748 9.3005
R16724 gnd.n2761 gnd.n2749 9.3005
R16725 gnd.n2758 gnd.n2750 9.3005
R16726 gnd.n2757 gnd.n2751 9.3005
R16727 gnd.n2756 gnd.n2752 9.3005
R16728 gnd.n2754 gnd.n2753 9.3005
R16729 gnd.n2453 gnd.n2452 9.3005
R16730 gnd.n2870 gnd.n2869 9.3005
R16731 gnd.n2871 gnd.n2451 9.3005
R16732 gnd.n2875 gnd.n2872 9.3005
R16733 gnd.n2874 gnd.n2873 9.3005
R16734 gnd.n2375 gnd.n2374 9.3005
R16735 gnd.n2950 gnd.n2949 9.3005
R16736 gnd.n2707 gnd.n2608 9.3005
R16737 gnd.n2610 gnd.n2609 9.3005
R16738 gnd.n2654 gnd.n2652 9.3005
R16739 gnd.n2655 gnd.n2651 9.3005
R16740 gnd.n2658 gnd.n2647 9.3005
R16741 gnd.n2659 gnd.n2646 9.3005
R16742 gnd.n2662 gnd.n2645 9.3005
R16743 gnd.n2663 gnd.n2644 9.3005
R16744 gnd.n2666 gnd.n2643 9.3005
R16745 gnd.n2667 gnd.n2642 9.3005
R16746 gnd.n2670 gnd.n2641 9.3005
R16747 gnd.n2671 gnd.n2640 9.3005
R16748 gnd.n2674 gnd.n2639 9.3005
R16749 gnd.n2675 gnd.n2638 9.3005
R16750 gnd.n2678 gnd.n2637 9.3005
R16751 gnd.n2679 gnd.n2636 9.3005
R16752 gnd.n2682 gnd.n2635 9.3005
R16753 gnd.n2683 gnd.n2634 9.3005
R16754 gnd.n2686 gnd.n2633 9.3005
R16755 gnd.n2687 gnd.n2632 9.3005
R16756 gnd.n2690 gnd.n2631 9.3005
R16757 gnd.n2691 gnd.n2630 9.3005
R16758 gnd.n2694 gnd.n2629 9.3005
R16759 gnd.n2696 gnd.n2628 9.3005
R16760 gnd.n2697 gnd.n2627 9.3005
R16761 gnd.n2698 gnd.n2626 9.3005
R16762 gnd.n2699 gnd.n2625 9.3005
R16763 gnd.n2706 gnd.n2705 9.3005
R16764 gnd.n2715 gnd.n2714 9.3005
R16765 gnd.n2716 gnd.n2602 9.3005
R16766 gnd.n2718 gnd.n2717 9.3005
R16767 gnd.n2593 gnd.n2592 9.3005
R16768 gnd.n2731 gnd.n2730 9.3005
R16769 gnd.n2732 gnd.n2591 9.3005
R16770 gnd.n2734 gnd.n2733 9.3005
R16771 gnd.n2580 gnd.n2579 9.3005
R16772 gnd.n2777 gnd.n2776 9.3005
R16773 gnd.n2778 gnd.n2534 9.3005
R16774 gnd.n2782 gnd.n2780 9.3005
R16775 gnd.n2781 gnd.n2513 9.3005
R16776 gnd.n2800 gnd.n2512 9.3005
R16777 gnd.n2803 gnd.n2802 9.3005
R16778 gnd.n2506 gnd.n2505 9.3005
R16779 gnd.n2814 gnd.n2812 9.3005
R16780 gnd.n2813 gnd.n2487 9.3005
R16781 gnd.n2831 gnd.n2486 9.3005
R16782 gnd.n2834 gnd.n2833 9.3005
R16783 gnd.n2481 gnd.n2476 9.3005
R16784 gnd.n2844 gnd.n2843 9.3005
R16785 gnd.n2479 gnd.n2459 9.3005
R16786 gnd.n2865 gnd.n2460 9.3005
R16787 gnd.n2864 gnd.n2863 9.3005
R16788 gnd.n2462 gnd.n2438 9.3005
R16789 gnd.n2896 gnd.n2895 9.3005
R16790 gnd.n2898 gnd.n2383 9.3005
R16791 gnd.n2945 gnd.n2384 9.3005
R16792 gnd.n2944 gnd.n2385 9.3005
R16793 gnd.n2943 gnd.n2386 9.3005
R16794 gnd.n2909 gnd.n2387 9.3005
R16795 gnd.n2911 gnd.n2405 9.3005
R16796 gnd.n2931 gnd.n2406 9.3005
R16797 gnd.n2930 gnd.n2407 9.3005
R16798 gnd.n2929 gnd.n2408 9.3005
R16799 gnd.n2920 gnd.n2409 9.3005
R16800 gnd.n2921 gnd.n2320 9.3005
R16801 gnd.n2987 gnd.n2986 9.3005
R16802 gnd.n2988 gnd.n2313 9.3005
R16803 gnd.n2998 gnd.n2997 9.3005
R16804 gnd.n3000 gnd.n2309 9.3005
R16805 gnd.n3010 gnd.n2310 9.3005
R16806 gnd.n3009 gnd.n3008 9.3005
R16807 gnd.n3006 gnd.n2288 9.3005
R16808 gnd.n3032 gnd.n2289 9.3005
R16809 gnd.n3031 gnd.n3030 9.3005
R16810 gnd.n2291 gnd.n2265 9.3005
R16811 gnd.n3072 gnd.n3071 9.3005
R16812 gnd.n3073 gnd.n2258 9.3005
R16813 gnd.n3084 gnd.n3083 9.3005
R16814 gnd.n3086 gnd.n2254 9.3005
R16815 gnd.n3096 gnd.n2255 9.3005
R16816 gnd.n3095 gnd.n3094 9.3005
R16817 gnd.n3092 gnd.n2233 9.3005
R16818 gnd.n3118 gnd.n2234 9.3005
R16819 gnd.n3117 gnd.n3116 9.3005
R16820 gnd.n2236 gnd.n2211 9.3005
R16821 gnd.n3162 gnd.n3161 9.3005
R16822 gnd.n3163 gnd.n2204 9.3005
R16823 gnd.n3173 gnd.n3172 9.3005
R16824 gnd.n3431 gnd.n2200 9.3005
R16825 gnd.n3439 gnd.n2201 9.3005
R16826 gnd.n3438 gnd.n3437 9.3005
R16827 gnd.n2182 gnd.n2181 9.3005
R16828 gnd.n3462 gnd.n3461 9.3005
R16829 gnd.n2604 gnd.n2603 9.3005
R16830 gnd.n6119 gnd.n657 9.3005
R16831 gnd.n6121 gnd.n6120 9.3005
R16832 gnd.n653 gnd.n652 9.3005
R16833 gnd.n6128 gnd.n6127 9.3005
R16834 gnd.n6129 gnd.n651 9.3005
R16835 gnd.n6131 gnd.n6130 9.3005
R16836 gnd.n647 gnd.n646 9.3005
R16837 gnd.n6138 gnd.n6137 9.3005
R16838 gnd.n6139 gnd.n645 9.3005
R16839 gnd.n6141 gnd.n6140 9.3005
R16840 gnd.n641 gnd.n640 9.3005
R16841 gnd.n6148 gnd.n6147 9.3005
R16842 gnd.n6149 gnd.n639 9.3005
R16843 gnd.n6151 gnd.n6150 9.3005
R16844 gnd.n635 gnd.n634 9.3005
R16845 gnd.n6158 gnd.n6157 9.3005
R16846 gnd.n6159 gnd.n633 9.3005
R16847 gnd.n6161 gnd.n6160 9.3005
R16848 gnd.n629 gnd.n628 9.3005
R16849 gnd.n6168 gnd.n6167 9.3005
R16850 gnd.n6169 gnd.n627 9.3005
R16851 gnd.n6171 gnd.n6170 9.3005
R16852 gnd.n623 gnd.n622 9.3005
R16853 gnd.n6178 gnd.n6177 9.3005
R16854 gnd.n6179 gnd.n621 9.3005
R16855 gnd.n6181 gnd.n6180 9.3005
R16856 gnd.n617 gnd.n616 9.3005
R16857 gnd.n6188 gnd.n6187 9.3005
R16858 gnd.n6189 gnd.n615 9.3005
R16859 gnd.n6191 gnd.n6190 9.3005
R16860 gnd.n611 gnd.n610 9.3005
R16861 gnd.n6198 gnd.n6197 9.3005
R16862 gnd.n6199 gnd.n609 9.3005
R16863 gnd.n6201 gnd.n6200 9.3005
R16864 gnd.n605 gnd.n604 9.3005
R16865 gnd.n6208 gnd.n6207 9.3005
R16866 gnd.n6209 gnd.n603 9.3005
R16867 gnd.n6211 gnd.n6210 9.3005
R16868 gnd.n599 gnd.n598 9.3005
R16869 gnd.n6218 gnd.n6217 9.3005
R16870 gnd.n6219 gnd.n597 9.3005
R16871 gnd.n6221 gnd.n6220 9.3005
R16872 gnd.n593 gnd.n592 9.3005
R16873 gnd.n6228 gnd.n6227 9.3005
R16874 gnd.n6229 gnd.n591 9.3005
R16875 gnd.n6231 gnd.n6230 9.3005
R16876 gnd.n587 gnd.n586 9.3005
R16877 gnd.n6238 gnd.n6237 9.3005
R16878 gnd.n6239 gnd.n585 9.3005
R16879 gnd.n6241 gnd.n6240 9.3005
R16880 gnd.n581 gnd.n580 9.3005
R16881 gnd.n6248 gnd.n6247 9.3005
R16882 gnd.n6249 gnd.n579 9.3005
R16883 gnd.n6251 gnd.n6250 9.3005
R16884 gnd.n575 gnd.n574 9.3005
R16885 gnd.n6258 gnd.n6257 9.3005
R16886 gnd.n6259 gnd.n573 9.3005
R16887 gnd.n6261 gnd.n6260 9.3005
R16888 gnd.n569 gnd.n568 9.3005
R16889 gnd.n6268 gnd.n6267 9.3005
R16890 gnd.n6269 gnd.n567 9.3005
R16891 gnd.n6271 gnd.n6270 9.3005
R16892 gnd.n563 gnd.n562 9.3005
R16893 gnd.n6278 gnd.n6277 9.3005
R16894 gnd.n6279 gnd.n561 9.3005
R16895 gnd.n6281 gnd.n6280 9.3005
R16896 gnd.n557 gnd.n556 9.3005
R16897 gnd.n6288 gnd.n6287 9.3005
R16898 gnd.n6289 gnd.n555 9.3005
R16899 gnd.n6291 gnd.n6290 9.3005
R16900 gnd.n551 gnd.n550 9.3005
R16901 gnd.n6298 gnd.n6297 9.3005
R16902 gnd.n6299 gnd.n549 9.3005
R16903 gnd.n6301 gnd.n6300 9.3005
R16904 gnd.n545 gnd.n544 9.3005
R16905 gnd.n6308 gnd.n6307 9.3005
R16906 gnd.n6309 gnd.n543 9.3005
R16907 gnd.n6311 gnd.n6310 9.3005
R16908 gnd.n539 gnd.n538 9.3005
R16909 gnd.n6318 gnd.n6317 9.3005
R16910 gnd.n6319 gnd.n537 9.3005
R16911 gnd.n6321 gnd.n6320 9.3005
R16912 gnd.n533 gnd.n532 9.3005
R16913 gnd.n6328 gnd.n6327 9.3005
R16914 gnd.n6329 gnd.n531 9.3005
R16915 gnd.n6331 gnd.n6330 9.3005
R16916 gnd.n527 gnd.n526 9.3005
R16917 gnd.n6338 gnd.n6337 9.3005
R16918 gnd.n6339 gnd.n525 9.3005
R16919 gnd.n6341 gnd.n6340 9.3005
R16920 gnd.n521 gnd.n520 9.3005
R16921 gnd.n6348 gnd.n6347 9.3005
R16922 gnd.n6349 gnd.n519 9.3005
R16923 gnd.n6351 gnd.n6350 9.3005
R16924 gnd.n515 gnd.n514 9.3005
R16925 gnd.n6358 gnd.n6357 9.3005
R16926 gnd.n6359 gnd.n513 9.3005
R16927 gnd.n6361 gnd.n6360 9.3005
R16928 gnd.n509 gnd.n508 9.3005
R16929 gnd.n6368 gnd.n6367 9.3005
R16930 gnd.n6369 gnd.n507 9.3005
R16931 gnd.n6371 gnd.n6370 9.3005
R16932 gnd.n503 gnd.n502 9.3005
R16933 gnd.n6378 gnd.n6377 9.3005
R16934 gnd.n6379 gnd.n501 9.3005
R16935 gnd.n6381 gnd.n6380 9.3005
R16936 gnd.n497 gnd.n496 9.3005
R16937 gnd.n6388 gnd.n6387 9.3005
R16938 gnd.n6389 gnd.n495 9.3005
R16939 gnd.n6391 gnd.n6390 9.3005
R16940 gnd.n491 gnd.n490 9.3005
R16941 gnd.n6398 gnd.n6397 9.3005
R16942 gnd.n6399 gnd.n489 9.3005
R16943 gnd.n6401 gnd.n6400 9.3005
R16944 gnd.n485 gnd.n484 9.3005
R16945 gnd.n6408 gnd.n6407 9.3005
R16946 gnd.n6409 gnd.n483 9.3005
R16947 gnd.n6411 gnd.n6410 9.3005
R16948 gnd.n479 gnd.n478 9.3005
R16949 gnd.n6418 gnd.n6417 9.3005
R16950 gnd.n6419 gnd.n477 9.3005
R16951 gnd.n6421 gnd.n6420 9.3005
R16952 gnd.n473 gnd.n472 9.3005
R16953 gnd.n6428 gnd.n6427 9.3005
R16954 gnd.n6429 gnd.n471 9.3005
R16955 gnd.n6431 gnd.n6430 9.3005
R16956 gnd.n467 gnd.n466 9.3005
R16957 gnd.n6438 gnd.n6437 9.3005
R16958 gnd.n6439 gnd.n465 9.3005
R16959 gnd.n6441 gnd.n6440 9.3005
R16960 gnd.n461 gnd.n460 9.3005
R16961 gnd.n6448 gnd.n6447 9.3005
R16962 gnd.n6449 gnd.n459 9.3005
R16963 gnd.n6451 gnd.n6450 9.3005
R16964 gnd.n455 gnd.n454 9.3005
R16965 gnd.n6458 gnd.n6457 9.3005
R16966 gnd.n6459 gnd.n453 9.3005
R16967 gnd.n6461 gnd.n6460 9.3005
R16968 gnd.n449 gnd.n448 9.3005
R16969 gnd.n6468 gnd.n6467 9.3005
R16970 gnd.n6469 gnd.n447 9.3005
R16971 gnd.n6471 gnd.n6470 9.3005
R16972 gnd.n443 gnd.n442 9.3005
R16973 gnd.n6478 gnd.n6477 9.3005
R16974 gnd.n6479 gnd.n441 9.3005
R16975 gnd.n6481 gnd.n6480 9.3005
R16976 gnd.n437 gnd.n436 9.3005
R16977 gnd.n6488 gnd.n6487 9.3005
R16978 gnd.n6489 gnd.n435 9.3005
R16979 gnd.n6491 gnd.n6490 9.3005
R16980 gnd.n431 gnd.n430 9.3005
R16981 gnd.n6498 gnd.n6497 9.3005
R16982 gnd.n6499 gnd.n429 9.3005
R16983 gnd.n6501 gnd.n6500 9.3005
R16984 gnd.n425 gnd.n424 9.3005
R16985 gnd.n6508 gnd.n6507 9.3005
R16986 gnd.n6509 gnd.n423 9.3005
R16987 gnd.n6511 gnd.n6510 9.3005
R16988 gnd.n419 gnd.n418 9.3005
R16989 gnd.n6518 gnd.n6517 9.3005
R16990 gnd.n6519 gnd.n417 9.3005
R16991 gnd.n6521 gnd.n6520 9.3005
R16992 gnd.n413 gnd.n412 9.3005
R16993 gnd.n6528 gnd.n6527 9.3005
R16994 gnd.n6529 gnd.n411 9.3005
R16995 gnd.n6531 gnd.n6530 9.3005
R16996 gnd.n407 gnd.n406 9.3005
R16997 gnd.n6538 gnd.n6537 9.3005
R16998 gnd.n6541 gnd.n6540 9.3005
R16999 gnd.n401 gnd.n400 9.3005
R17000 gnd.n6548 gnd.n6547 9.3005
R17001 gnd.n6549 gnd.n399 9.3005
R17002 gnd.n6551 gnd.n6550 9.3005
R17003 gnd.n395 gnd.n394 9.3005
R17004 gnd.n6558 gnd.n6557 9.3005
R17005 gnd.n6559 gnd.n393 9.3005
R17006 gnd.n6561 gnd.n6560 9.3005
R17007 gnd.n389 gnd.n388 9.3005
R17008 gnd.n6568 gnd.n6567 9.3005
R17009 gnd.n6569 gnd.n387 9.3005
R17010 gnd.n6571 gnd.n6570 9.3005
R17011 gnd.n383 gnd.n382 9.3005
R17012 gnd.n6578 gnd.n6577 9.3005
R17013 gnd.n6579 gnd.n381 9.3005
R17014 gnd.n6581 gnd.n6580 9.3005
R17015 gnd.n377 gnd.n376 9.3005
R17016 gnd.n6588 gnd.n6587 9.3005
R17017 gnd.n6589 gnd.n375 9.3005
R17018 gnd.n6591 gnd.n6590 9.3005
R17019 gnd.n371 gnd.n370 9.3005
R17020 gnd.n6598 gnd.n6597 9.3005
R17021 gnd.n6599 gnd.n369 9.3005
R17022 gnd.n6601 gnd.n6600 9.3005
R17023 gnd.n365 gnd.n364 9.3005
R17024 gnd.n6608 gnd.n6607 9.3005
R17025 gnd.n6609 gnd.n363 9.3005
R17026 gnd.n6611 gnd.n6610 9.3005
R17027 gnd.n359 gnd.n358 9.3005
R17028 gnd.n6618 gnd.n6617 9.3005
R17029 gnd.n6619 gnd.n357 9.3005
R17030 gnd.n6621 gnd.n6620 9.3005
R17031 gnd.n353 gnd.n352 9.3005
R17032 gnd.n6628 gnd.n6627 9.3005
R17033 gnd.n6629 gnd.n351 9.3005
R17034 gnd.n6631 gnd.n6630 9.3005
R17035 gnd.n347 gnd.n346 9.3005
R17036 gnd.n6638 gnd.n6637 9.3005
R17037 gnd.n6639 gnd.n345 9.3005
R17038 gnd.n6641 gnd.n6640 9.3005
R17039 gnd.n341 gnd.n340 9.3005
R17040 gnd.n6648 gnd.n6647 9.3005
R17041 gnd.n6649 gnd.n339 9.3005
R17042 gnd.n6651 gnd.n6650 9.3005
R17043 gnd.n335 gnd.n334 9.3005
R17044 gnd.n6658 gnd.n6657 9.3005
R17045 gnd.n6659 gnd.n333 9.3005
R17046 gnd.n6661 gnd.n6660 9.3005
R17047 gnd.n329 gnd.n328 9.3005
R17048 gnd.n6668 gnd.n6667 9.3005
R17049 gnd.n6669 gnd.n327 9.3005
R17050 gnd.n6671 gnd.n6670 9.3005
R17051 gnd.n323 gnd.n322 9.3005
R17052 gnd.n6678 gnd.n6677 9.3005
R17053 gnd.n6679 gnd.n321 9.3005
R17054 gnd.n6681 gnd.n6680 9.3005
R17055 gnd.n317 gnd.n316 9.3005
R17056 gnd.n6688 gnd.n6687 9.3005
R17057 gnd.n6689 gnd.n315 9.3005
R17058 gnd.n6691 gnd.n6690 9.3005
R17059 gnd.n311 gnd.n310 9.3005
R17060 gnd.n6698 gnd.n6697 9.3005
R17061 gnd.n6699 gnd.n309 9.3005
R17062 gnd.n6701 gnd.n6700 9.3005
R17063 gnd.n305 gnd.n304 9.3005
R17064 gnd.n6708 gnd.n6707 9.3005
R17065 gnd.n6709 gnd.n303 9.3005
R17066 gnd.n6711 gnd.n6710 9.3005
R17067 gnd.n299 gnd.n298 9.3005
R17068 gnd.n6718 gnd.n6717 9.3005
R17069 gnd.n6719 gnd.n297 9.3005
R17070 gnd.n6721 gnd.n6720 9.3005
R17071 gnd.n293 gnd.n292 9.3005
R17072 gnd.n6728 gnd.n6727 9.3005
R17073 gnd.n6729 gnd.n291 9.3005
R17074 gnd.n6731 gnd.n6730 9.3005
R17075 gnd.n287 gnd.n286 9.3005
R17076 gnd.n6738 gnd.n6737 9.3005
R17077 gnd.n6739 gnd.n285 9.3005
R17078 gnd.n6743 gnd.n6740 9.3005
R17079 gnd.n6742 gnd.n6741 9.3005
R17080 gnd.n281 gnd.n280 9.3005
R17081 gnd.n6751 gnd.n6750 9.3005
R17082 gnd.n6539 gnd.n405 9.3005
R17083 gnd.n7000 gnd.n89 9.3005
R17084 gnd.n6999 gnd.n91 9.3005
R17085 gnd.n95 gnd.n92 9.3005
R17086 gnd.n6994 gnd.n96 9.3005
R17087 gnd.n6993 gnd.n97 9.3005
R17088 gnd.n6992 gnd.n98 9.3005
R17089 gnd.n102 gnd.n99 9.3005
R17090 gnd.n6987 gnd.n103 9.3005
R17091 gnd.n6986 gnd.n104 9.3005
R17092 gnd.n6985 gnd.n105 9.3005
R17093 gnd.n109 gnd.n106 9.3005
R17094 gnd.n6980 gnd.n110 9.3005
R17095 gnd.n6979 gnd.n111 9.3005
R17096 gnd.n6978 gnd.n112 9.3005
R17097 gnd.n116 gnd.n113 9.3005
R17098 gnd.n6973 gnd.n117 9.3005
R17099 gnd.n6972 gnd.n118 9.3005
R17100 gnd.n6968 gnd.n119 9.3005
R17101 gnd.n123 gnd.n120 9.3005
R17102 gnd.n6963 gnd.n124 9.3005
R17103 gnd.n6962 gnd.n125 9.3005
R17104 gnd.n6961 gnd.n126 9.3005
R17105 gnd.n130 gnd.n127 9.3005
R17106 gnd.n6956 gnd.n131 9.3005
R17107 gnd.n6955 gnd.n132 9.3005
R17108 gnd.n6954 gnd.n133 9.3005
R17109 gnd.n137 gnd.n134 9.3005
R17110 gnd.n6949 gnd.n138 9.3005
R17111 gnd.n6948 gnd.n139 9.3005
R17112 gnd.n6947 gnd.n140 9.3005
R17113 gnd.n144 gnd.n141 9.3005
R17114 gnd.n6942 gnd.n145 9.3005
R17115 gnd.n6941 gnd.n146 9.3005
R17116 gnd.n6940 gnd.n147 9.3005
R17117 gnd.n151 gnd.n148 9.3005
R17118 gnd.n6935 gnd.n152 9.3005
R17119 gnd.n6934 gnd.n6933 9.3005
R17120 gnd.n6932 gnd.n155 9.3005
R17121 gnd.n7002 gnd.n7001 9.3005
R17122 gnd.n5466 gnd.n5465 9.3005
R17123 gnd.n1261 gnd.n1260 9.3005
R17124 gnd.n5480 gnd.n5479 9.3005
R17125 gnd.n5481 gnd.n1259 9.3005
R17126 gnd.n5524 gnd.n5482 9.3005
R17127 gnd.n5523 gnd.n5483 9.3005
R17128 gnd.n5522 gnd.n5484 9.3005
R17129 gnd.n5520 gnd.n5485 9.3005
R17130 gnd.n5519 gnd.n5486 9.3005
R17131 gnd.n5518 gnd.n5487 9.3005
R17132 gnd.n5516 gnd.n5488 9.3005
R17133 gnd.n5515 gnd.n5489 9.3005
R17134 gnd.n5513 gnd.n5490 9.3005
R17135 gnd.n5512 gnd.n5491 9.3005
R17136 gnd.n5511 gnd.n5492 9.3005
R17137 gnd.n5509 gnd.n5493 9.3005
R17138 gnd.n5508 gnd.n5494 9.3005
R17139 gnd.n5505 gnd.n5495 9.3005
R17140 gnd.n5504 gnd.n5496 9.3005
R17141 gnd.n5502 gnd.n5497 9.3005
R17142 gnd.n5501 gnd.n5499 9.3005
R17143 gnd.n5498 gnd.n237 9.3005
R17144 gnd.n6781 gnd.n238 9.3005
R17145 gnd.n6780 gnd.n239 9.3005
R17146 gnd.n6779 gnd.n240 9.3005
R17147 gnd.n6775 gnd.n241 9.3005
R17148 gnd.n6774 gnd.n242 9.3005
R17149 gnd.n6771 gnd.n243 9.3005
R17150 gnd.n6770 gnd.n244 9.3005
R17151 gnd.n6766 gnd.n245 9.3005
R17152 gnd.n6765 gnd.n246 9.3005
R17153 gnd.n269 gnd.n247 9.3005
R17154 gnd.n268 gnd.n248 9.3005
R17155 gnd.n264 gnd.n249 9.3005
R17156 gnd.n263 gnd.n250 9.3005
R17157 gnd.n260 gnd.n251 9.3005
R17158 gnd.n259 gnd.n252 9.3005
R17159 gnd.n257 gnd.n253 9.3005
R17160 gnd.n256 gnd.n255 9.3005
R17161 gnd.n254 gnd.n159 9.3005
R17162 gnd.n6929 gnd.n158 9.3005
R17163 gnd.n6931 gnd.n6930 9.3005
R17164 gnd.n5464 gnd.n1266 9.3005
R17165 gnd.n5453 gnd.n1271 9.3005
R17166 gnd.n5455 gnd.n5454 9.3005
R17167 gnd.n5452 gnd.n1273 9.3005
R17168 gnd.n5451 gnd.n5450 9.3005
R17169 gnd.n1275 gnd.n1274 9.3005
R17170 gnd.n5444 gnd.n5443 9.3005
R17171 gnd.n5442 gnd.n1277 9.3005
R17172 gnd.n5441 gnd.n5440 9.3005
R17173 gnd.n1279 gnd.n1278 9.3005
R17174 gnd.n5434 gnd.n5433 9.3005
R17175 gnd.n5432 gnd.n1281 9.3005
R17176 gnd.n5431 gnd.n5430 9.3005
R17177 gnd.n1283 gnd.n1282 9.3005
R17178 gnd.n5424 gnd.n5423 9.3005
R17179 gnd.n5422 gnd.n1285 9.3005
R17180 gnd.n5421 gnd.n5420 9.3005
R17181 gnd.n1287 gnd.n1286 9.3005
R17182 gnd.n5414 gnd.n5413 9.3005
R17183 gnd.n5412 gnd.n1289 9.3005
R17184 gnd.n1291 gnd.n1290 9.3005
R17185 gnd.n5399 gnd.n5354 9.3005
R17186 gnd.n5401 gnd.n5400 9.3005
R17187 gnd.n5398 gnd.n5356 9.3005
R17188 gnd.n5397 gnd.n5396 9.3005
R17189 gnd.n5358 gnd.n5357 9.3005
R17190 gnd.n5390 gnd.n5389 9.3005
R17191 gnd.n5388 gnd.n5360 9.3005
R17192 gnd.n5387 gnd.n5386 9.3005
R17193 gnd.n5362 gnd.n5361 9.3005
R17194 gnd.n5380 gnd.n5379 9.3005
R17195 gnd.n5378 gnd.n5364 9.3005
R17196 gnd.n5377 gnd.n5376 9.3005
R17197 gnd.n5366 gnd.n5365 9.3005
R17198 gnd.n5370 gnd.n5369 9.3005
R17199 gnd.n5368 gnd.n5367 9.3005
R17200 gnd.n1270 gnd.n1267 9.3005
R17201 gnd.n5463 gnd.n5462 9.3005
R17202 gnd.n5704 gnd.n1134 9.3005
R17203 gnd.n5703 gnd.n1135 9.3005
R17204 gnd.n1255 gnd.n1136 9.3005
R17205 gnd.n5547 gnd.n5546 9.3005
R17206 gnd.n5548 gnd.n1254 9.3005
R17207 gnd.n5552 gnd.n5549 9.3005
R17208 gnd.n5551 gnd.n5550 9.3005
R17209 gnd.n1228 gnd.n1227 9.3005
R17210 gnd.n5578 gnd.n5577 9.3005
R17211 gnd.n5579 gnd.n1226 9.3005
R17212 gnd.n5584 gnd.n5580 9.3005
R17213 gnd.n5583 gnd.n5582 9.3005
R17214 gnd.n5581 gnd.n1198 9.3005
R17215 gnd.n5615 gnd.n1199 9.3005
R17216 gnd.n5616 gnd.n214 9.3005
R17217 gnd.n6800 gnd.n213 9.3005
R17218 gnd.n6802 gnd.n6801 9.3005
R17219 gnd.n200 gnd.n199 9.3005
R17220 gnd.n6815 gnd.n6814 9.3005
R17221 gnd.n6816 gnd.n198 9.3005
R17222 gnd.n6818 gnd.n6817 9.3005
R17223 gnd.n184 gnd.n183 9.3005
R17224 gnd.n6831 gnd.n6830 9.3005
R17225 gnd.n6832 gnd.n182 9.3005
R17226 gnd.n6834 gnd.n6833 9.3005
R17227 gnd.n166 gnd.n165 9.3005
R17228 gnd.n6921 gnd.n6920 9.3005
R17229 gnd.n6922 gnd.n164 9.3005
R17230 gnd.n6924 gnd.n6923 9.3005
R17231 gnd.n88 gnd.n87 9.3005
R17232 gnd.n7004 gnd.n7003 9.3005
R17233 gnd.n5705 gnd.n1133 9.3005
R17234 gnd.n6799 gnd.n6798 9.3005
R17235 gnd.n3962 gnd.n3961 9.3005
R17236 gnd.n3966 gnd.n3963 9.3005
R17237 gnd.n3965 gnd.n3964 9.3005
R17238 gnd.n1986 gnd.n1985 9.3005
R17239 gnd.n4026 gnd.n4025 9.3005
R17240 gnd.n4027 gnd.n1984 9.3005
R17241 gnd.n4029 gnd.n4028 9.3005
R17242 gnd.n1982 gnd.n1981 9.3005
R17243 gnd.n4034 gnd.n4033 9.3005
R17244 gnd.n4035 gnd.n1980 9.3005
R17245 gnd.n4037 gnd.n4036 9.3005
R17246 gnd.n1978 gnd.n1977 9.3005
R17247 gnd.n4042 gnd.n4041 9.3005
R17248 gnd.n4043 gnd.n1976 9.3005
R17249 gnd.n4045 gnd.n4044 9.3005
R17250 gnd.n1974 gnd.n1973 9.3005
R17251 gnd.n4050 gnd.n4049 9.3005
R17252 gnd.n4051 gnd.n1972 9.3005
R17253 gnd.n4053 gnd.n4052 9.3005
R17254 gnd.n1968 gnd.n1967 9.3005
R17255 gnd.n4193 gnd.n4192 9.3005
R17256 gnd.n4194 gnd.n1966 9.3005
R17257 gnd.n4196 gnd.n4195 9.3005
R17258 gnd.n1962 gnd.n1961 9.3005
R17259 gnd.n4207 gnd.n4206 9.3005
R17260 gnd.n4208 gnd.n1960 9.3005
R17261 gnd.n4210 gnd.n4209 9.3005
R17262 gnd.n1954 gnd.n1953 9.3005
R17263 gnd.n4221 gnd.n4220 9.3005
R17264 gnd.n4222 gnd.n1952 9.3005
R17265 gnd.n4224 gnd.n4223 9.3005
R17266 gnd.n1946 gnd.n1945 9.3005
R17267 gnd.n4235 gnd.n4234 9.3005
R17268 gnd.n4236 gnd.n1944 9.3005
R17269 gnd.n4238 gnd.n4237 9.3005
R17270 gnd.n1669 gnd.n1668 9.3005
R17271 gnd.n4424 gnd.n4423 9.3005
R17272 gnd.n4425 gnd.n1667 9.3005
R17273 gnd.n4427 gnd.n4426 9.3005
R17274 gnd.n1651 gnd.n1650 9.3005
R17275 gnd.n4480 gnd.n4479 9.3005
R17276 gnd.n4481 gnd.n1649 9.3005
R17277 gnd.n4483 gnd.n4482 9.3005
R17278 gnd.n1630 gnd.n1629 9.3005
R17279 gnd.n4511 gnd.n4510 9.3005
R17280 gnd.n4512 gnd.n1628 9.3005
R17281 gnd.n4516 gnd.n4513 9.3005
R17282 gnd.n4515 gnd.n4514 9.3005
R17283 gnd.n1610 gnd.n1609 9.3005
R17284 gnd.n4541 gnd.n4540 9.3005
R17285 gnd.n4542 gnd.n1608 9.3005
R17286 gnd.n4554 gnd.n4543 9.3005
R17287 gnd.n4553 gnd.n4544 9.3005
R17288 gnd.n4552 gnd.n4545 9.3005
R17289 gnd.n4547 gnd.n4546 9.3005
R17290 gnd.n1563 gnd.n1562 9.3005
R17291 gnd.n4625 gnd.n4624 9.3005
R17292 gnd.n4626 gnd.n1561 9.3005
R17293 gnd.n4628 gnd.n4627 9.3005
R17294 gnd.n1540 gnd.n1539 9.3005
R17295 gnd.n4665 gnd.n4664 9.3005
R17296 gnd.n4666 gnd.n1538 9.3005
R17297 gnd.n4668 gnd.n4667 9.3005
R17298 gnd.n1518 gnd.n1517 9.3005
R17299 gnd.n4719 gnd.n4718 9.3005
R17300 gnd.n4720 gnd.n1516 9.3005
R17301 gnd.n4722 gnd.n4721 9.3005
R17302 gnd.n1499 gnd.n1498 9.3005
R17303 gnd.n4744 gnd.n4743 9.3005
R17304 gnd.n4745 gnd.n1497 9.3005
R17305 gnd.n4747 gnd.n4746 9.3005
R17306 gnd.n1477 gnd.n1476 9.3005
R17307 gnd.n4803 gnd.n4802 9.3005
R17308 gnd.n4804 gnd.n1475 9.3005
R17309 gnd.n4806 gnd.n4805 9.3005
R17310 gnd.n1455 gnd.n1454 9.3005
R17311 gnd.n4832 gnd.n4831 9.3005
R17312 gnd.n4833 gnd.n1453 9.3005
R17313 gnd.n4837 gnd.n4834 9.3005
R17314 gnd.n4836 gnd.n4835 9.3005
R17315 gnd.n1427 gnd.n1426 9.3005
R17316 gnd.n4887 gnd.n4886 9.3005
R17317 gnd.n4888 gnd.n1425 9.3005
R17318 gnd.n4890 gnd.n4889 9.3005
R17319 gnd.n1410 gnd.n1409 9.3005
R17320 gnd.n4913 gnd.n4912 9.3005
R17321 gnd.n4914 gnd.n1408 9.3005
R17322 gnd.n4919 gnd.n4915 9.3005
R17323 gnd.n4918 gnd.n4917 9.3005
R17324 gnd.n4916 gnd.n1346 9.3005
R17325 gnd.n5189 gnd.n1347 9.3005
R17326 gnd.n5188 gnd.n1348 9.3005
R17327 gnd.n5187 gnd.n1349 9.3005
R17328 gnd.n1357 gnd.n1350 9.3005
R17329 gnd.n1358 gnd.n1356 9.3005
R17330 gnd.n5177 gnd.n1359 9.3005
R17331 gnd.n5176 gnd.n1360 9.3005
R17332 gnd.n5175 gnd.n1361 9.3005
R17333 gnd.n1370 gnd.n1362 9.3005
R17334 gnd.n5166 gnd.n1371 9.3005
R17335 gnd.n5165 gnd.n1372 9.3005
R17336 gnd.n5164 gnd.n1373 9.3005
R17337 gnd.n5152 gnd.n1374 9.3005
R17338 gnd.n5155 gnd.n5154 9.3005
R17339 gnd.n5153 gnd.n1111 9.3005
R17340 gnd.n5720 gnd.n1112 9.3005
R17341 gnd.n5719 gnd.n1113 9.3005
R17342 gnd.n5718 gnd.n1114 9.3005
R17343 gnd.n1120 gnd.n1115 9.3005
R17344 gnd.n5712 gnd.n1121 9.3005
R17345 gnd.n5711 gnd.n1122 9.3005
R17346 gnd.n5710 gnd.n1123 9.3005
R17347 gnd.n5530 gnd.n1124 9.3005
R17348 gnd.n5532 gnd.n5531 9.3005
R17349 gnd.n5536 gnd.n5535 9.3005
R17350 gnd.n5537 gnd.n5529 9.3005
R17351 gnd.n5541 gnd.n5538 9.3005
R17352 gnd.n5540 gnd.n5539 9.3005
R17353 gnd.n1238 gnd.n1237 9.3005
R17354 gnd.n5567 gnd.n5566 9.3005
R17355 gnd.n5568 gnd.n1236 9.3005
R17356 gnd.n5572 gnd.n5569 9.3005
R17357 gnd.n5571 gnd.n5570 9.3005
R17358 gnd.n1210 gnd.n1209 9.3005
R17359 gnd.n5599 gnd.n5598 9.3005
R17360 gnd.n5600 gnd.n1208 9.3005
R17361 gnd.n5610 gnd.n5601 9.3005
R17362 gnd.n5609 gnd.n5602 9.3005
R17363 gnd.n5655 gnd.n5647 9.3005
R17364 gnd.n5654 gnd.n5648 9.3005
R17365 gnd.n5651 gnd.n5650 9.3005
R17366 gnd.n5649 gnd.n272 9.3005
R17367 gnd.n6760 gnd.n273 9.3005
R17368 gnd.n6759 gnd.n274 9.3005
R17369 gnd.n6758 gnd.n275 9.3005
R17370 gnd.n278 gnd.n276 9.3005
R17371 gnd.n6754 gnd.n279 9.3005
R17372 gnd.n6753 gnd.n6752 9.3005
R17373 gnd.n3926 gnd.n3925 9.3005
R17374 gnd.n3637 gnd.n3633 9.3005
R17375 gnd.n3636 gnd.n3635 9.3005
R17376 gnd.n3634 gnd.n2084 9.3005
R17377 gnd.n3815 gnd.n2085 9.3005
R17378 gnd.n3816 gnd.n2083 9.3005
R17379 gnd.n3819 gnd.n3818 9.3005
R17380 gnd.n3820 gnd.n2082 9.3005
R17381 gnd.n3823 gnd.n3822 9.3005
R17382 gnd.n3821 gnd.n2074 9.3005
R17383 gnd.n3843 gnd.n2075 9.3005
R17384 gnd.n3842 gnd.n2076 9.3005
R17385 gnd.n3841 gnd.n2077 9.3005
R17386 gnd.n2066 gnd.n2065 9.3005
R17387 gnd.n3876 gnd.n3875 9.3005
R17388 gnd.n3877 gnd.n2064 9.3005
R17389 gnd.n3881 gnd.n3878 9.3005
R17390 gnd.n3880 gnd.n3879 9.3005
R17391 gnd.n2053 gnd.n2052 9.3005
R17392 gnd.n3923 gnd.n3922 9.3005
R17393 gnd.n3924 gnd.n2051 9.3005
R17394 gnd.n3639 gnd.n3638 9.3005
R17395 gnd.n3631 gnd.n3630 9.3005
R17396 gnd.n3627 gnd.n3587 9.3005
R17397 gnd.n3626 gnd.n3623 9.3005
R17398 gnd.n3622 gnd.n3588 9.3005
R17399 gnd.n3621 gnd.n3620 9.3005
R17400 gnd.n3617 gnd.n3589 9.3005
R17401 gnd.n3616 gnd.n3613 9.3005
R17402 gnd.n3612 gnd.n3590 9.3005
R17403 gnd.n3611 gnd.n3610 9.3005
R17404 gnd.n3607 gnd.n3591 9.3005
R17405 gnd.n3606 gnd.n3603 9.3005
R17406 gnd.n3602 gnd.n3592 9.3005
R17407 gnd.n3601 gnd.n3600 9.3005
R17408 gnd.n3597 gnd.n3593 9.3005
R17409 gnd.n3596 gnd.n3594 9.3005
R17410 gnd.n2103 gnd.n2102 9.3005
R17411 gnd.n3789 gnd.n3788 9.3005
R17412 gnd.n3632 gnd.n3586 9.3005
R17413 gnd.n3641 gnd.n3640 9.3005
R17414 gnd.n3801 gnd.n3800 9.3005
R17415 gnd.n3799 gnd.n2101 9.3005
R17416 gnd.n3798 gnd.n3797 9.3005
R17417 gnd.n3796 gnd.n3791 9.3005
R17418 gnd.n3794 gnd.n3793 9.3005
R17419 gnd.n3792 gnd.n846 9.3005
R17420 gnd.n5938 gnd.n847 9.3005
R17421 gnd.n5937 gnd.n848 9.3005
R17422 gnd.n5936 gnd.n849 9.3005
R17423 gnd.n867 gnd.n850 9.3005
R17424 gnd.n5926 gnd.n868 9.3005
R17425 gnd.n5925 gnd.n869 9.3005
R17426 gnd.n5924 gnd.n870 9.3005
R17427 gnd.n888 gnd.n871 9.3005
R17428 gnd.n5914 gnd.n889 9.3005
R17429 gnd.n5913 gnd.n890 9.3005
R17430 gnd.n5912 gnd.n891 9.3005
R17431 gnd.n3912 gnd.n892 9.3005
R17432 gnd.n3914 gnd.n3913 9.3005
R17433 gnd.n3915 gnd.n2032 9.3005
R17434 gnd.n3932 gnd.n2031 9.3005
R17435 gnd.n3940 gnd.n3933 9.3005
R17436 gnd.n3939 gnd.n3934 9.3005
R17437 gnd.n3938 gnd.n3936 9.3005
R17438 gnd.n3935 gnd.n915 9.3005
R17439 gnd.n5900 gnd.n916 9.3005
R17440 gnd.n5899 gnd.n917 9.3005
R17441 gnd.n5898 gnd.n918 9.3005
R17442 gnd.n934 gnd.n919 9.3005
R17443 gnd.n5888 gnd.n935 9.3005
R17444 gnd.n5887 gnd.n936 9.3005
R17445 gnd.n5886 gnd.n937 9.3005
R17446 gnd.n956 gnd.n938 9.3005
R17447 gnd.n5876 gnd.n957 9.3005
R17448 gnd.n5875 gnd.n958 9.3005
R17449 gnd.n5874 gnd.n959 9.3005
R17450 gnd.n977 gnd.n960 9.3005
R17451 gnd.n5864 gnd.n978 9.3005
R17452 gnd.n5863 gnd.n979 9.3005
R17453 gnd.n5862 gnd.n980 9.3005
R17454 gnd.n998 gnd.n981 9.3005
R17455 gnd.n5852 gnd.n5851 9.3005
R17456 gnd.n3790 gnd.n2100 9.3005
R17457 gnd.n1812 gnd.n1808 9.3005
R17458 gnd.n1845 gnd.n1842 9.3005
R17459 gnd.n1846 gnd.n1841 9.3005
R17460 gnd.n1849 gnd.n1840 9.3005
R17461 gnd.n1850 gnd.n1839 9.3005
R17462 gnd.n1853 gnd.n1838 9.3005
R17463 gnd.n1854 gnd.n1837 9.3005
R17464 gnd.n1857 gnd.n1836 9.3005
R17465 gnd.n1858 gnd.n1835 9.3005
R17466 gnd.n1861 gnd.n1834 9.3005
R17467 gnd.n1862 gnd.n1833 9.3005
R17468 gnd.n1865 gnd.n1832 9.3005
R17469 gnd.n1866 gnd.n1831 9.3005
R17470 gnd.n1867 gnd.n1830 9.3005
R17471 gnd.n1829 gnd.n1826 9.3005
R17472 gnd.n1828 gnd.n1827 9.3005
R17473 gnd.n4343 gnd.n4342 9.3005
R17474 gnd.n1814 gnd.n1813 9.3005
R17475 gnd.n1873 gnd.n1871 9.3005
R17476 gnd.n4335 gnd.n1874 9.3005
R17477 gnd.n4334 gnd.n1875 9.3005
R17478 gnd.n4333 gnd.n1876 9.3005
R17479 gnd.n1880 gnd.n1877 9.3005
R17480 gnd.n4328 gnd.n1881 9.3005
R17481 gnd.n4327 gnd.n1882 9.3005
R17482 gnd.n4326 gnd.n1883 9.3005
R17483 gnd.n1887 gnd.n1884 9.3005
R17484 gnd.n4321 gnd.n1888 9.3005
R17485 gnd.n4320 gnd.n1889 9.3005
R17486 gnd.n4319 gnd.n1890 9.3005
R17487 gnd.n1894 gnd.n1891 9.3005
R17488 gnd.n4314 gnd.n1895 9.3005
R17489 gnd.n4313 gnd.n1896 9.3005
R17490 gnd.n4312 gnd.n1897 9.3005
R17491 gnd.n1902 gnd.n1900 9.3005
R17492 gnd.n4307 gnd.n4306 9.3005
R17493 gnd.n4344 gnd.n1807 9.3005
R17494 gnd.n3704 gnd.n3703 9.3005
R17495 gnd.n3702 gnd.n3690 9.3005
R17496 gnd.n3701 gnd.n3700 9.3005
R17497 gnd.n3699 gnd.n3691 9.3005
R17498 gnd.n3697 gnd.n3692 9.3005
R17499 gnd.n3696 gnd.n3694 9.3005
R17500 gnd.n3693 gnd.n2080 9.3005
R17501 gnd.n3827 gnd.n2081 9.3005
R17502 gnd.n3828 gnd.n2079 9.3005
R17503 gnd.n3830 gnd.n3829 9.3005
R17504 gnd.n3831 gnd.n2078 9.3005
R17505 gnd.n3837 gnd.n3832 9.3005
R17506 gnd.n3836 gnd.n3833 9.3005
R17507 gnd.n3835 gnd.n3834 9.3005
R17508 gnd.n2063 gnd.n2062 9.3005
R17509 gnd.n3886 gnd.n3885 9.3005
R17510 gnd.n3887 gnd.n2061 9.3005
R17511 gnd.n3891 gnd.n3888 9.3005
R17512 gnd.n3890 gnd.n3889 9.3005
R17513 gnd.n2035 gnd.n2033 9.3005
R17514 gnd.n3931 gnd.n3930 9.3005
R17515 gnd.n2047 gnd.n2034 9.3005
R17516 gnd.n2046 gnd.n2036 9.3005
R17517 gnd.n2045 gnd.n2037 9.3005
R17518 gnd.n2043 gnd.n2038 9.3005
R17519 gnd.n2042 gnd.n2039 9.3005
R17520 gnd.n2041 gnd.n2040 9.3005
R17521 gnd.n2004 gnd.n2003 9.3005
R17522 gnd.n3980 gnd.n3979 9.3005
R17523 gnd.n3981 gnd.n2002 9.3005
R17524 gnd.n3983 gnd.n3982 9.3005
R17525 gnd.n3984 gnd.n2001 9.3005
R17526 gnd.n3988 gnd.n3987 9.3005
R17527 gnd.n3989 gnd.n2000 9.3005
R17528 gnd.n3994 gnd.n3990 9.3005
R17529 gnd.n3995 gnd.n1999 9.3005
R17530 gnd.n3999 gnd.n3998 9.3005
R17531 gnd.n4000 gnd.n1998 9.3005
R17532 gnd.n4003 gnd.n4002 9.3005
R17533 gnd.n4001 gnd.n1904 9.3005
R17534 gnd.n4303 gnd.n1903 9.3005
R17535 gnd.n4305 gnd.n4304 9.3005
R17536 gnd.n3705 gnd.n3688 9.3005
R17537 gnd.n3712 gnd.n3711 9.3005
R17538 gnd.n3713 gnd.n3682 9.3005
R17539 gnd.n3716 gnd.n3681 9.3005
R17540 gnd.n3717 gnd.n3680 9.3005
R17541 gnd.n3720 gnd.n3679 9.3005
R17542 gnd.n3721 gnd.n3678 9.3005
R17543 gnd.n3724 gnd.n3677 9.3005
R17544 gnd.n3725 gnd.n3676 9.3005
R17545 gnd.n3728 gnd.n3675 9.3005
R17546 gnd.n3729 gnd.n3674 9.3005
R17547 gnd.n3732 gnd.n3673 9.3005
R17548 gnd.n3733 gnd.n3672 9.3005
R17549 gnd.n3736 gnd.n3671 9.3005
R17550 gnd.n3737 gnd.n3670 9.3005
R17551 gnd.n3740 gnd.n3669 9.3005
R17552 gnd.n3741 gnd.n3668 9.3005
R17553 gnd.n3744 gnd.n3667 9.3005
R17554 gnd.n3745 gnd.n3666 9.3005
R17555 gnd.n3748 gnd.n3665 9.3005
R17556 gnd.n3750 gnd.n3662 9.3005
R17557 gnd.n3753 gnd.n3661 9.3005
R17558 gnd.n3754 gnd.n3660 9.3005
R17559 gnd.n3757 gnd.n3659 9.3005
R17560 gnd.n3758 gnd.n3658 9.3005
R17561 gnd.n3761 gnd.n3657 9.3005
R17562 gnd.n3762 gnd.n3656 9.3005
R17563 gnd.n3765 gnd.n3655 9.3005
R17564 gnd.n3766 gnd.n3654 9.3005
R17565 gnd.n3769 gnd.n3653 9.3005
R17566 gnd.n3770 gnd.n3652 9.3005
R17567 gnd.n3773 gnd.n3651 9.3005
R17568 gnd.n3774 gnd.n3650 9.3005
R17569 gnd.n3777 gnd.n3649 9.3005
R17570 gnd.n3779 gnd.n3648 9.3005
R17571 gnd.n3780 gnd.n3647 9.3005
R17572 gnd.n3781 gnd.n3646 9.3005
R17573 gnd.n3782 gnd.n3645 9.3005
R17574 gnd.n3710 gnd.n3687 9.3005
R17575 gnd.n3709 gnd.n3708 9.3005
R17576 gnd.n3806 gnd.n3805 9.3005
R17577 gnd.n3807 gnd.n2091 9.3005
R17578 gnd.n3810 gnd.n3809 9.3005
R17579 gnd.n3808 gnd.n834 9.3005
R17580 gnd.n5944 gnd.n835 9.3005
R17581 gnd.n5943 gnd.n836 9.3005
R17582 gnd.n5942 gnd.n837 9.3005
R17583 gnd.n856 gnd.n838 9.3005
R17584 gnd.n5932 gnd.n857 9.3005
R17585 gnd.n5931 gnd.n858 9.3005
R17586 gnd.n5930 gnd.n859 9.3005
R17587 gnd.n878 gnd.n860 9.3005
R17588 gnd.n5920 gnd.n879 9.3005
R17589 gnd.n5919 gnd.n880 9.3005
R17590 gnd.n5918 gnd.n881 9.3005
R17591 gnd.n906 gnd.n900 9.3005
R17592 gnd.n5894 gnd.n925 9.3005
R17593 gnd.n5893 gnd.n926 9.3005
R17594 gnd.n5892 gnd.n927 9.3005
R17595 gnd.n945 gnd.n928 9.3005
R17596 gnd.n5882 gnd.n946 9.3005
R17597 gnd.n5881 gnd.n947 9.3005
R17598 gnd.n5880 gnd.n948 9.3005
R17599 gnd.n966 gnd.n949 9.3005
R17600 gnd.n5870 gnd.n967 9.3005
R17601 gnd.n5869 gnd.n968 9.3005
R17602 gnd.n5868 gnd.n969 9.3005
R17603 gnd.n988 gnd.n970 9.3005
R17604 gnd.n5858 gnd.n989 9.3005
R17605 gnd.n5857 gnd.n990 9.3005
R17606 gnd.n5856 gnd.n991 9.3005
R17607 gnd.n2093 gnd.n2092 9.3005
R17608 gnd.n5905 gnd.n5904 9.3005
R17609 gnd.n3852 gnd.n3849 9.3005
R17610 gnd.n3856 gnd.n3855 9.3005
R17611 gnd.n3857 gnd.n3848 9.3005
R17612 gnd.n3859 gnd.n3858 9.3005
R17613 gnd.n2072 gnd.n2071 9.3005
R17614 gnd.n3864 gnd.n3863 9.3005
R17615 gnd.n3865 gnd.n2070 9.3005
R17616 gnd.n3870 gnd.n3866 9.3005
R17617 gnd.n3869 gnd.n3867 9.3005
R17618 gnd.n3851 gnd.n3850 9.3005
R17619 gnd.n5950 gnd.n824 9.3005
R17620 gnd.n5951 gnd.n823 9.3005
R17621 gnd.n822 gnd.n818 9.3005
R17622 gnd.n5957 gnd.n817 9.3005
R17623 gnd.n5958 gnd.n816 9.3005
R17624 gnd.n5959 gnd.n815 9.3005
R17625 gnd.n814 gnd.n810 9.3005
R17626 gnd.n5965 gnd.n809 9.3005
R17627 gnd.n5966 gnd.n808 9.3005
R17628 gnd.n5967 gnd.n807 9.3005
R17629 gnd.n806 gnd.n802 9.3005
R17630 gnd.n5973 gnd.n801 9.3005
R17631 gnd.n5974 gnd.n800 9.3005
R17632 gnd.n5975 gnd.n799 9.3005
R17633 gnd.n798 gnd.n794 9.3005
R17634 gnd.n5981 gnd.n793 9.3005
R17635 gnd.n5982 gnd.n792 9.3005
R17636 gnd.n5983 gnd.n791 9.3005
R17637 gnd.n790 gnd.n786 9.3005
R17638 gnd.n5989 gnd.n785 9.3005
R17639 gnd.n5990 gnd.n784 9.3005
R17640 gnd.n5991 gnd.n783 9.3005
R17641 gnd.n782 gnd.n778 9.3005
R17642 gnd.n5997 gnd.n777 9.3005
R17643 gnd.n5998 gnd.n776 9.3005
R17644 gnd.n5999 gnd.n775 9.3005
R17645 gnd.n774 gnd.n770 9.3005
R17646 gnd.n6005 gnd.n769 9.3005
R17647 gnd.n6006 gnd.n768 9.3005
R17648 gnd.n6007 gnd.n767 9.3005
R17649 gnd.n766 gnd.n762 9.3005
R17650 gnd.n6013 gnd.n761 9.3005
R17651 gnd.n6014 gnd.n760 9.3005
R17652 gnd.n6015 gnd.n759 9.3005
R17653 gnd.n758 gnd.n754 9.3005
R17654 gnd.n6021 gnd.n753 9.3005
R17655 gnd.n6022 gnd.n752 9.3005
R17656 gnd.n6023 gnd.n751 9.3005
R17657 gnd.n750 gnd.n746 9.3005
R17658 gnd.n6029 gnd.n745 9.3005
R17659 gnd.n6030 gnd.n744 9.3005
R17660 gnd.n6031 gnd.n743 9.3005
R17661 gnd.n742 gnd.n738 9.3005
R17662 gnd.n6037 gnd.n737 9.3005
R17663 gnd.n6038 gnd.n736 9.3005
R17664 gnd.n6039 gnd.n735 9.3005
R17665 gnd.n734 gnd.n730 9.3005
R17666 gnd.n6045 gnd.n729 9.3005
R17667 gnd.n6046 gnd.n728 9.3005
R17668 gnd.n6047 gnd.n727 9.3005
R17669 gnd.n726 gnd.n722 9.3005
R17670 gnd.n6053 gnd.n721 9.3005
R17671 gnd.n6054 gnd.n720 9.3005
R17672 gnd.n6055 gnd.n719 9.3005
R17673 gnd.n718 gnd.n714 9.3005
R17674 gnd.n6061 gnd.n713 9.3005
R17675 gnd.n6062 gnd.n712 9.3005
R17676 gnd.n6063 gnd.n711 9.3005
R17677 gnd.n710 gnd.n706 9.3005
R17678 gnd.n6069 gnd.n705 9.3005
R17679 gnd.n6070 gnd.n704 9.3005
R17680 gnd.n6071 gnd.n703 9.3005
R17681 gnd.n702 gnd.n698 9.3005
R17682 gnd.n6077 gnd.n697 9.3005
R17683 gnd.n6078 gnd.n696 9.3005
R17684 gnd.n6079 gnd.n695 9.3005
R17685 gnd.n694 gnd.n690 9.3005
R17686 gnd.n6085 gnd.n689 9.3005
R17687 gnd.n6086 gnd.n688 9.3005
R17688 gnd.n6087 gnd.n687 9.3005
R17689 gnd.n686 gnd.n682 9.3005
R17690 gnd.n6093 gnd.n681 9.3005
R17691 gnd.n6094 gnd.n680 9.3005
R17692 gnd.n6095 gnd.n679 9.3005
R17693 gnd.n678 gnd.n674 9.3005
R17694 gnd.n6101 gnd.n673 9.3005
R17695 gnd.n6102 gnd.n672 9.3005
R17696 gnd.n6103 gnd.n671 9.3005
R17697 gnd.n670 gnd.n666 9.3005
R17698 gnd.n6109 gnd.n665 9.3005
R17699 gnd.n6110 gnd.n664 9.3005
R17700 gnd.n6111 gnd.n663 9.3005
R17701 gnd.n659 gnd.n658 9.3005
R17702 gnd.n6118 gnd.n6117 9.3005
R17703 gnd.n5949 gnd.n825 9.3005
R17704 gnd.n5039 gnd.n5038 9.3005
R17705 gnd.n5019 gnd.n5017 9.3005
R17706 gnd.n5046 gnd.n5045 9.3005
R17707 gnd.n5013 gnd.n5012 9.3005
R17708 gnd.n5058 gnd.n5057 9.3005
R17709 gnd.n5010 gnd.n5008 9.3005
R17710 gnd.n5065 gnd.n5064 9.3005
R17711 gnd.n5004 gnd.n5003 9.3005
R17712 gnd.n5077 gnd.n5076 9.3005
R17713 gnd.n5001 gnd.n4999 9.3005
R17714 gnd.n5084 gnd.n5083 9.3005
R17715 gnd.n4995 gnd.n4994 9.3005
R17716 gnd.n5096 gnd.n5095 9.3005
R17717 gnd.n4992 gnd.n4990 9.3005
R17718 gnd.n5105 gnd.n5104 9.3005
R17719 gnd.n5103 gnd.n4984 9.3005
R17720 gnd.n5114 gnd.n4983 9.3005
R17721 gnd.n5117 gnd.n5116 9.3005
R17722 gnd.n5022 gnd.n5021 9.3005
R17723 gnd.n5107 gnd.n5106 9.3005
R17724 gnd.n5094 gnd.n4989 9.3005
R17725 gnd.n5093 gnd.n5092 9.3005
R17726 gnd.n5000 gnd.n4996 9.3005
R17727 gnd.n5086 gnd.n5085 9.3005
R17728 gnd.n5075 gnd.n4998 9.3005
R17729 gnd.n5074 gnd.n5073 9.3005
R17730 gnd.n5009 gnd.n5005 9.3005
R17731 gnd.n5067 gnd.n5066 9.3005
R17732 gnd.n5056 gnd.n5007 9.3005
R17733 gnd.n5055 gnd.n5054 9.3005
R17734 gnd.n5018 gnd.n5014 9.3005
R17735 gnd.n5048 gnd.n5047 9.3005
R17736 gnd.n5037 gnd.n5016 9.3005
R17737 gnd.n5036 gnd.n5035 9.3005
R17738 gnd.n5024 gnd.n5023 9.3005
R17739 gnd.n4991 gnd.n4987 9.3005
R17740 gnd.n5113 gnd.n5112 9.3005
R17741 gnd.n4981 gnd.n4980 9.3005
R17742 gnd.n5124 gnd.n5123 9.3005
R17743 gnd.n5125 gnd.n4979 9.3005
R17744 gnd.n5127 gnd.n5126 9.3005
R17745 gnd.n4977 gnd.n4976 9.3005
R17746 gnd.n5137 gnd.n5136 9.3005
R17747 gnd.n5138 gnd.n4975 9.3005
R17748 gnd.n5140 gnd.n5139 9.3005
R17749 gnd.n4973 gnd.n4972 9.3005
R17750 gnd.n5146 gnd.n5145 9.3005
R17751 gnd.n4276 gnd.n1927 9.3005
R17752 gnd.n4275 gnd.n4274 9.3005
R17753 gnd.n4273 gnd.n1931 9.3005
R17754 gnd.n4272 gnd.n4271 9.3005
R17755 gnd.n4270 gnd.n1932 9.3005
R17756 gnd.n4269 gnd.n4268 9.3005
R17757 gnd.n4267 gnd.n1936 9.3005
R17758 gnd.n4266 gnd.n4265 9.3005
R17759 gnd.n4264 gnd.n1937 9.3005
R17760 gnd.n4263 gnd.n4262 9.3005
R17761 gnd.n4261 gnd.n1941 9.3005
R17762 gnd.n4260 gnd.n4259 9.3005
R17763 gnd.n4258 gnd.n1942 9.3005
R17764 gnd.n4257 gnd.n4256 9.3005
R17765 gnd.n4255 gnd.n4247 9.3005
R17766 gnd.n4254 gnd.n4253 9.3005
R17767 gnd.n4252 gnd.n4248 9.3005
R17768 gnd.n1643 gnd.n1642 9.3005
R17769 gnd.n4490 gnd.n4489 9.3005
R17770 gnd.n4491 gnd.n1641 9.3005
R17771 gnd.n4493 gnd.n4492 9.3005
R17772 gnd.n1623 gnd.n1622 9.3005
R17773 gnd.n4523 gnd.n4522 9.3005
R17774 gnd.n4524 gnd.n1621 9.3005
R17775 gnd.n4526 gnd.n4525 9.3005
R17776 gnd.n1597 gnd.n1596 9.3005
R17777 gnd.n4568 gnd.n4567 9.3005
R17778 gnd.n4569 gnd.n1594 9.3005
R17779 gnd.n4573 gnd.n4572 9.3005
R17780 gnd.n4571 gnd.n1595 9.3005
R17781 gnd.n4570 gnd.n1583 9.3005
R17782 gnd.n1581 gnd.n1580 9.3005
R17783 gnd.n4598 gnd.n4597 9.3005
R17784 gnd.n4599 gnd.n1579 9.3005
R17785 gnd.n4601 gnd.n4600 9.3005
R17786 gnd.n1555 gnd.n1553 9.3005
R17787 gnd.n4649 gnd.n4648 9.3005
R17788 gnd.n4647 gnd.n1554 9.3005
R17789 gnd.n4646 gnd.n4645 9.3005
R17790 gnd.n1532 gnd.n1530 9.3005
R17791 gnd.n4705 gnd.n4704 9.3005
R17792 gnd.n4703 gnd.n1531 9.3005
R17793 gnd.n4702 gnd.n4701 9.3005
R17794 gnd.n4700 gnd.n1533 9.3005
R17795 gnd.n4699 gnd.n4698 9.3005
R17796 gnd.n4697 gnd.n4688 9.3005
R17797 gnd.n4696 gnd.n4695 9.3005
R17798 gnd.n4694 gnd.n4689 9.3005
R17799 gnd.n4693 gnd.n4692 9.3005
R17800 gnd.n1470 gnd.n1469 9.3005
R17801 gnd.n4813 gnd.n4812 9.3005
R17802 gnd.n4814 gnd.n1467 9.3005
R17803 gnd.n4817 gnd.n4816 9.3005
R17804 gnd.n4815 gnd.n1468 9.3005
R17805 gnd.n1442 gnd.n1441 9.3005
R17806 gnd.n4852 gnd.n4851 9.3005
R17807 gnd.n4853 gnd.n1439 9.3005
R17808 gnd.n4872 gnd.n4871 9.3005
R17809 gnd.n4870 gnd.n1440 9.3005
R17810 gnd.n4869 gnd.n4868 9.3005
R17811 gnd.n4867 gnd.n4854 9.3005
R17812 gnd.n4866 gnd.n4865 9.3005
R17813 gnd.n4864 gnd.n4861 9.3005
R17814 gnd.n4863 gnd.n4862 9.3005
R17815 gnd.n1391 gnd.n1390 9.3005
R17816 gnd.n4943 gnd.n4942 9.3005
R17817 gnd.n4944 gnd.n1389 9.3005
R17818 gnd.n4947 gnd.n4946 9.3005
R17819 gnd.n4945 gnd.n1387 9.3005
R17820 gnd.n4952 gnd.n1386 9.3005
R17821 gnd.n4954 gnd.n4953 9.3005
R17822 gnd.n4955 gnd.n1385 9.3005
R17823 gnd.n4957 gnd.n4956 9.3005
R17824 gnd.n4960 gnd.n1384 9.3005
R17825 gnd.n4962 gnd.n4961 9.3005
R17826 gnd.n4963 gnd.n1383 9.3005
R17827 gnd.n4965 gnd.n4964 9.3005
R17828 gnd.n4968 gnd.n1382 9.3005
R17829 gnd.n4970 gnd.n4969 9.3005
R17830 gnd.n4971 gnd.n1380 9.3005
R17831 gnd.n5149 gnd.n5148 9.3005
R17832 gnd.n5147 gnd.n1381 9.3005
R17833 gnd.n4278 gnd.n4277 9.3005
R17834 gnd.n4281 gnd.n4280 9.3005
R17835 gnd.n4282 gnd.n1922 9.3005
R17836 gnd.n4284 gnd.n4283 9.3005
R17837 gnd.n4286 gnd.n4285 9.3005
R17838 gnd.n4287 gnd.n1915 9.3005
R17839 gnd.n4289 gnd.n4288 9.3005
R17840 gnd.n4290 gnd.n1914 9.3005
R17841 gnd.n4292 gnd.n4291 9.3005
R17842 gnd.n4293 gnd.n1908 9.3005
R17843 gnd.n4279 gnd.n1926 9.3005
R17844 gnd.n2019 gnd.n2018 9.3005
R17845 gnd.n3951 gnd.n3950 9.3005
R17846 gnd.n3952 gnd.n2017 9.3005
R17847 gnd.n3954 gnd.n3953 9.3005
R17848 gnd.n2007 gnd.n2006 9.3005
R17849 gnd.n3972 gnd.n3971 9.3005
R17850 gnd.n3973 gnd.n2005 9.3005
R17851 gnd.n3975 gnd.n3974 9.3005
R17852 gnd.n1991 gnd.n1989 9.3005
R17853 gnd.n4020 gnd.n4019 9.3005
R17854 gnd.n4018 gnd.n1990 9.3005
R17855 gnd.n4017 gnd.n4016 9.3005
R17856 gnd.n4015 gnd.n1992 9.3005
R17857 gnd.n4014 gnd.n4013 9.3005
R17858 gnd.n4012 gnd.n1995 9.3005
R17859 gnd.n4011 gnd.n4010 9.3005
R17860 gnd.n4009 gnd.n1996 9.3005
R17861 gnd.n4008 gnd.n4007 9.3005
R17862 gnd.n1907 gnd.n1905 9.3005
R17863 gnd.n4299 gnd.n4298 9.3005
R17864 gnd.n4297 gnd.n1906 9.3005
R17865 gnd.n4295 gnd.n4294 9.3005
R17866 gnd.n1910 gnd.n1909 9.3005
R17867 gnd.n4145 gnd.n4144 9.3005
R17868 gnd.n4147 gnd.n4146 9.3005
R17869 gnd.n4125 gnd.n4124 9.3005
R17870 gnd.n4153 gnd.n4152 9.3005
R17871 gnd.n4155 gnd.n4154 9.3005
R17872 gnd.n4115 gnd.n4114 9.3005
R17873 gnd.n4161 gnd.n4160 9.3005
R17874 gnd.n4163 gnd.n4162 9.3005
R17875 gnd.n4102 gnd.n4101 9.3005
R17876 gnd.n4169 gnd.n4168 9.3005
R17877 gnd.n4171 gnd.n4170 9.3005
R17878 gnd.n4092 gnd.n4091 9.3005
R17879 gnd.n4177 gnd.n4176 9.3005
R17880 gnd.n4179 gnd.n4178 9.3005
R17881 gnd.n4077 gnd.n4075 9.3005
R17882 gnd.n4185 gnd.n4184 9.3005
R17883 gnd.n4186 gnd.n4074 9.3005
R17884 gnd.n4079 gnd.n1000 9.3005
R17885 gnd.n4078 gnd.n4076 9.3005
R17886 gnd.n4183 gnd.n4182 9.3005
R17887 gnd.n4181 gnd.n4180 9.3005
R17888 gnd.n4087 gnd.n4086 9.3005
R17889 gnd.n4175 gnd.n4174 9.3005
R17890 gnd.n4173 gnd.n4172 9.3005
R17891 gnd.n4098 gnd.n4097 9.3005
R17892 gnd.n4167 gnd.n4166 9.3005
R17893 gnd.n4165 gnd.n4164 9.3005
R17894 gnd.n4109 gnd.n4108 9.3005
R17895 gnd.n4159 gnd.n4158 9.3005
R17896 gnd.n4157 gnd.n4156 9.3005
R17897 gnd.n4121 gnd.n4120 9.3005
R17898 gnd.n4151 gnd.n4150 9.3005
R17899 gnd.n4149 gnd.n4148 9.3005
R17900 gnd.n4134 gnd.n4133 9.3005
R17901 gnd.n4143 gnd.n4142 9.3005
R17902 gnd.n5846 gnd.n1001 9.3005
R17903 gnd.n5845 gnd.n5844 9.3005
R17904 gnd.n5843 gnd.n1005 9.3005
R17905 gnd.n5842 gnd.n5841 9.3005
R17906 gnd.n5840 gnd.n1006 9.3005
R17907 gnd.n5839 gnd.n5838 9.3005
R17908 gnd.n5837 gnd.n1010 9.3005
R17909 gnd.n5836 gnd.n5835 9.3005
R17910 gnd.n5834 gnd.n1011 9.3005
R17911 gnd.n5833 gnd.n5832 9.3005
R17912 gnd.n5831 gnd.n1015 9.3005
R17913 gnd.n5830 gnd.n5829 9.3005
R17914 gnd.n5828 gnd.n1016 9.3005
R17915 gnd.n5827 gnd.n5826 9.3005
R17916 gnd.n5825 gnd.n1020 9.3005
R17917 gnd.n5824 gnd.n5823 9.3005
R17918 gnd.n5822 gnd.n1021 9.3005
R17919 gnd.n5821 gnd.n5820 9.3005
R17920 gnd.n5819 gnd.n1025 9.3005
R17921 gnd.n5818 gnd.n5817 9.3005
R17922 gnd.n5816 gnd.n1026 9.3005
R17923 gnd.n5815 gnd.n5814 9.3005
R17924 gnd.n5813 gnd.n1030 9.3005
R17925 gnd.n5812 gnd.n5811 9.3005
R17926 gnd.n5810 gnd.n1031 9.3005
R17927 gnd.n5809 gnd.n5808 9.3005
R17928 gnd.n5807 gnd.n1035 9.3005
R17929 gnd.n5806 gnd.n5805 9.3005
R17930 gnd.n5804 gnd.n1036 9.3005
R17931 gnd.n5803 gnd.n5802 9.3005
R17932 gnd.n5801 gnd.n1040 9.3005
R17933 gnd.n5800 gnd.n5799 9.3005
R17934 gnd.n5798 gnd.n1041 9.3005
R17935 gnd.n5797 gnd.n5796 9.3005
R17936 gnd.n5795 gnd.n1045 9.3005
R17937 gnd.n5794 gnd.n5793 9.3005
R17938 gnd.n5792 gnd.n1046 9.3005
R17939 gnd.n5791 gnd.n5790 9.3005
R17940 gnd.n5789 gnd.n1050 9.3005
R17941 gnd.n5788 gnd.n5787 9.3005
R17942 gnd.n5786 gnd.n1051 9.3005
R17943 gnd.n5785 gnd.n5784 9.3005
R17944 gnd.n5783 gnd.n1055 9.3005
R17945 gnd.n5782 gnd.n5781 9.3005
R17946 gnd.n5780 gnd.n1056 9.3005
R17947 gnd.n5779 gnd.n5778 9.3005
R17948 gnd.n5777 gnd.n1060 9.3005
R17949 gnd.n5776 gnd.n5775 9.3005
R17950 gnd.n5774 gnd.n1061 9.3005
R17951 gnd.n5773 gnd.n5772 9.3005
R17952 gnd.n5771 gnd.n1065 9.3005
R17953 gnd.n5770 gnd.n5769 9.3005
R17954 gnd.n5768 gnd.n1066 9.3005
R17955 gnd.n5767 gnd.n5766 9.3005
R17956 gnd.n5765 gnd.n1070 9.3005
R17957 gnd.n5764 gnd.n5763 9.3005
R17958 gnd.n5762 gnd.n1071 9.3005
R17959 gnd.n5761 gnd.n5760 9.3005
R17960 gnd.n5759 gnd.n1075 9.3005
R17961 gnd.n5758 gnd.n5757 9.3005
R17962 gnd.n5756 gnd.n1076 9.3005
R17963 gnd.n5755 gnd.n5754 9.3005
R17964 gnd.n5753 gnd.n1080 9.3005
R17965 gnd.n5752 gnd.n5751 9.3005
R17966 gnd.n5750 gnd.n1081 9.3005
R17967 gnd.n5749 gnd.n5748 9.3005
R17968 gnd.n5747 gnd.n1085 9.3005
R17969 gnd.n5746 gnd.n5745 9.3005
R17970 gnd.n5744 gnd.n1086 9.3005
R17971 gnd.n5743 gnd.n5742 9.3005
R17972 gnd.n5741 gnd.n1090 9.3005
R17973 gnd.n5740 gnd.n5739 9.3005
R17974 gnd.n5738 gnd.n1091 9.3005
R17975 gnd.n5737 gnd.n5736 9.3005
R17976 gnd.n5735 gnd.n1095 9.3005
R17977 gnd.n5734 gnd.n5733 9.3005
R17978 gnd.n5732 gnd.n1096 9.3005
R17979 gnd.n5731 gnd.n5730 9.3005
R17980 gnd.n5729 gnd.n1100 9.3005
R17981 gnd.n5728 gnd.n5727 9.3005
R17982 gnd.n5726 gnd.n1101 9.3005
R17983 gnd.n5725 gnd.n1104 9.3005
R17984 gnd.n5848 gnd.n5847 9.3005
R17985 gnd.n1146 gnd.n1144 9.3005
R17986 gnd.n5699 gnd.n5698 9.3005
R17987 gnd.n5697 gnd.n1145 9.3005
R17988 gnd.n5696 gnd.n5695 9.3005
R17989 gnd.n5694 gnd.n1147 9.3005
R17990 gnd.n5693 gnd.n5692 9.3005
R17991 gnd.n5691 gnd.n1151 9.3005
R17992 gnd.n5690 gnd.n5689 9.3005
R17993 gnd.n5688 gnd.n1152 9.3005
R17994 gnd.n5687 gnd.n5686 9.3005
R17995 gnd.n5685 gnd.n1156 9.3005
R17996 gnd.n5684 gnd.n5683 9.3005
R17997 gnd.n5682 gnd.n1157 9.3005
R17998 gnd.n5681 gnd.n5680 9.3005
R17999 gnd.n5679 gnd.n1161 9.3005
R18000 gnd.n5678 gnd.n5677 9.3005
R18001 gnd.n5676 gnd.n1162 9.3005
R18002 gnd.n5675 gnd.n5674 9.3005
R18003 gnd.n5673 gnd.n1166 9.3005
R18004 gnd.n5672 gnd.n5671 9.3005
R18005 gnd.n5670 gnd.n1167 9.3005
R18006 gnd.n5669 gnd.n5668 9.3005
R18007 gnd.n229 gnd.n228 9.3005
R18008 gnd.n6791 gnd.n6790 9.3005
R18009 gnd.n6792 gnd.n227 9.3005
R18010 gnd.n6794 gnd.n6793 9.3005
R18011 gnd.n207 gnd.n206 9.3005
R18012 gnd.n6807 gnd.n6806 9.3005
R18013 gnd.n6808 gnd.n205 9.3005
R18014 gnd.n6810 gnd.n6809 9.3005
R18015 gnd.n192 gnd.n191 9.3005
R18016 gnd.n6823 gnd.n6822 9.3005
R18017 gnd.n6824 gnd.n190 9.3005
R18018 gnd.n6826 gnd.n6825 9.3005
R18019 gnd.n175 gnd.n174 9.3005
R18020 gnd.n6839 gnd.n6838 9.3005
R18021 gnd.n6840 gnd.n172 9.3005
R18022 gnd.n6916 gnd.n6915 9.3005
R18023 gnd.n6914 gnd.n173 9.3005
R18024 gnd.n6913 gnd.n6912 9.3005
R18025 gnd.n6911 gnd.n6841 9.3005
R18026 gnd.n6910 gnd.n6909 9.3005
R18027 gnd.n5027 gnd.n5026 9.3005
R18028 gnd.n6906 gnd.n6843 9.3005
R18029 gnd.n6905 gnd.n6904 9.3005
R18030 gnd.n6903 gnd.n6848 9.3005
R18031 gnd.n6902 gnd.n6901 9.3005
R18032 gnd.n6900 gnd.n6849 9.3005
R18033 gnd.n6899 gnd.n6898 9.3005
R18034 gnd.n6897 gnd.n6856 9.3005
R18035 gnd.n6896 gnd.n6895 9.3005
R18036 gnd.n6894 gnd.n6857 9.3005
R18037 gnd.n6893 gnd.n6892 9.3005
R18038 gnd.n6891 gnd.n6864 9.3005
R18039 gnd.n6890 gnd.n6889 9.3005
R18040 gnd.n6888 gnd.n6865 9.3005
R18041 gnd.n6887 gnd.n6886 9.3005
R18042 gnd.n6885 gnd.n6872 9.3005
R18043 gnd.n6884 gnd.n6883 9.3005
R18044 gnd.n6882 gnd.n6873 9.3005
R18045 gnd.n6881 gnd.n78 9.3005
R18046 gnd.n6908 gnd.n6907 9.3005
R18047 gnd.n5471 gnd.n5470 9.3005
R18048 gnd.n5472 gnd.n1262 9.3005
R18049 gnd.n5475 gnd.n5474 9.3005
R18050 gnd.n5473 gnd.n1263 9.3005
R18051 gnd.n1247 gnd.n1246 9.3005
R18052 gnd.n5557 gnd.n5556 9.3005
R18053 gnd.n5558 gnd.n1244 9.3005
R18054 gnd.n5561 gnd.n5560 9.3005
R18055 gnd.n5559 gnd.n1245 9.3005
R18056 gnd.n1218 gnd.n1217 9.3005
R18057 gnd.n5589 gnd.n5588 9.3005
R18058 gnd.n5590 gnd.n1215 9.3005
R18059 gnd.n5593 gnd.n5592 9.3005
R18060 gnd.n5591 gnd.n1216 9.3005
R18061 gnd.n1192 gnd.n1191 9.3005
R18062 gnd.n5622 gnd.n5621 9.3005
R18063 gnd.n5623 gnd.n1188 9.3005
R18064 gnd.n5626 gnd.n5625 9.3005
R18065 gnd.n5624 gnd.n1190 9.3005
R18066 gnd.n1189 gnd.n51 9.3005
R18067 gnd.n7040 gnd.n52 9.3005
R18068 gnd.n7039 gnd.n7038 9.3005
R18069 gnd.n7037 gnd.n53 9.3005
R18070 gnd.n7036 gnd.n7035 9.3005
R18071 gnd.n7034 gnd.n57 9.3005
R18072 gnd.n7033 gnd.n7032 9.3005
R18073 gnd.n7031 gnd.n58 9.3005
R18074 gnd.n7030 gnd.n7029 9.3005
R18075 gnd.n7028 gnd.n62 9.3005
R18076 gnd.n7027 gnd.n7026 9.3005
R18077 gnd.n7025 gnd.n63 9.3005
R18078 gnd.n7024 gnd.n7023 9.3005
R18079 gnd.n7022 gnd.n67 9.3005
R18080 gnd.n7021 gnd.n7020 9.3005
R18081 gnd.n7019 gnd.n68 9.3005
R18082 gnd.n7018 gnd.n7017 9.3005
R18083 gnd.n7016 gnd.n72 9.3005
R18084 gnd.n7015 gnd.n7014 9.3005
R18085 gnd.n7013 gnd.n73 9.3005
R18086 gnd.n7012 gnd.n7011 9.3005
R18087 gnd.n7010 gnd.n77 9.3005
R18088 gnd.n7009 gnd.n7008 9.3005
R18089 gnd.n1265 gnd.n1264 9.3005
R18090 gnd.t10 gnd.n2295 9.24152
R18091 gnd.n2197 gnd.t172 9.24152
R18092 gnd.n3454 gnd.t168 9.24152
R18093 gnd.n3991 gnd.t45 9.24152
R18094 gnd.t93 gnd.n1251 9.24152
R18095 gnd.t55 gnd.t10 8.92286
R18096 gnd.n4459 gnd.n4458 8.92286
R18097 gnd.n4585 gnd.n1589 8.92286
R18098 gnd.n4630 gnd.n1559 8.92286
R18099 gnd.t248 gnd.n1549 8.92286
R18100 gnd.n4741 gnd.t109 8.92286
R18101 gnd.n4753 gnd.n1493 8.92286
R18102 gnd.n4822 gnd.n4821 8.92286
R18103 gnd.n4924 gnd.n1401 8.92286
R18104 gnd.t205 gnd.n1341 8.92286
R18105 gnd.n3424 gnd.n3399 8.92171
R18106 gnd.n3392 gnd.n3367 8.92171
R18107 gnd.n3360 gnd.n3335 8.92171
R18108 gnd.n3329 gnd.n3304 8.92171
R18109 gnd.n3297 gnd.n3272 8.92171
R18110 gnd.n3265 gnd.n3240 8.92171
R18111 gnd.n3233 gnd.n3208 8.92171
R18112 gnd.n3202 gnd.n3177 8.92171
R18113 gnd.n5214 gnd.n5196 8.72777
R18114 gnd.n2927 gnd.t12 8.60421
R18115 gnd.n2359 gnd.n2347 8.43467
R18116 gnd.n38 gnd.n26 8.43467
R18117 gnd.n3925 gnd.n0 8.41456
R18118 gnd.n7041 gnd.n7040 8.41456
R18119 gnd.t208 gnd.n1674 8.28555
R18120 gnd.t227 gnd.n1646 8.28555
R18121 gnd.n1626 gnd.t125 8.28555
R18122 gnd.n4435 gnd.n1605 8.28555
R18123 gnd.n4622 gnd.t246 8.28555
R18124 gnd.n4651 gnd.n1542 8.28555
R18125 gnd.n4732 gnd.n1507 8.28555
R18126 gnd.n1488 gnd.t249 8.28555
R18127 gnd.n4787 gnd.n1458 8.28555
R18128 gnd.t108 gnd.n1429 8.28555
R18129 gnd.n3425 gnd.n3397 8.14595
R18130 gnd.n3393 gnd.n3365 8.14595
R18131 gnd.n3361 gnd.n3333 8.14595
R18132 gnd.n3330 gnd.n3302 8.14595
R18133 gnd.n3298 gnd.n3270 8.14595
R18134 gnd.n3266 gnd.n3238 8.14595
R18135 gnd.n3234 gnd.n3206 8.14595
R18136 gnd.n3203 gnd.n3175 8.14595
R18137 gnd.n3430 gnd.n3429 7.97301
R18138 gnd.t18 gnd.n2442 7.9669
R18139 gnd.n6882 gnd.n6881 7.75808
R18140 gnd.n5112 gnd.n4987 7.75808
R18141 gnd.n4142 gnd.n4133 7.75808
R18142 gnd.n3641 gnd.n3586 7.75808
R18143 gnd.n4467 gnd.t154 7.64824
R18144 gnd.n4498 gnd.n4497 7.64824
R18145 gnd.n4435 gnd.n1601 7.64824
R18146 gnd.n4662 gnd.n1542 7.64824
R18147 gnd.n4732 gnd.n1506 7.64824
R18148 gnd.n4787 gnd.n1449 7.64824
R18149 gnd.n4900 gnd.n1417 7.64824
R18150 gnd.n2836 gnd.t24 7.32958
R18151 gnd.n1696 gnd.n1695 7.30353
R18152 gnd.n5213 gnd.n5212 7.30353
R18153 gnd.n2796 gnd.n2515 7.01093
R18154 gnd.n2518 gnd.n2516 7.01093
R18155 gnd.n2806 gnd.n2805 7.01093
R18156 gnd.n2817 gnd.n2499 7.01093
R18157 gnd.n2816 gnd.n2502 7.01093
R18158 gnd.n2827 gnd.n2490 7.01093
R18159 gnd.n2493 gnd.n2491 7.01093
R18160 gnd.n2837 gnd.n2836 7.01093
R18161 gnd.n2847 gnd.n2471 7.01093
R18162 gnd.n2846 gnd.n2474 7.01093
R18163 gnd.n2855 gnd.n2465 7.01093
R18164 gnd.n2867 gnd.n2455 7.01093
R18165 gnd.n2877 gnd.n2440 7.01093
R18166 gnd.n2893 gnd.n2892 7.01093
R18167 gnd.n2442 gnd.n2379 7.01093
R18168 gnd.n2947 gnd.n2380 7.01093
R18169 gnd.n2941 gnd.n2940 7.01093
R18170 gnd.n2429 gnd.n2391 7.01093
R18171 gnd.n2933 gnd.n2402 7.01093
R18172 gnd.n2420 gnd.n2415 7.01093
R18173 gnd.n2927 gnd.n2926 7.01093
R18174 gnd.n2973 gnd.n2330 7.01093
R18175 gnd.n2972 gnd.n2971 7.01093
R18176 gnd.n2984 gnd.n2983 7.01093
R18177 gnd.n2323 gnd.n2315 7.01093
R18178 gnd.n3013 gnd.n2303 7.01093
R18179 gnd.n3012 gnd.n2306 7.01093
R18180 gnd.n3023 gnd.n2295 7.01093
R18181 gnd.n2296 gnd.n2284 7.01093
R18182 gnd.n3034 gnd.n2285 7.01093
R18183 gnd.n3058 gnd.n2276 7.01093
R18184 gnd.n3057 gnd.n2267 7.01093
R18185 gnd.n3081 gnd.n3080 7.01093
R18186 gnd.n3099 gnd.n2248 7.01093
R18187 gnd.n3098 gnd.n2251 7.01093
R18188 gnd.n3109 gnd.n2240 7.01093
R18189 gnd.n2241 gnd.n2228 7.01093
R18190 gnd.n3120 gnd.n2229 7.01093
R18191 gnd.n3147 gnd.n2213 7.01093
R18192 gnd.n3159 gnd.n3158 7.01093
R18193 gnd.n3141 gnd.n2206 7.01093
R18194 gnd.n3170 gnd.n3169 7.01093
R18195 gnd.n3442 gnd.n2194 7.01093
R18196 gnd.n3441 gnd.n2197 7.01093
R18197 gnd.n3454 gnd.n2186 7.01093
R18198 gnd.n2187 gnd.n2179 7.01093
R18199 gnd.n3464 gnd.n2105 7.01093
R18200 gnd.n4585 gnd.n4584 7.01093
R18201 gnd.n4604 gnd.n1559 7.01093
R18202 gnd.n4631 gnd.t248 7.01093
R18203 gnd.t109 gnd.n4740 7.01093
R18204 gnd.n4753 gnd.n4752 7.01093
R18205 gnd.n4822 gnd.n1462 7.01093
R18206 gnd.n4924 gnd.n4923 7.01093
R18207 gnd.n4939 gnd.t205 7.01093
R18208 gnd.n2474 gnd.t23 6.69227
R18209 gnd.n2306 gnd.t55 6.69227
R18210 gnd.n3148 gnd.t17 6.69227
R18211 gnd.n1646 gnd.t121 6.69227
R18212 gnd.n4859 gnd.t274 6.69227
R18213 gnd.n5343 gnd.n5342 6.5566
R18214 gnd.n1802 gnd.n1801 6.5566
R18215 gnd.n4355 gnd.n1737 6.5566
R18216 gnd.n5221 gnd.n5220 6.5566
R18217 gnd.n3079 gnd.n2248 6.37362
R18218 gnd.n4449 gnd.n4448 6.37362
R18219 gnd.n4537 gnd.n4536 6.37362
R18220 gnd.n4549 gnd.t66 6.37362
R18221 gnd.n4670 gnd.n1536 6.37362
R18222 gnd.n4682 gnd.n1523 6.37362
R18223 gnd.n4759 gnd.t106 6.37362
R18224 gnd.n4848 gnd.n1445 6.37362
R18225 gnd.n4772 gnd.n1432 6.37362
R18226 gnd.n4283 gnd.n1921 6.20656
R18227 gnd.n6971 gnd.n6968 6.20656
R18228 gnd.n3749 gnd.n3748 6.20656
R18229 gnd.n5135 gnd.n4975 6.20656
R18230 gnd.t53 gnd.n2903 6.05496
R18231 gnd.n2904 gnd.t21 6.05496
R18232 gnd.t251 gnd.n2330 6.05496
R18233 gnd.t20 gnd.n3068 6.05496
R18234 gnd.n3427 gnd.n3397 5.81868
R18235 gnd.n3395 gnd.n3365 5.81868
R18236 gnd.n3363 gnd.n3333 5.81868
R18237 gnd.n3332 gnd.n3302 5.81868
R18238 gnd.n3300 gnd.n3270 5.81868
R18239 gnd.n3268 gnd.n3238 5.81868
R18240 gnd.n3236 gnd.n3206 5.81868
R18241 gnd.n3205 gnd.n3175 5.81868
R18242 gnd.n1676 gnd.n1665 5.73631
R18243 gnd.n4467 gnd.n1660 5.73631
R18244 gnd.n4548 gnd.n1572 5.73631
R18245 gnd.n1573 gnd.n1565 5.73631
R18246 gnd.n1489 gnd.n1479 5.73631
R18247 gnd.n4760 gnd.n1481 5.73631
R18248 gnd.n4940 gnd.n1393 5.73631
R18249 gnd.n5192 gnd.n1341 5.73631
R18250 gnd.n5352 gnd.n1292 5.62001
R18251 gnd.n4350 gnd.n1806 5.62001
R18252 gnd.n4351 gnd.n4350 5.62001
R18253 gnd.n5352 gnd.n1293 5.62001
R18254 gnd.n2655 gnd.n2650 5.4308
R18255 gnd.n3472 gnd.n2172 5.4308
R18256 gnd.n2971 gnd.t19 5.41765
R18257 gnd.t11 gnd.n2994 5.41765
R18258 gnd.t260 gnd.n2260 5.41765
R18259 gnd.t119 gnd.n4528 5.41765
R18260 gnd.n4779 gnd.t103 5.41765
R18261 gnd.n1647 gnd.t227 5.09899
R18262 gnd.n4518 gnd.n1626 5.09899
R18263 gnd.n4530 gnd.n4529 5.09899
R18264 gnd.n4575 gnd.t253 5.09899
R18265 gnd.n4591 gnd.t66 5.09899
R18266 gnd.n4708 gnd.n1527 5.09899
R18267 gnd.n4716 gnd.n1520 5.09899
R18268 gnd.t106 gnd.n1472 5.09899
R18269 gnd.n4819 gnd.t76 5.09899
R18270 gnd.n4875 gnd.n1436 5.09899
R18271 gnd.n4884 gnd.n1429 5.09899
R18272 gnd.n3425 gnd.n3424 5.04292
R18273 gnd.n3393 gnd.n3392 5.04292
R18274 gnd.n3361 gnd.n3360 5.04292
R18275 gnd.n3330 gnd.n3329 5.04292
R18276 gnd.n3298 gnd.n3297 5.04292
R18277 gnd.n3266 gnd.n3265 5.04292
R18278 gnd.n3234 gnd.n3233 5.04292
R18279 gnd.n3203 gnd.n3202 5.04292
R18280 gnd.n2371 gnd.n2370 4.82753
R18281 gnd.n50 gnd.n49 4.82753
R18282 gnd.n2934 gnd.t14 4.78034
R18283 gnd.n2285 gnd.t15 4.78034
R18284 gnd.t269 gnd.n4216 4.78034
R18285 gnd.n5170 gnd.t41 4.78034
R18286 gnd.n2376 gnd.n2373 4.74817
R18287 gnd.n2426 gnd.n2336 4.74817
R18288 gnd.n2413 gnd.n2335 4.74817
R18289 gnd.n2334 gnd.n2333 4.74817
R18290 gnd.n2422 gnd.n2373 4.74817
R18291 gnd.n2423 gnd.n2336 4.74817
R18292 gnd.n2425 gnd.n2335 4.74817
R18293 gnd.n2412 gnd.n2334 4.74817
R18294 gnd.n1182 gnd.n220 4.74817
R18295 gnd.n5635 gnd.n219 4.74817
R18296 gnd.n5633 gnd.n218 4.74817
R18297 gnd.n6785 gnd.n217 4.74817
R18298 gnd.n221 gnd.n216 4.74817
R18299 gnd.n5617 gnd.n220 4.74817
R18300 gnd.n1183 gnd.n219 4.74817
R18301 gnd.n5636 gnd.n218 4.74817
R18302 gnd.n5632 gnd.n217 4.74817
R18303 gnd.n6786 gnd.n216 4.74817
R18304 gnd.n3868 gnd.n2059 4.74817
R18305 gnd.n3907 gnd.n3898 4.74817
R18306 gnd.n3905 gnd.n3904 4.74817
R18307 gnd.n3900 gnd.n3899 4.74817
R18308 gnd.n3960 gnd.n2011 4.74817
R18309 gnd.n5605 gnd.n5603 4.74817
R18310 gnd.n5641 gnd.n1173 4.74817
R18311 gnd.n5663 gnd.n5643 4.74817
R18312 gnd.n5661 gnd.n5660 4.74817
R18313 gnd.n5656 gnd.n5646 4.74817
R18314 gnd.n5608 gnd.n5603 4.74817
R18315 gnd.n5604 gnd.n1173 4.74817
R18316 gnd.n5643 gnd.n5642 4.74817
R18317 gnd.n5662 gnd.n5661 4.74817
R18318 gnd.n5646 gnd.n5644 4.74817
R18319 gnd.n5908 gnd.n898 4.74817
R18320 gnd.n5906 gnd.n899 4.74817
R18321 gnd.n2026 gnd.n904 4.74817
R18322 gnd.n3946 gnd.n903 4.74817
R18323 gnd.n905 gnd.n902 4.74817
R18324 gnd.n898 gnd.n882 4.74817
R18325 gnd.n5907 gnd.n5906 4.74817
R18326 gnd.n3911 gnd.n904 4.74817
R18327 gnd.n2027 gnd.n903 4.74817
R18328 gnd.n3945 gnd.n902 4.74817
R18329 gnd.n3896 gnd.n2059 4.74817
R18330 gnd.n3898 gnd.n3897 4.74817
R18331 gnd.n3906 gnd.n3905 4.74817
R18332 gnd.n3901 gnd.n3900 4.74817
R18333 gnd.n2013 gnd.n2011 4.74817
R18334 gnd.n2359 gnd.n2358 4.7074
R18335 gnd.n38 gnd.n37 4.7074
R18336 gnd.n2371 gnd.n2359 4.65959
R18337 gnd.n50 gnd.n38 4.65959
R18338 gnd.n5411 gnd.n5410 4.6132
R18339 gnd.n4346 gnd.n4345 4.6132
R18340 gnd.n4420 gnd.n4419 4.46168
R18341 gnd.n4465 gnd.n1653 4.46168
R18342 gnd.n4459 gnd.t192 4.46168
R18343 gnd.n4593 gnd.n4591 4.46168
R18344 gnd.n4621 gnd.n1567 4.46168
R18345 gnd.n4767 gnd.n1486 4.46168
R18346 gnd.n4810 gnd.n1472 4.46168
R18347 gnd.n4948 gnd.n1343 4.46168
R18348 gnd.n5209 gnd.n5196 4.46111
R18349 gnd.n3410 gnd.n3406 4.38594
R18350 gnd.n3378 gnd.n3374 4.38594
R18351 gnd.n3346 gnd.n3342 4.38594
R18352 gnd.n3315 gnd.n3311 4.38594
R18353 gnd.n3283 gnd.n3279 4.38594
R18354 gnd.n3251 gnd.n3247 4.38594
R18355 gnd.n3219 gnd.n3215 4.38594
R18356 gnd.n3188 gnd.n3184 4.38594
R18357 gnd.n3421 gnd.n3399 4.26717
R18358 gnd.n3389 gnd.n3367 4.26717
R18359 gnd.n3357 gnd.n3335 4.26717
R18360 gnd.n3326 gnd.n3304 4.26717
R18361 gnd.n3294 gnd.n3272 4.26717
R18362 gnd.n3262 gnd.n3240 4.26717
R18363 gnd.n3230 gnd.n3208 4.26717
R18364 gnd.n3199 gnd.n3177 4.26717
R18365 gnd.n2878 gnd.t16 4.14303
R18366 gnd.n3109 gnd.t13 4.14303
R18367 gnd.t157 gnd.n986 4.14303
R18368 gnd.t150 gnd.n1138 4.14303
R18369 gnd.n3429 gnd.n3428 4.08274
R18370 gnd.n5342 gnd.n5341 4.05904
R18371 gnd.n1801 gnd.n1800 4.05904
R18372 gnd.n4358 gnd.n1737 4.05904
R18373 gnd.n5222 gnd.n5221 4.05904
R18374 gnd.n15 gnd.n7 3.99943
R18375 gnd.n4508 gnd.n4507 3.82437
R18376 gnd.t250 gnd.n1599 3.82437
R18377 gnd.n4641 gnd.n1556 3.82437
R18378 gnd.n4725 gnd.n4724 3.82437
R18379 gnd.n4839 gnd.t242 3.82437
R18380 gnd.n4893 gnd.n4892 3.82437
R18381 gnd.t147 gnd.n1334 3.82437
R18382 gnd.n3429 gnd.n3301 3.70378
R18383 gnd.n2951 gnd.n2372 3.65935
R18384 gnd.n15 gnd.n14 3.60163
R18385 gnd.t25 gnd.n3079 3.50571
R18386 gnd.n4410 gnd.n1700 3.50571
R18387 gnd.n5349 gnd.n1313 3.50571
R18388 gnd.n3420 gnd.n3401 3.49141
R18389 gnd.n3388 gnd.n3369 3.49141
R18390 gnd.n3356 gnd.n3337 3.49141
R18391 gnd.n3325 gnd.n3306 3.49141
R18392 gnd.n3293 gnd.n3274 3.49141
R18393 gnd.n3261 gnd.n3242 3.49141
R18394 gnd.n3229 gnd.n3210 3.49141
R18395 gnd.n3198 gnd.n3179 3.49141
R18396 gnd.n4245 gnd.t136 3.18706
R18397 gnd.n4487 gnd.n1645 3.18706
R18398 gnd.n4576 gnd.n4575 3.18706
R18399 gnd.t246 gnd.n4621 3.18706
R18400 gnd.n4632 gnd.n4631 3.18706
R18401 gnd.n4740 gnd.n4739 3.18706
R18402 gnd.n4767 gnd.t249 3.18706
R18403 gnd.n4820 gnd.n4819 3.18706
R18404 gnd.n4909 gnd.n4907 3.18706
R18405 gnd.t195 gnd.n1401 3.18706
R18406 gnd.n2457 gnd.t16 2.8684
R18407 gnd.n4429 gnd.t276 2.8684
R18408 gnd.t62 gnd.n4939 2.8684
R18409 gnd.n2360 gnd.t85 2.82907
R18410 gnd.n2360 gnd.t87 2.82907
R18411 gnd.n2362 gnd.t110 2.82907
R18412 gnd.n2362 gnd.t280 2.82907
R18413 gnd.n2364 gnd.t80 2.82907
R18414 gnd.n2364 gnd.t283 2.82907
R18415 gnd.n2366 gnd.t254 2.82907
R18416 gnd.n2366 gnd.t7 2.82907
R18417 gnd.n2368 gnd.t259 2.82907
R18418 gnd.n2368 gnd.t26 2.82907
R18419 gnd.n2337 gnd.t9 2.82907
R18420 gnd.n2337 gnd.t44 2.82907
R18421 gnd.n2339 gnd.t84 2.82907
R18422 gnd.n2339 gnd.t3 2.82907
R18423 gnd.n2341 gnd.t30 2.82907
R18424 gnd.n2341 gnd.t35 2.82907
R18425 gnd.n2343 gnd.t70 2.82907
R18426 gnd.n2343 gnd.t282 2.82907
R18427 gnd.n2345 gnd.t123 2.82907
R18428 gnd.n2345 gnd.t1 2.82907
R18429 gnd.n2348 gnd.t81 2.82907
R18430 gnd.n2348 gnd.t241 2.82907
R18431 gnd.n2350 gnd.t271 2.82907
R18432 gnd.n2350 gnd.t75 2.82907
R18433 gnd.n2352 gnd.t31 2.82907
R18434 gnd.n2352 gnd.t257 2.82907
R18435 gnd.n2354 gnd.t107 2.82907
R18436 gnd.n2354 gnd.t124 2.82907
R18437 gnd.n2356 gnd.t48 2.82907
R18438 gnd.n2356 gnd.t100 2.82907
R18439 gnd.n47 gnd.t28 2.82907
R18440 gnd.n47 gnd.t86 2.82907
R18441 gnd.n45 gnd.t40 2.82907
R18442 gnd.n45 gnd.t68 2.82907
R18443 gnd.n43 gnd.t111 2.82907
R18444 gnd.n43 gnd.t114 2.82907
R18445 gnd.n41 gnd.t127 2.82907
R18446 gnd.n41 gnd.t267 2.82907
R18447 gnd.n39 gnd.t59 2.82907
R18448 gnd.n39 gnd.t268 2.82907
R18449 gnd.n24 gnd.t266 2.82907
R18450 gnd.n24 gnd.t128 2.82907
R18451 gnd.n22 gnd.t33 2.82907
R18452 gnd.n22 gnd.t243 2.82907
R18453 gnd.n20 gnd.t273 2.82907
R18454 gnd.n20 gnd.t5 2.82907
R18455 gnd.n18 gnd.t37 2.82907
R18456 gnd.n18 gnd.t89 2.82907
R18457 gnd.n16 gnd.t39 2.82907
R18458 gnd.n16 gnd.t58 2.82907
R18459 gnd.n35 gnd.t272 2.82907
R18460 gnd.n35 gnd.t52 2.82907
R18461 gnd.n33 gnd.t244 2.82907
R18462 gnd.n33 gnd.t74 2.82907
R18463 gnd.n31 gnd.t73 2.82907
R18464 gnd.n31 gnd.t77 2.82907
R18465 gnd.n29 gnd.t130 2.82907
R18466 gnd.n29 gnd.t92 2.82907
R18467 gnd.n27 gnd.t126 2.82907
R18468 gnd.n27 gnd.t129 2.82907
R18469 gnd.n3417 gnd.n3416 2.71565
R18470 gnd.n3385 gnd.n3384 2.71565
R18471 gnd.n3353 gnd.n3352 2.71565
R18472 gnd.n3322 gnd.n3321 2.71565
R18473 gnd.n3290 gnd.n3289 2.71565
R18474 gnd.n3258 gnd.n3257 2.71565
R18475 gnd.n3226 gnd.n3225 2.71565
R18476 gnd.n3195 gnd.n3194 2.71565
R18477 gnd.t154 gnd.n4466 2.54975
R18478 gnd.t192 gnd.n1655 2.54975
R18479 gnd.n4485 gnd.n1647 2.54975
R18480 gnd.t125 gnd.n1618 2.54975
R18481 gnd.n4557 gnd.n4556 2.54975
R18482 gnd.n4652 gnd.n1549 2.54975
R18483 gnd.n4741 gnd.n1501 2.54975
R18484 gnd.n4829 gnd.n4828 2.54975
R18485 gnd.n4874 gnd.t108 2.54975
R18486 gnd.n4910 gnd.n1412 2.54975
R18487 gnd.n4931 gnd.t230 2.54975
R18488 gnd.n2951 gnd.n2373 2.27742
R18489 gnd.n2951 gnd.n2336 2.27742
R18490 gnd.n2951 gnd.n2335 2.27742
R18491 gnd.n2951 gnd.n2334 2.27742
R18492 gnd.n6799 gnd.n220 2.27742
R18493 gnd.n6799 gnd.n219 2.27742
R18494 gnd.n6799 gnd.n218 2.27742
R18495 gnd.n6799 gnd.n217 2.27742
R18496 gnd.n6799 gnd.n216 2.27742
R18497 gnd.n5603 gnd.n215 2.27742
R18498 gnd.n1173 gnd.n215 2.27742
R18499 gnd.n5643 gnd.n215 2.27742
R18500 gnd.n5661 gnd.n215 2.27742
R18501 gnd.n5646 gnd.n215 2.27742
R18502 gnd.n5905 gnd.n898 2.27742
R18503 gnd.n5906 gnd.n5905 2.27742
R18504 gnd.n5905 gnd.n904 2.27742
R18505 gnd.n5905 gnd.n903 2.27742
R18506 gnd.n5905 gnd.n902 2.27742
R18507 gnd.n2059 gnd.n901 2.27742
R18508 gnd.n3898 gnd.n901 2.27742
R18509 gnd.n3905 gnd.n901 2.27742
R18510 gnd.n3900 gnd.n901 2.27742
R18511 gnd.n2011 gnd.n901 2.27742
R18512 gnd.n2805 gnd.t132 2.23109
R18513 gnd.n2428 gnd.t14 2.23109
R18514 gnd.t90 gnd.n1567 2.23109
R18515 gnd.t278 gnd.n1486 2.23109
R18516 gnd.n3413 gnd.n3403 1.93989
R18517 gnd.n3381 gnd.n3371 1.93989
R18518 gnd.n3349 gnd.n3339 1.93989
R18519 gnd.n3318 gnd.n3308 1.93989
R18520 gnd.n3286 gnd.n3276 1.93989
R18521 gnd.n3254 gnd.n3244 1.93989
R18522 gnd.n3222 gnd.n3212 1.93989
R18523 gnd.n3191 gnd.n3181 1.93989
R18524 gnd.n1676 gnd.t208 1.91244
R18525 gnd.n4496 gnd.n4495 1.91244
R18526 gnd.n4565 gnd.n4563 1.91244
R18527 gnd.n4661 gnd.n1544 1.91244
R18528 gnd.t245 gnd.n4641 1.91244
R18529 gnd.n4725 gnd.t239 1.91244
R18530 gnd.n1514 gnd.n1513 1.91244
R18531 gnd.n4842 gnd.n4841 1.91244
R18532 gnd.n4857 gnd.n4856 1.91244
R18533 gnd.n1404 gnd.t230 1.91244
R18534 gnd.t255 gnd.n2816 1.59378
R18535 gnd.n2995 gnd.t11 1.59378
R18536 gnd.n2269 gnd.t260 1.59378
R18537 gnd.n4498 gnd.t121 1.59378
R18538 gnd.t98 gnd.n1589 1.59378
R18539 gnd.n4821 gnd.t264 1.59378
R18540 gnd.n4900 gnd.t274 1.59378
R18541 gnd.n4421 gnd.n1671 1.27512
R18542 gnd.t139 gnd.n4465 1.27512
R18543 gnd.n4477 gnd.n4476 1.27512
R18544 gnd.n4508 gnd.t105 1.27512
R18545 gnd.n4583 gnd.n1584 1.27512
R18546 gnd.n4605 gnd.n1577 1.27512
R18547 gnd.n4750 gnd.n4749 1.27512
R18548 gnd.n4808 gnd.n1473 1.27512
R18549 gnd.n4892 gnd.t247 1.27512
R18550 gnd.n4922 gnd.n4921 1.27512
R18551 gnd.n4931 gnd.t161 1.27512
R18552 gnd.n5282 gnd.n1334 1.27512
R18553 gnd.t217 gnd.n1313 1.27512
R18554 gnd.n2658 gnd.n2650 1.16414
R18555 gnd.n3475 gnd.n2172 1.16414
R18556 gnd.n3412 gnd.n3405 1.16414
R18557 gnd.n3380 gnd.n3373 1.16414
R18558 gnd.n3348 gnd.n3341 1.16414
R18559 gnd.n3317 gnd.n3310 1.16414
R18560 gnd.n3285 gnd.n3278 1.16414
R18561 gnd.n3253 gnd.n3246 1.16414
R18562 gnd.n3221 gnd.n3214 1.16414
R18563 gnd.n3190 gnd.n3183 1.16414
R18564 gnd.n5410 gnd.n1289 0.970197
R18565 gnd.n4346 gnd.n1807 0.970197
R18566 gnd.n3396 gnd.n3364 0.962709
R18567 gnd.n3428 gnd.n3396 0.962709
R18568 gnd.n3269 gnd.n3237 0.962709
R18569 gnd.n3301 gnd.n3269 0.962709
R18570 gnd.n2904 gnd.t53 0.956468
R18571 gnd.n3069 gnd.t20 0.956468
R18572 gnd.t60 gnd.n840 0.956468
R18573 gnd.n5934 gnd.t47 0.956468
R18574 gnd.n4023 gnd.t8 0.956468
R18575 gnd.n3985 gnd.t43 0.956468
R18576 gnd.n4242 gnd.t64 0.956468
R18577 gnd.n5183 gnd.t101 0.956468
R18578 gnd.n5575 gnd.t38 0.956468
R18579 gnd.n1222 gnd.t57 0.956468
R18580 gnd.n266 gnd.t51 0.956468
R18581 gnd.t78 gnd.n177 0.956468
R18582 gnd.n2367 gnd.n2365 0.773756
R18583 gnd.n46 gnd.n44 0.773756
R18584 gnd.n2370 gnd.n2369 0.773756
R18585 gnd.n2369 gnd.n2367 0.773756
R18586 gnd.n2365 gnd.n2363 0.773756
R18587 gnd.n2363 gnd.n2361 0.773756
R18588 gnd.n42 gnd.n40 0.773756
R18589 gnd.n44 gnd.n42 0.773756
R18590 gnd.n48 gnd.n46 0.773756
R18591 gnd.n49 gnd.n48 0.773756
R18592 gnd.n2 gnd.n1 0.672012
R18593 gnd.n3 gnd.n2 0.672012
R18594 gnd.n4 gnd.n3 0.672012
R18595 gnd.n5 gnd.n4 0.672012
R18596 gnd.n6 gnd.n5 0.672012
R18597 gnd.n7 gnd.n6 0.672012
R18598 gnd.n9 gnd.n8 0.672012
R18599 gnd.n10 gnd.n9 0.672012
R18600 gnd.n11 gnd.n10 0.672012
R18601 gnd.n12 gnd.n11 0.672012
R18602 gnd.n13 gnd.n12 0.672012
R18603 gnd.n14 gnd.n13 0.672012
R18604 gnd.n4520 gnd.n1625 0.637812
R18605 gnd.n4528 gnd.n1612 0.637812
R18606 gnd.n4672 gnd.n4671 0.637812
R18607 gnd.n4715 gnd.n4714 0.637812
R18608 gnd.n4780 gnd.n4779 0.637812
R18609 gnd.n4883 gnd.n4881 0.637812
R18610 gnd.n2347 gnd.n2346 0.573776
R18611 gnd.n2346 gnd.n2344 0.573776
R18612 gnd.n2344 gnd.n2342 0.573776
R18613 gnd.n2342 gnd.n2340 0.573776
R18614 gnd.n2340 gnd.n2338 0.573776
R18615 gnd.n2358 gnd.n2357 0.573776
R18616 gnd.n2357 gnd.n2355 0.573776
R18617 gnd.n2355 gnd.n2353 0.573776
R18618 gnd.n2353 gnd.n2351 0.573776
R18619 gnd.n2351 gnd.n2349 0.573776
R18620 gnd.n19 gnd.n17 0.573776
R18621 gnd.n21 gnd.n19 0.573776
R18622 gnd.n23 gnd.n21 0.573776
R18623 gnd.n25 gnd.n23 0.573776
R18624 gnd.n26 gnd.n25 0.573776
R18625 gnd.n30 gnd.n28 0.573776
R18626 gnd.n32 gnd.n30 0.573776
R18627 gnd.n34 gnd.n32 0.573776
R18628 gnd.n36 gnd.n34 0.573776
R18629 gnd.n37 gnd.n36 0.573776
R18630 gnd gnd.n0 0.551497
R18631 gnd.n6799 gnd.n215 0.548625
R18632 gnd.n5905 gnd.n901 0.548625
R18633 gnd.n3640 gnd.n3639 0.532512
R18634 gnd.n3790 gnd.n3789 0.532512
R18635 gnd.n6909 gnd.n6908 0.532512
R18636 gnd.n7009 gnd.n78 0.532512
R18637 gnd.n5849 gnd.n5848 0.523366
R18638 gnd.n5025 gnd.n1104 0.523366
R18639 gnd.n7003 gnd.n7002 0.520317
R18640 gnd.n6932 gnd.n6931 0.520317
R18641 gnd.n5464 gnd.n5463 0.520317
R18642 gnd.n5368 gnd.n1133 0.520317
R18643 gnd.n1828 gnd.n991 0.520317
R18644 gnd.n4306 gnd.n4305 0.520317
R18645 gnd.n3709 gnd.n3688 0.520317
R18646 gnd.n3645 gnd.n2092 0.520317
R18647 gnd.n5147 gnd.n5146 0.489829
R18648 gnd.n4279 gnd.n4278 0.489829
R18649 gnd.n3132 gnd.n2176 0.486781
R18650 gnd.n2707 gnd.n2706 0.48678
R18651 gnd.n3449 gnd.n2130 0.480683
R18652 gnd.n2791 gnd.n2790 0.480683
R18653 gnd.n6119 gnd.n6118 0.480683
R18654 gnd.n6539 gnd.n6538 0.480683
R18655 gnd.n6752 gnd.n6751 0.480683
R18656 gnd.n3850 gnd.n825 0.480683
R18657 gnd.n7042 gnd.n7041 0.470187
R18658 gnd.n5851 gnd.n5850 0.432431
R18659 gnd.n5028 gnd.n5027 0.432431
R18660 gnd.n4286 gnd.n1921 0.388379
R18661 gnd.n3409 gnd.n3408 0.388379
R18662 gnd.n3377 gnd.n3376 0.388379
R18663 gnd.n3345 gnd.n3344 0.388379
R18664 gnd.n3314 gnd.n3313 0.388379
R18665 gnd.n3282 gnd.n3281 0.388379
R18666 gnd.n3250 gnd.n3249 0.388379
R18667 gnd.n3218 gnd.n3217 0.388379
R18668 gnd.n3187 gnd.n3186 0.388379
R18669 gnd.n6972 gnd.n6971 0.388379
R18670 gnd.n3750 gnd.n3749 0.388379
R18671 gnd.n5136 gnd.n5135 0.388379
R18672 gnd.n7042 gnd.n15 0.374463
R18673 gnd.n2231 gnd.t17 0.319156
R18674 gnd.n3872 gnd.t69 0.319156
R18675 gnd.n5910 gnd.t6 0.319156
R18676 gnd.t34 gnd.n2021 0.319156
R18677 gnd.t83 gnd.n3956 0.319156
R18678 gnd.n4204 gnd.t201 0.319156
R18679 gnd.t112 gnd.t245 0.319156
R18680 gnd.t96 gnd.t239 0.319156
R18681 gnd.t182 gnd.n5157 0.319156
R18682 gnd.n5506 gnd.t88 0.319156
R18683 gnd.n5639 gnd.t72 0.319156
R18684 gnd.n6777 gnd.t32 0.319156
R18685 gnd.t67 gnd.n209 0.319156
R18686 gnd.n2625 gnd.n2603 0.311721
R18687 gnd.n4297 gnd.n4296 0.302329
R18688 gnd.n5115 gnd.n1264 0.302329
R18689 gnd gnd.n7042 0.295112
R18690 gnd.n3520 gnd.n3519 0.268793
R18691 gnd.n3519 gnd.n3518 0.241354
R18692 gnd.n5411 gnd.n1290 0.229039
R18693 gnd.n5412 gnd.n5411 0.229039
R18694 gnd.n4345 gnd.n1812 0.229039
R18695 gnd.n4345 gnd.n4344 0.229039
R18696 gnd.n2779 gnd.n2578 0.206293
R18697 gnd.n3426 gnd.n3398 0.155672
R18698 gnd.n3419 gnd.n3398 0.155672
R18699 gnd.n3419 gnd.n3418 0.155672
R18700 gnd.n3418 gnd.n3402 0.155672
R18701 gnd.n3411 gnd.n3402 0.155672
R18702 gnd.n3411 gnd.n3410 0.155672
R18703 gnd.n3394 gnd.n3366 0.155672
R18704 gnd.n3387 gnd.n3366 0.155672
R18705 gnd.n3387 gnd.n3386 0.155672
R18706 gnd.n3386 gnd.n3370 0.155672
R18707 gnd.n3379 gnd.n3370 0.155672
R18708 gnd.n3379 gnd.n3378 0.155672
R18709 gnd.n3362 gnd.n3334 0.155672
R18710 gnd.n3355 gnd.n3334 0.155672
R18711 gnd.n3355 gnd.n3354 0.155672
R18712 gnd.n3354 gnd.n3338 0.155672
R18713 gnd.n3347 gnd.n3338 0.155672
R18714 gnd.n3347 gnd.n3346 0.155672
R18715 gnd.n3331 gnd.n3303 0.155672
R18716 gnd.n3324 gnd.n3303 0.155672
R18717 gnd.n3324 gnd.n3323 0.155672
R18718 gnd.n3323 gnd.n3307 0.155672
R18719 gnd.n3316 gnd.n3307 0.155672
R18720 gnd.n3316 gnd.n3315 0.155672
R18721 gnd.n3299 gnd.n3271 0.155672
R18722 gnd.n3292 gnd.n3271 0.155672
R18723 gnd.n3292 gnd.n3291 0.155672
R18724 gnd.n3291 gnd.n3275 0.155672
R18725 gnd.n3284 gnd.n3275 0.155672
R18726 gnd.n3284 gnd.n3283 0.155672
R18727 gnd.n3267 gnd.n3239 0.155672
R18728 gnd.n3260 gnd.n3239 0.155672
R18729 gnd.n3260 gnd.n3259 0.155672
R18730 gnd.n3259 gnd.n3243 0.155672
R18731 gnd.n3252 gnd.n3243 0.155672
R18732 gnd.n3252 gnd.n3251 0.155672
R18733 gnd.n3235 gnd.n3207 0.155672
R18734 gnd.n3228 gnd.n3207 0.155672
R18735 gnd.n3228 gnd.n3227 0.155672
R18736 gnd.n3227 gnd.n3211 0.155672
R18737 gnd.n3220 gnd.n3211 0.155672
R18738 gnd.n3220 gnd.n3219 0.155672
R18739 gnd.n3204 gnd.n3176 0.155672
R18740 gnd.n3197 gnd.n3176 0.155672
R18741 gnd.n3197 gnd.n3196 0.155672
R18742 gnd.n3196 gnd.n3180 0.155672
R18743 gnd.n3189 gnd.n3180 0.155672
R18744 gnd.n3189 gnd.n3188 0.155672
R18745 gnd.n3551 gnd.n2130 0.152939
R18746 gnd.n3551 gnd.n3550 0.152939
R18747 gnd.n3550 gnd.n3549 0.152939
R18748 gnd.n3549 gnd.n2132 0.152939
R18749 gnd.n2133 gnd.n2132 0.152939
R18750 gnd.n2134 gnd.n2133 0.152939
R18751 gnd.n2135 gnd.n2134 0.152939
R18752 gnd.n2136 gnd.n2135 0.152939
R18753 gnd.n2137 gnd.n2136 0.152939
R18754 gnd.n2138 gnd.n2137 0.152939
R18755 gnd.n2139 gnd.n2138 0.152939
R18756 gnd.n2140 gnd.n2139 0.152939
R18757 gnd.n2141 gnd.n2140 0.152939
R18758 gnd.n2142 gnd.n2141 0.152939
R18759 gnd.n3521 gnd.n2142 0.152939
R18760 gnd.n3521 gnd.n3520 0.152939
R18761 gnd.n2792 gnd.n2791 0.152939
R18762 gnd.n2792 gnd.n2496 0.152939
R18763 gnd.n2820 gnd.n2496 0.152939
R18764 gnd.n2821 gnd.n2820 0.152939
R18765 gnd.n2822 gnd.n2821 0.152939
R18766 gnd.n2823 gnd.n2822 0.152939
R18767 gnd.n2823 gnd.n2468 0.152939
R18768 gnd.n2850 gnd.n2468 0.152939
R18769 gnd.n2851 gnd.n2850 0.152939
R18770 gnd.n2852 gnd.n2851 0.152939
R18771 gnd.n2852 gnd.n2446 0.152939
R18772 gnd.n2881 gnd.n2446 0.152939
R18773 gnd.n2882 gnd.n2881 0.152939
R18774 gnd.n2883 gnd.n2882 0.152939
R18775 gnd.n2884 gnd.n2883 0.152939
R18776 gnd.n2886 gnd.n2884 0.152939
R18777 gnd.n2886 gnd.n2885 0.152939
R18778 gnd.n2885 gnd.n2395 0.152939
R18779 gnd.n2396 gnd.n2395 0.152939
R18780 gnd.n2397 gnd.n2396 0.152939
R18781 gnd.n2416 gnd.n2397 0.152939
R18782 gnd.n2417 gnd.n2416 0.152939
R18783 gnd.n2417 gnd.n2327 0.152939
R18784 gnd.n2976 gnd.n2327 0.152939
R18785 gnd.n2977 gnd.n2976 0.152939
R18786 gnd.n2978 gnd.n2977 0.152939
R18787 gnd.n2979 gnd.n2978 0.152939
R18788 gnd.n2979 gnd.n2300 0.152939
R18789 gnd.n3016 gnd.n2300 0.152939
R18790 gnd.n3017 gnd.n3016 0.152939
R18791 gnd.n3018 gnd.n3017 0.152939
R18792 gnd.n3019 gnd.n3018 0.152939
R18793 gnd.n3019 gnd.n2273 0.152939
R18794 gnd.n3061 gnd.n2273 0.152939
R18795 gnd.n3062 gnd.n3061 0.152939
R18796 gnd.n3063 gnd.n3062 0.152939
R18797 gnd.n3064 gnd.n3063 0.152939
R18798 gnd.n3064 gnd.n2245 0.152939
R18799 gnd.n3102 gnd.n2245 0.152939
R18800 gnd.n3103 gnd.n3102 0.152939
R18801 gnd.n3104 gnd.n3103 0.152939
R18802 gnd.n3105 gnd.n3104 0.152939
R18803 gnd.n3105 gnd.n2218 0.152939
R18804 gnd.n3151 gnd.n2218 0.152939
R18805 gnd.n3152 gnd.n3151 0.152939
R18806 gnd.n3153 gnd.n3152 0.152939
R18807 gnd.n3154 gnd.n3153 0.152939
R18808 gnd.n3154 gnd.n2191 0.152939
R18809 gnd.n3445 gnd.n2191 0.152939
R18810 gnd.n3446 gnd.n3445 0.152939
R18811 gnd.n3447 gnd.n3446 0.152939
R18812 gnd.n3448 gnd.n3447 0.152939
R18813 gnd.n3449 gnd.n3448 0.152939
R18814 gnd.n2790 gnd.n2520 0.152939
R18815 gnd.n2541 gnd.n2520 0.152939
R18816 gnd.n2542 gnd.n2541 0.152939
R18817 gnd.n2548 gnd.n2542 0.152939
R18818 gnd.n2549 gnd.n2548 0.152939
R18819 gnd.n2550 gnd.n2549 0.152939
R18820 gnd.n2550 gnd.n2539 0.152939
R18821 gnd.n2558 gnd.n2539 0.152939
R18822 gnd.n2559 gnd.n2558 0.152939
R18823 gnd.n2560 gnd.n2559 0.152939
R18824 gnd.n2560 gnd.n2537 0.152939
R18825 gnd.n2568 gnd.n2537 0.152939
R18826 gnd.n2569 gnd.n2568 0.152939
R18827 gnd.n2570 gnd.n2569 0.152939
R18828 gnd.n2570 gnd.n2535 0.152939
R18829 gnd.n2578 gnd.n2535 0.152939
R18830 gnd.n3518 gnd.n2147 0.152939
R18831 gnd.n2149 gnd.n2147 0.152939
R18832 gnd.n2150 gnd.n2149 0.152939
R18833 gnd.n2151 gnd.n2150 0.152939
R18834 gnd.n2152 gnd.n2151 0.152939
R18835 gnd.n2153 gnd.n2152 0.152939
R18836 gnd.n2154 gnd.n2153 0.152939
R18837 gnd.n2155 gnd.n2154 0.152939
R18838 gnd.n2156 gnd.n2155 0.152939
R18839 gnd.n2157 gnd.n2156 0.152939
R18840 gnd.n2158 gnd.n2157 0.152939
R18841 gnd.n2159 gnd.n2158 0.152939
R18842 gnd.n2160 gnd.n2159 0.152939
R18843 gnd.n2161 gnd.n2160 0.152939
R18844 gnd.n2162 gnd.n2161 0.152939
R18845 gnd.n2163 gnd.n2162 0.152939
R18846 gnd.n2164 gnd.n2163 0.152939
R18847 gnd.n2165 gnd.n2164 0.152939
R18848 gnd.n2166 gnd.n2165 0.152939
R18849 gnd.n2167 gnd.n2166 0.152939
R18850 gnd.n2168 gnd.n2167 0.152939
R18851 gnd.n2169 gnd.n2168 0.152939
R18852 gnd.n2173 gnd.n2169 0.152939
R18853 gnd.n2174 gnd.n2173 0.152939
R18854 gnd.n2175 gnd.n2174 0.152939
R18855 gnd.n2176 gnd.n2175 0.152939
R18856 gnd.n2953 gnd.n2952 0.152939
R18857 gnd.n2954 gnd.n2953 0.152939
R18858 gnd.n2955 gnd.n2954 0.152939
R18859 gnd.n2956 gnd.n2955 0.152939
R18860 gnd.n2957 gnd.n2956 0.152939
R18861 gnd.n2958 gnd.n2957 0.152939
R18862 gnd.n2958 gnd.n2281 0.152939
R18863 gnd.n3037 gnd.n2281 0.152939
R18864 gnd.n3038 gnd.n3037 0.152939
R18865 gnd.n3039 gnd.n3038 0.152939
R18866 gnd.n3040 gnd.n3039 0.152939
R18867 gnd.n3041 gnd.n3040 0.152939
R18868 gnd.n3042 gnd.n3041 0.152939
R18869 gnd.n3043 gnd.n3042 0.152939
R18870 gnd.n3044 gnd.n3043 0.152939
R18871 gnd.n3045 gnd.n3044 0.152939
R18872 gnd.n3045 gnd.n2225 0.152939
R18873 gnd.n3123 gnd.n2225 0.152939
R18874 gnd.n3124 gnd.n3123 0.152939
R18875 gnd.n3125 gnd.n3124 0.152939
R18876 gnd.n3126 gnd.n3125 0.152939
R18877 gnd.n3127 gnd.n3126 0.152939
R18878 gnd.n3128 gnd.n3127 0.152939
R18879 gnd.n3129 gnd.n3128 0.152939
R18880 gnd.n3130 gnd.n3129 0.152939
R18881 gnd.n3131 gnd.n3130 0.152939
R18882 gnd.n3133 gnd.n3131 0.152939
R18883 gnd.n3133 gnd.n3132 0.152939
R18884 gnd.n2708 gnd.n2707 0.152939
R18885 gnd.n2708 gnd.n2598 0.152939
R18886 gnd.n2723 gnd.n2598 0.152939
R18887 gnd.n2724 gnd.n2723 0.152939
R18888 gnd.n2725 gnd.n2724 0.152939
R18889 gnd.n2725 gnd.n2586 0.152939
R18890 gnd.n2739 gnd.n2586 0.152939
R18891 gnd.n2740 gnd.n2739 0.152939
R18892 gnd.n2741 gnd.n2740 0.152939
R18893 gnd.n2742 gnd.n2741 0.152939
R18894 gnd.n2743 gnd.n2742 0.152939
R18895 gnd.n2744 gnd.n2743 0.152939
R18896 gnd.n2745 gnd.n2744 0.152939
R18897 gnd.n2746 gnd.n2745 0.152939
R18898 gnd.n2747 gnd.n2746 0.152939
R18899 gnd.n2748 gnd.n2747 0.152939
R18900 gnd.n2749 gnd.n2748 0.152939
R18901 gnd.n2750 gnd.n2749 0.152939
R18902 gnd.n2751 gnd.n2750 0.152939
R18903 gnd.n2752 gnd.n2751 0.152939
R18904 gnd.n2753 gnd.n2752 0.152939
R18905 gnd.n2753 gnd.n2452 0.152939
R18906 gnd.n2870 gnd.n2452 0.152939
R18907 gnd.n2871 gnd.n2870 0.152939
R18908 gnd.n2872 gnd.n2871 0.152939
R18909 gnd.n2873 gnd.n2872 0.152939
R18910 gnd.n2873 gnd.n2374 0.152939
R18911 gnd.n2950 gnd.n2374 0.152939
R18912 gnd.n2626 gnd.n2625 0.152939
R18913 gnd.n2627 gnd.n2626 0.152939
R18914 gnd.n2628 gnd.n2627 0.152939
R18915 gnd.n2629 gnd.n2628 0.152939
R18916 gnd.n2630 gnd.n2629 0.152939
R18917 gnd.n2631 gnd.n2630 0.152939
R18918 gnd.n2632 gnd.n2631 0.152939
R18919 gnd.n2633 gnd.n2632 0.152939
R18920 gnd.n2634 gnd.n2633 0.152939
R18921 gnd.n2635 gnd.n2634 0.152939
R18922 gnd.n2636 gnd.n2635 0.152939
R18923 gnd.n2637 gnd.n2636 0.152939
R18924 gnd.n2638 gnd.n2637 0.152939
R18925 gnd.n2639 gnd.n2638 0.152939
R18926 gnd.n2640 gnd.n2639 0.152939
R18927 gnd.n2641 gnd.n2640 0.152939
R18928 gnd.n2642 gnd.n2641 0.152939
R18929 gnd.n2643 gnd.n2642 0.152939
R18930 gnd.n2644 gnd.n2643 0.152939
R18931 gnd.n2645 gnd.n2644 0.152939
R18932 gnd.n2646 gnd.n2645 0.152939
R18933 gnd.n2647 gnd.n2646 0.152939
R18934 gnd.n2651 gnd.n2647 0.152939
R18935 gnd.n2652 gnd.n2651 0.152939
R18936 gnd.n2652 gnd.n2609 0.152939
R18937 gnd.n2706 gnd.n2609 0.152939
R18938 gnd.n6120 gnd.n6119 0.152939
R18939 gnd.n6120 gnd.n652 0.152939
R18940 gnd.n6128 gnd.n652 0.152939
R18941 gnd.n6129 gnd.n6128 0.152939
R18942 gnd.n6130 gnd.n6129 0.152939
R18943 gnd.n6130 gnd.n646 0.152939
R18944 gnd.n6138 gnd.n646 0.152939
R18945 gnd.n6139 gnd.n6138 0.152939
R18946 gnd.n6140 gnd.n6139 0.152939
R18947 gnd.n6140 gnd.n640 0.152939
R18948 gnd.n6148 gnd.n640 0.152939
R18949 gnd.n6149 gnd.n6148 0.152939
R18950 gnd.n6150 gnd.n6149 0.152939
R18951 gnd.n6150 gnd.n634 0.152939
R18952 gnd.n6158 gnd.n634 0.152939
R18953 gnd.n6159 gnd.n6158 0.152939
R18954 gnd.n6160 gnd.n6159 0.152939
R18955 gnd.n6160 gnd.n628 0.152939
R18956 gnd.n6168 gnd.n628 0.152939
R18957 gnd.n6169 gnd.n6168 0.152939
R18958 gnd.n6170 gnd.n6169 0.152939
R18959 gnd.n6170 gnd.n622 0.152939
R18960 gnd.n6178 gnd.n622 0.152939
R18961 gnd.n6179 gnd.n6178 0.152939
R18962 gnd.n6180 gnd.n6179 0.152939
R18963 gnd.n6180 gnd.n616 0.152939
R18964 gnd.n6188 gnd.n616 0.152939
R18965 gnd.n6189 gnd.n6188 0.152939
R18966 gnd.n6190 gnd.n6189 0.152939
R18967 gnd.n6190 gnd.n610 0.152939
R18968 gnd.n6198 gnd.n610 0.152939
R18969 gnd.n6199 gnd.n6198 0.152939
R18970 gnd.n6200 gnd.n6199 0.152939
R18971 gnd.n6200 gnd.n604 0.152939
R18972 gnd.n6208 gnd.n604 0.152939
R18973 gnd.n6209 gnd.n6208 0.152939
R18974 gnd.n6210 gnd.n6209 0.152939
R18975 gnd.n6210 gnd.n598 0.152939
R18976 gnd.n6218 gnd.n598 0.152939
R18977 gnd.n6219 gnd.n6218 0.152939
R18978 gnd.n6220 gnd.n6219 0.152939
R18979 gnd.n6220 gnd.n592 0.152939
R18980 gnd.n6228 gnd.n592 0.152939
R18981 gnd.n6229 gnd.n6228 0.152939
R18982 gnd.n6230 gnd.n6229 0.152939
R18983 gnd.n6230 gnd.n586 0.152939
R18984 gnd.n6238 gnd.n586 0.152939
R18985 gnd.n6239 gnd.n6238 0.152939
R18986 gnd.n6240 gnd.n6239 0.152939
R18987 gnd.n6240 gnd.n580 0.152939
R18988 gnd.n6248 gnd.n580 0.152939
R18989 gnd.n6249 gnd.n6248 0.152939
R18990 gnd.n6250 gnd.n6249 0.152939
R18991 gnd.n6250 gnd.n574 0.152939
R18992 gnd.n6258 gnd.n574 0.152939
R18993 gnd.n6259 gnd.n6258 0.152939
R18994 gnd.n6260 gnd.n6259 0.152939
R18995 gnd.n6260 gnd.n568 0.152939
R18996 gnd.n6268 gnd.n568 0.152939
R18997 gnd.n6269 gnd.n6268 0.152939
R18998 gnd.n6270 gnd.n6269 0.152939
R18999 gnd.n6270 gnd.n562 0.152939
R19000 gnd.n6278 gnd.n562 0.152939
R19001 gnd.n6279 gnd.n6278 0.152939
R19002 gnd.n6280 gnd.n6279 0.152939
R19003 gnd.n6280 gnd.n556 0.152939
R19004 gnd.n6288 gnd.n556 0.152939
R19005 gnd.n6289 gnd.n6288 0.152939
R19006 gnd.n6290 gnd.n6289 0.152939
R19007 gnd.n6290 gnd.n550 0.152939
R19008 gnd.n6298 gnd.n550 0.152939
R19009 gnd.n6299 gnd.n6298 0.152939
R19010 gnd.n6300 gnd.n6299 0.152939
R19011 gnd.n6300 gnd.n544 0.152939
R19012 gnd.n6308 gnd.n544 0.152939
R19013 gnd.n6309 gnd.n6308 0.152939
R19014 gnd.n6310 gnd.n6309 0.152939
R19015 gnd.n6310 gnd.n538 0.152939
R19016 gnd.n6318 gnd.n538 0.152939
R19017 gnd.n6319 gnd.n6318 0.152939
R19018 gnd.n6320 gnd.n6319 0.152939
R19019 gnd.n6320 gnd.n532 0.152939
R19020 gnd.n6328 gnd.n532 0.152939
R19021 gnd.n6329 gnd.n6328 0.152939
R19022 gnd.n6330 gnd.n6329 0.152939
R19023 gnd.n6330 gnd.n526 0.152939
R19024 gnd.n6338 gnd.n526 0.152939
R19025 gnd.n6339 gnd.n6338 0.152939
R19026 gnd.n6340 gnd.n6339 0.152939
R19027 gnd.n6340 gnd.n520 0.152939
R19028 gnd.n6348 gnd.n520 0.152939
R19029 gnd.n6349 gnd.n6348 0.152939
R19030 gnd.n6350 gnd.n6349 0.152939
R19031 gnd.n6350 gnd.n514 0.152939
R19032 gnd.n6358 gnd.n514 0.152939
R19033 gnd.n6359 gnd.n6358 0.152939
R19034 gnd.n6360 gnd.n6359 0.152939
R19035 gnd.n6360 gnd.n508 0.152939
R19036 gnd.n6368 gnd.n508 0.152939
R19037 gnd.n6369 gnd.n6368 0.152939
R19038 gnd.n6370 gnd.n6369 0.152939
R19039 gnd.n6370 gnd.n502 0.152939
R19040 gnd.n6378 gnd.n502 0.152939
R19041 gnd.n6379 gnd.n6378 0.152939
R19042 gnd.n6380 gnd.n6379 0.152939
R19043 gnd.n6380 gnd.n496 0.152939
R19044 gnd.n6388 gnd.n496 0.152939
R19045 gnd.n6389 gnd.n6388 0.152939
R19046 gnd.n6390 gnd.n6389 0.152939
R19047 gnd.n6390 gnd.n490 0.152939
R19048 gnd.n6398 gnd.n490 0.152939
R19049 gnd.n6399 gnd.n6398 0.152939
R19050 gnd.n6400 gnd.n6399 0.152939
R19051 gnd.n6400 gnd.n484 0.152939
R19052 gnd.n6408 gnd.n484 0.152939
R19053 gnd.n6409 gnd.n6408 0.152939
R19054 gnd.n6410 gnd.n6409 0.152939
R19055 gnd.n6410 gnd.n478 0.152939
R19056 gnd.n6418 gnd.n478 0.152939
R19057 gnd.n6419 gnd.n6418 0.152939
R19058 gnd.n6420 gnd.n6419 0.152939
R19059 gnd.n6420 gnd.n472 0.152939
R19060 gnd.n6428 gnd.n472 0.152939
R19061 gnd.n6429 gnd.n6428 0.152939
R19062 gnd.n6430 gnd.n6429 0.152939
R19063 gnd.n6430 gnd.n466 0.152939
R19064 gnd.n6438 gnd.n466 0.152939
R19065 gnd.n6439 gnd.n6438 0.152939
R19066 gnd.n6440 gnd.n6439 0.152939
R19067 gnd.n6440 gnd.n460 0.152939
R19068 gnd.n6448 gnd.n460 0.152939
R19069 gnd.n6449 gnd.n6448 0.152939
R19070 gnd.n6450 gnd.n6449 0.152939
R19071 gnd.n6450 gnd.n454 0.152939
R19072 gnd.n6458 gnd.n454 0.152939
R19073 gnd.n6459 gnd.n6458 0.152939
R19074 gnd.n6460 gnd.n6459 0.152939
R19075 gnd.n6460 gnd.n448 0.152939
R19076 gnd.n6468 gnd.n448 0.152939
R19077 gnd.n6469 gnd.n6468 0.152939
R19078 gnd.n6470 gnd.n6469 0.152939
R19079 gnd.n6470 gnd.n442 0.152939
R19080 gnd.n6478 gnd.n442 0.152939
R19081 gnd.n6479 gnd.n6478 0.152939
R19082 gnd.n6480 gnd.n6479 0.152939
R19083 gnd.n6480 gnd.n436 0.152939
R19084 gnd.n6488 gnd.n436 0.152939
R19085 gnd.n6489 gnd.n6488 0.152939
R19086 gnd.n6490 gnd.n6489 0.152939
R19087 gnd.n6490 gnd.n430 0.152939
R19088 gnd.n6498 gnd.n430 0.152939
R19089 gnd.n6499 gnd.n6498 0.152939
R19090 gnd.n6500 gnd.n6499 0.152939
R19091 gnd.n6500 gnd.n424 0.152939
R19092 gnd.n6508 gnd.n424 0.152939
R19093 gnd.n6509 gnd.n6508 0.152939
R19094 gnd.n6510 gnd.n6509 0.152939
R19095 gnd.n6510 gnd.n418 0.152939
R19096 gnd.n6518 gnd.n418 0.152939
R19097 gnd.n6519 gnd.n6518 0.152939
R19098 gnd.n6520 gnd.n6519 0.152939
R19099 gnd.n6520 gnd.n412 0.152939
R19100 gnd.n6528 gnd.n412 0.152939
R19101 gnd.n6529 gnd.n6528 0.152939
R19102 gnd.n6530 gnd.n6529 0.152939
R19103 gnd.n6530 gnd.n406 0.152939
R19104 gnd.n6538 gnd.n406 0.152939
R19105 gnd.n6540 gnd.n6539 0.152939
R19106 gnd.n6540 gnd.n400 0.152939
R19107 gnd.n6548 gnd.n400 0.152939
R19108 gnd.n6549 gnd.n6548 0.152939
R19109 gnd.n6550 gnd.n6549 0.152939
R19110 gnd.n6550 gnd.n394 0.152939
R19111 gnd.n6558 gnd.n394 0.152939
R19112 gnd.n6559 gnd.n6558 0.152939
R19113 gnd.n6560 gnd.n6559 0.152939
R19114 gnd.n6560 gnd.n388 0.152939
R19115 gnd.n6568 gnd.n388 0.152939
R19116 gnd.n6569 gnd.n6568 0.152939
R19117 gnd.n6570 gnd.n6569 0.152939
R19118 gnd.n6570 gnd.n382 0.152939
R19119 gnd.n6578 gnd.n382 0.152939
R19120 gnd.n6579 gnd.n6578 0.152939
R19121 gnd.n6580 gnd.n6579 0.152939
R19122 gnd.n6580 gnd.n376 0.152939
R19123 gnd.n6588 gnd.n376 0.152939
R19124 gnd.n6589 gnd.n6588 0.152939
R19125 gnd.n6590 gnd.n6589 0.152939
R19126 gnd.n6590 gnd.n370 0.152939
R19127 gnd.n6598 gnd.n370 0.152939
R19128 gnd.n6599 gnd.n6598 0.152939
R19129 gnd.n6600 gnd.n6599 0.152939
R19130 gnd.n6600 gnd.n364 0.152939
R19131 gnd.n6608 gnd.n364 0.152939
R19132 gnd.n6609 gnd.n6608 0.152939
R19133 gnd.n6610 gnd.n6609 0.152939
R19134 gnd.n6610 gnd.n358 0.152939
R19135 gnd.n6618 gnd.n358 0.152939
R19136 gnd.n6619 gnd.n6618 0.152939
R19137 gnd.n6620 gnd.n6619 0.152939
R19138 gnd.n6620 gnd.n352 0.152939
R19139 gnd.n6628 gnd.n352 0.152939
R19140 gnd.n6629 gnd.n6628 0.152939
R19141 gnd.n6630 gnd.n6629 0.152939
R19142 gnd.n6630 gnd.n346 0.152939
R19143 gnd.n6638 gnd.n346 0.152939
R19144 gnd.n6639 gnd.n6638 0.152939
R19145 gnd.n6640 gnd.n6639 0.152939
R19146 gnd.n6640 gnd.n340 0.152939
R19147 gnd.n6648 gnd.n340 0.152939
R19148 gnd.n6649 gnd.n6648 0.152939
R19149 gnd.n6650 gnd.n6649 0.152939
R19150 gnd.n6650 gnd.n334 0.152939
R19151 gnd.n6658 gnd.n334 0.152939
R19152 gnd.n6659 gnd.n6658 0.152939
R19153 gnd.n6660 gnd.n6659 0.152939
R19154 gnd.n6660 gnd.n328 0.152939
R19155 gnd.n6668 gnd.n328 0.152939
R19156 gnd.n6669 gnd.n6668 0.152939
R19157 gnd.n6670 gnd.n6669 0.152939
R19158 gnd.n6670 gnd.n322 0.152939
R19159 gnd.n6678 gnd.n322 0.152939
R19160 gnd.n6679 gnd.n6678 0.152939
R19161 gnd.n6680 gnd.n6679 0.152939
R19162 gnd.n6680 gnd.n316 0.152939
R19163 gnd.n6688 gnd.n316 0.152939
R19164 gnd.n6689 gnd.n6688 0.152939
R19165 gnd.n6690 gnd.n6689 0.152939
R19166 gnd.n6690 gnd.n310 0.152939
R19167 gnd.n6698 gnd.n310 0.152939
R19168 gnd.n6699 gnd.n6698 0.152939
R19169 gnd.n6700 gnd.n6699 0.152939
R19170 gnd.n6700 gnd.n304 0.152939
R19171 gnd.n6708 gnd.n304 0.152939
R19172 gnd.n6709 gnd.n6708 0.152939
R19173 gnd.n6710 gnd.n6709 0.152939
R19174 gnd.n6710 gnd.n298 0.152939
R19175 gnd.n6718 gnd.n298 0.152939
R19176 gnd.n6719 gnd.n6718 0.152939
R19177 gnd.n6720 gnd.n6719 0.152939
R19178 gnd.n6720 gnd.n292 0.152939
R19179 gnd.n6728 gnd.n292 0.152939
R19180 gnd.n6729 gnd.n6728 0.152939
R19181 gnd.n6730 gnd.n6729 0.152939
R19182 gnd.n6730 gnd.n286 0.152939
R19183 gnd.n6738 gnd.n286 0.152939
R19184 gnd.n6739 gnd.n6738 0.152939
R19185 gnd.n6740 gnd.n6739 0.152939
R19186 gnd.n6741 gnd.n6740 0.152939
R19187 gnd.n6741 gnd.n280 0.152939
R19188 gnd.n6751 gnd.n280 0.152939
R19189 gnd.n5648 gnd.n5647 0.152939
R19190 gnd.n5650 gnd.n5648 0.152939
R19191 gnd.n5650 gnd.n5649 0.152939
R19192 gnd.n5649 gnd.n273 0.152939
R19193 gnd.n274 gnd.n273 0.152939
R19194 gnd.n275 gnd.n274 0.152939
R19195 gnd.n278 gnd.n275 0.152939
R19196 gnd.n279 gnd.n278 0.152939
R19197 gnd.n6752 gnd.n279 0.152939
R19198 gnd.n6800 gnd.n6799 0.152939
R19199 gnd.n6801 gnd.n6800 0.152939
R19200 gnd.n6801 gnd.n199 0.152939
R19201 gnd.n6815 gnd.n199 0.152939
R19202 gnd.n6816 gnd.n6815 0.152939
R19203 gnd.n6817 gnd.n6816 0.152939
R19204 gnd.n6817 gnd.n183 0.152939
R19205 gnd.n6831 gnd.n183 0.152939
R19206 gnd.n6832 gnd.n6831 0.152939
R19207 gnd.n6833 gnd.n6832 0.152939
R19208 gnd.n6833 gnd.n165 0.152939
R19209 gnd.n6921 gnd.n165 0.152939
R19210 gnd.n6922 gnd.n6921 0.152939
R19211 gnd.n6923 gnd.n6922 0.152939
R19212 gnd.n6923 gnd.n88 0.152939
R19213 gnd.n7003 gnd.n88 0.152939
R19214 gnd.n7002 gnd.n89 0.152939
R19215 gnd.n91 gnd.n89 0.152939
R19216 gnd.n95 gnd.n91 0.152939
R19217 gnd.n96 gnd.n95 0.152939
R19218 gnd.n97 gnd.n96 0.152939
R19219 gnd.n98 gnd.n97 0.152939
R19220 gnd.n102 gnd.n98 0.152939
R19221 gnd.n103 gnd.n102 0.152939
R19222 gnd.n104 gnd.n103 0.152939
R19223 gnd.n105 gnd.n104 0.152939
R19224 gnd.n109 gnd.n105 0.152939
R19225 gnd.n110 gnd.n109 0.152939
R19226 gnd.n111 gnd.n110 0.152939
R19227 gnd.n112 gnd.n111 0.152939
R19228 gnd.n116 gnd.n112 0.152939
R19229 gnd.n117 gnd.n116 0.152939
R19230 gnd.n118 gnd.n117 0.152939
R19231 gnd.n119 gnd.n118 0.152939
R19232 gnd.n123 gnd.n119 0.152939
R19233 gnd.n124 gnd.n123 0.152939
R19234 gnd.n125 gnd.n124 0.152939
R19235 gnd.n126 gnd.n125 0.152939
R19236 gnd.n130 gnd.n126 0.152939
R19237 gnd.n131 gnd.n130 0.152939
R19238 gnd.n132 gnd.n131 0.152939
R19239 gnd.n133 gnd.n132 0.152939
R19240 gnd.n137 gnd.n133 0.152939
R19241 gnd.n138 gnd.n137 0.152939
R19242 gnd.n139 gnd.n138 0.152939
R19243 gnd.n140 gnd.n139 0.152939
R19244 gnd.n144 gnd.n140 0.152939
R19245 gnd.n145 gnd.n144 0.152939
R19246 gnd.n146 gnd.n145 0.152939
R19247 gnd.n147 gnd.n146 0.152939
R19248 gnd.n151 gnd.n147 0.152939
R19249 gnd.n152 gnd.n151 0.152939
R19250 gnd.n6933 gnd.n152 0.152939
R19251 gnd.n6933 gnd.n6932 0.152939
R19252 gnd.n5465 gnd.n5464 0.152939
R19253 gnd.n5465 gnd.n1260 0.152939
R19254 gnd.n5480 gnd.n1260 0.152939
R19255 gnd.n5481 gnd.n5480 0.152939
R19256 gnd.n5482 gnd.n5481 0.152939
R19257 gnd.n5483 gnd.n5482 0.152939
R19258 gnd.n5484 gnd.n5483 0.152939
R19259 gnd.n5485 gnd.n5484 0.152939
R19260 gnd.n5486 gnd.n5485 0.152939
R19261 gnd.n5487 gnd.n5486 0.152939
R19262 gnd.n5488 gnd.n5487 0.152939
R19263 gnd.n5489 gnd.n5488 0.152939
R19264 gnd.n5490 gnd.n5489 0.152939
R19265 gnd.n5491 gnd.n5490 0.152939
R19266 gnd.n5492 gnd.n5491 0.152939
R19267 gnd.n5493 gnd.n5492 0.152939
R19268 gnd.n5494 gnd.n5493 0.152939
R19269 gnd.n5495 gnd.n5494 0.152939
R19270 gnd.n5496 gnd.n5495 0.152939
R19271 gnd.n5497 gnd.n5496 0.152939
R19272 gnd.n5499 gnd.n5497 0.152939
R19273 gnd.n5499 gnd.n5498 0.152939
R19274 gnd.n5498 gnd.n238 0.152939
R19275 gnd.n239 gnd.n238 0.152939
R19276 gnd.n240 gnd.n239 0.152939
R19277 gnd.n241 gnd.n240 0.152939
R19278 gnd.n242 gnd.n241 0.152939
R19279 gnd.n243 gnd.n242 0.152939
R19280 gnd.n244 gnd.n243 0.152939
R19281 gnd.n245 gnd.n244 0.152939
R19282 gnd.n246 gnd.n245 0.152939
R19283 gnd.n247 gnd.n246 0.152939
R19284 gnd.n248 gnd.n247 0.152939
R19285 gnd.n249 gnd.n248 0.152939
R19286 gnd.n250 gnd.n249 0.152939
R19287 gnd.n251 gnd.n250 0.152939
R19288 gnd.n252 gnd.n251 0.152939
R19289 gnd.n253 gnd.n252 0.152939
R19290 gnd.n255 gnd.n253 0.152939
R19291 gnd.n255 gnd.n254 0.152939
R19292 gnd.n254 gnd.n158 0.152939
R19293 gnd.n6931 gnd.n158 0.152939
R19294 gnd.n5369 gnd.n5368 0.152939
R19295 gnd.n5369 gnd.n5365 0.152939
R19296 gnd.n5377 gnd.n5365 0.152939
R19297 gnd.n5378 gnd.n5377 0.152939
R19298 gnd.n5379 gnd.n5378 0.152939
R19299 gnd.n5379 gnd.n5361 0.152939
R19300 gnd.n5387 gnd.n5361 0.152939
R19301 gnd.n5388 gnd.n5387 0.152939
R19302 gnd.n5389 gnd.n5388 0.152939
R19303 gnd.n5389 gnd.n5357 0.152939
R19304 gnd.n5397 gnd.n5357 0.152939
R19305 gnd.n5398 gnd.n5397 0.152939
R19306 gnd.n5400 gnd.n5398 0.152939
R19307 gnd.n5400 gnd.n5399 0.152939
R19308 gnd.n5399 gnd.n1290 0.152939
R19309 gnd.n5413 gnd.n5412 0.152939
R19310 gnd.n5413 gnd.n1286 0.152939
R19311 gnd.n5421 gnd.n1286 0.152939
R19312 gnd.n5422 gnd.n5421 0.152939
R19313 gnd.n5423 gnd.n5422 0.152939
R19314 gnd.n5423 gnd.n1282 0.152939
R19315 gnd.n5431 gnd.n1282 0.152939
R19316 gnd.n5432 gnd.n5431 0.152939
R19317 gnd.n5433 gnd.n5432 0.152939
R19318 gnd.n5433 gnd.n1278 0.152939
R19319 gnd.n5441 gnd.n1278 0.152939
R19320 gnd.n5442 gnd.n5441 0.152939
R19321 gnd.n5443 gnd.n5442 0.152939
R19322 gnd.n5443 gnd.n1274 0.152939
R19323 gnd.n5451 gnd.n1274 0.152939
R19324 gnd.n5452 gnd.n5451 0.152939
R19325 gnd.n5454 gnd.n5452 0.152939
R19326 gnd.n5454 gnd.n5453 0.152939
R19327 gnd.n5453 gnd.n1267 0.152939
R19328 gnd.n5463 gnd.n1267 0.152939
R19329 gnd.n1134 gnd.n1133 0.152939
R19330 gnd.n1135 gnd.n1134 0.152939
R19331 gnd.n1255 gnd.n1135 0.152939
R19332 gnd.n5547 gnd.n1255 0.152939
R19333 gnd.n5548 gnd.n5547 0.152939
R19334 gnd.n5549 gnd.n5548 0.152939
R19335 gnd.n5550 gnd.n5549 0.152939
R19336 gnd.n5550 gnd.n1227 0.152939
R19337 gnd.n5578 gnd.n1227 0.152939
R19338 gnd.n5579 gnd.n5578 0.152939
R19339 gnd.n5580 gnd.n5579 0.152939
R19340 gnd.n5582 gnd.n5580 0.152939
R19341 gnd.n5582 gnd.n5581 0.152939
R19342 gnd.n5581 gnd.n1199 0.152939
R19343 gnd.n1199 gnd.n214 0.152939
R19344 gnd.n6799 gnd.n214 0.152939
R19345 gnd.n3963 gnd.n3962 0.152939
R19346 gnd.n3964 gnd.n3963 0.152939
R19347 gnd.n3964 gnd.n1985 0.152939
R19348 gnd.n4026 gnd.n1985 0.152939
R19349 gnd.n4027 gnd.n4026 0.152939
R19350 gnd.n4028 gnd.n4027 0.152939
R19351 gnd.n4028 gnd.n1981 0.152939
R19352 gnd.n4034 gnd.n1981 0.152939
R19353 gnd.n4035 gnd.n4034 0.152939
R19354 gnd.n4036 gnd.n4035 0.152939
R19355 gnd.n4036 gnd.n1977 0.152939
R19356 gnd.n4042 gnd.n1977 0.152939
R19357 gnd.n4043 gnd.n4042 0.152939
R19358 gnd.n4044 gnd.n4043 0.152939
R19359 gnd.n4044 gnd.n1973 0.152939
R19360 gnd.n4050 gnd.n1973 0.152939
R19361 gnd.n4051 gnd.n4050 0.152939
R19362 gnd.n4052 gnd.n4051 0.152939
R19363 gnd.n4052 gnd.n1967 0.152939
R19364 gnd.n4193 gnd.n1967 0.152939
R19365 gnd.n4194 gnd.n4193 0.152939
R19366 gnd.n4195 gnd.n4194 0.152939
R19367 gnd.n4195 gnd.n1961 0.152939
R19368 gnd.n4207 gnd.n1961 0.152939
R19369 gnd.n4208 gnd.n4207 0.152939
R19370 gnd.n4209 gnd.n4208 0.152939
R19371 gnd.n4209 gnd.n1953 0.152939
R19372 gnd.n4221 gnd.n1953 0.152939
R19373 gnd.n4222 gnd.n4221 0.152939
R19374 gnd.n4223 gnd.n4222 0.152939
R19375 gnd.n4223 gnd.n1945 0.152939
R19376 gnd.n4235 gnd.n1945 0.152939
R19377 gnd.n4236 gnd.n4235 0.152939
R19378 gnd.n4237 gnd.n4236 0.152939
R19379 gnd.n4237 gnd.n1668 0.152939
R19380 gnd.n4424 gnd.n1668 0.152939
R19381 gnd.n4425 gnd.n4424 0.152939
R19382 gnd.n4426 gnd.n4425 0.152939
R19383 gnd.n4426 gnd.n1650 0.152939
R19384 gnd.n4480 gnd.n1650 0.152939
R19385 gnd.n4481 gnd.n4480 0.152939
R19386 gnd.n4482 gnd.n4481 0.152939
R19387 gnd.n4482 gnd.n1629 0.152939
R19388 gnd.n4511 gnd.n1629 0.152939
R19389 gnd.n4512 gnd.n4511 0.152939
R19390 gnd.n4513 gnd.n4512 0.152939
R19391 gnd.n4514 gnd.n4513 0.152939
R19392 gnd.n4514 gnd.n1609 0.152939
R19393 gnd.n4541 gnd.n1609 0.152939
R19394 gnd.n4542 gnd.n4541 0.152939
R19395 gnd.n4543 gnd.n4542 0.152939
R19396 gnd.n4544 gnd.n4543 0.152939
R19397 gnd.n4545 gnd.n4544 0.152939
R19398 gnd.n4546 gnd.n4545 0.152939
R19399 gnd.n4546 gnd.n1562 0.152939
R19400 gnd.n4625 gnd.n1562 0.152939
R19401 gnd.n4626 gnd.n4625 0.152939
R19402 gnd.n4627 gnd.n4626 0.152939
R19403 gnd.n4627 gnd.n1539 0.152939
R19404 gnd.n4665 gnd.n1539 0.152939
R19405 gnd.n4666 gnd.n4665 0.152939
R19406 gnd.n4667 gnd.n4666 0.152939
R19407 gnd.n4667 gnd.n1517 0.152939
R19408 gnd.n4719 gnd.n1517 0.152939
R19409 gnd.n4720 gnd.n4719 0.152939
R19410 gnd.n4721 gnd.n4720 0.152939
R19411 gnd.n4721 gnd.n1498 0.152939
R19412 gnd.n4744 gnd.n1498 0.152939
R19413 gnd.n4745 gnd.n4744 0.152939
R19414 gnd.n4746 gnd.n4745 0.152939
R19415 gnd.n4746 gnd.n1476 0.152939
R19416 gnd.n4803 gnd.n1476 0.152939
R19417 gnd.n4804 gnd.n4803 0.152939
R19418 gnd.n4805 gnd.n4804 0.152939
R19419 gnd.n4805 gnd.n1454 0.152939
R19420 gnd.n4832 gnd.n1454 0.152939
R19421 gnd.n4833 gnd.n4832 0.152939
R19422 gnd.n4834 gnd.n4833 0.152939
R19423 gnd.n4835 gnd.n4834 0.152939
R19424 gnd.n4835 gnd.n1426 0.152939
R19425 gnd.n4887 gnd.n1426 0.152939
R19426 gnd.n4888 gnd.n4887 0.152939
R19427 gnd.n4889 gnd.n4888 0.152939
R19428 gnd.n4889 gnd.n1409 0.152939
R19429 gnd.n4913 gnd.n1409 0.152939
R19430 gnd.n4914 gnd.n4913 0.152939
R19431 gnd.n4915 gnd.n4914 0.152939
R19432 gnd.n4917 gnd.n4915 0.152939
R19433 gnd.n4917 gnd.n4916 0.152939
R19434 gnd.n4916 gnd.n1347 0.152939
R19435 gnd.n1348 gnd.n1347 0.152939
R19436 gnd.n1349 gnd.n1348 0.152939
R19437 gnd.n1357 gnd.n1349 0.152939
R19438 gnd.n1358 gnd.n1357 0.152939
R19439 gnd.n1359 gnd.n1358 0.152939
R19440 gnd.n1360 gnd.n1359 0.152939
R19441 gnd.n1361 gnd.n1360 0.152939
R19442 gnd.n1370 gnd.n1361 0.152939
R19443 gnd.n1371 gnd.n1370 0.152939
R19444 gnd.n1372 gnd.n1371 0.152939
R19445 gnd.n1373 gnd.n1372 0.152939
R19446 gnd.n5152 gnd.n1373 0.152939
R19447 gnd.n5154 gnd.n5152 0.152939
R19448 gnd.n5154 gnd.n5153 0.152939
R19449 gnd.n5153 gnd.n1112 0.152939
R19450 gnd.n1113 gnd.n1112 0.152939
R19451 gnd.n1114 gnd.n1113 0.152939
R19452 gnd.n1120 gnd.n1114 0.152939
R19453 gnd.n1121 gnd.n1120 0.152939
R19454 gnd.n1122 gnd.n1121 0.152939
R19455 gnd.n1123 gnd.n1122 0.152939
R19456 gnd.n5530 gnd.n1123 0.152939
R19457 gnd.n5531 gnd.n5530 0.152939
R19458 gnd.n5536 gnd.n5531 0.152939
R19459 gnd.n5537 gnd.n5536 0.152939
R19460 gnd.n5538 gnd.n5537 0.152939
R19461 gnd.n5539 gnd.n5538 0.152939
R19462 gnd.n5539 gnd.n1237 0.152939
R19463 gnd.n5567 gnd.n1237 0.152939
R19464 gnd.n5568 gnd.n5567 0.152939
R19465 gnd.n5569 gnd.n5568 0.152939
R19466 gnd.n5570 gnd.n5569 0.152939
R19467 gnd.n5570 gnd.n1209 0.152939
R19468 gnd.n5599 gnd.n1209 0.152939
R19469 gnd.n5600 gnd.n5599 0.152939
R19470 gnd.n5601 gnd.n5600 0.152939
R19471 gnd.n5602 gnd.n5601 0.152939
R19472 gnd.n3639 gnd.n3633 0.152939
R19473 gnd.n3635 gnd.n3633 0.152939
R19474 gnd.n3635 gnd.n3634 0.152939
R19475 gnd.n3634 gnd.n2085 0.152939
R19476 gnd.n2085 gnd.n2083 0.152939
R19477 gnd.n3819 gnd.n2083 0.152939
R19478 gnd.n3820 gnd.n3819 0.152939
R19479 gnd.n3822 gnd.n3820 0.152939
R19480 gnd.n3822 gnd.n3821 0.152939
R19481 gnd.n3821 gnd.n2075 0.152939
R19482 gnd.n2076 gnd.n2075 0.152939
R19483 gnd.n2077 gnd.n2076 0.152939
R19484 gnd.n2077 gnd.n2065 0.152939
R19485 gnd.n3876 gnd.n2065 0.152939
R19486 gnd.n3877 gnd.n3876 0.152939
R19487 gnd.n3878 gnd.n3877 0.152939
R19488 gnd.n3879 gnd.n3878 0.152939
R19489 gnd.n3879 gnd.n2052 0.152939
R19490 gnd.n3923 gnd.n2052 0.152939
R19491 gnd.n3924 gnd.n3923 0.152939
R19492 gnd.n3789 gnd.n2102 0.152939
R19493 gnd.n3594 gnd.n2102 0.152939
R19494 gnd.n3594 gnd.n3593 0.152939
R19495 gnd.n3601 gnd.n3593 0.152939
R19496 gnd.n3602 gnd.n3601 0.152939
R19497 gnd.n3603 gnd.n3602 0.152939
R19498 gnd.n3603 gnd.n3591 0.152939
R19499 gnd.n3611 gnd.n3591 0.152939
R19500 gnd.n3612 gnd.n3611 0.152939
R19501 gnd.n3613 gnd.n3612 0.152939
R19502 gnd.n3613 gnd.n3589 0.152939
R19503 gnd.n3621 gnd.n3589 0.152939
R19504 gnd.n3622 gnd.n3621 0.152939
R19505 gnd.n3623 gnd.n3622 0.152939
R19506 gnd.n3623 gnd.n3587 0.152939
R19507 gnd.n3631 gnd.n3587 0.152939
R19508 gnd.n3632 gnd.n3631 0.152939
R19509 gnd.n3640 gnd.n3632 0.152939
R19510 gnd.n3800 gnd.n3790 0.152939
R19511 gnd.n3800 gnd.n3799 0.152939
R19512 gnd.n3799 gnd.n3798 0.152939
R19513 gnd.n3798 gnd.n3791 0.152939
R19514 gnd.n3793 gnd.n3791 0.152939
R19515 gnd.n3793 gnd.n3792 0.152939
R19516 gnd.n3792 gnd.n847 0.152939
R19517 gnd.n848 gnd.n847 0.152939
R19518 gnd.n849 gnd.n848 0.152939
R19519 gnd.n867 gnd.n849 0.152939
R19520 gnd.n868 gnd.n867 0.152939
R19521 gnd.n869 gnd.n868 0.152939
R19522 gnd.n870 gnd.n869 0.152939
R19523 gnd.n888 gnd.n870 0.152939
R19524 gnd.n889 gnd.n888 0.152939
R19525 gnd.n890 gnd.n889 0.152939
R19526 gnd.n891 gnd.n890 0.152939
R19527 gnd.n3912 gnd.n891 0.152939
R19528 gnd.n3913 gnd.n3912 0.152939
R19529 gnd.n3913 gnd.n2032 0.152939
R19530 gnd.n3932 gnd.n2032 0.152939
R19531 gnd.n3933 gnd.n3932 0.152939
R19532 gnd.n3934 gnd.n3933 0.152939
R19533 gnd.n3936 gnd.n3934 0.152939
R19534 gnd.n3936 gnd.n3935 0.152939
R19535 gnd.n3935 gnd.n916 0.152939
R19536 gnd.n917 gnd.n916 0.152939
R19537 gnd.n918 gnd.n917 0.152939
R19538 gnd.n934 gnd.n918 0.152939
R19539 gnd.n935 gnd.n934 0.152939
R19540 gnd.n936 gnd.n935 0.152939
R19541 gnd.n937 gnd.n936 0.152939
R19542 gnd.n956 gnd.n937 0.152939
R19543 gnd.n957 gnd.n956 0.152939
R19544 gnd.n958 gnd.n957 0.152939
R19545 gnd.n959 gnd.n958 0.152939
R19546 gnd.n977 gnd.n959 0.152939
R19547 gnd.n978 gnd.n977 0.152939
R19548 gnd.n979 gnd.n978 0.152939
R19549 gnd.n980 gnd.n979 0.152939
R19550 gnd.n998 gnd.n980 0.152939
R19551 gnd.n5851 gnd.n998 0.152939
R19552 gnd.n5905 gnd.n900 0.152939
R19553 gnd.n925 gnd.n900 0.152939
R19554 gnd.n926 gnd.n925 0.152939
R19555 gnd.n927 gnd.n926 0.152939
R19556 gnd.n945 gnd.n927 0.152939
R19557 gnd.n946 gnd.n945 0.152939
R19558 gnd.n947 gnd.n946 0.152939
R19559 gnd.n948 gnd.n947 0.152939
R19560 gnd.n966 gnd.n948 0.152939
R19561 gnd.n967 gnd.n966 0.152939
R19562 gnd.n968 gnd.n967 0.152939
R19563 gnd.n969 gnd.n968 0.152939
R19564 gnd.n988 gnd.n969 0.152939
R19565 gnd.n989 gnd.n988 0.152939
R19566 gnd.n990 gnd.n989 0.152939
R19567 gnd.n991 gnd.n990 0.152939
R19568 gnd.n1829 gnd.n1828 0.152939
R19569 gnd.n1830 gnd.n1829 0.152939
R19570 gnd.n1831 gnd.n1830 0.152939
R19571 gnd.n1832 gnd.n1831 0.152939
R19572 gnd.n1833 gnd.n1832 0.152939
R19573 gnd.n1834 gnd.n1833 0.152939
R19574 gnd.n1835 gnd.n1834 0.152939
R19575 gnd.n1836 gnd.n1835 0.152939
R19576 gnd.n1837 gnd.n1836 0.152939
R19577 gnd.n1838 gnd.n1837 0.152939
R19578 gnd.n1839 gnd.n1838 0.152939
R19579 gnd.n1840 gnd.n1839 0.152939
R19580 gnd.n1841 gnd.n1840 0.152939
R19581 gnd.n1842 gnd.n1841 0.152939
R19582 gnd.n1842 gnd.n1812 0.152939
R19583 gnd.n4344 gnd.n4343 0.152939
R19584 gnd.n4343 gnd.n1813 0.152939
R19585 gnd.n1873 gnd.n1813 0.152939
R19586 gnd.n1874 gnd.n1873 0.152939
R19587 gnd.n1875 gnd.n1874 0.152939
R19588 gnd.n1876 gnd.n1875 0.152939
R19589 gnd.n1880 gnd.n1876 0.152939
R19590 gnd.n1881 gnd.n1880 0.152939
R19591 gnd.n1882 gnd.n1881 0.152939
R19592 gnd.n1883 gnd.n1882 0.152939
R19593 gnd.n1887 gnd.n1883 0.152939
R19594 gnd.n1888 gnd.n1887 0.152939
R19595 gnd.n1889 gnd.n1888 0.152939
R19596 gnd.n1890 gnd.n1889 0.152939
R19597 gnd.n1894 gnd.n1890 0.152939
R19598 gnd.n1895 gnd.n1894 0.152939
R19599 gnd.n1896 gnd.n1895 0.152939
R19600 gnd.n1897 gnd.n1896 0.152939
R19601 gnd.n1902 gnd.n1897 0.152939
R19602 gnd.n4306 gnd.n1902 0.152939
R19603 gnd.n3703 gnd.n3688 0.152939
R19604 gnd.n3703 gnd.n3702 0.152939
R19605 gnd.n3702 gnd.n3701 0.152939
R19606 gnd.n3701 gnd.n3691 0.152939
R19607 gnd.n3692 gnd.n3691 0.152939
R19608 gnd.n3694 gnd.n3692 0.152939
R19609 gnd.n3694 gnd.n3693 0.152939
R19610 gnd.n3693 gnd.n2081 0.152939
R19611 gnd.n2081 gnd.n2079 0.152939
R19612 gnd.n3830 gnd.n2079 0.152939
R19613 gnd.n3831 gnd.n3830 0.152939
R19614 gnd.n3832 gnd.n3831 0.152939
R19615 gnd.n3833 gnd.n3832 0.152939
R19616 gnd.n3834 gnd.n3833 0.152939
R19617 gnd.n3834 gnd.n2062 0.152939
R19618 gnd.n3886 gnd.n2062 0.152939
R19619 gnd.n3887 gnd.n3886 0.152939
R19620 gnd.n3888 gnd.n3887 0.152939
R19621 gnd.n3889 gnd.n3888 0.152939
R19622 gnd.n3889 gnd.n2033 0.152939
R19623 gnd.n3931 gnd.n2033 0.152939
R19624 gnd.n3931 gnd.n2034 0.152939
R19625 gnd.n2036 gnd.n2034 0.152939
R19626 gnd.n2037 gnd.n2036 0.152939
R19627 gnd.n2038 gnd.n2037 0.152939
R19628 gnd.n2039 gnd.n2038 0.152939
R19629 gnd.n2040 gnd.n2039 0.152939
R19630 gnd.n2040 gnd.n2003 0.152939
R19631 gnd.n3980 gnd.n2003 0.152939
R19632 gnd.n3981 gnd.n3980 0.152939
R19633 gnd.n3982 gnd.n3981 0.152939
R19634 gnd.n3982 gnd.n2001 0.152939
R19635 gnd.n3988 gnd.n2001 0.152939
R19636 gnd.n3989 gnd.n3988 0.152939
R19637 gnd.n3990 gnd.n3989 0.152939
R19638 gnd.n3990 gnd.n1999 0.152939
R19639 gnd.n3999 gnd.n1999 0.152939
R19640 gnd.n4000 gnd.n3999 0.152939
R19641 gnd.n4002 gnd.n4000 0.152939
R19642 gnd.n4002 gnd.n4001 0.152939
R19643 gnd.n4001 gnd.n1903 0.152939
R19644 gnd.n4305 gnd.n1903 0.152939
R19645 gnd.n3646 gnd.n3645 0.152939
R19646 gnd.n3647 gnd.n3646 0.152939
R19647 gnd.n3648 gnd.n3647 0.152939
R19648 gnd.n3649 gnd.n3648 0.152939
R19649 gnd.n3650 gnd.n3649 0.152939
R19650 gnd.n3651 gnd.n3650 0.152939
R19651 gnd.n3652 gnd.n3651 0.152939
R19652 gnd.n3653 gnd.n3652 0.152939
R19653 gnd.n3654 gnd.n3653 0.152939
R19654 gnd.n3655 gnd.n3654 0.152939
R19655 gnd.n3656 gnd.n3655 0.152939
R19656 gnd.n3657 gnd.n3656 0.152939
R19657 gnd.n3658 gnd.n3657 0.152939
R19658 gnd.n3659 gnd.n3658 0.152939
R19659 gnd.n3660 gnd.n3659 0.152939
R19660 gnd.n3661 gnd.n3660 0.152939
R19661 gnd.n3662 gnd.n3661 0.152939
R19662 gnd.n3665 gnd.n3662 0.152939
R19663 gnd.n3666 gnd.n3665 0.152939
R19664 gnd.n3667 gnd.n3666 0.152939
R19665 gnd.n3668 gnd.n3667 0.152939
R19666 gnd.n3669 gnd.n3668 0.152939
R19667 gnd.n3670 gnd.n3669 0.152939
R19668 gnd.n3671 gnd.n3670 0.152939
R19669 gnd.n3672 gnd.n3671 0.152939
R19670 gnd.n3673 gnd.n3672 0.152939
R19671 gnd.n3674 gnd.n3673 0.152939
R19672 gnd.n3675 gnd.n3674 0.152939
R19673 gnd.n3676 gnd.n3675 0.152939
R19674 gnd.n3677 gnd.n3676 0.152939
R19675 gnd.n3678 gnd.n3677 0.152939
R19676 gnd.n3679 gnd.n3678 0.152939
R19677 gnd.n3680 gnd.n3679 0.152939
R19678 gnd.n3681 gnd.n3680 0.152939
R19679 gnd.n3682 gnd.n3681 0.152939
R19680 gnd.n3711 gnd.n3682 0.152939
R19681 gnd.n3711 gnd.n3710 0.152939
R19682 gnd.n3710 gnd.n3709 0.152939
R19683 gnd.n3806 gnd.n2092 0.152939
R19684 gnd.n3807 gnd.n3806 0.152939
R19685 gnd.n3809 gnd.n3807 0.152939
R19686 gnd.n3809 gnd.n3808 0.152939
R19687 gnd.n3808 gnd.n835 0.152939
R19688 gnd.n836 gnd.n835 0.152939
R19689 gnd.n837 gnd.n836 0.152939
R19690 gnd.n856 gnd.n837 0.152939
R19691 gnd.n857 gnd.n856 0.152939
R19692 gnd.n858 gnd.n857 0.152939
R19693 gnd.n859 gnd.n858 0.152939
R19694 gnd.n878 gnd.n859 0.152939
R19695 gnd.n879 gnd.n878 0.152939
R19696 gnd.n880 gnd.n879 0.152939
R19697 gnd.n881 gnd.n880 0.152939
R19698 gnd.n5905 gnd.n881 0.152939
R19699 gnd.n3850 gnd.n3849 0.152939
R19700 gnd.n3856 gnd.n3849 0.152939
R19701 gnd.n3857 gnd.n3856 0.152939
R19702 gnd.n3858 gnd.n3857 0.152939
R19703 gnd.n3858 gnd.n2071 0.152939
R19704 gnd.n3864 gnd.n2071 0.152939
R19705 gnd.n3865 gnd.n3864 0.152939
R19706 gnd.n3866 gnd.n3865 0.152939
R19707 gnd.n3867 gnd.n3866 0.152939
R19708 gnd.n6118 gnd.n658 0.152939
R19709 gnd.n663 gnd.n658 0.152939
R19710 gnd.n664 gnd.n663 0.152939
R19711 gnd.n665 gnd.n664 0.152939
R19712 gnd.n670 gnd.n665 0.152939
R19713 gnd.n671 gnd.n670 0.152939
R19714 gnd.n672 gnd.n671 0.152939
R19715 gnd.n673 gnd.n672 0.152939
R19716 gnd.n678 gnd.n673 0.152939
R19717 gnd.n679 gnd.n678 0.152939
R19718 gnd.n680 gnd.n679 0.152939
R19719 gnd.n681 gnd.n680 0.152939
R19720 gnd.n686 gnd.n681 0.152939
R19721 gnd.n687 gnd.n686 0.152939
R19722 gnd.n688 gnd.n687 0.152939
R19723 gnd.n689 gnd.n688 0.152939
R19724 gnd.n694 gnd.n689 0.152939
R19725 gnd.n695 gnd.n694 0.152939
R19726 gnd.n696 gnd.n695 0.152939
R19727 gnd.n697 gnd.n696 0.152939
R19728 gnd.n702 gnd.n697 0.152939
R19729 gnd.n703 gnd.n702 0.152939
R19730 gnd.n704 gnd.n703 0.152939
R19731 gnd.n705 gnd.n704 0.152939
R19732 gnd.n710 gnd.n705 0.152939
R19733 gnd.n711 gnd.n710 0.152939
R19734 gnd.n712 gnd.n711 0.152939
R19735 gnd.n713 gnd.n712 0.152939
R19736 gnd.n718 gnd.n713 0.152939
R19737 gnd.n719 gnd.n718 0.152939
R19738 gnd.n720 gnd.n719 0.152939
R19739 gnd.n721 gnd.n720 0.152939
R19740 gnd.n726 gnd.n721 0.152939
R19741 gnd.n727 gnd.n726 0.152939
R19742 gnd.n728 gnd.n727 0.152939
R19743 gnd.n729 gnd.n728 0.152939
R19744 gnd.n734 gnd.n729 0.152939
R19745 gnd.n735 gnd.n734 0.152939
R19746 gnd.n736 gnd.n735 0.152939
R19747 gnd.n737 gnd.n736 0.152939
R19748 gnd.n742 gnd.n737 0.152939
R19749 gnd.n743 gnd.n742 0.152939
R19750 gnd.n744 gnd.n743 0.152939
R19751 gnd.n745 gnd.n744 0.152939
R19752 gnd.n750 gnd.n745 0.152939
R19753 gnd.n751 gnd.n750 0.152939
R19754 gnd.n752 gnd.n751 0.152939
R19755 gnd.n753 gnd.n752 0.152939
R19756 gnd.n758 gnd.n753 0.152939
R19757 gnd.n759 gnd.n758 0.152939
R19758 gnd.n760 gnd.n759 0.152939
R19759 gnd.n761 gnd.n760 0.152939
R19760 gnd.n766 gnd.n761 0.152939
R19761 gnd.n767 gnd.n766 0.152939
R19762 gnd.n768 gnd.n767 0.152939
R19763 gnd.n769 gnd.n768 0.152939
R19764 gnd.n774 gnd.n769 0.152939
R19765 gnd.n775 gnd.n774 0.152939
R19766 gnd.n776 gnd.n775 0.152939
R19767 gnd.n777 gnd.n776 0.152939
R19768 gnd.n782 gnd.n777 0.152939
R19769 gnd.n783 gnd.n782 0.152939
R19770 gnd.n784 gnd.n783 0.152939
R19771 gnd.n785 gnd.n784 0.152939
R19772 gnd.n790 gnd.n785 0.152939
R19773 gnd.n791 gnd.n790 0.152939
R19774 gnd.n792 gnd.n791 0.152939
R19775 gnd.n793 gnd.n792 0.152939
R19776 gnd.n798 gnd.n793 0.152939
R19777 gnd.n799 gnd.n798 0.152939
R19778 gnd.n800 gnd.n799 0.152939
R19779 gnd.n801 gnd.n800 0.152939
R19780 gnd.n806 gnd.n801 0.152939
R19781 gnd.n807 gnd.n806 0.152939
R19782 gnd.n808 gnd.n807 0.152939
R19783 gnd.n809 gnd.n808 0.152939
R19784 gnd.n814 gnd.n809 0.152939
R19785 gnd.n815 gnd.n814 0.152939
R19786 gnd.n816 gnd.n815 0.152939
R19787 gnd.n817 gnd.n816 0.152939
R19788 gnd.n822 gnd.n817 0.152939
R19789 gnd.n823 gnd.n822 0.152939
R19790 gnd.n824 gnd.n823 0.152939
R19791 gnd.n825 gnd.n824 0.152939
R19792 gnd.n5124 gnd.n4980 0.152939
R19793 gnd.n5125 gnd.n5124 0.152939
R19794 gnd.n5126 gnd.n5125 0.152939
R19795 gnd.n5126 gnd.n4976 0.152939
R19796 gnd.n5137 gnd.n4976 0.152939
R19797 gnd.n5138 gnd.n5137 0.152939
R19798 gnd.n5139 gnd.n5138 0.152939
R19799 gnd.n5139 gnd.n4972 0.152939
R19800 gnd.n5146 gnd.n4972 0.152939
R19801 gnd.n4278 gnd.n1927 0.152939
R19802 gnd.n4274 gnd.n1927 0.152939
R19803 gnd.n4274 gnd.n4273 0.152939
R19804 gnd.n4273 gnd.n4272 0.152939
R19805 gnd.n4272 gnd.n1932 0.152939
R19806 gnd.n4268 gnd.n1932 0.152939
R19807 gnd.n4268 gnd.n4267 0.152939
R19808 gnd.n4267 gnd.n4266 0.152939
R19809 gnd.n4266 gnd.n1937 0.152939
R19810 gnd.n4262 gnd.n1937 0.152939
R19811 gnd.n4262 gnd.n4261 0.152939
R19812 gnd.n4261 gnd.n4260 0.152939
R19813 gnd.n4260 gnd.n1942 0.152939
R19814 gnd.n4256 gnd.n1942 0.152939
R19815 gnd.n4256 gnd.n4255 0.152939
R19816 gnd.n4255 gnd.n4254 0.152939
R19817 gnd.n4254 gnd.n4248 0.152939
R19818 gnd.n4248 gnd.n1642 0.152939
R19819 gnd.n4490 gnd.n1642 0.152939
R19820 gnd.n4491 gnd.n4490 0.152939
R19821 gnd.n4492 gnd.n4491 0.152939
R19822 gnd.n4492 gnd.n1622 0.152939
R19823 gnd.n4523 gnd.n1622 0.152939
R19824 gnd.n4524 gnd.n4523 0.152939
R19825 gnd.n4525 gnd.n4524 0.152939
R19826 gnd.n4525 gnd.n1596 0.152939
R19827 gnd.n4568 gnd.n1596 0.152939
R19828 gnd.n4569 gnd.n4568 0.152939
R19829 gnd.n4572 gnd.n4569 0.152939
R19830 gnd.n4572 gnd.n4571 0.152939
R19831 gnd.n4571 gnd.n4570 0.152939
R19832 gnd.n4570 gnd.n1580 0.152939
R19833 gnd.n4598 gnd.n1580 0.152939
R19834 gnd.n4599 gnd.n4598 0.152939
R19835 gnd.n4600 gnd.n4599 0.152939
R19836 gnd.n4600 gnd.n1555 0.152939
R19837 gnd.n4648 gnd.n1555 0.152939
R19838 gnd.n4648 gnd.n4647 0.152939
R19839 gnd.n4647 gnd.n4646 0.152939
R19840 gnd.n4646 gnd.n1532 0.152939
R19841 gnd.n4704 gnd.n1532 0.152939
R19842 gnd.n4704 gnd.n4703 0.152939
R19843 gnd.n4703 gnd.n4702 0.152939
R19844 gnd.n4702 gnd.n1533 0.152939
R19845 gnd.n4698 gnd.n1533 0.152939
R19846 gnd.n4698 gnd.n4697 0.152939
R19847 gnd.n4697 gnd.n4696 0.152939
R19848 gnd.n4696 gnd.n4689 0.152939
R19849 gnd.n4692 gnd.n4689 0.152939
R19850 gnd.n4692 gnd.n1469 0.152939
R19851 gnd.n4813 gnd.n1469 0.152939
R19852 gnd.n4814 gnd.n4813 0.152939
R19853 gnd.n4816 gnd.n4814 0.152939
R19854 gnd.n4816 gnd.n4815 0.152939
R19855 gnd.n4815 gnd.n1441 0.152939
R19856 gnd.n4852 gnd.n1441 0.152939
R19857 gnd.n4853 gnd.n4852 0.152939
R19858 gnd.n4871 gnd.n4853 0.152939
R19859 gnd.n4871 gnd.n4870 0.152939
R19860 gnd.n4870 gnd.n4869 0.152939
R19861 gnd.n4869 gnd.n4854 0.152939
R19862 gnd.n4865 gnd.n4854 0.152939
R19863 gnd.n4865 gnd.n4864 0.152939
R19864 gnd.n4864 gnd.n4863 0.152939
R19865 gnd.n4863 gnd.n1390 0.152939
R19866 gnd.n4943 gnd.n1390 0.152939
R19867 gnd.n4944 gnd.n4943 0.152939
R19868 gnd.n4946 gnd.n4944 0.152939
R19869 gnd.n4946 gnd.n4945 0.152939
R19870 gnd.n4945 gnd.n1386 0.152939
R19871 gnd.n4954 gnd.n1386 0.152939
R19872 gnd.n4955 gnd.n4954 0.152939
R19873 gnd.n4956 gnd.n4955 0.152939
R19874 gnd.n4956 gnd.n1384 0.152939
R19875 gnd.n4962 gnd.n1384 0.152939
R19876 gnd.n4963 gnd.n4962 0.152939
R19877 gnd.n4964 gnd.n4963 0.152939
R19878 gnd.n4964 gnd.n1382 0.152939
R19879 gnd.n4970 gnd.n1382 0.152939
R19880 gnd.n4971 gnd.n4970 0.152939
R19881 gnd.n5148 gnd.n4971 0.152939
R19882 gnd.n5148 gnd.n5147 0.152939
R19883 gnd.n4291 gnd.n1908 0.152939
R19884 gnd.n4291 gnd.n4290 0.152939
R19885 gnd.n4290 gnd.n4289 0.152939
R19886 gnd.n4289 gnd.n1915 0.152939
R19887 gnd.n4285 gnd.n1915 0.152939
R19888 gnd.n4285 gnd.n4284 0.152939
R19889 gnd.n4284 gnd.n1922 0.152939
R19890 gnd.n4280 gnd.n1922 0.152939
R19891 gnd.n4280 gnd.n4279 0.152939
R19892 gnd.n3951 gnd.n2018 0.152939
R19893 gnd.n3952 gnd.n3951 0.152939
R19894 gnd.n3953 gnd.n3952 0.152939
R19895 gnd.n3953 gnd.n2006 0.152939
R19896 gnd.n3972 gnd.n2006 0.152939
R19897 gnd.n3973 gnd.n3972 0.152939
R19898 gnd.n3974 gnd.n3973 0.152939
R19899 gnd.n3974 gnd.n1991 0.152939
R19900 gnd.n4019 gnd.n1991 0.152939
R19901 gnd.n4019 gnd.n4018 0.152939
R19902 gnd.n4018 gnd.n4017 0.152939
R19903 gnd.n4017 gnd.n1992 0.152939
R19904 gnd.n4013 gnd.n1992 0.152939
R19905 gnd.n4013 gnd.n4012 0.152939
R19906 gnd.n4012 gnd.n4011 0.152939
R19907 gnd.n4011 gnd.n1996 0.152939
R19908 gnd.n4007 gnd.n1996 0.152939
R19909 gnd.n4007 gnd.n1907 0.152939
R19910 gnd.n4298 gnd.n1907 0.152939
R19911 gnd.n4298 gnd.n4297 0.152939
R19912 gnd.n5848 gnd.n1001 0.152939
R19913 gnd.n5844 gnd.n1001 0.152939
R19914 gnd.n5844 gnd.n5843 0.152939
R19915 gnd.n5843 gnd.n5842 0.152939
R19916 gnd.n5842 gnd.n1006 0.152939
R19917 gnd.n5838 gnd.n1006 0.152939
R19918 gnd.n5838 gnd.n5837 0.152939
R19919 gnd.n5837 gnd.n5836 0.152939
R19920 gnd.n5836 gnd.n1011 0.152939
R19921 gnd.n5832 gnd.n1011 0.152939
R19922 gnd.n5832 gnd.n5831 0.152939
R19923 gnd.n5831 gnd.n5830 0.152939
R19924 gnd.n5830 gnd.n1016 0.152939
R19925 gnd.n5826 gnd.n1016 0.152939
R19926 gnd.n5826 gnd.n5825 0.152939
R19927 gnd.n5825 gnd.n5824 0.152939
R19928 gnd.n5824 gnd.n1021 0.152939
R19929 gnd.n5820 gnd.n1021 0.152939
R19930 gnd.n5820 gnd.n5819 0.152939
R19931 gnd.n5819 gnd.n5818 0.152939
R19932 gnd.n5818 gnd.n1026 0.152939
R19933 gnd.n5814 gnd.n1026 0.152939
R19934 gnd.n5814 gnd.n5813 0.152939
R19935 gnd.n5813 gnd.n5812 0.152939
R19936 gnd.n5812 gnd.n1031 0.152939
R19937 gnd.n5808 gnd.n1031 0.152939
R19938 gnd.n5808 gnd.n5807 0.152939
R19939 gnd.n5807 gnd.n5806 0.152939
R19940 gnd.n5806 gnd.n1036 0.152939
R19941 gnd.n5802 gnd.n1036 0.152939
R19942 gnd.n5802 gnd.n5801 0.152939
R19943 gnd.n5801 gnd.n5800 0.152939
R19944 gnd.n5800 gnd.n1041 0.152939
R19945 gnd.n5796 gnd.n1041 0.152939
R19946 gnd.n5796 gnd.n5795 0.152939
R19947 gnd.n5795 gnd.n5794 0.152939
R19948 gnd.n5794 gnd.n1046 0.152939
R19949 gnd.n5790 gnd.n1046 0.152939
R19950 gnd.n5790 gnd.n5789 0.152939
R19951 gnd.n5789 gnd.n5788 0.152939
R19952 gnd.n5788 gnd.n1051 0.152939
R19953 gnd.n5784 gnd.n1051 0.152939
R19954 gnd.n5784 gnd.n5783 0.152939
R19955 gnd.n5783 gnd.n5782 0.152939
R19956 gnd.n5782 gnd.n1056 0.152939
R19957 gnd.n5778 gnd.n1056 0.152939
R19958 gnd.n5778 gnd.n5777 0.152939
R19959 gnd.n5777 gnd.n5776 0.152939
R19960 gnd.n5776 gnd.n1061 0.152939
R19961 gnd.n5772 gnd.n1061 0.152939
R19962 gnd.n5772 gnd.n5771 0.152939
R19963 gnd.n5771 gnd.n5770 0.152939
R19964 gnd.n5770 gnd.n1066 0.152939
R19965 gnd.n5766 gnd.n1066 0.152939
R19966 gnd.n5766 gnd.n5765 0.152939
R19967 gnd.n5765 gnd.n5764 0.152939
R19968 gnd.n5764 gnd.n1071 0.152939
R19969 gnd.n5760 gnd.n1071 0.152939
R19970 gnd.n5760 gnd.n5759 0.152939
R19971 gnd.n5759 gnd.n5758 0.152939
R19972 gnd.n5758 gnd.n1076 0.152939
R19973 gnd.n5754 gnd.n1076 0.152939
R19974 gnd.n5754 gnd.n5753 0.152939
R19975 gnd.n5753 gnd.n5752 0.152939
R19976 gnd.n5752 gnd.n1081 0.152939
R19977 gnd.n5748 gnd.n1081 0.152939
R19978 gnd.n5748 gnd.n5747 0.152939
R19979 gnd.n5747 gnd.n5746 0.152939
R19980 gnd.n5746 gnd.n1086 0.152939
R19981 gnd.n5742 gnd.n1086 0.152939
R19982 gnd.n5742 gnd.n5741 0.152939
R19983 gnd.n5741 gnd.n5740 0.152939
R19984 gnd.n5740 gnd.n1091 0.152939
R19985 gnd.n5736 gnd.n1091 0.152939
R19986 gnd.n5736 gnd.n5735 0.152939
R19987 gnd.n5735 gnd.n5734 0.152939
R19988 gnd.n5734 gnd.n1096 0.152939
R19989 gnd.n5730 gnd.n1096 0.152939
R19990 gnd.n5730 gnd.n5729 0.152939
R19991 gnd.n5729 gnd.n5728 0.152939
R19992 gnd.n5728 gnd.n1101 0.152939
R19993 gnd.n1104 gnd.n1101 0.152939
R19994 gnd.n5027 gnd.n1146 0.152939
R19995 gnd.n5698 gnd.n1146 0.152939
R19996 gnd.n5698 gnd.n5697 0.152939
R19997 gnd.n5697 gnd.n5696 0.152939
R19998 gnd.n5696 gnd.n1147 0.152939
R19999 gnd.n5692 gnd.n1147 0.152939
R20000 gnd.n5692 gnd.n5691 0.152939
R20001 gnd.n5691 gnd.n5690 0.152939
R20002 gnd.n5690 gnd.n1152 0.152939
R20003 gnd.n5686 gnd.n1152 0.152939
R20004 gnd.n5686 gnd.n5685 0.152939
R20005 gnd.n5685 gnd.n5684 0.152939
R20006 gnd.n5684 gnd.n1157 0.152939
R20007 gnd.n5680 gnd.n1157 0.152939
R20008 gnd.n5680 gnd.n5679 0.152939
R20009 gnd.n5679 gnd.n5678 0.152939
R20010 gnd.n5678 gnd.n1162 0.152939
R20011 gnd.n5674 gnd.n1162 0.152939
R20012 gnd.n5674 gnd.n5673 0.152939
R20013 gnd.n5673 gnd.n5672 0.152939
R20014 gnd.n5672 gnd.n1167 0.152939
R20015 gnd.n5668 gnd.n1167 0.152939
R20016 gnd.n5668 gnd.n228 0.152939
R20017 gnd.n6791 gnd.n228 0.152939
R20018 gnd.n6792 gnd.n6791 0.152939
R20019 gnd.n6793 gnd.n6792 0.152939
R20020 gnd.n6793 gnd.n206 0.152939
R20021 gnd.n6807 gnd.n206 0.152939
R20022 gnd.n6808 gnd.n6807 0.152939
R20023 gnd.n6809 gnd.n6808 0.152939
R20024 gnd.n6809 gnd.n191 0.152939
R20025 gnd.n6823 gnd.n191 0.152939
R20026 gnd.n6824 gnd.n6823 0.152939
R20027 gnd.n6825 gnd.n6824 0.152939
R20028 gnd.n6825 gnd.n174 0.152939
R20029 gnd.n6839 gnd.n174 0.152939
R20030 gnd.n6840 gnd.n6839 0.152939
R20031 gnd.n6915 gnd.n6840 0.152939
R20032 gnd.n6915 gnd.n6914 0.152939
R20033 gnd.n6914 gnd.n6913 0.152939
R20034 gnd.n6913 gnd.n6841 0.152939
R20035 gnd.n6909 gnd.n6841 0.152939
R20036 gnd.n6908 gnd.n6843 0.152939
R20037 gnd.n6904 gnd.n6843 0.152939
R20038 gnd.n6904 gnd.n6903 0.152939
R20039 gnd.n6903 gnd.n6902 0.152939
R20040 gnd.n6902 gnd.n6849 0.152939
R20041 gnd.n6898 gnd.n6849 0.152939
R20042 gnd.n6898 gnd.n6897 0.152939
R20043 gnd.n6897 gnd.n6896 0.152939
R20044 gnd.n6896 gnd.n6857 0.152939
R20045 gnd.n6892 gnd.n6857 0.152939
R20046 gnd.n6892 gnd.n6891 0.152939
R20047 gnd.n6891 gnd.n6890 0.152939
R20048 gnd.n6890 gnd.n6865 0.152939
R20049 gnd.n6886 gnd.n6865 0.152939
R20050 gnd.n6886 gnd.n6885 0.152939
R20051 gnd.n6885 gnd.n6884 0.152939
R20052 gnd.n6884 gnd.n6873 0.152939
R20053 gnd.n6873 gnd.n78 0.152939
R20054 gnd.n5471 gnd.n1264 0.152939
R20055 gnd.n5472 gnd.n5471 0.152939
R20056 gnd.n5474 gnd.n5472 0.152939
R20057 gnd.n5474 gnd.n5473 0.152939
R20058 gnd.n5473 gnd.n1246 0.152939
R20059 gnd.n5557 gnd.n1246 0.152939
R20060 gnd.n5558 gnd.n5557 0.152939
R20061 gnd.n5560 gnd.n5558 0.152939
R20062 gnd.n5560 gnd.n5559 0.152939
R20063 gnd.n5559 gnd.n1217 0.152939
R20064 gnd.n5589 gnd.n1217 0.152939
R20065 gnd.n5590 gnd.n5589 0.152939
R20066 gnd.n5592 gnd.n5590 0.152939
R20067 gnd.n5592 gnd.n5591 0.152939
R20068 gnd.n5591 gnd.n1191 0.152939
R20069 gnd.n5622 gnd.n1191 0.152939
R20070 gnd.n5623 gnd.n5622 0.152939
R20071 gnd.n5625 gnd.n5623 0.152939
R20072 gnd.n5625 gnd.n5624 0.152939
R20073 gnd.n5624 gnd.n51 0.152939
R20074 gnd.n7040 gnd.n51 0.152939
R20075 gnd.n7040 gnd.n7039 0.152939
R20076 gnd.n7039 gnd.n53 0.152939
R20077 gnd.n7035 gnd.n53 0.152939
R20078 gnd.n7035 gnd.n7034 0.152939
R20079 gnd.n7034 gnd.n7033 0.152939
R20080 gnd.n7033 gnd.n58 0.152939
R20081 gnd.n7029 gnd.n58 0.152939
R20082 gnd.n7029 gnd.n7028 0.152939
R20083 gnd.n7028 gnd.n7027 0.152939
R20084 gnd.n7027 gnd.n63 0.152939
R20085 gnd.n7023 gnd.n63 0.152939
R20086 gnd.n7023 gnd.n7022 0.152939
R20087 gnd.n7022 gnd.n7021 0.152939
R20088 gnd.n7021 gnd.n68 0.152939
R20089 gnd.n7017 gnd.n68 0.152939
R20090 gnd.n7017 gnd.n7016 0.152939
R20091 gnd.n7016 gnd.n7015 0.152939
R20092 gnd.n7015 gnd.n73 0.152939
R20093 gnd.n7011 gnd.n73 0.152939
R20094 gnd.n7011 gnd.n7010 0.152939
R20095 gnd.n7010 gnd.n7009 0.152939
R20096 gnd.n5115 gnd.n4980 0.151415
R20097 gnd.n4296 gnd.n1908 0.151415
R20098 gnd.n3925 gnd.n3924 0.145814
R20099 gnd.n3925 gnd.n2018 0.145814
R20100 gnd.n2372 gnd.n0 0.127478
R20101 gnd.n5647 gnd.n215 0.10111
R20102 gnd.n3867 gnd.n901 0.10111
R20103 gnd.n2952 gnd.n2951 0.0767195
R20104 gnd.n2951 gnd.n2950 0.0767195
R20105 gnd.n5850 gnd.n5849 0.063
R20106 gnd.n5028 gnd.n5025 0.063
R20107 gnd.n3962 gnd.n901 0.0523293
R20108 gnd.n5602 gnd.n215 0.0523293
R20109 gnd.n3519 gnd.n2146 0.0477147
R20110 gnd.n2715 gnd.n2603 0.0442063
R20111 gnd.n2716 gnd.n2715 0.0442063
R20112 gnd.n2717 gnd.n2716 0.0442063
R20113 gnd.n2717 gnd.n2592 0.0442063
R20114 gnd.n2731 gnd.n2592 0.0442063
R20115 gnd.n2732 gnd.n2731 0.0442063
R20116 gnd.n2733 gnd.n2732 0.0442063
R20117 gnd.n2733 gnd.n2579 0.0442063
R20118 gnd.n2777 gnd.n2579 0.0442063
R20119 gnd.n2778 gnd.n2777 0.0442063
R20120 gnd.n2780 gnd.n2513 0.0344674
R20121 gnd.n5116 gnd.n5114 0.0344674
R20122 gnd.n4295 gnd.n1909 0.0344674
R20123 gnd.n2800 gnd.n2799 0.0269946
R20124 gnd.n2802 gnd.n2801 0.0269946
R20125 gnd.n2508 gnd.n2506 0.0269946
R20126 gnd.n2812 gnd.n2810 0.0269946
R20127 gnd.n2811 gnd.n2487 0.0269946
R20128 gnd.n2831 gnd.n2830 0.0269946
R20129 gnd.n2833 gnd.n2832 0.0269946
R20130 gnd.n2482 gnd.n2481 0.0269946
R20131 gnd.n2843 gnd.n2477 0.0269946
R20132 gnd.n2842 gnd.n2479 0.0269946
R20133 gnd.n2478 gnd.n2460 0.0269946
R20134 gnd.n2863 gnd.n2461 0.0269946
R20135 gnd.n2862 gnd.n2462 0.0269946
R20136 gnd.n2896 gnd.n2437 0.0269946
R20137 gnd.n2898 gnd.n2897 0.0269946
R20138 gnd.n2899 gnd.n2384 0.0269946
R20139 gnd.n2432 gnd.n2385 0.0269946
R20140 gnd.n2434 gnd.n2386 0.0269946
R20141 gnd.n2909 gnd.n2908 0.0269946
R20142 gnd.n2911 gnd.n2910 0.0269946
R20143 gnd.n2912 gnd.n2406 0.0269946
R20144 gnd.n2914 gnd.n2407 0.0269946
R20145 gnd.n2917 gnd.n2408 0.0269946
R20146 gnd.n2920 gnd.n2919 0.0269946
R20147 gnd.n2922 gnd.n2921 0.0269946
R20148 gnd.n2987 gnd.n2319 0.0269946
R20149 gnd.n2989 gnd.n2988 0.0269946
R20150 gnd.n2998 gnd.n2312 0.0269946
R20151 gnd.n3000 gnd.n2999 0.0269946
R20152 gnd.n3001 gnd.n2310 0.0269946
R20153 gnd.n3008 gnd.n3004 0.0269946
R20154 gnd.n3007 gnd.n3006 0.0269946
R20155 gnd.n3005 gnd.n2289 0.0269946
R20156 gnd.n3030 gnd.n2290 0.0269946
R20157 gnd.n3029 gnd.n2291 0.0269946
R20158 gnd.n3072 gnd.n2264 0.0269946
R20159 gnd.n3074 gnd.n3073 0.0269946
R20160 gnd.n3084 gnd.n2257 0.0269946
R20161 gnd.n3086 gnd.n3085 0.0269946
R20162 gnd.n3087 gnd.n2255 0.0269946
R20163 gnd.n3094 gnd.n3090 0.0269946
R20164 gnd.n3093 gnd.n3092 0.0269946
R20165 gnd.n3091 gnd.n2234 0.0269946
R20166 gnd.n3116 gnd.n2235 0.0269946
R20167 gnd.n3115 gnd.n2236 0.0269946
R20168 gnd.n3162 gnd.n2210 0.0269946
R20169 gnd.n3164 gnd.n3163 0.0269946
R20170 gnd.n3173 gnd.n2203 0.0269946
R20171 gnd.n3432 gnd.n2201 0.0269946
R20172 gnd.n3437 gnd.n3435 0.0269946
R20173 gnd.n3436 gnd.n2182 0.0269946
R20174 gnd.n3461 gnd.n3460 0.0269946
R20175 gnd.n5025 gnd.n5024 0.0246168
R20176 gnd.n5849 gnd.n1000 0.0246168
R20177 gnd.n2780 gnd.n2779 0.0202011
R20178 gnd.n5024 gnd.n5022 0.0174837
R20179 gnd.n5036 gnd.n5022 0.0174837
R20180 gnd.n5038 gnd.n5036 0.0174837
R20181 gnd.n5038 gnd.n5037 0.0174837
R20182 gnd.n5037 gnd.n5017 0.0174837
R20183 gnd.n5047 gnd.n5017 0.0174837
R20184 gnd.n5047 gnd.n5046 0.0174837
R20185 gnd.n5046 gnd.n5018 0.0174837
R20186 gnd.n5018 gnd.n5013 0.0174837
R20187 gnd.n5055 gnd.n5013 0.0174837
R20188 gnd.n5057 gnd.n5055 0.0174837
R20189 gnd.n5057 gnd.n5056 0.0174837
R20190 gnd.n5056 gnd.n5008 0.0174837
R20191 gnd.n5066 gnd.n5008 0.0174837
R20192 gnd.n5066 gnd.n5065 0.0174837
R20193 gnd.n5065 gnd.n5009 0.0174837
R20194 gnd.n5009 gnd.n5004 0.0174837
R20195 gnd.n5074 gnd.n5004 0.0174837
R20196 gnd.n5076 gnd.n5074 0.0174837
R20197 gnd.n5076 gnd.n5075 0.0174837
R20198 gnd.n5075 gnd.n4999 0.0174837
R20199 gnd.n5085 gnd.n4999 0.0174837
R20200 gnd.n5085 gnd.n5084 0.0174837
R20201 gnd.n5084 gnd.n5000 0.0174837
R20202 gnd.n5000 gnd.n4995 0.0174837
R20203 gnd.n5093 gnd.n4995 0.0174837
R20204 gnd.n5095 gnd.n5093 0.0174837
R20205 gnd.n5095 gnd.n5094 0.0174837
R20206 gnd.n5094 gnd.n4990 0.0174837
R20207 gnd.n5106 gnd.n4990 0.0174837
R20208 gnd.n5106 gnd.n5105 0.0174837
R20209 gnd.n5105 gnd.n4991 0.0174837
R20210 gnd.n4991 gnd.n4984 0.0174837
R20211 gnd.n5113 gnd.n4984 0.0174837
R20212 gnd.n5114 gnd.n5113 0.0174837
R20213 gnd.n4074 gnd.n1000 0.0174837
R20214 gnd.n4076 gnd.n4074 0.0174837
R20215 gnd.n4184 gnd.n4076 0.0174837
R20216 gnd.n4184 gnd.n4183 0.0174837
R20217 gnd.n4183 gnd.n4077 0.0174837
R20218 gnd.n4180 gnd.n4077 0.0174837
R20219 gnd.n4180 gnd.n4179 0.0174837
R20220 gnd.n4179 gnd.n4087 0.0174837
R20221 gnd.n4176 gnd.n4087 0.0174837
R20222 gnd.n4176 gnd.n4175 0.0174837
R20223 gnd.n4175 gnd.n4092 0.0174837
R20224 gnd.n4172 gnd.n4092 0.0174837
R20225 gnd.n4172 gnd.n4171 0.0174837
R20226 gnd.n4171 gnd.n4098 0.0174837
R20227 gnd.n4168 gnd.n4098 0.0174837
R20228 gnd.n4168 gnd.n4167 0.0174837
R20229 gnd.n4167 gnd.n4102 0.0174837
R20230 gnd.n4164 gnd.n4102 0.0174837
R20231 gnd.n4164 gnd.n4163 0.0174837
R20232 gnd.n4163 gnd.n4109 0.0174837
R20233 gnd.n4160 gnd.n4109 0.0174837
R20234 gnd.n4160 gnd.n4159 0.0174837
R20235 gnd.n4159 gnd.n4115 0.0174837
R20236 gnd.n4156 gnd.n4115 0.0174837
R20237 gnd.n4156 gnd.n4155 0.0174837
R20238 gnd.n4155 gnd.n4121 0.0174837
R20239 gnd.n4152 gnd.n4121 0.0174837
R20240 gnd.n4152 gnd.n4151 0.0174837
R20241 gnd.n4151 gnd.n4125 0.0174837
R20242 gnd.n4148 gnd.n4125 0.0174837
R20243 gnd.n4148 gnd.n4147 0.0174837
R20244 gnd.n4147 gnd.n4134 0.0174837
R20245 gnd.n4144 gnd.n4134 0.0174837
R20246 gnd.n4144 gnd.n4143 0.0174837
R20247 gnd.n4143 gnd.n1909 0.0174837
R20248 gnd.n2779 gnd.n2778 0.0148637
R20249 gnd.n3430 gnd.n3174 0.0144266
R20250 gnd.n3431 gnd.n3430 0.0130679
R20251 gnd.n2799 gnd.n2513 0.00797283
R20252 gnd.n2801 gnd.n2800 0.00797283
R20253 gnd.n2802 gnd.n2508 0.00797283
R20254 gnd.n2810 gnd.n2506 0.00797283
R20255 gnd.n2812 gnd.n2811 0.00797283
R20256 gnd.n2830 gnd.n2487 0.00797283
R20257 gnd.n2832 gnd.n2831 0.00797283
R20258 gnd.n2833 gnd.n2482 0.00797283
R20259 gnd.n2481 gnd.n2477 0.00797283
R20260 gnd.n2843 gnd.n2842 0.00797283
R20261 gnd.n2479 gnd.n2478 0.00797283
R20262 gnd.n2461 gnd.n2460 0.00797283
R20263 gnd.n2863 gnd.n2862 0.00797283
R20264 gnd.n2462 gnd.n2437 0.00797283
R20265 gnd.n2897 gnd.n2896 0.00797283
R20266 gnd.n2899 gnd.n2898 0.00797283
R20267 gnd.n2432 gnd.n2384 0.00797283
R20268 gnd.n2434 gnd.n2385 0.00797283
R20269 gnd.n2908 gnd.n2386 0.00797283
R20270 gnd.n2910 gnd.n2909 0.00797283
R20271 gnd.n2912 gnd.n2911 0.00797283
R20272 gnd.n2914 gnd.n2406 0.00797283
R20273 gnd.n2917 gnd.n2407 0.00797283
R20274 gnd.n2919 gnd.n2408 0.00797283
R20275 gnd.n2922 gnd.n2920 0.00797283
R20276 gnd.n2921 gnd.n2319 0.00797283
R20277 gnd.n2989 gnd.n2987 0.00797283
R20278 gnd.n2988 gnd.n2312 0.00797283
R20279 gnd.n2999 gnd.n2998 0.00797283
R20280 gnd.n3001 gnd.n3000 0.00797283
R20281 gnd.n3004 gnd.n2310 0.00797283
R20282 gnd.n3008 gnd.n3007 0.00797283
R20283 gnd.n3006 gnd.n3005 0.00797283
R20284 gnd.n2290 gnd.n2289 0.00797283
R20285 gnd.n3030 gnd.n3029 0.00797283
R20286 gnd.n2291 gnd.n2264 0.00797283
R20287 gnd.n3074 gnd.n3072 0.00797283
R20288 gnd.n3073 gnd.n2257 0.00797283
R20289 gnd.n3085 gnd.n3084 0.00797283
R20290 gnd.n3087 gnd.n3086 0.00797283
R20291 gnd.n3090 gnd.n2255 0.00797283
R20292 gnd.n3094 gnd.n3093 0.00797283
R20293 gnd.n3092 gnd.n3091 0.00797283
R20294 gnd.n2235 gnd.n2234 0.00797283
R20295 gnd.n3116 gnd.n3115 0.00797283
R20296 gnd.n2236 gnd.n2210 0.00797283
R20297 gnd.n3164 gnd.n3162 0.00797283
R20298 gnd.n3163 gnd.n2203 0.00797283
R20299 gnd.n3174 gnd.n3173 0.00797283
R20300 gnd.n3432 gnd.n3431 0.00797283
R20301 gnd.n3435 gnd.n2201 0.00797283
R20302 gnd.n3437 gnd.n3436 0.00797283
R20303 gnd.n3460 gnd.n2182 0.00797283
R20304 gnd.n3461 gnd.n2146 0.00797283
R20305 gnd.n5499 gnd.n1167 0.00614909
R20306 gnd.n3932 gnd.n3931 0.00614909
R20307 gnd.n5116 gnd.n5115 0.000839674
R20308 gnd.n4296 gnd.n4295 0.000839674
R20309 commonsourceibias.n25 commonsourceibias.t46 230.006
R20310 commonsourceibias.n91 commonsourceibias.t62 230.006
R20311 commonsourceibias.n154 commonsourceibias.t54 230.006
R20312 commonsourceibias.n258 commonsourceibias.t16 230.006
R20313 commonsourceibias.n217 commonsourceibias.t75 230.006
R20314 commonsourceibias.n355 commonsourceibias.t65 230.006
R20315 commonsourceibias.n70 commonsourceibias.t32 207.983
R20316 commonsourceibias.n136 commonsourceibias.t71 207.983
R20317 commonsourceibias.n199 commonsourceibias.t61 207.983
R20318 commonsourceibias.n304 commonsourceibias.t2 207.983
R20319 commonsourceibias.n338 commonsourceibias.t84 207.983
R20320 commonsourceibias.n401 commonsourceibias.t73 207.983
R20321 commonsourceibias.n10 commonsourceibias.t14 168.701
R20322 commonsourceibias.n63 commonsourceibias.t24 168.701
R20323 commonsourceibias.n57 commonsourceibias.t30 168.701
R20324 commonsourceibias.n16 commonsourceibias.t20 168.701
R20325 commonsourceibias.n49 commonsourceibias.t36 168.701
R20326 commonsourceibias.n43 commonsourceibias.t44 168.701
R20327 commonsourceibias.n19 commonsourceibias.t26 168.701
R20328 commonsourceibias.n21 commonsourceibias.t34 168.701
R20329 commonsourceibias.n23 commonsourceibias.t10 168.701
R20330 commonsourceibias.n26 commonsourceibias.t40 168.701
R20331 commonsourceibias.n1 commonsourceibias.t81 168.701
R20332 commonsourceibias.n129 commonsourceibias.t55 168.701
R20333 commonsourceibias.n123 commonsourceibias.t53 168.701
R20334 commonsourceibias.n7 commonsourceibias.t76 168.701
R20335 commonsourceibias.n115 commonsourceibias.t86 168.701
R20336 commonsourceibias.n109 commonsourceibias.t50 168.701
R20337 commonsourceibias.n85 commonsourceibias.t69 168.701
R20338 commonsourceibias.n87 commonsourceibias.t67 168.701
R20339 commonsourceibias.n89 commonsourceibias.t78 168.701
R20340 commonsourceibias.n92 commonsourceibias.t64 168.701
R20341 commonsourceibias.n155 commonsourceibias.t57 168.701
R20342 commonsourceibias.n152 commonsourceibias.t68 168.701
R20343 commonsourceibias.n150 commonsourceibias.t58 168.701
R20344 commonsourceibias.n148 commonsourceibias.t60 168.701
R20345 commonsourceibias.n172 commonsourceibias.t91 168.701
R20346 commonsourceibias.n178 commonsourceibias.t77 168.701
R20347 commonsourceibias.n145 commonsourceibias.t66 168.701
R20348 commonsourceibias.n186 commonsourceibias.t95 168.701
R20349 commonsourceibias.n192 commonsourceibias.t49 168.701
R20350 commonsourceibias.n139 commonsourceibias.t72 168.701
R20351 commonsourceibias.n259 commonsourceibias.t8 168.701
R20352 commonsourceibias.n256 commonsourceibias.t18 168.701
R20353 commonsourceibias.n254 commonsourceibias.t4 168.701
R20354 commonsourceibias.n252 commonsourceibias.t42 168.701
R20355 commonsourceibias.n276 commonsourceibias.t12 168.701
R20356 commonsourceibias.n282 commonsourceibias.t6 168.701
R20357 commonsourceibias.n284 commonsourceibias.t28 168.701
R20358 commonsourceibias.n291 commonsourceibias.t0 168.701
R20359 commonsourceibias.n297 commonsourceibias.t38 168.701
R20360 commonsourceibias.n244 commonsourceibias.t22 168.701
R20361 commonsourceibias.n203 commonsourceibias.t92 168.701
R20362 commonsourceibias.n331 commonsourceibias.t51 168.701
R20363 commonsourceibias.n325 commonsourceibias.t63 168.701
R20364 commonsourceibias.n318 commonsourceibias.t88 168.701
R20365 commonsourceibias.n316 commonsourceibias.t48 168.701
R20366 commonsourceibias.n218 commonsourceibias.t59 168.701
R20367 commonsourceibias.n215 commonsourceibias.t90 168.701
R20368 commonsourceibias.n213 commonsourceibias.t80 168.701
R20369 commonsourceibias.n211 commonsourceibias.t83 168.701
R20370 commonsourceibias.n235 commonsourceibias.t94 168.701
R20371 commonsourceibias.n356 commonsourceibias.t52 168.701
R20372 commonsourceibias.n353 commonsourceibias.t82 168.701
R20373 commonsourceibias.n351 commonsourceibias.t70 168.701
R20374 commonsourceibias.n349 commonsourceibias.t74 168.701
R20375 commonsourceibias.n373 commonsourceibias.t87 168.701
R20376 commonsourceibias.n379 commonsourceibias.t89 168.701
R20377 commonsourceibias.n381 commonsourceibias.t79 168.701
R20378 commonsourceibias.n388 commonsourceibias.t56 168.701
R20379 commonsourceibias.n394 commonsourceibias.t93 168.701
R20380 commonsourceibias.n341 commonsourceibias.t85 168.701
R20381 commonsourceibias.n27 commonsourceibias.n24 161.3
R20382 commonsourceibias.n29 commonsourceibias.n28 161.3
R20383 commonsourceibias.n31 commonsourceibias.n30 161.3
R20384 commonsourceibias.n32 commonsourceibias.n22 161.3
R20385 commonsourceibias.n34 commonsourceibias.n33 161.3
R20386 commonsourceibias.n36 commonsourceibias.n35 161.3
R20387 commonsourceibias.n37 commonsourceibias.n20 161.3
R20388 commonsourceibias.n39 commonsourceibias.n38 161.3
R20389 commonsourceibias.n41 commonsourceibias.n40 161.3
R20390 commonsourceibias.n42 commonsourceibias.n18 161.3
R20391 commonsourceibias.n45 commonsourceibias.n44 161.3
R20392 commonsourceibias.n46 commonsourceibias.n17 161.3
R20393 commonsourceibias.n48 commonsourceibias.n47 161.3
R20394 commonsourceibias.n50 commonsourceibias.n15 161.3
R20395 commonsourceibias.n52 commonsourceibias.n51 161.3
R20396 commonsourceibias.n53 commonsourceibias.n14 161.3
R20397 commonsourceibias.n55 commonsourceibias.n54 161.3
R20398 commonsourceibias.n56 commonsourceibias.n13 161.3
R20399 commonsourceibias.n59 commonsourceibias.n58 161.3
R20400 commonsourceibias.n60 commonsourceibias.n12 161.3
R20401 commonsourceibias.n62 commonsourceibias.n61 161.3
R20402 commonsourceibias.n64 commonsourceibias.n11 161.3
R20403 commonsourceibias.n66 commonsourceibias.n65 161.3
R20404 commonsourceibias.n68 commonsourceibias.n67 161.3
R20405 commonsourceibias.n69 commonsourceibias.n9 161.3
R20406 commonsourceibias.n93 commonsourceibias.n90 161.3
R20407 commonsourceibias.n95 commonsourceibias.n94 161.3
R20408 commonsourceibias.n97 commonsourceibias.n96 161.3
R20409 commonsourceibias.n98 commonsourceibias.n88 161.3
R20410 commonsourceibias.n100 commonsourceibias.n99 161.3
R20411 commonsourceibias.n102 commonsourceibias.n101 161.3
R20412 commonsourceibias.n103 commonsourceibias.n86 161.3
R20413 commonsourceibias.n105 commonsourceibias.n104 161.3
R20414 commonsourceibias.n107 commonsourceibias.n106 161.3
R20415 commonsourceibias.n108 commonsourceibias.n84 161.3
R20416 commonsourceibias.n111 commonsourceibias.n110 161.3
R20417 commonsourceibias.n112 commonsourceibias.n8 161.3
R20418 commonsourceibias.n114 commonsourceibias.n113 161.3
R20419 commonsourceibias.n116 commonsourceibias.n6 161.3
R20420 commonsourceibias.n118 commonsourceibias.n117 161.3
R20421 commonsourceibias.n119 commonsourceibias.n5 161.3
R20422 commonsourceibias.n121 commonsourceibias.n120 161.3
R20423 commonsourceibias.n122 commonsourceibias.n4 161.3
R20424 commonsourceibias.n125 commonsourceibias.n124 161.3
R20425 commonsourceibias.n126 commonsourceibias.n3 161.3
R20426 commonsourceibias.n128 commonsourceibias.n127 161.3
R20427 commonsourceibias.n130 commonsourceibias.n2 161.3
R20428 commonsourceibias.n132 commonsourceibias.n131 161.3
R20429 commonsourceibias.n134 commonsourceibias.n133 161.3
R20430 commonsourceibias.n135 commonsourceibias.n0 161.3
R20431 commonsourceibias.n198 commonsourceibias.n138 161.3
R20432 commonsourceibias.n197 commonsourceibias.n196 161.3
R20433 commonsourceibias.n195 commonsourceibias.n194 161.3
R20434 commonsourceibias.n193 commonsourceibias.n140 161.3
R20435 commonsourceibias.n191 commonsourceibias.n190 161.3
R20436 commonsourceibias.n189 commonsourceibias.n141 161.3
R20437 commonsourceibias.n188 commonsourceibias.n187 161.3
R20438 commonsourceibias.n185 commonsourceibias.n142 161.3
R20439 commonsourceibias.n184 commonsourceibias.n183 161.3
R20440 commonsourceibias.n182 commonsourceibias.n143 161.3
R20441 commonsourceibias.n181 commonsourceibias.n180 161.3
R20442 commonsourceibias.n179 commonsourceibias.n144 161.3
R20443 commonsourceibias.n177 commonsourceibias.n176 161.3
R20444 commonsourceibias.n175 commonsourceibias.n146 161.3
R20445 commonsourceibias.n174 commonsourceibias.n173 161.3
R20446 commonsourceibias.n171 commonsourceibias.n147 161.3
R20447 commonsourceibias.n170 commonsourceibias.n169 161.3
R20448 commonsourceibias.n168 commonsourceibias.n167 161.3
R20449 commonsourceibias.n166 commonsourceibias.n149 161.3
R20450 commonsourceibias.n165 commonsourceibias.n164 161.3
R20451 commonsourceibias.n163 commonsourceibias.n162 161.3
R20452 commonsourceibias.n161 commonsourceibias.n151 161.3
R20453 commonsourceibias.n160 commonsourceibias.n159 161.3
R20454 commonsourceibias.n158 commonsourceibias.n157 161.3
R20455 commonsourceibias.n156 commonsourceibias.n153 161.3
R20456 commonsourceibias.n303 commonsourceibias.n243 161.3
R20457 commonsourceibias.n302 commonsourceibias.n301 161.3
R20458 commonsourceibias.n300 commonsourceibias.n299 161.3
R20459 commonsourceibias.n298 commonsourceibias.n245 161.3
R20460 commonsourceibias.n296 commonsourceibias.n295 161.3
R20461 commonsourceibias.n294 commonsourceibias.n246 161.3
R20462 commonsourceibias.n293 commonsourceibias.n292 161.3
R20463 commonsourceibias.n290 commonsourceibias.n247 161.3
R20464 commonsourceibias.n289 commonsourceibias.n288 161.3
R20465 commonsourceibias.n287 commonsourceibias.n248 161.3
R20466 commonsourceibias.n286 commonsourceibias.n285 161.3
R20467 commonsourceibias.n283 commonsourceibias.n249 161.3
R20468 commonsourceibias.n281 commonsourceibias.n280 161.3
R20469 commonsourceibias.n279 commonsourceibias.n250 161.3
R20470 commonsourceibias.n278 commonsourceibias.n277 161.3
R20471 commonsourceibias.n275 commonsourceibias.n251 161.3
R20472 commonsourceibias.n274 commonsourceibias.n273 161.3
R20473 commonsourceibias.n272 commonsourceibias.n271 161.3
R20474 commonsourceibias.n270 commonsourceibias.n253 161.3
R20475 commonsourceibias.n269 commonsourceibias.n268 161.3
R20476 commonsourceibias.n267 commonsourceibias.n266 161.3
R20477 commonsourceibias.n265 commonsourceibias.n255 161.3
R20478 commonsourceibias.n264 commonsourceibias.n263 161.3
R20479 commonsourceibias.n262 commonsourceibias.n261 161.3
R20480 commonsourceibias.n260 commonsourceibias.n257 161.3
R20481 commonsourceibias.n237 commonsourceibias.n236 161.3
R20482 commonsourceibias.n234 commonsourceibias.n210 161.3
R20483 commonsourceibias.n233 commonsourceibias.n232 161.3
R20484 commonsourceibias.n231 commonsourceibias.n230 161.3
R20485 commonsourceibias.n229 commonsourceibias.n212 161.3
R20486 commonsourceibias.n228 commonsourceibias.n227 161.3
R20487 commonsourceibias.n226 commonsourceibias.n225 161.3
R20488 commonsourceibias.n224 commonsourceibias.n214 161.3
R20489 commonsourceibias.n223 commonsourceibias.n222 161.3
R20490 commonsourceibias.n221 commonsourceibias.n220 161.3
R20491 commonsourceibias.n219 commonsourceibias.n216 161.3
R20492 commonsourceibias.n313 commonsourceibias.n209 161.3
R20493 commonsourceibias.n337 commonsourceibias.n202 161.3
R20494 commonsourceibias.n336 commonsourceibias.n335 161.3
R20495 commonsourceibias.n334 commonsourceibias.n333 161.3
R20496 commonsourceibias.n332 commonsourceibias.n204 161.3
R20497 commonsourceibias.n330 commonsourceibias.n329 161.3
R20498 commonsourceibias.n328 commonsourceibias.n205 161.3
R20499 commonsourceibias.n327 commonsourceibias.n326 161.3
R20500 commonsourceibias.n324 commonsourceibias.n206 161.3
R20501 commonsourceibias.n323 commonsourceibias.n322 161.3
R20502 commonsourceibias.n321 commonsourceibias.n207 161.3
R20503 commonsourceibias.n320 commonsourceibias.n319 161.3
R20504 commonsourceibias.n317 commonsourceibias.n208 161.3
R20505 commonsourceibias.n315 commonsourceibias.n314 161.3
R20506 commonsourceibias.n400 commonsourceibias.n340 161.3
R20507 commonsourceibias.n399 commonsourceibias.n398 161.3
R20508 commonsourceibias.n397 commonsourceibias.n396 161.3
R20509 commonsourceibias.n395 commonsourceibias.n342 161.3
R20510 commonsourceibias.n393 commonsourceibias.n392 161.3
R20511 commonsourceibias.n391 commonsourceibias.n343 161.3
R20512 commonsourceibias.n390 commonsourceibias.n389 161.3
R20513 commonsourceibias.n387 commonsourceibias.n344 161.3
R20514 commonsourceibias.n386 commonsourceibias.n385 161.3
R20515 commonsourceibias.n384 commonsourceibias.n345 161.3
R20516 commonsourceibias.n383 commonsourceibias.n382 161.3
R20517 commonsourceibias.n380 commonsourceibias.n346 161.3
R20518 commonsourceibias.n378 commonsourceibias.n377 161.3
R20519 commonsourceibias.n376 commonsourceibias.n347 161.3
R20520 commonsourceibias.n375 commonsourceibias.n374 161.3
R20521 commonsourceibias.n372 commonsourceibias.n348 161.3
R20522 commonsourceibias.n371 commonsourceibias.n370 161.3
R20523 commonsourceibias.n369 commonsourceibias.n368 161.3
R20524 commonsourceibias.n367 commonsourceibias.n350 161.3
R20525 commonsourceibias.n366 commonsourceibias.n365 161.3
R20526 commonsourceibias.n364 commonsourceibias.n363 161.3
R20527 commonsourceibias.n362 commonsourceibias.n352 161.3
R20528 commonsourceibias.n361 commonsourceibias.n360 161.3
R20529 commonsourceibias.n359 commonsourceibias.n358 161.3
R20530 commonsourceibias.n357 commonsourceibias.n354 161.3
R20531 commonsourceibias.n80 commonsourceibias.n78 81.5057
R20532 commonsourceibias.n240 commonsourceibias.n238 81.5057
R20533 commonsourceibias.n80 commonsourceibias.n79 80.9324
R20534 commonsourceibias.n82 commonsourceibias.n81 80.9324
R20535 commonsourceibias.n77 commonsourceibias.n76 80.9324
R20536 commonsourceibias.n75 commonsourceibias.n74 80.9324
R20537 commonsourceibias.n73 commonsourceibias.n72 80.9324
R20538 commonsourceibias.n307 commonsourceibias.n306 80.9324
R20539 commonsourceibias.n309 commonsourceibias.n308 80.9324
R20540 commonsourceibias.n311 commonsourceibias.n310 80.9324
R20541 commonsourceibias.n242 commonsourceibias.n241 80.9324
R20542 commonsourceibias.n240 commonsourceibias.n239 80.9324
R20543 commonsourceibias.n71 commonsourceibias.n70 80.6037
R20544 commonsourceibias.n137 commonsourceibias.n136 80.6037
R20545 commonsourceibias.n200 commonsourceibias.n199 80.6037
R20546 commonsourceibias.n305 commonsourceibias.n304 80.6037
R20547 commonsourceibias.n339 commonsourceibias.n338 80.6037
R20548 commonsourceibias.n402 commonsourceibias.n401 80.6037
R20549 commonsourceibias.n65 commonsourceibias.n64 56.5617
R20550 commonsourceibias.n51 commonsourceibias.n50 56.5617
R20551 commonsourceibias.n42 commonsourceibias.n41 56.5617
R20552 commonsourceibias.n28 commonsourceibias.n27 56.5617
R20553 commonsourceibias.n131 commonsourceibias.n130 56.5617
R20554 commonsourceibias.n117 commonsourceibias.n116 56.5617
R20555 commonsourceibias.n108 commonsourceibias.n107 56.5617
R20556 commonsourceibias.n94 commonsourceibias.n93 56.5617
R20557 commonsourceibias.n157 commonsourceibias.n156 56.5617
R20558 commonsourceibias.n171 commonsourceibias.n170 56.5617
R20559 commonsourceibias.n180 commonsourceibias.n179 56.5617
R20560 commonsourceibias.n194 commonsourceibias.n193 56.5617
R20561 commonsourceibias.n261 commonsourceibias.n260 56.5617
R20562 commonsourceibias.n275 commonsourceibias.n274 56.5617
R20563 commonsourceibias.n285 commonsourceibias.n283 56.5617
R20564 commonsourceibias.n299 commonsourceibias.n298 56.5617
R20565 commonsourceibias.n333 commonsourceibias.n332 56.5617
R20566 commonsourceibias.n319 commonsourceibias.n317 56.5617
R20567 commonsourceibias.n220 commonsourceibias.n219 56.5617
R20568 commonsourceibias.n234 commonsourceibias.n233 56.5617
R20569 commonsourceibias.n358 commonsourceibias.n357 56.5617
R20570 commonsourceibias.n372 commonsourceibias.n371 56.5617
R20571 commonsourceibias.n382 commonsourceibias.n380 56.5617
R20572 commonsourceibias.n396 commonsourceibias.n395 56.5617
R20573 commonsourceibias.n56 commonsourceibias.n55 56.0773
R20574 commonsourceibias.n37 commonsourceibias.n36 56.0773
R20575 commonsourceibias.n122 commonsourceibias.n121 56.0773
R20576 commonsourceibias.n103 commonsourceibias.n102 56.0773
R20577 commonsourceibias.n166 commonsourceibias.n165 56.0773
R20578 commonsourceibias.n185 commonsourceibias.n184 56.0773
R20579 commonsourceibias.n270 commonsourceibias.n269 56.0773
R20580 commonsourceibias.n290 commonsourceibias.n289 56.0773
R20581 commonsourceibias.n324 commonsourceibias.n323 56.0773
R20582 commonsourceibias.n229 commonsourceibias.n228 56.0773
R20583 commonsourceibias.n367 commonsourceibias.n366 56.0773
R20584 commonsourceibias.n387 commonsourceibias.n386 56.0773
R20585 commonsourceibias.n70 commonsourceibias.n69 46.0096
R20586 commonsourceibias.n136 commonsourceibias.n135 46.0096
R20587 commonsourceibias.n199 commonsourceibias.n198 46.0096
R20588 commonsourceibias.n304 commonsourceibias.n303 46.0096
R20589 commonsourceibias.n338 commonsourceibias.n337 46.0096
R20590 commonsourceibias.n401 commonsourceibias.n400 46.0096
R20591 commonsourceibias.n58 commonsourceibias.n12 41.5458
R20592 commonsourceibias.n33 commonsourceibias.n32 41.5458
R20593 commonsourceibias.n124 commonsourceibias.n3 41.5458
R20594 commonsourceibias.n99 commonsourceibias.n98 41.5458
R20595 commonsourceibias.n162 commonsourceibias.n161 41.5458
R20596 commonsourceibias.n187 commonsourceibias.n141 41.5458
R20597 commonsourceibias.n266 commonsourceibias.n265 41.5458
R20598 commonsourceibias.n292 commonsourceibias.n246 41.5458
R20599 commonsourceibias.n326 commonsourceibias.n205 41.5458
R20600 commonsourceibias.n225 commonsourceibias.n224 41.5458
R20601 commonsourceibias.n363 commonsourceibias.n362 41.5458
R20602 commonsourceibias.n389 commonsourceibias.n343 41.5458
R20603 commonsourceibias.n48 commonsourceibias.n17 40.577
R20604 commonsourceibias.n44 commonsourceibias.n17 40.577
R20605 commonsourceibias.n114 commonsourceibias.n8 40.577
R20606 commonsourceibias.n110 commonsourceibias.n8 40.577
R20607 commonsourceibias.n173 commonsourceibias.n146 40.577
R20608 commonsourceibias.n177 commonsourceibias.n146 40.577
R20609 commonsourceibias.n277 commonsourceibias.n250 40.577
R20610 commonsourceibias.n281 commonsourceibias.n250 40.577
R20611 commonsourceibias.n315 commonsourceibias.n209 40.577
R20612 commonsourceibias.n236 commonsourceibias.n209 40.577
R20613 commonsourceibias.n374 commonsourceibias.n347 40.577
R20614 commonsourceibias.n378 commonsourceibias.n347 40.577
R20615 commonsourceibias.n62 commonsourceibias.n12 39.6083
R20616 commonsourceibias.n32 commonsourceibias.n31 39.6083
R20617 commonsourceibias.n128 commonsourceibias.n3 39.6083
R20618 commonsourceibias.n98 commonsourceibias.n97 39.6083
R20619 commonsourceibias.n161 commonsourceibias.n160 39.6083
R20620 commonsourceibias.n191 commonsourceibias.n141 39.6083
R20621 commonsourceibias.n265 commonsourceibias.n264 39.6083
R20622 commonsourceibias.n296 commonsourceibias.n246 39.6083
R20623 commonsourceibias.n330 commonsourceibias.n205 39.6083
R20624 commonsourceibias.n224 commonsourceibias.n223 39.6083
R20625 commonsourceibias.n362 commonsourceibias.n361 39.6083
R20626 commonsourceibias.n393 commonsourceibias.n343 39.6083
R20627 commonsourceibias.n26 commonsourceibias.n25 33.0515
R20628 commonsourceibias.n92 commonsourceibias.n91 33.0515
R20629 commonsourceibias.n155 commonsourceibias.n154 33.0515
R20630 commonsourceibias.n259 commonsourceibias.n258 33.0515
R20631 commonsourceibias.n218 commonsourceibias.n217 33.0515
R20632 commonsourceibias.n356 commonsourceibias.n355 33.0515
R20633 commonsourceibias.n25 commonsourceibias.n24 28.5514
R20634 commonsourceibias.n91 commonsourceibias.n90 28.5514
R20635 commonsourceibias.n154 commonsourceibias.n153 28.5514
R20636 commonsourceibias.n258 commonsourceibias.n257 28.5514
R20637 commonsourceibias.n217 commonsourceibias.n216 28.5514
R20638 commonsourceibias.n355 commonsourceibias.n354 28.5514
R20639 commonsourceibias.n69 commonsourceibias.n68 26.0455
R20640 commonsourceibias.n135 commonsourceibias.n134 26.0455
R20641 commonsourceibias.n198 commonsourceibias.n197 26.0455
R20642 commonsourceibias.n303 commonsourceibias.n302 26.0455
R20643 commonsourceibias.n337 commonsourceibias.n336 26.0455
R20644 commonsourceibias.n400 commonsourceibias.n399 26.0455
R20645 commonsourceibias.n55 commonsourceibias.n14 25.0767
R20646 commonsourceibias.n38 commonsourceibias.n37 25.0767
R20647 commonsourceibias.n121 commonsourceibias.n5 25.0767
R20648 commonsourceibias.n104 commonsourceibias.n103 25.0767
R20649 commonsourceibias.n167 commonsourceibias.n166 25.0767
R20650 commonsourceibias.n184 commonsourceibias.n143 25.0767
R20651 commonsourceibias.n271 commonsourceibias.n270 25.0767
R20652 commonsourceibias.n289 commonsourceibias.n248 25.0767
R20653 commonsourceibias.n323 commonsourceibias.n207 25.0767
R20654 commonsourceibias.n230 commonsourceibias.n229 25.0767
R20655 commonsourceibias.n368 commonsourceibias.n367 25.0767
R20656 commonsourceibias.n386 commonsourceibias.n345 25.0767
R20657 commonsourceibias.n51 commonsourceibias.n16 24.3464
R20658 commonsourceibias.n41 commonsourceibias.n19 24.3464
R20659 commonsourceibias.n117 commonsourceibias.n7 24.3464
R20660 commonsourceibias.n107 commonsourceibias.n85 24.3464
R20661 commonsourceibias.n170 commonsourceibias.n148 24.3464
R20662 commonsourceibias.n180 commonsourceibias.n145 24.3464
R20663 commonsourceibias.n274 commonsourceibias.n252 24.3464
R20664 commonsourceibias.n285 commonsourceibias.n284 24.3464
R20665 commonsourceibias.n319 commonsourceibias.n318 24.3464
R20666 commonsourceibias.n233 commonsourceibias.n211 24.3464
R20667 commonsourceibias.n371 commonsourceibias.n349 24.3464
R20668 commonsourceibias.n382 commonsourceibias.n381 24.3464
R20669 commonsourceibias.n65 commonsourceibias.n10 23.8546
R20670 commonsourceibias.n27 commonsourceibias.n26 23.8546
R20671 commonsourceibias.n131 commonsourceibias.n1 23.8546
R20672 commonsourceibias.n93 commonsourceibias.n92 23.8546
R20673 commonsourceibias.n156 commonsourceibias.n155 23.8546
R20674 commonsourceibias.n194 commonsourceibias.n139 23.8546
R20675 commonsourceibias.n260 commonsourceibias.n259 23.8546
R20676 commonsourceibias.n299 commonsourceibias.n244 23.8546
R20677 commonsourceibias.n333 commonsourceibias.n203 23.8546
R20678 commonsourceibias.n219 commonsourceibias.n218 23.8546
R20679 commonsourceibias.n357 commonsourceibias.n356 23.8546
R20680 commonsourceibias.n396 commonsourceibias.n341 23.8546
R20681 commonsourceibias.n64 commonsourceibias.n63 16.9689
R20682 commonsourceibias.n28 commonsourceibias.n23 16.9689
R20683 commonsourceibias.n130 commonsourceibias.n129 16.9689
R20684 commonsourceibias.n94 commonsourceibias.n89 16.9689
R20685 commonsourceibias.n157 commonsourceibias.n152 16.9689
R20686 commonsourceibias.n193 commonsourceibias.n192 16.9689
R20687 commonsourceibias.n261 commonsourceibias.n256 16.9689
R20688 commonsourceibias.n298 commonsourceibias.n297 16.9689
R20689 commonsourceibias.n332 commonsourceibias.n331 16.9689
R20690 commonsourceibias.n220 commonsourceibias.n215 16.9689
R20691 commonsourceibias.n358 commonsourceibias.n353 16.9689
R20692 commonsourceibias.n395 commonsourceibias.n394 16.9689
R20693 commonsourceibias.n50 commonsourceibias.n49 16.477
R20694 commonsourceibias.n43 commonsourceibias.n42 16.477
R20695 commonsourceibias.n116 commonsourceibias.n115 16.477
R20696 commonsourceibias.n109 commonsourceibias.n108 16.477
R20697 commonsourceibias.n172 commonsourceibias.n171 16.477
R20698 commonsourceibias.n179 commonsourceibias.n178 16.477
R20699 commonsourceibias.n276 commonsourceibias.n275 16.477
R20700 commonsourceibias.n283 commonsourceibias.n282 16.477
R20701 commonsourceibias.n317 commonsourceibias.n316 16.477
R20702 commonsourceibias.n235 commonsourceibias.n234 16.477
R20703 commonsourceibias.n373 commonsourceibias.n372 16.477
R20704 commonsourceibias.n380 commonsourceibias.n379 16.477
R20705 commonsourceibias.n57 commonsourceibias.n56 15.9852
R20706 commonsourceibias.n36 commonsourceibias.n21 15.9852
R20707 commonsourceibias.n123 commonsourceibias.n122 15.9852
R20708 commonsourceibias.n102 commonsourceibias.n87 15.9852
R20709 commonsourceibias.n165 commonsourceibias.n150 15.9852
R20710 commonsourceibias.n186 commonsourceibias.n185 15.9852
R20711 commonsourceibias.n269 commonsourceibias.n254 15.9852
R20712 commonsourceibias.n291 commonsourceibias.n290 15.9852
R20713 commonsourceibias.n325 commonsourceibias.n324 15.9852
R20714 commonsourceibias.n228 commonsourceibias.n213 15.9852
R20715 commonsourceibias.n366 commonsourceibias.n351 15.9852
R20716 commonsourceibias.n388 commonsourceibias.n387 15.9852
R20717 commonsourceibias.n73 commonsourceibias.n71 13.2057
R20718 commonsourceibias.n307 commonsourceibias.n305 13.2057
R20719 commonsourceibias.n404 commonsourceibias.n201 11.9876
R20720 commonsourceibias.n404 commonsourceibias.n403 10.3347
R20721 commonsourceibias.n112 commonsourceibias.n83 9.50363
R20722 commonsourceibias.n313 commonsourceibias.n312 9.50363
R20723 commonsourceibias.n201 commonsourceibias.n137 8.732
R20724 commonsourceibias.n403 commonsourceibias.n339 8.732
R20725 commonsourceibias.n58 commonsourceibias.n57 8.60764
R20726 commonsourceibias.n33 commonsourceibias.n21 8.60764
R20727 commonsourceibias.n124 commonsourceibias.n123 8.60764
R20728 commonsourceibias.n99 commonsourceibias.n87 8.60764
R20729 commonsourceibias.n162 commonsourceibias.n150 8.60764
R20730 commonsourceibias.n187 commonsourceibias.n186 8.60764
R20731 commonsourceibias.n266 commonsourceibias.n254 8.60764
R20732 commonsourceibias.n292 commonsourceibias.n291 8.60764
R20733 commonsourceibias.n326 commonsourceibias.n325 8.60764
R20734 commonsourceibias.n225 commonsourceibias.n213 8.60764
R20735 commonsourceibias.n363 commonsourceibias.n351 8.60764
R20736 commonsourceibias.n389 commonsourceibias.n388 8.60764
R20737 commonsourceibias.n49 commonsourceibias.n48 8.11581
R20738 commonsourceibias.n44 commonsourceibias.n43 8.11581
R20739 commonsourceibias.n115 commonsourceibias.n114 8.11581
R20740 commonsourceibias.n110 commonsourceibias.n109 8.11581
R20741 commonsourceibias.n173 commonsourceibias.n172 8.11581
R20742 commonsourceibias.n178 commonsourceibias.n177 8.11581
R20743 commonsourceibias.n277 commonsourceibias.n276 8.11581
R20744 commonsourceibias.n282 commonsourceibias.n281 8.11581
R20745 commonsourceibias.n316 commonsourceibias.n315 8.11581
R20746 commonsourceibias.n236 commonsourceibias.n235 8.11581
R20747 commonsourceibias.n374 commonsourceibias.n373 8.11581
R20748 commonsourceibias.n379 commonsourceibias.n378 8.11581
R20749 commonsourceibias.n63 commonsourceibias.n62 7.62397
R20750 commonsourceibias.n31 commonsourceibias.n23 7.62397
R20751 commonsourceibias.n129 commonsourceibias.n128 7.62397
R20752 commonsourceibias.n97 commonsourceibias.n89 7.62397
R20753 commonsourceibias.n160 commonsourceibias.n152 7.62397
R20754 commonsourceibias.n192 commonsourceibias.n191 7.62397
R20755 commonsourceibias.n264 commonsourceibias.n256 7.62397
R20756 commonsourceibias.n297 commonsourceibias.n296 7.62397
R20757 commonsourceibias.n331 commonsourceibias.n330 7.62397
R20758 commonsourceibias.n223 commonsourceibias.n215 7.62397
R20759 commonsourceibias.n361 commonsourceibias.n353 7.62397
R20760 commonsourceibias.n394 commonsourceibias.n393 7.62397
R20761 commonsourceibias.n201 commonsourceibias.n200 5.00473
R20762 commonsourceibias.n403 commonsourceibias.n402 5.00473
R20763 commonsourceibias commonsourceibias.n404 3.87639
R20764 commonsourceibias.n78 commonsourceibias.t41 2.82907
R20765 commonsourceibias.n78 commonsourceibias.t47 2.82907
R20766 commonsourceibias.n79 commonsourceibias.t35 2.82907
R20767 commonsourceibias.n79 commonsourceibias.t11 2.82907
R20768 commonsourceibias.n81 commonsourceibias.t45 2.82907
R20769 commonsourceibias.n81 commonsourceibias.t27 2.82907
R20770 commonsourceibias.n76 commonsourceibias.t21 2.82907
R20771 commonsourceibias.n76 commonsourceibias.t37 2.82907
R20772 commonsourceibias.n74 commonsourceibias.t25 2.82907
R20773 commonsourceibias.n74 commonsourceibias.t31 2.82907
R20774 commonsourceibias.n72 commonsourceibias.t33 2.82907
R20775 commonsourceibias.n72 commonsourceibias.t15 2.82907
R20776 commonsourceibias.n306 commonsourceibias.t23 2.82907
R20777 commonsourceibias.n306 commonsourceibias.t3 2.82907
R20778 commonsourceibias.n308 commonsourceibias.t1 2.82907
R20779 commonsourceibias.n308 commonsourceibias.t39 2.82907
R20780 commonsourceibias.n310 commonsourceibias.t7 2.82907
R20781 commonsourceibias.n310 commonsourceibias.t29 2.82907
R20782 commonsourceibias.n241 commonsourceibias.t43 2.82907
R20783 commonsourceibias.n241 commonsourceibias.t13 2.82907
R20784 commonsourceibias.n239 commonsourceibias.t19 2.82907
R20785 commonsourceibias.n239 commonsourceibias.t5 2.82907
R20786 commonsourceibias.n238 commonsourceibias.t17 2.82907
R20787 commonsourceibias.n238 commonsourceibias.t9 2.82907
R20788 commonsourceibias.n68 commonsourceibias.n10 0.738255
R20789 commonsourceibias.n134 commonsourceibias.n1 0.738255
R20790 commonsourceibias.n197 commonsourceibias.n139 0.738255
R20791 commonsourceibias.n302 commonsourceibias.n244 0.738255
R20792 commonsourceibias.n336 commonsourceibias.n203 0.738255
R20793 commonsourceibias.n399 commonsourceibias.n341 0.738255
R20794 commonsourceibias.n75 commonsourceibias.n73 0.573776
R20795 commonsourceibias.n77 commonsourceibias.n75 0.573776
R20796 commonsourceibias.n82 commonsourceibias.n80 0.573776
R20797 commonsourceibias.n242 commonsourceibias.n240 0.573776
R20798 commonsourceibias.n311 commonsourceibias.n309 0.573776
R20799 commonsourceibias.n309 commonsourceibias.n307 0.573776
R20800 commonsourceibias.n83 commonsourceibias.n77 0.287138
R20801 commonsourceibias.n83 commonsourceibias.n82 0.287138
R20802 commonsourceibias.n312 commonsourceibias.n242 0.287138
R20803 commonsourceibias.n312 commonsourceibias.n311 0.287138
R20804 commonsourceibias.n71 commonsourceibias.n9 0.285035
R20805 commonsourceibias.n137 commonsourceibias.n0 0.285035
R20806 commonsourceibias.n200 commonsourceibias.n138 0.285035
R20807 commonsourceibias.n305 commonsourceibias.n243 0.285035
R20808 commonsourceibias.n339 commonsourceibias.n202 0.285035
R20809 commonsourceibias.n402 commonsourceibias.n340 0.285035
R20810 commonsourceibias.n16 commonsourceibias.n14 0.246418
R20811 commonsourceibias.n38 commonsourceibias.n19 0.246418
R20812 commonsourceibias.n7 commonsourceibias.n5 0.246418
R20813 commonsourceibias.n104 commonsourceibias.n85 0.246418
R20814 commonsourceibias.n167 commonsourceibias.n148 0.246418
R20815 commonsourceibias.n145 commonsourceibias.n143 0.246418
R20816 commonsourceibias.n271 commonsourceibias.n252 0.246418
R20817 commonsourceibias.n284 commonsourceibias.n248 0.246418
R20818 commonsourceibias.n318 commonsourceibias.n207 0.246418
R20819 commonsourceibias.n230 commonsourceibias.n211 0.246418
R20820 commonsourceibias.n368 commonsourceibias.n349 0.246418
R20821 commonsourceibias.n381 commonsourceibias.n345 0.246418
R20822 commonsourceibias.n67 commonsourceibias.n9 0.189894
R20823 commonsourceibias.n67 commonsourceibias.n66 0.189894
R20824 commonsourceibias.n66 commonsourceibias.n11 0.189894
R20825 commonsourceibias.n61 commonsourceibias.n11 0.189894
R20826 commonsourceibias.n61 commonsourceibias.n60 0.189894
R20827 commonsourceibias.n60 commonsourceibias.n59 0.189894
R20828 commonsourceibias.n59 commonsourceibias.n13 0.189894
R20829 commonsourceibias.n54 commonsourceibias.n13 0.189894
R20830 commonsourceibias.n54 commonsourceibias.n53 0.189894
R20831 commonsourceibias.n53 commonsourceibias.n52 0.189894
R20832 commonsourceibias.n52 commonsourceibias.n15 0.189894
R20833 commonsourceibias.n47 commonsourceibias.n15 0.189894
R20834 commonsourceibias.n47 commonsourceibias.n46 0.189894
R20835 commonsourceibias.n46 commonsourceibias.n45 0.189894
R20836 commonsourceibias.n45 commonsourceibias.n18 0.189894
R20837 commonsourceibias.n40 commonsourceibias.n18 0.189894
R20838 commonsourceibias.n40 commonsourceibias.n39 0.189894
R20839 commonsourceibias.n39 commonsourceibias.n20 0.189894
R20840 commonsourceibias.n35 commonsourceibias.n20 0.189894
R20841 commonsourceibias.n35 commonsourceibias.n34 0.189894
R20842 commonsourceibias.n34 commonsourceibias.n22 0.189894
R20843 commonsourceibias.n30 commonsourceibias.n22 0.189894
R20844 commonsourceibias.n30 commonsourceibias.n29 0.189894
R20845 commonsourceibias.n29 commonsourceibias.n24 0.189894
R20846 commonsourceibias.n111 commonsourceibias.n84 0.189894
R20847 commonsourceibias.n106 commonsourceibias.n84 0.189894
R20848 commonsourceibias.n106 commonsourceibias.n105 0.189894
R20849 commonsourceibias.n105 commonsourceibias.n86 0.189894
R20850 commonsourceibias.n101 commonsourceibias.n86 0.189894
R20851 commonsourceibias.n101 commonsourceibias.n100 0.189894
R20852 commonsourceibias.n100 commonsourceibias.n88 0.189894
R20853 commonsourceibias.n96 commonsourceibias.n88 0.189894
R20854 commonsourceibias.n96 commonsourceibias.n95 0.189894
R20855 commonsourceibias.n95 commonsourceibias.n90 0.189894
R20856 commonsourceibias.n133 commonsourceibias.n0 0.189894
R20857 commonsourceibias.n133 commonsourceibias.n132 0.189894
R20858 commonsourceibias.n132 commonsourceibias.n2 0.189894
R20859 commonsourceibias.n127 commonsourceibias.n2 0.189894
R20860 commonsourceibias.n127 commonsourceibias.n126 0.189894
R20861 commonsourceibias.n126 commonsourceibias.n125 0.189894
R20862 commonsourceibias.n125 commonsourceibias.n4 0.189894
R20863 commonsourceibias.n120 commonsourceibias.n4 0.189894
R20864 commonsourceibias.n120 commonsourceibias.n119 0.189894
R20865 commonsourceibias.n119 commonsourceibias.n118 0.189894
R20866 commonsourceibias.n118 commonsourceibias.n6 0.189894
R20867 commonsourceibias.n113 commonsourceibias.n6 0.189894
R20868 commonsourceibias.n196 commonsourceibias.n138 0.189894
R20869 commonsourceibias.n196 commonsourceibias.n195 0.189894
R20870 commonsourceibias.n195 commonsourceibias.n140 0.189894
R20871 commonsourceibias.n190 commonsourceibias.n140 0.189894
R20872 commonsourceibias.n190 commonsourceibias.n189 0.189894
R20873 commonsourceibias.n189 commonsourceibias.n188 0.189894
R20874 commonsourceibias.n188 commonsourceibias.n142 0.189894
R20875 commonsourceibias.n183 commonsourceibias.n142 0.189894
R20876 commonsourceibias.n183 commonsourceibias.n182 0.189894
R20877 commonsourceibias.n182 commonsourceibias.n181 0.189894
R20878 commonsourceibias.n181 commonsourceibias.n144 0.189894
R20879 commonsourceibias.n176 commonsourceibias.n144 0.189894
R20880 commonsourceibias.n176 commonsourceibias.n175 0.189894
R20881 commonsourceibias.n175 commonsourceibias.n174 0.189894
R20882 commonsourceibias.n174 commonsourceibias.n147 0.189894
R20883 commonsourceibias.n169 commonsourceibias.n147 0.189894
R20884 commonsourceibias.n169 commonsourceibias.n168 0.189894
R20885 commonsourceibias.n168 commonsourceibias.n149 0.189894
R20886 commonsourceibias.n164 commonsourceibias.n149 0.189894
R20887 commonsourceibias.n164 commonsourceibias.n163 0.189894
R20888 commonsourceibias.n163 commonsourceibias.n151 0.189894
R20889 commonsourceibias.n159 commonsourceibias.n151 0.189894
R20890 commonsourceibias.n159 commonsourceibias.n158 0.189894
R20891 commonsourceibias.n158 commonsourceibias.n153 0.189894
R20892 commonsourceibias.n262 commonsourceibias.n257 0.189894
R20893 commonsourceibias.n263 commonsourceibias.n262 0.189894
R20894 commonsourceibias.n263 commonsourceibias.n255 0.189894
R20895 commonsourceibias.n267 commonsourceibias.n255 0.189894
R20896 commonsourceibias.n268 commonsourceibias.n267 0.189894
R20897 commonsourceibias.n268 commonsourceibias.n253 0.189894
R20898 commonsourceibias.n272 commonsourceibias.n253 0.189894
R20899 commonsourceibias.n273 commonsourceibias.n272 0.189894
R20900 commonsourceibias.n273 commonsourceibias.n251 0.189894
R20901 commonsourceibias.n278 commonsourceibias.n251 0.189894
R20902 commonsourceibias.n279 commonsourceibias.n278 0.189894
R20903 commonsourceibias.n280 commonsourceibias.n279 0.189894
R20904 commonsourceibias.n280 commonsourceibias.n249 0.189894
R20905 commonsourceibias.n286 commonsourceibias.n249 0.189894
R20906 commonsourceibias.n287 commonsourceibias.n286 0.189894
R20907 commonsourceibias.n288 commonsourceibias.n287 0.189894
R20908 commonsourceibias.n288 commonsourceibias.n247 0.189894
R20909 commonsourceibias.n293 commonsourceibias.n247 0.189894
R20910 commonsourceibias.n294 commonsourceibias.n293 0.189894
R20911 commonsourceibias.n295 commonsourceibias.n294 0.189894
R20912 commonsourceibias.n295 commonsourceibias.n245 0.189894
R20913 commonsourceibias.n300 commonsourceibias.n245 0.189894
R20914 commonsourceibias.n301 commonsourceibias.n300 0.189894
R20915 commonsourceibias.n301 commonsourceibias.n243 0.189894
R20916 commonsourceibias.n221 commonsourceibias.n216 0.189894
R20917 commonsourceibias.n222 commonsourceibias.n221 0.189894
R20918 commonsourceibias.n222 commonsourceibias.n214 0.189894
R20919 commonsourceibias.n226 commonsourceibias.n214 0.189894
R20920 commonsourceibias.n227 commonsourceibias.n226 0.189894
R20921 commonsourceibias.n227 commonsourceibias.n212 0.189894
R20922 commonsourceibias.n231 commonsourceibias.n212 0.189894
R20923 commonsourceibias.n232 commonsourceibias.n231 0.189894
R20924 commonsourceibias.n232 commonsourceibias.n210 0.189894
R20925 commonsourceibias.n237 commonsourceibias.n210 0.189894
R20926 commonsourceibias.n314 commonsourceibias.n208 0.189894
R20927 commonsourceibias.n320 commonsourceibias.n208 0.189894
R20928 commonsourceibias.n321 commonsourceibias.n320 0.189894
R20929 commonsourceibias.n322 commonsourceibias.n321 0.189894
R20930 commonsourceibias.n322 commonsourceibias.n206 0.189894
R20931 commonsourceibias.n327 commonsourceibias.n206 0.189894
R20932 commonsourceibias.n328 commonsourceibias.n327 0.189894
R20933 commonsourceibias.n329 commonsourceibias.n328 0.189894
R20934 commonsourceibias.n329 commonsourceibias.n204 0.189894
R20935 commonsourceibias.n334 commonsourceibias.n204 0.189894
R20936 commonsourceibias.n335 commonsourceibias.n334 0.189894
R20937 commonsourceibias.n335 commonsourceibias.n202 0.189894
R20938 commonsourceibias.n359 commonsourceibias.n354 0.189894
R20939 commonsourceibias.n360 commonsourceibias.n359 0.189894
R20940 commonsourceibias.n360 commonsourceibias.n352 0.189894
R20941 commonsourceibias.n364 commonsourceibias.n352 0.189894
R20942 commonsourceibias.n365 commonsourceibias.n364 0.189894
R20943 commonsourceibias.n365 commonsourceibias.n350 0.189894
R20944 commonsourceibias.n369 commonsourceibias.n350 0.189894
R20945 commonsourceibias.n370 commonsourceibias.n369 0.189894
R20946 commonsourceibias.n370 commonsourceibias.n348 0.189894
R20947 commonsourceibias.n375 commonsourceibias.n348 0.189894
R20948 commonsourceibias.n376 commonsourceibias.n375 0.189894
R20949 commonsourceibias.n377 commonsourceibias.n376 0.189894
R20950 commonsourceibias.n377 commonsourceibias.n346 0.189894
R20951 commonsourceibias.n383 commonsourceibias.n346 0.189894
R20952 commonsourceibias.n384 commonsourceibias.n383 0.189894
R20953 commonsourceibias.n385 commonsourceibias.n384 0.189894
R20954 commonsourceibias.n385 commonsourceibias.n344 0.189894
R20955 commonsourceibias.n390 commonsourceibias.n344 0.189894
R20956 commonsourceibias.n391 commonsourceibias.n390 0.189894
R20957 commonsourceibias.n392 commonsourceibias.n391 0.189894
R20958 commonsourceibias.n392 commonsourceibias.n342 0.189894
R20959 commonsourceibias.n397 commonsourceibias.n342 0.189894
R20960 commonsourceibias.n398 commonsourceibias.n397 0.189894
R20961 commonsourceibias.n398 commonsourceibias.n340 0.189894
R20962 commonsourceibias.n112 commonsourceibias.n111 0.170955
R20963 commonsourceibias.n113 commonsourceibias.n112 0.170955
R20964 commonsourceibias.n313 commonsourceibias.n237 0.170955
R20965 commonsourceibias.n314 commonsourceibias.n313 0.170955
R20966 plus.n46 plus.t9 252.611
R20967 plus.n9 plus.t11 252.611
R20968 plus.n76 plus.t4 243.97
R20969 plus.n72 plus.t12 231.093
R20970 plus.n35 plus.t7 231.093
R20971 plus.n76 plus.n75 223.454
R20972 plus.n78 plus.n77 223.454
R20973 plus.n47 plus.t5 187.445
R20974 plus.n44 plus.t18 187.445
R20975 plus.n42 plus.t17 187.445
R20976 plus.n59 plus.t13 187.445
R20977 plus.n65 plus.t14 187.445
R20978 plus.n38 plus.t10 187.445
R20979 plus.n1 plus.t6 187.445
R20980 plus.n28 plus.t16 187.445
R20981 plus.n22 plus.t15 187.445
R20982 plus.n5 plus.t20 187.445
R20983 plus.n7 plus.t19 187.445
R20984 plus.n10 plus.t8 187.445
R20985 plus.n73 plus.n72 161.3
R20986 plus.n71 plus.n37 161.3
R20987 plus.n70 plus.n69 161.3
R20988 plus.n68 plus.n67 161.3
R20989 plus.n66 plus.n39 161.3
R20990 plus.n64 plus.n63 161.3
R20991 plus.n62 plus.n40 161.3
R20992 plus.n61 plus.n60 161.3
R20993 plus.n58 plus.n41 161.3
R20994 plus.n57 plus.n56 161.3
R20995 plus.n55 plus.n54 161.3
R20996 plus.n53 plus.n43 161.3
R20997 plus.n52 plus.n51 161.3
R20998 plus.n50 plus.n49 161.3
R20999 plus.n48 plus.n45 161.3
R21000 plus.n11 plus.n8 161.3
R21001 plus.n13 plus.n12 161.3
R21002 plus.n15 plus.n14 161.3
R21003 plus.n16 plus.n6 161.3
R21004 plus.n18 plus.n17 161.3
R21005 plus.n20 plus.n19 161.3
R21006 plus.n21 plus.n4 161.3
R21007 plus.n24 plus.n23 161.3
R21008 plus.n25 plus.n3 161.3
R21009 plus.n27 plus.n26 161.3
R21010 plus.n29 plus.n2 161.3
R21011 plus.n31 plus.n30 161.3
R21012 plus.n33 plus.n32 161.3
R21013 plus.n34 plus.n0 161.3
R21014 plus.n36 plus.n35 161.3
R21015 plus.n49 plus.n48 56.5617
R21016 plus.n58 plus.n57 56.5617
R21017 plus.n67 plus.n66 56.5617
R21018 plus.n30 plus.n29 56.5617
R21019 plus.n21 plus.n20 56.5617
R21020 plus.n12 plus.n11 56.5617
R21021 plus.n71 plus.n70 46.3896
R21022 plus.n34 plus.n33 46.3896
R21023 plus.n46 plus.n45 42.8164
R21024 plus.n9 plus.n8 42.8164
R21025 plus.n54 plus.n53 42.5146
R21026 plus.n60 plus.n40 42.5146
R21027 plus.n23 plus.n3 42.5146
R21028 plus.n17 plus.n16 42.5146
R21029 plus.n53 plus.n52 38.6395
R21030 plus.n64 plus.n40 38.6395
R21031 plus.n27 plus.n3 38.6395
R21032 plus.n16 plus.n15 38.6395
R21033 plus.n47 plus.n46 38.2514
R21034 plus.n10 plus.n9 38.2514
R21035 plus.n74 plus.n73 31.491
R21036 plus.n49 plus.n44 19.9199
R21037 plus.n66 plus.n65 19.9199
R21038 plus.n29 plus.n28 19.9199
R21039 plus.n12 plus.n7 19.9199
R21040 plus.n75 plus.t1 19.8005
R21041 plus.n75 plus.t2 19.8005
R21042 plus.n77 plus.t0 19.8005
R21043 plus.n77 plus.t3 19.8005
R21044 plus.n57 plus.n42 17.9525
R21045 plus.n59 plus.n58 17.9525
R21046 plus.n22 plus.n21 17.9525
R21047 plus.n20 plus.n5 17.9525
R21048 plus.n48 plus.n47 15.9852
R21049 plus.n67 plus.n38 15.9852
R21050 plus.n30 plus.n1 15.9852
R21051 plus.n11 plus.n10 15.9852
R21052 plus.n72 plus.n71 15.3369
R21053 plus.n35 plus.n34 15.3369
R21054 plus plus.n79 14.0959
R21055 plus.n74 plus.n36 11.9494
R21056 plus.n70 plus.n38 8.60764
R21057 plus.n33 plus.n1 8.60764
R21058 plus.n54 plus.n42 6.6403
R21059 plus.n60 plus.n59 6.6403
R21060 plus.n23 plus.n22 6.6403
R21061 plus.n17 plus.n5 6.6403
R21062 plus.n79 plus.n78 5.40567
R21063 plus.n52 plus.n44 4.67295
R21064 plus.n65 plus.n64 4.67295
R21065 plus.n28 plus.n27 4.67295
R21066 plus.n15 plus.n7 4.67295
R21067 plus.n79 plus.n74 1.188
R21068 plus.n78 plus.n76 0.716017
R21069 plus.n50 plus.n45 0.189894
R21070 plus.n51 plus.n50 0.189894
R21071 plus.n51 plus.n43 0.189894
R21072 plus.n55 plus.n43 0.189894
R21073 plus.n56 plus.n55 0.189894
R21074 plus.n56 plus.n41 0.189894
R21075 plus.n61 plus.n41 0.189894
R21076 plus.n62 plus.n61 0.189894
R21077 plus.n63 plus.n62 0.189894
R21078 plus.n63 plus.n39 0.189894
R21079 plus.n68 plus.n39 0.189894
R21080 plus.n69 plus.n68 0.189894
R21081 plus.n69 plus.n37 0.189894
R21082 plus.n73 plus.n37 0.189894
R21083 plus.n36 plus.n0 0.189894
R21084 plus.n32 plus.n0 0.189894
R21085 plus.n32 plus.n31 0.189894
R21086 plus.n31 plus.n2 0.189894
R21087 plus.n26 plus.n2 0.189894
R21088 plus.n26 plus.n25 0.189894
R21089 plus.n25 plus.n24 0.189894
R21090 plus.n24 plus.n4 0.189894
R21091 plus.n19 plus.n4 0.189894
R21092 plus.n19 plus.n18 0.189894
R21093 plus.n18 plus.n6 0.189894
R21094 plus.n14 plus.n6 0.189894
R21095 plus.n14 plus.n13 0.189894
R21096 plus.n13 plus.n8 0.189894
R21097 a_n2903_n3924.n0 a_n2903_n3924.t37 214.981
R21098 a_n2903_n3924.n2 a_n2903_n3924.t2 214.452
R21099 a_n2903_n3924.n11 a_n2903_n3924.t38 214.321
R21100 a_n2903_n3924.n12 a_n2903_n3924.t36 214.321
R21101 a_n2903_n3924.n13 a_n2903_n3924.t1 214.321
R21102 a_n2903_n3924.n14 a_n2903_n3924.t0 214.321
R21103 a_n2903_n3924.n15 a_n2903_n3924.t3 214.321
R21104 a_n2903_n3924.n0 a_n2903_n3924.t39 214.321
R21105 a_n2903_n3924.n1 a_n2903_n3924.t31 55.8337
R21106 a_n2903_n3924.n3 a_n2903_n3924.t6 55.8337
R21107 a_n2903_n3924.n10 a_n2903_n3924.t11 55.8337
R21108 a_n2903_n3924.n34 a_n2903_n3924.t28 55.8335
R21109 a_n2903_n3924.n32 a_n2903_n3924.t9 55.8335
R21110 a_n2903_n3924.n25 a_n2903_n3924.t13 55.8335
R21111 a_n2903_n3924.n24 a_n2903_n3924.t29 55.8335
R21112 a_n2903_n3924.n17 a_n2903_n3924.t33 55.8335
R21113 a_n2903_n3924.n36 a_n2903_n3924.n35 53.0052
R21114 a_n2903_n3924.n38 a_n2903_n3924.n37 53.0052
R21115 a_n2903_n3924.n5 a_n2903_n3924.n4 53.0052
R21116 a_n2903_n3924.n7 a_n2903_n3924.n6 53.0052
R21117 a_n2903_n3924.n9 a_n2903_n3924.n8 53.0052
R21118 a_n2903_n3924.n31 a_n2903_n3924.n30 53.0051
R21119 a_n2903_n3924.n29 a_n2903_n3924.n28 53.0051
R21120 a_n2903_n3924.n27 a_n2903_n3924.n26 53.0051
R21121 a_n2903_n3924.n23 a_n2903_n3924.n22 53.0051
R21122 a_n2903_n3924.n21 a_n2903_n3924.n20 53.0051
R21123 a_n2903_n3924.n19 a_n2903_n3924.n18 53.0051
R21124 a_n2903_n3924.n40 a_n2903_n3924.n39 53.0051
R21125 a_n2903_n3924.n16 a_n2903_n3924.n10 12.2417
R21126 a_n2903_n3924.n34 a_n2903_n3924.n33 12.2417
R21127 a_n2903_n3924.n17 a_n2903_n3924.n16 5.16214
R21128 a_n2903_n3924.n33 a_n2903_n3924.n32 5.16214
R21129 a_n2903_n3924.n35 a_n2903_n3924.t26 2.82907
R21130 a_n2903_n3924.n35 a_n2903_n3924.t30 2.82907
R21131 a_n2903_n3924.n37 a_n2903_n3924.t23 2.82907
R21132 a_n2903_n3924.n37 a_n2903_n3924.t27 2.82907
R21133 a_n2903_n3924.n4 a_n2903_n3924.t8 2.82907
R21134 a_n2903_n3924.n4 a_n2903_n3924.t10 2.82907
R21135 a_n2903_n3924.n6 a_n2903_n3924.t19 2.82907
R21136 a_n2903_n3924.n6 a_n2903_n3924.t7 2.82907
R21137 a_n2903_n3924.n8 a_n2903_n3924.t14 2.82907
R21138 a_n2903_n3924.n8 a_n2903_n3924.t17 2.82907
R21139 a_n2903_n3924.n30 a_n2903_n3924.t4 2.82907
R21140 a_n2903_n3924.n30 a_n2903_n3924.t12 2.82907
R21141 a_n2903_n3924.n28 a_n2903_n3924.t18 2.82907
R21142 a_n2903_n3924.n28 a_n2903_n3924.t5 2.82907
R21143 a_n2903_n3924.n26 a_n2903_n3924.t15 2.82907
R21144 a_n2903_n3924.n26 a_n2903_n3924.t16 2.82907
R21145 a_n2903_n3924.n22 a_n2903_n3924.t21 2.82907
R21146 a_n2903_n3924.n22 a_n2903_n3924.t32 2.82907
R21147 a_n2903_n3924.n20 a_n2903_n3924.t25 2.82907
R21148 a_n2903_n3924.n20 a_n2903_n3924.t20 2.82907
R21149 a_n2903_n3924.n18 a_n2903_n3924.t34 2.82907
R21150 a_n2903_n3924.n18 a_n2903_n3924.t24 2.82907
R21151 a_n2903_n3924.t35 a_n2903_n3924.n40 2.82907
R21152 a_n2903_n3924.n40 a_n2903_n3924.t22 2.82907
R21153 a_n2903_n3924.n33 a_n2903_n3924.n2 1.95694
R21154 a_n2903_n3924.n16 a_n2903_n3924.n0 1.95694
R21155 a_n2903_n3924.n0 a_n2903_n3924.n15 0.684366
R21156 a_n2903_n3924.n15 a_n2903_n3924.n14 0.672012
R21157 a_n2903_n3924.n14 a_n2903_n3924.n13 0.672012
R21158 a_n2903_n3924.n13 a_n2903_n3924.n12 0.672012
R21159 a_n2903_n3924.n12 a_n2903_n3924.n11 0.672012
R21160 a_n2903_n3924.n11 a_n2903_n3924.n2 0.541924
R21161 a_n2903_n3924.n19 a_n2903_n3924.n17 0.530672
R21162 a_n2903_n3924.n21 a_n2903_n3924.n19 0.530672
R21163 a_n2903_n3924.n23 a_n2903_n3924.n21 0.530672
R21164 a_n2903_n3924.n24 a_n2903_n3924.n23 0.530672
R21165 a_n2903_n3924.n27 a_n2903_n3924.n25 0.530672
R21166 a_n2903_n3924.n29 a_n2903_n3924.n27 0.530672
R21167 a_n2903_n3924.n31 a_n2903_n3924.n29 0.530672
R21168 a_n2903_n3924.n32 a_n2903_n3924.n31 0.530672
R21169 a_n2903_n3924.n10 a_n2903_n3924.n9 0.530672
R21170 a_n2903_n3924.n9 a_n2903_n3924.n7 0.530672
R21171 a_n2903_n3924.n7 a_n2903_n3924.n5 0.530672
R21172 a_n2903_n3924.n5 a_n2903_n3924.n3 0.530672
R21173 a_n2903_n3924.n39 a_n2903_n3924.n1 0.530672
R21174 a_n2903_n3924.n39 a_n2903_n3924.n38 0.530672
R21175 a_n2903_n3924.n38 a_n2903_n3924.n36 0.530672
R21176 a_n2903_n3924.n36 a_n2903_n3924.n34 0.530672
R21177 a_n2903_n3924.n25 a_n2903_n3924.n24 0.235414
R21178 a_n2903_n3924.n3 a_n2903_n3924.n1 0.235414
R21179 outputibias.n27 outputibias.n1 289.615
R21180 outputibias.n58 outputibias.n32 289.615
R21181 outputibias.n90 outputibias.n64 289.615
R21182 outputibias.n122 outputibias.n96 289.615
R21183 outputibias.n28 outputibias.n27 185
R21184 outputibias.n26 outputibias.n25 185
R21185 outputibias.n5 outputibias.n4 185
R21186 outputibias.n20 outputibias.n19 185
R21187 outputibias.n18 outputibias.n17 185
R21188 outputibias.n9 outputibias.n8 185
R21189 outputibias.n12 outputibias.n11 185
R21190 outputibias.n59 outputibias.n58 185
R21191 outputibias.n57 outputibias.n56 185
R21192 outputibias.n36 outputibias.n35 185
R21193 outputibias.n51 outputibias.n50 185
R21194 outputibias.n49 outputibias.n48 185
R21195 outputibias.n40 outputibias.n39 185
R21196 outputibias.n43 outputibias.n42 185
R21197 outputibias.n91 outputibias.n90 185
R21198 outputibias.n89 outputibias.n88 185
R21199 outputibias.n68 outputibias.n67 185
R21200 outputibias.n83 outputibias.n82 185
R21201 outputibias.n81 outputibias.n80 185
R21202 outputibias.n72 outputibias.n71 185
R21203 outputibias.n75 outputibias.n74 185
R21204 outputibias.n123 outputibias.n122 185
R21205 outputibias.n121 outputibias.n120 185
R21206 outputibias.n100 outputibias.n99 185
R21207 outputibias.n115 outputibias.n114 185
R21208 outputibias.n113 outputibias.n112 185
R21209 outputibias.n104 outputibias.n103 185
R21210 outputibias.n107 outputibias.n106 185
R21211 outputibias.n0 outputibias.t8 178.945
R21212 outputibias.n133 outputibias.t10 177.018
R21213 outputibias.n132 outputibias.t11 177.018
R21214 outputibias.n0 outputibias.t9 177.018
R21215 outputibias.t5 outputibias.n10 147.661
R21216 outputibias.t7 outputibias.n41 147.661
R21217 outputibias.t1 outputibias.n73 147.661
R21218 outputibias.t3 outputibias.n105 147.661
R21219 outputibias.n128 outputibias.t4 132.363
R21220 outputibias.n128 outputibias.t6 130.436
R21221 outputibias.n129 outputibias.t0 130.436
R21222 outputibias.n130 outputibias.t2 130.436
R21223 outputibias.n27 outputibias.n26 104.615
R21224 outputibias.n26 outputibias.n4 104.615
R21225 outputibias.n19 outputibias.n4 104.615
R21226 outputibias.n19 outputibias.n18 104.615
R21227 outputibias.n18 outputibias.n8 104.615
R21228 outputibias.n11 outputibias.n8 104.615
R21229 outputibias.n58 outputibias.n57 104.615
R21230 outputibias.n57 outputibias.n35 104.615
R21231 outputibias.n50 outputibias.n35 104.615
R21232 outputibias.n50 outputibias.n49 104.615
R21233 outputibias.n49 outputibias.n39 104.615
R21234 outputibias.n42 outputibias.n39 104.615
R21235 outputibias.n90 outputibias.n89 104.615
R21236 outputibias.n89 outputibias.n67 104.615
R21237 outputibias.n82 outputibias.n67 104.615
R21238 outputibias.n82 outputibias.n81 104.615
R21239 outputibias.n81 outputibias.n71 104.615
R21240 outputibias.n74 outputibias.n71 104.615
R21241 outputibias.n122 outputibias.n121 104.615
R21242 outputibias.n121 outputibias.n99 104.615
R21243 outputibias.n114 outputibias.n99 104.615
R21244 outputibias.n114 outputibias.n113 104.615
R21245 outputibias.n113 outputibias.n103 104.615
R21246 outputibias.n106 outputibias.n103 104.615
R21247 outputibias.n63 outputibias.n31 95.6354
R21248 outputibias.n63 outputibias.n62 94.6732
R21249 outputibias.n95 outputibias.n94 94.6732
R21250 outputibias.n127 outputibias.n126 94.6732
R21251 outputibias.n11 outputibias.t5 52.3082
R21252 outputibias.n42 outputibias.t7 52.3082
R21253 outputibias.n74 outputibias.t1 52.3082
R21254 outputibias.n106 outputibias.t3 52.3082
R21255 outputibias.n12 outputibias.n10 15.6674
R21256 outputibias.n43 outputibias.n41 15.6674
R21257 outputibias.n75 outputibias.n73 15.6674
R21258 outputibias.n107 outputibias.n105 15.6674
R21259 outputibias.n13 outputibias.n9 12.8005
R21260 outputibias.n44 outputibias.n40 12.8005
R21261 outputibias.n76 outputibias.n72 12.8005
R21262 outputibias.n108 outputibias.n104 12.8005
R21263 outputibias.n17 outputibias.n16 12.0247
R21264 outputibias.n48 outputibias.n47 12.0247
R21265 outputibias.n80 outputibias.n79 12.0247
R21266 outputibias.n112 outputibias.n111 12.0247
R21267 outputibias.n20 outputibias.n7 11.249
R21268 outputibias.n51 outputibias.n38 11.249
R21269 outputibias.n83 outputibias.n70 11.249
R21270 outputibias.n115 outputibias.n102 11.249
R21271 outputibias.n21 outputibias.n5 10.4732
R21272 outputibias.n52 outputibias.n36 10.4732
R21273 outputibias.n84 outputibias.n68 10.4732
R21274 outputibias.n116 outputibias.n100 10.4732
R21275 outputibias.n25 outputibias.n24 9.69747
R21276 outputibias.n56 outputibias.n55 9.69747
R21277 outputibias.n88 outputibias.n87 9.69747
R21278 outputibias.n120 outputibias.n119 9.69747
R21279 outputibias.n31 outputibias.n30 9.45567
R21280 outputibias.n62 outputibias.n61 9.45567
R21281 outputibias.n94 outputibias.n93 9.45567
R21282 outputibias.n126 outputibias.n125 9.45567
R21283 outputibias.n30 outputibias.n29 9.3005
R21284 outputibias.n3 outputibias.n2 9.3005
R21285 outputibias.n24 outputibias.n23 9.3005
R21286 outputibias.n22 outputibias.n21 9.3005
R21287 outputibias.n7 outputibias.n6 9.3005
R21288 outputibias.n16 outputibias.n15 9.3005
R21289 outputibias.n14 outputibias.n13 9.3005
R21290 outputibias.n61 outputibias.n60 9.3005
R21291 outputibias.n34 outputibias.n33 9.3005
R21292 outputibias.n55 outputibias.n54 9.3005
R21293 outputibias.n53 outputibias.n52 9.3005
R21294 outputibias.n38 outputibias.n37 9.3005
R21295 outputibias.n47 outputibias.n46 9.3005
R21296 outputibias.n45 outputibias.n44 9.3005
R21297 outputibias.n93 outputibias.n92 9.3005
R21298 outputibias.n66 outputibias.n65 9.3005
R21299 outputibias.n87 outputibias.n86 9.3005
R21300 outputibias.n85 outputibias.n84 9.3005
R21301 outputibias.n70 outputibias.n69 9.3005
R21302 outputibias.n79 outputibias.n78 9.3005
R21303 outputibias.n77 outputibias.n76 9.3005
R21304 outputibias.n125 outputibias.n124 9.3005
R21305 outputibias.n98 outputibias.n97 9.3005
R21306 outputibias.n119 outputibias.n118 9.3005
R21307 outputibias.n117 outputibias.n116 9.3005
R21308 outputibias.n102 outputibias.n101 9.3005
R21309 outputibias.n111 outputibias.n110 9.3005
R21310 outputibias.n109 outputibias.n108 9.3005
R21311 outputibias.n28 outputibias.n3 8.92171
R21312 outputibias.n59 outputibias.n34 8.92171
R21313 outputibias.n91 outputibias.n66 8.92171
R21314 outputibias.n123 outputibias.n98 8.92171
R21315 outputibias.n29 outputibias.n1 8.14595
R21316 outputibias.n60 outputibias.n32 8.14595
R21317 outputibias.n92 outputibias.n64 8.14595
R21318 outputibias.n124 outputibias.n96 8.14595
R21319 outputibias.n31 outputibias.n1 5.81868
R21320 outputibias.n62 outputibias.n32 5.81868
R21321 outputibias.n94 outputibias.n64 5.81868
R21322 outputibias.n126 outputibias.n96 5.81868
R21323 outputibias.n131 outputibias.n130 5.20947
R21324 outputibias.n29 outputibias.n28 5.04292
R21325 outputibias.n60 outputibias.n59 5.04292
R21326 outputibias.n92 outputibias.n91 5.04292
R21327 outputibias.n124 outputibias.n123 5.04292
R21328 outputibias.n131 outputibias.n127 4.42209
R21329 outputibias.n14 outputibias.n10 4.38594
R21330 outputibias.n45 outputibias.n41 4.38594
R21331 outputibias.n77 outputibias.n73 4.38594
R21332 outputibias.n109 outputibias.n105 4.38594
R21333 outputibias.n132 outputibias.n131 4.28454
R21334 outputibias.n25 outputibias.n3 4.26717
R21335 outputibias.n56 outputibias.n34 4.26717
R21336 outputibias.n88 outputibias.n66 4.26717
R21337 outputibias.n120 outputibias.n98 4.26717
R21338 outputibias.n24 outputibias.n5 3.49141
R21339 outputibias.n55 outputibias.n36 3.49141
R21340 outputibias.n87 outputibias.n68 3.49141
R21341 outputibias.n119 outputibias.n100 3.49141
R21342 outputibias.n21 outputibias.n20 2.71565
R21343 outputibias.n52 outputibias.n51 2.71565
R21344 outputibias.n84 outputibias.n83 2.71565
R21345 outputibias.n116 outputibias.n115 2.71565
R21346 outputibias.n17 outputibias.n7 1.93989
R21347 outputibias.n48 outputibias.n38 1.93989
R21348 outputibias.n80 outputibias.n70 1.93989
R21349 outputibias.n112 outputibias.n102 1.93989
R21350 outputibias.n130 outputibias.n129 1.9266
R21351 outputibias.n129 outputibias.n128 1.9266
R21352 outputibias.n133 outputibias.n132 1.92658
R21353 outputibias.n134 outputibias.n133 1.29913
R21354 outputibias.n16 outputibias.n9 1.16414
R21355 outputibias.n47 outputibias.n40 1.16414
R21356 outputibias.n79 outputibias.n72 1.16414
R21357 outputibias.n111 outputibias.n104 1.16414
R21358 outputibias.n127 outputibias.n95 0.962709
R21359 outputibias.n95 outputibias.n63 0.962709
R21360 outputibias.n13 outputibias.n12 0.388379
R21361 outputibias.n44 outputibias.n43 0.388379
R21362 outputibias.n76 outputibias.n75 0.388379
R21363 outputibias.n108 outputibias.n107 0.388379
R21364 outputibias.n134 outputibias.n0 0.337251
R21365 outputibias outputibias.n134 0.302375
R21366 outputibias.n30 outputibias.n2 0.155672
R21367 outputibias.n23 outputibias.n2 0.155672
R21368 outputibias.n23 outputibias.n22 0.155672
R21369 outputibias.n22 outputibias.n6 0.155672
R21370 outputibias.n15 outputibias.n6 0.155672
R21371 outputibias.n15 outputibias.n14 0.155672
R21372 outputibias.n61 outputibias.n33 0.155672
R21373 outputibias.n54 outputibias.n33 0.155672
R21374 outputibias.n54 outputibias.n53 0.155672
R21375 outputibias.n53 outputibias.n37 0.155672
R21376 outputibias.n46 outputibias.n37 0.155672
R21377 outputibias.n46 outputibias.n45 0.155672
R21378 outputibias.n93 outputibias.n65 0.155672
R21379 outputibias.n86 outputibias.n65 0.155672
R21380 outputibias.n86 outputibias.n85 0.155672
R21381 outputibias.n85 outputibias.n69 0.155672
R21382 outputibias.n78 outputibias.n69 0.155672
R21383 outputibias.n78 outputibias.n77 0.155672
R21384 outputibias.n125 outputibias.n97 0.155672
R21385 outputibias.n118 outputibias.n97 0.155672
R21386 outputibias.n118 outputibias.n117 0.155672
R21387 outputibias.n117 outputibias.n101 0.155672
R21388 outputibias.n110 outputibias.n101 0.155672
R21389 outputibias.n110 outputibias.n109 0.155672
R21390 output.n41 output.n15 289.615
R21391 output.n72 output.n46 289.615
R21392 output.n104 output.n78 289.615
R21393 output.n136 output.n110 289.615
R21394 output.n77 output.n45 197.26
R21395 output.n77 output.n76 196.298
R21396 output.n109 output.n108 196.298
R21397 output.n141 output.n140 196.298
R21398 output.n42 output.n41 185
R21399 output.n40 output.n39 185
R21400 output.n19 output.n18 185
R21401 output.n34 output.n33 185
R21402 output.n32 output.n31 185
R21403 output.n23 output.n22 185
R21404 output.n26 output.n25 185
R21405 output.n73 output.n72 185
R21406 output.n71 output.n70 185
R21407 output.n50 output.n49 185
R21408 output.n65 output.n64 185
R21409 output.n63 output.n62 185
R21410 output.n54 output.n53 185
R21411 output.n57 output.n56 185
R21412 output.n105 output.n104 185
R21413 output.n103 output.n102 185
R21414 output.n82 output.n81 185
R21415 output.n97 output.n96 185
R21416 output.n95 output.n94 185
R21417 output.n86 output.n85 185
R21418 output.n89 output.n88 185
R21419 output.n137 output.n136 185
R21420 output.n135 output.n134 185
R21421 output.n114 output.n113 185
R21422 output.n129 output.n128 185
R21423 output.n127 output.n126 185
R21424 output.n118 output.n117 185
R21425 output.n121 output.n120 185
R21426 output.t19 output.n24 147.661
R21427 output.t18 output.n55 147.661
R21428 output.t17 output.n87 147.661
R21429 output.t16 output.n119 147.661
R21430 output.n41 output.n40 104.615
R21431 output.n40 output.n18 104.615
R21432 output.n33 output.n18 104.615
R21433 output.n33 output.n32 104.615
R21434 output.n32 output.n22 104.615
R21435 output.n25 output.n22 104.615
R21436 output.n72 output.n71 104.615
R21437 output.n71 output.n49 104.615
R21438 output.n64 output.n49 104.615
R21439 output.n64 output.n63 104.615
R21440 output.n63 output.n53 104.615
R21441 output.n56 output.n53 104.615
R21442 output.n104 output.n103 104.615
R21443 output.n103 output.n81 104.615
R21444 output.n96 output.n81 104.615
R21445 output.n96 output.n95 104.615
R21446 output.n95 output.n85 104.615
R21447 output.n88 output.n85 104.615
R21448 output.n136 output.n135 104.615
R21449 output.n135 output.n113 104.615
R21450 output.n128 output.n113 104.615
R21451 output.n128 output.n127 104.615
R21452 output.n127 output.n117 104.615
R21453 output.n120 output.n117 104.615
R21454 output.n1 output.t12 77.056
R21455 output.n14 output.t14 76.6694
R21456 output.n1 output.n0 72.7095
R21457 output.n3 output.n2 72.7095
R21458 output.n5 output.n4 72.7095
R21459 output.n7 output.n6 72.7095
R21460 output.n9 output.n8 72.7095
R21461 output.n11 output.n10 72.7095
R21462 output.n13 output.n12 72.7095
R21463 output.n25 output.t19 52.3082
R21464 output.n56 output.t18 52.3082
R21465 output.n88 output.t17 52.3082
R21466 output.n120 output.t16 52.3082
R21467 output.n26 output.n24 15.6674
R21468 output.n57 output.n55 15.6674
R21469 output.n89 output.n87 15.6674
R21470 output.n121 output.n119 15.6674
R21471 output.n27 output.n23 12.8005
R21472 output.n58 output.n54 12.8005
R21473 output.n90 output.n86 12.8005
R21474 output.n122 output.n118 12.8005
R21475 output.n31 output.n30 12.0247
R21476 output.n62 output.n61 12.0247
R21477 output.n94 output.n93 12.0247
R21478 output.n126 output.n125 12.0247
R21479 output.n34 output.n21 11.249
R21480 output.n65 output.n52 11.249
R21481 output.n97 output.n84 11.249
R21482 output.n129 output.n116 11.249
R21483 output.n35 output.n19 10.4732
R21484 output.n66 output.n50 10.4732
R21485 output.n98 output.n82 10.4732
R21486 output.n130 output.n114 10.4732
R21487 output.n39 output.n38 9.69747
R21488 output.n70 output.n69 9.69747
R21489 output.n102 output.n101 9.69747
R21490 output.n134 output.n133 9.69747
R21491 output.n45 output.n44 9.45567
R21492 output.n76 output.n75 9.45567
R21493 output.n108 output.n107 9.45567
R21494 output.n140 output.n139 9.45567
R21495 output.n44 output.n43 9.3005
R21496 output.n17 output.n16 9.3005
R21497 output.n38 output.n37 9.3005
R21498 output.n36 output.n35 9.3005
R21499 output.n21 output.n20 9.3005
R21500 output.n30 output.n29 9.3005
R21501 output.n28 output.n27 9.3005
R21502 output.n75 output.n74 9.3005
R21503 output.n48 output.n47 9.3005
R21504 output.n69 output.n68 9.3005
R21505 output.n67 output.n66 9.3005
R21506 output.n52 output.n51 9.3005
R21507 output.n61 output.n60 9.3005
R21508 output.n59 output.n58 9.3005
R21509 output.n107 output.n106 9.3005
R21510 output.n80 output.n79 9.3005
R21511 output.n101 output.n100 9.3005
R21512 output.n99 output.n98 9.3005
R21513 output.n84 output.n83 9.3005
R21514 output.n93 output.n92 9.3005
R21515 output.n91 output.n90 9.3005
R21516 output.n139 output.n138 9.3005
R21517 output.n112 output.n111 9.3005
R21518 output.n133 output.n132 9.3005
R21519 output.n131 output.n130 9.3005
R21520 output.n116 output.n115 9.3005
R21521 output.n125 output.n124 9.3005
R21522 output.n123 output.n122 9.3005
R21523 output.n42 output.n17 8.92171
R21524 output.n73 output.n48 8.92171
R21525 output.n105 output.n80 8.92171
R21526 output.n137 output.n112 8.92171
R21527 output output.n141 8.15037
R21528 output.n43 output.n15 8.14595
R21529 output.n74 output.n46 8.14595
R21530 output.n106 output.n78 8.14595
R21531 output.n138 output.n110 8.14595
R21532 output.n45 output.n15 5.81868
R21533 output.n76 output.n46 5.81868
R21534 output.n108 output.n78 5.81868
R21535 output.n140 output.n110 5.81868
R21536 output.n43 output.n42 5.04292
R21537 output.n74 output.n73 5.04292
R21538 output.n106 output.n105 5.04292
R21539 output.n138 output.n137 5.04292
R21540 output.n28 output.n24 4.38594
R21541 output.n59 output.n55 4.38594
R21542 output.n91 output.n87 4.38594
R21543 output.n123 output.n119 4.38594
R21544 output.n39 output.n17 4.26717
R21545 output.n70 output.n48 4.26717
R21546 output.n102 output.n80 4.26717
R21547 output.n134 output.n112 4.26717
R21548 output.n0 output.t3 3.9605
R21549 output.n0 output.t7 3.9605
R21550 output.n2 output.t10 3.9605
R21551 output.n2 output.t15 3.9605
R21552 output.n4 output.t0 3.9605
R21553 output.n4 output.t5 3.9605
R21554 output.n6 output.t9 3.9605
R21555 output.n6 output.t1 3.9605
R21556 output.n8 output.t4 3.9605
R21557 output.n8 output.t2 3.9605
R21558 output.n10 output.t8 3.9605
R21559 output.n10 output.t11 3.9605
R21560 output.n12 output.t13 3.9605
R21561 output.n12 output.t6 3.9605
R21562 output.n38 output.n19 3.49141
R21563 output.n69 output.n50 3.49141
R21564 output.n101 output.n82 3.49141
R21565 output.n133 output.n114 3.49141
R21566 output.n35 output.n34 2.71565
R21567 output.n66 output.n65 2.71565
R21568 output.n98 output.n97 2.71565
R21569 output.n130 output.n129 2.71565
R21570 output.n31 output.n21 1.93989
R21571 output.n62 output.n52 1.93989
R21572 output.n94 output.n84 1.93989
R21573 output.n126 output.n116 1.93989
R21574 output.n30 output.n23 1.16414
R21575 output.n61 output.n54 1.16414
R21576 output.n93 output.n86 1.16414
R21577 output.n125 output.n118 1.16414
R21578 output.n141 output.n109 0.962709
R21579 output.n109 output.n77 0.962709
R21580 output.n27 output.n26 0.388379
R21581 output.n58 output.n57 0.388379
R21582 output.n90 output.n89 0.388379
R21583 output.n122 output.n121 0.388379
R21584 output.n14 output.n13 0.387128
R21585 output.n13 output.n11 0.387128
R21586 output.n11 output.n9 0.387128
R21587 output.n9 output.n7 0.387128
R21588 output.n7 output.n5 0.387128
R21589 output.n5 output.n3 0.387128
R21590 output.n3 output.n1 0.387128
R21591 output.n44 output.n16 0.155672
R21592 output.n37 output.n16 0.155672
R21593 output.n37 output.n36 0.155672
R21594 output.n36 output.n20 0.155672
R21595 output.n29 output.n20 0.155672
R21596 output.n29 output.n28 0.155672
R21597 output.n75 output.n47 0.155672
R21598 output.n68 output.n47 0.155672
R21599 output.n68 output.n67 0.155672
R21600 output.n67 output.n51 0.155672
R21601 output.n60 output.n51 0.155672
R21602 output.n60 output.n59 0.155672
R21603 output.n107 output.n79 0.155672
R21604 output.n100 output.n79 0.155672
R21605 output.n100 output.n99 0.155672
R21606 output.n99 output.n83 0.155672
R21607 output.n92 output.n83 0.155672
R21608 output.n92 output.n91 0.155672
R21609 output.n139 output.n111 0.155672
R21610 output.n132 output.n111 0.155672
R21611 output.n132 output.n131 0.155672
R21612 output.n131 output.n115 0.155672
R21613 output.n124 output.n115 0.155672
R21614 output.n124 output.n123 0.155672
R21615 output output.n14 0.126227
R21616 minus.n46 minus.t20 252.611
R21617 minus.n9 minus.t13 252.611
R21618 minus.n78 minus.t3 243.255
R21619 minus.n72 minus.t15 231.093
R21620 minus.n35 minus.t17 231.093
R21621 minus.n77 minus.n75 224.169
R21622 minus.n77 minus.n76 223.454
R21623 minus.n38 minus.t12 187.445
R21624 minus.n65 minus.t7 187.445
R21625 minus.n59 minus.t6 187.445
R21626 minus.n42 minus.t11 187.445
R21627 minus.n44 minus.t10 187.445
R21628 minus.n47 minus.t16 187.445
R21629 minus.n10 minus.t9 187.445
R21630 minus.n7 minus.t8 187.445
R21631 minus.n5 minus.t5 187.445
R21632 minus.n22 minus.t18 187.445
R21633 minus.n28 minus.t19 187.445
R21634 minus.n1 minus.t14 187.445
R21635 minus.n48 minus.n45 161.3
R21636 minus.n50 minus.n49 161.3
R21637 minus.n52 minus.n51 161.3
R21638 minus.n53 minus.n43 161.3
R21639 minus.n55 minus.n54 161.3
R21640 minus.n57 minus.n56 161.3
R21641 minus.n58 minus.n41 161.3
R21642 minus.n61 minus.n60 161.3
R21643 minus.n62 minus.n40 161.3
R21644 minus.n64 minus.n63 161.3
R21645 minus.n66 minus.n39 161.3
R21646 minus.n68 minus.n67 161.3
R21647 minus.n70 minus.n69 161.3
R21648 minus.n71 minus.n37 161.3
R21649 minus.n73 minus.n72 161.3
R21650 minus.n36 minus.n35 161.3
R21651 minus.n34 minus.n0 161.3
R21652 minus.n33 minus.n32 161.3
R21653 minus.n31 minus.n30 161.3
R21654 minus.n29 minus.n2 161.3
R21655 minus.n27 minus.n26 161.3
R21656 minus.n25 minus.n3 161.3
R21657 minus.n24 minus.n23 161.3
R21658 minus.n21 minus.n4 161.3
R21659 minus.n20 minus.n19 161.3
R21660 minus.n18 minus.n17 161.3
R21661 minus.n16 minus.n6 161.3
R21662 minus.n15 minus.n14 161.3
R21663 minus.n13 minus.n12 161.3
R21664 minus.n11 minus.n8 161.3
R21665 minus.n67 minus.n66 56.5617
R21666 minus.n58 minus.n57 56.5617
R21667 minus.n49 minus.n48 56.5617
R21668 minus.n12 minus.n11 56.5617
R21669 minus.n21 minus.n20 56.5617
R21670 minus.n30 minus.n29 56.5617
R21671 minus.n71 minus.n70 46.3896
R21672 minus.n34 minus.n33 46.3896
R21673 minus.n46 minus.n45 42.8164
R21674 minus.n9 minus.n8 42.8164
R21675 minus.n60 minus.n40 42.5146
R21676 minus.n54 minus.n53 42.5146
R21677 minus.n17 minus.n16 42.5146
R21678 minus.n23 minus.n3 42.5146
R21679 minus.n64 minus.n40 38.6395
R21680 minus.n53 minus.n52 38.6395
R21681 minus.n16 minus.n15 38.6395
R21682 minus.n27 minus.n3 38.6395
R21683 minus.n47 minus.n46 38.2514
R21684 minus.n10 minus.n9 38.2514
R21685 minus.n74 minus.n73 31.7069
R21686 minus.n66 minus.n65 19.9199
R21687 minus.n49 minus.n44 19.9199
R21688 minus.n12 minus.n7 19.9199
R21689 minus.n29 minus.n28 19.9199
R21690 minus.n76 minus.t2 19.8005
R21691 minus.n76 minus.t0 19.8005
R21692 minus.n75 minus.t1 19.8005
R21693 minus.n75 minus.t4 19.8005
R21694 minus.n59 minus.n58 17.9525
R21695 minus.n57 minus.n42 17.9525
R21696 minus.n20 minus.n5 17.9525
R21697 minus.n22 minus.n21 17.9525
R21698 minus.n67 minus.n38 15.9852
R21699 minus.n48 minus.n47 15.9852
R21700 minus.n11 minus.n10 15.9852
R21701 minus.n30 minus.n1 15.9852
R21702 minus.n72 minus.n71 15.3369
R21703 minus.n35 minus.n34 15.3369
R21704 minus.n74 minus.n36 12.1653
R21705 minus minus.n79 11.2237
R21706 minus.n70 minus.n38 8.60764
R21707 minus.n33 minus.n1 8.60764
R21708 minus.n60 minus.n59 6.6403
R21709 minus.n54 minus.n42 6.6403
R21710 minus.n17 minus.n5 6.6403
R21711 minus.n23 minus.n22 6.6403
R21712 minus.n79 minus.n78 4.80222
R21713 minus.n65 minus.n64 4.67295
R21714 minus.n52 minus.n44 4.67295
R21715 minus.n15 minus.n7 4.67295
R21716 minus.n28 minus.n27 4.67295
R21717 minus.n79 minus.n74 0.972091
R21718 minus.n78 minus.n77 0.716017
R21719 minus.n73 minus.n37 0.189894
R21720 minus.n69 minus.n37 0.189894
R21721 minus.n69 minus.n68 0.189894
R21722 minus.n68 minus.n39 0.189894
R21723 minus.n63 minus.n39 0.189894
R21724 minus.n63 minus.n62 0.189894
R21725 minus.n62 minus.n61 0.189894
R21726 minus.n61 minus.n41 0.189894
R21727 minus.n56 minus.n41 0.189894
R21728 minus.n56 minus.n55 0.189894
R21729 minus.n55 minus.n43 0.189894
R21730 minus.n51 minus.n43 0.189894
R21731 minus.n51 minus.n50 0.189894
R21732 minus.n50 minus.n45 0.189894
R21733 minus.n13 minus.n8 0.189894
R21734 minus.n14 minus.n13 0.189894
R21735 minus.n14 minus.n6 0.189894
R21736 minus.n18 minus.n6 0.189894
R21737 minus.n19 minus.n18 0.189894
R21738 minus.n19 minus.n4 0.189894
R21739 minus.n24 minus.n4 0.189894
R21740 minus.n25 minus.n24 0.189894
R21741 minus.n26 minus.n25 0.189894
R21742 minus.n26 minus.n2 0.189894
R21743 minus.n31 minus.n2 0.189894
R21744 minus.n32 minus.n31 0.189894
R21745 minus.n32 minus.n0 0.189894
R21746 minus.n36 minus.n0 0.189894
R21747 a_n2318_8322.n9 a_n2318_8322.t7 74.6477
R21748 a_n2318_8322.t26 a_n2318_8322.n22 74.6477
R21749 a_n2318_8322.n1 a_n2318_8322.t25 74.6474
R21750 a_n2318_8322.n16 a_n2318_8322.t12 74.2899
R21751 a_n2318_8322.n6 a_n2318_8322.t15 74.2899
R21752 a_n2318_8322.n10 a_n2318_8322.t5 74.2899
R21753 a_n2318_8322.n11 a_n2318_8322.t8 74.2899
R21754 a_n2318_8322.n14 a_n2318_8322.t9 74.2899
R21755 a_n2318_8322.n22 a_n2318_8322.n21 70.6783
R21756 a_n2318_8322.n20 a_n2318_8322.n19 70.6783
R21757 a_n2318_8322.n18 a_n2318_8322.n17 70.6783
R21758 a_n2318_8322.n1 a_n2318_8322.n0 70.6783
R21759 a_n2318_8322.n3 a_n2318_8322.n2 70.6783
R21760 a_n2318_8322.n5 a_n2318_8322.n4 70.6783
R21761 a_n2318_8322.n9 a_n2318_8322.n8 70.6783
R21762 a_n2318_8322.n13 a_n2318_8322.n12 70.6783
R21763 a_n2318_8322.n16 a_n2318_8322.n15 23.4712
R21764 a_n2318_8322.n7 a_n2318_8322.t2 9.69317
R21765 a_n2318_8322.n15 a_n2318_8322.n14 6.95632
R21766 a_n2318_8322.n7 a_n2318_8322.n6 6.19447
R21767 a_n2318_8322.n15 a_n2318_8322.n7 5.3452
R21768 a_n2318_8322.n21 a_n2318_8322.t14 3.61217
R21769 a_n2318_8322.n21 a_n2318_8322.t13 3.61217
R21770 a_n2318_8322.n19 a_n2318_8322.t23 3.61217
R21771 a_n2318_8322.n19 a_n2318_8322.t18 3.61217
R21772 a_n2318_8322.n17 a_n2318_8322.t21 3.61217
R21773 a_n2318_8322.n17 a_n2318_8322.t20 3.61217
R21774 a_n2318_8322.n0 a_n2318_8322.t22 3.61217
R21775 a_n2318_8322.n0 a_n2318_8322.t19 3.61217
R21776 a_n2318_8322.n2 a_n2318_8322.t17 3.61217
R21777 a_n2318_8322.n2 a_n2318_8322.t27 3.61217
R21778 a_n2318_8322.n4 a_n2318_8322.t24 3.61217
R21779 a_n2318_8322.n4 a_n2318_8322.t16 3.61217
R21780 a_n2318_8322.n8 a_n2318_8322.t10 3.61217
R21781 a_n2318_8322.n8 a_n2318_8322.t11 3.61217
R21782 a_n2318_8322.n12 a_n2318_8322.t6 3.61217
R21783 a_n2318_8322.n12 a_n2318_8322.t4 3.61217
R21784 a_n2318_8322.n6 a_n2318_8322.n5 0.358259
R21785 a_n2318_8322.n5 a_n2318_8322.n3 0.358259
R21786 a_n2318_8322.n3 a_n2318_8322.n1 0.358259
R21787 a_n2318_8322.n14 a_n2318_8322.n13 0.358259
R21788 a_n2318_8322.n13 a_n2318_8322.n11 0.358259
R21789 a_n2318_8322.n10 a_n2318_8322.n9 0.358259
R21790 a_n2318_8322.n18 a_n2318_8322.n16 0.358259
R21791 a_n2318_8322.n20 a_n2318_8322.n18 0.358259
R21792 a_n2318_8322.n22 a_n2318_8322.n20 0.358259
R21793 a_n2318_8322.n11 a_n2318_8322.n10 0.101793
R21794 a_n2318_8322.t3 a_n2318_8322.t0 0.0788333
R21795 a_n2318_8322.t1 a_n2318_8322.t3 0.0631667
R21796 a_n2318_8322.t2 a_n2318_8322.t1 0.0471944
R21797 a_n2318_8322.t2 a_n2318_8322.t0 0.0453889
R21798 diffpairibias.n0 diffpairibias.t18 436.822
R21799 diffpairibias.n21 diffpairibias.t19 435.479
R21800 diffpairibias.n20 diffpairibias.t16 435.479
R21801 diffpairibias.n19 diffpairibias.t17 435.479
R21802 diffpairibias.n18 diffpairibias.t21 435.479
R21803 diffpairibias.n0 diffpairibias.t22 435.479
R21804 diffpairibias.n1 diffpairibias.t20 435.479
R21805 diffpairibias.n2 diffpairibias.t23 435.479
R21806 diffpairibias.n10 diffpairibias.t0 377.536
R21807 diffpairibias.n10 diffpairibias.t8 376.193
R21808 diffpairibias.n11 diffpairibias.t10 376.193
R21809 diffpairibias.n12 diffpairibias.t6 376.193
R21810 diffpairibias.n13 diffpairibias.t2 376.193
R21811 diffpairibias.n14 diffpairibias.t12 376.193
R21812 diffpairibias.n15 diffpairibias.t4 376.193
R21813 diffpairibias.n16 diffpairibias.t14 376.193
R21814 diffpairibias.n3 diffpairibias.t1 113.368
R21815 diffpairibias.n3 diffpairibias.t9 112.698
R21816 diffpairibias.n4 diffpairibias.t11 112.698
R21817 diffpairibias.n5 diffpairibias.t7 112.698
R21818 diffpairibias.n6 diffpairibias.t3 112.698
R21819 diffpairibias.n7 diffpairibias.t13 112.698
R21820 diffpairibias.n8 diffpairibias.t5 112.698
R21821 diffpairibias.n9 diffpairibias.t15 112.698
R21822 diffpairibias.n17 diffpairibias.n16 4.77242
R21823 diffpairibias.n17 diffpairibias.n9 4.30807
R21824 diffpairibias.n18 diffpairibias.n17 4.13945
R21825 diffpairibias.n16 diffpairibias.n15 1.34352
R21826 diffpairibias.n15 diffpairibias.n14 1.34352
R21827 diffpairibias.n14 diffpairibias.n13 1.34352
R21828 diffpairibias.n13 diffpairibias.n12 1.34352
R21829 diffpairibias.n12 diffpairibias.n11 1.34352
R21830 diffpairibias.n11 diffpairibias.n10 1.34352
R21831 diffpairibias.n2 diffpairibias.n1 1.34352
R21832 diffpairibias.n1 diffpairibias.n0 1.34352
R21833 diffpairibias.n19 diffpairibias.n18 1.34352
R21834 diffpairibias.n20 diffpairibias.n19 1.34352
R21835 diffpairibias.n21 diffpairibias.n20 1.34352
R21836 diffpairibias.n22 diffpairibias.n21 0.862419
R21837 diffpairibias diffpairibias.n22 0.684875
R21838 diffpairibias.n9 diffpairibias.n8 0.672012
R21839 diffpairibias.n8 diffpairibias.n7 0.672012
R21840 diffpairibias.n7 diffpairibias.n6 0.672012
R21841 diffpairibias.n6 diffpairibias.n5 0.672012
R21842 diffpairibias.n5 diffpairibias.n4 0.672012
R21843 diffpairibias.n4 diffpairibias.n3 0.672012
R21844 diffpairibias.n22 diffpairibias.n2 0.190907
C0 CSoutput outputibias 0.032386f
C1 vdd CSoutput 0.116834p
C2 minus diffpairibias 3.46e-19
C3 commonsourceibias output 0.006808f
C4 CSoutput minus 2.50162f
C5 vdd plus 0.085153f
C6 commonsourceibias outputibias 0.003832f
C7 plus diffpairibias 2.47e-19
C8 vdd commonsourceibias 0.004218f
C9 CSoutput plus 0.837031f
C10 commonsourceibias diffpairibias 0.052851f
C11 CSoutput commonsourceibias 29.0223f
C12 minus plus 8.791639f
C13 minus commonsourceibias 0.323289f
C14 plus commonsourceibias 0.277692f
C15 output outputibias 2.34152f
C16 vdd output 7.23429f
C17 CSoutput output 6.13571f
C18 diffpairibias gnd 48.96854f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.118807p
C22 plus gnd 31.831968f
C23 minus gnd 25.730589f
C24 CSoutput gnd 88.0566f
C25 vdd gnd 0.442491p
C26 diffpairibias.t18 gnd 0.087401f
C27 diffpairibias.t22 gnd 0.087239f
C28 diffpairibias.n0 gnd 0.102784f
C29 diffpairibias.t20 gnd 0.087239f
C30 diffpairibias.n1 gnd 0.050171f
C31 diffpairibias.t23 gnd 0.087239f
C32 diffpairibias.n2 gnd 0.039841f
C33 diffpairibias.t1 gnd 0.083757f
C34 diffpairibias.t9 gnd 0.083392f
C35 diffpairibias.n3 gnd 0.131682f
C36 diffpairibias.t11 gnd 0.083392f
C37 diffpairibias.n4 gnd 0.07027f
C38 diffpairibias.t7 gnd 0.083392f
C39 diffpairibias.n5 gnd 0.07027f
C40 diffpairibias.t3 gnd 0.083392f
C41 diffpairibias.n6 gnd 0.07027f
C42 diffpairibias.t13 gnd 0.083392f
C43 diffpairibias.n7 gnd 0.07027f
C44 diffpairibias.t5 gnd 0.083392f
C45 diffpairibias.n8 gnd 0.07027f
C46 diffpairibias.t15 gnd 0.083392f
C47 diffpairibias.n9 gnd 0.099771f
C48 diffpairibias.t0 gnd 0.08427f
C49 diffpairibias.t8 gnd 0.084123f
C50 diffpairibias.n10 gnd 0.091784f
C51 diffpairibias.t10 gnd 0.084123f
C52 diffpairibias.n11 gnd 0.050681f
C53 diffpairibias.t6 gnd 0.084123f
C54 diffpairibias.n12 gnd 0.050681f
C55 diffpairibias.t2 gnd 0.084123f
C56 diffpairibias.n13 gnd 0.050681f
C57 diffpairibias.t12 gnd 0.084123f
C58 diffpairibias.n14 gnd 0.050681f
C59 diffpairibias.t4 gnd 0.084123f
C60 diffpairibias.n15 gnd 0.050681f
C61 diffpairibias.t14 gnd 0.084123f
C62 diffpairibias.n16 gnd 0.059977f
C63 diffpairibias.n17 gnd 0.226448f
C64 diffpairibias.t21 gnd 0.087239f
C65 diffpairibias.n18 gnd 0.050181f
C66 diffpairibias.t17 gnd 0.087239f
C67 diffpairibias.n19 gnd 0.050171f
C68 diffpairibias.t16 gnd 0.087239f
C69 diffpairibias.n20 gnd 0.050171f
C70 diffpairibias.t19 gnd 0.087239f
C71 diffpairibias.n21 gnd 0.045859f
C72 diffpairibias.n22 gnd 0.046268f
C73 a_n2318_8322.t0 gnd 39.618103f
C74 a_n2318_8322.t2 gnd 27.7211f
C75 a_n2318_8322.t3 gnd 19.739399f
C76 a_n2318_8322.t1 gnd 39.618103f
C77 a_n2318_8322.t25 gnd 0.897207f
C78 a_n2318_8322.t22 gnd 0.09582f
C79 a_n2318_8322.t19 gnd 0.09582f
C80 a_n2318_8322.n0 gnd 0.674956f
C81 a_n2318_8322.n1 gnd 0.754166f
C82 a_n2318_8322.t17 gnd 0.09582f
C83 a_n2318_8322.t27 gnd 0.09582f
C84 a_n2318_8322.n2 gnd 0.674956f
C85 a_n2318_8322.n3 gnd 0.383181f
C86 a_n2318_8322.t24 gnd 0.09582f
C87 a_n2318_8322.t16 gnd 0.09582f
C88 a_n2318_8322.n4 gnd 0.674956f
C89 a_n2318_8322.n5 gnd 0.383181f
C90 a_n2318_8322.t15 gnd 0.895423f
C91 a_n2318_8322.n6 gnd 0.881475f
C92 a_n2318_8322.n7 gnd 3.12946f
C93 a_n2318_8322.t7 gnd 0.89721f
C94 a_n2318_8322.t10 gnd 0.09582f
C95 a_n2318_8322.t11 gnd 0.09582f
C96 a_n2318_8322.n8 gnd 0.674956f
C97 a_n2318_8322.n9 gnd 0.754164f
C98 a_n2318_8322.t5 gnd 0.895423f
C99 a_n2318_8322.n10 gnd 0.379506f
C100 a_n2318_8322.t8 gnd 0.895423f
C101 a_n2318_8322.n11 gnd 0.379506f
C102 a_n2318_8322.t6 gnd 0.09582f
C103 a_n2318_8322.t4 gnd 0.09582f
C104 a_n2318_8322.n12 gnd 0.674956f
C105 a_n2318_8322.n13 gnd 0.383181f
C106 a_n2318_8322.t9 gnd 0.895423f
C107 a_n2318_8322.n14 gnd 1.07467f
C108 a_n2318_8322.n15 gnd 1.82686f
C109 a_n2318_8322.t12 gnd 0.895423f
C110 a_n2318_8322.n16 gnd 1.5519f
C111 a_n2318_8322.t21 gnd 0.09582f
C112 a_n2318_8322.t20 gnd 0.09582f
C113 a_n2318_8322.n17 gnd 0.674956f
C114 a_n2318_8322.n18 gnd 0.383181f
C115 a_n2318_8322.t23 gnd 0.09582f
C116 a_n2318_8322.t18 gnd 0.09582f
C117 a_n2318_8322.n19 gnd 0.674956f
C118 a_n2318_8322.n20 gnd 0.383181f
C119 a_n2318_8322.t14 gnd 0.09582f
C120 a_n2318_8322.t13 gnd 0.09582f
C121 a_n2318_8322.n21 gnd 0.674956f
C122 a_n2318_8322.n22 gnd 0.754164f
C123 a_n2318_8322.t26 gnd 0.89721f
C124 minus.n0 gnd 0.03064f
C125 minus.t14 gnd 0.515204f
C126 minus.n1 gnd 0.208372f
C127 minus.n2 gnd 0.03064f
C128 minus.t19 gnd 0.515204f
C129 minus.n3 gnd 0.024903f
C130 minus.n4 gnd 0.03064f
C131 minus.t18 gnd 0.515204f
C132 minus.t5 gnd 0.515204f
C133 minus.n5 gnd 0.208372f
C134 minus.n6 gnd 0.03064f
C135 minus.t8 gnd 0.515204f
C136 minus.n7 gnd 0.208372f
C137 minus.n8 gnd 0.131525f
C138 minus.t9 gnd 0.515204f
C139 minus.t13 gnd 0.578439f
C140 minus.n9 gnd 0.241768f
C141 minus.n10 gnd 0.240637f
C142 minus.n11 gnd 0.038113f
C143 minus.n12 gnd 0.03582f
C144 minus.n13 gnd 0.03064f
C145 minus.n14 gnd 0.03064f
C146 minus.n15 gnd 0.038381f
C147 minus.n16 gnd 0.024903f
C148 minus.n17 gnd 0.039417f
C149 minus.n18 gnd 0.03064f
C150 minus.n19 gnd 0.03064f
C151 minus.n20 gnd 0.036966f
C152 minus.n21 gnd 0.036966f
C153 minus.n22 gnd 0.208372f
C154 minus.n23 gnd 0.039417f
C155 minus.n24 gnd 0.03064f
C156 minus.n25 gnd 0.03064f
C157 minus.n26 gnd 0.03064f
C158 minus.n27 gnd 0.038381f
C159 minus.n28 gnd 0.208372f
C160 minus.n29 gnd 0.03582f
C161 minus.n30 gnd 0.038113f
C162 minus.n31 gnd 0.03064f
C163 minus.n32 gnd 0.03064f
C164 minus.n33 gnd 0.039904f
C165 minus.n34 gnd 0.01269f
C166 minus.t17 gnd 0.557193f
C167 minus.n35 gnd 0.242015f
C168 minus.n36 gnd 0.360024f
C169 minus.n37 gnd 0.03064f
C170 minus.t15 gnd 0.557193f
C171 minus.t12 gnd 0.515204f
C172 minus.n38 gnd 0.208372f
C173 minus.n39 gnd 0.03064f
C174 minus.t7 gnd 0.515204f
C175 minus.n40 gnd 0.024903f
C176 minus.n41 gnd 0.03064f
C177 minus.t6 gnd 0.515204f
C178 minus.t11 gnd 0.515204f
C179 minus.n42 gnd 0.208372f
C180 minus.n43 gnd 0.03064f
C181 minus.t10 gnd 0.515204f
C182 minus.n44 gnd 0.208372f
C183 minus.n45 gnd 0.131525f
C184 minus.t16 gnd 0.515204f
C185 minus.t20 gnd 0.578439f
C186 minus.n46 gnd 0.241768f
C187 minus.n47 gnd 0.240637f
C188 minus.n48 gnd 0.038113f
C189 minus.n49 gnd 0.03582f
C190 minus.n50 gnd 0.03064f
C191 minus.n51 gnd 0.03064f
C192 minus.n52 gnd 0.038381f
C193 minus.n53 gnd 0.024903f
C194 minus.n54 gnd 0.039417f
C195 minus.n55 gnd 0.03064f
C196 minus.n56 gnd 0.03064f
C197 minus.n57 gnd 0.036966f
C198 minus.n58 gnd 0.036966f
C199 minus.n59 gnd 0.208372f
C200 minus.n60 gnd 0.039417f
C201 minus.n61 gnd 0.03064f
C202 minus.n62 gnd 0.03064f
C203 minus.n63 gnd 0.03064f
C204 minus.n64 gnd 0.038381f
C205 minus.n65 gnd 0.208372f
C206 minus.n66 gnd 0.03582f
C207 minus.n67 gnd 0.038113f
C208 minus.n68 gnd 0.03064f
C209 minus.n69 gnd 0.03064f
C210 minus.n70 gnd 0.039904f
C211 minus.n71 gnd 0.01269f
C212 minus.n72 gnd 0.242015f
C213 minus.n73 gnd 0.954724f
C214 minus.n74 gnd 1.43503f
C215 minus.t1 gnd 0.009445f
C216 minus.t4 gnd 0.009445f
C217 minus.n75 gnd 0.031059f
C218 minus.t2 gnd 0.009445f
C219 minus.t0 gnd 0.009445f
C220 minus.n76 gnd 0.030633f
C221 minus.n77 gnd 0.261439f
C222 minus.t3 gnd 0.052572f
C223 minus.n78 gnd 0.142665f
C224 minus.n79 gnd 1.72784f
C225 output.t12 gnd 0.464308f
C226 output.t3 gnd 0.044422f
C227 output.t7 gnd 0.044422f
C228 output.n0 gnd 0.364624f
C229 output.n1 gnd 0.614102f
C230 output.t10 gnd 0.044422f
C231 output.t15 gnd 0.044422f
C232 output.n2 gnd 0.364624f
C233 output.n3 gnd 0.350265f
C234 output.t0 gnd 0.044422f
C235 output.t5 gnd 0.044422f
C236 output.n4 gnd 0.364624f
C237 output.n5 gnd 0.350265f
C238 output.t9 gnd 0.044422f
C239 output.t1 gnd 0.044422f
C240 output.n6 gnd 0.364624f
C241 output.n7 gnd 0.350265f
C242 output.t4 gnd 0.044422f
C243 output.t2 gnd 0.044422f
C244 output.n8 gnd 0.364624f
C245 output.n9 gnd 0.350265f
C246 output.t8 gnd 0.044422f
C247 output.t11 gnd 0.044422f
C248 output.n10 gnd 0.364624f
C249 output.n11 gnd 0.350265f
C250 output.t13 gnd 0.044422f
C251 output.t6 gnd 0.044422f
C252 output.n12 gnd 0.364624f
C253 output.n13 gnd 0.350265f
C254 output.t14 gnd 0.462979f
C255 output.n14 gnd 0.28994f
C256 output.n15 gnd 0.015803f
C257 output.n16 gnd 0.011243f
C258 output.n17 gnd 0.006041f
C259 output.n18 gnd 0.01428f
C260 output.n19 gnd 0.006397f
C261 output.n20 gnd 0.011243f
C262 output.n21 gnd 0.006041f
C263 output.n22 gnd 0.01428f
C264 output.n23 gnd 0.006397f
C265 output.n24 gnd 0.048111f
C266 output.t19 gnd 0.023274f
C267 output.n25 gnd 0.01071f
C268 output.n26 gnd 0.008435f
C269 output.n27 gnd 0.006041f
C270 output.n28 gnd 0.267512f
C271 output.n29 gnd 0.011243f
C272 output.n30 gnd 0.006041f
C273 output.n31 gnd 0.006397f
C274 output.n32 gnd 0.01428f
C275 output.n33 gnd 0.01428f
C276 output.n34 gnd 0.006397f
C277 output.n35 gnd 0.006041f
C278 output.n36 gnd 0.011243f
C279 output.n37 gnd 0.011243f
C280 output.n38 gnd 0.006041f
C281 output.n39 gnd 0.006397f
C282 output.n40 gnd 0.01428f
C283 output.n41 gnd 0.030913f
C284 output.n42 gnd 0.006397f
C285 output.n43 gnd 0.006041f
C286 output.n44 gnd 0.025987f
C287 output.n45 gnd 0.097665f
C288 output.n46 gnd 0.015803f
C289 output.n47 gnd 0.011243f
C290 output.n48 gnd 0.006041f
C291 output.n49 gnd 0.01428f
C292 output.n50 gnd 0.006397f
C293 output.n51 gnd 0.011243f
C294 output.n52 gnd 0.006041f
C295 output.n53 gnd 0.01428f
C296 output.n54 gnd 0.006397f
C297 output.n55 gnd 0.048111f
C298 output.t18 gnd 0.023274f
C299 output.n56 gnd 0.01071f
C300 output.n57 gnd 0.008435f
C301 output.n58 gnd 0.006041f
C302 output.n59 gnd 0.267512f
C303 output.n60 gnd 0.011243f
C304 output.n61 gnd 0.006041f
C305 output.n62 gnd 0.006397f
C306 output.n63 gnd 0.01428f
C307 output.n64 gnd 0.01428f
C308 output.n65 gnd 0.006397f
C309 output.n66 gnd 0.006041f
C310 output.n67 gnd 0.011243f
C311 output.n68 gnd 0.011243f
C312 output.n69 gnd 0.006041f
C313 output.n70 gnd 0.006397f
C314 output.n71 gnd 0.01428f
C315 output.n72 gnd 0.030913f
C316 output.n73 gnd 0.006397f
C317 output.n74 gnd 0.006041f
C318 output.n75 gnd 0.025987f
C319 output.n76 gnd 0.09306f
C320 output.n77 gnd 1.65264f
C321 output.n78 gnd 0.015803f
C322 output.n79 gnd 0.011243f
C323 output.n80 gnd 0.006041f
C324 output.n81 gnd 0.01428f
C325 output.n82 gnd 0.006397f
C326 output.n83 gnd 0.011243f
C327 output.n84 gnd 0.006041f
C328 output.n85 gnd 0.01428f
C329 output.n86 gnd 0.006397f
C330 output.n87 gnd 0.048111f
C331 output.t17 gnd 0.023274f
C332 output.n88 gnd 0.01071f
C333 output.n89 gnd 0.008435f
C334 output.n90 gnd 0.006041f
C335 output.n91 gnd 0.267512f
C336 output.n92 gnd 0.011243f
C337 output.n93 gnd 0.006041f
C338 output.n94 gnd 0.006397f
C339 output.n95 gnd 0.01428f
C340 output.n96 gnd 0.01428f
C341 output.n97 gnd 0.006397f
C342 output.n98 gnd 0.006041f
C343 output.n99 gnd 0.011243f
C344 output.n100 gnd 0.011243f
C345 output.n101 gnd 0.006041f
C346 output.n102 gnd 0.006397f
C347 output.n103 gnd 0.01428f
C348 output.n104 gnd 0.030913f
C349 output.n105 gnd 0.006397f
C350 output.n106 gnd 0.006041f
C351 output.n107 gnd 0.025987f
C352 output.n108 gnd 0.09306f
C353 output.n109 gnd 0.713089f
C354 output.n110 gnd 0.015803f
C355 output.n111 gnd 0.011243f
C356 output.n112 gnd 0.006041f
C357 output.n113 gnd 0.01428f
C358 output.n114 gnd 0.006397f
C359 output.n115 gnd 0.011243f
C360 output.n116 gnd 0.006041f
C361 output.n117 gnd 0.01428f
C362 output.n118 gnd 0.006397f
C363 output.n119 gnd 0.048111f
C364 output.t16 gnd 0.023274f
C365 output.n120 gnd 0.01071f
C366 output.n121 gnd 0.008435f
C367 output.n122 gnd 0.006041f
C368 output.n123 gnd 0.267512f
C369 output.n124 gnd 0.011243f
C370 output.n125 gnd 0.006041f
C371 output.n126 gnd 0.006397f
C372 output.n127 gnd 0.01428f
C373 output.n128 gnd 0.01428f
C374 output.n129 gnd 0.006397f
C375 output.n130 gnd 0.006041f
C376 output.n131 gnd 0.011243f
C377 output.n132 gnd 0.011243f
C378 output.n133 gnd 0.006041f
C379 output.n134 gnd 0.006397f
C380 output.n135 gnd 0.01428f
C381 output.n136 gnd 0.030913f
C382 output.n137 gnd 0.006397f
C383 output.n138 gnd 0.006041f
C384 output.n139 gnd 0.025987f
C385 output.n140 gnd 0.09306f
C386 output.n141 gnd 1.67353f
C387 outputibias.t9 gnd 0.11477f
C388 outputibias.t8 gnd 0.115567f
C389 outputibias.n0 gnd 0.130108f
C390 outputibias.n1 gnd 0.001372f
C391 outputibias.n2 gnd 9.76e-19
C392 outputibias.n3 gnd 5.24e-19
C393 outputibias.n4 gnd 0.001239f
C394 outputibias.n5 gnd 5.55e-19
C395 outputibias.n6 gnd 9.76e-19
C396 outputibias.n7 gnd 5.24e-19
C397 outputibias.n8 gnd 0.001239f
C398 outputibias.n9 gnd 5.55e-19
C399 outputibias.n10 gnd 0.004176f
C400 outputibias.t5 gnd 0.00202f
C401 outputibias.n11 gnd 9.3e-19
C402 outputibias.n12 gnd 7.32e-19
C403 outputibias.n13 gnd 5.24e-19
C404 outputibias.n14 gnd 0.02322f
C405 outputibias.n15 gnd 9.76e-19
C406 outputibias.n16 gnd 5.24e-19
C407 outputibias.n17 gnd 5.55e-19
C408 outputibias.n18 gnd 0.001239f
C409 outputibias.n19 gnd 0.001239f
C410 outputibias.n20 gnd 5.55e-19
C411 outputibias.n21 gnd 5.24e-19
C412 outputibias.n22 gnd 9.76e-19
C413 outputibias.n23 gnd 9.76e-19
C414 outputibias.n24 gnd 5.24e-19
C415 outputibias.n25 gnd 5.55e-19
C416 outputibias.n26 gnd 0.001239f
C417 outputibias.n27 gnd 0.002683f
C418 outputibias.n28 gnd 5.55e-19
C419 outputibias.n29 gnd 5.24e-19
C420 outputibias.n30 gnd 0.002256f
C421 outputibias.n31 gnd 0.005781f
C422 outputibias.n32 gnd 0.001372f
C423 outputibias.n33 gnd 9.76e-19
C424 outputibias.n34 gnd 5.24e-19
C425 outputibias.n35 gnd 0.001239f
C426 outputibias.n36 gnd 5.55e-19
C427 outputibias.n37 gnd 9.76e-19
C428 outputibias.n38 gnd 5.24e-19
C429 outputibias.n39 gnd 0.001239f
C430 outputibias.n40 gnd 5.55e-19
C431 outputibias.n41 gnd 0.004176f
C432 outputibias.t7 gnd 0.00202f
C433 outputibias.n42 gnd 9.3e-19
C434 outputibias.n43 gnd 7.32e-19
C435 outputibias.n44 gnd 5.24e-19
C436 outputibias.n45 gnd 0.02322f
C437 outputibias.n46 gnd 9.76e-19
C438 outputibias.n47 gnd 5.24e-19
C439 outputibias.n48 gnd 5.55e-19
C440 outputibias.n49 gnd 0.001239f
C441 outputibias.n50 gnd 0.001239f
C442 outputibias.n51 gnd 5.55e-19
C443 outputibias.n52 gnd 5.24e-19
C444 outputibias.n53 gnd 9.76e-19
C445 outputibias.n54 gnd 9.76e-19
C446 outputibias.n55 gnd 5.24e-19
C447 outputibias.n56 gnd 5.55e-19
C448 outputibias.n57 gnd 0.001239f
C449 outputibias.n58 gnd 0.002683f
C450 outputibias.n59 gnd 5.55e-19
C451 outputibias.n60 gnd 5.24e-19
C452 outputibias.n61 gnd 0.002256f
C453 outputibias.n62 gnd 0.005197f
C454 outputibias.n63 gnd 0.121892f
C455 outputibias.n64 gnd 0.001372f
C456 outputibias.n65 gnd 9.76e-19
C457 outputibias.n66 gnd 5.24e-19
C458 outputibias.n67 gnd 0.001239f
C459 outputibias.n68 gnd 5.55e-19
C460 outputibias.n69 gnd 9.76e-19
C461 outputibias.n70 gnd 5.24e-19
C462 outputibias.n71 gnd 0.001239f
C463 outputibias.n72 gnd 5.55e-19
C464 outputibias.n73 gnd 0.004176f
C465 outputibias.t1 gnd 0.00202f
C466 outputibias.n74 gnd 9.3e-19
C467 outputibias.n75 gnd 7.32e-19
C468 outputibias.n76 gnd 5.24e-19
C469 outputibias.n77 gnd 0.02322f
C470 outputibias.n78 gnd 9.76e-19
C471 outputibias.n79 gnd 5.24e-19
C472 outputibias.n80 gnd 5.55e-19
C473 outputibias.n81 gnd 0.001239f
C474 outputibias.n82 gnd 0.001239f
C475 outputibias.n83 gnd 5.55e-19
C476 outputibias.n84 gnd 5.24e-19
C477 outputibias.n85 gnd 9.76e-19
C478 outputibias.n86 gnd 9.76e-19
C479 outputibias.n87 gnd 5.24e-19
C480 outputibias.n88 gnd 5.55e-19
C481 outputibias.n89 gnd 0.001239f
C482 outputibias.n90 gnd 0.002683f
C483 outputibias.n91 gnd 5.55e-19
C484 outputibias.n92 gnd 5.24e-19
C485 outputibias.n93 gnd 0.002256f
C486 outputibias.n94 gnd 0.005197f
C487 outputibias.n95 gnd 0.064513f
C488 outputibias.n96 gnd 0.001372f
C489 outputibias.n97 gnd 9.76e-19
C490 outputibias.n98 gnd 5.24e-19
C491 outputibias.n99 gnd 0.001239f
C492 outputibias.n100 gnd 5.55e-19
C493 outputibias.n101 gnd 9.76e-19
C494 outputibias.n102 gnd 5.24e-19
C495 outputibias.n103 gnd 0.001239f
C496 outputibias.n104 gnd 5.55e-19
C497 outputibias.n105 gnd 0.004176f
C498 outputibias.t3 gnd 0.00202f
C499 outputibias.n106 gnd 9.3e-19
C500 outputibias.n107 gnd 7.32e-19
C501 outputibias.n108 gnd 5.24e-19
C502 outputibias.n109 gnd 0.02322f
C503 outputibias.n110 gnd 9.76e-19
C504 outputibias.n111 gnd 5.24e-19
C505 outputibias.n112 gnd 5.55e-19
C506 outputibias.n113 gnd 0.001239f
C507 outputibias.n114 gnd 0.001239f
C508 outputibias.n115 gnd 5.55e-19
C509 outputibias.n116 gnd 5.24e-19
C510 outputibias.n117 gnd 9.76e-19
C511 outputibias.n118 gnd 9.76e-19
C512 outputibias.n119 gnd 5.24e-19
C513 outputibias.n120 gnd 5.55e-19
C514 outputibias.n121 gnd 0.001239f
C515 outputibias.n122 gnd 0.002683f
C516 outputibias.n123 gnd 5.55e-19
C517 outputibias.n124 gnd 5.24e-19
C518 outputibias.n125 gnd 0.002256f
C519 outputibias.n126 gnd 0.005197f
C520 outputibias.n127 gnd 0.084814f
C521 outputibias.t2 gnd 0.108319f
C522 outputibias.t0 gnd 0.108319f
C523 outputibias.t6 gnd 0.108319f
C524 outputibias.t4 gnd 0.109238f
C525 outputibias.n128 gnd 0.134674f
C526 outputibias.n129 gnd 0.07244f
C527 outputibias.n130 gnd 0.079818f
C528 outputibias.n131 gnd 0.164901f
C529 outputibias.t11 gnd 0.11477f
C530 outputibias.n132 gnd 0.067481f
C531 outputibias.t10 gnd 0.11477f
C532 outputibias.n133 gnd 0.065115f
C533 outputibias.n134 gnd 0.029159f
C534 a_n2903_n3924.n0 gnd 1.45586f
C535 a_n2903_n3924.t22 gnd 0.088483f
C536 a_n2903_n3924.t31 gnd 0.919619f
C537 a_n2903_n3924.n1 gnd 0.347657f
C538 a_n2903_n3924.t2 gnd 1.14306f
C539 a_n2903_n3924.n2 gnd 1.19083f
C540 a_n2903_n3924.t6 gnd 0.919619f
C541 a_n2903_n3924.n3 gnd 0.347657f
C542 a_n2903_n3924.t8 gnd 0.088483f
C543 a_n2903_n3924.t10 gnd 0.088483f
C544 a_n2903_n3924.n4 gnd 0.722655f
C545 a_n2903_n3924.n5 gnd 0.364177f
C546 a_n2903_n3924.t19 gnd 0.088483f
C547 a_n2903_n3924.t7 gnd 0.088483f
C548 a_n2903_n3924.n6 gnd 0.722655f
C549 a_n2903_n3924.n7 gnd 0.364177f
C550 a_n2903_n3924.t14 gnd 0.088483f
C551 a_n2903_n3924.t17 gnd 0.088483f
C552 a_n2903_n3924.n8 gnd 0.722655f
C553 a_n2903_n3924.n9 gnd 0.364177f
C554 a_n2903_n3924.t11 gnd 0.919619f
C555 a_n2903_n3924.n10 gnd 0.860834f
C556 a_n2903_n3924.t37 gnd 1.14419f
C557 a_n2903_n3924.t38 gnd 1.14261f
C558 a_n2903_n3924.n11 gnd 0.745791f
C559 a_n2903_n3924.t36 gnd 1.14261f
C560 a_n2903_n3924.n12 gnd 0.804757f
C561 a_n2903_n3924.t1 gnd 1.14261f
C562 a_n2903_n3924.n13 gnd 0.804757f
C563 a_n2903_n3924.t0 gnd 1.14261f
C564 a_n2903_n3924.n14 gnd 0.804757f
C565 a_n2903_n3924.t3 gnd 1.14261f
C566 a_n2903_n3924.n15 gnd 0.804757f
C567 a_n2903_n3924.t39 gnd 1.14261f
C568 a_n2903_n3924.n16 gnd 0.834168f
C569 a_n2903_n3924.t33 gnd 0.919616f
C570 a_n2903_n3924.n17 gnd 0.571219f
C571 a_n2903_n3924.t34 gnd 0.088483f
C572 a_n2903_n3924.t24 gnd 0.088483f
C573 a_n2903_n3924.n18 gnd 0.722654f
C574 a_n2903_n3924.n19 gnd 0.364178f
C575 a_n2903_n3924.t25 gnd 0.088483f
C576 a_n2903_n3924.t20 gnd 0.088483f
C577 a_n2903_n3924.n20 gnd 0.722654f
C578 a_n2903_n3924.n21 gnd 0.364178f
C579 a_n2903_n3924.t21 gnd 0.088483f
C580 a_n2903_n3924.t32 gnd 0.088483f
C581 a_n2903_n3924.n22 gnd 0.722654f
C582 a_n2903_n3924.n23 gnd 0.364178f
C583 a_n2903_n3924.t29 gnd 0.919616f
C584 a_n2903_n3924.n24 gnd 0.347661f
C585 a_n2903_n3924.t13 gnd 0.919616f
C586 a_n2903_n3924.n25 gnd 0.347661f
C587 a_n2903_n3924.t15 gnd 0.088483f
C588 a_n2903_n3924.t16 gnd 0.088483f
C589 a_n2903_n3924.n26 gnd 0.722654f
C590 a_n2903_n3924.n27 gnd 0.364178f
C591 a_n2903_n3924.t18 gnd 0.088483f
C592 a_n2903_n3924.t5 gnd 0.088483f
C593 a_n2903_n3924.n28 gnd 0.722654f
C594 a_n2903_n3924.n29 gnd 0.364178f
C595 a_n2903_n3924.t4 gnd 0.088483f
C596 a_n2903_n3924.t12 gnd 0.088483f
C597 a_n2903_n3924.n30 gnd 0.722654f
C598 a_n2903_n3924.n31 gnd 0.364178f
C599 a_n2903_n3924.t9 gnd 0.919616f
C600 a_n2903_n3924.n32 gnd 0.571219f
C601 a_n2903_n3924.n33 gnd 0.834168f
C602 a_n2903_n3924.t28 gnd 0.919616f
C603 a_n2903_n3924.n34 gnd 0.860837f
C604 a_n2903_n3924.t26 gnd 0.088483f
C605 a_n2903_n3924.t30 gnd 0.088483f
C606 a_n2903_n3924.n35 gnd 0.722655f
C607 a_n2903_n3924.n36 gnd 0.364177f
C608 a_n2903_n3924.t23 gnd 0.088483f
C609 a_n2903_n3924.t27 gnd 0.088483f
C610 a_n2903_n3924.n37 gnd 0.722655f
C611 a_n2903_n3924.n38 gnd 0.364177f
C612 a_n2903_n3924.n39 gnd 0.364176f
C613 a_n2903_n3924.n40 gnd 0.722656f
C614 a_n2903_n3924.t35 gnd 0.088483f
C615 plus.n0 gnd 0.022489f
C616 plus.t7 gnd 0.408961f
C617 plus.t6 gnd 0.378142f
C618 plus.n1 gnd 0.152937f
C619 plus.n2 gnd 0.022489f
C620 plus.t16 gnd 0.378142f
C621 plus.n3 gnd 0.018278f
C622 plus.n4 gnd 0.022489f
C623 plus.t15 gnd 0.378142f
C624 plus.t20 gnd 0.378142f
C625 plus.n5 gnd 0.152937f
C626 plus.n6 gnd 0.022489f
C627 plus.t19 gnd 0.378142f
C628 plus.n7 gnd 0.152937f
C629 plus.n8 gnd 0.096534f
C630 plus.t8 gnd 0.378142f
C631 plus.t11 gnd 0.424554f
C632 plus.n9 gnd 0.17745f
C633 plus.n10 gnd 0.176619f
C634 plus.n11 gnd 0.027974f
C635 plus.n12 gnd 0.02629f
C636 plus.n13 gnd 0.022489f
C637 plus.n14 gnd 0.022489f
C638 plus.n15 gnd 0.028171f
C639 plus.n16 gnd 0.018278f
C640 plus.n17 gnd 0.028931f
C641 plus.n18 gnd 0.022489f
C642 plus.n19 gnd 0.022489f
C643 plus.n20 gnd 0.027132f
C644 plus.n21 gnd 0.027132f
C645 plus.n22 gnd 0.152937f
C646 plus.n23 gnd 0.028931f
C647 plus.n24 gnd 0.022489f
C648 plus.n25 gnd 0.022489f
C649 plus.n26 gnd 0.022489f
C650 plus.n27 gnd 0.028171f
C651 plus.n28 gnd 0.152937f
C652 plus.n29 gnd 0.02629f
C653 plus.n30 gnd 0.027974f
C654 plus.n31 gnd 0.022489f
C655 plus.n32 gnd 0.022489f
C656 plus.n33 gnd 0.029288f
C657 plus.n34 gnd 0.009314f
C658 plus.n35 gnd 0.17763f
C659 plus.n36 gnd 0.258461f
C660 plus.n37 gnd 0.022489f
C661 plus.t10 gnd 0.378142f
C662 plus.n38 gnd 0.152937f
C663 plus.n39 gnd 0.022489f
C664 plus.t14 gnd 0.378142f
C665 plus.n40 gnd 0.018278f
C666 plus.n41 gnd 0.022489f
C667 plus.t13 gnd 0.378142f
C668 plus.t17 gnd 0.378142f
C669 plus.n42 gnd 0.152937f
C670 plus.n43 gnd 0.022489f
C671 plus.t18 gnd 0.378142f
C672 plus.n44 gnd 0.152937f
C673 plus.n45 gnd 0.096534f
C674 plus.t5 gnd 0.378142f
C675 plus.t9 gnd 0.424554f
C676 plus.n46 gnd 0.17745f
C677 plus.n47 gnd 0.176619f
C678 plus.n48 gnd 0.027974f
C679 plus.n49 gnd 0.02629f
C680 plus.n50 gnd 0.022489f
C681 plus.n51 gnd 0.022489f
C682 plus.n52 gnd 0.028171f
C683 plus.n53 gnd 0.018278f
C684 plus.n54 gnd 0.028931f
C685 plus.n55 gnd 0.022489f
C686 plus.n56 gnd 0.022489f
C687 plus.n57 gnd 0.027132f
C688 plus.n58 gnd 0.027132f
C689 plus.n59 gnd 0.152937f
C690 plus.n60 gnd 0.028931f
C691 plus.n61 gnd 0.022489f
C692 plus.n62 gnd 0.022489f
C693 plus.n63 gnd 0.022489f
C694 plus.n64 gnd 0.028171f
C695 plus.n65 gnd 0.152937f
C696 plus.n66 gnd 0.02629f
C697 plus.n67 gnd 0.027974f
C698 plus.n68 gnd 0.022489f
C699 plus.n69 gnd 0.022489f
C700 plus.n70 gnd 0.029288f
C701 plus.n71 gnd 0.009314f
C702 plus.t12 gnd 0.408961f
C703 plus.n72 gnd 0.17763f
C704 plus.n73 gnd 0.691723f
C705 plus.n74 gnd 1.04434f
C706 plus.t4 gnd 0.038822f
C707 plus.t1 gnd 0.006933f
C708 plus.t2 gnd 0.006933f
C709 plus.n75 gnd 0.022483f
C710 plus.n76 gnd 0.174542f
C711 plus.t0 gnd 0.006933f
C712 plus.t3 gnd 0.006933f
C713 plus.n77 gnd 0.022483f
C714 plus.n78 gnd 0.131015f
C715 plus.n79 gnd 2.30863f
C716 commonsourceibias.n0 gnd 0.010301f
C717 commonsourceibias.t71 gnd 0.155981f
C718 commonsourceibias.t81 gnd 0.144227f
C719 commonsourceibias.n1 gnd 0.057546f
C720 commonsourceibias.n2 gnd 0.00772f
C721 commonsourceibias.t55 gnd 0.144227f
C722 commonsourceibias.n3 gnd 0.006245f
C723 commonsourceibias.n4 gnd 0.00772f
C724 commonsourceibias.t53 gnd 0.144227f
C725 commonsourceibias.n5 gnd 0.007453f
C726 commonsourceibias.n6 gnd 0.00772f
C727 commonsourceibias.t76 gnd 0.144227f
C728 commonsourceibias.n7 gnd 0.057546f
C729 commonsourceibias.t86 gnd 0.144227f
C730 commonsourceibias.n8 gnd 0.006235f
C731 commonsourceibias.n9 gnd 0.010301f
C732 commonsourceibias.t32 gnd 0.155981f
C733 commonsourceibias.t14 gnd 0.144227f
C734 commonsourceibias.n10 gnd 0.057546f
C735 commonsourceibias.n11 gnd 0.00772f
C736 commonsourceibias.t24 gnd 0.144227f
C737 commonsourceibias.n12 gnd 0.006245f
C738 commonsourceibias.n13 gnd 0.00772f
C739 commonsourceibias.t30 gnd 0.144227f
C740 commonsourceibias.n14 gnd 0.007453f
C741 commonsourceibias.n15 gnd 0.00772f
C742 commonsourceibias.t20 gnd 0.144227f
C743 commonsourceibias.n16 gnd 0.057546f
C744 commonsourceibias.t36 gnd 0.144227f
C745 commonsourceibias.n17 gnd 0.006235f
C746 commonsourceibias.n18 gnd 0.00772f
C747 commonsourceibias.t44 gnd 0.144227f
C748 commonsourceibias.t26 gnd 0.144227f
C749 commonsourceibias.n19 gnd 0.057546f
C750 commonsourceibias.n20 gnd 0.00772f
C751 commonsourceibias.t34 gnd 0.144227f
C752 commonsourceibias.n21 gnd 0.057546f
C753 commonsourceibias.n22 gnd 0.00772f
C754 commonsourceibias.t10 gnd 0.144227f
C755 commonsourceibias.n23 gnd 0.057546f
C756 commonsourceibias.n24 gnd 0.038863f
C757 commonsourceibias.t40 gnd 0.144227f
C758 commonsourceibias.t46 gnd 0.162743f
C759 commonsourceibias.n25 gnd 0.066782f
C760 commonsourceibias.n26 gnd 0.069137f
C761 commonsourceibias.n27 gnd 0.009515f
C762 commonsourceibias.n28 gnd 0.010526f
C763 commonsourceibias.n29 gnd 0.00772f
C764 commonsourceibias.n30 gnd 0.00772f
C765 commonsourceibias.n31 gnd 0.010457f
C766 commonsourceibias.n32 gnd 0.006245f
C767 commonsourceibias.n33 gnd 0.010587f
C768 commonsourceibias.n34 gnd 0.00772f
C769 commonsourceibias.n35 gnd 0.00772f
C770 commonsourceibias.n36 gnd 0.010651f
C771 commonsourceibias.n37 gnd 0.009185f
C772 commonsourceibias.n38 gnd 0.007453f
C773 commonsourceibias.n39 gnd 0.00772f
C774 commonsourceibias.n40 gnd 0.00772f
C775 commonsourceibias.n41 gnd 0.009442f
C776 commonsourceibias.n42 gnd 0.010598f
C777 commonsourceibias.n43 gnd 0.057546f
C778 commonsourceibias.n44 gnd 0.010527f
C779 commonsourceibias.n45 gnd 0.00772f
C780 commonsourceibias.n46 gnd 0.00772f
C781 commonsourceibias.n47 gnd 0.00772f
C782 commonsourceibias.n48 gnd 0.010527f
C783 commonsourceibias.n49 gnd 0.057546f
C784 commonsourceibias.n50 gnd 0.010598f
C785 commonsourceibias.n51 gnd 0.009442f
C786 commonsourceibias.n52 gnd 0.00772f
C787 commonsourceibias.n53 gnd 0.00772f
C788 commonsourceibias.n54 gnd 0.00772f
C789 commonsourceibias.n55 gnd 0.009185f
C790 commonsourceibias.n56 gnd 0.010651f
C791 commonsourceibias.n57 gnd 0.057546f
C792 commonsourceibias.n58 gnd 0.010587f
C793 commonsourceibias.n59 gnd 0.00772f
C794 commonsourceibias.n60 gnd 0.00772f
C795 commonsourceibias.n61 gnd 0.00772f
C796 commonsourceibias.n62 gnd 0.010457f
C797 commonsourceibias.n63 gnd 0.057546f
C798 commonsourceibias.n64 gnd 0.010526f
C799 commonsourceibias.n65 gnd 0.009515f
C800 commonsourceibias.n66 gnd 0.00772f
C801 commonsourceibias.n67 gnd 0.00772f
C802 commonsourceibias.n68 gnd 0.007831f
C803 commonsourceibias.n69 gnd 0.008096f
C804 commonsourceibias.n70 gnd 0.068855f
C805 commonsourceibias.n71 gnd 0.076384f
C806 commonsourceibias.t33 gnd 0.016658f
C807 commonsourceibias.t15 gnd 0.016658f
C808 commonsourceibias.n72 gnd 0.147197f
C809 commonsourceibias.n73 gnd 0.12719f
C810 commonsourceibias.t25 gnd 0.016658f
C811 commonsourceibias.t31 gnd 0.016658f
C812 commonsourceibias.n74 gnd 0.147197f
C813 commonsourceibias.n75 gnd 0.067614f
C814 commonsourceibias.t21 gnd 0.016658f
C815 commonsourceibias.t37 gnd 0.016658f
C816 commonsourceibias.n76 gnd 0.147197f
C817 commonsourceibias.n77 gnd 0.056488f
C818 commonsourceibias.t41 gnd 0.016658f
C819 commonsourceibias.t47 gnd 0.016658f
C820 commonsourceibias.n78 gnd 0.14769f
C821 commonsourceibias.t35 gnd 0.016658f
C822 commonsourceibias.t11 gnd 0.016658f
C823 commonsourceibias.n79 gnd 0.147197f
C824 commonsourceibias.n80 gnd 0.13716f
C825 commonsourceibias.t45 gnd 0.016658f
C826 commonsourceibias.t27 gnd 0.016658f
C827 commonsourceibias.n81 gnd 0.147197f
C828 commonsourceibias.n82 gnd 0.056488f
C829 commonsourceibias.n83 gnd 0.068401f
C830 commonsourceibias.n84 gnd 0.00772f
C831 commonsourceibias.t50 gnd 0.144227f
C832 commonsourceibias.t69 gnd 0.144227f
C833 commonsourceibias.n85 gnd 0.057546f
C834 commonsourceibias.n86 gnd 0.00772f
C835 commonsourceibias.t67 gnd 0.144227f
C836 commonsourceibias.n87 gnd 0.057546f
C837 commonsourceibias.n88 gnd 0.00772f
C838 commonsourceibias.t78 gnd 0.144227f
C839 commonsourceibias.n89 gnd 0.057546f
C840 commonsourceibias.n90 gnd 0.038863f
C841 commonsourceibias.t64 gnd 0.144227f
C842 commonsourceibias.t62 gnd 0.162743f
C843 commonsourceibias.n91 gnd 0.066782f
C844 commonsourceibias.n92 gnd 0.069137f
C845 commonsourceibias.n93 gnd 0.009515f
C846 commonsourceibias.n94 gnd 0.010526f
C847 commonsourceibias.n95 gnd 0.00772f
C848 commonsourceibias.n96 gnd 0.00772f
C849 commonsourceibias.n97 gnd 0.010457f
C850 commonsourceibias.n98 gnd 0.006245f
C851 commonsourceibias.n99 gnd 0.010587f
C852 commonsourceibias.n100 gnd 0.00772f
C853 commonsourceibias.n101 gnd 0.00772f
C854 commonsourceibias.n102 gnd 0.010651f
C855 commonsourceibias.n103 gnd 0.009185f
C856 commonsourceibias.n104 gnd 0.007453f
C857 commonsourceibias.n105 gnd 0.00772f
C858 commonsourceibias.n106 gnd 0.00772f
C859 commonsourceibias.n107 gnd 0.009442f
C860 commonsourceibias.n108 gnd 0.010598f
C861 commonsourceibias.n109 gnd 0.057546f
C862 commonsourceibias.n110 gnd 0.010527f
C863 commonsourceibias.n111 gnd 0.007683f
C864 commonsourceibias.n112 gnd 0.055804f
C865 commonsourceibias.n113 gnd 0.007683f
C866 commonsourceibias.n114 gnd 0.010527f
C867 commonsourceibias.n115 gnd 0.057546f
C868 commonsourceibias.n116 gnd 0.010598f
C869 commonsourceibias.n117 gnd 0.009442f
C870 commonsourceibias.n118 gnd 0.00772f
C871 commonsourceibias.n119 gnd 0.00772f
C872 commonsourceibias.n120 gnd 0.00772f
C873 commonsourceibias.n121 gnd 0.009185f
C874 commonsourceibias.n122 gnd 0.010651f
C875 commonsourceibias.n123 gnd 0.057546f
C876 commonsourceibias.n124 gnd 0.010587f
C877 commonsourceibias.n125 gnd 0.00772f
C878 commonsourceibias.n126 gnd 0.00772f
C879 commonsourceibias.n127 gnd 0.00772f
C880 commonsourceibias.n128 gnd 0.010457f
C881 commonsourceibias.n129 gnd 0.057546f
C882 commonsourceibias.n130 gnd 0.010526f
C883 commonsourceibias.n131 gnd 0.009515f
C884 commonsourceibias.n132 gnd 0.00772f
C885 commonsourceibias.n133 gnd 0.00772f
C886 commonsourceibias.n134 gnd 0.007831f
C887 commonsourceibias.n135 gnd 0.008096f
C888 commonsourceibias.n136 gnd 0.068855f
C889 commonsourceibias.n137 gnd 0.04456f
C890 commonsourceibias.n138 gnd 0.010301f
C891 commonsourceibias.t72 gnd 0.144227f
C892 commonsourceibias.n139 gnd 0.057546f
C893 commonsourceibias.n140 gnd 0.00772f
C894 commonsourceibias.t49 gnd 0.144227f
C895 commonsourceibias.n141 gnd 0.006245f
C896 commonsourceibias.n142 gnd 0.00772f
C897 commonsourceibias.t95 gnd 0.144227f
C898 commonsourceibias.n143 gnd 0.007453f
C899 commonsourceibias.n144 gnd 0.00772f
C900 commonsourceibias.t66 gnd 0.144227f
C901 commonsourceibias.n145 gnd 0.057546f
C902 commonsourceibias.t77 gnd 0.144227f
C903 commonsourceibias.n146 gnd 0.006235f
C904 commonsourceibias.n147 gnd 0.00772f
C905 commonsourceibias.t91 gnd 0.144227f
C906 commonsourceibias.t60 gnd 0.144227f
C907 commonsourceibias.n148 gnd 0.057546f
C908 commonsourceibias.n149 gnd 0.00772f
C909 commonsourceibias.t58 gnd 0.144227f
C910 commonsourceibias.n150 gnd 0.057546f
C911 commonsourceibias.n151 gnd 0.00772f
C912 commonsourceibias.t68 gnd 0.144227f
C913 commonsourceibias.n152 gnd 0.057546f
C914 commonsourceibias.n153 gnd 0.038863f
C915 commonsourceibias.t57 gnd 0.144227f
C916 commonsourceibias.t54 gnd 0.162743f
C917 commonsourceibias.n154 gnd 0.066782f
C918 commonsourceibias.n155 gnd 0.069137f
C919 commonsourceibias.n156 gnd 0.009515f
C920 commonsourceibias.n157 gnd 0.010526f
C921 commonsourceibias.n158 gnd 0.00772f
C922 commonsourceibias.n159 gnd 0.00772f
C923 commonsourceibias.n160 gnd 0.010457f
C924 commonsourceibias.n161 gnd 0.006245f
C925 commonsourceibias.n162 gnd 0.010587f
C926 commonsourceibias.n163 gnd 0.00772f
C927 commonsourceibias.n164 gnd 0.00772f
C928 commonsourceibias.n165 gnd 0.010651f
C929 commonsourceibias.n166 gnd 0.009185f
C930 commonsourceibias.n167 gnd 0.007453f
C931 commonsourceibias.n168 gnd 0.00772f
C932 commonsourceibias.n169 gnd 0.00772f
C933 commonsourceibias.n170 gnd 0.009442f
C934 commonsourceibias.n171 gnd 0.010598f
C935 commonsourceibias.n172 gnd 0.057546f
C936 commonsourceibias.n173 gnd 0.010527f
C937 commonsourceibias.n174 gnd 0.00772f
C938 commonsourceibias.n175 gnd 0.00772f
C939 commonsourceibias.n176 gnd 0.00772f
C940 commonsourceibias.n177 gnd 0.010527f
C941 commonsourceibias.n178 gnd 0.057546f
C942 commonsourceibias.n179 gnd 0.010598f
C943 commonsourceibias.n180 gnd 0.009442f
C944 commonsourceibias.n181 gnd 0.00772f
C945 commonsourceibias.n182 gnd 0.00772f
C946 commonsourceibias.n183 gnd 0.00772f
C947 commonsourceibias.n184 gnd 0.009185f
C948 commonsourceibias.n185 gnd 0.010651f
C949 commonsourceibias.n186 gnd 0.057546f
C950 commonsourceibias.n187 gnd 0.010587f
C951 commonsourceibias.n188 gnd 0.00772f
C952 commonsourceibias.n189 gnd 0.00772f
C953 commonsourceibias.n190 gnd 0.00772f
C954 commonsourceibias.n191 gnd 0.010457f
C955 commonsourceibias.n192 gnd 0.057546f
C956 commonsourceibias.n193 gnd 0.010526f
C957 commonsourceibias.n194 gnd 0.009515f
C958 commonsourceibias.n195 gnd 0.00772f
C959 commonsourceibias.n196 gnd 0.00772f
C960 commonsourceibias.n197 gnd 0.007831f
C961 commonsourceibias.n198 gnd 0.008096f
C962 commonsourceibias.t61 gnd 0.155981f
C963 commonsourceibias.n199 gnd 0.068855f
C964 commonsourceibias.n200 gnd 0.023432f
C965 commonsourceibias.n201 gnd 0.388694f
C966 commonsourceibias.n202 gnd 0.010301f
C967 commonsourceibias.t84 gnd 0.155981f
C968 commonsourceibias.t92 gnd 0.144227f
C969 commonsourceibias.n203 gnd 0.057546f
C970 commonsourceibias.n204 gnd 0.00772f
C971 commonsourceibias.t51 gnd 0.144227f
C972 commonsourceibias.n205 gnd 0.006245f
C973 commonsourceibias.n206 gnd 0.00772f
C974 commonsourceibias.t63 gnd 0.144227f
C975 commonsourceibias.n207 gnd 0.007453f
C976 commonsourceibias.n208 gnd 0.00772f
C977 commonsourceibias.t48 gnd 0.144227f
C978 commonsourceibias.n209 gnd 0.006235f
C979 commonsourceibias.n210 gnd 0.00772f
C980 commonsourceibias.t94 gnd 0.144227f
C981 commonsourceibias.t83 gnd 0.144227f
C982 commonsourceibias.n211 gnd 0.057546f
C983 commonsourceibias.n212 gnd 0.00772f
C984 commonsourceibias.t80 gnd 0.144227f
C985 commonsourceibias.n213 gnd 0.057546f
C986 commonsourceibias.n214 gnd 0.00772f
C987 commonsourceibias.t90 gnd 0.144227f
C988 commonsourceibias.n215 gnd 0.057546f
C989 commonsourceibias.n216 gnd 0.038863f
C990 commonsourceibias.t59 gnd 0.144227f
C991 commonsourceibias.t75 gnd 0.162743f
C992 commonsourceibias.n217 gnd 0.066782f
C993 commonsourceibias.n218 gnd 0.069137f
C994 commonsourceibias.n219 gnd 0.009515f
C995 commonsourceibias.n220 gnd 0.010526f
C996 commonsourceibias.n221 gnd 0.00772f
C997 commonsourceibias.n222 gnd 0.00772f
C998 commonsourceibias.n223 gnd 0.010457f
C999 commonsourceibias.n224 gnd 0.006245f
C1000 commonsourceibias.n225 gnd 0.010587f
C1001 commonsourceibias.n226 gnd 0.00772f
C1002 commonsourceibias.n227 gnd 0.00772f
C1003 commonsourceibias.n228 gnd 0.010651f
C1004 commonsourceibias.n229 gnd 0.009185f
C1005 commonsourceibias.n230 gnd 0.007453f
C1006 commonsourceibias.n231 gnd 0.00772f
C1007 commonsourceibias.n232 gnd 0.00772f
C1008 commonsourceibias.n233 gnd 0.009442f
C1009 commonsourceibias.n234 gnd 0.010598f
C1010 commonsourceibias.n235 gnd 0.057546f
C1011 commonsourceibias.n236 gnd 0.010527f
C1012 commonsourceibias.n237 gnd 0.007683f
C1013 commonsourceibias.t17 gnd 0.016658f
C1014 commonsourceibias.t9 gnd 0.016658f
C1015 commonsourceibias.n238 gnd 0.14769f
C1016 commonsourceibias.t19 gnd 0.016658f
C1017 commonsourceibias.t5 gnd 0.016658f
C1018 commonsourceibias.n239 gnd 0.147197f
C1019 commonsourceibias.n240 gnd 0.13716f
C1020 commonsourceibias.t43 gnd 0.016658f
C1021 commonsourceibias.t13 gnd 0.016658f
C1022 commonsourceibias.n241 gnd 0.147197f
C1023 commonsourceibias.n242 gnd 0.056488f
C1024 commonsourceibias.n243 gnd 0.010301f
C1025 commonsourceibias.t22 gnd 0.144227f
C1026 commonsourceibias.n244 gnd 0.057546f
C1027 commonsourceibias.n245 gnd 0.00772f
C1028 commonsourceibias.t38 gnd 0.144227f
C1029 commonsourceibias.n246 gnd 0.006245f
C1030 commonsourceibias.n247 gnd 0.00772f
C1031 commonsourceibias.t0 gnd 0.144227f
C1032 commonsourceibias.n248 gnd 0.007453f
C1033 commonsourceibias.n249 gnd 0.00772f
C1034 commonsourceibias.t6 gnd 0.144227f
C1035 commonsourceibias.n250 gnd 0.006235f
C1036 commonsourceibias.n251 gnd 0.00772f
C1037 commonsourceibias.t12 gnd 0.144227f
C1038 commonsourceibias.t42 gnd 0.144227f
C1039 commonsourceibias.n252 gnd 0.057546f
C1040 commonsourceibias.n253 gnd 0.00772f
C1041 commonsourceibias.t4 gnd 0.144227f
C1042 commonsourceibias.n254 gnd 0.057546f
C1043 commonsourceibias.n255 gnd 0.00772f
C1044 commonsourceibias.t18 gnd 0.144227f
C1045 commonsourceibias.n256 gnd 0.057546f
C1046 commonsourceibias.n257 gnd 0.038863f
C1047 commonsourceibias.t8 gnd 0.144227f
C1048 commonsourceibias.t16 gnd 0.162743f
C1049 commonsourceibias.n258 gnd 0.066782f
C1050 commonsourceibias.n259 gnd 0.069137f
C1051 commonsourceibias.n260 gnd 0.009515f
C1052 commonsourceibias.n261 gnd 0.010526f
C1053 commonsourceibias.n262 gnd 0.00772f
C1054 commonsourceibias.n263 gnd 0.00772f
C1055 commonsourceibias.n264 gnd 0.010457f
C1056 commonsourceibias.n265 gnd 0.006245f
C1057 commonsourceibias.n266 gnd 0.010587f
C1058 commonsourceibias.n267 gnd 0.00772f
C1059 commonsourceibias.n268 gnd 0.00772f
C1060 commonsourceibias.n269 gnd 0.010651f
C1061 commonsourceibias.n270 gnd 0.009185f
C1062 commonsourceibias.n271 gnd 0.007453f
C1063 commonsourceibias.n272 gnd 0.00772f
C1064 commonsourceibias.n273 gnd 0.00772f
C1065 commonsourceibias.n274 gnd 0.009442f
C1066 commonsourceibias.n275 gnd 0.010598f
C1067 commonsourceibias.n276 gnd 0.057546f
C1068 commonsourceibias.n277 gnd 0.010527f
C1069 commonsourceibias.n278 gnd 0.00772f
C1070 commonsourceibias.n279 gnd 0.00772f
C1071 commonsourceibias.n280 gnd 0.00772f
C1072 commonsourceibias.n281 gnd 0.010527f
C1073 commonsourceibias.n282 gnd 0.057546f
C1074 commonsourceibias.n283 gnd 0.010598f
C1075 commonsourceibias.t28 gnd 0.144227f
C1076 commonsourceibias.n284 gnd 0.057546f
C1077 commonsourceibias.n285 gnd 0.009442f
C1078 commonsourceibias.n286 gnd 0.00772f
C1079 commonsourceibias.n287 gnd 0.00772f
C1080 commonsourceibias.n288 gnd 0.00772f
C1081 commonsourceibias.n289 gnd 0.009185f
C1082 commonsourceibias.n290 gnd 0.010651f
C1083 commonsourceibias.n291 gnd 0.057546f
C1084 commonsourceibias.n292 gnd 0.010587f
C1085 commonsourceibias.n293 gnd 0.00772f
C1086 commonsourceibias.n294 gnd 0.00772f
C1087 commonsourceibias.n295 gnd 0.00772f
C1088 commonsourceibias.n296 gnd 0.010457f
C1089 commonsourceibias.n297 gnd 0.057546f
C1090 commonsourceibias.n298 gnd 0.010526f
C1091 commonsourceibias.n299 gnd 0.009515f
C1092 commonsourceibias.n300 gnd 0.00772f
C1093 commonsourceibias.n301 gnd 0.00772f
C1094 commonsourceibias.n302 gnd 0.007831f
C1095 commonsourceibias.n303 gnd 0.008096f
C1096 commonsourceibias.t2 gnd 0.155981f
C1097 commonsourceibias.n304 gnd 0.068855f
C1098 commonsourceibias.n305 gnd 0.076384f
C1099 commonsourceibias.t23 gnd 0.016658f
C1100 commonsourceibias.t3 gnd 0.016658f
C1101 commonsourceibias.n306 gnd 0.147197f
C1102 commonsourceibias.n307 gnd 0.12719f
C1103 commonsourceibias.t1 gnd 0.016658f
C1104 commonsourceibias.t39 gnd 0.016658f
C1105 commonsourceibias.n308 gnd 0.147197f
C1106 commonsourceibias.n309 gnd 0.067614f
C1107 commonsourceibias.t7 gnd 0.016658f
C1108 commonsourceibias.t29 gnd 0.016658f
C1109 commonsourceibias.n310 gnd 0.147197f
C1110 commonsourceibias.n311 gnd 0.056488f
C1111 commonsourceibias.n312 gnd 0.068401f
C1112 commonsourceibias.n313 gnd 0.055804f
C1113 commonsourceibias.n314 gnd 0.007683f
C1114 commonsourceibias.n315 gnd 0.010527f
C1115 commonsourceibias.n316 gnd 0.057546f
C1116 commonsourceibias.n317 gnd 0.010598f
C1117 commonsourceibias.t88 gnd 0.144227f
C1118 commonsourceibias.n318 gnd 0.057546f
C1119 commonsourceibias.n319 gnd 0.009442f
C1120 commonsourceibias.n320 gnd 0.00772f
C1121 commonsourceibias.n321 gnd 0.00772f
C1122 commonsourceibias.n322 gnd 0.00772f
C1123 commonsourceibias.n323 gnd 0.009185f
C1124 commonsourceibias.n324 gnd 0.010651f
C1125 commonsourceibias.n325 gnd 0.057546f
C1126 commonsourceibias.n326 gnd 0.010587f
C1127 commonsourceibias.n327 gnd 0.00772f
C1128 commonsourceibias.n328 gnd 0.00772f
C1129 commonsourceibias.n329 gnd 0.00772f
C1130 commonsourceibias.n330 gnd 0.010457f
C1131 commonsourceibias.n331 gnd 0.057546f
C1132 commonsourceibias.n332 gnd 0.010526f
C1133 commonsourceibias.n333 gnd 0.009515f
C1134 commonsourceibias.n334 gnd 0.00772f
C1135 commonsourceibias.n335 gnd 0.00772f
C1136 commonsourceibias.n336 gnd 0.007831f
C1137 commonsourceibias.n337 gnd 0.008096f
C1138 commonsourceibias.n338 gnd 0.068855f
C1139 commonsourceibias.n339 gnd 0.04456f
C1140 commonsourceibias.n340 gnd 0.010301f
C1141 commonsourceibias.t85 gnd 0.144227f
C1142 commonsourceibias.n341 gnd 0.057546f
C1143 commonsourceibias.n342 gnd 0.00772f
C1144 commonsourceibias.t93 gnd 0.144227f
C1145 commonsourceibias.n343 gnd 0.006245f
C1146 commonsourceibias.n344 gnd 0.00772f
C1147 commonsourceibias.t56 gnd 0.144227f
C1148 commonsourceibias.n345 gnd 0.007453f
C1149 commonsourceibias.n346 gnd 0.00772f
C1150 commonsourceibias.t89 gnd 0.144227f
C1151 commonsourceibias.n347 gnd 0.006235f
C1152 commonsourceibias.n348 gnd 0.00772f
C1153 commonsourceibias.t87 gnd 0.144227f
C1154 commonsourceibias.t74 gnd 0.144227f
C1155 commonsourceibias.n349 gnd 0.057546f
C1156 commonsourceibias.n350 gnd 0.00772f
C1157 commonsourceibias.t70 gnd 0.144227f
C1158 commonsourceibias.n351 gnd 0.057546f
C1159 commonsourceibias.n352 gnd 0.00772f
C1160 commonsourceibias.t82 gnd 0.144227f
C1161 commonsourceibias.n353 gnd 0.057546f
C1162 commonsourceibias.n354 gnd 0.038863f
C1163 commonsourceibias.t52 gnd 0.144227f
C1164 commonsourceibias.t65 gnd 0.162743f
C1165 commonsourceibias.n355 gnd 0.066782f
C1166 commonsourceibias.n356 gnd 0.069137f
C1167 commonsourceibias.n357 gnd 0.009515f
C1168 commonsourceibias.n358 gnd 0.010526f
C1169 commonsourceibias.n359 gnd 0.00772f
C1170 commonsourceibias.n360 gnd 0.00772f
C1171 commonsourceibias.n361 gnd 0.010457f
C1172 commonsourceibias.n362 gnd 0.006245f
C1173 commonsourceibias.n363 gnd 0.010587f
C1174 commonsourceibias.n364 gnd 0.00772f
C1175 commonsourceibias.n365 gnd 0.00772f
C1176 commonsourceibias.n366 gnd 0.010651f
C1177 commonsourceibias.n367 gnd 0.009185f
C1178 commonsourceibias.n368 gnd 0.007453f
C1179 commonsourceibias.n369 gnd 0.00772f
C1180 commonsourceibias.n370 gnd 0.00772f
C1181 commonsourceibias.n371 gnd 0.009442f
C1182 commonsourceibias.n372 gnd 0.010598f
C1183 commonsourceibias.n373 gnd 0.057546f
C1184 commonsourceibias.n374 gnd 0.010527f
C1185 commonsourceibias.n375 gnd 0.00772f
C1186 commonsourceibias.n376 gnd 0.00772f
C1187 commonsourceibias.n377 gnd 0.00772f
C1188 commonsourceibias.n378 gnd 0.010527f
C1189 commonsourceibias.n379 gnd 0.057546f
C1190 commonsourceibias.n380 gnd 0.010598f
C1191 commonsourceibias.t79 gnd 0.144227f
C1192 commonsourceibias.n381 gnd 0.057546f
C1193 commonsourceibias.n382 gnd 0.009442f
C1194 commonsourceibias.n383 gnd 0.00772f
C1195 commonsourceibias.n384 gnd 0.00772f
C1196 commonsourceibias.n385 gnd 0.00772f
C1197 commonsourceibias.n386 gnd 0.009185f
C1198 commonsourceibias.n387 gnd 0.010651f
C1199 commonsourceibias.n388 gnd 0.057546f
C1200 commonsourceibias.n389 gnd 0.010587f
C1201 commonsourceibias.n390 gnd 0.00772f
C1202 commonsourceibias.n391 gnd 0.00772f
C1203 commonsourceibias.n392 gnd 0.00772f
C1204 commonsourceibias.n393 gnd 0.010457f
C1205 commonsourceibias.n394 gnd 0.057546f
C1206 commonsourceibias.n395 gnd 0.010526f
C1207 commonsourceibias.n396 gnd 0.009515f
C1208 commonsourceibias.n397 gnd 0.00772f
C1209 commonsourceibias.n398 gnd 0.00772f
C1210 commonsourceibias.n399 gnd 0.007831f
C1211 commonsourceibias.n400 gnd 0.008096f
C1212 commonsourceibias.t73 gnd 0.155981f
C1213 commonsourceibias.n401 gnd 0.068855f
C1214 commonsourceibias.n402 gnd 0.023432f
C1215 commonsourceibias.n403 gnd 0.212991f
C1216 commonsourceibias.n404 gnd 4.01312f
C1217 CSoutput.n0 gnd 0.044771f
C1218 CSoutput.t156 gnd 0.29615f
C1219 CSoutput.n1 gnd 0.133727f
C1220 CSoutput.n2 gnd 0.044771f
C1221 CSoutput.t161 gnd 0.29615f
C1222 CSoutput.n3 gnd 0.035485f
C1223 CSoutput.n4 gnd 0.044771f
C1224 CSoutput.t150 gnd 0.29615f
C1225 CSoutput.n5 gnd 0.030599f
C1226 CSoutput.n6 gnd 0.044771f
C1227 CSoutput.t159 gnd 0.29615f
C1228 CSoutput.t165 gnd 0.29615f
C1229 CSoutput.n7 gnd 0.132269f
C1230 CSoutput.n8 gnd 0.044771f
C1231 CSoutput.t163 gnd 0.29615f
C1232 CSoutput.n9 gnd 0.029174f
C1233 CSoutput.n10 gnd 0.044771f
C1234 CSoutput.t151 gnd 0.29615f
C1235 CSoutput.t162 gnd 0.29615f
C1236 CSoutput.n11 gnd 0.132269f
C1237 CSoutput.n12 gnd 0.044771f
C1238 CSoutput.t160 gnd 0.29615f
C1239 CSoutput.n13 gnd 0.030599f
C1240 CSoutput.n14 gnd 0.044771f
C1241 CSoutput.t149 gnd 0.29615f
C1242 CSoutput.t155 gnd 0.29615f
C1243 CSoutput.n15 gnd 0.132269f
C1244 CSoutput.n16 gnd 0.044771f
C1245 CSoutput.t158 gnd 0.29615f
C1246 CSoutput.n17 gnd 0.032681f
C1247 CSoutput.t145 gnd 0.353907f
C1248 CSoutput.t147 gnd 0.29615f
C1249 CSoutput.n18 gnd 0.168856f
C1250 CSoutput.n19 gnd 0.163849f
C1251 CSoutput.n20 gnd 0.190084f
C1252 CSoutput.n21 gnd 0.044771f
C1253 CSoutput.n22 gnd 0.037366f
C1254 CSoutput.n23 gnd 0.132269f
C1255 CSoutput.n24 gnd 0.03602f
C1256 CSoutput.n25 gnd 0.035485f
C1257 CSoutput.n26 gnd 0.044771f
C1258 CSoutput.n27 gnd 0.044771f
C1259 CSoutput.n28 gnd 0.037079f
C1260 CSoutput.n29 gnd 0.031481f
C1261 CSoutput.n30 gnd 0.135214f
C1262 CSoutput.n31 gnd 0.031915f
C1263 CSoutput.n32 gnd 0.044771f
C1264 CSoutput.n33 gnd 0.044771f
C1265 CSoutput.n34 gnd 0.044771f
C1266 CSoutput.n35 gnd 0.036684f
C1267 CSoutput.n36 gnd 0.132269f
C1268 CSoutput.n37 gnd 0.035083f
C1269 CSoutput.n38 gnd 0.036422f
C1270 CSoutput.n39 gnd 0.044771f
C1271 CSoutput.n40 gnd 0.044771f
C1272 CSoutput.n41 gnd 0.037359f
C1273 CSoutput.n42 gnd 0.034146f
C1274 CSoutput.n43 gnd 0.132269f
C1275 CSoutput.n44 gnd 0.035012f
C1276 CSoutput.n45 gnd 0.044771f
C1277 CSoutput.n46 gnd 0.044771f
C1278 CSoutput.n47 gnd 0.044771f
C1279 CSoutput.n48 gnd 0.035012f
C1280 CSoutput.n49 gnd 0.132269f
C1281 CSoutput.n50 gnd 0.034146f
C1282 CSoutput.n51 gnd 0.037359f
C1283 CSoutput.n52 gnd 0.044771f
C1284 CSoutput.n53 gnd 0.044771f
C1285 CSoutput.n54 gnd 0.036422f
C1286 CSoutput.n55 gnd 0.035083f
C1287 CSoutput.n56 gnd 0.132269f
C1288 CSoutput.n57 gnd 0.036684f
C1289 CSoutput.n58 gnd 0.044771f
C1290 CSoutput.n59 gnd 0.044771f
C1291 CSoutput.n60 gnd 0.044771f
C1292 CSoutput.n61 gnd 0.031915f
C1293 CSoutput.n62 gnd 0.135214f
C1294 CSoutput.n63 gnd 0.031481f
C1295 CSoutput.t144 gnd 0.29615f
C1296 CSoutput.n64 gnd 0.132269f
C1297 CSoutput.n65 gnd 0.037079f
C1298 CSoutput.n66 gnd 0.044771f
C1299 CSoutput.n67 gnd 0.044771f
C1300 CSoutput.n68 gnd 0.044771f
C1301 CSoutput.n69 gnd 0.03602f
C1302 CSoutput.n70 gnd 0.132269f
C1303 CSoutput.n71 gnd 0.037366f
C1304 CSoutput.n72 gnd 0.032681f
C1305 CSoutput.n73 gnd 0.044771f
C1306 CSoutput.n74 gnd 0.044771f
C1307 CSoutput.n75 gnd 0.033892f
C1308 CSoutput.n76 gnd 0.020129f
C1309 CSoutput.t148 gnd 0.332746f
C1310 CSoutput.n77 gnd 0.165295f
C1311 CSoutput.n78 gnd 0.707281f
C1312 CSoutput.t93 gnd 0.055846f
C1313 CSoutput.t41 gnd 0.055846f
C1314 CSoutput.n79 gnd 0.432374f
C1315 CSoutput.t105 gnd 0.055846f
C1316 CSoutput.t58 gnd 0.055846f
C1317 CSoutput.n80 gnd 0.431603f
C1318 CSoutput.n81 gnd 0.438077f
C1319 CSoutput.t22 gnd 0.055846f
C1320 CSoutput.t69 gnd 0.055846f
C1321 CSoutput.n82 gnd 0.431603f
C1322 CSoutput.n83 gnd 0.215866f
C1323 CSoutput.t25 gnd 0.055846f
C1324 CSoutput.t50 gnd 0.055846f
C1325 CSoutput.n84 gnd 0.431603f
C1326 CSoutput.n85 gnd 0.215866f
C1327 CSoutput.t110 gnd 0.055846f
C1328 CSoutput.t64 gnd 0.055846f
C1329 CSoutput.n86 gnd 0.431603f
C1330 CSoutput.n87 gnd 0.215866f
C1331 CSoutput.t28 gnd 0.055846f
C1332 CSoutput.t96 gnd 0.055846f
C1333 CSoutput.n88 gnd 0.431603f
C1334 CSoutput.n89 gnd 0.215866f
C1335 CSoutput.t36 gnd 0.055846f
C1336 CSoutput.t78 gnd 0.055846f
C1337 CSoutput.n90 gnd 0.431603f
C1338 CSoutput.n91 gnd 0.215866f
C1339 CSoutput.t53 gnd 0.055846f
C1340 CSoutput.t71 gnd 0.055846f
C1341 CSoutput.n92 gnd 0.431603f
C1342 CSoutput.n93 gnd 0.395848f
C1343 CSoutput.t19 gnd 0.055846f
C1344 CSoutput.t90 gnd 0.055846f
C1345 CSoutput.n94 gnd 0.432374f
C1346 CSoutput.t81 gnd 0.055846f
C1347 CSoutput.t59 gnd 0.055846f
C1348 CSoutput.n95 gnd 0.431603f
C1349 CSoutput.n96 gnd 0.438077f
C1350 CSoutput.t42 gnd 0.055846f
C1351 CSoutput.t103 gnd 0.055846f
C1352 CSoutput.n97 gnd 0.431603f
C1353 CSoutput.n98 gnd 0.215866f
C1354 CSoutput.t80 gnd 0.055846f
C1355 CSoutput.t77 gnd 0.055846f
C1356 CSoutput.n99 gnd 0.431603f
C1357 CSoutput.n100 gnd 0.215866f
C1358 CSoutput.t68 gnd 0.055846f
C1359 CSoutput.t38 gnd 0.055846f
C1360 CSoutput.n101 gnd 0.431603f
C1361 CSoutput.n102 gnd 0.215866f
C1362 CSoutput.t21 gnd 0.055846f
C1363 CSoutput.t67 gnd 0.055846f
C1364 CSoutput.n103 gnd 0.431603f
C1365 CSoutput.n104 gnd 0.215866f
C1366 CSoutput.t66 gnd 0.055846f
C1367 CSoutput.t37 gnd 0.055846f
C1368 CSoutput.n105 gnd 0.431603f
C1369 CSoutput.n106 gnd 0.215866f
C1370 CSoutput.t17 gnd 0.055846f
C1371 CSoutput.t18 gnd 0.055846f
C1372 CSoutput.n107 gnd 0.431603f
C1373 CSoutput.n108 gnd 0.32191f
C1374 CSoutput.n109 gnd 0.405927f
C1375 CSoutput.t32 gnd 0.055846f
C1376 CSoutput.t102 gnd 0.055846f
C1377 CSoutput.n110 gnd 0.432374f
C1378 CSoutput.t88 gnd 0.055846f
C1379 CSoutput.t70 gnd 0.055846f
C1380 CSoutput.n111 gnd 0.431603f
C1381 CSoutput.n112 gnd 0.438077f
C1382 CSoutput.t54 gnd 0.055846f
C1383 CSoutput.t111 gnd 0.055846f
C1384 CSoutput.n113 gnd 0.431603f
C1385 CSoutput.n114 gnd 0.215866f
C1386 CSoutput.t85 gnd 0.055846f
C1387 CSoutput.t86 gnd 0.055846f
C1388 CSoutput.n115 gnd 0.431603f
C1389 CSoutput.n116 gnd 0.215866f
C1390 CSoutput.t75 gnd 0.055846f
C1391 CSoutput.t52 gnd 0.055846f
C1392 CSoutput.n117 gnd 0.431603f
C1393 CSoutput.n118 gnd 0.215866f
C1394 CSoutput.t33 gnd 0.055846f
C1395 CSoutput.t76 gnd 0.055846f
C1396 CSoutput.n119 gnd 0.431603f
C1397 CSoutput.n120 gnd 0.215866f
C1398 CSoutput.t74 gnd 0.055846f
C1399 CSoutput.t49 gnd 0.055846f
C1400 CSoutput.n121 gnd 0.431603f
C1401 CSoutput.n122 gnd 0.215866f
C1402 CSoutput.t31 gnd 0.055846f
C1403 CSoutput.t30 gnd 0.055846f
C1404 CSoutput.n123 gnd 0.431603f
C1405 CSoutput.n124 gnd 0.32191f
C1406 CSoutput.n125 gnd 0.453722f
C1407 CSoutput.n126 gnd 7.80723f
C1408 CSoutput.n128 gnd 0.79199f
C1409 CSoutput.n129 gnd 0.593993f
C1410 CSoutput.n130 gnd 0.79199f
C1411 CSoutput.n131 gnd 0.79199f
C1412 CSoutput.n132 gnd 2.13228f
C1413 CSoutput.n133 gnd 0.79199f
C1414 CSoutput.n134 gnd 0.79199f
C1415 CSoutput.t164 gnd 0.989988f
C1416 CSoutput.n135 gnd 0.79199f
C1417 CSoutput.n136 gnd 0.79199f
C1418 CSoutput.n140 gnd 0.79199f
C1419 CSoutput.n144 gnd 0.79199f
C1420 CSoutput.n145 gnd 0.79199f
C1421 CSoutput.n147 gnd 0.79199f
C1422 CSoutput.n152 gnd 0.79199f
C1423 CSoutput.n154 gnd 0.79199f
C1424 CSoutput.n155 gnd 0.79199f
C1425 CSoutput.n157 gnd 0.79199f
C1426 CSoutput.n158 gnd 0.79199f
C1427 CSoutput.n160 gnd 0.79199f
C1428 CSoutput.t153 gnd 13.234099f
C1429 CSoutput.n162 gnd 0.79199f
C1430 CSoutput.n163 gnd 0.593993f
C1431 CSoutput.n164 gnd 0.79199f
C1432 CSoutput.n165 gnd 0.79199f
C1433 CSoutput.n166 gnd 2.13228f
C1434 CSoutput.n167 gnd 0.79199f
C1435 CSoutput.n168 gnd 0.79199f
C1436 CSoutput.t152 gnd 0.989988f
C1437 CSoutput.n169 gnd 0.79199f
C1438 CSoutput.n170 gnd 0.79199f
C1439 CSoutput.n174 gnd 0.79199f
C1440 CSoutput.n178 gnd 0.79199f
C1441 CSoutput.n179 gnd 0.79199f
C1442 CSoutput.n181 gnd 0.79199f
C1443 CSoutput.n186 gnd 0.79199f
C1444 CSoutput.n188 gnd 0.79199f
C1445 CSoutput.n189 gnd 0.79199f
C1446 CSoutput.n191 gnd 0.79199f
C1447 CSoutput.n192 gnd 0.79199f
C1448 CSoutput.n194 gnd 0.79199f
C1449 CSoutput.n195 gnd 0.593993f
C1450 CSoutput.n197 gnd 0.79199f
C1451 CSoutput.n198 gnd 0.593993f
C1452 CSoutput.n199 gnd 0.79199f
C1453 CSoutput.n200 gnd 0.79199f
C1454 CSoutput.n201 gnd 2.13228f
C1455 CSoutput.n202 gnd 0.79199f
C1456 CSoutput.n203 gnd 0.79199f
C1457 CSoutput.t146 gnd 0.989988f
C1458 CSoutput.n204 gnd 0.79199f
C1459 CSoutput.n205 gnd 2.13228f
C1460 CSoutput.n207 gnd 0.79199f
C1461 CSoutput.n208 gnd 0.79199f
C1462 CSoutput.n210 gnd 0.79199f
C1463 CSoutput.n211 gnd 0.79199f
C1464 CSoutput.t154 gnd 13.0184f
C1465 CSoutput.t157 gnd 13.234099f
C1466 CSoutput.n217 gnd 2.48459f
C1467 CSoutput.n218 gnd 10.1213f
C1468 CSoutput.n219 gnd 10.5448f
C1469 CSoutput.n224 gnd 2.69148f
C1470 CSoutput.n230 gnd 0.79199f
C1471 CSoutput.n232 gnd 0.79199f
C1472 CSoutput.n234 gnd 0.79199f
C1473 CSoutput.n236 gnd 0.79199f
C1474 CSoutput.n238 gnd 0.79199f
C1475 CSoutput.n244 gnd 0.79199f
C1476 CSoutput.n251 gnd 1.453f
C1477 CSoutput.n252 gnd 1.453f
C1478 CSoutput.n253 gnd 0.79199f
C1479 CSoutput.n254 gnd 0.79199f
C1480 CSoutput.n256 gnd 0.593993f
C1481 CSoutput.n257 gnd 0.508701f
C1482 CSoutput.n259 gnd 0.593993f
C1483 CSoutput.n260 gnd 0.508701f
C1484 CSoutput.n261 gnd 0.593993f
C1485 CSoutput.n263 gnd 0.79199f
C1486 CSoutput.n265 gnd 2.13228f
C1487 CSoutput.n266 gnd 2.48459f
C1488 CSoutput.n267 gnd 9.30901f
C1489 CSoutput.n269 gnd 0.593993f
C1490 CSoutput.n270 gnd 1.52838f
C1491 CSoutput.n271 gnd 0.593993f
C1492 CSoutput.n273 gnd 0.79199f
C1493 CSoutput.n275 gnd 2.13228f
C1494 CSoutput.n276 gnd 4.64445f
C1495 CSoutput.t40 gnd 0.055846f
C1496 CSoutput.t94 gnd 0.055846f
C1497 CSoutput.n277 gnd 0.432374f
C1498 CSoutput.t56 gnd 0.055846f
C1499 CSoutput.t106 gnd 0.055846f
C1500 CSoutput.n278 gnd 0.431603f
C1501 CSoutput.n279 gnd 0.438077f
C1502 CSoutput.t87 gnd 0.055846f
C1503 CSoutput.t20 gnd 0.055846f
C1504 CSoutput.n280 gnd 0.431603f
C1505 CSoutput.n281 gnd 0.215866f
C1506 CSoutput.t48 gnd 0.055846f
C1507 CSoutput.t26 gnd 0.055846f
C1508 CSoutput.n282 gnd 0.431603f
C1509 CSoutput.n283 gnd 0.215866f
C1510 CSoutput.t65 gnd 0.055846f
C1511 CSoutput.t44 gnd 0.055846f
C1512 CSoutput.n284 gnd 0.431603f
C1513 CSoutput.n285 gnd 0.215866f
C1514 CSoutput.t97 gnd 0.055846f
C1515 CSoutput.t29 gnd 0.055846f
C1516 CSoutput.n286 gnd 0.431603f
C1517 CSoutput.n287 gnd 0.215866f
C1518 CSoutput.t79 gnd 0.055846f
C1519 CSoutput.t34 gnd 0.055846f
C1520 CSoutput.n288 gnd 0.431603f
C1521 CSoutput.n289 gnd 0.215866f
C1522 CSoutput.t89 gnd 0.055846f
C1523 CSoutput.t51 gnd 0.055846f
C1524 CSoutput.n290 gnd 0.431603f
C1525 CSoutput.n291 gnd 0.395848f
C1526 CSoutput.t62 gnd 0.055846f
C1527 CSoutput.t82 gnd 0.055846f
C1528 CSoutput.n292 gnd 0.432374f
C1529 CSoutput.t16 gnd 0.055846f
C1530 CSoutput.t46 gnd 0.055846f
C1531 CSoutput.n293 gnd 0.431603f
C1532 CSoutput.n294 gnd 0.438077f
C1533 CSoutput.t47 gnd 0.055846f
C1534 CSoutput.t101 gnd 0.055846f
C1535 CSoutput.n295 gnd 0.431603f
C1536 CSoutput.n296 gnd 0.215866f
C1537 CSoutput.t43 gnd 0.055846f
C1538 CSoutput.t45 gnd 0.055846f
C1539 CSoutput.n297 gnd 0.431603f
C1540 CSoutput.n298 gnd 0.215866f
C1541 CSoutput.t99 gnd 0.055846f
C1542 CSoutput.t100 gnd 0.055846f
C1543 CSoutput.n299 gnd 0.431603f
C1544 CSoutput.n300 gnd 0.215866f
C1545 CSoutput.t24 gnd 0.055846f
C1546 CSoutput.t84 gnd 0.055846f
C1547 CSoutput.n301 gnd 0.431603f
C1548 CSoutput.n302 gnd 0.215866f
C1549 CSoutput.t98 gnd 0.055846f
C1550 CSoutput.t23 gnd 0.055846f
C1551 CSoutput.n303 gnd 0.431603f
C1552 CSoutput.n304 gnd 0.215866f
C1553 CSoutput.t63 gnd 0.055846f
C1554 CSoutput.t83 gnd 0.055846f
C1555 CSoutput.n305 gnd 0.431603f
C1556 CSoutput.n306 gnd 0.32191f
C1557 CSoutput.n307 gnd 0.405927f
C1558 CSoutput.t72 gnd 0.055846f
C1559 CSoutput.t91 gnd 0.055846f
C1560 CSoutput.n308 gnd 0.432374f
C1561 CSoutput.t27 gnd 0.055846f
C1562 CSoutput.t60 gnd 0.055846f
C1563 CSoutput.n309 gnd 0.431603f
C1564 CSoutput.n310 gnd 0.438077f
C1565 CSoutput.t61 gnd 0.055846f
C1566 CSoutput.t109 gnd 0.055846f
C1567 CSoutput.n311 gnd 0.431603f
C1568 CSoutput.n312 gnd 0.215866f
C1569 CSoutput.t55 gnd 0.055846f
C1570 CSoutput.t57 gnd 0.055846f
C1571 CSoutput.n313 gnd 0.431603f
C1572 CSoutput.n314 gnd 0.215866f
C1573 CSoutput.t107 gnd 0.055846f
C1574 CSoutput.t108 gnd 0.055846f
C1575 CSoutput.n315 gnd 0.431603f
C1576 CSoutput.n316 gnd 0.215866f
C1577 CSoutput.t39 gnd 0.055846f
C1578 CSoutput.t95 gnd 0.055846f
C1579 CSoutput.n317 gnd 0.431603f
C1580 CSoutput.n318 gnd 0.215866f
C1581 CSoutput.t104 gnd 0.055846f
C1582 CSoutput.t35 gnd 0.055846f
C1583 CSoutput.n319 gnd 0.431603f
C1584 CSoutput.n320 gnd 0.215866f
C1585 CSoutput.t73 gnd 0.055846f
C1586 CSoutput.t92 gnd 0.055846f
C1587 CSoutput.n321 gnd 0.431602f
C1588 CSoutput.n322 gnd 0.321912f
C1589 CSoutput.n323 gnd 0.453722f
C1590 CSoutput.n324 gnd 11.4378f
C1591 CSoutput.t122 gnd 0.048865f
C1592 CSoutput.t128 gnd 0.048865f
C1593 CSoutput.n325 gnd 0.433232f
C1594 CSoutput.t130 gnd 0.048865f
C1595 CSoutput.t131 gnd 0.048865f
C1596 CSoutput.n326 gnd 0.431786f
C1597 CSoutput.n327 gnd 0.402344f
C1598 CSoutput.t121 gnd 0.048865f
C1599 CSoutput.t113 gnd 0.048865f
C1600 CSoutput.n328 gnd 0.431786f
C1601 CSoutput.n329 gnd 0.198337f
C1602 CSoutput.t116 gnd 0.048865f
C1603 CSoutput.t135 gnd 0.048865f
C1604 CSoutput.n330 gnd 0.431786f
C1605 CSoutput.n331 gnd 0.198337f
C1606 CSoutput.t114 gnd 0.048865f
C1607 CSoutput.t141 gnd 0.048865f
C1608 CSoutput.n332 gnd 0.431786f
C1609 CSoutput.n333 gnd 0.198337f
C1610 CSoutput.t13 gnd 0.048865f
C1611 CSoutput.t117 gnd 0.048865f
C1612 CSoutput.n334 gnd 0.431786f
C1613 CSoutput.n335 gnd 0.365773f
C1614 CSoutput.t137 gnd 0.048865f
C1615 CSoutput.t9 gnd 0.048865f
C1616 CSoutput.n336 gnd 0.433232f
C1617 CSoutput.t14 gnd 0.048865f
C1618 CSoutput.t8 gnd 0.048865f
C1619 CSoutput.n337 gnd 0.431786f
C1620 CSoutput.n338 gnd 0.402344f
C1621 CSoutput.t120 gnd 0.048865f
C1622 CSoutput.t142 gnd 0.048865f
C1623 CSoutput.n339 gnd 0.431786f
C1624 CSoutput.n340 gnd 0.198337f
C1625 CSoutput.t2 gnd 0.048865f
C1626 CSoutput.t6 gnd 0.048865f
C1627 CSoutput.n341 gnd 0.431786f
C1628 CSoutput.n342 gnd 0.198337f
C1629 CSoutput.t134 gnd 0.048865f
C1630 CSoutput.t139 gnd 0.048865f
C1631 CSoutput.n343 gnd 0.431786f
C1632 CSoutput.n344 gnd 0.198337f
C1633 CSoutput.t129 gnd 0.048865f
C1634 CSoutput.t132 gnd 0.048865f
C1635 CSoutput.n345 gnd 0.431786f
C1636 CSoutput.n346 gnd 0.301118f
C1637 CSoutput.n347 gnd 0.5595f
C1638 CSoutput.n348 gnd 11.5935f
C1639 CSoutput.t133 gnd 0.048865f
C1640 CSoutput.t11 gnd 0.048865f
C1641 CSoutput.n349 gnd 0.433232f
C1642 CSoutput.t115 gnd 0.048865f
C1643 CSoutput.t118 gnd 0.048865f
C1644 CSoutput.n350 gnd 0.431786f
C1645 CSoutput.n351 gnd 0.402344f
C1646 CSoutput.t136 gnd 0.048865f
C1647 CSoutput.t140 gnd 0.048865f
C1648 CSoutput.n352 gnd 0.431786f
C1649 CSoutput.n353 gnd 0.198337f
C1650 CSoutput.t127 gnd 0.048865f
C1651 CSoutput.t5 gnd 0.048865f
C1652 CSoutput.n354 gnd 0.431786f
C1653 CSoutput.n355 gnd 0.198337f
C1654 CSoutput.t124 gnd 0.048865f
C1655 CSoutput.t125 gnd 0.048865f
C1656 CSoutput.n356 gnd 0.431786f
C1657 CSoutput.n357 gnd 0.198337f
C1658 CSoutput.t123 gnd 0.048865f
C1659 CSoutput.t12 gnd 0.048865f
C1660 CSoutput.n358 gnd 0.431786f
C1661 CSoutput.n359 gnd 0.365773f
C1662 CSoutput.t10 gnd 0.048865f
C1663 CSoutput.t138 gnd 0.048865f
C1664 CSoutput.n360 gnd 0.433232f
C1665 CSoutput.t1 gnd 0.048865f
C1666 CSoutput.t3 gnd 0.048865f
C1667 CSoutput.n361 gnd 0.431786f
C1668 CSoutput.n362 gnd 0.402344f
C1669 CSoutput.t7 gnd 0.048865f
C1670 CSoutput.t119 gnd 0.048865f
C1671 CSoutput.n363 gnd 0.431786f
C1672 CSoutput.n364 gnd 0.198337f
C1673 CSoutput.t143 gnd 0.048865f
C1674 CSoutput.t4 gnd 0.048865f
C1675 CSoutput.n365 gnd 0.431786f
C1676 CSoutput.n366 gnd 0.198337f
C1677 CSoutput.t0 gnd 0.048865f
C1678 CSoutput.t112 gnd 0.048865f
C1679 CSoutput.n367 gnd 0.431786f
C1680 CSoutput.n368 gnd 0.198337f
C1681 CSoutput.t15 gnd 0.048865f
C1682 CSoutput.t126 gnd 0.048865f
C1683 CSoutput.n369 gnd 0.431786f
C1684 CSoutput.n370 gnd 0.301118f
C1685 CSoutput.n371 gnd 0.5595f
C1686 CSoutput.n372 gnd 6.51617f
C1687 CSoutput.n373 gnd 14.2994f
C1688 a_n7636_8799.n0 gnd 2.71862f
C1689 a_n7636_8799.n1 gnd 1.64714f
C1690 a_n7636_8799.n2 gnd 3.76849f
C1691 a_n7636_8799.n3 gnd 0.205533f
C1692 a_n7636_8799.n4 gnd 0.287271f
C1693 a_n7636_8799.n5 gnd 0.205533f
C1694 a_n7636_8799.n6 gnd 0.205533f
C1695 a_n7636_8799.n7 gnd 0.205533f
C1696 a_n7636_8799.n8 gnd 0.27078f
C1697 a_n7636_8799.n9 gnd 0.205533f
C1698 a_n7636_8799.n10 gnd 0.287271f
C1699 a_n7636_8799.n11 gnd 0.205533f
C1700 a_n7636_8799.n12 gnd 0.205533f
C1701 a_n7636_8799.n13 gnd 0.205533f
C1702 a_n7636_8799.n14 gnd 0.27078f
C1703 a_n7636_8799.n15 gnd 0.205533f
C1704 a_n7636_8799.n16 gnd 0.45021f
C1705 a_n7636_8799.n17 gnd 0.205533f
C1706 a_n7636_8799.n18 gnd 0.205533f
C1707 a_n7636_8799.n19 gnd 0.205533f
C1708 a_n7636_8799.n20 gnd 0.27078f
C1709 a_n7636_8799.n21 gnd 0.322163f
C1710 a_n7636_8799.n22 gnd 0.205533f
C1711 a_n7636_8799.n23 gnd 0.205533f
C1712 a_n7636_8799.n24 gnd 0.205533f
C1713 a_n7636_8799.n25 gnd 0.205533f
C1714 a_n7636_8799.n26 gnd 0.235888f
C1715 a_n7636_8799.n27 gnd 0.322163f
C1716 a_n7636_8799.n28 gnd 0.205533f
C1717 a_n7636_8799.n29 gnd 0.205533f
C1718 a_n7636_8799.n30 gnd 0.205533f
C1719 a_n7636_8799.n31 gnd 0.205533f
C1720 a_n7636_8799.n32 gnd 0.235888f
C1721 a_n7636_8799.n33 gnd 0.322163f
C1722 a_n7636_8799.n34 gnd 0.205533f
C1723 a_n7636_8799.n35 gnd 0.205533f
C1724 a_n7636_8799.n36 gnd 0.205533f
C1725 a_n7636_8799.n37 gnd 0.205533f
C1726 a_n7636_8799.n38 gnd 0.398827f
C1727 a_n7636_8799.n39 gnd 1.50639f
C1728 a_n7636_8799.n40 gnd 2.51925f
C1729 a_n7636_8799.n41 gnd 0.008525f
C1730 a_n7636_8799.n42 gnd 0.001144f
C1731 a_n7636_8799.n44 gnd 0.007655f
C1732 a_n7636_8799.n45 gnd 0.011571f
C1733 a_n7636_8799.n46 gnd 0.007958f
C1734 a_n7636_8799.n48 gnd 3.98e-19
C1735 a_n7636_8799.n49 gnd 0.008247f
C1736 a_n7636_8799.n50 gnd 0.01139f
C1737 a_n7636_8799.n51 gnd 0.007339f
C1738 a_n7636_8799.n52 gnd 0.008525f
C1739 a_n7636_8799.n53 gnd 0.001144f
C1740 a_n7636_8799.n55 gnd 0.007655f
C1741 a_n7636_8799.n56 gnd 0.011571f
C1742 a_n7636_8799.n57 gnd 0.007958f
C1743 a_n7636_8799.n59 gnd 3.98e-19
C1744 a_n7636_8799.n60 gnd 0.008247f
C1745 a_n7636_8799.n61 gnd 0.01139f
C1746 a_n7636_8799.n62 gnd 0.007339f
C1747 a_n7636_8799.n63 gnd 0.008525f
C1748 a_n7636_8799.n64 gnd 0.001144f
C1749 a_n7636_8799.n66 gnd 0.007655f
C1750 a_n7636_8799.n67 gnd 0.011571f
C1751 a_n7636_8799.n68 gnd 0.007958f
C1752 a_n7636_8799.n70 gnd 3.98e-19
C1753 a_n7636_8799.n71 gnd 0.008247f
C1754 a_n7636_8799.n72 gnd 0.01139f
C1755 a_n7636_8799.n73 gnd 0.007339f
C1756 a_n7636_8799.n74 gnd 0.001144f
C1757 a_n7636_8799.n76 gnd 0.007655f
C1758 a_n7636_8799.n77 gnd 0.011571f
C1759 a_n7636_8799.n78 gnd 0.007958f
C1760 a_n7636_8799.n80 gnd 3.98e-19
C1761 a_n7636_8799.n81 gnd 0.008247f
C1762 a_n7636_8799.n82 gnd 0.01139f
C1763 a_n7636_8799.n83 gnd 0.007339f
C1764 a_n7636_8799.n84 gnd 0.247442f
C1765 a_n7636_8799.n85 gnd 0.001144f
C1766 a_n7636_8799.n87 gnd 0.007655f
C1767 a_n7636_8799.n88 gnd 0.011571f
C1768 a_n7636_8799.n89 gnd 0.007958f
C1769 a_n7636_8799.n91 gnd 3.98e-19
C1770 a_n7636_8799.n92 gnd 0.008247f
C1771 a_n7636_8799.n93 gnd 0.01139f
C1772 a_n7636_8799.n94 gnd 0.007339f
C1773 a_n7636_8799.n95 gnd 0.247442f
C1774 a_n7636_8799.n96 gnd 0.001144f
C1775 a_n7636_8799.n98 gnd 0.007655f
C1776 a_n7636_8799.n99 gnd 0.011571f
C1777 a_n7636_8799.n100 gnd 0.007958f
C1778 a_n7636_8799.n102 gnd 3.98e-19
C1779 a_n7636_8799.n103 gnd 0.008247f
C1780 a_n7636_8799.n104 gnd 0.01139f
C1781 a_n7636_8799.n105 gnd 0.007339f
C1782 a_n7636_8799.n106 gnd 0.247442f
C1783 a_n7636_8799.t19 gnd 0.14256f
C1784 a_n7636_8799.t13 gnd 0.14256f
C1785 a_n7636_8799.t20 gnd 0.14256f
C1786 a_n7636_8799.n107 gnd 1.12439f
C1787 a_n7636_8799.t15 gnd 0.14256f
C1788 a_n7636_8799.t8 gnd 0.14256f
C1789 a_n7636_8799.n108 gnd 1.12439f
C1790 a_n7636_8799.t12 gnd 0.14256f
C1791 a_n7636_8799.t18 gnd 0.14256f
C1792 a_n7636_8799.n109 gnd 1.12254f
C1793 a_n7636_8799.t9 gnd 0.14256f
C1794 a_n7636_8799.t11 gnd 0.14256f
C1795 a_n7636_8799.n110 gnd 1.12254f
C1796 a_n7636_8799.t7 gnd 0.14256f
C1797 a_n7636_8799.t10 gnd 0.14256f
C1798 a_n7636_8799.n111 gnd 1.12254f
C1799 a_n7636_8799.n112 gnd 3.15297f
C1800 a_n7636_8799.t23 gnd 0.11088f
C1801 a_n7636_8799.t5 gnd 0.11088f
C1802 a_n7636_8799.n113 gnd 0.982662f
C1803 a_n7636_8799.t29 gnd 0.11088f
C1804 a_n7636_8799.t3 gnd 0.11088f
C1805 a_n7636_8799.n114 gnd 0.979773f
C1806 a_n7636_8799.t2 gnd 0.11088f
C1807 a_n7636_8799.t22 gnd 0.11088f
C1808 a_n7636_8799.n115 gnd 0.982661f
C1809 a_n7636_8799.t31 gnd 0.11088f
C1810 a_n7636_8799.t26 gnd 0.11088f
C1811 a_n7636_8799.n116 gnd 0.979772f
C1812 a_n7636_8799.t24 gnd 0.11088f
C1813 a_n7636_8799.t25 gnd 0.11088f
C1814 a_n7636_8799.n117 gnd 0.982661f
C1815 a_n7636_8799.t0 gnd 0.11088f
C1816 a_n7636_8799.t28 gnd 0.11088f
C1817 a_n7636_8799.n118 gnd 0.979772f
C1818 a_n7636_8799.t4 gnd 0.11088f
C1819 a_n7636_8799.t30 gnd 0.11088f
C1820 a_n7636_8799.n119 gnd 0.979773f
C1821 a_n7636_8799.t1 gnd 0.11088f
C1822 a_n7636_8799.t27 gnd 0.11088f
C1823 a_n7636_8799.n120 gnd 0.979773f
C1824 a_n7636_8799.t73 gnd 0.591119f
C1825 a_n7636_8799.n121 gnd 0.264275f
C1826 a_n7636_8799.t32 gnd 0.591119f
C1827 a_n7636_8799.t58 gnd 0.591119f
C1828 a_n7636_8799.n122 gnd 0.267549f
C1829 a_n7636_8799.t57 gnd 0.591119f
C1830 a_n7636_8799.t68 gnd 0.591119f
C1831 a_n7636_8799.t94 gnd 0.591119f
C1832 a_n7636_8799.n123 gnd 0.26961f
C1833 a_n7636_8799.t110 gnd 0.591119f
C1834 a_n7636_8799.t113 gnd 0.591119f
C1835 a_n7636_8799.n124 gnd 0.263213f
C1836 a_n7636_8799.t112 gnd 0.602307f
C1837 a_n7636_8799.n125 gnd 0.247823f
C1838 a_n7636_8799.n126 gnd 0.01166f
C1839 a_n7636_8799.t69 gnd 0.591119f
C1840 a_n7636_8799.n127 gnd 0.264005f
C1841 a_n7636_8799.n128 gnd 0.267534f
C1842 a_n7636_8799.t67 gnd 0.591119f
C1843 a_n7636_8799.n129 gnd 0.264094f
C1844 a_n7636_8799.n130 gnd 0.258778f
C1845 a_n7636_8799.t91 gnd 0.591119f
C1846 a_n7636_8799.n131 gnd 0.263847f
C1847 a_n7636_8799.n132 gnd 0.27004f
C1848 a_n7636_8799.t89 gnd 0.591119f
C1849 a_n7636_8799.n133 gnd 0.267418f
C1850 a_n7636_8799.n134 gnd 0.26353f
C1851 a_n7636_8799.t55 gnd 0.591119f
C1852 a_n7636_8799.n135 gnd 0.259095f
C1853 a_n7636_8799.t111 gnd 0.591119f
C1854 a_n7636_8799.n136 gnd 0.267533f
C1855 a_n7636_8799.t41 gnd 0.602297f
C1856 a_n7636_8799.t84 gnd 0.591119f
C1857 a_n7636_8799.n137 gnd 0.264275f
C1858 a_n7636_8799.t40 gnd 0.591119f
C1859 a_n7636_8799.t63 gnd 0.591119f
C1860 a_n7636_8799.n138 gnd 0.267549f
C1861 a_n7636_8799.t66 gnd 0.591119f
C1862 a_n7636_8799.t75 gnd 0.591119f
C1863 a_n7636_8799.t106 gnd 0.591119f
C1864 a_n7636_8799.n139 gnd 0.26961f
C1865 a_n7636_8799.t122 gnd 0.591119f
C1866 a_n7636_8799.t125 gnd 0.591119f
C1867 a_n7636_8799.n140 gnd 0.263213f
C1868 a_n7636_8799.t126 gnd 0.602307f
C1869 a_n7636_8799.n141 gnd 0.247823f
C1870 a_n7636_8799.n142 gnd 0.01166f
C1871 a_n7636_8799.t77 gnd 0.591119f
C1872 a_n7636_8799.n143 gnd 0.264005f
C1873 a_n7636_8799.n144 gnd 0.267534f
C1874 a_n7636_8799.t76 gnd 0.591119f
C1875 a_n7636_8799.n145 gnd 0.264094f
C1876 a_n7636_8799.n146 gnd 0.258778f
C1877 a_n7636_8799.t105 gnd 0.591119f
C1878 a_n7636_8799.n147 gnd 0.263847f
C1879 a_n7636_8799.n148 gnd 0.27004f
C1880 a_n7636_8799.t101 gnd 0.591119f
C1881 a_n7636_8799.n149 gnd 0.267418f
C1882 a_n7636_8799.n150 gnd 0.26353f
C1883 a_n7636_8799.t62 gnd 0.591119f
C1884 a_n7636_8799.n151 gnd 0.259095f
C1885 a_n7636_8799.t124 gnd 0.591119f
C1886 a_n7636_8799.n152 gnd 0.267533f
C1887 a_n7636_8799.t53 gnd 0.602297f
C1888 a_n7636_8799.n153 gnd 0.890291f
C1889 a_n7636_8799.t85 gnd 0.591119f
C1890 a_n7636_8799.n154 gnd 0.264275f
C1891 a_n7636_8799.t74 gnd 0.591119f
C1892 a_n7636_8799.t118 gnd 0.591119f
C1893 a_n7636_8799.n155 gnd 0.267549f
C1894 a_n7636_8799.t93 gnd 0.591119f
C1895 a_n7636_8799.t33 gnd 0.591119f
C1896 a_n7636_8799.t65 gnd 0.591119f
C1897 a_n7636_8799.n156 gnd 0.26961f
C1898 a_n7636_8799.t115 gnd 0.591119f
C1899 a_n7636_8799.t72 gnd 0.591119f
C1900 a_n7636_8799.n157 gnd 0.263213f
C1901 a_n7636_8799.t90 gnd 0.602307f
C1902 a_n7636_8799.n158 gnd 0.247823f
C1903 a_n7636_8799.n159 gnd 0.01166f
C1904 a_n7636_8799.t107 gnd 0.591119f
C1905 a_n7636_8799.n160 gnd 0.264005f
C1906 a_n7636_8799.n161 gnd 0.267534f
C1907 a_n7636_8799.t47 gnd 0.591119f
C1908 a_n7636_8799.n162 gnd 0.264094f
C1909 a_n7636_8799.n163 gnd 0.258778f
C1910 a_n7636_8799.t79 gnd 0.591119f
C1911 a_n7636_8799.n164 gnd 0.263847f
C1912 a_n7636_8799.n165 gnd 0.27004f
C1913 a_n7636_8799.t121 gnd 0.591119f
C1914 a_n7636_8799.n166 gnd 0.267418f
C1915 a_n7636_8799.n167 gnd 0.26353f
C1916 a_n7636_8799.t38 gnd 0.591119f
C1917 a_n7636_8799.n168 gnd 0.259095f
C1918 a_n7636_8799.t50 gnd 0.591119f
C1919 a_n7636_8799.n169 gnd 0.267533f
C1920 a_n7636_8799.t102 gnd 0.602297f
C1921 a_n7636_8799.n170 gnd 1.55447f
C1922 a_n7636_8799.t71 gnd 0.591119f
C1923 a_n7636_8799.t52 gnd 0.591119f
C1924 a_n7636_8799.t116 gnd 0.591119f
C1925 a_n7636_8799.n171 gnd 0.26714f
C1926 a_n7636_8799.t83 gnd 0.591119f
C1927 a_n7636_8799.t82 gnd 0.591119f
C1928 a_n7636_8799.t34 gnd 0.591119f
C1929 a_n7636_8799.n172 gnd 0.264094f
C1930 a_n7636_8799.t88 gnd 0.591119f
C1931 a_n7636_8799.t86 gnd 0.591119f
C1932 a_n7636_8799.t36 gnd 0.591119f
C1933 a_n7636_8799.n173 gnd 0.267549f
C1934 a_n7636_8799.t35 gnd 0.591119f
C1935 a_n7636_8799.t104 gnd 0.591119f
C1936 a_n7636_8799.t48 gnd 0.591119f
C1937 a_n7636_8799.n174 gnd 0.26353f
C1938 a_n7636_8799.t39 gnd 0.591119f
C1939 a_n7636_8799.t108 gnd 0.591119f
C1940 a_n7636_8799.t70 gnd 0.591119f
C1941 a_n7636_8799.n175 gnd 0.267533f
C1942 a_n7636_8799.t51 gnd 0.602307f
C1943 a_n7636_8799.n176 gnd 0.247823f
C1944 a_n7636_8799.n177 gnd 0.264275f
C1945 a_n7636_8799.n178 gnd 0.259095f
C1946 a_n7636_8799.n179 gnd 0.267418f
C1947 a_n7636_8799.n180 gnd 0.27004f
C1948 a_n7636_8799.n181 gnd 0.263847f
C1949 a_n7636_8799.n182 gnd 0.258778f
C1950 a_n7636_8799.n183 gnd 0.267534f
C1951 a_n7636_8799.n184 gnd 0.26961f
C1952 a_n7636_8799.n185 gnd 0.263213f
C1953 a_n7636_8799.n186 gnd 0.258619f
C1954 a_n7636_8799.t81 gnd 0.591119f
C1955 a_n7636_8799.t61 gnd 0.591119f
C1956 a_n7636_8799.t127 gnd 0.591119f
C1957 a_n7636_8799.n187 gnd 0.26714f
C1958 a_n7636_8799.t97 gnd 0.591119f
C1959 a_n7636_8799.t96 gnd 0.591119f
C1960 a_n7636_8799.t42 gnd 0.591119f
C1961 a_n7636_8799.n188 gnd 0.264094f
C1962 a_n7636_8799.t100 gnd 0.591119f
C1963 a_n7636_8799.t98 gnd 0.591119f
C1964 a_n7636_8799.t44 gnd 0.591119f
C1965 a_n7636_8799.n189 gnd 0.267549f
C1966 a_n7636_8799.t43 gnd 0.591119f
C1967 a_n7636_8799.t119 gnd 0.591119f
C1968 a_n7636_8799.t59 gnd 0.591119f
C1969 a_n7636_8799.n190 gnd 0.26353f
C1970 a_n7636_8799.t45 gnd 0.591119f
C1971 a_n7636_8799.t120 gnd 0.591119f
C1972 a_n7636_8799.t80 gnd 0.591119f
C1973 a_n7636_8799.n191 gnd 0.267533f
C1974 a_n7636_8799.t60 gnd 0.602307f
C1975 a_n7636_8799.n192 gnd 0.247823f
C1976 a_n7636_8799.n193 gnd 0.264275f
C1977 a_n7636_8799.n194 gnd 0.259095f
C1978 a_n7636_8799.n195 gnd 0.267418f
C1979 a_n7636_8799.n196 gnd 0.27004f
C1980 a_n7636_8799.n197 gnd 0.263847f
C1981 a_n7636_8799.n198 gnd 0.258778f
C1982 a_n7636_8799.n199 gnd 0.267534f
C1983 a_n7636_8799.n200 gnd 0.26961f
C1984 a_n7636_8799.n201 gnd 0.263213f
C1985 a_n7636_8799.n202 gnd 0.258619f
C1986 a_n7636_8799.n203 gnd 0.890291f
C1987 a_n7636_8799.t103 gnd 0.591119f
C1988 a_n7636_8799.t49 gnd 0.591119f
C1989 a_n7636_8799.t87 gnd 0.591119f
C1990 a_n7636_8799.n204 gnd 0.26714f
C1991 a_n7636_8799.t37 gnd 0.591119f
C1992 a_n7636_8799.t56 gnd 0.591119f
C1993 a_n7636_8799.t123 gnd 0.591119f
C1994 a_n7636_8799.n205 gnd 0.264094f
C1995 a_n7636_8799.t95 gnd 0.591119f
C1996 a_n7636_8799.t117 gnd 0.591119f
C1997 a_n7636_8799.t78 gnd 0.591119f
C1998 a_n7636_8799.n206 gnd 0.267549f
C1999 a_n7636_8799.t99 gnd 0.591119f
C2000 a_n7636_8799.t46 gnd 0.591119f
C2001 a_n7636_8799.t114 gnd 0.591119f
C2002 a_n7636_8799.n207 gnd 0.26353f
C2003 a_n7636_8799.t64 gnd 0.591119f
C2004 a_n7636_8799.t109 gnd 0.591119f
C2005 a_n7636_8799.t54 gnd 0.591119f
C2006 a_n7636_8799.n208 gnd 0.267533f
C2007 a_n7636_8799.t92 gnd 0.602307f
C2008 a_n7636_8799.n209 gnd 0.247823f
C2009 a_n7636_8799.n210 gnd 0.264275f
C2010 a_n7636_8799.n211 gnd 0.259095f
C2011 a_n7636_8799.n212 gnd 0.267418f
C2012 a_n7636_8799.n213 gnd 0.27004f
C2013 a_n7636_8799.n214 gnd 0.263847f
C2014 a_n7636_8799.n215 gnd 0.258778f
C2015 a_n7636_8799.n216 gnd 0.267534f
C2016 a_n7636_8799.n217 gnd 0.26961f
C2017 a_n7636_8799.n218 gnd 0.263213f
C2018 a_n7636_8799.n219 gnd 0.258619f
C2019 a_n7636_8799.n220 gnd 1.20614f
C2020 a_n7636_8799.n221 gnd 13.8223f
C2021 a_n7636_8799.n222 gnd 4.32613f
C2022 a_n7636_8799.n223 gnd 6.27519f
C2023 a_n7636_8799.t14 gnd 0.14256f
C2024 a_n7636_8799.t17 gnd 0.14256f
C2025 a_n7636_8799.n224 gnd 1.12254f
C2026 a_n7636_8799.t16 gnd 0.14256f
C2027 a_n7636_8799.t21 gnd 0.14256f
C2028 a_n7636_8799.n225 gnd 1.12254f
C2029 a_n7636_8799.n226 gnd 1.00902f
C2030 a_n7636_8799.n227 gnd 1.12254f
C2031 a_n7636_8799.t6 gnd 0.14256f
C2032 vdd.t230 gnd 0.037018f
C2033 vdd.t213 gnd 0.037018f
C2034 vdd.n0 gnd 0.291968f
C2035 vdd.t195 gnd 0.037018f
C2036 vdd.t225 gnd 0.037018f
C2037 vdd.n1 gnd 0.291486f
C2038 vdd.n2 gnd 0.268806f
C2039 vdd.t210 gnd 0.037018f
C2040 vdd.t234 gnd 0.037018f
C2041 vdd.n3 gnd 0.291486f
C2042 vdd.n4 gnd 0.135945f
C2043 vdd.t236 gnd 0.037018f
C2044 vdd.t218 gnd 0.037018f
C2045 vdd.n5 gnd 0.291486f
C2046 vdd.n6 gnd 0.127559f
C2047 vdd.t239 gnd 0.037018f
C2048 vdd.t208 gnd 0.037018f
C2049 vdd.n7 gnd 0.291968f
C2050 vdd.t216 gnd 0.037018f
C2051 vdd.t232 gnd 0.037018f
C2052 vdd.n8 gnd 0.291486f
C2053 vdd.n9 gnd 0.268806f
C2054 vdd.t223 gnd 0.037018f
C2055 vdd.t198 gnd 0.037018f
C2056 vdd.n10 gnd 0.291486f
C2057 vdd.n11 gnd 0.135945f
C2058 vdd.t205 gnd 0.037018f
C2059 vdd.t221 gnd 0.037018f
C2060 vdd.n12 gnd 0.291486f
C2061 vdd.n13 gnd 0.127559f
C2062 vdd.n14 gnd 0.090182f
C2063 vdd.t253 gnd 0.020566f
C2064 vdd.t175 gnd 0.020566f
C2065 vdd.n15 gnd 0.189298f
C2066 vdd.t117 gnd 0.020566f
C2067 vdd.t249 gnd 0.020566f
C2068 vdd.n16 gnd 0.188744f
C2069 vdd.n17 gnd 0.328474f
C2070 vdd.t247 gnd 0.020566f
C2071 vdd.t144 gnd 0.020566f
C2072 vdd.n18 gnd 0.188744f
C2073 vdd.n19 gnd 0.135894f
C2074 vdd.t118 gnd 0.020566f
C2075 vdd.t174 gnd 0.020566f
C2076 vdd.n20 gnd 0.189298f
C2077 vdd.t254 gnd 0.020566f
C2078 vdd.t122 gnd 0.020566f
C2079 vdd.n21 gnd 0.188744f
C2080 vdd.n22 gnd 0.328474f
C2081 vdd.t176 gnd 0.020566f
C2082 vdd.t248 gnd 0.020566f
C2083 vdd.n23 gnd 0.188744f
C2084 vdd.n24 gnd 0.135894f
C2085 vdd.t250 gnd 0.020566f
C2086 vdd.t145 gnd 0.020566f
C2087 vdd.n25 gnd 0.188744f
C2088 vdd.t251 gnd 0.020566f
C2089 vdd.t252 gnd 0.020566f
C2090 vdd.n26 gnd 0.188744f
C2091 vdd.n27 gnd 21.5184f
C2092 vdd.n28 gnd 7.98329f
C2093 vdd.n29 gnd 0.005609f
C2094 vdd.n30 gnd 0.005205f
C2095 vdd.n31 gnd 0.002879f
C2096 vdd.n32 gnd 0.006611f
C2097 vdd.n33 gnd 0.002797f
C2098 vdd.n34 gnd 0.002961f
C2099 vdd.n35 gnd 0.005205f
C2100 vdd.n36 gnd 0.002797f
C2101 vdd.n37 gnd 0.006611f
C2102 vdd.n38 gnd 0.002961f
C2103 vdd.n39 gnd 0.005205f
C2104 vdd.n40 gnd 0.002797f
C2105 vdd.n41 gnd 0.004958f
C2106 vdd.n42 gnd 0.004973f
C2107 vdd.t187 gnd 0.014203f
C2108 vdd.n43 gnd 0.031601f
C2109 vdd.n44 gnd 0.164461f
C2110 vdd.n45 gnd 0.002797f
C2111 vdd.n46 gnd 0.002961f
C2112 vdd.n47 gnd 0.006611f
C2113 vdd.n48 gnd 0.006611f
C2114 vdd.n49 gnd 0.002961f
C2115 vdd.n50 gnd 0.002797f
C2116 vdd.n51 gnd 0.005205f
C2117 vdd.n52 gnd 0.005205f
C2118 vdd.n53 gnd 0.002797f
C2119 vdd.n54 gnd 0.002961f
C2120 vdd.n55 gnd 0.006611f
C2121 vdd.n56 gnd 0.006611f
C2122 vdd.n57 gnd 0.002961f
C2123 vdd.n58 gnd 0.002797f
C2124 vdd.n59 gnd 0.005205f
C2125 vdd.n60 gnd 0.005205f
C2126 vdd.n61 gnd 0.002797f
C2127 vdd.n62 gnd 0.002961f
C2128 vdd.n63 gnd 0.006611f
C2129 vdd.n64 gnd 0.006611f
C2130 vdd.n65 gnd 0.01563f
C2131 vdd.n66 gnd 0.002879f
C2132 vdd.n67 gnd 0.002797f
C2133 vdd.n68 gnd 0.013453f
C2134 vdd.n69 gnd 0.009392f
C2135 vdd.t156 gnd 0.032905f
C2136 vdd.t137 gnd 0.032905f
C2137 vdd.n70 gnd 0.226146f
C2138 vdd.n71 gnd 0.177829f
C2139 vdd.t107 gnd 0.032905f
C2140 vdd.t257 gnd 0.032905f
C2141 vdd.n72 gnd 0.226146f
C2142 vdd.n73 gnd 0.143507f
C2143 vdd.t143 gnd 0.032905f
C2144 vdd.t125 gnd 0.032905f
C2145 vdd.n74 gnd 0.226146f
C2146 vdd.n75 gnd 0.143507f
C2147 vdd.t171 gnd 0.032905f
C2148 vdd.t141 gnd 0.032905f
C2149 vdd.n76 gnd 0.226146f
C2150 vdd.n77 gnd 0.143507f
C2151 vdd.t99 gnd 0.032905f
C2152 vdd.t264 gnd 0.032905f
C2153 vdd.n78 gnd 0.226146f
C2154 vdd.n79 gnd 0.143507f
C2155 vdd.t260 gnd 0.032905f
C2156 vdd.t95 gnd 0.032905f
C2157 vdd.n80 gnd 0.226146f
C2158 vdd.n81 gnd 0.143507f
C2159 vdd.t128 gnd 0.032905f
C2160 vdd.t10 gnd 0.032905f
C2161 vdd.n82 gnd 0.226146f
C2162 vdd.n83 gnd 0.143507f
C2163 vdd.n84 gnd 0.005609f
C2164 vdd.n85 gnd 0.005205f
C2165 vdd.n86 gnd 0.002879f
C2166 vdd.n87 gnd 0.006611f
C2167 vdd.n88 gnd 0.002797f
C2168 vdd.n89 gnd 0.002961f
C2169 vdd.n90 gnd 0.005205f
C2170 vdd.n91 gnd 0.002797f
C2171 vdd.n92 gnd 0.006611f
C2172 vdd.n93 gnd 0.002961f
C2173 vdd.n94 gnd 0.005205f
C2174 vdd.n95 gnd 0.002797f
C2175 vdd.n96 gnd 0.004958f
C2176 vdd.n97 gnd 0.004973f
C2177 vdd.t151 gnd 0.014203f
C2178 vdd.n98 gnd 0.031601f
C2179 vdd.n99 gnd 0.164461f
C2180 vdd.n100 gnd 0.002797f
C2181 vdd.n101 gnd 0.002961f
C2182 vdd.n102 gnd 0.006611f
C2183 vdd.n103 gnd 0.006611f
C2184 vdd.n104 gnd 0.002961f
C2185 vdd.n105 gnd 0.002797f
C2186 vdd.n106 gnd 0.005205f
C2187 vdd.n107 gnd 0.005205f
C2188 vdd.n108 gnd 0.002797f
C2189 vdd.n109 gnd 0.002961f
C2190 vdd.n110 gnd 0.006611f
C2191 vdd.n111 gnd 0.006611f
C2192 vdd.n112 gnd 0.002961f
C2193 vdd.n113 gnd 0.002797f
C2194 vdd.n114 gnd 0.005205f
C2195 vdd.n115 gnd 0.005205f
C2196 vdd.n116 gnd 0.002797f
C2197 vdd.n117 gnd 0.002961f
C2198 vdd.n118 gnd 0.006611f
C2199 vdd.n119 gnd 0.006611f
C2200 vdd.n120 gnd 0.01563f
C2201 vdd.n121 gnd 0.002879f
C2202 vdd.n122 gnd 0.002797f
C2203 vdd.n123 gnd 0.013453f
C2204 vdd.n124 gnd 0.009098f
C2205 vdd.n125 gnd 0.10677f
C2206 vdd.n126 gnd 0.005609f
C2207 vdd.n127 gnd 0.005205f
C2208 vdd.n128 gnd 0.002879f
C2209 vdd.n129 gnd 0.006611f
C2210 vdd.n130 gnd 0.002797f
C2211 vdd.n131 gnd 0.002961f
C2212 vdd.n132 gnd 0.005205f
C2213 vdd.n133 gnd 0.002797f
C2214 vdd.n134 gnd 0.006611f
C2215 vdd.n135 gnd 0.002961f
C2216 vdd.n136 gnd 0.005205f
C2217 vdd.n137 gnd 0.002797f
C2218 vdd.n138 gnd 0.004958f
C2219 vdd.n139 gnd 0.004973f
C2220 vdd.t162 gnd 0.014203f
C2221 vdd.n140 gnd 0.031601f
C2222 vdd.n141 gnd 0.164461f
C2223 vdd.n142 gnd 0.002797f
C2224 vdd.n143 gnd 0.002961f
C2225 vdd.n144 gnd 0.006611f
C2226 vdd.n145 gnd 0.006611f
C2227 vdd.n146 gnd 0.002961f
C2228 vdd.n147 gnd 0.002797f
C2229 vdd.n148 gnd 0.005205f
C2230 vdd.n149 gnd 0.005205f
C2231 vdd.n150 gnd 0.002797f
C2232 vdd.n151 gnd 0.002961f
C2233 vdd.n152 gnd 0.006611f
C2234 vdd.n153 gnd 0.006611f
C2235 vdd.n154 gnd 0.002961f
C2236 vdd.n155 gnd 0.002797f
C2237 vdd.n156 gnd 0.005205f
C2238 vdd.n157 gnd 0.005205f
C2239 vdd.n158 gnd 0.002797f
C2240 vdd.n159 gnd 0.002961f
C2241 vdd.n160 gnd 0.006611f
C2242 vdd.n161 gnd 0.006611f
C2243 vdd.n162 gnd 0.01563f
C2244 vdd.n163 gnd 0.002879f
C2245 vdd.n164 gnd 0.002797f
C2246 vdd.n165 gnd 0.013453f
C2247 vdd.n166 gnd 0.009392f
C2248 vdd.t182 gnd 0.032905f
C2249 vdd.t164 gnd 0.032905f
C2250 vdd.n167 gnd 0.226146f
C2251 vdd.n168 gnd 0.177829f
C2252 vdd.t103 gnd 0.032905f
C2253 vdd.t101 gnd 0.032905f
C2254 vdd.n169 gnd 0.226146f
C2255 vdd.n170 gnd 0.143507f
C2256 vdd.t262 gnd 0.032905f
C2257 vdd.t12 gnd 0.032905f
C2258 vdd.n171 gnd 0.226146f
C2259 vdd.n172 gnd 0.143507f
C2260 vdd.t97 gnd 0.032905f
C2261 vdd.t180 gnd 0.032905f
C2262 vdd.n173 gnd 0.226146f
C2263 vdd.n174 gnd 0.143507f
C2264 vdd.t116 gnd 0.032905f
C2265 vdd.t255 gnd 0.032905f
C2266 vdd.n175 gnd 0.226146f
C2267 vdd.n176 gnd 0.143507f
C2268 vdd.t265 gnd 0.032905f
C2269 vdd.t1 gnd 0.032905f
C2270 vdd.n177 gnd 0.226146f
C2271 vdd.n178 gnd 0.143507f
C2272 vdd.t242 gnd 0.032905f
C2273 vdd.t160 gnd 0.032905f
C2274 vdd.n179 gnd 0.226146f
C2275 vdd.n180 gnd 0.143507f
C2276 vdd.n181 gnd 0.005609f
C2277 vdd.n182 gnd 0.005205f
C2278 vdd.n183 gnd 0.002879f
C2279 vdd.n184 gnd 0.006611f
C2280 vdd.n185 gnd 0.002797f
C2281 vdd.n186 gnd 0.002961f
C2282 vdd.n187 gnd 0.005205f
C2283 vdd.n188 gnd 0.002797f
C2284 vdd.n189 gnd 0.006611f
C2285 vdd.n190 gnd 0.002961f
C2286 vdd.n191 gnd 0.005205f
C2287 vdd.n192 gnd 0.002797f
C2288 vdd.n193 gnd 0.004958f
C2289 vdd.n194 gnd 0.004973f
C2290 vdd.t191 gnd 0.014203f
C2291 vdd.n195 gnd 0.031601f
C2292 vdd.n196 gnd 0.164461f
C2293 vdd.n197 gnd 0.002797f
C2294 vdd.n198 gnd 0.002961f
C2295 vdd.n199 gnd 0.006611f
C2296 vdd.n200 gnd 0.006611f
C2297 vdd.n201 gnd 0.002961f
C2298 vdd.n202 gnd 0.002797f
C2299 vdd.n203 gnd 0.005205f
C2300 vdd.n204 gnd 0.005205f
C2301 vdd.n205 gnd 0.002797f
C2302 vdd.n206 gnd 0.002961f
C2303 vdd.n207 gnd 0.006611f
C2304 vdd.n208 gnd 0.006611f
C2305 vdd.n209 gnd 0.002961f
C2306 vdd.n210 gnd 0.002797f
C2307 vdd.n211 gnd 0.005205f
C2308 vdd.n212 gnd 0.005205f
C2309 vdd.n213 gnd 0.002797f
C2310 vdd.n214 gnd 0.002961f
C2311 vdd.n215 gnd 0.006611f
C2312 vdd.n216 gnd 0.006611f
C2313 vdd.n217 gnd 0.01563f
C2314 vdd.n218 gnd 0.002879f
C2315 vdd.n219 gnd 0.002797f
C2316 vdd.n220 gnd 0.013453f
C2317 vdd.n221 gnd 0.009098f
C2318 vdd.n222 gnd 0.063517f
C2319 vdd.n223 gnd 0.22887f
C2320 vdd.n224 gnd 0.005609f
C2321 vdd.n225 gnd 0.005205f
C2322 vdd.n226 gnd 0.002879f
C2323 vdd.n227 gnd 0.006611f
C2324 vdd.n228 gnd 0.002797f
C2325 vdd.n229 gnd 0.002961f
C2326 vdd.n230 gnd 0.005205f
C2327 vdd.n231 gnd 0.002797f
C2328 vdd.n232 gnd 0.006611f
C2329 vdd.n233 gnd 0.002961f
C2330 vdd.n234 gnd 0.005205f
C2331 vdd.n235 gnd 0.002797f
C2332 vdd.n236 gnd 0.004958f
C2333 vdd.n237 gnd 0.004973f
C2334 vdd.t168 gnd 0.014203f
C2335 vdd.n238 gnd 0.031601f
C2336 vdd.n239 gnd 0.164461f
C2337 vdd.n240 gnd 0.002797f
C2338 vdd.n241 gnd 0.002961f
C2339 vdd.n242 gnd 0.006611f
C2340 vdd.n243 gnd 0.006611f
C2341 vdd.n244 gnd 0.002961f
C2342 vdd.n245 gnd 0.002797f
C2343 vdd.n246 gnd 0.005205f
C2344 vdd.n247 gnd 0.005205f
C2345 vdd.n248 gnd 0.002797f
C2346 vdd.n249 gnd 0.002961f
C2347 vdd.n250 gnd 0.006611f
C2348 vdd.n251 gnd 0.006611f
C2349 vdd.n252 gnd 0.002961f
C2350 vdd.n253 gnd 0.002797f
C2351 vdd.n254 gnd 0.005205f
C2352 vdd.n255 gnd 0.005205f
C2353 vdd.n256 gnd 0.002797f
C2354 vdd.n257 gnd 0.002961f
C2355 vdd.n258 gnd 0.006611f
C2356 vdd.n259 gnd 0.006611f
C2357 vdd.n260 gnd 0.01563f
C2358 vdd.n261 gnd 0.002879f
C2359 vdd.n262 gnd 0.002797f
C2360 vdd.n263 gnd 0.013453f
C2361 vdd.n264 gnd 0.009392f
C2362 vdd.t3 gnd 0.032905f
C2363 vdd.t163 gnd 0.032905f
C2364 vdd.n265 gnd 0.226146f
C2365 vdd.n266 gnd 0.177829f
C2366 vdd.t115 gnd 0.032905f
C2367 vdd.t114 gnd 0.032905f
C2368 vdd.n267 gnd 0.226146f
C2369 vdd.n268 gnd 0.143507f
C2370 vdd.t94 gnd 0.032905f
C2371 vdd.t112 gnd 0.032905f
C2372 vdd.n269 gnd 0.226146f
C2373 vdd.n270 gnd 0.143507f
C2374 vdd.t135 gnd 0.032905f
C2375 vdd.t159 gnd 0.032905f
C2376 vdd.n271 gnd 0.226146f
C2377 vdd.n272 gnd 0.143507f
C2378 vdd.t154 gnd 0.032905f
C2379 vdd.t184 gnd 0.032905f
C2380 vdd.n273 gnd 0.226146f
C2381 vdd.n274 gnd 0.143507f
C2382 vdd.t106 gnd 0.032905f
C2383 vdd.t104 gnd 0.032905f
C2384 vdd.n275 gnd 0.226146f
C2385 vdd.n276 gnd 0.143507f
C2386 vdd.t127 gnd 0.032905f
C2387 vdd.t167 gnd 0.032905f
C2388 vdd.n277 gnd 0.226146f
C2389 vdd.n278 gnd 0.143507f
C2390 vdd.n279 gnd 0.005609f
C2391 vdd.n280 gnd 0.005205f
C2392 vdd.n281 gnd 0.002879f
C2393 vdd.n282 gnd 0.006611f
C2394 vdd.n283 gnd 0.002797f
C2395 vdd.n284 gnd 0.002961f
C2396 vdd.n285 gnd 0.005205f
C2397 vdd.n286 gnd 0.002797f
C2398 vdd.n287 gnd 0.006611f
C2399 vdd.n288 gnd 0.002961f
C2400 vdd.n289 gnd 0.005205f
C2401 vdd.n290 gnd 0.002797f
C2402 vdd.n291 gnd 0.004958f
C2403 vdd.n292 gnd 0.004973f
C2404 vdd.t244 gnd 0.014203f
C2405 vdd.n293 gnd 0.031601f
C2406 vdd.n294 gnd 0.164461f
C2407 vdd.n295 gnd 0.002797f
C2408 vdd.n296 gnd 0.002961f
C2409 vdd.n297 gnd 0.006611f
C2410 vdd.n298 gnd 0.006611f
C2411 vdd.n299 gnd 0.002961f
C2412 vdd.n300 gnd 0.002797f
C2413 vdd.n301 gnd 0.005205f
C2414 vdd.n302 gnd 0.005205f
C2415 vdd.n303 gnd 0.002797f
C2416 vdd.n304 gnd 0.002961f
C2417 vdd.n305 gnd 0.006611f
C2418 vdd.n306 gnd 0.006611f
C2419 vdd.n307 gnd 0.002961f
C2420 vdd.n308 gnd 0.002797f
C2421 vdd.n309 gnd 0.005205f
C2422 vdd.n310 gnd 0.005205f
C2423 vdd.n311 gnd 0.002797f
C2424 vdd.n312 gnd 0.002961f
C2425 vdd.n313 gnd 0.006611f
C2426 vdd.n314 gnd 0.006611f
C2427 vdd.n315 gnd 0.01563f
C2428 vdd.n316 gnd 0.002879f
C2429 vdd.n317 gnd 0.002797f
C2430 vdd.n318 gnd 0.013453f
C2431 vdd.n319 gnd 0.009098f
C2432 vdd.n320 gnd 0.063517f
C2433 vdd.n321 gnd 0.256304f
C2434 vdd.n322 gnd 0.007855f
C2435 vdd.n323 gnd 0.01022f
C2436 vdd.n324 gnd 0.008226f
C2437 vdd.n325 gnd 0.008226f
C2438 vdd.n326 gnd 0.01022f
C2439 vdd.n327 gnd 0.01022f
C2440 vdd.n328 gnd 0.746807f
C2441 vdd.n329 gnd 0.01022f
C2442 vdd.n330 gnd 0.01022f
C2443 vdd.n331 gnd 0.01022f
C2444 vdd.n332 gnd 0.809476f
C2445 vdd.n333 gnd 0.01022f
C2446 vdd.n334 gnd 0.01022f
C2447 vdd.n335 gnd 0.01022f
C2448 vdd.n336 gnd 0.01022f
C2449 vdd.n337 gnd 0.008226f
C2450 vdd.n338 gnd 0.01022f
C2451 vdd.t183 gnd 0.522243f
C2452 vdd.n339 gnd 0.01022f
C2453 vdd.n340 gnd 0.01022f
C2454 vdd.n341 gnd 0.01022f
C2455 vdd.t0 gnd 0.522243f
C2456 vdd.n342 gnd 0.01022f
C2457 vdd.n343 gnd 0.01022f
C2458 vdd.n344 gnd 0.01022f
C2459 vdd.n345 gnd 0.01022f
C2460 vdd.n346 gnd 0.01022f
C2461 vdd.n347 gnd 0.008226f
C2462 vdd.n348 gnd 0.01022f
C2463 vdd.n349 gnd 0.590134f
C2464 vdd.n350 gnd 0.01022f
C2465 vdd.n351 gnd 0.01022f
C2466 vdd.n352 gnd 0.01022f
C2467 vdd.t9 gnd 0.522243f
C2468 vdd.n353 gnd 0.01022f
C2469 vdd.n354 gnd 0.01022f
C2470 vdd.n355 gnd 0.01022f
C2471 vdd.n356 gnd 0.01022f
C2472 vdd.n357 gnd 0.01022f
C2473 vdd.n358 gnd 0.008226f
C2474 vdd.n359 gnd 0.01022f
C2475 vdd.t150 gnd 0.522243f
C2476 vdd.n360 gnd 0.01022f
C2477 vdd.n361 gnd 0.01022f
C2478 vdd.n362 gnd 0.01022f
C2479 vdd.n363 gnd 0.88259f
C2480 vdd.n364 gnd 0.01022f
C2481 vdd.n365 gnd 0.01022f
C2482 vdd.n366 gnd 0.01022f
C2483 vdd.n367 gnd 0.01022f
C2484 vdd.n368 gnd 0.01022f
C2485 vdd.n369 gnd 0.006828f
C2486 vdd.n370 gnd 0.023274f
C2487 vdd.t51 gnd 0.522243f
C2488 vdd.n371 gnd 0.01022f
C2489 vdd.n372 gnd 0.023274f
C2490 vdd.n404 gnd 0.01022f
C2491 vdd.t53 gnd 0.125739f
C2492 vdd.t52 gnd 0.13438f
C2493 vdd.t50 gnd 0.164213f
C2494 vdd.n405 gnd 0.210498f
C2495 vdd.n406 gnd 0.177679f
C2496 vdd.n407 gnd 0.013491f
C2497 vdd.n408 gnd 0.01022f
C2498 vdd.n409 gnd 0.008226f
C2499 vdd.n410 gnd 0.01022f
C2500 vdd.n411 gnd 0.008226f
C2501 vdd.n412 gnd 0.01022f
C2502 vdd.n413 gnd 0.008226f
C2503 vdd.n414 gnd 0.01022f
C2504 vdd.n415 gnd 0.008226f
C2505 vdd.n416 gnd 0.01022f
C2506 vdd.n417 gnd 0.008226f
C2507 vdd.n418 gnd 0.01022f
C2508 vdd.t86 gnd 0.125739f
C2509 vdd.t85 gnd 0.13438f
C2510 vdd.t84 gnd 0.164213f
C2511 vdd.n419 gnd 0.210498f
C2512 vdd.n420 gnd 0.177679f
C2513 vdd.n421 gnd 0.008226f
C2514 vdd.n422 gnd 0.01022f
C2515 vdd.n423 gnd 0.008226f
C2516 vdd.n424 gnd 0.01022f
C2517 vdd.n425 gnd 0.008226f
C2518 vdd.n426 gnd 0.01022f
C2519 vdd.n427 gnd 0.008226f
C2520 vdd.n428 gnd 0.01022f
C2521 vdd.n429 gnd 0.008226f
C2522 vdd.n430 gnd 0.01022f
C2523 vdd.t92 gnd 0.125739f
C2524 vdd.t91 gnd 0.13438f
C2525 vdd.t90 gnd 0.164213f
C2526 vdd.n431 gnd 0.210498f
C2527 vdd.n432 gnd 0.177679f
C2528 vdd.n433 gnd 0.017604f
C2529 vdd.n434 gnd 0.01022f
C2530 vdd.n435 gnd 0.008226f
C2531 vdd.n436 gnd 0.01022f
C2532 vdd.n437 gnd 0.008226f
C2533 vdd.n438 gnd 0.01022f
C2534 vdd.n439 gnd 0.008226f
C2535 vdd.n440 gnd 0.01022f
C2536 vdd.n441 gnd 0.008226f
C2537 vdd.n442 gnd 0.01022f
C2538 vdd.n443 gnd 0.023274f
C2539 vdd.n444 gnd 0.023433f
C2540 vdd.n445 gnd 0.023433f
C2541 vdd.n446 gnd 0.006828f
C2542 vdd.n447 gnd 0.008226f
C2543 vdd.n448 gnd 0.01022f
C2544 vdd.n449 gnd 0.01022f
C2545 vdd.n450 gnd 0.008226f
C2546 vdd.n451 gnd 0.01022f
C2547 vdd.n452 gnd 0.01022f
C2548 vdd.n453 gnd 0.01022f
C2549 vdd.n454 gnd 0.01022f
C2550 vdd.n455 gnd 0.01022f
C2551 vdd.n456 gnd 0.008226f
C2552 vdd.n457 gnd 0.008226f
C2553 vdd.n458 gnd 0.01022f
C2554 vdd.n459 gnd 0.01022f
C2555 vdd.n460 gnd 0.008226f
C2556 vdd.n461 gnd 0.01022f
C2557 vdd.n462 gnd 0.01022f
C2558 vdd.n463 gnd 0.01022f
C2559 vdd.n464 gnd 0.01022f
C2560 vdd.n465 gnd 0.01022f
C2561 vdd.n466 gnd 0.008226f
C2562 vdd.n467 gnd 0.008226f
C2563 vdd.n468 gnd 0.01022f
C2564 vdd.n469 gnd 0.01022f
C2565 vdd.n470 gnd 0.008226f
C2566 vdd.n471 gnd 0.01022f
C2567 vdd.n472 gnd 0.01022f
C2568 vdd.n473 gnd 0.01022f
C2569 vdd.n474 gnd 0.01022f
C2570 vdd.n475 gnd 0.01022f
C2571 vdd.n476 gnd 0.008226f
C2572 vdd.n477 gnd 0.008226f
C2573 vdd.n478 gnd 0.01022f
C2574 vdd.n479 gnd 0.01022f
C2575 vdd.n480 gnd 0.008226f
C2576 vdd.n481 gnd 0.01022f
C2577 vdd.n482 gnd 0.01022f
C2578 vdd.n483 gnd 0.01022f
C2579 vdd.n484 gnd 0.01022f
C2580 vdd.n485 gnd 0.01022f
C2581 vdd.n486 gnd 0.008226f
C2582 vdd.n487 gnd 0.008226f
C2583 vdd.n488 gnd 0.01022f
C2584 vdd.n489 gnd 0.01022f
C2585 vdd.n490 gnd 0.006869f
C2586 vdd.n491 gnd 0.01022f
C2587 vdd.n492 gnd 0.01022f
C2588 vdd.n493 gnd 0.01022f
C2589 vdd.n494 gnd 0.01022f
C2590 vdd.n495 gnd 0.01022f
C2591 vdd.n496 gnd 0.006869f
C2592 vdd.n497 gnd 0.008226f
C2593 vdd.n498 gnd 0.01022f
C2594 vdd.n499 gnd 0.01022f
C2595 vdd.n500 gnd 0.008226f
C2596 vdd.n501 gnd 0.01022f
C2597 vdd.n502 gnd 0.01022f
C2598 vdd.n503 gnd 0.01022f
C2599 vdd.n504 gnd 0.01022f
C2600 vdd.n505 gnd 0.01022f
C2601 vdd.n506 gnd 0.008226f
C2602 vdd.n507 gnd 0.008226f
C2603 vdd.n508 gnd 0.01022f
C2604 vdd.n509 gnd 0.01022f
C2605 vdd.n510 gnd 0.008226f
C2606 vdd.n511 gnd 0.01022f
C2607 vdd.n512 gnd 0.01022f
C2608 vdd.n513 gnd 0.01022f
C2609 vdd.n514 gnd 0.01022f
C2610 vdd.n515 gnd 0.01022f
C2611 vdd.n516 gnd 0.008226f
C2612 vdd.n517 gnd 0.008226f
C2613 vdd.n518 gnd 0.01022f
C2614 vdd.n519 gnd 0.01022f
C2615 vdd.n520 gnd 0.008226f
C2616 vdd.n521 gnd 0.01022f
C2617 vdd.n522 gnd 0.01022f
C2618 vdd.n523 gnd 0.01022f
C2619 vdd.n524 gnd 0.01022f
C2620 vdd.n525 gnd 0.01022f
C2621 vdd.n526 gnd 0.008226f
C2622 vdd.n527 gnd 0.008226f
C2623 vdd.n528 gnd 0.01022f
C2624 vdd.n529 gnd 0.01022f
C2625 vdd.n530 gnd 0.008226f
C2626 vdd.n531 gnd 0.01022f
C2627 vdd.n532 gnd 0.01022f
C2628 vdd.n533 gnd 0.01022f
C2629 vdd.n534 gnd 0.01022f
C2630 vdd.n535 gnd 0.01022f
C2631 vdd.n536 gnd 0.008226f
C2632 vdd.n537 gnd 0.008226f
C2633 vdd.n538 gnd 0.01022f
C2634 vdd.n539 gnd 0.01022f
C2635 vdd.n540 gnd 0.008226f
C2636 vdd.n541 gnd 0.01022f
C2637 vdd.n542 gnd 0.01022f
C2638 vdd.n543 gnd 0.01022f
C2639 vdd.n544 gnd 0.01022f
C2640 vdd.n545 gnd 0.01022f
C2641 vdd.n546 gnd 0.005594f
C2642 vdd.n547 gnd 0.017604f
C2643 vdd.n548 gnd 0.01022f
C2644 vdd.n549 gnd 0.01022f
C2645 vdd.n550 gnd 0.008144f
C2646 vdd.n551 gnd 0.01022f
C2647 vdd.n552 gnd 0.01022f
C2648 vdd.n553 gnd 0.01022f
C2649 vdd.n554 gnd 0.01022f
C2650 vdd.n555 gnd 0.01022f
C2651 vdd.n556 gnd 0.008226f
C2652 vdd.n557 gnd 0.008226f
C2653 vdd.n558 gnd 0.01022f
C2654 vdd.n559 gnd 0.01022f
C2655 vdd.n560 gnd 0.008226f
C2656 vdd.n561 gnd 0.01022f
C2657 vdd.n562 gnd 0.01022f
C2658 vdd.n563 gnd 0.01022f
C2659 vdd.n564 gnd 0.01022f
C2660 vdd.n565 gnd 0.01022f
C2661 vdd.n566 gnd 0.008226f
C2662 vdd.n567 gnd 0.008226f
C2663 vdd.n568 gnd 0.01022f
C2664 vdd.n569 gnd 0.01022f
C2665 vdd.n570 gnd 0.008226f
C2666 vdd.n571 gnd 0.01022f
C2667 vdd.n572 gnd 0.01022f
C2668 vdd.n573 gnd 0.01022f
C2669 vdd.n574 gnd 0.01022f
C2670 vdd.n575 gnd 0.01022f
C2671 vdd.n576 gnd 0.008226f
C2672 vdd.n577 gnd 0.008226f
C2673 vdd.n578 gnd 0.01022f
C2674 vdd.n579 gnd 0.01022f
C2675 vdd.n580 gnd 0.008226f
C2676 vdd.n581 gnd 0.01022f
C2677 vdd.n582 gnd 0.01022f
C2678 vdd.n583 gnd 0.01022f
C2679 vdd.n584 gnd 0.01022f
C2680 vdd.n585 gnd 0.01022f
C2681 vdd.n586 gnd 0.008226f
C2682 vdd.n587 gnd 0.008226f
C2683 vdd.n588 gnd 0.01022f
C2684 vdd.n589 gnd 0.01022f
C2685 vdd.n590 gnd 0.008226f
C2686 vdd.n591 gnd 0.01022f
C2687 vdd.n592 gnd 0.01022f
C2688 vdd.n593 gnd 0.01022f
C2689 vdd.n594 gnd 0.01022f
C2690 vdd.n595 gnd 0.01022f
C2691 vdd.n596 gnd 0.008226f
C2692 vdd.n597 gnd 0.01022f
C2693 vdd.n598 gnd 0.008226f
C2694 vdd.n599 gnd 0.004319f
C2695 vdd.n600 gnd 0.01022f
C2696 vdd.n601 gnd 0.01022f
C2697 vdd.n602 gnd 0.008226f
C2698 vdd.n603 gnd 0.01022f
C2699 vdd.n604 gnd 0.008226f
C2700 vdd.n605 gnd 0.01022f
C2701 vdd.n606 gnd 0.008226f
C2702 vdd.n607 gnd 0.01022f
C2703 vdd.n608 gnd 0.008226f
C2704 vdd.n609 gnd 0.01022f
C2705 vdd.n610 gnd 0.008226f
C2706 vdd.n611 gnd 0.01022f
C2707 vdd.n612 gnd 0.01022f
C2708 vdd.n613 gnd 0.569244f
C2709 vdd.t96 gnd 0.522243f
C2710 vdd.n614 gnd 0.01022f
C2711 vdd.n615 gnd 0.008226f
C2712 vdd.n616 gnd 0.01022f
C2713 vdd.n617 gnd 0.008226f
C2714 vdd.n618 gnd 0.01022f
C2715 vdd.t93 gnd 0.522243f
C2716 vdd.n619 gnd 0.01022f
C2717 vdd.n620 gnd 0.008226f
C2718 vdd.n621 gnd 0.01022f
C2719 vdd.n622 gnd 0.008226f
C2720 vdd.n623 gnd 0.01022f
C2721 vdd.t100 gnd 0.522243f
C2722 vdd.n624 gnd 0.652803f
C2723 vdd.n625 gnd 0.01022f
C2724 vdd.n626 gnd 0.008226f
C2725 vdd.n627 gnd 0.01022f
C2726 vdd.n628 gnd 0.008226f
C2727 vdd.n629 gnd 0.01022f
C2728 vdd.t102 gnd 0.522243f
C2729 vdd.n630 gnd 0.01022f
C2730 vdd.n631 gnd 0.008226f
C2731 vdd.n632 gnd 0.01022f
C2732 vdd.n633 gnd 0.008226f
C2733 vdd.n634 gnd 0.01022f
C2734 vdd.n635 gnd 0.725917f
C2735 vdd.n636 gnd 0.866923f
C2736 vdd.t136 gnd 0.522243f
C2737 vdd.n637 gnd 0.01022f
C2738 vdd.n638 gnd 0.008226f
C2739 vdd.n639 gnd 0.01022f
C2740 vdd.n640 gnd 0.008226f
C2741 vdd.n641 gnd 0.01022f
C2742 vdd.n642 gnd 0.548355f
C2743 vdd.n643 gnd 0.01022f
C2744 vdd.n644 gnd 0.008226f
C2745 vdd.n645 gnd 0.01022f
C2746 vdd.n646 gnd 0.008226f
C2747 vdd.n647 gnd 0.01022f
C2748 vdd.n648 gnd 1.04449f
C2749 vdd.t161 gnd 0.522243f
C2750 vdd.n649 gnd 0.01022f
C2751 vdd.n650 gnd 0.008226f
C2752 vdd.n651 gnd 0.01022f
C2753 vdd.n652 gnd 0.008226f
C2754 vdd.n653 gnd 0.01022f
C2755 vdd.t26 gnd 0.522243f
C2756 vdd.n654 gnd 0.01022f
C2757 vdd.n655 gnd 0.008226f
C2758 vdd.n656 gnd 0.023433f
C2759 vdd.n657 gnd 0.023433f
C2760 vdd.n658 gnd 9.118349f
C2761 vdd.n659 gnd 0.579689f
C2762 vdd.n660 gnd 0.023433f
C2763 vdd.n661 gnd 0.00879f
C2764 vdd.n662 gnd 0.008226f
C2765 vdd.n667 gnd 0.006541f
C2766 vdd.n668 gnd 0.008226f
C2767 vdd.n669 gnd 0.01022f
C2768 vdd.n670 gnd 0.01022f
C2769 vdd.n671 gnd 0.01022f
C2770 vdd.n672 gnd 0.01022f
C2771 vdd.n673 gnd 0.01022f
C2772 vdd.n674 gnd 0.008226f
C2773 vdd.n675 gnd 0.01022f
C2774 vdd.n676 gnd 0.01022f
C2775 vdd.n677 gnd 0.01022f
C2776 vdd.n678 gnd 0.01022f
C2777 vdd.n679 gnd 0.01022f
C2778 vdd.n680 gnd 0.008226f
C2779 vdd.n681 gnd 0.01022f
C2780 vdd.n682 gnd 0.01022f
C2781 vdd.n683 gnd 0.01022f
C2782 vdd.n684 gnd 0.01022f
C2783 vdd.n685 gnd 0.01022f
C2784 vdd.t44 gnd 0.125739f
C2785 vdd.t45 gnd 0.13438f
C2786 vdd.t43 gnd 0.164213f
C2787 vdd.n686 gnd 0.210498f
C2788 vdd.n687 gnd 0.176857f
C2789 vdd.n688 gnd 0.016782f
C2790 vdd.n689 gnd 0.01022f
C2791 vdd.n690 gnd 0.01022f
C2792 vdd.n691 gnd 0.01022f
C2793 vdd.n692 gnd 0.01022f
C2794 vdd.n693 gnd 0.01022f
C2795 vdd.n694 gnd 0.008226f
C2796 vdd.n695 gnd 0.01022f
C2797 vdd.n696 gnd 0.01022f
C2798 vdd.n697 gnd 0.01022f
C2799 vdd.n698 gnd 0.01022f
C2800 vdd.n699 gnd 0.01022f
C2801 vdd.n700 gnd 0.008226f
C2802 vdd.n701 gnd 0.01022f
C2803 vdd.n702 gnd 0.01022f
C2804 vdd.n703 gnd 0.01022f
C2805 vdd.n704 gnd 0.01022f
C2806 vdd.n705 gnd 0.01022f
C2807 vdd.n706 gnd 0.008226f
C2808 vdd.n707 gnd 0.01022f
C2809 vdd.n708 gnd 0.01022f
C2810 vdd.n709 gnd 0.01022f
C2811 vdd.n710 gnd 0.01022f
C2812 vdd.n711 gnd 0.01022f
C2813 vdd.n712 gnd 0.008226f
C2814 vdd.n713 gnd 0.01022f
C2815 vdd.n714 gnd 0.01022f
C2816 vdd.n715 gnd 0.01022f
C2817 vdd.n716 gnd 0.01022f
C2818 vdd.n717 gnd 0.01022f
C2819 vdd.n718 gnd 0.008226f
C2820 vdd.n719 gnd 0.01022f
C2821 vdd.n720 gnd 0.01022f
C2822 vdd.n721 gnd 0.01022f
C2823 vdd.n722 gnd 0.008144f
C2824 vdd.t34 gnd 0.125739f
C2825 vdd.t35 gnd 0.13438f
C2826 vdd.t33 gnd 0.164213f
C2827 vdd.n723 gnd 0.210498f
C2828 vdd.n724 gnd 0.176857f
C2829 vdd.n725 gnd 0.01022f
C2830 vdd.n726 gnd 0.008226f
C2831 vdd.n728 gnd 0.01022f
C2832 vdd.n730 gnd 0.01022f
C2833 vdd.n731 gnd 0.01022f
C2834 vdd.n732 gnd 0.008226f
C2835 vdd.n733 gnd 0.01022f
C2836 vdd.n734 gnd 0.01022f
C2837 vdd.n735 gnd 0.01022f
C2838 vdd.n736 gnd 0.01022f
C2839 vdd.n737 gnd 0.01022f
C2840 vdd.n738 gnd 0.008226f
C2841 vdd.n739 gnd 0.01022f
C2842 vdd.n740 gnd 0.01022f
C2843 vdd.n741 gnd 0.01022f
C2844 vdd.n742 gnd 0.01022f
C2845 vdd.n743 gnd 0.01022f
C2846 vdd.n744 gnd 0.008226f
C2847 vdd.n745 gnd 0.01022f
C2848 vdd.n746 gnd 0.01022f
C2849 vdd.n747 gnd 0.01022f
C2850 vdd.n748 gnd 0.006541f
C2851 vdd.n753 gnd 0.00695f
C2852 vdd.n754 gnd 0.00695f
C2853 vdd.n755 gnd 0.00695f
C2854 vdd.n756 gnd 8.90946f
C2855 vdd.n757 gnd 0.00695f
C2856 vdd.n758 gnd 0.00695f
C2857 vdd.n759 gnd 0.00695f
C2858 vdd.n761 gnd 0.00695f
C2859 vdd.n762 gnd 0.00695f
C2860 vdd.n764 gnd 0.00695f
C2861 vdd.n765 gnd 0.005059f
C2862 vdd.n767 gnd 0.00695f
C2863 vdd.t20 gnd 0.280846f
C2864 vdd.t19 gnd 0.28748f
C2865 vdd.t17 gnd 0.183347f
C2866 vdd.n768 gnd 0.099089f
C2867 vdd.n769 gnd 0.056206f
C2868 vdd.n770 gnd 0.009933f
C2869 vdd.n771 gnd 0.016087f
C2870 vdd.n773 gnd 0.00695f
C2871 vdd.n774 gnd 0.71025f
C2872 vdd.n775 gnd 0.015224f
C2873 vdd.n776 gnd 0.015224f
C2874 vdd.n777 gnd 0.00695f
C2875 vdd.n778 gnd 0.016255f
C2876 vdd.n779 gnd 0.00695f
C2877 vdd.n780 gnd 0.00695f
C2878 vdd.n781 gnd 0.00695f
C2879 vdd.n782 gnd 0.00695f
C2880 vdd.n783 gnd 0.00695f
C2881 vdd.n785 gnd 0.00695f
C2882 vdd.n786 gnd 0.00695f
C2883 vdd.n788 gnd 0.00695f
C2884 vdd.n789 gnd 0.00695f
C2885 vdd.n791 gnd 0.00695f
C2886 vdd.n792 gnd 0.00695f
C2887 vdd.n794 gnd 0.00695f
C2888 vdd.n795 gnd 0.00695f
C2889 vdd.n797 gnd 0.00695f
C2890 vdd.n798 gnd 0.00695f
C2891 vdd.n800 gnd 0.00695f
C2892 vdd.n801 gnd 0.005059f
C2893 vdd.n803 gnd 0.00695f
C2894 vdd.t89 gnd 0.280846f
C2895 vdd.t88 gnd 0.28748f
C2896 vdd.t87 gnd 0.183347f
C2897 vdd.n804 gnd 0.099089f
C2898 vdd.n805 gnd 0.056206f
C2899 vdd.n806 gnd 0.009933f
C2900 vdd.n807 gnd 0.00695f
C2901 vdd.n808 gnd 0.00695f
C2902 vdd.t18 gnd 0.355125f
C2903 vdd.n809 gnd 0.00695f
C2904 vdd.n810 gnd 0.00695f
C2905 vdd.n811 gnd 0.00695f
C2906 vdd.n812 gnd 0.00695f
C2907 vdd.n813 gnd 0.00695f
C2908 vdd.n814 gnd 0.71025f
C2909 vdd.n815 gnd 0.00695f
C2910 vdd.n816 gnd 0.00695f
C2911 vdd.n817 gnd 0.600579f
C2912 vdd.n818 gnd 0.00695f
C2913 vdd.n819 gnd 0.00695f
C2914 vdd.n820 gnd 0.00695f
C2915 vdd.n821 gnd 0.00695f
C2916 vdd.n822 gnd 0.694583f
C2917 vdd.n823 gnd 0.00695f
C2918 vdd.n824 gnd 0.00695f
C2919 vdd.n825 gnd 0.00695f
C2920 vdd.n826 gnd 0.00695f
C2921 vdd.n827 gnd 0.00695f
C2922 vdd.n828 gnd 0.71025f
C2923 vdd.n829 gnd 0.00695f
C2924 vdd.n830 gnd 0.00695f
C2925 vdd.t226 gnd 0.355125f
C2926 vdd.n831 gnd 0.00695f
C2927 vdd.n832 gnd 0.00695f
C2928 vdd.n833 gnd 0.00695f
C2929 vdd.t199 gnd 0.355125f
C2930 vdd.n834 gnd 0.00695f
C2931 vdd.n835 gnd 0.00695f
C2932 vdd.n836 gnd 0.00695f
C2933 vdd.n837 gnd 0.00695f
C2934 vdd.n838 gnd 0.00695f
C2935 vdd.t40 gnd 0.297678f
C2936 vdd.n839 gnd 0.00695f
C2937 vdd.n840 gnd 0.00695f
C2938 vdd.n841 gnd 0.569244f
C2939 vdd.n842 gnd 0.00695f
C2940 vdd.t41 gnd 0.28748f
C2941 vdd.t39 gnd 0.183347f
C2942 vdd.t42 gnd 0.28748f
C2943 vdd.n843 gnd 0.161576f
C2944 vdd.n844 gnd 0.00695f
C2945 vdd.n845 gnd 0.00695f
C2946 vdd.n846 gnd 0.454351f
C2947 vdd.n847 gnd 0.00695f
C2948 vdd.n848 gnd 0.00695f
C2949 vdd.t201 gnd 0.104449f
C2950 vdd.n849 gnd 0.412572f
C2951 vdd.n850 gnd 0.00695f
C2952 vdd.n851 gnd 0.00695f
C2953 vdd.n852 gnd 0.00695f
C2954 vdd.n853 gnd 0.611024f
C2955 vdd.n854 gnd 0.00695f
C2956 vdd.n855 gnd 0.00695f
C2957 vdd.t211 gnd 0.355125f
C2958 vdd.n856 gnd 0.00695f
C2959 vdd.n857 gnd 0.00695f
C2960 vdd.n858 gnd 0.00695f
C2961 vdd.t207 gnd 0.355125f
C2962 vdd.n859 gnd 0.00695f
C2963 vdd.n860 gnd 0.00695f
C2964 vdd.t227 gnd 0.355125f
C2965 vdd.n861 gnd 0.00695f
C2966 vdd.n862 gnd 0.00695f
C2967 vdd.n863 gnd 0.00695f
C2968 vdd.t192 gnd 0.282011f
C2969 vdd.n864 gnd 0.00695f
C2970 vdd.n865 gnd 0.00695f
C2971 vdd.n866 gnd 0.584912f
C2972 vdd.n867 gnd 0.00695f
C2973 vdd.n868 gnd 0.00695f
C2974 vdd.n869 gnd 0.00695f
C2975 vdd.t228 gnd 0.355125f
C2976 vdd.n870 gnd 0.00695f
C2977 vdd.n871 gnd 0.00695f
C2978 vdd.t238 gnd 0.297678f
C2979 vdd.n872 gnd 0.428239f
C2980 vdd.n873 gnd 0.00695f
C2981 vdd.n874 gnd 0.00695f
C2982 vdd.n875 gnd 0.00695f
C2983 vdd.n876 gnd 0.370792f
C2984 vdd.n877 gnd 0.00695f
C2985 vdd.n878 gnd 0.00695f
C2986 vdd.t231 gnd 0.355125f
C2987 vdd.n879 gnd 0.00695f
C2988 vdd.n880 gnd 0.00695f
C2989 vdd.n881 gnd 0.00695f
C2990 vdd.n882 gnd 0.71025f
C2991 vdd.n883 gnd 0.00695f
C2992 vdd.n884 gnd 0.00695f
C2993 vdd.t196 gnd 0.240232f
C2994 vdd.t215 gnd 0.339458f
C2995 vdd.n885 gnd 0.00695f
C2996 vdd.n886 gnd 0.00695f
C2997 vdd.n887 gnd 0.00695f
C2998 vdd.n888 gnd 0.532687f
C2999 vdd.n889 gnd 0.00695f
C3000 vdd.n890 gnd 0.00695f
C3001 vdd.n891 gnd 0.00695f
C3002 vdd.n892 gnd 0.00695f
C3003 vdd.n893 gnd 0.00695f
C3004 vdd.t68 gnd 0.355125f
C3005 vdd.n894 gnd 0.00695f
C3006 vdd.n895 gnd 0.00695f
C3007 vdd.t197 gnd 0.355125f
C3008 vdd.n896 gnd 0.00695f
C3009 vdd.n897 gnd 0.015224f
C3010 vdd.n898 gnd 0.015224f
C3011 vdd.n899 gnd 0.846033f
C3012 vdd.n900 gnd 0.00695f
C3013 vdd.n901 gnd 0.00695f
C3014 vdd.t222 gnd 0.355125f
C3015 vdd.n902 gnd 0.015224f
C3016 vdd.n903 gnd 0.00695f
C3017 vdd.n904 gnd 0.00695f
C3018 vdd.t235 gnd 0.647581f
C3019 vdd.n922 gnd 0.016255f
C3020 vdd.n940 gnd 0.015224f
C3021 vdd.n941 gnd 0.00695f
C3022 vdd.n942 gnd 0.015224f
C3023 vdd.t83 gnd 0.280846f
C3024 vdd.t82 gnd 0.28748f
C3025 vdd.t81 gnd 0.183347f
C3026 vdd.n943 gnd 0.099089f
C3027 vdd.n944 gnd 0.056206f
C3028 vdd.n945 gnd 0.016087f
C3029 vdd.n946 gnd 0.00695f
C3030 vdd.n947 gnd 0.376015f
C3031 vdd.n948 gnd 0.015224f
C3032 vdd.n949 gnd 0.00695f
C3033 vdd.n950 gnd 0.016255f
C3034 vdd.n951 gnd 0.00695f
C3035 vdd.t66 gnd 0.280846f
C3036 vdd.t65 gnd 0.28748f
C3037 vdd.t63 gnd 0.183347f
C3038 vdd.n952 gnd 0.099089f
C3039 vdd.n953 gnd 0.056206f
C3040 vdd.n954 gnd 0.009933f
C3041 vdd.n955 gnd 0.00695f
C3042 vdd.n956 gnd 0.00695f
C3043 vdd.t64 gnd 0.355125f
C3044 vdd.n957 gnd 0.00695f
C3045 vdd.t233 gnd 0.355125f
C3046 vdd.n958 gnd 0.00695f
C3047 vdd.n959 gnd 0.00695f
C3048 vdd.n960 gnd 0.00695f
C3049 vdd.n961 gnd 0.00695f
C3050 vdd.n962 gnd 0.00695f
C3051 vdd.n963 gnd 0.71025f
C3052 vdd.n964 gnd 0.00695f
C3053 vdd.n965 gnd 0.00695f
C3054 vdd.t209 gnd 0.355125f
C3055 vdd.n966 gnd 0.00695f
C3056 vdd.n967 gnd 0.00695f
C3057 vdd.n968 gnd 0.00695f
C3058 vdd.n969 gnd 0.00695f
C3059 vdd.n970 gnd 0.470018f
C3060 vdd.n971 gnd 0.00695f
C3061 vdd.n972 gnd 0.00695f
C3062 vdd.n973 gnd 0.00695f
C3063 vdd.n974 gnd 0.00695f
C3064 vdd.n975 gnd 0.00695f
C3065 vdd.n976 gnd 0.626691f
C3066 vdd.n977 gnd 0.00695f
C3067 vdd.n978 gnd 0.00695f
C3068 vdd.t224 gnd 0.339458f
C3069 vdd.t193 gnd 0.240232f
C3070 vdd.n979 gnd 0.00695f
C3071 vdd.n980 gnd 0.00695f
C3072 vdd.n981 gnd 0.00695f
C3073 vdd.t214 gnd 0.355125f
C3074 vdd.n982 gnd 0.00695f
C3075 vdd.n983 gnd 0.00695f
C3076 vdd.t194 gnd 0.355125f
C3077 vdd.n984 gnd 0.00695f
C3078 vdd.n985 gnd 0.00695f
C3079 vdd.n986 gnd 0.00695f
C3080 vdd.t212 gnd 0.297678f
C3081 vdd.n987 gnd 0.00695f
C3082 vdd.n988 gnd 0.00695f
C3083 vdd.n989 gnd 0.569244f
C3084 vdd.n990 gnd 0.00695f
C3085 vdd.n991 gnd 0.00695f
C3086 vdd.n992 gnd 0.00695f
C3087 vdd.t229 gnd 0.355125f
C3088 vdd.n993 gnd 0.00695f
C3089 vdd.n994 gnd 0.00695f
C3090 vdd.t202 gnd 0.282011f
C3091 vdd.n995 gnd 0.412572f
C3092 vdd.n996 gnd 0.00695f
C3093 vdd.n997 gnd 0.00695f
C3094 vdd.n998 gnd 0.00695f
C3095 vdd.n999 gnd 0.611024f
C3096 vdd.n1000 gnd 0.00695f
C3097 vdd.n1001 gnd 0.00695f
C3098 vdd.t237 gnd 0.355125f
C3099 vdd.n1002 gnd 0.00695f
C3100 vdd.n1003 gnd 0.00695f
C3101 vdd.n1004 gnd 0.00695f
C3102 vdd.n1005 gnd 0.71025f
C3103 vdd.n1006 gnd 0.00695f
C3104 vdd.n1007 gnd 0.00695f
C3105 vdd.t206 gnd 0.355125f
C3106 vdd.n1008 gnd 0.00695f
C3107 vdd.n1009 gnd 0.00695f
C3108 vdd.n1010 gnd 0.00695f
C3109 vdd.t200 gnd 0.104449f
C3110 vdd.n1011 gnd 0.00695f
C3111 vdd.n1012 gnd 0.00695f
C3112 vdd.n1013 gnd 0.00695f
C3113 vdd.t73 gnd 0.28748f
C3114 vdd.t71 gnd 0.183347f
C3115 vdd.t74 gnd 0.28748f
C3116 vdd.n1014 gnd 0.161576f
C3117 vdd.n1015 gnd 0.00695f
C3118 vdd.n1016 gnd 0.00695f
C3119 vdd.t219 gnd 0.355125f
C3120 vdd.n1017 gnd 0.00695f
C3121 vdd.n1018 gnd 0.00695f
C3122 vdd.t72 gnd 0.297678f
C3123 vdd.n1019 gnd 0.605801f
C3124 vdd.n1020 gnd 0.00695f
C3125 vdd.n1021 gnd 0.00695f
C3126 vdd.n1022 gnd 0.00695f
C3127 vdd.n1023 gnd 0.370792f
C3128 vdd.n1024 gnd 0.00695f
C3129 vdd.n1025 gnd 0.00695f
C3130 vdd.n1026 gnd 0.49613f
C3131 vdd.n1027 gnd 0.00695f
C3132 vdd.n1028 gnd 0.00695f
C3133 vdd.n1029 gnd 0.00695f
C3134 vdd.n1030 gnd 0.71025f
C3135 vdd.n1031 gnd 0.00695f
C3136 vdd.n1032 gnd 0.00695f
C3137 vdd.t203 gnd 0.355125f
C3138 vdd.n1033 gnd 0.00695f
C3139 vdd.n1034 gnd 0.00695f
C3140 vdd.n1035 gnd 0.00695f
C3141 vdd.n1036 gnd 0.71025f
C3142 vdd.n1037 gnd 0.00695f
C3143 vdd.n1038 gnd 0.00695f
C3144 vdd.n1039 gnd 0.00695f
C3145 vdd.n1040 gnd 0.00695f
C3146 vdd.n1041 gnd 0.00695f
C3147 vdd.t22 gnd 0.355125f
C3148 vdd.n1042 gnd 0.00695f
C3149 vdd.n1043 gnd 0.00695f
C3150 vdd.n1044 gnd 0.00695f
C3151 vdd.n1045 gnd 0.015224f
C3152 vdd.n1046 gnd 0.015224f
C3153 vdd.n1047 gnd 1.00271f
C3154 vdd.n1048 gnd 0.00695f
C3155 vdd.n1049 gnd 0.00695f
C3156 vdd.n1050 gnd 0.464796f
C3157 vdd.n1051 gnd 0.015224f
C3158 vdd.n1052 gnd 0.00695f
C3159 vdd.n1053 gnd 0.00695f
C3160 vdd.n1054 gnd 9.118349f
C3161 vdd.n1087 gnd 0.016255f
C3162 vdd.n1088 gnd 0.00695f
C3163 vdd.n1089 gnd 0.00695f
C3164 vdd.n1090 gnd 0.00695f
C3165 vdd.n1091 gnd 0.006541f
C3166 vdd.n1094 gnd 0.023433f
C3167 vdd.n1095 gnd 0.006828f
C3168 vdd.n1096 gnd 0.008226f
C3169 vdd.n1098 gnd 0.01022f
C3170 vdd.n1099 gnd 0.01022f
C3171 vdd.n1100 gnd 0.008226f
C3172 vdd.n1102 gnd 0.01022f
C3173 vdd.n1103 gnd 0.01022f
C3174 vdd.n1104 gnd 0.01022f
C3175 vdd.n1105 gnd 0.01022f
C3176 vdd.n1106 gnd 0.01022f
C3177 vdd.n1107 gnd 0.008226f
C3178 vdd.n1109 gnd 0.01022f
C3179 vdd.n1110 gnd 0.01022f
C3180 vdd.n1111 gnd 0.01022f
C3181 vdd.n1112 gnd 0.01022f
C3182 vdd.n1113 gnd 0.01022f
C3183 vdd.n1114 gnd 0.008226f
C3184 vdd.n1116 gnd 0.01022f
C3185 vdd.n1117 gnd 0.01022f
C3186 vdd.n1118 gnd 0.01022f
C3187 vdd.n1119 gnd 0.01022f
C3188 vdd.n1120 gnd 0.006869f
C3189 vdd.t80 gnd 0.125739f
C3190 vdd.t79 gnd 0.13438f
C3191 vdd.t78 gnd 0.164213f
C3192 vdd.n1121 gnd 0.210498f
C3193 vdd.n1122 gnd 0.176857f
C3194 vdd.n1124 gnd 0.01022f
C3195 vdd.n1125 gnd 0.01022f
C3196 vdd.n1126 gnd 0.008226f
C3197 vdd.n1127 gnd 0.01022f
C3198 vdd.n1129 gnd 0.01022f
C3199 vdd.n1130 gnd 0.01022f
C3200 vdd.n1131 gnd 0.01022f
C3201 vdd.n1132 gnd 0.01022f
C3202 vdd.n1133 gnd 0.008226f
C3203 vdd.n1135 gnd 0.01022f
C3204 vdd.n1136 gnd 0.01022f
C3205 vdd.n1137 gnd 0.01022f
C3206 vdd.n1138 gnd 0.01022f
C3207 vdd.n1139 gnd 0.01022f
C3208 vdd.n1140 gnd 0.008226f
C3209 vdd.n1142 gnd 0.01022f
C3210 vdd.n1143 gnd 0.01022f
C3211 vdd.n1144 gnd 0.01022f
C3212 vdd.n1145 gnd 0.01022f
C3213 vdd.n1146 gnd 0.01022f
C3214 vdd.n1147 gnd 0.008226f
C3215 vdd.n1149 gnd 0.01022f
C3216 vdd.n1150 gnd 0.01022f
C3217 vdd.n1151 gnd 0.01022f
C3218 vdd.n1152 gnd 0.01022f
C3219 vdd.n1153 gnd 0.01022f
C3220 vdd.n1154 gnd 0.008226f
C3221 vdd.n1156 gnd 0.01022f
C3222 vdd.n1157 gnd 0.01022f
C3223 vdd.n1158 gnd 0.01022f
C3224 vdd.n1159 gnd 0.01022f
C3225 vdd.n1160 gnd 0.008144f
C3226 vdd.t62 gnd 0.125739f
C3227 vdd.t61 gnd 0.13438f
C3228 vdd.t60 gnd 0.164213f
C3229 vdd.n1161 gnd 0.210498f
C3230 vdd.n1162 gnd 0.176857f
C3231 vdd.n1164 gnd 0.01022f
C3232 vdd.n1165 gnd 0.01022f
C3233 vdd.n1166 gnd 0.008226f
C3234 vdd.n1167 gnd 0.01022f
C3235 vdd.n1169 gnd 0.01022f
C3236 vdd.n1170 gnd 0.01022f
C3237 vdd.n1171 gnd 0.01022f
C3238 vdd.n1172 gnd 0.01022f
C3239 vdd.n1173 gnd 0.008226f
C3240 vdd.n1175 gnd 0.01022f
C3241 vdd.n1176 gnd 0.01022f
C3242 vdd.n1177 gnd 0.01022f
C3243 vdd.n1178 gnd 0.01022f
C3244 vdd.n1179 gnd 0.01022f
C3245 vdd.n1180 gnd 0.008226f
C3246 vdd.n1182 gnd 0.01022f
C3247 vdd.n1183 gnd 0.01022f
C3248 vdd.n1184 gnd 0.01022f
C3249 vdd.n1185 gnd 0.01022f
C3250 vdd.n1186 gnd 0.01022f
C3251 vdd.n1187 gnd 0.008226f
C3252 vdd.n1189 gnd 0.01022f
C3253 vdd.n1190 gnd 0.01022f
C3254 vdd.n1191 gnd 0.006541f
C3255 vdd.n1192 gnd 0.008226f
C3256 vdd.n1193 gnd 0.00695f
C3257 vdd.n1194 gnd 0.00695f
C3258 vdd.n1195 gnd 0.00695f
C3259 vdd.n1196 gnd 0.00695f
C3260 vdd.n1197 gnd 0.00695f
C3261 vdd.n1198 gnd 0.00695f
C3262 vdd.n1199 gnd 0.00695f
C3263 vdd.n1200 gnd 0.00695f
C3264 vdd.n1201 gnd 0.00695f
C3265 vdd.n1202 gnd 0.00695f
C3266 vdd.n1203 gnd 0.00695f
C3267 vdd.n1204 gnd 0.00695f
C3268 vdd.n1205 gnd 0.00695f
C3269 vdd.n1206 gnd 0.00695f
C3270 vdd.n1207 gnd 0.00695f
C3271 vdd.n1208 gnd 0.00695f
C3272 vdd.n1209 gnd 0.00695f
C3273 vdd.n1210 gnd 0.00695f
C3274 vdd.n1211 gnd 0.00695f
C3275 vdd.n1212 gnd 0.00695f
C3276 vdd.n1213 gnd 0.00695f
C3277 vdd.n1214 gnd 0.00695f
C3278 vdd.n1215 gnd 0.00695f
C3279 vdd.n1216 gnd 0.00695f
C3280 vdd.n1217 gnd 0.00695f
C3281 vdd.n1218 gnd 0.00695f
C3282 vdd.n1219 gnd 0.00695f
C3283 vdd.n1220 gnd 0.00695f
C3284 vdd.n1221 gnd 0.00695f
C3285 vdd.n1222 gnd 0.00695f
C3286 vdd.n1223 gnd 0.00695f
C3287 vdd.t23 gnd 0.280846f
C3288 vdd.t24 gnd 0.28748f
C3289 vdd.t21 gnd 0.183347f
C3290 vdd.n1224 gnd 0.099089f
C3291 vdd.n1225 gnd 0.056206f
C3292 vdd.n1226 gnd 0.009933f
C3293 vdd.n1227 gnd 0.00695f
C3294 vdd.n1228 gnd 0.00695f
C3295 vdd.n1229 gnd 0.00695f
C3296 vdd.n1230 gnd 0.00695f
C3297 vdd.n1231 gnd 0.00695f
C3298 vdd.n1232 gnd 0.00695f
C3299 vdd.n1233 gnd 0.00695f
C3300 vdd.n1234 gnd 0.00695f
C3301 vdd.n1235 gnd 0.00695f
C3302 vdd.n1236 gnd 0.00695f
C3303 vdd.n1237 gnd 0.00695f
C3304 vdd.n1238 gnd 0.00695f
C3305 vdd.n1239 gnd 0.00695f
C3306 vdd.n1240 gnd 0.00695f
C3307 vdd.n1241 gnd 0.00695f
C3308 vdd.n1242 gnd 0.00695f
C3309 vdd.n1243 gnd 0.00695f
C3310 vdd.t37 gnd 0.280846f
C3311 vdd.t38 gnd 0.28748f
C3312 vdd.t36 gnd 0.183347f
C3313 vdd.n1244 gnd 0.099089f
C3314 vdd.n1245 gnd 0.056206f
C3315 vdd.n1246 gnd 0.00695f
C3316 vdd.n1247 gnd 0.00695f
C3317 vdd.n1248 gnd 0.00695f
C3318 vdd.n1249 gnd 0.00695f
C3319 vdd.n1250 gnd 0.00695f
C3320 vdd.n1251 gnd 0.00695f
C3321 vdd.n1252 gnd 0.00695f
C3322 vdd.n1253 gnd 0.00695f
C3323 vdd.n1254 gnd 0.00695f
C3324 vdd.n1255 gnd 0.00695f
C3325 vdd.n1256 gnd 0.00695f
C3326 vdd.n1257 gnd 0.00695f
C3327 vdd.n1258 gnd 0.00695f
C3328 vdd.n1259 gnd 0.00695f
C3329 vdd.n1260 gnd 0.00695f
C3330 vdd.n1261 gnd 0.00695f
C3331 vdd.n1262 gnd 0.00695f
C3332 vdd.n1263 gnd 0.00695f
C3333 vdd.n1264 gnd 0.00695f
C3334 vdd.n1265 gnd 0.00695f
C3335 vdd.n1266 gnd 0.00695f
C3336 vdd.n1267 gnd 0.00695f
C3337 vdd.n1268 gnd 0.00695f
C3338 vdd.n1269 gnd 0.00695f
C3339 vdd.n1270 gnd 0.00695f
C3340 vdd.n1271 gnd 0.00695f
C3341 vdd.n1272 gnd 0.005059f
C3342 vdd.n1273 gnd 0.009933f
C3343 vdd.n1274 gnd 0.005366f
C3344 vdd.n1275 gnd 0.00695f
C3345 vdd.n1276 gnd 0.00695f
C3346 vdd.n1277 gnd 0.00695f
C3347 vdd.n1278 gnd 0.016255f
C3348 vdd.n1279 gnd 0.016255f
C3349 vdd.n1280 gnd 0.015224f
C3350 vdd.n1281 gnd 0.015224f
C3351 vdd.n1282 gnd 0.00695f
C3352 vdd.n1283 gnd 0.00695f
C3353 vdd.n1284 gnd 0.00695f
C3354 vdd.n1285 gnd 0.00695f
C3355 vdd.n1286 gnd 0.00695f
C3356 vdd.n1287 gnd 0.00695f
C3357 vdd.n1288 gnd 0.00695f
C3358 vdd.n1289 gnd 0.00695f
C3359 vdd.n1290 gnd 0.00695f
C3360 vdd.n1291 gnd 0.00695f
C3361 vdd.n1292 gnd 0.00695f
C3362 vdd.n1293 gnd 0.00695f
C3363 vdd.n1294 gnd 0.00695f
C3364 vdd.n1295 gnd 0.00695f
C3365 vdd.n1296 gnd 0.00695f
C3366 vdd.n1297 gnd 0.00695f
C3367 vdd.n1298 gnd 0.00695f
C3368 vdd.n1299 gnd 0.00695f
C3369 vdd.n1300 gnd 0.00695f
C3370 vdd.n1301 gnd 0.00695f
C3371 vdd.n1302 gnd 0.00695f
C3372 vdd.n1303 gnd 0.00695f
C3373 vdd.n1304 gnd 0.00695f
C3374 vdd.n1305 gnd 0.00695f
C3375 vdd.n1306 gnd 0.00695f
C3376 vdd.n1307 gnd 0.00695f
C3377 vdd.n1308 gnd 0.00695f
C3378 vdd.n1309 gnd 0.423016f
C3379 vdd.n1310 gnd 0.00695f
C3380 vdd.n1311 gnd 0.00695f
C3381 vdd.n1312 gnd 0.00695f
C3382 vdd.n1313 gnd 0.00695f
C3383 vdd.n1314 gnd 0.00695f
C3384 vdd.n1315 gnd 0.00695f
C3385 vdd.n1316 gnd 0.00695f
C3386 vdd.n1317 gnd 0.00695f
C3387 vdd.n1318 gnd 0.00695f
C3388 vdd.n1319 gnd 0.00695f
C3389 vdd.n1320 gnd 0.00695f
C3390 vdd.n1321 gnd 0.00695f
C3391 vdd.n1322 gnd 0.00695f
C3392 vdd.n1323 gnd 0.00695f
C3393 vdd.n1324 gnd 0.00695f
C3394 vdd.n1325 gnd 0.00695f
C3395 vdd.n1326 gnd 0.00695f
C3396 vdd.n1327 gnd 0.00695f
C3397 vdd.n1328 gnd 0.00695f
C3398 vdd.n1329 gnd 0.00695f
C3399 vdd.n1330 gnd 0.224564f
C3400 vdd.n1331 gnd 0.00695f
C3401 vdd.n1332 gnd 0.00695f
C3402 vdd.n1333 gnd 0.00695f
C3403 vdd.n1334 gnd 0.00695f
C3404 vdd.n1335 gnd 0.00695f
C3405 vdd.n1336 gnd 0.00695f
C3406 vdd.n1337 gnd 0.00695f
C3407 vdd.n1338 gnd 0.00695f
C3408 vdd.n1339 gnd 0.00695f
C3409 vdd.n1340 gnd 0.00695f
C3410 vdd.n1341 gnd 0.00695f
C3411 vdd.n1342 gnd 0.00695f
C3412 vdd.n1343 gnd 0.00695f
C3413 vdd.n1344 gnd 0.00695f
C3414 vdd.n1345 gnd 0.00695f
C3415 vdd.n1346 gnd 0.00695f
C3416 vdd.n1347 gnd 0.00695f
C3417 vdd.n1348 gnd 0.00695f
C3418 vdd.n1349 gnd 0.00695f
C3419 vdd.n1350 gnd 0.00695f
C3420 vdd.n1351 gnd 0.00695f
C3421 vdd.n1352 gnd 0.00695f
C3422 vdd.n1353 gnd 0.00695f
C3423 vdd.n1354 gnd 0.00695f
C3424 vdd.n1355 gnd 0.00695f
C3425 vdd.n1356 gnd 0.00695f
C3426 vdd.n1357 gnd 0.00695f
C3427 vdd.n1358 gnd 0.015224f
C3428 vdd.n1359 gnd 0.015224f
C3429 vdd.n1360 gnd 0.016255f
C3430 vdd.n1361 gnd 0.00695f
C3431 vdd.n1362 gnd 0.00695f
C3432 vdd.n1363 gnd 0.005366f
C3433 vdd.n1364 gnd 0.00695f
C3434 vdd.n1365 gnd 0.00695f
C3435 vdd.n1366 gnd 0.005059f
C3436 vdd.n1367 gnd 0.00695f
C3437 vdd.n1368 gnd 0.00695f
C3438 vdd.n1369 gnd 0.00695f
C3439 vdd.n1370 gnd 0.00695f
C3440 vdd.n1371 gnd 0.00695f
C3441 vdd.n1372 gnd 0.00695f
C3442 vdd.n1373 gnd 0.00695f
C3443 vdd.n1374 gnd 0.00695f
C3444 vdd.n1375 gnd 0.00695f
C3445 vdd.n1376 gnd 0.00695f
C3446 vdd.n1377 gnd 0.00695f
C3447 vdd.n1378 gnd 0.00695f
C3448 vdd.n1379 gnd 0.00695f
C3449 vdd.n1380 gnd 0.00695f
C3450 vdd.n1381 gnd 0.00695f
C3451 vdd.n1382 gnd 0.00695f
C3452 vdd.n1383 gnd 0.00695f
C3453 vdd.n1384 gnd 0.00695f
C3454 vdd.n1385 gnd 0.00695f
C3455 vdd.n1386 gnd 0.00695f
C3456 vdd.n1387 gnd 0.00695f
C3457 vdd.n1388 gnd 0.00695f
C3458 vdd.n1389 gnd 0.00695f
C3459 vdd.n1390 gnd 0.00695f
C3460 vdd.n1391 gnd 0.00695f
C3461 vdd.n1392 gnd 0.00695f
C3462 vdd.n1393 gnd 0.027855f
C3463 vdd.n1395 gnd 0.023433f
C3464 vdd.n1396 gnd 0.008226f
C3465 vdd.n1398 gnd 0.01022f
C3466 vdd.n1399 gnd 0.008226f
C3467 vdd.n1400 gnd 0.01022f
C3468 vdd.n1402 gnd 0.01022f
C3469 vdd.n1403 gnd 0.01022f
C3470 vdd.n1405 gnd 0.01022f
C3471 vdd.n1406 gnd 0.006828f
C3472 vdd.n1407 gnd 0.579689f
C3473 vdd.n1408 gnd 0.01022f
C3474 vdd.n1409 gnd 0.023433f
C3475 vdd.n1410 gnd 0.008226f
C3476 vdd.n1411 gnd 0.01022f
C3477 vdd.n1412 gnd 0.008226f
C3478 vdd.n1413 gnd 0.01022f
C3479 vdd.n1414 gnd 1.04449f
C3480 vdd.n1415 gnd 0.01022f
C3481 vdd.n1416 gnd 0.008226f
C3482 vdd.n1417 gnd 0.008226f
C3483 vdd.n1418 gnd 0.01022f
C3484 vdd.n1419 gnd 0.008226f
C3485 vdd.n1420 gnd 0.01022f
C3486 vdd.t169 gnd 0.522243f
C3487 vdd.n1421 gnd 0.01022f
C3488 vdd.n1422 gnd 0.008226f
C3489 vdd.n1423 gnd 0.01022f
C3490 vdd.n1424 gnd 0.008226f
C3491 vdd.n1425 gnd 0.01022f
C3492 vdd.t188 gnd 0.522243f
C3493 vdd.n1426 gnd 0.01022f
C3494 vdd.n1427 gnd 0.008226f
C3495 vdd.n1428 gnd 0.01022f
C3496 vdd.n1429 gnd 0.008226f
C3497 vdd.n1430 gnd 0.01022f
C3498 vdd.t6 gnd 0.522243f
C3499 vdd.n1431 gnd 0.725917f
C3500 vdd.n1432 gnd 0.01022f
C3501 vdd.n1433 gnd 0.008226f
C3502 vdd.n1434 gnd 0.01022f
C3503 vdd.n1435 gnd 0.008226f
C3504 vdd.n1436 gnd 0.01022f
C3505 vdd.n1437 gnd 0.830366f
C3506 vdd.n1438 gnd 0.01022f
C3507 vdd.n1439 gnd 0.008226f
C3508 vdd.n1440 gnd 0.01022f
C3509 vdd.n1441 gnd 0.008226f
C3510 vdd.n1442 gnd 0.01022f
C3511 vdd.n1443 gnd 0.652803f
C3512 vdd.t146 gnd 0.522243f
C3513 vdd.n1444 gnd 0.01022f
C3514 vdd.n1445 gnd 0.008226f
C3515 vdd.n1446 gnd 0.01022f
C3516 vdd.n1447 gnd 0.008226f
C3517 vdd.n1448 gnd 0.01022f
C3518 vdd.t152 gnd 0.522243f
C3519 vdd.n1449 gnd 0.01022f
C3520 vdd.n1450 gnd 0.008226f
C3521 vdd.n1451 gnd 0.01022f
C3522 vdd.n1452 gnd 0.008226f
C3523 vdd.n1453 gnd 0.01022f
C3524 vdd.t172 gnd 0.522243f
C3525 vdd.n1454 gnd 0.569244f
C3526 vdd.n1455 gnd 0.01022f
C3527 vdd.n1456 gnd 0.008226f
C3528 vdd.n1457 gnd 0.01022f
C3529 vdd.n1458 gnd 0.008226f
C3530 vdd.n1459 gnd 0.01022f
C3531 vdd.t130 gnd 0.522243f
C3532 vdd.n1460 gnd 0.01022f
C3533 vdd.n1461 gnd 0.008226f
C3534 vdd.n1462 gnd 0.01022f
C3535 vdd.n1463 gnd 0.008226f
C3536 vdd.n1464 gnd 0.01022f
C3537 vdd.n1465 gnd 0.809476f
C3538 vdd.n1466 gnd 0.866923f
C3539 vdd.t148 gnd 0.522243f
C3540 vdd.n1467 gnd 0.01022f
C3541 vdd.n1468 gnd 0.008226f
C3542 vdd.n1469 gnd 0.01022f
C3543 vdd.n1470 gnd 0.008226f
C3544 vdd.n1471 gnd 0.01022f
C3545 vdd.n1472 gnd 0.631914f
C3546 vdd.n1473 gnd 0.01022f
C3547 vdd.n1474 gnd 0.008226f
C3548 vdd.n1475 gnd 0.01022f
C3549 vdd.n1476 gnd 0.008226f
C3550 vdd.n1477 gnd 0.01022f
C3551 vdd.t123 gnd 0.522243f
C3552 vdd.t138 gnd 0.522243f
C3553 vdd.n1478 gnd 0.01022f
C3554 vdd.n1479 gnd 0.008226f
C3555 vdd.n1480 gnd 0.01022f
C3556 vdd.n1481 gnd 0.008226f
C3557 vdd.n1482 gnd 0.01022f
C3558 vdd.t133 gnd 0.522243f
C3559 vdd.n1483 gnd 0.01022f
C3560 vdd.n1484 gnd 0.008226f
C3561 vdd.n1485 gnd 0.01022f
C3562 vdd.n1486 gnd 0.008226f
C3563 vdd.n1487 gnd 0.01022f
C3564 vdd.t110 gnd 0.522243f
C3565 vdd.n1488 gnd 0.767697f
C3566 vdd.n1489 gnd 0.01022f
C3567 vdd.n1490 gnd 0.008226f
C3568 vdd.n1491 gnd 0.01022f
C3569 vdd.n1492 gnd 0.008226f
C3570 vdd.n1493 gnd 0.01022f
C3571 vdd.n1494 gnd 1.04449f
C3572 vdd.n1495 gnd 0.01022f
C3573 vdd.n1496 gnd 0.008226f
C3574 vdd.n1497 gnd 0.01022f
C3575 vdd.n1498 gnd 0.008226f
C3576 vdd.n1499 gnd 0.01022f
C3577 vdd.n1500 gnd 0.88259f
C3578 vdd.n1501 gnd 0.01022f
C3579 vdd.n1502 gnd 0.008226f
C3580 vdd.n1503 gnd 0.023274f
C3581 vdd.n1504 gnd 0.006828f
C3582 vdd.n1505 gnd 0.023274f
C3583 vdd.n1506 gnd 1.37872f
C3584 vdd.n1507 gnd 0.023274f
C3585 vdd.n1508 gnd 0.006828f
C3586 vdd.n1509 gnd 0.01022f
C3587 vdd.t55 gnd 0.125739f
C3588 vdd.t56 gnd 0.13438f
C3589 vdd.t54 gnd 0.164213f
C3590 vdd.n1510 gnd 0.210498f
C3591 vdd.n1511 gnd 0.177679f
C3592 vdd.n1512 gnd 0.013491f
C3593 vdd.n1513 gnd 0.01022f
C3594 vdd.n1544 gnd 0.01022f
C3595 vdd.n1545 gnd 0.01022f
C3596 vdd.n1546 gnd 0.023433f
C3597 vdd.n1547 gnd 0.008226f
C3598 vdd.n1548 gnd 0.01022f
C3599 vdd.n1549 gnd 0.01022f
C3600 vdd.n1550 gnd 0.01022f
C3601 vdd.n1551 gnd 0.01022f
C3602 vdd.n1552 gnd 0.008226f
C3603 vdd.n1553 gnd 0.01022f
C3604 vdd.n1554 gnd 0.01022f
C3605 vdd.n1555 gnd 0.01022f
C3606 vdd.n1556 gnd 0.01022f
C3607 vdd.n1557 gnd 0.01022f
C3608 vdd.n1558 gnd 0.008226f
C3609 vdd.n1559 gnd 0.01022f
C3610 vdd.n1560 gnd 0.01022f
C3611 vdd.n1561 gnd 0.01022f
C3612 vdd.n1562 gnd 0.01022f
C3613 vdd.n1563 gnd 0.01022f
C3614 vdd.n1564 gnd 0.008226f
C3615 vdd.n1565 gnd 0.01022f
C3616 vdd.n1566 gnd 0.01022f
C3617 vdd.n1567 gnd 0.01022f
C3618 vdd.n1568 gnd 0.01022f
C3619 vdd.n1569 gnd 0.01022f
C3620 vdd.n1570 gnd 0.006869f
C3621 vdd.n1571 gnd 0.01022f
C3622 vdd.n1572 gnd 0.01022f
C3623 vdd.n1573 gnd 0.01022f
C3624 vdd.n1574 gnd 0.008226f
C3625 vdd.n1575 gnd 0.01022f
C3626 vdd.n1576 gnd 0.01022f
C3627 vdd.n1577 gnd 0.01022f
C3628 vdd.n1578 gnd 0.01022f
C3629 vdd.n1579 gnd 0.01022f
C3630 vdd.n1580 gnd 0.008226f
C3631 vdd.n1581 gnd 0.01022f
C3632 vdd.n1582 gnd 0.01022f
C3633 vdd.n1583 gnd 0.01022f
C3634 vdd.n1584 gnd 0.01022f
C3635 vdd.n1585 gnd 0.01022f
C3636 vdd.n1586 gnd 0.008226f
C3637 vdd.n1587 gnd 0.01022f
C3638 vdd.n1588 gnd 0.01022f
C3639 vdd.n1589 gnd 0.01022f
C3640 vdd.n1590 gnd 0.01022f
C3641 vdd.n1591 gnd 0.01022f
C3642 vdd.n1592 gnd 0.008226f
C3643 vdd.n1593 gnd 0.01022f
C3644 vdd.n1594 gnd 0.01022f
C3645 vdd.n1595 gnd 0.01022f
C3646 vdd.n1596 gnd 0.01022f
C3647 vdd.n1597 gnd 0.01022f
C3648 vdd.n1598 gnd 0.008226f
C3649 vdd.n1599 gnd 0.01022f
C3650 vdd.n1600 gnd 0.01022f
C3651 vdd.n1601 gnd 0.01022f
C3652 vdd.n1602 gnd 0.01022f
C3653 vdd.n1603 gnd 0.008144f
C3654 vdd.n1604 gnd 0.01022f
C3655 vdd.n1605 gnd 0.01022f
C3656 vdd.n1606 gnd 0.01022f
C3657 vdd.n1607 gnd 0.01022f
C3658 vdd.n1608 gnd 0.01022f
C3659 vdd.n1609 gnd 0.008226f
C3660 vdd.n1610 gnd 0.01022f
C3661 vdd.n1611 gnd 0.01022f
C3662 vdd.n1612 gnd 0.01022f
C3663 vdd.n1613 gnd 0.01022f
C3664 vdd.n1614 gnd 0.01022f
C3665 vdd.n1615 gnd 0.008226f
C3666 vdd.n1616 gnd 0.01022f
C3667 vdd.n1617 gnd 0.01022f
C3668 vdd.n1618 gnd 0.01022f
C3669 vdd.n1619 gnd 0.01022f
C3670 vdd.n1620 gnd 0.01022f
C3671 vdd.n1621 gnd 0.008226f
C3672 vdd.n1622 gnd 0.01022f
C3673 vdd.n1623 gnd 0.01022f
C3674 vdd.n1624 gnd 0.01022f
C3675 vdd.n1625 gnd 0.01022f
C3676 vdd.n1626 gnd 0.01022f
C3677 vdd.n1627 gnd 0.008226f
C3678 vdd.n1628 gnd 0.01022f
C3679 vdd.n1629 gnd 0.01022f
C3680 vdd.n1630 gnd 0.01022f
C3681 vdd.n1631 gnd 0.01022f
C3682 vdd.n1632 gnd 0.01022f
C3683 vdd.n1633 gnd 0.004319f
C3684 vdd.n1634 gnd 0.01022f
C3685 vdd.n1635 gnd 0.008226f
C3686 vdd.n1636 gnd 0.008226f
C3687 vdd.n1637 gnd 0.008226f
C3688 vdd.n1638 gnd 0.01022f
C3689 vdd.n1639 gnd 0.01022f
C3690 vdd.n1640 gnd 0.01022f
C3691 vdd.n1641 gnd 0.008226f
C3692 vdd.n1642 gnd 0.008226f
C3693 vdd.n1643 gnd 0.008226f
C3694 vdd.n1644 gnd 0.01022f
C3695 vdd.n1645 gnd 0.01022f
C3696 vdd.n1646 gnd 0.01022f
C3697 vdd.n1647 gnd 0.008226f
C3698 vdd.n1648 gnd 0.008226f
C3699 vdd.n1649 gnd 0.008226f
C3700 vdd.n1650 gnd 0.01022f
C3701 vdd.n1651 gnd 0.01022f
C3702 vdd.n1652 gnd 0.01022f
C3703 vdd.n1653 gnd 0.008226f
C3704 vdd.n1654 gnd 0.008226f
C3705 vdd.n1655 gnd 0.008226f
C3706 vdd.n1656 gnd 0.01022f
C3707 vdd.n1657 gnd 0.01022f
C3708 vdd.n1658 gnd 0.01022f
C3709 vdd.n1659 gnd 0.008226f
C3710 vdd.n1660 gnd 0.008226f
C3711 vdd.n1661 gnd 0.008226f
C3712 vdd.n1662 gnd 0.01022f
C3713 vdd.n1663 gnd 0.01022f
C3714 vdd.n1664 gnd 0.01022f
C3715 vdd.n1665 gnd 0.01022f
C3716 vdd.t48 gnd 0.125739f
C3717 vdd.t49 gnd 0.13438f
C3718 vdd.t46 gnd 0.164213f
C3719 vdd.n1666 gnd 0.210498f
C3720 vdd.n1667 gnd 0.177679f
C3721 vdd.n1668 gnd 0.017604f
C3722 vdd.n1669 gnd 0.005594f
C3723 vdd.n1670 gnd 0.008226f
C3724 vdd.n1671 gnd 0.01022f
C3725 vdd.n1672 gnd 0.01022f
C3726 vdd.n1673 gnd 0.01022f
C3727 vdd.n1674 gnd 0.008226f
C3728 vdd.n1675 gnd 0.008226f
C3729 vdd.n1676 gnd 0.008226f
C3730 vdd.n1677 gnd 0.01022f
C3731 vdd.n1678 gnd 0.01022f
C3732 vdd.n1679 gnd 0.01022f
C3733 vdd.n1680 gnd 0.008226f
C3734 vdd.n1681 gnd 0.008226f
C3735 vdd.n1682 gnd 0.008226f
C3736 vdd.n1683 gnd 0.01022f
C3737 vdd.n1684 gnd 0.01022f
C3738 vdd.n1685 gnd 0.01022f
C3739 vdd.n1686 gnd 0.008226f
C3740 vdd.n1687 gnd 0.008226f
C3741 vdd.n1688 gnd 0.008226f
C3742 vdd.n1689 gnd 0.01022f
C3743 vdd.n1690 gnd 0.01022f
C3744 vdd.n1691 gnd 0.01022f
C3745 vdd.n1692 gnd 0.008226f
C3746 vdd.n1693 gnd 0.008226f
C3747 vdd.n1694 gnd 0.008226f
C3748 vdd.n1695 gnd 0.01022f
C3749 vdd.n1696 gnd 0.01022f
C3750 vdd.n1697 gnd 0.01022f
C3751 vdd.n1698 gnd 0.008226f
C3752 vdd.n1699 gnd 0.006869f
C3753 vdd.n1700 gnd 0.01022f
C3754 vdd.n1701 gnd 0.01022f
C3755 vdd.t58 gnd 0.125739f
C3756 vdd.t59 gnd 0.13438f
C3757 vdd.t57 gnd 0.164213f
C3758 vdd.n1702 gnd 0.210498f
C3759 vdd.n1703 gnd 0.177679f
C3760 vdd.n1704 gnd 0.017604f
C3761 vdd.n1705 gnd 0.01022f
C3762 vdd.n1706 gnd 0.01022f
C3763 vdd.n1707 gnd 0.01022f
C3764 vdd.n1708 gnd 0.008226f
C3765 vdd.n1709 gnd 0.008226f
C3766 vdd.n1710 gnd 0.008226f
C3767 vdd.n1711 gnd 0.01022f
C3768 vdd.n1712 gnd 0.01022f
C3769 vdd.n1713 gnd 0.01022f
C3770 vdd.n1714 gnd 0.008226f
C3771 vdd.n1715 gnd 0.008226f
C3772 vdd.n1716 gnd 0.008226f
C3773 vdd.n1717 gnd 0.01022f
C3774 vdd.n1718 gnd 0.01022f
C3775 vdd.n1719 gnd 0.01022f
C3776 vdd.n1720 gnd 0.008226f
C3777 vdd.n1721 gnd 0.008226f
C3778 vdd.n1722 gnd 0.008226f
C3779 vdd.n1723 gnd 0.01022f
C3780 vdd.n1724 gnd 0.01022f
C3781 vdd.n1725 gnd 0.01022f
C3782 vdd.n1726 gnd 0.008226f
C3783 vdd.n1727 gnd 0.008226f
C3784 vdd.n1728 gnd 0.008226f
C3785 vdd.n1729 gnd 0.01022f
C3786 vdd.n1730 gnd 0.01022f
C3787 vdd.n1731 gnd 0.01022f
C3788 vdd.n1732 gnd 0.008226f
C3789 vdd.n1733 gnd 0.006828f
C3790 vdd.n1734 gnd 0.023433f
C3791 vdd.n1736 gnd 2.30831f
C3792 vdd.n1737 gnd 0.023433f
C3793 vdd.n1738 gnd 0.003907f
C3794 vdd.n1739 gnd 0.023433f
C3795 vdd.n1740 gnd 0.023274f
C3796 vdd.n1741 gnd 0.01022f
C3797 vdd.n1742 gnd 0.008226f
C3798 vdd.n1743 gnd 0.01022f
C3799 vdd.t47 gnd 0.522243f
C3800 vdd.n1744 gnd 0.684138f
C3801 vdd.n1745 gnd 0.01022f
C3802 vdd.n1746 gnd 0.008226f
C3803 vdd.n1747 gnd 0.01022f
C3804 vdd.n1748 gnd 0.01022f
C3805 vdd.n1749 gnd 0.01022f
C3806 vdd.n1750 gnd 0.008226f
C3807 vdd.n1751 gnd 0.01022f
C3808 vdd.n1752 gnd 1.04449f
C3809 vdd.n1753 gnd 0.01022f
C3810 vdd.n1754 gnd 0.008226f
C3811 vdd.n1755 gnd 0.01022f
C3812 vdd.n1756 gnd 0.01022f
C3813 vdd.n1757 gnd 0.01022f
C3814 vdd.n1758 gnd 0.008226f
C3815 vdd.n1759 gnd 0.01022f
C3816 vdd.n1760 gnd 0.866923f
C3817 vdd.t108 gnd 0.522243f
C3818 vdd.n1761 gnd 0.600579f
C3819 vdd.n1762 gnd 0.01022f
C3820 vdd.n1763 gnd 0.008226f
C3821 vdd.n1764 gnd 0.01022f
C3822 vdd.n1765 gnd 0.01022f
C3823 vdd.n1766 gnd 0.01022f
C3824 vdd.n1767 gnd 0.008226f
C3825 vdd.n1768 gnd 0.01022f
C3826 vdd.n1769 gnd 0.621469f
C3827 vdd.n1770 gnd 0.01022f
C3828 vdd.n1771 gnd 0.008226f
C3829 vdd.n1772 gnd 0.01022f
C3830 vdd.n1773 gnd 0.01022f
C3831 vdd.n1774 gnd 0.01022f
C3832 vdd.n1775 gnd 0.008226f
C3833 vdd.n1776 gnd 0.01022f
C3834 vdd.n1777 gnd 0.590134f
C3835 vdd.n1778 gnd 0.799031f
C3836 vdd.n1779 gnd 0.01022f
C3837 vdd.n1780 gnd 0.008226f
C3838 vdd.n1781 gnd 0.01022f
C3839 vdd.n1782 gnd 0.01022f
C3840 vdd.n1783 gnd 0.01022f
C3841 vdd.n1784 gnd 0.008226f
C3842 vdd.n1785 gnd 0.01022f
C3843 vdd.n1786 gnd 0.866923f
C3844 vdd.n1787 gnd 0.01022f
C3845 vdd.n1788 gnd 0.008226f
C3846 vdd.n1789 gnd 0.01022f
C3847 vdd.n1790 gnd 0.01022f
C3848 vdd.n1791 gnd 0.01022f
C3849 vdd.n1792 gnd 0.008226f
C3850 vdd.n1793 gnd 0.01022f
C3851 vdd.t4 gnd 0.522243f
C3852 vdd.n1794 gnd 0.757252f
C3853 vdd.n1795 gnd 0.01022f
C3854 vdd.n1796 gnd 0.008226f
C3855 vdd.n1797 gnd 0.01022f
C3856 vdd.n1798 gnd 0.01022f
C3857 vdd.n1799 gnd 0.01022f
C3858 vdd.n1800 gnd 0.008226f
C3859 vdd.n1801 gnd 0.01022f
C3860 vdd.n1802 gnd 0.579689f
C3861 vdd.n1803 gnd 0.01022f
C3862 vdd.n1804 gnd 0.008226f
C3863 vdd.n1805 gnd 0.01022f
C3864 vdd.n1806 gnd 0.01022f
C3865 vdd.n1807 gnd 0.01022f
C3866 vdd.n1808 gnd 0.008226f
C3867 vdd.n1809 gnd 0.01022f
C3868 vdd.n1810 gnd 0.746807f
C3869 vdd.n1811 gnd 0.642358f
C3870 vdd.n1812 gnd 0.01022f
C3871 vdd.n1813 gnd 0.008226f
C3872 vdd.n1814 gnd 0.007855f
C3873 vdd.n1815 gnd 0.005609f
C3874 vdd.n1816 gnd 0.005205f
C3875 vdd.n1817 gnd 0.002879f
C3876 vdd.n1818 gnd 0.006611f
C3877 vdd.n1819 gnd 0.002797f
C3878 vdd.n1820 gnd 0.002961f
C3879 vdd.n1821 gnd 0.005205f
C3880 vdd.n1822 gnd 0.002797f
C3881 vdd.n1823 gnd 0.006611f
C3882 vdd.n1824 gnd 0.002961f
C3883 vdd.n1825 gnd 0.005205f
C3884 vdd.n1826 gnd 0.002797f
C3885 vdd.n1827 gnd 0.004958f
C3886 vdd.n1828 gnd 0.004973f
C3887 vdd.t186 gnd 0.014203f
C3888 vdd.n1829 gnd 0.031601f
C3889 vdd.n1830 gnd 0.164461f
C3890 vdd.n1831 gnd 0.002797f
C3891 vdd.n1832 gnd 0.002961f
C3892 vdd.n1833 gnd 0.006611f
C3893 vdd.n1834 gnd 0.006611f
C3894 vdd.n1835 gnd 0.002961f
C3895 vdd.n1836 gnd 0.002797f
C3896 vdd.n1837 gnd 0.005205f
C3897 vdd.n1838 gnd 0.005205f
C3898 vdd.n1839 gnd 0.002797f
C3899 vdd.n1840 gnd 0.002961f
C3900 vdd.n1841 gnd 0.006611f
C3901 vdd.n1842 gnd 0.006611f
C3902 vdd.n1843 gnd 0.002961f
C3903 vdd.n1844 gnd 0.002797f
C3904 vdd.n1845 gnd 0.005205f
C3905 vdd.n1846 gnd 0.005205f
C3906 vdd.n1847 gnd 0.002797f
C3907 vdd.n1848 gnd 0.002961f
C3908 vdd.n1849 gnd 0.006611f
C3909 vdd.n1850 gnd 0.006611f
C3910 vdd.n1851 gnd 0.01563f
C3911 vdd.n1852 gnd 0.002879f
C3912 vdd.n1853 gnd 0.002797f
C3913 vdd.n1854 gnd 0.013453f
C3914 vdd.n1855 gnd 0.009392f
C3915 vdd.t8 gnd 0.032905f
C3916 vdd.t261 gnd 0.032905f
C3917 vdd.n1856 gnd 0.226146f
C3918 vdd.n1857 gnd 0.177829f
C3919 vdd.t147 gnd 0.032905f
C3920 vdd.t263 gnd 0.032905f
C3921 vdd.n1858 gnd 0.226146f
C3922 vdd.n1859 gnd 0.143507f
C3923 vdd.t153 gnd 0.032905f
C3924 vdd.t246 gnd 0.032905f
C3925 vdd.n1860 gnd 0.226146f
C3926 vdd.n1861 gnd 0.143507f
C3927 vdd.t142 gnd 0.032905f
C3928 vdd.t173 gnd 0.032905f
C3929 vdd.n1862 gnd 0.226146f
C3930 vdd.n1863 gnd 0.143507f
C3931 vdd.t5 gnd 0.032905f
C3932 vdd.t179 gnd 0.032905f
C3933 vdd.n1864 gnd 0.226146f
C3934 vdd.n1865 gnd 0.143507f
C3935 vdd.t157 gnd 0.032905f
C3936 vdd.t139 gnd 0.032905f
C3937 vdd.n1866 gnd 0.226146f
C3938 vdd.n1867 gnd 0.143507f
C3939 vdd.t120 gnd 0.032905f
C3940 vdd.t134 gnd 0.032905f
C3941 vdd.n1868 gnd 0.226146f
C3942 vdd.n1869 gnd 0.143507f
C3943 vdd.n1870 gnd 0.005609f
C3944 vdd.n1871 gnd 0.005205f
C3945 vdd.n1872 gnd 0.002879f
C3946 vdd.n1873 gnd 0.006611f
C3947 vdd.n1874 gnd 0.002797f
C3948 vdd.n1875 gnd 0.002961f
C3949 vdd.n1876 gnd 0.005205f
C3950 vdd.n1877 gnd 0.002797f
C3951 vdd.n1878 gnd 0.006611f
C3952 vdd.n1879 gnd 0.002961f
C3953 vdd.n1880 gnd 0.005205f
C3954 vdd.n1881 gnd 0.002797f
C3955 vdd.n1882 gnd 0.004958f
C3956 vdd.n1883 gnd 0.004973f
C3957 vdd.t129 gnd 0.014203f
C3958 vdd.n1884 gnd 0.031601f
C3959 vdd.n1885 gnd 0.164461f
C3960 vdd.n1886 gnd 0.002797f
C3961 vdd.n1887 gnd 0.002961f
C3962 vdd.n1888 gnd 0.006611f
C3963 vdd.n1889 gnd 0.006611f
C3964 vdd.n1890 gnd 0.002961f
C3965 vdd.n1891 gnd 0.002797f
C3966 vdd.n1892 gnd 0.005205f
C3967 vdd.n1893 gnd 0.005205f
C3968 vdd.n1894 gnd 0.002797f
C3969 vdd.n1895 gnd 0.002961f
C3970 vdd.n1896 gnd 0.006611f
C3971 vdd.n1897 gnd 0.006611f
C3972 vdd.n1898 gnd 0.002961f
C3973 vdd.n1899 gnd 0.002797f
C3974 vdd.n1900 gnd 0.005205f
C3975 vdd.n1901 gnd 0.005205f
C3976 vdd.n1902 gnd 0.002797f
C3977 vdd.n1903 gnd 0.002961f
C3978 vdd.n1904 gnd 0.006611f
C3979 vdd.n1905 gnd 0.006611f
C3980 vdd.n1906 gnd 0.01563f
C3981 vdd.n1907 gnd 0.002879f
C3982 vdd.n1908 gnd 0.002797f
C3983 vdd.n1909 gnd 0.013453f
C3984 vdd.n1910 gnd 0.009098f
C3985 vdd.n1911 gnd 0.10677f
C3986 vdd.n1912 gnd 0.005609f
C3987 vdd.n1913 gnd 0.005205f
C3988 vdd.n1914 gnd 0.002879f
C3989 vdd.n1915 gnd 0.006611f
C3990 vdd.n1916 gnd 0.002797f
C3991 vdd.n1917 gnd 0.002961f
C3992 vdd.n1918 gnd 0.005205f
C3993 vdd.n1919 gnd 0.002797f
C3994 vdd.n1920 gnd 0.006611f
C3995 vdd.n1921 gnd 0.002961f
C3996 vdd.n1922 gnd 0.005205f
C3997 vdd.n1923 gnd 0.002797f
C3998 vdd.n1924 gnd 0.004958f
C3999 vdd.n1925 gnd 0.004973f
C4000 vdd.t243 gnd 0.014203f
C4001 vdd.n1926 gnd 0.031601f
C4002 vdd.n1927 gnd 0.164461f
C4003 vdd.n1928 gnd 0.002797f
C4004 vdd.n1929 gnd 0.002961f
C4005 vdd.n1930 gnd 0.006611f
C4006 vdd.n1931 gnd 0.006611f
C4007 vdd.n1932 gnd 0.002961f
C4008 vdd.n1933 gnd 0.002797f
C4009 vdd.n1934 gnd 0.005205f
C4010 vdd.n1935 gnd 0.005205f
C4011 vdd.n1936 gnd 0.002797f
C4012 vdd.n1937 gnd 0.002961f
C4013 vdd.n1938 gnd 0.006611f
C4014 vdd.n1939 gnd 0.006611f
C4015 vdd.n1940 gnd 0.002961f
C4016 vdd.n1941 gnd 0.002797f
C4017 vdd.n1942 gnd 0.005205f
C4018 vdd.n1943 gnd 0.005205f
C4019 vdd.n1944 gnd 0.002797f
C4020 vdd.n1945 gnd 0.002961f
C4021 vdd.n1946 gnd 0.006611f
C4022 vdd.n1947 gnd 0.006611f
C4023 vdd.n1948 gnd 0.01563f
C4024 vdd.n1949 gnd 0.002879f
C4025 vdd.n1950 gnd 0.002797f
C4026 vdd.n1951 gnd 0.013453f
C4027 vdd.n1952 gnd 0.009392f
C4028 vdd.t7 gnd 0.032905f
C4029 vdd.t189 gnd 0.032905f
C4030 vdd.n1953 gnd 0.226146f
C4031 vdd.n1954 gnd 0.177829f
C4032 vdd.t181 gnd 0.032905f
C4033 vdd.t241 gnd 0.032905f
C4034 vdd.n1955 gnd 0.226146f
C4035 vdd.n1956 gnd 0.143507f
C4036 vdd.t177 gnd 0.032905f
C4037 vdd.t14 gnd 0.032905f
C4038 vdd.n1957 gnd 0.226146f
C4039 vdd.n1958 gnd 0.143507f
C4040 vdd.t185 gnd 0.032905f
C4041 vdd.t245 gnd 0.032905f
C4042 vdd.n1959 gnd 0.226146f
C4043 vdd.n1960 gnd 0.143507f
C4044 vdd.t165 gnd 0.032905f
C4045 vdd.t149 gnd 0.032905f
C4046 vdd.n1961 gnd 0.226146f
C4047 vdd.n1962 gnd 0.143507f
C4048 vdd.t132 gnd 0.032905f
C4049 vdd.t178 gnd 0.032905f
C4050 vdd.n1963 gnd 0.226146f
C4051 vdd.n1964 gnd 0.143507f
C4052 vdd.t119 gnd 0.032905f
C4053 vdd.t166 gnd 0.032905f
C4054 vdd.n1965 gnd 0.226146f
C4055 vdd.n1966 gnd 0.143507f
C4056 vdd.n1967 gnd 0.005609f
C4057 vdd.n1968 gnd 0.005205f
C4058 vdd.n1969 gnd 0.002879f
C4059 vdd.n1970 gnd 0.006611f
C4060 vdd.n1971 gnd 0.002797f
C4061 vdd.n1972 gnd 0.002961f
C4062 vdd.n1973 gnd 0.005205f
C4063 vdd.n1974 gnd 0.002797f
C4064 vdd.n1975 gnd 0.006611f
C4065 vdd.n1976 gnd 0.002961f
C4066 vdd.n1977 gnd 0.005205f
C4067 vdd.n1978 gnd 0.002797f
C4068 vdd.n1979 gnd 0.004958f
C4069 vdd.n1980 gnd 0.004973f
C4070 vdd.t155 gnd 0.014203f
C4071 vdd.n1981 gnd 0.031601f
C4072 vdd.n1982 gnd 0.164461f
C4073 vdd.n1983 gnd 0.002797f
C4074 vdd.n1984 gnd 0.002961f
C4075 vdd.n1985 gnd 0.006611f
C4076 vdd.n1986 gnd 0.006611f
C4077 vdd.n1987 gnd 0.002961f
C4078 vdd.n1988 gnd 0.002797f
C4079 vdd.n1989 gnd 0.005205f
C4080 vdd.n1990 gnd 0.005205f
C4081 vdd.n1991 gnd 0.002797f
C4082 vdd.n1992 gnd 0.002961f
C4083 vdd.n1993 gnd 0.006611f
C4084 vdd.n1994 gnd 0.006611f
C4085 vdd.n1995 gnd 0.002961f
C4086 vdd.n1996 gnd 0.002797f
C4087 vdd.n1997 gnd 0.005205f
C4088 vdd.n1998 gnd 0.005205f
C4089 vdd.n1999 gnd 0.002797f
C4090 vdd.n2000 gnd 0.002961f
C4091 vdd.n2001 gnd 0.006611f
C4092 vdd.n2002 gnd 0.006611f
C4093 vdd.n2003 gnd 0.01563f
C4094 vdd.n2004 gnd 0.002879f
C4095 vdd.n2005 gnd 0.002797f
C4096 vdd.n2006 gnd 0.013453f
C4097 vdd.n2007 gnd 0.009098f
C4098 vdd.n2008 gnd 0.063517f
C4099 vdd.n2009 gnd 0.22887f
C4100 vdd.n2010 gnd 0.005609f
C4101 vdd.n2011 gnd 0.005205f
C4102 vdd.n2012 gnd 0.002879f
C4103 vdd.n2013 gnd 0.006611f
C4104 vdd.n2014 gnd 0.002797f
C4105 vdd.n2015 gnd 0.002961f
C4106 vdd.n2016 gnd 0.005205f
C4107 vdd.n2017 gnd 0.002797f
C4108 vdd.n2018 gnd 0.006611f
C4109 vdd.n2019 gnd 0.002961f
C4110 vdd.n2020 gnd 0.005205f
C4111 vdd.n2021 gnd 0.002797f
C4112 vdd.n2022 gnd 0.004958f
C4113 vdd.n2023 gnd 0.004973f
C4114 vdd.t170 gnd 0.014203f
C4115 vdd.n2024 gnd 0.031601f
C4116 vdd.n2025 gnd 0.164461f
C4117 vdd.n2026 gnd 0.002797f
C4118 vdd.n2027 gnd 0.002961f
C4119 vdd.n2028 gnd 0.006611f
C4120 vdd.n2029 gnd 0.006611f
C4121 vdd.n2030 gnd 0.002961f
C4122 vdd.n2031 gnd 0.002797f
C4123 vdd.n2032 gnd 0.005205f
C4124 vdd.n2033 gnd 0.005205f
C4125 vdd.n2034 gnd 0.002797f
C4126 vdd.n2035 gnd 0.002961f
C4127 vdd.n2036 gnd 0.006611f
C4128 vdd.n2037 gnd 0.006611f
C4129 vdd.n2038 gnd 0.002961f
C4130 vdd.n2039 gnd 0.002797f
C4131 vdd.n2040 gnd 0.005205f
C4132 vdd.n2041 gnd 0.005205f
C4133 vdd.n2042 gnd 0.002797f
C4134 vdd.n2043 gnd 0.002961f
C4135 vdd.n2044 gnd 0.006611f
C4136 vdd.n2045 gnd 0.006611f
C4137 vdd.n2046 gnd 0.01563f
C4138 vdd.n2047 gnd 0.002879f
C4139 vdd.n2048 gnd 0.002797f
C4140 vdd.n2049 gnd 0.013453f
C4141 vdd.n2050 gnd 0.009392f
C4142 vdd.t121 gnd 0.032905f
C4143 vdd.t259 gnd 0.032905f
C4144 vdd.n2051 gnd 0.226146f
C4145 vdd.n2052 gnd 0.177829f
C4146 vdd.t240 gnd 0.032905f
C4147 vdd.t16 gnd 0.032905f
C4148 vdd.n2053 gnd 0.226146f
C4149 vdd.n2054 gnd 0.143507f
C4150 vdd.t256 gnd 0.032905f
C4151 vdd.t113 gnd 0.032905f
C4152 vdd.n2055 gnd 0.226146f
C4153 vdd.n2056 gnd 0.143507f
C4154 vdd.t131 gnd 0.032905f
C4155 vdd.t266 gnd 0.032905f
C4156 vdd.n2057 gnd 0.226146f
C4157 vdd.n2058 gnd 0.143507f
C4158 vdd.t267 gnd 0.032905f
C4159 vdd.t190 gnd 0.032905f
C4160 vdd.n2059 gnd 0.226146f
C4161 vdd.n2060 gnd 0.143507f
C4162 vdd.t124 gnd 0.032905f
C4163 vdd.t258 gnd 0.032905f
C4164 vdd.n2061 gnd 0.226146f
C4165 vdd.n2062 gnd 0.143507f
C4166 vdd.t111 gnd 0.032905f
C4167 vdd.t158 gnd 0.032905f
C4168 vdd.n2063 gnd 0.226146f
C4169 vdd.n2064 gnd 0.143507f
C4170 vdd.n2065 gnd 0.005609f
C4171 vdd.n2066 gnd 0.005205f
C4172 vdd.n2067 gnd 0.002879f
C4173 vdd.n2068 gnd 0.006611f
C4174 vdd.n2069 gnd 0.002797f
C4175 vdd.n2070 gnd 0.002961f
C4176 vdd.n2071 gnd 0.005205f
C4177 vdd.n2072 gnd 0.002797f
C4178 vdd.n2073 gnd 0.006611f
C4179 vdd.n2074 gnd 0.002961f
C4180 vdd.n2075 gnd 0.005205f
C4181 vdd.n2076 gnd 0.002797f
C4182 vdd.n2077 gnd 0.004958f
C4183 vdd.n2078 gnd 0.004973f
C4184 vdd.t109 gnd 0.014203f
C4185 vdd.n2079 gnd 0.031601f
C4186 vdd.n2080 gnd 0.164461f
C4187 vdd.n2081 gnd 0.002797f
C4188 vdd.n2082 gnd 0.002961f
C4189 vdd.n2083 gnd 0.006611f
C4190 vdd.n2084 gnd 0.006611f
C4191 vdd.n2085 gnd 0.002961f
C4192 vdd.n2086 gnd 0.002797f
C4193 vdd.n2087 gnd 0.005205f
C4194 vdd.n2088 gnd 0.005205f
C4195 vdd.n2089 gnd 0.002797f
C4196 vdd.n2090 gnd 0.002961f
C4197 vdd.n2091 gnd 0.006611f
C4198 vdd.n2092 gnd 0.006611f
C4199 vdd.n2093 gnd 0.002961f
C4200 vdd.n2094 gnd 0.002797f
C4201 vdd.n2095 gnd 0.005205f
C4202 vdd.n2096 gnd 0.005205f
C4203 vdd.n2097 gnd 0.002797f
C4204 vdd.n2098 gnd 0.002961f
C4205 vdd.n2099 gnd 0.006611f
C4206 vdd.n2100 gnd 0.006611f
C4207 vdd.n2101 gnd 0.01563f
C4208 vdd.n2102 gnd 0.002879f
C4209 vdd.n2103 gnd 0.002797f
C4210 vdd.n2104 gnd 0.013453f
C4211 vdd.n2105 gnd 0.009098f
C4212 vdd.n2106 gnd 0.063517f
C4213 vdd.n2107 gnd 0.256304f
C4214 vdd.n2108 gnd 2.56833f
C4215 vdd.n2109 gnd 0.602843f
C4216 vdd.n2110 gnd 0.007855f
C4217 vdd.n2111 gnd 0.01022f
C4218 vdd.n2112 gnd 0.008226f
C4219 vdd.n2113 gnd 0.01022f
C4220 vdd.n2114 gnd 0.819921f
C4221 vdd.n2115 gnd 0.01022f
C4222 vdd.n2116 gnd 0.008226f
C4223 vdd.n2117 gnd 0.01022f
C4224 vdd.n2118 gnd 0.01022f
C4225 vdd.n2119 gnd 0.01022f
C4226 vdd.n2120 gnd 0.008226f
C4227 vdd.n2121 gnd 0.01022f
C4228 vdd.t13 gnd 0.522243f
C4229 vdd.n2122 gnd 0.866923f
C4230 vdd.n2123 gnd 0.01022f
C4231 vdd.n2124 gnd 0.008226f
C4232 vdd.n2125 gnd 0.01022f
C4233 vdd.n2126 gnd 0.01022f
C4234 vdd.n2127 gnd 0.01022f
C4235 vdd.n2128 gnd 0.008226f
C4236 vdd.n2129 gnd 0.01022f
C4237 vdd.n2130 gnd 0.736362f
C4238 vdd.n2131 gnd 0.01022f
C4239 vdd.n2132 gnd 0.008226f
C4240 vdd.n2133 gnd 0.01022f
C4241 vdd.n2134 gnd 0.01022f
C4242 vdd.n2135 gnd 0.01022f
C4243 vdd.n2136 gnd 0.008226f
C4244 vdd.n2137 gnd 0.01022f
C4245 vdd.n2138 gnd 0.866923f
C4246 vdd.t15 gnd 0.522243f
C4247 vdd.n2139 gnd 0.5588f
C4248 vdd.n2140 gnd 0.01022f
C4249 vdd.n2141 gnd 0.008226f
C4250 vdd.n2142 gnd 0.01022f
C4251 vdd.n2143 gnd 0.01022f
C4252 vdd.n2144 gnd 0.01022f
C4253 vdd.n2145 gnd 0.008226f
C4254 vdd.n2146 gnd 0.01022f
C4255 vdd.n2147 gnd 0.663248f
C4256 vdd.n2148 gnd 0.01022f
C4257 vdd.n2149 gnd 0.008226f
C4258 vdd.n2150 gnd 0.01022f
C4259 vdd.n2151 gnd 0.01022f
C4260 vdd.n2152 gnd 0.01022f
C4261 vdd.n2153 gnd 0.008226f
C4262 vdd.n2154 gnd 0.01022f
C4263 vdd.n2155 gnd 0.548355f
C4264 vdd.n2156 gnd 0.84081f
C4265 vdd.n2157 gnd 0.01022f
C4266 vdd.n2158 gnd 0.008226f
C4267 vdd.n2159 gnd 0.01022f
C4268 vdd.n2160 gnd 0.01022f
C4269 vdd.n2161 gnd 0.01022f
C4270 vdd.n2162 gnd 0.008226f
C4271 vdd.n2163 gnd 0.01022f
C4272 vdd.n2164 gnd 1.01837f
C4273 vdd.n2165 gnd 0.01022f
C4274 vdd.n2166 gnd 0.008226f
C4275 vdd.n2167 gnd 0.01022f
C4276 vdd.n2168 gnd 0.01022f
C4277 vdd.n2169 gnd 0.023274f
C4278 vdd.n2170 gnd 0.01022f
C4279 vdd.n2171 gnd 0.01022f
C4280 vdd.n2172 gnd 0.008226f
C4281 vdd.n2173 gnd 0.01022f
C4282 vdd.t30 gnd 0.522243f
C4283 vdd.n2174 gnd 0.987038f
C4284 vdd.n2175 gnd 0.01022f
C4285 vdd.n2176 gnd 0.008226f
C4286 vdd.n2177 gnd 0.01022f
C4287 vdd.n2178 gnd 0.01022f
C4288 vdd.n2179 gnd 0.023274f
C4289 vdd.n2180 gnd 0.006828f
C4290 vdd.n2181 gnd 0.023274f
C4291 vdd.n2182 gnd 1.37872f
C4292 vdd.n2183 gnd 0.023274f
C4293 vdd.n2184 gnd 0.023433f
C4294 vdd.n2185 gnd 0.003907f
C4295 vdd.t32 gnd 0.125739f
C4296 vdd.t31 gnd 0.13438f
C4297 vdd.t29 gnd 0.164213f
C4298 vdd.n2186 gnd 0.210498f
C4299 vdd.n2187 gnd 0.176857f
C4300 vdd.n2188 gnd 0.012668f
C4301 vdd.n2189 gnd 0.004319f
C4302 vdd.n2190 gnd 0.00879f
C4303 vdd.n2191 gnd 0.772928f
C4304 vdd.n2193 gnd 0.008226f
C4305 vdd.n2194 gnd 0.008226f
C4306 vdd.n2195 gnd 0.01022f
C4307 vdd.n2197 gnd 0.01022f
C4308 vdd.n2198 gnd 0.01022f
C4309 vdd.n2199 gnd 0.008226f
C4310 vdd.n2200 gnd 0.008226f
C4311 vdd.n2201 gnd 0.008226f
C4312 vdd.n2202 gnd 0.01022f
C4313 vdd.n2204 gnd 0.01022f
C4314 vdd.n2205 gnd 0.01022f
C4315 vdd.n2206 gnd 0.008226f
C4316 vdd.n2207 gnd 0.008226f
C4317 vdd.n2208 gnd 0.008226f
C4318 vdd.n2209 gnd 0.01022f
C4319 vdd.n2211 gnd 0.01022f
C4320 vdd.n2212 gnd 0.01022f
C4321 vdd.n2213 gnd 0.008226f
C4322 vdd.n2214 gnd 0.008226f
C4323 vdd.n2215 gnd 0.008226f
C4324 vdd.n2216 gnd 0.01022f
C4325 vdd.n2218 gnd 0.01022f
C4326 vdd.n2219 gnd 0.01022f
C4327 vdd.n2220 gnd 0.008226f
C4328 vdd.n2221 gnd 0.01022f
C4329 vdd.n2222 gnd 0.01022f
C4330 vdd.n2223 gnd 0.01022f
C4331 vdd.n2224 gnd 0.016782f
C4332 vdd.n2225 gnd 0.005594f
C4333 vdd.n2226 gnd 0.008226f
C4334 vdd.n2227 gnd 0.01022f
C4335 vdd.n2229 gnd 0.01022f
C4336 vdd.n2230 gnd 0.01022f
C4337 vdd.n2231 gnd 0.008226f
C4338 vdd.n2232 gnd 0.008226f
C4339 vdd.n2233 gnd 0.008226f
C4340 vdd.n2234 gnd 0.01022f
C4341 vdd.n2236 gnd 0.01022f
C4342 vdd.n2237 gnd 0.01022f
C4343 vdd.n2238 gnd 0.008226f
C4344 vdd.n2239 gnd 0.008226f
C4345 vdd.n2240 gnd 0.008226f
C4346 vdd.n2241 gnd 0.01022f
C4347 vdd.n2243 gnd 0.01022f
C4348 vdd.n2244 gnd 0.01022f
C4349 vdd.n2245 gnd 0.008226f
C4350 vdd.n2246 gnd 0.008226f
C4351 vdd.n2247 gnd 0.008226f
C4352 vdd.n2248 gnd 0.01022f
C4353 vdd.n2250 gnd 0.01022f
C4354 vdd.n2251 gnd 0.01022f
C4355 vdd.n2252 gnd 0.008226f
C4356 vdd.n2253 gnd 0.008226f
C4357 vdd.n2254 gnd 0.008226f
C4358 vdd.n2255 gnd 0.01022f
C4359 vdd.n2257 gnd 0.01022f
C4360 vdd.n2258 gnd 0.01022f
C4361 vdd.n2259 gnd 0.008226f
C4362 vdd.n2260 gnd 0.01022f
C4363 vdd.n2261 gnd 0.01022f
C4364 vdd.n2262 gnd 0.01022f
C4365 vdd.n2263 gnd 0.016782f
C4366 vdd.n2264 gnd 0.006869f
C4367 vdd.n2265 gnd 0.008226f
C4368 vdd.n2266 gnd 0.01022f
C4369 vdd.n2268 gnd 0.01022f
C4370 vdd.n2269 gnd 0.01022f
C4371 vdd.n2270 gnd 0.008226f
C4372 vdd.n2271 gnd 0.008226f
C4373 vdd.n2272 gnd 0.008226f
C4374 vdd.n2273 gnd 0.01022f
C4375 vdd.n2275 gnd 0.01022f
C4376 vdd.n2276 gnd 0.01022f
C4377 vdd.n2277 gnd 0.008226f
C4378 vdd.n2278 gnd 0.008226f
C4379 vdd.n2279 gnd 0.008226f
C4380 vdd.n2280 gnd 0.01022f
C4381 vdd.n2282 gnd 0.01022f
C4382 vdd.n2283 gnd 0.01022f
C4383 vdd.n2284 gnd 0.008226f
C4384 vdd.n2285 gnd 0.008226f
C4385 vdd.n2286 gnd 0.008226f
C4386 vdd.n2287 gnd 0.01022f
C4387 vdd.n2289 gnd 0.01022f
C4388 vdd.n2290 gnd 0.008226f
C4389 vdd.n2291 gnd 0.008226f
C4390 vdd.n2292 gnd 0.01022f
C4391 vdd.n2294 gnd 0.01022f
C4392 vdd.n2295 gnd 0.01022f
C4393 vdd.n2296 gnd 0.008226f
C4394 vdd.n2297 gnd 0.00879f
C4395 vdd.n2298 gnd 0.772928f
C4396 vdd.n2299 gnd 0.027855f
C4397 vdd.n2300 gnd 0.00695f
C4398 vdd.n2301 gnd 0.00695f
C4399 vdd.n2302 gnd 0.00695f
C4400 vdd.n2303 gnd 0.00695f
C4401 vdd.n2304 gnd 0.00695f
C4402 vdd.n2305 gnd 0.00695f
C4403 vdd.n2306 gnd 0.00695f
C4404 vdd.n2307 gnd 0.00695f
C4405 vdd.n2308 gnd 0.00695f
C4406 vdd.n2309 gnd 0.00695f
C4407 vdd.n2310 gnd 0.00695f
C4408 vdd.n2311 gnd 0.00695f
C4409 vdd.n2312 gnd 0.00695f
C4410 vdd.n2313 gnd 0.00695f
C4411 vdd.n2314 gnd 0.00695f
C4412 vdd.n2315 gnd 0.00695f
C4413 vdd.n2316 gnd 0.00695f
C4414 vdd.n2317 gnd 0.00695f
C4415 vdd.n2318 gnd 0.00695f
C4416 vdd.n2319 gnd 0.00695f
C4417 vdd.n2320 gnd 0.00695f
C4418 vdd.n2321 gnd 0.00695f
C4419 vdd.n2322 gnd 0.00695f
C4420 vdd.n2323 gnd 0.00695f
C4421 vdd.n2324 gnd 0.00695f
C4422 vdd.n2325 gnd 0.00695f
C4423 vdd.n2326 gnd 0.00695f
C4424 vdd.n2327 gnd 0.00695f
C4425 vdd.n2328 gnd 0.00695f
C4426 vdd.n2329 gnd 0.00695f
C4427 vdd.n2330 gnd 0.00695f
C4428 vdd.n2331 gnd 0.016255f
C4429 vdd.n2332 gnd 0.016255f
C4430 vdd.n2334 gnd 8.90946f
C4431 vdd.n2336 gnd 0.016255f
C4432 vdd.n2337 gnd 0.016255f
C4433 vdd.n2338 gnd 0.015224f
C4434 vdd.n2339 gnd 0.00695f
C4435 vdd.n2340 gnd 0.00695f
C4436 vdd.n2341 gnd 0.71025f
C4437 vdd.n2342 gnd 0.00695f
C4438 vdd.n2343 gnd 0.00695f
C4439 vdd.n2344 gnd 0.00695f
C4440 vdd.n2345 gnd 0.00695f
C4441 vdd.n2346 gnd 0.00695f
C4442 vdd.n2347 gnd 0.600579f
C4443 vdd.n2348 gnd 0.00695f
C4444 vdd.n2349 gnd 0.00695f
C4445 vdd.n2350 gnd 0.00695f
C4446 vdd.n2351 gnd 0.00695f
C4447 vdd.n2352 gnd 0.00695f
C4448 vdd.n2353 gnd 0.71025f
C4449 vdd.n2354 gnd 0.00695f
C4450 vdd.n2355 gnd 0.00695f
C4451 vdd.n2356 gnd 0.00695f
C4452 vdd.n2357 gnd 0.00695f
C4453 vdd.n2358 gnd 0.00695f
C4454 vdd.n2359 gnd 0.694583f
C4455 vdd.n2360 gnd 0.00695f
C4456 vdd.n2361 gnd 0.00695f
C4457 vdd.n2362 gnd 0.00695f
C4458 vdd.n2363 gnd 0.00695f
C4459 vdd.n2364 gnd 0.00695f
C4460 vdd.n2365 gnd 0.71025f
C4461 vdd.n2366 gnd 0.00695f
C4462 vdd.n2367 gnd 0.00695f
C4463 vdd.n2368 gnd 0.00695f
C4464 vdd.n2369 gnd 0.00695f
C4465 vdd.n2370 gnd 0.00695f
C4466 vdd.n2371 gnd 0.569244f
C4467 vdd.n2372 gnd 0.00695f
C4468 vdd.n2373 gnd 0.00695f
C4469 vdd.n2374 gnd 0.005928f
C4470 vdd.n2375 gnd 0.020133f
C4471 vdd.n2376 gnd 0.004497f
C4472 vdd.n2377 gnd 0.00695f
C4473 vdd.n2378 gnd 0.412572f
C4474 vdd.n2379 gnd 0.00695f
C4475 vdd.n2380 gnd 0.00695f
C4476 vdd.n2381 gnd 0.00695f
C4477 vdd.n2382 gnd 0.00695f
C4478 vdd.n2383 gnd 0.00695f
C4479 vdd.n2384 gnd 0.454351f
C4480 vdd.n2385 gnd 0.00695f
C4481 vdd.n2386 gnd 0.00695f
C4482 vdd.n2387 gnd 0.00695f
C4483 vdd.n2388 gnd 0.00695f
C4484 vdd.n2389 gnd 0.00695f
C4485 vdd.n2390 gnd 0.611024f
C4486 vdd.n2391 gnd 0.00695f
C4487 vdd.n2392 gnd 0.00695f
C4488 vdd.n2393 gnd 0.00695f
C4489 vdd.n2394 gnd 0.00695f
C4490 vdd.n2395 gnd 0.00695f
C4491 vdd.n2396 gnd 0.584912f
C4492 vdd.n2397 gnd 0.00695f
C4493 vdd.n2398 gnd 0.00695f
C4494 vdd.n2399 gnd 0.00695f
C4495 vdd.n2400 gnd 0.00695f
C4496 vdd.n2401 gnd 0.00695f
C4497 vdd.n2402 gnd 0.428239f
C4498 vdd.n2403 gnd 0.00695f
C4499 vdd.n2404 gnd 0.00695f
C4500 vdd.n2405 gnd 0.00695f
C4501 vdd.n2406 gnd 0.00695f
C4502 vdd.n2407 gnd 0.00695f
C4503 vdd.n2408 gnd 0.224564f
C4504 vdd.n2409 gnd 0.00695f
C4505 vdd.n2410 gnd 0.00695f
C4506 vdd.n2411 gnd 0.00695f
C4507 vdd.n2412 gnd 0.00695f
C4508 vdd.n2413 gnd 0.00695f
C4509 vdd.n2414 gnd 0.370792f
C4510 vdd.n2415 gnd 0.00695f
C4511 vdd.n2416 gnd 0.00695f
C4512 vdd.n2417 gnd 0.00695f
C4513 vdd.n2418 gnd 0.00695f
C4514 vdd.n2419 gnd 0.00695f
C4515 vdd.n2420 gnd 0.71025f
C4516 vdd.n2421 gnd 0.00695f
C4517 vdd.n2422 gnd 0.00695f
C4518 vdd.n2423 gnd 0.00695f
C4519 vdd.n2424 gnd 0.00695f
C4520 vdd.n2425 gnd 0.00695f
C4521 vdd.n2426 gnd 0.00695f
C4522 vdd.n2427 gnd 0.00695f
C4523 vdd.n2428 gnd 0.532687f
C4524 vdd.n2429 gnd 0.00695f
C4525 vdd.n2430 gnd 0.00695f
C4526 vdd.n2431 gnd 0.00695f
C4527 vdd.n2432 gnd 0.00695f
C4528 vdd.n2433 gnd 0.00695f
C4529 vdd.n2434 gnd 0.00695f
C4530 vdd.n2435 gnd 0.443906f
C4531 vdd.n2436 gnd 0.00695f
C4532 vdd.n2437 gnd 0.00695f
C4533 vdd.n2438 gnd 0.00695f
C4534 vdd.n2439 gnd 0.016087f
C4535 vdd.n2440 gnd 0.015392f
C4536 vdd.n2441 gnd 0.00695f
C4537 vdd.n2442 gnd 0.00695f
C4538 vdd.n2443 gnd 0.005366f
C4539 vdd.n2444 gnd 0.00695f
C4540 vdd.n2445 gnd 0.00695f
C4541 vdd.n2446 gnd 0.005059f
C4542 vdd.n2447 gnd 0.00695f
C4543 vdd.n2448 gnd 0.00695f
C4544 vdd.n2449 gnd 0.00695f
C4545 vdd.n2450 gnd 0.00695f
C4546 vdd.n2451 gnd 0.00695f
C4547 vdd.n2452 gnd 0.00695f
C4548 vdd.n2453 gnd 0.00695f
C4549 vdd.n2454 gnd 0.00695f
C4550 vdd.n2455 gnd 0.00695f
C4551 vdd.n2456 gnd 0.00695f
C4552 vdd.n2457 gnd 0.00695f
C4553 vdd.n2458 gnd 0.00695f
C4554 vdd.n2459 gnd 0.00695f
C4555 vdd.n2460 gnd 0.00695f
C4556 vdd.n2461 gnd 0.00695f
C4557 vdd.n2462 gnd 0.00695f
C4558 vdd.n2463 gnd 0.00695f
C4559 vdd.n2464 gnd 0.00695f
C4560 vdd.n2465 gnd 0.00695f
C4561 vdd.n2466 gnd 0.00695f
C4562 vdd.n2467 gnd 0.00695f
C4563 vdd.n2468 gnd 0.00695f
C4564 vdd.n2469 gnd 0.00695f
C4565 vdd.n2470 gnd 0.00695f
C4566 vdd.n2471 gnd 0.00695f
C4567 vdd.n2472 gnd 0.00695f
C4568 vdd.n2473 gnd 0.00695f
C4569 vdd.n2474 gnd 0.00695f
C4570 vdd.n2475 gnd 0.00695f
C4571 vdd.n2476 gnd 0.00695f
C4572 vdd.n2477 gnd 0.00695f
C4573 vdd.n2478 gnd 0.00695f
C4574 vdd.n2479 gnd 0.00695f
C4575 vdd.n2480 gnd 0.00695f
C4576 vdd.n2481 gnd 0.00695f
C4577 vdd.n2482 gnd 0.00695f
C4578 vdd.n2483 gnd 0.00695f
C4579 vdd.n2484 gnd 0.00695f
C4580 vdd.n2485 gnd 0.00695f
C4581 vdd.n2486 gnd 0.00695f
C4582 vdd.n2487 gnd 0.00695f
C4583 vdd.n2488 gnd 0.00695f
C4584 vdd.n2489 gnd 0.00695f
C4585 vdd.n2490 gnd 0.00695f
C4586 vdd.n2491 gnd 0.00695f
C4587 vdd.n2492 gnd 0.00695f
C4588 vdd.n2493 gnd 0.00695f
C4589 vdd.n2494 gnd 0.00695f
C4590 vdd.n2495 gnd 0.00695f
C4591 vdd.n2496 gnd 0.00695f
C4592 vdd.n2497 gnd 0.00695f
C4593 vdd.n2498 gnd 0.00695f
C4594 vdd.n2499 gnd 0.00695f
C4595 vdd.n2500 gnd 0.00695f
C4596 vdd.n2501 gnd 0.00695f
C4597 vdd.n2502 gnd 0.00695f
C4598 vdd.n2503 gnd 0.00695f
C4599 vdd.n2504 gnd 0.00695f
C4600 vdd.n2505 gnd 0.00695f
C4601 vdd.n2506 gnd 0.00695f
C4602 vdd.n2507 gnd 0.016255f
C4603 vdd.n2508 gnd 0.015224f
C4604 vdd.n2509 gnd 0.015224f
C4605 vdd.n2510 gnd 0.846033f
C4606 vdd.n2511 gnd 0.015224f
C4607 vdd.n2512 gnd 0.016255f
C4608 vdd.n2513 gnd 0.015392f
C4609 vdd.n2514 gnd 0.00695f
C4610 vdd.n2515 gnd 0.00695f
C4611 vdd.n2516 gnd 0.00695f
C4612 vdd.n2517 gnd 0.005366f
C4613 vdd.n2518 gnd 0.009933f
C4614 vdd.n2519 gnd 0.005059f
C4615 vdd.n2520 gnd 0.00695f
C4616 vdd.n2521 gnd 0.00695f
C4617 vdd.n2522 gnd 0.00695f
C4618 vdd.n2523 gnd 0.00695f
C4619 vdd.n2524 gnd 0.00695f
C4620 vdd.n2525 gnd 0.00695f
C4621 vdd.n2526 gnd 0.00695f
C4622 vdd.n2527 gnd 0.00695f
C4623 vdd.n2528 gnd 0.00695f
C4624 vdd.n2529 gnd 0.00695f
C4625 vdd.n2530 gnd 0.00695f
C4626 vdd.n2531 gnd 0.00695f
C4627 vdd.n2532 gnd 0.00695f
C4628 vdd.n2533 gnd 0.00695f
C4629 vdd.n2534 gnd 0.00695f
C4630 vdd.n2535 gnd 0.00695f
C4631 vdd.n2536 gnd 0.00695f
C4632 vdd.n2537 gnd 0.00695f
C4633 vdd.n2538 gnd 0.00695f
C4634 vdd.n2539 gnd 0.00695f
C4635 vdd.n2540 gnd 0.00695f
C4636 vdd.n2541 gnd 0.00695f
C4637 vdd.n2542 gnd 0.00695f
C4638 vdd.n2543 gnd 0.00695f
C4639 vdd.n2544 gnd 0.00695f
C4640 vdd.n2545 gnd 0.00695f
C4641 vdd.n2546 gnd 0.00695f
C4642 vdd.n2547 gnd 0.00695f
C4643 vdd.n2548 gnd 0.00695f
C4644 vdd.n2549 gnd 0.00695f
C4645 vdd.n2550 gnd 0.00695f
C4646 vdd.n2551 gnd 0.00695f
C4647 vdd.n2552 gnd 0.00695f
C4648 vdd.n2553 gnd 0.00695f
C4649 vdd.n2554 gnd 0.00695f
C4650 vdd.n2555 gnd 0.00695f
C4651 vdd.n2556 gnd 0.00695f
C4652 vdd.n2557 gnd 0.00695f
C4653 vdd.n2558 gnd 0.00695f
C4654 vdd.n2559 gnd 0.00695f
C4655 vdd.n2560 gnd 0.00695f
C4656 vdd.n2561 gnd 0.00695f
C4657 vdd.n2562 gnd 0.00695f
C4658 vdd.n2563 gnd 0.00695f
C4659 vdd.n2564 gnd 0.00695f
C4660 vdd.n2565 gnd 0.00695f
C4661 vdd.n2566 gnd 0.00695f
C4662 vdd.n2567 gnd 0.00695f
C4663 vdd.n2568 gnd 0.00695f
C4664 vdd.n2569 gnd 0.00695f
C4665 vdd.n2570 gnd 0.00695f
C4666 vdd.n2571 gnd 0.00695f
C4667 vdd.n2572 gnd 0.00695f
C4668 vdd.n2573 gnd 0.00695f
C4669 vdd.n2574 gnd 0.00695f
C4670 vdd.n2575 gnd 0.00695f
C4671 vdd.n2576 gnd 0.00695f
C4672 vdd.n2577 gnd 0.00695f
C4673 vdd.n2578 gnd 0.00695f
C4674 vdd.n2579 gnd 0.00695f
C4675 vdd.n2580 gnd 0.016255f
C4676 vdd.n2581 gnd 0.016255f
C4677 vdd.n2582 gnd 0.866923f
C4678 vdd.t217 gnd 3.08123f
C4679 vdd.t204 gnd 3.08123f
C4680 vdd.n2615 gnd 0.016255f
C4681 vdd.t220 gnd 0.647581f
C4682 vdd.n2616 gnd 0.00695f
C4683 vdd.n2617 gnd 0.00695f
C4684 vdd.t69 gnd 0.280846f
C4685 vdd.t70 gnd 0.28748f
C4686 vdd.t67 gnd 0.183347f
C4687 vdd.n2618 gnd 0.099089f
C4688 vdd.n2619 gnd 0.056206f
C4689 vdd.n2620 gnd 0.00695f
C4690 vdd.t76 gnd 0.280846f
C4691 vdd.t77 gnd 0.28748f
C4692 vdd.t75 gnd 0.183347f
C4693 vdd.n2621 gnd 0.099089f
C4694 vdd.n2622 gnd 0.056206f
C4695 vdd.n2623 gnd 0.009933f
C4696 vdd.n2624 gnd 0.00695f
C4697 vdd.n2625 gnd 0.00695f
C4698 vdd.n2626 gnd 0.00695f
C4699 vdd.n2627 gnd 0.00695f
C4700 vdd.n2628 gnd 0.00695f
C4701 vdd.n2629 gnd 0.00695f
C4702 vdd.n2630 gnd 0.00695f
C4703 vdd.n2631 gnd 0.00695f
C4704 vdd.n2632 gnd 0.00695f
C4705 vdd.n2633 gnd 0.00695f
C4706 vdd.n2634 gnd 0.00695f
C4707 vdd.n2635 gnd 0.00695f
C4708 vdd.n2636 gnd 0.00695f
C4709 vdd.n2637 gnd 0.00695f
C4710 vdd.n2638 gnd 0.00695f
C4711 vdd.n2639 gnd 0.00695f
C4712 vdd.n2640 gnd 0.00695f
C4713 vdd.n2641 gnd 0.00695f
C4714 vdd.n2642 gnd 0.00695f
C4715 vdd.n2643 gnd 0.00695f
C4716 vdd.n2644 gnd 0.00695f
C4717 vdd.n2645 gnd 0.00695f
C4718 vdd.n2646 gnd 0.00695f
C4719 vdd.n2647 gnd 0.00695f
C4720 vdd.n2648 gnd 0.00695f
C4721 vdd.n2649 gnd 0.00695f
C4722 vdd.n2650 gnd 0.00695f
C4723 vdd.n2651 gnd 0.00695f
C4724 vdd.n2652 gnd 0.00695f
C4725 vdd.n2653 gnd 0.00695f
C4726 vdd.n2654 gnd 0.00695f
C4727 vdd.n2655 gnd 0.00695f
C4728 vdd.n2656 gnd 0.00695f
C4729 vdd.n2657 gnd 0.00695f
C4730 vdd.n2658 gnd 0.00695f
C4731 vdd.n2659 gnd 0.00695f
C4732 vdd.n2660 gnd 0.00695f
C4733 vdd.n2661 gnd 0.00695f
C4734 vdd.n2662 gnd 0.00695f
C4735 vdd.n2663 gnd 0.00695f
C4736 vdd.n2664 gnd 0.00695f
C4737 vdd.n2665 gnd 0.00695f
C4738 vdd.n2666 gnd 0.00695f
C4739 vdd.n2667 gnd 0.00695f
C4740 vdd.n2668 gnd 0.00695f
C4741 vdd.n2669 gnd 0.00695f
C4742 vdd.n2670 gnd 0.00695f
C4743 vdd.n2671 gnd 0.00695f
C4744 vdd.n2672 gnd 0.00695f
C4745 vdd.n2673 gnd 0.00695f
C4746 vdd.n2674 gnd 0.00695f
C4747 vdd.n2675 gnd 0.00695f
C4748 vdd.n2676 gnd 0.00695f
C4749 vdd.n2677 gnd 0.00695f
C4750 vdd.n2678 gnd 0.00695f
C4751 vdd.n2679 gnd 0.00695f
C4752 vdd.n2680 gnd 0.00695f
C4753 vdd.n2681 gnd 0.00695f
C4754 vdd.n2682 gnd 0.005059f
C4755 vdd.n2683 gnd 0.00695f
C4756 vdd.n2684 gnd 0.00695f
C4757 vdd.n2685 gnd 0.005366f
C4758 vdd.n2686 gnd 0.00695f
C4759 vdd.n2687 gnd 0.00695f
C4760 vdd.n2688 gnd 0.016255f
C4761 vdd.n2689 gnd 0.015224f
C4762 vdd.n2690 gnd 0.015224f
C4763 vdd.n2691 gnd 0.00695f
C4764 vdd.n2692 gnd 0.00695f
C4765 vdd.n2693 gnd 0.00695f
C4766 vdd.n2694 gnd 0.00695f
C4767 vdd.n2695 gnd 0.00695f
C4768 vdd.n2696 gnd 0.00695f
C4769 vdd.n2697 gnd 0.00695f
C4770 vdd.n2698 gnd 0.00695f
C4771 vdd.n2699 gnd 0.00695f
C4772 vdd.n2700 gnd 0.00695f
C4773 vdd.n2701 gnd 0.00695f
C4774 vdd.n2702 gnd 0.00695f
C4775 vdd.n2703 gnd 0.00695f
C4776 vdd.n2704 gnd 0.00695f
C4777 vdd.n2705 gnd 0.00695f
C4778 vdd.n2706 gnd 0.00695f
C4779 vdd.n2707 gnd 0.00695f
C4780 vdd.n2708 gnd 0.00695f
C4781 vdd.n2709 gnd 0.00695f
C4782 vdd.n2710 gnd 0.00695f
C4783 vdd.n2711 gnd 0.00695f
C4784 vdd.n2712 gnd 0.00695f
C4785 vdd.n2713 gnd 0.00695f
C4786 vdd.n2714 gnd 0.00695f
C4787 vdd.n2715 gnd 0.00695f
C4788 vdd.n2716 gnd 0.00695f
C4789 vdd.n2717 gnd 0.00695f
C4790 vdd.n2718 gnd 0.00695f
C4791 vdd.n2719 gnd 0.00695f
C4792 vdd.n2720 gnd 0.00695f
C4793 vdd.n2721 gnd 0.00695f
C4794 vdd.n2722 gnd 0.00695f
C4795 vdd.n2723 gnd 0.00695f
C4796 vdd.n2724 gnd 0.00695f
C4797 vdd.n2725 gnd 0.00695f
C4798 vdd.n2726 gnd 0.00695f
C4799 vdd.n2727 gnd 0.00695f
C4800 vdd.n2728 gnd 0.00695f
C4801 vdd.n2729 gnd 0.00695f
C4802 vdd.n2730 gnd 0.00695f
C4803 vdd.n2731 gnd 0.00695f
C4804 vdd.n2732 gnd 0.00695f
C4805 vdd.n2733 gnd 0.00695f
C4806 vdd.n2734 gnd 0.00695f
C4807 vdd.n2735 gnd 0.00695f
C4808 vdd.n2736 gnd 0.00695f
C4809 vdd.n2737 gnd 0.00695f
C4810 vdd.n2738 gnd 0.00695f
C4811 vdd.n2739 gnd 0.00695f
C4812 vdd.n2740 gnd 0.00695f
C4813 vdd.n2741 gnd 0.00695f
C4814 vdd.n2742 gnd 0.00695f
C4815 vdd.n2743 gnd 0.00695f
C4816 vdd.n2744 gnd 0.00695f
C4817 vdd.n2745 gnd 0.00695f
C4818 vdd.n2746 gnd 0.00695f
C4819 vdd.n2747 gnd 0.00695f
C4820 vdd.n2748 gnd 0.00695f
C4821 vdd.n2749 gnd 0.00695f
C4822 vdd.n2750 gnd 0.00695f
C4823 vdd.n2751 gnd 0.00695f
C4824 vdd.n2752 gnd 0.00695f
C4825 vdd.n2753 gnd 0.00695f
C4826 vdd.n2754 gnd 0.00695f
C4827 vdd.n2755 gnd 0.00695f
C4828 vdd.n2756 gnd 0.00695f
C4829 vdd.n2757 gnd 0.00695f
C4830 vdd.n2758 gnd 0.00695f
C4831 vdd.n2759 gnd 0.00695f
C4832 vdd.n2760 gnd 0.00695f
C4833 vdd.n2761 gnd 0.00695f
C4834 vdd.n2762 gnd 0.00695f
C4835 vdd.n2763 gnd 0.00695f
C4836 vdd.n2764 gnd 0.224564f
C4837 vdd.n2765 gnd 0.00695f
C4838 vdd.n2766 gnd 0.00695f
C4839 vdd.n2767 gnd 0.00695f
C4840 vdd.n2768 gnd 0.00695f
C4841 vdd.n2769 gnd 0.00695f
C4842 vdd.n2770 gnd 0.00695f
C4843 vdd.n2771 gnd 0.00695f
C4844 vdd.n2772 gnd 0.00695f
C4845 vdd.n2773 gnd 0.00695f
C4846 vdd.n2774 gnd 0.00695f
C4847 vdd.n2775 gnd 0.00695f
C4848 vdd.n2776 gnd 0.00695f
C4849 vdd.n2777 gnd 0.00695f
C4850 vdd.n2778 gnd 0.00695f
C4851 vdd.n2779 gnd 0.443906f
C4852 vdd.n2780 gnd 0.00695f
C4853 vdd.n2781 gnd 0.00695f
C4854 vdd.n2782 gnd 0.00695f
C4855 vdd.n2783 gnd 0.015224f
C4856 vdd.n2784 gnd 0.015224f
C4857 vdd.n2785 gnd 0.016255f
C4858 vdd.n2786 gnd 0.016255f
C4859 vdd.n2787 gnd 0.00695f
C4860 vdd.n2788 gnd 0.00695f
C4861 vdd.n2789 gnd 0.00695f
C4862 vdd.n2790 gnd 0.005366f
C4863 vdd.n2791 gnd 0.009933f
C4864 vdd.n2792 gnd 0.005059f
C4865 vdd.n2793 gnd 0.00695f
C4866 vdd.n2794 gnd 0.00695f
C4867 vdd.n2795 gnd 0.00695f
C4868 vdd.n2796 gnd 0.00695f
C4869 vdd.n2797 gnd 0.00695f
C4870 vdd.n2798 gnd 0.00695f
C4871 vdd.n2799 gnd 0.00695f
C4872 vdd.n2800 gnd 0.00695f
C4873 vdd.n2801 gnd 0.00695f
C4874 vdd.n2802 gnd 0.00695f
C4875 vdd.n2803 gnd 0.00695f
C4876 vdd.n2804 gnd 0.00695f
C4877 vdd.n2805 gnd 0.00695f
C4878 vdd.n2806 gnd 0.00695f
C4879 vdd.n2807 gnd 0.00695f
C4880 vdd.n2808 gnd 0.00695f
C4881 vdd.n2809 gnd 0.00695f
C4882 vdd.n2810 gnd 0.00695f
C4883 vdd.n2811 gnd 0.00695f
C4884 vdd.n2812 gnd 0.00695f
C4885 vdd.n2813 gnd 0.00695f
C4886 vdd.n2814 gnd 0.00695f
C4887 vdd.n2815 gnd 0.00695f
C4888 vdd.n2816 gnd 0.00695f
C4889 vdd.n2817 gnd 0.00695f
C4890 vdd.n2818 gnd 0.00695f
C4891 vdd.n2819 gnd 0.00695f
C4892 vdd.n2820 gnd 0.00695f
C4893 vdd.n2821 gnd 0.00695f
C4894 vdd.n2822 gnd 0.00695f
C4895 vdd.n2823 gnd 0.00695f
C4896 vdd.n2824 gnd 0.00695f
C4897 vdd.n2825 gnd 0.00695f
C4898 vdd.n2826 gnd 0.00695f
C4899 vdd.n2827 gnd 0.00695f
C4900 vdd.n2828 gnd 0.00695f
C4901 vdd.n2829 gnd 0.00695f
C4902 vdd.n2830 gnd 0.00695f
C4903 vdd.n2831 gnd 0.00695f
C4904 vdd.n2832 gnd 0.00695f
C4905 vdd.n2833 gnd 0.00695f
C4906 vdd.n2834 gnd 0.00695f
C4907 vdd.n2835 gnd 0.00695f
C4908 vdd.n2836 gnd 0.00695f
C4909 vdd.n2837 gnd 0.00695f
C4910 vdd.n2838 gnd 0.00695f
C4911 vdd.n2839 gnd 0.00695f
C4912 vdd.n2840 gnd 0.00695f
C4913 vdd.n2841 gnd 0.00695f
C4914 vdd.n2842 gnd 0.00695f
C4915 vdd.n2843 gnd 0.00695f
C4916 vdd.n2844 gnd 0.00695f
C4917 vdd.n2845 gnd 0.00695f
C4918 vdd.n2846 gnd 0.00695f
C4919 vdd.n2847 gnd 0.00695f
C4920 vdd.n2848 gnd 0.00695f
C4921 vdd.n2849 gnd 0.00695f
C4922 vdd.n2850 gnd 0.00695f
C4923 vdd.n2851 gnd 0.00695f
C4924 vdd.n2852 gnd 0.016255f
C4925 vdd.n2853 gnd 0.016255f
C4926 vdd.n2855 gnd 0.866923f
C4927 vdd.n2857 gnd 0.016255f
C4928 vdd.n2858 gnd 0.016255f
C4929 vdd.n2859 gnd 0.015224f
C4930 vdd.n2860 gnd 0.00695f
C4931 vdd.n2861 gnd 0.00695f
C4932 vdd.n2862 gnd 0.376015f
C4933 vdd.n2863 gnd 0.00695f
C4934 vdd.n2864 gnd 0.00695f
C4935 vdd.n2865 gnd 0.00695f
C4936 vdd.n2866 gnd 0.00695f
C4937 vdd.n2867 gnd 0.00695f
C4938 vdd.n2868 gnd 0.423016f
C4939 vdd.n2869 gnd 0.00695f
C4940 vdd.n2870 gnd 0.00695f
C4941 vdd.n2871 gnd 0.00695f
C4942 vdd.n2872 gnd 0.00695f
C4943 vdd.n2873 gnd 0.00695f
C4944 vdd.n2874 gnd 0.71025f
C4945 vdd.n2875 gnd 0.00695f
C4946 vdd.n2876 gnd 0.00695f
C4947 vdd.n2877 gnd 0.00695f
C4948 vdd.n2878 gnd 0.00695f
C4949 vdd.n2879 gnd 0.00695f
C4950 vdd.n2880 gnd 0.470018f
C4951 vdd.n2881 gnd 0.00695f
C4952 vdd.n2882 gnd 0.00695f
C4953 vdd.n2883 gnd 0.00695f
C4954 vdd.n2884 gnd 0.00695f
C4955 vdd.n2885 gnd 0.00695f
C4956 vdd.n2886 gnd 0.626691f
C4957 vdd.n2887 gnd 0.00695f
C4958 vdd.n2888 gnd 0.00695f
C4959 vdd.n2889 gnd 0.00695f
C4960 vdd.n2890 gnd 0.00695f
C4961 vdd.n2891 gnd 0.00695f
C4962 vdd.n2892 gnd 0.569244f
C4963 vdd.n2893 gnd 0.00695f
C4964 vdd.n2894 gnd 0.00695f
C4965 vdd.n2895 gnd 0.00695f
C4966 vdd.n2896 gnd 0.00695f
C4967 vdd.n2897 gnd 0.00695f
C4968 vdd.n2898 gnd 0.412572f
C4969 vdd.n2899 gnd 0.00695f
C4970 vdd.n2900 gnd 0.00695f
C4971 vdd.n2901 gnd 0.00695f
C4972 vdd.n2902 gnd 0.00695f
C4973 vdd.n2903 gnd 0.00695f
C4974 vdd.n2904 gnd 0.224564f
C4975 vdd.n2905 gnd 0.00695f
C4976 vdd.n2906 gnd 0.00695f
C4977 vdd.n2907 gnd 0.00695f
C4978 vdd.n2908 gnd 0.00695f
C4979 vdd.n2909 gnd 0.00695f
C4980 vdd.n2910 gnd 0.611024f
C4981 vdd.n2911 gnd 0.00695f
C4982 vdd.n2912 gnd 0.00695f
C4983 vdd.n2913 gnd 0.00695f
C4984 vdd.n2914 gnd 0.00695f
C4985 vdd.n2915 gnd 0.00695f
C4986 vdd.n2916 gnd 0.71025f
C4987 vdd.n2917 gnd 0.00695f
C4988 vdd.n2918 gnd 0.00695f
C4989 vdd.n2919 gnd 0.004497f
C4990 vdd.n2920 gnd 0.020133f
C4991 vdd.n2921 gnd 0.005928f
C4992 vdd.n2922 gnd 0.00695f
C4993 vdd.n2923 gnd 0.605801f
C4994 vdd.n2924 gnd 0.00695f
C4995 vdd.n2925 gnd 0.00695f
C4996 vdd.n2926 gnd 0.00695f
C4997 vdd.n2927 gnd 0.00695f
C4998 vdd.n2928 gnd 0.00695f
C4999 vdd.n2929 gnd 0.49613f
C5000 vdd.n2930 gnd 0.00695f
C5001 vdd.n2931 gnd 0.00695f
C5002 vdd.n2932 gnd 0.00695f
C5003 vdd.n2933 gnd 0.00695f
C5004 vdd.n2934 gnd 0.00695f
C5005 vdd.n2935 gnd 0.370792f
C5006 vdd.n2936 gnd 0.00695f
C5007 vdd.n2937 gnd 0.00695f
C5008 vdd.n2938 gnd 0.00695f
C5009 vdd.n2939 gnd 0.00695f
C5010 vdd.n2940 gnd 0.00695f
C5011 vdd.n2941 gnd 0.71025f
C5012 vdd.n2942 gnd 0.00695f
C5013 vdd.n2943 gnd 0.00695f
C5014 vdd.n2944 gnd 0.00695f
C5015 vdd.n2945 gnd 0.00695f
C5016 vdd.n2946 gnd 0.00695f
C5017 vdd.n2947 gnd 0.00695f
C5018 vdd.n2949 gnd 0.00695f
C5019 vdd.n2950 gnd 0.00695f
C5020 vdd.n2952 gnd 0.00695f
C5021 vdd.n2953 gnd 0.00695f
C5022 vdd.n2956 gnd 0.00695f
C5023 vdd.n2957 gnd 0.00695f
C5024 vdd.n2958 gnd 0.00695f
C5025 vdd.n2959 gnd 0.00695f
C5026 vdd.n2961 gnd 0.00695f
C5027 vdd.n2962 gnd 0.00695f
C5028 vdd.n2963 gnd 0.00695f
C5029 vdd.n2964 gnd 0.00695f
C5030 vdd.n2965 gnd 0.00695f
C5031 vdd.n2966 gnd 0.00695f
C5032 vdd.n2968 gnd 0.00695f
C5033 vdd.n2969 gnd 0.00695f
C5034 vdd.n2970 gnd 0.00695f
C5035 vdd.n2971 gnd 0.00695f
C5036 vdd.n2972 gnd 0.00695f
C5037 vdd.n2973 gnd 0.00695f
C5038 vdd.n2975 gnd 0.00695f
C5039 vdd.n2976 gnd 0.00695f
C5040 vdd.n2977 gnd 0.00695f
C5041 vdd.n2978 gnd 0.00695f
C5042 vdd.n2979 gnd 0.00695f
C5043 vdd.n2980 gnd 0.00695f
C5044 vdd.n2982 gnd 0.00695f
C5045 vdd.n2983 gnd 0.016255f
C5046 vdd.n2984 gnd 0.016255f
C5047 vdd.n2985 gnd 0.015224f
C5048 vdd.n2986 gnd 0.00695f
C5049 vdd.n2987 gnd 0.00695f
C5050 vdd.n2988 gnd 0.00695f
C5051 vdd.n2989 gnd 0.00695f
C5052 vdd.n2990 gnd 0.00695f
C5053 vdd.n2991 gnd 0.00695f
C5054 vdd.n2992 gnd 0.71025f
C5055 vdd.n2993 gnd 0.00695f
C5056 vdd.n2994 gnd 0.00695f
C5057 vdd.n2995 gnd 0.00695f
C5058 vdd.n2996 gnd 0.00695f
C5059 vdd.n2997 gnd 0.00695f
C5060 vdd.n2998 gnd 0.464796f
C5061 vdd.n2999 gnd 0.00695f
C5062 vdd.n3000 gnd 0.00695f
C5063 vdd.n3001 gnd 0.00695f
C5064 vdd.n3002 gnd 0.016087f
C5065 vdd.n3004 gnd 0.016255f
C5066 vdd.n3005 gnd 0.015392f
C5067 vdd.n3006 gnd 0.00695f
C5068 vdd.n3007 gnd 0.005366f
C5069 vdd.n3008 gnd 0.00695f
C5070 vdd.n3010 gnd 0.00695f
C5071 vdd.n3011 gnd 0.00695f
C5072 vdd.n3012 gnd 0.00695f
C5073 vdd.n3013 gnd 0.00695f
C5074 vdd.n3014 gnd 0.00695f
C5075 vdd.n3015 gnd 0.00695f
C5076 vdd.n3017 gnd 0.00695f
C5077 vdd.n3018 gnd 0.00695f
C5078 vdd.n3019 gnd 0.00695f
C5079 vdd.n3020 gnd 0.00695f
C5080 vdd.n3021 gnd 0.00695f
C5081 vdd.n3022 gnd 0.00695f
C5082 vdd.n3024 gnd 0.00695f
C5083 vdd.n3025 gnd 0.00695f
C5084 vdd.n3026 gnd 0.00695f
C5085 vdd.n3027 gnd 0.00695f
C5086 vdd.n3028 gnd 0.00695f
C5087 vdd.n3029 gnd 0.00695f
C5088 vdd.n3031 gnd 0.00695f
C5089 vdd.n3032 gnd 0.00695f
C5090 vdd.n3033 gnd 0.00695f
C5091 vdd.n3034 gnd 0.776915f
C5092 vdd.n3035 gnd 0.023869f
C5093 vdd.n3036 gnd 0.00695f
C5094 vdd.n3037 gnd 0.00695f
C5095 vdd.n3039 gnd 0.00695f
C5096 vdd.n3040 gnd 0.00695f
C5097 vdd.n3041 gnd 0.00695f
C5098 vdd.n3042 gnd 0.00695f
C5099 vdd.n3043 gnd 0.00695f
C5100 vdd.n3044 gnd 0.00695f
C5101 vdd.n3046 gnd 0.00695f
C5102 vdd.n3047 gnd 0.00695f
C5103 vdd.n3048 gnd 0.00695f
C5104 vdd.n3049 gnd 0.00695f
C5105 vdd.n3050 gnd 0.00695f
C5106 vdd.n3051 gnd 0.00695f
C5107 vdd.n3053 gnd 0.00695f
C5108 vdd.n3054 gnd 0.00695f
C5109 vdd.n3055 gnd 0.00695f
C5110 vdd.n3056 gnd 0.00695f
C5111 vdd.n3057 gnd 0.00695f
C5112 vdd.n3058 gnd 0.00695f
C5113 vdd.n3060 gnd 0.00695f
C5114 vdd.n3061 gnd 0.00695f
C5115 vdd.n3063 gnd 0.00695f
C5116 vdd.n3064 gnd 0.00695f
C5117 vdd.n3065 gnd 0.016255f
C5118 vdd.n3066 gnd 0.015224f
C5119 vdd.n3067 gnd 0.015224f
C5120 vdd.n3068 gnd 1.00271f
C5121 vdd.n3069 gnd 0.015224f
C5122 vdd.n3070 gnd 0.016255f
C5123 vdd.n3071 gnd 0.015392f
C5124 vdd.n3072 gnd 0.00695f
C5125 vdd.n3073 gnd 0.005366f
C5126 vdd.n3074 gnd 0.00695f
C5127 vdd.n3076 gnd 0.00695f
C5128 vdd.n3077 gnd 0.00695f
C5129 vdd.n3078 gnd 0.00695f
C5130 vdd.n3079 gnd 0.00695f
C5131 vdd.n3080 gnd 0.00695f
C5132 vdd.n3081 gnd 0.00695f
C5133 vdd.n3083 gnd 0.00695f
C5134 vdd.n3084 gnd 0.00695f
C5135 vdd.n3085 gnd 0.00695f
C5136 vdd.n3086 gnd 0.00695f
C5137 vdd.n3087 gnd 0.00695f
C5138 vdd.n3088 gnd 0.00695f
C5139 vdd.n3090 gnd 0.00695f
C5140 vdd.n3091 gnd 0.00695f
C5141 vdd.n3092 gnd 0.00695f
C5142 vdd.n3093 gnd 0.00695f
C5143 vdd.n3094 gnd 0.00695f
C5144 vdd.n3095 gnd 0.00695f
C5145 vdd.n3097 gnd 0.00695f
C5146 vdd.n3098 gnd 0.00695f
C5147 vdd.n3100 gnd 0.00695f
C5148 vdd.n3101 gnd 0.023869f
C5149 vdd.n3102 gnd 0.776915f
C5150 vdd.n3103 gnd 0.00879f
C5151 vdd.n3104 gnd 0.003907f
C5152 vdd.t27 gnd 0.125739f
C5153 vdd.t28 gnd 0.13438f
C5154 vdd.t25 gnd 0.164213f
C5155 vdd.n3105 gnd 0.210498f
C5156 vdd.n3106 gnd 0.176857f
C5157 vdd.n3107 gnd 0.012668f
C5158 vdd.n3108 gnd 0.01022f
C5159 vdd.n3109 gnd 0.004319f
C5160 vdd.n3110 gnd 0.008226f
C5161 vdd.n3111 gnd 0.01022f
C5162 vdd.n3112 gnd 0.01022f
C5163 vdd.n3113 gnd 0.008226f
C5164 vdd.n3114 gnd 0.008226f
C5165 vdd.n3115 gnd 0.01022f
C5166 vdd.n3117 gnd 0.01022f
C5167 vdd.n3118 gnd 0.008226f
C5168 vdd.n3119 gnd 0.008226f
C5169 vdd.n3120 gnd 0.008226f
C5170 vdd.n3121 gnd 0.01022f
C5171 vdd.n3123 gnd 0.01022f
C5172 vdd.n3125 gnd 0.01022f
C5173 vdd.n3126 gnd 0.008226f
C5174 vdd.n3127 gnd 0.008226f
C5175 vdd.n3128 gnd 0.008226f
C5176 vdd.n3129 gnd 0.01022f
C5177 vdd.n3131 gnd 0.01022f
C5178 vdd.n3133 gnd 0.01022f
C5179 vdd.n3134 gnd 0.008226f
C5180 vdd.n3135 gnd 0.008226f
C5181 vdd.n3136 gnd 0.008226f
C5182 vdd.n3137 gnd 0.01022f
C5183 vdd.n3139 gnd 0.01022f
C5184 vdd.n3140 gnd 0.01022f
C5185 vdd.n3141 gnd 0.008226f
C5186 vdd.n3142 gnd 0.008226f
C5187 vdd.n3143 gnd 0.01022f
C5188 vdd.n3144 gnd 0.01022f
C5189 vdd.n3146 gnd 0.01022f
C5190 vdd.n3147 gnd 0.008226f
C5191 vdd.n3148 gnd 0.01022f
C5192 vdd.n3149 gnd 0.01022f
C5193 vdd.n3150 gnd 0.01022f
C5194 vdd.n3151 gnd 0.016782f
C5195 vdd.n3152 gnd 0.005594f
C5196 vdd.n3153 gnd 0.01022f
C5197 vdd.n3155 gnd 0.01022f
C5198 vdd.n3157 gnd 0.01022f
C5199 vdd.n3158 gnd 0.008226f
C5200 vdd.n3159 gnd 0.008226f
C5201 vdd.n3160 gnd 0.008226f
C5202 vdd.n3161 gnd 0.01022f
C5203 vdd.n3163 gnd 0.01022f
C5204 vdd.n3165 gnd 0.01022f
C5205 vdd.n3166 gnd 0.008226f
C5206 vdd.n3167 gnd 0.008226f
C5207 vdd.n3168 gnd 0.008226f
C5208 vdd.n3169 gnd 0.01022f
C5209 vdd.n3171 gnd 0.01022f
C5210 vdd.n3173 gnd 0.01022f
C5211 vdd.n3174 gnd 0.008226f
C5212 vdd.n3175 gnd 0.008226f
C5213 vdd.n3176 gnd 0.008226f
C5214 vdd.n3177 gnd 0.01022f
C5215 vdd.n3179 gnd 0.01022f
C5216 vdd.n3181 gnd 0.01022f
C5217 vdd.n3182 gnd 0.008226f
C5218 vdd.n3183 gnd 0.008226f
C5219 vdd.n3184 gnd 0.008226f
C5220 vdd.n3185 gnd 0.01022f
C5221 vdd.n3187 gnd 0.01022f
C5222 vdd.n3189 gnd 0.01022f
C5223 vdd.n3190 gnd 0.008226f
C5224 vdd.n3191 gnd 0.008226f
C5225 vdd.n3192 gnd 0.006869f
C5226 vdd.n3193 gnd 0.01022f
C5227 vdd.n3195 gnd 0.01022f
C5228 vdd.n3197 gnd 0.01022f
C5229 vdd.n3198 gnd 0.006869f
C5230 vdd.n3199 gnd 0.008226f
C5231 vdd.n3200 gnd 0.008226f
C5232 vdd.n3201 gnd 0.01022f
C5233 vdd.n3203 gnd 0.01022f
C5234 vdd.n3205 gnd 0.01022f
C5235 vdd.n3206 gnd 0.008226f
C5236 vdd.n3207 gnd 0.008226f
C5237 vdd.n3208 gnd 0.008226f
C5238 vdd.n3209 gnd 0.01022f
C5239 vdd.n3211 gnd 0.01022f
C5240 vdd.n3213 gnd 0.01022f
C5241 vdd.n3214 gnd 0.008226f
C5242 vdd.n3215 gnd 0.008226f
C5243 vdd.n3216 gnd 0.008226f
C5244 vdd.n3217 gnd 0.01022f
C5245 vdd.n3219 gnd 0.01022f
C5246 vdd.n3220 gnd 0.01022f
C5247 vdd.n3221 gnd 0.008226f
C5248 vdd.n3222 gnd 0.008226f
C5249 vdd.n3223 gnd 0.01022f
C5250 vdd.n3224 gnd 0.01022f
C5251 vdd.n3225 gnd 0.008226f
C5252 vdd.n3226 gnd 0.008226f
C5253 vdd.n3227 gnd 0.01022f
C5254 vdd.n3228 gnd 0.01022f
C5255 vdd.n3230 gnd 0.01022f
C5256 vdd.n3231 gnd 0.008226f
C5257 vdd.n3232 gnd 0.006828f
C5258 vdd.n3233 gnd 0.023433f
C5259 vdd.n3234 gnd 0.023274f
C5260 vdd.n3235 gnd 0.006828f
C5261 vdd.n3236 gnd 0.023274f
C5262 vdd.n3237 gnd 1.37872f
C5263 vdd.n3238 gnd 0.023274f
C5264 vdd.n3239 gnd 0.006828f
C5265 vdd.n3240 gnd 0.023274f
C5266 vdd.n3241 gnd 0.01022f
C5267 vdd.n3242 gnd 0.01022f
C5268 vdd.n3243 gnd 0.008226f
C5269 vdd.n3244 gnd 0.01022f
C5270 vdd.n3245 gnd 0.987038f
C5271 vdd.n3246 gnd 0.01022f
C5272 vdd.n3247 gnd 0.008226f
C5273 vdd.n3248 gnd 0.01022f
C5274 vdd.n3249 gnd 0.01022f
C5275 vdd.n3250 gnd 0.01022f
C5276 vdd.n3251 gnd 0.008226f
C5277 vdd.n3252 gnd 0.01022f
C5278 vdd.n3253 gnd 1.01837f
C5279 vdd.n3254 gnd 0.01022f
C5280 vdd.n3255 gnd 0.008226f
C5281 vdd.n3256 gnd 0.01022f
C5282 vdd.n3257 gnd 0.01022f
C5283 vdd.n3258 gnd 0.01022f
C5284 vdd.n3259 gnd 0.008226f
C5285 vdd.n3260 gnd 0.01022f
C5286 vdd.t2 gnd 0.522243f
C5287 vdd.n3261 gnd 0.84081f
C5288 vdd.n3262 gnd 0.01022f
C5289 vdd.n3263 gnd 0.008226f
C5290 vdd.n3264 gnd 0.01022f
C5291 vdd.n3265 gnd 0.01022f
C5292 vdd.n3266 gnd 0.01022f
C5293 vdd.n3267 gnd 0.008226f
C5294 vdd.n3268 gnd 0.01022f
C5295 vdd.n3269 gnd 0.663248f
C5296 vdd.n3270 gnd 0.01022f
C5297 vdd.n3271 gnd 0.008226f
C5298 vdd.n3272 gnd 0.01022f
C5299 vdd.n3273 gnd 0.01022f
C5300 vdd.n3274 gnd 0.01022f
C5301 vdd.n3275 gnd 0.008226f
C5302 vdd.n3276 gnd 0.01022f
C5303 vdd.n3277 gnd 0.830366f
C5304 vdd.n3278 gnd 0.5588f
C5305 vdd.n3279 gnd 0.01022f
C5306 vdd.n3280 gnd 0.008226f
C5307 vdd.n3281 gnd 0.01022f
C5308 vdd.n3282 gnd 0.01022f
C5309 vdd.n3283 gnd 0.01022f
C5310 vdd.n3284 gnd 0.008226f
C5311 vdd.n3285 gnd 0.01022f
C5312 vdd.n3286 gnd 0.736362f
C5313 vdd.n3287 gnd 0.01022f
C5314 vdd.n3288 gnd 0.008226f
C5315 vdd.n3289 gnd 0.01022f
C5316 vdd.n3290 gnd 0.01022f
C5317 vdd.n3291 gnd 0.01022f
C5318 vdd.n3292 gnd 0.01022f
C5319 vdd.n3293 gnd 0.01022f
C5320 vdd.n3294 gnd 0.008226f
C5321 vdd.n3295 gnd 0.008226f
C5322 vdd.n3296 gnd 0.01022f
C5323 vdd.t11 gnd 0.522243f
C5324 vdd.n3297 gnd 0.866923f
C5325 vdd.n3298 gnd 0.01022f
C5326 vdd.n3299 gnd 0.008226f
C5327 vdd.n3300 gnd 0.01022f
C5328 vdd.n3301 gnd 0.01022f
C5329 vdd.n3302 gnd 0.01022f
C5330 vdd.n3303 gnd 0.008226f
C5331 vdd.n3304 gnd 0.01022f
C5332 vdd.n3305 gnd 0.819921f
C5333 vdd.n3306 gnd 0.01022f
C5334 vdd.n3307 gnd 0.01022f
C5335 vdd.n3308 gnd 0.008226f
C5336 vdd.n3309 gnd 0.008226f
C5337 vdd.n3310 gnd 0.008226f
C5338 vdd.n3311 gnd 0.01022f
C5339 vdd.n3312 gnd 0.01022f
C5340 vdd.n3313 gnd 0.01022f
C5341 vdd.n3314 gnd 0.01022f
C5342 vdd.n3315 gnd 0.008226f
C5343 vdd.n3316 gnd 0.008226f
C5344 vdd.n3317 gnd 0.008226f
C5345 vdd.n3318 gnd 0.01022f
C5346 vdd.n3319 gnd 0.01022f
C5347 vdd.n3320 gnd 0.01022f
C5348 vdd.n3321 gnd 0.01022f
C5349 vdd.n3322 gnd 0.008226f
C5350 vdd.n3323 gnd 0.008226f
C5351 vdd.n3324 gnd 0.008226f
C5352 vdd.n3325 gnd 0.01022f
C5353 vdd.n3326 gnd 0.01022f
C5354 vdd.n3327 gnd 0.01022f
C5355 vdd.n3328 gnd 0.866923f
C5356 vdd.n3329 gnd 0.01022f
C5357 vdd.n3330 gnd 0.008226f
C5358 vdd.n3331 gnd 0.008226f
C5359 vdd.n3332 gnd 0.008226f
C5360 vdd.n3333 gnd 0.01022f
C5361 vdd.n3334 gnd 0.01022f
C5362 vdd.n3335 gnd 0.01022f
C5363 vdd.n3336 gnd 0.01022f
C5364 vdd.n3337 gnd 0.008226f
C5365 vdd.n3338 gnd 0.008226f
C5366 vdd.n3339 gnd 0.006828f
C5367 vdd.n3340 gnd 0.023274f
C5368 vdd.n3341 gnd 0.023433f
C5369 vdd.n3342 gnd 0.003907f
C5370 vdd.n3343 gnd 0.023433f
C5371 vdd.n3345 gnd 2.30831f
C5372 vdd.n3346 gnd 1.37872f
C5373 vdd.n3347 gnd 0.684138f
C5374 vdd.n3348 gnd 0.01022f
C5375 vdd.n3349 gnd 0.008226f
C5376 vdd.n3350 gnd 0.008226f
C5377 vdd.n3351 gnd 0.008226f
C5378 vdd.n3352 gnd 0.01022f
C5379 vdd.n3353 gnd 1.04449f
C5380 vdd.n3354 gnd 1.04449f
C5381 vdd.n3355 gnd 0.600579f
C5382 vdd.n3356 gnd 0.01022f
C5383 vdd.n3357 gnd 0.008226f
C5384 vdd.n3358 gnd 0.008226f
C5385 vdd.n3359 gnd 0.008226f
C5386 vdd.n3360 gnd 0.01022f
C5387 vdd.n3361 gnd 0.621469f
C5388 vdd.n3362 gnd 0.767697f
C5389 vdd.t126 gnd 0.522243f
C5390 vdd.n3363 gnd 0.799031f
C5391 vdd.n3364 gnd 0.01022f
C5392 vdd.n3365 gnd 0.008226f
C5393 vdd.n3366 gnd 0.008226f
C5394 vdd.n3367 gnd 0.008226f
C5395 vdd.n3368 gnd 0.01022f
C5396 vdd.n3369 gnd 0.866923f
C5397 vdd.t105 gnd 0.522243f
C5398 vdd.n3370 gnd 0.631914f
C5399 vdd.n3371 gnd 0.757252f
C5400 vdd.n3372 gnd 0.01022f
C5401 vdd.n3373 gnd 0.008226f
C5402 vdd.n3374 gnd 0.008226f
C5403 vdd.n3375 gnd 0.008226f
C5404 vdd.n3376 gnd 0.01022f
C5405 vdd.n3377 gnd 0.579689f
C5406 vdd.t98 gnd 0.522243f
C5407 vdd.n3378 gnd 0.866923f
C5408 vdd.t140 gnd 0.522243f
C5409 vdd.n3379 gnd 0.642358f
C5410 vdd.n3380 gnd 0.01022f
C5411 vdd.n3381 gnd 0.008226f
C5412 vdd.n3382 gnd 0.007855f
C5413 vdd.n3383 gnd 0.602843f
C5414 vdd.n3384 gnd 2.55694f
C5415 a_n2140_13878.t16 gnd 0.186868f
C5416 a_n2140_13878.t15 gnd 0.186868f
C5417 a_n2140_13878.t10 gnd 0.186868f
C5418 a_n2140_13878.n0 gnd 1.47299f
C5419 a_n2140_13878.t7 gnd 0.186868f
C5420 a_n2140_13878.t9 gnd 0.186868f
C5421 a_n2140_13878.n1 gnd 1.47143f
C5422 a_n2140_13878.n2 gnd 2.05603f
C5423 a_n2140_13878.t17 gnd 0.186868f
C5424 a_n2140_13878.t8 gnd 0.186868f
C5425 a_n2140_13878.n3 gnd 1.47143f
C5426 a_n2140_13878.n4 gnd 1.00289f
C5427 a_n2140_13878.t14 gnd 0.186868f
C5428 a_n2140_13878.t6 gnd 0.186868f
C5429 a_n2140_13878.n5 gnd 1.47143f
C5430 a_n2140_13878.n6 gnd 4.06212f
C5431 a_n2140_13878.t2 gnd 1.74974f
C5432 a_n2140_13878.t21 gnd 0.186868f
C5433 a_n2140_13878.t22 gnd 0.186868f
C5434 a_n2140_13878.n7 gnd 1.3163f
C5435 a_n2140_13878.n8 gnd 1.47077f
C5436 a_n2140_13878.t23 gnd 1.74626f
C5437 a_n2140_13878.n9 gnd 0.740113f
C5438 a_n2140_13878.t3 gnd 1.74626f
C5439 a_n2140_13878.n10 gnd 0.740113f
C5440 a_n2140_13878.t0 gnd 0.186868f
C5441 a_n2140_13878.t4 gnd 0.186868f
C5442 a_n2140_13878.n11 gnd 1.3163f
C5443 a_n2140_13878.n12 gnd 0.74728f
C5444 a_n2140_13878.t1 gnd 1.74626f
C5445 a_n2140_13878.n13 gnd 2.09583f
C5446 a_n2140_13878.n14 gnd 2.85974f
C5447 a_n2140_13878.t11 gnd 0.186868f
C5448 a_n2140_13878.t12 gnd 0.186868f
C5449 a_n2140_13878.n15 gnd 1.47142f
C5450 a_n2140_13878.n16 gnd 2.01665f
C5451 a_n2140_13878.t18 gnd 0.186868f
C5452 a_n2140_13878.t19 gnd 0.186868f
C5453 a_n2140_13878.n17 gnd 1.47143f
C5454 a_n2140_13878.n18 gnd 0.651951f
C5455 a_n2140_13878.t5 gnd 0.186868f
C5456 a_n2140_13878.t13 gnd 0.186868f
C5457 a_n2140_13878.n19 gnd 1.47143f
C5458 a_n2140_13878.n20 gnd 1.32263f
C5459 a_n2140_13878.n21 gnd 1.47386f
C5460 a_n2140_13878.t20 gnd 0.186868f
C5461 a_n2318_13878.n0 gnd 2.73227f
C5462 a_n2318_13878.n1 gnd 3.94723f
C5463 a_n2318_13878.n2 gnd 3.81658f
C5464 a_n2318_13878.n3 gnd 0.652811f
C5465 a_n2318_13878.n4 gnd 0.210856f
C5466 a_n2318_13878.n5 gnd 0.210856f
C5467 a_n2318_13878.n6 gnd 0.729399f
C5468 a_n2318_13878.n7 gnd 0.210856f
C5469 a_n2318_13878.n8 gnd 0.433021f
C5470 a_n2318_13878.n9 gnd 0.652788f
C5471 a_n2318_13878.n10 gnd 0.200068f
C5472 a_n2318_13878.n11 gnd 0.147354f
C5473 a_n2318_13878.n12 gnd 0.231593f
C5474 a_n2318_13878.n13 gnd 0.178879f
C5475 a_n2318_13878.n14 gnd 0.200068f
C5476 a_n2318_13878.n15 gnd 1.09189f
C5477 a_n2318_13878.n16 gnd 0.147354f
C5478 a_n2318_13878.n17 gnd 0.705502f
C5479 a_n2318_13878.n18 gnd 0.50033f
C5480 a_n2318_13878.n19 gnd 0.210856f
C5481 a_n2318_13878.n20 gnd 0.210856f
C5482 a_n2318_13878.n21 gnd 0.433358f
C5483 a_n2318_13878.n22 gnd 0.210856f
C5484 a_n2318_13878.n23 gnd 0.210856f
C5485 a_n2318_13878.n24 gnd 1.73596f
C5486 a_n2318_13878.n25 gnd 2.03016f
C5487 a_n2318_13878.n26 gnd 1.73596f
C5488 a_n2318_13878.n27 gnd 1.85287f
C5489 a_n2318_13878.n28 gnd 3.14412f
C5490 a_n2318_13878.n29 gnd 0.278541f
C5491 a_n2318_13878.n30 gnd 0.742063f
C5492 a_n2318_13878.n31 gnd 0.004739f
C5493 a_n2318_13878.n32 gnd 0.01025f
C5494 a_n2318_13878.n33 gnd 0.01025f
C5495 a_n2318_13878.n34 gnd 0.004739f
C5496 a_n2318_13878.n35 gnd 0.278541f
C5497 a_n2318_13878.n36 gnd 0.278541f
C5498 a_n2318_13878.n37 gnd 0.433358f
C5499 a_n2318_13878.n38 gnd 0.004739f
C5500 a_n2318_13878.n39 gnd 0.01025f
C5501 a_n2318_13878.n40 gnd 0.01025f
C5502 a_n2318_13878.n41 gnd 0.004739f
C5503 a_n2318_13878.n42 gnd 0.278541f
C5504 a_n2318_13878.n43 gnd 0.008164f
C5505 a_n2318_13878.n44 gnd 0.278541f
C5506 a_n2318_13878.n45 gnd 0.008164f
C5507 a_n2318_13878.n46 gnd 0.278541f
C5508 a_n2318_13878.n47 gnd 0.008164f
C5509 a_n2318_13878.n48 gnd 0.278541f
C5510 a_n2318_13878.n49 gnd 0.008164f
C5511 a_n2318_13878.n50 gnd 0.278541f
C5512 a_n2318_13878.n51 gnd 0.278541f
C5513 a_n2318_13878.n52 gnd 0.004739f
C5514 a_n2318_13878.n53 gnd 0.01025f
C5515 a_n2318_13878.n54 gnd 0.01025f
C5516 a_n2318_13878.n55 gnd 0.004739f
C5517 a_n2318_13878.n56 gnd 0.278541f
C5518 a_n2318_13878.n57 gnd 0.278541f
C5519 a_n2318_13878.n58 gnd 0.004739f
C5520 a_n2318_13878.n59 gnd 0.01025f
C5521 a_n2318_13878.n60 gnd 0.105428f
C5522 a_n2318_13878.n61 gnd 0.01025f
C5523 a_n2318_13878.n62 gnd 0.004739f
C5524 a_n2318_13878.n63 gnd 0.278541f
C5525 a_n2318_13878.t5 gnd 0.146252f
C5526 a_n2318_13878.t6 gnd 0.691694f
C5527 a_n2318_13878.t0 gnd 0.680295f
C5528 a_n2318_13878.t4 gnd 0.680295f
C5529 a_n2318_13878.n64 gnd 0.297177f
C5530 a_n2318_13878.t28 gnd 0.680295f
C5531 a_n2318_13878.t2 gnd 0.680295f
C5532 a_n2318_13878.t26 gnd 0.680295f
C5533 a_n2318_13878.n65 gnd 0.297177f
C5534 a_n2318_13878.t22 gnd 0.680295f
C5535 a_n2318_13878.t14 gnd 0.691694f
C5536 a_n2318_13878.t41 gnd 0.113752f
C5537 a_n2318_13878.t43 gnd 0.113752f
C5538 a_n2318_13878.n66 gnd 1.00811f
C5539 a_n2318_13878.t44 gnd 0.113752f
C5540 a_n2318_13878.t46 gnd 0.113752f
C5541 a_n2318_13878.n67 gnd 1.00515f
C5542 a_n2318_13878.t40 gnd 0.113752f
C5543 a_n2318_13878.t37 gnd 0.113752f
C5544 a_n2318_13878.n68 gnd 1.00811f
C5545 a_n2318_13878.t33 gnd 0.113752f
C5546 a_n2318_13878.t32 gnd 0.113752f
C5547 a_n2318_13878.n69 gnd 1.00515f
C5548 a_n2318_13878.t39 gnd 0.113752f
C5549 a_n2318_13878.t42 gnd 0.113752f
C5550 a_n2318_13878.n70 gnd 1.00515f
C5551 a_n2318_13878.t45 gnd 0.113752f
C5552 a_n2318_13878.t47 gnd 0.113752f
C5553 a_n2318_13878.n71 gnd 1.00515f
C5554 a_n2318_13878.t38 gnd 0.113752f
C5555 a_n2318_13878.t34 gnd 0.113752f
C5556 a_n2318_13878.n72 gnd 1.00811f
C5557 a_n2318_13878.t35 gnd 0.113752f
C5558 a_n2318_13878.t36 gnd 0.113752f
C5559 a_n2318_13878.n73 gnd 1.00515f
C5560 a_n2318_13878.t78 gnd 0.691694f
C5561 a_n2318_13878.t59 gnd 0.680295f
C5562 a_n2318_13878.t63 gnd 0.680295f
C5563 a_n2318_13878.n74 gnd 0.297177f
C5564 a_n2318_13878.t53 gnd 0.680295f
C5565 a_n2318_13878.t68 gnd 0.680295f
C5566 a_n2318_13878.t75 gnd 0.680295f
C5567 a_n2318_13878.n75 gnd 0.297177f
C5568 a_n2318_13878.t76 gnd 0.680295f
C5569 a_n2318_13878.t50 gnd 0.691694f
C5570 a_n2318_13878.t17 gnd 1.36943f
C5571 a_n2318_13878.t25 gnd 0.146252f
C5572 a_n2318_13878.t9 gnd 0.146252f
C5573 a_n2318_13878.n76 gnd 1.0302f
C5574 a_n2318_13878.t13 gnd 0.146252f
C5575 a_n2318_13878.t31 gnd 0.146252f
C5576 a_n2318_13878.n77 gnd 1.0302f
C5577 a_n2318_13878.t11 gnd 0.146252f
C5578 a_n2318_13878.t21 gnd 0.146252f
C5579 a_n2318_13878.n78 gnd 1.0302f
C5580 a_n2318_13878.t19 gnd 1.3667f
C5581 a_n2318_13878.t10 gnd 0.680295f
C5582 a_n2318_13878.n79 gnd 0.297177f
C5583 a_n2318_13878.t12 gnd 0.680295f
C5584 a_n2318_13878.t16 gnd 0.691694f
C5585 a_n2318_13878.t24 gnd 0.680295f
C5586 a_n2318_13878.t57 gnd 0.680295f
C5587 a_n2318_13878.n80 gnd 0.297177f
C5588 a_n2318_13878.t71 gnd 0.680295f
C5589 a_n2318_13878.t74 gnd 0.691694f
C5590 a_n2318_13878.t52 gnd 0.680295f
C5591 a_n2318_13878.n81 gnd 0.2996f
C5592 a_n2318_13878.t72 gnd 0.680295f
C5593 a_n2318_13878.n82 gnd 0.297177f
C5594 a_n2318_13878.n83 gnd 0.292702f
C5595 a_n2318_13878.t49 gnd 0.680295f
C5596 a_n2318_13878.n84 gnd 0.292702f
C5597 a_n2318_13878.t66 gnd 0.680295f
C5598 a_n2318_13878.n85 gnd 0.2996f
C5599 a_n2318_13878.t51 gnd 0.691694f
C5600 a_n2318_13878.n86 gnd 0.2996f
C5601 a_n2318_13878.t8 gnd 0.680295f
C5602 a_n2318_13878.n87 gnd 0.297177f
C5603 a_n2318_13878.n88 gnd 0.292702f
C5604 a_n2318_13878.t30 gnd 0.680295f
C5605 a_n2318_13878.n89 gnd 0.292702f
C5606 a_n2318_13878.t20 gnd 0.680295f
C5607 a_n2318_13878.n90 gnd 0.2996f
C5608 a_n2318_13878.t18 gnd 0.691694f
C5609 a_n2318_13878.n91 gnd 1.17031f
C5610 a_n2318_13878.t56 gnd 0.680295f
C5611 a_n2318_13878.n92 gnd 0.295302f
C5612 a_n2318_13878.t62 gnd 0.680295f
C5613 a_n2318_13878.n93 gnd 0.295302f
C5614 a_n2318_13878.t55 gnd 0.680295f
C5615 a_n2318_13878.n94 gnd 0.295302f
C5616 a_n2318_13878.t67 gnd 0.680295f
C5617 a_n2318_13878.n95 gnd 0.295302f
C5618 a_n2318_13878.t58 gnd 0.680295f
C5619 a_n2318_13878.n96 gnd 0.28994f
C5620 a_n2318_13878.t79 gnd 0.680295f
C5621 a_n2318_13878.n97 gnd 0.299101f
C5622 a_n2318_13878.t60 gnd 0.691694f
C5623 a_n2318_13878.t69 gnd 0.680295f
C5624 a_n2318_13878.n98 gnd 0.28994f
C5625 a_n2318_13878.t54 gnd 0.680295f
C5626 a_n2318_13878.n99 gnd 0.299101f
C5627 a_n2318_13878.t64 gnd 0.691694f
C5628 a_n2318_13878.t73 gnd 0.680295f
C5629 a_n2318_13878.n100 gnd 0.28994f
C5630 a_n2318_13878.t61 gnd 0.680295f
C5631 a_n2318_13878.n101 gnd 0.299101f
C5632 a_n2318_13878.t77 gnd 0.691694f
C5633 a_n2318_13878.t65 gnd 0.680295f
C5634 a_n2318_13878.n102 gnd 0.28994f
C5635 a_n2318_13878.t48 gnd 0.680295f
C5636 a_n2318_13878.n103 gnd 0.299101f
C5637 a_n2318_13878.t70 gnd 0.691694f
C5638 a_n2318_13878.n104 gnd 1.41607f
C5639 a_n2318_13878.n105 gnd 0.2996f
C5640 a_n2318_13878.n106 gnd 0.292702f
C5641 a_n2318_13878.n107 gnd 0.292702f
C5642 a_n2318_13878.n108 gnd 0.2996f
C5643 a_n2318_13878.n109 gnd 0.2996f
C5644 a_n2318_13878.n110 gnd 0.292702f
C5645 a_n2318_13878.n111 gnd 0.292702f
C5646 a_n2318_13878.n112 gnd 0.2996f
C5647 a_n2318_13878.n113 gnd 0.839379f
C5648 a_n2318_13878.t7 gnd 1.36671f
C5649 a_n2318_13878.t15 gnd 1.36943f
C5650 a_n2318_13878.t27 gnd 0.146252f
C5651 a_n2318_13878.t23 gnd 0.146252f
C5652 a_n2318_13878.n114 gnd 1.0302f
C5653 a_n2318_13878.t29 gnd 0.146252f
C5654 a_n2318_13878.t3 gnd 0.146252f
C5655 a_n2318_13878.n115 gnd 1.0302f
C5656 a_n2318_13878.n116 gnd 1.0302f
C5657 a_n2318_13878.t1 gnd 0.146252f
.ends

