* NGSPICE file created from opamp17.ext - technology: sky130A

.subckt opamp17 gnd CSoutput output vdd plus minus commonsourceibias outputibias diffpairibias
X0 gnd.t330 commonsourceibias.t28 commonsourceibias.t29 gnd.t268 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X1 a_n2804_13878.t7 a_n2982_13878.t72 vdd.t227 vdd.t226 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X2 a_n2804_13878.t31 a_n2982_13878.t62 a_n2982_13878.t63 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 vdd.t144 a_n8300_8799.t48 CSoutput.t71 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X4 commonsourceibias.t27 commonsourceibias.t26 gnd.t329 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X5 CSoutput.t70 a_n8300_8799.t49 vdd.t145 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X6 a_n3827_n3924.t50 diffpairibias.t20 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X7 gnd.t328 commonsourceibias.t24 commonsourceibias.t25 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 a_n2982_8322.t37 a_n2982_13878.t73 a_n8300_8799.t26 vdd.t224 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X9 commonsourceibias.t23 commonsourceibias.t22 gnd.t327 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X10 gnd.t326 commonsourceibias.t48 CSoutput.t143 gnd.t263 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X11 gnd.t150 gnd.t148 gnd.t149 gnd.t73 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X12 gnd.t153 gnd.t151 gnd.t152 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X13 gnd.t147 gnd.t146 plus.t4 gnd.t73 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X14 CSoutput.t69 a_n8300_8799.t50 vdd.t237 vdd.t112 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X15 a_n8300_8799.t2 plus.t5 a_n3827_n3924.t3 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X16 minus.t4 gnd.t143 gnd.t145 gnd.t144 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X17 vdd.t238 a_n8300_8799.t51 CSoutput.t68 vdd.t4 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X18 gnd.t142 gnd.t140 gnd.t141 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X19 output.t19 outputibias.t8 gnd.t181 gnd.t180 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X20 a_n8300_8799.t29 a_n2982_13878.t74 a_n2982_8322.t36 vdd.t210 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X21 vdd.t230 a_n8300_8799.t52 CSoutput.t67 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X22 vdd.t231 a_n8300_8799.t53 CSoutput.t66 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X23 commonsourceibias.t21 commonsourceibias.t20 gnd.t325 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X24 a_n8300_8799.t21 a_n2982_13878.t75 a_n2982_8322.t35 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X25 gnd.t139 gnd.t136 gnd.t138 gnd.t137 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X26 gnd.t135 gnd.t132 gnd.t134 gnd.t133 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X27 a_n8300_8799.t10 plus.t6 a_n3827_n3924.t22 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X28 gnd.t324 commonsourceibias.t49 CSoutput.t142 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X29 CSoutput.t141 commonsourceibias.t50 gnd.t323 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X30 gnd.t322 commonsourceibias.t18 commonsourceibias.t19 gnd.t263 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X31 a_n3827_n3924.t49 diffpairibias.t21 gnd.t197 gnd.t196 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X32 a_n3827_n3924.t9 minus.t5 a_n2982_13878.t4 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X33 commonsourceibias.t17 commonsourceibias.t16 gnd.t321 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X34 CSoutput.t65 a_n8300_8799.t54 vdd.t135 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X35 a_n3827_n3924.t5 plus.t7 a_n8300_8799.t4 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X36 vdd.t136 a_n8300_8799.t55 CSoutput.t64 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X37 a_n2982_13878.t5 minus.t6 a_n3827_n3924.t12 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X38 a_n3827_n3924.t0 plus.t8 a_n8300_8799.t0 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X39 a_n3827_n3924.t38 minus.t7 a_n2982_13878.t20 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X40 gnd.t320 commonsourceibias.t14 commonsourceibias.t15 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X41 CSoutput.t140 commonsourceibias.t51 gnd.t319 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X42 a_n2804_13878.t30 a_n2982_13878.t58 a_n2982_13878.t59 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X43 a_n2982_13878.t23 a_n2982_13878.t22 a_n2804_13878.t29 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X44 output.t18 outputibias.t9 gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X45 CSoutput.t63 a_n8300_8799.t56 vdd.t113 vdd.t112 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X46 a_n3827_n3924.t8 minus.t8 a_n2982_13878.t3 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X47 vdd.t85 vdd.t83 vdd.t84 vdd.t60 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X48 vdd.t114 a_n8300_8799.t57 CSoutput.t62 vdd.t4 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X49 diffpairibias.t19 diffpairibias.t18 gnd.t191 gnd.t190 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X50 a_n2982_13878.t29 a_n2982_13878.t28 a_n2804_13878.t28 vdd.t209 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X51 CSoutput.t139 commonsourceibias.t52 gnd.t318 gnd.t279 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 CSoutput.t138 commonsourceibias.t53 gnd.t317 gnd.t252 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X53 a_n8300_8799.t35 a_n2982_13878.t76 a_n2982_8322.t34 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X54 CSoutput.t61 a_n8300_8799.t58 vdd.t120 vdd.t119 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X55 a_n2982_13878.t18 minus.t9 a_n3827_n3924.t36 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X56 a_n2982_13878.t31 a_n2982_13878.t30 a_n2804_13878.t27 vdd.t225 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X57 gnd.t131 gnd.t129 gnd.t130 gnd.t50 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X58 gnd.t128 gnd.t126 plus.t3 gnd.t127 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X59 vdd.t122 a_n8300_8799.t59 CSoutput.t60 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X60 vdd.t129 a_n8300_8799.t60 CSoutput.t59 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X61 a_n8300_8799.t25 a_n2982_13878.t77 a_n2982_8322.t33 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X62 diffpairibias.t17 diffpairibias.t16 gnd.t332 gnd.t331 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X63 CSoutput.t58 a_n8300_8799.t61 vdd.t131 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X64 gnd.t125 gnd.t123 gnd.t124 gnd.t50 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X65 a_n8300_8799.t22 a_n2982_13878.t78 a_n2982_8322.t32 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X66 CSoutput.t144 a_n2982_8322.t5 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X67 a_n2982_8322.t31 a_n2982_13878.t79 a_n8300_8799.t34 vdd.t225 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X68 CSoutput.t137 commonsourceibias.t54 gnd.t316 gnd.t252 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X69 vdd.t82 vdd.t80 vdd.t81 vdd.t47 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X70 CSoutput.t57 a_n8300_8799.t62 vdd.t87 vdd.t86 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X71 plus.t2 gnd.t120 gnd.t122 gnd.t121 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X72 output.t15 CSoutput.t145 vdd.t163 gnd.t186 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X73 gnd.t315 commonsourceibias.t55 CSoutput.t136 gnd.t241 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X74 CSoutput.t146 a_n2982_8322.t4 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X75 CSoutput.t135 commonsourceibias.t56 gnd.t314 gnd.t254 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X76 a_n8300_8799.t17 plus.t9 a_n3827_n3924.t33 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X77 gnd.t313 commonsourceibias.t57 CSoutput.t134 gnd.t229 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X78 gnd.t119 gnd.t117 gnd.t118 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X79 a_n3827_n3924.t48 diffpairibias.t22 gnd.t203 gnd.t202 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X80 vdd.t89 a_n8300_8799.t63 CSoutput.t56 vdd.t88 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X81 a_n3827_n3924.t16 minus.t10 a_n2982_13878.t8 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X82 vdd.t95 a_n8300_8799.t64 CSoutput.t55 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X83 CSoutput.t133 commonsourceibias.t58 gnd.t312 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X84 a_n2982_13878.t57 a_n2982_13878.t56 a_n2804_13878.t26 vdd.t224 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X85 vdd.t97 a_n8300_8799.t65 CSoutput.t54 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 a_n8300_8799.t41 a_n2982_13878.t80 a_n2982_8322.t30 vdd.t213 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X87 a_n2982_13878.t35 a_n2982_13878.t34 a_n2804_13878.t25 vdd.t176 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X88 a_n2982_13878.t7 minus.t11 a_n3827_n3924.t15 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X89 a_n3827_n3924.t17 plus.t10 a_n8300_8799.t8 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X90 outputibias.t7 outputibias.t6 gnd.t208 gnd.t207 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X91 commonsourceibias.t43 commonsourceibias.t42 gnd.t311 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X92 gnd.t310 commonsourceibias.t59 CSoutput.t132 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X93 CSoutput.t131 commonsourceibias.t60 gnd.t309 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 gnd.t116 gnd.t114 gnd.t115 gnd.t58 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X95 outputibias.t5 outputibias.t4 gnd.t165 gnd.t164 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X96 diffpairibias.t15 diffpairibias.t14 gnd.t22 gnd.t21 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X97 a_n3827_n3924.t35 minus.t12 a_n2982_13878.t17 gnd.t183 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X98 vdd.t79 vdd.t77 vdd.t78 vdd.t67 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X99 CSoutput.t53 a_n8300_8799.t66 vdd.t148 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X100 vdd.t76 vdd.t73 vdd.t75 vdd.t74 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X101 CSoutput.t52 a_n8300_8799.t67 vdd.t150 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X102 a_n2804_13878.t24 a_n2982_13878.t68 a_n2982_13878.t69 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X103 vdd.t241 a_n8300_8799.t68 CSoutput.t51 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X104 vdd.t223 a_n2982_13878.t81 a_n2982_8322.t13 vdd.t222 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X105 gnd.t308 commonsourceibias.t40 commonsourceibias.t41 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X106 a_n2982_13878.t39 a_n2982_13878.t38 a_n2804_13878.t23 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X107 vdd.t72 vdd.t70 vdd.t71 vdd.t47 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X108 output.t14 CSoutput.t147 vdd.t106 gnd.t27 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X109 CSoutput.t130 commonsourceibias.t61 gnd.t307 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X110 a_n2982_8322.t12 a_n2982_13878.t82 vdd.t221 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X111 a_n3827_n3924.t47 diffpairibias.t23 gnd.t17 gnd.t16 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X112 CSoutput.t50 a_n8300_8799.t69 vdd.t242 vdd.t86 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X113 gnd.t306 commonsourceibias.t62 CSoutput.t129 gnd.t268 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X114 a_n2982_13878.t11 minus.t13 a_n3827_n3924.t21 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X115 commonsourceibias.t39 commonsourceibias.t38 gnd.t305 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X116 a_n3827_n3924.t32 plus.t11 a_n8300_8799.t16 gnd.t187 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X117 vdd.t219 a_n2982_13878.t83 a_n2804_13878.t6 vdd.t218 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X118 gnd.t304 commonsourceibias.t63 CSoutput.t128 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X119 gnd.t113 gnd.t111 minus.t3 gnd.t112 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X120 gnd.t110 gnd.t108 gnd.t109 gnd.t58 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X121 gnd.t107 gnd.t105 gnd.t106 gnd.t36 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X122 gnd.t303 commonsourceibias.t36 commonsourceibias.t37 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X123 vdd.t69 vdd.t66 vdd.t68 vdd.t67 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X124 a_n2804_13878.t22 a_n2982_13878.t52 a_n2982_13878.t53 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X125 vdd.t232 a_n8300_8799.t70 CSoutput.t49 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X126 vdd.t233 a_n8300_8799.t71 CSoutput.t48 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X127 a_n2982_8322.t29 a_n2982_13878.t84 a_n8300_8799.t37 vdd.t203 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X128 CSoutput.t127 commonsourceibias.t64 gnd.t302 gnd.t254 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X129 a_n8300_8799.t9 plus.t12 a_n3827_n3924.t19 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X130 vdd.t65 vdd.t63 vdd.t64 vdd.t29 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X131 commonsourceibias.t33 commonsourceibias.t32 gnd.t301 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X132 vdd.t62 vdd.t59 vdd.t61 vdd.t60 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X133 a_n2982_8322.t11 a_n2982_13878.t85 vdd.t216 vdd.t215 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X134 gnd.t300 commonsourceibias.t65 CSoutput.t126 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X135 a_n2982_13878.t21 minus.t14 a_n3827_n3924.t40 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X136 a_n8300_8799.t40 a_n2982_13878.t86 a_n2982_8322.t28 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X137 CSoutput.t47 a_n8300_8799.t72 vdd.t159 vdd.t92 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X138 diffpairibias.t13 diffpairibias.t12 gnd.t173 gnd.t172 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X139 vdd.t160 a_n8300_8799.t73 CSoutput.t46 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X140 a_n2982_13878.t67 a_n2982_13878.t66 a_n2804_13878.t21 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X141 a_n8300_8799.t28 a_n2982_13878.t87 a_n2982_8322.t27 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X142 a_n2804_13878.t20 a_n2982_13878.t44 a_n2982_13878.t45 vdd.t213 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X143 a_n8300_8799.t6 plus.t13 a_n3827_n3924.t11 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X144 gnd.t299 commonsourceibias.t66 CSoutput.t125 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X145 output.t13 CSoutput.t148 vdd.t107 gnd.t28 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X146 a_n3827_n3924.t6 minus.t15 a_n2982_13878.t1 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X147 vdd.t109 CSoutput.t149 output.t12 gnd.t154 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X148 gnd.t298 commonsourceibias.t67 CSoutput.t124 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X149 a_n3827_n3924.t26 minus.t16 a_n2982_13878.t13 gnd.t30 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X150 vdd.t58 vdd.t56 vdd.t57 vdd.t15 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X151 CSoutput.t45 a_n8300_8799.t74 vdd.t164 vdd.t119 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X152 a_n2982_13878.t71 minus.t17 a_n3827_n3924.t57 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X153 vdd.t212 a_n2982_13878.t88 a_n2982_8322.t10 vdd.t211 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X154 a_n2804_13878.t19 a_n2982_13878.t46 a_n2982_13878.t47 vdd.t210 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X155 vdd.t165 a_n8300_8799.t75 CSoutput.t44 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X156 a_n2982_13878.t37 a_n2982_13878.t36 a_n2804_13878.t18 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X157 gnd.t104 gnd.t102 gnd.t103 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X158 vdd.t110 CSoutput.t150 output.t11 gnd.t155 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X159 CSoutput.t123 commonsourceibias.t68 gnd.t297 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X160 gnd.t296 commonsourceibias.t69 CSoutput.t122 gnd.t241 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X161 gnd.t295 commonsourceibias.t70 CSoutput.t121 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X162 vdd.t161 a_n8300_8799.t76 CSoutput.t43 vdd.t90 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X163 a_n3827_n3924.t46 diffpairibias.t24 gnd.t201 gnd.t200 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X164 a_n3827_n3924.t45 diffpairibias.t25 gnd.t179 gnd.t178 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X165 a_n2982_13878.t9 minus.t18 a_n3827_n3924.t18 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X166 vdd.t162 a_n8300_8799.t77 CSoutput.t42 vdd.t88 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X167 gnd.t101 gnd.t99 gnd.t100 gnd.t36 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X168 gnd.t98 gnd.t96 minus.t2 gnd.t97 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X169 vdd.t55 vdd.t53 vdd.t54 vdd.t29 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X170 a_n2804_13878.t17 a_n2982_13878.t64 a_n2982_13878.t65 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X171 a_n2982_8322.t26 a_n2982_13878.t89 a_n8300_8799.t38 vdd.t209 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X172 CSoutput.t41 a_n8300_8799.t78 vdd.t166 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X173 vdd.t111 CSoutput.t151 output.t10 gnd.t156 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X174 a_n2982_13878.t15 minus.t19 a_n3827_n3924.t31 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X175 CSoutput.t120 commonsourceibias.t71 gnd.t294 gnd.t279 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X176 output.t9 CSoutput.t152 vdd.t170 gnd.t205 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X177 gnd.t95 gnd.t93 gnd.t94 gnd.t50 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X178 gnd.t293 commonsourceibias.t72 CSoutput.t119 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X179 diffpairibias.t11 diffpairibias.t10 gnd.t7 gnd.t6 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X180 a_n2804_13878.t5 a_n2982_13878.t90 vdd.t208 vdd.t207 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X181 vdd.t206 a_n2982_13878.t91 a_n2804_13878.t4 vdd.t205 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X182 CSoutput.t40 a_n8300_8799.t79 vdd.t167 vdd.t119 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X183 gnd.t292 commonsourceibias.t73 CSoutput.t118 gnd.t263 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X184 a_n3827_n3924.t53 plus.t14 a_n8300_8799.t45 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X185 CSoutput.t117 commonsourceibias.t74 gnd.t291 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X186 vdd.t151 a_n8300_8799.t80 CSoutput.t39 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X187 output.t8 CSoutput.t153 vdd.t171 gnd.t206 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X188 vdd.t152 a_n8300_8799.t81 CSoutput.t38 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X189 CSoutput.t37 a_n8300_8799.t82 vdd.t99 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X190 a_n3827_n3924.t7 minus.t20 a_n2982_13878.t2 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X191 a_n2804_13878.t16 a_n2982_13878.t54 a_n2982_13878.t55 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X192 diffpairibias.t9 diffpairibias.t8 gnd.t24 gnd.t23 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X193 a_n3827_n3924.t54 plus.t15 a_n8300_8799.t46 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X194 gnd.t290 commonsourceibias.t75 CSoutput.t116 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X195 CSoutput.t154 a_n2982_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X196 a_n3827_n3924.t1 minus.t21 a_n2982_13878.t0 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X197 a_n8300_8799.t47 plus.t16 a_n3827_n3924.t56 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X198 gnd.t92 gnd.t90 gnd.t91 gnd.t36 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X199 vdd.t100 a_n8300_8799.t83 CSoutput.t36 vdd.t90 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X200 commonsourceibias.t31 commonsourceibias.t30 gnd.t289 gnd.t279 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X201 a_n2982_8322.t25 a_n2982_13878.t92 a_n8300_8799.t24 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X202 CSoutput.t35 a_n8300_8799.t84 vdd.t3 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X203 a_n2982_13878.t61 a_n2982_13878.t60 a_n2804_13878.t15 vdd.t203 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X204 diffpairibias.t7 diffpairibias.t6 gnd.t19 gnd.t18 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X205 vdd.t5 a_n8300_8799.t85 CSoutput.t34 vdd.t4 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X206 a_n2804_13878.t14 a_n2982_13878.t26 a_n2982_13878.t27 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X207 vdd.t52 vdd.t50 vdd.t51 vdd.t33 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X208 vdd.t201 a_n2982_13878.t93 a_n2982_8322.t9 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X209 vdd.t228 a_n8300_8799.t86 CSoutput.t33 vdd.t88 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X210 gnd.t89 gnd.t86 gnd.t88 gnd.t87 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X211 CSoutput.t115 commonsourceibias.t76 gnd.t288 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X212 CSoutput.t155 a_n2982_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X213 output.t17 outputibias.t10 gnd.t171 gnd.t170 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X214 gnd.t85 gnd.t83 gnd.t84 gnd.t58 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X215 commonsourceibias.t5 commonsourceibias.t4 gnd.t287 gnd.t252 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X216 CSoutput.t32 a_n8300_8799.t87 vdd.t229 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X217 gnd.t82 gnd.t79 gnd.t81 gnd.t80 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X218 a_n2804_13878.t3 a_n2982_13878.t94 vdd.t199 vdd.t198 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X219 vdd.t49 vdd.t46 vdd.t48 vdd.t47 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X220 vdd.t45 vdd.t43 vdd.t44 vdd.t33 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X221 vdd.t8 CSoutput.t156 output.t7 gnd.t9 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X222 CSoutput.t114 commonsourceibias.t77 gnd.t286 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X223 plus.t1 gnd.t76 gnd.t78 gnd.t77 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X224 gnd.t285 commonsourceibias.t78 CSoutput.t113 gnd.t268 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X225 output.t16 outputibias.t11 gnd.t161 gnd.t160 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X226 CSoutput.t31 a_n8300_8799.t88 vdd.t146 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X227 gnd.t284 commonsourceibias.t2 commonsourceibias.t3 gnd.t229 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X228 gnd.t75 gnd.t72 gnd.t74 gnd.t73 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X229 gnd.t283 commonsourceibias.t79 CSoutput.t112 gnd.t241 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X230 CSoutput.t111 commonsourceibias.t80 gnd.t282 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X231 gnd.t71 gnd.t69 minus.t1 gnd.t70 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X232 CSoutput.t110 commonsourceibias.t81 gnd.t281 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X233 gnd.t68 gnd.t65 gnd.t67 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X234 gnd.t64 gnd.t61 gnd.t63 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X235 CSoutput.t109 commonsourceibias.t82 gnd.t280 gnd.t279 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X236 gnd.t278 commonsourceibias.t83 CSoutput.t108 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X237 vdd.t42 vdd.t40 vdd.t41 vdd.t19 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X238 vdd.t147 a_n8300_8799.t89 CSoutput.t30 vdd.t115 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X239 a_n3827_n3924.t44 diffpairibias.t26 gnd.t189 gnd.t188 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X240 commonsourceibias.t1 commonsourceibias.t0 gnd.t277 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X241 vdd.t197 a_n2982_13878.t95 a_n2982_8322.t8 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X242 a_n2982_8322.t24 a_n2982_13878.t96 a_n8300_8799.t19 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X243 CSoutput.t107 commonsourceibias.t84 gnd.t276 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X244 gnd.t275 commonsourceibias.t85 CSoutput.t106 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X245 CSoutput.t105 commonsourceibias.t86 gnd.t274 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X246 gnd.t273 commonsourceibias.t87 CSoutput.t104 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X247 gnd.t272 commonsourceibias.t88 CSoutput.t103 gnd.t229 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X248 CSoutput.t102 commonsourceibias.t89 gnd.t271 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X249 gnd.t60 gnd.t57 gnd.t59 gnd.t58 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X250 a_n3827_n3924.t23 plus.t17 a_n8300_8799.t11 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X251 vdd.t39 vdd.t36 vdd.t38 vdd.t37 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X252 vdd.t239 a_n8300_8799.t90 CSoutput.t29 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X253 a_n8300_8799.t12 plus.t18 a_n3827_n3924.t24 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X254 CSoutput.t28 a_n8300_8799.t91 vdd.t240 vdd.t86 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X255 a_n3827_n3924.t13 minus.t22 a_n2982_13878.t6 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X256 a_n2804_13878.t13 a_n2982_13878.t48 a_n2982_13878.t49 vdd.t189 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X257 CSoutput.t27 a_n8300_8799.t92 vdd.t234 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X258 CSoutput.t101 commonsourceibias.t90 gnd.t270 gnd.t254 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X259 a_n2982_8322.t23 a_n2982_13878.t97 a_n8300_8799.t32 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X260 vdd.t35 vdd.t32 vdd.t34 vdd.t33 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X261 gnd.t269 commonsourceibias.t91 CSoutput.t100 gnd.t268 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X262 diffpairibias.t5 diffpairibias.t4 gnd.t177 gnd.t176 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X263 CSoutput.t99 commonsourceibias.t92 gnd.t267 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X264 a_n3827_n3924.t37 minus.t23 a_n2982_13878.t19 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X265 a_n8300_8799.t44 plus.t19 a_n3827_n3924.t52 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X266 output.t6 CSoutput.t157 vdd.t9 gnd.t10 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X267 CSoutput.t26 a_n8300_8799.t93 vdd.t235 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X268 gnd.t265 commonsourceibias.t93 CSoutput.t98 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X269 CSoutput.t25 a_n8300_8799.t94 vdd.t137 vdd.t92 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X270 a_n3827_n3924.t43 diffpairibias.t27 gnd.t163 gnd.t162 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X271 vdd.t31 vdd.t28 vdd.t30 vdd.t29 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X272 gnd.t264 commonsourceibias.t94 CSoutput.t97 gnd.t263 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X273 a_n2982_8322.t7 a_n2982_13878.t98 vdd.t193 vdd.t192 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X274 gnd.t262 commonsourceibias.t95 CSoutput.t96 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X275 CSoutput.t95 commonsourceibias.t96 gnd.t261 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X276 CSoutput.t24 a_n8300_8799.t95 vdd.t138 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X277 outputibias.t3 outputibias.t2 gnd.t195 gnd.t194 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X278 gnd.t260 commonsourceibias.t6 commonsourceibias.t7 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X279 a_n3827_n3924.t10 plus.t20 a_n8300_8799.t5 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X280 vdd.t116 a_n8300_8799.t96 CSoutput.t23 vdd.t115 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X281 CSoutput.t22 a_n8300_8799.t97 vdd.t118 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X282 vdd.t191 a_n2982_13878.t99 a_n2804_13878.t2 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X283 vdd.t123 a_n8300_8799.t98 CSoutput.t21 vdd.t115 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X284 CSoutput.t20 a_n8300_8799.t99 vdd.t124 vdd.t112 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X285 gnd.t259 commonsourceibias.t97 CSoutput.t94 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X286 CSoutput.t93 commonsourceibias.t98 gnd.t257 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X287 CSoutput.t92 commonsourceibias.t99 gnd.t253 gnd.t252 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X288 gnd.t256 commonsourceibias.t100 CSoutput.t91 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X289 commonsourceibias.t13 commonsourceibias.t12 gnd.t255 gnd.t254 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X290 gnd.t251 commonsourceibias.t101 CSoutput.t90 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X291 a_n8300_8799.t1 plus.t21 a_n3827_n3924.t2 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X292 gnd.t250 commonsourceibias.t10 commonsourceibias.t11 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X293 a_n3827_n3924.t34 minus.t24 a_n2982_13878.t16 gnd.t187 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X294 a_n2982_8322.t22 a_n2982_13878.t100 a_n8300_8799.t31 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X295 a_n8300_8799.t36 a_n2982_13878.t101 a_n2982_8322.t21 vdd.t189 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X296 gnd.t249 commonsourceibias.t102 CSoutput.t89 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X297 a_n2804_13878.t1 a_n2982_13878.t102 vdd.t188 vdd.t187 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X298 CSoutput.t88 commonsourceibias.t103 gnd.t247 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X299 vdd.t27 vdd.t25 vdd.t26 vdd.t11 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X300 vdd.t132 a_n8300_8799.t100 CSoutput.t19 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X301 CSoutput.t18 a_n8300_8799.t101 vdd.t133 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X302 vdd.t125 CSoutput.t158 output.t5 gnd.t166 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X303 a_n2982_13878.t41 a_n2982_13878.t40 a_n2804_13878.t12 vdd.t177 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X304 gnd.t246 commonsourceibias.t8 commonsourceibias.t9 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X305 a_n8300_8799.t39 a_n2982_13878.t103 a_n2982_8322.t20 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X306 a_n8300_8799.t3 plus.t22 a_n3827_n3924.t4 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X307 CSoutput.t87 commonsourceibias.t104 gnd.t245 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X308 a_n8300_8799.t30 a_n2982_13878.t104 a_n2982_8322.t19 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X309 a_n2982_8322.t18 a_n2982_13878.t105 a_n8300_8799.t23 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X310 a_n2982_13878.t14 minus.t25 a_n3827_n3924.t28 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X311 vdd.t91 a_n8300_8799.t102 CSoutput.t17 vdd.t90 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X312 CSoutput.t16 a_n8300_8799.t103 vdd.t93 vdd.t92 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X313 CSoutput.t86 commonsourceibias.t105 gnd.t243 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X314 gnd.t244 commonsourceibias.t106 CSoutput.t85 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X315 CSoutput.t15 a_n8300_8799.t104 vdd.t102 vdd.t101 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X316 CSoutput.t14 a_n8300_8799.t105 vdd.t103 vdd.t101 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X317 a_n2804_13878.t11 a_n2982_13878.t50 a_n2982_13878.t51 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X318 vdd.t139 a_n8300_8799.t106 CSoutput.t13 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X319 gnd.t242 commonsourceibias.t46 commonsourceibias.t47 gnd.t241 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X320 gnd.t240 commonsourceibias.t44 commonsourceibias.t45 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X321 a_n3827_n3924.t14 plus.t23 a_n8300_8799.t7 gnd.t30 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X322 a_n8300_8799.t14 plus.t24 a_n3827_n3924.t29 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X323 a_n3827_n3924.t42 diffpairibias.t28 gnd.t193 gnd.t192 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X324 vdd.t141 a_n8300_8799.t107 CSoutput.t12 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X325 CSoutput.t84 commonsourceibias.t107 gnd.t238 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X326 gnd.t236 commonsourceibias.t108 CSoutput.t83 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X327 CSoutput.t11 a_n8300_8799.t108 vdd.t154 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X328 a_n2982_13878.t33 a_n2982_13878.t32 a_n2804_13878.t10 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X329 output.t4 CSoutput.t159 vdd.t126 gnd.t167 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X330 a_n8300_8799.t27 a_n2982_13878.t106 a_n2982_8322.t17 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X331 vdd.t155 a_n8300_8799.t109 CSoutput.t10 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X332 CSoutput.t9 a_n8300_8799.t110 vdd.t243 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X333 a_n3827_n3924.t27 plus.t25 a_n8300_8799.t13 gnd.t183 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X334 vdd.t24 vdd.t22 vdd.t23 vdd.t19 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X335 gnd.t56 gnd.t53 gnd.t55 gnd.t54 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X336 gnd.t234 commonsourceibias.t109 CSoutput.t82 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X337 gnd.t45 gnd.t42 gnd.t44 gnd.t43 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X338 diffpairibias.t3 diffpairibias.t2 gnd.t159 gnd.t158 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X339 CSoutput.t8 a_n8300_8799.t111 vdd.t236 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X340 CSoutput.t81 commonsourceibias.t110 gnd.t232 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X341 output.t3 CSoutput.t160 vdd.t127 gnd.t168 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X342 a_n2982_8322.t16 a_n2982_13878.t107 a_n8300_8799.t33 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X343 vdd.t142 CSoutput.t161 output.t2 gnd.t175 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X344 gnd.t230 commonsourceibias.t111 CSoutput.t80 gnd.t229 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X345 vdd.t168 a_n8300_8799.t112 CSoutput.t7 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X346 gnd.t52 gnd.t49 gnd.t51 gnd.t50 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X347 CSoutput.t162 a_n2982_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X348 CSoutput.t6 a_n8300_8799.t113 vdd.t156 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X349 diffpairibias.t1 diffpairibias.t0 gnd.t210 gnd.t209 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X350 gnd.t48 gnd.t46 plus.t0 gnd.t47 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X351 a_n8300_8799.t18 plus.t26 a_n3827_n3924.t39 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X352 CSoutput.t79 commonsourceibias.t112 gnd.t228 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X353 outputibias.t1 outputibias.t0 gnd.t334 gnd.t333 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X354 minus.t0 gnd.t39 gnd.t41 gnd.t40 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X355 CSoutput.t163 a_n2982_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X356 vdd.t179 a_n2982_13878.t108 a_n2804_13878.t0 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X357 CSoutput.t5 a_n8300_8799.t114 vdd.t108 vdd.t101 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X358 gnd.t226 commonsourceibias.t113 CSoutput.t78 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X359 vdd.t1 a_n8300_8799.t115 CSoutput.t4 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X360 gnd.t38 gnd.t35 gnd.t37 gnd.t36 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X361 a_n2982_8322.t15 a_n2982_13878.t109 a_n8300_8799.t42 vdd.t177 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X362 a_n2982_13878.t10 minus.t26 a_n3827_n3924.t20 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X363 vdd.t104 CSoutput.t164 output.t1 gnd.t25 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X364 a_n2982_8322.t14 a_n2982_13878.t110 a_n8300_8799.t20 vdd.t176 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X365 CSoutput.t77 commonsourceibias.t114 gnd.t224 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X366 vdd.t157 a_n8300_8799.t116 CSoutput.t3 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X367 vdd.t7 a_n8300_8799.t117 CSoutput.t2 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X368 CSoutput.t1 a_n8300_8799.t118 vdd.t158 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X369 gnd.t222 commonsourceibias.t115 CSoutput.t76 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X370 commonsourceibias.t35 commonsourceibias.t34 gnd.t220 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X371 CSoutput.t75 commonsourceibias.t116 gnd.t218 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X372 a_n3827_n3924.t51 plus.t27 a_n8300_8799.t43 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X373 vdd.t21 vdd.t18 vdd.t20 vdd.t19 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X374 a_n2982_8322.t6 a_n2982_13878.t111 vdd.t175 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X375 a_n2982_13878.t12 minus.t27 a_n3827_n3924.t25 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X376 a_n2804_13878.t9 a_n2982_13878.t42 a_n2982_13878.t43 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X377 vdd.t105 CSoutput.t165 output.t0 gnd.t26 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X378 vdd.t17 vdd.t14 vdd.t16 vdd.t15 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X379 a_n3827_n3924.t41 diffpairibias.t29 gnd.t199 gnd.t198 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X380 a_n2982_13878.t70 minus.t28 a_n3827_n3924.t55 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X381 vdd.t13 vdd.t10 vdd.t12 vdd.t11 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X382 CSoutput.t0 a_n8300_8799.t119 vdd.t169 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X383 CSoutput.t74 commonsourceibias.t117 gnd.t214 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X384 CSoutput.t73 commonsourceibias.t118 gnd.t216 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X385 a_n3827_n3924.t30 plus.t28 a_n8300_8799.t15 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X386 gnd.t212 commonsourceibias.t119 CSoutput.t72 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X387 a_n2982_13878.t25 a_n2982_13878.t24 a_n2804_13878.t8 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 commonsourceibias.n25 commonsourceibias.t16 230.006
R1 commonsourceibias.n91 commonsourceibias.t96 230.006
R2 commonsourceibias.n218 commonsourceibias.t118 230.006
R3 commonsourceibias.n154 commonsourceibias.t98 230.006
R4 commonsourceibias.n322 commonsourceibias.t46 230.006
R5 commonsourceibias.n281 commonsourceibias.t69 230.006
R6 commonsourceibias.n483 commonsourceibias.t55 230.006
R7 commonsourceibias.n419 commonsourceibias.t79 230.006
R8 commonsourceibias.n70 commonsourceibias.t2 207.983
R9 commonsourceibias.n136 commonsourceibias.t57 207.983
R10 commonsourceibias.n263 commonsourceibias.t111 207.983
R11 commonsourceibias.n199 commonsourceibias.t88 207.983
R12 commonsourceibias.n368 commonsourceibias.t38 207.983
R13 commonsourceibias.n402 commonsourceibias.t114 207.983
R14 commonsourceibias.n529 commonsourceibias.t51 207.983
R15 commonsourceibias.n465 commonsourceibias.t74 207.983
R16 commonsourceibias.n10 commonsourceibias.t42 168.701
R17 commonsourceibias.n63 commonsourceibias.t44 168.701
R18 commonsourceibias.n57 commonsourceibias.t32 168.701
R19 commonsourceibias.n16 commonsourceibias.t24 168.701
R20 commonsourceibias.n49 commonsourceibias.t4 168.701
R21 commonsourceibias.n43 commonsourceibias.t14 168.701
R22 commonsourceibias.n19 commonsourceibias.t22 168.701
R23 commonsourceibias.n21 commonsourceibias.t36 168.701
R24 commonsourceibias.n23 commonsourceibias.t26 168.701
R25 commonsourceibias.n26 commonsourceibias.t8 168.701
R26 commonsourceibias.n1 commonsourceibias.t110 168.701
R27 commonsourceibias.n129 commonsourceibias.t70 168.701
R28 commonsourceibias.n123 commonsourceibias.t117 168.701
R29 commonsourceibias.n7 commonsourceibias.t85 168.701
R30 commonsourceibias.n115 commonsourceibias.t54 168.701
R31 commonsourceibias.n109 commonsourceibias.t97 168.701
R32 commonsourceibias.n85 commonsourceibias.t86 168.701
R33 commonsourceibias.n87 commonsourceibias.t115 168.701
R34 commonsourceibias.n89 commonsourceibias.t80 168.701
R35 commonsourceibias.n92 commonsourceibias.t66 168.701
R36 commonsourceibias.n219 commonsourceibias.t75 168.701
R37 commonsourceibias.n216 commonsourceibias.t60 168.701
R38 commonsourceibias.n214 commonsourceibias.t49 168.701
R39 commonsourceibias.n212 commonsourceibias.t84 168.701
R40 commonsourceibias.n236 commonsourceibias.t93 168.701
R41 commonsourceibias.n242 commonsourceibias.t53 168.701
R42 commonsourceibias.n209 commonsourceibias.t119 168.701
R43 commonsourceibias.n250 commonsourceibias.t104 168.701
R44 commonsourceibias.n256 commonsourceibias.t59 168.701
R45 commonsourceibias.n203 commonsourceibias.t50 168.701
R46 commonsourceibias.n139 commonsourceibias.t105 168.701
R47 commonsourceibias.n192 commonsourceibias.t101 168.701
R48 commonsourceibias.n186 commonsourceibias.t89 168.701
R49 commonsourceibias.n145 commonsourceibias.t106 168.701
R50 commonsourceibias.n178 commonsourceibias.t99 168.701
R51 commonsourceibias.n172 commonsourceibias.t87 168.701
R52 commonsourceibias.n148 commonsourceibias.t107 168.701
R53 commonsourceibias.n150 commonsourceibias.t100 168.701
R54 commonsourceibias.n152 commonsourceibias.t112 168.701
R55 commonsourceibias.n155 commonsourceibias.t108 168.701
R56 commonsourceibias.n323 commonsourceibias.t0 168.701
R57 commonsourceibias.n320 commonsourceibias.t6 168.701
R58 commonsourceibias.n318 commonsourceibias.t20 168.701
R59 commonsourceibias.n316 commonsourceibias.t10 168.701
R60 commonsourceibias.n340 commonsourceibias.t34 168.701
R61 commonsourceibias.n346 commonsourceibias.t40 168.701
R62 commonsourceibias.n348 commonsourceibias.t12 168.701
R63 commonsourceibias.n355 commonsourceibias.t18 168.701
R64 commonsourceibias.n361 commonsourceibias.t30 168.701
R65 commonsourceibias.n308 commonsourceibias.t28 168.701
R66 commonsourceibias.n267 commonsourceibias.t78 168.701
R67 commonsourceibias.n395 commonsourceibias.t52 168.701
R68 commonsourceibias.n389 commonsourceibias.t94 168.701
R69 commonsourceibias.n382 commonsourceibias.t64 168.701
R70 commonsourceibias.n380 commonsourceibias.t113 168.701
R71 commonsourceibias.n282 commonsourceibias.t58 168.701
R72 commonsourceibias.n279 commonsourceibias.t63 168.701
R73 commonsourceibias.n277 commonsourceibias.t92 168.701
R74 commonsourceibias.n275 commonsourceibias.t65 168.701
R75 commonsourceibias.n299 commonsourceibias.t76 168.701
R76 commonsourceibias.n484 commonsourceibias.t68 168.701
R77 commonsourceibias.n481 commonsourceibias.t72 168.701
R78 commonsourceibias.n479 commonsourceibias.t61 168.701
R79 commonsourceibias.n477 commonsourceibias.t109 168.701
R80 commonsourceibias.n501 commonsourceibias.t77 168.701
R81 commonsourceibias.n507 commonsourceibias.t67 168.701
R82 commonsourceibias.n509 commonsourceibias.t56 168.701
R83 commonsourceibias.n516 commonsourceibias.t48 168.701
R84 commonsourceibias.n522 commonsourceibias.t71 168.701
R85 commonsourceibias.n469 commonsourceibias.t62 168.701
R86 commonsourceibias.n420 commonsourceibias.t116 168.701
R87 commonsourceibias.n417 commonsourceibias.t102 168.701
R88 commonsourceibias.n415 commonsourceibias.t81 168.701
R89 commonsourceibias.n413 commonsourceibias.t95 168.701
R90 commonsourceibias.n437 commonsourceibias.t103 168.701
R91 commonsourceibias.n443 commonsourceibias.t83 168.701
R92 commonsourceibias.n445 commonsourceibias.t90 168.701
R93 commonsourceibias.n452 commonsourceibias.t73 168.701
R94 commonsourceibias.n458 commonsourceibias.t82 168.701
R95 commonsourceibias.n405 commonsourceibias.t91 168.701
R96 commonsourceibias.n27 commonsourceibias.n24 161.3
R97 commonsourceibias.n29 commonsourceibias.n28 161.3
R98 commonsourceibias.n31 commonsourceibias.n30 161.3
R99 commonsourceibias.n32 commonsourceibias.n22 161.3
R100 commonsourceibias.n34 commonsourceibias.n33 161.3
R101 commonsourceibias.n36 commonsourceibias.n35 161.3
R102 commonsourceibias.n37 commonsourceibias.n20 161.3
R103 commonsourceibias.n39 commonsourceibias.n38 161.3
R104 commonsourceibias.n41 commonsourceibias.n40 161.3
R105 commonsourceibias.n42 commonsourceibias.n18 161.3
R106 commonsourceibias.n45 commonsourceibias.n44 161.3
R107 commonsourceibias.n46 commonsourceibias.n17 161.3
R108 commonsourceibias.n48 commonsourceibias.n47 161.3
R109 commonsourceibias.n50 commonsourceibias.n15 161.3
R110 commonsourceibias.n52 commonsourceibias.n51 161.3
R111 commonsourceibias.n53 commonsourceibias.n14 161.3
R112 commonsourceibias.n55 commonsourceibias.n54 161.3
R113 commonsourceibias.n56 commonsourceibias.n13 161.3
R114 commonsourceibias.n59 commonsourceibias.n58 161.3
R115 commonsourceibias.n60 commonsourceibias.n12 161.3
R116 commonsourceibias.n62 commonsourceibias.n61 161.3
R117 commonsourceibias.n64 commonsourceibias.n11 161.3
R118 commonsourceibias.n66 commonsourceibias.n65 161.3
R119 commonsourceibias.n68 commonsourceibias.n67 161.3
R120 commonsourceibias.n69 commonsourceibias.n9 161.3
R121 commonsourceibias.n93 commonsourceibias.n90 161.3
R122 commonsourceibias.n95 commonsourceibias.n94 161.3
R123 commonsourceibias.n97 commonsourceibias.n96 161.3
R124 commonsourceibias.n98 commonsourceibias.n88 161.3
R125 commonsourceibias.n100 commonsourceibias.n99 161.3
R126 commonsourceibias.n102 commonsourceibias.n101 161.3
R127 commonsourceibias.n103 commonsourceibias.n86 161.3
R128 commonsourceibias.n105 commonsourceibias.n104 161.3
R129 commonsourceibias.n107 commonsourceibias.n106 161.3
R130 commonsourceibias.n108 commonsourceibias.n84 161.3
R131 commonsourceibias.n111 commonsourceibias.n110 161.3
R132 commonsourceibias.n112 commonsourceibias.n8 161.3
R133 commonsourceibias.n114 commonsourceibias.n113 161.3
R134 commonsourceibias.n116 commonsourceibias.n6 161.3
R135 commonsourceibias.n118 commonsourceibias.n117 161.3
R136 commonsourceibias.n119 commonsourceibias.n5 161.3
R137 commonsourceibias.n121 commonsourceibias.n120 161.3
R138 commonsourceibias.n122 commonsourceibias.n4 161.3
R139 commonsourceibias.n125 commonsourceibias.n124 161.3
R140 commonsourceibias.n126 commonsourceibias.n3 161.3
R141 commonsourceibias.n128 commonsourceibias.n127 161.3
R142 commonsourceibias.n130 commonsourceibias.n2 161.3
R143 commonsourceibias.n132 commonsourceibias.n131 161.3
R144 commonsourceibias.n134 commonsourceibias.n133 161.3
R145 commonsourceibias.n135 commonsourceibias.n0 161.3
R146 commonsourceibias.n262 commonsourceibias.n202 161.3
R147 commonsourceibias.n261 commonsourceibias.n260 161.3
R148 commonsourceibias.n259 commonsourceibias.n258 161.3
R149 commonsourceibias.n257 commonsourceibias.n204 161.3
R150 commonsourceibias.n255 commonsourceibias.n254 161.3
R151 commonsourceibias.n253 commonsourceibias.n205 161.3
R152 commonsourceibias.n252 commonsourceibias.n251 161.3
R153 commonsourceibias.n249 commonsourceibias.n206 161.3
R154 commonsourceibias.n248 commonsourceibias.n247 161.3
R155 commonsourceibias.n246 commonsourceibias.n207 161.3
R156 commonsourceibias.n245 commonsourceibias.n244 161.3
R157 commonsourceibias.n243 commonsourceibias.n208 161.3
R158 commonsourceibias.n241 commonsourceibias.n240 161.3
R159 commonsourceibias.n239 commonsourceibias.n210 161.3
R160 commonsourceibias.n238 commonsourceibias.n237 161.3
R161 commonsourceibias.n235 commonsourceibias.n211 161.3
R162 commonsourceibias.n234 commonsourceibias.n233 161.3
R163 commonsourceibias.n232 commonsourceibias.n231 161.3
R164 commonsourceibias.n230 commonsourceibias.n213 161.3
R165 commonsourceibias.n229 commonsourceibias.n228 161.3
R166 commonsourceibias.n227 commonsourceibias.n226 161.3
R167 commonsourceibias.n225 commonsourceibias.n215 161.3
R168 commonsourceibias.n224 commonsourceibias.n223 161.3
R169 commonsourceibias.n222 commonsourceibias.n221 161.3
R170 commonsourceibias.n220 commonsourceibias.n217 161.3
R171 commonsourceibias.n156 commonsourceibias.n153 161.3
R172 commonsourceibias.n158 commonsourceibias.n157 161.3
R173 commonsourceibias.n160 commonsourceibias.n159 161.3
R174 commonsourceibias.n161 commonsourceibias.n151 161.3
R175 commonsourceibias.n163 commonsourceibias.n162 161.3
R176 commonsourceibias.n165 commonsourceibias.n164 161.3
R177 commonsourceibias.n166 commonsourceibias.n149 161.3
R178 commonsourceibias.n168 commonsourceibias.n167 161.3
R179 commonsourceibias.n170 commonsourceibias.n169 161.3
R180 commonsourceibias.n171 commonsourceibias.n147 161.3
R181 commonsourceibias.n174 commonsourceibias.n173 161.3
R182 commonsourceibias.n175 commonsourceibias.n146 161.3
R183 commonsourceibias.n177 commonsourceibias.n176 161.3
R184 commonsourceibias.n179 commonsourceibias.n144 161.3
R185 commonsourceibias.n181 commonsourceibias.n180 161.3
R186 commonsourceibias.n182 commonsourceibias.n143 161.3
R187 commonsourceibias.n184 commonsourceibias.n183 161.3
R188 commonsourceibias.n185 commonsourceibias.n142 161.3
R189 commonsourceibias.n188 commonsourceibias.n187 161.3
R190 commonsourceibias.n189 commonsourceibias.n141 161.3
R191 commonsourceibias.n191 commonsourceibias.n190 161.3
R192 commonsourceibias.n193 commonsourceibias.n140 161.3
R193 commonsourceibias.n195 commonsourceibias.n194 161.3
R194 commonsourceibias.n197 commonsourceibias.n196 161.3
R195 commonsourceibias.n198 commonsourceibias.n138 161.3
R196 commonsourceibias.n367 commonsourceibias.n307 161.3
R197 commonsourceibias.n366 commonsourceibias.n365 161.3
R198 commonsourceibias.n364 commonsourceibias.n363 161.3
R199 commonsourceibias.n362 commonsourceibias.n309 161.3
R200 commonsourceibias.n360 commonsourceibias.n359 161.3
R201 commonsourceibias.n358 commonsourceibias.n310 161.3
R202 commonsourceibias.n357 commonsourceibias.n356 161.3
R203 commonsourceibias.n354 commonsourceibias.n311 161.3
R204 commonsourceibias.n353 commonsourceibias.n352 161.3
R205 commonsourceibias.n351 commonsourceibias.n312 161.3
R206 commonsourceibias.n350 commonsourceibias.n349 161.3
R207 commonsourceibias.n347 commonsourceibias.n313 161.3
R208 commonsourceibias.n345 commonsourceibias.n344 161.3
R209 commonsourceibias.n343 commonsourceibias.n314 161.3
R210 commonsourceibias.n342 commonsourceibias.n341 161.3
R211 commonsourceibias.n339 commonsourceibias.n315 161.3
R212 commonsourceibias.n338 commonsourceibias.n337 161.3
R213 commonsourceibias.n336 commonsourceibias.n335 161.3
R214 commonsourceibias.n334 commonsourceibias.n317 161.3
R215 commonsourceibias.n333 commonsourceibias.n332 161.3
R216 commonsourceibias.n331 commonsourceibias.n330 161.3
R217 commonsourceibias.n329 commonsourceibias.n319 161.3
R218 commonsourceibias.n328 commonsourceibias.n327 161.3
R219 commonsourceibias.n326 commonsourceibias.n325 161.3
R220 commonsourceibias.n324 commonsourceibias.n321 161.3
R221 commonsourceibias.n301 commonsourceibias.n300 161.3
R222 commonsourceibias.n298 commonsourceibias.n274 161.3
R223 commonsourceibias.n297 commonsourceibias.n296 161.3
R224 commonsourceibias.n295 commonsourceibias.n294 161.3
R225 commonsourceibias.n293 commonsourceibias.n276 161.3
R226 commonsourceibias.n292 commonsourceibias.n291 161.3
R227 commonsourceibias.n290 commonsourceibias.n289 161.3
R228 commonsourceibias.n288 commonsourceibias.n278 161.3
R229 commonsourceibias.n287 commonsourceibias.n286 161.3
R230 commonsourceibias.n285 commonsourceibias.n284 161.3
R231 commonsourceibias.n283 commonsourceibias.n280 161.3
R232 commonsourceibias.n377 commonsourceibias.n273 161.3
R233 commonsourceibias.n401 commonsourceibias.n266 161.3
R234 commonsourceibias.n400 commonsourceibias.n399 161.3
R235 commonsourceibias.n398 commonsourceibias.n397 161.3
R236 commonsourceibias.n396 commonsourceibias.n268 161.3
R237 commonsourceibias.n394 commonsourceibias.n393 161.3
R238 commonsourceibias.n392 commonsourceibias.n269 161.3
R239 commonsourceibias.n391 commonsourceibias.n390 161.3
R240 commonsourceibias.n388 commonsourceibias.n270 161.3
R241 commonsourceibias.n387 commonsourceibias.n386 161.3
R242 commonsourceibias.n385 commonsourceibias.n271 161.3
R243 commonsourceibias.n384 commonsourceibias.n383 161.3
R244 commonsourceibias.n381 commonsourceibias.n272 161.3
R245 commonsourceibias.n379 commonsourceibias.n378 161.3
R246 commonsourceibias.n528 commonsourceibias.n468 161.3
R247 commonsourceibias.n527 commonsourceibias.n526 161.3
R248 commonsourceibias.n525 commonsourceibias.n524 161.3
R249 commonsourceibias.n523 commonsourceibias.n470 161.3
R250 commonsourceibias.n521 commonsourceibias.n520 161.3
R251 commonsourceibias.n519 commonsourceibias.n471 161.3
R252 commonsourceibias.n518 commonsourceibias.n517 161.3
R253 commonsourceibias.n515 commonsourceibias.n472 161.3
R254 commonsourceibias.n514 commonsourceibias.n513 161.3
R255 commonsourceibias.n512 commonsourceibias.n473 161.3
R256 commonsourceibias.n511 commonsourceibias.n510 161.3
R257 commonsourceibias.n508 commonsourceibias.n474 161.3
R258 commonsourceibias.n506 commonsourceibias.n505 161.3
R259 commonsourceibias.n504 commonsourceibias.n475 161.3
R260 commonsourceibias.n503 commonsourceibias.n502 161.3
R261 commonsourceibias.n500 commonsourceibias.n476 161.3
R262 commonsourceibias.n499 commonsourceibias.n498 161.3
R263 commonsourceibias.n497 commonsourceibias.n496 161.3
R264 commonsourceibias.n495 commonsourceibias.n478 161.3
R265 commonsourceibias.n494 commonsourceibias.n493 161.3
R266 commonsourceibias.n492 commonsourceibias.n491 161.3
R267 commonsourceibias.n490 commonsourceibias.n480 161.3
R268 commonsourceibias.n489 commonsourceibias.n488 161.3
R269 commonsourceibias.n487 commonsourceibias.n486 161.3
R270 commonsourceibias.n485 commonsourceibias.n482 161.3
R271 commonsourceibias.n464 commonsourceibias.n404 161.3
R272 commonsourceibias.n463 commonsourceibias.n462 161.3
R273 commonsourceibias.n461 commonsourceibias.n460 161.3
R274 commonsourceibias.n459 commonsourceibias.n406 161.3
R275 commonsourceibias.n457 commonsourceibias.n456 161.3
R276 commonsourceibias.n455 commonsourceibias.n407 161.3
R277 commonsourceibias.n454 commonsourceibias.n453 161.3
R278 commonsourceibias.n451 commonsourceibias.n408 161.3
R279 commonsourceibias.n450 commonsourceibias.n449 161.3
R280 commonsourceibias.n448 commonsourceibias.n409 161.3
R281 commonsourceibias.n447 commonsourceibias.n446 161.3
R282 commonsourceibias.n444 commonsourceibias.n410 161.3
R283 commonsourceibias.n442 commonsourceibias.n441 161.3
R284 commonsourceibias.n440 commonsourceibias.n411 161.3
R285 commonsourceibias.n439 commonsourceibias.n438 161.3
R286 commonsourceibias.n436 commonsourceibias.n412 161.3
R287 commonsourceibias.n435 commonsourceibias.n434 161.3
R288 commonsourceibias.n433 commonsourceibias.n432 161.3
R289 commonsourceibias.n431 commonsourceibias.n414 161.3
R290 commonsourceibias.n430 commonsourceibias.n429 161.3
R291 commonsourceibias.n428 commonsourceibias.n427 161.3
R292 commonsourceibias.n426 commonsourceibias.n416 161.3
R293 commonsourceibias.n425 commonsourceibias.n424 161.3
R294 commonsourceibias.n423 commonsourceibias.n422 161.3
R295 commonsourceibias.n421 commonsourceibias.n418 161.3
R296 commonsourceibias.n80 commonsourceibias.n78 81.5057
R297 commonsourceibias.n304 commonsourceibias.n302 81.5057
R298 commonsourceibias.n80 commonsourceibias.n79 80.9324
R299 commonsourceibias.n82 commonsourceibias.n81 80.9324
R300 commonsourceibias.n77 commonsourceibias.n76 80.9324
R301 commonsourceibias.n75 commonsourceibias.n74 80.9324
R302 commonsourceibias.n73 commonsourceibias.n72 80.9324
R303 commonsourceibias.n371 commonsourceibias.n370 80.9324
R304 commonsourceibias.n373 commonsourceibias.n372 80.9324
R305 commonsourceibias.n375 commonsourceibias.n374 80.9324
R306 commonsourceibias.n306 commonsourceibias.n305 80.9324
R307 commonsourceibias.n304 commonsourceibias.n303 80.9324
R308 commonsourceibias.n71 commonsourceibias.n70 80.6037
R309 commonsourceibias.n137 commonsourceibias.n136 80.6037
R310 commonsourceibias.n264 commonsourceibias.n263 80.6037
R311 commonsourceibias.n200 commonsourceibias.n199 80.6037
R312 commonsourceibias.n369 commonsourceibias.n368 80.6037
R313 commonsourceibias.n403 commonsourceibias.n402 80.6037
R314 commonsourceibias.n530 commonsourceibias.n529 80.6037
R315 commonsourceibias.n466 commonsourceibias.n465 80.6037
R316 commonsourceibias.n65 commonsourceibias.n64 56.5617
R317 commonsourceibias.n51 commonsourceibias.n50 56.5617
R318 commonsourceibias.n42 commonsourceibias.n41 56.5617
R319 commonsourceibias.n28 commonsourceibias.n27 56.5617
R320 commonsourceibias.n131 commonsourceibias.n130 56.5617
R321 commonsourceibias.n117 commonsourceibias.n116 56.5617
R322 commonsourceibias.n108 commonsourceibias.n107 56.5617
R323 commonsourceibias.n94 commonsourceibias.n93 56.5617
R324 commonsourceibias.n221 commonsourceibias.n220 56.5617
R325 commonsourceibias.n235 commonsourceibias.n234 56.5617
R326 commonsourceibias.n244 commonsourceibias.n243 56.5617
R327 commonsourceibias.n258 commonsourceibias.n257 56.5617
R328 commonsourceibias.n194 commonsourceibias.n193 56.5617
R329 commonsourceibias.n180 commonsourceibias.n179 56.5617
R330 commonsourceibias.n171 commonsourceibias.n170 56.5617
R331 commonsourceibias.n157 commonsourceibias.n156 56.5617
R332 commonsourceibias.n325 commonsourceibias.n324 56.5617
R333 commonsourceibias.n339 commonsourceibias.n338 56.5617
R334 commonsourceibias.n349 commonsourceibias.n347 56.5617
R335 commonsourceibias.n363 commonsourceibias.n362 56.5617
R336 commonsourceibias.n397 commonsourceibias.n396 56.5617
R337 commonsourceibias.n383 commonsourceibias.n381 56.5617
R338 commonsourceibias.n284 commonsourceibias.n283 56.5617
R339 commonsourceibias.n298 commonsourceibias.n297 56.5617
R340 commonsourceibias.n486 commonsourceibias.n485 56.5617
R341 commonsourceibias.n500 commonsourceibias.n499 56.5617
R342 commonsourceibias.n510 commonsourceibias.n508 56.5617
R343 commonsourceibias.n524 commonsourceibias.n523 56.5617
R344 commonsourceibias.n422 commonsourceibias.n421 56.5617
R345 commonsourceibias.n436 commonsourceibias.n435 56.5617
R346 commonsourceibias.n446 commonsourceibias.n444 56.5617
R347 commonsourceibias.n460 commonsourceibias.n459 56.5617
R348 commonsourceibias.n56 commonsourceibias.n55 56.0773
R349 commonsourceibias.n37 commonsourceibias.n36 56.0773
R350 commonsourceibias.n122 commonsourceibias.n121 56.0773
R351 commonsourceibias.n103 commonsourceibias.n102 56.0773
R352 commonsourceibias.n230 commonsourceibias.n229 56.0773
R353 commonsourceibias.n249 commonsourceibias.n248 56.0773
R354 commonsourceibias.n185 commonsourceibias.n184 56.0773
R355 commonsourceibias.n166 commonsourceibias.n165 56.0773
R356 commonsourceibias.n334 commonsourceibias.n333 56.0773
R357 commonsourceibias.n354 commonsourceibias.n353 56.0773
R358 commonsourceibias.n388 commonsourceibias.n387 56.0773
R359 commonsourceibias.n293 commonsourceibias.n292 56.0773
R360 commonsourceibias.n495 commonsourceibias.n494 56.0773
R361 commonsourceibias.n515 commonsourceibias.n514 56.0773
R362 commonsourceibias.n431 commonsourceibias.n430 56.0773
R363 commonsourceibias.n451 commonsourceibias.n450 56.0773
R364 commonsourceibias.n70 commonsourceibias.n69 46.0096
R365 commonsourceibias.n136 commonsourceibias.n135 46.0096
R366 commonsourceibias.n263 commonsourceibias.n262 46.0096
R367 commonsourceibias.n199 commonsourceibias.n198 46.0096
R368 commonsourceibias.n368 commonsourceibias.n367 46.0096
R369 commonsourceibias.n402 commonsourceibias.n401 46.0096
R370 commonsourceibias.n529 commonsourceibias.n528 46.0096
R371 commonsourceibias.n465 commonsourceibias.n464 46.0096
R372 commonsourceibias.n58 commonsourceibias.n12 41.5458
R373 commonsourceibias.n33 commonsourceibias.n32 41.5458
R374 commonsourceibias.n124 commonsourceibias.n3 41.5458
R375 commonsourceibias.n99 commonsourceibias.n98 41.5458
R376 commonsourceibias.n226 commonsourceibias.n225 41.5458
R377 commonsourceibias.n251 commonsourceibias.n205 41.5458
R378 commonsourceibias.n187 commonsourceibias.n141 41.5458
R379 commonsourceibias.n162 commonsourceibias.n161 41.5458
R380 commonsourceibias.n330 commonsourceibias.n329 41.5458
R381 commonsourceibias.n356 commonsourceibias.n310 41.5458
R382 commonsourceibias.n390 commonsourceibias.n269 41.5458
R383 commonsourceibias.n289 commonsourceibias.n288 41.5458
R384 commonsourceibias.n491 commonsourceibias.n490 41.5458
R385 commonsourceibias.n517 commonsourceibias.n471 41.5458
R386 commonsourceibias.n427 commonsourceibias.n426 41.5458
R387 commonsourceibias.n453 commonsourceibias.n407 41.5458
R388 commonsourceibias.n48 commonsourceibias.n17 40.577
R389 commonsourceibias.n44 commonsourceibias.n17 40.577
R390 commonsourceibias.n114 commonsourceibias.n8 40.577
R391 commonsourceibias.n110 commonsourceibias.n8 40.577
R392 commonsourceibias.n237 commonsourceibias.n210 40.577
R393 commonsourceibias.n241 commonsourceibias.n210 40.577
R394 commonsourceibias.n177 commonsourceibias.n146 40.577
R395 commonsourceibias.n173 commonsourceibias.n146 40.577
R396 commonsourceibias.n341 commonsourceibias.n314 40.577
R397 commonsourceibias.n345 commonsourceibias.n314 40.577
R398 commonsourceibias.n379 commonsourceibias.n273 40.577
R399 commonsourceibias.n300 commonsourceibias.n273 40.577
R400 commonsourceibias.n502 commonsourceibias.n475 40.577
R401 commonsourceibias.n506 commonsourceibias.n475 40.577
R402 commonsourceibias.n438 commonsourceibias.n411 40.577
R403 commonsourceibias.n442 commonsourceibias.n411 40.577
R404 commonsourceibias.n62 commonsourceibias.n12 39.6083
R405 commonsourceibias.n32 commonsourceibias.n31 39.6083
R406 commonsourceibias.n128 commonsourceibias.n3 39.6083
R407 commonsourceibias.n98 commonsourceibias.n97 39.6083
R408 commonsourceibias.n225 commonsourceibias.n224 39.6083
R409 commonsourceibias.n255 commonsourceibias.n205 39.6083
R410 commonsourceibias.n191 commonsourceibias.n141 39.6083
R411 commonsourceibias.n161 commonsourceibias.n160 39.6083
R412 commonsourceibias.n329 commonsourceibias.n328 39.6083
R413 commonsourceibias.n360 commonsourceibias.n310 39.6083
R414 commonsourceibias.n394 commonsourceibias.n269 39.6083
R415 commonsourceibias.n288 commonsourceibias.n287 39.6083
R416 commonsourceibias.n490 commonsourceibias.n489 39.6083
R417 commonsourceibias.n521 commonsourceibias.n471 39.6083
R418 commonsourceibias.n426 commonsourceibias.n425 39.6083
R419 commonsourceibias.n457 commonsourceibias.n407 39.6083
R420 commonsourceibias.n26 commonsourceibias.n25 33.0515
R421 commonsourceibias.n92 commonsourceibias.n91 33.0515
R422 commonsourceibias.n155 commonsourceibias.n154 33.0515
R423 commonsourceibias.n219 commonsourceibias.n218 33.0515
R424 commonsourceibias.n323 commonsourceibias.n322 33.0515
R425 commonsourceibias.n282 commonsourceibias.n281 33.0515
R426 commonsourceibias.n484 commonsourceibias.n483 33.0515
R427 commonsourceibias.n420 commonsourceibias.n419 33.0515
R428 commonsourceibias.n25 commonsourceibias.n24 28.5514
R429 commonsourceibias.n91 commonsourceibias.n90 28.5514
R430 commonsourceibias.n218 commonsourceibias.n217 28.5514
R431 commonsourceibias.n154 commonsourceibias.n153 28.5514
R432 commonsourceibias.n322 commonsourceibias.n321 28.5514
R433 commonsourceibias.n281 commonsourceibias.n280 28.5514
R434 commonsourceibias.n483 commonsourceibias.n482 28.5514
R435 commonsourceibias.n419 commonsourceibias.n418 28.5514
R436 commonsourceibias.n69 commonsourceibias.n68 26.0455
R437 commonsourceibias.n135 commonsourceibias.n134 26.0455
R438 commonsourceibias.n262 commonsourceibias.n261 26.0455
R439 commonsourceibias.n198 commonsourceibias.n197 26.0455
R440 commonsourceibias.n367 commonsourceibias.n366 26.0455
R441 commonsourceibias.n401 commonsourceibias.n400 26.0455
R442 commonsourceibias.n528 commonsourceibias.n527 26.0455
R443 commonsourceibias.n464 commonsourceibias.n463 26.0455
R444 commonsourceibias.n55 commonsourceibias.n14 25.0767
R445 commonsourceibias.n38 commonsourceibias.n37 25.0767
R446 commonsourceibias.n121 commonsourceibias.n5 25.0767
R447 commonsourceibias.n104 commonsourceibias.n103 25.0767
R448 commonsourceibias.n231 commonsourceibias.n230 25.0767
R449 commonsourceibias.n248 commonsourceibias.n207 25.0767
R450 commonsourceibias.n184 commonsourceibias.n143 25.0767
R451 commonsourceibias.n167 commonsourceibias.n166 25.0767
R452 commonsourceibias.n335 commonsourceibias.n334 25.0767
R453 commonsourceibias.n353 commonsourceibias.n312 25.0767
R454 commonsourceibias.n387 commonsourceibias.n271 25.0767
R455 commonsourceibias.n294 commonsourceibias.n293 25.0767
R456 commonsourceibias.n496 commonsourceibias.n495 25.0767
R457 commonsourceibias.n514 commonsourceibias.n473 25.0767
R458 commonsourceibias.n432 commonsourceibias.n431 25.0767
R459 commonsourceibias.n450 commonsourceibias.n409 25.0767
R460 commonsourceibias.n51 commonsourceibias.n16 24.3464
R461 commonsourceibias.n41 commonsourceibias.n19 24.3464
R462 commonsourceibias.n117 commonsourceibias.n7 24.3464
R463 commonsourceibias.n107 commonsourceibias.n85 24.3464
R464 commonsourceibias.n234 commonsourceibias.n212 24.3464
R465 commonsourceibias.n244 commonsourceibias.n209 24.3464
R466 commonsourceibias.n180 commonsourceibias.n145 24.3464
R467 commonsourceibias.n170 commonsourceibias.n148 24.3464
R468 commonsourceibias.n338 commonsourceibias.n316 24.3464
R469 commonsourceibias.n349 commonsourceibias.n348 24.3464
R470 commonsourceibias.n383 commonsourceibias.n382 24.3464
R471 commonsourceibias.n297 commonsourceibias.n275 24.3464
R472 commonsourceibias.n499 commonsourceibias.n477 24.3464
R473 commonsourceibias.n510 commonsourceibias.n509 24.3464
R474 commonsourceibias.n435 commonsourceibias.n413 24.3464
R475 commonsourceibias.n446 commonsourceibias.n445 24.3464
R476 commonsourceibias.n65 commonsourceibias.n10 23.8546
R477 commonsourceibias.n27 commonsourceibias.n26 23.8546
R478 commonsourceibias.n131 commonsourceibias.n1 23.8546
R479 commonsourceibias.n93 commonsourceibias.n92 23.8546
R480 commonsourceibias.n220 commonsourceibias.n219 23.8546
R481 commonsourceibias.n258 commonsourceibias.n203 23.8546
R482 commonsourceibias.n194 commonsourceibias.n139 23.8546
R483 commonsourceibias.n156 commonsourceibias.n155 23.8546
R484 commonsourceibias.n324 commonsourceibias.n323 23.8546
R485 commonsourceibias.n363 commonsourceibias.n308 23.8546
R486 commonsourceibias.n397 commonsourceibias.n267 23.8546
R487 commonsourceibias.n283 commonsourceibias.n282 23.8546
R488 commonsourceibias.n485 commonsourceibias.n484 23.8546
R489 commonsourceibias.n524 commonsourceibias.n469 23.8546
R490 commonsourceibias.n421 commonsourceibias.n420 23.8546
R491 commonsourceibias.n460 commonsourceibias.n405 23.8546
R492 commonsourceibias.n64 commonsourceibias.n63 16.9689
R493 commonsourceibias.n28 commonsourceibias.n23 16.9689
R494 commonsourceibias.n130 commonsourceibias.n129 16.9689
R495 commonsourceibias.n94 commonsourceibias.n89 16.9689
R496 commonsourceibias.n221 commonsourceibias.n216 16.9689
R497 commonsourceibias.n257 commonsourceibias.n256 16.9689
R498 commonsourceibias.n193 commonsourceibias.n192 16.9689
R499 commonsourceibias.n157 commonsourceibias.n152 16.9689
R500 commonsourceibias.n325 commonsourceibias.n320 16.9689
R501 commonsourceibias.n362 commonsourceibias.n361 16.9689
R502 commonsourceibias.n396 commonsourceibias.n395 16.9689
R503 commonsourceibias.n284 commonsourceibias.n279 16.9689
R504 commonsourceibias.n486 commonsourceibias.n481 16.9689
R505 commonsourceibias.n523 commonsourceibias.n522 16.9689
R506 commonsourceibias.n422 commonsourceibias.n417 16.9689
R507 commonsourceibias.n459 commonsourceibias.n458 16.9689
R508 commonsourceibias.n50 commonsourceibias.n49 16.477
R509 commonsourceibias.n43 commonsourceibias.n42 16.477
R510 commonsourceibias.n116 commonsourceibias.n115 16.477
R511 commonsourceibias.n109 commonsourceibias.n108 16.477
R512 commonsourceibias.n236 commonsourceibias.n235 16.477
R513 commonsourceibias.n243 commonsourceibias.n242 16.477
R514 commonsourceibias.n179 commonsourceibias.n178 16.477
R515 commonsourceibias.n172 commonsourceibias.n171 16.477
R516 commonsourceibias.n340 commonsourceibias.n339 16.477
R517 commonsourceibias.n347 commonsourceibias.n346 16.477
R518 commonsourceibias.n381 commonsourceibias.n380 16.477
R519 commonsourceibias.n299 commonsourceibias.n298 16.477
R520 commonsourceibias.n501 commonsourceibias.n500 16.477
R521 commonsourceibias.n508 commonsourceibias.n507 16.477
R522 commonsourceibias.n437 commonsourceibias.n436 16.477
R523 commonsourceibias.n444 commonsourceibias.n443 16.477
R524 commonsourceibias.n57 commonsourceibias.n56 15.9852
R525 commonsourceibias.n36 commonsourceibias.n21 15.9852
R526 commonsourceibias.n123 commonsourceibias.n122 15.9852
R527 commonsourceibias.n102 commonsourceibias.n87 15.9852
R528 commonsourceibias.n229 commonsourceibias.n214 15.9852
R529 commonsourceibias.n250 commonsourceibias.n249 15.9852
R530 commonsourceibias.n186 commonsourceibias.n185 15.9852
R531 commonsourceibias.n165 commonsourceibias.n150 15.9852
R532 commonsourceibias.n333 commonsourceibias.n318 15.9852
R533 commonsourceibias.n355 commonsourceibias.n354 15.9852
R534 commonsourceibias.n389 commonsourceibias.n388 15.9852
R535 commonsourceibias.n292 commonsourceibias.n277 15.9852
R536 commonsourceibias.n494 commonsourceibias.n479 15.9852
R537 commonsourceibias.n516 commonsourceibias.n515 15.9852
R538 commonsourceibias.n430 commonsourceibias.n415 15.9852
R539 commonsourceibias.n452 commonsourceibias.n451 15.9852
R540 commonsourceibias.n73 commonsourceibias.n71 13.2057
R541 commonsourceibias.n371 commonsourceibias.n369 13.2057
R542 commonsourceibias.n532 commonsourceibias.n265 10.4122
R543 commonsourceibias.n112 commonsourceibias.n83 9.50363
R544 commonsourceibias.n377 commonsourceibias.n376 9.50363
R545 commonsourceibias.n201 commonsourceibias.n137 8.7339
R546 commonsourceibias.n467 commonsourceibias.n403 8.7339
R547 commonsourceibias.n58 commonsourceibias.n57 8.60764
R548 commonsourceibias.n33 commonsourceibias.n21 8.60764
R549 commonsourceibias.n124 commonsourceibias.n123 8.60764
R550 commonsourceibias.n99 commonsourceibias.n87 8.60764
R551 commonsourceibias.n226 commonsourceibias.n214 8.60764
R552 commonsourceibias.n251 commonsourceibias.n250 8.60764
R553 commonsourceibias.n187 commonsourceibias.n186 8.60764
R554 commonsourceibias.n162 commonsourceibias.n150 8.60764
R555 commonsourceibias.n330 commonsourceibias.n318 8.60764
R556 commonsourceibias.n356 commonsourceibias.n355 8.60764
R557 commonsourceibias.n390 commonsourceibias.n389 8.60764
R558 commonsourceibias.n289 commonsourceibias.n277 8.60764
R559 commonsourceibias.n491 commonsourceibias.n479 8.60764
R560 commonsourceibias.n517 commonsourceibias.n516 8.60764
R561 commonsourceibias.n427 commonsourceibias.n415 8.60764
R562 commonsourceibias.n453 commonsourceibias.n452 8.60764
R563 commonsourceibias.n532 commonsourceibias.n531 8.46921
R564 commonsourceibias.n49 commonsourceibias.n48 8.11581
R565 commonsourceibias.n44 commonsourceibias.n43 8.11581
R566 commonsourceibias.n115 commonsourceibias.n114 8.11581
R567 commonsourceibias.n110 commonsourceibias.n109 8.11581
R568 commonsourceibias.n237 commonsourceibias.n236 8.11581
R569 commonsourceibias.n242 commonsourceibias.n241 8.11581
R570 commonsourceibias.n178 commonsourceibias.n177 8.11581
R571 commonsourceibias.n173 commonsourceibias.n172 8.11581
R572 commonsourceibias.n341 commonsourceibias.n340 8.11581
R573 commonsourceibias.n346 commonsourceibias.n345 8.11581
R574 commonsourceibias.n380 commonsourceibias.n379 8.11581
R575 commonsourceibias.n300 commonsourceibias.n299 8.11581
R576 commonsourceibias.n502 commonsourceibias.n501 8.11581
R577 commonsourceibias.n507 commonsourceibias.n506 8.11581
R578 commonsourceibias.n438 commonsourceibias.n437 8.11581
R579 commonsourceibias.n443 commonsourceibias.n442 8.11581
R580 commonsourceibias.n63 commonsourceibias.n62 7.62397
R581 commonsourceibias.n31 commonsourceibias.n23 7.62397
R582 commonsourceibias.n129 commonsourceibias.n128 7.62397
R583 commonsourceibias.n97 commonsourceibias.n89 7.62397
R584 commonsourceibias.n224 commonsourceibias.n216 7.62397
R585 commonsourceibias.n256 commonsourceibias.n255 7.62397
R586 commonsourceibias.n192 commonsourceibias.n191 7.62397
R587 commonsourceibias.n160 commonsourceibias.n152 7.62397
R588 commonsourceibias.n328 commonsourceibias.n320 7.62397
R589 commonsourceibias.n361 commonsourceibias.n360 7.62397
R590 commonsourceibias.n395 commonsourceibias.n394 7.62397
R591 commonsourceibias.n287 commonsourceibias.n279 7.62397
R592 commonsourceibias.n489 commonsourceibias.n481 7.62397
R593 commonsourceibias.n522 commonsourceibias.n521 7.62397
R594 commonsourceibias.n425 commonsourceibias.n417 7.62397
R595 commonsourceibias.n458 commonsourceibias.n457 7.62397
R596 commonsourceibias.n265 commonsourceibias.n264 5.00473
R597 commonsourceibias.n201 commonsourceibias.n200 5.00473
R598 commonsourceibias.n531 commonsourceibias.n530 5.00473
R599 commonsourceibias.n467 commonsourceibias.n466 5.00473
R600 commonsourceibias commonsourceibias.n532 3.87639
R601 commonsourceibias.n265 commonsourceibias.n201 3.72967
R602 commonsourceibias.n531 commonsourceibias.n467 3.72967
R603 commonsourceibias.n78 commonsourceibias.t9 2.82907
R604 commonsourceibias.n78 commonsourceibias.t17 2.82907
R605 commonsourceibias.n79 commonsourceibias.t37 2.82907
R606 commonsourceibias.n79 commonsourceibias.t27 2.82907
R607 commonsourceibias.n81 commonsourceibias.t15 2.82907
R608 commonsourceibias.n81 commonsourceibias.t23 2.82907
R609 commonsourceibias.n76 commonsourceibias.t25 2.82907
R610 commonsourceibias.n76 commonsourceibias.t5 2.82907
R611 commonsourceibias.n74 commonsourceibias.t45 2.82907
R612 commonsourceibias.n74 commonsourceibias.t33 2.82907
R613 commonsourceibias.n72 commonsourceibias.t3 2.82907
R614 commonsourceibias.n72 commonsourceibias.t43 2.82907
R615 commonsourceibias.n370 commonsourceibias.t29 2.82907
R616 commonsourceibias.n370 commonsourceibias.t39 2.82907
R617 commonsourceibias.n372 commonsourceibias.t19 2.82907
R618 commonsourceibias.n372 commonsourceibias.t31 2.82907
R619 commonsourceibias.n374 commonsourceibias.t41 2.82907
R620 commonsourceibias.n374 commonsourceibias.t13 2.82907
R621 commonsourceibias.n305 commonsourceibias.t11 2.82907
R622 commonsourceibias.n305 commonsourceibias.t35 2.82907
R623 commonsourceibias.n303 commonsourceibias.t7 2.82907
R624 commonsourceibias.n303 commonsourceibias.t21 2.82907
R625 commonsourceibias.n302 commonsourceibias.t47 2.82907
R626 commonsourceibias.n302 commonsourceibias.t1 2.82907
R627 commonsourceibias.n68 commonsourceibias.n10 0.738255
R628 commonsourceibias.n134 commonsourceibias.n1 0.738255
R629 commonsourceibias.n261 commonsourceibias.n203 0.738255
R630 commonsourceibias.n197 commonsourceibias.n139 0.738255
R631 commonsourceibias.n366 commonsourceibias.n308 0.738255
R632 commonsourceibias.n400 commonsourceibias.n267 0.738255
R633 commonsourceibias.n527 commonsourceibias.n469 0.738255
R634 commonsourceibias.n463 commonsourceibias.n405 0.738255
R635 commonsourceibias.n75 commonsourceibias.n73 0.573776
R636 commonsourceibias.n77 commonsourceibias.n75 0.573776
R637 commonsourceibias.n82 commonsourceibias.n80 0.573776
R638 commonsourceibias.n306 commonsourceibias.n304 0.573776
R639 commonsourceibias.n375 commonsourceibias.n373 0.573776
R640 commonsourceibias.n373 commonsourceibias.n371 0.573776
R641 commonsourceibias.n83 commonsourceibias.n77 0.287138
R642 commonsourceibias.n83 commonsourceibias.n82 0.287138
R643 commonsourceibias.n376 commonsourceibias.n306 0.287138
R644 commonsourceibias.n376 commonsourceibias.n375 0.287138
R645 commonsourceibias.n71 commonsourceibias.n9 0.285035
R646 commonsourceibias.n137 commonsourceibias.n0 0.285035
R647 commonsourceibias.n264 commonsourceibias.n202 0.285035
R648 commonsourceibias.n200 commonsourceibias.n138 0.285035
R649 commonsourceibias.n369 commonsourceibias.n307 0.285035
R650 commonsourceibias.n403 commonsourceibias.n266 0.285035
R651 commonsourceibias.n530 commonsourceibias.n468 0.285035
R652 commonsourceibias.n466 commonsourceibias.n404 0.285035
R653 commonsourceibias.n16 commonsourceibias.n14 0.246418
R654 commonsourceibias.n38 commonsourceibias.n19 0.246418
R655 commonsourceibias.n7 commonsourceibias.n5 0.246418
R656 commonsourceibias.n104 commonsourceibias.n85 0.246418
R657 commonsourceibias.n231 commonsourceibias.n212 0.246418
R658 commonsourceibias.n209 commonsourceibias.n207 0.246418
R659 commonsourceibias.n145 commonsourceibias.n143 0.246418
R660 commonsourceibias.n167 commonsourceibias.n148 0.246418
R661 commonsourceibias.n335 commonsourceibias.n316 0.246418
R662 commonsourceibias.n348 commonsourceibias.n312 0.246418
R663 commonsourceibias.n382 commonsourceibias.n271 0.246418
R664 commonsourceibias.n294 commonsourceibias.n275 0.246418
R665 commonsourceibias.n496 commonsourceibias.n477 0.246418
R666 commonsourceibias.n509 commonsourceibias.n473 0.246418
R667 commonsourceibias.n432 commonsourceibias.n413 0.246418
R668 commonsourceibias.n445 commonsourceibias.n409 0.246418
R669 commonsourceibias.n67 commonsourceibias.n9 0.189894
R670 commonsourceibias.n67 commonsourceibias.n66 0.189894
R671 commonsourceibias.n66 commonsourceibias.n11 0.189894
R672 commonsourceibias.n61 commonsourceibias.n11 0.189894
R673 commonsourceibias.n61 commonsourceibias.n60 0.189894
R674 commonsourceibias.n60 commonsourceibias.n59 0.189894
R675 commonsourceibias.n59 commonsourceibias.n13 0.189894
R676 commonsourceibias.n54 commonsourceibias.n13 0.189894
R677 commonsourceibias.n54 commonsourceibias.n53 0.189894
R678 commonsourceibias.n53 commonsourceibias.n52 0.189894
R679 commonsourceibias.n52 commonsourceibias.n15 0.189894
R680 commonsourceibias.n47 commonsourceibias.n15 0.189894
R681 commonsourceibias.n47 commonsourceibias.n46 0.189894
R682 commonsourceibias.n46 commonsourceibias.n45 0.189894
R683 commonsourceibias.n45 commonsourceibias.n18 0.189894
R684 commonsourceibias.n40 commonsourceibias.n18 0.189894
R685 commonsourceibias.n40 commonsourceibias.n39 0.189894
R686 commonsourceibias.n39 commonsourceibias.n20 0.189894
R687 commonsourceibias.n35 commonsourceibias.n20 0.189894
R688 commonsourceibias.n35 commonsourceibias.n34 0.189894
R689 commonsourceibias.n34 commonsourceibias.n22 0.189894
R690 commonsourceibias.n30 commonsourceibias.n22 0.189894
R691 commonsourceibias.n30 commonsourceibias.n29 0.189894
R692 commonsourceibias.n29 commonsourceibias.n24 0.189894
R693 commonsourceibias.n111 commonsourceibias.n84 0.189894
R694 commonsourceibias.n106 commonsourceibias.n84 0.189894
R695 commonsourceibias.n106 commonsourceibias.n105 0.189894
R696 commonsourceibias.n105 commonsourceibias.n86 0.189894
R697 commonsourceibias.n101 commonsourceibias.n86 0.189894
R698 commonsourceibias.n101 commonsourceibias.n100 0.189894
R699 commonsourceibias.n100 commonsourceibias.n88 0.189894
R700 commonsourceibias.n96 commonsourceibias.n88 0.189894
R701 commonsourceibias.n96 commonsourceibias.n95 0.189894
R702 commonsourceibias.n95 commonsourceibias.n90 0.189894
R703 commonsourceibias.n133 commonsourceibias.n0 0.189894
R704 commonsourceibias.n133 commonsourceibias.n132 0.189894
R705 commonsourceibias.n132 commonsourceibias.n2 0.189894
R706 commonsourceibias.n127 commonsourceibias.n2 0.189894
R707 commonsourceibias.n127 commonsourceibias.n126 0.189894
R708 commonsourceibias.n126 commonsourceibias.n125 0.189894
R709 commonsourceibias.n125 commonsourceibias.n4 0.189894
R710 commonsourceibias.n120 commonsourceibias.n4 0.189894
R711 commonsourceibias.n120 commonsourceibias.n119 0.189894
R712 commonsourceibias.n119 commonsourceibias.n118 0.189894
R713 commonsourceibias.n118 commonsourceibias.n6 0.189894
R714 commonsourceibias.n113 commonsourceibias.n6 0.189894
R715 commonsourceibias.n260 commonsourceibias.n202 0.189894
R716 commonsourceibias.n260 commonsourceibias.n259 0.189894
R717 commonsourceibias.n259 commonsourceibias.n204 0.189894
R718 commonsourceibias.n254 commonsourceibias.n204 0.189894
R719 commonsourceibias.n254 commonsourceibias.n253 0.189894
R720 commonsourceibias.n253 commonsourceibias.n252 0.189894
R721 commonsourceibias.n252 commonsourceibias.n206 0.189894
R722 commonsourceibias.n247 commonsourceibias.n206 0.189894
R723 commonsourceibias.n247 commonsourceibias.n246 0.189894
R724 commonsourceibias.n246 commonsourceibias.n245 0.189894
R725 commonsourceibias.n245 commonsourceibias.n208 0.189894
R726 commonsourceibias.n240 commonsourceibias.n208 0.189894
R727 commonsourceibias.n240 commonsourceibias.n239 0.189894
R728 commonsourceibias.n239 commonsourceibias.n238 0.189894
R729 commonsourceibias.n238 commonsourceibias.n211 0.189894
R730 commonsourceibias.n233 commonsourceibias.n211 0.189894
R731 commonsourceibias.n233 commonsourceibias.n232 0.189894
R732 commonsourceibias.n232 commonsourceibias.n213 0.189894
R733 commonsourceibias.n228 commonsourceibias.n213 0.189894
R734 commonsourceibias.n228 commonsourceibias.n227 0.189894
R735 commonsourceibias.n227 commonsourceibias.n215 0.189894
R736 commonsourceibias.n223 commonsourceibias.n215 0.189894
R737 commonsourceibias.n223 commonsourceibias.n222 0.189894
R738 commonsourceibias.n222 commonsourceibias.n217 0.189894
R739 commonsourceibias.n196 commonsourceibias.n138 0.189894
R740 commonsourceibias.n196 commonsourceibias.n195 0.189894
R741 commonsourceibias.n195 commonsourceibias.n140 0.189894
R742 commonsourceibias.n190 commonsourceibias.n140 0.189894
R743 commonsourceibias.n190 commonsourceibias.n189 0.189894
R744 commonsourceibias.n189 commonsourceibias.n188 0.189894
R745 commonsourceibias.n188 commonsourceibias.n142 0.189894
R746 commonsourceibias.n183 commonsourceibias.n142 0.189894
R747 commonsourceibias.n183 commonsourceibias.n182 0.189894
R748 commonsourceibias.n182 commonsourceibias.n181 0.189894
R749 commonsourceibias.n181 commonsourceibias.n144 0.189894
R750 commonsourceibias.n176 commonsourceibias.n144 0.189894
R751 commonsourceibias.n176 commonsourceibias.n175 0.189894
R752 commonsourceibias.n175 commonsourceibias.n174 0.189894
R753 commonsourceibias.n174 commonsourceibias.n147 0.189894
R754 commonsourceibias.n169 commonsourceibias.n147 0.189894
R755 commonsourceibias.n169 commonsourceibias.n168 0.189894
R756 commonsourceibias.n168 commonsourceibias.n149 0.189894
R757 commonsourceibias.n164 commonsourceibias.n149 0.189894
R758 commonsourceibias.n164 commonsourceibias.n163 0.189894
R759 commonsourceibias.n163 commonsourceibias.n151 0.189894
R760 commonsourceibias.n159 commonsourceibias.n151 0.189894
R761 commonsourceibias.n159 commonsourceibias.n158 0.189894
R762 commonsourceibias.n158 commonsourceibias.n153 0.189894
R763 commonsourceibias.n326 commonsourceibias.n321 0.189894
R764 commonsourceibias.n327 commonsourceibias.n326 0.189894
R765 commonsourceibias.n327 commonsourceibias.n319 0.189894
R766 commonsourceibias.n331 commonsourceibias.n319 0.189894
R767 commonsourceibias.n332 commonsourceibias.n331 0.189894
R768 commonsourceibias.n332 commonsourceibias.n317 0.189894
R769 commonsourceibias.n336 commonsourceibias.n317 0.189894
R770 commonsourceibias.n337 commonsourceibias.n336 0.189894
R771 commonsourceibias.n337 commonsourceibias.n315 0.189894
R772 commonsourceibias.n342 commonsourceibias.n315 0.189894
R773 commonsourceibias.n343 commonsourceibias.n342 0.189894
R774 commonsourceibias.n344 commonsourceibias.n343 0.189894
R775 commonsourceibias.n344 commonsourceibias.n313 0.189894
R776 commonsourceibias.n350 commonsourceibias.n313 0.189894
R777 commonsourceibias.n351 commonsourceibias.n350 0.189894
R778 commonsourceibias.n352 commonsourceibias.n351 0.189894
R779 commonsourceibias.n352 commonsourceibias.n311 0.189894
R780 commonsourceibias.n357 commonsourceibias.n311 0.189894
R781 commonsourceibias.n358 commonsourceibias.n357 0.189894
R782 commonsourceibias.n359 commonsourceibias.n358 0.189894
R783 commonsourceibias.n359 commonsourceibias.n309 0.189894
R784 commonsourceibias.n364 commonsourceibias.n309 0.189894
R785 commonsourceibias.n365 commonsourceibias.n364 0.189894
R786 commonsourceibias.n365 commonsourceibias.n307 0.189894
R787 commonsourceibias.n285 commonsourceibias.n280 0.189894
R788 commonsourceibias.n286 commonsourceibias.n285 0.189894
R789 commonsourceibias.n286 commonsourceibias.n278 0.189894
R790 commonsourceibias.n290 commonsourceibias.n278 0.189894
R791 commonsourceibias.n291 commonsourceibias.n290 0.189894
R792 commonsourceibias.n291 commonsourceibias.n276 0.189894
R793 commonsourceibias.n295 commonsourceibias.n276 0.189894
R794 commonsourceibias.n296 commonsourceibias.n295 0.189894
R795 commonsourceibias.n296 commonsourceibias.n274 0.189894
R796 commonsourceibias.n301 commonsourceibias.n274 0.189894
R797 commonsourceibias.n378 commonsourceibias.n272 0.189894
R798 commonsourceibias.n384 commonsourceibias.n272 0.189894
R799 commonsourceibias.n385 commonsourceibias.n384 0.189894
R800 commonsourceibias.n386 commonsourceibias.n385 0.189894
R801 commonsourceibias.n386 commonsourceibias.n270 0.189894
R802 commonsourceibias.n391 commonsourceibias.n270 0.189894
R803 commonsourceibias.n392 commonsourceibias.n391 0.189894
R804 commonsourceibias.n393 commonsourceibias.n392 0.189894
R805 commonsourceibias.n393 commonsourceibias.n268 0.189894
R806 commonsourceibias.n398 commonsourceibias.n268 0.189894
R807 commonsourceibias.n399 commonsourceibias.n398 0.189894
R808 commonsourceibias.n399 commonsourceibias.n266 0.189894
R809 commonsourceibias.n487 commonsourceibias.n482 0.189894
R810 commonsourceibias.n488 commonsourceibias.n487 0.189894
R811 commonsourceibias.n488 commonsourceibias.n480 0.189894
R812 commonsourceibias.n492 commonsourceibias.n480 0.189894
R813 commonsourceibias.n493 commonsourceibias.n492 0.189894
R814 commonsourceibias.n493 commonsourceibias.n478 0.189894
R815 commonsourceibias.n497 commonsourceibias.n478 0.189894
R816 commonsourceibias.n498 commonsourceibias.n497 0.189894
R817 commonsourceibias.n498 commonsourceibias.n476 0.189894
R818 commonsourceibias.n503 commonsourceibias.n476 0.189894
R819 commonsourceibias.n504 commonsourceibias.n503 0.189894
R820 commonsourceibias.n505 commonsourceibias.n504 0.189894
R821 commonsourceibias.n505 commonsourceibias.n474 0.189894
R822 commonsourceibias.n511 commonsourceibias.n474 0.189894
R823 commonsourceibias.n512 commonsourceibias.n511 0.189894
R824 commonsourceibias.n513 commonsourceibias.n512 0.189894
R825 commonsourceibias.n513 commonsourceibias.n472 0.189894
R826 commonsourceibias.n518 commonsourceibias.n472 0.189894
R827 commonsourceibias.n519 commonsourceibias.n518 0.189894
R828 commonsourceibias.n520 commonsourceibias.n519 0.189894
R829 commonsourceibias.n520 commonsourceibias.n470 0.189894
R830 commonsourceibias.n525 commonsourceibias.n470 0.189894
R831 commonsourceibias.n526 commonsourceibias.n525 0.189894
R832 commonsourceibias.n526 commonsourceibias.n468 0.189894
R833 commonsourceibias.n423 commonsourceibias.n418 0.189894
R834 commonsourceibias.n424 commonsourceibias.n423 0.189894
R835 commonsourceibias.n424 commonsourceibias.n416 0.189894
R836 commonsourceibias.n428 commonsourceibias.n416 0.189894
R837 commonsourceibias.n429 commonsourceibias.n428 0.189894
R838 commonsourceibias.n429 commonsourceibias.n414 0.189894
R839 commonsourceibias.n433 commonsourceibias.n414 0.189894
R840 commonsourceibias.n434 commonsourceibias.n433 0.189894
R841 commonsourceibias.n434 commonsourceibias.n412 0.189894
R842 commonsourceibias.n439 commonsourceibias.n412 0.189894
R843 commonsourceibias.n440 commonsourceibias.n439 0.189894
R844 commonsourceibias.n441 commonsourceibias.n440 0.189894
R845 commonsourceibias.n441 commonsourceibias.n410 0.189894
R846 commonsourceibias.n447 commonsourceibias.n410 0.189894
R847 commonsourceibias.n448 commonsourceibias.n447 0.189894
R848 commonsourceibias.n449 commonsourceibias.n448 0.189894
R849 commonsourceibias.n449 commonsourceibias.n408 0.189894
R850 commonsourceibias.n454 commonsourceibias.n408 0.189894
R851 commonsourceibias.n455 commonsourceibias.n454 0.189894
R852 commonsourceibias.n456 commonsourceibias.n455 0.189894
R853 commonsourceibias.n456 commonsourceibias.n406 0.189894
R854 commonsourceibias.n461 commonsourceibias.n406 0.189894
R855 commonsourceibias.n462 commonsourceibias.n461 0.189894
R856 commonsourceibias.n462 commonsourceibias.n404 0.189894
R857 commonsourceibias.n112 commonsourceibias.n111 0.170955
R858 commonsourceibias.n113 commonsourceibias.n112 0.170955
R859 commonsourceibias.n377 commonsourceibias.n301 0.170955
R860 commonsourceibias.n378 commonsourceibias.n377 0.170955
R861 gnd.n7003 gnd.n536 1868.32
R862 gnd.n6323 gnd.n6276 939.716
R863 gnd.n7356 gnd.n172 838.452
R864 gnd.n7324 gnd.n170 838.452
R865 gnd.n3268 gnd.n3156 838.452
R866 gnd.n5527 gnd.n3270 838.452
R867 gnd.n6047 gnd.n2636 838.452
R868 gnd.n5967 gnd.n2634 838.452
R869 gnd.n4153 gnd.n2379 838.452
R870 gnd.n4109 gnd.n4108 838.452
R871 gnd.n7358 gnd.n167 783.196
R872 gnd.n383 gnd.n169 783.196
R873 gnd.n5530 gnd.n5529 783.196
R874 gnd.n5647 gnd.n3202 783.196
R875 gnd.n6049 gnd.n2631 783.196
R876 gnd.n2842 gnd.n2633 783.196
R877 gnd.n6154 gnd.n2452 783.196
R878 gnd.n6274 gnd.n2383 783.196
R879 gnd.n6338 gnd.n1045 766.379
R880 gnd.n2340 gnd.n1042 766.379
R881 gnd.n1504 gnd.n1403 766.379
R882 gnd.n1502 gnd.n1405 766.379
R883 gnd.n6322 gnd.n1039 756.769
R884 gnd.n6333 gnd.n6332 756.769
R885 gnd.n1749 gnd.n1365 756.769
R886 gnd.n1735 gnd.n1355 756.769
R887 gnd.n6028 gnd.n2666 711.122
R888 gnd.n5716 gnd.n3092 711.122
R889 gnd.n6032 gnd.n2648 711.122
R890 gnd.n5718 gnd.n3087 711.122
R891 gnd.n6545 gnd.n809 670.282
R892 gnd.n7002 gnd.n537 670.282
R893 gnd.n7214 gnd.n7213 670.282
R894 gnd.n4068 gnd.n977 670.282
R895 gnd.n812 gnd.n809 585
R896 gnd.n6543 gnd.n809 585
R897 gnd.n6541 gnd.n6540 585
R898 gnd.n6542 gnd.n6541 585
R899 gnd.n6539 gnd.n811 585
R900 gnd.n811 gnd.n810 585
R901 gnd.n6538 gnd.n6537 585
R902 gnd.n6537 gnd.n6536 585
R903 gnd.n817 gnd.n816 585
R904 gnd.n6535 gnd.n817 585
R905 gnd.n6533 gnd.n6532 585
R906 gnd.n6534 gnd.n6533 585
R907 gnd.n6531 gnd.n819 585
R908 gnd.n819 gnd.n818 585
R909 gnd.n6530 gnd.n6529 585
R910 gnd.n6529 gnd.n6528 585
R911 gnd.n825 gnd.n824 585
R912 gnd.n6527 gnd.n825 585
R913 gnd.n6525 gnd.n6524 585
R914 gnd.n6526 gnd.n6525 585
R915 gnd.n6523 gnd.n827 585
R916 gnd.n827 gnd.n826 585
R917 gnd.n6522 gnd.n6521 585
R918 gnd.n6521 gnd.n6520 585
R919 gnd.n833 gnd.n832 585
R920 gnd.n6519 gnd.n833 585
R921 gnd.n6517 gnd.n6516 585
R922 gnd.n6518 gnd.n6517 585
R923 gnd.n6515 gnd.n835 585
R924 gnd.n835 gnd.n834 585
R925 gnd.n6514 gnd.n6513 585
R926 gnd.n6513 gnd.n6512 585
R927 gnd.n841 gnd.n840 585
R928 gnd.n6511 gnd.n841 585
R929 gnd.n6509 gnd.n6508 585
R930 gnd.n6510 gnd.n6509 585
R931 gnd.n6507 gnd.n843 585
R932 gnd.n843 gnd.n842 585
R933 gnd.n6506 gnd.n6505 585
R934 gnd.n6505 gnd.n6504 585
R935 gnd.n849 gnd.n848 585
R936 gnd.n6503 gnd.n849 585
R937 gnd.n6501 gnd.n6500 585
R938 gnd.n6502 gnd.n6501 585
R939 gnd.n6499 gnd.n851 585
R940 gnd.n851 gnd.n850 585
R941 gnd.n6498 gnd.n6497 585
R942 gnd.n6497 gnd.n6496 585
R943 gnd.n857 gnd.n856 585
R944 gnd.n6495 gnd.n857 585
R945 gnd.n6493 gnd.n6492 585
R946 gnd.n6494 gnd.n6493 585
R947 gnd.n6491 gnd.n859 585
R948 gnd.n859 gnd.n858 585
R949 gnd.n6490 gnd.n6489 585
R950 gnd.n6489 gnd.n6488 585
R951 gnd.n865 gnd.n864 585
R952 gnd.n6487 gnd.n865 585
R953 gnd.n6485 gnd.n6484 585
R954 gnd.n6486 gnd.n6485 585
R955 gnd.n6483 gnd.n867 585
R956 gnd.n867 gnd.n866 585
R957 gnd.n6482 gnd.n6481 585
R958 gnd.n6481 gnd.n6480 585
R959 gnd.n873 gnd.n872 585
R960 gnd.n6479 gnd.n873 585
R961 gnd.n6477 gnd.n6476 585
R962 gnd.n6478 gnd.n6477 585
R963 gnd.n6475 gnd.n875 585
R964 gnd.n875 gnd.n874 585
R965 gnd.n6474 gnd.n6473 585
R966 gnd.n6473 gnd.n6472 585
R967 gnd.n881 gnd.n880 585
R968 gnd.n6471 gnd.n881 585
R969 gnd.n6469 gnd.n6468 585
R970 gnd.n6470 gnd.n6469 585
R971 gnd.n6467 gnd.n883 585
R972 gnd.n883 gnd.n882 585
R973 gnd.n6466 gnd.n6465 585
R974 gnd.n6465 gnd.n6464 585
R975 gnd.n889 gnd.n888 585
R976 gnd.n6463 gnd.n889 585
R977 gnd.n6461 gnd.n6460 585
R978 gnd.n6462 gnd.n6461 585
R979 gnd.n6459 gnd.n891 585
R980 gnd.n891 gnd.n890 585
R981 gnd.n6458 gnd.n6457 585
R982 gnd.n6457 gnd.n6456 585
R983 gnd.n897 gnd.n896 585
R984 gnd.n6455 gnd.n897 585
R985 gnd.n6453 gnd.n6452 585
R986 gnd.n6454 gnd.n6453 585
R987 gnd.n6451 gnd.n899 585
R988 gnd.n899 gnd.n898 585
R989 gnd.n6450 gnd.n6449 585
R990 gnd.n6449 gnd.n6448 585
R991 gnd.n905 gnd.n904 585
R992 gnd.n6447 gnd.n905 585
R993 gnd.n6445 gnd.n6444 585
R994 gnd.n6446 gnd.n6445 585
R995 gnd.n6443 gnd.n907 585
R996 gnd.n907 gnd.n906 585
R997 gnd.n6442 gnd.n6441 585
R998 gnd.n6441 gnd.n6440 585
R999 gnd.n913 gnd.n912 585
R1000 gnd.n6439 gnd.n913 585
R1001 gnd.n6437 gnd.n6436 585
R1002 gnd.n6438 gnd.n6437 585
R1003 gnd.n6435 gnd.n915 585
R1004 gnd.n915 gnd.n914 585
R1005 gnd.n6434 gnd.n6433 585
R1006 gnd.n6433 gnd.n6432 585
R1007 gnd.n921 gnd.n920 585
R1008 gnd.n6431 gnd.n921 585
R1009 gnd.n6429 gnd.n6428 585
R1010 gnd.n6430 gnd.n6429 585
R1011 gnd.n6427 gnd.n923 585
R1012 gnd.n923 gnd.n922 585
R1013 gnd.n6426 gnd.n6425 585
R1014 gnd.n6425 gnd.n6424 585
R1015 gnd.n929 gnd.n928 585
R1016 gnd.n6423 gnd.n929 585
R1017 gnd.n6421 gnd.n6420 585
R1018 gnd.n6422 gnd.n6421 585
R1019 gnd.n6419 gnd.n931 585
R1020 gnd.n931 gnd.n930 585
R1021 gnd.n6418 gnd.n6417 585
R1022 gnd.n6417 gnd.n6416 585
R1023 gnd.n937 gnd.n936 585
R1024 gnd.n6415 gnd.n937 585
R1025 gnd.n6413 gnd.n6412 585
R1026 gnd.n6414 gnd.n6413 585
R1027 gnd.n6411 gnd.n939 585
R1028 gnd.n939 gnd.n938 585
R1029 gnd.n6410 gnd.n6409 585
R1030 gnd.n6409 gnd.n6408 585
R1031 gnd.n945 gnd.n944 585
R1032 gnd.n6407 gnd.n945 585
R1033 gnd.n6405 gnd.n6404 585
R1034 gnd.n6406 gnd.n6405 585
R1035 gnd.n6403 gnd.n947 585
R1036 gnd.n947 gnd.n946 585
R1037 gnd.n6402 gnd.n6401 585
R1038 gnd.n6401 gnd.n6400 585
R1039 gnd.n953 gnd.n952 585
R1040 gnd.n6399 gnd.n953 585
R1041 gnd.n6397 gnd.n6396 585
R1042 gnd.n6398 gnd.n6397 585
R1043 gnd.n6395 gnd.n955 585
R1044 gnd.n955 gnd.n954 585
R1045 gnd.n6394 gnd.n6393 585
R1046 gnd.n6393 gnd.n6392 585
R1047 gnd.n961 gnd.n960 585
R1048 gnd.n6391 gnd.n961 585
R1049 gnd.n6389 gnd.n6388 585
R1050 gnd.n6390 gnd.n6389 585
R1051 gnd.n6387 gnd.n963 585
R1052 gnd.n963 gnd.n962 585
R1053 gnd.n6386 gnd.n6385 585
R1054 gnd.n6385 gnd.n6384 585
R1055 gnd.n969 gnd.n968 585
R1056 gnd.n6383 gnd.n969 585
R1057 gnd.n6381 gnd.n6380 585
R1058 gnd.n6382 gnd.n6381 585
R1059 gnd.n6379 gnd.n971 585
R1060 gnd.n971 gnd.n970 585
R1061 gnd.n6378 gnd.n6377 585
R1062 gnd.n6377 gnd.n6376 585
R1063 gnd.n6546 gnd.n6545 585
R1064 gnd.n6545 gnd.n6544 585
R1065 gnd.n807 gnd.n806 585
R1066 gnd.n806 gnd.n805 585
R1067 gnd.n6551 gnd.n6550 585
R1068 gnd.n6552 gnd.n6551 585
R1069 gnd.n804 gnd.n803 585
R1070 gnd.n6553 gnd.n804 585
R1071 gnd.n6556 gnd.n6555 585
R1072 gnd.n6555 gnd.n6554 585
R1073 gnd.n801 gnd.n800 585
R1074 gnd.n800 gnd.n799 585
R1075 gnd.n6561 gnd.n6560 585
R1076 gnd.n6562 gnd.n6561 585
R1077 gnd.n798 gnd.n797 585
R1078 gnd.n6563 gnd.n798 585
R1079 gnd.n6566 gnd.n6565 585
R1080 gnd.n6565 gnd.n6564 585
R1081 gnd.n795 gnd.n794 585
R1082 gnd.n794 gnd.n793 585
R1083 gnd.n6571 gnd.n6570 585
R1084 gnd.n6572 gnd.n6571 585
R1085 gnd.n792 gnd.n791 585
R1086 gnd.n6573 gnd.n792 585
R1087 gnd.n6576 gnd.n6575 585
R1088 gnd.n6575 gnd.n6574 585
R1089 gnd.n789 gnd.n788 585
R1090 gnd.n788 gnd.n787 585
R1091 gnd.n6581 gnd.n6580 585
R1092 gnd.n6582 gnd.n6581 585
R1093 gnd.n786 gnd.n785 585
R1094 gnd.n6583 gnd.n786 585
R1095 gnd.n6586 gnd.n6585 585
R1096 gnd.n6585 gnd.n6584 585
R1097 gnd.n783 gnd.n782 585
R1098 gnd.n782 gnd.n781 585
R1099 gnd.n6591 gnd.n6590 585
R1100 gnd.n6592 gnd.n6591 585
R1101 gnd.n780 gnd.n779 585
R1102 gnd.n6593 gnd.n780 585
R1103 gnd.n6596 gnd.n6595 585
R1104 gnd.n6595 gnd.n6594 585
R1105 gnd.n777 gnd.n776 585
R1106 gnd.n776 gnd.n775 585
R1107 gnd.n6601 gnd.n6600 585
R1108 gnd.n6602 gnd.n6601 585
R1109 gnd.n774 gnd.n773 585
R1110 gnd.n6603 gnd.n774 585
R1111 gnd.n6606 gnd.n6605 585
R1112 gnd.n6605 gnd.n6604 585
R1113 gnd.n771 gnd.n770 585
R1114 gnd.n770 gnd.n769 585
R1115 gnd.n6611 gnd.n6610 585
R1116 gnd.n6612 gnd.n6611 585
R1117 gnd.n768 gnd.n767 585
R1118 gnd.n6613 gnd.n768 585
R1119 gnd.n6616 gnd.n6615 585
R1120 gnd.n6615 gnd.n6614 585
R1121 gnd.n765 gnd.n764 585
R1122 gnd.n764 gnd.n763 585
R1123 gnd.n6621 gnd.n6620 585
R1124 gnd.n6622 gnd.n6621 585
R1125 gnd.n762 gnd.n761 585
R1126 gnd.n6623 gnd.n762 585
R1127 gnd.n6626 gnd.n6625 585
R1128 gnd.n6625 gnd.n6624 585
R1129 gnd.n759 gnd.n758 585
R1130 gnd.n758 gnd.n757 585
R1131 gnd.n6631 gnd.n6630 585
R1132 gnd.n6632 gnd.n6631 585
R1133 gnd.n756 gnd.n755 585
R1134 gnd.n6633 gnd.n756 585
R1135 gnd.n6636 gnd.n6635 585
R1136 gnd.n6635 gnd.n6634 585
R1137 gnd.n753 gnd.n752 585
R1138 gnd.n752 gnd.n751 585
R1139 gnd.n6641 gnd.n6640 585
R1140 gnd.n6642 gnd.n6641 585
R1141 gnd.n750 gnd.n749 585
R1142 gnd.n6643 gnd.n750 585
R1143 gnd.n6646 gnd.n6645 585
R1144 gnd.n6645 gnd.n6644 585
R1145 gnd.n747 gnd.n746 585
R1146 gnd.n746 gnd.n745 585
R1147 gnd.n6651 gnd.n6650 585
R1148 gnd.n6652 gnd.n6651 585
R1149 gnd.n744 gnd.n743 585
R1150 gnd.n6653 gnd.n744 585
R1151 gnd.n6656 gnd.n6655 585
R1152 gnd.n6655 gnd.n6654 585
R1153 gnd.n741 gnd.n740 585
R1154 gnd.n740 gnd.n739 585
R1155 gnd.n6661 gnd.n6660 585
R1156 gnd.n6662 gnd.n6661 585
R1157 gnd.n738 gnd.n737 585
R1158 gnd.n6663 gnd.n738 585
R1159 gnd.n6666 gnd.n6665 585
R1160 gnd.n6665 gnd.n6664 585
R1161 gnd.n735 gnd.n734 585
R1162 gnd.n734 gnd.n733 585
R1163 gnd.n6671 gnd.n6670 585
R1164 gnd.n6672 gnd.n6671 585
R1165 gnd.n732 gnd.n731 585
R1166 gnd.n6673 gnd.n732 585
R1167 gnd.n6676 gnd.n6675 585
R1168 gnd.n6675 gnd.n6674 585
R1169 gnd.n729 gnd.n728 585
R1170 gnd.n728 gnd.n727 585
R1171 gnd.n6681 gnd.n6680 585
R1172 gnd.n6682 gnd.n6681 585
R1173 gnd.n726 gnd.n725 585
R1174 gnd.n6683 gnd.n726 585
R1175 gnd.n6686 gnd.n6685 585
R1176 gnd.n6685 gnd.n6684 585
R1177 gnd.n723 gnd.n722 585
R1178 gnd.n722 gnd.n721 585
R1179 gnd.n6691 gnd.n6690 585
R1180 gnd.n6692 gnd.n6691 585
R1181 gnd.n720 gnd.n719 585
R1182 gnd.n6693 gnd.n720 585
R1183 gnd.n6696 gnd.n6695 585
R1184 gnd.n6695 gnd.n6694 585
R1185 gnd.n717 gnd.n716 585
R1186 gnd.n716 gnd.n715 585
R1187 gnd.n6701 gnd.n6700 585
R1188 gnd.n6702 gnd.n6701 585
R1189 gnd.n714 gnd.n713 585
R1190 gnd.n6703 gnd.n714 585
R1191 gnd.n6706 gnd.n6705 585
R1192 gnd.n6705 gnd.n6704 585
R1193 gnd.n711 gnd.n710 585
R1194 gnd.n710 gnd.n709 585
R1195 gnd.n6711 gnd.n6710 585
R1196 gnd.n6712 gnd.n6711 585
R1197 gnd.n708 gnd.n707 585
R1198 gnd.n6713 gnd.n708 585
R1199 gnd.n6716 gnd.n6715 585
R1200 gnd.n6715 gnd.n6714 585
R1201 gnd.n705 gnd.n704 585
R1202 gnd.n704 gnd.n703 585
R1203 gnd.n6721 gnd.n6720 585
R1204 gnd.n6722 gnd.n6721 585
R1205 gnd.n702 gnd.n701 585
R1206 gnd.n6723 gnd.n702 585
R1207 gnd.n6726 gnd.n6725 585
R1208 gnd.n6725 gnd.n6724 585
R1209 gnd.n699 gnd.n698 585
R1210 gnd.n698 gnd.n697 585
R1211 gnd.n6731 gnd.n6730 585
R1212 gnd.n6732 gnd.n6731 585
R1213 gnd.n696 gnd.n695 585
R1214 gnd.n6733 gnd.n696 585
R1215 gnd.n6736 gnd.n6735 585
R1216 gnd.n6735 gnd.n6734 585
R1217 gnd.n693 gnd.n692 585
R1218 gnd.n692 gnd.n691 585
R1219 gnd.n6741 gnd.n6740 585
R1220 gnd.n6742 gnd.n6741 585
R1221 gnd.n690 gnd.n689 585
R1222 gnd.n6743 gnd.n690 585
R1223 gnd.n6746 gnd.n6745 585
R1224 gnd.n6745 gnd.n6744 585
R1225 gnd.n687 gnd.n686 585
R1226 gnd.n686 gnd.n685 585
R1227 gnd.n6751 gnd.n6750 585
R1228 gnd.n6752 gnd.n6751 585
R1229 gnd.n684 gnd.n683 585
R1230 gnd.n6753 gnd.n684 585
R1231 gnd.n6756 gnd.n6755 585
R1232 gnd.n6755 gnd.n6754 585
R1233 gnd.n681 gnd.n680 585
R1234 gnd.n680 gnd.n679 585
R1235 gnd.n6761 gnd.n6760 585
R1236 gnd.n6762 gnd.n6761 585
R1237 gnd.n678 gnd.n677 585
R1238 gnd.n6763 gnd.n678 585
R1239 gnd.n6766 gnd.n6765 585
R1240 gnd.n6765 gnd.n6764 585
R1241 gnd.n675 gnd.n674 585
R1242 gnd.n674 gnd.n673 585
R1243 gnd.n6771 gnd.n6770 585
R1244 gnd.n6772 gnd.n6771 585
R1245 gnd.n672 gnd.n671 585
R1246 gnd.n6773 gnd.n672 585
R1247 gnd.n6776 gnd.n6775 585
R1248 gnd.n6775 gnd.n6774 585
R1249 gnd.n669 gnd.n668 585
R1250 gnd.n668 gnd.n667 585
R1251 gnd.n6781 gnd.n6780 585
R1252 gnd.n6782 gnd.n6781 585
R1253 gnd.n666 gnd.n665 585
R1254 gnd.n6783 gnd.n666 585
R1255 gnd.n6786 gnd.n6785 585
R1256 gnd.n6785 gnd.n6784 585
R1257 gnd.n663 gnd.n662 585
R1258 gnd.n662 gnd.n661 585
R1259 gnd.n6791 gnd.n6790 585
R1260 gnd.n6792 gnd.n6791 585
R1261 gnd.n660 gnd.n659 585
R1262 gnd.n6793 gnd.n660 585
R1263 gnd.n6796 gnd.n6795 585
R1264 gnd.n6795 gnd.n6794 585
R1265 gnd.n657 gnd.n656 585
R1266 gnd.n656 gnd.n655 585
R1267 gnd.n6801 gnd.n6800 585
R1268 gnd.n6802 gnd.n6801 585
R1269 gnd.n654 gnd.n653 585
R1270 gnd.n6803 gnd.n654 585
R1271 gnd.n6806 gnd.n6805 585
R1272 gnd.n6805 gnd.n6804 585
R1273 gnd.n651 gnd.n650 585
R1274 gnd.n650 gnd.n649 585
R1275 gnd.n6811 gnd.n6810 585
R1276 gnd.n6812 gnd.n6811 585
R1277 gnd.n648 gnd.n647 585
R1278 gnd.n6813 gnd.n648 585
R1279 gnd.n6816 gnd.n6815 585
R1280 gnd.n6815 gnd.n6814 585
R1281 gnd.n645 gnd.n644 585
R1282 gnd.n644 gnd.n643 585
R1283 gnd.n6821 gnd.n6820 585
R1284 gnd.n6822 gnd.n6821 585
R1285 gnd.n642 gnd.n641 585
R1286 gnd.n6823 gnd.n642 585
R1287 gnd.n6826 gnd.n6825 585
R1288 gnd.n6825 gnd.n6824 585
R1289 gnd.n639 gnd.n638 585
R1290 gnd.n638 gnd.n637 585
R1291 gnd.n6831 gnd.n6830 585
R1292 gnd.n6832 gnd.n6831 585
R1293 gnd.n636 gnd.n635 585
R1294 gnd.n6833 gnd.n636 585
R1295 gnd.n6836 gnd.n6835 585
R1296 gnd.n6835 gnd.n6834 585
R1297 gnd.n633 gnd.n632 585
R1298 gnd.n632 gnd.n631 585
R1299 gnd.n6841 gnd.n6840 585
R1300 gnd.n6842 gnd.n6841 585
R1301 gnd.n630 gnd.n629 585
R1302 gnd.n6843 gnd.n630 585
R1303 gnd.n6846 gnd.n6845 585
R1304 gnd.n6845 gnd.n6844 585
R1305 gnd.n627 gnd.n626 585
R1306 gnd.n626 gnd.n625 585
R1307 gnd.n6851 gnd.n6850 585
R1308 gnd.n6852 gnd.n6851 585
R1309 gnd.n624 gnd.n623 585
R1310 gnd.n6853 gnd.n624 585
R1311 gnd.n6856 gnd.n6855 585
R1312 gnd.n6855 gnd.n6854 585
R1313 gnd.n621 gnd.n620 585
R1314 gnd.n620 gnd.n619 585
R1315 gnd.n6861 gnd.n6860 585
R1316 gnd.n6862 gnd.n6861 585
R1317 gnd.n618 gnd.n617 585
R1318 gnd.n6863 gnd.n618 585
R1319 gnd.n6866 gnd.n6865 585
R1320 gnd.n6865 gnd.n6864 585
R1321 gnd.n615 gnd.n614 585
R1322 gnd.n614 gnd.n613 585
R1323 gnd.n6871 gnd.n6870 585
R1324 gnd.n6872 gnd.n6871 585
R1325 gnd.n612 gnd.n611 585
R1326 gnd.n6873 gnd.n612 585
R1327 gnd.n6876 gnd.n6875 585
R1328 gnd.n6875 gnd.n6874 585
R1329 gnd.n609 gnd.n608 585
R1330 gnd.n608 gnd.n607 585
R1331 gnd.n6881 gnd.n6880 585
R1332 gnd.n6882 gnd.n6881 585
R1333 gnd.n606 gnd.n605 585
R1334 gnd.n6883 gnd.n606 585
R1335 gnd.n6886 gnd.n6885 585
R1336 gnd.n6885 gnd.n6884 585
R1337 gnd.n603 gnd.n602 585
R1338 gnd.n602 gnd.n601 585
R1339 gnd.n6891 gnd.n6890 585
R1340 gnd.n6892 gnd.n6891 585
R1341 gnd.n600 gnd.n599 585
R1342 gnd.n6893 gnd.n600 585
R1343 gnd.n6896 gnd.n6895 585
R1344 gnd.n6895 gnd.n6894 585
R1345 gnd.n597 gnd.n596 585
R1346 gnd.n596 gnd.n595 585
R1347 gnd.n6901 gnd.n6900 585
R1348 gnd.n6902 gnd.n6901 585
R1349 gnd.n594 gnd.n593 585
R1350 gnd.n6903 gnd.n594 585
R1351 gnd.n6906 gnd.n6905 585
R1352 gnd.n6905 gnd.n6904 585
R1353 gnd.n591 gnd.n590 585
R1354 gnd.n590 gnd.n589 585
R1355 gnd.n6911 gnd.n6910 585
R1356 gnd.n6912 gnd.n6911 585
R1357 gnd.n588 gnd.n587 585
R1358 gnd.n6913 gnd.n588 585
R1359 gnd.n6916 gnd.n6915 585
R1360 gnd.n6915 gnd.n6914 585
R1361 gnd.n585 gnd.n584 585
R1362 gnd.n584 gnd.n583 585
R1363 gnd.n6921 gnd.n6920 585
R1364 gnd.n6922 gnd.n6921 585
R1365 gnd.n582 gnd.n581 585
R1366 gnd.n6923 gnd.n582 585
R1367 gnd.n6926 gnd.n6925 585
R1368 gnd.n6925 gnd.n6924 585
R1369 gnd.n579 gnd.n578 585
R1370 gnd.n578 gnd.n577 585
R1371 gnd.n6931 gnd.n6930 585
R1372 gnd.n6932 gnd.n6931 585
R1373 gnd.n576 gnd.n575 585
R1374 gnd.n6933 gnd.n576 585
R1375 gnd.n6936 gnd.n6935 585
R1376 gnd.n6935 gnd.n6934 585
R1377 gnd.n573 gnd.n572 585
R1378 gnd.n572 gnd.n571 585
R1379 gnd.n6941 gnd.n6940 585
R1380 gnd.n6942 gnd.n6941 585
R1381 gnd.n570 gnd.n569 585
R1382 gnd.n6943 gnd.n570 585
R1383 gnd.n6946 gnd.n6945 585
R1384 gnd.n6945 gnd.n6944 585
R1385 gnd.n567 gnd.n566 585
R1386 gnd.n566 gnd.n565 585
R1387 gnd.n6951 gnd.n6950 585
R1388 gnd.n6952 gnd.n6951 585
R1389 gnd.n564 gnd.n563 585
R1390 gnd.n6953 gnd.n564 585
R1391 gnd.n6956 gnd.n6955 585
R1392 gnd.n6955 gnd.n6954 585
R1393 gnd.n561 gnd.n560 585
R1394 gnd.n560 gnd.n559 585
R1395 gnd.n6961 gnd.n6960 585
R1396 gnd.n6962 gnd.n6961 585
R1397 gnd.n558 gnd.n557 585
R1398 gnd.n6963 gnd.n558 585
R1399 gnd.n6966 gnd.n6965 585
R1400 gnd.n6965 gnd.n6964 585
R1401 gnd.n555 gnd.n554 585
R1402 gnd.n554 gnd.n553 585
R1403 gnd.n6971 gnd.n6970 585
R1404 gnd.n6972 gnd.n6971 585
R1405 gnd.n552 gnd.n551 585
R1406 gnd.n6973 gnd.n552 585
R1407 gnd.n6976 gnd.n6975 585
R1408 gnd.n6975 gnd.n6974 585
R1409 gnd.n549 gnd.n548 585
R1410 gnd.n548 gnd.n547 585
R1411 gnd.n6981 gnd.n6980 585
R1412 gnd.n6982 gnd.n6981 585
R1413 gnd.n546 gnd.n545 585
R1414 gnd.n6983 gnd.n546 585
R1415 gnd.n6986 gnd.n6985 585
R1416 gnd.n6985 gnd.n6984 585
R1417 gnd.n543 gnd.n542 585
R1418 gnd.n542 gnd.n541 585
R1419 gnd.n6992 gnd.n6991 585
R1420 gnd.n6993 gnd.n6992 585
R1421 gnd.n540 gnd.n539 585
R1422 gnd.n6994 gnd.n540 585
R1423 gnd.n6997 gnd.n6996 585
R1424 gnd.n6996 gnd.n6995 585
R1425 gnd.n6998 gnd.n537 585
R1426 gnd.n537 gnd.n536 585
R1427 gnd.n412 gnd.n411 585
R1428 gnd.n7205 gnd.n411 585
R1429 gnd.n7208 gnd.n7207 585
R1430 gnd.n7207 gnd.n7206 585
R1431 gnd.n415 gnd.n414 585
R1432 gnd.n7204 gnd.n415 585
R1433 gnd.n7202 gnd.n7201 585
R1434 gnd.n7203 gnd.n7202 585
R1435 gnd.n418 gnd.n417 585
R1436 gnd.n417 gnd.n416 585
R1437 gnd.n7197 gnd.n7196 585
R1438 gnd.n7196 gnd.n7195 585
R1439 gnd.n421 gnd.n420 585
R1440 gnd.n7194 gnd.n421 585
R1441 gnd.n7192 gnd.n7191 585
R1442 gnd.n7193 gnd.n7192 585
R1443 gnd.n424 gnd.n423 585
R1444 gnd.n423 gnd.n422 585
R1445 gnd.n7187 gnd.n7186 585
R1446 gnd.n7186 gnd.n7185 585
R1447 gnd.n427 gnd.n426 585
R1448 gnd.n7184 gnd.n427 585
R1449 gnd.n7182 gnd.n7181 585
R1450 gnd.n7183 gnd.n7182 585
R1451 gnd.n430 gnd.n429 585
R1452 gnd.n429 gnd.n428 585
R1453 gnd.n7177 gnd.n7176 585
R1454 gnd.n7176 gnd.n7175 585
R1455 gnd.n433 gnd.n432 585
R1456 gnd.n7174 gnd.n433 585
R1457 gnd.n7172 gnd.n7171 585
R1458 gnd.n7173 gnd.n7172 585
R1459 gnd.n436 gnd.n435 585
R1460 gnd.n435 gnd.n434 585
R1461 gnd.n7167 gnd.n7166 585
R1462 gnd.n7166 gnd.n7165 585
R1463 gnd.n439 gnd.n438 585
R1464 gnd.n7164 gnd.n439 585
R1465 gnd.n7162 gnd.n7161 585
R1466 gnd.n7163 gnd.n7162 585
R1467 gnd.n442 gnd.n441 585
R1468 gnd.n441 gnd.n440 585
R1469 gnd.n7157 gnd.n7156 585
R1470 gnd.n7156 gnd.n7155 585
R1471 gnd.n445 gnd.n444 585
R1472 gnd.n7154 gnd.n445 585
R1473 gnd.n7152 gnd.n7151 585
R1474 gnd.n7153 gnd.n7152 585
R1475 gnd.n448 gnd.n447 585
R1476 gnd.n447 gnd.n446 585
R1477 gnd.n7147 gnd.n7146 585
R1478 gnd.n7146 gnd.n7145 585
R1479 gnd.n451 gnd.n450 585
R1480 gnd.n7144 gnd.n451 585
R1481 gnd.n7142 gnd.n7141 585
R1482 gnd.n7143 gnd.n7142 585
R1483 gnd.n454 gnd.n453 585
R1484 gnd.n453 gnd.n452 585
R1485 gnd.n7137 gnd.n7136 585
R1486 gnd.n7136 gnd.n7135 585
R1487 gnd.n457 gnd.n456 585
R1488 gnd.n7134 gnd.n457 585
R1489 gnd.n7132 gnd.n7131 585
R1490 gnd.n7133 gnd.n7132 585
R1491 gnd.n460 gnd.n459 585
R1492 gnd.n459 gnd.n458 585
R1493 gnd.n7127 gnd.n7126 585
R1494 gnd.n7126 gnd.n7125 585
R1495 gnd.n463 gnd.n462 585
R1496 gnd.n7124 gnd.n463 585
R1497 gnd.n7122 gnd.n7121 585
R1498 gnd.n7123 gnd.n7122 585
R1499 gnd.n466 gnd.n465 585
R1500 gnd.n465 gnd.n464 585
R1501 gnd.n7117 gnd.n7116 585
R1502 gnd.n7116 gnd.n7115 585
R1503 gnd.n469 gnd.n468 585
R1504 gnd.n7114 gnd.n469 585
R1505 gnd.n7112 gnd.n7111 585
R1506 gnd.n7113 gnd.n7112 585
R1507 gnd.n472 gnd.n471 585
R1508 gnd.n471 gnd.n470 585
R1509 gnd.n7107 gnd.n7106 585
R1510 gnd.n7106 gnd.n7105 585
R1511 gnd.n475 gnd.n474 585
R1512 gnd.n7104 gnd.n475 585
R1513 gnd.n7102 gnd.n7101 585
R1514 gnd.n7103 gnd.n7102 585
R1515 gnd.n478 gnd.n477 585
R1516 gnd.n477 gnd.n476 585
R1517 gnd.n7097 gnd.n7096 585
R1518 gnd.n7096 gnd.n7095 585
R1519 gnd.n481 gnd.n480 585
R1520 gnd.n7094 gnd.n481 585
R1521 gnd.n7092 gnd.n7091 585
R1522 gnd.n7093 gnd.n7092 585
R1523 gnd.n484 gnd.n483 585
R1524 gnd.n483 gnd.n482 585
R1525 gnd.n7087 gnd.n7086 585
R1526 gnd.n7086 gnd.n7085 585
R1527 gnd.n487 gnd.n486 585
R1528 gnd.n7084 gnd.n487 585
R1529 gnd.n7082 gnd.n7081 585
R1530 gnd.n7083 gnd.n7082 585
R1531 gnd.n490 gnd.n489 585
R1532 gnd.n489 gnd.n488 585
R1533 gnd.n7077 gnd.n7076 585
R1534 gnd.n7076 gnd.n7075 585
R1535 gnd.n493 gnd.n492 585
R1536 gnd.n7074 gnd.n493 585
R1537 gnd.n7072 gnd.n7071 585
R1538 gnd.n7073 gnd.n7072 585
R1539 gnd.n496 gnd.n495 585
R1540 gnd.n495 gnd.n494 585
R1541 gnd.n7067 gnd.n7066 585
R1542 gnd.n7066 gnd.n7065 585
R1543 gnd.n499 gnd.n498 585
R1544 gnd.n7064 gnd.n499 585
R1545 gnd.n7062 gnd.n7061 585
R1546 gnd.n7063 gnd.n7062 585
R1547 gnd.n502 gnd.n501 585
R1548 gnd.n501 gnd.n500 585
R1549 gnd.n7057 gnd.n7056 585
R1550 gnd.n7056 gnd.n7055 585
R1551 gnd.n505 gnd.n504 585
R1552 gnd.n7054 gnd.n505 585
R1553 gnd.n7052 gnd.n7051 585
R1554 gnd.n7053 gnd.n7052 585
R1555 gnd.n508 gnd.n507 585
R1556 gnd.n507 gnd.n506 585
R1557 gnd.n7047 gnd.n7046 585
R1558 gnd.n7046 gnd.n7045 585
R1559 gnd.n511 gnd.n510 585
R1560 gnd.n7044 gnd.n511 585
R1561 gnd.n7042 gnd.n7041 585
R1562 gnd.n7043 gnd.n7042 585
R1563 gnd.n514 gnd.n513 585
R1564 gnd.n513 gnd.n512 585
R1565 gnd.n7037 gnd.n7036 585
R1566 gnd.n7036 gnd.n7035 585
R1567 gnd.n517 gnd.n516 585
R1568 gnd.n7034 gnd.n517 585
R1569 gnd.n7032 gnd.n7031 585
R1570 gnd.n7033 gnd.n7032 585
R1571 gnd.n520 gnd.n519 585
R1572 gnd.n519 gnd.n518 585
R1573 gnd.n7027 gnd.n7026 585
R1574 gnd.n7026 gnd.n7025 585
R1575 gnd.n523 gnd.n522 585
R1576 gnd.n7024 gnd.n523 585
R1577 gnd.n7022 gnd.n7021 585
R1578 gnd.n7023 gnd.n7022 585
R1579 gnd.n526 gnd.n525 585
R1580 gnd.n525 gnd.n524 585
R1581 gnd.n7017 gnd.n7016 585
R1582 gnd.n7016 gnd.n7015 585
R1583 gnd.n529 gnd.n528 585
R1584 gnd.n7014 gnd.n529 585
R1585 gnd.n7012 gnd.n7011 585
R1586 gnd.n7013 gnd.n7012 585
R1587 gnd.n532 gnd.n531 585
R1588 gnd.n531 gnd.n530 585
R1589 gnd.n7007 gnd.n7006 585
R1590 gnd.n7006 gnd.n7005 585
R1591 gnd.n535 gnd.n534 585
R1592 gnd.n7004 gnd.n535 585
R1593 gnd.n7002 gnd.n7001 585
R1594 gnd.n7003 gnd.n7002 585
R1595 gnd.n6047 gnd.n6046 585
R1596 gnd.n6048 gnd.n6047 585
R1597 gnd.n2622 gnd.n2621 585
R1598 gnd.n6041 gnd.n2622 585
R1599 gnd.n6056 gnd.n6055 585
R1600 gnd.n6055 gnd.n6054 585
R1601 gnd.n6057 gnd.n2617 585
R1602 gnd.n4352 gnd.n2617 585
R1603 gnd.n6059 gnd.n6058 585
R1604 gnd.n6060 gnd.n6059 585
R1605 gnd.n2602 gnd.n2601 585
R1606 gnd.n4346 gnd.n2602 585
R1607 gnd.n6068 gnd.n6067 585
R1608 gnd.n6067 gnd.n6066 585
R1609 gnd.n6069 gnd.n2597 585
R1610 gnd.n4363 gnd.n2597 585
R1611 gnd.n6071 gnd.n6070 585
R1612 gnd.n6072 gnd.n6071 585
R1613 gnd.n2581 gnd.n2580 585
R1614 gnd.n4339 gnd.n2581 585
R1615 gnd.n6080 gnd.n6079 585
R1616 gnd.n6079 gnd.n6078 585
R1617 gnd.n6081 gnd.n2576 585
R1618 gnd.n4331 gnd.n2576 585
R1619 gnd.n6083 gnd.n6082 585
R1620 gnd.n6084 gnd.n6083 585
R1621 gnd.n2563 gnd.n2562 585
R1622 gnd.n4325 gnd.n2563 585
R1623 gnd.n6092 gnd.n6091 585
R1624 gnd.n6091 gnd.n6090 585
R1625 gnd.n6093 gnd.n2557 585
R1626 gnd.n4317 gnd.n2557 585
R1627 gnd.n6095 gnd.n6094 585
R1628 gnd.n6096 gnd.n6095 585
R1629 gnd.n2558 gnd.n2556 585
R1630 gnd.n4289 gnd.n2556 585
R1631 gnd.n4271 gnd.n4270 585
R1632 gnd.n4270 gnd.n4022 585
R1633 gnd.n4272 gnd.n4032 585
R1634 gnd.n4281 gnd.n4032 585
R1635 gnd.n4274 gnd.n4273 585
R1636 gnd.n4275 gnd.n4274 585
R1637 gnd.n4039 gnd.n4038 585
R1638 gnd.n4259 gnd.n4038 585
R1639 gnd.n4247 gnd.n4246 585
R1640 gnd.n4248 gnd.n4247 585
R1641 gnd.n4057 gnd.n4055 585
R1642 gnd.n4251 gnd.n4055 585
R1643 gnd.n2536 gnd.n2535 585
R1644 gnd.n4240 gnd.n2536 585
R1645 gnd.n6106 gnd.n6105 585
R1646 gnd.n6105 gnd.n6104 585
R1647 gnd.n6107 gnd.n2531 585
R1648 gnd.n4189 gnd.n2531 585
R1649 gnd.n6109 gnd.n6108 585
R1650 gnd.n6110 gnd.n6109 585
R1651 gnd.n2515 gnd.n2514 585
R1652 gnd.n4195 gnd.n2515 585
R1653 gnd.n6118 gnd.n6117 585
R1654 gnd.n6117 gnd.n6116 585
R1655 gnd.n6119 gnd.n2510 585
R1656 gnd.n4201 gnd.n2510 585
R1657 gnd.n6121 gnd.n6120 585
R1658 gnd.n6122 gnd.n6121 585
R1659 gnd.n2495 gnd.n2494 585
R1660 gnd.n4207 gnd.n2495 585
R1661 gnd.n6130 gnd.n6129 585
R1662 gnd.n6129 gnd.n6128 585
R1663 gnd.n6131 gnd.n2490 585
R1664 gnd.n4172 gnd.n2490 585
R1665 gnd.n6133 gnd.n6132 585
R1666 gnd.n6134 gnd.n6133 585
R1667 gnd.n2476 gnd.n2475 585
R1668 gnd.n2479 gnd.n2476 585
R1669 gnd.n6142 gnd.n6141 585
R1670 gnd.n6141 gnd.n6140 585
R1671 gnd.n6143 gnd.n2469 585
R1672 gnd.n2469 gnd.n2467 585
R1673 gnd.n6145 gnd.n6144 585
R1674 gnd.n6146 gnd.n6145 585
R1675 gnd.n2471 gnd.n2468 585
R1676 gnd.n2468 gnd.n2464 585
R1677 gnd.n2470 gnd.n2455 585
R1678 gnd.n6152 gnd.n2455 585
R1679 gnd.n4108 gnd.n2449 585
R1680 gnd.n4108 gnd.n2380 585
R1681 gnd.n4110 gnd.n4109 585
R1682 gnd.n4112 gnd.n4111 585
R1683 gnd.n4114 gnd.n4113 585
R1684 gnd.n4118 gnd.n4106 585
R1685 gnd.n4120 gnd.n4119 585
R1686 gnd.n4122 gnd.n4121 585
R1687 gnd.n4124 gnd.n4123 585
R1688 gnd.n4128 gnd.n4104 585
R1689 gnd.n4130 gnd.n4129 585
R1690 gnd.n4132 gnd.n4131 585
R1691 gnd.n4134 gnd.n4133 585
R1692 gnd.n4138 gnd.n4102 585
R1693 gnd.n4140 gnd.n4139 585
R1694 gnd.n4142 gnd.n4141 585
R1695 gnd.n4144 gnd.n4143 585
R1696 gnd.n4099 gnd.n4098 585
R1697 gnd.n4148 gnd.n4100 585
R1698 gnd.n4149 gnd.n4095 585
R1699 gnd.n4150 gnd.n2379 585
R1700 gnd.n6276 gnd.n2379 585
R1701 gnd.n5968 gnd.n5967 585
R1702 gnd.n5969 gnd.n2737 585
R1703 gnd.n5970 gnd.n2732 585
R1704 gnd.n2750 gnd.n2721 585
R1705 gnd.n5977 gnd.n2720 585
R1706 gnd.n5978 gnd.n2719 585
R1707 gnd.n2747 gnd.n2713 585
R1708 gnd.n5985 gnd.n2712 585
R1709 gnd.n5986 gnd.n2711 585
R1710 gnd.n2745 gnd.n2703 585
R1711 gnd.n5993 gnd.n2702 585
R1712 gnd.n5994 gnd.n2701 585
R1713 gnd.n2742 gnd.n2695 585
R1714 gnd.n6001 gnd.n2694 585
R1715 gnd.n6002 gnd.n2693 585
R1716 gnd.n2740 gnd.n2685 585
R1717 gnd.n6009 gnd.n2684 585
R1718 gnd.n6010 gnd.n2683 585
R1719 gnd.n2682 gnd.n2636 585
R1720 gnd.n5965 gnd.n2636 585
R1721 gnd.n2642 gnd.n2634 585
R1722 gnd.n6048 gnd.n2634 585
R1723 gnd.n6040 gnd.n6039 585
R1724 gnd.n6041 gnd.n6040 585
R1725 gnd.n2641 gnd.n2625 585
R1726 gnd.n6054 gnd.n2625 585
R1727 gnd.n4355 gnd.n4353 585
R1728 gnd.n4353 gnd.n4352 585
R1729 gnd.n4356 gnd.n2615 585
R1730 gnd.n6060 gnd.n2615 585
R1731 gnd.n4357 gnd.n4004 585
R1732 gnd.n4346 gnd.n4004 585
R1733 gnd.n4001 gnd.n2604 585
R1734 gnd.n6066 gnd.n2604 585
R1735 gnd.n4362 gnd.n4361 585
R1736 gnd.n4363 gnd.n4362 585
R1737 gnd.n4000 gnd.n2595 585
R1738 gnd.n6072 gnd.n2595 585
R1739 gnd.n4338 gnd.n4337 585
R1740 gnd.n4339 gnd.n4338 585
R1741 gnd.n4007 gnd.n2584 585
R1742 gnd.n6078 gnd.n2584 585
R1743 gnd.n4333 gnd.n4332 585
R1744 gnd.n4332 gnd.n4331 585
R1745 gnd.n4009 gnd.n2575 585
R1746 gnd.n6084 gnd.n2575 585
R1747 gnd.n4324 gnd.n4323 585
R1748 gnd.n4325 gnd.n4324 585
R1749 gnd.n4013 gnd.n2565 585
R1750 gnd.n6090 gnd.n2565 585
R1751 gnd.n4319 gnd.n4318 585
R1752 gnd.n4318 gnd.n4317 585
R1753 gnd.n4015 gnd.n2554 585
R1754 gnd.n6096 gnd.n2554 585
R1755 gnd.n4288 gnd.n4287 585
R1756 gnd.n4289 gnd.n4288 585
R1757 gnd.n4025 gnd.n4024 585
R1758 gnd.n4024 gnd.n4022 585
R1759 gnd.n4283 gnd.n4282 585
R1760 gnd.n4282 gnd.n4281 585
R1761 gnd.n4028 gnd.n4027 585
R1762 gnd.n4275 gnd.n4028 585
R1763 gnd.n4258 gnd.n4257 585
R1764 gnd.n4259 gnd.n4258 585
R1765 gnd.n4048 gnd.n4047 585
R1766 gnd.n4248 gnd.n4047 585
R1767 gnd.n4253 gnd.n4252 585
R1768 gnd.n4252 gnd.n4251 585
R1769 gnd.n4051 gnd.n4050 585
R1770 gnd.n4240 gnd.n4051 585
R1771 gnd.n4186 gnd.n2539 585
R1772 gnd.n6104 gnd.n2539 585
R1773 gnd.n4191 gnd.n4190 585
R1774 gnd.n4190 gnd.n4189 585
R1775 gnd.n4192 gnd.n2529 585
R1776 gnd.n6110 gnd.n2529 585
R1777 gnd.n4194 gnd.n4193 585
R1778 gnd.n4195 gnd.n4194 585
R1779 gnd.n4079 gnd.n2518 585
R1780 gnd.n6116 gnd.n2518 585
R1781 gnd.n4203 gnd.n4202 585
R1782 gnd.n4202 gnd.n4201 585
R1783 gnd.n4204 gnd.n2508 585
R1784 gnd.n6122 gnd.n2508 585
R1785 gnd.n4206 gnd.n4205 585
R1786 gnd.n4207 gnd.n4206 585
R1787 gnd.n4075 gnd.n2498 585
R1788 gnd.n6128 gnd.n2498 585
R1789 gnd.n4171 gnd.n4170 585
R1790 gnd.n4172 gnd.n4171 585
R1791 gnd.n4090 gnd.n2488 585
R1792 gnd.n6134 gnd.n2488 585
R1793 gnd.n4165 gnd.n4164 585
R1794 gnd.n4164 gnd.n2479 585
R1795 gnd.n4163 gnd.n2478 585
R1796 gnd.n6140 gnd.n2478 585
R1797 gnd.n4162 gnd.n4161 585
R1798 gnd.n4161 gnd.n2467 585
R1799 gnd.n4092 gnd.n2466 585
R1800 gnd.n6146 gnd.n2466 585
R1801 gnd.n4157 gnd.n4156 585
R1802 gnd.n4156 gnd.n2464 585
R1803 gnd.n4155 gnd.n2454 585
R1804 gnd.n6152 gnd.n2454 585
R1805 gnd.n4154 gnd.n4153 585
R1806 gnd.n4153 gnd.n2380 585
R1807 gnd.n6338 gnd.n6337 585
R1808 gnd.n6339 gnd.n6338 585
R1809 gnd.n1046 gnd.n1044 585
R1810 gnd.n1044 gnd.n1040 585
R1811 gnd.n1026 gnd.n1025 585
R1812 gnd.n2332 gnd.n1026 585
R1813 gnd.n6349 gnd.n6348 585
R1814 gnd.n6348 gnd.n6347 585
R1815 gnd.n6350 gnd.n1020 585
R1816 gnd.n1989 gnd.n1020 585
R1817 gnd.n6352 gnd.n6351 585
R1818 gnd.n6353 gnd.n6352 585
R1819 gnd.n1021 gnd.n1019 585
R1820 gnd.n1019 gnd.n1015 585
R1821 gnd.n1000 gnd.n999 585
R1822 gnd.n1004 gnd.n1000 585
R1823 gnd.n6363 gnd.n6362 585
R1824 gnd.n6362 gnd.n6361 585
R1825 gnd.n6364 gnd.n994 585
R1826 gnd.n1998 gnd.n994 585
R1827 gnd.n6366 gnd.n6365 585
R1828 gnd.n6367 gnd.n6366 585
R1829 gnd.n995 gnd.n993 585
R1830 gnd.n993 gnd.n989 585
R1831 gnd.n2043 gnd.n2042 585
R1832 gnd.n2042 gnd.n980 585
R1833 gnd.n2041 gnd.n1158 585
R1834 gnd.n2041 gnd.n978 585
R1835 gnd.n2040 gnd.n1160 585
R1836 gnd.n2040 gnd.n2039 585
R1837 gnd.n2029 gnd.n1159 585
R1838 gnd.n1171 gnd.n1159 585
R1839 gnd.n2028 gnd.n2027 585
R1840 gnd.n2027 gnd.n2026 585
R1841 gnd.n1167 gnd.n1165 585
R1842 gnd.n2013 gnd.n1167 585
R1843 gnd.n1963 gnd.n1188 585
R1844 gnd.n1188 gnd.n1179 585
R1845 gnd.n1965 gnd.n1964 585
R1846 gnd.n1966 gnd.n1965 585
R1847 gnd.n1189 gnd.n1187 585
R1848 gnd.n1195 gnd.n1187 585
R1849 gnd.n1942 gnd.n1941 585
R1850 gnd.n1943 gnd.n1942 585
R1851 gnd.n1206 gnd.n1205 585
R1852 gnd.n1205 gnd.n1201 585
R1853 gnd.n1932 gnd.n1931 585
R1854 gnd.n1933 gnd.n1932 585
R1855 gnd.n1217 gnd.n1216 585
R1856 gnd.n1221 gnd.n1216 585
R1857 gnd.n1910 gnd.n1233 585
R1858 gnd.n1575 gnd.n1233 585
R1859 gnd.n1912 gnd.n1911 585
R1860 gnd.n1913 gnd.n1912 585
R1861 gnd.n1234 gnd.n1232 585
R1862 gnd.n1232 gnd.n1228 585
R1863 gnd.n1901 gnd.n1900 585
R1864 gnd.n1902 gnd.n1901 585
R1865 gnd.n1242 gnd.n1241 585
R1866 gnd.n1583 gnd.n1241 585
R1867 gnd.n1879 gnd.n1258 585
R1868 gnd.n1258 gnd.n1246 585
R1869 gnd.n1881 gnd.n1880 585
R1870 gnd.n1882 gnd.n1881 585
R1871 gnd.n1259 gnd.n1257 585
R1872 gnd.n1257 gnd.n1253 585
R1873 gnd.n1870 gnd.n1869 585
R1874 gnd.n1871 gnd.n1870 585
R1875 gnd.n1267 gnd.n1266 585
R1876 gnd.n1272 gnd.n1266 585
R1877 gnd.n1848 gnd.n1284 585
R1878 gnd.n1284 gnd.n1271 585
R1879 gnd.n1850 gnd.n1849 585
R1880 gnd.n1851 gnd.n1850 585
R1881 gnd.n1285 gnd.n1283 585
R1882 gnd.n1283 gnd.n1279 585
R1883 gnd.n1839 gnd.n1838 585
R1884 gnd.n1840 gnd.n1839 585
R1885 gnd.n1292 gnd.n1291 585
R1886 gnd.n1297 gnd.n1291 585
R1887 gnd.n1817 gnd.n1310 585
R1888 gnd.n1310 gnd.n1296 585
R1889 gnd.n1819 gnd.n1818 585
R1890 gnd.n1820 gnd.n1819 585
R1891 gnd.n1311 gnd.n1309 585
R1892 gnd.n1309 gnd.n1305 585
R1893 gnd.n1808 gnd.n1807 585
R1894 gnd.n1809 gnd.n1808 585
R1895 gnd.n1318 gnd.n1317 585
R1896 gnd.n1323 gnd.n1317 585
R1897 gnd.n1786 gnd.n1336 585
R1898 gnd.n1336 gnd.n1322 585
R1899 gnd.n1788 gnd.n1787 585
R1900 gnd.n1789 gnd.n1788 585
R1901 gnd.n1337 gnd.n1335 585
R1902 gnd.n1335 gnd.n1331 585
R1903 gnd.n1777 gnd.n1776 585
R1904 gnd.n1778 gnd.n1777 585
R1905 gnd.n1345 gnd.n1344 585
R1906 gnd.n1667 gnd.n1344 585
R1907 gnd.n1755 gnd.n1361 585
R1908 gnd.n1361 gnd.n1349 585
R1909 gnd.n1757 gnd.n1756 585
R1910 gnd.n1758 gnd.n1757 585
R1911 gnd.n1362 gnd.n1360 585
R1912 gnd.n1360 gnd.n1356 585
R1913 gnd.n1746 gnd.n1745 585
R1914 gnd.n1747 gnd.n1746 585
R1915 gnd.n1369 gnd.n1368 585
R1916 gnd.n1368 gnd.n1366 585
R1917 gnd.n1740 gnd.n1739 585
R1918 gnd.n1739 gnd.n1738 585
R1919 gnd.n1373 gnd.n1372 585
R1920 gnd.n1381 gnd.n1373 585
R1921 gnd.n1534 gnd.n1533 585
R1922 gnd.n1535 gnd.n1534 585
R1923 gnd.n1383 gnd.n1382 585
R1924 gnd.n1382 gnd.n1380 585
R1925 gnd.n1529 gnd.n1528 585
R1926 gnd.n1528 gnd.n1527 585
R1927 gnd.n1386 gnd.n1385 585
R1928 gnd.n1387 gnd.n1386 585
R1929 gnd.n1518 gnd.n1517 585
R1930 gnd.n1519 gnd.n1518 585
R1931 gnd.n1395 gnd.n1394 585
R1932 gnd.n1394 gnd.n1393 585
R1933 gnd.n1513 gnd.n1512 585
R1934 gnd.n1512 gnd.n1511 585
R1935 gnd.n1398 gnd.n1397 585
R1936 gnd.n1399 gnd.n1398 585
R1937 gnd.n1502 gnd.n1501 585
R1938 gnd.n1503 gnd.n1502 585
R1939 gnd.n1498 gnd.n1405 585
R1940 gnd.n1497 gnd.n1496 585
R1941 gnd.n1494 gnd.n1407 585
R1942 gnd.n1494 gnd.n1404 585
R1943 gnd.n1493 gnd.n1492 585
R1944 gnd.n1491 gnd.n1490 585
R1945 gnd.n1489 gnd.n1412 585
R1946 gnd.n1487 gnd.n1486 585
R1947 gnd.n1485 gnd.n1413 585
R1948 gnd.n1484 gnd.n1483 585
R1949 gnd.n1481 gnd.n1418 585
R1950 gnd.n1479 gnd.n1478 585
R1951 gnd.n1477 gnd.n1419 585
R1952 gnd.n1476 gnd.n1475 585
R1953 gnd.n1473 gnd.n1424 585
R1954 gnd.n1471 gnd.n1470 585
R1955 gnd.n1469 gnd.n1425 585
R1956 gnd.n1468 gnd.n1467 585
R1957 gnd.n1465 gnd.n1430 585
R1958 gnd.n1463 gnd.n1462 585
R1959 gnd.n1461 gnd.n1431 585
R1960 gnd.n1460 gnd.n1459 585
R1961 gnd.n1457 gnd.n1436 585
R1962 gnd.n1455 gnd.n1454 585
R1963 gnd.n1452 gnd.n1437 585
R1964 gnd.n1451 gnd.n1450 585
R1965 gnd.n1448 gnd.n1446 585
R1966 gnd.n1444 gnd.n1403 585
R1967 gnd.n2340 gnd.n2339 585
R1968 gnd.n1070 gnd.n1069 585
R1969 gnd.n1146 gnd.n1145 585
R1970 gnd.n1144 gnd.n1143 585
R1971 gnd.n1142 gnd.n1141 585
R1972 gnd.n1135 gnd.n1075 585
R1973 gnd.n1137 gnd.n1136 585
R1974 gnd.n1134 gnd.n1133 585
R1975 gnd.n1132 gnd.n1131 585
R1976 gnd.n1125 gnd.n1077 585
R1977 gnd.n1127 gnd.n1126 585
R1978 gnd.n1124 gnd.n1123 585
R1979 gnd.n1122 gnd.n1121 585
R1980 gnd.n1115 gnd.n1079 585
R1981 gnd.n1117 gnd.n1116 585
R1982 gnd.n1114 gnd.n1113 585
R1983 gnd.n1112 gnd.n1111 585
R1984 gnd.n1105 gnd.n1081 585
R1985 gnd.n1107 gnd.n1106 585
R1986 gnd.n1104 gnd.n1103 585
R1987 gnd.n1102 gnd.n1101 585
R1988 gnd.n1095 gnd.n1083 585
R1989 gnd.n1097 gnd.n1096 585
R1990 gnd.n1094 gnd.n1093 585
R1991 gnd.n1092 gnd.n1091 585
R1992 gnd.n1086 gnd.n1085 585
R1993 gnd.n1087 gnd.n1045 585
R1994 gnd.n6323 gnd.n1045 585
R1995 gnd.n2336 gnd.n1042 585
R1996 gnd.n6339 gnd.n1042 585
R1997 gnd.n2335 gnd.n2334 585
R1998 gnd.n2334 gnd.n1040 585
R1999 gnd.n2333 gnd.n1150 585
R2000 gnd.n2333 gnd.n2332 585
R2001 gnd.n1988 gnd.n1028 585
R2002 gnd.n6347 gnd.n1028 585
R2003 gnd.n1991 gnd.n1990 585
R2004 gnd.n1990 gnd.n1989 585
R2005 gnd.n1992 gnd.n1017 585
R2006 gnd.n6353 gnd.n1017 585
R2007 gnd.n1994 gnd.n1993 585
R2008 gnd.n1994 gnd.n1015 585
R2009 gnd.n1996 gnd.n1995 585
R2010 gnd.n1995 gnd.n1004 585
R2011 gnd.n1997 gnd.n1002 585
R2012 gnd.n6361 gnd.n1002 585
R2013 gnd.n2000 gnd.n1999 585
R2014 gnd.n1999 gnd.n1998 585
R2015 gnd.n2001 gnd.n991 585
R2016 gnd.n6367 gnd.n991 585
R2017 gnd.n2003 gnd.n2002 585
R2018 gnd.n2003 gnd.n989 585
R2019 gnd.n2004 gnd.n1976 585
R2020 gnd.n2004 gnd.n980 585
R2021 gnd.n2006 gnd.n2005 585
R2022 gnd.n2005 gnd.n978 585
R2023 gnd.n2007 gnd.n1161 585
R2024 gnd.n2039 gnd.n1161 585
R2025 gnd.n2009 gnd.n2008 585
R2026 gnd.n2008 gnd.n1171 585
R2027 gnd.n2010 gnd.n1169 585
R2028 gnd.n2026 gnd.n1169 585
R2029 gnd.n2012 gnd.n2011 585
R2030 gnd.n2013 gnd.n2012 585
R2031 gnd.n1182 gnd.n1181 585
R2032 gnd.n1181 gnd.n1179 585
R2033 gnd.n1968 gnd.n1967 585
R2034 gnd.n1967 gnd.n1966 585
R2035 gnd.n1185 gnd.n1184 585
R2036 gnd.n1195 gnd.n1185 585
R2037 gnd.n1569 gnd.n1203 585
R2038 gnd.n1943 gnd.n1203 585
R2039 gnd.n1571 gnd.n1570 585
R2040 gnd.n1570 gnd.n1201 585
R2041 gnd.n1572 gnd.n1215 585
R2042 gnd.n1933 gnd.n1215 585
R2043 gnd.n1574 gnd.n1573 585
R2044 gnd.n1574 gnd.n1221 585
R2045 gnd.n1577 gnd.n1576 585
R2046 gnd.n1576 gnd.n1575 585
R2047 gnd.n1578 gnd.n1230 585
R2048 gnd.n1913 gnd.n1230 585
R2049 gnd.n1580 gnd.n1579 585
R2050 gnd.n1579 gnd.n1228 585
R2051 gnd.n1581 gnd.n1240 585
R2052 gnd.n1902 gnd.n1240 585
R2053 gnd.n1584 gnd.n1582 585
R2054 gnd.n1584 gnd.n1583 585
R2055 gnd.n1586 gnd.n1585 585
R2056 gnd.n1585 gnd.n1246 585
R2057 gnd.n1587 gnd.n1255 585
R2058 gnd.n1882 gnd.n1255 585
R2059 gnd.n1590 gnd.n1589 585
R2060 gnd.n1589 gnd.n1253 585
R2061 gnd.n1591 gnd.n1265 585
R2062 gnd.n1871 gnd.n1265 585
R2063 gnd.n1594 gnd.n1593 585
R2064 gnd.n1593 gnd.n1272 585
R2065 gnd.n1592 gnd.n1559 585
R2066 gnd.n1592 gnd.n1271 585
R2067 gnd.n1646 gnd.n1281 585
R2068 gnd.n1851 gnd.n1281 585
R2069 gnd.n1648 gnd.n1647 585
R2070 gnd.n1647 gnd.n1279 585
R2071 gnd.n1649 gnd.n1290 585
R2072 gnd.n1840 gnd.n1290 585
R2073 gnd.n1651 gnd.n1650 585
R2074 gnd.n1651 gnd.n1297 585
R2075 gnd.n1653 gnd.n1652 585
R2076 gnd.n1652 gnd.n1296 585
R2077 gnd.n1654 gnd.n1307 585
R2078 gnd.n1820 gnd.n1307 585
R2079 gnd.n1656 gnd.n1655 585
R2080 gnd.n1655 gnd.n1305 585
R2081 gnd.n1657 gnd.n1316 585
R2082 gnd.n1809 gnd.n1316 585
R2083 gnd.n1659 gnd.n1658 585
R2084 gnd.n1659 gnd.n1323 585
R2085 gnd.n1661 gnd.n1660 585
R2086 gnd.n1660 gnd.n1322 585
R2087 gnd.n1662 gnd.n1333 585
R2088 gnd.n1789 gnd.n1333 585
R2089 gnd.n1664 gnd.n1663 585
R2090 gnd.n1663 gnd.n1331 585
R2091 gnd.n1665 gnd.n1343 585
R2092 gnd.n1778 gnd.n1343 585
R2093 gnd.n1668 gnd.n1666 585
R2094 gnd.n1668 gnd.n1667 585
R2095 gnd.n1670 gnd.n1669 585
R2096 gnd.n1669 gnd.n1349 585
R2097 gnd.n1671 gnd.n1358 585
R2098 gnd.n1758 gnd.n1358 585
R2099 gnd.n1673 gnd.n1672 585
R2100 gnd.n1672 gnd.n1356 585
R2101 gnd.n1674 gnd.n1367 585
R2102 gnd.n1747 gnd.n1367 585
R2103 gnd.n1675 gnd.n1375 585
R2104 gnd.n1375 gnd.n1366 585
R2105 gnd.n1677 gnd.n1676 585
R2106 gnd.n1738 gnd.n1677 585
R2107 gnd.n1376 gnd.n1374 585
R2108 gnd.n1381 gnd.n1374 585
R2109 gnd.n1537 gnd.n1536 585
R2110 gnd.n1536 gnd.n1535 585
R2111 gnd.n1379 gnd.n1378 585
R2112 gnd.n1380 gnd.n1379 585
R2113 gnd.n1526 gnd.n1525 585
R2114 gnd.n1527 gnd.n1526 585
R2115 gnd.n1389 gnd.n1388 585
R2116 gnd.n1388 gnd.n1387 585
R2117 gnd.n1521 gnd.n1520 585
R2118 gnd.n1520 gnd.n1519 585
R2119 gnd.n1392 gnd.n1391 585
R2120 gnd.n1393 gnd.n1392 585
R2121 gnd.n1510 gnd.n1509 585
R2122 gnd.n1511 gnd.n1510 585
R2123 gnd.n1401 gnd.n1400 585
R2124 gnd.n1400 gnd.n1399 585
R2125 gnd.n1505 gnd.n1504 585
R2126 gnd.n1504 gnd.n1503 585
R2127 gnd.n7356 gnd.n7355 585
R2128 gnd.n7357 gnd.n7356 585
R2129 gnd.n159 gnd.n158 585
R2130 gnd.n168 gnd.n159 585
R2131 gnd.n7365 gnd.n7364 585
R2132 gnd.n7364 gnd.n7363 585
R2133 gnd.n7366 gnd.n154 585
R2134 gnd.n154 gnd.n153 585
R2135 gnd.n7368 gnd.n7367 585
R2136 gnd.n7369 gnd.n7368 585
R2137 gnd.n140 gnd.n139 585
R2138 gnd.n143 gnd.n140 585
R2139 gnd.n7377 gnd.n7376 585
R2140 gnd.n7376 gnd.n7375 585
R2141 gnd.n7378 gnd.n135 585
R2142 gnd.n7340 gnd.n135 585
R2143 gnd.n7380 gnd.n7379 585
R2144 gnd.n7381 gnd.n7380 585
R2145 gnd.n119 gnd.n118 585
R2146 gnd.n7248 gnd.n119 585
R2147 gnd.n7389 gnd.n7388 585
R2148 gnd.n7388 gnd.n7387 585
R2149 gnd.n7390 gnd.n114 585
R2150 gnd.n7241 gnd.n114 585
R2151 gnd.n7392 gnd.n7391 585
R2152 gnd.n7393 gnd.n7392 585
R2153 gnd.n101 gnd.n100 585
R2154 gnd.n7233 gnd.n101 585
R2155 gnd.n7401 gnd.n7400 585
R2156 gnd.n7400 gnd.n7399 585
R2157 gnd.n7402 gnd.n95 585
R2158 gnd.n7226 gnd.n95 585
R2159 gnd.n7404 gnd.n7403 585
R2160 gnd.n7405 gnd.n7404 585
R2161 gnd.n96 gnd.n94 585
R2162 gnd.n5442 gnd.n94 585
R2163 gnd.n5454 gnd.n5453 585
R2164 gnd.n5453 gnd.n5452 585
R2165 gnd.n5455 gnd.n76 585
R2166 gnd.n7413 gnd.n76 585
R2167 gnd.n5457 gnd.n5456 585
R2168 gnd.n5458 gnd.n5457 585
R2169 gnd.n3381 gnd.n3380 585
R2170 gnd.n3380 gnd.n3378 585
R2171 gnd.n5423 gnd.n5422 585
R2172 gnd.n5424 gnd.n5423 585
R2173 gnd.n3360 gnd.n3359 585
R2174 gnd.n5467 gnd.n3360 585
R2175 gnd.n5474 gnd.n5473 585
R2176 gnd.n5473 gnd.n5472 585
R2177 gnd.n5475 gnd.n3355 585
R2178 gnd.n5415 gnd.n3355 585
R2179 gnd.n5477 gnd.n5476 585
R2180 gnd.n5478 gnd.n5477 585
R2181 gnd.n3343 gnd.n3342 585
R2182 gnd.n5403 gnd.n3343 585
R2183 gnd.n5486 gnd.n5485 585
R2184 gnd.n5485 gnd.n5484 585
R2185 gnd.n5487 gnd.n3338 585
R2186 gnd.n5396 gnd.n3338 585
R2187 gnd.n5489 gnd.n5488 585
R2188 gnd.n5490 gnd.n5489 585
R2189 gnd.n3323 gnd.n3322 585
R2190 gnd.n5388 gnd.n3323 585
R2191 gnd.n5498 gnd.n5497 585
R2192 gnd.n5497 gnd.n5496 585
R2193 gnd.n5499 gnd.n3318 585
R2194 gnd.n5328 gnd.n3318 585
R2195 gnd.n5501 gnd.n5500 585
R2196 gnd.n5502 gnd.n5501 585
R2197 gnd.n3303 gnd.n3302 585
R2198 gnd.n5319 gnd.n3303 585
R2199 gnd.n5510 gnd.n5509 585
R2200 gnd.n5509 gnd.n5508 585
R2201 gnd.n5511 gnd.n3296 585
R2202 gnd.n5313 gnd.n3296 585
R2203 gnd.n5513 gnd.n5512 585
R2204 gnd.n5514 gnd.n5513 585
R2205 gnd.n3297 gnd.n3295 585
R2206 gnd.n5306 gnd.n3295 585
R2207 gnd.n3279 gnd.n3273 585
R2208 gnd.n5520 gnd.n3279 585
R2209 gnd.n5525 gnd.n3271 585
R2210 gnd.n5345 gnd.n3271 585
R2211 gnd.n5527 gnd.n5526 585
R2212 gnd.n5528 gnd.n5527 585
R2213 gnd.n3270 gnd.n3110 585
R2214 gnd.n5695 gnd.n3111 585
R2215 gnd.n5694 gnd.n3112 585
R2216 gnd.n3187 gnd.n3113 585
R2217 gnd.n5687 gnd.n3119 585
R2218 gnd.n5686 gnd.n3120 585
R2219 gnd.n3190 gnd.n3121 585
R2220 gnd.n5679 gnd.n3127 585
R2221 gnd.n5678 gnd.n3128 585
R2222 gnd.n3192 gnd.n3129 585
R2223 gnd.n5671 gnd.n3135 585
R2224 gnd.n5670 gnd.n3136 585
R2225 gnd.n3195 gnd.n3137 585
R2226 gnd.n5663 gnd.n3143 585
R2227 gnd.n5662 gnd.n3144 585
R2228 gnd.n3197 gnd.n3145 585
R2229 gnd.n5655 gnd.n3153 585
R2230 gnd.n5654 gnd.n5651 585
R2231 gnd.n3156 gnd.n3154 585
R2232 gnd.n5649 gnd.n3156 585
R2233 gnd.n7325 gnd.n7324 585
R2234 gnd.n7322 gnd.n7263 585
R2235 gnd.n7321 gnd.n7320 585
R2236 gnd.n7314 gnd.n7265 585
R2237 gnd.n7316 gnd.n7315 585
R2238 gnd.n7312 gnd.n7267 585
R2239 gnd.n7311 gnd.n7310 585
R2240 gnd.n7304 gnd.n7269 585
R2241 gnd.n7306 gnd.n7305 585
R2242 gnd.n7302 gnd.n7271 585
R2243 gnd.n7301 gnd.n7300 585
R2244 gnd.n7294 gnd.n7273 585
R2245 gnd.n7296 gnd.n7295 585
R2246 gnd.n7292 gnd.n7275 585
R2247 gnd.n7291 gnd.n7290 585
R2248 gnd.n7284 gnd.n7277 585
R2249 gnd.n7286 gnd.n7285 585
R2250 gnd.n7282 gnd.n7281 585
R2251 gnd.n7280 gnd.n172 585
R2252 gnd.n172 gnd.n171 585
R2253 gnd.n7328 gnd.n170 585
R2254 gnd.n7357 gnd.n170 585
R2255 gnd.n7330 gnd.n7329 585
R2256 gnd.n7329 gnd.n168 585
R2257 gnd.n7331 gnd.n161 585
R2258 gnd.n7363 gnd.n161 585
R2259 gnd.n7333 gnd.n7332 585
R2260 gnd.n7332 gnd.n153 585
R2261 gnd.n7334 gnd.n152 585
R2262 gnd.n7369 gnd.n152 585
R2263 gnd.n7336 gnd.n7335 585
R2264 gnd.n7335 gnd.n143 585
R2265 gnd.n7337 gnd.n142 585
R2266 gnd.n7375 gnd.n142 585
R2267 gnd.n7339 gnd.n7338 585
R2268 gnd.n7340 gnd.n7339 585
R2269 gnd.n388 gnd.n133 585
R2270 gnd.n7381 gnd.n133 585
R2271 gnd.n7250 gnd.n7249 585
R2272 gnd.n7249 gnd.n7248 585
R2273 gnd.n390 gnd.n122 585
R2274 gnd.n7387 gnd.n122 585
R2275 gnd.n7240 gnd.n7239 585
R2276 gnd.n7241 gnd.n7240 585
R2277 gnd.n393 gnd.n113 585
R2278 gnd.n7393 gnd.n113 585
R2279 gnd.n7235 gnd.n7234 585
R2280 gnd.n7234 gnd.n7233 585
R2281 gnd.n395 gnd.n103 585
R2282 gnd.n7399 gnd.n103 585
R2283 gnd.n5438 gnd.n397 585
R2284 gnd.n7226 gnd.n397 585
R2285 gnd.n5439 gnd.n92 585
R2286 gnd.n7405 gnd.n92 585
R2287 gnd.n5441 gnd.n5440 585
R2288 gnd.n5442 gnd.n5441 585
R2289 gnd.n72 gnd.n71 585
R2290 gnd.n5452 gnd.n72 585
R2291 gnd.n7415 gnd.n7414 585
R2292 gnd.n7414 gnd.n7413 585
R2293 gnd.n7416 gnd.n70 585
R2294 gnd.n5458 gnd.n70 585
R2295 gnd.n3388 gnd.n68 585
R2296 gnd.n3388 gnd.n3378 585
R2297 gnd.n5408 gnd.n3389 585
R2298 gnd.n5424 gnd.n3389 585
R2299 gnd.n5409 gnd.n3369 585
R2300 gnd.n5467 gnd.n3369 585
R2301 gnd.n3393 gnd.n3363 585
R2302 gnd.n5472 gnd.n3363 585
R2303 gnd.n5414 gnd.n5413 585
R2304 gnd.n5415 gnd.n5414 585
R2305 gnd.n3392 gnd.n3353 585
R2306 gnd.n5478 gnd.n3353 585
R2307 gnd.n5405 gnd.n5404 585
R2308 gnd.n5404 gnd.n5403 585
R2309 gnd.n3395 gnd.n3346 585
R2310 gnd.n5484 gnd.n3346 585
R2311 gnd.n5395 gnd.n5394 585
R2312 gnd.n5396 gnd.n5395 585
R2313 gnd.n3398 gnd.n3336 585
R2314 gnd.n5490 gnd.n3336 585
R2315 gnd.n5390 gnd.n5389 585
R2316 gnd.n5389 gnd.n5388 585
R2317 gnd.n3400 gnd.n3326 585
R2318 gnd.n5496 gnd.n3326 585
R2319 gnd.n5331 gnd.n5329 585
R2320 gnd.n5329 gnd.n5328 585
R2321 gnd.n5332 gnd.n3316 585
R2322 gnd.n5502 gnd.n3316 585
R2323 gnd.n5333 gnd.n5311 585
R2324 gnd.n5319 gnd.n5311 585
R2325 gnd.n5309 gnd.n3306 585
R2326 gnd.n5508 gnd.n3306 585
R2327 gnd.n5337 gnd.n5308 585
R2328 gnd.n5313 gnd.n5308 585
R2329 gnd.n5338 gnd.n3293 585
R2330 gnd.n5514 gnd.n3293 585
R2331 gnd.n5339 gnd.n5307 585
R2332 gnd.n5307 gnd.n5306 585
R2333 gnd.n3417 gnd.n3277 585
R2334 gnd.n5520 gnd.n3277 585
R2335 gnd.n5344 gnd.n5343 585
R2336 gnd.n5345 gnd.n5344 585
R2337 gnd.n3416 gnd.n3268 585
R2338 gnd.n5528 gnd.n3268 585
R2339 gnd.n1039 gnd.n1038 585
R2340 gnd.n1043 gnd.n1039 585
R2341 gnd.n6342 gnd.n6341 585
R2342 gnd.n6341 gnd.n6340 585
R2343 gnd.n6343 gnd.n1031 585
R2344 gnd.n2331 gnd.n1031 585
R2345 gnd.n6345 gnd.n6344 585
R2346 gnd.n6346 gnd.n6345 585
R2347 gnd.n1032 gnd.n1030 585
R2348 gnd.n1030 gnd.n1027 585
R2349 gnd.n1014 gnd.n1013 585
R2350 gnd.n1018 gnd.n1014 585
R2351 gnd.n6356 gnd.n6355 585
R2352 gnd.n6355 gnd.n6354 585
R2353 gnd.n6357 gnd.n1006 585
R2354 gnd.n1151 gnd.n1006 585
R2355 gnd.n6359 gnd.n6358 585
R2356 gnd.n6360 gnd.n6359 585
R2357 gnd.n1007 gnd.n1005 585
R2358 gnd.n1005 gnd.n1001 585
R2359 gnd.n988 gnd.n987 585
R2360 gnd.n992 gnd.n988 585
R2361 gnd.n6370 gnd.n6369 585
R2362 gnd.n6369 gnd.n6368 585
R2363 gnd.n6371 gnd.n982 585
R2364 gnd.n1154 gnd.n982 585
R2365 gnd.n6373 gnd.n6372 585
R2366 gnd.n6374 gnd.n6373 585
R2367 gnd.n983 gnd.n981 585
R2368 gnd.n2038 gnd.n981 585
R2369 gnd.n2022 gnd.n1174 585
R2370 gnd.n1174 gnd.n1173 585
R2371 gnd.n2024 gnd.n2023 585
R2372 gnd.n2025 gnd.n2024 585
R2373 gnd.n1175 gnd.n1172 585
R2374 gnd.n1172 gnd.n1168 585
R2375 gnd.n2016 gnd.n2015 585
R2376 gnd.n2015 gnd.n2014 585
R2377 gnd.n1178 gnd.n1177 585
R2378 gnd.n1186 gnd.n1178 585
R2379 gnd.n1951 gnd.n1950 585
R2380 gnd.n1952 gnd.n1951 585
R2381 gnd.n1197 gnd.n1196 585
R2382 gnd.n1204 gnd.n1196 585
R2383 gnd.n1946 gnd.n1945 585
R2384 gnd.n1945 gnd.n1944 585
R2385 gnd.n1200 gnd.n1199 585
R2386 gnd.n1934 gnd.n1200 585
R2387 gnd.n1921 gnd.n1223 585
R2388 gnd.n1223 gnd.n1214 585
R2389 gnd.n1923 gnd.n1922 585
R2390 gnd.n1924 gnd.n1923 585
R2391 gnd.n1224 gnd.n1222 585
R2392 gnd.n1231 gnd.n1222 585
R2393 gnd.n1916 gnd.n1915 585
R2394 gnd.n1915 gnd.n1914 585
R2395 gnd.n1227 gnd.n1226 585
R2396 gnd.n1903 gnd.n1227 585
R2397 gnd.n1890 gnd.n1248 585
R2398 gnd.n1248 gnd.n1239 585
R2399 gnd.n1892 gnd.n1891 585
R2400 gnd.n1893 gnd.n1892 585
R2401 gnd.n1249 gnd.n1247 585
R2402 gnd.n1256 gnd.n1247 585
R2403 gnd.n1885 gnd.n1884 585
R2404 gnd.n1884 gnd.n1883 585
R2405 gnd.n1252 gnd.n1251 585
R2406 gnd.n1872 gnd.n1252 585
R2407 gnd.n1859 gnd.n1274 585
R2408 gnd.n1274 gnd.n1264 585
R2409 gnd.n1861 gnd.n1860 585
R2410 gnd.n1862 gnd.n1861 585
R2411 gnd.n1275 gnd.n1273 585
R2412 gnd.n1282 gnd.n1273 585
R2413 gnd.n1854 gnd.n1853 585
R2414 gnd.n1853 gnd.n1852 585
R2415 gnd.n1278 gnd.n1277 585
R2416 gnd.n1841 gnd.n1278 585
R2417 gnd.n1828 gnd.n1300 585
R2418 gnd.n1300 gnd.n1299 585
R2419 gnd.n1830 gnd.n1829 585
R2420 gnd.n1831 gnd.n1830 585
R2421 gnd.n1301 gnd.n1298 585
R2422 gnd.n1308 gnd.n1298 585
R2423 gnd.n1823 gnd.n1822 585
R2424 gnd.n1822 gnd.n1821 585
R2425 gnd.n1304 gnd.n1303 585
R2426 gnd.n1810 gnd.n1304 585
R2427 gnd.n1797 gnd.n1326 585
R2428 gnd.n1326 gnd.n1325 585
R2429 gnd.n1799 gnd.n1798 585
R2430 gnd.n1800 gnd.n1799 585
R2431 gnd.n1327 gnd.n1324 585
R2432 gnd.n1334 gnd.n1324 585
R2433 gnd.n1792 gnd.n1791 585
R2434 gnd.n1791 gnd.n1790 585
R2435 gnd.n1330 gnd.n1329 585
R2436 gnd.n1779 gnd.n1330 585
R2437 gnd.n1766 gnd.n1351 585
R2438 gnd.n1351 gnd.n1342 585
R2439 gnd.n1768 gnd.n1767 585
R2440 gnd.n1769 gnd.n1768 585
R2441 gnd.n1352 gnd.n1350 585
R2442 gnd.n1359 gnd.n1350 585
R2443 gnd.n1761 gnd.n1760 585
R2444 gnd.n1760 gnd.n1759 585
R2445 gnd.n1355 gnd.n1354 585
R2446 gnd.n1748 gnd.n1355 585
R2447 gnd.n1735 gnd.n1734 585
R2448 gnd.n1733 gnd.n1686 585
R2449 gnd.n1732 gnd.n1685 585
R2450 gnd.n1737 gnd.n1685 585
R2451 gnd.n1731 gnd.n1730 585
R2452 gnd.n1729 gnd.n1728 585
R2453 gnd.n1727 gnd.n1726 585
R2454 gnd.n1725 gnd.n1724 585
R2455 gnd.n1723 gnd.n1722 585
R2456 gnd.n1721 gnd.n1720 585
R2457 gnd.n1719 gnd.n1718 585
R2458 gnd.n1717 gnd.n1716 585
R2459 gnd.n1715 gnd.n1714 585
R2460 gnd.n1713 gnd.n1712 585
R2461 gnd.n1711 gnd.n1710 585
R2462 gnd.n1709 gnd.n1708 585
R2463 gnd.n1707 gnd.n1706 585
R2464 gnd.n1702 gnd.n1365 585
R2465 gnd.n6332 gnd.n6331 585
R2466 gnd.n6325 gnd.n1053 585
R2467 gnd.n6327 gnd.n6326 585
R2468 gnd.n1056 gnd.n1055 585
R2469 gnd.n6297 gnd.n6296 585
R2470 gnd.n6299 gnd.n6298 585
R2471 gnd.n6301 gnd.n6300 585
R2472 gnd.n6303 gnd.n6302 585
R2473 gnd.n6305 gnd.n6304 585
R2474 gnd.n6307 gnd.n6306 585
R2475 gnd.n6309 gnd.n6308 585
R2476 gnd.n6311 gnd.n6310 585
R2477 gnd.n6313 gnd.n6312 585
R2478 gnd.n6316 gnd.n6315 585
R2479 gnd.n6314 gnd.n6286 585
R2480 gnd.n6320 gnd.n6283 585
R2481 gnd.n6322 gnd.n6321 585
R2482 gnd.n6323 gnd.n6322 585
R2483 gnd.n6334 gnd.n6333 585
R2484 gnd.n6333 gnd.n1043 585
R2485 gnd.n1049 gnd.n1041 585
R2486 gnd.n6340 gnd.n1041 585
R2487 gnd.n2330 gnd.n2329 585
R2488 gnd.n2331 gnd.n2330 585
R2489 gnd.n2324 gnd.n1029 585
R2490 gnd.n6346 gnd.n1029 585
R2491 gnd.n2323 gnd.n2322 585
R2492 gnd.n2322 gnd.n1027 585
R2493 gnd.n2321 gnd.n2319 585
R2494 gnd.n2321 gnd.n1018 585
R2495 gnd.n2061 gnd.n1016 585
R2496 gnd.n6354 gnd.n1016 585
R2497 gnd.n1153 gnd.n1152 585
R2498 gnd.n1152 gnd.n1151 585
R2499 gnd.n2055 gnd.n1003 585
R2500 gnd.n6360 gnd.n1003 585
R2501 gnd.n2054 gnd.n2053 585
R2502 gnd.n2053 gnd.n1001 585
R2503 gnd.n2052 gnd.n2050 585
R2504 gnd.n2052 gnd.n992 585
R2505 gnd.n2048 gnd.n990 585
R2506 gnd.n6368 gnd.n990 585
R2507 gnd.n1156 gnd.n1155 585
R2508 gnd.n1155 gnd.n1154 585
R2509 gnd.n2035 gnd.n979 585
R2510 gnd.n6374 gnd.n979 585
R2511 gnd.n2037 gnd.n2036 585
R2512 gnd.n2038 gnd.n2037 585
R2513 gnd.n1163 gnd.n1162 585
R2514 gnd.n1173 gnd.n1162 585
R2515 gnd.n1957 gnd.n1170 585
R2516 gnd.n2025 gnd.n1170 585
R2517 gnd.n1959 gnd.n1958 585
R2518 gnd.n1958 gnd.n1168 585
R2519 gnd.n1960 gnd.n1180 585
R2520 gnd.n2014 gnd.n1180 585
R2521 gnd.n1955 gnd.n1954 585
R2522 gnd.n1954 gnd.n1186 585
R2523 gnd.n1953 gnd.n1193 585
R2524 gnd.n1953 gnd.n1952 585
R2525 gnd.n1938 gnd.n1194 585
R2526 gnd.n1204 gnd.n1194 585
R2527 gnd.n1937 gnd.n1202 585
R2528 gnd.n1944 gnd.n1202 585
R2529 gnd.n1936 gnd.n1935 585
R2530 gnd.n1935 gnd.n1934 585
R2531 gnd.n1213 gnd.n1210 585
R2532 gnd.n1214 gnd.n1213 585
R2533 gnd.n1926 gnd.n1925 585
R2534 gnd.n1925 gnd.n1924 585
R2535 gnd.n1220 gnd.n1219 585
R2536 gnd.n1231 gnd.n1220 585
R2537 gnd.n1906 gnd.n1229 585
R2538 gnd.n1914 gnd.n1229 585
R2539 gnd.n1905 gnd.n1904 585
R2540 gnd.n1904 gnd.n1903 585
R2541 gnd.n1238 gnd.n1236 585
R2542 gnd.n1239 gnd.n1238 585
R2543 gnd.n1895 gnd.n1894 585
R2544 gnd.n1894 gnd.n1893 585
R2545 gnd.n1245 gnd.n1244 585
R2546 gnd.n1256 gnd.n1245 585
R2547 gnd.n1875 gnd.n1254 585
R2548 gnd.n1883 gnd.n1254 585
R2549 gnd.n1874 gnd.n1873 585
R2550 gnd.n1873 gnd.n1872 585
R2551 gnd.n1263 gnd.n1261 585
R2552 gnd.n1264 gnd.n1263 585
R2553 gnd.n1864 gnd.n1863 585
R2554 gnd.n1863 gnd.n1862 585
R2555 gnd.n1270 gnd.n1269 585
R2556 gnd.n1282 gnd.n1270 585
R2557 gnd.n1844 gnd.n1280 585
R2558 gnd.n1852 gnd.n1280 585
R2559 gnd.n1843 gnd.n1842 585
R2560 gnd.n1842 gnd.n1841 585
R2561 gnd.n1289 gnd.n1287 585
R2562 gnd.n1299 gnd.n1289 585
R2563 gnd.n1833 gnd.n1832 585
R2564 gnd.n1832 gnd.n1831 585
R2565 gnd.n1295 gnd.n1294 585
R2566 gnd.n1308 gnd.n1295 585
R2567 gnd.n1813 gnd.n1306 585
R2568 gnd.n1821 gnd.n1306 585
R2569 gnd.n1812 gnd.n1811 585
R2570 gnd.n1811 gnd.n1810 585
R2571 gnd.n1315 gnd.n1313 585
R2572 gnd.n1325 gnd.n1315 585
R2573 gnd.n1802 gnd.n1801 585
R2574 gnd.n1801 gnd.n1800 585
R2575 gnd.n1321 gnd.n1320 585
R2576 gnd.n1334 gnd.n1321 585
R2577 gnd.n1782 gnd.n1332 585
R2578 gnd.n1790 gnd.n1332 585
R2579 gnd.n1781 gnd.n1780 585
R2580 gnd.n1780 gnd.n1779 585
R2581 gnd.n1341 gnd.n1339 585
R2582 gnd.n1342 gnd.n1341 585
R2583 gnd.n1771 gnd.n1770 585
R2584 gnd.n1770 gnd.n1769 585
R2585 gnd.n1348 gnd.n1347 585
R2586 gnd.n1359 gnd.n1348 585
R2587 gnd.n1751 gnd.n1357 585
R2588 gnd.n1759 gnd.n1357 585
R2589 gnd.n1750 gnd.n1749 585
R2590 gnd.n1749 gnd.n1748 585
R2591 gnd.n5160 gnd.n5159 585
R2592 gnd.n5161 gnd.n5160 585
R2593 gnd.n4969 gnd.n3533 585
R2594 gnd.n3533 gnd.n3517 585
R2595 gnd.n4968 gnd.n4967 585
R2596 gnd.n4967 gnd.n3516 585
R2597 gnd.n4966 gnd.n3525 585
R2598 gnd.t97 gnd.n3525 585
R2599 gnd.n4965 gnd.n4964 585
R2600 gnd.n4964 gnd.n3523 585
R2601 gnd.n4963 gnd.n3535 585
R2602 gnd.n4963 gnd.n4962 585
R2603 gnd.n4953 gnd.n3536 585
R2604 gnd.n3540 gnd.n3536 585
R2605 gnd.n4955 gnd.n4954 585
R2606 gnd.n4956 gnd.n4955 585
R2607 gnd.n4952 gnd.n3542 585
R2608 gnd.n3547 gnd.n3542 585
R2609 gnd.n4951 gnd.n4950 585
R2610 gnd.n4950 gnd.n4949 585
R2611 gnd.n3544 gnd.n3543 585
R2612 gnd.n4911 gnd.n3544 585
R2613 gnd.n4936 gnd.n4935 585
R2614 gnd.n4937 gnd.n4936 585
R2615 gnd.n4934 gnd.n3557 585
R2616 gnd.n3557 gnd.n3554 585
R2617 gnd.n4933 gnd.n4932 585
R2618 gnd.n4932 gnd.n4931 585
R2619 gnd.n3559 gnd.n3558 585
R2620 gnd.n3560 gnd.n3559 585
R2621 gnd.n4899 gnd.n4898 585
R2622 gnd.n4900 gnd.n4899 585
R2623 gnd.n4897 gnd.n3570 585
R2624 gnd.n4893 gnd.n3570 585
R2625 gnd.n4896 gnd.n4895 585
R2626 gnd.n4895 gnd.n4894 585
R2627 gnd.n3572 gnd.n3571 585
R2628 gnd.n4881 gnd.n3572 585
R2629 gnd.n4870 gnd.n3589 585
R2630 gnd.n3589 gnd.n3583 585
R2631 gnd.n4872 gnd.n4871 585
R2632 gnd.n4873 gnd.n4872 585
R2633 gnd.n4869 gnd.n3588 585
R2634 gnd.n3594 gnd.n3588 585
R2635 gnd.n4868 gnd.n4867 585
R2636 gnd.n4867 gnd.n4866 585
R2637 gnd.n3591 gnd.n3590 585
R2638 gnd.n4843 gnd.n3591 585
R2639 gnd.n4855 gnd.n4854 585
R2640 gnd.n4856 gnd.n4855 585
R2641 gnd.n4853 gnd.n3604 585
R2642 gnd.n4849 gnd.n3604 585
R2643 gnd.n4852 gnd.n4851 585
R2644 gnd.n4851 gnd.n4850 585
R2645 gnd.n3606 gnd.n3605 585
R2646 gnd.n4838 gnd.n3606 585
R2647 gnd.n4824 gnd.n4823 585
R2648 gnd.n4823 gnd.n3611 585
R2649 gnd.n4825 gnd.n3623 585
R2650 gnd.n4787 gnd.n3623 585
R2651 gnd.n4827 gnd.n4826 585
R2652 gnd.n4828 gnd.n4827 585
R2653 gnd.n4822 gnd.n3622 585
R2654 gnd.n3622 gnd.n3619 585
R2655 gnd.n4821 gnd.n4820 585
R2656 gnd.n4820 gnd.n4819 585
R2657 gnd.n3625 gnd.n3624 585
R2658 gnd.n4778 gnd.n3625 585
R2659 gnd.n4764 gnd.n4763 585
R2660 gnd.n4763 gnd.n3634 585
R2661 gnd.n4765 gnd.n3645 585
R2662 gnd.n3645 gnd.n3643 585
R2663 gnd.n4767 gnd.n4766 585
R2664 gnd.n4768 gnd.n4767 585
R2665 gnd.n4762 gnd.n3644 585
R2666 gnd.n4757 gnd.n3644 585
R2667 gnd.n4761 gnd.n4760 585
R2668 gnd.n4760 gnd.n4759 585
R2669 gnd.n3647 gnd.n3646 585
R2670 gnd.n3648 gnd.n3647 585
R2671 gnd.n4746 gnd.n4745 585
R2672 gnd.n4747 gnd.n4746 585
R2673 gnd.n4744 gnd.n3656 585
R2674 gnd.n4740 gnd.n3656 585
R2675 gnd.n4743 gnd.n4742 585
R2676 gnd.n4742 gnd.n4741 585
R2677 gnd.n3658 gnd.n3657 585
R2678 gnd.n3664 gnd.n3658 585
R2679 gnd.n4732 gnd.n4731 585
R2680 gnd.n4733 gnd.n4732 585
R2681 gnd.n4730 gnd.n3666 585
R2682 gnd.n3666 gnd.n3663 585
R2683 gnd.n4729 gnd.n4728 585
R2684 gnd.n4728 gnd.n4727 585
R2685 gnd.n3668 gnd.n3667 585
R2686 gnd.n4633 gnd.n3668 585
R2687 gnd.n4705 gnd.n4704 585
R2688 gnd.n4706 gnd.n4705 585
R2689 gnd.n4703 gnd.n3682 585
R2690 gnd.n3682 gnd.n3679 585
R2691 gnd.n4702 gnd.n4701 585
R2692 gnd.n4701 gnd.n4700 585
R2693 gnd.n3684 gnd.n3683 585
R2694 gnd.n4642 gnd.n3684 585
R2695 gnd.n3707 gnd.n3706 585
R2696 gnd.n3707 gnd.n3692 585
R2697 gnd.n4650 gnd.n4649 585
R2698 gnd.n4649 gnd.n4648 585
R2699 gnd.n4651 gnd.n3704 585
R2700 gnd.n3704 gnd.n3702 585
R2701 gnd.n4653 gnd.n4652 585
R2702 gnd.n4654 gnd.n4653 585
R2703 gnd.n3705 gnd.n3703 585
R2704 gnd.n3703 gnd.n3699 585
R2705 gnd.n4625 gnd.n4624 585
R2706 gnd.n4626 gnd.n4625 585
R2707 gnd.n4623 gnd.n3713 585
R2708 gnd.n3719 gnd.n3713 585
R2709 gnd.n4622 gnd.n4621 585
R2710 gnd.n4621 gnd.n4620 585
R2711 gnd.n3715 gnd.n3714 585
R2712 gnd.n3728 gnd.n3715 585
R2713 gnd.n4609 gnd.n4608 585
R2714 gnd.n4610 gnd.n4609 585
R2715 gnd.n4607 gnd.n3729 585
R2716 gnd.n3729 gnd.n3725 585
R2717 gnd.n4606 gnd.n4605 585
R2718 gnd.n4605 gnd.n4604 585
R2719 gnd.n3731 gnd.n3730 585
R2720 gnd.n4536 gnd.n3731 585
R2721 gnd.n4563 gnd.n4562 585
R2722 gnd.n4563 gnd.n3740 585
R2723 gnd.n4565 gnd.n4564 585
R2724 gnd.n4564 gnd.n3739 585
R2725 gnd.n4566 gnd.n3751 585
R2726 gnd.n4551 gnd.n3751 585
R2727 gnd.n4568 gnd.n4567 585
R2728 gnd.n4569 gnd.n4568 585
R2729 gnd.n4561 gnd.n3750 585
R2730 gnd.n3750 gnd.n3747 585
R2731 gnd.n4560 gnd.n4559 585
R2732 gnd.n4559 gnd.n4558 585
R2733 gnd.n3753 gnd.n3752 585
R2734 gnd.n3759 gnd.n3753 585
R2735 gnd.n4529 gnd.n4528 585
R2736 gnd.n4530 gnd.n4529 585
R2737 gnd.n4527 gnd.n3761 585
R2738 gnd.n4515 gnd.n3761 585
R2739 gnd.n4526 gnd.n4525 585
R2740 gnd.n4525 gnd.n4524 585
R2741 gnd.n3767 gnd.n3762 585
R2742 gnd.n3769 gnd.n3767 585
R2743 gnd.n3766 gnd.n3765 585
R2744 gnd.n3766 gnd.n2989 585
R2745 gnd.n3764 gnd.n3763 585
R2746 gnd.n3763 gnd.n2987 585
R2747 gnd.n2973 gnd.n2972 585
R2748 gnd.n2977 gnd.n2973 585
R2749 gnd.n5843 gnd.n5842 585
R2750 gnd.n5842 gnd.n5841 585
R2751 gnd.n5844 gnd.n2951 585
R2752 gnd.n2974 gnd.n2951 585
R2753 gnd.n5909 gnd.n5908 585
R2754 gnd.n5907 gnd.n2950 585
R2755 gnd.n5906 gnd.n2949 585
R2756 gnd.n5911 gnd.n2949 585
R2757 gnd.n5905 gnd.n5904 585
R2758 gnd.n5903 gnd.n5902 585
R2759 gnd.n5901 gnd.n5900 585
R2760 gnd.n5899 gnd.n5898 585
R2761 gnd.n5897 gnd.n5896 585
R2762 gnd.n5895 gnd.n5894 585
R2763 gnd.n5893 gnd.n5892 585
R2764 gnd.n5891 gnd.n5890 585
R2765 gnd.n5889 gnd.n5888 585
R2766 gnd.n5887 gnd.n5886 585
R2767 gnd.n5885 gnd.n5884 585
R2768 gnd.n5883 gnd.n5882 585
R2769 gnd.n5881 gnd.n5880 585
R2770 gnd.n5879 gnd.n5878 585
R2771 gnd.n5877 gnd.n5876 585
R2772 gnd.n5875 gnd.n5874 585
R2773 gnd.n5873 gnd.n5872 585
R2774 gnd.n5871 gnd.n5870 585
R2775 gnd.n5869 gnd.n5868 585
R2776 gnd.n5867 gnd.n5866 585
R2777 gnd.n5865 gnd.n5864 585
R2778 gnd.n5863 gnd.n5862 585
R2779 gnd.n5861 gnd.n5860 585
R2780 gnd.n5859 gnd.n5858 585
R2781 gnd.n5857 gnd.n5856 585
R2782 gnd.n5855 gnd.n5854 585
R2783 gnd.n5853 gnd.n5852 585
R2784 gnd.n5851 gnd.n5850 585
R2785 gnd.n5849 gnd.n2913 585
R2786 gnd.n5914 gnd.n5913 585
R2787 gnd.n2915 gnd.n2912 585
R2788 gnd.n3775 gnd.n3774 585
R2789 gnd.n3777 gnd.n3776 585
R2790 gnd.n3780 gnd.n3779 585
R2791 gnd.n3782 gnd.n3781 585
R2792 gnd.n3784 gnd.n3783 585
R2793 gnd.n3786 gnd.n3785 585
R2794 gnd.n3788 gnd.n3787 585
R2795 gnd.n3790 gnd.n3789 585
R2796 gnd.n3792 gnd.n3791 585
R2797 gnd.n3794 gnd.n3793 585
R2798 gnd.n3796 gnd.n3795 585
R2799 gnd.n3798 gnd.n3797 585
R2800 gnd.n3800 gnd.n3799 585
R2801 gnd.n3802 gnd.n3801 585
R2802 gnd.n3804 gnd.n3803 585
R2803 gnd.n3806 gnd.n3805 585
R2804 gnd.n3808 gnd.n3807 585
R2805 gnd.n3810 gnd.n3809 585
R2806 gnd.n3812 gnd.n3811 585
R2807 gnd.n3814 gnd.n3813 585
R2808 gnd.n3816 gnd.n3815 585
R2809 gnd.n3818 gnd.n3817 585
R2810 gnd.n3820 gnd.n3819 585
R2811 gnd.n3822 gnd.n3821 585
R2812 gnd.n3824 gnd.n3823 585
R2813 gnd.n3826 gnd.n3825 585
R2814 gnd.n3828 gnd.n3827 585
R2815 gnd.n3830 gnd.n3829 585
R2816 gnd.n3832 gnd.n3831 585
R2817 gnd.n3834 gnd.n3833 585
R2818 gnd.n3836 gnd.n3835 585
R2819 gnd.n5041 gnd.n3531 585
R2820 gnd.n5042 gnd.n5040 585
R2821 gnd.n5044 gnd.n5043 585
R2822 gnd.n5046 gnd.n5037 585
R2823 gnd.n5048 gnd.n5047 585
R2824 gnd.n5049 gnd.n5036 585
R2825 gnd.n5051 gnd.n5050 585
R2826 gnd.n5053 gnd.n5034 585
R2827 gnd.n5055 gnd.n5054 585
R2828 gnd.n5056 gnd.n5033 585
R2829 gnd.n5058 gnd.n5057 585
R2830 gnd.n5060 gnd.n5031 585
R2831 gnd.n5062 gnd.n5061 585
R2832 gnd.n5063 gnd.n5030 585
R2833 gnd.n5065 gnd.n5064 585
R2834 gnd.n5067 gnd.n5028 585
R2835 gnd.n5069 gnd.n5068 585
R2836 gnd.n5070 gnd.n5027 585
R2837 gnd.n5072 gnd.n5071 585
R2838 gnd.n5074 gnd.n5025 585
R2839 gnd.n5076 gnd.n5075 585
R2840 gnd.n5077 gnd.n5024 585
R2841 gnd.n5079 gnd.n5078 585
R2842 gnd.n5081 gnd.n5022 585
R2843 gnd.n5083 gnd.n5082 585
R2844 gnd.n5084 gnd.n5021 585
R2845 gnd.n5086 gnd.n5085 585
R2846 gnd.n5088 gnd.n5019 585
R2847 gnd.n5090 gnd.n5089 585
R2848 gnd.n5092 gnd.n5016 585
R2849 gnd.n5094 gnd.n5093 585
R2850 gnd.n5096 gnd.n5015 585
R2851 gnd.n5097 gnd.n4991 585
R2852 gnd.n5100 gnd.n3231 585
R2853 gnd.n5102 gnd.n5101 585
R2854 gnd.n5104 gnd.n5013 585
R2855 gnd.n5106 gnd.n5105 585
R2856 gnd.n5108 gnd.n5010 585
R2857 gnd.n5110 gnd.n5109 585
R2858 gnd.n5112 gnd.n5008 585
R2859 gnd.n5114 gnd.n5113 585
R2860 gnd.n5115 gnd.n5007 585
R2861 gnd.n5117 gnd.n5116 585
R2862 gnd.n5119 gnd.n5005 585
R2863 gnd.n5121 gnd.n5120 585
R2864 gnd.n5122 gnd.n5004 585
R2865 gnd.n5124 gnd.n5123 585
R2866 gnd.n5126 gnd.n5002 585
R2867 gnd.n5128 gnd.n5127 585
R2868 gnd.n5129 gnd.n5001 585
R2869 gnd.n5131 gnd.n5130 585
R2870 gnd.n5133 gnd.n4999 585
R2871 gnd.n5135 gnd.n5134 585
R2872 gnd.n5136 gnd.n4998 585
R2873 gnd.n5138 gnd.n5137 585
R2874 gnd.n5140 gnd.n4996 585
R2875 gnd.n5142 gnd.n5141 585
R2876 gnd.n5143 gnd.n4995 585
R2877 gnd.n5145 gnd.n5144 585
R2878 gnd.n5147 gnd.n4993 585
R2879 gnd.n5149 gnd.n5148 585
R2880 gnd.n5150 gnd.n4992 585
R2881 gnd.n5152 gnd.n5151 585
R2882 gnd.n5154 gnd.n4989 585
R2883 gnd.n5156 gnd.n5155 585
R2884 gnd.n5157 gnd.n3534 585
R2885 gnd.n5162 gnd.n3530 585
R2886 gnd.n5162 gnd.n5161 585
R2887 gnd.n5164 gnd.n5163 585
R2888 gnd.n5163 gnd.n3517 585
R2889 gnd.n5165 gnd.n3528 585
R2890 gnd.n3528 gnd.n3516 585
R2891 gnd.n5167 gnd.n5166 585
R2892 gnd.t97 gnd.n5167 585
R2893 gnd.n3529 gnd.n3527 585
R2894 gnd.n3527 gnd.n3523 585
R2895 gnd.n4961 gnd.n4960 585
R2896 gnd.n4962 gnd.n4961 585
R2897 gnd.n4959 gnd.n3537 585
R2898 gnd.n3540 gnd.n3537 585
R2899 gnd.n4958 gnd.n4957 585
R2900 gnd.n4957 gnd.n4956 585
R2901 gnd.n3539 gnd.n3538 585
R2902 gnd.n3547 gnd.n3539 585
R2903 gnd.n4908 gnd.n3545 585
R2904 gnd.n4949 gnd.n3545 585
R2905 gnd.n4910 gnd.n4909 585
R2906 gnd.n4911 gnd.n4910 585
R2907 gnd.n4907 gnd.n3556 585
R2908 gnd.n4937 gnd.n3556 585
R2909 gnd.n4906 gnd.n4905 585
R2910 gnd.n4905 gnd.n3554 585
R2911 gnd.n4904 gnd.n3561 585
R2912 gnd.n4931 gnd.n3561 585
R2913 gnd.n4903 gnd.n4902 585
R2914 gnd.n4902 gnd.n3560 585
R2915 gnd.n4901 gnd.n3567 585
R2916 gnd.n4901 gnd.n4900 585
R2917 gnd.n4877 gnd.n3568 585
R2918 gnd.n4893 gnd.n3568 585
R2919 gnd.n4878 gnd.n3574 585
R2920 gnd.n4894 gnd.n3574 585
R2921 gnd.n4880 gnd.n4879 585
R2922 gnd.n4881 gnd.n4880 585
R2923 gnd.n4876 gnd.n3585 585
R2924 gnd.n3585 gnd.n3583 585
R2925 gnd.n4875 gnd.n4874 585
R2926 gnd.n4874 gnd.n4873 585
R2927 gnd.n3587 gnd.n3586 585
R2928 gnd.n3594 gnd.n3587 585
R2929 gnd.n4842 gnd.n3592 585
R2930 gnd.n4866 gnd.n3592 585
R2931 gnd.n4845 gnd.n4844 585
R2932 gnd.n4844 gnd.n4843 585
R2933 gnd.n4846 gnd.n3602 585
R2934 gnd.n4856 gnd.n3602 585
R2935 gnd.n4848 gnd.n4847 585
R2936 gnd.n4849 gnd.n4848 585
R2937 gnd.n4841 gnd.n3608 585
R2938 gnd.n4850 gnd.n3608 585
R2939 gnd.n4840 gnd.n4839 585
R2940 gnd.n4839 gnd.n4838 585
R2941 gnd.n3610 gnd.n3609 585
R2942 gnd.n3611 gnd.n3610 585
R2943 gnd.n4786 gnd.n4785 585
R2944 gnd.n4787 gnd.n4786 585
R2945 gnd.n4784 gnd.n3621 585
R2946 gnd.n4828 gnd.n3621 585
R2947 gnd.n4783 gnd.n4782 585
R2948 gnd.n4782 gnd.n3619 585
R2949 gnd.n4781 gnd.n3626 585
R2950 gnd.n4819 gnd.n3626 585
R2951 gnd.n4780 gnd.n4779 585
R2952 gnd.n4779 gnd.n4778 585
R2953 gnd.n3633 gnd.n3632 585
R2954 gnd.n3634 gnd.n3633 585
R2955 gnd.n4753 gnd.n4752 585
R2956 gnd.n4752 gnd.n3643 585
R2957 gnd.n4754 gnd.n3642 585
R2958 gnd.n4768 gnd.n3642 585
R2959 gnd.n4756 gnd.n4755 585
R2960 gnd.n4757 gnd.n4756 585
R2961 gnd.n4751 gnd.n3649 585
R2962 gnd.n4759 gnd.n3649 585
R2963 gnd.n4750 gnd.n4749 585
R2964 gnd.n4749 gnd.n3648 585
R2965 gnd.n4748 gnd.n3651 585
R2966 gnd.n4748 gnd.n4747 585
R2967 gnd.n4737 gnd.n3652 585
R2968 gnd.n4740 gnd.n3652 585
R2969 gnd.n4739 gnd.n4738 585
R2970 gnd.n4741 gnd.n4739 585
R2971 gnd.n4736 gnd.n3660 585
R2972 gnd.n3664 gnd.n3660 585
R2973 gnd.n4735 gnd.n4734 585
R2974 gnd.n4734 gnd.n4733 585
R2975 gnd.n3662 gnd.n3661 585
R2976 gnd.n3663 gnd.n3662 585
R2977 gnd.n4632 gnd.n3670 585
R2978 gnd.n4727 gnd.n3670 585
R2979 gnd.n4635 gnd.n4634 585
R2980 gnd.n4634 gnd.n4633 585
R2981 gnd.n4636 gnd.n3681 585
R2982 gnd.n4706 gnd.n3681 585
R2983 gnd.n4638 gnd.n4637 585
R2984 gnd.n4637 gnd.n3679 585
R2985 gnd.n4639 gnd.n3685 585
R2986 gnd.n4700 gnd.n3685 585
R2987 gnd.n4644 gnd.n4643 585
R2988 gnd.n4643 gnd.n4642 585
R2989 gnd.n4645 gnd.n3710 585
R2990 gnd.n3710 gnd.n3692 585
R2991 gnd.n4647 gnd.n4646 585
R2992 gnd.n4648 gnd.n4647 585
R2993 gnd.n4631 gnd.n3709 585
R2994 gnd.n3709 gnd.n3702 585
R2995 gnd.n4630 gnd.n3701 585
R2996 gnd.n4654 gnd.n3701 585
R2997 gnd.n4629 gnd.n4628 585
R2998 gnd.n4628 gnd.n3699 585
R2999 gnd.n4627 gnd.n3711 585
R3000 gnd.n4627 gnd.n4626 585
R3001 gnd.n4538 gnd.n3712 585
R3002 gnd.n3719 gnd.n3712 585
R3003 gnd.n4539 gnd.n3717 585
R3004 gnd.n4620 gnd.n3717 585
R3005 gnd.n4541 gnd.n4540 585
R3006 gnd.n4540 gnd.n3728 585
R3007 gnd.n4542 gnd.n3727 585
R3008 gnd.n4610 gnd.n3727 585
R3009 gnd.n4544 gnd.n4543 585
R3010 gnd.n4543 gnd.n3725 585
R3011 gnd.n4545 gnd.n3732 585
R3012 gnd.n4604 gnd.n3732 585
R3013 gnd.n4546 gnd.n4537 585
R3014 gnd.n4537 gnd.n4536 585
R3015 gnd.n4548 gnd.n4547 585
R3016 gnd.n4548 gnd.n3740 585
R3017 gnd.n4549 gnd.n4534 585
R3018 gnd.n4549 gnd.n3739 585
R3019 gnd.n4553 gnd.n4552 585
R3020 gnd.n4552 gnd.n4551 585
R3021 gnd.n4554 gnd.n3749 585
R3022 gnd.n4569 gnd.n3749 585
R3023 gnd.n4555 gnd.n3756 585
R3024 gnd.n3756 gnd.n3747 585
R3025 gnd.n4557 gnd.n4556 585
R3026 gnd.n4558 gnd.n4557 585
R3027 gnd.n4533 gnd.n3755 585
R3028 gnd.n3759 gnd.n3755 585
R3029 gnd.n4532 gnd.n4531 585
R3030 gnd.n4531 gnd.n4530 585
R3031 gnd.n3758 gnd.n3757 585
R3032 gnd.n4515 gnd.n3758 585
R3033 gnd.n3847 gnd.n3846 585
R3034 gnd.n4524 gnd.n3847 585
R3035 gnd.n3845 gnd.n3770 585
R3036 gnd.n3770 gnd.n3769 585
R3037 gnd.n3844 gnd.n3843 585
R3038 gnd.n3843 gnd.n2989 585
R3039 gnd.n3842 gnd.n3771 585
R3040 gnd.n3842 gnd.n2987 585
R3041 gnd.n3841 gnd.n3840 585
R3042 gnd.n3841 gnd.n2977 585
R3043 gnd.n3839 gnd.n2975 585
R3044 gnd.n5841 gnd.n2975 585
R3045 gnd.n3838 gnd.n3837 585
R3046 gnd.n3837 gnd.n2974 585
R3047 gnd.n6050 gnd.n6049 585
R3048 gnd.n6049 gnd.n6048 585
R3049 gnd.n6051 gnd.n2626 585
R3050 gnd.n6041 gnd.n2626 585
R3051 gnd.n6053 gnd.n6052 585
R3052 gnd.n6054 gnd.n6053 585
R3053 gnd.n2612 gnd.n2611 585
R3054 gnd.n4352 gnd.n2612 585
R3055 gnd.n6062 gnd.n6061 585
R3056 gnd.n6061 gnd.n6060 585
R3057 gnd.n6063 gnd.n2606 585
R3058 gnd.n4346 gnd.n2606 585
R3059 gnd.n6065 gnd.n6064 585
R3060 gnd.n6066 gnd.n6065 585
R3061 gnd.n2592 gnd.n2591 585
R3062 gnd.n4363 gnd.n2592 585
R3063 gnd.n6074 gnd.n6073 585
R3064 gnd.n6073 gnd.n6072 585
R3065 gnd.n6075 gnd.n2586 585
R3066 gnd.n4339 gnd.n2586 585
R3067 gnd.n6077 gnd.n6076 585
R3068 gnd.n6078 gnd.n6077 585
R3069 gnd.n2572 gnd.n2571 585
R3070 gnd.n4331 gnd.n2572 585
R3071 gnd.n6086 gnd.n6085 585
R3072 gnd.n6085 gnd.n6084 585
R3073 gnd.n6087 gnd.n2567 585
R3074 gnd.n4325 gnd.n2567 585
R3075 gnd.n6089 gnd.n6088 585
R3076 gnd.n6090 gnd.n6089 585
R3077 gnd.n2551 gnd.n2549 585
R3078 gnd.n4317 gnd.n2551 585
R3079 gnd.n6098 gnd.n6097 585
R3080 gnd.n6097 gnd.n6096 585
R3081 gnd.n2550 gnd.n2548 585
R3082 gnd.n4289 gnd.n2550 585
R3083 gnd.n4278 gnd.n4277 585
R3084 gnd.n4277 gnd.n4022 585
R3085 gnd.n4280 gnd.n4279 585
R3086 gnd.n4281 gnd.n4280 585
R3087 gnd.n4276 gnd.n4035 585
R3088 gnd.n4276 gnd.n4275 585
R3089 gnd.n4034 gnd.n4033 585
R3090 gnd.n4259 gnd.n4033 585
R3091 gnd.n4249 gnd.n4056 585
R3092 gnd.n4249 gnd.n4248 585
R3093 gnd.n4250 gnd.n2542 585
R3094 gnd.n4251 gnd.n4250 585
R3095 gnd.n6101 gnd.n2540 585
R3096 gnd.n4240 gnd.n2540 585
R3097 gnd.n6103 gnd.n6102 585
R3098 gnd.n6104 gnd.n6103 585
R3099 gnd.n2526 gnd.n2525 585
R3100 gnd.n4189 gnd.n2526 585
R3101 gnd.n6112 gnd.n6111 585
R3102 gnd.n6111 gnd.n6110 585
R3103 gnd.n6113 gnd.n2520 585
R3104 gnd.n4195 gnd.n2520 585
R3105 gnd.n6115 gnd.n6114 585
R3106 gnd.n6116 gnd.n6115 585
R3107 gnd.n2505 gnd.n2504 585
R3108 gnd.n4201 gnd.n2505 585
R3109 gnd.n6124 gnd.n6123 585
R3110 gnd.n6123 gnd.n6122 585
R3111 gnd.n6125 gnd.n2499 585
R3112 gnd.n4207 gnd.n2499 585
R3113 gnd.n6127 gnd.n6126 585
R3114 gnd.n6128 gnd.n6127 585
R3115 gnd.n2486 gnd.n2485 585
R3116 gnd.n4172 gnd.n2486 585
R3117 gnd.n6136 gnd.n6135 585
R3118 gnd.n6135 gnd.n6134 585
R3119 gnd.n6137 gnd.n2480 585
R3120 gnd.n2480 gnd.n2479 585
R3121 gnd.n6139 gnd.n6138 585
R3122 gnd.n6140 gnd.n6139 585
R3123 gnd.n2463 gnd.n2462 585
R3124 gnd.n2467 gnd.n2463 585
R3125 gnd.n6148 gnd.n6147 585
R3126 gnd.n6147 gnd.n6146 585
R3127 gnd.n6149 gnd.n2456 585
R3128 gnd.n2464 gnd.n2456 585
R3129 gnd.n6151 gnd.n6150 585
R3130 gnd.n6152 gnd.n6151 585
R3131 gnd.n2457 gnd.n2383 585
R3132 gnd.n2383 gnd.n2380 585
R3133 gnd.n6274 gnd.n6273 585
R3134 gnd.n6272 gnd.n2382 585
R3135 gnd.n6271 gnd.n2381 585
R3136 gnd.n6276 gnd.n2381 585
R3137 gnd.n6270 gnd.n6269 585
R3138 gnd.n6268 gnd.n6267 585
R3139 gnd.n6266 gnd.n6265 585
R3140 gnd.n6264 gnd.n6263 585
R3141 gnd.n6262 gnd.n6261 585
R3142 gnd.n6260 gnd.n6259 585
R3143 gnd.n6258 gnd.n6257 585
R3144 gnd.n6256 gnd.n6255 585
R3145 gnd.n6254 gnd.n6253 585
R3146 gnd.n6252 gnd.n6251 585
R3147 gnd.n6250 gnd.n6249 585
R3148 gnd.n6248 gnd.n6247 585
R3149 gnd.n6246 gnd.n6245 585
R3150 gnd.n6244 gnd.n6243 585
R3151 gnd.n6242 gnd.n6241 585
R3152 gnd.n6239 gnd.n6238 585
R3153 gnd.n6237 gnd.n6236 585
R3154 gnd.n6235 gnd.n6234 585
R3155 gnd.n6233 gnd.n6232 585
R3156 gnd.n6231 gnd.n6230 585
R3157 gnd.n6229 gnd.n6228 585
R3158 gnd.n6227 gnd.n6226 585
R3159 gnd.n6225 gnd.n6224 585
R3160 gnd.n6223 gnd.n6222 585
R3161 gnd.n6221 gnd.n6220 585
R3162 gnd.n6219 gnd.n6218 585
R3163 gnd.n6217 gnd.n6216 585
R3164 gnd.n6215 gnd.n6214 585
R3165 gnd.n6213 gnd.n6212 585
R3166 gnd.n6211 gnd.n6210 585
R3167 gnd.n6209 gnd.n6208 585
R3168 gnd.n6207 gnd.n6206 585
R3169 gnd.n6205 gnd.n6204 585
R3170 gnd.n6203 gnd.n6202 585
R3171 gnd.n6201 gnd.n6200 585
R3172 gnd.n6199 gnd.n6198 585
R3173 gnd.n6197 gnd.n6196 585
R3174 gnd.n6195 gnd.n6194 585
R3175 gnd.n6193 gnd.n6192 585
R3176 gnd.n6191 gnd.n6190 585
R3177 gnd.n6189 gnd.n6188 585
R3178 gnd.n6187 gnd.n6186 585
R3179 gnd.n6185 gnd.n6184 585
R3180 gnd.n6183 gnd.n6182 585
R3181 gnd.n6181 gnd.n6180 585
R3182 gnd.n6179 gnd.n6178 585
R3183 gnd.n6177 gnd.n6176 585
R3184 gnd.n6175 gnd.n6174 585
R3185 gnd.n6173 gnd.n6172 585
R3186 gnd.n6171 gnd.n6170 585
R3187 gnd.n6169 gnd.n6168 585
R3188 gnd.n6167 gnd.n6166 585
R3189 gnd.n6165 gnd.n6164 585
R3190 gnd.n6163 gnd.n6162 585
R3191 gnd.n6161 gnd.n6160 585
R3192 gnd.n2452 gnd.n2445 585
R3193 gnd.n2843 gnd.n2842 585
R3194 gnd.n2849 gnd.n2848 585
R3195 gnd.n2851 gnd.n2850 585
R3196 gnd.n2853 gnd.n2852 585
R3197 gnd.n2855 gnd.n2854 585
R3198 gnd.n2857 gnd.n2856 585
R3199 gnd.n2859 gnd.n2858 585
R3200 gnd.n2861 gnd.n2860 585
R3201 gnd.n2863 gnd.n2862 585
R3202 gnd.n2865 gnd.n2864 585
R3203 gnd.n2867 gnd.n2866 585
R3204 gnd.n2869 gnd.n2868 585
R3205 gnd.n2871 gnd.n2870 585
R3206 gnd.n2873 gnd.n2872 585
R3207 gnd.n2875 gnd.n2874 585
R3208 gnd.n2877 gnd.n2876 585
R3209 gnd.n2879 gnd.n2878 585
R3210 gnd.n2881 gnd.n2880 585
R3211 gnd.n2883 gnd.n2882 585
R3212 gnd.n2886 gnd.n2885 585
R3213 gnd.n2884 gnd.n2822 585
R3214 gnd.n2891 gnd.n2890 585
R3215 gnd.n2893 gnd.n2892 585
R3216 gnd.n2895 gnd.n2894 585
R3217 gnd.n2897 gnd.n2896 585
R3218 gnd.n2899 gnd.n2898 585
R3219 gnd.n2901 gnd.n2900 585
R3220 gnd.n2903 gnd.n2902 585
R3221 gnd.n2905 gnd.n2904 585
R3222 gnd.n2908 gnd.n2907 585
R3223 gnd.n2906 gnd.n2813 585
R3224 gnd.n5917 gnd.n5916 585
R3225 gnd.n5919 gnd.n5918 585
R3226 gnd.n5921 gnd.n5920 585
R3227 gnd.n5923 gnd.n5922 585
R3228 gnd.n5925 gnd.n5924 585
R3229 gnd.n5927 gnd.n5926 585
R3230 gnd.n5929 gnd.n5928 585
R3231 gnd.n5931 gnd.n5930 585
R3232 gnd.n5934 gnd.n5933 585
R3233 gnd.n5936 gnd.n5935 585
R3234 gnd.n5938 gnd.n5937 585
R3235 gnd.n5940 gnd.n5939 585
R3236 gnd.n5942 gnd.n5941 585
R3237 gnd.n5944 gnd.n5943 585
R3238 gnd.n5946 gnd.n5945 585
R3239 gnd.n5948 gnd.n5947 585
R3240 gnd.n5950 gnd.n5949 585
R3241 gnd.n5952 gnd.n5951 585
R3242 gnd.n5954 gnd.n5953 585
R3243 gnd.n5956 gnd.n5955 585
R3244 gnd.n5958 gnd.n5957 585
R3245 gnd.n5960 gnd.n5959 585
R3246 gnd.n5961 gnd.n2782 585
R3247 gnd.n5963 gnd.n5962 585
R3248 gnd.n2783 gnd.n2781 585
R3249 gnd.n2784 gnd.n2631 585
R3250 gnd.n5965 gnd.n2631 585
R3251 gnd.n6044 gnd.n2633 585
R3252 gnd.n6048 gnd.n2633 585
R3253 gnd.n6043 gnd.n6042 585
R3254 gnd.n6042 gnd.n6041 585
R3255 gnd.n2639 gnd.n2624 585
R3256 gnd.n6054 gnd.n2624 585
R3257 gnd.n4351 gnd.n4350 585
R3258 gnd.n4352 gnd.n4351 585
R3259 gnd.n4349 gnd.n2614 585
R3260 gnd.n6060 gnd.n2614 585
R3261 gnd.n4348 gnd.n4347 585
R3262 gnd.n4347 gnd.n4346 585
R3263 gnd.n4344 gnd.n2603 585
R3264 gnd.n6066 gnd.n2603 585
R3265 gnd.n4343 gnd.n3999 585
R3266 gnd.n4363 gnd.n3999 585
R3267 gnd.n4342 gnd.n2594 585
R3268 gnd.n6072 gnd.n2594 585
R3269 gnd.n4341 gnd.n4340 585
R3270 gnd.n4340 gnd.n4339 585
R3271 gnd.n4005 gnd.n2583 585
R3272 gnd.n6078 gnd.n2583 585
R3273 gnd.n4330 gnd.n4329 585
R3274 gnd.n4331 gnd.n4330 585
R3275 gnd.n4328 gnd.n2574 585
R3276 gnd.n6084 gnd.n2574 585
R3277 gnd.n4327 gnd.n4326 585
R3278 gnd.n4326 gnd.n4325 585
R3279 gnd.n4011 gnd.n2564 585
R3280 gnd.n6090 gnd.n2564 585
R3281 gnd.n4264 gnd.n4016 585
R3282 gnd.n4317 gnd.n4016 585
R3283 gnd.n4265 gnd.n2553 585
R3284 gnd.n6096 gnd.n2553 585
R3285 gnd.n4266 gnd.n4023 585
R3286 gnd.n4289 gnd.n4023 585
R3287 gnd.n4268 gnd.n4267 585
R3288 gnd.n4267 gnd.n4022 585
R3289 gnd.n4263 gnd.n4030 585
R3290 gnd.n4281 gnd.n4030 585
R3291 gnd.n4262 gnd.n4037 585
R3292 gnd.n4275 gnd.n4037 585
R3293 gnd.n4261 gnd.n4260 585
R3294 gnd.n4260 gnd.n4259 585
R3295 gnd.n4045 gnd.n4043 585
R3296 gnd.n4248 gnd.n4045 585
R3297 gnd.n4243 gnd.n4053 585
R3298 gnd.n4251 gnd.n4053 585
R3299 gnd.n4242 gnd.n4241 585
R3300 gnd.n4241 gnd.n4240 585
R3301 gnd.n4059 gnd.n2538 585
R3302 gnd.n6104 gnd.n2538 585
R3303 gnd.n4188 gnd.n4187 585
R3304 gnd.n4189 gnd.n4188 585
R3305 gnd.n4180 gnd.n2528 585
R3306 gnd.n6110 gnd.n2528 585
R3307 gnd.n4197 gnd.n4196 585
R3308 gnd.n4196 gnd.n4195 585
R3309 gnd.n4198 gnd.n2517 585
R3310 gnd.n6116 gnd.n2517 585
R3311 gnd.n4200 gnd.n4199 585
R3312 gnd.n4201 gnd.n4200 585
R3313 gnd.n4178 gnd.n2507 585
R3314 gnd.n6122 gnd.n2507 585
R3315 gnd.n4177 gnd.n4074 585
R3316 gnd.n4207 gnd.n4074 585
R3317 gnd.n4175 gnd.n2497 585
R3318 gnd.n6128 gnd.n2497 585
R3319 gnd.n4174 gnd.n4173 585
R3320 gnd.n4173 gnd.n4172 585
R3321 gnd.n4089 gnd.n2487 585
R3322 gnd.n6134 gnd.n2487 585
R3323 gnd.n4088 gnd.n4087 585
R3324 gnd.n4087 gnd.n2479 585
R3325 gnd.n4085 gnd.n2477 585
R3326 gnd.n6140 gnd.n2477 585
R3327 gnd.n4084 gnd.n4083 585
R3328 gnd.n4083 gnd.n2467 585
R3329 gnd.n4082 gnd.n2465 585
R3330 gnd.n6146 gnd.n2465 585
R3331 gnd.n4081 gnd.n2453 585
R3332 gnd.n2464 gnd.n2453 585
R3333 gnd.n6153 gnd.n2451 585
R3334 gnd.n6153 gnd.n6152 585
R3335 gnd.n6155 gnd.n6154 585
R3336 gnd.n6154 gnd.n2380 585
R3337 gnd.n7359 gnd.n7358 585
R3338 gnd.n7358 gnd.n7357 585
R3339 gnd.n7360 gnd.n162 585
R3340 gnd.n168 gnd.n162 585
R3341 gnd.n7362 gnd.n7361 585
R3342 gnd.n7363 gnd.n7362 585
R3343 gnd.n150 gnd.n149 585
R3344 gnd.n153 gnd.n150 585
R3345 gnd.n7371 gnd.n7370 585
R3346 gnd.n7370 gnd.n7369 585
R3347 gnd.n7372 gnd.n144 585
R3348 gnd.n144 gnd.n143 585
R3349 gnd.n7374 gnd.n7373 585
R3350 gnd.n7375 gnd.n7374 585
R3351 gnd.n130 gnd.n129 585
R3352 gnd.n7340 gnd.n130 585
R3353 gnd.n7383 gnd.n7382 585
R3354 gnd.n7382 gnd.n7381 585
R3355 gnd.n7384 gnd.n124 585
R3356 gnd.n7248 gnd.n124 585
R3357 gnd.n7386 gnd.n7385 585
R3358 gnd.n7387 gnd.n7386 585
R3359 gnd.n110 gnd.n109 585
R3360 gnd.n7241 gnd.n110 585
R3361 gnd.n7395 gnd.n7394 585
R3362 gnd.n7394 gnd.n7393 585
R3363 gnd.n7396 gnd.n105 585
R3364 gnd.n7233 gnd.n105 585
R3365 gnd.n7398 gnd.n7397 585
R3366 gnd.n7399 gnd.n7398 585
R3367 gnd.n89 gnd.n87 585
R3368 gnd.n7226 gnd.n89 585
R3369 gnd.n7407 gnd.n7406 585
R3370 gnd.n7406 gnd.n7405 585
R3371 gnd.n88 gnd.n80 585
R3372 gnd.n5442 gnd.n88 585
R3373 gnd.n7410 gnd.n78 585
R3374 gnd.n5452 gnd.n78 585
R3375 gnd.n7412 gnd.n7411 585
R3376 gnd.n7413 gnd.n7412 585
R3377 gnd.n3375 gnd.n77 585
R3378 gnd.n5458 gnd.n77 585
R3379 gnd.n3377 gnd.n3376 585
R3380 gnd.n3378 gnd.n3377 585
R3381 gnd.n3366 gnd.n3365 585
R3382 gnd.n5424 gnd.n3365 585
R3383 gnd.n5468 gnd.n3367 585
R3384 gnd.n5468 gnd.n5467 585
R3385 gnd.n5471 gnd.n5470 585
R3386 gnd.n5472 gnd.n5471 585
R3387 gnd.n5469 gnd.n3350 585
R3388 gnd.n5415 gnd.n3350 585
R3389 gnd.n5480 gnd.n5479 585
R3390 gnd.n5479 gnd.n5478 585
R3391 gnd.n5481 gnd.n3347 585
R3392 gnd.n5403 gnd.n3347 585
R3393 gnd.n5483 gnd.n5482 585
R3394 gnd.n5484 gnd.n5483 585
R3395 gnd.n3334 gnd.n3333 585
R3396 gnd.n5396 gnd.n3334 585
R3397 gnd.n5492 gnd.n5491 585
R3398 gnd.n5491 gnd.n5490 585
R3399 gnd.n5493 gnd.n3328 585
R3400 gnd.n5388 gnd.n3328 585
R3401 gnd.n5495 gnd.n5494 585
R3402 gnd.n5496 gnd.n5495 585
R3403 gnd.n3313 gnd.n3312 585
R3404 gnd.n5328 gnd.n3313 585
R3405 gnd.n5504 gnd.n5503 585
R3406 gnd.n5503 gnd.n5502 585
R3407 gnd.n5505 gnd.n3307 585
R3408 gnd.n5319 gnd.n3307 585
R3409 gnd.n5507 gnd.n5506 585
R3410 gnd.n5508 gnd.n5507 585
R3411 gnd.n3290 gnd.n3289 585
R3412 gnd.n5313 gnd.n3290 585
R3413 gnd.n5516 gnd.n5515 585
R3414 gnd.n5515 gnd.n5514 585
R3415 gnd.n5517 gnd.n3281 585
R3416 gnd.n5306 gnd.n3281 585
R3417 gnd.n5519 gnd.n5518 585
R3418 gnd.n5520 gnd.n5519 585
R3419 gnd.n3282 gnd.n3280 585
R3420 gnd.n5345 gnd.n3280 585
R3421 gnd.n3283 gnd.n3202 585
R3422 gnd.n5528 gnd.n3202 585
R3423 gnd.n5647 gnd.n5646 585
R3424 gnd.n5645 gnd.n3201 585
R3425 gnd.n5644 gnd.n3200 585
R3426 gnd.n5649 gnd.n3200 585
R3427 gnd.n5643 gnd.n5642 585
R3428 gnd.n5641 gnd.n5640 585
R3429 gnd.n5639 gnd.n5638 585
R3430 gnd.n5637 gnd.n5636 585
R3431 gnd.n5635 gnd.n5634 585
R3432 gnd.n5633 gnd.n5632 585
R3433 gnd.n5631 gnd.n5630 585
R3434 gnd.n5629 gnd.n5628 585
R3435 gnd.n5627 gnd.n5626 585
R3436 gnd.n5625 gnd.n5624 585
R3437 gnd.n5623 gnd.n5622 585
R3438 gnd.n5621 gnd.n5620 585
R3439 gnd.n5619 gnd.n5618 585
R3440 gnd.n5617 gnd.n5616 585
R3441 gnd.n5615 gnd.n5614 585
R3442 gnd.n5612 gnd.n5611 585
R3443 gnd.n5610 gnd.n5609 585
R3444 gnd.n5608 gnd.n5607 585
R3445 gnd.n5606 gnd.n5605 585
R3446 gnd.n5604 gnd.n5603 585
R3447 gnd.n5602 gnd.n5601 585
R3448 gnd.n5600 gnd.n5599 585
R3449 gnd.n5598 gnd.n5597 585
R3450 gnd.n5595 gnd.n5594 585
R3451 gnd.n5593 gnd.n5592 585
R3452 gnd.n5591 gnd.n5590 585
R3453 gnd.n5589 gnd.n5588 585
R3454 gnd.n5587 gnd.n5586 585
R3455 gnd.n5585 gnd.n5584 585
R3456 gnd.n5583 gnd.n5582 585
R3457 gnd.n5581 gnd.n5580 585
R3458 gnd.n5579 gnd.n5578 585
R3459 gnd.n5577 gnd.n5576 585
R3460 gnd.n5575 gnd.n5574 585
R3461 gnd.n5573 gnd.n5572 585
R3462 gnd.n5571 gnd.n5570 585
R3463 gnd.n5569 gnd.n5568 585
R3464 gnd.n5567 gnd.n5566 585
R3465 gnd.n5565 gnd.n5564 585
R3466 gnd.n5563 gnd.n5562 585
R3467 gnd.n5561 gnd.n5560 585
R3468 gnd.n5559 gnd.n5558 585
R3469 gnd.n5557 gnd.n5556 585
R3470 gnd.n5555 gnd.n5554 585
R3471 gnd.n5553 gnd.n5552 585
R3472 gnd.n5551 gnd.n5550 585
R3473 gnd.n5549 gnd.n5548 585
R3474 gnd.n5547 gnd.n5546 585
R3475 gnd.n5545 gnd.n5544 585
R3476 gnd.n5543 gnd.n5542 585
R3477 gnd.n5541 gnd.n5540 585
R3478 gnd.n5539 gnd.n5538 585
R3479 gnd.n5537 gnd.n5536 585
R3480 gnd.n5531 gnd.n5530 585
R3481 gnd.n384 gnd.n383 585
R3482 gnd.n381 gnd.n177 585
R3483 gnd.n380 gnd.n379 585
R3484 gnd.n373 gnd.n179 585
R3485 gnd.n375 gnd.n374 585
R3486 gnd.n371 gnd.n181 585
R3487 gnd.n370 gnd.n369 585
R3488 gnd.n363 gnd.n183 585
R3489 gnd.n365 gnd.n364 585
R3490 gnd.n361 gnd.n185 585
R3491 gnd.n360 gnd.n359 585
R3492 gnd.n353 gnd.n187 585
R3493 gnd.n355 gnd.n354 585
R3494 gnd.n351 gnd.n189 585
R3495 gnd.n350 gnd.n349 585
R3496 gnd.n343 gnd.n191 585
R3497 gnd.n345 gnd.n344 585
R3498 gnd.n341 gnd.n193 585
R3499 gnd.n340 gnd.n339 585
R3500 gnd.n333 gnd.n195 585
R3501 gnd.n335 gnd.n334 585
R3502 gnd.n331 gnd.n199 585
R3503 gnd.n330 gnd.n329 585
R3504 gnd.n323 gnd.n201 585
R3505 gnd.n325 gnd.n324 585
R3506 gnd.n321 gnd.n203 585
R3507 gnd.n320 gnd.n319 585
R3508 gnd.n313 gnd.n205 585
R3509 gnd.n315 gnd.n314 585
R3510 gnd.n311 gnd.n207 585
R3511 gnd.n310 gnd.n309 585
R3512 gnd.n303 gnd.n209 585
R3513 gnd.n305 gnd.n304 585
R3514 gnd.n301 gnd.n211 585
R3515 gnd.n300 gnd.n299 585
R3516 gnd.n293 gnd.n213 585
R3517 gnd.n295 gnd.n294 585
R3518 gnd.n291 gnd.n215 585
R3519 gnd.n290 gnd.n289 585
R3520 gnd.n283 gnd.n217 585
R3521 gnd.n285 gnd.n284 585
R3522 gnd.n281 gnd.n280 585
R3523 gnd.n279 gnd.n222 585
R3524 gnd.n273 gnd.n223 585
R3525 gnd.n275 gnd.n274 585
R3526 gnd.n270 gnd.n225 585
R3527 gnd.n269 gnd.n268 585
R3528 gnd.n262 gnd.n227 585
R3529 gnd.n264 gnd.n263 585
R3530 gnd.n260 gnd.n229 585
R3531 gnd.n259 gnd.n258 585
R3532 gnd.n252 gnd.n231 585
R3533 gnd.n254 gnd.n253 585
R3534 gnd.n250 gnd.n233 585
R3535 gnd.n249 gnd.n248 585
R3536 gnd.n242 gnd.n235 585
R3537 gnd.n244 gnd.n243 585
R3538 gnd.n240 gnd.n239 585
R3539 gnd.n238 gnd.n167 585
R3540 gnd.n171 gnd.n167 585
R3541 gnd.n7353 gnd.n169 585
R3542 gnd.n7357 gnd.n169 585
R3543 gnd.n7352 gnd.n7351 585
R3544 gnd.n7351 gnd.n168 585
R3545 gnd.n7350 gnd.n160 585
R3546 gnd.n7363 gnd.n160 585
R3547 gnd.n7349 gnd.n7348 585
R3548 gnd.n7348 gnd.n153 585
R3549 gnd.n7347 gnd.n151 585
R3550 gnd.n7369 gnd.n151 585
R3551 gnd.n7346 gnd.n7345 585
R3552 gnd.n7345 gnd.n143 585
R3553 gnd.n7343 gnd.n141 585
R3554 gnd.n7375 gnd.n141 585
R3555 gnd.n7342 gnd.n7341 585
R3556 gnd.n7341 gnd.n7340 585
R3557 gnd.n387 gnd.n132 585
R3558 gnd.n7381 gnd.n132 585
R3559 gnd.n7247 gnd.n7246 585
R3560 gnd.n7248 gnd.n7247 585
R3561 gnd.n7244 gnd.n121 585
R3562 gnd.n7387 gnd.n121 585
R3563 gnd.n7243 gnd.n7242 585
R3564 gnd.n7242 gnd.n7241 585
R3565 gnd.n391 gnd.n112 585
R3566 gnd.n7393 gnd.n112 585
R3567 gnd.n7232 gnd.n7231 585
R3568 gnd.n7233 gnd.n7232 585
R3569 gnd.n7229 gnd.n102 585
R3570 gnd.n7399 gnd.n102 585
R3571 gnd.n7228 gnd.n7227 585
R3572 gnd.n7227 gnd.n7226 585
R3573 gnd.n396 gnd.n91 585
R3574 gnd.n7405 gnd.n91 585
R3575 gnd.n5433 gnd.n5432 585
R3576 gnd.n5442 gnd.n5433 585
R3577 gnd.n5430 gnd.n3385 585
R3578 gnd.n5452 gnd.n3385 585
R3579 gnd.n5429 gnd.n74 585
R3580 gnd.n7413 gnd.n74 585
R3581 gnd.n5428 gnd.n3379 585
R3582 gnd.n5458 gnd.n3379 585
R3583 gnd.n5427 gnd.n5426 585
R3584 gnd.n5426 gnd.n3378 585
R3585 gnd.n5425 gnd.n3386 585
R3586 gnd.n5425 gnd.n5424 585
R3587 gnd.n5419 gnd.n3368 585
R3588 gnd.n5467 gnd.n3368 585
R3589 gnd.n5418 gnd.n3362 585
R3590 gnd.n5472 gnd.n3362 585
R3591 gnd.n5417 gnd.n5416 585
R3592 gnd.n5416 gnd.n5415 585
R3593 gnd.n3391 gnd.n3352 585
R3594 gnd.n5478 gnd.n3352 585
R3595 gnd.n5402 gnd.n5401 585
R3596 gnd.n5403 gnd.n5402 585
R3597 gnd.n5399 gnd.n3345 585
R3598 gnd.n5484 gnd.n3345 585
R3599 gnd.n5398 gnd.n5397 585
R3600 gnd.n5397 gnd.n5396 585
R3601 gnd.n3397 gnd.n3335 585
R3602 gnd.n5490 gnd.n3335 585
R3603 gnd.n5324 gnd.n3401 585
R3604 gnd.n5388 gnd.n3401 585
R3605 gnd.n5325 gnd.n3325 585
R3606 gnd.n5496 gnd.n3325 585
R3607 gnd.n5327 gnd.n5326 585
R3608 gnd.n5328 gnd.n5327 585
R3609 gnd.n5322 gnd.n3315 585
R3610 gnd.n5502 gnd.n3315 585
R3611 gnd.n5321 gnd.n5320 585
R3612 gnd.n5320 gnd.n5319 585
R3613 gnd.n5316 gnd.n3305 585
R3614 gnd.n5508 gnd.n3305 585
R3615 gnd.n5315 gnd.n5314 585
R3616 gnd.n5314 gnd.n5313 585
R3617 gnd.n5312 gnd.n3292 585
R3618 gnd.n5514 gnd.n3292 585
R3619 gnd.n3276 gnd.n3275 585
R3620 gnd.n5306 gnd.n3276 585
R3621 gnd.n5522 gnd.n5521 585
R3622 gnd.n5521 gnd.n5520 585
R3623 gnd.n5523 gnd.n3265 585
R3624 gnd.n5345 gnd.n3265 585
R3625 gnd.n5529 gnd.n3266 585
R3626 gnd.n5529 gnd.n5528 585
R3627 gnd.n977 gnd.n976 585
R3628 gnd.n2489 gnd.n977 585
R3629 gnd.n7213 gnd.n7212 585
R3630 gnd.n7213 gnd.n134 585
R3631 gnd.n7215 gnd.n7214 585
R3632 gnd.n7214 gnd.n131 585
R3633 gnd.n7216 gnd.n406 585
R3634 gnd.n406 gnd.n123 585
R3635 gnd.n7218 gnd.n7217 585
R3636 gnd.n7218 gnd.n120 585
R3637 gnd.n7219 gnd.n405 585
R3638 gnd.n7219 gnd.n392 585
R3639 gnd.n7221 gnd.n7220 585
R3640 gnd.n7220 gnd.n111 585
R3641 gnd.n7222 gnd.n399 585
R3642 gnd.n399 gnd.n104 585
R3643 gnd.n7224 gnd.n7223 585
R3644 gnd.n7225 gnd.n7224 585
R3645 gnd.n400 gnd.n398 585
R3646 gnd.n398 gnd.n93 585
R3647 gnd.n5447 gnd.n5444 585
R3648 gnd.n5444 gnd.n90 585
R3649 gnd.n5450 gnd.n5449 585
R3650 gnd.n5451 gnd.n5450 585
R3651 gnd.n5446 gnd.n5443 585
R3652 gnd.n5443 gnd.n75 585
R3653 gnd.n3374 gnd.n3373 585
R3654 gnd.n3374 gnd.n73 585
R3655 gnd.n5461 gnd.n5460 585
R3656 gnd.n5460 gnd.n5459 585
R3657 gnd.n5463 gnd.n3371 585
R3658 gnd.n3390 gnd.n3371 585
R3659 gnd.n5465 gnd.n5464 585
R3660 gnd.n5466 gnd.n5465 585
R3661 gnd.n5374 gnd.n3370 585
R3662 gnd.n3370 gnd.n3364 585
R3663 gnd.n5376 gnd.n5375 585
R3664 gnd.n5375 gnd.n3361 585
R3665 gnd.n5378 gnd.n5371 585
R3666 gnd.n5371 gnd.n3354 585
R3667 gnd.n5380 gnd.n5379 585
R3668 gnd.n5380 gnd.n3351 585
R3669 gnd.n5381 gnd.n5370 585
R3670 gnd.n5381 gnd.n3396 585
R3671 gnd.n5383 gnd.n5382 585
R3672 gnd.n5382 gnd.n3344 585
R3673 gnd.n5384 gnd.n3403 585
R3674 gnd.n3403 gnd.n3337 585
R3675 gnd.n5386 gnd.n5385 585
R3676 gnd.n5387 gnd.n5386 585
R3677 gnd.n3404 gnd.n3402 585
R3678 gnd.n3402 gnd.n3327 585
R3679 gnd.n5364 gnd.n5363 585
R3680 gnd.n5363 gnd.n3324 585
R3681 gnd.n5362 gnd.n3406 585
R3682 gnd.n5362 gnd.n3317 585
R3683 gnd.n5361 gnd.n5360 585
R3684 gnd.n5361 gnd.n3314 585
R3685 gnd.n3408 gnd.n3407 585
R3686 gnd.n5318 gnd.n3407 585
R3687 gnd.n5356 gnd.n5355 585
R3688 gnd.n5355 gnd.n3304 585
R3689 gnd.n5354 gnd.n3410 585
R3690 gnd.n5354 gnd.n3294 585
R3691 gnd.n5353 gnd.n5352 585
R3692 gnd.n5353 gnd.n3291 585
R3693 gnd.n3412 gnd.n3411 585
R3694 gnd.n3411 gnd.n3278 585
R3695 gnd.n5348 gnd.n5347 585
R3696 gnd.n5347 gnd.n5346 585
R3697 gnd.n3415 gnd.n3414 585
R3698 gnd.n3415 gnd.n3269 585
R3699 gnd.n5289 gnd.n5288 585
R3700 gnd.n5289 gnd.n3267 585
R3701 gnd.n5290 gnd.n5285 585
R3702 gnd.n5290 gnd.n3199 585
R3703 gnd.n5292 gnd.n5291 585
R3704 gnd.n5291 gnd.n3157 585
R3705 gnd.n5293 gnd.n3447 585
R3706 gnd.n3447 gnd.n3445 585
R3707 gnd.n5295 gnd.n5294 585
R3708 gnd.n5296 gnd.n5295 585
R3709 gnd.n3448 gnd.n3446 585
R3710 gnd.n3446 gnd.n3090 585
R3711 gnd.n5279 gnd.n3089 585
R3712 gnd.n5717 gnd.n3089 585
R3713 gnd.n5278 gnd.n5277 585
R3714 gnd.n5277 gnd.n3088 585
R3715 gnd.n5276 gnd.n3450 585
R3716 gnd.n5276 gnd.n5275 585
R3717 gnd.n5263 gnd.n3451 585
R3718 gnd.n3452 gnd.n3451 585
R3719 gnd.n5265 gnd.n5264 585
R3720 gnd.n5266 gnd.n5265 585
R3721 gnd.n3460 gnd.n3459 585
R3722 gnd.n3459 gnd.n3458 585
R3723 gnd.n5257 gnd.n5256 585
R3724 gnd.n5256 gnd.n5255 585
R3725 gnd.n3463 gnd.n3462 585
R3726 gnd.n3470 gnd.n3463 585
R3727 gnd.n5245 gnd.n5244 585
R3728 gnd.n5246 gnd.n5245 585
R3729 gnd.n3472 gnd.n3471 585
R3730 gnd.n3471 gnd.n3469 585
R3731 gnd.n5240 gnd.n5239 585
R3732 gnd.n5239 gnd.n5238 585
R3733 gnd.n3475 gnd.n3474 585
R3734 gnd.n3476 gnd.n3475 585
R3735 gnd.n5228 gnd.n5227 585
R3736 gnd.n5229 gnd.n5228 585
R3737 gnd.n3484 gnd.n3483 585
R3738 gnd.n3483 gnd.n3482 585
R3739 gnd.n5223 gnd.n5222 585
R3740 gnd.n5222 gnd.n5221 585
R3741 gnd.n3487 gnd.n3486 585
R3742 gnd.n3488 gnd.n3487 585
R3743 gnd.n5211 gnd.n5210 585
R3744 gnd.n5212 gnd.n5211 585
R3745 gnd.n3496 gnd.n3495 585
R3746 gnd.n3495 gnd.n3494 585
R3747 gnd.n5206 gnd.n5205 585
R3748 gnd.n5205 gnd.n5204 585
R3749 gnd.n3499 gnd.n3498 585
R3750 gnd.n3500 gnd.n3499 585
R3751 gnd.n5194 gnd.n5193 585
R3752 gnd.n5195 gnd.n5194 585
R3753 gnd.n3507 gnd.n3506 585
R3754 gnd.n5185 gnd.n3506 585
R3755 gnd.n5189 gnd.n5188 585
R3756 gnd.n5188 gnd.n5187 585
R3757 gnd.n3510 gnd.n3509 585
R3758 gnd.n3532 gnd.n3510 585
R3759 gnd.n5176 gnd.n5175 585
R3760 gnd.n5177 gnd.n5176 585
R3761 gnd.n3519 gnd.n3518 585
R3762 gnd.n3526 gnd.n3518 585
R3763 gnd.n5171 gnd.n5170 585
R3764 gnd.n5170 gnd.n5169 585
R3765 gnd.n3522 gnd.n3521 585
R3766 gnd.t144 gnd.n3522 585
R3767 gnd.n4945 gnd.n3549 585
R3768 gnd.n3549 gnd.n3541 585
R3769 gnd.n4947 gnd.n4946 585
R3770 gnd.n4948 gnd.n4947 585
R3771 gnd.n3550 gnd.n3548 585
R3772 gnd.n4913 gnd.n3548 585
R3773 gnd.n4940 gnd.n4939 585
R3774 gnd.n4939 gnd.n4938 585
R3775 gnd.n3553 gnd.n3552 585
R3776 gnd.n4930 gnd.n3553 585
R3777 gnd.n4889 gnd.n3578 585
R3778 gnd.n3578 gnd.n3569 585
R3779 gnd.n4891 gnd.n4890 585
R3780 gnd.n4892 gnd.n4891 585
R3781 gnd.n3579 gnd.n3577 585
R3782 gnd.n3577 gnd.n3573 585
R3783 gnd.n4884 gnd.n4883 585
R3784 gnd.n4883 gnd.n4882 585
R3785 gnd.n3582 gnd.n3581 585
R3786 gnd.n4794 gnd.n3582 585
R3787 gnd.n4864 gnd.n4863 585
R3788 gnd.n4865 gnd.n4864 585
R3789 gnd.n3597 gnd.n3596 585
R3790 gnd.n3603 gnd.n3596 585
R3791 gnd.n4859 gnd.n4858 585
R3792 gnd.n4858 gnd.n4857 585
R3793 gnd.n3600 gnd.n3599 585
R3794 gnd.n3607 gnd.n3600 585
R3795 gnd.n4836 gnd.n4835 585
R3796 gnd.n4837 gnd.n4836 585
R3797 gnd.n3615 gnd.n3614 585
R3798 gnd.n4788 gnd.n3614 585
R3799 gnd.n4831 gnd.n4830 585
R3800 gnd.n4830 gnd.n4829 585
R3801 gnd.n3618 gnd.n3617 585
R3802 gnd.n4818 gnd.n3618 585
R3803 gnd.n4776 gnd.n4775 585
R3804 gnd.n4777 gnd.n4776 585
R3805 gnd.n3637 gnd.n3636 585
R3806 gnd.n4679 gnd.n3636 585
R3807 gnd.n4771 gnd.n4770 585
R3808 gnd.n4770 gnd.n4769 585
R3809 gnd.n3640 gnd.n3639 585
R3810 gnd.n4758 gnd.n3640 585
R3811 gnd.n4719 gnd.n4718 585
R3812 gnd.n4719 gnd.n3655 585
R3813 gnd.n4720 gnd.n4715 585
R3814 gnd.n4720 gnd.n3653 585
R3815 gnd.n4722 gnd.n4721 585
R3816 gnd.n4721 gnd.n3659 585
R3817 gnd.n4723 gnd.n3674 585
R3818 gnd.n3674 gnd.n3665 585
R3819 gnd.n4725 gnd.n4724 585
R3820 gnd.n4726 gnd.n4725 585
R3821 gnd.n3675 gnd.n3673 585
R3822 gnd.n3673 gnd.n3669 585
R3823 gnd.n4709 gnd.n4708 585
R3824 gnd.n4708 gnd.n4707 585
R3825 gnd.n3678 gnd.n3677 585
R3826 gnd.n4699 gnd.n3678 585
R3827 gnd.n4662 gnd.n3694 585
R3828 gnd.n4641 gnd.n3694 585
R3829 gnd.n4664 gnd.n4663 585
R3830 gnd.n4665 gnd.n4664 585
R3831 gnd.n3695 gnd.n3693 585
R3832 gnd.n3708 gnd.n3693 585
R3833 gnd.n4657 gnd.n4656 585
R3834 gnd.n4656 gnd.n4655 585
R3835 gnd.n3698 gnd.n3697 585
R3836 gnd.n4589 gnd.n3698 585
R3837 gnd.n4618 gnd.n4617 585
R3838 gnd.n4619 gnd.n4618 585
R3839 gnd.n3721 gnd.n3720 585
R3840 gnd.n3720 gnd.n3716 585
R3841 gnd.n4613 gnd.n4612 585
R3842 gnd.n4612 gnd.n4611 585
R3843 gnd.n3724 gnd.n3723 585
R3844 gnd.n4603 gnd.n3724 585
R3845 gnd.n4578 gnd.n3742 585
R3846 gnd.n4535 gnd.n3742 585
R3847 gnd.n4580 gnd.n4579 585
R3848 gnd.n4581 gnd.n4580 585
R3849 gnd.n3743 gnd.n3741 585
R3850 gnd.n4550 gnd.n3741 585
R3851 gnd.n4573 gnd.n4572 585
R3852 gnd.n4572 gnd.n4571 585
R3853 gnd.n3746 gnd.n3745 585
R3854 gnd.n3754 gnd.n3746 585
R3855 gnd.n4520 gnd.n4516 585
R3856 gnd.n4516 gnd.n3760 585
R3857 gnd.n4522 gnd.n4521 585
R3858 gnd.n4523 gnd.n4522 585
R3859 gnd.n2986 gnd.n2985 585
R3860 gnd.n3768 gnd.n2986 585
R3861 gnd.n5836 gnd.n5835 585
R3862 gnd.n5835 gnd.n5834 585
R3863 gnd.n5837 gnd.n2980 585
R3864 gnd.n4500 gnd.n2980 585
R3865 gnd.n5839 gnd.n5838 585
R3866 gnd.n5840 gnd.n5839 585
R3867 gnd.n2981 gnd.n2979 585
R3868 gnd.n2979 gnd.n2948 585
R3869 gnd.n4488 gnd.n3859 585
R3870 gnd.n3859 gnd.n2916 585
R3871 gnd.n4490 gnd.n4489 585
R3872 gnd.n4491 gnd.n4490 585
R3873 gnd.n3860 gnd.n3858 585
R3874 gnd.n3866 gnd.n3858 585
R3875 gnd.n4482 gnd.n4481 585
R3876 gnd.n4481 gnd.n4480 585
R3877 gnd.n3863 gnd.n3862 585
R3878 gnd.n3864 gnd.n3863 585
R3879 gnd.n4460 gnd.n4459 585
R3880 gnd.n4461 gnd.n4460 585
R3881 gnd.n3877 gnd.n3876 585
R3882 gnd.n3876 gnd.n3874 585
R3883 gnd.n4455 gnd.n4454 585
R3884 gnd.n4454 gnd.n4453 585
R3885 gnd.n3880 gnd.n3879 585
R3886 gnd.n3881 gnd.n3880 585
R3887 gnd.n4444 gnd.n4443 585
R3888 gnd.n4445 gnd.n4444 585
R3889 gnd.n3891 gnd.n3890 585
R3890 gnd.n3890 gnd.n3888 585
R3891 gnd.n4439 gnd.n4438 585
R3892 gnd.n4438 gnd.n4437 585
R3893 gnd.n3894 gnd.n3893 585
R3894 gnd.n3895 gnd.n3894 585
R3895 gnd.n4428 gnd.n4427 585
R3896 gnd.n4429 gnd.n4428 585
R3897 gnd.n3905 gnd.n3904 585
R3898 gnd.n3904 gnd.n3902 585
R3899 gnd.n4423 gnd.n4422 585
R3900 gnd.n4422 gnd.n4421 585
R3901 gnd.n3908 gnd.n3907 585
R3902 gnd.n3917 gnd.n3908 585
R3903 gnd.n4412 gnd.n4411 585
R3904 gnd.n4413 gnd.n4412 585
R3905 gnd.n3919 gnd.n3918 585
R3906 gnd.n3918 gnd.n3915 585
R3907 gnd.n4407 gnd.n4406 585
R3908 gnd.n4406 gnd.n4405 585
R3909 gnd.n3922 gnd.n3921 585
R3910 gnd.n3923 gnd.n3922 585
R3911 gnd.n4396 gnd.n4395 585
R3912 gnd.n4397 gnd.n4396 585
R3913 gnd.n3983 gnd.n3982 585
R3914 gnd.n3982 gnd.n3929 585
R3915 gnd.n4391 gnd.n4390 585
R3916 gnd.n4390 gnd.n2663 585
R3917 gnd.n4389 gnd.n3985 585
R3918 gnd.n4389 gnd.n2649 585
R3919 gnd.n4388 gnd.n4386 585
R3920 gnd.n4388 gnd.n4387 585
R3921 gnd.n3987 gnd.n3986 585
R3922 gnd.n3986 gnd.n2752 585
R3923 gnd.n4382 gnd.n4381 585
R3924 gnd.n4381 gnd.n2738 585
R3925 gnd.n4380 gnd.n3989 585
R3926 gnd.n4380 gnd.n2635 585
R3927 gnd.n4379 gnd.n4378 585
R3928 gnd.n4379 gnd.n2632 585
R3929 gnd.n3991 gnd.n3990 585
R3930 gnd.n3990 gnd.n2640 585
R3931 gnd.n4374 gnd.n4373 585
R3932 gnd.n4373 gnd.n2623 585
R3933 gnd.n4372 gnd.n3993 585
R3934 gnd.n4372 gnd.n2616 585
R3935 gnd.n4371 gnd.n4370 585
R3936 gnd.n4371 gnd.n2613 585
R3937 gnd.n3995 gnd.n3994 585
R3938 gnd.n3994 gnd.n2605 585
R3939 gnd.n4366 gnd.n4365 585
R3940 gnd.n4365 gnd.n4364 585
R3941 gnd.n3998 gnd.n3997 585
R3942 gnd.n3998 gnd.n2596 585
R3943 gnd.n4306 gnd.n4305 585
R3944 gnd.n4305 gnd.n2593 585
R3945 gnd.n4307 gnd.n4300 585
R3946 gnd.n4300 gnd.n2585 585
R3947 gnd.n4309 gnd.n4308 585
R3948 gnd.n4309 gnd.n2582 585
R3949 gnd.n4310 gnd.n4299 585
R3950 gnd.n4310 gnd.n4010 585
R3951 gnd.n4312 gnd.n4311 585
R3952 gnd.n4311 gnd.n2573 585
R3953 gnd.n4313 gnd.n4018 585
R3954 gnd.n4018 gnd.n2566 585
R3955 gnd.n4315 gnd.n4314 585
R3956 gnd.n4316 gnd.n4315 585
R3957 gnd.n4294 gnd.n4017 585
R3958 gnd.n4017 gnd.n2555 585
R3959 gnd.n4293 gnd.n4292 585
R3960 gnd.n4292 gnd.n2552 585
R3961 gnd.n4291 gnd.n4021 585
R3962 gnd.n4291 gnd.n4290 585
R3963 gnd.n4227 gnd.n4020 585
R3964 gnd.n4031 gnd.n4020 585
R3965 gnd.n4229 gnd.n4225 585
R3966 gnd.n4225 gnd.n4029 585
R3967 gnd.n4231 gnd.n4230 585
R3968 gnd.n4231 gnd.n4036 585
R3969 gnd.n4232 gnd.n4224 585
R3970 gnd.n4232 gnd.n4046 585
R3971 gnd.n4234 gnd.n4233 585
R3972 gnd.n4233 gnd.n4054 585
R3973 gnd.n4236 gnd.n4061 585
R3974 gnd.n4061 gnd.n4052 585
R3975 gnd.n4238 gnd.n4237 585
R3976 gnd.n4239 gnd.n4238 585
R3977 gnd.n4222 gnd.n4060 585
R3978 gnd.n4060 gnd.n2537 585
R3979 gnd.n4221 gnd.n4220 585
R3980 gnd.n4220 gnd.n2530 585
R3981 gnd.n4219 gnd.n4062 585
R3982 gnd.n4219 gnd.n2527 585
R3983 gnd.n4218 gnd.n4217 585
R3984 gnd.n4218 gnd.n2519 585
R3985 gnd.n4065 gnd.n4064 585
R3986 gnd.n4064 gnd.n2516 585
R3987 gnd.n4212 gnd.n4211 585
R3988 gnd.n4211 gnd.n2509 585
R3989 gnd.n4210 gnd.n4067 585
R3990 gnd.n4210 gnd.n2506 585
R3991 gnd.n4209 gnd.n4073 585
R3992 gnd.n4209 gnd.n4208 585
R3993 gnd.n4069 gnd.n4068 585
R3994 gnd.n4068 gnd.n2496 585
R3995 gnd.n5716 gnd.n5715 585
R3996 gnd.n5717 gnd.n5716 585
R3997 gnd.n3093 gnd.n3091 585
R3998 gnd.n3091 gnd.n3088 585
R3999 gnd.n5273 gnd.n5272 585
R4000 gnd.n5275 gnd.n5273 585
R4001 gnd.n3454 gnd.n3453 585
R4002 gnd.n3453 gnd.n3452 585
R4003 gnd.n5268 gnd.n5267 585
R4004 gnd.n5267 gnd.n5266 585
R4005 gnd.n3457 gnd.n3456 585
R4006 gnd.n3458 gnd.n3457 585
R4007 gnd.n5253 gnd.n5252 585
R4008 gnd.n5255 gnd.n5253 585
R4009 gnd.n3465 gnd.n3464 585
R4010 gnd.n3470 gnd.n3464 585
R4011 gnd.n5248 gnd.n5247 585
R4012 gnd.n5247 gnd.n5246 585
R4013 gnd.n3468 gnd.n3467 585
R4014 gnd.n3469 gnd.n3468 585
R4015 gnd.n5236 gnd.n5235 585
R4016 gnd.n5238 gnd.n5236 585
R4017 gnd.n3478 gnd.n3477 585
R4018 gnd.n3477 gnd.n3476 585
R4019 gnd.n5231 gnd.n5230 585
R4020 gnd.n5230 gnd.n5229 585
R4021 gnd.n3481 gnd.n3480 585
R4022 gnd.n3482 gnd.n3481 585
R4023 gnd.n5219 gnd.n5218 585
R4024 gnd.n5221 gnd.n5219 585
R4025 gnd.n3490 gnd.n3489 585
R4026 gnd.n3489 gnd.n3488 585
R4027 gnd.n5214 gnd.n5213 585
R4028 gnd.n5213 gnd.n5212 585
R4029 gnd.n3493 gnd.n3492 585
R4030 gnd.n3494 gnd.n3493 585
R4031 gnd.n5202 gnd.n5201 585
R4032 gnd.n5204 gnd.n5202 585
R4033 gnd.n3502 gnd.n3501 585
R4034 gnd.n3501 gnd.n3500 585
R4035 gnd.n5197 gnd.n5196 585
R4036 gnd.n5196 gnd.n5195 585
R4037 gnd.n3505 gnd.n3504 585
R4038 gnd.n5185 gnd.n3505 585
R4039 gnd.n5184 gnd.n5183 585
R4040 gnd.n5187 gnd.n5184 585
R4041 gnd.n3512 gnd.n3511 585
R4042 gnd.n3532 gnd.n3511 585
R4043 gnd.n5179 gnd.n5178 585
R4044 gnd.n5178 gnd.n5177 585
R4045 gnd.n3515 gnd.n3514 585
R4046 gnd.n3526 gnd.n3515 585
R4047 gnd.n4918 gnd.n3524 585
R4048 gnd.n5169 gnd.n3524 585
R4049 gnd.n4917 gnd.n4916 585
R4050 gnd.n4916 gnd.t144 585
R4051 gnd.n4922 gnd.n4915 585
R4052 gnd.n4915 gnd.n3541 585
R4053 gnd.n4923 gnd.n3546 585
R4054 gnd.n4948 gnd.n3546 585
R4055 gnd.n4924 gnd.n4914 585
R4056 gnd.n4914 gnd.n4913 585
R4057 gnd.n3564 gnd.n3555 585
R4058 gnd.n4938 gnd.n3555 585
R4059 gnd.n4929 gnd.n4928 585
R4060 gnd.n4930 gnd.n4929 585
R4061 gnd.n3563 gnd.n3562 585
R4062 gnd.n3569 gnd.n3562 585
R4063 gnd.n4799 gnd.n3575 585
R4064 gnd.n4892 gnd.n3575 585
R4065 gnd.n4800 gnd.n4798 585
R4066 gnd.n4798 gnd.n3573 585
R4067 gnd.n4796 gnd.n3584 585
R4068 gnd.n4882 gnd.n3584 585
R4069 gnd.n4804 gnd.n4795 585
R4070 gnd.n4795 gnd.n4794 585
R4071 gnd.n4805 gnd.n3593 585
R4072 gnd.n4865 gnd.n3593 585
R4073 gnd.n4806 gnd.n4793 585
R4074 gnd.n4793 gnd.n3603 585
R4075 gnd.n4791 gnd.n3601 585
R4076 gnd.n4857 gnd.n3601 585
R4077 gnd.n4810 gnd.n4790 585
R4078 gnd.n4790 gnd.n3607 585
R4079 gnd.n4811 gnd.n3612 585
R4080 gnd.n4837 gnd.n3612 585
R4081 gnd.n4812 gnd.n4789 585
R4082 gnd.n4789 gnd.n4788 585
R4083 gnd.n3629 gnd.n3620 585
R4084 gnd.n4829 gnd.n3620 585
R4085 gnd.n4817 gnd.n4816 585
R4086 gnd.n4818 gnd.n4817 585
R4087 gnd.n3628 gnd.n3627 585
R4088 gnd.n4777 gnd.n3627 585
R4089 gnd.n4681 gnd.n4680 585
R4090 gnd.n4680 gnd.n4679 585
R4091 gnd.n4678 gnd.n3641 585
R4092 gnd.n4769 gnd.n3641 585
R4093 gnd.n4685 gnd.n3650 585
R4094 gnd.n4758 gnd.n3650 585
R4095 gnd.n4686 gnd.n4677 585
R4096 gnd.n4677 gnd.n3655 585
R4097 gnd.n4687 gnd.n4676 585
R4098 gnd.n4676 gnd.n3653 585
R4099 gnd.n4675 gnd.n4673 585
R4100 gnd.n4675 gnd.n3659 585
R4101 gnd.n4691 gnd.n4672 585
R4102 gnd.n4672 gnd.n3665 585
R4103 gnd.n4692 gnd.n3671 585
R4104 gnd.n4726 gnd.n3671 585
R4105 gnd.n4693 gnd.n4671 585
R4106 gnd.n4671 gnd.n3669 585
R4107 gnd.n3688 gnd.n3680 585
R4108 gnd.n4707 gnd.n3680 585
R4109 gnd.n4698 gnd.n4697 585
R4110 gnd.n4699 gnd.n4698 585
R4111 gnd.n3687 gnd.n3686 585
R4112 gnd.n4641 gnd.n3686 585
R4113 gnd.n4667 gnd.n4666 585
R4114 gnd.n4666 gnd.n4665 585
R4115 gnd.n3691 gnd.n3690 585
R4116 gnd.n3708 gnd.n3691 585
R4117 gnd.n4591 gnd.n3700 585
R4118 gnd.n4655 gnd.n3700 585
R4119 gnd.n4594 gnd.n4590 585
R4120 gnd.n4590 gnd.n4589 585
R4121 gnd.n4595 gnd.n3718 585
R4122 gnd.n4619 gnd.n3718 585
R4123 gnd.n4596 gnd.n4587 585
R4124 gnd.n4587 gnd.n3716 585
R4125 gnd.n3735 gnd.n3726 585
R4126 gnd.n4611 gnd.n3726 585
R4127 gnd.n4601 gnd.n4600 585
R4128 gnd.n4603 gnd.n4601 585
R4129 gnd.n3734 gnd.n3733 585
R4130 gnd.n4535 gnd.n3733 585
R4131 gnd.n4583 gnd.n4582 585
R4132 gnd.n4582 gnd.n4581 585
R4133 gnd.n3738 gnd.n3737 585
R4134 gnd.n4550 gnd.n3738 585
R4135 gnd.n4508 gnd.n3748 585
R4136 gnd.n4571 gnd.n3748 585
R4137 gnd.n4509 gnd.n4507 585
R4138 gnd.n4507 gnd.n3754 585
R4139 gnd.n3851 gnd.n3849 585
R4140 gnd.n3849 gnd.n3760 585
R4141 gnd.n4514 gnd.n4513 585
R4142 gnd.n4523 gnd.n4514 585
R4143 gnd.n3850 gnd.n3848 585
R4144 gnd.n3848 gnd.n3768 585
R4145 gnd.n4503 gnd.n2988 585
R4146 gnd.n5834 gnd.n2988 585
R4147 gnd.n4502 gnd.n4501 585
R4148 gnd.n4501 gnd.n4500 585
R4149 gnd.n4499 gnd.n2976 585
R4150 gnd.n5840 gnd.n2976 585
R4151 gnd.n4493 gnd.n3853 585
R4152 gnd.n4493 gnd.n2948 585
R4153 gnd.n4495 gnd.n4494 585
R4154 gnd.n4494 gnd.n2916 585
R4155 gnd.n4492 gnd.n3855 585
R4156 gnd.n4492 gnd.n4491 585
R4157 gnd.n3951 gnd.n3856 585
R4158 gnd.n3866 gnd.n3856 585
R4159 gnd.n3952 gnd.n3865 585
R4160 gnd.n4480 gnd.n3865 585
R4161 gnd.n3949 gnd.n3948 585
R4162 gnd.n3948 gnd.n3864 585
R4163 gnd.n3956 gnd.n3875 585
R4164 gnd.n4461 gnd.n3875 585
R4165 gnd.n3957 gnd.n3947 585
R4166 gnd.n3947 gnd.n3874 585
R4167 gnd.n3958 gnd.n3882 585
R4168 gnd.n4453 gnd.n3882 585
R4169 gnd.n3945 gnd.n3944 585
R4170 gnd.n3944 gnd.n3881 585
R4171 gnd.n3962 gnd.n3889 585
R4172 gnd.n4445 gnd.n3889 585
R4173 gnd.n3963 gnd.n3943 585
R4174 gnd.n3943 gnd.n3888 585
R4175 gnd.n3964 gnd.n3896 585
R4176 gnd.n4437 gnd.n3896 585
R4177 gnd.n3941 gnd.n3940 585
R4178 gnd.n3940 gnd.n3895 585
R4179 gnd.n3968 gnd.n3903 585
R4180 gnd.n4429 gnd.n3903 585
R4181 gnd.n3969 gnd.n3939 585
R4182 gnd.n3939 gnd.n3902 585
R4183 gnd.n3970 gnd.n3909 585
R4184 gnd.n4421 gnd.n3909 585
R4185 gnd.n3937 gnd.n3936 585
R4186 gnd.n3936 gnd.n3917 585
R4187 gnd.n3974 gnd.n3916 585
R4188 gnd.n4413 gnd.n3916 585
R4189 gnd.n3975 gnd.n3935 585
R4190 gnd.n3935 gnd.n3915 585
R4191 gnd.n3976 gnd.n3924 585
R4192 gnd.n4405 gnd.n3924 585
R4193 gnd.n3932 gnd.n3930 585
R4194 gnd.n3930 gnd.n3923 585
R4195 gnd.n3981 gnd.n3980 585
R4196 gnd.n4397 gnd.n3981 585
R4197 gnd.n3931 gnd.n2666 585
R4198 gnd.n3929 gnd.n2666 585
R4199 gnd.n6028 gnd.n6027 585
R4200 gnd.n6026 gnd.n2665 585
R4201 gnd.n2668 gnd.n2664 585
R4202 gnd.n6030 gnd.n2664 585
R4203 gnd.n6022 gnd.n2670 585
R4204 gnd.n6021 gnd.n2671 585
R4205 gnd.n6020 gnd.n2672 585
R4206 gnd.n2675 gnd.n2673 585
R4207 gnd.n6015 gnd.n2676 585
R4208 gnd.n6014 gnd.n2677 585
R4209 gnd.n6013 gnd.n2678 585
R4210 gnd.n2687 gnd.n2679 585
R4211 gnd.n6006 gnd.n2688 585
R4212 gnd.n6005 gnd.n2689 585
R4213 gnd.n2691 gnd.n2690 585
R4214 gnd.n5998 gnd.n2697 585
R4215 gnd.n5997 gnd.n2698 585
R4216 gnd.n2705 gnd.n2699 585
R4217 gnd.n5990 gnd.n2706 585
R4218 gnd.n5989 gnd.n2707 585
R4219 gnd.n2709 gnd.n2708 585
R4220 gnd.n5982 gnd.n2715 585
R4221 gnd.n5981 gnd.n2716 585
R4222 gnd.n2723 gnd.n2717 585
R4223 gnd.n5974 gnd.n2724 585
R4224 gnd.n5973 gnd.n2725 585
R4225 gnd.n2730 gnd.n2729 585
R4226 gnd.n2661 gnd.n2646 585
R4227 gnd.n6034 gnd.n2647 585
R4228 gnd.n6033 gnd.n6032 585
R4229 gnd.n5719 gnd.n5718 585
R4230 gnd.n5718 gnd.n5717 585
R4231 gnd.n5720 gnd.n3086 585
R4232 gnd.n3088 gnd.n3086 585
R4233 gnd.n5274 gnd.n3084 585
R4234 gnd.n5275 gnd.n5274 585
R4235 gnd.n5724 gnd.n3083 585
R4236 gnd.n3452 gnd.n3083 585
R4237 gnd.n5725 gnd.n3082 585
R4238 gnd.n5266 gnd.n3082 585
R4239 gnd.n5726 gnd.n3081 585
R4240 gnd.n3458 gnd.n3081 585
R4241 gnd.n5254 gnd.n3079 585
R4242 gnd.n5255 gnd.n5254 585
R4243 gnd.n5730 gnd.n3078 585
R4244 gnd.n3470 gnd.n3078 585
R4245 gnd.n5731 gnd.n3077 585
R4246 gnd.n5246 gnd.n3077 585
R4247 gnd.n5732 gnd.n3076 585
R4248 gnd.n3469 gnd.n3076 585
R4249 gnd.n5237 gnd.n3074 585
R4250 gnd.n5238 gnd.n5237 585
R4251 gnd.n5736 gnd.n3073 585
R4252 gnd.n3476 gnd.n3073 585
R4253 gnd.n5737 gnd.n3072 585
R4254 gnd.n5229 gnd.n3072 585
R4255 gnd.n5738 gnd.n3071 585
R4256 gnd.n3482 gnd.n3071 585
R4257 gnd.n5220 gnd.n3069 585
R4258 gnd.n5221 gnd.n5220 585
R4259 gnd.n5742 gnd.n3068 585
R4260 gnd.n3488 gnd.n3068 585
R4261 gnd.n5743 gnd.n3067 585
R4262 gnd.n5212 gnd.n3067 585
R4263 gnd.n5744 gnd.n3066 585
R4264 gnd.n3494 gnd.n3066 585
R4265 gnd.n5203 gnd.n3064 585
R4266 gnd.n5204 gnd.n5203 585
R4267 gnd.n5748 gnd.n3063 585
R4268 gnd.n3500 gnd.n3063 585
R4269 gnd.n5749 gnd.n3062 585
R4270 gnd.n5195 gnd.n3062 585
R4271 gnd.n5750 gnd.n3061 585
R4272 gnd.n5185 gnd.n3061 585
R4273 gnd.n5186 gnd.n3059 585
R4274 gnd.n5187 gnd.n5186 585
R4275 gnd.n5754 gnd.n3058 585
R4276 gnd.n3532 gnd.n3058 585
R4277 gnd.n5755 gnd.n3057 585
R4278 gnd.n5177 gnd.n3057 585
R4279 gnd.n5756 gnd.n3056 585
R4280 gnd.n3526 gnd.n3056 585
R4281 gnd.n5168 gnd.n3054 585
R4282 gnd.n5169 gnd.n5168 585
R4283 gnd.n5760 gnd.n3053 585
R4284 gnd.t144 gnd.n3053 585
R4285 gnd.n5761 gnd.n3052 585
R4286 gnd.n3541 gnd.n3052 585
R4287 gnd.n5762 gnd.n3051 585
R4288 gnd.n4948 gnd.n3051 585
R4289 gnd.n4912 gnd.n3049 585
R4290 gnd.n4913 gnd.n4912 585
R4291 gnd.n5766 gnd.n3048 585
R4292 gnd.n4938 gnd.n3048 585
R4293 gnd.n5767 gnd.n3047 585
R4294 gnd.n4930 gnd.n3047 585
R4295 gnd.n5768 gnd.n3046 585
R4296 gnd.n3569 gnd.n3046 585
R4297 gnd.n3576 gnd.n3044 585
R4298 gnd.n4892 gnd.n3576 585
R4299 gnd.n5772 gnd.n3043 585
R4300 gnd.n3573 gnd.n3043 585
R4301 gnd.n5773 gnd.n3042 585
R4302 gnd.n4882 gnd.n3042 585
R4303 gnd.n5774 gnd.n3041 585
R4304 gnd.n4794 gnd.n3041 585
R4305 gnd.n3595 gnd.n3039 585
R4306 gnd.n4865 gnd.n3595 585
R4307 gnd.n5778 gnd.n3038 585
R4308 gnd.n3603 gnd.n3038 585
R4309 gnd.n5779 gnd.n3037 585
R4310 gnd.n4857 gnd.n3037 585
R4311 gnd.n5780 gnd.n3036 585
R4312 gnd.n3607 gnd.n3036 585
R4313 gnd.n3613 gnd.n3034 585
R4314 gnd.n4837 gnd.n3613 585
R4315 gnd.n5784 gnd.n3033 585
R4316 gnd.n4788 gnd.n3033 585
R4317 gnd.n5785 gnd.n3032 585
R4318 gnd.n4829 gnd.n3032 585
R4319 gnd.n5786 gnd.n3031 585
R4320 gnd.n4818 gnd.n3031 585
R4321 gnd.n3635 gnd.n3029 585
R4322 gnd.n4777 gnd.n3635 585
R4323 gnd.n5790 gnd.n3028 585
R4324 gnd.n4679 gnd.n3028 585
R4325 gnd.n5791 gnd.n3027 585
R4326 gnd.n4769 gnd.n3027 585
R4327 gnd.n5792 gnd.n3026 585
R4328 gnd.n4758 gnd.n3026 585
R4329 gnd.n3654 gnd.n3024 585
R4330 gnd.n3655 gnd.n3654 585
R4331 gnd.n5796 gnd.n3023 585
R4332 gnd.n3653 gnd.n3023 585
R4333 gnd.n5797 gnd.n3022 585
R4334 gnd.n3659 gnd.n3022 585
R4335 gnd.n5798 gnd.n3021 585
R4336 gnd.n3665 gnd.n3021 585
R4337 gnd.n3672 gnd.n3019 585
R4338 gnd.n4726 gnd.n3672 585
R4339 gnd.n5802 gnd.n3018 585
R4340 gnd.n3669 gnd.n3018 585
R4341 gnd.n5803 gnd.n3017 585
R4342 gnd.n4707 gnd.n3017 585
R4343 gnd.n5804 gnd.n3016 585
R4344 gnd.n4699 gnd.n3016 585
R4345 gnd.n4640 gnd.n3014 585
R4346 gnd.n4641 gnd.n4640 585
R4347 gnd.n5808 gnd.n3013 585
R4348 gnd.n4665 gnd.n3013 585
R4349 gnd.n5809 gnd.n3012 585
R4350 gnd.n3708 gnd.n3012 585
R4351 gnd.n5810 gnd.n3011 585
R4352 gnd.n4655 gnd.n3011 585
R4353 gnd.n4588 gnd.n3009 585
R4354 gnd.n4589 gnd.n4588 585
R4355 gnd.n5814 gnd.n3008 585
R4356 gnd.n4619 gnd.n3008 585
R4357 gnd.n5815 gnd.n3007 585
R4358 gnd.n3716 gnd.n3007 585
R4359 gnd.n5816 gnd.n3006 585
R4360 gnd.n4611 gnd.n3006 585
R4361 gnd.n4602 gnd.n3004 585
R4362 gnd.n4603 gnd.n4602 585
R4363 gnd.n5820 gnd.n3003 585
R4364 gnd.n4535 gnd.n3003 585
R4365 gnd.n5821 gnd.n3002 585
R4366 gnd.n4581 gnd.n3002 585
R4367 gnd.n5822 gnd.n3001 585
R4368 gnd.n4550 gnd.n3001 585
R4369 gnd.n4570 gnd.n2999 585
R4370 gnd.n4571 gnd.n4570 585
R4371 gnd.n5826 gnd.n2998 585
R4372 gnd.n3754 gnd.n2998 585
R4373 gnd.n5827 gnd.n2997 585
R4374 gnd.n3760 gnd.n2997 585
R4375 gnd.n5828 gnd.n2996 585
R4376 gnd.n4523 gnd.n2996 585
R4377 gnd.n2993 gnd.n2991 585
R4378 gnd.n3768 gnd.n2991 585
R4379 gnd.n5833 gnd.n5832 585
R4380 gnd.n5834 gnd.n5833 585
R4381 gnd.n2992 gnd.n2990 585
R4382 gnd.n4500 gnd.n2990 585
R4383 gnd.n4469 gnd.n2978 585
R4384 gnd.n5840 gnd.n2978 585
R4385 gnd.n4472 gnd.n4468 585
R4386 gnd.n4468 gnd.n2948 585
R4387 gnd.n4473 gnd.n4467 585
R4388 gnd.n4467 gnd.n2916 585
R4389 gnd.n4474 gnd.n3857 585
R4390 gnd.n4491 gnd.n3857 585
R4391 gnd.n3870 gnd.n3868 585
R4392 gnd.n3868 gnd.n3866 585
R4393 gnd.n4479 gnd.n4478 585
R4394 gnd.n4480 gnd.n4479 585
R4395 gnd.n3869 gnd.n3867 585
R4396 gnd.n3867 gnd.n3864 585
R4397 gnd.n4463 gnd.n4462 585
R4398 gnd.n4462 gnd.n4461 585
R4399 gnd.n3873 gnd.n3872 585
R4400 gnd.n3874 gnd.n3873 585
R4401 gnd.n4452 gnd.n4451 585
R4402 gnd.n4453 gnd.n4452 585
R4403 gnd.n3884 gnd.n3883 585
R4404 gnd.n3883 gnd.n3881 585
R4405 gnd.n4447 gnd.n4446 585
R4406 gnd.n4446 gnd.n4445 585
R4407 gnd.n3887 gnd.n3886 585
R4408 gnd.n3888 gnd.n3887 585
R4409 gnd.n4436 gnd.n4435 585
R4410 gnd.n4437 gnd.n4436 585
R4411 gnd.n3898 gnd.n3897 585
R4412 gnd.n3897 gnd.n3895 585
R4413 gnd.n4431 gnd.n4430 585
R4414 gnd.n4430 gnd.n4429 585
R4415 gnd.n3901 gnd.n3900 585
R4416 gnd.n3902 gnd.n3901 585
R4417 gnd.n4420 gnd.n4419 585
R4418 gnd.n4421 gnd.n4420 585
R4419 gnd.n3911 gnd.n3910 585
R4420 gnd.n3917 gnd.n3910 585
R4421 gnd.n4415 gnd.n4414 585
R4422 gnd.n4414 gnd.n4413 585
R4423 gnd.n3914 gnd.n3913 585
R4424 gnd.n3915 gnd.n3914 585
R4425 gnd.n4404 gnd.n4403 585
R4426 gnd.n4405 gnd.n4404 585
R4427 gnd.n3926 gnd.n3925 585
R4428 gnd.n3925 gnd.n3923 585
R4429 gnd.n4399 gnd.n4398 585
R4430 gnd.n4398 gnd.n4397 585
R4431 gnd.n3928 gnd.n2648 585
R4432 gnd.n3929 gnd.n2648 585
R4433 gnd.n5658 gnd.n3148 585
R4434 gnd.n5297 gnd.n3148 585
R4435 gnd.n5659 gnd.n3147 585
R4436 gnd.n3440 gnd.n3141 585
R4437 gnd.n5666 gnd.n3140 585
R4438 gnd.n5667 gnd.n3139 585
R4439 gnd.n3437 gnd.n3133 585
R4440 gnd.n5674 gnd.n3132 585
R4441 gnd.n5675 gnd.n3131 585
R4442 gnd.n3435 gnd.n3125 585
R4443 gnd.n5682 gnd.n3124 585
R4444 gnd.n5683 gnd.n3123 585
R4445 gnd.n3432 gnd.n3117 585
R4446 gnd.n5690 gnd.n3116 585
R4447 gnd.n5691 gnd.n3115 585
R4448 gnd.n3430 gnd.n3108 585
R4449 gnd.n5698 gnd.n3107 585
R4450 gnd.n5699 gnd.n3106 585
R4451 gnd.n3427 gnd.n3103 585
R4452 gnd.n5704 gnd.n3102 585
R4453 gnd.n5705 gnd.n3101 585
R4454 gnd.n5706 gnd.n3100 585
R4455 gnd.n3424 gnd.n3098 585
R4456 gnd.n5710 gnd.n3097 585
R4457 gnd.n5711 gnd.n3096 585
R4458 gnd.n5712 gnd.n3092 585
R4459 gnd.n5300 gnd.n3087 585
R4460 gnd.n5301 gnd.n5299 585
R4461 gnd.n3422 gnd.n3421 585
R4462 gnd.n3443 gnd.n3442 585
R4463 gnd.n3772 gnd.t148 543.808
R4464 gnd.n5017 gnd.t151 543.808
R4465 gnd.n5846 gnd.t72 543.808
R4466 gnd.n5011 gnd.t61 543.808
R4467 gnd.n5160 gnd.n3534 458.866
R4468 gnd.n5162 gnd.n3531 458.866
R4469 gnd.n3837 gnd.n3836 458.866
R4470 gnd.n5909 gnd.n2951 458.866
R4471 gnd.n6544 gnd.n6543 439.709
R4472 gnd.n2726 gnd.t79 371.625
R4473 gnd.n5652 gnd.t49 371.625
R4474 gnd.n2733 gnd.t65 371.625
R4475 gnd.n3221 gnd.t123 371.625
R4476 gnd.n3244 gnd.t129 371.625
R4477 gnd.n5532 gnd.t93 371.625
R4478 gnd.n175 gnd.t90 371.625
R4479 gnd.n197 gnd.t99 371.625
R4480 gnd.n219 gnd.t105 371.625
R4481 gnd.n7261 gnd.t35 371.625
R4482 gnd.n2402 gnd.t83 371.625
R4483 gnd.n2424 gnd.t108 371.625
R4484 gnd.n2446 gnd.t114 371.625
R4485 gnd.n4096 gnd.t57 371.625
R4486 gnd.n2803 gnd.t102 371.625
R4487 gnd.n2844 gnd.t117 371.625
R4488 gnd.n2823 gnd.t140 371.625
R4489 gnd.n3149 gnd.t53 371.625
R4490 gnd.n1703 gnd.t86 323.425
R4491 gnd.n1051 gnd.t132 323.425
R4492 gnd.n2310 gnd.n2284 289.615
R4493 gnd.n2278 gnd.n2252 289.615
R4494 gnd.n2246 gnd.n2220 289.615
R4495 gnd.n2215 gnd.n2189 289.615
R4496 gnd.n2183 gnd.n2157 289.615
R4497 gnd.n2151 gnd.n2125 289.615
R4498 gnd.n2119 gnd.n2093 289.615
R4499 gnd.n2088 gnd.n2062 289.615
R4500 gnd.n1440 gnd.t136 279.217
R4501 gnd.n1072 gnd.t42 279.217
R4502 gnd.n2958 gnd.t48 260.649
R4503 gnd.n4981 gnd.t71 260.649
R4504 gnd.n5911 gnd.n5910 256.663
R4505 gnd.n5911 gnd.n2917 256.663
R4506 gnd.n5911 gnd.n2918 256.663
R4507 gnd.n5911 gnd.n2919 256.663
R4508 gnd.n5911 gnd.n2920 256.663
R4509 gnd.n5911 gnd.n2921 256.663
R4510 gnd.n5911 gnd.n2922 256.663
R4511 gnd.n5911 gnd.n2923 256.663
R4512 gnd.n5911 gnd.n2924 256.663
R4513 gnd.n5911 gnd.n2925 256.663
R4514 gnd.n5911 gnd.n2926 256.663
R4515 gnd.n5911 gnd.n2927 256.663
R4516 gnd.n5911 gnd.n2928 256.663
R4517 gnd.n5911 gnd.n2929 256.663
R4518 gnd.n5911 gnd.n2930 256.663
R4519 gnd.n5911 gnd.n2931 256.663
R4520 gnd.n5914 gnd.n2914 256.663
R4521 gnd.n5912 gnd.n5911 256.663
R4522 gnd.n5911 gnd.n2932 256.663
R4523 gnd.n5911 gnd.n2933 256.663
R4524 gnd.n5911 gnd.n2934 256.663
R4525 gnd.n5911 gnd.n2935 256.663
R4526 gnd.n5911 gnd.n2936 256.663
R4527 gnd.n5911 gnd.n2937 256.663
R4528 gnd.n5911 gnd.n2938 256.663
R4529 gnd.n5911 gnd.n2939 256.663
R4530 gnd.n5911 gnd.n2940 256.663
R4531 gnd.n5911 gnd.n2941 256.663
R4532 gnd.n5911 gnd.n2942 256.663
R4533 gnd.n5911 gnd.n2943 256.663
R4534 gnd.n5911 gnd.n2944 256.663
R4535 gnd.n5911 gnd.n2945 256.663
R4536 gnd.n5911 gnd.n2946 256.663
R4537 gnd.n5911 gnd.n2947 256.663
R4538 gnd.n5039 gnd.n4991 256.663
R4539 gnd.n5045 gnd.n4991 256.663
R4540 gnd.n5038 gnd.n4991 256.663
R4541 gnd.n5052 gnd.n4991 256.663
R4542 gnd.n5035 gnd.n4991 256.663
R4543 gnd.n5059 gnd.n4991 256.663
R4544 gnd.n5032 gnd.n4991 256.663
R4545 gnd.n5066 gnd.n4991 256.663
R4546 gnd.n5029 gnd.n4991 256.663
R4547 gnd.n5073 gnd.n4991 256.663
R4548 gnd.n5026 gnd.n4991 256.663
R4549 gnd.n5080 gnd.n4991 256.663
R4550 gnd.n5023 gnd.n4991 256.663
R4551 gnd.n5087 gnd.n4991 256.663
R4552 gnd.n5020 gnd.n4991 256.663
R4553 gnd.n5095 gnd.n4991 256.663
R4554 gnd.n5098 gnd.n3231 256.663
R4555 gnd.n5099 gnd.n4991 256.663
R4556 gnd.n5103 gnd.n4991 256.663
R4557 gnd.n5014 gnd.n4991 256.663
R4558 gnd.n5111 gnd.n4991 256.663
R4559 gnd.n5009 gnd.n4991 256.663
R4560 gnd.n5118 gnd.n4991 256.663
R4561 gnd.n5006 gnd.n4991 256.663
R4562 gnd.n5125 gnd.n4991 256.663
R4563 gnd.n5003 gnd.n4991 256.663
R4564 gnd.n5132 gnd.n4991 256.663
R4565 gnd.n5000 gnd.n4991 256.663
R4566 gnd.n5139 gnd.n4991 256.663
R4567 gnd.n4997 gnd.n4991 256.663
R4568 gnd.n5146 gnd.n4991 256.663
R4569 gnd.n4994 gnd.n4991 256.663
R4570 gnd.n5153 gnd.n4991 256.663
R4571 gnd.n4991 gnd.n4990 256.663
R4572 gnd.n6276 gnd.n2370 242.672
R4573 gnd.n6276 gnd.n2371 242.672
R4574 gnd.n6276 gnd.n2372 242.672
R4575 gnd.n6276 gnd.n2373 242.672
R4576 gnd.n6276 gnd.n2374 242.672
R4577 gnd.n6276 gnd.n2375 242.672
R4578 gnd.n6276 gnd.n2376 242.672
R4579 gnd.n6276 gnd.n2377 242.672
R4580 gnd.n6276 gnd.n2378 242.672
R4581 gnd.n5966 gnd.n5965 242.672
R4582 gnd.n5965 gnd.n2751 242.672
R4583 gnd.n5965 gnd.n2749 242.672
R4584 gnd.n5965 gnd.n2748 242.672
R4585 gnd.n5965 gnd.n2746 242.672
R4586 gnd.n5965 gnd.n2744 242.672
R4587 gnd.n5965 gnd.n2743 242.672
R4588 gnd.n5965 gnd.n2741 242.672
R4589 gnd.n5965 gnd.n2739 242.672
R4590 gnd.n1495 gnd.n1404 242.672
R4591 gnd.n1408 gnd.n1404 242.672
R4592 gnd.n1488 gnd.n1404 242.672
R4593 gnd.n1482 gnd.n1404 242.672
R4594 gnd.n1480 gnd.n1404 242.672
R4595 gnd.n1474 gnd.n1404 242.672
R4596 gnd.n1472 gnd.n1404 242.672
R4597 gnd.n1466 gnd.n1404 242.672
R4598 gnd.n1464 gnd.n1404 242.672
R4599 gnd.n1458 gnd.n1404 242.672
R4600 gnd.n1456 gnd.n1404 242.672
R4601 gnd.n1449 gnd.n1404 242.672
R4602 gnd.n1447 gnd.n1404 242.672
R4603 gnd.n6323 gnd.n2341 242.672
R4604 gnd.n6323 gnd.n1068 242.672
R4605 gnd.n6323 gnd.n1067 242.672
R4606 gnd.n6323 gnd.n1066 242.672
R4607 gnd.n6323 gnd.n1065 242.672
R4608 gnd.n6323 gnd.n1064 242.672
R4609 gnd.n6323 gnd.n1063 242.672
R4610 gnd.n6323 gnd.n1062 242.672
R4611 gnd.n6323 gnd.n1061 242.672
R4612 gnd.n6323 gnd.n1060 242.672
R4613 gnd.n6323 gnd.n1059 242.672
R4614 gnd.n6323 gnd.n1058 242.672
R4615 gnd.n6323 gnd.n1057 242.672
R4616 gnd.n5649 gnd.n3186 242.672
R4617 gnd.n5649 gnd.n3188 242.672
R4618 gnd.n5649 gnd.n3189 242.672
R4619 gnd.n5649 gnd.n3191 242.672
R4620 gnd.n5649 gnd.n3193 242.672
R4621 gnd.n5649 gnd.n3194 242.672
R4622 gnd.n5649 gnd.n3196 242.672
R4623 gnd.n5649 gnd.n3198 242.672
R4624 gnd.n5650 gnd.n5649 242.672
R4625 gnd.n7323 gnd.n171 242.672
R4626 gnd.n7264 gnd.n171 242.672
R4627 gnd.n7313 gnd.n171 242.672
R4628 gnd.n7268 gnd.n171 242.672
R4629 gnd.n7303 gnd.n171 242.672
R4630 gnd.n7272 gnd.n171 242.672
R4631 gnd.n7293 gnd.n171 242.672
R4632 gnd.n7276 gnd.n171 242.672
R4633 gnd.n7283 gnd.n171 242.672
R4634 gnd.n1737 gnd.n1736 242.672
R4635 gnd.n1737 gnd.n1678 242.672
R4636 gnd.n1737 gnd.n1679 242.672
R4637 gnd.n1737 gnd.n1680 242.672
R4638 gnd.n1737 gnd.n1681 242.672
R4639 gnd.n1737 gnd.n1682 242.672
R4640 gnd.n1737 gnd.n1683 242.672
R4641 gnd.n1737 gnd.n1684 242.672
R4642 gnd.n6323 gnd.n1050 242.672
R4643 gnd.n6324 gnd.n6323 242.672
R4644 gnd.n6323 gnd.n6277 242.672
R4645 gnd.n6323 gnd.n6278 242.672
R4646 gnd.n6323 gnd.n6279 242.672
R4647 gnd.n6323 gnd.n6280 242.672
R4648 gnd.n6323 gnd.n6281 242.672
R4649 gnd.n6323 gnd.n6282 242.672
R4650 gnd.n6276 gnd.n6275 242.672
R4651 gnd.n6276 gnd.n2342 242.672
R4652 gnd.n6276 gnd.n2343 242.672
R4653 gnd.n6276 gnd.n2344 242.672
R4654 gnd.n6276 gnd.n2345 242.672
R4655 gnd.n6276 gnd.n2346 242.672
R4656 gnd.n6276 gnd.n2347 242.672
R4657 gnd.n6276 gnd.n2348 242.672
R4658 gnd.n6276 gnd.n2349 242.672
R4659 gnd.n6276 gnd.n2350 242.672
R4660 gnd.n6276 gnd.n2351 242.672
R4661 gnd.n6276 gnd.n2352 242.672
R4662 gnd.n6276 gnd.n2353 242.672
R4663 gnd.n6276 gnd.n2354 242.672
R4664 gnd.n6276 gnd.n2355 242.672
R4665 gnd.n6276 gnd.n2356 242.672
R4666 gnd.n6276 gnd.n2357 242.672
R4667 gnd.n6276 gnd.n2358 242.672
R4668 gnd.n6276 gnd.n2359 242.672
R4669 gnd.n6276 gnd.n2360 242.672
R4670 gnd.n6276 gnd.n2361 242.672
R4671 gnd.n6276 gnd.n2362 242.672
R4672 gnd.n6276 gnd.n2363 242.672
R4673 gnd.n6276 gnd.n2364 242.672
R4674 gnd.n6276 gnd.n2365 242.672
R4675 gnd.n6276 gnd.n2366 242.672
R4676 gnd.n6276 gnd.n2367 242.672
R4677 gnd.n6276 gnd.n2368 242.672
R4678 gnd.n6276 gnd.n2369 242.672
R4679 gnd.n5965 gnd.n2753 242.672
R4680 gnd.n5965 gnd.n2754 242.672
R4681 gnd.n5965 gnd.n2755 242.672
R4682 gnd.n5965 gnd.n2756 242.672
R4683 gnd.n5965 gnd.n2757 242.672
R4684 gnd.n5965 gnd.n2758 242.672
R4685 gnd.n5965 gnd.n2759 242.672
R4686 gnd.n5965 gnd.n2760 242.672
R4687 gnd.n5965 gnd.n2761 242.672
R4688 gnd.n5965 gnd.n2762 242.672
R4689 gnd.n5965 gnd.n2763 242.672
R4690 gnd.n5965 gnd.n2764 242.672
R4691 gnd.n5965 gnd.n2765 242.672
R4692 gnd.n5965 gnd.n2766 242.672
R4693 gnd.n5965 gnd.n2767 242.672
R4694 gnd.n5965 gnd.n2768 242.672
R4695 gnd.n5915 gnd.n2814 242.672
R4696 gnd.n5965 gnd.n2769 242.672
R4697 gnd.n5965 gnd.n2770 242.672
R4698 gnd.n5965 gnd.n2771 242.672
R4699 gnd.n5965 gnd.n2772 242.672
R4700 gnd.n5965 gnd.n2773 242.672
R4701 gnd.n5965 gnd.n2774 242.672
R4702 gnd.n5965 gnd.n2775 242.672
R4703 gnd.n5965 gnd.n2776 242.672
R4704 gnd.n5965 gnd.n2777 242.672
R4705 gnd.n5965 gnd.n2778 242.672
R4706 gnd.n5965 gnd.n2779 242.672
R4707 gnd.n5965 gnd.n2780 242.672
R4708 gnd.n5965 gnd.n5964 242.672
R4709 gnd.n5649 gnd.n5648 242.672
R4710 gnd.n5649 gnd.n3158 242.672
R4711 gnd.n5649 gnd.n3159 242.672
R4712 gnd.n5649 gnd.n3160 242.672
R4713 gnd.n5649 gnd.n3161 242.672
R4714 gnd.n5649 gnd.n3162 242.672
R4715 gnd.n5649 gnd.n3163 242.672
R4716 gnd.n5649 gnd.n3164 242.672
R4717 gnd.n5649 gnd.n3165 242.672
R4718 gnd.n5649 gnd.n3166 242.672
R4719 gnd.n5649 gnd.n3167 242.672
R4720 gnd.n5649 gnd.n3168 242.672
R4721 gnd.n5649 gnd.n3169 242.672
R4722 gnd.n5596 gnd.n3232 242.672
R4723 gnd.n5649 gnd.n3170 242.672
R4724 gnd.n5649 gnd.n3171 242.672
R4725 gnd.n5649 gnd.n3172 242.672
R4726 gnd.n5649 gnd.n3173 242.672
R4727 gnd.n5649 gnd.n3174 242.672
R4728 gnd.n5649 gnd.n3175 242.672
R4729 gnd.n5649 gnd.n3176 242.672
R4730 gnd.n5649 gnd.n3177 242.672
R4731 gnd.n5649 gnd.n3178 242.672
R4732 gnd.n5649 gnd.n3179 242.672
R4733 gnd.n5649 gnd.n3180 242.672
R4734 gnd.n5649 gnd.n3181 242.672
R4735 gnd.n5649 gnd.n3182 242.672
R4736 gnd.n5649 gnd.n3183 242.672
R4737 gnd.n5649 gnd.n3184 242.672
R4738 gnd.n5649 gnd.n3185 242.672
R4739 gnd.n382 gnd.n171 242.672
R4740 gnd.n178 gnd.n171 242.672
R4741 gnd.n372 gnd.n171 242.672
R4742 gnd.n182 gnd.n171 242.672
R4743 gnd.n362 gnd.n171 242.672
R4744 gnd.n186 gnd.n171 242.672
R4745 gnd.n352 gnd.n171 242.672
R4746 gnd.n190 gnd.n171 242.672
R4747 gnd.n342 gnd.n171 242.672
R4748 gnd.n194 gnd.n171 242.672
R4749 gnd.n332 gnd.n171 242.672
R4750 gnd.n200 gnd.n171 242.672
R4751 gnd.n322 gnd.n171 242.672
R4752 gnd.n204 gnd.n171 242.672
R4753 gnd.n312 gnd.n171 242.672
R4754 gnd.n208 gnd.n171 242.672
R4755 gnd.n302 gnd.n171 242.672
R4756 gnd.n212 gnd.n171 242.672
R4757 gnd.n292 gnd.n171 242.672
R4758 gnd.n216 gnd.n171 242.672
R4759 gnd.n282 gnd.n171 242.672
R4760 gnd.n272 gnd.n171 242.672
R4761 gnd.n271 gnd.n171 242.672
R4762 gnd.n226 gnd.n171 242.672
R4763 gnd.n261 gnd.n171 242.672
R4764 gnd.n230 gnd.n171 242.672
R4765 gnd.n251 gnd.n171 242.672
R4766 gnd.n234 gnd.n171 242.672
R4767 gnd.n241 gnd.n171 242.672
R4768 gnd.n6030 gnd.n6029 242.672
R4769 gnd.n6030 gnd.n2650 242.672
R4770 gnd.n6030 gnd.n2651 242.672
R4771 gnd.n6030 gnd.n2652 242.672
R4772 gnd.n6030 gnd.n2653 242.672
R4773 gnd.n6030 gnd.n2654 242.672
R4774 gnd.n6030 gnd.n2655 242.672
R4775 gnd.n6030 gnd.n2656 242.672
R4776 gnd.n6030 gnd.n2657 242.672
R4777 gnd.n6030 gnd.n2658 242.672
R4778 gnd.n6030 gnd.n2659 242.672
R4779 gnd.n6030 gnd.n2660 242.672
R4780 gnd.n6030 gnd.n2662 242.672
R4781 gnd.n6031 gnd.n6030 242.672
R4782 gnd.n5297 gnd.n3441 242.672
R4783 gnd.n5297 gnd.n3439 242.672
R4784 gnd.n5297 gnd.n3438 242.672
R4785 gnd.n5297 gnd.n3436 242.672
R4786 gnd.n5297 gnd.n3434 242.672
R4787 gnd.n5297 gnd.n3433 242.672
R4788 gnd.n5297 gnd.n3431 242.672
R4789 gnd.n5297 gnd.n3429 242.672
R4790 gnd.n5297 gnd.n3428 242.672
R4791 gnd.n5297 gnd.n3426 242.672
R4792 gnd.n5297 gnd.n3425 242.672
R4793 gnd.n5297 gnd.n3423 242.672
R4794 gnd.n5298 gnd.n5297 242.672
R4795 gnd.n5297 gnd.n3444 242.672
R4796 gnd.n240 gnd.n167 240.244
R4797 gnd.n243 gnd.n242 240.244
R4798 gnd.n250 gnd.n249 240.244
R4799 gnd.n253 gnd.n252 240.244
R4800 gnd.n260 gnd.n259 240.244
R4801 gnd.n263 gnd.n262 240.244
R4802 gnd.n270 gnd.n269 240.244
R4803 gnd.n274 gnd.n273 240.244
R4804 gnd.n281 gnd.n222 240.244
R4805 gnd.n284 gnd.n283 240.244
R4806 gnd.n291 gnd.n290 240.244
R4807 gnd.n294 gnd.n293 240.244
R4808 gnd.n301 gnd.n300 240.244
R4809 gnd.n304 gnd.n303 240.244
R4810 gnd.n311 gnd.n310 240.244
R4811 gnd.n314 gnd.n313 240.244
R4812 gnd.n321 gnd.n320 240.244
R4813 gnd.n324 gnd.n323 240.244
R4814 gnd.n331 gnd.n330 240.244
R4815 gnd.n334 gnd.n333 240.244
R4816 gnd.n341 gnd.n340 240.244
R4817 gnd.n344 gnd.n343 240.244
R4818 gnd.n351 gnd.n350 240.244
R4819 gnd.n354 gnd.n353 240.244
R4820 gnd.n361 gnd.n360 240.244
R4821 gnd.n364 gnd.n363 240.244
R4822 gnd.n371 gnd.n370 240.244
R4823 gnd.n374 gnd.n373 240.244
R4824 gnd.n381 gnd.n380 240.244
R4825 gnd.n5529 gnd.n3265 240.244
R4826 gnd.n5521 gnd.n3265 240.244
R4827 gnd.n5521 gnd.n3276 240.244
R4828 gnd.n3292 gnd.n3276 240.244
R4829 gnd.n5314 gnd.n3292 240.244
R4830 gnd.n5314 gnd.n3305 240.244
R4831 gnd.n5320 gnd.n3305 240.244
R4832 gnd.n5320 gnd.n3315 240.244
R4833 gnd.n5327 gnd.n3315 240.244
R4834 gnd.n5327 gnd.n3325 240.244
R4835 gnd.n3401 gnd.n3325 240.244
R4836 gnd.n3401 gnd.n3335 240.244
R4837 gnd.n5397 gnd.n3335 240.244
R4838 gnd.n5397 gnd.n3345 240.244
R4839 gnd.n5402 gnd.n3345 240.244
R4840 gnd.n5402 gnd.n3352 240.244
R4841 gnd.n5416 gnd.n3352 240.244
R4842 gnd.n5416 gnd.n3362 240.244
R4843 gnd.n3368 gnd.n3362 240.244
R4844 gnd.n5425 gnd.n3368 240.244
R4845 gnd.n5426 gnd.n5425 240.244
R4846 gnd.n5426 gnd.n3379 240.244
R4847 gnd.n3379 gnd.n74 240.244
R4848 gnd.n3385 gnd.n74 240.244
R4849 gnd.n5433 gnd.n3385 240.244
R4850 gnd.n5433 gnd.n91 240.244
R4851 gnd.n7227 gnd.n91 240.244
R4852 gnd.n7227 gnd.n102 240.244
R4853 gnd.n7232 gnd.n102 240.244
R4854 gnd.n7232 gnd.n112 240.244
R4855 gnd.n7242 gnd.n112 240.244
R4856 gnd.n7242 gnd.n121 240.244
R4857 gnd.n7247 gnd.n121 240.244
R4858 gnd.n7247 gnd.n132 240.244
R4859 gnd.n7341 gnd.n132 240.244
R4860 gnd.n7341 gnd.n141 240.244
R4861 gnd.n7345 gnd.n141 240.244
R4862 gnd.n7345 gnd.n151 240.244
R4863 gnd.n7348 gnd.n151 240.244
R4864 gnd.n7348 gnd.n160 240.244
R4865 gnd.n7351 gnd.n160 240.244
R4866 gnd.n7351 gnd.n169 240.244
R4867 gnd.n3201 gnd.n3200 240.244
R4868 gnd.n5642 gnd.n3200 240.244
R4869 gnd.n5640 gnd.n5639 240.244
R4870 gnd.n5636 gnd.n5635 240.244
R4871 gnd.n5632 gnd.n5631 240.244
R4872 gnd.n5628 gnd.n5627 240.244
R4873 gnd.n5624 gnd.n5623 240.244
R4874 gnd.n5620 gnd.n5619 240.244
R4875 gnd.n5616 gnd.n5615 240.244
R4876 gnd.n5611 gnd.n5610 240.244
R4877 gnd.n5607 gnd.n5606 240.244
R4878 gnd.n5603 gnd.n5602 240.244
R4879 gnd.n5599 gnd.n5598 240.244
R4880 gnd.n5594 gnd.n5593 240.244
R4881 gnd.n5590 gnd.n5589 240.244
R4882 gnd.n5586 gnd.n5585 240.244
R4883 gnd.n5582 gnd.n5581 240.244
R4884 gnd.n5578 gnd.n5577 240.244
R4885 gnd.n5574 gnd.n5573 240.244
R4886 gnd.n5570 gnd.n5569 240.244
R4887 gnd.n5566 gnd.n5565 240.244
R4888 gnd.n5562 gnd.n5561 240.244
R4889 gnd.n5558 gnd.n5557 240.244
R4890 gnd.n5554 gnd.n5553 240.244
R4891 gnd.n5550 gnd.n5549 240.244
R4892 gnd.n5546 gnd.n5545 240.244
R4893 gnd.n5542 gnd.n5541 240.244
R4894 gnd.n5538 gnd.n5537 240.244
R4895 gnd.n3280 gnd.n3202 240.244
R4896 gnd.n5519 gnd.n3280 240.244
R4897 gnd.n5519 gnd.n3281 240.244
R4898 gnd.n5515 gnd.n3281 240.244
R4899 gnd.n5515 gnd.n3290 240.244
R4900 gnd.n5507 gnd.n3290 240.244
R4901 gnd.n5507 gnd.n3307 240.244
R4902 gnd.n5503 gnd.n3307 240.244
R4903 gnd.n5503 gnd.n3313 240.244
R4904 gnd.n5495 gnd.n3313 240.244
R4905 gnd.n5495 gnd.n3328 240.244
R4906 gnd.n5491 gnd.n3328 240.244
R4907 gnd.n5491 gnd.n3334 240.244
R4908 gnd.n5483 gnd.n3334 240.244
R4909 gnd.n5483 gnd.n3347 240.244
R4910 gnd.n5479 gnd.n3347 240.244
R4911 gnd.n5479 gnd.n3350 240.244
R4912 gnd.n5471 gnd.n3350 240.244
R4913 gnd.n5471 gnd.n5468 240.244
R4914 gnd.n5468 gnd.n3365 240.244
R4915 gnd.n3377 gnd.n3365 240.244
R4916 gnd.n3377 gnd.n77 240.244
R4917 gnd.n7412 gnd.n77 240.244
R4918 gnd.n7412 gnd.n78 240.244
R4919 gnd.n88 gnd.n78 240.244
R4920 gnd.n7406 gnd.n88 240.244
R4921 gnd.n7406 gnd.n89 240.244
R4922 gnd.n7398 gnd.n89 240.244
R4923 gnd.n7398 gnd.n105 240.244
R4924 gnd.n7394 gnd.n105 240.244
R4925 gnd.n7394 gnd.n110 240.244
R4926 gnd.n7386 gnd.n110 240.244
R4927 gnd.n7386 gnd.n124 240.244
R4928 gnd.n7382 gnd.n124 240.244
R4929 gnd.n7382 gnd.n130 240.244
R4930 gnd.n7374 gnd.n130 240.244
R4931 gnd.n7374 gnd.n144 240.244
R4932 gnd.n7370 gnd.n144 240.244
R4933 gnd.n7370 gnd.n150 240.244
R4934 gnd.n7362 gnd.n150 240.244
R4935 gnd.n7362 gnd.n162 240.244
R4936 gnd.n7358 gnd.n162 240.244
R4937 gnd.n2781 gnd.n2631 240.244
R4938 gnd.n5963 gnd.n2782 240.244
R4939 gnd.n5959 gnd.n5958 240.244
R4940 gnd.n5955 gnd.n5954 240.244
R4941 gnd.n5951 gnd.n5950 240.244
R4942 gnd.n5947 gnd.n5946 240.244
R4943 gnd.n5943 gnd.n5942 240.244
R4944 gnd.n5939 gnd.n5938 240.244
R4945 gnd.n5935 gnd.n5934 240.244
R4946 gnd.n5930 gnd.n5929 240.244
R4947 gnd.n5926 gnd.n5925 240.244
R4948 gnd.n5922 gnd.n5921 240.244
R4949 gnd.n5918 gnd.n5917 240.244
R4950 gnd.n2907 gnd.n2906 240.244
R4951 gnd.n2904 gnd.n2903 240.244
R4952 gnd.n2900 gnd.n2899 240.244
R4953 gnd.n2896 gnd.n2895 240.244
R4954 gnd.n2892 gnd.n2891 240.244
R4955 gnd.n2885 gnd.n2884 240.244
R4956 gnd.n2882 gnd.n2881 240.244
R4957 gnd.n2878 gnd.n2877 240.244
R4958 gnd.n2874 gnd.n2873 240.244
R4959 gnd.n2870 gnd.n2869 240.244
R4960 gnd.n2866 gnd.n2865 240.244
R4961 gnd.n2862 gnd.n2861 240.244
R4962 gnd.n2858 gnd.n2857 240.244
R4963 gnd.n2854 gnd.n2853 240.244
R4964 gnd.n2850 gnd.n2849 240.244
R4965 gnd.n6154 gnd.n6153 240.244
R4966 gnd.n6153 gnd.n2453 240.244
R4967 gnd.n2465 gnd.n2453 240.244
R4968 gnd.n4083 gnd.n2465 240.244
R4969 gnd.n4083 gnd.n2477 240.244
R4970 gnd.n4087 gnd.n2477 240.244
R4971 gnd.n4087 gnd.n2487 240.244
R4972 gnd.n4173 gnd.n2487 240.244
R4973 gnd.n4173 gnd.n2497 240.244
R4974 gnd.n4074 gnd.n2497 240.244
R4975 gnd.n4074 gnd.n2507 240.244
R4976 gnd.n4200 gnd.n2507 240.244
R4977 gnd.n4200 gnd.n2517 240.244
R4978 gnd.n4196 gnd.n2517 240.244
R4979 gnd.n4196 gnd.n2528 240.244
R4980 gnd.n4188 gnd.n2528 240.244
R4981 gnd.n4188 gnd.n2538 240.244
R4982 gnd.n4241 gnd.n2538 240.244
R4983 gnd.n4241 gnd.n4053 240.244
R4984 gnd.n4053 gnd.n4045 240.244
R4985 gnd.n4260 gnd.n4045 240.244
R4986 gnd.n4260 gnd.n4037 240.244
R4987 gnd.n4037 gnd.n4030 240.244
R4988 gnd.n4267 gnd.n4030 240.244
R4989 gnd.n4267 gnd.n4023 240.244
R4990 gnd.n4023 gnd.n2553 240.244
R4991 gnd.n4016 gnd.n2553 240.244
R4992 gnd.n4016 gnd.n2564 240.244
R4993 gnd.n4326 gnd.n2564 240.244
R4994 gnd.n4326 gnd.n2574 240.244
R4995 gnd.n4330 gnd.n2574 240.244
R4996 gnd.n4330 gnd.n2583 240.244
R4997 gnd.n4340 gnd.n2583 240.244
R4998 gnd.n4340 gnd.n2594 240.244
R4999 gnd.n3999 gnd.n2594 240.244
R5000 gnd.n3999 gnd.n2603 240.244
R5001 gnd.n4347 gnd.n2603 240.244
R5002 gnd.n4347 gnd.n2614 240.244
R5003 gnd.n4351 gnd.n2614 240.244
R5004 gnd.n4351 gnd.n2624 240.244
R5005 gnd.n6042 gnd.n2624 240.244
R5006 gnd.n6042 gnd.n2633 240.244
R5007 gnd.n2382 gnd.n2381 240.244
R5008 gnd.n6269 gnd.n2381 240.244
R5009 gnd.n6267 gnd.n6266 240.244
R5010 gnd.n6263 gnd.n6262 240.244
R5011 gnd.n6259 gnd.n6258 240.244
R5012 gnd.n6255 gnd.n6254 240.244
R5013 gnd.n6251 gnd.n6250 240.244
R5014 gnd.n6247 gnd.n6246 240.244
R5015 gnd.n6243 gnd.n6242 240.244
R5016 gnd.n6238 gnd.n6237 240.244
R5017 gnd.n6234 gnd.n6233 240.244
R5018 gnd.n6230 gnd.n6229 240.244
R5019 gnd.n6226 gnd.n6225 240.244
R5020 gnd.n6222 gnd.n6221 240.244
R5021 gnd.n6218 gnd.n6217 240.244
R5022 gnd.n6214 gnd.n6213 240.244
R5023 gnd.n6210 gnd.n6209 240.244
R5024 gnd.n6206 gnd.n6205 240.244
R5025 gnd.n6202 gnd.n6201 240.244
R5026 gnd.n6198 gnd.n6197 240.244
R5027 gnd.n6194 gnd.n6193 240.244
R5028 gnd.n6190 gnd.n6189 240.244
R5029 gnd.n6186 gnd.n6185 240.244
R5030 gnd.n6182 gnd.n6181 240.244
R5031 gnd.n6178 gnd.n6177 240.244
R5032 gnd.n6174 gnd.n6173 240.244
R5033 gnd.n6170 gnd.n6169 240.244
R5034 gnd.n6166 gnd.n6165 240.244
R5035 gnd.n6162 gnd.n6161 240.244
R5036 gnd.n6151 gnd.n2383 240.244
R5037 gnd.n6151 gnd.n2456 240.244
R5038 gnd.n6147 gnd.n2456 240.244
R5039 gnd.n6147 gnd.n2463 240.244
R5040 gnd.n6139 gnd.n2463 240.244
R5041 gnd.n6139 gnd.n2480 240.244
R5042 gnd.n6135 gnd.n2480 240.244
R5043 gnd.n6135 gnd.n2486 240.244
R5044 gnd.n6127 gnd.n2486 240.244
R5045 gnd.n6127 gnd.n2499 240.244
R5046 gnd.n6123 gnd.n2499 240.244
R5047 gnd.n6123 gnd.n2505 240.244
R5048 gnd.n6115 gnd.n2505 240.244
R5049 gnd.n6115 gnd.n2520 240.244
R5050 gnd.n6111 gnd.n2520 240.244
R5051 gnd.n6111 gnd.n2526 240.244
R5052 gnd.n6103 gnd.n2526 240.244
R5053 gnd.n6103 gnd.n2540 240.244
R5054 gnd.n4250 gnd.n2540 240.244
R5055 gnd.n4250 gnd.n4249 240.244
R5056 gnd.n4249 gnd.n4033 240.244
R5057 gnd.n4276 gnd.n4033 240.244
R5058 gnd.n4280 gnd.n4276 240.244
R5059 gnd.n4280 gnd.n4277 240.244
R5060 gnd.n4277 gnd.n2550 240.244
R5061 gnd.n6097 gnd.n2550 240.244
R5062 gnd.n6097 gnd.n2551 240.244
R5063 gnd.n6089 gnd.n2551 240.244
R5064 gnd.n6089 gnd.n2567 240.244
R5065 gnd.n6085 gnd.n2567 240.244
R5066 gnd.n6085 gnd.n2572 240.244
R5067 gnd.n6077 gnd.n2572 240.244
R5068 gnd.n6077 gnd.n2586 240.244
R5069 gnd.n6073 gnd.n2586 240.244
R5070 gnd.n6073 gnd.n2592 240.244
R5071 gnd.n6065 gnd.n2592 240.244
R5072 gnd.n6065 gnd.n2606 240.244
R5073 gnd.n6061 gnd.n2606 240.244
R5074 gnd.n6061 gnd.n2612 240.244
R5075 gnd.n6053 gnd.n2612 240.244
R5076 gnd.n6053 gnd.n2626 240.244
R5077 gnd.n6049 gnd.n2626 240.244
R5078 gnd.n6322 gnd.n6283 240.244
R5079 gnd.n6315 gnd.n6314 240.244
R5080 gnd.n6312 gnd.n6311 240.244
R5081 gnd.n6308 gnd.n6307 240.244
R5082 gnd.n6304 gnd.n6303 240.244
R5083 gnd.n6300 gnd.n6299 240.244
R5084 gnd.n6296 gnd.n1056 240.244
R5085 gnd.n6326 gnd.n6325 240.244
R5086 gnd.n1749 gnd.n1357 240.244
R5087 gnd.n1357 gnd.n1348 240.244
R5088 gnd.n1770 gnd.n1348 240.244
R5089 gnd.n1770 gnd.n1341 240.244
R5090 gnd.n1780 gnd.n1341 240.244
R5091 gnd.n1780 gnd.n1332 240.244
R5092 gnd.n1332 gnd.n1321 240.244
R5093 gnd.n1801 gnd.n1321 240.244
R5094 gnd.n1801 gnd.n1315 240.244
R5095 gnd.n1811 gnd.n1315 240.244
R5096 gnd.n1811 gnd.n1306 240.244
R5097 gnd.n1306 gnd.n1295 240.244
R5098 gnd.n1832 gnd.n1295 240.244
R5099 gnd.n1832 gnd.n1289 240.244
R5100 gnd.n1842 gnd.n1289 240.244
R5101 gnd.n1842 gnd.n1280 240.244
R5102 gnd.n1280 gnd.n1270 240.244
R5103 gnd.n1863 gnd.n1270 240.244
R5104 gnd.n1863 gnd.n1263 240.244
R5105 gnd.n1873 gnd.n1263 240.244
R5106 gnd.n1873 gnd.n1254 240.244
R5107 gnd.n1254 gnd.n1245 240.244
R5108 gnd.n1894 gnd.n1245 240.244
R5109 gnd.n1894 gnd.n1238 240.244
R5110 gnd.n1904 gnd.n1238 240.244
R5111 gnd.n1904 gnd.n1229 240.244
R5112 gnd.n1229 gnd.n1220 240.244
R5113 gnd.n1925 gnd.n1220 240.244
R5114 gnd.n1925 gnd.n1213 240.244
R5115 gnd.n1935 gnd.n1213 240.244
R5116 gnd.n1935 gnd.n1202 240.244
R5117 gnd.n1202 gnd.n1194 240.244
R5118 gnd.n1953 gnd.n1194 240.244
R5119 gnd.n1954 gnd.n1953 240.244
R5120 gnd.n1954 gnd.n1180 240.244
R5121 gnd.n1958 gnd.n1180 240.244
R5122 gnd.n1958 gnd.n1170 240.244
R5123 gnd.n1170 gnd.n1162 240.244
R5124 gnd.n2037 gnd.n1162 240.244
R5125 gnd.n2037 gnd.n979 240.244
R5126 gnd.n1155 gnd.n979 240.244
R5127 gnd.n1155 gnd.n990 240.244
R5128 gnd.n2052 gnd.n990 240.244
R5129 gnd.n2053 gnd.n2052 240.244
R5130 gnd.n2053 gnd.n1003 240.244
R5131 gnd.n1152 gnd.n1003 240.244
R5132 gnd.n1152 gnd.n1016 240.244
R5133 gnd.n2321 gnd.n1016 240.244
R5134 gnd.n2322 gnd.n2321 240.244
R5135 gnd.n2322 gnd.n1029 240.244
R5136 gnd.n2330 gnd.n1029 240.244
R5137 gnd.n2330 gnd.n1041 240.244
R5138 gnd.n6333 gnd.n1041 240.244
R5139 gnd.n1686 gnd.n1685 240.244
R5140 gnd.n1730 gnd.n1685 240.244
R5141 gnd.n1728 gnd.n1727 240.244
R5142 gnd.n1724 gnd.n1723 240.244
R5143 gnd.n1720 gnd.n1719 240.244
R5144 gnd.n1716 gnd.n1715 240.244
R5145 gnd.n1712 gnd.n1711 240.244
R5146 gnd.n1708 gnd.n1707 240.244
R5147 gnd.n1760 gnd.n1355 240.244
R5148 gnd.n1760 gnd.n1350 240.244
R5149 gnd.n1768 gnd.n1350 240.244
R5150 gnd.n1768 gnd.n1351 240.244
R5151 gnd.n1351 gnd.n1330 240.244
R5152 gnd.n1791 gnd.n1330 240.244
R5153 gnd.n1791 gnd.n1324 240.244
R5154 gnd.n1799 gnd.n1324 240.244
R5155 gnd.n1799 gnd.n1326 240.244
R5156 gnd.n1326 gnd.n1304 240.244
R5157 gnd.n1822 gnd.n1304 240.244
R5158 gnd.n1822 gnd.n1298 240.244
R5159 gnd.n1830 gnd.n1298 240.244
R5160 gnd.n1830 gnd.n1300 240.244
R5161 gnd.n1300 gnd.n1278 240.244
R5162 gnd.n1853 gnd.n1278 240.244
R5163 gnd.n1853 gnd.n1273 240.244
R5164 gnd.n1861 gnd.n1273 240.244
R5165 gnd.n1861 gnd.n1274 240.244
R5166 gnd.n1274 gnd.n1252 240.244
R5167 gnd.n1884 gnd.n1252 240.244
R5168 gnd.n1884 gnd.n1247 240.244
R5169 gnd.n1892 gnd.n1247 240.244
R5170 gnd.n1892 gnd.n1248 240.244
R5171 gnd.n1248 gnd.n1227 240.244
R5172 gnd.n1915 gnd.n1227 240.244
R5173 gnd.n1915 gnd.n1222 240.244
R5174 gnd.n1923 gnd.n1222 240.244
R5175 gnd.n1923 gnd.n1223 240.244
R5176 gnd.n1223 gnd.n1200 240.244
R5177 gnd.n1945 gnd.n1200 240.244
R5178 gnd.n1945 gnd.n1196 240.244
R5179 gnd.n1951 gnd.n1196 240.244
R5180 gnd.n1951 gnd.n1178 240.244
R5181 gnd.n2015 gnd.n1178 240.244
R5182 gnd.n2015 gnd.n1172 240.244
R5183 gnd.n2024 gnd.n1172 240.244
R5184 gnd.n2024 gnd.n1174 240.244
R5185 gnd.n1174 gnd.n981 240.244
R5186 gnd.n6373 gnd.n981 240.244
R5187 gnd.n6373 gnd.n982 240.244
R5188 gnd.n6369 gnd.n982 240.244
R5189 gnd.n6369 gnd.n988 240.244
R5190 gnd.n1005 gnd.n988 240.244
R5191 gnd.n6359 gnd.n1005 240.244
R5192 gnd.n6359 gnd.n1006 240.244
R5193 gnd.n6355 gnd.n1006 240.244
R5194 gnd.n6355 gnd.n1014 240.244
R5195 gnd.n1030 gnd.n1014 240.244
R5196 gnd.n6345 gnd.n1030 240.244
R5197 gnd.n6345 gnd.n1031 240.244
R5198 gnd.n6341 gnd.n1031 240.244
R5199 gnd.n6341 gnd.n1039 240.244
R5200 gnd.n7282 gnd.n172 240.244
R5201 gnd.n7285 gnd.n7284 240.244
R5202 gnd.n7292 gnd.n7291 240.244
R5203 gnd.n7295 gnd.n7294 240.244
R5204 gnd.n7302 gnd.n7301 240.244
R5205 gnd.n7305 gnd.n7304 240.244
R5206 gnd.n7312 gnd.n7311 240.244
R5207 gnd.n7315 gnd.n7314 240.244
R5208 gnd.n7322 gnd.n7321 240.244
R5209 gnd.n5344 gnd.n3268 240.244
R5210 gnd.n5344 gnd.n3277 240.244
R5211 gnd.n5307 gnd.n3277 240.244
R5212 gnd.n5307 gnd.n3293 240.244
R5213 gnd.n5308 gnd.n3293 240.244
R5214 gnd.n5308 gnd.n3306 240.244
R5215 gnd.n5311 gnd.n3306 240.244
R5216 gnd.n5311 gnd.n3316 240.244
R5217 gnd.n5329 gnd.n3316 240.244
R5218 gnd.n5329 gnd.n3326 240.244
R5219 gnd.n5389 gnd.n3326 240.244
R5220 gnd.n5389 gnd.n3336 240.244
R5221 gnd.n5395 gnd.n3336 240.244
R5222 gnd.n5395 gnd.n3346 240.244
R5223 gnd.n5404 gnd.n3346 240.244
R5224 gnd.n5404 gnd.n3353 240.244
R5225 gnd.n5414 gnd.n3353 240.244
R5226 gnd.n5414 gnd.n3363 240.244
R5227 gnd.n3369 gnd.n3363 240.244
R5228 gnd.n3389 gnd.n3369 240.244
R5229 gnd.n3389 gnd.n3388 240.244
R5230 gnd.n3388 gnd.n70 240.244
R5231 gnd.n7414 gnd.n70 240.244
R5232 gnd.n7414 gnd.n72 240.244
R5233 gnd.n5441 gnd.n72 240.244
R5234 gnd.n5441 gnd.n92 240.244
R5235 gnd.n397 gnd.n92 240.244
R5236 gnd.n397 gnd.n103 240.244
R5237 gnd.n7234 gnd.n103 240.244
R5238 gnd.n7234 gnd.n113 240.244
R5239 gnd.n7240 gnd.n113 240.244
R5240 gnd.n7240 gnd.n122 240.244
R5241 gnd.n7249 gnd.n122 240.244
R5242 gnd.n7249 gnd.n133 240.244
R5243 gnd.n7339 gnd.n133 240.244
R5244 gnd.n7339 gnd.n142 240.244
R5245 gnd.n7335 gnd.n142 240.244
R5246 gnd.n7335 gnd.n152 240.244
R5247 gnd.n7332 gnd.n152 240.244
R5248 gnd.n7332 gnd.n161 240.244
R5249 gnd.n7329 gnd.n161 240.244
R5250 gnd.n7329 gnd.n170 240.244
R5251 gnd.n3112 gnd.n3111 240.244
R5252 gnd.n3187 gnd.n3119 240.244
R5253 gnd.n3190 gnd.n3120 240.244
R5254 gnd.n3128 gnd.n3127 240.244
R5255 gnd.n3192 gnd.n3135 240.244
R5256 gnd.n3195 gnd.n3136 240.244
R5257 gnd.n3144 gnd.n3143 240.244
R5258 gnd.n3197 gnd.n3153 240.244
R5259 gnd.n5651 gnd.n3156 240.244
R5260 gnd.n5527 gnd.n3271 240.244
R5261 gnd.n3279 gnd.n3271 240.244
R5262 gnd.n3295 gnd.n3279 240.244
R5263 gnd.n5513 gnd.n3295 240.244
R5264 gnd.n5513 gnd.n3296 240.244
R5265 gnd.n5509 gnd.n3296 240.244
R5266 gnd.n5509 gnd.n3303 240.244
R5267 gnd.n5501 gnd.n3303 240.244
R5268 gnd.n5501 gnd.n3318 240.244
R5269 gnd.n5497 gnd.n3318 240.244
R5270 gnd.n5497 gnd.n3323 240.244
R5271 gnd.n5489 gnd.n3323 240.244
R5272 gnd.n5489 gnd.n3338 240.244
R5273 gnd.n5485 gnd.n3338 240.244
R5274 gnd.n5485 gnd.n3343 240.244
R5275 gnd.n5477 gnd.n3343 240.244
R5276 gnd.n5477 gnd.n3355 240.244
R5277 gnd.n5473 gnd.n3355 240.244
R5278 gnd.n5473 gnd.n3360 240.244
R5279 gnd.n5423 gnd.n3360 240.244
R5280 gnd.n5423 gnd.n3380 240.244
R5281 gnd.n5457 gnd.n3380 240.244
R5282 gnd.n5457 gnd.n76 240.244
R5283 gnd.n5453 gnd.n76 240.244
R5284 gnd.n5453 gnd.n94 240.244
R5285 gnd.n7404 gnd.n94 240.244
R5286 gnd.n7404 gnd.n95 240.244
R5287 gnd.n7400 gnd.n95 240.244
R5288 gnd.n7400 gnd.n101 240.244
R5289 gnd.n7392 gnd.n101 240.244
R5290 gnd.n7392 gnd.n114 240.244
R5291 gnd.n7388 gnd.n114 240.244
R5292 gnd.n7388 gnd.n119 240.244
R5293 gnd.n7380 gnd.n119 240.244
R5294 gnd.n7380 gnd.n135 240.244
R5295 gnd.n7376 gnd.n135 240.244
R5296 gnd.n7376 gnd.n140 240.244
R5297 gnd.n7368 gnd.n140 240.244
R5298 gnd.n7368 gnd.n154 240.244
R5299 gnd.n7364 gnd.n154 240.244
R5300 gnd.n7364 gnd.n159 240.244
R5301 gnd.n7356 gnd.n159 240.244
R5302 gnd.n1085 gnd.n1045 240.244
R5303 gnd.n1093 gnd.n1092 240.244
R5304 gnd.n1096 gnd.n1095 240.244
R5305 gnd.n1103 gnd.n1102 240.244
R5306 gnd.n1106 gnd.n1105 240.244
R5307 gnd.n1113 gnd.n1112 240.244
R5308 gnd.n1116 gnd.n1115 240.244
R5309 gnd.n1123 gnd.n1122 240.244
R5310 gnd.n1126 gnd.n1125 240.244
R5311 gnd.n1133 gnd.n1132 240.244
R5312 gnd.n1136 gnd.n1135 240.244
R5313 gnd.n1143 gnd.n1142 240.244
R5314 gnd.n1145 gnd.n1069 240.244
R5315 gnd.n1504 gnd.n1400 240.244
R5316 gnd.n1510 gnd.n1400 240.244
R5317 gnd.n1510 gnd.n1392 240.244
R5318 gnd.n1520 gnd.n1392 240.244
R5319 gnd.n1520 gnd.n1388 240.244
R5320 gnd.n1526 gnd.n1388 240.244
R5321 gnd.n1526 gnd.n1379 240.244
R5322 gnd.n1536 gnd.n1379 240.244
R5323 gnd.n1536 gnd.n1374 240.244
R5324 gnd.n1677 gnd.n1374 240.244
R5325 gnd.n1677 gnd.n1375 240.244
R5326 gnd.n1375 gnd.n1367 240.244
R5327 gnd.n1672 gnd.n1367 240.244
R5328 gnd.n1672 gnd.n1358 240.244
R5329 gnd.n1669 gnd.n1358 240.244
R5330 gnd.n1669 gnd.n1668 240.244
R5331 gnd.n1668 gnd.n1343 240.244
R5332 gnd.n1663 gnd.n1343 240.244
R5333 gnd.n1663 gnd.n1333 240.244
R5334 gnd.n1660 gnd.n1333 240.244
R5335 gnd.n1660 gnd.n1659 240.244
R5336 gnd.n1659 gnd.n1316 240.244
R5337 gnd.n1655 gnd.n1316 240.244
R5338 gnd.n1655 gnd.n1307 240.244
R5339 gnd.n1652 gnd.n1307 240.244
R5340 gnd.n1652 gnd.n1651 240.244
R5341 gnd.n1651 gnd.n1290 240.244
R5342 gnd.n1647 gnd.n1290 240.244
R5343 gnd.n1647 gnd.n1281 240.244
R5344 gnd.n1592 gnd.n1281 240.244
R5345 gnd.n1593 gnd.n1592 240.244
R5346 gnd.n1593 gnd.n1265 240.244
R5347 gnd.n1589 gnd.n1265 240.244
R5348 gnd.n1589 gnd.n1255 240.244
R5349 gnd.n1585 gnd.n1255 240.244
R5350 gnd.n1585 gnd.n1584 240.244
R5351 gnd.n1584 gnd.n1240 240.244
R5352 gnd.n1579 gnd.n1240 240.244
R5353 gnd.n1579 gnd.n1230 240.244
R5354 gnd.n1576 gnd.n1230 240.244
R5355 gnd.n1576 gnd.n1574 240.244
R5356 gnd.n1574 gnd.n1215 240.244
R5357 gnd.n1570 gnd.n1215 240.244
R5358 gnd.n1570 gnd.n1203 240.244
R5359 gnd.n1203 gnd.n1185 240.244
R5360 gnd.n1967 gnd.n1185 240.244
R5361 gnd.n1967 gnd.n1181 240.244
R5362 gnd.n2012 gnd.n1181 240.244
R5363 gnd.n2012 gnd.n1169 240.244
R5364 gnd.n2008 gnd.n1169 240.244
R5365 gnd.n2008 gnd.n1161 240.244
R5366 gnd.n2005 gnd.n1161 240.244
R5367 gnd.n2005 gnd.n2004 240.244
R5368 gnd.n2004 gnd.n2003 240.244
R5369 gnd.n2003 gnd.n991 240.244
R5370 gnd.n1999 gnd.n991 240.244
R5371 gnd.n1999 gnd.n1002 240.244
R5372 gnd.n1995 gnd.n1002 240.244
R5373 gnd.n1995 gnd.n1994 240.244
R5374 gnd.n1994 gnd.n1017 240.244
R5375 gnd.n1990 gnd.n1017 240.244
R5376 gnd.n1990 gnd.n1028 240.244
R5377 gnd.n2333 gnd.n1028 240.244
R5378 gnd.n2334 gnd.n2333 240.244
R5379 gnd.n2334 gnd.n1042 240.244
R5380 gnd.n1496 gnd.n1494 240.244
R5381 gnd.n1494 gnd.n1493 240.244
R5382 gnd.n1490 gnd.n1489 240.244
R5383 gnd.n1487 gnd.n1413 240.244
R5384 gnd.n1483 gnd.n1481 240.244
R5385 gnd.n1479 gnd.n1419 240.244
R5386 gnd.n1475 gnd.n1473 240.244
R5387 gnd.n1471 gnd.n1425 240.244
R5388 gnd.n1467 gnd.n1465 240.244
R5389 gnd.n1463 gnd.n1431 240.244
R5390 gnd.n1459 gnd.n1457 240.244
R5391 gnd.n1455 gnd.n1437 240.244
R5392 gnd.n1450 gnd.n1448 240.244
R5393 gnd.n1502 gnd.n1398 240.244
R5394 gnd.n1512 gnd.n1398 240.244
R5395 gnd.n1512 gnd.n1394 240.244
R5396 gnd.n1518 gnd.n1394 240.244
R5397 gnd.n1518 gnd.n1386 240.244
R5398 gnd.n1528 gnd.n1386 240.244
R5399 gnd.n1528 gnd.n1382 240.244
R5400 gnd.n1534 gnd.n1382 240.244
R5401 gnd.n1534 gnd.n1373 240.244
R5402 gnd.n1739 gnd.n1373 240.244
R5403 gnd.n1739 gnd.n1368 240.244
R5404 gnd.n1746 gnd.n1368 240.244
R5405 gnd.n1746 gnd.n1360 240.244
R5406 gnd.n1757 gnd.n1360 240.244
R5407 gnd.n1757 gnd.n1361 240.244
R5408 gnd.n1361 gnd.n1344 240.244
R5409 gnd.n1777 gnd.n1344 240.244
R5410 gnd.n1777 gnd.n1335 240.244
R5411 gnd.n1788 gnd.n1335 240.244
R5412 gnd.n1788 gnd.n1336 240.244
R5413 gnd.n1336 gnd.n1317 240.244
R5414 gnd.n1808 gnd.n1317 240.244
R5415 gnd.n1808 gnd.n1309 240.244
R5416 gnd.n1819 gnd.n1309 240.244
R5417 gnd.n1819 gnd.n1310 240.244
R5418 gnd.n1310 gnd.n1291 240.244
R5419 gnd.n1839 gnd.n1291 240.244
R5420 gnd.n1839 gnd.n1283 240.244
R5421 gnd.n1850 gnd.n1283 240.244
R5422 gnd.n1850 gnd.n1284 240.244
R5423 gnd.n1284 gnd.n1266 240.244
R5424 gnd.n1870 gnd.n1266 240.244
R5425 gnd.n1870 gnd.n1257 240.244
R5426 gnd.n1881 gnd.n1257 240.244
R5427 gnd.n1881 gnd.n1258 240.244
R5428 gnd.n1258 gnd.n1241 240.244
R5429 gnd.n1901 gnd.n1241 240.244
R5430 gnd.n1901 gnd.n1232 240.244
R5431 gnd.n1912 gnd.n1232 240.244
R5432 gnd.n1912 gnd.n1233 240.244
R5433 gnd.n1233 gnd.n1216 240.244
R5434 gnd.n1932 gnd.n1216 240.244
R5435 gnd.n1932 gnd.n1205 240.244
R5436 gnd.n1942 gnd.n1205 240.244
R5437 gnd.n1942 gnd.n1187 240.244
R5438 gnd.n1965 gnd.n1187 240.244
R5439 gnd.n1965 gnd.n1188 240.244
R5440 gnd.n1188 gnd.n1167 240.244
R5441 gnd.n2027 gnd.n1167 240.244
R5442 gnd.n2027 gnd.n1159 240.244
R5443 gnd.n2040 gnd.n1159 240.244
R5444 gnd.n2041 gnd.n2040 240.244
R5445 gnd.n2042 gnd.n2041 240.244
R5446 gnd.n2042 gnd.n993 240.244
R5447 gnd.n6366 gnd.n993 240.244
R5448 gnd.n6366 gnd.n994 240.244
R5449 gnd.n6362 gnd.n994 240.244
R5450 gnd.n6362 gnd.n1000 240.244
R5451 gnd.n1019 gnd.n1000 240.244
R5452 gnd.n6352 gnd.n1019 240.244
R5453 gnd.n6352 gnd.n1020 240.244
R5454 gnd.n6348 gnd.n1020 240.244
R5455 gnd.n6348 gnd.n1026 240.244
R5456 gnd.n1044 gnd.n1026 240.244
R5457 gnd.n6338 gnd.n1044 240.244
R5458 gnd.n2683 gnd.n2636 240.244
R5459 gnd.n2740 gnd.n2684 240.244
R5460 gnd.n2694 gnd.n2693 240.244
R5461 gnd.n2742 gnd.n2701 240.244
R5462 gnd.n2745 gnd.n2702 240.244
R5463 gnd.n2712 gnd.n2711 240.244
R5464 gnd.n2747 gnd.n2719 240.244
R5465 gnd.n2750 gnd.n2720 240.244
R5466 gnd.n2737 gnd.n2732 240.244
R5467 gnd.n4153 gnd.n2454 240.244
R5468 gnd.n4156 gnd.n2454 240.244
R5469 gnd.n4156 gnd.n2466 240.244
R5470 gnd.n4161 gnd.n2466 240.244
R5471 gnd.n4161 gnd.n2478 240.244
R5472 gnd.n4164 gnd.n2478 240.244
R5473 gnd.n4164 gnd.n2488 240.244
R5474 gnd.n4171 gnd.n2488 240.244
R5475 gnd.n4171 gnd.n2498 240.244
R5476 gnd.n4206 gnd.n2498 240.244
R5477 gnd.n4206 gnd.n2508 240.244
R5478 gnd.n4202 gnd.n2508 240.244
R5479 gnd.n4202 gnd.n2518 240.244
R5480 gnd.n4194 gnd.n2518 240.244
R5481 gnd.n4194 gnd.n2529 240.244
R5482 gnd.n4190 gnd.n2529 240.244
R5483 gnd.n4190 gnd.n2539 240.244
R5484 gnd.n4051 gnd.n2539 240.244
R5485 gnd.n4252 gnd.n4051 240.244
R5486 gnd.n4252 gnd.n4047 240.244
R5487 gnd.n4258 gnd.n4047 240.244
R5488 gnd.n4258 gnd.n4028 240.244
R5489 gnd.n4282 gnd.n4028 240.244
R5490 gnd.n4282 gnd.n4024 240.244
R5491 gnd.n4288 gnd.n4024 240.244
R5492 gnd.n4288 gnd.n2554 240.244
R5493 gnd.n4318 gnd.n2554 240.244
R5494 gnd.n4318 gnd.n2565 240.244
R5495 gnd.n4324 gnd.n2565 240.244
R5496 gnd.n4324 gnd.n2575 240.244
R5497 gnd.n4332 gnd.n2575 240.244
R5498 gnd.n4332 gnd.n2584 240.244
R5499 gnd.n4338 gnd.n2584 240.244
R5500 gnd.n4338 gnd.n2595 240.244
R5501 gnd.n4362 gnd.n2595 240.244
R5502 gnd.n4362 gnd.n2604 240.244
R5503 gnd.n4004 gnd.n2604 240.244
R5504 gnd.n4004 gnd.n2615 240.244
R5505 gnd.n4353 gnd.n2615 240.244
R5506 gnd.n4353 gnd.n2625 240.244
R5507 gnd.n6040 gnd.n2625 240.244
R5508 gnd.n6040 gnd.n2634 240.244
R5509 gnd.n4113 gnd.n4112 240.244
R5510 gnd.n4119 gnd.n4118 240.244
R5511 gnd.n4123 gnd.n4122 240.244
R5512 gnd.n4129 gnd.n4128 240.244
R5513 gnd.n4133 gnd.n4132 240.244
R5514 gnd.n4139 gnd.n4138 240.244
R5515 gnd.n4143 gnd.n4142 240.244
R5516 gnd.n4100 gnd.n4099 240.244
R5517 gnd.n4095 gnd.n2379 240.244
R5518 gnd.n4108 gnd.n2455 240.244
R5519 gnd.n2468 gnd.n2455 240.244
R5520 gnd.n6145 gnd.n2468 240.244
R5521 gnd.n6145 gnd.n2469 240.244
R5522 gnd.n6141 gnd.n2469 240.244
R5523 gnd.n6141 gnd.n2476 240.244
R5524 gnd.n6133 gnd.n2476 240.244
R5525 gnd.n6133 gnd.n2490 240.244
R5526 gnd.n6129 gnd.n2490 240.244
R5527 gnd.n6129 gnd.n2495 240.244
R5528 gnd.n6121 gnd.n2495 240.244
R5529 gnd.n6121 gnd.n2510 240.244
R5530 gnd.n6117 gnd.n2510 240.244
R5531 gnd.n6117 gnd.n2515 240.244
R5532 gnd.n6109 gnd.n2515 240.244
R5533 gnd.n6109 gnd.n2531 240.244
R5534 gnd.n6105 gnd.n2531 240.244
R5535 gnd.n6105 gnd.n2536 240.244
R5536 gnd.n4055 gnd.n2536 240.244
R5537 gnd.n4247 gnd.n4055 240.244
R5538 gnd.n4247 gnd.n4038 240.244
R5539 gnd.n4274 gnd.n4038 240.244
R5540 gnd.n4274 gnd.n4032 240.244
R5541 gnd.n4270 gnd.n4032 240.244
R5542 gnd.n4270 gnd.n2556 240.244
R5543 gnd.n6095 gnd.n2556 240.244
R5544 gnd.n6095 gnd.n2557 240.244
R5545 gnd.n6091 gnd.n2557 240.244
R5546 gnd.n6091 gnd.n2563 240.244
R5547 gnd.n6083 gnd.n2563 240.244
R5548 gnd.n6083 gnd.n2576 240.244
R5549 gnd.n6079 gnd.n2576 240.244
R5550 gnd.n6079 gnd.n2581 240.244
R5551 gnd.n6071 gnd.n2581 240.244
R5552 gnd.n6071 gnd.n2597 240.244
R5553 gnd.n6067 gnd.n2597 240.244
R5554 gnd.n6067 gnd.n2602 240.244
R5555 gnd.n6059 gnd.n2602 240.244
R5556 gnd.n6059 gnd.n2617 240.244
R5557 gnd.n6055 gnd.n2617 240.244
R5558 gnd.n6055 gnd.n2622 240.244
R5559 gnd.n6047 gnd.n2622 240.244
R5560 gnd.n6545 gnd.n806 240.244
R5561 gnd.n6551 gnd.n806 240.244
R5562 gnd.n6551 gnd.n804 240.244
R5563 gnd.n6555 gnd.n804 240.244
R5564 gnd.n6555 gnd.n800 240.244
R5565 gnd.n6561 gnd.n800 240.244
R5566 gnd.n6561 gnd.n798 240.244
R5567 gnd.n6565 gnd.n798 240.244
R5568 gnd.n6565 gnd.n794 240.244
R5569 gnd.n6571 gnd.n794 240.244
R5570 gnd.n6571 gnd.n792 240.244
R5571 gnd.n6575 gnd.n792 240.244
R5572 gnd.n6575 gnd.n788 240.244
R5573 gnd.n6581 gnd.n788 240.244
R5574 gnd.n6581 gnd.n786 240.244
R5575 gnd.n6585 gnd.n786 240.244
R5576 gnd.n6585 gnd.n782 240.244
R5577 gnd.n6591 gnd.n782 240.244
R5578 gnd.n6591 gnd.n780 240.244
R5579 gnd.n6595 gnd.n780 240.244
R5580 gnd.n6595 gnd.n776 240.244
R5581 gnd.n6601 gnd.n776 240.244
R5582 gnd.n6601 gnd.n774 240.244
R5583 gnd.n6605 gnd.n774 240.244
R5584 gnd.n6605 gnd.n770 240.244
R5585 gnd.n6611 gnd.n770 240.244
R5586 gnd.n6611 gnd.n768 240.244
R5587 gnd.n6615 gnd.n768 240.244
R5588 gnd.n6615 gnd.n764 240.244
R5589 gnd.n6621 gnd.n764 240.244
R5590 gnd.n6621 gnd.n762 240.244
R5591 gnd.n6625 gnd.n762 240.244
R5592 gnd.n6625 gnd.n758 240.244
R5593 gnd.n6631 gnd.n758 240.244
R5594 gnd.n6631 gnd.n756 240.244
R5595 gnd.n6635 gnd.n756 240.244
R5596 gnd.n6635 gnd.n752 240.244
R5597 gnd.n6641 gnd.n752 240.244
R5598 gnd.n6641 gnd.n750 240.244
R5599 gnd.n6645 gnd.n750 240.244
R5600 gnd.n6645 gnd.n746 240.244
R5601 gnd.n6651 gnd.n746 240.244
R5602 gnd.n6651 gnd.n744 240.244
R5603 gnd.n6655 gnd.n744 240.244
R5604 gnd.n6655 gnd.n740 240.244
R5605 gnd.n6661 gnd.n740 240.244
R5606 gnd.n6661 gnd.n738 240.244
R5607 gnd.n6665 gnd.n738 240.244
R5608 gnd.n6665 gnd.n734 240.244
R5609 gnd.n6671 gnd.n734 240.244
R5610 gnd.n6671 gnd.n732 240.244
R5611 gnd.n6675 gnd.n732 240.244
R5612 gnd.n6675 gnd.n728 240.244
R5613 gnd.n6681 gnd.n728 240.244
R5614 gnd.n6681 gnd.n726 240.244
R5615 gnd.n6685 gnd.n726 240.244
R5616 gnd.n6685 gnd.n722 240.244
R5617 gnd.n6691 gnd.n722 240.244
R5618 gnd.n6691 gnd.n720 240.244
R5619 gnd.n6695 gnd.n720 240.244
R5620 gnd.n6695 gnd.n716 240.244
R5621 gnd.n6701 gnd.n716 240.244
R5622 gnd.n6701 gnd.n714 240.244
R5623 gnd.n6705 gnd.n714 240.244
R5624 gnd.n6705 gnd.n710 240.244
R5625 gnd.n6711 gnd.n710 240.244
R5626 gnd.n6711 gnd.n708 240.244
R5627 gnd.n6715 gnd.n708 240.244
R5628 gnd.n6715 gnd.n704 240.244
R5629 gnd.n6721 gnd.n704 240.244
R5630 gnd.n6721 gnd.n702 240.244
R5631 gnd.n6725 gnd.n702 240.244
R5632 gnd.n6725 gnd.n698 240.244
R5633 gnd.n6731 gnd.n698 240.244
R5634 gnd.n6731 gnd.n696 240.244
R5635 gnd.n6735 gnd.n696 240.244
R5636 gnd.n6735 gnd.n692 240.244
R5637 gnd.n6741 gnd.n692 240.244
R5638 gnd.n6741 gnd.n690 240.244
R5639 gnd.n6745 gnd.n690 240.244
R5640 gnd.n6745 gnd.n686 240.244
R5641 gnd.n6751 gnd.n686 240.244
R5642 gnd.n6751 gnd.n684 240.244
R5643 gnd.n6755 gnd.n684 240.244
R5644 gnd.n6755 gnd.n680 240.244
R5645 gnd.n6761 gnd.n680 240.244
R5646 gnd.n6761 gnd.n678 240.244
R5647 gnd.n6765 gnd.n678 240.244
R5648 gnd.n6765 gnd.n674 240.244
R5649 gnd.n6771 gnd.n674 240.244
R5650 gnd.n6771 gnd.n672 240.244
R5651 gnd.n6775 gnd.n672 240.244
R5652 gnd.n6775 gnd.n668 240.244
R5653 gnd.n6781 gnd.n668 240.244
R5654 gnd.n6781 gnd.n666 240.244
R5655 gnd.n6785 gnd.n666 240.244
R5656 gnd.n6785 gnd.n662 240.244
R5657 gnd.n6791 gnd.n662 240.244
R5658 gnd.n6791 gnd.n660 240.244
R5659 gnd.n6795 gnd.n660 240.244
R5660 gnd.n6795 gnd.n656 240.244
R5661 gnd.n6801 gnd.n656 240.244
R5662 gnd.n6801 gnd.n654 240.244
R5663 gnd.n6805 gnd.n654 240.244
R5664 gnd.n6805 gnd.n650 240.244
R5665 gnd.n6811 gnd.n650 240.244
R5666 gnd.n6811 gnd.n648 240.244
R5667 gnd.n6815 gnd.n648 240.244
R5668 gnd.n6815 gnd.n644 240.244
R5669 gnd.n6821 gnd.n644 240.244
R5670 gnd.n6821 gnd.n642 240.244
R5671 gnd.n6825 gnd.n642 240.244
R5672 gnd.n6825 gnd.n638 240.244
R5673 gnd.n6831 gnd.n638 240.244
R5674 gnd.n6831 gnd.n636 240.244
R5675 gnd.n6835 gnd.n636 240.244
R5676 gnd.n6835 gnd.n632 240.244
R5677 gnd.n6841 gnd.n632 240.244
R5678 gnd.n6841 gnd.n630 240.244
R5679 gnd.n6845 gnd.n630 240.244
R5680 gnd.n6845 gnd.n626 240.244
R5681 gnd.n6851 gnd.n626 240.244
R5682 gnd.n6851 gnd.n624 240.244
R5683 gnd.n6855 gnd.n624 240.244
R5684 gnd.n6855 gnd.n620 240.244
R5685 gnd.n6861 gnd.n620 240.244
R5686 gnd.n6861 gnd.n618 240.244
R5687 gnd.n6865 gnd.n618 240.244
R5688 gnd.n6865 gnd.n614 240.244
R5689 gnd.n6871 gnd.n614 240.244
R5690 gnd.n6871 gnd.n612 240.244
R5691 gnd.n6875 gnd.n612 240.244
R5692 gnd.n6875 gnd.n608 240.244
R5693 gnd.n6881 gnd.n608 240.244
R5694 gnd.n6881 gnd.n606 240.244
R5695 gnd.n6885 gnd.n606 240.244
R5696 gnd.n6885 gnd.n602 240.244
R5697 gnd.n6891 gnd.n602 240.244
R5698 gnd.n6891 gnd.n600 240.244
R5699 gnd.n6895 gnd.n600 240.244
R5700 gnd.n6895 gnd.n596 240.244
R5701 gnd.n6901 gnd.n596 240.244
R5702 gnd.n6901 gnd.n594 240.244
R5703 gnd.n6905 gnd.n594 240.244
R5704 gnd.n6905 gnd.n590 240.244
R5705 gnd.n6911 gnd.n590 240.244
R5706 gnd.n6911 gnd.n588 240.244
R5707 gnd.n6915 gnd.n588 240.244
R5708 gnd.n6915 gnd.n584 240.244
R5709 gnd.n6921 gnd.n584 240.244
R5710 gnd.n6921 gnd.n582 240.244
R5711 gnd.n6925 gnd.n582 240.244
R5712 gnd.n6925 gnd.n578 240.244
R5713 gnd.n6931 gnd.n578 240.244
R5714 gnd.n6931 gnd.n576 240.244
R5715 gnd.n6935 gnd.n576 240.244
R5716 gnd.n6935 gnd.n572 240.244
R5717 gnd.n6941 gnd.n572 240.244
R5718 gnd.n6941 gnd.n570 240.244
R5719 gnd.n6945 gnd.n570 240.244
R5720 gnd.n6945 gnd.n566 240.244
R5721 gnd.n6951 gnd.n566 240.244
R5722 gnd.n6951 gnd.n564 240.244
R5723 gnd.n6955 gnd.n564 240.244
R5724 gnd.n6955 gnd.n560 240.244
R5725 gnd.n6961 gnd.n560 240.244
R5726 gnd.n6961 gnd.n558 240.244
R5727 gnd.n6965 gnd.n558 240.244
R5728 gnd.n6965 gnd.n554 240.244
R5729 gnd.n6971 gnd.n554 240.244
R5730 gnd.n6971 gnd.n552 240.244
R5731 gnd.n6975 gnd.n552 240.244
R5732 gnd.n6975 gnd.n548 240.244
R5733 gnd.n6981 gnd.n548 240.244
R5734 gnd.n6981 gnd.n546 240.244
R5735 gnd.n6985 gnd.n546 240.244
R5736 gnd.n6985 gnd.n542 240.244
R5737 gnd.n6992 gnd.n542 240.244
R5738 gnd.n6992 gnd.n540 240.244
R5739 gnd.n6996 gnd.n540 240.244
R5740 gnd.n6996 gnd.n537 240.244
R5741 gnd.n7002 gnd.n535 240.244
R5742 gnd.n7006 gnd.n535 240.244
R5743 gnd.n7006 gnd.n531 240.244
R5744 gnd.n7012 gnd.n531 240.244
R5745 gnd.n7012 gnd.n529 240.244
R5746 gnd.n7016 gnd.n529 240.244
R5747 gnd.n7016 gnd.n525 240.244
R5748 gnd.n7022 gnd.n525 240.244
R5749 gnd.n7022 gnd.n523 240.244
R5750 gnd.n7026 gnd.n523 240.244
R5751 gnd.n7026 gnd.n519 240.244
R5752 gnd.n7032 gnd.n519 240.244
R5753 gnd.n7032 gnd.n517 240.244
R5754 gnd.n7036 gnd.n517 240.244
R5755 gnd.n7036 gnd.n513 240.244
R5756 gnd.n7042 gnd.n513 240.244
R5757 gnd.n7042 gnd.n511 240.244
R5758 gnd.n7046 gnd.n511 240.244
R5759 gnd.n7046 gnd.n507 240.244
R5760 gnd.n7052 gnd.n507 240.244
R5761 gnd.n7052 gnd.n505 240.244
R5762 gnd.n7056 gnd.n505 240.244
R5763 gnd.n7056 gnd.n501 240.244
R5764 gnd.n7062 gnd.n501 240.244
R5765 gnd.n7062 gnd.n499 240.244
R5766 gnd.n7066 gnd.n499 240.244
R5767 gnd.n7066 gnd.n495 240.244
R5768 gnd.n7072 gnd.n495 240.244
R5769 gnd.n7072 gnd.n493 240.244
R5770 gnd.n7076 gnd.n493 240.244
R5771 gnd.n7076 gnd.n489 240.244
R5772 gnd.n7082 gnd.n489 240.244
R5773 gnd.n7082 gnd.n487 240.244
R5774 gnd.n7086 gnd.n487 240.244
R5775 gnd.n7086 gnd.n483 240.244
R5776 gnd.n7092 gnd.n483 240.244
R5777 gnd.n7092 gnd.n481 240.244
R5778 gnd.n7096 gnd.n481 240.244
R5779 gnd.n7096 gnd.n477 240.244
R5780 gnd.n7102 gnd.n477 240.244
R5781 gnd.n7102 gnd.n475 240.244
R5782 gnd.n7106 gnd.n475 240.244
R5783 gnd.n7106 gnd.n471 240.244
R5784 gnd.n7112 gnd.n471 240.244
R5785 gnd.n7112 gnd.n469 240.244
R5786 gnd.n7116 gnd.n469 240.244
R5787 gnd.n7116 gnd.n465 240.244
R5788 gnd.n7122 gnd.n465 240.244
R5789 gnd.n7122 gnd.n463 240.244
R5790 gnd.n7126 gnd.n463 240.244
R5791 gnd.n7126 gnd.n459 240.244
R5792 gnd.n7132 gnd.n459 240.244
R5793 gnd.n7132 gnd.n457 240.244
R5794 gnd.n7136 gnd.n457 240.244
R5795 gnd.n7136 gnd.n453 240.244
R5796 gnd.n7142 gnd.n453 240.244
R5797 gnd.n7142 gnd.n451 240.244
R5798 gnd.n7146 gnd.n451 240.244
R5799 gnd.n7146 gnd.n447 240.244
R5800 gnd.n7152 gnd.n447 240.244
R5801 gnd.n7152 gnd.n445 240.244
R5802 gnd.n7156 gnd.n445 240.244
R5803 gnd.n7156 gnd.n441 240.244
R5804 gnd.n7162 gnd.n441 240.244
R5805 gnd.n7162 gnd.n439 240.244
R5806 gnd.n7166 gnd.n439 240.244
R5807 gnd.n7166 gnd.n435 240.244
R5808 gnd.n7172 gnd.n435 240.244
R5809 gnd.n7172 gnd.n433 240.244
R5810 gnd.n7176 gnd.n433 240.244
R5811 gnd.n7176 gnd.n429 240.244
R5812 gnd.n7182 gnd.n429 240.244
R5813 gnd.n7182 gnd.n427 240.244
R5814 gnd.n7186 gnd.n427 240.244
R5815 gnd.n7186 gnd.n423 240.244
R5816 gnd.n7192 gnd.n423 240.244
R5817 gnd.n7192 gnd.n421 240.244
R5818 gnd.n7196 gnd.n421 240.244
R5819 gnd.n7196 gnd.n417 240.244
R5820 gnd.n7202 gnd.n417 240.244
R5821 gnd.n7202 gnd.n415 240.244
R5822 gnd.n7207 gnd.n415 240.244
R5823 gnd.n7207 gnd.n411 240.244
R5824 gnd.n7213 gnd.n411 240.244
R5825 gnd.n4209 gnd.n4068 240.244
R5826 gnd.n4210 gnd.n4209 240.244
R5827 gnd.n4211 gnd.n4210 240.244
R5828 gnd.n4211 gnd.n4064 240.244
R5829 gnd.n4218 gnd.n4064 240.244
R5830 gnd.n4219 gnd.n4218 240.244
R5831 gnd.n4220 gnd.n4219 240.244
R5832 gnd.n4220 gnd.n4060 240.244
R5833 gnd.n4238 gnd.n4060 240.244
R5834 gnd.n4238 gnd.n4061 240.244
R5835 gnd.n4233 gnd.n4061 240.244
R5836 gnd.n4233 gnd.n4232 240.244
R5837 gnd.n4232 gnd.n4231 240.244
R5838 gnd.n4231 gnd.n4225 240.244
R5839 gnd.n4225 gnd.n4020 240.244
R5840 gnd.n4291 gnd.n4020 240.244
R5841 gnd.n4292 gnd.n4291 240.244
R5842 gnd.n4292 gnd.n4017 240.244
R5843 gnd.n4315 gnd.n4017 240.244
R5844 gnd.n4315 gnd.n4018 240.244
R5845 gnd.n4311 gnd.n4018 240.244
R5846 gnd.n4311 gnd.n4310 240.244
R5847 gnd.n4310 gnd.n4309 240.244
R5848 gnd.n4309 gnd.n4300 240.244
R5849 gnd.n4305 gnd.n4300 240.244
R5850 gnd.n4305 gnd.n3998 240.244
R5851 gnd.n4365 gnd.n3998 240.244
R5852 gnd.n4365 gnd.n3994 240.244
R5853 gnd.n4371 gnd.n3994 240.244
R5854 gnd.n4372 gnd.n4371 240.244
R5855 gnd.n4373 gnd.n4372 240.244
R5856 gnd.n4373 gnd.n3990 240.244
R5857 gnd.n4379 gnd.n3990 240.244
R5858 gnd.n4380 gnd.n4379 240.244
R5859 gnd.n4381 gnd.n4380 240.244
R5860 gnd.n4381 gnd.n3986 240.244
R5861 gnd.n4388 gnd.n3986 240.244
R5862 gnd.n4389 gnd.n4388 240.244
R5863 gnd.n4390 gnd.n4389 240.244
R5864 gnd.n4390 gnd.n3982 240.244
R5865 gnd.n4396 gnd.n3982 240.244
R5866 gnd.n4396 gnd.n3922 240.244
R5867 gnd.n4406 gnd.n3922 240.244
R5868 gnd.n4406 gnd.n3918 240.244
R5869 gnd.n4412 gnd.n3918 240.244
R5870 gnd.n4412 gnd.n3908 240.244
R5871 gnd.n4422 gnd.n3908 240.244
R5872 gnd.n4422 gnd.n3904 240.244
R5873 gnd.n4428 gnd.n3904 240.244
R5874 gnd.n4428 gnd.n3894 240.244
R5875 gnd.n4438 gnd.n3894 240.244
R5876 gnd.n4438 gnd.n3890 240.244
R5877 gnd.n4444 gnd.n3890 240.244
R5878 gnd.n4444 gnd.n3880 240.244
R5879 gnd.n4454 gnd.n3880 240.244
R5880 gnd.n4454 gnd.n3876 240.244
R5881 gnd.n4460 gnd.n3876 240.244
R5882 gnd.n4460 gnd.n3863 240.244
R5883 gnd.n4481 gnd.n3863 240.244
R5884 gnd.n4481 gnd.n3858 240.244
R5885 gnd.n4490 gnd.n3858 240.244
R5886 gnd.n4490 gnd.n3859 240.244
R5887 gnd.n3859 gnd.n2979 240.244
R5888 gnd.n5839 gnd.n2979 240.244
R5889 gnd.n5839 gnd.n2980 240.244
R5890 gnd.n5835 gnd.n2980 240.244
R5891 gnd.n5835 gnd.n2986 240.244
R5892 gnd.n4522 gnd.n2986 240.244
R5893 gnd.n4522 gnd.n4516 240.244
R5894 gnd.n4516 gnd.n3746 240.244
R5895 gnd.n4572 gnd.n3746 240.244
R5896 gnd.n4572 gnd.n3741 240.244
R5897 gnd.n4580 gnd.n3741 240.244
R5898 gnd.n4580 gnd.n3742 240.244
R5899 gnd.n3742 gnd.n3724 240.244
R5900 gnd.n4612 gnd.n3724 240.244
R5901 gnd.n4612 gnd.n3720 240.244
R5902 gnd.n4618 gnd.n3720 240.244
R5903 gnd.n4618 gnd.n3698 240.244
R5904 gnd.n4656 gnd.n3698 240.244
R5905 gnd.n4656 gnd.n3693 240.244
R5906 gnd.n4664 gnd.n3693 240.244
R5907 gnd.n4664 gnd.n3694 240.244
R5908 gnd.n3694 gnd.n3678 240.244
R5909 gnd.n4708 gnd.n3678 240.244
R5910 gnd.n4708 gnd.n3673 240.244
R5911 gnd.n4725 gnd.n3673 240.244
R5912 gnd.n4725 gnd.n3674 240.244
R5913 gnd.n4721 gnd.n3674 240.244
R5914 gnd.n4721 gnd.n4720 240.244
R5915 gnd.n4720 gnd.n4719 240.244
R5916 gnd.n4719 gnd.n3640 240.244
R5917 gnd.n4770 gnd.n3640 240.244
R5918 gnd.n4770 gnd.n3636 240.244
R5919 gnd.n4776 gnd.n3636 240.244
R5920 gnd.n4776 gnd.n3618 240.244
R5921 gnd.n4830 gnd.n3618 240.244
R5922 gnd.n4830 gnd.n3614 240.244
R5923 gnd.n4836 gnd.n3614 240.244
R5924 gnd.n4836 gnd.n3600 240.244
R5925 gnd.n4858 gnd.n3600 240.244
R5926 gnd.n4858 gnd.n3596 240.244
R5927 gnd.n4864 gnd.n3596 240.244
R5928 gnd.n4864 gnd.n3582 240.244
R5929 gnd.n4883 gnd.n3582 240.244
R5930 gnd.n4883 gnd.n3577 240.244
R5931 gnd.n4891 gnd.n3577 240.244
R5932 gnd.n4891 gnd.n3578 240.244
R5933 gnd.n3578 gnd.n3553 240.244
R5934 gnd.n4939 gnd.n3553 240.244
R5935 gnd.n4939 gnd.n3548 240.244
R5936 gnd.n4947 gnd.n3548 240.244
R5937 gnd.n4947 gnd.n3549 240.244
R5938 gnd.n3549 gnd.n3522 240.244
R5939 gnd.n5170 gnd.n3522 240.244
R5940 gnd.n5170 gnd.n3518 240.244
R5941 gnd.n5176 gnd.n3518 240.244
R5942 gnd.n5176 gnd.n3510 240.244
R5943 gnd.n5188 gnd.n3510 240.244
R5944 gnd.n5188 gnd.n3506 240.244
R5945 gnd.n5194 gnd.n3506 240.244
R5946 gnd.n5194 gnd.n3499 240.244
R5947 gnd.n5205 gnd.n3499 240.244
R5948 gnd.n5205 gnd.n3495 240.244
R5949 gnd.n5211 gnd.n3495 240.244
R5950 gnd.n5211 gnd.n3487 240.244
R5951 gnd.n5222 gnd.n3487 240.244
R5952 gnd.n5222 gnd.n3483 240.244
R5953 gnd.n5228 gnd.n3483 240.244
R5954 gnd.n5228 gnd.n3475 240.244
R5955 gnd.n5239 gnd.n3475 240.244
R5956 gnd.n5239 gnd.n3471 240.244
R5957 gnd.n5245 gnd.n3471 240.244
R5958 gnd.n5245 gnd.n3463 240.244
R5959 gnd.n5256 gnd.n3463 240.244
R5960 gnd.n5256 gnd.n3459 240.244
R5961 gnd.n5265 gnd.n3459 240.244
R5962 gnd.n5265 gnd.n3451 240.244
R5963 gnd.n5276 gnd.n3451 240.244
R5964 gnd.n5277 gnd.n5276 240.244
R5965 gnd.n5277 gnd.n3089 240.244
R5966 gnd.n3446 gnd.n3089 240.244
R5967 gnd.n5295 gnd.n3446 240.244
R5968 gnd.n5295 gnd.n3447 240.244
R5969 gnd.n5291 gnd.n3447 240.244
R5970 gnd.n5291 gnd.n5290 240.244
R5971 gnd.n5290 gnd.n5289 240.244
R5972 gnd.n5289 gnd.n3415 240.244
R5973 gnd.n5347 gnd.n3415 240.244
R5974 gnd.n5347 gnd.n3411 240.244
R5975 gnd.n5353 gnd.n3411 240.244
R5976 gnd.n5354 gnd.n5353 240.244
R5977 gnd.n5355 gnd.n5354 240.244
R5978 gnd.n5355 gnd.n3407 240.244
R5979 gnd.n5361 gnd.n3407 240.244
R5980 gnd.n5362 gnd.n5361 240.244
R5981 gnd.n5363 gnd.n5362 240.244
R5982 gnd.n5363 gnd.n3402 240.244
R5983 gnd.n5386 gnd.n3402 240.244
R5984 gnd.n5386 gnd.n3403 240.244
R5985 gnd.n5382 gnd.n3403 240.244
R5986 gnd.n5382 gnd.n5381 240.244
R5987 gnd.n5381 gnd.n5380 240.244
R5988 gnd.n5380 gnd.n5371 240.244
R5989 gnd.n5375 gnd.n5371 240.244
R5990 gnd.n5375 gnd.n3370 240.244
R5991 gnd.n5465 gnd.n3370 240.244
R5992 gnd.n5465 gnd.n3371 240.244
R5993 gnd.n5460 gnd.n3371 240.244
R5994 gnd.n5460 gnd.n3374 240.244
R5995 gnd.n5443 gnd.n3374 240.244
R5996 gnd.n5450 gnd.n5443 240.244
R5997 gnd.n5450 gnd.n5444 240.244
R5998 gnd.n5444 gnd.n398 240.244
R5999 gnd.n7224 gnd.n398 240.244
R6000 gnd.n7224 gnd.n399 240.244
R6001 gnd.n7220 gnd.n399 240.244
R6002 gnd.n7220 gnd.n7219 240.244
R6003 gnd.n7219 gnd.n7218 240.244
R6004 gnd.n7218 gnd.n406 240.244
R6005 gnd.n7214 gnd.n406 240.244
R6006 gnd.n6541 gnd.n809 240.244
R6007 gnd.n6541 gnd.n811 240.244
R6008 gnd.n6537 gnd.n811 240.244
R6009 gnd.n6537 gnd.n817 240.244
R6010 gnd.n6533 gnd.n817 240.244
R6011 gnd.n6533 gnd.n819 240.244
R6012 gnd.n6529 gnd.n819 240.244
R6013 gnd.n6529 gnd.n825 240.244
R6014 gnd.n6525 gnd.n825 240.244
R6015 gnd.n6525 gnd.n827 240.244
R6016 gnd.n6521 gnd.n827 240.244
R6017 gnd.n6521 gnd.n833 240.244
R6018 gnd.n6517 gnd.n833 240.244
R6019 gnd.n6517 gnd.n835 240.244
R6020 gnd.n6513 gnd.n835 240.244
R6021 gnd.n6513 gnd.n841 240.244
R6022 gnd.n6509 gnd.n841 240.244
R6023 gnd.n6509 gnd.n843 240.244
R6024 gnd.n6505 gnd.n843 240.244
R6025 gnd.n6505 gnd.n849 240.244
R6026 gnd.n6501 gnd.n849 240.244
R6027 gnd.n6501 gnd.n851 240.244
R6028 gnd.n6497 gnd.n851 240.244
R6029 gnd.n6497 gnd.n857 240.244
R6030 gnd.n6493 gnd.n857 240.244
R6031 gnd.n6493 gnd.n859 240.244
R6032 gnd.n6489 gnd.n859 240.244
R6033 gnd.n6489 gnd.n865 240.244
R6034 gnd.n6485 gnd.n865 240.244
R6035 gnd.n6485 gnd.n867 240.244
R6036 gnd.n6481 gnd.n867 240.244
R6037 gnd.n6481 gnd.n873 240.244
R6038 gnd.n6477 gnd.n873 240.244
R6039 gnd.n6477 gnd.n875 240.244
R6040 gnd.n6473 gnd.n875 240.244
R6041 gnd.n6473 gnd.n881 240.244
R6042 gnd.n6469 gnd.n881 240.244
R6043 gnd.n6469 gnd.n883 240.244
R6044 gnd.n6465 gnd.n883 240.244
R6045 gnd.n6465 gnd.n889 240.244
R6046 gnd.n6461 gnd.n889 240.244
R6047 gnd.n6461 gnd.n891 240.244
R6048 gnd.n6457 gnd.n891 240.244
R6049 gnd.n6457 gnd.n897 240.244
R6050 gnd.n6453 gnd.n897 240.244
R6051 gnd.n6453 gnd.n899 240.244
R6052 gnd.n6449 gnd.n899 240.244
R6053 gnd.n6449 gnd.n905 240.244
R6054 gnd.n6445 gnd.n905 240.244
R6055 gnd.n6445 gnd.n907 240.244
R6056 gnd.n6441 gnd.n907 240.244
R6057 gnd.n6441 gnd.n913 240.244
R6058 gnd.n6437 gnd.n913 240.244
R6059 gnd.n6437 gnd.n915 240.244
R6060 gnd.n6433 gnd.n915 240.244
R6061 gnd.n6433 gnd.n921 240.244
R6062 gnd.n6429 gnd.n921 240.244
R6063 gnd.n6429 gnd.n923 240.244
R6064 gnd.n6425 gnd.n923 240.244
R6065 gnd.n6425 gnd.n929 240.244
R6066 gnd.n6421 gnd.n929 240.244
R6067 gnd.n6421 gnd.n931 240.244
R6068 gnd.n6417 gnd.n931 240.244
R6069 gnd.n6417 gnd.n937 240.244
R6070 gnd.n6413 gnd.n937 240.244
R6071 gnd.n6413 gnd.n939 240.244
R6072 gnd.n6409 gnd.n939 240.244
R6073 gnd.n6409 gnd.n945 240.244
R6074 gnd.n6405 gnd.n945 240.244
R6075 gnd.n6405 gnd.n947 240.244
R6076 gnd.n6401 gnd.n947 240.244
R6077 gnd.n6401 gnd.n953 240.244
R6078 gnd.n6397 gnd.n953 240.244
R6079 gnd.n6397 gnd.n955 240.244
R6080 gnd.n6393 gnd.n955 240.244
R6081 gnd.n6393 gnd.n961 240.244
R6082 gnd.n6389 gnd.n961 240.244
R6083 gnd.n6389 gnd.n963 240.244
R6084 gnd.n6385 gnd.n963 240.244
R6085 gnd.n6385 gnd.n969 240.244
R6086 gnd.n6381 gnd.n969 240.244
R6087 gnd.n6381 gnd.n971 240.244
R6088 gnd.n6377 gnd.n971 240.244
R6089 gnd.n6377 gnd.n977 240.244
R6090 gnd.n3981 gnd.n2666 240.244
R6091 gnd.n3981 gnd.n3930 240.244
R6092 gnd.n3930 gnd.n3924 240.244
R6093 gnd.n3935 gnd.n3924 240.244
R6094 gnd.n3935 gnd.n3916 240.244
R6095 gnd.n3936 gnd.n3916 240.244
R6096 gnd.n3936 gnd.n3909 240.244
R6097 gnd.n3939 gnd.n3909 240.244
R6098 gnd.n3939 gnd.n3903 240.244
R6099 gnd.n3940 gnd.n3903 240.244
R6100 gnd.n3940 gnd.n3896 240.244
R6101 gnd.n3943 gnd.n3896 240.244
R6102 gnd.n3943 gnd.n3889 240.244
R6103 gnd.n3944 gnd.n3889 240.244
R6104 gnd.n3944 gnd.n3882 240.244
R6105 gnd.n3947 gnd.n3882 240.244
R6106 gnd.n3947 gnd.n3875 240.244
R6107 gnd.n3948 gnd.n3875 240.244
R6108 gnd.n3948 gnd.n3865 240.244
R6109 gnd.n3865 gnd.n3856 240.244
R6110 gnd.n4492 gnd.n3856 240.244
R6111 gnd.n4494 gnd.n4492 240.244
R6112 gnd.n4494 gnd.n4493 240.244
R6113 gnd.n4493 gnd.n2976 240.244
R6114 gnd.n4501 gnd.n2976 240.244
R6115 gnd.n4501 gnd.n2988 240.244
R6116 gnd.n3848 gnd.n2988 240.244
R6117 gnd.n4514 gnd.n3848 240.244
R6118 gnd.n4514 gnd.n3849 240.244
R6119 gnd.n4507 gnd.n3849 240.244
R6120 gnd.n4507 gnd.n3748 240.244
R6121 gnd.n3748 gnd.n3738 240.244
R6122 gnd.n4582 gnd.n3738 240.244
R6123 gnd.n4582 gnd.n3733 240.244
R6124 gnd.n4601 gnd.n3733 240.244
R6125 gnd.n4601 gnd.n3726 240.244
R6126 gnd.n4587 gnd.n3726 240.244
R6127 gnd.n4587 gnd.n3718 240.244
R6128 gnd.n4590 gnd.n3718 240.244
R6129 gnd.n4590 gnd.n3700 240.244
R6130 gnd.n3700 gnd.n3691 240.244
R6131 gnd.n4666 gnd.n3691 240.244
R6132 gnd.n4666 gnd.n3686 240.244
R6133 gnd.n4698 gnd.n3686 240.244
R6134 gnd.n4698 gnd.n3680 240.244
R6135 gnd.n4671 gnd.n3680 240.244
R6136 gnd.n4671 gnd.n3671 240.244
R6137 gnd.n4672 gnd.n3671 240.244
R6138 gnd.n4675 gnd.n4672 240.244
R6139 gnd.n4676 gnd.n4675 240.244
R6140 gnd.n4677 gnd.n4676 240.244
R6141 gnd.n4677 gnd.n3650 240.244
R6142 gnd.n3650 gnd.n3641 240.244
R6143 gnd.n4680 gnd.n3641 240.244
R6144 gnd.n4680 gnd.n3627 240.244
R6145 gnd.n4817 gnd.n3627 240.244
R6146 gnd.n4817 gnd.n3620 240.244
R6147 gnd.n4789 gnd.n3620 240.244
R6148 gnd.n4789 gnd.n3612 240.244
R6149 gnd.n4790 gnd.n3612 240.244
R6150 gnd.n4790 gnd.n3601 240.244
R6151 gnd.n4793 gnd.n3601 240.244
R6152 gnd.n4793 gnd.n3593 240.244
R6153 gnd.n4795 gnd.n3593 240.244
R6154 gnd.n4795 gnd.n3584 240.244
R6155 gnd.n4798 gnd.n3584 240.244
R6156 gnd.n4798 gnd.n3575 240.244
R6157 gnd.n3575 gnd.n3562 240.244
R6158 gnd.n4929 gnd.n3562 240.244
R6159 gnd.n4929 gnd.n3555 240.244
R6160 gnd.n4914 gnd.n3555 240.244
R6161 gnd.n4914 gnd.n3546 240.244
R6162 gnd.n4915 gnd.n3546 240.244
R6163 gnd.n4916 gnd.n4915 240.244
R6164 gnd.n4916 gnd.n3524 240.244
R6165 gnd.n3524 gnd.n3515 240.244
R6166 gnd.n5178 gnd.n3515 240.244
R6167 gnd.n5178 gnd.n3511 240.244
R6168 gnd.n5184 gnd.n3511 240.244
R6169 gnd.n5184 gnd.n3505 240.244
R6170 gnd.n5196 gnd.n3505 240.244
R6171 gnd.n5196 gnd.n3501 240.244
R6172 gnd.n5202 gnd.n3501 240.244
R6173 gnd.n5202 gnd.n3493 240.244
R6174 gnd.n5213 gnd.n3493 240.244
R6175 gnd.n5213 gnd.n3489 240.244
R6176 gnd.n5219 gnd.n3489 240.244
R6177 gnd.n5219 gnd.n3481 240.244
R6178 gnd.n5230 gnd.n3481 240.244
R6179 gnd.n5230 gnd.n3477 240.244
R6180 gnd.n5236 gnd.n3477 240.244
R6181 gnd.n5236 gnd.n3468 240.244
R6182 gnd.n5247 gnd.n3468 240.244
R6183 gnd.n5247 gnd.n3464 240.244
R6184 gnd.n5253 gnd.n3464 240.244
R6185 gnd.n5253 gnd.n3457 240.244
R6186 gnd.n5267 gnd.n3457 240.244
R6187 gnd.n5267 gnd.n3453 240.244
R6188 gnd.n5273 gnd.n3453 240.244
R6189 gnd.n5273 gnd.n3091 240.244
R6190 gnd.n5716 gnd.n3091 240.244
R6191 gnd.n2665 gnd.n2664 240.244
R6192 gnd.n2670 gnd.n2664 240.244
R6193 gnd.n2672 gnd.n2671 240.244
R6194 gnd.n2676 gnd.n2675 240.244
R6195 gnd.n2678 gnd.n2677 240.244
R6196 gnd.n2688 gnd.n2687 240.244
R6197 gnd.n2690 gnd.n2689 240.244
R6198 gnd.n2698 gnd.n2697 240.244
R6199 gnd.n2706 gnd.n2705 240.244
R6200 gnd.n2708 gnd.n2707 240.244
R6201 gnd.n2716 gnd.n2715 240.244
R6202 gnd.n2724 gnd.n2723 240.244
R6203 gnd.n2729 gnd.n2725 240.244
R6204 gnd.n2661 gnd.n2647 240.244
R6205 gnd.n4398 gnd.n2648 240.244
R6206 gnd.n4398 gnd.n3925 240.244
R6207 gnd.n4404 gnd.n3925 240.244
R6208 gnd.n4404 gnd.n3914 240.244
R6209 gnd.n4414 gnd.n3914 240.244
R6210 gnd.n4414 gnd.n3910 240.244
R6211 gnd.n4420 gnd.n3910 240.244
R6212 gnd.n4420 gnd.n3901 240.244
R6213 gnd.n4430 gnd.n3901 240.244
R6214 gnd.n4430 gnd.n3897 240.244
R6215 gnd.n4436 gnd.n3897 240.244
R6216 gnd.n4436 gnd.n3887 240.244
R6217 gnd.n4446 gnd.n3887 240.244
R6218 gnd.n4446 gnd.n3883 240.244
R6219 gnd.n4452 gnd.n3883 240.244
R6220 gnd.n4452 gnd.n3873 240.244
R6221 gnd.n4462 gnd.n3873 240.244
R6222 gnd.n4462 gnd.n3867 240.244
R6223 gnd.n4479 gnd.n3867 240.244
R6224 gnd.n4479 gnd.n3868 240.244
R6225 gnd.n3868 gnd.n3857 240.244
R6226 gnd.n4467 gnd.n3857 240.244
R6227 gnd.n4468 gnd.n4467 240.244
R6228 gnd.n4468 gnd.n2978 240.244
R6229 gnd.n2990 gnd.n2978 240.244
R6230 gnd.n5833 gnd.n2990 240.244
R6231 gnd.n5833 gnd.n2991 240.244
R6232 gnd.n2996 gnd.n2991 240.244
R6233 gnd.n2997 gnd.n2996 240.244
R6234 gnd.n2998 gnd.n2997 240.244
R6235 gnd.n4570 gnd.n2998 240.244
R6236 gnd.n4570 gnd.n3001 240.244
R6237 gnd.n3002 gnd.n3001 240.244
R6238 gnd.n3003 gnd.n3002 240.244
R6239 gnd.n4602 gnd.n3003 240.244
R6240 gnd.n4602 gnd.n3006 240.244
R6241 gnd.n3007 gnd.n3006 240.244
R6242 gnd.n3008 gnd.n3007 240.244
R6243 gnd.n4588 gnd.n3008 240.244
R6244 gnd.n4588 gnd.n3011 240.244
R6245 gnd.n3012 gnd.n3011 240.244
R6246 gnd.n3013 gnd.n3012 240.244
R6247 gnd.n4640 gnd.n3013 240.244
R6248 gnd.n4640 gnd.n3016 240.244
R6249 gnd.n3017 gnd.n3016 240.244
R6250 gnd.n3018 gnd.n3017 240.244
R6251 gnd.n3672 gnd.n3018 240.244
R6252 gnd.n3672 gnd.n3021 240.244
R6253 gnd.n3022 gnd.n3021 240.244
R6254 gnd.n3023 gnd.n3022 240.244
R6255 gnd.n3654 gnd.n3023 240.244
R6256 gnd.n3654 gnd.n3026 240.244
R6257 gnd.n3027 gnd.n3026 240.244
R6258 gnd.n3028 gnd.n3027 240.244
R6259 gnd.n3635 gnd.n3028 240.244
R6260 gnd.n3635 gnd.n3031 240.244
R6261 gnd.n3032 gnd.n3031 240.244
R6262 gnd.n3033 gnd.n3032 240.244
R6263 gnd.n3613 gnd.n3033 240.244
R6264 gnd.n3613 gnd.n3036 240.244
R6265 gnd.n3037 gnd.n3036 240.244
R6266 gnd.n3038 gnd.n3037 240.244
R6267 gnd.n3595 gnd.n3038 240.244
R6268 gnd.n3595 gnd.n3041 240.244
R6269 gnd.n3042 gnd.n3041 240.244
R6270 gnd.n3043 gnd.n3042 240.244
R6271 gnd.n3576 gnd.n3043 240.244
R6272 gnd.n3576 gnd.n3046 240.244
R6273 gnd.n3047 gnd.n3046 240.244
R6274 gnd.n3048 gnd.n3047 240.244
R6275 gnd.n4912 gnd.n3048 240.244
R6276 gnd.n4912 gnd.n3051 240.244
R6277 gnd.n3052 gnd.n3051 240.244
R6278 gnd.n3053 gnd.n3052 240.244
R6279 gnd.n5168 gnd.n3053 240.244
R6280 gnd.n5168 gnd.n3056 240.244
R6281 gnd.n3057 gnd.n3056 240.244
R6282 gnd.n3058 gnd.n3057 240.244
R6283 gnd.n5186 gnd.n3058 240.244
R6284 gnd.n5186 gnd.n3061 240.244
R6285 gnd.n3062 gnd.n3061 240.244
R6286 gnd.n3063 gnd.n3062 240.244
R6287 gnd.n5203 gnd.n3063 240.244
R6288 gnd.n5203 gnd.n3066 240.244
R6289 gnd.n3067 gnd.n3066 240.244
R6290 gnd.n3068 gnd.n3067 240.244
R6291 gnd.n5220 gnd.n3068 240.244
R6292 gnd.n5220 gnd.n3071 240.244
R6293 gnd.n3072 gnd.n3071 240.244
R6294 gnd.n3073 gnd.n3072 240.244
R6295 gnd.n5237 gnd.n3073 240.244
R6296 gnd.n5237 gnd.n3076 240.244
R6297 gnd.n3077 gnd.n3076 240.244
R6298 gnd.n3078 gnd.n3077 240.244
R6299 gnd.n5254 gnd.n3078 240.244
R6300 gnd.n5254 gnd.n3081 240.244
R6301 gnd.n3082 gnd.n3081 240.244
R6302 gnd.n3083 gnd.n3082 240.244
R6303 gnd.n5274 gnd.n3083 240.244
R6304 gnd.n5274 gnd.n3086 240.244
R6305 gnd.n5718 gnd.n3086 240.244
R6306 gnd.n3097 gnd.n3096 240.244
R6307 gnd.n3424 gnd.n3100 240.244
R6308 gnd.n3102 gnd.n3101 240.244
R6309 gnd.n3427 gnd.n3106 240.244
R6310 gnd.n3430 gnd.n3107 240.244
R6311 gnd.n3116 gnd.n3115 240.244
R6312 gnd.n3432 gnd.n3123 240.244
R6313 gnd.n3435 gnd.n3124 240.244
R6314 gnd.n3132 gnd.n3131 240.244
R6315 gnd.n3437 gnd.n3139 240.244
R6316 gnd.n3440 gnd.n3140 240.244
R6317 gnd.n3148 gnd.n3147 240.244
R6318 gnd.n3443 gnd.n3148 240.244
R6319 gnd.n5299 gnd.n3422 240.244
R6320 gnd.n2958 gnd.n2957 240.132
R6321 gnd.n4981 gnd.n4980 240.132
R6322 gnd.n6544 gnd.n805 225.874
R6323 gnd.n6552 gnd.n805 225.874
R6324 gnd.n6553 gnd.n6552 225.874
R6325 gnd.n6554 gnd.n6553 225.874
R6326 gnd.n6554 gnd.n799 225.874
R6327 gnd.n6562 gnd.n799 225.874
R6328 gnd.n6563 gnd.n6562 225.874
R6329 gnd.n6564 gnd.n6563 225.874
R6330 gnd.n6564 gnd.n793 225.874
R6331 gnd.n6572 gnd.n793 225.874
R6332 gnd.n6573 gnd.n6572 225.874
R6333 gnd.n6574 gnd.n6573 225.874
R6334 gnd.n6574 gnd.n787 225.874
R6335 gnd.n6582 gnd.n787 225.874
R6336 gnd.n6583 gnd.n6582 225.874
R6337 gnd.n6584 gnd.n6583 225.874
R6338 gnd.n6584 gnd.n781 225.874
R6339 gnd.n6592 gnd.n781 225.874
R6340 gnd.n6593 gnd.n6592 225.874
R6341 gnd.n6594 gnd.n6593 225.874
R6342 gnd.n6594 gnd.n775 225.874
R6343 gnd.n6602 gnd.n775 225.874
R6344 gnd.n6603 gnd.n6602 225.874
R6345 gnd.n6604 gnd.n6603 225.874
R6346 gnd.n6604 gnd.n769 225.874
R6347 gnd.n6612 gnd.n769 225.874
R6348 gnd.n6613 gnd.n6612 225.874
R6349 gnd.n6614 gnd.n6613 225.874
R6350 gnd.n6614 gnd.n763 225.874
R6351 gnd.n6622 gnd.n763 225.874
R6352 gnd.n6623 gnd.n6622 225.874
R6353 gnd.n6624 gnd.n6623 225.874
R6354 gnd.n6624 gnd.n757 225.874
R6355 gnd.n6632 gnd.n757 225.874
R6356 gnd.n6633 gnd.n6632 225.874
R6357 gnd.n6634 gnd.n6633 225.874
R6358 gnd.n6634 gnd.n751 225.874
R6359 gnd.n6642 gnd.n751 225.874
R6360 gnd.n6643 gnd.n6642 225.874
R6361 gnd.n6644 gnd.n6643 225.874
R6362 gnd.n6644 gnd.n745 225.874
R6363 gnd.n6652 gnd.n745 225.874
R6364 gnd.n6653 gnd.n6652 225.874
R6365 gnd.n6654 gnd.n6653 225.874
R6366 gnd.n6654 gnd.n739 225.874
R6367 gnd.n6662 gnd.n739 225.874
R6368 gnd.n6663 gnd.n6662 225.874
R6369 gnd.n6664 gnd.n6663 225.874
R6370 gnd.n6664 gnd.n733 225.874
R6371 gnd.n6672 gnd.n733 225.874
R6372 gnd.n6673 gnd.n6672 225.874
R6373 gnd.n6674 gnd.n6673 225.874
R6374 gnd.n6674 gnd.n727 225.874
R6375 gnd.n6682 gnd.n727 225.874
R6376 gnd.n6683 gnd.n6682 225.874
R6377 gnd.n6684 gnd.n6683 225.874
R6378 gnd.n6684 gnd.n721 225.874
R6379 gnd.n6692 gnd.n721 225.874
R6380 gnd.n6693 gnd.n6692 225.874
R6381 gnd.n6694 gnd.n6693 225.874
R6382 gnd.n6694 gnd.n715 225.874
R6383 gnd.n6702 gnd.n715 225.874
R6384 gnd.n6703 gnd.n6702 225.874
R6385 gnd.n6704 gnd.n6703 225.874
R6386 gnd.n6704 gnd.n709 225.874
R6387 gnd.n6712 gnd.n709 225.874
R6388 gnd.n6713 gnd.n6712 225.874
R6389 gnd.n6714 gnd.n6713 225.874
R6390 gnd.n6714 gnd.n703 225.874
R6391 gnd.n6722 gnd.n703 225.874
R6392 gnd.n6723 gnd.n6722 225.874
R6393 gnd.n6724 gnd.n6723 225.874
R6394 gnd.n6724 gnd.n697 225.874
R6395 gnd.n6732 gnd.n697 225.874
R6396 gnd.n6733 gnd.n6732 225.874
R6397 gnd.n6734 gnd.n6733 225.874
R6398 gnd.n6734 gnd.n691 225.874
R6399 gnd.n6742 gnd.n691 225.874
R6400 gnd.n6743 gnd.n6742 225.874
R6401 gnd.n6744 gnd.n6743 225.874
R6402 gnd.n6744 gnd.n685 225.874
R6403 gnd.n6752 gnd.n685 225.874
R6404 gnd.n6753 gnd.n6752 225.874
R6405 gnd.n6754 gnd.n6753 225.874
R6406 gnd.n6754 gnd.n679 225.874
R6407 gnd.n6762 gnd.n679 225.874
R6408 gnd.n6763 gnd.n6762 225.874
R6409 gnd.n6764 gnd.n6763 225.874
R6410 gnd.n6764 gnd.n673 225.874
R6411 gnd.n6772 gnd.n673 225.874
R6412 gnd.n6773 gnd.n6772 225.874
R6413 gnd.n6774 gnd.n6773 225.874
R6414 gnd.n6774 gnd.n667 225.874
R6415 gnd.n6782 gnd.n667 225.874
R6416 gnd.n6783 gnd.n6782 225.874
R6417 gnd.n6784 gnd.n6783 225.874
R6418 gnd.n6784 gnd.n661 225.874
R6419 gnd.n6792 gnd.n661 225.874
R6420 gnd.n6793 gnd.n6792 225.874
R6421 gnd.n6794 gnd.n6793 225.874
R6422 gnd.n6794 gnd.n655 225.874
R6423 gnd.n6802 gnd.n655 225.874
R6424 gnd.n6803 gnd.n6802 225.874
R6425 gnd.n6804 gnd.n6803 225.874
R6426 gnd.n6804 gnd.n649 225.874
R6427 gnd.n6812 gnd.n649 225.874
R6428 gnd.n6813 gnd.n6812 225.874
R6429 gnd.n6814 gnd.n6813 225.874
R6430 gnd.n6814 gnd.n643 225.874
R6431 gnd.n6822 gnd.n643 225.874
R6432 gnd.n6823 gnd.n6822 225.874
R6433 gnd.n6824 gnd.n6823 225.874
R6434 gnd.n6824 gnd.n637 225.874
R6435 gnd.n6832 gnd.n637 225.874
R6436 gnd.n6833 gnd.n6832 225.874
R6437 gnd.n6834 gnd.n6833 225.874
R6438 gnd.n6834 gnd.n631 225.874
R6439 gnd.n6842 gnd.n631 225.874
R6440 gnd.n6843 gnd.n6842 225.874
R6441 gnd.n6844 gnd.n6843 225.874
R6442 gnd.n6844 gnd.n625 225.874
R6443 gnd.n6852 gnd.n625 225.874
R6444 gnd.n6853 gnd.n6852 225.874
R6445 gnd.n6854 gnd.n6853 225.874
R6446 gnd.n6854 gnd.n619 225.874
R6447 gnd.n6862 gnd.n619 225.874
R6448 gnd.n6863 gnd.n6862 225.874
R6449 gnd.n6864 gnd.n6863 225.874
R6450 gnd.n6864 gnd.n613 225.874
R6451 gnd.n6872 gnd.n613 225.874
R6452 gnd.n6873 gnd.n6872 225.874
R6453 gnd.n6874 gnd.n6873 225.874
R6454 gnd.n6874 gnd.n607 225.874
R6455 gnd.n6882 gnd.n607 225.874
R6456 gnd.n6883 gnd.n6882 225.874
R6457 gnd.n6884 gnd.n6883 225.874
R6458 gnd.n6884 gnd.n601 225.874
R6459 gnd.n6892 gnd.n601 225.874
R6460 gnd.n6893 gnd.n6892 225.874
R6461 gnd.n6894 gnd.n6893 225.874
R6462 gnd.n6894 gnd.n595 225.874
R6463 gnd.n6902 gnd.n595 225.874
R6464 gnd.n6903 gnd.n6902 225.874
R6465 gnd.n6904 gnd.n6903 225.874
R6466 gnd.n6904 gnd.n589 225.874
R6467 gnd.n6912 gnd.n589 225.874
R6468 gnd.n6913 gnd.n6912 225.874
R6469 gnd.n6914 gnd.n6913 225.874
R6470 gnd.n6914 gnd.n583 225.874
R6471 gnd.n6922 gnd.n583 225.874
R6472 gnd.n6923 gnd.n6922 225.874
R6473 gnd.n6924 gnd.n6923 225.874
R6474 gnd.n6924 gnd.n577 225.874
R6475 gnd.n6932 gnd.n577 225.874
R6476 gnd.n6933 gnd.n6932 225.874
R6477 gnd.n6934 gnd.n6933 225.874
R6478 gnd.n6934 gnd.n571 225.874
R6479 gnd.n6942 gnd.n571 225.874
R6480 gnd.n6943 gnd.n6942 225.874
R6481 gnd.n6944 gnd.n6943 225.874
R6482 gnd.n6944 gnd.n565 225.874
R6483 gnd.n6952 gnd.n565 225.874
R6484 gnd.n6953 gnd.n6952 225.874
R6485 gnd.n6954 gnd.n6953 225.874
R6486 gnd.n6954 gnd.n559 225.874
R6487 gnd.n6962 gnd.n559 225.874
R6488 gnd.n6963 gnd.n6962 225.874
R6489 gnd.n6964 gnd.n6963 225.874
R6490 gnd.n6964 gnd.n553 225.874
R6491 gnd.n6972 gnd.n553 225.874
R6492 gnd.n6973 gnd.n6972 225.874
R6493 gnd.n6974 gnd.n6973 225.874
R6494 gnd.n6974 gnd.n547 225.874
R6495 gnd.n6982 gnd.n547 225.874
R6496 gnd.n6983 gnd.n6982 225.874
R6497 gnd.n6984 gnd.n6983 225.874
R6498 gnd.n6984 gnd.n541 225.874
R6499 gnd.n6993 gnd.n541 225.874
R6500 gnd.n6994 gnd.n6993 225.874
R6501 gnd.n6995 gnd.n6994 225.874
R6502 gnd.n6995 gnd.n536 225.874
R6503 gnd.n1440 gnd.t139 224.174
R6504 gnd.n1072 gnd.t44 224.174
R6505 gnd.n3232 gnd.n3169 199.319
R6506 gnd.n3232 gnd.n3170 199.319
R6507 gnd.n2814 gnd.n2769 199.319
R6508 gnd.n2814 gnd.n2768 199.319
R6509 gnd.n2959 gnd.n2956 186.49
R6510 gnd.n4982 gnd.n4979 186.49
R6511 gnd.n2311 gnd.n2310 185
R6512 gnd.n2309 gnd.n2308 185
R6513 gnd.n2288 gnd.n2287 185
R6514 gnd.n2303 gnd.n2302 185
R6515 gnd.n2301 gnd.n2300 185
R6516 gnd.n2292 gnd.n2291 185
R6517 gnd.n2295 gnd.n2294 185
R6518 gnd.n2279 gnd.n2278 185
R6519 gnd.n2277 gnd.n2276 185
R6520 gnd.n2256 gnd.n2255 185
R6521 gnd.n2271 gnd.n2270 185
R6522 gnd.n2269 gnd.n2268 185
R6523 gnd.n2260 gnd.n2259 185
R6524 gnd.n2263 gnd.n2262 185
R6525 gnd.n2247 gnd.n2246 185
R6526 gnd.n2245 gnd.n2244 185
R6527 gnd.n2224 gnd.n2223 185
R6528 gnd.n2239 gnd.n2238 185
R6529 gnd.n2237 gnd.n2236 185
R6530 gnd.n2228 gnd.n2227 185
R6531 gnd.n2231 gnd.n2230 185
R6532 gnd.n2216 gnd.n2215 185
R6533 gnd.n2214 gnd.n2213 185
R6534 gnd.n2193 gnd.n2192 185
R6535 gnd.n2208 gnd.n2207 185
R6536 gnd.n2206 gnd.n2205 185
R6537 gnd.n2197 gnd.n2196 185
R6538 gnd.n2200 gnd.n2199 185
R6539 gnd.n2184 gnd.n2183 185
R6540 gnd.n2182 gnd.n2181 185
R6541 gnd.n2161 gnd.n2160 185
R6542 gnd.n2176 gnd.n2175 185
R6543 gnd.n2174 gnd.n2173 185
R6544 gnd.n2165 gnd.n2164 185
R6545 gnd.n2168 gnd.n2167 185
R6546 gnd.n2152 gnd.n2151 185
R6547 gnd.n2150 gnd.n2149 185
R6548 gnd.n2129 gnd.n2128 185
R6549 gnd.n2144 gnd.n2143 185
R6550 gnd.n2142 gnd.n2141 185
R6551 gnd.n2133 gnd.n2132 185
R6552 gnd.n2136 gnd.n2135 185
R6553 gnd.n2120 gnd.n2119 185
R6554 gnd.n2118 gnd.n2117 185
R6555 gnd.n2097 gnd.n2096 185
R6556 gnd.n2112 gnd.n2111 185
R6557 gnd.n2110 gnd.n2109 185
R6558 gnd.n2101 gnd.n2100 185
R6559 gnd.n2104 gnd.n2103 185
R6560 gnd.n2089 gnd.n2088 185
R6561 gnd.n2087 gnd.n2086 185
R6562 gnd.n2066 gnd.n2065 185
R6563 gnd.n2081 gnd.n2080 185
R6564 gnd.n2079 gnd.n2078 185
R6565 gnd.n2070 gnd.n2069 185
R6566 gnd.n2073 gnd.n2072 185
R6567 gnd.n7004 gnd.n7003 183.87
R6568 gnd.n7005 gnd.n7004 183.87
R6569 gnd.n7005 gnd.n530 183.87
R6570 gnd.n7013 gnd.n530 183.87
R6571 gnd.n7014 gnd.n7013 183.87
R6572 gnd.n7015 gnd.n7014 183.87
R6573 gnd.n7015 gnd.n524 183.87
R6574 gnd.n7023 gnd.n524 183.87
R6575 gnd.n7024 gnd.n7023 183.87
R6576 gnd.n7025 gnd.n7024 183.87
R6577 gnd.n7025 gnd.n518 183.87
R6578 gnd.n7033 gnd.n518 183.87
R6579 gnd.n7034 gnd.n7033 183.87
R6580 gnd.n7035 gnd.n7034 183.87
R6581 gnd.n7035 gnd.n512 183.87
R6582 gnd.n7043 gnd.n512 183.87
R6583 gnd.n7044 gnd.n7043 183.87
R6584 gnd.n7045 gnd.n7044 183.87
R6585 gnd.n7045 gnd.n506 183.87
R6586 gnd.n7053 gnd.n506 183.87
R6587 gnd.n7054 gnd.n7053 183.87
R6588 gnd.n7055 gnd.n7054 183.87
R6589 gnd.n7055 gnd.n500 183.87
R6590 gnd.n7063 gnd.n500 183.87
R6591 gnd.n7064 gnd.n7063 183.87
R6592 gnd.n7065 gnd.n7064 183.87
R6593 gnd.n7065 gnd.n494 183.87
R6594 gnd.n7073 gnd.n494 183.87
R6595 gnd.n7074 gnd.n7073 183.87
R6596 gnd.n7075 gnd.n7074 183.87
R6597 gnd.n7075 gnd.n488 183.87
R6598 gnd.n7083 gnd.n488 183.87
R6599 gnd.n7084 gnd.n7083 183.87
R6600 gnd.n7085 gnd.n7084 183.87
R6601 gnd.n7085 gnd.n482 183.87
R6602 gnd.n7093 gnd.n482 183.87
R6603 gnd.n7094 gnd.n7093 183.87
R6604 gnd.n7095 gnd.n7094 183.87
R6605 gnd.n7095 gnd.n476 183.87
R6606 gnd.n7103 gnd.n476 183.87
R6607 gnd.n7104 gnd.n7103 183.87
R6608 gnd.n7105 gnd.n7104 183.87
R6609 gnd.n7105 gnd.n470 183.87
R6610 gnd.n7113 gnd.n470 183.87
R6611 gnd.n7114 gnd.n7113 183.87
R6612 gnd.n7115 gnd.n7114 183.87
R6613 gnd.n7115 gnd.n464 183.87
R6614 gnd.n7123 gnd.n464 183.87
R6615 gnd.n7124 gnd.n7123 183.87
R6616 gnd.n7125 gnd.n7124 183.87
R6617 gnd.n7125 gnd.n458 183.87
R6618 gnd.n7133 gnd.n458 183.87
R6619 gnd.n7134 gnd.n7133 183.87
R6620 gnd.n7135 gnd.n7134 183.87
R6621 gnd.n7135 gnd.n452 183.87
R6622 gnd.n7143 gnd.n452 183.87
R6623 gnd.n7144 gnd.n7143 183.87
R6624 gnd.n7145 gnd.n7144 183.87
R6625 gnd.n7145 gnd.n446 183.87
R6626 gnd.n7153 gnd.n446 183.87
R6627 gnd.n7154 gnd.n7153 183.87
R6628 gnd.n7155 gnd.n7154 183.87
R6629 gnd.n7155 gnd.n440 183.87
R6630 gnd.n7163 gnd.n440 183.87
R6631 gnd.n7164 gnd.n7163 183.87
R6632 gnd.n7165 gnd.n7164 183.87
R6633 gnd.n7165 gnd.n434 183.87
R6634 gnd.n7173 gnd.n434 183.87
R6635 gnd.n7174 gnd.n7173 183.87
R6636 gnd.n7175 gnd.n7174 183.87
R6637 gnd.n7175 gnd.n428 183.87
R6638 gnd.n7183 gnd.n428 183.87
R6639 gnd.n7184 gnd.n7183 183.87
R6640 gnd.n7185 gnd.n7184 183.87
R6641 gnd.n7185 gnd.n422 183.87
R6642 gnd.n7193 gnd.n422 183.87
R6643 gnd.n7194 gnd.n7193 183.87
R6644 gnd.n7195 gnd.n7194 183.87
R6645 gnd.n7195 gnd.n416 183.87
R6646 gnd.n7203 gnd.n416 183.87
R6647 gnd.n7204 gnd.n7203 183.87
R6648 gnd.n7206 gnd.n7204 183.87
R6649 gnd.n7206 gnd.n7205 183.87
R6650 gnd.n1441 gnd.t138 178.987
R6651 gnd.n1073 gnd.t45 178.987
R6652 gnd.n5596 gnd.n3231 171.457
R6653 gnd.n5915 gnd.n5914 171.457
R6654 gnd.n1 gnd.t1 170.774
R6655 gnd.n9 gnd.t163 170.103
R6656 gnd.n8 gnd.t17 170.103
R6657 gnd.n7 gnd.t193 170.103
R6658 gnd.n6 gnd.t179 170.103
R6659 gnd.n5 gnd.t199 170.103
R6660 gnd.n4 gnd.t201 170.103
R6661 gnd.n3 gnd.t197 170.103
R6662 gnd.n2 gnd.t203 170.103
R6663 gnd.n1 gnd.t189 170.103
R6664 gnd.n5155 gnd.n5154 163.367
R6665 gnd.n5152 gnd.n4992 163.367
R6666 gnd.n5148 gnd.n5147 163.367
R6667 gnd.n5145 gnd.n4995 163.367
R6668 gnd.n5141 gnd.n5140 163.367
R6669 gnd.n5138 gnd.n4998 163.367
R6670 gnd.n5134 gnd.n5133 163.367
R6671 gnd.n5131 gnd.n5001 163.367
R6672 gnd.n5127 gnd.n5126 163.367
R6673 gnd.n5124 gnd.n5004 163.367
R6674 gnd.n5120 gnd.n5119 163.367
R6675 gnd.n5117 gnd.n5007 163.367
R6676 gnd.n5113 gnd.n5112 163.367
R6677 gnd.n5110 gnd.n5010 163.367
R6678 gnd.n5105 gnd.n5104 163.367
R6679 gnd.n5102 gnd.n5100 163.367
R6680 gnd.n5097 gnd.n5096 163.367
R6681 gnd.n5094 gnd.n5016 163.367
R6682 gnd.n5089 gnd.n5088 163.367
R6683 gnd.n5086 gnd.n5021 163.367
R6684 gnd.n5082 gnd.n5081 163.367
R6685 gnd.n5079 gnd.n5024 163.367
R6686 gnd.n5075 gnd.n5074 163.367
R6687 gnd.n5072 gnd.n5027 163.367
R6688 gnd.n5068 gnd.n5067 163.367
R6689 gnd.n5065 gnd.n5030 163.367
R6690 gnd.n5061 gnd.n5060 163.367
R6691 gnd.n5058 gnd.n5033 163.367
R6692 gnd.n5054 gnd.n5053 163.367
R6693 gnd.n5051 gnd.n5036 163.367
R6694 gnd.n5047 gnd.n5046 163.367
R6695 gnd.n5044 gnd.n5040 163.367
R6696 gnd.n3837 gnd.n2975 163.367
R6697 gnd.n3841 gnd.n2975 163.367
R6698 gnd.n3842 gnd.n3841 163.367
R6699 gnd.n3843 gnd.n3842 163.367
R6700 gnd.n3843 gnd.n3770 163.367
R6701 gnd.n3847 gnd.n3770 163.367
R6702 gnd.n3847 gnd.n3758 163.367
R6703 gnd.n4531 gnd.n3758 163.367
R6704 gnd.n4531 gnd.n3755 163.367
R6705 gnd.n4557 gnd.n3755 163.367
R6706 gnd.n4557 gnd.n3756 163.367
R6707 gnd.n3756 gnd.n3749 163.367
R6708 gnd.n4552 gnd.n3749 163.367
R6709 gnd.n4552 gnd.n4549 163.367
R6710 gnd.n4549 gnd.n4548 163.367
R6711 gnd.n4548 gnd.n4537 163.367
R6712 gnd.n4537 gnd.n3732 163.367
R6713 gnd.n4543 gnd.n3732 163.367
R6714 gnd.n4543 gnd.n3727 163.367
R6715 gnd.n4540 gnd.n3727 163.367
R6716 gnd.n4540 gnd.n3717 163.367
R6717 gnd.n3717 gnd.n3712 163.367
R6718 gnd.n4627 gnd.n3712 163.367
R6719 gnd.n4628 gnd.n4627 163.367
R6720 gnd.n4628 gnd.n3701 163.367
R6721 gnd.n3709 gnd.n3701 163.367
R6722 gnd.n4647 gnd.n3709 163.367
R6723 gnd.n4647 gnd.n3710 163.367
R6724 gnd.n4643 gnd.n3710 163.367
R6725 gnd.n4643 gnd.n3685 163.367
R6726 gnd.n4637 gnd.n3685 163.367
R6727 gnd.n4637 gnd.n3681 163.367
R6728 gnd.n4634 gnd.n3681 163.367
R6729 gnd.n4634 gnd.n3670 163.367
R6730 gnd.n3670 gnd.n3662 163.367
R6731 gnd.n4734 gnd.n3662 163.367
R6732 gnd.n4734 gnd.n3660 163.367
R6733 gnd.n4739 gnd.n3660 163.367
R6734 gnd.n4739 gnd.n3652 163.367
R6735 gnd.n4748 gnd.n3652 163.367
R6736 gnd.n4749 gnd.n4748 163.367
R6737 gnd.n4749 gnd.n3649 163.367
R6738 gnd.n4756 gnd.n3649 163.367
R6739 gnd.n4756 gnd.n3642 163.367
R6740 gnd.n4752 gnd.n3642 163.367
R6741 gnd.n4752 gnd.n3633 163.367
R6742 gnd.n4779 gnd.n3633 163.367
R6743 gnd.n4779 gnd.n3626 163.367
R6744 gnd.n4782 gnd.n3626 163.367
R6745 gnd.n4782 gnd.n3621 163.367
R6746 gnd.n4786 gnd.n3621 163.367
R6747 gnd.n4786 gnd.n3610 163.367
R6748 gnd.n4839 gnd.n3610 163.367
R6749 gnd.n4839 gnd.n3608 163.367
R6750 gnd.n4848 gnd.n3608 163.367
R6751 gnd.n4848 gnd.n3602 163.367
R6752 gnd.n4844 gnd.n3602 163.367
R6753 gnd.n4844 gnd.n3592 163.367
R6754 gnd.n3592 gnd.n3587 163.367
R6755 gnd.n4874 gnd.n3587 163.367
R6756 gnd.n4874 gnd.n3585 163.367
R6757 gnd.n4880 gnd.n3585 163.367
R6758 gnd.n4880 gnd.n3574 163.367
R6759 gnd.n3574 gnd.n3568 163.367
R6760 gnd.n4901 gnd.n3568 163.367
R6761 gnd.n4902 gnd.n4901 163.367
R6762 gnd.n4902 gnd.n3561 163.367
R6763 gnd.n4905 gnd.n3561 163.367
R6764 gnd.n4905 gnd.n3556 163.367
R6765 gnd.n4910 gnd.n3556 163.367
R6766 gnd.n4910 gnd.n3545 163.367
R6767 gnd.n3545 gnd.n3539 163.367
R6768 gnd.n4957 gnd.n3539 163.367
R6769 gnd.n4957 gnd.n3537 163.367
R6770 gnd.n4961 gnd.n3537 163.367
R6771 gnd.n4961 gnd.n3527 163.367
R6772 gnd.n5167 gnd.n3527 163.367
R6773 gnd.n5167 gnd.n3528 163.367
R6774 gnd.n5163 gnd.n3528 163.367
R6775 gnd.n5163 gnd.n5162 163.367
R6776 gnd.n2950 gnd.n2949 163.367
R6777 gnd.n5904 gnd.n2949 163.367
R6778 gnd.n5902 gnd.n5901 163.367
R6779 gnd.n5898 gnd.n5897 163.367
R6780 gnd.n5894 gnd.n5893 163.367
R6781 gnd.n5890 gnd.n5889 163.367
R6782 gnd.n5886 gnd.n5885 163.367
R6783 gnd.n5882 gnd.n5881 163.367
R6784 gnd.n5878 gnd.n5877 163.367
R6785 gnd.n5874 gnd.n5873 163.367
R6786 gnd.n5870 gnd.n5869 163.367
R6787 gnd.n5866 gnd.n5865 163.367
R6788 gnd.n5862 gnd.n5861 163.367
R6789 gnd.n5858 gnd.n5857 163.367
R6790 gnd.n5854 gnd.n5853 163.367
R6791 gnd.n5850 gnd.n5849 163.367
R6792 gnd.n5913 gnd.n2915 163.367
R6793 gnd.n3776 gnd.n3775 163.367
R6794 gnd.n3781 gnd.n3780 163.367
R6795 gnd.n3785 gnd.n3784 163.367
R6796 gnd.n3789 gnd.n3788 163.367
R6797 gnd.n3793 gnd.n3792 163.367
R6798 gnd.n3797 gnd.n3796 163.367
R6799 gnd.n3801 gnd.n3800 163.367
R6800 gnd.n3805 gnd.n3804 163.367
R6801 gnd.n3809 gnd.n3808 163.367
R6802 gnd.n3813 gnd.n3812 163.367
R6803 gnd.n3817 gnd.n3816 163.367
R6804 gnd.n3821 gnd.n3820 163.367
R6805 gnd.n3825 gnd.n3824 163.367
R6806 gnd.n3829 gnd.n3828 163.367
R6807 gnd.n3833 gnd.n3832 163.367
R6808 gnd.n5842 gnd.n2951 163.367
R6809 gnd.n5842 gnd.n2973 163.367
R6810 gnd.n3763 gnd.n2973 163.367
R6811 gnd.n3766 gnd.n3763 163.367
R6812 gnd.n3767 gnd.n3766 163.367
R6813 gnd.n4525 gnd.n3767 163.367
R6814 gnd.n4525 gnd.n3761 163.367
R6815 gnd.n4529 gnd.n3761 163.367
R6816 gnd.n4529 gnd.n3753 163.367
R6817 gnd.n4559 gnd.n3753 163.367
R6818 gnd.n4559 gnd.n3750 163.367
R6819 gnd.n4568 gnd.n3750 163.367
R6820 gnd.n4568 gnd.n3751 163.367
R6821 gnd.n4564 gnd.n3751 163.367
R6822 gnd.n4564 gnd.n4563 163.367
R6823 gnd.n4563 gnd.n3731 163.367
R6824 gnd.n4605 gnd.n3731 163.367
R6825 gnd.n4605 gnd.n3729 163.367
R6826 gnd.n4609 gnd.n3729 163.367
R6827 gnd.n4609 gnd.n3715 163.367
R6828 gnd.n4621 gnd.n3715 163.367
R6829 gnd.n4621 gnd.n3713 163.367
R6830 gnd.n4625 gnd.n3713 163.367
R6831 gnd.n4625 gnd.n3703 163.367
R6832 gnd.n4653 gnd.n3703 163.367
R6833 gnd.n4653 gnd.n3704 163.367
R6834 gnd.n4649 gnd.n3704 163.367
R6835 gnd.n4649 gnd.n3707 163.367
R6836 gnd.n3707 gnd.n3684 163.367
R6837 gnd.n4701 gnd.n3684 163.367
R6838 gnd.n4701 gnd.n3682 163.367
R6839 gnd.n4705 gnd.n3682 163.367
R6840 gnd.n4705 gnd.n3668 163.367
R6841 gnd.n4728 gnd.n3668 163.367
R6842 gnd.n4728 gnd.n3666 163.367
R6843 gnd.n4732 gnd.n3666 163.367
R6844 gnd.n4732 gnd.n3658 163.367
R6845 gnd.n4742 gnd.n3658 163.367
R6846 gnd.n4742 gnd.n3656 163.367
R6847 gnd.n4746 gnd.n3656 163.367
R6848 gnd.n4746 gnd.n3647 163.367
R6849 gnd.n4760 gnd.n3647 163.367
R6850 gnd.n4760 gnd.n3644 163.367
R6851 gnd.n4767 gnd.n3644 163.367
R6852 gnd.n4767 gnd.n3645 163.367
R6853 gnd.n4763 gnd.n3645 163.367
R6854 gnd.n4763 gnd.n3625 163.367
R6855 gnd.n4820 gnd.n3625 163.367
R6856 gnd.n4820 gnd.n3622 163.367
R6857 gnd.n4827 gnd.n3622 163.367
R6858 gnd.n4827 gnd.n3623 163.367
R6859 gnd.n4823 gnd.n3623 163.367
R6860 gnd.n4823 gnd.n3606 163.367
R6861 gnd.n4851 gnd.n3606 163.367
R6862 gnd.n4851 gnd.n3604 163.367
R6863 gnd.n4855 gnd.n3604 163.367
R6864 gnd.n4855 gnd.n3591 163.367
R6865 gnd.n4867 gnd.n3591 163.367
R6866 gnd.n4867 gnd.n3588 163.367
R6867 gnd.n4872 gnd.n3588 163.367
R6868 gnd.n4872 gnd.n3589 163.367
R6869 gnd.n3589 gnd.n3572 163.367
R6870 gnd.n4895 gnd.n3572 163.367
R6871 gnd.n4895 gnd.n3570 163.367
R6872 gnd.n4899 gnd.n3570 163.367
R6873 gnd.n4899 gnd.n3559 163.367
R6874 gnd.n4932 gnd.n3559 163.367
R6875 gnd.n4932 gnd.n3557 163.367
R6876 gnd.n4936 gnd.n3557 163.367
R6877 gnd.n4936 gnd.n3544 163.367
R6878 gnd.n4950 gnd.n3544 163.367
R6879 gnd.n4950 gnd.n3542 163.367
R6880 gnd.n4955 gnd.n3542 163.367
R6881 gnd.n4955 gnd.n3536 163.367
R6882 gnd.n4963 gnd.n3536 163.367
R6883 gnd.n4964 gnd.n4963 163.367
R6884 gnd.n4964 gnd.n3525 163.367
R6885 gnd.n4967 gnd.n3525 163.367
R6886 gnd.n4967 gnd.n3533 163.367
R6887 gnd.n5160 gnd.n3533 163.367
R6888 gnd.n7205 gnd.n171 160.351
R6889 gnd.n4988 gnd.n4987 156.462
R6890 gnd.n2251 gnd.n2219 153.042
R6891 gnd.n2315 gnd.n2314 152.079
R6892 gnd.n2283 gnd.n2282 152.079
R6893 gnd.n2251 gnd.n2250 152.079
R6894 gnd.n2964 gnd.n2963 152
R6895 gnd.n2965 gnd.n2954 152
R6896 gnd.n2967 gnd.n2966 152
R6897 gnd.n2969 gnd.n2952 152
R6898 gnd.n2971 gnd.n2970 152
R6899 gnd.n4986 gnd.n4970 152
R6900 gnd.n4978 gnd.n4971 152
R6901 gnd.n4977 gnd.n4976 152
R6902 gnd.n4975 gnd.n4972 152
R6903 gnd.n4973 gnd.t69 150.546
R6904 gnd.t171 gnd.n2293 147.661
R6905 gnd.t32 gnd.n2261 147.661
R6906 gnd.t181 gnd.n2229 147.661
R6907 gnd.t161 gnd.n2198 147.661
R6908 gnd.t208 gnd.n2166 147.661
R6909 gnd.t334 gnd.n2134 147.661
R6910 gnd.t195 gnd.n2102 147.661
R6911 gnd.t165 gnd.n2071 147.661
R6912 gnd.n5099 gnd.n5098 143.351
R6913 gnd.n2931 gnd.n2914 143.351
R6914 gnd.n5912 gnd.n2914 143.351
R6915 gnd.n2961 gnd.t126 130.484
R6916 gnd.n2970 gnd.t46 126.766
R6917 gnd.n2968 gnd.t120 126.766
R6918 gnd.n2954 gnd.t146 126.766
R6919 gnd.n2962 gnd.t76 126.766
R6920 gnd.n4974 gnd.t143 126.766
R6921 gnd.n4976 gnd.t96 126.766
R6922 gnd.n4985 gnd.t39 126.766
R6923 gnd.n4987 gnd.t111 126.766
R6924 gnd.n2310 gnd.n2309 104.615
R6925 gnd.n2309 gnd.n2287 104.615
R6926 gnd.n2302 gnd.n2287 104.615
R6927 gnd.n2302 gnd.n2301 104.615
R6928 gnd.n2301 gnd.n2291 104.615
R6929 gnd.n2294 gnd.n2291 104.615
R6930 gnd.n2278 gnd.n2277 104.615
R6931 gnd.n2277 gnd.n2255 104.615
R6932 gnd.n2270 gnd.n2255 104.615
R6933 gnd.n2270 gnd.n2269 104.615
R6934 gnd.n2269 gnd.n2259 104.615
R6935 gnd.n2262 gnd.n2259 104.615
R6936 gnd.n2246 gnd.n2245 104.615
R6937 gnd.n2245 gnd.n2223 104.615
R6938 gnd.n2238 gnd.n2223 104.615
R6939 gnd.n2238 gnd.n2237 104.615
R6940 gnd.n2237 gnd.n2227 104.615
R6941 gnd.n2230 gnd.n2227 104.615
R6942 gnd.n2215 gnd.n2214 104.615
R6943 gnd.n2214 gnd.n2192 104.615
R6944 gnd.n2207 gnd.n2192 104.615
R6945 gnd.n2207 gnd.n2206 104.615
R6946 gnd.n2206 gnd.n2196 104.615
R6947 gnd.n2199 gnd.n2196 104.615
R6948 gnd.n2183 gnd.n2182 104.615
R6949 gnd.n2182 gnd.n2160 104.615
R6950 gnd.n2175 gnd.n2160 104.615
R6951 gnd.n2175 gnd.n2174 104.615
R6952 gnd.n2174 gnd.n2164 104.615
R6953 gnd.n2167 gnd.n2164 104.615
R6954 gnd.n2151 gnd.n2150 104.615
R6955 gnd.n2150 gnd.n2128 104.615
R6956 gnd.n2143 gnd.n2128 104.615
R6957 gnd.n2143 gnd.n2142 104.615
R6958 gnd.n2142 gnd.n2132 104.615
R6959 gnd.n2135 gnd.n2132 104.615
R6960 gnd.n2119 gnd.n2118 104.615
R6961 gnd.n2118 gnd.n2096 104.615
R6962 gnd.n2111 gnd.n2096 104.615
R6963 gnd.n2111 gnd.n2110 104.615
R6964 gnd.n2110 gnd.n2100 104.615
R6965 gnd.n2103 gnd.n2100 104.615
R6966 gnd.n2088 gnd.n2087 104.615
R6967 gnd.n2087 gnd.n2065 104.615
R6968 gnd.n2080 gnd.n2065 104.615
R6969 gnd.n2080 gnd.n2079 104.615
R6970 gnd.n2079 gnd.n2069 104.615
R6971 gnd.n2072 gnd.n2069 104.615
R6972 gnd.n1703 gnd.t89 100.632
R6973 gnd.n1051 gnd.t134 100.632
R6974 gnd.n243 gnd.n241 99.6594
R6975 gnd.n249 gnd.n234 99.6594
R6976 gnd.n253 gnd.n251 99.6594
R6977 gnd.n259 gnd.n230 99.6594
R6978 gnd.n263 gnd.n261 99.6594
R6979 gnd.n269 gnd.n226 99.6594
R6980 gnd.n274 gnd.n271 99.6594
R6981 gnd.n272 gnd.n222 99.6594
R6982 gnd.n284 gnd.n282 99.6594
R6983 gnd.n290 gnd.n216 99.6594
R6984 gnd.n294 gnd.n292 99.6594
R6985 gnd.n300 gnd.n212 99.6594
R6986 gnd.n304 gnd.n302 99.6594
R6987 gnd.n310 gnd.n208 99.6594
R6988 gnd.n314 gnd.n312 99.6594
R6989 gnd.n320 gnd.n204 99.6594
R6990 gnd.n324 gnd.n322 99.6594
R6991 gnd.n330 gnd.n200 99.6594
R6992 gnd.n334 gnd.n332 99.6594
R6993 gnd.n340 gnd.n194 99.6594
R6994 gnd.n344 gnd.n342 99.6594
R6995 gnd.n350 gnd.n190 99.6594
R6996 gnd.n354 gnd.n352 99.6594
R6997 gnd.n360 gnd.n186 99.6594
R6998 gnd.n364 gnd.n362 99.6594
R6999 gnd.n370 gnd.n182 99.6594
R7000 gnd.n374 gnd.n372 99.6594
R7001 gnd.n380 gnd.n178 99.6594
R7002 gnd.n383 gnd.n382 99.6594
R7003 gnd.n5648 gnd.n5647 99.6594
R7004 gnd.n5642 gnd.n3158 99.6594
R7005 gnd.n5639 gnd.n3159 99.6594
R7006 gnd.n5635 gnd.n3160 99.6594
R7007 gnd.n5631 gnd.n3161 99.6594
R7008 gnd.n5627 gnd.n3162 99.6594
R7009 gnd.n5623 gnd.n3163 99.6594
R7010 gnd.n5619 gnd.n3164 99.6594
R7011 gnd.n5615 gnd.n3165 99.6594
R7012 gnd.n5610 gnd.n3166 99.6594
R7013 gnd.n5606 gnd.n3167 99.6594
R7014 gnd.n5602 gnd.n3168 99.6594
R7015 gnd.n5598 gnd.n3169 99.6594
R7016 gnd.n5593 gnd.n3171 99.6594
R7017 gnd.n5589 gnd.n3172 99.6594
R7018 gnd.n5585 gnd.n3173 99.6594
R7019 gnd.n5581 gnd.n3174 99.6594
R7020 gnd.n5577 gnd.n3175 99.6594
R7021 gnd.n5573 gnd.n3176 99.6594
R7022 gnd.n5569 gnd.n3177 99.6594
R7023 gnd.n5565 gnd.n3178 99.6594
R7024 gnd.n5561 gnd.n3179 99.6594
R7025 gnd.n5557 gnd.n3180 99.6594
R7026 gnd.n5553 gnd.n3181 99.6594
R7027 gnd.n5549 gnd.n3182 99.6594
R7028 gnd.n5545 gnd.n3183 99.6594
R7029 gnd.n5541 gnd.n3184 99.6594
R7030 gnd.n5537 gnd.n3185 99.6594
R7031 gnd.n5964 gnd.n5963 99.6594
R7032 gnd.n5959 gnd.n2780 99.6594
R7033 gnd.n5955 gnd.n2779 99.6594
R7034 gnd.n5951 gnd.n2778 99.6594
R7035 gnd.n5947 gnd.n2777 99.6594
R7036 gnd.n5943 gnd.n2776 99.6594
R7037 gnd.n5939 gnd.n2775 99.6594
R7038 gnd.n5935 gnd.n2774 99.6594
R7039 gnd.n5930 gnd.n2773 99.6594
R7040 gnd.n5926 gnd.n2772 99.6594
R7041 gnd.n5922 gnd.n2771 99.6594
R7042 gnd.n5918 gnd.n2770 99.6594
R7043 gnd.n2906 gnd.n2768 99.6594
R7044 gnd.n2904 gnd.n2767 99.6594
R7045 gnd.n2900 gnd.n2766 99.6594
R7046 gnd.n2896 gnd.n2765 99.6594
R7047 gnd.n2892 gnd.n2764 99.6594
R7048 gnd.n2884 gnd.n2763 99.6594
R7049 gnd.n2882 gnd.n2762 99.6594
R7050 gnd.n2878 gnd.n2761 99.6594
R7051 gnd.n2874 gnd.n2760 99.6594
R7052 gnd.n2870 gnd.n2759 99.6594
R7053 gnd.n2866 gnd.n2758 99.6594
R7054 gnd.n2862 gnd.n2757 99.6594
R7055 gnd.n2858 gnd.n2756 99.6594
R7056 gnd.n2854 gnd.n2755 99.6594
R7057 gnd.n2850 gnd.n2754 99.6594
R7058 gnd.n2842 gnd.n2753 99.6594
R7059 gnd.n6275 gnd.n6274 99.6594
R7060 gnd.n6269 gnd.n2342 99.6594
R7061 gnd.n6266 gnd.n2343 99.6594
R7062 gnd.n6262 gnd.n2344 99.6594
R7063 gnd.n6258 gnd.n2345 99.6594
R7064 gnd.n6254 gnd.n2346 99.6594
R7065 gnd.n6250 gnd.n2347 99.6594
R7066 gnd.n6246 gnd.n2348 99.6594
R7067 gnd.n6242 gnd.n2349 99.6594
R7068 gnd.n6237 gnd.n2350 99.6594
R7069 gnd.n6233 gnd.n2351 99.6594
R7070 gnd.n6229 gnd.n2352 99.6594
R7071 gnd.n6225 gnd.n2353 99.6594
R7072 gnd.n6221 gnd.n2354 99.6594
R7073 gnd.n6217 gnd.n2355 99.6594
R7074 gnd.n6213 gnd.n2356 99.6594
R7075 gnd.n6209 gnd.n2357 99.6594
R7076 gnd.n6205 gnd.n2358 99.6594
R7077 gnd.n6201 gnd.n2359 99.6594
R7078 gnd.n6197 gnd.n2360 99.6594
R7079 gnd.n6193 gnd.n2361 99.6594
R7080 gnd.n6189 gnd.n2362 99.6594
R7081 gnd.n6185 gnd.n2363 99.6594
R7082 gnd.n6181 gnd.n2364 99.6594
R7083 gnd.n6177 gnd.n2365 99.6594
R7084 gnd.n6173 gnd.n2366 99.6594
R7085 gnd.n6169 gnd.n2367 99.6594
R7086 gnd.n6165 gnd.n2368 99.6594
R7087 gnd.n6161 gnd.n2369 99.6594
R7088 gnd.n6314 gnd.n6282 99.6594
R7089 gnd.n6312 gnd.n6281 99.6594
R7090 gnd.n6308 gnd.n6280 99.6594
R7091 gnd.n6304 gnd.n6279 99.6594
R7092 gnd.n6300 gnd.n6278 99.6594
R7093 gnd.n6296 gnd.n6277 99.6594
R7094 gnd.n6326 gnd.n6324 99.6594
R7095 gnd.n6332 gnd.n1050 99.6594
R7096 gnd.n1736 gnd.n1735 99.6594
R7097 gnd.n1730 gnd.n1678 99.6594
R7098 gnd.n1727 gnd.n1679 99.6594
R7099 gnd.n1723 gnd.n1680 99.6594
R7100 gnd.n1719 gnd.n1681 99.6594
R7101 gnd.n1715 gnd.n1682 99.6594
R7102 gnd.n1711 gnd.n1683 99.6594
R7103 gnd.n1707 gnd.n1684 99.6594
R7104 gnd.n7285 gnd.n7283 99.6594
R7105 gnd.n7291 gnd.n7276 99.6594
R7106 gnd.n7295 gnd.n7293 99.6594
R7107 gnd.n7301 gnd.n7272 99.6594
R7108 gnd.n7305 gnd.n7303 99.6594
R7109 gnd.n7311 gnd.n7268 99.6594
R7110 gnd.n7315 gnd.n7313 99.6594
R7111 gnd.n7321 gnd.n7264 99.6594
R7112 gnd.n7324 gnd.n7323 99.6594
R7113 gnd.n3270 gnd.n3186 99.6594
R7114 gnd.n3188 gnd.n3112 99.6594
R7115 gnd.n3189 gnd.n3119 99.6594
R7116 gnd.n3191 gnd.n3190 99.6594
R7117 gnd.n3193 gnd.n3128 99.6594
R7118 gnd.n3194 gnd.n3135 99.6594
R7119 gnd.n3196 gnd.n3195 99.6594
R7120 gnd.n3198 gnd.n3144 99.6594
R7121 gnd.n5650 gnd.n3153 99.6594
R7122 gnd.n1092 gnd.n1057 99.6594
R7123 gnd.n1096 gnd.n1058 99.6594
R7124 gnd.n1102 gnd.n1059 99.6594
R7125 gnd.n1106 gnd.n1060 99.6594
R7126 gnd.n1112 gnd.n1061 99.6594
R7127 gnd.n1116 gnd.n1062 99.6594
R7128 gnd.n1122 gnd.n1063 99.6594
R7129 gnd.n1126 gnd.n1064 99.6594
R7130 gnd.n1132 gnd.n1065 99.6594
R7131 gnd.n1136 gnd.n1066 99.6594
R7132 gnd.n1142 gnd.n1067 99.6594
R7133 gnd.n1145 gnd.n1068 99.6594
R7134 gnd.n2341 gnd.n2340 99.6594
R7135 gnd.n1495 gnd.n1405 99.6594
R7136 gnd.n1493 gnd.n1408 99.6594
R7137 gnd.n1489 gnd.n1488 99.6594
R7138 gnd.n1482 gnd.n1413 99.6594
R7139 gnd.n1481 gnd.n1480 99.6594
R7140 gnd.n1474 gnd.n1419 99.6594
R7141 gnd.n1473 gnd.n1472 99.6594
R7142 gnd.n1466 gnd.n1425 99.6594
R7143 gnd.n1465 gnd.n1464 99.6594
R7144 gnd.n1458 gnd.n1431 99.6594
R7145 gnd.n1457 gnd.n1456 99.6594
R7146 gnd.n1449 gnd.n1437 99.6594
R7147 gnd.n1448 gnd.n1447 99.6594
R7148 gnd.n2739 gnd.n2684 99.6594
R7149 gnd.n2741 gnd.n2693 99.6594
R7150 gnd.n2743 gnd.n2742 99.6594
R7151 gnd.n2744 gnd.n2702 99.6594
R7152 gnd.n2746 gnd.n2711 99.6594
R7153 gnd.n2748 gnd.n2747 99.6594
R7154 gnd.n2749 gnd.n2720 99.6594
R7155 gnd.n2751 gnd.n2732 99.6594
R7156 gnd.n5967 gnd.n5966 99.6594
R7157 gnd.n4109 gnd.n2370 99.6594
R7158 gnd.n4113 gnd.n2371 99.6594
R7159 gnd.n4119 gnd.n2372 99.6594
R7160 gnd.n4123 gnd.n2373 99.6594
R7161 gnd.n4129 gnd.n2374 99.6594
R7162 gnd.n4133 gnd.n2375 99.6594
R7163 gnd.n4139 gnd.n2376 99.6594
R7164 gnd.n4143 gnd.n2377 99.6594
R7165 gnd.n4100 gnd.n2378 99.6594
R7166 gnd.n4112 gnd.n2370 99.6594
R7167 gnd.n4118 gnd.n2371 99.6594
R7168 gnd.n4122 gnd.n2372 99.6594
R7169 gnd.n4128 gnd.n2373 99.6594
R7170 gnd.n4132 gnd.n2374 99.6594
R7171 gnd.n4138 gnd.n2375 99.6594
R7172 gnd.n4142 gnd.n2376 99.6594
R7173 gnd.n4099 gnd.n2377 99.6594
R7174 gnd.n4095 gnd.n2378 99.6594
R7175 gnd.n5966 gnd.n2737 99.6594
R7176 gnd.n2751 gnd.n2750 99.6594
R7177 gnd.n2749 gnd.n2719 99.6594
R7178 gnd.n2748 gnd.n2712 99.6594
R7179 gnd.n2746 gnd.n2745 99.6594
R7180 gnd.n2744 gnd.n2701 99.6594
R7181 gnd.n2743 gnd.n2694 99.6594
R7182 gnd.n2741 gnd.n2740 99.6594
R7183 gnd.n2739 gnd.n2683 99.6594
R7184 gnd.n1496 gnd.n1495 99.6594
R7185 gnd.n1490 gnd.n1408 99.6594
R7186 gnd.n1488 gnd.n1487 99.6594
R7187 gnd.n1483 gnd.n1482 99.6594
R7188 gnd.n1480 gnd.n1479 99.6594
R7189 gnd.n1475 gnd.n1474 99.6594
R7190 gnd.n1472 gnd.n1471 99.6594
R7191 gnd.n1467 gnd.n1466 99.6594
R7192 gnd.n1464 gnd.n1463 99.6594
R7193 gnd.n1459 gnd.n1458 99.6594
R7194 gnd.n1456 gnd.n1455 99.6594
R7195 gnd.n1450 gnd.n1449 99.6594
R7196 gnd.n1447 gnd.n1403 99.6594
R7197 gnd.n2341 gnd.n1069 99.6594
R7198 gnd.n1143 gnd.n1068 99.6594
R7199 gnd.n1135 gnd.n1067 99.6594
R7200 gnd.n1133 gnd.n1066 99.6594
R7201 gnd.n1125 gnd.n1065 99.6594
R7202 gnd.n1123 gnd.n1064 99.6594
R7203 gnd.n1115 gnd.n1063 99.6594
R7204 gnd.n1113 gnd.n1062 99.6594
R7205 gnd.n1105 gnd.n1061 99.6594
R7206 gnd.n1103 gnd.n1060 99.6594
R7207 gnd.n1095 gnd.n1059 99.6594
R7208 gnd.n1093 gnd.n1058 99.6594
R7209 gnd.n1085 gnd.n1057 99.6594
R7210 gnd.n3186 gnd.n3111 99.6594
R7211 gnd.n3188 gnd.n3187 99.6594
R7212 gnd.n3189 gnd.n3120 99.6594
R7213 gnd.n3191 gnd.n3127 99.6594
R7214 gnd.n3193 gnd.n3192 99.6594
R7215 gnd.n3194 gnd.n3136 99.6594
R7216 gnd.n3196 gnd.n3143 99.6594
R7217 gnd.n3198 gnd.n3197 99.6594
R7218 gnd.n5651 gnd.n5650 99.6594
R7219 gnd.n7323 gnd.n7322 99.6594
R7220 gnd.n7314 gnd.n7264 99.6594
R7221 gnd.n7313 gnd.n7312 99.6594
R7222 gnd.n7304 gnd.n7268 99.6594
R7223 gnd.n7303 gnd.n7302 99.6594
R7224 gnd.n7294 gnd.n7272 99.6594
R7225 gnd.n7293 gnd.n7292 99.6594
R7226 gnd.n7284 gnd.n7276 99.6594
R7227 gnd.n7283 gnd.n7282 99.6594
R7228 gnd.n1736 gnd.n1686 99.6594
R7229 gnd.n1728 gnd.n1678 99.6594
R7230 gnd.n1724 gnd.n1679 99.6594
R7231 gnd.n1720 gnd.n1680 99.6594
R7232 gnd.n1716 gnd.n1681 99.6594
R7233 gnd.n1712 gnd.n1682 99.6594
R7234 gnd.n1708 gnd.n1683 99.6594
R7235 gnd.n1684 gnd.n1365 99.6594
R7236 gnd.n6325 gnd.n1050 99.6594
R7237 gnd.n6324 gnd.n1056 99.6594
R7238 gnd.n6299 gnd.n6277 99.6594
R7239 gnd.n6303 gnd.n6278 99.6594
R7240 gnd.n6307 gnd.n6279 99.6594
R7241 gnd.n6311 gnd.n6280 99.6594
R7242 gnd.n6315 gnd.n6281 99.6594
R7243 gnd.n6283 gnd.n6282 99.6594
R7244 gnd.n6275 gnd.n2382 99.6594
R7245 gnd.n6267 gnd.n2342 99.6594
R7246 gnd.n6263 gnd.n2343 99.6594
R7247 gnd.n6259 gnd.n2344 99.6594
R7248 gnd.n6255 gnd.n2345 99.6594
R7249 gnd.n6251 gnd.n2346 99.6594
R7250 gnd.n6247 gnd.n2347 99.6594
R7251 gnd.n6243 gnd.n2348 99.6594
R7252 gnd.n6238 gnd.n2349 99.6594
R7253 gnd.n6234 gnd.n2350 99.6594
R7254 gnd.n6230 gnd.n2351 99.6594
R7255 gnd.n6226 gnd.n2352 99.6594
R7256 gnd.n6222 gnd.n2353 99.6594
R7257 gnd.n6218 gnd.n2354 99.6594
R7258 gnd.n6214 gnd.n2355 99.6594
R7259 gnd.n6210 gnd.n2356 99.6594
R7260 gnd.n6206 gnd.n2357 99.6594
R7261 gnd.n6202 gnd.n2358 99.6594
R7262 gnd.n6198 gnd.n2359 99.6594
R7263 gnd.n6194 gnd.n2360 99.6594
R7264 gnd.n6190 gnd.n2361 99.6594
R7265 gnd.n6186 gnd.n2362 99.6594
R7266 gnd.n6182 gnd.n2363 99.6594
R7267 gnd.n6178 gnd.n2364 99.6594
R7268 gnd.n6174 gnd.n2365 99.6594
R7269 gnd.n6170 gnd.n2366 99.6594
R7270 gnd.n6166 gnd.n2367 99.6594
R7271 gnd.n6162 gnd.n2368 99.6594
R7272 gnd.n2452 gnd.n2369 99.6594
R7273 gnd.n2849 gnd.n2753 99.6594
R7274 gnd.n2853 gnd.n2754 99.6594
R7275 gnd.n2857 gnd.n2755 99.6594
R7276 gnd.n2861 gnd.n2756 99.6594
R7277 gnd.n2865 gnd.n2757 99.6594
R7278 gnd.n2869 gnd.n2758 99.6594
R7279 gnd.n2873 gnd.n2759 99.6594
R7280 gnd.n2877 gnd.n2760 99.6594
R7281 gnd.n2881 gnd.n2761 99.6594
R7282 gnd.n2885 gnd.n2762 99.6594
R7283 gnd.n2891 gnd.n2763 99.6594
R7284 gnd.n2895 gnd.n2764 99.6594
R7285 gnd.n2899 gnd.n2765 99.6594
R7286 gnd.n2903 gnd.n2766 99.6594
R7287 gnd.n2907 gnd.n2767 99.6594
R7288 gnd.n5917 gnd.n2769 99.6594
R7289 gnd.n5921 gnd.n2770 99.6594
R7290 gnd.n5925 gnd.n2771 99.6594
R7291 gnd.n5929 gnd.n2772 99.6594
R7292 gnd.n5934 gnd.n2773 99.6594
R7293 gnd.n5938 gnd.n2774 99.6594
R7294 gnd.n5942 gnd.n2775 99.6594
R7295 gnd.n5946 gnd.n2776 99.6594
R7296 gnd.n5950 gnd.n2777 99.6594
R7297 gnd.n5954 gnd.n2778 99.6594
R7298 gnd.n5958 gnd.n2779 99.6594
R7299 gnd.n2782 gnd.n2780 99.6594
R7300 gnd.n5964 gnd.n2781 99.6594
R7301 gnd.n5648 gnd.n3201 99.6594
R7302 gnd.n5640 gnd.n3158 99.6594
R7303 gnd.n5636 gnd.n3159 99.6594
R7304 gnd.n5632 gnd.n3160 99.6594
R7305 gnd.n5628 gnd.n3161 99.6594
R7306 gnd.n5624 gnd.n3162 99.6594
R7307 gnd.n5620 gnd.n3163 99.6594
R7308 gnd.n5616 gnd.n3164 99.6594
R7309 gnd.n5611 gnd.n3165 99.6594
R7310 gnd.n5607 gnd.n3166 99.6594
R7311 gnd.n5603 gnd.n3167 99.6594
R7312 gnd.n5599 gnd.n3168 99.6594
R7313 gnd.n5594 gnd.n3170 99.6594
R7314 gnd.n5590 gnd.n3171 99.6594
R7315 gnd.n5586 gnd.n3172 99.6594
R7316 gnd.n5582 gnd.n3173 99.6594
R7317 gnd.n5578 gnd.n3174 99.6594
R7318 gnd.n5574 gnd.n3175 99.6594
R7319 gnd.n5570 gnd.n3176 99.6594
R7320 gnd.n5566 gnd.n3177 99.6594
R7321 gnd.n5562 gnd.n3178 99.6594
R7322 gnd.n5558 gnd.n3179 99.6594
R7323 gnd.n5554 gnd.n3180 99.6594
R7324 gnd.n5550 gnd.n3181 99.6594
R7325 gnd.n5546 gnd.n3182 99.6594
R7326 gnd.n5542 gnd.n3183 99.6594
R7327 gnd.n5538 gnd.n3184 99.6594
R7328 gnd.n5530 gnd.n3185 99.6594
R7329 gnd.n382 gnd.n381 99.6594
R7330 gnd.n373 gnd.n178 99.6594
R7331 gnd.n372 gnd.n371 99.6594
R7332 gnd.n363 gnd.n182 99.6594
R7333 gnd.n362 gnd.n361 99.6594
R7334 gnd.n353 gnd.n186 99.6594
R7335 gnd.n352 gnd.n351 99.6594
R7336 gnd.n343 gnd.n190 99.6594
R7337 gnd.n342 gnd.n341 99.6594
R7338 gnd.n333 gnd.n194 99.6594
R7339 gnd.n332 gnd.n331 99.6594
R7340 gnd.n323 gnd.n200 99.6594
R7341 gnd.n322 gnd.n321 99.6594
R7342 gnd.n313 gnd.n204 99.6594
R7343 gnd.n312 gnd.n311 99.6594
R7344 gnd.n303 gnd.n208 99.6594
R7345 gnd.n302 gnd.n301 99.6594
R7346 gnd.n293 gnd.n212 99.6594
R7347 gnd.n292 gnd.n291 99.6594
R7348 gnd.n283 gnd.n216 99.6594
R7349 gnd.n282 gnd.n281 99.6594
R7350 gnd.n273 gnd.n272 99.6594
R7351 gnd.n271 gnd.n270 99.6594
R7352 gnd.n262 gnd.n226 99.6594
R7353 gnd.n261 gnd.n260 99.6594
R7354 gnd.n252 gnd.n230 99.6594
R7355 gnd.n251 gnd.n250 99.6594
R7356 gnd.n242 gnd.n234 99.6594
R7357 gnd.n241 gnd.n240 99.6594
R7358 gnd.n6029 gnd.n6028 99.6594
R7359 gnd.n2670 gnd.n2650 99.6594
R7360 gnd.n2672 gnd.n2651 99.6594
R7361 gnd.n2676 gnd.n2652 99.6594
R7362 gnd.n2678 gnd.n2653 99.6594
R7363 gnd.n2688 gnd.n2654 99.6594
R7364 gnd.n2690 gnd.n2655 99.6594
R7365 gnd.n2698 gnd.n2656 99.6594
R7366 gnd.n2706 gnd.n2657 99.6594
R7367 gnd.n2708 gnd.n2658 99.6594
R7368 gnd.n2716 gnd.n2659 99.6594
R7369 gnd.n2724 gnd.n2660 99.6594
R7370 gnd.n2729 gnd.n2662 99.6594
R7371 gnd.n6031 gnd.n2647 99.6594
R7372 gnd.n6029 gnd.n2665 99.6594
R7373 gnd.n2671 gnd.n2650 99.6594
R7374 gnd.n2675 gnd.n2651 99.6594
R7375 gnd.n2677 gnd.n2652 99.6594
R7376 gnd.n2687 gnd.n2653 99.6594
R7377 gnd.n2689 gnd.n2654 99.6594
R7378 gnd.n2697 gnd.n2655 99.6594
R7379 gnd.n2705 gnd.n2656 99.6594
R7380 gnd.n2707 gnd.n2657 99.6594
R7381 gnd.n2715 gnd.n2658 99.6594
R7382 gnd.n2723 gnd.n2659 99.6594
R7383 gnd.n2725 gnd.n2660 99.6594
R7384 gnd.n2662 gnd.n2661 99.6594
R7385 gnd.n6032 gnd.n6031 99.6594
R7386 gnd.n3423 gnd.n3096 99.6594
R7387 gnd.n3425 gnd.n3424 99.6594
R7388 gnd.n3426 gnd.n3101 99.6594
R7389 gnd.n3428 gnd.n3427 99.6594
R7390 gnd.n3429 gnd.n3107 99.6594
R7391 gnd.n3431 gnd.n3115 99.6594
R7392 gnd.n3433 gnd.n3432 99.6594
R7393 gnd.n3434 gnd.n3124 99.6594
R7394 gnd.n3436 gnd.n3131 99.6594
R7395 gnd.n3438 gnd.n3437 99.6594
R7396 gnd.n3439 gnd.n3140 99.6594
R7397 gnd.n3441 gnd.n3147 99.6594
R7398 gnd.n3444 gnd.n3443 99.6594
R7399 gnd.n5299 gnd.n5298 99.6594
R7400 gnd.n3441 gnd.n3440 99.6594
R7401 gnd.n3439 gnd.n3139 99.6594
R7402 gnd.n3438 gnd.n3132 99.6594
R7403 gnd.n3436 gnd.n3435 99.6594
R7404 gnd.n3434 gnd.n3123 99.6594
R7405 gnd.n3433 gnd.n3116 99.6594
R7406 gnd.n3431 gnd.n3430 99.6594
R7407 gnd.n3429 gnd.n3106 99.6594
R7408 gnd.n3428 gnd.n3102 99.6594
R7409 gnd.n3426 gnd.n3100 99.6594
R7410 gnd.n3425 gnd.n3097 99.6594
R7411 gnd.n3423 gnd.n3092 99.6594
R7412 gnd.n5298 gnd.n3087 99.6594
R7413 gnd.n3444 gnd.n3422 99.6594
R7414 gnd.n2726 gnd.t82 98.63
R7415 gnd.n5652 gnd.t52 98.63
R7416 gnd.n2733 gnd.t67 98.63
R7417 gnd.n3221 gnd.t125 98.63
R7418 gnd.n3244 gnd.t131 98.63
R7419 gnd.n5532 gnd.t95 98.63
R7420 gnd.n175 gnd.t91 98.63
R7421 gnd.n197 gnd.t100 98.63
R7422 gnd.n219 gnd.t106 98.63
R7423 gnd.n7261 gnd.t37 98.63
R7424 gnd.n2402 gnd.t85 98.63
R7425 gnd.n2424 gnd.t110 98.63
R7426 gnd.n2446 gnd.t116 98.63
R7427 gnd.n4096 gnd.t60 98.63
R7428 gnd.n2803 gnd.t103 98.63
R7429 gnd.n2844 gnd.t118 98.63
R7430 gnd.n2823 gnd.t141 98.63
R7431 gnd.n3149 gnd.t55 98.63
R7432 gnd.n3772 gnd.t150 88.9408
R7433 gnd.n5017 gnd.t152 88.9408
R7434 gnd.n5846 gnd.t75 88.933
R7435 gnd.n5011 gnd.t63 88.933
R7436 gnd.n2961 gnd.n2960 81.8399
R7437 gnd.n1704 gnd.t88 74.8376
R7438 gnd.n1052 gnd.t135 74.8376
R7439 gnd.n3773 gnd.t149 72.8438
R7440 gnd.n5018 gnd.t153 72.8438
R7441 gnd.n2962 gnd.n2955 72.8411
R7442 gnd.n2968 gnd.n2953 72.8411
R7443 gnd.n4985 gnd.n4984 72.8411
R7444 gnd.n2727 gnd.t81 72.836
R7445 gnd.n5847 gnd.t74 72.836
R7446 gnd.n5012 gnd.t64 72.836
R7447 gnd.n5653 gnd.t51 72.836
R7448 gnd.n2734 gnd.t68 72.836
R7449 gnd.n3222 gnd.t124 72.836
R7450 gnd.n3245 gnd.t130 72.836
R7451 gnd.n5533 gnd.t94 72.836
R7452 gnd.n176 gnd.t92 72.836
R7453 gnd.n198 gnd.t101 72.836
R7454 gnd.n220 gnd.t107 72.836
R7455 gnd.n7262 gnd.t38 72.836
R7456 gnd.n2403 gnd.t84 72.836
R7457 gnd.n2425 gnd.t109 72.836
R7458 gnd.n2447 gnd.t115 72.836
R7459 gnd.n4097 gnd.t59 72.836
R7460 gnd.n2804 gnd.t104 72.836
R7461 gnd.n2845 gnd.t119 72.836
R7462 gnd.n2824 gnd.t142 72.836
R7463 gnd.n3150 gnd.t56 72.836
R7464 gnd.n5155 gnd.n4990 71.676
R7465 gnd.n5153 gnd.n5152 71.676
R7466 gnd.n5148 gnd.n4994 71.676
R7467 gnd.n5146 gnd.n5145 71.676
R7468 gnd.n5141 gnd.n4997 71.676
R7469 gnd.n5139 gnd.n5138 71.676
R7470 gnd.n5134 gnd.n5000 71.676
R7471 gnd.n5132 gnd.n5131 71.676
R7472 gnd.n5127 gnd.n5003 71.676
R7473 gnd.n5125 gnd.n5124 71.676
R7474 gnd.n5120 gnd.n5006 71.676
R7475 gnd.n5118 gnd.n5117 71.676
R7476 gnd.n5113 gnd.n5009 71.676
R7477 gnd.n5111 gnd.n5110 71.676
R7478 gnd.n5105 gnd.n5014 71.676
R7479 gnd.n5103 gnd.n5102 71.676
R7480 gnd.n5098 gnd.n5097 71.676
R7481 gnd.n5095 gnd.n5094 71.676
R7482 gnd.n5089 gnd.n5020 71.676
R7483 gnd.n5087 gnd.n5086 71.676
R7484 gnd.n5082 gnd.n5023 71.676
R7485 gnd.n5080 gnd.n5079 71.676
R7486 gnd.n5075 gnd.n5026 71.676
R7487 gnd.n5073 gnd.n5072 71.676
R7488 gnd.n5068 gnd.n5029 71.676
R7489 gnd.n5066 gnd.n5065 71.676
R7490 gnd.n5061 gnd.n5032 71.676
R7491 gnd.n5059 gnd.n5058 71.676
R7492 gnd.n5054 gnd.n5035 71.676
R7493 gnd.n5052 gnd.n5051 71.676
R7494 gnd.n5047 gnd.n5038 71.676
R7495 gnd.n5045 gnd.n5044 71.676
R7496 gnd.n5039 gnd.n3531 71.676
R7497 gnd.n5910 gnd.n5909 71.676
R7498 gnd.n5904 gnd.n2917 71.676
R7499 gnd.n5901 gnd.n2918 71.676
R7500 gnd.n5897 gnd.n2919 71.676
R7501 gnd.n5893 gnd.n2920 71.676
R7502 gnd.n5889 gnd.n2921 71.676
R7503 gnd.n5885 gnd.n2922 71.676
R7504 gnd.n5881 gnd.n2923 71.676
R7505 gnd.n5877 gnd.n2924 71.676
R7506 gnd.n5873 gnd.n2925 71.676
R7507 gnd.n5869 gnd.n2926 71.676
R7508 gnd.n5865 gnd.n2927 71.676
R7509 gnd.n5861 gnd.n2928 71.676
R7510 gnd.n5857 gnd.n2929 71.676
R7511 gnd.n5853 gnd.n2930 71.676
R7512 gnd.n5849 gnd.n2931 71.676
R7513 gnd.n2932 gnd.n2915 71.676
R7514 gnd.n3776 gnd.n2933 71.676
R7515 gnd.n3781 gnd.n2934 71.676
R7516 gnd.n3785 gnd.n2935 71.676
R7517 gnd.n3789 gnd.n2936 71.676
R7518 gnd.n3793 gnd.n2937 71.676
R7519 gnd.n3797 gnd.n2938 71.676
R7520 gnd.n3801 gnd.n2939 71.676
R7521 gnd.n3805 gnd.n2940 71.676
R7522 gnd.n3809 gnd.n2941 71.676
R7523 gnd.n3813 gnd.n2942 71.676
R7524 gnd.n3817 gnd.n2943 71.676
R7525 gnd.n3821 gnd.n2944 71.676
R7526 gnd.n3825 gnd.n2945 71.676
R7527 gnd.n3829 gnd.n2946 71.676
R7528 gnd.n3833 gnd.n2947 71.676
R7529 gnd.n5910 gnd.n2950 71.676
R7530 gnd.n5902 gnd.n2917 71.676
R7531 gnd.n5898 gnd.n2918 71.676
R7532 gnd.n5894 gnd.n2919 71.676
R7533 gnd.n5890 gnd.n2920 71.676
R7534 gnd.n5886 gnd.n2921 71.676
R7535 gnd.n5882 gnd.n2922 71.676
R7536 gnd.n5878 gnd.n2923 71.676
R7537 gnd.n5874 gnd.n2924 71.676
R7538 gnd.n5870 gnd.n2925 71.676
R7539 gnd.n5866 gnd.n2926 71.676
R7540 gnd.n5862 gnd.n2927 71.676
R7541 gnd.n5858 gnd.n2928 71.676
R7542 gnd.n5854 gnd.n2929 71.676
R7543 gnd.n5850 gnd.n2930 71.676
R7544 gnd.n5913 gnd.n5912 71.676
R7545 gnd.n3775 gnd.n2932 71.676
R7546 gnd.n3780 gnd.n2933 71.676
R7547 gnd.n3784 gnd.n2934 71.676
R7548 gnd.n3788 gnd.n2935 71.676
R7549 gnd.n3792 gnd.n2936 71.676
R7550 gnd.n3796 gnd.n2937 71.676
R7551 gnd.n3800 gnd.n2938 71.676
R7552 gnd.n3804 gnd.n2939 71.676
R7553 gnd.n3808 gnd.n2940 71.676
R7554 gnd.n3812 gnd.n2941 71.676
R7555 gnd.n3816 gnd.n2942 71.676
R7556 gnd.n3820 gnd.n2943 71.676
R7557 gnd.n3824 gnd.n2944 71.676
R7558 gnd.n3828 gnd.n2945 71.676
R7559 gnd.n3832 gnd.n2946 71.676
R7560 gnd.n3836 gnd.n2947 71.676
R7561 gnd.n5040 gnd.n5039 71.676
R7562 gnd.n5046 gnd.n5045 71.676
R7563 gnd.n5038 gnd.n5036 71.676
R7564 gnd.n5053 gnd.n5052 71.676
R7565 gnd.n5035 gnd.n5033 71.676
R7566 gnd.n5060 gnd.n5059 71.676
R7567 gnd.n5032 gnd.n5030 71.676
R7568 gnd.n5067 gnd.n5066 71.676
R7569 gnd.n5029 gnd.n5027 71.676
R7570 gnd.n5074 gnd.n5073 71.676
R7571 gnd.n5026 gnd.n5024 71.676
R7572 gnd.n5081 gnd.n5080 71.676
R7573 gnd.n5023 gnd.n5021 71.676
R7574 gnd.n5088 gnd.n5087 71.676
R7575 gnd.n5020 gnd.n5016 71.676
R7576 gnd.n5096 gnd.n5095 71.676
R7577 gnd.n5100 gnd.n5099 71.676
R7578 gnd.n5104 gnd.n5103 71.676
R7579 gnd.n5014 gnd.n5010 71.676
R7580 gnd.n5112 gnd.n5111 71.676
R7581 gnd.n5009 gnd.n5007 71.676
R7582 gnd.n5119 gnd.n5118 71.676
R7583 gnd.n5006 gnd.n5004 71.676
R7584 gnd.n5126 gnd.n5125 71.676
R7585 gnd.n5003 gnd.n5001 71.676
R7586 gnd.n5133 gnd.n5132 71.676
R7587 gnd.n5000 gnd.n4998 71.676
R7588 gnd.n5140 gnd.n5139 71.676
R7589 gnd.n4997 gnd.n4995 71.676
R7590 gnd.n5147 gnd.n5146 71.676
R7591 gnd.n4994 gnd.n4992 71.676
R7592 gnd.n5154 gnd.n5153 71.676
R7593 gnd.n4990 gnd.n3534 71.676
R7594 gnd.n10 gnd.t24 69.1507
R7595 gnd.n18 gnd.t22 68.4792
R7596 gnd.n17 gnd.t210 68.4792
R7597 gnd.n16 gnd.t7 68.4792
R7598 gnd.n15 gnd.t173 68.4792
R7599 gnd.n14 gnd.t19 68.4792
R7600 gnd.n13 gnd.t159 68.4792
R7601 gnd.n12 gnd.t332 68.4792
R7602 gnd.n11 gnd.t177 68.4792
R7603 gnd.n10 gnd.t191 68.4792
R7604 gnd.n1503 gnd.n1404 64.369
R7605 gnd.n6276 gnd.n2380 63.0944
R7606 gnd.n7357 gnd.n171 63.0944
R7607 gnd.n3778 gnd.n3773 59.5399
R7608 gnd.n5091 gnd.n5018 59.5399
R7609 gnd.n5848 gnd.n5847 59.5399
R7610 gnd.n5107 gnd.n5012 59.5399
R7611 gnd.n5845 gnd.n2971 59.1804
R7612 gnd.n6323 gnd.n1043 57.3586
R7613 gnd.n1632 gnd.t305 56.407
R7614 gnd.n1597 gnd.t319 56.407
R7615 gnd.n1608 gnd.t291 56.407
R7616 gnd.n1620 gnd.t224 56.407
R7617 gnd.n56 gnd.t284 56.407
R7618 gnd.n21 gnd.t230 56.407
R7619 gnd.n32 gnd.t272 56.407
R7620 gnd.n44 gnd.t313 56.407
R7621 gnd.n1641 gnd.t242 55.8337
R7622 gnd.n1606 gnd.t315 55.8337
R7623 gnd.n1617 gnd.t283 55.8337
R7624 gnd.n1629 gnd.t296 55.8337
R7625 gnd.n65 gnd.t321 55.8337
R7626 gnd.n30 gnd.t216 55.8337
R7627 gnd.n41 gnd.t257 55.8337
R7628 gnd.n53 gnd.t261 55.8337
R7629 gnd.n2959 gnd.n2958 54.358
R7630 gnd.n4982 gnd.n4981 54.358
R7631 gnd.n1632 gnd.n1631 53.0052
R7632 gnd.n1634 gnd.n1633 53.0052
R7633 gnd.n1636 gnd.n1635 53.0052
R7634 gnd.n1638 gnd.n1637 53.0052
R7635 gnd.n1640 gnd.n1639 53.0052
R7636 gnd.n1597 gnd.n1596 53.0052
R7637 gnd.n1599 gnd.n1598 53.0052
R7638 gnd.n1601 gnd.n1600 53.0052
R7639 gnd.n1603 gnd.n1602 53.0052
R7640 gnd.n1605 gnd.n1604 53.0052
R7641 gnd.n1608 gnd.n1607 53.0052
R7642 gnd.n1610 gnd.n1609 53.0052
R7643 gnd.n1612 gnd.n1611 53.0052
R7644 gnd.n1614 gnd.n1613 53.0052
R7645 gnd.n1616 gnd.n1615 53.0052
R7646 gnd.n1620 gnd.n1619 53.0052
R7647 gnd.n1622 gnd.n1621 53.0052
R7648 gnd.n1624 gnd.n1623 53.0052
R7649 gnd.n1626 gnd.n1625 53.0052
R7650 gnd.n1628 gnd.n1627 53.0052
R7651 gnd.n64 gnd.n63 53.0052
R7652 gnd.n62 gnd.n61 53.0052
R7653 gnd.n60 gnd.n59 53.0052
R7654 gnd.n58 gnd.n57 53.0052
R7655 gnd.n56 gnd.n55 53.0052
R7656 gnd.n29 gnd.n28 53.0052
R7657 gnd.n27 gnd.n26 53.0052
R7658 gnd.n25 gnd.n24 53.0052
R7659 gnd.n23 gnd.n22 53.0052
R7660 gnd.n21 gnd.n20 53.0052
R7661 gnd.n40 gnd.n39 53.0052
R7662 gnd.n38 gnd.n37 53.0052
R7663 gnd.n36 gnd.n35 53.0052
R7664 gnd.n34 gnd.n33 53.0052
R7665 gnd.n32 gnd.n31 53.0052
R7666 gnd.n52 gnd.n51 53.0052
R7667 gnd.n50 gnd.n49 53.0052
R7668 gnd.n48 gnd.n47 53.0052
R7669 gnd.n46 gnd.n45 53.0052
R7670 gnd.n44 gnd.n43 53.0052
R7671 gnd.n4973 gnd.n4972 52.4801
R7672 gnd.n2294 gnd.t171 52.3082
R7673 gnd.n2262 gnd.t32 52.3082
R7674 gnd.n2230 gnd.t181 52.3082
R7675 gnd.n2199 gnd.t161 52.3082
R7676 gnd.n2167 gnd.t208 52.3082
R7677 gnd.n2135 gnd.t334 52.3082
R7678 gnd.n2103 gnd.t195 52.3082
R7679 gnd.n2072 gnd.t165 52.3082
R7680 gnd.n2124 gnd.n2092 51.4173
R7681 gnd.n2188 gnd.n2187 50.455
R7682 gnd.n2156 gnd.n2155 50.455
R7683 gnd.n2124 gnd.n2123 50.455
R7684 gnd.n1441 gnd.n1440 45.1884
R7685 gnd.n1073 gnd.n1072 45.1884
R7686 gnd.n5158 gnd.n4988 44.3322
R7687 gnd.n2962 gnd.n2961 44.3189
R7688 gnd.n2728 gnd.n2727 42.4732
R7689 gnd.n3151 gnd.n3150 42.4732
R7690 gnd.n5654 gnd.n5653 42.2793
R7691 gnd.n1453 gnd.n1441 42.2793
R7692 gnd.n1074 gnd.n1073 42.2793
R7693 gnd.n1706 gnd.n1704 42.2793
R7694 gnd.n1053 gnd.n1052 42.2793
R7695 gnd.n5969 gnd.n2734 42.2793
R7696 gnd.n5613 gnd.n3222 42.2793
R7697 gnd.n5576 gnd.n3245 42.2793
R7698 gnd.n5536 gnd.n5533 42.2793
R7699 gnd.n177 gnd.n176 42.2793
R7700 gnd.n199 gnd.n198 42.2793
R7701 gnd.n221 gnd.n220 42.2793
R7702 gnd.n7263 gnd.n7262 42.2793
R7703 gnd.n6240 gnd.n2403 42.2793
R7704 gnd.n6200 gnd.n2425 42.2793
R7705 gnd.n6160 gnd.n2447 42.2793
R7706 gnd.n4149 gnd.n4097 42.2793
R7707 gnd.n5932 gnd.n2804 42.2793
R7708 gnd.n2848 gnd.n2845 42.2793
R7709 gnd.n2890 gnd.n2824 42.2793
R7710 gnd.n2960 gnd.n2959 41.6274
R7711 gnd.n4983 gnd.n4982 41.6274
R7712 gnd.n2969 gnd.n2968 40.8975
R7713 gnd.n4986 gnd.n4985 40.8975
R7714 gnd.n6543 gnd.n6542 40.1465
R7715 gnd.n6542 gnd.n810 40.1465
R7716 gnd.n6536 gnd.n810 40.1465
R7717 gnd.n6536 gnd.n6535 40.1465
R7718 gnd.n6535 gnd.n6534 40.1465
R7719 gnd.n6534 gnd.n818 40.1465
R7720 gnd.n6528 gnd.n818 40.1465
R7721 gnd.n6528 gnd.n6527 40.1465
R7722 gnd.n6527 gnd.n6526 40.1465
R7723 gnd.n6526 gnd.n826 40.1465
R7724 gnd.n6520 gnd.n826 40.1465
R7725 gnd.n6520 gnd.n6519 40.1465
R7726 gnd.n6519 gnd.n6518 40.1465
R7727 gnd.n6518 gnd.n834 40.1465
R7728 gnd.n6512 gnd.n834 40.1465
R7729 gnd.n6512 gnd.n6511 40.1465
R7730 gnd.n6511 gnd.n6510 40.1465
R7731 gnd.n6510 gnd.n842 40.1465
R7732 gnd.n6504 gnd.n842 40.1465
R7733 gnd.n6504 gnd.n6503 40.1465
R7734 gnd.n6503 gnd.n6502 40.1465
R7735 gnd.n6502 gnd.n850 40.1465
R7736 gnd.n6496 gnd.n850 40.1465
R7737 gnd.n6496 gnd.n6495 40.1465
R7738 gnd.n6495 gnd.n6494 40.1465
R7739 gnd.n6494 gnd.n858 40.1465
R7740 gnd.n6488 gnd.n858 40.1465
R7741 gnd.n6488 gnd.n6487 40.1465
R7742 gnd.n6487 gnd.n6486 40.1465
R7743 gnd.n6486 gnd.n866 40.1465
R7744 gnd.n6480 gnd.n866 40.1465
R7745 gnd.n6480 gnd.n6479 40.1465
R7746 gnd.n6479 gnd.n6478 40.1465
R7747 gnd.n6478 gnd.n874 40.1465
R7748 gnd.n6472 gnd.n874 40.1465
R7749 gnd.n6472 gnd.n6471 40.1465
R7750 gnd.n6471 gnd.n6470 40.1465
R7751 gnd.n6470 gnd.n882 40.1465
R7752 gnd.n6464 gnd.n882 40.1465
R7753 gnd.n6464 gnd.n6463 40.1465
R7754 gnd.n6463 gnd.n6462 40.1465
R7755 gnd.n6462 gnd.n890 40.1465
R7756 gnd.n6456 gnd.n890 40.1465
R7757 gnd.n6456 gnd.n6455 40.1465
R7758 gnd.n6455 gnd.n6454 40.1465
R7759 gnd.n6454 gnd.n898 40.1465
R7760 gnd.n6448 gnd.n898 40.1465
R7761 gnd.n6448 gnd.n6447 40.1465
R7762 gnd.n6447 gnd.n6446 40.1465
R7763 gnd.n6446 gnd.n906 40.1465
R7764 gnd.n6440 gnd.n906 40.1465
R7765 gnd.n6440 gnd.n6439 40.1465
R7766 gnd.n6439 gnd.n6438 40.1465
R7767 gnd.n6438 gnd.n914 40.1465
R7768 gnd.n6432 gnd.n914 40.1465
R7769 gnd.n6432 gnd.n6431 40.1465
R7770 gnd.n6431 gnd.n6430 40.1465
R7771 gnd.n6430 gnd.n922 40.1465
R7772 gnd.n6424 gnd.n922 40.1465
R7773 gnd.n6424 gnd.n6423 40.1465
R7774 gnd.n6423 gnd.n6422 40.1465
R7775 gnd.n6422 gnd.n930 40.1465
R7776 gnd.n6416 gnd.n930 40.1465
R7777 gnd.n6416 gnd.n6415 40.1465
R7778 gnd.n6415 gnd.n6414 40.1465
R7779 gnd.n6414 gnd.n938 40.1465
R7780 gnd.n6408 gnd.n938 40.1465
R7781 gnd.n6408 gnd.n6407 40.1465
R7782 gnd.n6407 gnd.n6406 40.1465
R7783 gnd.n6406 gnd.n946 40.1465
R7784 gnd.n6400 gnd.n946 40.1465
R7785 gnd.n6400 gnd.n6399 40.1465
R7786 gnd.n6399 gnd.n6398 40.1465
R7787 gnd.n6398 gnd.n954 40.1465
R7788 gnd.n6392 gnd.n954 40.1465
R7789 gnd.n6392 gnd.n6391 40.1465
R7790 gnd.n6391 gnd.n6390 40.1465
R7791 gnd.n6390 gnd.n962 40.1465
R7792 gnd.n6384 gnd.n962 40.1465
R7793 gnd.n6384 gnd.n6383 40.1465
R7794 gnd.n6383 gnd.n6382 40.1465
R7795 gnd.n6382 gnd.n970 40.1465
R7796 gnd.n6376 gnd.n970 40.1465
R7797 gnd.n2968 gnd.n2967 35.055
R7798 gnd.n2963 gnd.n2962 35.055
R7799 gnd.n4975 gnd.n4974 35.055
R7800 gnd.n4985 gnd.n4971 35.055
R7801 gnd.n1503 gnd.n1399 31.8661
R7802 gnd.n1511 gnd.n1399 31.8661
R7803 gnd.n1519 gnd.n1393 31.8661
R7804 gnd.n1519 gnd.n1387 31.8661
R7805 gnd.n1527 gnd.n1387 31.8661
R7806 gnd.n1527 gnd.n1380 31.8661
R7807 gnd.n1535 gnd.n1380 31.8661
R7808 gnd.n1535 gnd.n1381 31.8661
R7809 gnd.n1747 gnd.n1366 31.8661
R7810 gnd.n6152 gnd.n2380 31.8661
R7811 gnd.n6146 gnd.n2464 31.8661
R7812 gnd.n6146 gnd.n2467 31.8661
R7813 gnd.n6140 gnd.n2467 31.8661
R7814 gnd.n6140 gnd.n2479 31.8661
R7815 gnd.n2738 gnd.n2635 31.8661
R7816 gnd.n4387 gnd.n2752 31.8661
R7817 gnd.n4387 gnd.n2649 31.8661
R7818 gnd.n3929 gnd.n2663 31.8661
R7819 gnd.n4397 gnd.n3929 31.8661
R7820 gnd.n4405 gnd.n3923 31.8661
R7821 gnd.n4405 gnd.n3915 31.8661
R7822 gnd.n4413 gnd.n3915 31.8661
R7823 gnd.n4413 gnd.n3917 31.8661
R7824 gnd.n4421 gnd.n3902 31.8661
R7825 gnd.n4429 gnd.n3902 31.8661
R7826 gnd.n4429 gnd.n3895 31.8661
R7827 gnd.n4437 gnd.n3895 31.8661
R7828 gnd.n4445 gnd.n3888 31.8661
R7829 gnd.n4445 gnd.n3881 31.8661
R7830 gnd.n4453 gnd.n3881 31.8661
R7831 gnd.n4461 gnd.n3874 31.8661
R7832 gnd.n4461 gnd.n3864 31.8661
R7833 gnd.n4480 gnd.n3864 31.8661
R7834 gnd.n4480 gnd.n3866 31.8661
R7835 gnd.n4491 gnd.n2916 31.8661
R7836 gnd.n5187 gnd.n5185 31.8661
R7837 gnd.n5195 gnd.n3500 31.8661
R7838 gnd.n5204 gnd.n3500 31.8661
R7839 gnd.n5204 gnd.n3494 31.8661
R7840 gnd.n5212 gnd.n3494 31.8661
R7841 gnd.n5221 gnd.n3488 31.8661
R7842 gnd.n5221 gnd.n3482 31.8661
R7843 gnd.n5229 gnd.n3482 31.8661
R7844 gnd.n5238 gnd.n3476 31.8661
R7845 gnd.n5238 gnd.n3469 31.8661
R7846 gnd.n5246 gnd.n3469 31.8661
R7847 gnd.n5246 gnd.n3470 31.8661
R7848 gnd.n5255 gnd.n3458 31.8661
R7849 gnd.n5266 gnd.n3458 31.8661
R7850 gnd.n5266 gnd.n3452 31.8661
R7851 gnd.n5275 gnd.n3452 31.8661
R7852 gnd.n5717 gnd.n3088 31.8661
R7853 gnd.n5717 gnd.n3090 31.8661
R7854 gnd.n5296 gnd.n3445 31.8661
R7855 gnd.n3445 gnd.n3157 31.8661
R7856 gnd.n3267 gnd.n3199 31.8661
R7857 gnd.n7375 gnd.n143 31.8661
R7858 gnd.n7369 gnd.n143 31.8661
R7859 gnd.n7369 gnd.n153 31.8661
R7860 gnd.n7363 gnd.n153 31.8661
R7861 gnd.n7357 gnd.n168 31.8661
R7862 gnd.n4172 gnd.n2489 31.5474
R7863 gnd.n7381 gnd.n134 31.5474
R7864 gnd.n5041 gnd.n3530 29.8151
R7865 gnd.n3838 gnd.n3835 29.8151
R7866 gnd.n4453 gnd.t188 27.0862
R7867 gnd.t209 gnd.n3488 27.0862
R7868 gnd.n5911 gnd.n2948 26.4489
R7869 gnd.n4991 gnd.n3532 26.4489
R7870 gnd.n2727 gnd.n2726 25.7944
R7871 gnd.n5653 gnd.n5652 25.7944
R7872 gnd.n1704 gnd.n1703 25.7944
R7873 gnd.n1052 gnd.n1051 25.7944
R7874 gnd.n2734 gnd.n2733 25.7944
R7875 gnd.n3222 gnd.n3221 25.7944
R7876 gnd.n3245 gnd.n3244 25.7944
R7877 gnd.n5533 gnd.n5532 25.7944
R7878 gnd.n176 gnd.n175 25.7944
R7879 gnd.n198 gnd.n197 25.7944
R7880 gnd.n220 gnd.n219 25.7944
R7881 gnd.n7262 gnd.n7261 25.7944
R7882 gnd.n2403 gnd.n2402 25.7944
R7883 gnd.n2425 gnd.n2424 25.7944
R7884 gnd.n2447 gnd.n2446 25.7944
R7885 gnd.n4097 gnd.n4096 25.7944
R7886 gnd.n2804 gnd.n2803 25.7944
R7887 gnd.n2845 gnd.n2844 25.7944
R7888 gnd.n2824 gnd.n2823 25.7944
R7889 gnd.n3150 gnd.n3149 25.7944
R7890 gnd.n1748 gnd.n1356 24.8557
R7891 gnd.n1359 gnd.n1349 24.8557
R7892 gnd.n1778 gnd.n1342 24.8557
R7893 gnd.n1779 gnd.n1331 24.8557
R7894 gnd.n1334 gnd.n1322 24.8557
R7895 gnd.n1800 gnd.n1323 24.8557
R7896 gnd.n1821 gnd.n1820 24.8557
R7897 gnd.n1308 gnd.n1296 24.8557
R7898 gnd.n1831 gnd.n1297 24.8557
R7899 gnd.n1841 gnd.n1279 24.8557
R7900 gnd.n1852 gnd.n1851 24.8557
R7901 gnd.n1862 gnd.n1272 24.8557
R7902 gnd.n1871 gnd.n1264 24.8557
R7903 gnd.n1872 gnd.n1253 24.8557
R7904 gnd.n1883 gnd.n1882 24.8557
R7905 gnd.n1902 gnd.n1239 24.8557
R7906 gnd.n1914 gnd.n1913 24.8557
R7907 gnd.n1575 gnd.n1231 24.8557
R7908 gnd.n1924 gnd.n1221 24.8557
R7909 gnd.n1933 gnd.n1214 24.8557
R7910 gnd.n1944 gnd.n1943 24.8557
R7911 gnd.n1204 gnd.n1195 24.8557
R7912 gnd.n1186 gnd.n1179 24.8557
R7913 gnd.n2014 gnd.n2013 24.8557
R7914 gnd.n2026 gnd.n1168 24.8557
R7915 gnd.n2025 gnd.n1171 24.8557
R7916 gnd.n2038 gnd.n978 24.8557
R7917 gnd.n6374 gnd.n980 24.8557
R7918 gnd.n6368 gnd.n6367 24.8557
R7919 gnd.n6361 gnd.n1001 24.8557
R7920 gnd.n6360 gnd.n1004 24.8557
R7921 gnd.n6354 gnd.n6353 24.8557
R7922 gnd.n1989 gnd.n1018 24.8557
R7923 gnd.n6347 gnd.n1027 24.8557
R7924 gnd.n6340 gnd.n6339 24.8557
R7925 gnd.n4397 gnd.t80 24.537
R7926 gnd.t23 gnd.n3888 24.537
R7927 gnd.n5229 gnd.t162 24.537
R7928 gnd.t54 gnd.n3088 24.537
R7929 gnd.n6376 gnd.n6375 24.0881
R7930 gnd.n6030 gnd.n2663 23.8997
R7931 gnd.n5297 gnd.n3090 23.8997
R7932 gnd.n1769 gnd.t164 23.2624
R7933 gnd.n1759 gnd.t87 22.6251
R7934 gnd.n5841 gnd.n2974 21.6691
R7935 gnd.n4551 gnd.n3739 21.6691
R7936 gnd.n4610 gnd.n3728 21.6691
R7937 gnd.n4654 gnd.n3702 21.6691
R7938 gnd.n4733 gnd.n3663 21.6691
R7939 gnd.n4741 gnd.n4740 21.6691
R7940 gnd.n4759 gnd.n3648 21.6691
R7941 gnd.n4768 gnd.n3643 21.6691
R7942 gnd.n4850 gnd.n4849 21.6691
R7943 gnd.n4873 gnd.n3583 21.6691
R7944 gnd.n4931 gnd.n3560 21.6691
R7945 gnd.n1738 gnd.t160 21.3504
R7946 gnd.n5840 gnd.n2977 21.0318
R7947 gnd.n5834 gnd.n2987 21.0318
R7948 gnd.n4648 gnd.n3708 21.0318
R7949 gnd.n4641 gnd.n3692 21.0318
R7950 gnd.n4788 gnd.n3611 21.0318
R7951 gnd.n4838 gnd.n3607 21.0318
R7952 gnd.n5169 gnd.t97 21.0318
R7953 gnd.n5177 gnd.n3516 21.0318
R7954 gnd.t154 gnd.n989 20.7131
R7955 gnd.n1966 gnd.t27 20.0758
R7956 gnd.n6134 gnd.t241 20.0758
R7957 gnd.n7340 gnd.t215 20.0758
R7958 gnd.n2957 gnd.t122 19.8005
R7959 gnd.n2957 gnd.t147 19.8005
R7960 gnd.n2956 gnd.t78 19.8005
R7961 gnd.n2956 gnd.t128 19.8005
R7962 gnd.n4980 gnd.t145 19.8005
R7963 gnd.n4980 gnd.t98 19.8005
R7964 gnd.n4979 gnd.t41 19.8005
R7965 gnd.n4979 gnd.t113 19.8005
R7966 gnd.n5965 gnd.n2752 19.7572
R7967 gnd.n4524 gnd.n4523 19.7572
R7968 gnd.n4589 gnd.n3699 19.7572
R7969 gnd.n4707 gnd.n3679 19.7572
R7970 gnd.n4818 gnd.n3619 19.7572
R7971 gnd.n4856 gnd.n3603 19.7572
R7972 gnd.n3541 gnd.n3540 19.7572
R7973 gnd.n5649 gnd.n3157 19.7572
R7974 gnd.n2953 gnd.n2952 19.5087
R7975 gnd.n2966 gnd.n2953 19.5087
R7976 gnd.n2964 gnd.n2955 19.5087
R7977 gnd.n4984 gnd.n4978 19.5087
R7978 gnd.t175 gnd.n1228 19.4385
R7979 gnd.n3917 gnd.t0 19.4385
R7980 gnd.n5255 gnd.t21 19.4385
R7981 gnd.n4399 gnd.n3928 19.3944
R7982 gnd.n4399 gnd.n3926 19.3944
R7983 gnd.n4403 gnd.n3926 19.3944
R7984 gnd.n4403 gnd.n3913 19.3944
R7985 gnd.n4415 gnd.n3913 19.3944
R7986 gnd.n4415 gnd.n3911 19.3944
R7987 gnd.n4419 gnd.n3911 19.3944
R7988 gnd.n4419 gnd.n3900 19.3944
R7989 gnd.n4431 gnd.n3900 19.3944
R7990 gnd.n4431 gnd.n3898 19.3944
R7991 gnd.n4435 gnd.n3898 19.3944
R7992 gnd.n4435 gnd.n3886 19.3944
R7993 gnd.n4447 gnd.n3886 19.3944
R7994 gnd.n4447 gnd.n3884 19.3944
R7995 gnd.n4451 gnd.n3884 19.3944
R7996 gnd.n4451 gnd.n3872 19.3944
R7997 gnd.n4463 gnd.n3872 19.3944
R7998 gnd.n4463 gnd.n3869 19.3944
R7999 gnd.n4478 gnd.n3869 19.3944
R8000 gnd.n4478 gnd.n3870 19.3944
R8001 gnd.n4474 gnd.n3870 19.3944
R8002 gnd.n4474 gnd.n4473 19.3944
R8003 gnd.n4473 gnd.n4472 19.3944
R8004 gnd.n4472 gnd.n4469 19.3944
R8005 gnd.n4469 gnd.n2992 19.3944
R8006 gnd.n5832 gnd.n2992 19.3944
R8007 gnd.n5832 gnd.n2993 19.3944
R8008 gnd.n5828 gnd.n2993 19.3944
R8009 gnd.n5828 gnd.n5827 19.3944
R8010 gnd.n5827 gnd.n5826 19.3944
R8011 gnd.n5826 gnd.n2999 19.3944
R8012 gnd.n5822 gnd.n2999 19.3944
R8013 gnd.n5822 gnd.n5821 19.3944
R8014 gnd.n5821 gnd.n5820 19.3944
R8015 gnd.n5820 gnd.n3004 19.3944
R8016 gnd.n5816 gnd.n3004 19.3944
R8017 gnd.n5816 gnd.n5815 19.3944
R8018 gnd.n5815 gnd.n5814 19.3944
R8019 gnd.n5814 gnd.n3009 19.3944
R8020 gnd.n5810 gnd.n3009 19.3944
R8021 gnd.n5810 gnd.n5809 19.3944
R8022 gnd.n5809 gnd.n5808 19.3944
R8023 gnd.n5808 gnd.n3014 19.3944
R8024 gnd.n5804 gnd.n3014 19.3944
R8025 gnd.n5804 gnd.n5803 19.3944
R8026 gnd.n5803 gnd.n5802 19.3944
R8027 gnd.n5802 gnd.n3019 19.3944
R8028 gnd.n5798 gnd.n3019 19.3944
R8029 gnd.n5798 gnd.n5797 19.3944
R8030 gnd.n5797 gnd.n5796 19.3944
R8031 gnd.n5796 gnd.n3024 19.3944
R8032 gnd.n5792 gnd.n3024 19.3944
R8033 gnd.n5792 gnd.n5791 19.3944
R8034 gnd.n5791 gnd.n5790 19.3944
R8035 gnd.n5790 gnd.n3029 19.3944
R8036 gnd.n5786 gnd.n3029 19.3944
R8037 gnd.n5786 gnd.n5785 19.3944
R8038 gnd.n5785 gnd.n5784 19.3944
R8039 gnd.n5784 gnd.n3034 19.3944
R8040 gnd.n5780 gnd.n3034 19.3944
R8041 gnd.n5780 gnd.n5779 19.3944
R8042 gnd.n5779 gnd.n5778 19.3944
R8043 gnd.n5778 gnd.n3039 19.3944
R8044 gnd.n5774 gnd.n3039 19.3944
R8045 gnd.n5774 gnd.n5773 19.3944
R8046 gnd.n5773 gnd.n5772 19.3944
R8047 gnd.n5772 gnd.n3044 19.3944
R8048 gnd.n5768 gnd.n3044 19.3944
R8049 gnd.n5768 gnd.n5767 19.3944
R8050 gnd.n5767 gnd.n5766 19.3944
R8051 gnd.n5766 gnd.n3049 19.3944
R8052 gnd.n5762 gnd.n3049 19.3944
R8053 gnd.n5762 gnd.n5761 19.3944
R8054 gnd.n5761 gnd.n5760 19.3944
R8055 gnd.n5760 gnd.n3054 19.3944
R8056 gnd.n5756 gnd.n3054 19.3944
R8057 gnd.n5756 gnd.n5755 19.3944
R8058 gnd.n5755 gnd.n5754 19.3944
R8059 gnd.n5754 gnd.n3059 19.3944
R8060 gnd.n5750 gnd.n3059 19.3944
R8061 gnd.n5750 gnd.n5749 19.3944
R8062 gnd.n5749 gnd.n5748 19.3944
R8063 gnd.n5748 gnd.n3064 19.3944
R8064 gnd.n5744 gnd.n3064 19.3944
R8065 gnd.n5744 gnd.n5743 19.3944
R8066 gnd.n5743 gnd.n5742 19.3944
R8067 gnd.n5742 gnd.n3069 19.3944
R8068 gnd.n5738 gnd.n3069 19.3944
R8069 gnd.n5738 gnd.n5737 19.3944
R8070 gnd.n5737 gnd.n5736 19.3944
R8071 gnd.n5736 gnd.n3074 19.3944
R8072 gnd.n5732 gnd.n3074 19.3944
R8073 gnd.n5732 gnd.n5731 19.3944
R8074 gnd.n5731 gnd.n5730 19.3944
R8075 gnd.n5730 gnd.n3079 19.3944
R8076 gnd.n5726 gnd.n3079 19.3944
R8077 gnd.n5726 gnd.n5725 19.3944
R8078 gnd.n5725 gnd.n5724 19.3944
R8079 gnd.n5724 gnd.n3084 19.3944
R8080 gnd.n5720 gnd.n3084 19.3944
R8081 gnd.n5720 gnd.n5719 19.3944
R8082 gnd.n2730 gnd.n2646 19.3944
R8083 gnd.n6034 gnd.n2646 19.3944
R8084 gnd.n6034 gnd.n6033 19.3944
R8085 gnd.n6027 gnd.n6026 19.3944
R8086 gnd.n6026 gnd.n2668 19.3944
R8087 gnd.n6022 gnd.n2668 19.3944
R8088 gnd.n6022 gnd.n6021 19.3944
R8089 gnd.n6021 gnd.n6020 19.3944
R8090 gnd.n6020 gnd.n2673 19.3944
R8091 gnd.n6015 gnd.n2673 19.3944
R8092 gnd.n6015 gnd.n6014 19.3944
R8093 gnd.n6014 gnd.n6013 19.3944
R8094 gnd.n6013 gnd.n2679 19.3944
R8095 gnd.n6006 gnd.n2679 19.3944
R8096 gnd.n6006 gnd.n6005 19.3944
R8097 gnd.n6005 gnd.n2691 19.3944
R8098 gnd.n5998 gnd.n2691 19.3944
R8099 gnd.n5998 gnd.n5997 19.3944
R8100 gnd.n5997 gnd.n2699 19.3944
R8101 gnd.n5990 gnd.n2699 19.3944
R8102 gnd.n5990 gnd.n5989 19.3944
R8103 gnd.n5989 gnd.n2709 19.3944
R8104 gnd.n5982 gnd.n2709 19.3944
R8105 gnd.n5982 gnd.n5981 19.3944
R8106 gnd.n5981 gnd.n2717 19.3944
R8107 gnd.n5974 gnd.n2717 19.3944
R8108 gnd.n5974 gnd.n5973 19.3944
R8109 gnd.n5695 gnd.n3110 19.3944
R8110 gnd.n5695 gnd.n5694 19.3944
R8111 gnd.n5694 gnd.n3113 19.3944
R8112 gnd.n5687 gnd.n3113 19.3944
R8113 gnd.n5687 gnd.n5686 19.3944
R8114 gnd.n5686 gnd.n3121 19.3944
R8115 gnd.n5679 gnd.n3121 19.3944
R8116 gnd.n5679 gnd.n5678 19.3944
R8117 gnd.n5678 gnd.n3129 19.3944
R8118 gnd.n5671 gnd.n3129 19.3944
R8119 gnd.n5671 gnd.n5670 19.3944
R8120 gnd.n5670 gnd.n3137 19.3944
R8121 gnd.n5663 gnd.n3137 19.3944
R8122 gnd.n5663 gnd.n5662 19.3944
R8123 gnd.n5662 gnd.n3145 19.3944
R8124 gnd.n5655 gnd.n3145 19.3944
R8125 gnd.n1498 gnd.n1497 19.3944
R8126 gnd.n1497 gnd.n1407 19.3944
R8127 gnd.n1492 gnd.n1407 19.3944
R8128 gnd.n1492 gnd.n1491 19.3944
R8129 gnd.n1491 gnd.n1412 19.3944
R8130 gnd.n1486 gnd.n1412 19.3944
R8131 gnd.n1486 gnd.n1485 19.3944
R8132 gnd.n1485 gnd.n1484 19.3944
R8133 gnd.n1484 gnd.n1418 19.3944
R8134 gnd.n1478 gnd.n1418 19.3944
R8135 gnd.n1478 gnd.n1477 19.3944
R8136 gnd.n1477 gnd.n1476 19.3944
R8137 gnd.n1476 gnd.n1424 19.3944
R8138 gnd.n1470 gnd.n1424 19.3944
R8139 gnd.n1470 gnd.n1469 19.3944
R8140 gnd.n1469 gnd.n1468 19.3944
R8141 gnd.n1468 gnd.n1430 19.3944
R8142 gnd.n1462 gnd.n1430 19.3944
R8143 gnd.n1462 gnd.n1461 19.3944
R8144 gnd.n1461 gnd.n1460 19.3944
R8145 gnd.n1460 gnd.n1436 19.3944
R8146 gnd.n1454 gnd.n1436 19.3944
R8147 gnd.n1452 gnd.n1451 19.3944
R8148 gnd.n1451 gnd.n1446 19.3944
R8149 gnd.n1446 gnd.n1444 19.3944
R8150 gnd.n1146 gnd.n1144 19.3944
R8151 gnd.n1146 gnd.n1070 19.3944
R8152 gnd.n2339 gnd.n1070 19.3944
R8153 gnd.n1087 gnd.n1086 19.3944
R8154 gnd.n1091 gnd.n1086 19.3944
R8155 gnd.n1094 gnd.n1091 19.3944
R8156 gnd.n1097 gnd.n1094 19.3944
R8157 gnd.n1097 gnd.n1083 19.3944
R8158 gnd.n1101 gnd.n1083 19.3944
R8159 gnd.n1104 gnd.n1101 19.3944
R8160 gnd.n1107 gnd.n1104 19.3944
R8161 gnd.n1107 gnd.n1081 19.3944
R8162 gnd.n1111 gnd.n1081 19.3944
R8163 gnd.n1114 gnd.n1111 19.3944
R8164 gnd.n1117 gnd.n1114 19.3944
R8165 gnd.n1117 gnd.n1079 19.3944
R8166 gnd.n1121 gnd.n1079 19.3944
R8167 gnd.n1124 gnd.n1121 19.3944
R8168 gnd.n1127 gnd.n1124 19.3944
R8169 gnd.n1127 gnd.n1077 19.3944
R8170 gnd.n1131 gnd.n1077 19.3944
R8171 gnd.n1134 gnd.n1131 19.3944
R8172 gnd.n1137 gnd.n1134 19.3944
R8173 gnd.n1137 gnd.n1075 19.3944
R8174 gnd.n1141 gnd.n1075 19.3944
R8175 gnd.n1751 gnd.n1750 19.3944
R8176 gnd.n1751 gnd.n1347 19.3944
R8177 gnd.n1771 gnd.n1347 19.3944
R8178 gnd.n1771 gnd.n1339 19.3944
R8179 gnd.n1781 gnd.n1339 19.3944
R8180 gnd.n1782 gnd.n1781 19.3944
R8181 gnd.n1782 gnd.n1320 19.3944
R8182 gnd.n1802 gnd.n1320 19.3944
R8183 gnd.n1802 gnd.n1313 19.3944
R8184 gnd.n1812 gnd.n1313 19.3944
R8185 gnd.n1813 gnd.n1812 19.3944
R8186 gnd.n1813 gnd.n1294 19.3944
R8187 gnd.n1833 gnd.n1294 19.3944
R8188 gnd.n1833 gnd.n1287 19.3944
R8189 gnd.n1843 gnd.n1287 19.3944
R8190 gnd.n1844 gnd.n1843 19.3944
R8191 gnd.n1844 gnd.n1269 19.3944
R8192 gnd.n1864 gnd.n1269 19.3944
R8193 gnd.n1864 gnd.n1261 19.3944
R8194 gnd.n1874 gnd.n1261 19.3944
R8195 gnd.n1875 gnd.n1874 19.3944
R8196 gnd.n1875 gnd.n1244 19.3944
R8197 gnd.n1895 gnd.n1244 19.3944
R8198 gnd.n1895 gnd.n1236 19.3944
R8199 gnd.n1905 gnd.n1236 19.3944
R8200 gnd.n1906 gnd.n1905 19.3944
R8201 gnd.n1906 gnd.n1219 19.3944
R8202 gnd.n1926 gnd.n1219 19.3944
R8203 gnd.n1926 gnd.n1210 19.3944
R8204 gnd.n1936 gnd.n1210 19.3944
R8205 gnd.n1937 gnd.n1936 19.3944
R8206 gnd.n1938 gnd.n1937 19.3944
R8207 gnd.n1938 gnd.n1193 19.3944
R8208 gnd.n1955 gnd.n1193 19.3944
R8209 gnd.n1960 gnd.n1955 19.3944
R8210 gnd.n1960 gnd.n1959 19.3944
R8211 gnd.n1959 gnd.n1957 19.3944
R8212 gnd.n1957 gnd.n1163 19.3944
R8213 gnd.n2036 gnd.n1163 19.3944
R8214 gnd.n2036 gnd.n2035 19.3944
R8215 gnd.n2035 gnd.n1156 19.3944
R8216 gnd.n2048 gnd.n1156 19.3944
R8217 gnd.n2050 gnd.n2048 19.3944
R8218 gnd.n2054 gnd.n2050 19.3944
R8219 gnd.n2055 gnd.n2054 19.3944
R8220 gnd.n2055 gnd.n1153 19.3944
R8221 gnd.n2061 gnd.n1153 19.3944
R8222 gnd.n2319 gnd.n2061 19.3944
R8223 gnd.n2323 gnd.n2319 19.3944
R8224 gnd.n2324 gnd.n2323 19.3944
R8225 gnd.n2329 gnd.n2324 19.3944
R8226 gnd.n2329 gnd.n1049 19.3944
R8227 gnd.n6334 gnd.n1049 19.3944
R8228 gnd.n1734 gnd.n1733 19.3944
R8229 gnd.n1733 gnd.n1732 19.3944
R8230 gnd.n1732 gnd.n1731 19.3944
R8231 gnd.n1731 gnd.n1729 19.3944
R8232 gnd.n1729 gnd.n1726 19.3944
R8233 gnd.n1726 gnd.n1725 19.3944
R8234 gnd.n1725 gnd.n1722 19.3944
R8235 gnd.n1722 gnd.n1721 19.3944
R8236 gnd.n1721 gnd.n1718 19.3944
R8237 gnd.n1718 gnd.n1717 19.3944
R8238 gnd.n1717 gnd.n1714 19.3944
R8239 gnd.n1714 gnd.n1713 19.3944
R8240 gnd.n1713 gnd.n1710 19.3944
R8241 gnd.n1710 gnd.n1709 19.3944
R8242 gnd.n1761 gnd.n1354 19.3944
R8243 gnd.n1761 gnd.n1352 19.3944
R8244 gnd.n1767 gnd.n1352 19.3944
R8245 gnd.n1767 gnd.n1766 19.3944
R8246 gnd.n1766 gnd.n1329 19.3944
R8247 gnd.n1792 gnd.n1329 19.3944
R8248 gnd.n1792 gnd.n1327 19.3944
R8249 gnd.n1798 gnd.n1327 19.3944
R8250 gnd.n1798 gnd.n1797 19.3944
R8251 gnd.n1797 gnd.n1303 19.3944
R8252 gnd.n1823 gnd.n1303 19.3944
R8253 gnd.n1823 gnd.n1301 19.3944
R8254 gnd.n1829 gnd.n1301 19.3944
R8255 gnd.n1829 gnd.n1828 19.3944
R8256 gnd.n1828 gnd.n1277 19.3944
R8257 gnd.n1854 gnd.n1277 19.3944
R8258 gnd.n1854 gnd.n1275 19.3944
R8259 gnd.n1860 gnd.n1275 19.3944
R8260 gnd.n1860 gnd.n1859 19.3944
R8261 gnd.n1859 gnd.n1251 19.3944
R8262 gnd.n1885 gnd.n1251 19.3944
R8263 gnd.n1885 gnd.n1249 19.3944
R8264 gnd.n1891 gnd.n1249 19.3944
R8265 gnd.n1891 gnd.n1890 19.3944
R8266 gnd.n1890 gnd.n1226 19.3944
R8267 gnd.n1916 gnd.n1226 19.3944
R8268 gnd.n1916 gnd.n1224 19.3944
R8269 gnd.n1922 gnd.n1224 19.3944
R8270 gnd.n1922 gnd.n1921 19.3944
R8271 gnd.n1921 gnd.n1199 19.3944
R8272 gnd.n1946 gnd.n1199 19.3944
R8273 gnd.n1946 gnd.n1197 19.3944
R8274 gnd.n1950 gnd.n1197 19.3944
R8275 gnd.n1950 gnd.n1177 19.3944
R8276 gnd.n2016 gnd.n1177 19.3944
R8277 gnd.n2016 gnd.n1175 19.3944
R8278 gnd.n2023 gnd.n1175 19.3944
R8279 gnd.n2023 gnd.n2022 19.3944
R8280 gnd.n2022 gnd.n983 19.3944
R8281 gnd.n6372 gnd.n983 19.3944
R8282 gnd.n6372 gnd.n6371 19.3944
R8283 gnd.n6371 gnd.n6370 19.3944
R8284 gnd.n6370 gnd.n987 19.3944
R8285 gnd.n1007 gnd.n987 19.3944
R8286 gnd.n6358 gnd.n1007 19.3944
R8287 gnd.n6358 gnd.n6357 19.3944
R8288 gnd.n6357 gnd.n6356 19.3944
R8289 gnd.n6356 gnd.n1013 19.3944
R8290 gnd.n1032 gnd.n1013 19.3944
R8291 gnd.n6344 gnd.n1032 19.3944
R8292 gnd.n6344 gnd.n6343 19.3944
R8293 gnd.n6343 gnd.n6342 19.3944
R8294 gnd.n6342 gnd.n1038 19.3944
R8295 gnd.n6321 gnd.n6320 19.3944
R8296 gnd.n6320 gnd.n6286 19.3944
R8297 gnd.n6316 gnd.n6286 19.3944
R8298 gnd.n6316 gnd.n6313 19.3944
R8299 gnd.n6313 gnd.n6310 19.3944
R8300 gnd.n6310 gnd.n6309 19.3944
R8301 gnd.n6309 gnd.n6306 19.3944
R8302 gnd.n6306 gnd.n6305 19.3944
R8303 gnd.n6305 gnd.n6302 19.3944
R8304 gnd.n6302 gnd.n6301 19.3944
R8305 gnd.n6301 gnd.n6298 19.3944
R8306 gnd.n6298 gnd.n6297 19.3944
R8307 gnd.n6297 gnd.n1055 19.3944
R8308 gnd.n6327 gnd.n1055 19.3944
R8309 gnd.n1505 gnd.n1401 19.3944
R8310 gnd.n1509 gnd.n1401 19.3944
R8311 gnd.n1509 gnd.n1391 19.3944
R8312 gnd.n1521 gnd.n1391 19.3944
R8313 gnd.n1521 gnd.n1389 19.3944
R8314 gnd.n1525 gnd.n1389 19.3944
R8315 gnd.n1525 gnd.n1378 19.3944
R8316 gnd.n1537 gnd.n1378 19.3944
R8317 gnd.n1537 gnd.n1376 19.3944
R8318 gnd.n1676 gnd.n1376 19.3944
R8319 gnd.n1676 gnd.n1675 19.3944
R8320 gnd.n1675 gnd.n1674 19.3944
R8321 gnd.n1674 gnd.n1673 19.3944
R8322 gnd.n1673 gnd.n1671 19.3944
R8323 gnd.n1671 gnd.n1670 19.3944
R8324 gnd.n1670 gnd.n1666 19.3944
R8325 gnd.n1666 gnd.n1665 19.3944
R8326 gnd.n1665 gnd.n1664 19.3944
R8327 gnd.n1664 gnd.n1662 19.3944
R8328 gnd.n1662 gnd.n1661 19.3944
R8329 gnd.n1661 gnd.n1658 19.3944
R8330 gnd.n1658 gnd.n1657 19.3944
R8331 gnd.n1657 gnd.n1656 19.3944
R8332 gnd.n1656 gnd.n1654 19.3944
R8333 gnd.n1654 gnd.n1653 19.3944
R8334 gnd.n1653 gnd.n1650 19.3944
R8335 gnd.n1650 gnd.n1649 19.3944
R8336 gnd.n1649 gnd.n1648 19.3944
R8337 gnd.n1648 gnd.n1646 19.3944
R8338 gnd.n1594 gnd.n1559 19.3944
R8339 gnd.n1591 gnd.n1590 19.3944
R8340 gnd.n1587 gnd.n1586 19.3944
R8341 gnd.n1582 gnd.n1581 19.3944
R8342 gnd.n1581 gnd.n1580 19.3944
R8343 gnd.n1580 gnd.n1578 19.3944
R8344 gnd.n1578 gnd.n1577 19.3944
R8345 gnd.n1577 gnd.n1573 19.3944
R8346 gnd.n1573 gnd.n1572 19.3944
R8347 gnd.n1572 gnd.n1571 19.3944
R8348 gnd.n1571 gnd.n1569 19.3944
R8349 gnd.n1569 gnd.n1184 19.3944
R8350 gnd.n1968 gnd.n1184 19.3944
R8351 gnd.n1968 gnd.n1182 19.3944
R8352 gnd.n2011 gnd.n1182 19.3944
R8353 gnd.n2011 gnd.n2010 19.3944
R8354 gnd.n2010 gnd.n2009 19.3944
R8355 gnd.n2009 gnd.n2007 19.3944
R8356 gnd.n2007 gnd.n2006 19.3944
R8357 gnd.n2006 gnd.n1976 19.3944
R8358 gnd.n2002 gnd.n1976 19.3944
R8359 gnd.n2002 gnd.n2001 19.3944
R8360 gnd.n2001 gnd.n2000 19.3944
R8361 gnd.n2000 gnd.n1997 19.3944
R8362 gnd.n1997 gnd.n1996 19.3944
R8363 gnd.n1996 gnd.n1993 19.3944
R8364 gnd.n1993 gnd.n1992 19.3944
R8365 gnd.n1992 gnd.n1991 19.3944
R8366 gnd.n1991 gnd.n1988 19.3944
R8367 gnd.n1988 gnd.n1150 19.3944
R8368 gnd.n2335 gnd.n1150 19.3944
R8369 gnd.n2336 gnd.n2335 19.3944
R8370 gnd.n1501 gnd.n1397 19.3944
R8371 gnd.n1513 gnd.n1397 19.3944
R8372 gnd.n1513 gnd.n1395 19.3944
R8373 gnd.n1517 gnd.n1395 19.3944
R8374 gnd.n1517 gnd.n1385 19.3944
R8375 gnd.n1529 gnd.n1385 19.3944
R8376 gnd.n1529 gnd.n1383 19.3944
R8377 gnd.n1533 gnd.n1383 19.3944
R8378 gnd.n1533 gnd.n1372 19.3944
R8379 gnd.n1740 gnd.n1372 19.3944
R8380 gnd.n1740 gnd.n1369 19.3944
R8381 gnd.n1745 gnd.n1369 19.3944
R8382 gnd.n1745 gnd.n1362 19.3944
R8383 gnd.n1756 gnd.n1362 19.3944
R8384 gnd.n1756 gnd.n1755 19.3944
R8385 gnd.n1755 gnd.n1345 19.3944
R8386 gnd.n1776 gnd.n1345 19.3944
R8387 gnd.n1776 gnd.n1337 19.3944
R8388 gnd.n1787 gnd.n1337 19.3944
R8389 gnd.n1787 gnd.n1786 19.3944
R8390 gnd.n1786 gnd.n1318 19.3944
R8391 gnd.n1807 gnd.n1318 19.3944
R8392 gnd.n1807 gnd.n1311 19.3944
R8393 gnd.n1818 gnd.n1311 19.3944
R8394 gnd.n1818 gnd.n1817 19.3944
R8395 gnd.n1817 gnd.n1292 19.3944
R8396 gnd.n1838 gnd.n1292 19.3944
R8397 gnd.n1838 gnd.n1285 19.3944
R8398 gnd.n1849 gnd.n1285 19.3944
R8399 gnd.n1849 gnd.n1848 19.3944
R8400 gnd.n1848 gnd.n1267 19.3944
R8401 gnd.n1869 gnd.n1267 19.3944
R8402 gnd.n1869 gnd.n1259 19.3944
R8403 gnd.n1880 gnd.n1259 19.3944
R8404 gnd.n1880 gnd.n1879 19.3944
R8405 gnd.n1879 gnd.n1242 19.3944
R8406 gnd.n1900 gnd.n1242 19.3944
R8407 gnd.n1900 gnd.n1234 19.3944
R8408 gnd.n1911 gnd.n1234 19.3944
R8409 gnd.n1911 gnd.n1910 19.3944
R8410 gnd.n1910 gnd.n1217 19.3944
R8411 gnd.n1931 gnd.n1217 19.3944
R8412 gnd.n1931 gnd.n1206 19.3944
R8413 gnd.n1941 gnd.n1206 19.3944
R8414 gnd.n1941 gnd.n1189 19.3944
R8415 gnd.n1964 gnd.n1189 19.3944
R8416 gnd.n1964 gnd.n1963 19.3944
R8417 gnd.n1963 gnd.n1165 19.3944
R8418 gnd.n2028 gnd.n1165 19.3944
R8419 gnd.n2029 gnd.n2028 19.3944
R8420 gnd.n2029 gnd.n1160 19.3944
R8421 gnd.n1160 gnd.n1158 19.3944
R8422 gnd.n2043 gnd.n1158 19.3944
R8423 gnd.n2043 gnd.n995 19.3944
R8424 gnd.n6365 gnd.n995 19.3944
R8425 gnd.n6365 gnd.n6364 19.3944
R8426 gnd.n6364 gnd.n6363 19.3944
R8427 gnd.n6363 gnd.n999 19.3944
R8428 gnd.n1021 gnd.n999 19.3944
R8429 gnd.n6351 gnd.n1021 19.3944
R8430 gnd.n6351 gnd.n6350 19.3944
R8431 gnd.n6350 gnd.n6349 19.3944
R8432 gnd.n6349 gnd.n1025 19.3944
R8433 gnd.n1046 gnd.n1025 19.3944
R8434 gnd.n6337 gnd.n1046 19.3944
R8435 gnd.n6010 gnd.n2682 19.3944
R8436 gnd.n6010 gnd.n6009 19.3944
R8437 gnd.n6009 gnd.n2685 19.3944
R8438 gnd.n6002 gnd.n2685 19.3944
R8439 gnd.n6002 gnd.n6001 19.3944
R8440 gnd.n6001 gnd.n2695 19.3944
R8441 gnd.n5994 gnd.n2695 19.3944
R8442 gnd.n5994 gnd.n5993 19.3944
R8443 gnd.n5993 gnd.n2703 19.3944
R8444 gnd.n5986 gnd.n2703 19.3944
R8445 gnd.n5986 gnd.n5985 19.3944
R8446 gnd.n5985 gnd.n2713 19.3944
R8447 gnd.n5978 gnd.n2713 19.3944
R8448 gnd.n5978 gnd.n5977 19.3944
R8449 gnd.n5977 gnd.n2721 19.3944
R8450 gnd.n5970 gnd.n2721 19.3944
R8451 gnd.n7001 gnd.n534 19.3944
R8452 gnd.n7007 gnd.n534 19.3944
R8453 gnd.n7007 gnd.n532 19.3944
R8454 gnd.n7011 gnd.n532 19.3944
R8455 gnd.n7011 gnd.n528 19.3944
R8456 gnd.n7017 gnd.n528 19.3944
R8457 gnd.n7017 gnd.n526 19.3944
R8458 gnd.n7021 gnd.n526 19.3944
R8459 gnd.n7021 gnd.n522 19.3944
R8460 gnd.n7027 gnd.n522 19.3944
R8461 gnd.n7027 gnd.n520 19.3944
R8462 gnd.n7031 gnd.n520 19.3944
R8463 gnd.n7031 gnd.n516 19.3944
R8464 gnd.n7037 gnd.n516 19.3944
R8465 gnd.n7037 gnd.n514 19.3944
R8466 gnd.n7041 gnd.n514 19.3944
R8467 gnd.n7041 gnd.n510 19.3944
R8468 gnd.n7047 gnd.n510 19.3944
R8469 gnd.n7047 gnd.n508 19.3944
R8470 gnd.n7051 gnd.n508 19.3944
R8471 gnd.n7051 gnd.n504 19.3944
R8472 gnd.n7057 gnd.n504 19.3944
R8473 gnd.n7057 gnd.n502 19.3944
R8474 gnd.n7061 gnd.n502 19.3944
R8475 gnd.n7061 gnd.n498 19.3944
R8476 gnd.n7067 gnd.n498 19.3944
R8477 gnd.n7067 gnd.n496 19.3944
R8478 gnd.n7071 gnd.n496 19.3944
R8479 gnd.n7071 gnd.n492 19.3944
R8480 gnd.n7077 gnd.n492 19.3944
R8481 gnd.n7077 gnd.n490 19.3944
R8482 gnd.n7081 gnd.n490 19.3944
R8483 gnd.n7081 gnd.n486 19.3944
R8484 gnd.n7087 gnd.n486 19.3944
R8485 gnd.n7087 gnd.n484 19.3944
R8486 gnd.n7091 gnd.n484 19.3944
R8487 gnd.n7091 gnd.n480 19.3944
R8488 gnd.n7097 gnd.n480 19.3944
R8489 gnd.n7097 gnd.n478 19.3944
R8490 gnd.n7101 gnd.n478 19.3944
R8491 gnd.n7101 gnd.n474 19.3944
R8492 gnd.n7107 gnd.n474 19.3944
R8493 gnd.n7107 gnd.n472 19.3944
R8494 gnd.n7111 gnd.n472 19.3944
R8495 gnd.n7111 gnd.n468 19.3944
R8496 gnd.n7117 gnd.n468 19.3944
R8497 gnd.n7117 gnd.n466 19.3944
R8498 gnd.n7121 gnd.n466 19.3944
R8499 gnd.n7121 gnd.n462 19.3944
R8500 gnd.n7127 gnd.n462 19.3944
R8501 gnd.n7127 gnd.n460 19.3944
R8502 gnd.n7131 gnd.n460 19.3944
R8503 gnd.n7131 gnd.n456 19.3944
R8504 gnd.n7137 gnd.n456 19.3944
R8505 gnd.n7137 gnd.n454 19.3944
R8506 gnd.n7141 gnd.n454 19.3944
R8507 gnd.n7141 gnd.n450 19.3944
R8508 gnd.n7147 gnd.n450 19.3944
R8509 gnd.n7147 gnd.n448 19.3944
R8510 gnd.n7151 gnd.n448 19.3944
R8511 gnd.n7151 gnd.n444 19.3944
R8512 gnd.n7157 gnd.n444 19.3944
R8513 gnd.n7157 gnd.n442 19.3944
R8514 gnd.n7161 gnd.n442 19.3944
R8515 gnd.n7161 gnd.n438 19.3944
R8516 gnd.n7167 gnd.n438 19.3944
R8517 gnd.n7167 gnd.n436 19.3944
R8518 gnd.n7171 gnd.n436 19.3944
R8519 gnd.n7171 gnd.n432 19.3944
R8520 gnd.n7177 gnd.n432 19.3944
R8521 gnd.n7177 gnd.n430 19.3944
R8522 gnd.n7181 gnd.n430 19.3944
R8523 gnd.n7181 gnd.n426 19.3944
R8524 gnd.n7187 gnd.n426 19.3944
R8525 gnd.n7187 gnd.n424 19.3944
R8526 gnd.n7191 gnd.n424 19.3944
R8527 gnd.n7191 gnd.n420 19.3944
R8528 gnd.n7197 gnd.n420 19.3944
R8529 gnd.n7197 gnd.n418 19.3944
R8530 gnd.n7201 gnd.n418 19.3944
R8531 gnd.n7201 gnd.n414 19.3944
R8532 gnd.n7208 gnd.n414 19.3944
R8533 gnd.n7208 gnd.n412 19.3944
R8534 gnd.n7212 gnd.n412 19.3944
R8535 gnd.n6546 gnd.n807 19.3944
R8536 gnd.n6550 gnd.n807 19.3944
R8537 gnd.n6550 gnd.n803 19.3944
R8538 gnd.n6556 gnd.n803 19.3944
R8539 gnd.n6556 gnd.n801 19.3944
R8540 gnd.n6560 gnd.n801 19.3944
R8541 gnd.n6560 gnd.n797 19.3944
R8542 gnd.n6566 gnd.n797 19.3944
R8543 gnd.n6566 gnd.n795 19.3944
R8544 gnd.n6570 gnd.n795 19.3944
R8545 gnd.n6570 gnd.n791 19.3944
R8546 gnd.n6576 gnd.n791 19.3944
R8547 gnd.n6576 gnd.n789 19.3944
R8548 gnd.n6580 gnd.n789 19.3944
R8549 gnd.n6580 gnd.n785 19.3944
R8550 gnd.n6586 gnd.n785 19.3944
R8551 gnd.n6586 gnd.n783 19.3944
R8552 gnd.n6590 gnd.n783 19.3944
R8553 gnd.n6590 gnd.n779 19.3944
R8554 gnd.n6596 gnd.n779 19.3944
R8555 gnd.n6596 gnd.n777 19.3944
R8556 gnd.n6600 gnd.n777 19.3944
R8557 gnd.n6600 gnd.n773 19.3944
R8558 gnd.n6606 gnd.n773 19.3944
R8559 gnd.n6606 gnd.n771 19.3944
R8560 gnd.n6610 gnd.n771 19.3944
R8561 gnd.n6610 gnd.n767 19.3944
R8562 gnd.n6616 gnd.n767 19.3944
R8563 gnd.n6616 gnd.n765 19.3944
R8564 gnd.n6620 gnd.n765 19.3944
R8565 gnd.n6620 gnd.n761 19.3944
R8566 gnd.n6626 gnd.n761 19.3944
R8567 gnd.n6626 gnd.n759 19.3944
R8568 gnd.n6630 gnd.n759 19.3944
R8569 gnd.n6630 gnd.n755 19.3944
R8570 gnd.n6636 gnd.n755 19.3944
R8571 gnd.n6636 gnd.n753 19.3944
R8572 gnd.n6640 gnd.n753 19.3944
R8573 gnd.n6640 gnd.n749 19.3944
R8574 gnd.n6646 gnd.n749 19.3944
R8575 gnd.n6646 gnd.n747 19.3944
R8576 gnd.n6650 gnd.n747 19.3944
R8577 gnd.n6650 gnd.n743 19.3944
R8578 gnd.n6656 gnd.n743 19.3944
R8579 gnd.n6656 gnd.n741 19.3944
R8580 gnd.n6660 gnd.n741 19.3944
R8581 gnd.n6660 gnd.n737 19.3944
R8582 gnd.n6666 gnd.n737 19.3944
R8583 gnd.n6666 gnd.n735 19.3944
R8584 gnd.n6670 gnd.n735 19.3944
R8585 gnd.n6670 gnd.n731 19.3944
R8586 gnd.n6676 gnd.n731 19.3944
R8587 gnd.n6676 gnd.n729 19.3944
R8588 gnd.n6680 gnd.n729 19.3944
R8589 gnd.n6680 gnd.n725 19.3944
R8590 gnd.n6686 gnd.n725 19.3944
R8591 gnd.n6686 gnd.n723 19.3944
R8592 gnd.n6690 gnd.n723 19.3944
R8593 gnd.n6690 gnd.n719 19.3944
R8594 gnd.n6696 gnd.n719 19.3944
R8595 gnd.n6696 gnd.n717 19.3944
R8596 gnd.n6700 gnd.n717 19.3944
R8597 gnd.n6700 gnd.n713 19.3944
R8598 gnd.n6706 gnd.n713 19.3944
R8599 gnd.n6706 gnd.n711 19.3944
R8600 gnd.n6710 gnd.n711 19.3944
R8601 gnd.n6710 gnd.n707 19.3944
R8602 gnd.n6716 gnd.n707 19.3944
R8603 gnd.n6716 gnd.n705 19.3944
R8604 gnd.n6720 gnd.n705 19.3944
R8605 gnd.n6720 gnd.n701 19.3944
R8606 gnd.n6726 gnd.n701 19.3944
R8607 gnd.n6726 gnd.n699 19.3944
R8608 gnd.n6730 gnd.n699 19.3944
R8609 gnd.n6730 gnd.n695 19.3944
R8610 gnd.n6736 gnd.n695 19.3944
R8611 gnd.n6736 gnd.n693 19.3944
R8612 gnd.n6740 gnd.n693 19.3944
R8613 gnd.n6740 gnd.n689 19.3944
R8614 gnd.n6746 gnd.n689 19.3944
R8615 gnd.n6746 gnd.n687 19.3944
R8616 gnd.n6750 gnd.n687 19.3944
R8617 gnd.n6750 gnd.n683 19.3944
R8618 gnd.n6756 gnd.n683 19.3944
R8619 gnd.n6756 gnd.n681 19.3944
R8620 gnd.n6760 gnd.n681 19.3944
R8621 gnd.n6760 gnd.n677 19.3944
R8622 gnd.n6766 gnd.n677 19.3944
R8623 gnd.n6766 gnd.n675 19.3944
R8624 gnd.n6770 gnd.n675 19.3944
R8625 gnd.n6770 gnd.n671 19.3944
R8626 gnd.n6776 gnd.n671 19.3944
R8627 gnd.n6776 gnd.n669 19.3944
R8628 gnd.n6780 gnd.n669 19.3944
R8629 gnd.n6780 gnd.n665 19.3944
R8630 gnd.n6786 gnd.n665 19.3944
R8631 gnd.n6786 gnd.n663 19.3944
R8632 gnd.n6790 gnd.n663 19.3944
R8633 gnd.n6790 gnd.n659 19.3944
R8634 gnd.n6796 gnd.n659 19.3944
R8635 gnd.n6796 gnd.n657 19.3944
R8636 gnd.n6800 gnd.n657 19.3944
R8637 gnd.n6800 gnd.n653 19.3944
R8638 gnd.n6806 gnd.n653 19.3944
R8639 gnd.n6806 gnd.n651 19.3944
R8640 gnd.n6810 gnd.n651 19.3944
R8641 gnd.n6810 gnd.n647 19.3944
R8642 gnd.n6816 gnd.n647 19.3944
R8643 gnd.n6816 gnd.n645 19.3944
R8644 gnd.n6820 gnd.n645 19.3944
R8645 gnd.n6820 gnd.n641 19.3944
R8646 gnd.n6826 gnd.n641 19.3944
R8647 gnd.n6826 gnd.n639 19.3944
R8648 gnd.n6830 gnd.n639 19.3944
R8649 gnd.n6830 gnd.n635 19.3944
R8650 gnd.n6836 gnd.n635 19.3944
R8651 gnd.n6836 gnd.n633 19.3944
R8652 gnd.n6840 gnd.n633 19.3944
R8653 gnd.n6840 gnd.n629 19.3944
R8654 gnd.n6846 gnd.n629 19.3944
R8655 gnd.n6846 gnd.n627 19.3944
R8656 gnd.n6850 gnd.n627 19.3944
R8657 gnd.n6850 gnd.n623 19.3944
R8658 gnd.n6856 gnd.n623 19.3944
R8659 gnd.n6856 gnd.n621 19.3944
R8660 gnd.n6860 gnd.n621 19.3944
R8661 gnd.n6860 gnd.n617 19.3944
R8662 gnd.n6866 gnd.n617 19.3944
R8663 gnd.n6866 gnd.n615 19.3944
R8664 gnd.n6870 gnd.n615 19.3944
R8665 gnd.n6870 gnd.n611 19.3944
R8666 gnd.n6876 gnd.n611 19.3944
R8667 gnd.n6876 gnd.n609 19.3944
R8668 gnd.n6880 gnd.n609 19.3944
R8669 gnd.n6880 gnd.n605 19.3944
R8670 gnd.n6886 gnd.n605 19.3944
R8671 gnd.n6886 gnd.n603 19.3944
R8672 gnd.n6890 gnd.n603 19.3944
R8673 gnd.n6890 gnd.n599 19.3944
R8674 gnd.n6896 gnd.n599 19.3944
R8675 gnd.n6896 gnd.n597 19.3944
R8676 gnd.n6900 gnd.n597 19.3944
R8677 gnd.n6900 gnd.n593 19.3944
R8678 gnd.n6906 gnd.n593 19.3944
R8679 gnd.n6906 gnd.n591 19.3944
R8680 gnd.n6910 gnd.n591 19.3944
R8681 gnd.n6910 gnd.n587 19.3944
R8682 gnd.n6916 gnd.n587 19.3944
R8683 gnd.n6916 gnd.n585 19.3944
R8684 gnd.n6920 gnd.n585 19.3944
R8685 gnd.n6920 gnd.n581 19.3944
R8686 gnd.n6926 gnd.n581 19.3944
R8687 gnd.n6926 gnd.n579 19.3944
R8688 gnd.n6930 gnd.n579 19.3944
R8689 gnd.n6930 gnd.n575 19.3944
R8690 gnd.n6936 gnd.n575 19.3944
R8691 gnd.n6936 gnd.n573 19.3944
R8692 gnd.n6940 gnd.n573 19.3944
R8693 gnd.n6940 gnd.n569 19.3944
R8694 gnd.n6946 gnd.n569 19.3944
R8695 gnd.n6946 gnd.n567 19.3944
R8696 gnd.n6950 gnd.n567 19.3944
R8697 gnd.n6950 gnd.n563 19.3944
R8698 gnd.n6956 gnd.n563 19.3944
R8699 gnd.n6956 gnd.n561 19.3944
R8700 gnd.n6960 gnd.n561 19.3944
R8701 gnd.n6960 gnd.n557 19.3944
R8702 gnd.n6966 gnd.n557 19.3944
R8703 gnd.n6966 gnd.n555 19.3944
R8704 gnd.n6970 gnd.n555 19.3944
R8705 gnd.n6970 gnd.n551 19.3944
R8706 gnd.n6976 gnd.n551 19.3944
R8707 gnd.n6976 gnd.n549 19.3944
R8708 gnd.n6980 gnd.n549 19.3944
R8709 gnd.n6980 gnd.n545 19.3944
R8710 gnd.n6986 gnd.n545 19.3944
R8711 gnd.n6986 gnd.n543 19.3944
R8712 gnd.n6991 gnd.n543 19.3944
R8713 gnd.n6991 gnd.n539 19.3944
R8714 gnd.n6997 gnd.n539 19.3944
R8715 gnd.n6998 gnd.n6997 19.3944
R8716 gnd.n5646 gnd.n5645 19.3944
R8717 gnd.n5645 gnd.n5644 19.3944
R8718 gnd.n5644 gnd.n5643 19.3944
R8719 gnd.n5643 gnd.n5641 19.3944
R8720 gnd.n5641 gnd.n5638 19.3944
R8721 gnd.n5638 gnd.n5637 19.3944
R8722 gnd.n5637 gnd.n5634 19.3944
R8723 gnd.n5634 gnd.n5633 19.3944
R8724 gnd.n5633 gnd.n5630 19.3944
R8725 gnd.n5630 gnd.n5629 19.3944
R8726 gnd.n5629 gnd.n5626 19.3944
R8727 gnd.n5626 gnd.n5625 19.3944
R8728 gnd.n5625 gnd.n5622 19.3944
R8729 gnd.n5622 gnd.n5621 19.3944
R8730 gnd.n5621 gnd.n5618 19.3944
R8731 gnd.n5618 gnd.n5617 19.3944
R8732 gnd.n5617 gnd.n5614 19.3944
R8733 gnd.n5612 gnd.n5609 19.3944
R8734 gnd.n5609 gnd.n5608 19.3944
R8735 gnd.n5608 gnd.n5605 19.3944
R8736 gnd.n5605 gnd.n5604 19.3944
R8737 gnd.n5604 gnd.n5601 19.3944
R8738 gnd.n5601 gnd.n5600 19.3944
R8739 gnd.n5600 gnd.n5597 19.3944
R8740 gnd.n5595 gnd.n5592 19.3944
R8741 gnd.n5592 gnd.n5591 19.3944
R8742 gnd.n5591 gnd.n5588 19.3944
R8743 gnd.n5588 gnd.n5587 19.3944
R8744 gnd.n5587 gnd.n5584 19.3944
R8745 gnd.n5584 gnd.n5583 19.3944
R8746 gnd.n5583 gnd.n5580 19.3944
R8747 gnd.n5580 gnd.n5579 19.3944
R8748 gnd.n5575 gnd.n5572 19.3944
R8749 gnd.n5572 gnd.n5571 19.3944
R8750 gnd.n5571 gnd.n5568 19.3944
R8751 gnd.n5568 gnd.n5567 19.3944
R8752 gnd.n5567 gnd.n5564 19.3944
R8753 gnd.n5564 gnd.n5563 19.3944
R8754 gnd.n5563 gnd.n5560 19.3944
R8755 gnd.n5560 gnd.n5559 19.3944
R8756 gnd.n5559 gnd.n5556 19.3944
R8757 gnd.n5556 gnd.n5555 19.3944
R8758 gnd.n5555 gnd.n5552 19.3944
R8759 gnd.n5552 gnd.n5551 19.3944
R8760 gnd.n5551 gnd.n5548 19.3944
R8761 gnd.n5548 gnd.n5547 19.3944
R8762 gnd.n5547 gnd.n5544 19.3944
R8763 gnd.n5544 gnd.n5543 19.3944
R8764 gnd.n5543 gnd.n5540 19.3944
R8765 gnd.n5540 gnd.n5539 19.3944
R8766 gnd.n5523 gnd.n3266 19.3944
R8767 gnd.n5523 gnd.n5522 19.3944
R8768 gnd.n5522 gnd.n3275 19.3944
R8769 gnd.n5312 gnd.n3275 19.3944
R8770 gnd.n5315 gnd.n5312 19.3944
R8771 gnd.n5316 gnd.n5315 19.3944
R8772 gnd.n5321 gnd.n5316 19.3944
R8773 gnd.n5322 gnd.n5321 19.3944
R8774 gnd.n5326 gnd.n5322 19.3944
R8775 gnd.n5326 gnd.n5325 19.3944
R8776 gnd.n5325 gnd.n5324 19.3944
R8777 gnd.n5324 gnd.n3397 19.3944
R8778 gnd.n5398 gnd.n3397 19.3944
R8779 gnd.n5399 gnd.n5398 19.3944
R8780 gnd.n5401 gnd.n5399 19.3944
R8781 gnd.n5401 gnd.n3391 19.3944
R8782 gnd.n5417 gnd.n3391 19.3944
R8783 gnd.n5418 gnd.n5417 19.3944
R8784 gnd.n5419 gnd.n5418 19.3944
R8785 gnd.n5419 gnd.n3386 19.3944
R8786 gnd.n5427 gnd.n3386 19.3944
R8787 gnd.n5428 gnd.n5427 19.3944
R8788 gnd.n5429 gnd.n5428 19.3944
R8789 gnd.n5430 gnd.n5429 19.3944
R8790 gnd.n5432 gnd.n5430 19.3944
R8791 gnd.n5432 gnd.n396 19.3944
R8792 gnd.n7228 gnd.n396 19.3944
R8793 gnd.n7229 gnd.n7228 19.3944
R8794 gnd.n7231 gnd.n7229 19.3944
R8795 gnd.n7231 gnd.n391 19.3944
R8796 gnd.n7243 gnd.n391 19.3944
R8797 gnd.n7244 gnd.n7243 19.3944
R8798 gnd.n7246 gnd.n7244 19.3944
R8799 gnd.n7246 gnd.n387 19.3944
R8800 gnd.n7342 gnd.n387 19.3944
R8801 gnd.n7343 gnd.n7342 19.3944
R8802 gnd.n7346 gnd.n7343 19.3944
R8803 gnd.n7347 gnd.n7346 19.3944
R8804 gnd.n7349 gnd.n7347 19.3944
R8805 gnd.n7350 gnd.n7349 19.3944
R8806 gnd.n7352 gnd.n7350 19.3944
R8807 gnd.n7353 gnd.n7352 19.3944
R8808 gnd.n5526 gnd.n5525 19.3944
R8809 gnd.n5525 gnd.n3273 19.3944
R8810 gnd.n3297 gnd.n3273 19.3944
R8811 gnd.n5512 gnd.n3297 19.3944
R8812 gnd.n5512 gnd.n5511 19.3944
R8813 gnd.n5511 gnd.n5510 19.3944
R8814 gnd.n5510 gnd.n3302 19.3944
R8815 gnd.n5500 gnd.n3302 19.3944
R8816 gnd.n5500 gnd.n5499 19.3944
R8817 gnd.n5499 gnd.n5498 19.3944
R8818 gnd.n5498 gnd.n3322 19.3944
R8819 gnd.n5488 gnd.n3322 19.3944
R8820 gnd.n5488 gnd.n5487 19.3944
R8821 gnd.n5487 gnd.n5486 19.3944
R8822 gnd.n5486 gnd.n3342 19.3944
R8823 gnd.n5476 gnd.n3342 19.3944
R8824 gnd.n5476 gnd.n5475 19.3944
R8825 gnd.n5475 gnd.n5474 19.3944
R8826 gnd.n5474 gnd.n3359 19.3944
R8827 gnd.n5422 gnd.n3359 19.3944
R8828 gnd.n5422 gnd.n3381 19.3944
R8829 gnd.n5456 gnd.n3381 19.3944
R8830 gnd.n5456 gnd.n5455 19.3944
R8831 gnd.n5455 gnd.n5454 19.3944
R8832 gnd.n5454 gnd.n96 19.3944
R8833 gnd.n7403 gnd.n96 19.3944
R8834 gnd.n7403 gnd.n7402 19.3944
R8835 gnd.n7402 gnd.n7401 19.3944
R8836 gnd.n7401 gnd.n100 19.3944
R8837 gnd.n7391 gnd.n100 19.3944
R8838 gnd.n7391 gnd.n7390 19.3944
R8839 gnd.n7390 gnd.n7389 19.3944
R8840 gnd.n7389 gnd.n118 19.3944
R8841 gnd.n7379 gnd.n118 19.3944
R8842 gnd.n7379 gnd.n7378 19.3944
R8843 gnd.n7378 gnd.n7377 19.3944
R8844 gnd.n7377 gnd.n139 19.3944
R8845 gnd.n7367 gnd.n139 19.3944
R8846 gnd.n7367 gnd.n7366 19.3944
R8847 gnd.n7366 gnd.n7365 19.3944
R8848 gnd.n7365 gnd.n158 19.3944
R8849 gnd.n7355 gnd.n158 19.3944
R8850 gnd.n335 gnd.n195 19.3944
R8851 gnd.n339 gnd.n195 19.3944
R8852 gnd.n339 gnd.n193 19.3944
R8853 gnd.n345 gnd.n193 19.3944
R8854 gnd.n345 gnd.n191 19.3944
R8855 gnd.n349 gnd.n191 19.3944
R8856 gnd.n349 gnd.n189 19.3944
R8857 gnd.n355 gnd.n189 19.3944
R8858 gnd.n355 gnd.n187 19.3944
R8859 gnd.n359 gnd.n187 19.3944
R8860 gnd.n359 gnd.n185 19.3944
R8861 gnd.n365 gnd.n185 19.3944
R8862 gnd.n365 gnd.n183 19.3944
R8863 gnd.n369 gnd.n183 19.3944
R8864 gnd.n369 gnd.n181 19.3944
R8865 gnd.n375 gnd.n181 19.3944
R8866 gnd.n375 gnd.n179 19.3944
R8867 gnd.n379 gnd.n179 19.3944
R8868 gnd.n285 gnd.n217 19.3944
R8869 gnd.n289 gnd.n217 19.3944
R8870 gnd.n289 gnd.n215 19.3944
R8871 gnd.n295 gnd.n215 19.3944
R8872 gnd.n295 gnd.n213 19.3944
R8873 gnd.n299 gnd.n213 19.3944
R8874 gnd.n299 gnd.n211 19.3944
R8875 gnd.n305 gnd.n211 19.3944
R8876 gnd.n305 gnd.n209 19.3944
R8877 gnd.n309 gnd.n209 19.3944
R8878 gnd.n309 gnd.n207 19.3944
R8879 gnd.n315 gnd.n207 19.3944
R8880 gnd.n315 gnd.n205 19.3944
R8881 gnd.n319 gnd.n205 19.3944
R8882 gnd.n319 gnd.n203 19.3944
R8883 gnd.n325 gnd.n203 19.3944
R8884 gnd.n325 gnd.n201 19.3944
R8885 gnd.n329 gnd.n201 19.3944
R8886 gnd.n239 gnd.n238 19.3944
R8887 gnd.n244 gnd.n239 19.3944
R8888 gnd.n244 gnd.n235 19.3944
R8889 gnd.n248 gnd.n235 19.3944
R8890 gnd.n248 gnd.n233 19.3944
R8891 gnd.n254 gnd.n233 19.3944
R8892 gnd.n254 gnd.n231 19.3944
R8893 gnd.n258 gnd.n231 19.3944
R8894 gnd.n258 gnd.n229 19.3944
R8895 gnd.n264 gnd.n229 19.3944
R8896 gnd.n264 gnd.n227 19.3944
R8897 gnd.n268 gnd.n227 19.3944
R8898 gnd.n268 gnd.n225 19.3944
R8899 gnd.n275 gnd.n225 19.3944
R8900 gnd.n275 gnd.n223 19.3944
R8901 gnd.n279 gnd.n223 19.3944
R8902 gnd.n280 gnd.n279 19.3944
R8903 gnd.n7281 gnd.n7280 19.3944
R8904 gnd.n7286 gnd.n7281 19.3944
R8905 gnd.n7286 gnd.n7277 19.3944
R8906 gnd.n7290 gnd.n7277 19.3944
R8907 gnd.n7290 gnd.n7275 19.3944
R8908 gnd.n7296 gnd.n7275 19.3944
R8909 gnd.n7296 gnd.n7273 19.3944
R8910 gnd.n7300 gnd.n7273 19.3944
R8911 gnd.n7300 gnd.n7271 19.3944
R8912 gnd.n7306 gnd.n7271 19.3944
R8913 gnd.n7306 gnd.n7269 19.3944
R8914 gnd.n7310 gnd.n7269 19.3944
R8915 gnd.n7310 gnd.n7267 19.3944
R8916 gnd.n7316 gnd.n7267 19.3944
R8917 gnd.n7316 gnd.n7265 19.3944
R8918 gnd.n7320 gnd.n7265 19.3944
R8919 gnd.n5343 gnd.n3416 19.3944
R8920 gnd.n5343 gnd.n3417 19.3944
R8921 gnd.n5339 gnd.n3417 19.3944
R8922 gnd.n5339 gnd.n5338 19.3944
R8923 gnd.n5338 gnd.n5337 19.3944
R8924 gnd.n5337 gnd.n5309 19.3944
R8925 gnd.n5333 gnd.n5309 19.3944
R8926 gnd.n5333 gnd.n5332 19.3944
R8927 gnd.n5332 gnd.n5331 19.3944
R8928 gnd.n5331 gnd.n3400 19.3944
R8929 gnd.n5390 gnd.n3400 19.3944
R8930 gnd.n5390 gnd.n3398 19.3944
R8931 gnd.n5394 gnd.n3398 19.3944
R8932 gnd.n5394 gnd.n3395 19.3944
R8933 gnd.n5405 gnd.n3395 19.3944
R8934 gnd.n5405 gnd.n3392 19.3944
R8935 gnd.n5413 gnd.n3392 19.3944
R8936 gnd.n5413 gnd.n3393 19.3944
R8937 gnd.n5409 gnd.n3393 19.3944
R8938 gnd.n5409 gnd.n5408 19.3944
R8939 gnd.n5408 gnd.n68 19.3944
R8940 gnd.n7416 gnd.n68 19.3944
R8941 gnd.n7416 gnd.n7415 19.3944
R8942 gnd.n7415 gnd.n71 19.3944
R8943 gnd.n5440 gnd.n71 19.3944
R8944 gnd.n5440 gnd.n5439 19.3944
R8945 gnd.n5439 gnd.n5438 19.3944
R8946 gnd.n5438 gnd.n395 19.3944
R8947 gnd.n7235 gnd.n395 19.3944
R8948 gnd.n7235 gnd.n393 19.3944
R8949 gnd.n7239 gnd.n393 19.3944
R8950 gnd.n7239 gnd.n390 19.3944
R8951 gnd.n7250 gnd.n390 19.3944
R8952 gnd.n7250 gnd.n388 19.3944
R8953 gnd.n7338 gnd.n388 19.3944
R8954 gnd.n7338 gnd.n7337 19.3944
R8955 gnd.n7337 gnd.n7336 19.3944
R8956 gnd.n7336 gnd.n7334 19.3944
R8957 gnd.n7334 gnd.n7333 19.3944
R8958 gnd.n7333 gnd.n7331 19.3944
R8959 gnd.n7331 gnd.n7330 19.3944
R8960 gnd.n7330 gnd.n7328 19.3944
R8961 gnd.n3283 gnd.n3282 19.3944
R8962 gnd.n5518 gnd.n3282 19.3944
R8963 gnd.n5518 gnd.n5517 19.3944
R8964 gnd.n5517 gnd.n5516 19.3944
R8965 gnd.n5516 gnd.n3289 19.3944
R8966 gnd.n5506 gnd.n3289 19.3944
R8967 gnd.n5506 gnd.n5505 19.3944
R8968 gnd.n5505 gnd.n5504 19.3944
R8969 gnd.n5504 gnd.n3312 19.3944
R8970 gnd.n5494 gnd.n3312 19.3944
R8971 gnd.n5494 gnd.n5493 19.3944
R8972 gnd.n5493 gnd.n5492 19.3944
R8973 gnd.n5492 gnd.n3333 19.3944
R8974 gnd.n5482 gnd.n3333 19.3944
R8975 gnd.n5482 gnd.n5481 19.3944
R8976 gnd.n5481 gnd.n5480 19.3944
R8977 gnd.n5470 gnd.n5469 19.3944
R8978 gnd.n3367 gnd.n3366 19.3944
R8979 gnd.n3376 gnd.n3375 19.3944
R8980 gnd.n7411 gnd.n7410 19.3944
R8981 gnd.n7407 gnd.n80 19.3944
R8982 gnd.n7407 gnd.n87 19.3944
R8983 gnd.n7397 gnd.n87 19.3944
R8984 gnd.n7397 gnd.n7396 19.3944
R8985 gnd.n7396 gnd.n7395 19.3944
R8986 gnd.n7395 gnd.n109 19.3944
R8987 gnd.n7385 gnd.n109 19.3944
R8988 gnd.n7385 gnd.n7384 19.3944
R8989 gnd.n7384 gnd.n7383 19.3944
R8990 gnd.n7383 gnd.n129 19.3944
R8991 gnd.n7373 gnd.n129 19.3944
R8992 gnd.n7373 gnd.n7372 19.3944
R8993 gnd.n7372 gnd.n7371 19.3944
R8994 gnd.n7371 gnd.n149 19.3944
R8995 gnd.n7361 gnd.n149 19.3944
R8996 gnd.n7361 gnd.n7360 19.3944
R8997 gnd.n7360 gnd.n7359 19.3944
R8998 gnd.n4073 gnd.n4069 19.3944
R8999 gnd.n4073 gnd.n4067 19.3944
R9000 gnd.n4212 gnd.n4067 19.3944
R9001 gnd.n4212 gnd.n4065 19.3944
R9002 gnd.n4217 gnd.n4065 19.3944
R9003 gnd.n4217 gnd.n4062 19.3944
R9004 gnd.n4221 gnd.n4062 19.3944
R9005 gnd.n4222 gnd.n4221 19.3944
R9006 gnd.n4237 gnd.n4236 19.3944
R9007 gnd.n4234 gnd.n4224 19.3944
R9008 gnd.n4230 gnd.n4229 19.3944
R9009 gnd.n4227 gnd.n4021 19.3944
R9010 gnd.n4294 gnd.n4293 19.3944
R9011 gnd.n4314 gnd.n4294 19.3944
R9012 gnd.n4314 gnd.n4313 19.3944
R9013 gnd.n4313 gnd.n4312 19.3944
R9014 gnd.n4312 gnd.n4299 19.3944
R9015 gnd.n4308 gnd.n4299 19.3944
R9016 gnd.n4308 gnd.n4307 19.3944
R9017 gnd.n4307 gnd.n4306 19.3944
R9018 gnd.n4306 gnd.n3997 19.3944
R9019 gnd.n4366 gnd.n3997 19.3944
R9020 gnd.n4366 gnd.n3995 19.3944
R9021 gnd.n4370 gnd.n3995 19.3944
R9022 gnd.n4370 gnd.n3993 19.3944
R9023 gnd.n4374 gnd.n3993 19.3944
R9024 gnd.n4374 gnd.n3991 19.3944
R9025 gnd.n4378 gnd.n3991 19.3944
R9026 gnd.n4378 gnd.n3989 19.3944
R9027 gnd.n4382 gnd.n3989 19.3944
R9028 gnd.n4382 gnd.n3987 19.3944
R9029 gnd.n4386 gnd.n3987 19.3944
R9030 gnd.n4386 gnd.n3985 19.3944
R9031 gnd.n4391 gnd.n3985 19.3944
R9032 gnd.n4391 gnd.n3983 19.3944
R9033 gnd.n4395 gnd.n3983 19.3944
R9034 gnd.n4395 gnd.n3921 19.3944
R9035 gnd.n4407 gnd.n3921 19.3944
R9036 gnd.n4407 gnd.n3919 19.3944
R9037 gnd.n4411 gnd.n3919 19.3944
R9038 gnd.n4411 gnd.n3907 19.3944
R9039 gnd.n4423 gnd.n3907 19.3944
R9040 gnd.n4423 gnd.n3905 19.3944
R9041 gnd.n4427 gnd.n3905 19.3944
R9042 gnd.n4427 gnd.n3893 19.3944
R9043 gnd.n4439 gnd.n3893 19.3944
R9044 gnd.n4439 gnd.n3891 19.3944
R9045 gnd.n4443 gnd.n3891 19.3944
R9046 gnd.n4443 gnd.n3879 19.3944
R9047 gnd.n4455 gnd.n3879 19.3944
R9048 gnd.n4455 gnd.n3877 19.3944
R9049 gnd.n4459 gnd.n3877 19.3944
R9050 gnd.n4459 gnd.n3862 19.3944
R9051 gnd.n4482 gnd.n3862 19.3944
R9052 gnd.n4482 gnd.n3860 19.3944
R9053 gnd.n4489 gnd.n3860 19.3944
R9054 gnd.n4489 gnd.n4488 19.3944
R9055 gnd.n4488 gnd.n2981 19.3944
R9056 gnd.n5838 gnd.n2981 19.3944
R9057 gnd.n5838 gnd.n5837 19.3944
R9058 gnd.n5837 gnd.n5836 19.3944
R9059 gnd.n5836 gnd.n2985 19.3944
R9060 gnd.n4521 gnd.n2985 19.3944
R9061 gnd.n4521 gnd.n4520 19.3944
R9062 gnd.n4520 gnd.n3745 19.3944
R9063 gnd.n4573 gnd.n3745 19.3944
R9064 gnd.n4573 gnd.n3743 19.3944
R9065 gnd.n4579 gnd.n3743 19.3944
R9066 gnd.n4579 gnd.n4578 19.3944
R9067 gnd.n4578 gnd.n3723 19.3944
R9068 gnd.n4613 gnd.n3723 19.3944
R9069 gnd.n4613 gnd.n3721 19.3944
R9070 gnd.n4617 gnd.n3721 19.3944
R9071 gnd.n4617 gnd.n3697 19.3944
R9072 gnd.n4657 gnd.n3697 19.3944
R9073 gnd.n4657 gnd.n3695 19.3944
R9074 gnd.n4663 gnd.n3695 19.3944
R9075 gnd.n4663 gnd.n4662 19.3944
R9076 gnd.n4662 gnd.n3677 19.3944
R9077 gnd.n4709 gnd.n3677 19.3944
R9078 gnd.n4709 gnd.n3675 19.3944
R9079 gnd.n4724 gnd.n3675 19.3944
R9080 gnd.n4724 gnd.n4723 19.3944
R9081 gnd.n4723 gnd.n4722 19.3944
R9082 gnd.n4722 gnd.n4715 19.3944
R9083 gnd.n4718 gnd.n4715 19.3944
R9084 gnd.n4718 gnd.n3639 19.3944
R9085 gnd.n4771 gnd.n3639 19.3944
R9086 gnd.n4771 gnd.n3637 19.3944
R9087 gnd.n4775 gnd.n3637 19.3944
R9088 gnd.n4775 gnd.n3617 19.3944
R9089 gnd.n4831 gnd.n3617 19.3944
R9090 gnd.n4831 gnd.n3615 19.3944
R9091 gnd.n4835 gnd.n3615 19.3944
R9092 gnd.n4835 gnd.n3599 19.3944
R9093 gnd.n4859 gnd.n3599 19.3944
R9094 gnd.n4859 gnd.n3597 19.3944
R9095 gnd.n4863 gnd.n3597 19.3944
R9096 gnd.n4863 gnd.n3581 19.3944
R9097 gnd.n4884 gnd.n3581 19.3944
R9098 gnd.n4884 gnd.n3579 19.3944
R9099 gnd.n4890 gnd.n3579 19.3944
R9100 gnd.n4890 gnd.n4889 19.3944
R9101 gnd.n4889 gnd.n3552 19.3944
R9102 gnd.n4940 gnd.n3552 19.3944
R9103 gnd.n4940 gnd.n3550 19.3944
R9104 gnd.n4946 gnd.n3550 19.3944
R9105 gnd.n4946 gnd.n4945 19.3944
R9106 gnd.n4945 gnd.n3521 19.3944
R9107 gnd.n5171 gnd.n3521 19.3944
R9108 gnd.n5171 gnd.n3519 19.3944
R9109 gnd.n5175 gnd.n3519 19.3944
R9110 gnd.n5175 gnd.n3509 19.3944
R9111 gnd.n5189 gnd.n3509 19.3944
R9112 gnd.n5189 gnd.n3507 19.3944
R9113 gnd.n5193 gnd.n3507 19.3944
R9114 gnd.n5193 gnd.n3498 19.3944
R9115 gnd.n5206 gnd.n3498 19.3944
R9116 gnd.n5206 gnd.n3496 19.3944
R9117 gnd.n5210 gnd.n3496 19.3944
R9118 gnd.n5210 gnd.n3486 19.3944
R9119 gnd.n5223 gnd.n3486 19.3944
R9120 gnd.n5223 gnd.n3484 19.3944
R9121 gnd.n5227 gnd.n3484 19.3944
R9122 gnd.n5227 gnd.n3474 19.3944
R9123 gnd.n5240 gnd.n3474 19.3944
R9124 gnd.n5240 gnd.n3472 19.3944
R9125 gnd.n5244 gnd.n3472 19.3944
R9126 gnd.n5244 gnd.n3462 19.3944
R9127 gnd.n5257 gnd.n3462 19.3944
R9128 gnd.n5257 gnd.n3460 19.3944
R9129 gnd.n5264 gnd.n3460 19.3944
R9130 gnd.n5264 gnd.n5263 19.3944
R9131 gnd.n5263 gnd.n3450 19.3944
R9132 gnd.n5278 gnd.n3450 19.3944
R9133 gnd.n5279 gnd.n5278 19.3944
R9134 gnd.n5279 gnd.n3448 19.3944
R9135 gnd.n5294 gnd.n3448 19.3944
R9136 gnd.n5294 gnd.n5293 19.3944
R9137 gnd.n5293 gnd.n5292 19.3944
R9138 gnd.n5292 gnd.n5285 19.3944
R9139 gnd.n5288 gnd.n5285 19.3944
R9140 gnd.n5288 gnd.n3414 19.3944
R9141 gnd.n5348 gnd.n3414 19.3944
R9142 gnd.n5348 gnd.n3412 19.3944
R9143 gnd.n5352 gnd.n3412 19.3944
R9144 gnd.n5352 gnd.n3410 19.3944
R9145 gnd.n5356 gnd.n3410 19.3944
R9146 gnd.n5356 gnd.n3408 19.3944
R9147 gnd.n5360 gnd.n3408 19.3944
R9148 gnd.n5360 gnd.n3406 19.3944
R9149 gnd.n5364 gnd.n3406 19.3944
R9150 gnd.n5364 gnd.n3404 19.3944
R9151 gnd.n5385 gnd.n3404 19.3944
R9152 gnd.n5385 gnd.n5384 19.3944
R9153 gnd.n5384 gnd.n5383 19.3944
R9154 gnd.n5383 gnd.n5370 19.3944
R9155 gnd.n5379 gnd.n5370 19.3944
R9156 gnd.n5379 gnd.n5378 19.3944
R9157 gnd.n5376 gnd.n5374 19.3944
R9158 gnd.n5464 gnd.n5463 19.3944
R9159 gnd.n5461 gnd.n3373 19.3944
R9160 gnd.n5449 gnd.n5446 19.3944
R9161 gnd.n5447 gnd.n400 19.3944
R9162 gnd.n7223 gnd.n400 19.3944
R9163 gnd.n7223 gnd.n7222 19.3944
R9164 gnd.n7222 gnd.n7221 19.3944
R9165 gnd.n7221 gnd.n405 19.3944
R9166 gnd.n7217 gnd.n405 19.3944
R9167 gnd.n7217 gnd.n7216 19.3944
R9168 gnd.n7216 gnd.n7215 19.3944
R9169 gnd.n6273 gnd.n6272 19.3944
R9170 gnd.n6272 gnd.n6271 19.3944
R9171 gnd.n6271 gnd.n6270 19.3944
R9172 gnd.n6270 gnd.n6268 19.3944
R9173 gnd.n6268 gnd.n6265 19.3944
R9174 gnd.n6265 gnd.n6264 19.3944
R9175 gnd.n6264 gnd.n6261 19.3944
R9176 gnd.n6261 gnd.n6260 19.3944
R9177 gnd.n6260 gnd.n6257 19.3944
R9178 gnd.n6257 gnd.n6256 19.3944
R9179 gnd.n6256 gnd.n6253 19.3944
R9180 gnd.n6253 gnd.n6252 19.3944
R9181 gnd.n6252 gnd.n6249 19.3944
R9182 gnd.n6249 gnd.n6248 19.3944
R9183 gnd.n6248 gnd.n6245 19.3944
R9184 gnd.n6245 gnd.n6244 19.3944
R9185 gnd.n6244 gnd.n6241 19.3944
R9186 gnd.n6239 gnd.n6236 19.3944
R9187 gnd.n6236 gnd.n6235 19.3944
R9188 gnd.n6235 gnd.n6232 19.3944
R9189 gnd.n6232 gnd.n6231 19.3944
R9190 gnd.n6231 gnd.n6228 19.3944
R9191 gnd.n6228 gnd.n6227 19.3944
R9192 gnd.n6227 gnd.n6224 19.3944
R9193 gnd.n6224 gnd.n6223 19.3944
R9194 gnd.n6223 gnd.n6220 19.3944
R9195 gnd.n6220 gnd.n6219 19.3944
R9196 gnd.n6219 gnd.n6216 19.3944
R9197 gnd.n6216 gnd.n6215 19.3944
R9198 gnd.n6215 gnd.n6212 19.3944
R9199 gnd.n6212 gnd.n6211 19.3944
R9200 gnd.n6211 gnd.n6208 19.3944
R9201 gnd.n6208 gnd.n6207 19.3944
R9202 gnd.n6207 gnd.n6204 19.3944
R9203 gnd.n6204 gnd.n6203 19.3944
R9204 gnd.n6199 gnd.n6196 19.3944
R9205 gnd.n6196 gnd.n6195 19.3944
R9206 gnd.n6195 gnd.n6192 19.3944
R9207 gnd.n6192 gnd.n6191 19.3944
R9208 gnd.n6191 gnd.n6188 19.3944
R9209 gnd.n6188 gnd.n6187 19.3944
R9210 gnd.n6187 gnd.n6184 19.3944
R9211 gnd.n6184 gnd.n6183 19.3944
R9212 gnd.n6183 gnd.n6180 19.3944
R9213 gnd.n6180 gnd.n6179 19.3944
R9214 gnd.n6179 gnd.n6176 19.3944
R9215 gnd.n6176 gnd.n6175 19.3944
R9216 gnd.n6175 gnd.n6172 19.3944
R9217 gnd.n6172 gnd.n6171 19.3944
R9218 gnd.n6171 gnd.n6168 19.3944
R9219 gnd.n6168 gnd.n6167 19.3944
R9220 gnd.n6167 gnd.n6164 19.3944
R9221 gnd.n6164 gnd.n6163 19.3944
R9222 gnd.n4111 gnd.n4110 19.3944
R9223 gnd.n4114 gnd.n4111 19.3944
R9224 gnd.n4114 gnd.n4106 19.3944
R9225 gnd.n4120 gnd.n4106 19.3944
R9226 gnd.n4121 gnd.n4120 19.3944
R9227 gnd.n4124 gnd.n4121 19.3944
R9228 gnd.n4124 gnd.n4104 19.3944
R9229 gnd.n4130 gnd.n4104 19.3944
R9230 gnd.n4131 gnd.n4130 19.3944
R9231 gnd.n4134 gnd.n4131 19.3944
R9232 gnd.n4134 gnd.n4102 19.3944
R9233 gnd.n4140 gnd.n4102 19.3944
R9234 gnd.n4141 gnd.n4140 19.3944
R9235 gnd.n4144 gnd.n4141 19.3944
R9236 gnd.n4144 gnd.n4098 19.3944
R9237 gnd.n4148 gnd.n4098 19.3944
R9238 gnd.n4155 gnd.n4154 19.3944
R9239 gnd.n4157 gnd.n4155 19.3944
R9240 gnd.n4157 gnd.n4092 19.3944
R9241 gnd.n4162 gnd.n4092 19.3944
R9242 gnd.n4163 gnd.n4162 19.3944
R9243 gnd.n4165 gnd.n4163 19.3944
R9244 gnd.n4165 gnd.n4090 19.3944
R9245 gnd.n4170 gnd.n4090 19.3944
R9246 gnd.n4170 gnd.n4075 19.3944
R9247 gnd.n4205 gnd.n4075 19.3944
R9248 gnd.n4205 gnd.n4204 19.3944
R9249 gnd.n4204 gnd.n4203 19.3944
R9250 gnd.n4203 gnd.n4079 19.3944
R9251 gnd.n4193 gnd.n4079 19.3944
R9252 gnd.n4193 gnd.n4192 19.3944
R9253 gnd.n4192 gnd.n4191 19.3944
R9254 gnd.n4191 gnd.n4186 19.3944
R9255 gnd.n4186 gnd.n4050 19.3944
R9256 gnd.n4253 gnd.n4050 19.3944
R9257 gnd.n4253 gnd.n4048 19.3944
R9258 gnd.n4257 gnd.n4048 19.3944
R9259 gnd.n4257 gnd.n4027 19.3944
R9260 gnd.n4283 gnd.n4027 19.3944
R9261 gnd.n4283 gnd.n4025 19.3944
R9262 gnd.n4287 gnd.n4025 19.3944
R9263 gnd.n4287 gnd.n4015 19.3944
R9264 gnd.n4319 gnd.n4015 19.3944
R9265 gnd.n4319 gnd.n4013 19.3944
R9266 gnd.n4323 gnd.n4013 19.3944
R9267 gnd.n4323 gnd.n4009 19.3944
R9268 gnd.n4333 gnd.n4009 19.3944
R9269 gnd.n4333 gnd.n4007 19.3944
R9270 gnd.n4337 gnd.n4007 19.3944
R9271 gnd.n4337 gnd.n4000 19.3944
R9272 gnd.n4361 gnd.n4000 19.3944
R9273 gnd.n4361 gnd.n4001 19.3944
R9274 gnd.n4357 gnd.n4001 19.3944
R9275 gnd.n4357 gnd.n4356 19.3944
R9276 gnd.n4356 gnd.n4355 19.3944
R9277 gnd.n4355 gnd.n2641 19.3944
R9278 gnd.n6039 gnd.n2641 19.3944
R9279 gnd.n6039 gnd.n2642 19.3944
R9280 gnd.n6155 gnd.n2451 19.3944
R9281 gnd.n4081 gnd.n2451 19.3944
R9282 gnd.n4082 gnd.n4081 19.3944
R9283 gnd.n4084 gnd.n4082 19.3944
R9284 gnd.n4085 gnd.n4084 19.3944
R9285 gnd.n4088 gnd.n4085 19.3944
R9286 gnd.n4089 gnd.n4088 19.3944
R9287 gnd.n4174 gnd.n4089 19.3944
R9288 gnd.n4175 gnd.n4174 19.3944
R9289 gnd.n4177 gnd.n4175 19.3944
R9290 gnd.n4178 gnd.n4177 19.3944
R9291 gnd.n4199 gnd.n4178 19.3944
R9292 gnd.n4199 gnd.n4198 19.3944
R9293 gnd.n4198 gnd.n4197 19.3944
R9294 gnd.n4197 gnd.n4180 19.3944
R9295 gnd.n4187 gnd.n4180 19.3944
R9296 gnd.n4187 gnd.n4059 19.3944
R9297 gnd.n4242 gnd.n4059 19.3944
R9298 gnd.n4243 gnd.n4242 19.3944
R9299 gnd.n4243 gnd.n4043 19.3944
R9300 gnd.n4261 gnd.n4043 19.3944
R9301 gnd.n4262 gnd.n4261 19.3944
R9302 gnd.n4263 gnd.n4262 19.3944
R9303 gnd.n4268 gnd.n4263 19.3944
R9304 gnd.n4268 gnd.n4266 19.3944
R9305 gnd.n4266 gnd.n4265 19.3944
R9306 gnd.n4265 gnd.n4264 19.3944
R9307 gnd.n4264 gnd.n4011 19.3944
R9308 gnd.n4327 gnd.n4011 19.3944
R9309 gnd.n4328 gnd.n4327 19.3944
R9310 gnd.n4329 gnd.n4328 19.3944
R9311 gnd.n4329 gnd.n4005 19.3944
R9312 gnd.n4341 gnd.n4005 19.3944
R9313 gnd.n4342 gnd.n4341 19.3944
R9314 gnd.n4343 gnd.n4342 19.3944
R9315 gnd.n4344 gnd.n4343 19.3944
R9316 gnd.n4348 gnd.n4344 19.3944
R9317 gnd.n4349 gnd.n4348 19.3944
R9318 gnd.n4350 gnd.n4349 19.3944
R9319 gnd.n4350 gnd.n2639 19.3944
R9320 gnd.n6043 gnd.n2639 19.3944
R9321 gnd.n6044 gnd.n6043 19.3944
R9322 gnd.n2470 gnd.n2449 19.3944
R9323 gnd.n2471 gnd.n2470 19.3944
R9324 gnd.n6144 gnd.n2471 19.3944
R9325 gnd.n6144 gnd.n6143 19.3944
R9326 gnd.n6143 gnd.n6142 19.3944
R9327 gnd.n6142 gnd.n2475 19.3944
R9328 gnd.n6132 gnd.n2475 19.3944
R9329 gnd.n6132 gnd.n6131 19.3944
R9330 gnd.n6131 gnd.n6130 19.3944
R9331 gnd.n6130 gnd.n2494 19.3944
R9332 gnd.n6120 gnd.n2494 19.3944
R9333 gnd.n6120 gnd.n6119 19.3944
R9334 gnd.n6119 gnd.n6118 19.3944
R9335 gnd.n6118 gnd.n2514 19.3944
R9336 gnd.n6108 gnd.n2514 19.3944
R9337 gnd.n6108 gnd.n6107 19.3944
R9338 gnd.n6107 gnd.n6106 19.3944
R9339 gnd.n6106 gnd.n2535 19.3944
R9340 gnd.n4057 gnd.n2535 19.3944
R9341 gnd.n4246 gnd.n4057 19.3944
R9342 gnd.n4246 gnd.n4039 19.3944
R9343 gnd.n4273 gnd.n4039 19.3944
R9344 gnd.n4273 gnd.n4272 19.3944
R9345 gnd.n4272 gnd.n4271 19.3944
R9346 gnd.n4271 gnd.n2558 19.3944
R9347 gnd.n6094 gnd.n2558 19.3944
R9348 gnd.n6094 gnd.n6093 19.3944
R9349 gnd.n6093 gnd.n6092 19.3944
R9350 gnd.n6092 gnd.n2562 19.3944
R9351 gnd.n6082 gnd.n2562 19.3944
R9352 gnd.n6082 gnd.n6081 19.3944
R9353 gnd.n6081 gnd.n6080 19.3944
R9354 gnd.n6080 gnd.n2580 19.3944
R9355 gnd.n6070 gnd.n2580 19.3944
R9356 gnd.n6070 gnd.n6069 19.3944
R9357 gnd.n6069 gnd.n6068 19.3944
R9358 gnd.n6068 gnd.n2601 19.3944
R9359 gnd.n6058 gnd.n2601 19.3944
R9360 gnd.n6058 gnd.n6057 19.3944
R9361 gnd.n6057 gnd.n6056 19.3944
R9362 gnd.n6056 gnd.n2621 19.3944
R9363 gnd.n6046 gnd.n2621 19.3944
R9364 gnd.n2784 gnd.n2783 19.3944
R9365 gnd.n5962 gnd.n2783 19.3944
R9366 gnd.n5962 gnd.n5961 19.3944
R9367 gnd.n5961 gnd.n5960 19.3944
R9368 gnd.n5960 gnd.n5957 19.3944
R9369 gnd.n5957 gnd.n5956 19.3944
R9370 gnd.n5956 gnd.n5953 19.3944
R9371 gnd.n5953 gnd.n5952 19.3944
R9372 gnd.n5952 gnd.n5949 19.3944
R9373 gnd.n5949 gnd.n5948 19.3944
R9374 gnd.n5948 gnd.n5945 19.3944
R9375 gnd.n5945 gnd.n5944 19.3944
R9376 gnd.n5944 gnd.n5941 19.3944
R9377 gnd.n5941 gnd.n5940 19.3944
R9378 gnd.n5940 gnd.n5937 19.3944
R9379 gnd.n5937 gnd.n5936 19.3944
R9380 gnd.n5936 gnd.n5933 19.3944
R9381 gnd.n2886 gnd.n2822 19.3944
R9382 gnd.n2886 gnd.n2883 19.3944
R9383 gnd.n2883 gnd.n2880 19.3944
R9384 gnd.n2880 gnd.n2879 19.3944
R9385 gnd.n2879 gnd.n2876 19.3944
R9386 gnd.n2876 gnd.n2875 19.3944
R9387 gnd.n2875 gnd.n2872 19.3944
R9388 gnd.n2872 gnd.n2871 19.3944
R9389 gnd.n2871 gnd.n2868 19.3944
R9390 gnd.n2868 gnd.n2867 19.3944
R9391 gnd.n2867 gnd.n2864 19.3944
R9392 gnd.n2864 gnd.n2863 19.3944
R9393 gnd.n2863 gnd.n2860 19.3944
R9394 gnd.n2860 gnd.n2859 19.3944
R9395 gnd.n2859 gnd.n2856 19.3944
R9396 gnd.n2856 gnd.n2855 19.3944
R9397 gnd.n2855 gnd.n2852 19.3944
R9398 gnd.n2852 gnd.n2851 19.3944
R9399 gnd.n2908 gnd.n2813 19.3944
R9400 gnd.n2908 gnd.n2905 19.3944
R9401 gnd.n2905 gnd.n2902 19.3944
R9402 gnd.n2902 gnd.n2901 19.3944
R9403 gnd.n2901 gnd.n2898 19.3944
R9404 gnd.n2898 gnd.n2897 19.3944
R9405 gnd.n2897 gnd.n2894 19.3944
R9406 gnd.n2894 gnd.n2893 19.3944
R9407 gnd.n5931 gnd.n5928 19.3944
R9408 gnd.n5928 gnd.n5927 19.3944
R9409 gnd.n5927 gnd.n5924 19.3944
R9410 gnd.n5924 gnd.n5923 19.3944
R9411 gnd.n5923 gnd.n5920 19.3944
R9412 gnd.n5920 gnd.n5919 19.3944
R9413 gnd.n5919 gnd.n5916 19.3944
R9414 gnd.n6150 gnd.n2457 19.3944
R9415 gnd.n6150 gnd.n6149 19.3944
R9416 gnd.n6149 gnd.n6148 19.3944
R9417 gnd.n6148 gnd.n2462 19.3944
R9418 gnd.n6138 gnd.n2462 19.3944
R9419 gnd.n6138 gnd.n6137 19.3944
R9420 gnd.n6137 gnd.n6136 19.3944
R9421 gnd.n6136 gnd.n2485 19.3944
R9422 gnd.n6126 gnd.n2485 19.3944
R9423 gnd.n6126 gnd.n6125 19.3944
R9424 gnd.n6125 gnd.n6124 19.3944
R9425 gnd.n6124 gnd.n2504 19.3944
R9426 gnd.n6114 gnd.n2504 19.3944
R9427 gnd.n6114 gnd.n6113 19.3944
R9428 gnd.n6113 gnd.n6112 19.3944
R9429 gnd.n6112 gnd.n2525 19.3944
R9430 gnd.n6102 gnd.n6101 19.3944
R9431 gnd.n4056 gnd.n2542 19.3944
R9432 gnd.n4035 gnd.n4034 19.3944
R9433 gnd.n4279 gnd.n4278 19.3944
R9434 gnd.n6098 gnd.n2548 19.3944
R9435 gnd.n6098 gnd.n2549 19.3944
R9436 gnd.n6088 gnd.n2549 19.3944
R9437 gnd.n6088 gnd.n6087 19.3944
R9438 gnd.n6087 gnd.n6086 19.3944
R9439 gnd.n6086 gnd.n2571 19.3944
R9440 gnd.n6076 gnd.n2571 19.3944
R9441 gnd.n6076 gnd.n6075 19.3944
R9442 gnd.n6075 gnd.n6074 19.3944
R9443 gnd.n6074 gnd.n2591 19.3944
R9444 gnd.n6064 gnd.n2591 19.3944
R9445 gnd.n6064 gnd.n6063 19.3944
R9446 gnd.n6063 gnd.n6062 19.3944
R9447 gnd.n6062 gnd.n2611 19.3944
R9448 gnd.n6052 gnd.n2611 19.3944
R9449 gnd.n6052 gnd.n6051 19.3944
R9450 gnd.n6051 gnd.n6050 19.3944
R9451 gnd.n6540 gnd.n812 19.3944
R9452 gnd.n6540 gnd.n6539 19.3944
R9453 gnd.n6539 gnd.n6538 19.3944
R9454 gnd.n6538 gnd.n816 19.3944
R9455 gnd.n6532 gnd.n816 19.3944
R9456 gnd.n6532 gnd.n6531 19.3944
R9457 gnd.n6531 gnd.n6530 19.3944
R9458 gnd.n6530 gnd.n824 19.3944
R9459 gnd.n6524 gnd.n824 19.3944
R9460 gnd.n6524 gnd.n6523 19.3944
R9461 gnd.n6523 gnd.n6522 19.3944
R9462 gnd.n6522 gnd.n832 19.3944
R9463 gnd.n6516 gnd.n832 19.3944
R9464 gnd.n6516 gnd.n6515 19.3944
R9465 gnd.n6515 gnd.n6514 19.3944
R9466 gnd.n6514 gnd.n840 19.3944
R9467 gnd.n6508 gnd.n840 19.3944
R9468 gnd.n6508 gnd.n6507 19.3944
R9469 gnd.n6507 gnd.n6506 19.3944
R9470 gnd.n6506 gnd.n848 19.3944
R9471 gnd.n6500 gnd.n848 19.3944
R9472 gnd.n6500 gnd.n6499 19.3944
R9473 gnd.n6499 gnd.n6498 19.3944
R9474 gnd.n6498 gnd.n856 19.3944
R9475 gnd.n6492 gnd.n856 19.3944
R9476 gnd.n6492 gnd.n6491 19.3944
R9477 gnd.n6491 gnd.n6490 19.3944
R9478 gnd.n6490 gnd.n864 19.3944
R9479 gnd.n6484 gnd.n864 19.3944
R9480 gnd.n6484 gnd.n6483 19.3944
R9481 gnd.n6483 gnd.n6482 19.3944
R9482 gnd.n6482 gnd.n872 19.3944
R9483 gnd.n6476 gnd.n872 19.3944
R9484 gnd.n6476 gnd.n6475 19.3944
R9485 gnd.n6475 gnd.n6474 19.3944
R9486 gnd.n6474 gnd.n880 19.3944
R9487 gnd.n6468 gnd.n880 19.3944
R9488 gnd.n6468 gnd.n6467 19.3944
R9489 gnd.n6467 gnd.n6466 19.3944
R9490 gnd.n6466 gnd.n888 19.3944
R9491 gnd.n6460 gnd.n888 19.3944
R9492 gnd.n6460 gnd.n6459 19.3944
R9493 gnd.n6459 gnd.n6458 19.3944
R9494 gnd.n6458 gnd.n896 19.3944
R9495 gnd.n6452 gnd.n896 19.3944
R9496 gnd.n6452 gnd.n6451 19.3944
R9497 gnd.n6451 gnd.n6450 19.3944
R9498 gnd.n6450 gnd.n904 19.3944
R9499 gnd.n6444 gnd.n904 19.3944
R9500 gnd.n6444 gnd.n6443 19.3944
R9501 gnd.n6443 gnd.n6442 19.3944
R9502 gnd.n6442 gnd.n912 19.3944
R9503 gnd.n6436 gnd.n912 19.3944
R9504 gnd.n6436 gnd.n6435 19.3944
R9505 gnd.n6435 gnd.n6434 19.3944
R9506 gnd.n6434 gnd.n920 19.3944
R9507 gnd.n6428 gnd.n920 19.3944
R9508 gnd.n6428 gnd.n6427 19.3944
R9509 gnd.n6427 gnd.n6426 19.3944
R9510 gnd.n6426 gnd.n928 19.3944
R9511 gnd.n6420 gnd.n928 19.3944
R9512 gnd.n6420 gnd.n6419 19.3944
R9513 gnd.n6419 gnd.n6418 19.3944
R9514 gnd.n6418 gnd.n936 19.3944
R9515 gnd.n6412 gnd.n936 19.3944
R9516 gnd.n6412 gnd.n6411 19.3944
R9517 gnd.n6411 gnd.n6410 19.3944
R9518 gnd.n6410 gnd.n944 19.3944
R9519 gnd.n6404 gnd.n944 19.3944
R9520 gnd.n6404 gnd.n6403 19.3944
R9521 gnd.n6403 gnd.n6402 19.3944
R9522 gnd.n6402 gnd.n952 19.3944
R9523 gnd.n6396 gnd.n952 19.3944
R9524 gnd.n6396 gnd.n6395 19.3944
R9525 gnd.n6395 gnd.n6394 19.3944
R9526 gnd.n6394 gnd.n960 19.3944
R9527 gnd.n6388 gnd.n960 19.3944
R9528 gnd.n6388 gnd.n6387 19.3944
R9529 gnd.n6387 gnd.n6386 19.3944
R9530 gnd.n6386 gnd.n968 19.3944
R9531 gnd.n6380 gnd.n968 19.3944
R9532 gnd.n6380 gnd.n6379 19.3944
R9533 gnd.n6379 gnd.n6378 19.3944
R9534 gnd.n6378 gnd.n976 19.3944
R9535 gnd.n3980 gnd.n3931 19.3944
R9536 gnd.n3980 gnd.n3932 19.3944
R9537 gnd.n3976 gnd.n3932 19.3944
R9538 gnd.n3976 gnd.n3975 19.3944
R9539 gnd.n3975 gnd.n3974 19.3944
R9540 gnd.n3974 gnd.n3937 19.3944
R9541 gnd.n3970 gnd.n3937 19.3944
R9542 gnd.n3970 gnd.n3969 19.3944
R9543 gnd.n3969 gnd.n3968 19.3944
R9544 gnd.n3968 gnd.n3941 19.3944
R9545 gnd.n3964 gnd.n3941 19.3944
R9546 gnd.n3964 gnd.n3963 19.3944
R9547 gnd.n3963 gnd.n3962 19.3944
R9548 gnd.n3962 gnd.n3945 19.3944
R9549 gnd.n3958 gnd.n3945 19.3944
R9550 gnd.n3958 gnd.n3957 19.3944
R9551 gnd.n3957 gnd.n3956 19.3944
R9552 gnd.n3956 gnd.n3949 19.3944
R9553 gnd.n3952 gnd.n3949 19.3944
R9554 gnd.n3952 gnd.n3951 19.3944
R9555 gnd.n3951 gnd.n3855 19.3944
R9556 gnd.n4495 gnd.n3855 19.3944
R9557 gnd.n4495 gnd.n3853 19.3944
R9558 gnd.n4499 gnd.n3853 19.3944
R9559 gnd.n4502 gnd.n4499 19.3944
R9560 gnd.n4503 gnd.n4502 19.3944
R9561 gnd.n4503 gnd.n3850 19.3944
R9562 gnd.n4513 gnd.n3850 19.3944
R9563 gnd.n4513 gnd.n3851 19.3944
R9564 gnd.n4509 gnd.n3851 19.3944
R9565 gnd.n4509 gnd.n4508 19.3944
R9566 gnd.n4508 gnd.n3737 19.3944
R9567 gnd.n4583 gnd.n3737 19.3944
R9568 gnd.n4583 gnd.n3734 19.3944
R9569 gnd.n4600 gnd.n3734 19.3944
R9570 gnd.n4600 gnd.n3735 19.3944
R9571 gnd.n4596 gnd.n3735 19.3944
R9572 gnd.n4596 gnd.n4595 19.3944
R9573 gnd.n4595 gnd.n4594 19.3944
R9574 gnd.n4594 gnd.n4591 19.3944
R9575 gnd.n4591 gnd.n3690 19.3944
R9576 gnd.n4667 gnd.n3690 19.3944
R9577 gnd.n4667 gnd.n3687 19.3944
R9578 gnd.n4697 gnd.n3687 19.3944
R9579 gnd.n4697 gnd.n3688 19.3944
R9580 gnd.n4693 gnd.n3688 19.3944
R9581 gnd.n4693 gnd.n4692 19.3944
R9582 gnd.n4692 gnd.n4691 19.3944
R9583 gnd.n4691 gnd.n4673 19.3944
R9584 gnd.n4687 gnd.n4673 19.3944
R9585 gnd.n4687 gnd.n4686 19.3944
R9586 gnd.n4686 gnd.n4685 19.3944
R9587 gnd.n4685 gnd.n4678 19.3944
R9588 gnd.n4681 gnd.n4678 19.3944
R9589 gnd.n4681 gnd.n3628 19.3944
R9590 gnd.n4816 gnd.n3628 19.3944
R9591 gnd.n4816 gnd.n3629 19.3944
R9592 gnd.n4812 gnd.n3629 19.3944
R9593 gnd.n4812 gnd.n4811 19.3944
R9594 gnd.n4811 gnd.n4810 19.3944
R9595 gnd.n4810 gnd.n4791 19.3944
R9596 gnd.n4806 gnd.n4791 19.3944
R9597 gnd.n4806 gnd.n4805 19.3944
R9598 gnd.n4805 gnd.n4804 19.3944
R9599 gnd.n4804 gnd.n4796 19.3944
R9600 gnd.n4800 gnd.n4796 19.3944
R9601 gnd.n4800 gnd.n4799 19.3944
R9602 gnd.n4799 gnd.n3563 19.3944
R9603 gnd.n4928 gnd.n3563 19.3944
R9604 gnd.n4928 gnd.n3564 19.3944
R9605 gnd.n4924 gnd.n3564 19.3944
R9606 gnd.n4924 gnd.n4923 19.3944
R9607 gnd.n4923 gnd.n4922 19.3944
R9608 gnd.n4922 gnd.n4917 19.3944
R9609 gnd.n4918 gnd.n4917 19.3944
R9610 gnd.n4918 gnd.n3514 19.3944
R9611 gnd.n5179 gnd.n3514 19.3944
R9612 gnd.n5179 gnd.n3512 19.3944
R9613 gnd.n5183 gnd.n3512 19.3944
R9614 gnd.n5183 gnd.n3504 19.3944
R9615 gnd.n5197 gnd.n3504 19.3944
R9616 gnd.n5197 gnd.n3502 19.3944
R9617 gnd.n5201 gnd.n3502 19.3944
R9618 gnd.n5201 gnd.n3492 19.3944
R9619 gnd.n5214 gnd.n3492 19.3944
R9620 gnd.n5214 gnd.n3490 19.3944
R9621 gnd.n5218 gnd.n3490 19.3944
R9622 gnd.n5218 gnd.n3480 19.3944
R9623 gnd.n5231 gnd.n3480 19.3944
R9624 gnd.n5231 gnd.n3478 19.3944
R9625 gnd.n5235 gnd.n3478 19.3944
R9626 gnd.n5235 gnd.n3467 19.3944
R9627 gnd.n5248 gnd.n3467 19.3944
R9628 gnd.n5248 gnd.n3465 19.3944
R9629 gnd.n5252 gnd.n3465 19.3944
R9630 gnd.n5252 gnd.n3456 19.3944
R9631 gnd.n5268 gnd.n3456 19.3944
R9632 gnd.n5268 gnd.n3454 19.3944
R9633 gnd.n5272 gnd.n3454 19.3944
R9634 gnd.n5272 gnd.n3093 19.3944
R9635 gnd.n5715 gnd.n3093 19.3944
R9636 gnd.n5712 gnd.n5711 19.3944
R9637 gnd.n5711 gnd.n5710 19.3944
R9638 gnd.n5710 gnd.n3098 19.3944
R9639 gnd.n5706 gnd.n3098 19.3944
R9640 gnd.n5706 gnd.n5705 19.3944
R9641 gnd.n5705 gnd.n5704 19.3944
R9642 gnd.n5704 gnd.n3103 19.3944
R9643 gnd.n5699 gnd.n3103 19.3944
R9644 gnd.n5699 gnd.n5698 19.3944
R9645 gnd.n5698 gnd.n3108 19.3944
R9646 gnd.n5691 gnd.n3108 19.3944
R9647 gnd.n5691 gnd.n5690 19.3944
R9648 gnd.n5690 gnd.n3117 19.3944
R9649 gnd.n5683 gnd.n3117 19.3944
R9650 gnd.n5683 gnd.n5682 19.3944
R9651 gnd.n5682 gnd.n3125 19.3944
R9652 gnd.n5675 gnd.n3125 19.3944
R9653 gnd.n5675 gnd.n5674 19.3944
R9654 gnd.n5674 gnd.n3133 19.3944
R9655 gnd.n5667 gnd.n3133 19.3944
R9656 gnd.n5667 gnd.n5666 19.3944
R9657 gnd.n5666 gnd.n3141 19.3944
R9658 gnd.n5659 gnd.n3141 19.3944
R9659 gnd.n5659 gnd.n5658 19.3944
R9660 gnd.n3442 gnd.n3421 19.3944
R9661 gnd.n5301 gnd.n3421 19.3944
R9662 gnd.n5301 gnd.n5300 19.3944
R9663 gnd.n4172 gnd.n2496 19.1199
R9664 gnd.n4207 gnd.n2506 19.1199
R9665 gnd.n6122 gnd.n2509 19.1199
R9666 gnd.n4201 gnd.n2516 19.1199
R9667 gnd.n6116 gnd.n2519 19.1199
R9668 gnd.n6110 gnd.n2530 19.1199
R9669 gnd.n4189 gnd.n2537 19.1199
R9670 gnd.n4240 gnd.n4052 19.1199
R9671 gnd.n4251 gnd.n4054 19.1199
R9672 gnd.n4248 gnd.n4046 19.1199
R9673 gnd.n4259 gnd.n4036 19.1199
R9674 gnd.n4281 gnd.n4031 19.1199
R9675 gnd.n4290 gnd.n4022 19.1199
R9676 gnd.n4289 gnd.n2552 19.1199
R9677 gnd.n6096 gnd.n2555 19.1199
R9678 gnd.n4317 gnd.n4316 19.1199
R9679 gnd.n6090 gnd.n2566 19.1199
R9680 gnd.n4325 gnd.n2573 19.1199
R9681 gnd.n4331 gnd.n2582 19.1199
R9682 gnd.n6078 gnd.n2585 19.1199
R9683 gnd.n4339 gnd.n2593 19.1199
R9684 gnd.n6072 gnd.n2596 19.1199
R9685 gnd.n4364 gnd.n4363 19.1199
R9686 gnd.n6066 gnd.n2605 19.1199
R9687 gnd.n4346 gnd.n2613 19.1199
R9688 gnd.n6060 gnd.n2616 19.1199
R9689 gnd.n4352 gnd.n2623 19.1199
R9690 gnd.n6041 gnd.n2632 19.1199
R9691 gnd.n6048 gnd.n2635 19.1199
R9692 gnd.n4530 gnd.t77 19.1199
R9693 gnd.n4956 gnd.t70 19.1199
R9694 gnd.n5528 gnd.n3267 19.1199
R9695 gnd.n5345 gnd.n3269 19.1199
R9696 gnd.n5306 gnd.n3278 19.1199
R9697 gnd.n5514 gnd.n3291 19.1199
R9698 gnd.n5313 gnd.n3294 19.1199
R9699 gnd.n5508 gnd.n3304 19.1199
R9700 gnd.n5319 gnd.n5318 19.1199
R9701 gnd.n5502 gnd.n3314 19.1199
R9702 gnd.n5328 gnd.n3317 19.1199
R9703 gnd.n5496 gnd.n3324 19.1199
R9704 gnd.n5388 gnd.n3327 19.1199
R9705 gnd.n5396 gnd.n3337 19.1199
R9706 gnd.n5484 gnd.n3344 19.1199
R9707 gnd.n5403 gnd.n3396 19.1199
R9708 gnd.n5478 gnd.n3351 19.1199
R9709 gnd.n5415 gnd.n3354 19.1199
R9710 gnd.n5472 gnd.n3361 19.1199
R9711 gnd.n5467 gnd.n3364 19.1199
R9712 gnd.n3390 gnd.n3378 19.1199
R9713 gnd.n5459 gnd.n5458 19.1199
R9714 gnd.n7413 gnd.n73 19.1199
R9715 gnd.n5452 gnd.n75 19.1199
R9716 gnd.n7405 gnd.n90 19.1199
R9717 gnd.n7226 gnd.n93 19.1199
R9718 gnd.n7233 gnd.n104 19.1199
R9719 gnd.n7393 gnd.n111 19.1199
R9720 gnd.n7241 gnd.n392 19.1199
R9721 gnd.n7387 gnd.n120 19.1199
R9722 gnd.n7381 gnd.n131 19.1199
R9723 gnd.t206 gnd.n1271 18.8012
R9724 gnd.n1893 gnd.t31 18.8012
R9725 gnd.n4239 gnd.t233 18.8012
R9726 gnd.n5451 gnd.t237 18.8012
R9727 gnd.n1737 gnd.n1366 18.4825
R9728 gnd.n4620 gnd.n3716 18.4825
R9729 gnd.n4794 gnd.n3594 18.4825
R9730 gnd.n5597 gnd.n5596 18.4247
R9731 gnd.n5916 gnd.n5915 18.4247
R9732 gnd.n5655 gnd.n5654 18.2308
R9733 gnd.n5970 gnd.n5969 18.2308
R9734 gnd.n7320 gnd.n7263 18.2308
R9735 gnd.n4149 gnd.n4148 18.2308
R9736 gnd.n1809 gnd.t155 18.1639
R9737 gnd.n4208 gnd.t217 18.1639
R9738 gnd.t235 gnd.n123 18.1639
R9739 gnd.n5845 gnd.n5844 17.6395
R9740 gnd.n5159 gnd.n5158 17.6395
R9741 gnd.n1790 gnd.t168 17.5266
R9742 gnd.n4642 gnd.t200 17.5266
R9743 gnd.n4787 gnd.t18 17.5266
R9744 gnd.n1299 gnd.t26 16.8893
R9745 gnd.n6152 gnd.t58 16.8893
R9746 gnd.n4491 gnd.t190 16.8893
R9747 gnd.n4604 gnd.t196 16.8893
R9748 gnd.n4894 gnd.t172 16.8893
R9749 gnd.n5185 gnd.t16 16.8893
R9750 gnd.n168 gnd.t36 16.8893
R9751 gnd.n5579 gnd.n5576 16.6793
R9752 gnd.n329 gnd.n199 16.6793
R9753 gnd.n6203 gnd.n6200 16.6793
R9754 gnd.n2893 gnd.n2890 16.6793
R9755 gnd.n4569 gnd.t15 16.5706
R9756 gnd.t12 gnd.n3554 16.5706
R9757 gnd.t137 gnd.n1393 16.2519
R9758 gnd.n1256 gnd.t28 16.2519
R9759 gnd.n3773 gnd.n3772 16.0975
R9760 gnd.n5018 gnd.n5017 16.0975
R9761 gnd.n5847 gnd.n5846 16.0975
R9762 gnd.n5012 gnd.n5011 16.0975
R9763 gnd.n4581 gnd.n3740 15.9333
R9764 gnd.n4727 gnd.t204 15.9333
R9765 gnd.n4747 gnd.n3653 15.9333
R9766 gnd.n4747 gnd.n3655 15.9333
R9767 gnd.t5 gnd.n3634 15.9333
R9768 gnd.n4900 gnd.n3569 15.9333
R9769 gnd.n2295 gnd.n2293 15.6674
R9770 gnd.n2263 gnd.n2261 15.6674
R9771 gnd.n2231 gnd.n2229 15.6674
R9772 gnd.n2200 gnd.n2198 15.6674
R9773 gnd.n2168 gnd.n2166 15.6674
R9774 gnd.n2136 gnd.n2134 15.6674
R9775 gnd.n2104 gnd.n2102 15.6674
R9776 gnd.n2073 gnd.n2071 15.6674
R9777 gnd.n1511 gnd.t137 15.6146
R9778 gnd.n2332 gnd.t43 15.6146
R9779 gnd.t133 gnd.n1040 15.6146
R9780 gnd.n5536 gnd.n5531 15.3217
R9781 gnd.n384 gnd.n177 15.3217
R9782 gnd.n6160 gnd.n2445 15.3217
R9783 gnd.n2848 gnd.n2843 15.3217
R9784 gnd.n4633 gnd.t184 15.296
R9785 gnd.n4778 gnd.t13 15.296
R9786 gnd.n4974 gnd.n4973 15.0827
R9787 gnd.n2960 gnd.n2955 15.0481
R9788 gnd.n4984 gnd.n4983 15.0481
R9789 gnd.n1173 gnd.t167 14.9773
R9790 gnd.n2464 gnd.t58 14.9773
R9791 gnd.n6054 gnd.t66 14.9773
R9792 gnd.n3866 gnd.t190 14.9773
R9793 gnd.n5195 gnd.t16 14.9773
R9794 gnd.n5520 gnd.t50 14.9773
R9795 gnd.n7363 gnd.t36 14.9773
R9796 gnd.t73 gnd.n2989 14.6587
R9797 gnd.t30 gnd.n3747 14.6587
R9798 gnd.n4571 gnd.n4569 14.6587
R9799 gnd.n4611 gnd.n3725 14.6587
R9800 gnd.n4882 gnd.n4881 14.6587
R9801 gnd.n4938 gnd.n3554 14.6587
R9802 gnd.n4937 gnd.t4 14.6587
R9803 gnd.t62 gnd.n3523 14.6587
R9804 gnd.t207 gnd.n992 14.34
R9805 gnd.n1151 gnd.t25 14.34
R9806 gnd.t180 gnd.n1305 13.7027
R9807 gnd.n1706 gnd.n1702 13.5763
R9808 gnd.n6331 gnd.n1053 13.5763
R9809 gnd.n1738 gnd.n1737 13.384
R9810 gnd.n3760 gnd.n3759 13.384
R9811 gnd.n4620 gnd.n4619 13.384
R9812 gnd.n4727 gnd.n3669 13.384
R9813 gnd.t157 gnd.n3659 13.384
R9814 gnd.n4758 gnd.t183 13.384
R9815 gnd.n4777 gnd.n3634 13.384
R9816 gnd.n4865 gnd.n3594 13.384
R9817 gnd.n4949 gnd.n4948 13.384
R9818 gnd.n2971 gnd.n2952 13.1884
R9819 gnd.n2966 gnd.n2965 13.1884
R9820 gnd.n2965 gnd.n2964 13.1884
R9821 gnd.n4977 gnd.n4972 13.1884
R9822 gnd.n4978 gnd.n4977 13.1884
R9823 gnd.n2967 gnd.n2954 13.146
R9824 gnd.n2963 gnd.n2954 13.146
R9825 gnd.n4976 gnd.n4975 13.146
R9826 gnd.n4976 gnd.n4971 13.146
R9827 gnd.n2296 gnd.n2292 12.8005
R9828 gnd.n2264 gnd.n2260 12.8005
R9829 gnd.n2232 gnd.n2228 12.8005
R9830 gnd.n2201 gnd.n2197 12.8005
R9831 gnd.n2169 gnd.n2165 12.8005
R9832 gnd.n2137 gnd.n2133 12.8005
R9833 gnd.n2105 gnd.n2101 12.8005
R9834 gnd.n2074 gnd.n2070 12.8005
R9835 gnd.n6128 gnd.n2496 12.7467
R9836 gnd.n4208 gnd.n4207 12.7467
R9837 gnd.n6122 gnd.n2506 12.7467
R9838 gnd.n6116 gnd.n2516 12.7467
R9839 gnd.n4195 gnd.n2519 12.7467
R9840 gnd.n6110 gnd.n2527 12.7467
R9841 gnd.n4189 gnd.n2530 12.7467
R9842 gnd.n6104 gnd.n2537 12.7467
R9843 gnd.n4240 gnd.n4239 12.7467
R9844 gnd.n4251 gnd.n4052 12.7467
R9845 gnd.n4259 gnd.n4046 12.7467
R9846 gnd.n4275 gnd.n4036 12.7467
R9847 gnd.n4281 gnd.n4029 12.7467
R9848 gnd.n4031 gnd.n4022 12.7467
R9849 gnd.n6096 gnd.n2552 12.7467
R9850 gnd.n4317 gnd.n2555 12.7467
R9851 gnd.n4325 gnd.n2566 12.7467
R9852 gnd.n6084 gnd.n2573 12.7467
R9853 gnd.n4331 gnd.n4010 12.7467
R9854 gnd.n6078 gnd.n2582 12.7467
R9855 gnd.n6072 gnd.n2593 12.7467
R9856 gnd.n4363 gnd.n2596 12.7467
R9857 gnd.n4346 gnd.n2605 12.7467
R9858 gnd.n6060 gnd.n2613 12.7467
R9859 gnd.n4352 gnd.n2616 12.7467
R9860 gnd.n6054 gnd.n2623 12.7467
R9861 gnd.n6041 gnd.n2640 12.7467
R9862 gnd.n6048 gnd.n2632 12.7467
R9863 gnd.n5528 gnd.n3269 12.7467
R9864 gnd.n5346 gnd.n5345 12.7467
R9865 gnd.n5520 gnd.n3278 12.7467
R9866 gnd.n5306 gnd.n3291 12.7467
R9867 gnd.n5514 gnd.n3294 12.7467
R9868 gnd.n5313 gnd.n3304 12.7467
R9869 gnd.n5319 gnd.n3314 12.7467
R9870 gnd.n5502 gnd.n3317 12.7467
R9871 gnd.n5496 gnd.n3327 12.7467
R9872 gnd.n5388 gnd.n5387 12.7467
R9873 gnd.n5490 gnd.n3337 12.7467
R9874 gnd.n5396 gnd.n3344 12.7467
R9875 gnd.n5403 gnd.n3351 12.7467
R9876 gnd.n5478 gnd.n3354 12.7467
R9877 gnd.n5472 gnd.n3364 12.7467
R9878 gnd.n5467 gnd.n5466 12.7467
R9879 gnd.n5424 gnd.n3390 12.7467
R9880 gnd.n5459 gnd.n3378 12.7467
R9881 gnd.n7413 gnd.n75 12.7467
R9882 gnd.n5452 gnd.n5451 12.7467
R9883 gnd.n5442 gnd.n90 12.7467
R9884 gnd.n7405 gnd.n93 12.7467
R9885 gnd.n7226 gnd.n7225 12.7467
R9886 gnd.n7399 gnd.n104 12.7467
R9887 gnd.n7233 gnd.n111 12.7467
R9888 gnd.n7241 gnd.n120 12.7467
R9889 gnd.n7387 gnd.n123 12.7467
R9890 gnd.n7248 gnd.n131 12.7467
R9891 gnd.n4290 gnd.t254 12.4281
R9892 gnd.n4421 gnd.t0 12.4281
R9893 gnd.n3470 gnd.t21 12.4281
R9894 gnd.t211 gnd.n3361 12.4281
R9895 gnd.n1709 gnd.n1706 12.4126
R9896 gnd.n6327 gnd.n1053 12.4126
R9897 gnd.n5908 gnd.n5845 12.1761
R9898 gnd.n5158 gnd.n5157 12.1761
R9899 gnd.n5965 gnd.n2738 12.1094
R9900 gnd.n4524 gnd.n3768 12.1094
R9901 gnd.n4655 gnd.n3699 12.1094
R9902 gnd.n4699 gnd.n3679 12.1094
R9903 gnd.n4829 gnd.n3619 12.1094
R9904 gnd.n4857 gnd.n4856 12.1094
R9905 gnd.n3540 gnd.t144 12.1094
R9906 gnd.n5161 gnd.t40 12.1094
R9907 gnd.n5649 gnd.n3199 12.1094
R9908 gnd.n2300 gnd.n2299 12.0247
R9909 gnd.n2268 gnd.n2267 12.0247
R9910 gnd.n2236 gnd.n2235 12.0247
R9911 gnd.n2205 gnd.n2204 12.0247
R9912 gnd.n2173 gnd.n2172 12.0247
R9913 gnd.n2141 gnd.n2140 12.0247
R9914 gnd.n2109 gnd.n2108 12.0247
R9915 gnd.n2078 gnd.n2077 12.0247
R9916 gnd.t241 gnd.n2479 11.7908
R9917 gnd.t268 gnd.n2585 11.7908
R9918 gnd.n6066 gnd.t223 11.7908
R9919 gnd.n5508 gnd.t229 11.7908
R9920 gnd.t231 gnd.n3324 11.7908
R9921 gnd.n7375 gnd.t215 11.7908
R9922 gnd.n4535 gnd.t3 11.4721
R9923 gnd.n3719 gnd.t33 11.4721
R9924 gnd.n4866 gnd.t29 11.4721
R9925 gnd.n4892 gnd.t182 11.4721
R9926 gnd.n2303 gnd.n2290 11.249
R9927 gnd.n2271 gnd.n2258 11.249
R9928 gnd.n2239 gnd.n2226 11.249
R9929 gnd.n2208 gnd.n2195 11.249
R9930 gnd.n2176 gnd.n2163 11.249
R9931 gnd.n2144 gnd.n2131 11.249
R9932 gnd.n2112 gnd.n2099 11.249
R9933 gnd.n2081 gnd.n2068 11.249
R9934 gnd.n1810 gnd.t180 11.1535
R9935 gnd.n4195 gnd.t266 11.1535
R9936 gnd.n6090 gnd.t263 11.1535
R9937 gnd.n5484 gnd.t213 11.1535
R9938 gnd.n7399 gnd.t221 11.1535
R9939 gnd.n4665 gnd.n3692 10.8348
R9940 gnd.n4837 gnd.n3611 10.8348
R9941 gnd.n3526 gnd.n3516 10.8348
R9942 gnd.n5539 gnd.n5536 10.6672
R9943 gnd.n379 gnd.n177 10.6672
R9944 gnd.n6163 gnd.n6160 10.6672
R9945 gnd.n2851 gnd.n2848 10.6672
R9946 gnd.n5093 gnd.n5015 10.6151
R9947 gnd.n5093 gnd.n5092 10.6151
R9948 gnd.n5090 gnd.n5019 10.6151
R9949 gnd.n5085 gnd.n5019 10.6151
R9950 gnd.n5085 gnd.n5084 10.6151
R9951 gnd.n5084 gnd.n5083 10.6151
R9952 gnd.n5083 gnd.n5022 10.6151
R9953 gnd.n5078 gnd.n5022 10.6151
R9954 gnd.n5078 gnd.n5077 10.6151
R9955 gnd.n5077 gnd.n5076 10.6151
R9956 gnd.n5076 gnd.n5025 10.6151
R9957 gnd.n5071 gnd.n5025 10.6151
R9958 gnd.n5071 gnd.n5070 10.6151
R9959 gnd.n5070 gnd.n5069 10.6151
R9960 gnd.n5069 gnd.n5028 10.6151
R9961 gnd.n5064 gnd.n5028 10.6151
R9962 gnd.n5064 gnd.n5063 10.6151
R9963 gnd.n5063 gnd.n5062 10.6151
R9964 gnd.n5062 gnd.n5031 10.6151
R9965 gnd.n5057 gnd.n5031 10.6151
R9966 gnd.n5057 gnd.n5056 10.6151
R9967 gnd.n5056 gnd.n5055 10.6151
R9968 gnd.n5055 gnd.n5034 10.6151
R9969 gnd.n5050 gnd.n5034 10.6151
R9970 gnd.n5050 gnd.n5049 10.6151
R9971 gnd.n5049 gnd.n5048 10.6151
R9972 gnd.n5048 gnd.n5037 10.6151
R9973 gnd.n5043 gnd.n5037 10.6151
R9974 gnd.n5043 gnd.n5042 10.6151
R9975 gnd.n5042 gnd.n5041 10.6151
R9976 gnd.n3839 gnd.n3838 10.6151
R9977 gnd.n3840 gnd.n3839 10.6151
R9978 gnd.n3840 gnd.n3771 10.6151
R9979 gnd.n3844 gnd.n3771 10.6151
R9980 gnd.n3845 gnd.n3844 10.6151
R9981 gnd.n3846 gnd.n3845 10.6151
R9982 gnd.n3846 gnd.n3757 10.6151
R9983 gnd.n4532 gnd.n3757 10.6151
R9984 gnd.n4533 gnd.n4532 10.6151
R9985 gnd.n4556 gnd.n4533 10.6151
R9986 gnd.n4556 gnd.n4555 10.6151
R9987 gnd.n4555 gnd.n4554 10.6151
R9988 gnd.n4554 gnd.n4553 10.6151
R9989 gnd.n4553 gnd.n4534 10.6151
R9990 gnd.n4547 gnd.n4534 10.6151
R9991 gnd.n4547 gnd.n4546 10.6151
R9992 gnd.n4546 gnd.n4545 10.6151
R9993 gnd.n4545 gnd.n4544 10.6151
R9994 gnd.n4544 gnd.n4542 10.6151
R9995 gnd.n4542 gnd.n4541 10.6151
R9996 gnd.n4541 gnd.n4539 10.6151
R9997 gnd.n4539 gnd.n4538 10.6151
R9998 gnd.n4538 gnd.n3711 10.6151
R9999 gnd.n4629 gnd.n3711 10.6151
R10000 gnd.n4630 gnd.n4629 10.6151
R10001 gnd.n4631 gnd.n4630 10.6151
R10002 gnd.n4646 gnd.n4631 10.6151
R10003 gnd.n4646 gnd.n4645 10.6151
R10004 gnd.n4645 gnd.n4644 10.6151
R10005 gnd.n4644 gnd.n4639 10.6151
R10006 gnd.n4639 gnd.n4638 10.6151
R10007 gnd.n4638 gnd.n4636 10.6151
R10008 gnd.n4636 gnd.n4635 10.6151
R10009 gnd.n4635 gnd.n4632 10.6151
R10010 gnd.n4632 gnd.n3661 10.6151
R10011 gnd.n4735 gnd.n3661 10.6151
R10012 gnd.n4736 gnd.n4735 10.6151
R10013 gnd.n4738 gnd.n4736 10.6151
R10014 gnd.n4738 gnd.n4737 10.6151
R10015 gnd.n4737 gnd.n3651 10.6151
R10016 gnd.n4750 gnd.n3651 10.6151
R10017 gnd.n4751 gnd.n4750 10.6151
R10018 gnd.n4755 gnd.n4751 10.6151
R10019 gnd.n4755 gnd.n4754 10.6151
R10020 gnd.n4754 gnd.n4753 10.6151
R10021 gnd.n4753 gnd.n3632 10.6151
R10022 gnd.n4780 gnd.n3632 10.6151
R10023 gnd.n4781 gnd.n4780 10.6151
R10024 gnd.n4783 gnd.n4781 10.6151
R10025 gnd.n4784 gnd.n4783 10.6151
R10026 gnd.n4785 gnd.n4784 10.6151
R10027 gnd.n4785 gnd.n3609 10.6151
R10028 gnd.n4840 gnd.n3609 10.6151
R10029 gnd.n4841 gnd.n4840 10.6151
R10030 gnd.n4847 gnd.n4841 10.6151
R10031 gnd.n4847 gnd.n4846 10.6151
R10032 gnd.n4846 gnd.n4845 10.6151
R10033 gnd.n4845 gnd.n4842 10.6151
R10034 gnd.n4842 gnd.n3586 10.6151
R10035 gnd.n4875 gnd.n3586 10.6151
R10036 gnd.n4876 gnd.n4875 10.6151
R10037 gnd.n4879 gnd.n4876 10.6151
R10038 gnd.n4879 gnd.n4878 10.6151
R10039 gnd.n4878 gnd.n4877 10.6151
R10040 gnd.n4877 gnd.n3567 10.6151
R10041 gnd.n4903 gnd.n3567 10.6151
R10042 gnd.n4904 gnd.n4903 10.6151
R10043 gnd.n4906 gnd.n4904 10.6151
R10044 gnd.n4907 gnd.n4906 10.6151
R10045 gnd.n4909 gnd.n4907 10.6151
R10046 gnd.n4909 gnd.n4908 10.6151
R10047 gnd.n4908 gnd.n3538 10.6151
R10048 gnd.n4958 gnd.n3538 10.6151
R10049 gnd.n4959 gnd.n4958 10.6151
R10050 gnd.n4960 gnd.n4959 10.6151
R10051 gnd.n4960 gnd.n3529 10.6151
R10052 gnd.n5166 gnd.n3529 10.6151
R10053 gnd.n5166 gnd.n5165 10.6151
R10054 gnd.n5165 gnd.n5164 10.6151
R10055 gnd.n5164 gnd.n3530 10.6151
R10056 gnd.n3774 gnd.n2912 10.6151
R10057 gnd.n3777 gnd.n3774 10.6151
R10058 gnd.n3782 gnd.n3779 10.6151
R10059 gnd.n3783 gnd.n3782 10.6151
R10060 gnd.n3786 gnd.n3783 10.6151
R10061 gnd.n3787 gnd.n3786 10.6151
R10062 gnd.n3790 gnd.n3787 10.6151
R10063 gnd.n3791 gnd.n3790 10.6151
R10064 gnd.n3794 gnd.n3791 10.6151
R10065 gnd.n3795 gnd.n3794 10.6151
R10066 gnd.n3798 gnd.n3795 10.6151
R10067 gnd.n3799 gnd.n3798 10.6151
R10068 gnd.n3802 gnd.n3799 10.6151
R10069 gnd.n3803 gnd.n3802 10.6151
R10070 gnd.n3806 gnd.n3803 10.6151
R10071 gnd.n3807 gnd.n3806 10.6151
R10072 gnd.n3810 gnd.n3807 10.6151
R10073 gnd.n3811 gnd.n3810 10.6151
R10074 gnd.n3814 gnd.n3811 10.6151
R10075 gnd.n3815 gnd.n3814 10.6151
R10076 gnd.n3818 gnd.n3815 10.6151
R10077 gnd.n3819 gnd.n3818 10.6151
R10078 gnd.n3822 gnd.n3819 10.6151
R10079 gnd.n3823 gnd.n3822 10.6151
R10080 gnd.n3826 gnd.n3823 10.6151
R10081 gnd.n3827 gnd.n3826 10.6151
R10082 gnd.n3830 gnd.n3827 10.6151
R10083 gnd.n3831 gnd.n3830 10.6151
R10084 gnd.n3834 gnd.n3831 10.6151
R10085 gnd.n3835 gnd.n3834 10.6151
R10086 gnd.n5908 gnd.n5907 10.6151
R10087 gnd.n5907 gnd.n5906 10.6151
R10088 gnd.n5906 gnd.n5905 10.6151
R10089 gnd.n5905 gnd.n5903 10.6151
R10090 gnd.n5903 gnd.n5900 10.6151
R10091 gnd.n5900 gnd.n5899 10.6151
R10092 gnd.n5899 gnd.n5896 10.6151
R10093 gnd.n5896 gnd.n5895 10.6151
R10094 gnd.n5895 gnd.n5892 10.6151
R10095 gnd.n5892 gnd.n5891 10.6151
R10096 gnd.n5891 gnd.n5888 10.6151
R10097 gnd.n5888 gnd.n5887 10.6151
R10098 gnd.n5887 gnd.n5884 10.6151
R10099 gnd.n5884 gnd.n5883 10.6151
R10100 gnd.n5883 gnd.n5880 10.6151
R10101 gnd.n5880 gnd.n5879 10.6151
R10102 gnd.n5879 gnd.n5876 10.6151
R10103 gnd.n5876 gnd.n5875 10.6151
R10104 gnd.n5875 gnd.n5872 10.6151
R10105 gnd.n5872 gnd.n5871 10.6151
R10106 gnd.n5871 gnd.n5868 10.6151
R10107 gnd.n5868 gnd.n5867 10.6151
R10108 gnd.n5867 gnd.n5864 10.6151
R10109 gnd.n5864 gnd.n5863 10.6151
R10110 gnd.n5863 gnd.n5860 10.6151
R10111 gnd.n5860 gnd.n5859 10.6151
R10112 gnd.n5859 gnd.n5856 10.6151
R10113 gnd.n5856 gnd.n5855 10.6151
R10114 gnd.n5852 gnd.n5851 10.6151
R10115 gnd.n5851 gnd.n2913 10.6151
R10116 gnd.n5157 gnd.n5156 10.6151
R10117 gnd.n5156 gnd.n4989 10.6151
R10118 gnd.n5151 gnd.n4989 10.6151
R10119 gnd.n5151 gnd.n5150 10.6151
R10120 gnd.n5150 gnd.n5149 10.6151
R10121 gnd.n5149 gnd.n4993 10.6151
R10122 gnd.n5144 gnd.n4993 10.6151
R10123 gnd.n5144 gnd.n5143 10.6151
R10124 gnd.n5143 gnd.n5142 10.6151
R10125 gnd.n5142 gnd.n4996 10.6151
R10126 gnd.n5137 gnd.n4996 10.6151
R10127 gnd.n5137 gnd.n5136 10.6151
R10128 gnd.n5136 gnd.n5135 10.6151
R10129 gnd.n5135 gnd.n4999 10.6151
R10130 gnd.n5130 gnd.n4999 10.6151
R10131 gnd.n5130 gnd.n5129 10.6151
R10132 gnd.n5129 gnd.n5128 10.6151
R10133 gnd.n5128 gnd.n5002 10.6151
R10134 gnd.n5123 gnd.n5002 10.6151
R10135 gnd.n5123 gnd.n5122 10.6151
R10136 gnd.n5122 gnd.n5121 10.6151
R10137 gnd.n5121 gnd.n5005 10.6151
R10138 gnd.n5116 gnd.n5005 10.6151
R10139 gnd.n5116 gnd.n5115 10.6151
R10140 gnd.n5115 gnd.n5114 10.6151
R10141 gnd.n5114 gnd.n5008 10.6151
R10142 gnd.n5109 gnd.n5008 10.6151
R10143 gnd.n5109 gnd.n5108 10.6151
R10144 gnd.n5106 gnd.n5013 10.6151
R10145 gnd.n5101 gnd.n5013 10.6151
R10146 gnd.n5844 gnd.n5843 10.6151
R10147 gnd.n5843 gnd.n2972 10.6151
R10148 gnd.n3764 gnd.n2972 10.6151
R10149 gnd.n3765 gnd.n3764 10.6151
R10150 gnd.n3765 gnd.n3762 10.6151
R10151 gnd.n4526 gnd.n3762 10.6151
R10152 gnd.n4527 gnd.n4526 10.6151
R10153 gnd.n4528 gnd.n4527 10.6151
R10154 gnd.n4528 gnd.n3752 10.6151
R10155 gnd.n4560 gnd.n3752 10.6151
R10156 gnd.n4561 gnd.n4560 10.6151
R10157 gnd.n4567 gnd.n4561 10.6151
R10158 gnd.n4567 gnd.n4566 10.6151
R10159 gnd.n4566 gnd.n4565 10.6151
R10160 gnd.n4565 gnd.n4562 10.6151
R10161 gnd.n4562 gnd.n3730 10.6151
R10162 gnd.n4606 gnd.n3730 10.6151
R10163 gnd.n4607 gnd.n4606 10.6151
R10164 gnd.n4608 gnd.n4607 10.6151
R10165 gnd.n4608 gnd.n3714 10.6151
R10166 gnd.n4622 gnd.n3714 10.6151
R10167 gnd.n4623 gnd.n4622 10.6151
R10168 gnd.n4624 gnd.n4623 10.6151
R10169 gnd.n4624 gnd.n3705 10.6151
R10170 gnd.n4652 gnd.n3705 10.6151
R10171 gnd.n4652 gnd.n4651 10.6151
R10172 gnd.n4651 gnd.n4650 10.6151
R10173 gnd.n4650 gnd.n3706 10.6151
R10174 gnd.n3706 gnd.n3683 10.6151
R10175 gnd.n4702 gnd.n3683 10.6151
R10176 gnd.n4703 gnd.n4702 10.6151
R10177 gnd.n4704 gnd.n4703 10.6151
R10178 gnd.n4704 gnd.n3667 10.6151
R10179 gnd.n4729 gnd.n3667 10.6151
R10180 gnd.n4730 gnd.n4729 10.6151
R10181 gnd.n4731 gnd.n4730 10.6151
R10182 gnd.n4731 gnd.n3657 10.6151
R10183 gnd.n4743 gnd.n3657 10.6151
R10184 gnd.n4744 gnd.n4743 10.6151
R10185 gnd.n4745 gnd.n4744 10.6151
R10186 gnd.n4745 gnd.n3646 10.6151
R10187 gnd.n4761 gnd.n3646 10.6151
R10188 gnd.n4762 gnd.n4761 10.6151
R10189 gnd.n4766 gnd.n4762 10.6151
R10190 gnd.n4766 gnd.n4765 10.6151
R10191 gnd.n4765 gnd.n4764 10.6151
R10192 gnd.n4764 gnd.n3624 10.6151
R10193 gnd.n4821 gnd.n3624 10.6151
R10194 gnd.n4822 gnd.n4821 10.6151
R10195 gnd.n4826 gnd.n4822 10.6151
R10196 gnd.n4826 gnd.n4825 10.6151
R10197 gnd.n4825 gnd.n4824 10.6151
R10198 gnd.n4824 gnd.n3605 10.6151
R10199 gnd.n4852 gnd.n3605 10.6151
R10200 gnd.n4853 gnd.n4852 10.6151
R10201 gnd.n4854 gnd.n4853 10.6151
R10202 gnd.n4854 gnd.n3590 10.6151
R10203 gnd.n4868 gnd.n3590 10.6151
R10204 gnd.n4869 gnd.n4868 10.6151
R10205 gnd.n4871 gnd.n4869 10.6151
R10206 gnd.n4871 gnd.n4870 10.6151
R10207 gnd.n4870 gnd.n3571 10.6151
R10208 gnd.n4896 gnd.n3571 10.6151
R10209 gnd.n4897 gnd.n4896 10.6151
R10210 gnd.n4898 gnd.n4897 10.6151
R10211 gnd.n4898 gnd.n3558 10.6151
R10212 gnd.n4933 gnd.n3558 10.6151
R10213 gnd.n4934 gnd.n4933 10.6151
R10214 gnd.n4935 gnd.n4934 10.6151
R10215 gnd.n4935 gnd.n3543 10.6151
R10216 gnd.n4951 gnd.n3543 10.6151
R10217 gnd.n4952 gnd.n4951 10.6151
R10218 gnd.n4954 gnd.n4952 10.6151
R10219 gnd.n4954 gnd.n4953 10.6151
R10220 gnd.n4953 gnd.n3535 10.6151
R10221 gnd.n4965 gnd.n3535 10.6151
R10222 gnd.n4966 gnd.n4965 10.6151
R10223 gnd.n4968 gnd.n4966 10.6151
R10224 gnd.n4969 gnd.n4968 10.6151
R10225 gnd.n5159 gnd.n4969 10.6151
R10226 gnd.n1381 gnd.t160 10.5161
R10227 gnd.n1998 gnd.t207 10.5161
R10228 gnd.t25 gnd.n1015 10.5161
R10229 gnd.n4248 gnd.t219 10.5161
R10230 gnd.n4275 gnd.t225 10.5161
R10231 gnd.n5424 gnd.t252 10.5161
R10232 gnd.n5458 gnd.t258 10.5161
R10233 gnd.n2304 gnd.n2288 10.4732
R10234 gnd.n2272 gnd.n2256 10.4732
R10235 gnd.n2240 gnd.n2224 10.4732
R10236 gnd.n2209 gnd.n2193 10.4732
R10237 gnd.n2177 gnd.n2161 10.4732
R10238 gnd.n2145 gnd.n2129 10.4732
R10239 gnd.n2113 gnd.n2097 10.4732
R10240 gnd.n2082 gnd.n2066 10.4732
R10241 gnd.n4626 gnd.t33 10.1975
R10242 gnd.n4843 gnd.t29 10.1975
R10243 gnd.n2039 gnd.t167 9.87883
R10244 gnd.n4201 gnd.t248 9.87883
R10245 gnd.n6084 gnd.t279 9.87883
R10246 gnd.n5490 gnd.t239 9.87883
R10247 gnd.n7393 gnd.t227 9.87883
R10248 gnd.n2308 gnd.n2307 9.69747
R10249 gnd.n2276 gnd.n2275 9.69747
R10250 gnd.n2244 gnd.n2243 9.69747
R10251 gnd.n2213 gnd.n2212 9.69747
R10252 gnd.n2181 gnd.n2180 9.69747
R10253 gnd.n2149 gnd.n2148 9.69747
R10254 gnd.n2117 gnd.n2116 9.69747
R10255 gnd.n2086 gnd.n2085 9.69747
R10256 gnd.n3769 gnd.n3768 9.56018
R10257 gnd.n4603 gnd.t8 9.56018
R10258 gnd.n4700 gnd.n4699 9.56018
R10259 gnd.n4829 gnd.n4828 9.56018
R10260 gnd.t2 gnd.n3573 9.56018
R10261 gnd.n4962 gnd.t144 9.56018
R10262 gnd.t40 gnd.n3517 9.56018
R10263 gnd.n5161 gnd.n3532 9.56018
R10264 gnd.n2314 gnd.n2313 9.45567
R10265 gnd.n2282 gnd.n2281 9.45567
R10266 gnd.n2250 gnd.n2249 9.45567
R10267 gnd.n2219 gnd.n2218 9.45567
R10268 gnd.n2187 gnd.n2186 9.45567
R10269 gnd.n2155 gnd.n2154 9.45567
R10270 gnd.n2123 gnd.n2122 9.45567
R10271 gnd.n2092 gnd.n2091 9.45567
R10272 gnd.n5576 gnd.n5575 9.30959
R10273 gnd.n335 gnd.n199 9.30959
R10274 gnd.n6200 gnd.n6199 9.30959
R10275 gnd.n2890 gnd.n2822 9.30959
R10276 gnd.n2313 gnd.n2312 9.3005
R10277 gnd.n2286 gnd.n2285 9.3005
R10278 gnd.n2307 gnd.n2306 9.3005
R10279 gnd.n2305 gnd.n2304 9.3005
R10280 gnd.n2290 gnd.n2289 9.3005
R10281 gnd.n2299 gnd.n2298 9.3005
R10282 gnd.n2297 gnd.n2296 9.3005
R10283 gnd.n2281 gnd.n2280 9.3005
R10284 gnd.n2254 gnd.n2253 9.3005
R10285 gnd.n2275 gnd.n2274 9.3005
R10286 gnd.n2273 gnd.n2272 9.3005
R10287 gnd.n2258 gnd.n2257 9.3005
R10288 gnd.n2267 gnd.n2266 9.3005
R10289 gnd.n2265 gnd.n2264 9.3005
R10290 gnd.n2249 gnd.n2248 9.3005
R10291 gnd.n2222 gnd.n2221 9.3005
R10292 gnd.n2243 gnd.n2242 9.3005
R10293 gnd.n2241 gnd.n2240 9.3005
R10294 gnd.n2226 gnd.n2225 9.3005
R10295 gnd.n2235 gnd.n2234 9.3005
R10296 gnd.n2233 gnd.n2232 9.3005
R10297 gnd.n2218 gnd.n2217 9.3005
R10298 gnd.n2191 gnd.n2190 9.3005
R10299 gnd.n2212 gnd.n2211 9.3005
R10300 gnd.n2210 gnd.n2209 9.3005
R10301 gnd.n2195 gnd.n2194 9.3005
R10302 gnd.n2204 gnd.n2203 9.3005
R10303 gnd.n2202 gnd.n2201 9.3005
R10304 gnd.n2186 gnd.n2185 9.3005
R10305 gnd.n2159 gnd.n2158 9.3005
R10306 gnd.n2180 gnd.n2179 9.3005
R10307 gnd.n2178 gnd.n2177 9.3005
R10308 gnd.n2163 gnd.n2162 9.3005
R10309 gnd.n2172 gnd.n2171 9.3005
R10310 gnd.n2170 gnd.n2169 9.3005
R10311 gnd.n2154 gnd.n2153 9.3005
R10312 gnd.n2127 gnd.n2126 9.3005
R10313 gnd.n2148 gnd.n2147 9.3005
R10314 gnd.n2146 gnd.n2145 9.3005
R10315 gnd.n2131 gnd.n2130 9.3005
R10316 gnd.n2140 gnd.n2139 9.3005
R10317 gnd.n2138 gnd.n2137 9.3005
R10318 gnd.n2122 gnd.n2121 9.3005
R10319 gnd.n2095 gnd.n2094 9.3005
R10320 gnd.n2116 gnd.n2115 9.3005
R10321 gnd.n2114 gnd.n2113 9.3005
R10322 gnd.n2099 gnd.n2098 9.3005
R10323 gnd.n2108 gnd.n2107 9.3005
R10324 gnd.n2106 gnd.n2105 9.3005
R10325 gnd.n2091 gnd.n2090 9.3005
R10326 gnd.n2064 gnd.n2063 9.3005
R10327 gnd.n2085 gnd.n2084 9.3005
R10328 gnd.n2083 gnd.n2082 9.3005
R10329 gnd.n2068 gnd.n2067 9.3005
R10330 gnd.n2077 gnd.n2076 9.3005
R10331 gnd.n2075 gnd.n2074 9.3005
R10332 gnd.n6320 gnd.n6319 9.3005
R10333 gnd.n6318 gnd.n6286 9.3005
R10334 gnd.n6317 gnd.n6316 9.3005
R10335 gnd.n6313 gnd.n6287 9.3005
R10336 gnd.n6310 gnd.n6288 9.3005
R10337 gnd.n6309 gnd.n6289 9.3005
R10338 gnd.n6306 gnd.n6290 9.3005
R10339 gnd.n6305 gnd.n6291 9.3005
R10340 gnd.n6302 gnd.n6292 9.3005
R10341 gnd.n6301 gnd.n6293 9.3005
R10342 gnd.n6298 gnd.n6294 9.3005
R10343 gnd.n6297 gnd.n6295 9.3005
R10344 gnd.n1055 gnd.n1054 9.3005
R10345 gnd.n6328 gnd.n6327 9.3005
R10346 gnd.n6329 gnd.n1053 9.3005
R10347 gnd.n6331 gnd.n6330 9.3005
R10348 gnd.n6321 gnd.n6285 9.3005
R10349 gnd.n1762 gnd.n1761 9.3005
R10350 gnd.n1763 gnd.n1352 9.3005
R10351 gnd.n1767 gnd.n1764 9.3005
R10352 gnd.n1766 gnd.n1765 9.3005
R10353 gnd.n1329 gnd.n1328 9.3005
R10354 gnd.n1793 gnd.n1792 9.3005
R10355 gnd.n1794 gnd.n1327 9.3005
R10356 gnd.n1798 gnd.n1795 9.3005
R10357 gnd.n1797 gnd.n1796 9.3005
R10358 gnd.n1303 gnd.n1302 9.3005
R10359 gnd.n1824 gnd.n1823 9.3005
R10360 gnd.n1825 gnd.n1301 9.3005
R10361 gnd.n1829 gnd.n1826 9.3005
R10362 gnd.n1828 gnd.n1827 9.3005
R10363 gnd.n1277 gnd.n1276 9.3005
R10364 gnd.n1855 gnd.n1854 9.3005
R10365 gnd.n1856 gnd.n1275 9.3005
R10366 gnd.n1860 gnd.n1857 9.3005
R10367 gnd.n1859 gnd.n1858 9.3005
R10368 gnd.n1251 gnd.n1250 9.3005
R10369 gnd.n1886 gnd.n1885 9.3005
R10370 gnd.n1887 gnd.n1249 9.3005
R10371 gnd.n1891 gnd.n1888 9.3005
R10372 gnd.n1890 gnd.n1889 9.3005
R10373 gnd.n1226 gnd.n1225 9.3005
R10374 gnd.n1917 gnd.n1916 9.3005
R10375 gnd.n1918 gnd.n1224 9.3005
R10376 gnd.n1922 gnd.n1919 9.3005
R10377 gnd.n1921 gnd.n1920 9.3005
R10378 gnd.n1199 gnd.n1198 9.3005
R10379 gnd.n1947 gnd.n1946 9.3005
R10380 gnd.n1948 gnd.n1197 9.3005
R10381 gnd.n1950 gnd.n1949 9.3005
R10382 gnd.n1177 gnd.n1176 9.3005
R10383 gnd.n2017 gnd.n2016 9.3005
R10384 gnd.n2018 gnd.n1175 9.3005
R10385 gnd.n2023 gnd.n2019 9.3005
R10386 gnd.n2022 gnd.n2021 9.3005
R10387 gnd.n2020 gnd.n983 9.3005
R10388 gnd.n6372 gnd.n984 9.3005
R10389 gnd.n6371 gnd.n985 9.3005
R10390 gnd.n6370 gnd.n986 9.3005
R10391 gnd.n1008 gnd.n987 9.3005
R10392 gnd.n1009 gnd.n1007 9.3005
R10393 gnd.n6358 gnd.n1010 9.3005
R10394 gnd.n6357 gnd.n1011 9.3005
R10395 gnd.n6356 gnd.n1012 9.3005
R10396 gnd.n1033 gnd.n1013 9.3005
R10397 gnd.n1034 gnd.n1032 9.3005
R10398 gnd.n6344 gnd.n1035 9.3005
R10399 gnd.n6343 gnd.n1036 9.3005
R10400 gnd.n6342 gnd.n1037 9.3005
R10401 gnd.n6284 gnd.n1038 9.3005
R10402 gnd.n1354 gnd.n1353 9.3005
R10403 gnd.n1706 gnd.n1705 9.3005
R10404 gnd.n1709 gnd.n1701 9.3005
R10405 gnd.n1710 gnd.n1700 9.3005
R10406 gnd.n1713 gnd.n1699 9.3005
R10407 gnd.n1714 gnd.n1698 9.3005
R10408 gnd.n1717 gnd.n1697 9.3005
R10409 gnd.n1718 gnd.n1696 9.3005
R10410 gnd.n1721 gnd.n1695 9.3005
R10411 gnd.n1722 gnd.n1694 9.3005
R10412 gnd.n1725 gnd.n1693 9.3005
R10413 gnd.n1726 gnd.n1692 9.3005
R10414 gnd.n1729 gnd.n1691 9.3005
R10415 gnd.n1731 gnd.n1690 9.3005
R10416 gnd.n1732 gnd.n1689 9.3005
R10417 gnd.n1733 gnd.n1688 9.3005
R10418 gnd.n1734 gnd.n1687 9.3005
R10419 gnd.n1702 gnd.n1370 9.3005
R10420 gnd.n1752 gnd.n1751 9.3005
R10421 gnd.n1753 gnd.n1347 9.3005
R10422 gnd.n1772 gnd.n1771 9.3005
R10423 gnd.n1774 gnd.n1339 9.3005
R10424 gnd.n1781 gnd.n1340 9.3005
R10425 gnd.n1783 gnd.n1782 9.3005
R10426 gnd.n1784 gnd.n1320 9.3005
R10427 gnd.n1803 gnd.n1802 9.3005
R10428 gnd.n1805 gnd.n1313 9.3005
R10429 gnd.n1812 gnd.n1314 9.3005
R10430 gnd.n1814 gnd.n1813 9.3005
R10431 gnd.n1815 gnd.n1294 9.3005
R10432 gnd.n1834 gnd.n1833 9.3005
R10433 gnd.n1836 gnd.n1287 9.3005
R10434 gnd.n1843 gnd.n1288 9.3005
R10435 gnd.n1845 gnd.n1844 9.3005
R10436 gnd.n1846 gnd.n1269 9.3005
R10437 gnd.n1865 gnd.n1864 9.3005
R10438 gnd.n1867 gnd.n1261 9.3005
R10439 gnd.n1874 gnd.n1262 9.3005
R10440 gnd.n1876 gnd.n1875 9.3005
R10441 gnd.n1877 gnd.n1244 9.3005
R10442 gnd.n1896 gnd.n1895 9.3005
R10443 gnd.n1898 gnd.n1236 9.3005
R10444 gnd.n1905 gnd.n1237 9.3005
R10445 gnd.n1907 gnd.n1906 9.3005
R10446 gnd.n1908 gnd.n1219 9.3005
R10447 gnd.n1927 gnd.n1926 9.3005
R10448 gnd.n1929 gnd.n1210 9.3005
R10449 gnd.n1936 gnd.n1212 9.3005
R10450 gnd.n1937 gnd.n1207 9.3005
R10451 gnd.n1939 gnd.n1938 9.3005
R10452 gnd.n1208 gnd.n1193 9.3005
R10453 gnd.n1955 gnd.n1191 9.3005
R10454 gnd.n1961 gnd.n1960 9.3005
R10455 gnd.n1959 gnd.n1956 9.3005
R10456 gnd.n1957 gnd.n1164 9.3005
R10457 gnd.n2031 gnd.n1163 9.3005
R10458 gnd.n2036 gnd.n2034 9.3005
R10459 gnd.n2035 gnd.n1157 9.3005
R10460 gnd.n2045 gnd.n1156 9.3005
R10461 gnd.n2048 gnd.n2047 9.3005
R10462 gnd.n2050 gnd.n2049 9.3005
R10463 gnd.n2054 gnd.n2051 9.3005
R10464 gnd.n2056 gnd.n2055 9.3005
R10465 gnd.n2058 gnd.n1153 9.3005
R10466 gnd.n2061 gnd.n2060 9.3005
R10467 gnd.n2319 gnd.n2318 9.3005
R10468 gnd.n2323 gnd.n2320 9.3005
R10469 gnd.n2325 gnd.n2324 9.3005
R10470 gnd.n2329 gnd.n2328 9.3005
R10471 gnd.n1049 gnd.n1047 9.3005
R10472 gnd.n6335 gnd.n6334 9.3005
R10473 gnd.n1750 gnd.n1364 9.3005
R10474 gnd.n1089 gnd.n1086 9.3005
R10475 gnd.n1091 gnd.n1090 9.3005
R10476 gnd.n1094 gnd.n1084 9.3005
R10477 gnd.n1098 gnd.n1097 9.3005
R10478 gnd.n1099 gnd.n1083 9.3005
R10479 gnd.n1101 gnd.n1100 9.3005
R10480 gnd.n1104 gnd.n1082 9.3005
R10481 gnd.n1108 gnd.n1107 9.3005
R10482 gnd.n1109 gnd.n1081 9.3005
R10483 gnd.n1111 gnd.n1110 9.3005
R10484 gnd.n1114 gnd.n1080 9.3005
R10485 gnd.n1118 gnd.n1117 9.3005
R10486 gnd.n1119 gnd.n1079 9.3005
R10487 gnd.n1121 gnd.n1120 9.3005
R10488 gnd.n1124 gnd.n1078 9.3005
R10489 gnd.n1128 gnd.n1127 9.3005
R10490 gnd.n1129 gnd.n1077 9.3005
R10491 gnd.n1131 gnd.n1130 9.3005
R10492 gnd.n1134 gnd.n1076 9.3005
R10493 gnd.n1138 gnd.n1137 9.3005
R10494 gnd.n1139 gnd.n1075 9.3005
R10495 gnd.n1141 gnd.n1140 9.3005
R10496 gnd.n1144 gnd.n1071 9.3005
R10497 gnd.n1147 gnd.n1146 9.3005
R10498 gnd.n1148 gnd.n1070 9.3005
R10499 gnd.n2339 gnd.n2338 9.3005
R10500 gnd.n1088 gnd.n1087 9.3005
R10501 gnd.n1581 gnd.n1560 9.3005
R10502 gnd.n1580 gnd.n1562 9.3005
R10503 gnd.n1578 gnd.n1563 9.3005
R10504 gnd.n1577 gnd.n1564 9.3005
R10505 gnd.n1573 gnd.n1565 9.3005
R10506 gnd.n1572 gnd.n1566 9.3005
R10507 gnd.n1571 gnd.n1567 9.3005
R10508 gnd.n1569 gnd.n1568 9.3005
R10509 gnd.n1184 gnd.n1183 9.3005
R10510 gnd.n1969 gnd.n1968 9.3005
R10511 gnd.n1970 gnd.n1182 9.3005
R10512 gnd.n2011 gnd.n1971 9.3005
R10513 gnd.n2010 gnd.n1972 9.3005
R10514 gnd.n2009 gnd.n1973 9.3005
R10515 gnd.n2007 gnd.n1974 9.3005
R10516 gnd.n2006 gnd.n1975 9.3005
R10517 gnd.n1977 gnd.n1976 9.3005
R10518 gnd.n2002 gnd.n1978 9.3005
R10519 gnd.n2001 gnd.n1979 9.3005
R10520 gnd.n2000 gnd.n1980 9.3005
R10521 gnd.n1997 gnd.n1981 9.3005
R10522 gnd.n1996 gnd.n1982 9.3005
R10523 gnd.n1993 gnd.n1983 9.3005
R10524 gnd.n1992 gnd.n1984 9.3005
R10525 gnd.n1991 gnd.n1985 9.3005
R10526 gnd.n1988 gnd.n1987 9.3005
R10527 gnd.n1986 gnd.n1150 9.3005
R10528 gnd.n2335 gnd.n1149 9.3005
R10529 gnd.n2337 gnd.n2336 9.3005
R10530 gnd.n1507 gnd.n1401 9.3005
R10531 gnd.n1509 gnd.n1508 9.3005
R10532 gnd.n1391 gnd.n1390 9.3005
R10533 gnd.n1522 gnd.n1521 9.3005
R10534 gnd.n1523 gnd.n1389 9.3005
R10535 gnd.n1525 gnd.n1524 9.3005
R10536 gnd.n1378 gnd.n1377 9.3005
R10537 gnd.n1538 gnd.n1537 9.3005
R10538 gnd.n1539 gnd.n1376 9.3005
R10539 gnd.n1676 gnd.n1540 9.3005
R10540 gnd.n1675 gnd.n1541 9.3005
R10541 gnd.n1674 gnd.n1542 9.3005
R10542 gnd.n1673 gnd.n1543 9.3005
R10543 gnd.n1671 gnd.n1544 9.3005
R10544 gnd.n1670 gnd.n1545 9.3005
R10545 gnd.n1666 gnd.n1546 9.3005
R10546 gnd.n1665 gnd.n1547 9.3005
R10547 gnd.n1664 gnd.n1548 9.3005
R10548 gnd.n1662 gnd.n1549 9.3005
R10549 gnd.n1661 gnd.n1550 9.3005
R10550 gnd.n1658 gnd.n1551 9.3005
R10551 gnd.n1657 gnd.n1552 9.3005
R10552 gnd.n1656 gnd.n1553 9.3005
R10553 gnd.n1654 gnd.n1554 9.3005
R10554 gnd.n1653 gnd.n1555 9.3005
R10555 gnd.n1650 gnd.n1556 9.3005
R10556 gnd.n1649 gnd.n1557 9.3005
R10557 gnd.n1648 gnd.n1558 9.3005
R10558 gnd.n1506 gnd.n1505 9.3005
R10559 gnd.n1446 gnd.n1445 9.3005
R10560 gnd.n1451 gnd.n1443 9.3005
R10561 gnd.n1452 gnd.n1442 9.3005
R10562 gnd.n1454 gnd.n1439 9.3005
R10563 gnd.n1438 gnd.n1436 9.3005
R10564 gnd.n1460 gnd.n1435 9.3005
R10565 gnd.n1461 gnd.n1434 9.3005
R10566 gnd.n1462 gnd.n1433 9.3005
R10567 gnd.n1432 gnd.n1430 9.3005
R10568 gnd.n1468 gnd.n1429 9.3005
R10569 gnd.n1469 gnd.n1428 9.3005
R10570 gnd.n1470 gnd.n1427 9.3005
R10571 gnd.n1426 gnd.n1424 9.3005
R10572 gnd.n1476 gnd.n1423 9.3005
R10573 gnd.n1477 gnd.n1422 9.3005
R10574 gnd.n1478 gnd.n1421 9.3005
R10575 gnd.n1420 gnd.n1418 9.3005
R10576 gnd.n1484 gnd.n1417 9.3005
R10577 gnd.n1485 gnd.n1416 9.3005
R10578 gnd.n1486 gnd.n1415 9.3005
R10579 gnd.n1414 gnd.n1412 9.3005
R10580 gnd.n1491 gnd.n1411 9.3005
R10581 gnd.n1492 gnd.n1410 9.3005
R10582 gnd.n1409 gnd.n1407 9.3005
R10583 gnd.n1497 gnd.n1406 9.3005
R10584 gnd.n1499 gnd.n1498 9.3005
R10585 gnd.n1444 gnd.n1402 9.3005
R10586 gnd.n1397 gnd.n1396 9.3005
R10587 gnd.n1514 gnd.n1513 9.3005
R10588 gnd.n1515 gnd.n1395 9.3005
R10589 gnd.n1517 gnd.n1516 9.3005
R10590 gnd.n1385 gnd.n1384 9.3005
R10591 gnd.n1530 gnd.n1529 9.3005
R10592 gnd.n1531 gnd.n1383 9.3005
R10593 gnd.n1533 gnd.n1532 9.3005
R10594 gnd.n1372 gnd.n1371 9.3005
R10595 gnd.n1741 gnd.n1740 9.3005
R10596 gnd.n1743 gnd.n1369 9.3005
R10597 gnd.n1745 gnd.n1744 9.3005
R10598 gnd.n1363 gnd.n1362 9.3005
R10599 gnd.n1756 gnd.n1754 9.3005
R10600 gnd.n1755 gnd.n1346 9.3005
R10601 gnd.n1773 gnd.n1345 9.3005
R10602 gnd.n1776 gnd.n1775 9.3005
R10603 gnd.n1338 gnd.n1337 9.3005
R10604 gnd.n1787 gnd.n1785 9.3005
R10605 gnd.n1786 gnd.n1319 9.3005
R10606 gnd.n1804 gnd.n1318 9.3005
R10607 gnd.n1807 gnd.n1806 9.3005
R10608 gnd.n1312 gnd.n1311 9.3005
R10609 gnd.n1818 gnd.n1816 9.3005
R10610 gnd.n1817 gnd.n1293 9.3005
R10611 gnd.n1835 gnd.n1292 9.3005
R10612 gnd.n1838 gnd.n1837 9.3005
R10613 gnd.n1286 gnd.n1285 9.3005
R10614 gnd.n1849 gnd.n1847 9.3005
R10615 gnd.n1848 gnd.n1268 9.3005
R10616 gnd.n1866 gnd.n1267 9.3005
R10617 gnd.n1869 gnd.n1868 9.3005
R10618 gnd.n1260 gnd.n1259 9.3005
R10619 gnd.n1880 gnd.n1878 9.3005
R10620 gnd.n1879 gnd.n1243 9.3005
R10621 gnd.n1897 gnd.n1242 9.3005
R10622 gnd.n1900 gnd.n1899 9.3005
R10623 gnd.n1235 gnd.n1234 9.3005
R10624 gnd.n1911 gnd.n1909 9.3005
R10625 gnd.n1910 gnd.n1218 9.3005
R10626 gnd.n1928 gnd.n1217 9.3005
R10627 gnd.n1931 gnd.n1930 9.3005
R10628 gnd.n1211 gnd.n1206 9.3005
R10629 gnd.n1941 gnd.n1940 9.3005
R10630 gnd.n1209 gnd.n1189 9.3005
R10631 gnd.n1964 gnd.n1190 9.3005
R10632 gnd.n1963 gnd.n1962 9.3005
R10633 gnd.n1192 gnd.n1165 9.3005
R10634 gnd.n2028 gnd.n1166 9.3005
R10635 gnd.n2030 gnd.n2029 9.3005
R10636 gnd.n2032 gnd.n1160 9.3005
R10637 gnd.n2033 gnd.n1158 9.3005
R10638 gnd.n2044 gnd.n2043 9.3005
R10639 gnd.n2046 gnd.n995 9.3005
R10640 gnd.n6365 gnd.n996 9.3005
R10641 gnd.n6364 gnd.n997 9.3005
R10642 gnd.n6363 gnd.n998 9.3005
R10643 gnd.n2057 gnd.n999 9.3005
R10644 gnd.n2059 gnd.n1021 9.3005
R10645 gnd.n6351 gnd.n1022 9.3005
R10646 gnd.n6350 gnd.n1023 9.3005
R10647 gnd.n6349 gnd.n1024 9.3005
R10648 gnd.n2326 gnd.n1025 9.3005
R10649 gnd.n2327 gnd.n1046 9.3005
R10650 gnd.n6337 gnd.n6336 9.3005
R10651 gnd.n1501 gnd.n1500 9.3005
R10652 gnd.n6547 gnd.n6546 9.3005
R10653 gnd.n6548 gnd.n807 9.3005
R10654 gnd.n6550 gnd.n6549 9.3005
R10655 gnd.n803 gnd.n802 9.3005
R10656 gnd.n6557 gnd.n6556 9.3005
R10657 gnd.n6558 gnd.n801 9.3005
R10658 gnd.n6560 gnd.n6559 9.3005
R10659 gnd.n797 gnd.n796 9.3005
R10660 gnd.n6567 gnd.n6566 9.3005
R10661 gnd.n6568 gnd.n795 9.3005
R10662 gnd.n6570 gnd.n6569 9.3005
R10663 gnd.n791 gnd.n790 9.3005
R10664 gnd.n6577 gnd.n6576 9.3005
R10665 gnd.n6578 gnd.n789 9.3005
R10666 gnd.n6580 gnd.n6579 9.3005
R10667 gnd.n785 gnd.n784 9.3005
R10668 gnd.n6587 gnd.n6586 9.3005
R10669 gnd.n6588 gnd.n783 9.3005
R10670 gnd.n6590 gnd.n6589 9.3005
R10671 gnd.n779 gnd.n778 9.3005
R10672 gnd.n6597 gnd.n6596 9.3005
R10673 gnd.n6598 gnd.n777 9.3005
R10674 gnd.n6600 gnd.n6599 9.3005
R10675 gnd.n773 gnd.n772 9.3005
R10676 gnd.n6607 gnd.n6606 9.3005
R10677 gnd.n6608 gnd.n771 9.3005
R10678 gnd.n6610 gnd.n6609 9.3005
R10679 gnd.n767 gnd.n766 9.3005
R10680 gnd.n6617 gnd.n6616 9.3005
R10681 gnd.n6618 gnd.n765 9.3005
R10682 gnd.n6620 gnd.n6619 9.3005
R10683 gnd.n761 gnd.n760 9.3005
R10684 gnd.n6627 gnd.n6626 9.3005
R10685 gnd.n6628 gnd.n759 9.3005
R10686 gnd.n6630 gnd.n6629 9.3005
R10687 gnd.n755 gnd.n754 9.3005
R10688 gnd.n6637 gnd.n6636 9.3005
R10689 gnd.n6638 gnd.n753 9.3005
R10690 gnd.n6640 gnd.n6639 9.3005
R10691 gnd.n749 gnd.n748 9.3005
R10692 gnd.n6647 gnd.n6646 9.3005
R10693 gnd.n6648 gnd.n747 9.3005
R10694 gnd.n6650 gnd.n6649 9.3005
R10695 gnd.n743 gnd.n742 9.3005
R10696 gnd.n6657 gnd.n6656 9.3005
R10697 gnd.n6658 gnd.n741 9.3005
R10698 gnd.n6660 gnd.n6659 9.3005
R10699 gnd.n737 gnd.n736 9.3005
R10700 gnd.n6667 gnd.n6666 9.3005
R10701 gnd.n6668 gnd.n735 9.3005
R10702 gnd.n6670 gnd.n6669 9.3005
R10703 gnd.n731 gnd.n730 9.3005
R10704 gnd.n6677 gnd.n6676 9.3005
R10705 gnd.n6678 gnd.n729 9.3005
R10706 gnd.n6680 gnd.n6679 9.3005
R10707 gnd.n725 gnd.n724 9.3005
R10708 gnd.n6687 gnd.n6686 9.3005
R10709 gnd.n6688 gnd.n723 9.3005
R10710 gnd.n6690 gnd.n6689 9.3005
R10711 gnd.n719 gnd.n718 9.3005
R10712 gnd.n6697 gnd.n6696 9.3005
R10713 gnd.n6698 gnd.n717 9.3005
R10714 gnd.n6700 gnd.n6699 9.3005
R10715 gnd.n713 gnd.n712 9.3005
R10716 gnd.n6707 gnd.n6706 9.3005
R10717 gnd.n6708 gnd.n711 9.3005
R10718 gnd.n6710 gnd.n6709 9.3005
R10719 gnd.n707 gnd.n706 9.3005
R10720 gnd.n6717 gnd.n6716 9.3005
R10721 gnd.n6718 gnd.n705 9.3005
R10722 gnd.n6720 gnd.n6719 9.3005
R10723 gnd.n701 gnd.n700 9.3005
R10724 gnd.n6727 gnd.n6726 9.3005
R10725 gnd.n6728 gnd.n699 9.3005
R10726 gnd.n6730 gnd.n6729 9.3005
R10727 gnd.n695 gnd.n694 9.3005
R10728 gnd.n6737 gnd.n6736 9.3005
R10729 gnd.n6738 gnd.n693 9.3005
R10730 gnd.n6740 gnd.n6739 9.3005
R10731 gnd.n689 gnd.n688 9.3005
R10732 gnd.n6747 gnd.n6746 9.3005
R10733 gnd.n6748 gnd.n687 9.3005
R10734 gnd.n6750 gnd.n6749 9.3005
R10735 gnd.n683 gnd.n682 9.3005
R10736 gnd.n6757 gnd.n6756 9.3005
R10737 gnd.n6758 gnd.n681 9.3005
R10738 gnd.n6760 gnd.n6759 9.3005
R10739 gnd.n677 gnd.n676 9.3005
R10740 gnd.n6767 gnd.n6766 9.3005
R10741 gnd.n6768 gnd.n675 9.3005
R10742 gnd.n6770 gnd.n6769 9.3005
R10743 gnd.n671 gnd.n670 9.3005
R10744 gnd.n6777 gnd.n6776 9.3005
R10745 gnd.n6778 gnd.n669 9.3005
R10746 gnd.n6780 gnd.n6779 9.3005
R10747 gnd.n665 gnd.n664 9.3005
R10748 gnd.n6787 gnd.n6786 9.3005
R10749 gnd.n6788 gnd.n663 9.3005
R10750 gnd.n6790 gnd.n6789 9.3005
R10751 gnd.n659 gnd.n658 9.3005
R10752 gnd.n6797 gnd.n6796 9.3005
R10753 gnd.n6798 gnd.n657 9.3005
R10754 gnd.n6800 gnd.n6799 9.3005
R10755 gnd.n653 gnd.n652 9.3005
R10756 gnd.n6807 gnd.n6806 9.3005
R10757 gnd.n6808 gnd.n651 9.3005
R10758 gnd.n6810 gnd.n6809 9.3005
R10759 gnd.n647 gnd.n646 9.3005
R10760 gnd.n6817 gnd.n6816 9.3005
R10761 gnd.n6818 gnd.n645 9.3005
R10762 gnd.n6820 gnd.n6819 9.3005
R10763 gnd.n641 gnd.n640 9.3005
R10764 gnd.n6827 gnd.n6826 9.3005
R10765 gnd.n6828 gnd.n639 9.3005
R10766 gnd.n6830 gnd.n6829 9.3005
R10767 gnd.n635 gnd.n634 9.3005
R10768 gnd.n6837 gnd.n6836 9.3005
R10769 gnd.n6838 gnd.n633 9.3005
R10770 gnd.n6840 gnd.n6839 9.3005
R10771 gnd.n629 gnd.n628 9.3005
R10772 gnd.n6847 gnd.n6846 9.3005
R10773 gnd.n6848 gnd.n627 9.3005
R10774 gnd.n6850 gnd.n6849 9.3005
R10775 gnd.n623 gnd.n622 9.3005
R10776 gnd.n6857 gnd.n6856 9.3005
R10777 gnd.n6858 gnd.n621 9.3005
R10778 gnd.n6860 gnd.n6859 9.3005
R10779 gnd.n617 gnd.n616 9.3005
R10780 gnd.n6867 gnd.n6866 9.3005
R10781 gnd.n6868 gnd.n615 9.3005
R10782 gnd.n6870 gnd.n6869 9.3005
R10783 gnd.n611 gnd.n610 9.3005
R10784 gnd.n6877 gnd.n6876 9.3005
R10785 gnd.n6878 gnd.n609 9.3005
R10786 gnd.n6880 gnd.n6879 9.3005
R10787 gnd.n605 gnd.n604 9.3005
R10788 gnd.n6887 gnd.n6886 9.3005
R10789 gnd.n6888 gnd.n603 9.3005
R10790 gnd.n6890 gnd.n6889 9.3005
R10791 gnd.n599 gnd.n598 9.3005
R10792 gnd.n6897 gnd.n6896 9.3005
R10793 gnd.n6898 gnd.n597 9.3005
R10794 gnd.n6900 gnd.n6899 9.3005
R10795 gnd.n593 gnd.n592 9.3005
R10796 gnd.n6907 gnd.n6906 9.3005
R10797 gnd.n6908 gnd.n591 9.3005
R10798 gnd.n6910 gnd.n6909 9.3005
R10799 gnd.n587 gnd.n586 9.3005
R10800 gnd.n6917 gnd.n6916 9.3005
R10801 gnd.n6918 gnd.n585 9.3005
R10802 gnd.n6920 gnd.n6919 9.3005
R10803 gnd.n581 gnd.n580 9.3005
R10804 gnd.n6927 gnd.n6926 9.3005
R10805 gnd.n6928 gnd.n579 9.3005
R10806 gnd.n6930 gnd.n6929 9.3005
R10807 gnd.n575 gnd.n574 9.3005
R10808 gnd.n6937 gnd.n6936 9.3005
R10809 gnd.n6938 gnd.n573 9.3005
R10810 gnd.n6940 gnd.n6939 9.3005
R10811 gnd.n569 gnd.n568 9.3005
R10812 gnd.n6947 gnd.n6946 9.3005
R10813 gnd.n6948 gnd.n567 9.3005
R10814 gnd.n6950 gnd.n6949 9.3005
R10815 gnd.n563 gnd.n562 9.3005
R10816 gnd.n6957 gnd.n6956 9.3005
R10817 gnd.n6958 gnd.n561 9.3005
R10818 gnd.n6960 gnd.n6959 9.3005
R10819 gnd.n557 gnd.n556 9.3005
R10820 gnd.n6967 gnd.n6966 9.3005
R10821 gnd.n6968 gnd.n555 9.3005
R10822 gnd.n6970 gnd.n6969 9.3005
R10823 gnd.n551 gnd.n550 9.3005
R10824 gnd.n6977 gnd.n6976 9.3005
R10825 gnd.n6978 gnd.n549 9.3005
R10826 gnd.n6980 gnd.n6979 9.3005
R10827 gnd.n545 gnd.n544 9.3005
R10828 gnd.n6987 gnd.n6986 9.3005
R10829 gnd.n6988 gnd.n543 9.3005
R10830 gnd.n6991 gnd.n6990 9.3005
R10831 gnd.n6989 gnd.n539 9.3005
R10832 gnd.n6997 gnd.n538 9.3005
R10833 gnd.n6999 gnd.n6998 9.3005
R10834 gnd.n534 gnd.n533 9.3005
R10835 gnd.n7008 gnd.n7007 9.3005
R10836 gnd.n7009 gnd.n532 9.3005
R10837 gnd.n7011 gnd.n7010 9.3005
R10838 gnd.n528 gnd.n527 9.3005
R10839 gnd.n7018 gnd.n7017 9.3005
R10840 gnd.n7019 gnd.n526 9.3005
R10841 gnd.n7021 gnd.n7020 9.3005
R10842 gnd.n522 gnd.n521 9.3005
R10843 gnd.n7028 gnd.n7027 9.3005
R10844 gnd.n7029 gnd.n520 9.3005
R10845 gnd.n7031 gnd.n7030 9.3005
R10846 gnd.n516 gnd.n515 9.3005
R10847 gnd.n7038 gnd.n7037 9.3005
R10848 gnd.n7039 gnd.n514 9.3005
R10849 gnd.n7041 gnd.n7040 9.3005
R10850 gnd.n510 gnd.n509 9.3005
R10851 gnd.n7048 gnd.n7047 9.3005
R10852 gnd.n7049 gnd.n508 9.3005
R10853 gnd.n7051 gnd.n7050 9.3005
R10854 gnd.n504 gnd.n503 9.3005
R10855 gnd.n7058 gnd.n7057 9.3005
R10856 gnd.n7059 gnd.n502 9.3005
R10857 gnd.n7061 gnd.n7060 9.3005
R10858 gnd.n498 gnd.n497 9.3005
R10859 gnd.n7068 gnd.n7067 9.3005
R10860 gnd.n7069 gnd.n496 9.3005
R10861 gnd.n7071 gnd.n7070 9.3005
R10862 gnd.n492 gnd.n491 9.3005
R10863 gnd.n7078 gnd.n7077 9.3005
R10864 gnd.n7079 gnd.n490 9.3005
R10865 gnd.n7081 gnd.n7080 9.3005
R10866 gnd.n486 gnd.n485 9.3005
R10867 gnd.n7088 gnd.n7087 9.3005
R10868 gnd.n7089 gnd.n484 9.3005
R10869 gnd.n7091 gnd.n7090 9.3005
R10870 gnd.n480 gnd.n479 9.3005
R10871 gnd.n7098 gnd.n7097 9.3005
R10872 gnd.n7099 gnd.n478 9.3005
R10873 gnd.n7101 gnd.n7100 9.3005
R10874 gnd.n474 gnd.n473 9.3005
R10875 gnd.n7108 gnd.n7107 9.3005
R10876 gnd.n7109 gnd.n472 9.3005
R10877 gnd.n7111 gnd.n7110 9.3005
R10878 gnd.n468 gnd.n467 9.3005
R10879 gnd.n7118 gnd.n7117 9.3005
R10880 gnd.n7119 gnd.n466 9.3005
R10881 gnd.n7121 gnd.n7120 9.3005
R10882 gnd.n462 gnd.n461 9.3005
R10883 gnd.n7128 gnd.n7127 9.3005
R10884 gnd.n7129 gnd.n460 9.3005
R10885 gnd.n7131 gnd.n7130 9.3005
R10886 gnd.n456 gnd.n455 9.3005
R10887 gnd.n7138 gnd.n7137 9.3005
R10888 gnd.n7139 gnd.n454 9.3005
R10889 gnd.n7141 gnd.n7140 9.3005
R10890 gnd.n450 gnd.n449 9.3005
R10891 gnd.n7148 gnd.n7147 9.3005
R10892 gnd.n7149 gnd.n448 9.3005
R10893 gnd.n7151 gnd.n7150 9.3005
R10894 gnd.n444 gnd.n443 9.3005
R10895 gnd.n7158 gnd.n7157 9.3005
R10896 gnd.n7159 gnd.n442 9.3005
R10897 gnd.n7161 gnd.n7160 9.3005
R10898 gnd.n438 gnd.n437 9.3005
R10899 gnd.n7168 gnd.n7167 9.3005
R10900 gnd.n7169 gnd.n436 9.3005
R10901 gnd.n7171 gnd.n7170 9.3005
R10902 gnd.n432 gnd.n431 9.3005
R10903 gnd.n7178 gnd.n7177 9.3005
R10904 gnd.n7179 gnd.n430 9.3005
R10905 gnd.n7181 gnd.n7180 9.3005
R10906 gnd.n426 gnd.n425 9.3005
R10907 gnd.n7188 gnd.n7187 9.3005
R10908 gnd.n7189 gnd.n424 9.3005
R10909 gnd.n7191 gnd.n7190 9.3005
R10910 gnd.n420 gnd.n419 9.3005
R10911 gnd.n7198 gnd.n7197 9.3005
R10912 gnd.n7199 gnd.n418 9.3005
R10913 gnd.n7201 gnd.n7200 9.3005
R10914 gnd.n414 gnd.n413 9.3005
R10915 gnd.n7209 gnd.n7208 9.3005
R10916 gnd.n7210 gnd.n412 9.3005
R10917 gnd.n7212 gnd.n7211 9.3005
R10918 gnd.n7001 gnd.n7000 9.3005
R10919 gnd.n7417 gnd.n7416 9.3005
R10920 gnd.n7415 gnd.n69 9.3005
R10921 gnd.n5434 gnd.n71 9.3005
R10922 gnd.n5440 gnd.n5435 9.3005
R10923 gnd.n5439 gnd.n5436 9.3005
R10924 gnd.n5438 gnd.n5437 9.3005
R10925 gnd.n395 gnd.n394 9.3005
R10926 gnd.n7236 gnd.n7235 9.3005
R10927 gnd.n7237 gnd.n393 9.3005
R10928 gnd.n7239 gnd.n7238 9.3005
R10929 gnd.n390 gnd.n389 9.3005
R10930 gnd.n7251 gnd.n7250 9.3005
R10931 gnd.n7252 gnd.n388 9.3005
R10932 gnd.n7338 gnd.n7253 9.3005
R10933 gnd.n7337 gnd.n7254 9.3005
R10934 gnd.n7336 gnd.n7255 9.3005
R10935 gnd.n7334 gnd.n7256 9.3005
R10936 gnd.n7333 gnd.n7257 9.3005
R10937 gnd.n7331 gnd.n7258 9.3005
R10938 gnd.n7330 gnd.n7259 9.3005
R10939 gnd.n7328 gnd.n7327 9.3005
R10940 gnd.n7281 gnd.n7278 9.3005
R10941 gnd.n7287 gnd.n7286 9.3005
R10942 gnd.n7288 gnd.n7277 9.3005
R10943 gnd.n7290 gnd.n7289 9.3005
R10944 gnd.n7275 gnd.n7274 9.3005
R10945 gnd.n7297 gnd.n7296 9.3005
R10946 gnd.n7298 gnd.n7273 9.3005
R10947 gnd.n7300 gnd.n7299 9.3005
R10948 gnd.n7271 gnd.n7270 9.3005
R10949 gnd.n7307 gnd.n7306 9.3005
R10950 gnd.n7308 gnd.n7269 9.3005
R10951 gnd.n7310 gnd.n7309 9.3005
R10952 gnd.n7267 gnd.n7266 9.3005
R10953 gnd.n7317 gnd.n7316 9.3005
R10954 gnd.n7318 gnd.n7265 9.3005
R10955 gnd.n7320 gnd.n7319 9.3005
R10956 gnd.n7263 gnd.n7260 9.3005
R10957 gnd.n7326 gnd.n7325 9.3005
R10958 gnd.n7280 gnd.n7279 9.3005
R10959 gnd.n239 gnd.n236 9.3005
R10960 gnd.n245 gnd.n244 9.3005
R10961 gnd.n246 gnd.n235 9.3005
R10962 gnd.n248 gnd.n247 9.3005
R10963 gnd.n233 gnd.n232 9.3005
R10964 gnd.n255 gnd.n254 9.3005
R10965 gnd.n256 gnd.n231 9.3005
R10966 gnd.n258 gnd.n257 9.3005
R10967 gnd.n229 gnd.n228 9.3005
R10968 gnd.n265 gnd.n264 9.3005
R10969 gnd.n266 gnd.n227 9.3005
R10970 gnd.n268 gnd.n267 9.3005
R10971 gnd.n225 gnd.n224 9.3005
R10972 gnd.n276 gnd.n275 9.3005
R10973 gnd.n277 gnd.n223 9.3005
R10974 gnd.n279 gnd.n278 9.3005
R10975 gnd.n280 gnd.n218 9.3005
R10976 gnd.n286 gnd.n285 9.3005
R10977 gnd.n287 gnd.n217 9.3005
R10978 gnd.n289 gnd.n288 9.3005
R10979 gnd.n215 gnd.n214 9.3005
R10980 gnd.n296 gnd.n295 9.3005
R10981 gnd.n297 gnd.n213 9.3005
R10982 gnd.n299 gnd.n298 9.3005
R10983 gnd.n211 gnd.n210 9.3005
R10984 gnd.n306 gnd.n305 9.3005
R10985 gnd.n307 gnd.n209 9.3005
R10986 gnd.n309 gnd.n308 9.3005
R10987 gnd.n207 gnd.n206 9.3005
R10988 gnd.n316 gnd.n315 9.3005
R10989 gnd.n317 gnd.n205 9.3005
R10990 gnd.n319 gnd.n318 9.3005
R10991 gnd.n203 gnd.n202 9.3005
R10992 gnd.n326 gnd.n325 9.3005
R10993 gnd.n327 gnd.n201 9.3005
R10994 gnd.n329 gnd.n328 9.3005
R10995 gnd.n199 gnd.n196 9.3005
R10996 gnd.n336 gnd.n335 9.3005
R10997 gnd.n337 gnd.n195 9.3005
R10998 gnd.n339 gnd.n338 9.3005
R10999 gnd.n193 gnd.n192 9.3005
R11000 gnd.n346 gnd.n345 9.3005
R11001 gnd.n347 gnd.n191 9.3005
R11002 gnd.n349 gnd.n348 9.3005
R11003 gnd.n189 gnd.n188 9.3005
R11004 gnd.n356 gnd.n355 9.3005
R11005 gnd.n357 gnd.n187 9.3005
R11006 gnd.n359 gnd.n358 9.3005
R11007 gnd.n185 gnd.n184 9.3005
R11008 gnd.n366 gnd.n365 9.3005
R11009 gnd.n367 gnd.n183 9.3005
R11010 gnd.n369 gnd.n368 9.3005
R11011 gnd.n181 gnd.n180 9.3005
R11012 gnd.n376 gnd.n375 9.3005
R11013 gnd.n377 gnd.n179 9.3005
R11014 gnd.n379 gnd.n378 9.3005
R11015 gnd.n177 gnd.n174 9.3005
R11016 gnd.n385 gnd.n384 9.3005
R11017 gnd.n238 gnd.n237 9.3005
R11018 gnd.n5525 gnd.n5524 9.3005
R11019 gnd.n3274 gnd.n3273 9.3005
R11020 gnd.n3298 gnd.n3297 9.3005
R11021 gnd.n5512 gnd.n3299 9.3005
R11022 gnd.n5511 gnd.n3300 9.3005
R11023 gnd.n5510 gnd.n3301 9.3005
R11024 gnd.n5317 gnd.n3302 9.3005
R11025 gnd.n5500 gnd.n3319 9.3005
R11026 gnd.n5499 gnd.n3320 9.3005
R11027 gnd.n5498 gnd.n3321 9.3005
R11028 gnd.n5323 gnd.n3322 9.3005
R11029 gnd.n5488 gnd.n3339 9.3005
R11030 gnd.n5487 gnd.n3340 9.3005
R11031 gnd.n5486 gnd.n3341 9.3005
R11032 gnd.n5400 gnd.n3342 9.3005
R11033 gnd.n5476 gnd.n3356 9.3005
R11034 gnd.n5475 gnd.n3357 9.3005
R11035 gnd.n5474 gnd.n3358 9.3005
R11036 gnd.n5420 gnd.n3359 9.3005
R11037 gnd.n5422 gnd.n5421 9.3005
R11038 gnd.n3387 gnd.n3381 9.3005
R11039 gnd.n5456 gnd.n3382 9.3005
R11040 gnd.n5455 gnd.n3383 9.3005
R11041 gnd.n5454 gnd.n3384 9.3005
R11042 gnd.n5431 gnd.n96 9.3005
R11043 gnd.n7403 gnd.n97 9.3005
R11044 gnd.n7402 gnd.n98 9.3005
R11045 gnd.n7401 gnd.n99 9.3005
R11046 gnd.n7230 gnd.n100 9.3005
R11047 gnd.n7391 gnd.n115 9.3005
R11048 gnd.n7390 gnd.n116 9.3005
R11049 gnd.n7389 gnd.n117 9.3005
R11050 gnd.n7245 gnd.n118 9.3005
R11051 gnd.n7379 gnd.n136 9.3005
R11052 gnd.n7378 gnd.n137 9.3005
R11053 gnd.n7377 gnd.n138 9.3005
R11054 gnd.n7344 gnd.n139 9.3005
R11055 gnd.n7367 gnd.n155 9.3005
R11056 gnd.n7366 gnd.n156 9.3005
R11057 gnd.n7365 gnd.n157 9.3005
R11058 gnd.n173 gnd.n158 9.3005
R11059 gnd.n7355 gnd.n7354 9.3005
R11060 gnd.n5526 gnd.n3272 9.3005
R11061 gnd.n5524 gnd.n5523 9.3005
R11062 gnd.n5522 gnd.n3274 9.3005
R11063 gnd.n3298 gnd.n3275 9.3005
R11064 gnd.n5312 gnd.n3299 9.3005
R11065 gnd.n5315 gnd.n3300 9.3005
R11066 gnd.n5316 gnd.n3301 9.3005
R11067 gnd.n5321 gnd.n5317 9.3005
R11068 gnd.n5322 gnd.n3319 9.3005
R11069 gnd.n5326 gnd.n3320 9.3005
R11070 gnd.n5325 gnd.n3321 9.3005
R11071 gnd.n5324 gnd.n5323 9.3005
R11072 gnd.n3397 gnd.n3339 9.3005
R11073 gnd.n5398 gnd.n3340 9.3005
R11074 gnd.n5399 gnd.n3341 9.3005
R11075 gnd.n5401 gnd.n5400 9.3005
R11076 gnd.n3391 gnd.n3356 9.3005
R11077 gnd.n5417 gnd.n3357 9.3005
R11078 gnd.n5418 gnd.n3358 9.3005
R11079 gnd.n5420 gnd.n5419 9.3005
R11080 gnd.n5421 gnd.n3386 9.3005
R11081 gnd.n5427 gnd.n3387 9.3005
R11082 gnd.n5428 gnd.n3382 9.3005
R11083 gnd.n5429 gnd.n3383 9.3005
R11084 gnd.n5430 gnd.n3384 9.3005
R11085 gnd.n5432 gnd.n5431 9.3005
R11086 gnd.n396 gnd.n97 9.3005
R11087 gnd.n7228 gnd.n98 9.3005
R11088 gnd.n7229 gnd.n99 9.3005
R11089 gnd.n7231 gnd.n7230 9.3005
R11090 gnd.n391 gnd.n115 9.3005
R11091 gnd.n7243 gnd.n116 9.3005
R11092 gnd.n7244 gnd.n117 9.3005
R11093 gnd.n7246 gnd.n7245 9.3005
R11094 gnd.n387 gnd.n136 9.3005
R11095 gnd.n7342 gnd.n137 9.3005
R11096 gnd.n7343 gnd.n138 9.3005
R11097 gnd.n7346 gnd.n7344 9.3005
R11098 gnd.n7347 gnd.n155 9.3005
R11099 gnd.n7349 gnd.n156 9.3005
R11100 gnd.n7350 gnd.n157 9.3005
R11101 gnd.n7352 gnd.n173 9.3005
R11102 gnd.n7354 gnd.n7353 9.3005
R11103 gnd.n3272 gnd.n3266 9.3005
R11104 gnd.n5536 gnd.n5535 9.3005
R11105 gnd.n5539 gnd.n3264 9.3005
R11106 gnd.n5540 gnd.n3263 9.3005
R11107 gnd.n5543 gnd.n3262 9.3005
R11108 gnd.n5544 gnd.n3261 9.3005
R11109 gnd.n5547 gnd.n3260 9.3005
R11110 gnd.n5548 gnd.n3259 9.3005
R11111 gnd.n5551 gnd.n3258 9.3005
R11112 gnd.n5552 gnd.n3257 9.3005
R11113 gnd.n5555 gnd.n3256 9.3005
R11114 gnd.n5556 gnd.n3255 9.3005
R11115 gnd.n5559 gnd.n3254 9.3005
R11116 gnd.n5560 gnd.n3253 9.3005
R11117 gnd.n5563 gnd.n3252 9.3005
R11118 gnd.n5564 gnd.n3251 9.3005
R11119 gnd.n5567 gnd.n3250 9.3005
R11120 gnd.n5568 gnd.n3249 9.3005
R11121 gnd.n5571 gnd.n3248 9.3005
R11122 gnd.n5572 gnd.n3247 9.3005
R11123 gnd.n5575 gnd.n3246 9.3005
R11124 gnd.n5579 gnd.n3242 9.3005
R11125 gnd.n5580 gnd.n3241 9.3005
R11126 gnd.n5583 gnd.n3240 9.3005
R11127 gnd.n5584 gnd.n3239 9.3005
R11128 gnd.n5587 gnd.n3238 9.3005
R11129 gnd.n5588 gnd.n3237 9.3005
R11130 gnd.n5591 gnd.n3236 9.3005
R11131 gnd.n5592 gnd.n3235 9.3005
R11132 gnd.n5595 gnd.n3234 9.3005
R11133 gnd.n5597 gnd.n3230 9.3005
R11134 gnd.n5600 gnd.n3229 9.3005
R11135 gnd.n5601 gnd.n3228 9.3005
R11136 gnd.n5604 gnd.n3227 9.3005
R11137 gnd.n5605 gnd.n3226 9.3005
R11138 gnd.n5608 gnd.n3225 9.3005
R11139 gnd.n5609 gnd.n3224 9.3005
R11140 gnd.n5612 gnd.n3223 9.3005
R11141 gnd.n5614 gnd.n3220 9.3005
R11142 gnd.n5617 gnd.n3219 9.3005
R11143 gnd.n5618 gnd.n3218 9.3005
R11144 gnd.n5621 gnd.n3217 9.3005
R11145 gnd.n5622 gnd.n3216 9.3005
R11146 gnd.n5625 gnd.n3215 9.3005
R11147 gnd.n5626 gnd.n3214 9.3005
R11148 gnd.n5629 gnd.n3213 9.3005
R11149 gnd.n5630 gnd.n3212 9.3005
R11150 gnd.n5633 gnd.n3211 9.3005
R11151 gnd.n5634 gnd.n3210 9.3005
R11152 gnd.n5637 gnd.n3209 9.3005
R11153 gnd.n5638 gnd.n3208 9.3005
R11154 gnd.n5641 gnd.n3207 9.3005
R11155 gnd.n5643 gnd.n3206 9.3005
R11156 gnd.n5644 gnd.n3205 9.3005
R11157 gnd.n5645 gnd.n3204 9.3005
R11158 gnd.n5646 gnd.n3203 9.3005
R11159 gnd.n5576 gnd.n3243 9.3005
R11160 gnd.n5534 gnd.n5531 9.3005
R11161 gnd.n3285 gnd.n3282 9.3005
R11162 gnd.n5518 gnd.n3286 9.3005
R11163 gnd.n5517 gnd.n3287 9.3005
R11164 gnd.n5516 gnd.n3288 9.3005
R11165 gnd.n3308 gnd.n3289 9.3005
R11166 gnd.n5506 gnd.n3309 9.3005
R11167 gnd.n5505 gnd.n3310 9.3005
R11168 gnd.n5504 gnd.n3311 9.3005
R11169 gnd.n3329 gnd.n3312 9.3005
R11170 gnd.n5494 gnd.n3330 9.3005
R11171 gnd.n5493 gnd.n3331 9.3005
R11172 gnd.n5492 gnd.n3332 9.3005
R11173 gnd.n3348 gnd.n3333 9.3005
R11174 gnd.n5482 gnd.n3349 9.3005
R11175 gnd.n5481 gnd.n82 9.3005
R11176 gnd.n87 gnd.n81 9.3005
R11177 gnd.n7397 gnd.n106 9.3005
R11178 gnd.n7396 gnd.n107 9.3005
R11179 gnd.n7395 gnd.n108 9.3005
R11180 gnd.n125 gnd.n109 9.3005
R11181 gnd.n7385 gnd.n126 9.3005
R11182 gnd.n7384 gnd.n127 9.3005
R11183 gnd.n7383 gnd.n128 9.3005
R11184 gnd.n145 gnd.n129 9.3005
R11185 gnd.n7373 gnd.n146 9.3005
R11186 gnd.n7372 gnd.n147 9.3005
R11187 gnd.n7371 gnd.n148 9.3005
R11188 gnd.n163 gnd.n149 9.3005
R11189 gnd.n7361 gnd.n164 9.3005
R11190 gnd.n7360 gnd.n165 9.3005
R11191 gnd.n7359 gnd.n166 9.3005
R11192 gnd.n3284 gnd.n3283 9.3005
R11193 gnd.n7408 gnd.n7407 9.3005
R11194 gnd.n4295 gnd.n4294 9.3005
R11195 gnd.n4314 gnd.n4296 9.3005
R11196 gnd.n4313 gnd.n4297 9.3005
R11197 gnd.n4312 gnd.n4298 9.3005
R11198 gnd.n4301 gnd.n4299 9.3005
R11199 gnd.n4308 gnd.n4302 9.3005
R11200 gnd.n4307 gnd.n4303 9.3005
R11201 gnd.n4306 gnd.n4304 9.3005
R11202 gnd.n3997 gnd.n3996 9.3005
R11203 gnd.n4367 gnd.n4366 9.3005
R11204 gnd.n4368 gnd.n3995 9.3005
R11205 gnd.n4370 gnd.n4369 9.3005
R11206 gnd.n3993 gnd.n3992 9.3005
R11207 gnd.n4375 gnd.n4374 9.3005
R11208 gnd.n4376 gnd.n3991 9.3005
R11209 gnd.n4378 gnd.n4377 9.3005
R11210 gnd.n3989 gnd.n3988 9.3005
R11211 gnd.n4383 gnd.n4382 9.3005
R11212 gnd.n4384 gnd.n3987 9.3005
R11213 gnd.n4386 gnd.n4385 9.3005
R11214 gnd.n3985 gnd.n3984 9.3005
R11215 gnd.n4392 gnd.n4391 9.3005
R11216 gnd.n4393 gnd.n3983 9.3005
R11217 gnd.n4395 gnd.n4394 9.3005
R11218 gnd.n3921 gnd.n3920 9.3005
R11219 gnd.n4408 gnd.n4407 9.3005
R11220 gnd.n4409 gnd.n3919 9.3005
R11221 gnd.n4411 gnd.n4410 9.3005
R11222 gnd.n3907 gnd.n3906 9.3005
R11223 gnd.n4424 gnd.n4423 9.3005
R11224 gnd.n4425 gnd.n3905 9.3005
R11225 gnd.n4427 gnd.n4426 9.3005
R11226 gnd.n3893 gnd.n3892 9.3005
R11227 gnd.n4440 gnd.n4439 9.3005
R11228 gnd.n4441 gnd.n3891 9.3005
R11229 gnd.n4443 gnd.n4442 9.3005
R11230 gnd.n3879 gnd.n3878 9.3005
R11231 gnd.n4456 gnd.n4455 9.3005
R11232 gnd.n4457 gnd.n3877 9.3005
R11233 gnd.n4459 gnd.n4458 9.3005
R11234 gnd.n3862 gnd.n3861 9.3005
R11235 gnd.n4483 gnd.n4482 9.3005
R11236 gnd.n4484 gnd.n3860 9.3005
R11237 gnd.n4489 gnd.n4485 9.3005
R11238 gnd.n4488 gnd.n4487 9.3005
R11239 gnd.n4486 gnd.n2981 9.3005
R11240 gnd.n5838 gnd.n2982 9.3005
R11241 gnd.n5837 gnd.n2983 9.3005
R11242 gnd.n5836 gnd.n2984 9.3005
R11243 gnd.n4517 gnd.n2985 9.3005
R11244 gnd.n4521 gnd.n4518 9.3005
R11245 gnd.n4520 gnd.n4519 9.3005
R11246 gnd.n3745 gnd.n3744 9.3005
R11247 gnd.n4574 gnd.n4573 9.3005
R11248 gnd.n4575 gnd.n3743 9.3005
R11249 gnd.n4579 gnd.n4576 9.3005
R11250 gnd.n4578 gnd.n4577 9.3005
R11251 gnd.n3723 gnd.n3722 9.3005
R11252 gnd.n4614 gnd.n4613 9.3005
R11253 gnd.n4615 gnd.n3721 9.3005
R11254 gnd.n4617 gnd.n4616 9.3005
R11255 gnd.n3697 gnd.n3696 9.3005
R11256 gnd.n4658 gnd.n4657 9.3005
R11257 gnd.n4659 gnd.n3695 9.3005
R11258 gnd.n4663 gnd.n4660 9.3005
R11259 gnd.n4662 gnd.n4661 9.3005
R11260 gnd.n3677 gnd.n3676 9.3005
R11261 gnd.n4710 gnd.n4709 9.3005
R11262 gnd.n4711 gnd.n3675 9.3005
R11263 gnd.n4724 gnd.n4712 9.3005
R11264 gnd.n4723 gnd.n4713 9.3005
R11265 gnd.n4722 gnd.n4714 9.3005
R11266 gnd.n4716 gnd.n4715 9.3005
R11267 gnd.n4718 gnd.n4717 9.3005
R11268 gnd.n3639 gnd.n3638 9.3005
R11269 gnd.n4772 gnd.n4771 9.3005
R11270 gnd.n4773 gnd.n3637 9.3005
R11271 gnd.n4775 gnd.n4774 9.3005
R11272 gnd.n3617 gnd.n3616 9.3005
R11273 gnd.n4832 gnd.n4831 9.3005
R11274 gnd.n4833 gnd.n3615 9.3005
R11275 gnd.n4835 gnd.n4834 9.3005
R11276 gnd.n3599 gnd.n3598 9.3005
R11277 gnd.n4860 gnd.n4859 9.3005
R11278 gnd.n4861 gnd.n3597 9.3005
R11279 gnd.n4863 gnd.n4862 9.3005
R11280 gnd.n3581 gnd.n3580 9.3005
R11281 gnd.n4885 gnd.n4884 9.3005
R11282 gnd.n4886 gnd.n3579 9.3005
R11283 gnd.n4890 gnd.n4887 9.3005
R11284 gnd.n4889 gnd.n4888 9.3005
R11285 gnd.n3552 gnd.n3551 9.3005
R11286 gnd.n4941 gnd.n4940 9.3005
R11287 gnd.n4942 gnd.n3550 9.3005
R11288 gnd.n4946 gnd.n4943 9.3005
R11289 gnd.n4945 gnd.n4944 9.3005
R11290 gnd.n3521 gnd.n3520 9.3005
R11291 gnd.n5172 gnd.n5171 9.3005
R11292 gnd.n5173 gnd.n3519 9.3005
R11293 gnd.n5175 gnd.n5174 9.3005
R11294 gnd.n3509 gnd.n3508 9.3005
R11295 gnd.n5190 gnd.n5189 9.3005
R11296 gnd.n5191 gnd.n3507 9.3005
R11297 gnd.n5193 gnd.n5192 9.3005
R11298 gnd.n3498 gnd.n3497 9.3005
R11299 gnd.n5207 gnd.n5206 9.3005
R11300 gnd.n5208 gnd.n3496 9.3005
R11301 gnd.n5210 gnd.n5209 9.3005
R11302 gnd.n3486 gnd.n3485 9.3005
R11303 gnd.n5224 gnd.n5223 9.3005
R11304 gnd.n5225 gnd.n3484 9.3005
R11305 gnd.n5227 gnd.n5226 9.3005
R11306 gnd.n3474 gnd.n3473 9.3005
R11307 gnd.n5241 gnd.n5240 9.3005
R11308 gnd.n5242 gnd.n3472 9.3005
R11309 gnd.n5244 gnd.n5243 9.3005
R11310 gnd.n3462 gnd.n3461 9.3005
R11311 gnd.n5258 gnd.n5257 9.3005
R11312 gnd.n5259 gnd.n3460 9.3005
R11313 gnd.n5264 gnd.n5260 9.3005
R11314 gnd.n5263 gnd.n5262 9.3005
R11315 gnd.n5261 gnd.n3450 9.3005
R11316 gnd.n5278 gnd.n3449 9.3005
R11317 gnd.n5280 gnd.n5279 9.3005
R11318 gnd.n5281 gnd.n3448 9.3005
R11319 gnd.n5294 gnd.n5282 9.3005
R11320 gnd.n5293 gnd.n5283 9.3005
R11321 gnd.n5292 gnd.n5284 9.3005
R11322 gnd.n5286 gnd.n5285 9.3005
R11323 gnd.n5288 gnd.n5287 9.3005
R11324 gnd.n3414 gnd.n3413 9.3005
R11325 gnd.n5349 gnd.n5348 9.3005
R11326 gnd.n5350 gnd.n3412 9.3005
R11327 gnd.n5352 gnd.n5351 9.3005
R11328 gnd.n3410 gnd.n3409 9.3005
R11329 gnd.n5357 gnd.n5356 9.3005
R11330 gnd.n5358 gnd.n3408 9.3005
R11331 gnd.n5360 gnd.n5359 9.3005
R11332 gnd.n3406 gnd.n3405 9.3005
R11333 gnd.n5365 gnd.n5364 9.3005
R11334 gnd.n5366 gnd.n3404 9.3005
R11335 gnd.n5385 gnd.n5367 9.3005
R11336 gnd.n5384 gnd.n5368 9.3005
R11337 gnd.n5383 gnd.n5369 9.3005
R11338 gnd.n5372 gnd.n5370 9.3005
R11339 gnd.n5379 gnd.n5373 9.3005
R11340 gnd.n401 gnd.n400 9.3005
R11341 gnd.n7223 gnd.n402 9.3005
R11342 gnd.n7222 gnd.n403 9.3005
R11343 gnd.n7221 gnd.n404 9.3005
R11344 gnd.n407 gnd.n405 9.3005
R11345 gnd.n7217 gnd.n408 9.3005
R11346 gnd.n7216 gnd.n409 9.3005
R11347 gnd.n7215 gnd.n410 9.3005
R11348 gnd.n4257 gnd.n4256 9.3005
R11349 gnd.n4155 gnd.n4093 9.3005
R11350 gnd.n4158 gnd.n4157 9.3005
R11351 gnd.n4159 gnd.n4092 9.3005
R11352 gnd.n4162 gnd.n4160 9.3005
R11353 gnd.n4163 gnd.n4091 9.3005
R11354 gnd.n4166 gnd.n4165 9.3005
R11355 gnd.n4167 gnd.n4090 9.3005
R11356 gnd.n4170 gnd.n4169 9.3005
R11357 gnd.n4168 gnd.n4075 9.3005
R11358 gnd.n4205 gnd.n4076 9.3005
R11359 gnd.n4204 gnd.n4077 9.3005
R11360 gnd.n4203 gnd.n4078 9.3005
R11361 gnd.n4181 gnd.n4079 9.3005
R11362 gnd.n4193 gnd.n4182 9.3005
R11363 gnd.n4192 gnd.n4183 9.3005
R11364 gnd.n4191 gnd.n4184 9.3005
R11365 gnd.n4186 gnd.n4185 9.3005
R11366 gnd.n4050 gnd.n4049 9.3005
R11367 gnd.n4254 gnd.n4253 9.3005
R11368 gnd.n4255 gnd.n4048 9.3005
R11369 gnd.n4154 gnd.n4152 9.3005
R11370 gnd.n4148 gnd.n4147 9.3005
R11371 gnd.n4146 gnd.n4098 9.3005
R11372 gnd.n4145 gnd.n4144 9.3005
R11373 gnd.n4141 gnd.n4101 9.3005
R11374 gnd.n4140 gnd.n4137 9.3005
R11375 gnd.n4136 gnd.n4102 9.3005
R11376 gnd.n4135 gnd.n4134 9.3005
R11377 gnd.n4131 gnd.n4103 9.3005
R11378 gnd.n4130 gnd.n4127 9.3005
R11379 gnd.n4126 gnd.n4104 9.3005
R11380 gnd.n4125 gnd.n4124 9.3005
R11381 gnd.n4121 gnd.n4105 9.3005
R11382 gnd.n4120 gnd.n4117 9.3005
R11383 gnd.n4116 gnd.n4106 9.3005
R11384 gnd.n4115 gnd.n4114 9.3005
R11385 gnd.n4111 gnd.n4107 9.3005
R11386 gnd.n4110 gnd.n2448 9.3005
R11387 gnd.n4149 gnd.n4094 9.3005
R11388 gnd.n4151 gnd.n4150 9.3005
R11389 gnd.n5916 gnd.n2812 9.3005
R11390 gnd.n5919 gnd.n2811 9.3005
R11391 gnd.n5920 gnd.n2810 9.3005
R11392 gnd.n5923 gnd.n2809 9.3005
R11393 gnd.n5924 gnd.n2808 9.3005
R11394 gnd.n5927 gnd.n2807 9.3005
R11395 gnd.n5928 gnd.n2806 9.3005
R11396 gnd.n5931 gnd.n2805 9.3005
R11397 gnd.n5933 gnd.n2802 9.3005
R11398 gnd.n5936 gnd.n2801 9.3005
R11399 gnd.n5937 gnd.n2800 9.3005
R11400 gnd.n5940 gnd.n2799 9.3005
R11401 gnd.n5941 gnd.n2798 9.3005
R11402 gnd.n5944 gnd.n2797 9.3005
R11403 gnd.n5945 gnd.n2796 9.3005
R11404 gnd.n5948 gnd.n2795 9.3005
R11405 gnd.n5949 gnd.n2794 9.3005
R11406 gnd.n5952 gnd.n2793 9.3005
R11407 gnd.n5953 gnd.n2792 9.3005
R11408 gnd.n5956 gnd.n2791 9.3005
R11409 gnd.n5957 gnd.n2790 9.3005
R11410 gnd.n5960 gnd.n2789 9.3005
R11411 gnd.n5961 gnd.n2788 9.3005
R11412 gnd.n5962 gnd.n2787 9.3005
R11413 gnd.n2786 gnd.n2783 9.3005
R11414 gnd.n2785 gnd.n2784 9.3005
R11415 gnd.n2909 gnd.n2908 9.3005
R11416 gnd.n2905 gnd.n2815 9.3005
R11417 gnd.n2902 gnd.n2816 9.3005
R11418 gnd.n2901 gnd.n2817 9.3005
R11419 gnd.n2898 gnd.n2818 9.3005
R11420 gnd.n2897 gnd.n2819 9.3005
R11421 gnd.n2894 gnd.n2820 9.3005
R11422 gnd.n2893 gnd.n2821 9.3005
R11423 gnd.n2890 gnd.n2889 9.3005
R11424 gnd.n2888 gnd.n2822 9.3005
R11425 gnd.n2887 gnd.n2886 9.3005
R11426 gnd.n2883 gnd.n2825 9.3005
R11427 gnd.n2880 gnd.n2826 9.3005
R11428 gnd.n2879 gnd.n2827 9.3005
R11429 gnd.n2876 gnd.n2828 9.3005
R11430 gnd.n2875 gnd.n2829 9.3005
R11431 gnd.n2872 gnd.n2830 9.3005
R11432 gnd.n2871 gnd.n2831 9.3005
R11433 gnd.n2868 gnd.n2832 9.3005
R11434 gnd.n2867 gnd.n2833 9.3005
R11435 gnd.n2864 gnd.n2834 9.3005
R11436 gnd.n2863 gnd.n2835 9.3005
R11437 gnd.n2860 gnd.n2836 9.3005
R11438 gnd.n2859 gnd.n2837 9.3005
R11439 gnd.n2856 gnd.n2838 9.3005
R11440 gnd.n2855 gnd.n2839 9.3005
R11441 gnd.n2852 gnd.n2840 9.3005
R11442 gnd.n2851 gnd.n2841 9.3005
R11443 gnd.n2848 gnd.n2847 9.3005
R11444 gnd.n2846 gnd.n2843 9.3005
R11445 gnd.n2910 gnd.n2813 9.3005
R11446 gnd.n2470 gnd.n2450 9.3005
R11447 gnd.n4080 gnd.n2471 9.3005
R11448 gnd.n6144 gnd.n2472 9.3005
R11449 gnd.n6143 gnd.n2473 9.3005
R11450 gnd.n6142 gnd.n2474 9.3005
R11451 gnd.n4086 gnd.n2475 9.3005
R11452 gnd.n6132 gnd.n2491 9.3005
R11453 gnd.n6131 gnd.n2492 9.3005
R11454 gnd.n6130 gnd.n2493 9.3005
R11455 gnd.n4176 gnd.n2494 9.3005
R11456 gnd.n6120 gnd.n2511 9.3005
R11457 gnd.n6119 gnd.n2512 9.3005
R11458 gnd.n6118 gnd.n2513 9.3005
R11459 gnd.n4179 gnd.n2514 9.3005
R11460 gnd.n6108 gnd.n2532 9.3005
R11461 gnd.n6107 gnd.n2533 9.3005
R11462 gnd.n6106 gnd.n2534 9.3005
R11463 gnd.n4058 gnd.n2535 9.3005
R11464 gnd.n4244 gnd.n4057 9.3005
R11465 gnd.n4246 gnd.n4245 9.3005
R11466 gnd.n4044 gnd.n4039 9.3005
R11467 gnd.n4273 gnd.n4040 9.3005
R11468 gnd.n4272 gnd.n4041 9.3005
R11469 gnd.n4271 gnd.n4269 9.3005
R11470 gnd.n4042 gnd.n2558 9.3005
R11471 gnd.n6094 gnd.n2559 9.3005
R11472 gnd.n6093 gnd.n2560 9.3005
R11473 gnd.n6092 gnd.n2561 9.3005
R11474 gnd.n4012 gnd.n2562 9.3005
R11475 gnd.n6082 gnd.n2577 9.3005
R11476 gnd.n6081 gnd.n2578 9.3005
R11477 gnd.n6080 gnd.n2579 9.3005
R11478 gnd.n4006 gnd.n2580 9.3005
R11479 gnd.n6070 gnd.n2598 9.3005
R11480 gnd.n6069 gnd.n2599 9.3005
R11481 gnd.n6068 gnd.n2600 9.3005
R11482 gnd.n4345 gnd.n2601 9.3005
R11483 gnd.n6058 gnd.n2618 9.3005
R11484 gnd.n6057 gnd.n2619 9.3005
R11485 gnd.n6056 gnd.n2620 9.3005
R11486 gnd.n2637 gnd.n2621 9.3005
R11487 gnd.n6046 gnd.n6045 9.3005
R11488 gnd.n6156 gnd.n2449 9.3005
R11489 gnd.n2451 gnd.n2450 9.3005
R11490 gnd.n4081 gnd.n4080 9.3005
R11491 gnd.n4082 gnd.n2472 9.3005
R11492 gnd.n4084 gnd.n2473 9.3005
R11493 gnd.n4085 gnd.n2474 9.3005
R11494 gnd.n4088 gnd.n4086 9.3005
R11495 gnd.n4089 gnd.n2491 9.3005
R11496 gnd.n4174 gnd.n2492 9.3005
R11497 gnd.n4175 gnd.n2493 9.3005
R11498 gnd.n4177 gnd.n4176 9.3005
R11499 gnd.n4178 gnd.n2511 9.3005
R11500 gnd.n4199 gnd.n2512 9.3005
R11501 gnd.n4198 gnd.n2513 9.3005
R11502 gnd.n4197 gnd.n4179 9.3005
R11503 gnd.n4180 gnd.n2532 9.3005
R11504 gnd.n4187 gnd.n2533 9.3005
R11505 gnd.n4059 gnd.n2534 9.3005
R11506 gnd.n4242 gnd.n4058 9.3005
R11507 gnd.n4244 gnd.n4243 9.3005
R11508 gnd.n4245 gnd.n4043 9.3005
R11509 gnd.n4261 gnd.n4044 9.3005
R11510 gnd.n4262 gnd.n4040 9.3005
R11511 gnd.n4263 gnd.n4041 9.3005
R11512 gnd.n4269 gnd.n4268 9.3005
R11513 gnd.n4266 gnd.n4042 9.3005
R11514 gnd.n4265 gnd.n2559 9.3005
R11515 gnd.n4264 gnd.n2560 9.3005
R11516 gnd.n4011 gnd.n2561 9.3005
R11517 gnd.n4327 gnd.n4012 9.3005
R11518 gnd.n4328 gnd.n2577 9.3005
R11519 gnd.n4329 gnd.n2578 9.3005
R11520 gnd.n4005 gnd.n2579 9.3005
R11521 gnd.n4341 gnd.n4006 9.3005
R11522 gnd.n4342 gnd.n2598 9.3005
R11523 gnd.n4343 gnd.n2599 9.3005
R11524 gnd.n4344 gnd.n2600 9.3005
R11525 gnd.n4348 gnd.n4345 9.3005
R11526 gnd.n4349 gnd.n2618 9.3005
R11527 gnd.n4350 gnd.n2619 9.3005
R11528 gnd.n2639 gnd.n2620 9.3005
R11529 gnd.n6043 gnd.n2637 9.3005
R11530 gnd.n6045 gnd.n6044 9.3005
R11531 gnd.n6156 gnd.n6155 9.3005
R11532 gnd.n6160 gnd.n6159 9.3005
R11533 gnd.n6163 gnd.n2444 9.3005
R11534 gnd.n6164 gnd.n2443 9.3005
R11535 gnd.n6167 gnd.n2442 9.3005
R11536 gnd.n6168 gnd.n2441 9.3005
R11537 gnd.n6171 gnd.n2440 9.3005
R11538 gnd.n6172 gnd.n2439 9.3005
R11539 gnd.n6175 gnd.n2438 9.3005
R11540 gnd.n6176 gnd.n2437 9.3005
R11541 gnd.n6179 gnd.n2436 9.3005
R11542 gnd.n6180 gnd.n2435 9.3005
R11543 gnd.n6183 gnd.n2434 9.3005
R11544 gnd.n6184 gnd.n2433 9.3005
R11545 gnd.n6187 gnd.n2432 9.3005
R11546 gnd.n6188 gnd.n2431 9.3005
R11547 gnd.n6191 gnd.n2430 9.3005
R11548 gnd.n6192 gnd.n2429 9.3005
R11549 gnd.n6195 gnd.n2428 9.3005
R11550 gnd.n6196 gnd.n2427 9.3005
R11551 gnd.n6199 gnd.n2426 9.3005
R11552 gnd.n6203 gnd.n2422 9.3005
R11553 gnd.n6204 gnd.n2421 9.3005
R11554 gnd.n6207 gnd.n2420 9.3005
R11555 gnd.n6208 gnd.n2419 9.3005
R11556 gnd.n6211 gnd.n2418 9.3005
R11557 gnd.n6212 gnd.n2417 9.3005
R11558 gnd.n6215 gnd.n2416 9.3005
R11559 gnd.n6216 gnd.n2415 9.3005
R11560 gnd.n6219 gnd.n2414 9.3005
R11561 gnd.n6220 gnd.n2413 9.3005
R11562 gnd.n6223 gnd.n2412 9.3005
R11563 gnd.n6224 gnd.n2411 9.3005
R11564 gnd.n6227 gnd.n2410 9.3005
R11565 gnd.n6228 gnd.n2409 9.3005
R11566 gnd.n6231 gnd.n2408 9.3005
R11567 gnd.n6232 gnd.n2407 9.3005
R11568 gnd.n6235 gnd.n2406 9.3005
R11569 gnd.n6236 gnd.n2405 9.3005
R11570 gnd.n6239 gnd.n2404 9.3005
R11571 gnd.n6241 gnd.n2401 9.3005
R11572 gnd.n6244 gnd.n2400 9.3005
R11573 gnd.n6245 gnd.n2399 9.3005
R11574 gnd.n6248 gnd.n2398 9.3005
R11575 gnd.n6249 gnd.n2397 9.3005
R11576 gnd.n6252 gnd.n2396 9.3005
R11577 gnd.n6253 gnd.n2395 9.3005
R11578 gnd.n6256 gnd.n2394 9.3005
R11579 gnd.n6257 gnd.n2393 9.3005
R11580 gnd.n6260 gnd.n2392 9.3005
R11581 gnd.n6261 gnd.n2391 9.3005
R11582 gnd.n6264 gnd.n2390 9.3005
R11583 gnd.n6265 gnd.n2389 9.3005
R11584 gnd.n6268 gnd.n2388 9.3005
R11585 gnd.n6270 gnd.n2387 9.3005
R11586 gnd.n6271 gnd.n2386 9.3005
R11587 gnd.n6272 gnd.n2385 9.3005
R11588 gnd.n6273 gnd.n2384 9.3005
R11589 gnd.n6200 gnd.n2423 9.3005
R11590 gnd.n6158 gnd.n2445 9.3005
R11591 gnd.n6150 gnd.n2459 9.3005
R11592 gnd.n6149 gnd.n2460 9.3005
R11593 gnd.n6148 gnd.n2461 9.3005
R11594 gnd.n2481 gnd.n2462 9.3005
R11595 gnd.n6138 gnd.n2482 9.3005
R11596 gnd.n6137 gnd.n2483 9.3005
R11597 gnd.n6136 gnd.n2484 9.3005
R11598 gnd.n2500 gnd.n2485 9.3005
R11599 gnd.n6126 gnd.n2501 9.3005
R11600 gnd.n6125 gnd.n2502 9.3005
R11601 gnd.n6124 gnd.n2503 9.3005
R11602 gnd.n2521 gnd.n2504 9.3005
R11603 gnd.n6114 gnd.n2522 9.3005
R11604 gnd.n6113 gnd.n2523 9.3005
R11605 gnd.n6112 gnd.n2524 9.3005
R11606 gnd.n2549 gnd.n2543 9.3005
R11607 gnd.n6088 gnd.n2568 9.3005
R11608 gnd.n6087 gnd.n2569 9.3005
R11609 gnd.n6086 gnd.n2570 9.3005
R11610 gnd.n2587 gnd.n2571 9.3005
R11611 gnd.n6076 gnd.n2588 9.3005
R11612 gnd.n6075 gnd.n2589 9.3005
R11613 gnd.n6074 gnd.n2590 9.3005
R11614 gnd.n2607 gnd.n2591 9.3005
R11615 gnd.n6064 gnd.n2608 9.3005
R11616 gnd.n6063 gnd.n2609 9.3005
R11617 gnd.n6062 gnd.n2610 9.3005
R11618 gnd.n2627 gnd.n2611 9.3005
R11619 gnd.n6052 gnd.n2628 9.3005
R11620 gnd.n6051 gnd.n2629 9.3005
R11621 gnd.n6050 gnd.n2630 9.3005
R11622 gnd.n2458 gnd.n2457 9.3005
R11623 gnd.n6099 gnd.n6098 9.3005
R11624 gnd.n4073 gnd.n4072 9.3005
R11625 gnd.n4067 gnd.n4066 9.3005
R11626 gnd.n4213 gnd.n4212 9.3005
R11627 gnd.n4214 gnd.n4065 9.3005
R11628 gnd.n4217 gnd.n4216 9.3005
R11629 gnd.n4215 gnd.n4062 9.3005
R11630 gnd.n4221 gnd.n4063 9.3005
R11631 gnd.n4071 gnd.n4069 9.3005
R11632 gnd.n6378 gnd.n975 9.3005
R11633 gnd.n6379 gnd.n974 9.3005
R11634 gnd.n6380 gnd.n973 9.3005
R11635 gnd.n972 gnd.n968 9.3005
R11636 gnd.n6386 gnd.n967 9.3005
R11637 gnd.n6387 gnd.n966 9.3005
R11638 gnd.n6388 gnd.n965 9.3005
R11639 gnd.n964 gnd.n960 9.3005
R11640 gnd.n6394 gnd.n959 9.3005
R11641 gnd.n6395 gnd.n958 9.3005
R11642 gnd.n6396 gnd.n957 9.3005
R11643 gnd.n956 gnd.n952 9.3005
R11644 gnd.n6402 gnd.n951 9.3005
R11645 gnd.n6403 gnd.n950 9.3005
R11646 gnd.n6404 gnd.n949 9.3005
R11647 gnd.n948 gnd.n944 9.3005
R11648 gnd.n6410 gnd.n943 9.3005
R11649 gnd.n6411 gnd.n942 9.3005
R11650 gnd.n6412 gnd.n941 9.3005
R11651 gnd.n940 gnd.n936 9.3005
R11652 gnd.n6418 gnd.n935 9.3005
R11653 gnd.n6419 gnd.n934 9.3005
R11654 gnd.n6420 gnd.n933 9.3005
R11655 gnd.n932 gnd.n928 9.3005
R11656 gnd.n6426 gnd.n927 9.3005
R11657 gnd.n6427 gnd.n926 9.3005
R11658 gnd.n6428 gnd.n925 9.3005
R11659 gnd.n924 gnd.n920 9.3005
R11660 gnd.n6434 gnd.n919 9.3005
R11661 gnd.n6435 gnd.n918 9.3005
R11662 gnd.n6436 gnd.n917 9.3005
R11663 gnd.n916 gnd.n912 9.3005
R11664 gnd.n6442 gnd.n911 9.3005
R11665 gnd.n6443 gnd.n910 9.3005
R11666 gnd.n6444 gnd.n909 9.3005
R11667 gnd.n908 gnd.n904 9.3005
R11668 gnd.n6450 gnd.n903 9.3005
R11669 gnd.n6451 gnd.n902 9.3005
R11670 gnd.n6452 gnd.n901 9.3005
R11671 gnd.n900 gnd.n896 9.3005
R11672 gnd.n6458 gnd.n895 9.3005
R11673 gnd.n6459 gnd.n894 9.3005
R11674 gnd.n6460 gnd.n893 9.3005
R11675 gnd.n892 gnd.n888 9.3005
R11676 gnd.n6466 gnd.n887 9.3005
R11677 gnd.n6467 gnd.n886 9.3005
R11678 gnd.n6468 gnd.n885 9.3005
R11679 gnd.n884 gnd.n880 9.3005
R11680 gnd.n6474 gnd.n879 9.3005
R11681 gnd.n6475 gnd.n878 9.3005
R11682 gnd.n6476 gnd.n877 9.3005
R11683 gnd.n876 gnd.n872 9.3005
R11684 gnd.n6482 gnd.n871 9.3005
R11685 gnd.n6483 gnd.n870 9.3005
R11686 gnd.n6484 gnd.n869 9.3005
R11687 gnd.n868 gnd.n864 9.3005
R11688 gnd.n6490 gnd.n863 9.3005
R11689 gnd.n6491 gnd.n862 9.3005
R11690 gnd.n6492 gnd.n861 9.3005
R11691 gnd.n860 gnd.n856 9.3005
R11692 gnd.n6498 gnd.n855 9.3005
R11693 gnd.n6499 gnd.n854 9.3005
R11694 gnd.n6500 gnd.n853 9.3005
R11695 gnd.n852 gnd.n848 9.3005
R11696 gnd.n6506 gnd.n847 9.3005
R11697 gnd.n6507 gnd.n846 9.3005
R11698 gnd.n6508 gnd.n845 9.3005
R11699 gnd.n844 gnd.n840 9.3005
R11700 gnd.n6514 gnd.n839 9.3005
R11701 gnd.n6515 gnd.n838 9.3005
R11702 gnd.n6516 gnd.n837 9.3005
R11703 gnd.n836 gnd.n832 9.3005
R11704 gnd.n6522 gnd.n831 9.3005
R11705 gnd.n6523 gnd.n830 9.3005
R11706 gnd.n6524 gnd.n829 9.3005
R11707 gnd.n828 gnd.n824 9.3005
R11708 gnd.n6530 gnd.n823 9.3005
R11709 gnd.n6531 gnd.n822 9.3005
R11710 gnd.n6532 gnd.n821 9.3005
R11711 gnd.n820 gnd.n816 9.3005
R11712 gnd.n6538 gnd.n815 9.3005
R11713 gnd.n6539 gnd.n814 9.3005
R11714 gnd.n6540 gnd.n813 9.3005
R11715 gnd.n812 gnd.n808 9.3005
R11716 gnd.n4070 gnd.n976 9.3005
R11717 gnd.n5300 gnd.n3418 9.3005
R11718 gnd.n4400 gnd.n4399 9.3005
R11719 gnd.n4401 gnd.n3926 9.3005
R11720 gnd.n4403 gnd.n4402 9.3005
R11721 gnd.n3913 gnd.n3912 9.3005
R11722 gnd.n4416 gnd.n4415 9.3005
R11723 gnd.n4417 gnd.n3911 9.3005
R11724 gnd.n4419 gnd.n4418 9.3005
R11725 gnd.n3900 gnd.n3899 9.3005
R11726 gnd.n4432 gnd.n4431 9.3005
R11727 gnd.n4433 gnd.n3898 9.3005
R11728 gnd.n4435 gnd.n4434 9.3005
R11729 gnd.n3886 gnd.n3885 9.3005
R11730 gnd.n4448 gnd.n4447 9.3005
R11731 gnd.n4449 gnd.n3884 9.3005
R11732 gnd.n4451 gnd.n4450 9.3005
R11733 gnd.n3872 gnd.n3871 9.3005
R11734 gnd.n4464 gnd.n4463 9.3005
R11735 gnd.n4465 gnd.n3869 9.3005
R11736 gnd.n4478 gnd.n4477 9.3005
R11737 gnd.n4476 gnd.n3870 9.3005
R11738 gnd.n4475 gnd.n4474 9.3005
R11739 gnd.n4473 gnd.n4466 9.3005
R11740 gnd.n4472 gnd.n4471 9.3005
R11741 gnd.n4470 gnd.n4469 9.3005
R11742 gnd.n2994 gnd.n2992 9.3005
R11743 gnd.n5832 gnd.n5831 9.3005
R11744 gnd.n5830 gnd.n2993 9.3005
R11745 gnd.n5829 gnd.n5828 9.3005
R11746 gnd.n5827 gnd.n2995 9.3005
R11747 gnd.n5826 gnd.n5825 9.3005
R11748 gnd.n5824 gnd.n2999 9.3005
R11749 gnd.n5823 gnd.n5822 9.3005
R11750 gnd.n5821 gnd.n3000 9.3005
R11751 gnd.n5820 gnd.n5819 9.3005
R11752 gnd.n5818 gnd.n3004 9.3005
R11753 gnd.n5817 gnd.n5816 9.3005
R11754 gnd.n5815 gnd.n3005 9.3005
R11755 gnd.n5814 gnd.n5813 9.3005
R11756 gnd.n5812 gnd.n3009 9.3005
R11757 gnd.n5811 gnd.n5810 9.3005
R11758 gnd.n5809 gnd.n3010 9.3005
R11759 gnd.n5808 gnd.n5807 9.3005
R11760 gnd.n5806 gnd.n3014 9.3005
R11761 gnd.n5805 gnd.n5804 9.3005
R11762 gnd.n5803 gnd.n3015 9.3005
R11763 gnd.n5802 gnd.n5801 9.3005
R11764 gnd.n5800 gnd.n3019 9.3005
R11765 gnd.n5799 gnd.n5798 9.3005
R11766 gnd.n5797 gnd.n3020 9.3005
R11767 gnd.n5796 gnd.n5795 9.3005
R11768 gnd.n5794 gnd.n3024 9.3005
R11769 gnd.n5793 gnd.n5792 9.3005
R11770 gnd.n5791 gnd.n3025 9.3005
R11771 gnd.n5790 gnd.n5789 9.3005
R11772 gnd.n5788 gnd.n3029 9.3005
R11773 gnd.n5787 gnd.n5786 9.3005
R11774 gnd.n5785 gnd.n3030 9.3005
R11775 gnd.n5784 gnd.n5783 9.3005
R11776 gnd.n5782 gnd.n3034 9.3005
R11777 gnd.n5781 gnd.n5780 9.3005
R11778 gnd.n5779 gnd.n3035 9.3005
R11779 gnd.n5778 gnd.n5777 9.3005
R11780 gnd.n5776 gnd.n3039 9.3005
R11781 gnd.n5775 gnd.n5774 9.3005
R11782 gnd.n5773 gnd.n3040 9.3005
R11783 gnd.n5772 gnd.n5771 9.3005
R11784 gnd.n5770 gnd.n3044 9.3005
R11785 gnd.n5769 gnd.n5768 9.3005
R11786 gnd.n5767 gnd.n3045 9.3005
R11787 gnd.n5766 gnd.n5765 9.3005
R11788 gnd.n5764 gnd.n3049 9.3005
R11789 gnd.n5763 gnd.n5762 9.3005
R11790 gnd.n5761 gnd.n3050 9.3005
R11791 gnd.n5760 gnd.n5759 9.3005
R11792 gnd.n5758 gnd.n3054 9.3005
R11793 gnd.n5757 gnd.n5756 9.3005
R11794 gnd.n5755 gnd.n3055 9.3005
R11795 gnd.n5754 gnd.n5753 9.3005
R11796 gnd.n5752 gnd.n3059 9.3005
R11797 gnd.n5751 gnd.n5750 9.3005
R11798 gnd.n5749 gnd.n3060 9.3005
R11799 gnd.n5748 gnd.n5747 9.3005
R11800 gnd.n5746 gnd.n3064 9.3005
R11801 gnd.n5745 gnd.n5744 9.3005
R11802 gnd.n5743 gnd.n3065 9.3005
R11803 gnd.n5742 gnd.n5741 9.3005
R11804 gnd.n5740 gnd.n3069 9.3005
R11805 gnd.n5739 gnd.n5738 9.3005
R11806 gnd.n5737 gnd.n3070 9.3005
R11807 gnd.n5736 gnd.n5735 9.3005
R11808 gnd.n5734 gnd.n3074 9.3005
R11809 gnd.n5733 gnd.n5732 9.3005
R11810 gnd.n5731 gnd.n3075 9.3005
R11811 gnd.n5730 gnd.n5729 9.3005
R11812 gnd.n5728 gnd.n3079 9.3005
R11813 gnd.n5727 gnd.n5726 9.3005
R11814 gnd.n5725 gnd.n3080 9.3005
R11815 gnd.n5724 gnd.n5723 9.3005
R11816 gnd.n5722 gnd.n3084 9.3005
R11817 gnd.n5721 gnd.n5720 9.3005
R11818 gnd.n5719 gnd.n3085 9.3005
R11819 gnd.n3928 gnd.n3927 9.3005
R11820 gnd.n6033 gnd.n2644 9.3005
R11821 gnd.n4027 gnd.n4026 9.3005
R11822 gnd.n4284 gnd.n4283 9.3005
R11823 gnd.n4285 gnd.n4025 9.3005
R11824 gnd.n4287 gnd.n4286 9.3005
R11825 gnd.n4015 gnd.n4014 9.3005
R11826 gnd.n4320 gnd.n4319 9.3005
R11827 gnd.n4321 gnd.n4013 9.3005
R11828 gnd.n4323 gnd.n4322 9.3005
R11829 gnd.n4009 gnd.n4008 9.3005
R11830 gnd.n4334 gnd.n4333 9.3005
R11831 gnd.n4335 gnd.n4007 9.3005
R11832 gnd.n4337 gnd.n4336 9.3005
R11833 gnd.n4002 gnd.n4000 9.3005
R11834 gnd.n4361 gnd.n4360 9.3005
R11835 gnd.n4359 gnd.n4001 9.3005
R11836 gnd.n4358 gnd.n4357 9.3005
R11837 gnd.n4356 gnd.n4003 9.3005
R11838 gnd.n4355 gnd.n4354 9.3005
R11839 gnd.n2643 gnd.n2641 9.3005
R11840 gnd.n6039 gnd.n6038 9.3005
R11841 gnd.n6037 gnd.n2642 9.3005
R11842 gnd.n6011 gnd.n6010 9.3005
R11843 gnd.n6009 gnd.n6008 9.3005
R11844 gnd.n2686 gnd.n2685 9.3005
R11845 gnd.n6003 gnd.n6002 9.3005
R11846 gnd.n6001 gnd.n6000 9.3005
R11847 gnd.n2696 gnd.n2695 9.3005
R11848 gnd.n5995 gnd.n5994 9.3005
R11849 gnd.n5993 gnd.n5992 9.3005
R11850 gnd.n2704 gnd.n2703 9.3005
R11851 gnd.n5987 gnd.n5986 9.3005
R11852 gnd.n5985 gnd.n5984 9.3005
R11853 gnd.n2714 gnd.n2713 9.3005
R11854 gnd.n5979 gnd.n5978 9.3005
R11855 gnd.n5977 gnd.n5976 9.3005
R11856 gnd.n2722 gnd.n2721 9.3005
R11857 gnd.n5971 gnd.n5970 9.3005
R11858 gnd.n5969 gnd.n2736 9.3005
R11859 gnd.n5968 gnd.n2645 9.3005
R11860 gnd.n2682 gnd.n2680 9.3005
R11861 gnd.n6035 gnd.n6034 9.3005
R11862 gnd.n2735 gnd.n2646 9.3005
R11863 gnd.n2731 gnd.n2730 9.3005
R11864 gnd.n5973 gnd.n5972 9.3005
R11865 gnd.n5975 gnd.n5974 9.3005
R11866 gnd.n2718 gnd.n2717 9.3005
R11867 gnd.n5981 gnd.n5980 9.3005
R11868 gnd.n5983 gnd.n5982 9.3005
R11869 gnd.n2710 gnd.n2709 9.3005
R11870 gnd.n5989 gnd.n5988 9.3005
R11871 gnd.n5991 gnd.n5990 9.3005
R11872 gnd.n2700 gnd.n2699 9.3005
R11873 gnd.n5997 gnd.n5996 9.3005
R11874 gnd.n5999 gnd.n5998 9.3005
R11875 gnd.n2692 gnd.n2691 9.3005
R11876 gnd.n6005 gnd.n6004 9.3005
R11877 gnd.n6007 gnd.n6006 9.3005
R11878 gnd.n2681 gnd.n2679 9.3005
R11879 gnd.n6013 gnd.n6012 9.3005
R11880 gnd.n6014 gnd.n2674 9.3005
R11881 gnd.n6016 gnd.n6015 9.3005
R11882 gnd.n6018 gnd.n2673 9.3005
R11883 gnd.n6020 gnd.n6019 9.3005
R11884 gnd.n6021 gnd.n2669 9.3005
R11885 gnd.n6023 gnd.n6022 9.3005
R11886 gnd.n6024 gnd.n2668 9.3005
R11887 gnd.n6026 gnd.n6025 9.3005
R11888 gnd.n6027 gnd.n2667 9.3005
R11889 gnd.n3980 gnd.n3979 9.3005
R11890 gnd.n3978 gnd.n3932 9.3005
R11891 gnd.n3977 gnd.n3976 9.3005
R11892 gnd.n3975 gnd.n3934 9.3005
R11893 gnd.n3974 gnd.n3973 9.3005
R11894 gnd.n3972 gnd.n3937 9.3005
R11895 gnd.n3971 gnd.n3970 9.3005
R11896 gnd.n3969 gnd.n3938 9.3005
R11897 gnd.n3968 gnd.n3967 9.3005
R11898 gnd.n3966 gnd.n3941 9.3005
R11899 gnd.n3965 gnd.n3964 9.3005
R11900 gnd.n3963 gnd.n3942 9.3005
R11901 gnd.n3962 gnd.n3961 9.3005
R11902 gnd.n3960 gnd.n3945 9.3005
R11903 gnd.n3959 gnd.n3958 9.3005
R11904 gnd.n3957 gnd.n3946 9.3005
R11905 gnd.n3956 gnd.n3955 9.3005
R11906 gnd.n3954 gnd.n3949 9.3005
R11907 gnd.n3953 gnd.n3952 9.3005
R11908 gnd.n3951 gnd.n3950 9.3005
R11909 gnd.n3855 gnd.n3854 9.3005
R11910 gnd.n4496 gnd.n4495 9.3005
R11911 gnd.n4497 gnd.n3853 9.3005
R11912 gnd.n4499 gnd.n4498 9.3005
R11913 gnd.n4502 gnd.n3852 9.3005
R11914 gnd.n4504 gnd.n4503 9.3005
R11915 gnd.n4505 gnd.n3850 9.3005
R11916 gnd.n4513 gnd.n4512 9.3005
R11917 gnd.n4511 gnd.n3851 9.3005
R11918 gnd.n4510 gnd.n4509 9.3005
R11919 gnd.n4508 gnd.n4506 9.3005
R11920 gnd.n3737 gnd.n3736 9.3005
R11921 gnd.n4584 gnd.n4583 9.3005
R11922 gnd.n4585 gnd.n3734 9.3005
R11923 gnd.n4600 gnd.n4599 9.3005
R11924 gnd.n4598 gnd.n3735 9.3005
R11925 gnd.n4597 gnd.n4596 9.3005
R11926 gnd.n4595 gnd.n4586 9.3005
R11927 gnd.n4594 gnd.n4593 9.3005
R11928 gnd.n4592 gnd.n4591 9.3005
R11929 gnd.n3690 gnd.n3689 9.3005
R11930 gnd.n4668 gnd.n4667 9.3005
R11931 gnd.n4669 gnd.n3687 9.3005
R11932 gnd.n4697 gnd.n4696 9.3005
R11933 gnd.n4695 gnd.n3688 9.3005
R11934 gnd.n4694 gnd.n4693 9.3005
R11935 gnd.n4692 gnd.n4670 9.3005
R11936 gnd.n4691 gnd.n4690 9.3005
R11937 gnd.n4689 gnd.n4673 9.3005
R11938 gnd.n4688 gnd.n4687 9.3005
R11939 gnd.n4686 gnd.n4674 9.3005
R11940 gnd.n4685 gnd.n4684 9.3005
R11941 gnd.n4683 gnd.n4678 9.3005
R11942 gnd.n4682 gnd.n4681 9.3005
R11943 gnd.n3630 gnd.n3628 9.3005
R11944 gnd.n4816 gnd.n4815 9.3005
R11945 gnd.n4814 gnd.n3629 9.3005
R11946 gnd.n4813 gnd.n4812 9.3005
R11947 gnd.n4811 gnd.n3631 9.3005
R11948 gnd.n4810 gnd.n4809 9.3005
R11949 gnd.n4808 gnd.n4791 9.3005
R11950 gnd.n4807 gnd.n4806 9.3005
R11951 gnd.n4805 gnd.n4792 9.3005
R11952 gnd.n4804 gnd.n4803 9.3005
R11953 gnd.n4802 gnd.n4796 9.3005
R11954 gnd.n4801 gnd.n4800 9.3005
R11955 gnd.n4799 gnd.n4797 9.3005
R11956 gnd.n3565 gnd.n3563 9.3005
R11957 gnd.n4928 gnd.n4927 9.3005
R11958 gnd.n4926 gnd.n3564 9.3005
R11959 gnd.n4925 gnd.n4924 9.3005
R11960 gnd.n4923 gnd.n3566 9.3005
R11961 gnd.n4922 gnd.n4921 9.3005
R11962 gnd.n4920 gnd.n4917 9.3005
R11963 gnd.n4919 gnd.n4918 9.3005
R11964 gnd.n3514 gnd.n3513 9.3005
R11965 gnd.n5180 gnd.n5179 9.3005
R11966 gnd.n5181 gnd.n3512 9.3005
R11967 gnd.n5183 gnd.n5182 9.3005
R11968 gnd.n3504 gnd.n3503 9.3005
R11969 gnd.n5198 gnd.n5197 9.3005
R11970 gnd.n5199 gnd.n3502 9.3005
R11971 gnd.n5201 gnd.n5200 9.3005
R11972 gnd.n3492 gnd.n3491 9.3005
R11973 gnd.n5215 gnd.n5214 9.3005
R11974 gnd.n5216 gnd.n3490 9.3005
R11975 gnd.n5218 gnd.n5217 9.3005
R11976 gnd.n3480 gnd.n3479 9.3005
R11977 gnd.n5232 gnd.n5231 9.3005
R11978 gnd.n5233 gnd.n3478 9.3005
R11979 gnd.n5235 gnd.n5234 9.3005
R11980 gnd.n3467 gnd.n3466 9.3005
R11981 gnd.n5249 gnd.n5248 9.3005
R11982 gnd.n5250 gnd.n3465 9.3005
R11983 gnd.n5252 gnd.n5251 9.3005
R11984 gnd.n3456 gnd.n3455 9.3005
R11985 gnd.n5269 gnd.n5268 9.3005
R11986 gnd.n5270 gnd.n3454 9.3005
R11987 gnd.n5272 gnd.n5271 9.3005
R11988 gnd.n3094 gnd.n3093 9.3005
R11989 gnd.n5715 gnd.n5714 9.3005
R11990 gnd.n3933 gnd.n3931 9.3005
R11991 gnd.n5711 gnd.n3095 9.3005
R11992 gnd.n5710 gnd.n5709 9.3005
R11993 gnd.n5708 gnd.n3098 9.3005
R11994 gnd.n5707 gnd.n5706 9.3005
R11995 gnd.n5705 gnd.n3099 9.3005
R11996 gnd.n5704 gnd.n5703 9.3005
R11997 gnd.n5713 gnd.n5712 9.3005
R11998 gnd.n5656 gnd.n5655 9.3005
R11999 gnd.n3146 gnd.n3145 9.3005
R12000 gnd.n5662 gnd.n5661 9.3005
R12001 gnd.n5664 gnd.n5663 9.3005
R12002 gnd.n3138 gnd.n3137 9.3005
R12003 gnd.n5670 gnd.n5669 9.3005
R12004 gnd.n5672 gnd.n5671 9.3005
R12005 gnd.n3130 gnd.n3129 9.3005
R12006 gnd.n5678 gnd.n5677 9.3005
R12007 gnd.n5680 gnd.n5679 9.3005
R12008 gnd.n3122 gnd.n3121 9.3005
R12009 gnd.n5686 gnd.n5685 9.3005
R12010 gnd.n5688 gnd.n5687 9.3005
R12011 gnd.n3114 gnd.n3113 9.3005
R12012 gnd.n5694 gnd.n5693 9.3005
R12013 gnd.n5696 gnd.n5695 9.3005
R12014 gnd.n3110 gnd.n3105 9.3005
R12015 gnd.n5654 gnd.n3155 9.3005
R12016 gnd.n3419 gnd.n3154 9.3005
R12017 gnd.n5701 gnd.n3103 9.3005
R12018 gnd.n5700 gnd.n5699 9.3005
R12019 gnd.n5698 gnd.n5697 9.3005
R12020 gnd.n3109 gnd.n3108 9.3005
R12021 gnd.n5692 gnd.n5691 9.3005
R12022 gnd.n5690 gnd.n5689 9.3005
R12023 gnd.n3118 gnd.n3117 9.3005
R12024 gnd.n5684 gnd.n5683 9.3005
R12025 gnd.n5682 gnd.n5681 9.3005
R12026 gnd.n3126 gnd.n3125 9.3005
R12027 gnd.n5676 gnd.n5675 9.3005
R12028 gnd.n5674 gnd.n5673 9.3005
R12029 gnd.n3134 gnd.n3133 9.3005
R12030 gnd.n5668 gnd.n5667 9.3005
R12031 gnd.n5666 gnd.n5665 9.3005
R12032 gnd.n3142 gnd.n3141 9.3005
R12033 gnd.n5660 gnd.n5659 9.3005
R12034 gnd.n5658 gnd.n5657 9.3005
R12035 gnd.n3442 gnd.n3152 9.3005
R12036 gnd.n3421 gnd.n3420 9.3005
R12037 gnd.n5302 gnd.n5301 9.3005
R12038 gnd.n5343 gnd.n5342 9.3005
R12039 gnd.n5341 gnd.n3417 9.3005
R12040 gnd.n5340 gnd.n5339 9.3005
R12041 gnd.n5338 gnd.n5305 9.3005
R12042 gnd.n5337 gnd.n5336 9.3005
R12043 gnd.n5335 gnd.n5309 9.3005
R12044 gnd.n5334 gnd.n5333 9.3005
R12045 gnd.n5332 gnd.n5310 9.3005
R12046 gnd.n5331 gnd.n5330 9.3005
R12047 gnd.n3400 gnd.n3399 9.3005
R12048 gnd.n5391 gnd.n5390 9.3005
R12049 gnd.n5392 gnd.n3398 9.3005
R12050 gnd.n5394 gnd.n5393 9.3005
R12051 gnd.n3395 gnd.n3394 9.3005
R12052 gnd.n5406 gnd.n5405 9.3005
R12053 gnd.n5407 gnd.n3392 9.3005
R12054 gnd.n5413 gnd.n5412 9.3005
R12055 gnd.n5411 gnd.n3393 9.3005
R12056 gnd.n5410 gnd.n5409 9.3005
R12057 gnd.n5408 gnd.n67 9.3005
R12058 gnd.n5304 gnd.n3416 9.3005
R12059 gnd.n7418 gnd.n68 9.3005
R12060 gnd.t156 gnd.n1201 9.24152
R12061 gnd.n6346 gnd.t43 9.24152
R12062 gnd.n2331 gnd.t133 9.24152
R12063 gnd.n4010 gnd.t279 9.24152
R12064 gnd.n3759 gnd.t176 9.24152
R12065 gnd.n4913 gnd.t192 9.24152
R12066 gnd.n4949 gnd.t192 9.24152
R12067 gnd.n5387 gnd.t239 9.24152
R12068 gnd.t333 gnd.t156 8.92286
R12069 gnd.n4655 gnd.t14 8.92286
R12070 gnd.n4648 gnd.t185 8.92286
R12071 gnd.n4838 gnd.t187 8.92286
R12072 gnd.n4857 gnd.t174 8.92286
R12073 gnd.n2311 gnd.n2286 8.92171
R12074 gnd.n2279 gnd.n2254 8.92171
R12075 gnd.n2247 gnd.n2222 8.92171
R12076 gnd.n2216 gnd.n2191 8.92171
R12077 gnd.n2184 gnd.n2159 8.92171
R12078 gnd.n2152 gnd.n2127 8.92171
R12079 gnd.n2120 gnd.n2095 8.92171
R12080 gnd.n2089 gnd.n2064 8.92171
R12081 gnd.n4988 gnd.n4970 8.72777
R12082 gnd.t28 gnd.n1246 8.60421
R12083 gnd.t225 gnd.n4029 8.60421
R12084 gnd.t158 gnd.n3664 8.60421
R12085 gnd.n4757 gnd.t198 8.60421
R12086 gnd.n5466 gnd.t252 8.60421
R12087 gnd.n1618 gnd.n1606 8.43656
R12088 gnd.n42 gnd.n30 8.43656
R12089 gnd.n4530 gnd.n3760 8.28555
R12090 gnd.n4619 gnd.n3719 8.28555
R12091 gnd.n4633 gnd.n3669 8.28555
R12092 gnd.n4778 gnd.n4777 8.28555
R12093 gnd.n4866 gnd.n4865 8.28555
R12094 gnd.n4948 gnd.n3547 8.28555
R12095 gnd.n2312 gnd.n2284 8.14595
R12096 gnd.n2280 gnd.n2252 8.14595
R12097 gnd.n2248 gnd.n2220 8.14595
R12098 gnd.n2217 gnd.n2189 8.14595
R12099 gnd.n2185 gnd.n2157 8.14595
R12100 gnd.n2153 gnd.n2125 8.14595
R12101 gnd.n2121 gnd.n2093 8.14595
R12102 gnd.n2090 gnd.n2062 8.14595
R12103 gnd.n4256 gnd.n0 8.10675
R12104 gnd.n7419 gnd.n7418 8.10675
R12105 gnd.n2317 gnd.n2316 7.97301
R12106 gnd.n1840 gnd.t26 7.9669
R12107 gnd.t266 gnd.n2527 7.9669
R12108 gnd.n6030 gnd.n2649 7.9669
R12109 gnd.t202 gnd.n2987 7.9669
R12110 gnd.t97 gnd.t6 7.9669
R12111 gnd.n5297 gnd.n5296 7.9669
R12112 gnd.n7225 gnd.t221 7.9669
R12113 gnd.n7419 gnd.n66 7.78567
R12114 gnd.n5654 gnd.n3154 7.75808
R12115 gnd.n5969 gnd.n5968 7.75808
R12116 gnd.n7325 gnd.n7263 7.75808
R12117 gnd.n4150 gnd.n4149 7.75808
R12118 gnd.t8 gnd.n3725 7.64824
R12119 gnd.n4881 gnd.t2 7.64824
R12120 gnd.n1643 gnd.n1642 7.53171
R12121 gnd.t168 gnd.n1789 7.32958
R12122 gnd.t80 gnd.n3923 7.32958
R12123 gnd.n4437 gnd.t23 7.32958
R12124 gnd.t162 gnd.n3476 7.32958
R12125 gnd.n5275 gnd.t54 7.32958
R12126 gnd.n2970 gnd.n2969 7.30353
R12127 gnd.n4987 gnd.n4986 7.30353
R12128 gnd.n1748 gnd.n1747 7.01093
R12129 gnd.n1759 gnd.n1356 7.01093
R12130 gnd.n1758 gnd.n1359 7.01093
R12131 gnd.n1769 gnd.n1349 7.01093
R12132 gnd.n1667 gnd.n1342 7.01093
R12133 gnd.n1779 gnd.n1778 7.01093
R12134 gnd.n1790 gnd.n1331 7.01093
R12135 gnd.n1789 gnd.n1334 7.01093
R12136 gnd.n1800 gnd.n1322 7.01093
R12137 gnd.n1325 gnd.n1323 7.01093
R12138 gnd.n1810 gnd.n1809 7.01093
R12139 gnd.n1821 gnd.n1305 7.01093
R12140 gnd.n1831 gnd.n1296 7.01093
R12141 gnd.n1299 gnd.n1297 7.01093
R12142 gnd.n1841 gnd.n1840 7.01093
R12143 gnd.n1852 gnd.n1279 7.01093
R12144 gnd.n1862 gnd.n1271 7.01093
R12145 gnd.n1272 gnd.n1264 7.01093
R12146 gnd.n1883 gnd.n1253 7.01093
R12147 gnd.n1882 gnd.n1256 7.01093
R12148 gnd.n1893 gnd.n1246 7.01093
R12149 gnd.n1583 gnd.n1239 7.01093
R12150 gnd.n1903 gnd.n1902 7.01093
R12151 gnd.n1914 gnd.n1228 7.01093
R12152 gnd.n1913 gnd.n1231 7.01093
R12153 gnd.n1221 gnd.n1214 7.01093
R12154 gnd.n1934 gnd.n1933 7.01093
R12155 gnd.n1944 gnd.n1201 7.01093
R12156 gnd.n1943 gnd.n1204 7.01093
R12157 gnd.n1952 gnd.n1195 7.01093
R12158 gnd.n1966 gnd.n1186 7.01093
R12159 gnd.n2014 gnd.n1179 7.01093
R12160 gnd.n1173 gnd.n1171 7.01093
R12161 gnd.n2039 gnd.n2038 7.01093
R12162 gnd.n1154 gnd.n980 7.01093
R12163 gnd.n6368 gnd.n989 7.01093
R12164 gnd.n6367 gnd.n992 7.01093
R12165 gnd.n6361 gnd.n6360 7.01093
R12166 gnd.n1151 gnd.n1004 7.01093
R12167 gnd.n6354 gnd.n1015 7.01093
R12168 gnd.n6353 gnd.n1018 7.01093
R12169 gnd.n1989 gnd.n1027 7.01093
R12170 gnd.n6347 gnd.n6346 7.01093
R12171 gnd.n2332 gnd.n2331 7.01093
R12172 gnd.n6340 gnd.n1040 7.01093
R12173 gnd.n6339 gnd.n1043 7.01093
R12174 gnd.n3769 gnd.t73 7.01093
R12175 gnd.n4558 gnd.t30 7.01093
R12176 gnd.n4571 gnd.n3747 7.01093
R12177 gnd.n4611 gnd.n4610 7.01093
R12178 gnd.n4733 gnd.n3665 7.01093
R12179 gnd.n4769 gnd.n4768 7.01093
R12180 gnd.n4882 gnd.n3583 7.01093
R12181 gnd.n4938 gnd.n4937 7.01093
R12182 gnd.n4911 gnd.t4 7.01093
R12183 gnd.n4962 gnd.t62 7.01093
R12184 gnd.n1325 gnd.t155 6.69227
R12185 gnd.n1934 gnd.t333 6.69227
R12186 gnd.t186 gnd.n1001 6.69227
R12187 gnd.n5092 gnd.n5091 6.5566
R12188 gnd.n3778 gnd.n3777 6.5566
R12189 gnd.n5852 gnd.n5848 6.5566
R12190 gnd.n5107 gnd.n5106 6.5566
R12191 gnd.t127 gnd.n3754 6.37362
R12192 gnd.n4706 gnd.t184 6.37362
R12193 gnd.n4819 gnd.t13 6.37362
R12194 gnd.n2730 gnd.n2728 6.20656
R12195 gnd.n3442 gnd.n3151 6.20656
R12196 gnd.n1851 gnd.t194 6.05496
R12197 gnd.n1282 gnd.t206 6.05496
R12198 gnd.n1583 gnd.t31 6.05496
R12199 gnd.t166 gnd.n1168 6.05496
R12200 gnd.n3665 gnd.t158 6.05496
R12201 gnd.n4769 gnd.t198 6.05496
R12202 gnd.n2314 gnd.n2284 5.81868
R12203 gnd.n2282 gnd.n2252 5.81868
R12204 gnd.n2250 gnd.n2220 5.81868
R12205 gnd.n2219 gnd.n2189 5.81868
R12206 gnd.n2187 gnd.n2157 5.81868
R12207 gnd.n2155 gnd.n2125 5.81868
R12208 gnd.n2123 gnd.n2093 5.81868
R12209 gnd.n2092 gnd.n2062 5.81868
R12210 gnd.n4500 gnd.t121 5.73631
R12211 gnd.n4581 gnd.n3739 5.73631
R12212 gnd.n4536 gnd.n4535 5.73631
R12213 gnd.n4740 gnd.n3653 5.73631
R12214 gnd.n3655 gnd.n3648 5.73631
R12215 gnd.n4893 gnd.n4892 5.73631
R12216 gnd.n3569 gnd.n3560 5.73631
R12217 gnd.n5015 gnd.n3231 5.62001
R12218 gnd.n5914 gnd.n2912 5.62001
R12219 gnd.n5914 gnd.n2913 5.62001
R12220 gnd.n5101 gnd.n3231 5.62001
R12221 gnd.n1453 gnd.n1452 5.4308
R12222 gnd.n1144 gnd.n1074 5.4308
R12223 gnd.n1903 gnd.t175 5.41765
R12224 gnd.n1924 gnd.t10 5.41765
R12225 gnd.t170 gnd.n2025 5.41765
R12226 gnd.n5911 gnd.n2916 5.41765
R12227 gnd.t47 gnd.n2948 5.09899
R12228 gnd.t121 gnd.n2977 5.09899
R12229 gnd.n2312 gnd.n2311 5.04292
R12230 gnd.n2280 gnd.n2279 5.04292
R12231 gnd.n2248 gnd.n2247 5.04292
R12232 gnd.n2217 gnd.n2216 5.04292
R12233 gnd.n2185 gnd.n2184 5.04292
R12234 gnd.n2153 gnd.n2152 5.04292
R12235 gnd.n2121 gnd.n2120 5.04292
R12236 gnd.n2090 gnd.n2089 5.04292
R12237 gnd.n1872 gnd.t9 4.78034
R12238 gnd.n1952 gnd.t27 4.78034
R12239 gnd.t188 gnd.n3874 4.78034
R12240 gnd.n4536 gnd.t196 4.78034
R12241 gnd.t172 gnd.n4893 4.78034
R12242 gnd.n4991 gnd.t112 4.78034
R12243 gnd.n5212 gnd.t209 4.78034
R12244 gnd.n1646 gnd.n1645 4.74817
R12245 gnd.n1595 gnd.n1591 4.74817
R12246 gnd.n1588 gnd.n1587 4.74817
R12247 gnd.n1582 gnd.n1561 4.74817
R12248 gnd.n1645 gnd.n1559 4.74817
R12249 gnd.n1595 gnd.n1594 4.74817
R12250 gnd.n1590 gnd.n1588 4.74817
R12251 gnd.n1586 gnd.n1561 4.74817
R12252 gnd.n5469 gnd.n86 4.74817
R12253 gnd.n3367 gnd.n85 4.74817
R12254 gnd.n3376 gnd.n84 4.74817
R12255 gnd.n7411 gnd.n79 4.74817
R12256 gnd.n7409 gnd.n80 4.74817
R12257 gnd.n5480 gnd.n86 4.74817
R12258 gnd.n5470 gnd.n85 4.74817
R12259 gnd.n3366 gnd.n84 4.74817
R12260 gnd.n3375 gnd.n79 4.74817
R12261 gnd.n7410 gnd.n7409 4.74817
R12262 gnd.n4223 gnd.n4222 4.74817
R12263 gnd.n4235 gnd.n4234 4.74817
R12264 gnd.n4230 gnd.n4226 4.74817
R12265 gnd.n4228 gnd.n4227 4.74817
R12266 gnd.n4293 gnd.n4019 4.74817
R12267 gnd.n5377 gnd.n5376 4.74817
R12268 gnd.n5464 gnd.n3372 4.74817
R12269 gnd.n5462 gnd.n5461 4.74817
R12270 gnd.n5446 gnd.n5445 4.74817
R12271 gnd.n5448 gnd.n5447 4.74817
R12272 gnd.n5378 gnd.n5377 4.74817
R12273 gnd.n5374 gnd.n3372 4.74817
R12274 gnd.n5463 gnd.n5462 4.74817
R12275 gnd.n5445 gnd.n3373 4.74817
R12276 gnd.n5449 gnd.n5448 4.74817
R12277 gnd.n6102 gnd.n2541 4.74817
R12278 gnd.n6100 gnd.n2542 4.74817
R12279 gnd.n4034 gnd.n2547 4.74817
R12280 gnd.n4279 gnd.n2546 4.74817
R12281 gnd.n2548 gnd.n2545 4.74817
R12282 gnd.n2541 gnd.n2525 4.74817
R12283 gnd.n6101 gnd.n6100 4.74817
R12284 gnd.n4056 gnd.n2547 4.74817
R12285 gnd.n4035 gnd.n2546 4.74817
R12286 gnd.n4278 gnd.n2545 4.74817
R12287 gnd.n4237 gnd.n4223 4.74817
R12288 gnd.n4236 gnd.n4235 4.74817
R12289 gnd.n4226 gnd.n4224 4.74817
R12290 gnd.n4229 gnd.n4228 4.74817
R12291 gnd.n4021 gnd.n4019 4.74817
R12292 gnd.n1642 gnd.n1641 4.74296
R12293 gnd.n66 gnd.n65 4.74296
R12294 gnd.n1618 gnd.n1617 4.7074
R12295 gnd.n1630 gnd.n1629 4.7074
R12296 gnd.n42 gnd.n41 4.7074
R12297 gnd.n54 gnd.n53 4.7074
R12298 gnd.n1642 gnd.n1630 4.65959
R12299 gnd.n66 gnd.n54 4.65959
R12300 gnd.n5596 gnd.n3233 4.6132
R12301 gnd.n5915 gnd.n2911 4.6132
R12302 gnd.n2974 gnd.t47 4.46168
R12303 gnd.n4551 gnd.n4550 4.46168
R12304 gnd.t3 gnd.n3740 4.46168
R12305 gnd.n4604 gnd.n4603 4.46168
R12306 gnd.n4741 gnd.n3659 4.46168
R12307 gnd.n4759 gnd.n4758 4.46168
R12308 gnd.n4894 gnd.n3573 4.46168
R12309 gnd.n4900 gnd.t182 4.46168
R12310 gnd.n4931 gnd.n4930 4.46168
R12311 gnd.n4983 gnd.n4970 4.46111
R12312 gnd.n2297 gnd.n2293 4.38594
R12313 gnd.n2265 gnd.n2261 4.38594
R12314 gnd.n2233 gnd.n2229 4.38594
R12315 gnd.n2202 gnd.n2198 4.38594
R12316 gnd.n2170 gnd.n2166 4.38594
R12317 gnd.n2138 gnd.n2134 4.38594
R12318 gnd.n2106 gnd.n2102 4.38594
R12319 gnd.n2075 gnd.n2071 4.38594
R12320 gnd.n2308 gnd.n2286 4.26717
R12321 gnd.n2276 gnd.n2254 4.26717
R12322 gnd.n2244 gnd.n2222 4.26717
R12323 gnd.n2213 gnd.n2191 4.26717
R12324 gnd.n2181 gnd.n2159 4.26717
R12325 gnd.n2149 gnd.n2127 4.26717
R12326 gnd.n2117 gnd.n2095 4.26717
R12327 gnd.n2086 gnd.n2064 4.26717
R12328 gnd.t205 gnd.n1308 4.14303
R12329 gnd.n1154 gnd.t154 4.14303
R12330 gnd.n2640 gnd.t66 4.14303
R12331 gnd.n5346 gnd.t50 4.14303
R12332 gnd.n2316 gnd.n2315 4.08274
R12333 gnd.n5091 gnd.n5090 4.05904
R12334 gnd.n3779 gnd.n3778 4.05904
R12335 gnd.n5855 gnd.n5848 4.05904
R12336 gnd.n5108 gnd.n5107 4.05904
R12337 gnd.n19 gnd.n9 3.99943
R12338 gnd.n3664 gnd.t157 3.82437
R12339 gnd.t183 gnd.n4757 3.82437
R12340 gnd.n1644 gnd.n1643 3.81325
R12341 gnd.n1630 gnd.n1618 3.72967
R12342 gnd.n54 gnd.n42 3.72967
R12343 gnd.n2316 gnd.n2188 3.70378
R12344 gnd.n19 gnd.n18 3.60163
R12345 gnd.n6375 gnd.n978 3.50571
R12346 gnd.n6375 gnd.n6374 3.50571
R12347 gnd.n2307 gnd.n2288 3.49141
R12348 gnd.n2275 gnd.n2256 3.49141
R12349 gnd.n2243 gnd.n2224 3.49141
R12350 gnd.n2212 gnd.n2193 3.49141
R12351 gnd.n2180 gnd.n2161 3.49141
R12352 gnd.n2148 gnd.n2129 3.49141
R12353 gnd.n2116 gnd.n2097 3.49141
R12354 gnd.n2085 gnd.n2066 3.49141
R12355 gnd.n5614 gnd.n5613 3.29747
R12356 gnd.n5613 gnd.n5612 3.29747
R12357 gnd.n285 gnd.n221 3.29747
R12358 gnd.n280 gnd.n221 3.29747
R12359 gnd.n6241 gnd.n6240 3.29747
R12360 gnd.n6240 gnd.n6239 3.29747
R12361 gnd.n5933 gnd.n5932 3.29747
R12362 gnd.n5932 gnd.n5931 3.29747
R12363 gnd.n4558 gnd.n3754 3.18706
R12364 gnd.n4700 gnd.t34 3.18706
R12365 gnd.n4726 gnd.n3663 3.18706
R12366 gnd.n4679 gnd.n3643 3.18706
R12367 gnd.n4828 gnd.t169 3.18706
R12368 gnd.n4913 gnd.n4911 3.18706
R12369 gnd.n1820 gnd.t205 2.8684
R12370 gnd.t248 gnd.n2509 2.8684
R12371 gnd.n4500 gnd.t202 2.8684
R12372 gnd.t176 gnd.t127 2.8684
R12373 gnd.t6 gnd.n3526 2.8684
R12374 gnd.n392 gnd.t227 2.8684
R12375 gnd.n1631 gnd.t289 2.82907
R12376 gnd.n1631 gnd.t330 2.82907
R12377 gnd.n1633 gnd.t255 2.82907
R12378 gnd.n1633 gnd.t322 2.82907
R12379 gnd.n1635 gnd.t220 2.82907
R12380 gnd.n1635 gnd.t308 2.82907
R12381 gnd.n1637 gnd.t325 2.82907
R12382 gnd.n1637 gnd.t250 2.82907
R12383 gnd.n1639 gnd.t277 2.82907
R12384 gnd.n1639 gnd.t260 2.82907
R12385 gnd.n1596 gnd.t294 2.82907
R12386 gnd.n1596 gnd.t306 2.82907
R12387 gnd.n1598 gnd.t314 2.82907
R12388 gnd.n1598 gnd.t326 2.82907
R12389 gnd.n1600 gnd.t286 2.82907
R12390 gnd.n1600 gnd.t298 2.82907
R12391 gnd.n1602 gnd.t307 2.82907
R12392 gnd.n1602 gnd.t234 2.82907
R12393 gnd.n1604 gnd.t297 2.82907
R12394 gnd.n1604 gnd.t293 2.82907
R12395 gnd.n1607 gnd.t280 2.82907
R12396 gnd.n1607 gnd.t269 2.82907
R12397 gnd.n1609 gnd.t270 2.82907
R12398 gnd.n1609 gnd.t292 2.82907
R12399 gnd.n1611 gnd.t247 2.82907
R12400 gnd.n1611 gnd.t278 2.82907
R12401 gnd.n1613 gnd.t281 2.82907
R12402 gnd.n1613 gnd.t262 2.82907
R12403 gnd.n1615 gnd.t218 2.82907
R12404 gnd.n1615 gnd.t249 2.82907
R12405 gnd.n1619 gnd.t318 2.82907
R12406 gnd.n1619 gnd.t285 2.82907
R12407 gnd.n1621 gnd.t302 2.82907
R12408 gnd.n1621 gnd.t264 2.82907
R12409 gnd.n1623 gnd.t288 2.82907
R12410 gnd.n1623 gnd.t226 2.82907
R12411 gnd.n1625 gnd.t267 2.82907
R12412 gnd.n1625 gnd.t300 2.82907
R12413 gnd.n1627 gnd.t312 2.82907
R12414 gnd.n1627 gnd.t304 2.82907
R12415 gnd.n63 gnd.t329 2.82907
R12416 gnd.n63 gnd.t246 2.82907
R12417 gnd.n61 gnd.t327 2.82907
R12418 gnd.n61 gnd.t303 2.82907
R12419 gnd.n59 gnd.t287 2.82907
R12420 gnd.n59 gnd.t320 2.82907
R12421 gnd.n57 gnd.t301 2.82907
R12422 gnd.n57 gnd.t328 2.82907
R12423 gnd.n55 gnd.t311 2.82907
R12424 gnd.n55 gnd.t240 2.82907
R12425 gnd.n28 gnd.t309 2.82907
R12426 gnd.n28 gnd.t290 2.82907
R12427 gnd.n26 gnd.t276 2.82907
R12428 gnd.n26 gnd.t324 2.82907
R12429 gnd.n24 gnd.t317 2.82907
R12430 gnd.n24 gnd.t265 2.82907
R12431 gnd.n22 gnd.t245 2.82907
R12432 gnd.n22 gnd.t212 2.82907
R12433 gnd.n20 gnd.t323 2.82907
R12434 gnd.n20 gnd.t310 2.82907
R12435 gnd.n39 gnd.t228 2.82907
R12436 gnd.n39 gnd.t236 2.82907
R12437 gnd.n37 gnd.t238 2.82907
R12438 gnd.n37 gnd.t256 2.82907
R12439 gnd.n35 gnd.t253 2.82907
R12440 gnd.n35 gnd.t273 2.82907
R12441 gnd.n33 gnd.t271 2.82907
R12442 gnd.n33 gnd.t244 2.82907
R12443 gnd.n31 gnd.t243 2.82907
R12444 gnd.n31 gnd.t251 2.82907
R12445 gnd.n51 gnd.t282 2.82907
R12446 gnd.n51 gnd.t299 2.82907
R12447 gnd.n49 gnd.t274 2.82907
R12448 gnd.n49 gnd.t222 2.82907
R12449 gnd.n47 gnd.t316 2.82907
R12450 gnd.n47 gnd.t259 2.82907
R12451 gnd.n45 gnd.t214 2.82907
R12452 gnd.n45 gnd.t275 2.82907
R12453 gnd.n43 gnd.t232 2.82907
R12454 gnd.n43 gnd.t295 2.82907
R12455 gnd.n2304 gnd.n2303 2.71565
R12456 gnd.n2272 gnd.n2271 2.71565
R12457 gnd.n2240 gnd.n2239 2.71565
R12458 gnd.n2209 gnd.n2208 2.71565
R12459 gnd.n2177 gnd.n2176 2.71565
R12460 gnd.n2145 gnd.n2144 2.71565
R12461 gnd.n2113 gnd.n2112 2.71565
R12462 gnd.n2082 gnd.n2081 2.71565
R12463 gnd.n4515 gnd.t77 2.54975
R12464 gnd.t204 gnd.n4726 2.54975
R12465 gnd.n4679 gnd.t5 2.54975
R12466 gnd.n3547 gnd.t70 2.54975
R12467 gnd.n1645 gnd.n1644 2.27742
R12468 gnd.n1644 gnd.n1595 2.27742
R12469 gnd.n1644 gnd.n1588 2.27742
R12470 gnd.n1644 gnd.n1561 2.27742
R12471 gnd.n7408 gnd.n86 2.27742
R12472 gnd.n7408 gnd.n85 2.27742
R12473 gnd.n7408 gnd.n84 2.27742
R12474 gnd.n7408 gnd.n79 2.27742
R12475 gnd.n7409 gnd.n7408 2.27742
R12476 gnd.n5377 gnd.n83 2.27742
R12477 gnd.n3372 gnd.n83 2.27742
R12478 gnd.n5462 gnd.n83 2.27742
R12479 gnd.n5445 gnd.n83 2.27742
R12480 gnd.n5448 gnd.n83 2.27742
R12481 gnd.n6099 gnd.n2541 2.27742
R12482 gnd.n6100 gnd.n6099 2.27742
R12483 gnd.n6099 gnd.n2547 2.27742
R12484 gnd.n6099 gnd.n2546 2.27742
R12485 gnd.n6099 gnd.n2545 2.27742
R12486 gnd.n4223 gnd.n2544 2.27742
R12487 gnd.n4235 gnd.n2544 2.27742
R12488 gnd.n4226 gnd.n2544 2.27742
R12489 gnd.n4228 gnd.n2544 2.27742
R12490 gnd.n4019 gnd.n2544 2.27742
R12491 gnd.t87 gnd.n1758 2.23109
R12492 gnd.t9 gnd.n1871 2.23109
R12493 gnd.t219 gnd.n4054 2.23109
R12494 gnd.t258 gnd.n73 2.23109
R12495 gnd.n2300 gnd.n2290 1.93989
R12496 gnd.n2268 gnd.n2258 1.93989
R12497 gnd.n2236 gnd.n2226 1.93989
R12498 gnd.n2205 gnd.n2195 1.93989
R12499 gnd.n2173 gnd.n2163 1.93989
R12500 gnd.n2141 gnd.n2131 1.93989
R12501 gnd.n2109 gnd.n2099 1.93989
R12502 gnd.n2078 gnd.n2068 1.93989
R12503 gnd.n4523 gnd.n4515 1.91244
R12504 gnd.n3728 gnd.t11 1.91244
R12505 gnd.n4665 gnd.t185 1.91244
R12506 gnd.n4707 gnd.n4706 1.91244
R12507 gnd.n4819 gnd.n4818 1.91244
R12508 gnd.t187 gnd.n4837 1.91244
R12509 gnd.n4873 gnd.t20 1.91244
R12510 gnd.n4956 gnd.n3541 1.91244
R12511 gnd.n1667 gnd.t164 1.59378
R12512 gnd.n1575 gnd.t10 1.59378
R12513 gnd.n2026 gnd.t170 1.59378
R12514 gnd.n4316 gnd.t263 1.59378
R12515 gnd.n4589 gnd.t331 1.59378
R12516 gnd.t178 gnd.n3603 1.59378
R12517 gnd.n3396 gnd.t213 1.59378
R12518 gnd.t11 gnd.n3716 1.27512
R12519 gnd.n4794 gnd.t20 1.27512
R12520 gnd.n1454 gnd.n1453 1.16414
R12521 gnd.n1141 gnd.n1074 1.16414
R12522 gnd.n2299 gnd.n2292 1.16414
R12523 gnd.n2267 gnd.n2260 1.16414
R12524 gnd.n2235 gnd.n2228 1.16414
R12525 gnd.n2204 gnd.n2197 1.16414
R12526 gnd.n2172 gnd.n2165 1.16414
R12527 gnd.n2140 gnd.n2133 1.16414
R12528 gnd.n2108 gnd.n2101 1.16414
R12529 gnd.n2077 gnd.n2070 1.16414
R12530 gnd.n5596 gnd.n5595 0.970197
R12531 gnd.n5915 gnd.n2813 0.970197
R12532 gnd.n2283 gnd.n2251 0.962709
R12533 gnd.n2315 gnd.n2283 0.962709
R12534 gnd.n2156 gnd.n2124 0.962709
R12535 gnd.n2188 gnd.n2156 0.962709
R12536 gnd.t194 gnd.n1282 0.956468
R12537 gnd.n2013 gnd.t166 0.956468
R12538 gnd.n6128 gnd.t217 0.956468
R12539 gnd.n4339 gnd.t268 0.956468
R12540 gnd.n4364 gnd.t223 0.956468
R12541 gnd.t200 gnd.t34 0.956468
R12542 gnd.t18 gnd.t169 0.956468
R12543 gnd.n5318 gnd.t229 0.956468
R12544 gnd.n5328 gnd.t231 0.956468
R12545 gnd.n7248 gnd.t235 0.956468
R12546 gnd.n2 gnd.n1 0.672012
R12547 gnd.n3 gnd.n2 0.672012
R12548 gnd.n4 gnd.n3 0.672012
R12549 gnd.n5 gnd.n4 0.672012
R12550 gnd.n6 gnd.n5 0.672012
R12551 gnd.n7 gnd.n6 0.672012
R12552 gnd.n8 gnd.n7 0.672012
R12553 gnd.n9 gnd.n8 0.672012
R12554 gnd.n11 gnd.n10 0.672012
R12555 gnd.n12 gnd.n11 0.672012
R12556 gnd.n13 gnd.n12 0.672012
R12557 gnd.n14 gnd.n13 0.672012
R12558 gnd.n15 gnd.n14 0.672012
R12559 gnd.n16 gnd.n15 0.672012
R12560 gnd.n17 gnd.n16 0.672012
R12561 gnd.n18 gnd.n17 0.672012
R12562 gnd.n5841 gnd.n5840 0.637812
R12563 gnd.n5834 gnd.n2989 0.637812
R12564 gnd.n4550 gnd.t15 0.637812
R12565 gnd.t14 gnd.n4654 0.637812
R12566 gnd.n3708 gnd.n3702 0.637812
R12567 gnd.n4642 gnd.n4641 0.637812
R12568 gnd.n4788 gnd.n4787 0.637812
R12569 gnd.n4850 gnd.n3607 0.637812
R12570 gnd.n4849 gnd.t174 0.637812
R12571 gnd.n4930 gnd.t12 0.637812
R12572 gnd.n5169 gnd.n3523 0.637812
R12573 gnd.n5177 gnd.n3517 0.637812
R12574 gnd.n5187 gnd.t112 0.637812
R12575 gnd gnd.n0 0.624033
R12576 gnd.n1641 gnd.n1640 0.573776
R12577 gnd.n1640 gnd.n1638 0.573776
R12578 gnd.n1638 gnd.n1636 0.573776
R12579 gnd.n1636 gnd.n1634 0.573776
R12580 gnd.n1634 gnd.n1632 0.573776
R12581 gnd.n1606 gnd.n1605 0.573776
R12582 gnd.n1605 gnd.n1603 0.573776
R12583 gnd.n1603 gnd.n1601 0.573776
R12584 gnd.n1601 gnd.n1599 0.573776
R12585 gnd.n1599 gnd.n1597 0.573776
R12586 gnd.n1617 gnd.n1616 0.573776
R12587 gnd.n1616 gnd.n1614 0.573776
R12588 gnd.n1614 gnd.n1612 0.573776
R12589 gnd.n1612 gnd.n1610 0.573776
R12590 gnd.n1610 gnd.n1608 0.573776
R12591 gnd.n1629 gnd.n1628 0.573776
R12592 gnd.n1628 gnd.n1626 0.573776
R12593 gnd.n1626 gnd.n1624 0.573776
R12594 gnd.n1624 gnd.n1622 0.573776
R12595 gnd.n1622 gnd.n1620 0.573776
R12596 gnd.n58 gnd.n56 0.573776
R12597 gnd.n60 gnd.n58 0.573776
R12598 gnd.n62 gnd.n60 0.573776
R12599 gnd.n64 gnd.n62 0.573776
R12600 gnd.n65 gnd.n64 0.573776
R12601 gnd.n23 gnd.n21 0.573776
R12602 gnd.n25 gnd.n23 0.573776
R12603 gnd.n27 gnd.n25 0.573776
R12604 gnd.n29 gnd.n27 0.573776
R12605 gnd.n30 gnd.n29 0.573776
R12606 gnd.n34 gnd.n32 0.573776
R12607 gnd.n36 gnd.n34 0.573776
R12608 gnd.n38 gnd.n36 0.573776
R12609 gnd.n40 gnd.n38 0.573776
R12610 gnd.n41 gnd.n40 0.573776
R12611 gnd.n46 gnd.n44 0.573776
R12612 gnd.n48 gnd.n46 0.573776
R12613 gnd.n50 gnd.n48 0.573776
R12614 gnd.n52 gnd.n50 0.573776
R12615 gnd.n53 gnd.n52 0.573776
R12616 gnd.n7327 gnd.n7326 0.532512
R12617 gnd.n4152 gnd.n4151 0.532512
R12618 gnd.n237 gnd.n166 0.497451
R12619 gnd.n2785 gnd.n2630 0.497451
R12620 gnd.n3284 gnd.n3203 0.497451
R12621 gnd.n2458 gnd.n2384 0.497451
R12622 gnd.n2338 gnd.n2337 0.486781
R12623 gnd.n1506 gnd.n1402 0.48678
R12624 gnd.n6285 gnd.n6284 0.480683
R12625 gnd.n1687 gnd.n1353 0.480683
R12626 gnd.n7420 gnd.n7419 0.4705
R12627 gnd.n3418 gnd.n3085 0.451719
R12628 gnd.n3927 gnd.n2644 0.451719
R12629 gnd.n3933 gnd.n2667 0.451719
R12630 gnd.n5714 gnd.n5713 0.451719
R12631 gnd.n6547 gnd.n808 0.425805
R12632 gnd.n7000 gnd.n6999 0.425805
R12633 gnd.n7211 gnd.n410 0.425805
R12634 gnd.n4071 gnd.n4070 0.425805
R12635 gnd.n7408 gnd.n83 0.4255
R12636 gnd.n6099 gnd.n2544 0.4255
R12637 gnd.n5973 gnd.n2728 0.388379
R12638 gnd.n2296 gnd.n2295 0.388379
R12639 gnd.n2264 gnd.n2263 0.388379
R12640 gnd.n2232 gnd.n2231 0.388379
R12641 gnd.n2201 gnd.n2200 0.388379
R12642 gnd.n2169 gnd.n2168 0.388379
R12643 gnd.n2137 gnd.n2136 0.388379
R12644 gnd.n2105 gnd.n2104 0.388379
R12645 gnd.n2074 gnd.n2073 0.388379
R12646 gnd.n5658 gnd.n3151 0.388379
R12647 gnd.n7420 gnd.n19 0.374463
R12648 gnd gnd.n7420 0.367492
R12649 gnd.n1998 gnd.t186 0.319156
R12650 gnd.n6134 gnd.n2489 0.319156
R12651 gnd.n6104 gnd.t233 0.319156
R12652 gnd.t254 gnd.n4289 0.319156
R12653 gnd.n4626 gnd.t331 0.319156
R12654 gnd.n4843 gnd.t178 0.319156
R12655 gnd.n5415 gnd.t211 0.319156
R12656 gnd.t237 gnd.n5442 0.319156
R12657 gnd.n7340 gnd.n134 0.319156
R12658 gnd.n1500 gnd.n1499 0.311721
R12659 gnd.n6037 gnd.n6036 0.302329
R12660 gnd.n5304 gnd.n5303 0.302329
R12661 gnd.n7279 gnd.n386 0.293183
R12662 gnd.n6157 gnd.n2448 0.293183
R12663 gnd.n6330 gnd.n1048 0.268793
R12664 gnd.n386 gnd.n385 0.258122
R12665 gnd.n5534 gnd.n3104 0.258122
R12666 gnd.n2846 gnd.n2638 0.258122
R12667 gnd.n6158 gnd.n6157 0.258122
R12668 gnd.n1088 gnd.n1048 0.241354
R12669 gnd.n3233 gnd.n3230 0.229039
R12670 gnd.n3234 gnd.n3233 0.229039
R12671 gnd.n2911 gnd.n2812 0.229039
R12672 gnd.n2911 gnd.n2910 0.229039
R12673 gnd.n1742 gnd.n1370 0.206293
R12674 gnd.n2313 gnd.n2285 0.155672
R12675 gnd.n2306 gnd.n2285 0.155672
R12676 gnd.n2306 gnd.n2305 0.155672
R12677 gnd.n2305 gnd.n2289 0.155672
R12678 gnd.n2298 gnd.n2289 0.155672
R12679 gnd.n2298 gnd.n2297 0.155672
R12680 gnd.n2281 gnd.n2253 0.155672
R12681 gnd.n2274 gnd.n2253 0.155672
R12682 gnd.n2274 gnd.n2273 0.155672
R12683 gnd.n2273 gnd.n2257 0.155672
R12684 gnd.n2266 gnd.n2257 0.155672
R12685 gnd.n2266 gnd.n2265 0.155672
R12686 gnd.n2249 gnd.n2221 0.155672
R12687 gnd.n2242 gnd.n2221 0.155672
R12688 gnd.n2242 gnd.n2241 0.155672
R12689 gnd.n2241 gnd.n2225 0.155672
R12690 gnd.n2234 gnd.n2225 0.155672
R12691 gnd.n2234 gnd.n2233 0.155672
R12692 gnd.n2218 gnd.n2190 0.155672
R12693 gnd.n2211 gnd.n2190 0.155672
R12694 gnd.n2211 gnd.n2210 0.155672
R12695 gnd.n2210 gnd.n2194 0.155672
R12696 gnd.n2203 gnd.n2194 0.155672
R12697 gnd.n2203 gnd.n2202 0.155672
R12698 gnd.n2186 gnd.n2158 0.155672
R12699 gnd.n2179 gnd.n2158 0.155672
R12700 gnd.n2179 gnd.n2178 0.155672
R12701 gnd.n2178 gnd.n2162 0.155672
R12702 gnd.n2171 gnd.n2162 0.155672
R12703 gnd.n2171 gnd.n2170 0.155672
R12704 gnd.n2154 gnd.n2126 0.155672
R12705 gnd.n2147 gnd.n2126 0.155672
R12706 gnd.n2147 gnd.n2146 0.155672
R12707 gnd.n2146 gnd.n2130 0.155672
R12708 gnd.n2139 gnd.n2130 0.155672
R12709 gnd.n2139 gnd.n2138 0.155672
R12710 gnd.n2122 gnd.n2094 0.155672
R12711 gnd.n2115 gnd.n2094 0.155672
R12712 gnd.n2115 gnd.n2114 0.155672
R12713 gnd.n2114 gnd.n2098 0.155672
R12714 gnd.n2107 gnd.n2098 0.155672
R12715 gnd.n2107 gnd.n2106 0.155672
R12716 gnd.n2091 gnd.n2063 0.155672
R12717 gnd.n2084 gnd.n2063 0.155672
R12718 gnd.n2084 gnd.n2083 0.155672
R12719 gnd.n2083 gnd.n2067 0.155672
R12720 gnd.n2076 gnd.n2067 0.155672
R12721 gnd.n2076 gnd.n2075 0.155672
R12722 gnd.n6319 gnd.n6285 0.152939
R12723 gnd.n6319 gnd.n6318 0.152939
R12724 gnd.n6318 gnd.n6317 0.152939
R12725 gnd.n6317 gnd.n6287 0.152939
R12726 gnd.n6288 gnd.n6287 0.152939
R12727 gnd.n6289 gnd.n6288 0.152939
R12728 gnd.n6290 gnd.n6289 0.152939
R12729 gnd.n6291 gnd.n6290 0.152939
R12730 gnd.n6292 gnd.n6291 0.152939
R12731 gnd.n6293 gnd.n6292 0.152939
R12732 gnd.n6294 gnd.n6293 0.152939
R12733 gnd.n6295 gnd.n6294 0.152939
R12734 gnd.n6295 gnd.n1054 0.152939
R12735 gnd.n6328 gnd.n1054 0.152939
R12736 gnd.n6329 gnd.n6328 0.152939
R12737 gnd.n6330 gnd.n6329 0.152939
R12738 gnd.n1762 gnd.n1353 0.152939
R12739 gnd.n1763 gnd.n1762 0.152939
R12740 gnd.n1764 gnd.n1763 0.152939
R12741 gnd.n1765 gnd.n1764 0.152939
R12742 gnd.n1765 gnd.n1328 0.152939
R12743 gnd.n1793 gnd.n1328 0.152939
R12744 gnd.n1794 gnd.n1793 0.152939
R12745 gnd.n1795 gnd.n1794 0.152939
R12746 gnd.n1796 gnd.n1795 0.152939
R12747 gnd.n1796 gnd.n1302 0.152939
R12748 gnd.n1824 gnd.n1302 0.152939
R12749 gnd.n1825 gnd.n1824 0.152939
R12750 gnd.n1826 gnd.n1825 0.152939
R12751 gnd.n1827 gnd.n1826 0.152939
R12752 gnd.n1827 gnd.n1276 0.152939
R12753 gnd.n1855 gnd.n1276 0.152939
R12754 gnd.n1856 gnd.n1855 0.152939
R12755 gnd.n1857 gnd.n1856 0.152939
R12756 gnd.n1858 gnd.n1857 0.152939
R12757 gnd.n1858 gnd.n1250 0.152939
R12758 gnd.n1886 gnd.n1250 0.152939
R12759 gnd.n1887 gnd.n1886 0.152939
R12760 gnd.n1888 gnd.n1887 0.152939
R12761 gnd.n1889 gnd.n1888 0.152939
R12762 gnd.n1889 gnd.n1225 0.152939
R12763 gnd.n1917 gnd.n1225 0.152939
R12764 gnd.n1918 gnd.n1917 0.152939
R12765 gnd.n1919 gnd.n1918 0.152939
R12766 gnd.n1920 gnd.n1919 0.152939
R12767 gnd.n1920 gnd.n1198 0.152939
R12768 gnd.n1947 gnd.n1198 0.152939
R12769 gnd.n1948 gnd.n1947 0.152939
R12770 gnd.n1949 gnd.n1948 0.152939
R12771 gnd.n1949 gnd.n1176 0.152939
R12772 gnd.n2017 gnd.n1176 0.152939
R12773 gnd.n2018 gnd.n2017 0.152939
R12774 gnd.n2019 gnd.n2018 0.152939
R12775 gnd.n2021 gnd.n2019 0.152939
R12776 gnd.n2021 gnd.n2020 0.152939
R12777 gnd.n2020 gnd.n984 0.152939
R12778 gnd.n985 gnd.n984 0.152939
R12779 gnd.n986 gnd.n985 0.152939
R12780 gnd.n1008 gnd.n986 0.152939
R12781 gnd.n1009 gnd.n1008 0.152939
R12782 gnd.n1010 gnd.n1009 0.152939
R12783 gnd.n1011 gnd.n1010 0.152939
R12784 gnd.n1012 gnd.n1011 0.152939
R12785 gnd.n1033 gnd.n1012 0.152939
R12786 gnd.n1034 gnd.n1033 0.152939
R12787 gnd.n1035 gnd.n1034 0.152939
R12788 gnd.n1036 gnd.n1035 0.152939
R12789 gnd.n1037 gnd.n1036 0.152939
R12790 gnd.n6284 gnd.n1037 0.152939
R12791 gnd.n1688 gnd.n1687 0.152939
R12792 gnd.n1689 gnd.n1688 0.152939
R12793 gnd.n1690 gnd.n1689 0.152939
R12794 gnd.n1691 gnd.n1690 0.152939
R12795 gnd.n1692 gnd.n1691 0.152939
R12796 gnd.n1693 gnd.n1692 0.152939
R12797 gnd.n1694 gnd.n1693 0.152939
R12798 gnd.n1695 gnd.n1694 0.152939
R12799 gnd.n1696 gnd.n1695 0.152939
R12800 gnd.n1697 gnd.n1696 0.152939
R12801 gnd.n1698 gnd.n1697 0.152939
R12802 gnd.n1699 gnd.n1698 0.152939
R12803 gnd.n1700 gnd.n1699 0.152939
R12804 gnd.n1701 gnd.n1700 0.152939
R12805 gnd.n1705 gnd.n1701 0.152939
R12806 gnd.n1705 gnd.n1370 0.152939
R12807 gnd.n1089 gnd.n1088 0.152939
R12808 gnd.n1090 gnd.n1089 0.152939
R12809 gnd.n1090 gnd.n1084 0.152939
R12810 gnd.n1098 gnd.n1084 0.152939
R12811 gnd.n1099 gnd.n1098 0.152939
R12812 gnd.n1100 gnd.n1099 0.152939
R12813 gnd.n1100 gnd.n1082 0.152939
R12814 gnd.n1108 gnd.n1082 0.152939
R12815 gnd.n1109 gnd.n1108 0.152939
R12816 gnd.n1110 gnd.n1109 0.152939
R12817 gnd.n1110 gnd.n1080 0.152939
R12818 gnd.n1118 gnd.n1080 0.152939
R12819 gnd.n1119 gnd.n1118 0.152939
R12820 gnd.n1120 gnd.n1119 0.152939
R12821 gnd.n1120 gnd.n1078 0.152939
R12822 gnd.n1128 gnd.n1078 0.152939
R12823 gnd.n1129 gnd.n1128 0.152939
R12824 gnd.n1130 gnd.n1129 0.152939
R12825 gnd.n1130 gnd.n1076 0.152939
R12826 gnd.n1138 gnd.n1076 0.152939
R12827 gnd.n1139 gnd.n1138 0.152939
R12828 gnd.n1140 gnd.n1139 0.152939
R12829 gnd.n1140 gnd.n1071 0.152939
R12830 gnd.n1147 gnd.n1071 0.152939
R12831 gnd.n1148 gnd.n1147 0.152939
R12832 gnd.n2338 gnd.n1148 0.152939
R12833 gnd.n1562 gnd.n1560 0.152939
R12834 gnd.n1563 gnd.n1562 0.152939
R12835 gnd.n1564 gnd.n1563 0.152939
R12836 gnd.n1565 gnd.n1564 0.152939
R12837 gnd.n1566 gnd.n1565 0.152939
R12838 gnd.n1567 gnd.n1566 0.152939
R12839 gnd.n1568 gnd.n1567 0.152939
R12840 gnd.n1568 gnd.n1183 0.152939
R12841 gnd.n1969 gnd.n1183 0.152939
R12842 gnd.n1970 gnd.n1969 0.152939
R12843 gnd.n1971 gnd.n1970 0.152939
R12844 gnd.n1972 gnd.n1971 0.152939
R12845 gnd.n1973 gnd.n1972 0.152939
R12846 gnd.n1974 gnd.n1973 0.152939
R12847 gnd.n1975 gnd.n1974 0.152939
R12848 gnd.n1977 gnd.n1975 0.152939
R12849 gnd.n1978 gnd.n1977 0.152939
R12850 gnd.n1979 gnd.n1978 0.152939
R12851 gnd.n1980 gnd.n1979 0.152939
R12852 gnd.n1981 gnd.n1980 0.152939
R12853 gnd.n1982 gnd.n1981 0.152939
R12854 gnd.n1983 gnd.n1982 0.152939
R12855 gnd.n1984 gnd.n1983 0.152939
R12856 gnd.n1985 gnd.n1984 0.152939
R12857 gnd.n1987 gnd.n1985 0.152939
R12858 gnd.n1987 gnd.n1986 0.152939
R12859 gnd.n1986 gnd.n1149 0.152939
R12860 gnd.n2337 gnd.n1149 0.152939
R12861 gnd.n1507 gnd.n1506 0.152939
R12862 gnd.n1508 gnd.n1507 0.152939
R12863 gnd.n1508 gnd.n1390 0.152939
R12864 gnd.n1522 gnd.n1390 0.152939
R12865 gnd.n1523 gnd.n1522 0.152939
R12866 gnd.n1524 gnd.n1523 0.152939
R12867 gnd.n1524 gnd.n1377 0.152939
R12868 gnd.n1538 gnd.n1377 0.152939
R12869 gnd.n1539 gnd.n1538 0.152939
R12870 gnd.n1540 gnd.n1539 0.152939
R12871 gnd.n1541 gnd.n1540 0.152939
R12872 gnd.n1542 gnd.n1541 0.152939
R12873 gnd.n1543 gnd.n1542 0.152939
R12874 gnd.n1544 gnd.n1543 0.152939
R12875 gnd.n1545 gnd.n1544 0.152939
R12876 gnd.n1546 gnd.n1545 0.152939
R12877 gnd.n1547 gnd.n1546 0.152939
R12878 gnd.n1548 gnd.n1547 0.152939
R12879 gnd.n1549 gnd.n1548 0.152939
R12880 gnd.n1550 gnd.n1549 0.152939
R12881 gnd.n1551 gnd.n1550 0.152939
R12882 gnd.n1552 gnd.n1551 0.152939
R12883 gnd.n1553 gnd.n1552 0.152939
R12884 gnd.n1554 gnd.n1553 0.152939
R12885 gnd.n1555 gnd.n1554 0.152939
R12886 gnd.n1556 gnd.n1555 0.152939
R12887 gnd.n1557 gnd.n1556 0.152939
R12888 gnd.n1558 gnd.n1557 0.152939
R12889 gnd.n1499 gnd.n1406 0.152939
R12890 gnd.n1409 gnd.n1406 0.152939
R12891 gnd.n1410 gnd.n1409 0.152939
R12892 gnd.n1411 gnd.n1410 0.152939
R12893 gnd.n1414 gnd.n1411 0.152939
R12894 gnd.n1415 gnd.n1414 0.152939
R12895 gnd.n1416 gnd.n1415 0.152939
R12896 gnd.n1417 gnd.n1416 0.152939
R12897 gnd.n1420 gnd.n1417 0.152939
R12898 gnd.n1421 gnd.n1420 0.152939
R12899 gnd.n1422 gnd.n1421 0.152939
R12900 gnd.n1423 gnd.n1422 0.152939
R12901 gnd.n1426 gnd.n1423 0.152939
R12902 gnd.n1427 gnd.n1426 0.152939
R12903 gnd.n1428 gnd.n1427 0.152939
R12904 gnd.n1429 gnd.n1428 0.152939
R12905 gnd.n1432 gnd.n1429 0.152939
R12906 gnd.n1433 gnd.n1432 0.152939
R12907 gnd.n1434 gnd.n1433 0.152939
R12908 gnd.n1435 gnd.n1434 0.152939
R12909 gnd.n1438 gnd.n1435 0.152939
R12910 gnd.n1439 gnd.n1438 0.152939
R12911 gnd.n1442 gnd.n1439 0.152939
R12912 gnd.n1443 gnd.n1442 0.152939
R12913 gnd.n1445 gnd.n1443 0.152939
R12914 gnd.n1445 gnd.n1402 0.152939
R12915 gnd.n6548 gnd.n6547 0.152939
R12916 gnd.n6549 gnd.n6548 0.152939
R12917 gnd.n6549 gnd.n802 0.152939
R12918 gnd.n6557 gnd.n802 0.152939
R12919 gnd.n6558 gnd.n6557 0.152939
R12920 gnd.n6559 gnd.n6558 0.152939
R12921 gnd.n6559 gnd.n796 0.152939
R12922 gnd.n6567 gnd.n796 0.152939
R12923 gnd.n6568 gnd.n6567 0.152939
R12924 gnd.n6569 gnd.n6568 0.152939
R12925 gnd.n6569 gnd.n790 0.152939
R12926 gnd.n6577 gnd.n790 0.152939
R12927 gnd.n6578 gnd.n6577 0.152939
R12928 gnd.n6579 gnd.n6578 0.152939
R12929 gnd.n6579 gnd.n784 0.152939
R12930 gnd.n6587 gnd.n784 0.152939
R12931 gnd.n6588 gnd.n6587 0.152939
R12932 gnd.n6589 gnd.n6588 0.152939
R12933 gnd.n6589 gnd.n778 0.152939
R12934 gnd.n6597 gnd.n778 0.152939
R12935 gnd.n6598 gnd.n6597 0.152939
R12936 gnd.n6599 gnd.n6598 0.152939
R12937 gnd.n6599 gnd.n772 0.152939
R12938 gnd.n6607 gnd.n772 0.152939
R12939 gnd.n6608 gnd.n6607 0.152939
R12940 gnd.n6609 gnd.n6608 0.152939
R12941 gnd.n6609 gnd.n766 0.152939
R12942 gnd.n6617 gnd.n766 0.152939
R12943 gnd.n6618 gnd.n6617 0.152939
R12944 gnd.n6619 gnd.n6618 0.152939
R12945 gnd.n6619 gnd.n760 0.152939
R12946 gnd.n6627 gnd.n760 0.152939
R12947 gnd.n6628 gnd.n6627 0.152939
R12948 gnd.n6629 gnd.n6628 0.152939
R12949 gnd.n6629 gnd.n754 0.152939
R12950 gnd.n6637 gnd.n754 0.152939
R12951 gnd.n6638 gnd.n6637 0.152939
R12952 gnd.n6639 gnd.n6638 0.152939
R12953 gnd.n6639 gnd.n748 0.152939
R12954 gnd.n6647 gnd.n748 0.152939
R12955 gnd.n6648 gnd.n6647 0.152939
R12956 gnd.n6649 gnd.n6648 0.152939
R12957 gnd.n6649 gnd.n742 0.152939
R12958 gnd.n6657 gnd.n742 0.152939
R12959 gnd.n6658 gnd.n6657 0.152939
R12960 gnd.n6659 gnd.n6658 0.152939
R12961 gnd.n6659 gnd.n736 0.152939
R12962 gnd.n6667 gnd.n736 0.152939
R12963 gnd.n6668 gnd.n6667 0.152939
R12964 gnd.n6669 gnd.n6668 0.152939
R12965 gnd.n6669 gnd.n730 0.152939
R12966 gnd.n6677 gnd.n730 0.152939
R12967 gnd.n6678 gnd.n6677 0.152939
R12968 gnd.n6679 gnd.n6678 0.152939
R12969 gnd.n6679 gnd.n724 0.152939
R12970 gnd.n6687 gnd.n724 0.152939
R12971 gnd.n6688 gnd.n6687 0.152939
R12972 gnd.n6689 gnd.n6688 0.152939
R12973 gnd.n6689 gnd.n718 0.152939
R12974 gnd.n6697 gnd.n718 0.152939
R12975 gnd.n6698 gnd.n6697 0.152939
R12976 gnd.n6699 gnd.n6698 0.152939
R12977 gnd.n6699 gnd.n712 0.152939
R12978 gnd.n6707 gnd.n712 0.152939
R12979 gnd.n6708 gnd.n6707 0.152939
R12980 gnd.n6709 gnd.n6708 0.152939
R12981 gnd.n6709 gnd.n706 0.152939
R12982 gnd.n6717 gnd.n706 0.152939
R12983 gnd.n6718 gnd.n6717 0.152939
R12984 gnd.n6719 gnd.n6718 0.152939
R12985 gnd.n6719 gnd.n700 0.152939
R12986 gnd.n6727 gnd.n700 0.152939
R12987 gnd.n6728 gnd.n6727 0.152939
R12988 gnd.n6729 gnd.n6728 0.152939
R12989 gnd.n6729 gnd.n694 0.152939
R12990 gnd.n6737 gnd.n694 0.152939
R12991 gnd.n6738 gnd.n6737 0.152939
R12992 gnd.n6739 gnd.n6738 0.152939
R12993 gnd.n6739 gnd.n688 0.152939
R12994 gnd.n6747 gnd.n688 0.152939
R12995 gnd.n6748 gnd.n6747 0.152939
R12996 gnd.n6749 gnd.n6748 0.152939
R12997 gnd.n6749 gnd.n682 0.152939
R12998 gnd.n6757 gnd.n682 0.152939
R12999 gnd.n6758 gnd.n6757 0.152939
R13000 gnd.n6759 gnd.n6758 0.152939
R13001 gnd.n6759 gnd.n676 0.152939
R13002 gnd.n6767 gnd.n676 0.152939
R13003 gnd.n6768 gnd.n6767 0.152939
R13004 gnd.n6769 gnd.n6768 0.152939
R13005 gnd.n6769 gnd.n670 0.152939
R13006 gnd.n6777 gnd.n670 0.152939
R13007 gnd.n6778 gnd.n6777 0.152939
R13008 gnd.n6779 gnd.n6778 0.152939
R13009 gnd.n6779 gnd.n664 0.152939
R13010 gnd.n6787 gnd.n664 0.152939
R13011 gnd.n6788 gnd.n6787 0.152939
R13012 gnd.n6789 gnd.n6788 0.152939
R13013 gnd.n6789 gnd.n658 0.152939
R13014 gnd.n6797 gnd.n658 0.152939
R13015 gnd.n6798 gnd.n6797 0.152939
R13016 gnd.n6799 gnd.n6798 0.152939
R13017 gnd.n6799 gnd.n652 0.152939
R13018 gnd.n6807 gnd.n652 0.152939
R13019 gnd.n6808 gnd.n6807 0.152939
R13020 gnd.n6809 gnd.n6808 0.152939
R13021 gnd.n6809 gnd.n646 0.152939
R13022 gnd.n6817 gnd.n646 0.152939
R13023 gnd.n6818 gnd.n6817 0.152939
R13024 gnd.n6819 gnd.n6818 0.152939
R13025 gnd.n6819 gnd.n640 0.152939
R13026 gnd.n6827 gnd.n640 0.152939
R13027 gnd.n6828 gnd.n6827 0.152939
R13028 gnd.n6829 gnd.n6828 0.152939
R13029 gnd.n6829 gnd.n634 0.152939
R13030 gnd.n6837 gnd.n634 0.152939
R13031 gnd.n6838 gnd.n6837 0.152939
R13032 gnd.n6839 gnd.n6838 0.152939
R13033 gnd.n6839 gnd.n628 0.152939
R13034 gnd.n6847 gnd.n628 0.152939
R13035 gnd.n6848 gnd.n6847 0.152939
R13036 gnd.n6849 gnd.n6848 0.152939
R13037 gnd.n6849 gnd.n622 0.152939
R13038 gnd.n6857 gnd.n622 0.152939
R13039 gnd.n6858 gnd.n6857 0.152939
R13040 gnd.n6859 gnd.n6858 0.152939
R13041 gnd.n6859 gnd.n616 0.152939
R13042 gnd.n6867 gnd.n616 0.152939
R13043 gnd.n6868 gnd.n6867 0.152939
R13044 gnd.n6869 gnd.n6868 0.152939
R13045 gnd.n6869 gnd.n610 0.152939
R13046 gnd.n6877 gnd.n610 0.152939
R13047 gnd.n6878 gnd.n6877 0.152939
R13048 gnd.n6879 gnd.n6878 0.152939
R13049 gnd.n6879 gnd.n604 0.152939
R13050 gnd.n6887 gnd.n604 0.152939
R13051 gnd.n6888 gnd.n6887 0.152939
R13052 gnd.n6889 gnd.n6888 0.152939
R13053 gnd.n6889 gnd.n598 0.152939
R13054 gnd.n6897 gnd.n598 0.152939
R13055 gnd.n6898 gnd.n6897 0.152939
R13056 gnd.n6899 gnd.n6898 0.152939
R13057 gnd.n6899 gnd.n592 0.152939
R13058 gnd.n6907 gnd.n592 0.152939
R13059 gnd.n6908 gnd.n6907 0.152939
R13060 gnd.n6909 gnd.n6908 0.152939
R13061 gnd.n6909 gnd.n586 0.152939
R13062 gnd.n6917 gnd.n586 0.152939
R13063 gnd.n6918 gnd.n6917 0.152939
R13064 gnd.n6919 gnd.n6918 0.152939
R13065 gnd.n6919 gnd.n580 0.152939
R13066 gnd.n6927 gnd.n580 0.152939
R13067 gnd.n6928 gnd.n6927 0.152939
R13068 gnd.n6929 gnd.n6928 0.152939
R13069 gnd.n6929 gnd.n574 0.152939
R13070 gnd.n6937 gnd.n574 0.152939
R13071 gnd.n6938 gnd.n6937 0.152939
R13072 gnd.n6939 gnd.n6938 0.152939
R13073 gnd.n6939 gnd.n568 0.152939
R13074 gnd.n6947 gnd.n568 0.152939
R13075 gnd.n6948 gnd.n6947 0.152939
R13076 gnd.n6949 gnd.n6948 0.152939
R13077 gnd.n6949 gnd.n562 0.152939
R13078 gnd.n6957 gnd.n562 0.152939
R13079 gnd.n6958 gnd.n6957 0.152939
R13080 gnd.n6959 gnd.n6958 0.152939
R13081 gnd.n6959 gnd.n556 0.152939
R13082 gnd.n6967 gnd.n556 0.152939
R13083 gnd.n6968 gnd.n6967 0.152939
R13084 gnd.n6969 gnd.n6968 0.152939
R13085 gnd.n6969 gnd.n550 0.152939
R13086 gnd.n6977 gnd.n550 0.152939
R13087 gnd.n6978 gnd.n6977 0.152939
R13088 gnd.n6979 gnd.n6978 0.152939
R13089 gnd.n6979 gnd.n544 0.152939
R13090 gnd.n6987 gnd.n544 0.152939
R13091 gnd.n6988 gnd.n6987 0.152939
R13092 gnd.n6990 gnd.n6988 0.152939
R13093 gnd.n6990 gnd.n6989 0.152939
R13094 gnd.n6989 gnd.n538 0.152939
R13095 gnd.n6999 gnd.n538 0.152939
R13096 gnd.n7000 gnd.n533 0.152939
R13097 gnd.n7008 gnd.n533 0.152939
R13098 gnd.n7009 gnd.n7008 0.152939
R13099 gnd.n7010 gnd.n7009 0.152939
R13100 gnd.n7010 gnd.n527 0.152939
R13101 gnd.n7018 gnd.n527 0.152939
R13102 gnd.n7019 gnd.n7018 0.152939
R13103 gnd.n7020 gnd.n7019 0.152939
R13104 gnd.n7020 gnd.n521 0.152939
R13105 gnd.n7028 gnd.n521 0.152939
R13106 gnd.n7029 gnd.n7028 0.152939
R13107 gnd.n7030 gnd.n7029 0.152939
R13108 gnd.n7030 gnd.n515 0.152939
R13109 gnd.n7038 gnd.n515 0.152939
R13110 gnd.n7039 gnd.n7038 0.152939
R13111 gnd.n7040 gnd.n7039 0.152939
R13112 gnd.n7040 gnd.n509 0.152939
R13113 gnd.n7048 gnd.n509 0.152939
R13114 gnd.n7049 gnd.n7048 0.152939
R13115 gnd.n7050 gnd.n7049 0.152939
R13116 gnd.n7050 gnd.n503 0.152939
R13117 gnd.n7058 gnd.n503 0.152939
R13118 gnd.n7059 gnd.n7058 0.152939
R13119 gnd.n7060 gnd.n7059 0.152939
R13120 gnd.n7060 gnd.n497 0.152939
R13121 gnd.n7068 gnd.n497 0.152939
R13122 gnd.n7069 gnd.n7068 0.152939
R13123 gnd.n7070 gnd.n7069 0.152939
R13124 gnd.n7070 gnd.n491 0.152939
R13125 gnd.n7078 gnd.n491 0.152939
R13126 gnd.n7079 gnd.n7078 0.152939
R13127 gnd.n7080 gnd.n7079 0.152939
R13128 gnd.n7080 gnd.n485 0.152939
R13129 gnd.n7088 gnd.n485 0.152939
R13130 gnd.n7089 gnd.n7088 0.152939
R13131 gnd.n7090 gnd.n7089 0.152939
R13132 gnd.n7090 gnd.n479 0.152939
R13133 gnd.n7098 gnd.n479 0.152939
R13134 gnd.n7099 gnd.n7098 0.152939
R13135 gnd.n7100 gnd.n7099 0.152939
R13136 gnd.n7100 gnd.n473 0.152939
R13137 gnd.n7108 gnd.n473 0.152939
R13138 gnd.n7109 gnd.n7108 0.152939
R13139 gnd.n7110 gnd.n7109 0.152939
R13140 gnd.n7110 gnd.n467 0.152939
R13141 gnd.n7118 gnd.n467 0.152939
R13142 gnd.n7119 gnd.n7118 0.152939
R13143 gnd.n7120 gnd.n7119 0.152939
R13144 gnd.n7120 gnd.n461 0.152939
R13145 gnd.n7128 gnd.n461 0.152939
R13146 gnd.n7129 gnd.n7128 0.152939
R13147 gnd.n7130 gnd.n7129 0.152939
R13148 gnd.n7130 gnd.n455 0.152939
R13149 gnd.n7138 gnd.n455 0.152939
R13150 gnd.n7139 gnd.n7138 0.152939
R13151 gnd.n7140 gnd.n7139 0.152939
R13152 gnd.n7140 gnd.n449 0.152939
R13153 gnd.n7148 gnd.n449 0.152939
R13154 gnd.n7149 gnd.n7148 0.152939
R13155 gnd.n7150 gnd.n7149 0.152939
R13156 gnd.n7150 gnd.n443 0.152939
R13157 gnd.n7158 gnd.n443 0.152939
R13158 gnd.n7159 gnd.n7158 0.152939
R13159 gnd.n7160 gnd.n7159 0.152939
R13160 gnd.n7160 gnd.n437 0.152939
R13161 gnd.n7168 gnd.n437 0.152939
R13162 gnd.n7169 gnd.n7168 0.152939
R13163 gnd.n7170 gnd.n7169 0.152939
R13164 gnd.n7170 gnd.n431 0.152939
R13165 gnd.n7178 gnd.n431 0.152939
R13166 gnd.n7179 gnd.n7178 0.152939
R13167 gnd.n7180 gnd.n7179 0.152939
R13168 gnd.n7180 gnd.n425 0.152939
R13169 gnd.n7188 gnd.n425 0.152939
R13170 gnd.n7189 gnd.n7188 0.152939
R13171 gnd.n7190 gnd.n7189 0.152939
R13172 gnd.n7190 gnd.n419 0.152939
R13173 gnd.n7198 gnd.n419 0.152939
R13174 gnd.n7199 gnd.n7198 0.152939
R13175 gnd.n7200 gnd.n7199 0.152939
R13176 gnd.n7200 gnd.n413 0.152939
R13177 gnd.n7209 gnd.n413 0.152939
R13178 gnd.n7210 gnd.n7209 0.152939
R13179 gnd.n7211 gnd.n7210 0.152939
R13180 gnd.n402 gnd.n401 0.152939
R13181 gnd.n403 gnd.n402 0.152939
R13182 gnd.n404 gnd.n403 0.152939
R13183 gnd.n407 gnd.n404 0.152939
R13184 gnd.n408 gnd.n407 0.152939
R13185 gnd.n409 gnd.n408 0.152939
R13186 gnd.n410 gnd.n409 0.152939
R13187 gnd.n7408 gnd.n81 0.152939
R13188 gnd.n106 gnd.n81 0.152939
R13189 gnd.n107 gnd.n106 0.152939
R13190 gnd.n108 gnd.n107 0.152939
R13191 gnd.n125 gnd.n108 0.152939
R13192 gnd.n126 gnd.n125 0.152939
R13193 gnd.n127 gnd.n126 0.152939
R13194 gnd.n128 gnd.n127 0.152939
R13195 gnd.n145 gnd.n128 0.152939
R13196 gnd.n146 gnd.n145 0.152939
R13197 gnd.n147 gnd.n146 0.152939
R13198 gnd.n148 gnd.n147 0.152939
R13199 gnd.n163 gnd.n148 0.152939
R13200 gnd.n164 gnd.n163 0.152939
R13201 gnd.n165 gnd.n164 0.152939
R13202 gnd.n166 gnd.n165 0.152939
R13203 gnd.n7417 gnd.n69 0.152939
R13204 gnd.n5434 gnd.n69 0.152939
R13205 gnd.n5435 gnd.n5434 0.152939
R13206 gnd.n5436 gnd.n5435 0.152939
R13207 gnd.n5437 gnd.n5436 0.152939
R13208 gnd.n5437 gnd.n394 0.152939
R13209 gnd.n7236 gnd.n394 0.152939
R13210 gnd.n7237 gnd.n7236 0.152939
R13211 gnd.n7238 gnd.n7237 0.152939
R13212 gnd.n7238 gnd.n389 0.152939
R13213 gnd.n7251 gnd.n389 0.152939
R13214 gnd.n7252 gnd.n7251 0.152939
R13215 gnd.n7253 gnd.n7252 0.152939
R13216 gnd.n7254 gnd.n7253 0.152939
R13217 gnd.n7255 gnd.n7254 0.152939
R13218 gnd.n7256 gnd.n7255 0.152939
R13219 gnd.n7257 gnd.n7256 0.152939
R13220 gnd.n7258 gnd.n7257 0.152939
R13221 gnd.n7259 gnd.n7258 0.152939
R13222 gnd.n7327 gnd.n7259 0.152939
R13223 gnd.n7279 gnd.n7278 0.152939
R13224 gnd.n7287 gnd.n7278 0.152939
R13225 gnd.n7288 gnd.n7287 0.152939
R13226 gnd.n7289 gnd.n7288 0.152939
R13227 gnd.n7289 gnd.n7274 0.152939
R13228 gnd.n7297 gnd.n7274 0.152939
R13229 gnd.n7298 gnd.n7297 0.152939
R13230 gnd.n7299 gnd.n7298 0.152939
R13231 gnd.n7299 gnd.n7270 0.152939
R13232 gnd.n7307 gnd.n7270 0.152939
R13233 gnd.n7308 gnd.n7307 0.152939
R13234 gnd.n7309 gnd.n7308 0.152939
R13235 gnd.n7309 gnd.n7266 0.152939
R13236 gnd.n7317 gnd.n7266 0.152939
R13237 gnd.n7318 gnd.n7317 0.152939
R13238 gnd.n7319 gnd.n7318 0.152939
R13239 gnd.n7319 gnd.n7260 0.152939
R13240 gnd.n7326 gnd.n7260 0.152939
R13241 gnd.n237 gnd.n236 0.152939
R13242 gnd.n245 gnd.n236 0.152939
R13243 gnd.n246 gnd.n245 0.152939
R13244 gnd.n247 gnd.n246 0.152939
R13245 gnd.n247 gnd.n232 0.152939
R13246 gnd.n255 gnd.n232 0.152939
R13247 gnd.n256 gnd.n255 0.152939
R13248 gnd.n257 gnd.n256 0.152939
R13249 gnd.n257 gnd.n228 0.152939
R13250 gnd.n265 gnd.n228 0.152939
R13251 gnd.n266 gnd.n265 0.152939
R13252 gnd.n267 gnd.n266 0.152939
R13253 gnd.n267 gnd.n224 0.152939
R13254 gnd.n276 gnd.n224 0.152939
R13255 gnd.n277 gnd.n276 0.152939
R13256 gnd.n278 gnd.n277 0.152939
R13257 gnd.n278 gnd.n218 0.152939
R13258 gnd.n286 gnd.n218 0.152939
R13259 gnd.n287 gnd.n286 0.152939
R13260 gnd.n288 gnd.n287 0.152939
R13261 gnd.n288 gnd.n214 0.152939
R13262 gnd.n296 gnd.n214 0.152939
R13263 gnd.n297 gnd.n296 0.152939
R13264 gnd.n298 gnd.n297 0.152939
R13265 gnd.n298 gnd.n210 0.152939
R13266 gnd.n306 gnd.n210 0.152939
R13267 gnd.n307 gnd.n306 0.152939
R13268 gnd.n308 gnd.n307 0.152939
R13269 gnd.n308 gnd.n206 0.152939
R13270 gnd.n316 gnd.n206 0.152939
R13271 gnd.n317 gnd.n316 0.152939
R13272 gnd.n318 gnd.n317 0.152939
R13273 gnd.n318 gnd.n202 0.152939
R13274 gnd.n326 gnd.n202 0.152939
R13275 gnd.n327 gnd.n326 0.152939
R13276 gnd.n328 gnd.n327 0.152939
R13277 gnd.n328 gnd.n196 0.152939
R13278 gnd.n336 gnd.n196 0.152939
R13279 gnd.n337 gnd.n336 0.152939
R13280 gnd.n338 gnd.n337 0.152939
R13281 gnd.n338 gnd.n192 0.152939
R13282 gnd.n346 gnd.n192 0.152939
R13283 gnd.n347 gnd.n346 0.152939
R13284 gnd.n348 gnd.n347 0.152939
R13285 gnd.n348 gnd.n188 0.152939
R13286 gnd.n356 gnd.n188 0.152939
R13287 gnd.n357 gnd.n356 0.152939
R13288 gnd.n358 gnd.n357 0.152939
R13289 gnd.n358 gnd.n184 0.152939
R13290 gnd.n366 gnd.n184 0.152939
R13291 gnd.n367 gnd.n366 0.152939
R13292 gnd.n368 gnd.n367 0.152939
R13293 gnd.n368 gnd.n180 0.152939
R13294 gnd.n376 gnd.n180 0.152939
R13295 gnd.n377 gnd.n376 0.152939
R13296 gnd.n378 gnd.n377 0.152939
R13297 gnd.n378 gnd.n174 0.152939
R13298 gnd.n385 gnd.n174 0.152939
R13299 gnd.n3204 gnd.n3203 0.152939
R13300 gnd.n3205 gnd.n3204 0.152939
R13301 gnd.n3206 gnd.n3205 0.152939
R13302 gnd.n3207 gnd.n3206 0.152939
R13303 gnd.n3208 gnd.n3207 0.152939
R13304 gnd.n3209 gnd.n3208 0.152939
R13305 gnd.n3210 gnd.n3209 0.152939
R13306 gnd.n3211 gnd.n3210 0.152939
R13307 gnd.n3212 gnd.n3211 0.152939
R13308 gnd.n3213 gnd.n3212 0.152939
R13309 gnd.n3214 gnd.n3213 0.152939
R13310 gnd.n3215 gnd.n3214 0.152939
R13311 gnd.n3216 gnd.n3215 0.152939
R13312 gnd.n3217 gnd.n3216 0.152939
R13313 gnd.n3218 gnd.n3217 0.152939
R13314 gnd.n3219 gnd.n3218 0.152939
R13315 gnd.n3220 gnd.n3219 0.152939
R13316 gnd.n3223 gnd.n3220 0.152939
R13317 gnd.n3224 gnd.n3223 0.152939
R13318 gnd.n3225 gnd.n3224 0.152939
R13319 gnd.n3226 gnd.n3225 0.152939
R13320 gnd.n3227 gnd.n3226 0.152939
R13321 gnd.n3228 gnd.n3227 0.152939
R13322 gnd.n3229 gnd.n3228 0.152939
R13323 gnd.n3230 gnd.n3229 0.152939
R13324 gnd.n3235 gnd.n3234 0.152939
R13325 gnd.n3236 gnd.n3235 0.152939
R13326 gnd.n3237 gnd.n3236 0.152939
R13327 gnd.n3238 gnd.n3237 0.152939
R13328 gnd.n3239 gnd.n3238 0.152939
R13329 gnd.n3240 gnd.n3239 0.152939
R13330 gnd.n3241 gnd.n3240 0.152939
R13331 gnd.n3242 gnd.n3241 0.152939
R13332 gnd.n3243 gnd.n3242 0.152939
R13333 gnd.n3246 gnd.n3243 0.152939
R13334 gnd.n3247 gnd.n3246 0.152939
R13335 gnd.n3248 gnd.n3247 0.152939
R13336 gnd.n3249 gnd.n3248 0.152939
R13337 gnd.n3250 gnd.n3249 0.152939
R13338 gnd.n3251 gnd.n3250 0.152939
R13339 gnd.n3252 gnd.n3251 0.152939
R13340 gnd.n3253 gnd.n3252 0.152939
R13341 gnd.n3254 gnd.n3253 0.152939
R13342 gnd.n3255 gnd.n3254 0.152939
R13343 gnd.n3256 gnd.n3255 0.152939
R13344 gnd.n3257 gnd.n3256 0.152939
R13345 gnd.n3258 gnd.n3257 0.152939
R13346 gnd.n3259 gnd.n3258 0.152939
R13347 gnd.n3260 gnd.n3259 0.152939
R13348 gnd.n3261 gnd.n3260 0.152939
R13349 gnd.n3262 gnd.n3261 0.152939
R13350 gnd.n3263 gnd.n3262 0.152939
R13351 gnd.n3264 gnd.n3263 0.152939
R13352 gnd.n5535 gnd.n3264 0.152939
R13353 gnd.n5535 gnd.n5534 0.152939
R13354 gnd.n3285 gnd.n3284 0.152939
R13355 gnd.n3286 gnd.n3285 0.152939
R13356 gnd.n3287 gnd.n3286 0.152939
R13357 gnd.n3288 gnd.n3287 0.152939
R13358 gnd.n3308 gnd.n3288 0.152939
R13359 gnd.n3309 gnd.n3308 0.152939
R13360 gnd.n3310 gnd.n3309 0.152939
R13361 gnd.n3311 gnd.n3310 0.152939
R13362 gnd.n3329 gnd.n3311 0.152939
R13363 gnd.n3330 gnd.n3329 0.152939
R13364 gnd.n3331 gnd.n3330 0.152939
R13365 gnd.n3332 gnd.n3331 0.152939
R13366 gnd.n3348 gnd.n3332 0.152939
R13367 gnd.n3349 gnd.n3348 0.152939
R13368 gnd.n3349 gnd.n82 0.152939
R13369 gnd.n7408 gnd.n82 0.152939
R13370 gnd.n4296 gnd.n4295 0.152939
R13371 gnd.n4297 gnd.n4296 0.152939
R13372 gnd.n4298 gnd.n4297 0.152939
R13373 gnd.n4301 gnd.n4298 0.152939
R13374 gnd.n4302 gnd.n4301 0.152939
R13375 gnd.n4303 gnd.n4302 0.152939
R13376 gnd.n4304 gnd.n4303 0.152939
R13377 gnd.n4304 gnd.n3996 0.152939
R13378 gnd.n4367 gnd.n3996 0.152939
R13379 gnd.n4368 gnd.n4367 0.152939
R13380 gnd.n4369 gnd.n4368 0.152939
R13381 gnd.n4369 gnd.n3992 0.152939
R13382 gnd.n4375 gnd.n3992 0.152939
R13383 gnd.n4376 gnd.n4375 0.152939
R13384 gnd.n4377 gnd.n4376 0.152939
R13385 gnd.n4377 gnd.n3988 0.152939
R13386 gnd.n4383 gnd.n3988 0.152939
R13387 gnd.n4384 gnd.n4383 0.152939
R13388 gnd.n4385 gnd.n4384 0.152939
R13389 gnd.n4385 gnd.n3984 0.152939
R13390 gnd.n4392 gnd.n3984 0.152939
R13391 gnd.n4393 gnd.n4392 0.152939
R13392 gnd.n4394 gnd.n4393 0.152939
R13393 gnd.n4394 gnd.n3920 0.152939
R13394 gnd.n4408 gnd.n3920 0.152939
R13395 gnd.n4409 gnd.n4408 0.152939
R13396 gnd.n4410 gnd.n4409 0.152939
R13397 gnd.n4410 gnd.n3906 0.152939
R13398 gnd.n4424 gnd.n3906 0.152939
R13399 gnd.n4425 gnd.n4424 0.152939
R13400 gnd.n4426 gnd.n4425 0.152939
R13401 gnd.n4426 gnd.n3892 0.152939
R13402 gnd.n4440 gnd.n3892 0.152939
R13403 gnd.n4441 gnd.n4440 0.152939
R13404 gnd.n4442 gnd.n4441 0.152939
R13405 gnd.n4442 gnd.n3878 0.152939
R13406 gnd.n4456 gnd.n3878 0.152939
R13407 gnd.n4457 gnd.n4456 0.152939
R13408 gnd.n4458 gnd.n4457 0.152939
R13409 gnd.n4458 gnd.n3861 0.152939
R13410 gnd.n4483 gnd.n3861 0.152939
R13411 gnd.n4484 gnd.n4483 0.152939
R13412 gnd.n4485 gnd.n4484 0.152939
R13413 gnd.n4487 gnd.n4485 0.152939
R13414 gnd.n4487 gnd.n4486 0.152939
R13415 gnd.n4486 gnd.n2982 0.152939
R13416 gnd.n2983 gnd.n2982 0.152939
R13417 gnd.n2984 gnd.n2983 0.152939
R13418 gnd.n4517 gnd.n2984 0.152939
R13419 gnd.n4518 gnd.n4517 0.152939
R13420 gnd.n4519 gnd.n4518 0.152939
R13421 gnd.n4519 gnd.n3744 0.152939
R13422 gnd.n4574 gnd.n3744 0.152939
R13423 gnd.n4575 gnd.n4574 0.152939
R13424 gnd.n4576 gnd.n4575 0.152939
R13425 gnd.n4577 gnd.n4576 0.152939
R13426 gnd.n4577 gnd.n3722 0.152939
R13427 gnd.n4614 gnd.n3722 0.152939
R13428 gnd.n4615 gnd.n4614 0.152939
R13429 gnd.n4616 gnd.n4615 0.152939
R13430 gnd.n4616 gnd.n3696 0.152939
R13431 gnd.n4658 gnd.n3696 0.152939
R13432 gnd.n4659 gnd.n4658 0.152939
R13433 gnd.n4660 gnd.n4659 0.152939
R13434 gnd.n4661 gnd.n4660 0.152939
R13435 gnd.n4661 gnd.n3676 0.152939
R13436 gnd.n4710 gnd.n3676 0.152939
R13437 gnd.n4711 gnd.n4710 0.152939
R13438 gnd.n4712 gnd.n4711 0.152939
R13439 gnd.n4713 gnd.n4712 0.152939
R13440 gnd.n4714 gnd.n4713 0.152939
R13441 gnd.n4716 gnd.n4714 0.152939
R13442 gnd.n4717 gnd.n4716 0.152939
R13443 gnd.n4717 gnd.n3638 0.152939
R13444 gnd.n4772 gnd.n3638 0.152939
R13445 gnd.n4773 gnd.n4772 0.152939
R13446 gnd.n4774 gnd.n4773 0.152939
R13447 gnd.n4774 gnd.n3616 0.152939
R13448 gnd.n4832 gnd.n3616 0.152939
R13449 gnd.n4833 gnd.n4832 0.152939
R13450 gnd.n4834 gnd.n4833 0.152939
R13451 gnd.n4834 gnd.n3598 0.152939
R13452 gnd.n4860 gnd.n3598 0.152939
R13453 gnd.n4861 gnd.n4860 0.152939
R13454 gnd.n4862 gnd.n4861 0.152939
R13455 gnd.n4862 gnd.n3580 0.152939
R13456 gnd.n4885 gnd.n3580 0.152939
R13457 gnd.n4886 gnd.n4885 0.152939
R13458 gnd.n4887 gnd.n4886 0.152939
R13459 gnd.n4888 gnd.n4887 0.152939
R13460 gnd.n4888 gnd.n3551 0.152939
R13461 gnd.n4941 gnd.n3551 0.152939
R13462 gnd.n4942 gnd.n4941 0.152939
R13463 gnd.n4943 gnd.n4942 0.152939
R13464 gnd.n4944 gnd.n4943 0.152939
R13465 gnd.n4944 gnd.n3520 0.152939
R13466 gnd.n5172 gnd.n3520 0.152939
R13467 gnd.n5173 gnd.n5172 0.152939
R13468 gnd.n5174 gnd.n5173 0.152939
R13469 gnd.n5174 gnd.n3508 0.152939
R13470 gnd.n5190 gnd.n3508 0.152939
R13471 gnd.n5191 gnd.n5190 0.152939
R13472 gnd.n5192 gnd.n5191 0.152939
R13473 gnd.n5192 gnd.n3497 0.152939
R13474 gnd.n5207 gnd.n3497 0.152939
R13475 gnd.n5208 gnd.n5207 0.152939
R13476 gnd.n5209 gnd.n5208 0.152939
R13477 gnd.n5209 gnd.n3485 0.152939
R13478 gnd.n5224 gnd.n3485 0.152939
R13479 gnd.n5225 gnd.n5224 0.152939
R13480 gnd.n5226 gnd.n5225 0.152939
R13481 gnd.n5226 gnd.n3473 0.152939
R13482 gnd.n5241 gnd.n3473 0.152939
R13483 gnd.n5242 gnd.n5241 0.152939
R13484 gnd.n5243 gnd.n5242 0.152939
R13485 gnd.n5243 gnd.n3461 0.152939
R13486 gnd.n5258 gnd.n3461 0.152939
R13487 gnd.n5259 gnd.n5258 0.152939
R13488 gnd.n5260 gnd.n5259 0.152939
R13489 gnd.n5262 gnd.n5260 0.152939
R13490 gnd.n5262 gnd.n5261 0.152939
R13491 gnd.n5261 gnd.n3449 0.152939
R13492 gnd.n5280 gnd.n3449 0.152939
R13493 gnd.n5281 gnd.n5280 0.152939
R13494 gnd.n5282 gnd.n5281 0.152939
R13495 gnd.n5283 gnd.n5282 0.152939
R13496 gnd.n5284 gnd.n5283 0.152939
R13497 gnd.n5286 gnd.n5284 0.152939
R13498 gnd.n5287 gnd.n5286 0.152939
R13499 gnd.n5287 gnd.n3413 0.152939
R13500 gnd.n5349 gnd.n3413 0.152939
R13501 gnd.n5350 gnd.n5349 0.152939
R13502 gnd.n5351 gnd.n5350 0.152939
R13503 gnd.n5351 gnd.n3409 0.152939
R13504 gnd.n5357 gnd.n3409 0.152939
R13505 gnd.n5358 gnd.n5357 0.152939
R13506 gnd.n5359 gnd.n5358 0.152939
R13507 gnd.n5359 gnd.n3405 0.152939
R13508 gnd.n5365 gnd.n3405 0.152939
R13509 gnd.n5366 gnd.n5365 0.152939
R13510 gnd.n5367 gnd.n5366 0.152939
R13511 gnd.n5368 gnd.n5367 0.152939
R13512 gnd.n5369 gnd.n5368 0.152939
R13513 gnd.n5372 gnd.n5369 0.152939
R13514 gnd.n5373 gnd.n5372 0.152939
R13515 gnd.n4152 gnd.n4093 0.152939
R13516 gnd.n4158 gnd.n4093 0.152939
R13517 gnd.n4159 gnd.n4158 0.152939
R13518 gnd.n4160 gnd.n4159 0.152939
R13519 gnd.n4160 gnd.n4091 0.152939
R13520 gnd.n4166 gnd.n4091 0.152939
R13521 gnd.n4167 gnd.n4166 0.152939
R13522 gnd.n4169 gnd.n4167 0.152939
R13523 gnd.n4169 gnd.n4168 0.152939
R13524 gnd.n4168 gnd.n4076 0.152939
R13525 gnd.n4077 gnd.n4076 0.152939
R13526 gnd.n4078 gnd.n4077 0.152939
R13527 gnd.n4181 gnd.n4078 0.152939
R13528 gnd.n4182 gnd.n4181 0.152939
R13529 gnd.n4183 gnd.n4182 0.152939
R13530 gnd.n4184 gnd.n4183 0.152939
R13531 gnd.n4185 gnd.n4184 0.152939
R13532 gnd.n4185 gnd.n4049 0.152939
R13533 gnd.n4254 gnd.n4049 0.152939
R13534 gnd.n4255 gnd.n4254 0.152939
R13535 gnd.n4107 gnd.n2448 0.152939
R13536 gnd.n4115 gnd.n4107 0.152939
R13537 gnd.n4116 gnd.n4115 0.152939
R13538 gnd.n4117 gnd.n4116 0.152939
R13539 gnd.n4117 gnd.n4105 0.152939
R13540 gnd.n4125 gnd.n4105 0.152939
R13541 gnd.n4126 gnd.n4125 0.152939
R13542 gnd.n4127 gnd.n4126 0.152939
R13543 gnd.n4127 gnd.n4103 0.152939
R13544 gnd.n4135 gnd.n4103 0.152939
R13545 gnd.n4136 gnd.n4135 0.152939
R13546 gnd.n4137 gnd.n4136 0.152939
R13547 gnd.n4137 gnd.n4101 0.152939
R13548 gnd.n4145 gnd.n4101 0.152939
R13549 gnd.n4146 gnd.n4145 0.152939
R13550 gnd.n4147 gnd.n4146 0.152939
R13551 gnd.n4147 gnd.n4094 0.152939
R13552 gnd.n4151 gnd.n4094 0.152939
R13553 gnd.n6099 gnd.n2543 0.152939
R13554 gnd.n2568 gnd.n2543 0.152939
R13555 gnd.n2569 gnd.n2568 0.152939
R13556 gnd.n2570 gnd.n2569 0.152939
R13557 gnd.n2587 gnd.n2570 0.152939
R13558 gnd.n2588 gnd.n2587 0.152939
R13559 gnd.n2589 gnd.n2588 0.152939
R13560 gnd.n2590 gnd.n2589 0.152939
R13561 gnd.n2607 gnd.n2590 0.152939
R13562 gnd.n2608 gnd.n2607 0.152939
R13563 gnd.n2609 gnd.n2608 0.152939
R13564 gnd.n2610 gnd.n2609 0.152939
R13565 gnd.n2627 gnd.n2610 0.152939
R13566 gnd.n2628 gnd.n2627 0.152939
R13567 gnd.n2629 gnd.n2628 0.152939
R13568 gnd.n2630 gnd.n2629 0.152939
R13569 gnd.n2786 gnd.n2785 0.152939
R13570 gnd.n2787 gnd.n2786 0.152939
R13571 gnd.n2788 gnd.n2787 0.152939
R13572 gnd.n2789 gnd.n2788 0.152939
R13573 gnd.n2790 gnd.n2789 0.152939
R13574 gnd.n2791 gnd.n2790 0.152939
R13575 gnd.n2792 gnd.n2791 0.152939
R13576 gnd.n2793 gnd.n2792 0.152939
R13577 gnd.n2794 gnd.n2793 0.152939
R13578 gnd.n2795 gnd.n2794 0.152939
R13579 gnd.n2796 gnd.n2795 0.152939
R13580 gnd.n2797 gnd.n2796 0.152939
R13581 gnd.n2798 gnd.n2797 0.152939
R13582 gnd.n2799 gnd.n2798 0.152939
R13583 gnd.n2800 gnd.n2799 0.152939
R13584 gnd.n2801 gnd.n2800 0.152939
R13585 gnd.n2802 gnd.n2801 0.152939
R13586 gnd.n2805 gnd.n2802 0.152939
R13587 gnd.n2806 gnd.n2805 0.152939
R13588 gnd.n2807 gnd.n2806 0.152939
R13589 gnd.n2808 gnd.n2807 0.152939
R13590 gnd.n2809 gnd.n2808 0.152939
R13591 gnd.n2810 gnd.n2809 0.152939
R13592 gnd.n2811 gnd.n2810 0.152939
R13593 gnd.n2812 gnd.n2811 0.152939
R13594 gnd.n2910 gnd.n2909 0.152939
R13595 gnd.n2909 gnd.n2815 0.152939
R13596 gnd.n2816 gnd.n2815 0.152939
R13597 gnd.n2817 gnd.n2816 0.152939
R13598 gnd.n2818 gnd.n2817 0.152939
R13599 gnd.n2819 gnd.n2818 0.152939
R13600 gnd.n2820 gnd.n2819 0.152939
R13601 gnd.n2821 gnd.n2820 0.152939
R13602 gnd.n2889 gnd.n2821 0.152939
R13603 gnd.n2889 gnd.n2888 0.152939
R13604 gnd.n2888 gnd.n2887 0.152939
R13605 gnd.n2887 gnd.n2825 0.152939
R13606 gnd.n2826 gnd.n2825 0.152939
R13607 gnd.n2827 gnd.n2826 0.152939
R13608 gnd.n2828 gnd.n2827 0.152939
R13609 gnd.n2829 gnd.n2828 0.152939
R13610 gnd.n2830 gnd.n2829 0.152939
R13611 gnd.n2831 gnd.n2830 0.152939
R13612 gnd.n2832 gnd.n2831 0.152939
R13613 gnd.n2833 gnd.n2832 0.152939
R13614 gnd.n2834 gnd.n2833 0.152939
R13615 gnd.n2835 gnd.n2834 0.152939
R13616 gnd.n2836 gnd.n2835 0.152939
R13617 gnd.n2837 gnd.n2836 0.152939
R13618 gnd.n2838 gnd.n2837 0.152939
R13619 gnd.n2839 gnd.n2838 0.152939
R13620 gnd.n2840 gnd.n2839 0.152939
R13621 gnd.n2841 gnd.n2840 0.152939
R13622 gnd.n2847 gnd.n2841 0.152939
R13623 gnd.n2847 gnd.n2846 0.152939
R13624 gnd.n2385 gnd.n2384 0.152939
R13625 gnd.n2386 gnd.n2385 0.152939
R13626 gnd.n2387 gnd.n2386 0.152939
R13627 gnd.n2388 gnd.n2387 0.152939
R13628 gnd.n2389 gnd.n2388 0.152939
R13629 gnd.n2390 gnd.n2389 0.152939
R13630 gnd.n2391 gnd.n2390 0.152939
R13631 gnd.n2392 gnd.n2391 0.152939
R13632 gnd.n2393 gnd.n2392 0.152939
R13633 gnd.n2394 gnd.n2393 0.152939
R13634 gnd.n2395 gnd.n2394 0.152939
R13635 gnd.n2396 gnd.n2395 0.152939
R13636 gnd.n2397 gnd.n2396 0.152939
R13637 gnd.n2398 gnd.n2397 0.152939
R13638 gnd.n2399 gnd.n2398 0.152939
R13639 gnd.n2400 gnd.n2399 0.152939
R13640 gnd.n2401 gnd.n2400 0.152939
R13641 gnd.n2404 gnd.n2401 0.152939
R13642 gnd.n2405 gnd.n2404 0.152939
R13643 gnd.n2406 gnd.n2405 0.152939
R13644 gnd.n2407 gnd.n2406 0.152939
R13645 gnd.n2408 gnd.n2407 0.152939
R13646 gnd.n2409 gnd.n2408 0.152939
R13647 gnd.n2410 gnd.n2409 0.152939
R13648 gnd.n2411 gnd.n2410 0.152939
R13649 gnd.n2412 gnd.n2411 0.152939
R13650 gnd.n2413 gnd.n2412 0.152939
R13651 gnd.n2414 gnd.n2413 0.152939
R13652 gnd.n2415 gnd.n2414 0.152939
R13653 gnd.n2416 gnd.n2415 0.152939
R13654 gnd.n2417 gnd.n2416 0.152939
R13655 gnd.n2418 gnd.n2417 0.152939
R13656 gnd.n2419 gnd.n2418 0.152939
R13657 gnd.n2420 gnd.n2419 0.152939
R13658 gnd.n2421 gnd.n2420 0.152939
R13659 gnd.n2422 gnd.n2421 0.152939
R13660 gnd.n2423 gnd.n2422 0.152939
R13661 gnd.n2426 gnd.n2423 0.152939
R13662 gnd.n2427 gnd.n2426 0.152939
R13663 gnd.n2428 gnd.n2427 0.152939
R13664 gnd.n2429 gnd.n2428 0.152939
R13665 gnd.n2430 gnd.n2429 0.152939
R13666 gnd.n2431 gnd.n2430 0.152939
R13667 gnd.n2432 gnd.n2431 0.152939
R13668 gnd.n2433 gnd.n2432 0.152939
R13669 gnd.n2434 gnd.n2433 0.152939
R13670 gnd.n2435 gnd.n2434 0.152939
R13671 gnd.n2436 gnd.n2435 0.152939
R13672 gnd.n2437 gnd.n2436 0.152939
R13673 gnd.n2438 gnd.n2437 0.152939
R13674 gnd.n2439 gnd.n2438 0.152939
R13675 gnd.n2440 gnd.n2439 0.152939
R13676 gnd.n2441 gnd.n2440 0.152939
R13677 gnd.n2442 gnd.n2441 0.152939
R13678 gnd.n2443 gnd.n2442 0.152939
R13679 gnd.n2444 gnd.n2443 0.152939
R13680 gnd.n6159 gnd.n2444 0.152939
R13681 gnd.n6159 gnd.n6158 0.152939
R13682 gnd.n2459 gnd.n2458 0.152939
R13683 gnd.n2460 gnd.n2459 0.152939
R13684 gnd.n2461 gnd.n2460 0.152939
R13685 gnd.n2481 gnd.n2461 0.152939
R13686 gnd.n2482 gnd.n2481 0.152939
R13687 gnd.n2483 gnd.n2482 0.152939
R13688 gnd.n2484 gnd.n2483 0.152939
R13689 gnd.n2500 gnd.n2484 0.152939
R13690 gnd.n2501 gnd.n2500 0.152939
R13691 gnd.n2502 gnd.n2501 0.152939
R13692 gnd.n2503 gnd.n2502 0.152939
R13693 gnd.n2521 gnd.n2503 0.152939
R13694 gnd.n2522 gnd.n2521 0.152939
R13695 gnd.n2523 gnd.n2522 0.152939
R13696 gnd.n2524 gnd.n2523 0.152939
R13697 gnd.n6099 gnd.n2524 0.152939
R13698 gnd.n4072 gnd.n4071 0.152939
R13699 gnd.n4072 gnd.n4066 0.152939
R13700 gnd.n4213 gnd.n4066 0.152939
R13701 gnd.n4214 gnd.n4213 0.152939
R13702 gnd.n4216 gnd.n4214 0.152939
R13703 gnd.n4216 gnd.n4215 0.152939
R13704 gnd.n4215 gnd.n4063 0.152939
R13705 gnd.n813 gnd.n808 0.152939
R13706 gnd.n814 gnd.n813 0.152939
R13707 gnd.n815 gnd.n814 0.152939
R13708 gnd.n820 gnd.n815 0.152939
R13709 gnd.n821 gnd.n820 0.152939
R13710 gnd.n822 gnd.n821 0.152939
R13711 gnd.n823 gnd.n822 0.152939
R13712 gnd.n828 gnd.n823 0.152939
R13713 gnd.n829 gnd.n828 0.152939
R13714 gnd.n830 gnd.n829 0.152939
R13715 gnd.n831 gnd.n830 0.152939
R13716 gnd.n836 gnd.n831 0.152939
R13717 gnd.n837 gnd.n836 0.152939
R13718 gnd.n838 gnd.n837 0.152939
R13719 gnd.n839 gnd.n838 0.152939
R13720 gnd.n844 gnd.n839 0.152939
R13721 gnd.n845 gnd.n844 0.152939
R13722 gnd.n846 gnd.n845 0.152939
R13723 gnd.n847 gnd.n846 0.152939
R13724 gnd.n852 gnd.n847 0.152939
R13725 gnd.n853 gnd.n852 0.152939
R13726 gnd.n854 gnd.n853 0.152939
R13727 gnd.n855 gnd.n854 0.152939
R13728 gnd.n860 gnd.n855 0.152939
R13729 gnd.n861 gnd.n860 0.152939
R13730 gnd.n862 gnd.n861 0.152939
R13731 gnd.n863 gnd.n862 0.152939
R13732 gnd.n868 gnd.n863 0.152939
R13733 gnd.n869 gnd.n868 0.152939
R13734 gnd.n870 gnd.n869 0.152939
R13735 gnd.n871 gnd.n870 0.152939
R13736 gnd.n876 gnd.n871 0.152939
R13737 gnd.n877 gnd.n876 0.152939
R13738 gnd.n878 gnd.n877 0.152939
R13739 gnd.n879 gnd.n878 0.152939
R13740 gnd.n884 gnd.n879 0.152939
R13741 gnd.n885 gnd.n884 0.152939
R13742 gnd.n886 gnd.n885 0.152939
R13743 gnd.n887 gnd.n886 0.152939
R13744 gnd.n892 gnd.n887 0.152939
R13745 gnd.n893 gnd.n892 0.152939
R13746 gnd.n894 gnd.n893 0.152939
R13747 gnd.n895 gnd.n894 0.152939
R13748 gnd.n900 gnd.n895 0.152939
R13749 gnd.n901 gnd.n900 0.152939
R13750 gnd.n902 gnd.n901 0.152939
R13751 gnd.n903 gnd.n902 0.152939
R13752 gnd.n908 gnd.n903 0.152939
R13753 gnd.n909 gnd.n908 0.152939
R13754 gnd.n910 gnd.n909 0.152939
R13755 gnd.n911 gnd.n910 0.152939
R13756 gnd.n916 gnd.n911 0.152939
R13757 gnd.n917 gnd.n916 0.152939
R13758 gnd.n918 gnd.n917 0.152939
R13759 gnd.n919 gnd.n918 0.152939
R13760 gnd.n924 gnd.n919 0.152939
R13761 gnd.n925 gnd.n924 0.152939
R13762 gnd.n926 gnd.n925 0.152939
R13763 gnd.n927 gnd.n926 0.152939
R13764 gnd.n932 gnd.n927 0.152939
R13765 gnd.n933 gnd.n932 0.152939
R13766 gnd.n934 gnd.n933 0.152939
R13767 gnd.n935 gnd.n934 0.152939
R13768 gnd.n940 gnd.n935 0.152939
R13769 gnd.n941 gnd.n940 0.152939
R13770 gnd.n942 gnd.n941 0.152939
R13771 gnd.n943 gnd.n942 0.152939
R13772 gnd.n948 gnd.n943 0.152939
R13773 gnd.n949 gnd.n948 0.152939
R13774 gnd.n950 gnd.n949 0.152939
R13775 gnd.n951 gnd.n950 0.152939
R13776 gnd.n956 gnd.n951 0.152939
R13777 gnd.n957 gnd.n956 0.152939
R13778 gnd.n958 gnd.n957 0.152939
R13779 gnd.n959 gnd.n958 0.152939
R13780 gnd.n964 gnd.n959 0.152939
R13781 gnd.n965 gnd.n964 0.152939
R13782 gnd.n966 gnd.n965 0.152939
R13783 gnd.n967 gnd.n966 0.152939
R13784 gnd.n972 gnd.n967 0.152939
R13785 gnd.n973 gnd.n972 0.152939
R13786 gnd.n974 gnd.n973 0.152939
R13787 gnd.n975 gnd.n974 0.152939
R13788 gnd.n4070 gnd.n975 0.152939
R13789 gnd.n4400 gnd.n3927 0.152939
R13790 gnd.n4401 gnd.n4400 0.152939
R13791 gnd.n4402 gnd.n4401 0.152939
R13792 gnd.n4402 gnd.n3912 0.152939
R13793 gnd.n4416 gnd.n3912 0.152939
R13794 gnd.n4417 gnd.n4416 0.152939
R13795 gnd.n4418 gnd.n4417 0.152939
R13796 gnd.n4418 gnd.n3899 0.152939
R13797 gnd.n4432 gnd.n3899 0.152939
R13798 gnd.n4433 gnd.n4432 0.152939
R13799 gnd.n4434 gnd.n4433 0.152939
R13800 gnd.n4434 gnd.n3885 0.152939
R13801 gnd.n4448 gnd.n3885 0.152939
R13802 gnd.n4449 gnd.n4448 0.152939
R13803 gnd.n4450 gnd.n4449 0.152939
R13804 gnd.n4450 gnd.n3871 0.152939
R13805 gnd.n4464 gnd.n3871 0.152939
R13806 gnd.n4465 gnd.n4464 0.152939
R13807 gnd.n4477 gnd.n4465 0.152939
R13808 gnd.n4477 gnd.n4476 0.152939
R13809 gnd.n4476 gnd.n4475 0.152939
R13810 gnd.n4475 gnd.n4466 0.152939
R13811 gnd.n4471 gnd.n4466 0.152939
R13812 gnd.n4471 gnd.n4470 0.152939
R13813 gnd.n4470 gnd.n2994 0.152939
R13814 gnd.n5831 gnd.n2994 0.152939
R13815 gnd.n5831 gnd.n5830 0.152939
R13816 gnd.n5830 gnd.n5829 0.152939
R13817 gnd.n5829 gnd.n2995 0.152939
R13818 gnd.n5825 gnd.n2995 0.152939
R13819 gnd.n5825 gnd.n5824 0.152939
R13820 gnd.n5824 gnd.n5823 0.152939
R13821 gnd.n5823 gnd.n3000 0.152939
R13822 gnd.n5819 gnd.n3000 0.152939
R13823 gnd.n5819 gnd.n5818 0.152939
R13824 gnd.n5818 gnd.n5817 0.152939
R13825 gnd.n5817 gnd.n3005 0.152939
R13826 gnd.n5813 gnd.n3005 0.152939
R13827 gnd.n5813 gnd.n5812 0.152939
R13828 gnd.n5812 gnd.n5811 0.152939
R13829 gnd.n5811 gnd.n3010 0.152939
R13830 gnd.n5807 gnd.n3010 0.152939
R13831 gnd.n5807 gnd.n5806 0.152939
R13832 gnd.n5806 gnd.n5805 0.152939
R13833 gnd.n5805 gnd.n3015 0.152939
R13834 gnd.n5801 gnd.n3015 0.152939
R13835 gnd.n5801 gnd.n5800 0.152939
R13836 gnd.n5800 gnd.n5799 0.152939
R13837 gnd.n5799 gnd.n3020 0.152939
R13838 gnd.n5795 gnd.n3020 0.152939
R13839 gnd.n5795 gnd.n5794 0.152939
R13840 gnd.n5794 gnd.n5793 0.152939
R13841 gnd.n5793 gnd.n3025 0.152939
R13842 gnd.n5789 gnd.n3025 0.152939
R13843 gnd.n5789 gnd.n5788 0.152939
R13844 gnd.n5788 gnd.n5787 0.152939
R13845 gnd.n5787 gnd.n3030 0.152939
R13846 gnd.n5783 gnd.n3030 0.152939
R13847 gnd.n5783 gnd.n5782 0.152939
R13848 gnd.n5782 gnd.n5781 0.152939
R13849 gnd.n5781 gnd.n3035 0.152939
R13850 gnd.n5777 gnd.n3035 0.152939
R13851 gnd.n5777 gnd.n5776 0.152939
R13852 gnd.n5776 gnd.n5775 0.152939
R13853 gnd.n5775 gnd.n3040 0.152939
R13854 gnd.n5771 gnd.n3040 0.152939
R13855 gnd.n5771 gnd.n5770 0.152939
R13856 gnd.n5770 gnd.n5769 0.152939
R13857 gnd.n5769 gnd.n3045 0.152939
R13858 gnd.n5765 gnd.n3045 0.152939
R13859 gnd.n5765 gnd.n5764 0.152939
R13860 gnd.n5764 gnd.n5763 0.152939
R13861 gnd.n5763 gnd.n3050 0.152939
R13862 gnd.n5759 gnd.n3050 0.152939
R13863 gnd.n5759 gnd.n5758 0.152939
R13864 gnd.n5758 gnd.n5757 0.152939
R13865 gnd.n5757 gnd.n3055 0.152939
R13866 gnd.n5753 gnd.n3055 0.152939
R13867 gnd.n5753 gnd.n5752 0.152939
R13868 gnd.n5752 gnd.n5751 0.152939
R13869 gnd.n5751 gnd.n3060 0.152939
R13870 gnd.n5747 gnd.n3060 0.152939
R13871 gnd.n5747 gnd.n5746 0.152939
R13872 gnd.n5746 gnd.n5745 0.152939
R13873 gnd.n5745 gnd.n3065 0.152939
R13874 gnd.n5741 gnd.n3065 0.152939
R13875 gnd.n5741 gnd.n5740 0.152939
R13876 gnd.n5740 gnd.n5739 0.152939
R13877 gnd.n5739 gnd.n3070 0.152939
R13878 gnd.n5735 gnd.n3070 0.152939
R13879 gnd.n5735 gnd.n5734 0.152939
R13880 gnd.n5734 gnd.n5733 0.152939
R13881 gnd.n5733 gnd.n3075 0.152939
R13882 gnd.n5729 gnd.n3075 0.152939
R13883 gnd.n5729 gnd.n5728 0.152939
R13884 gnd.n5728 gnd.n5727 0.152939
R13885 gnd.n5727 gnd.n3080 0.152939
R13886 gnd.n5723 gnd.n3080 0.152939
R13887 gnd.n5723 gnd.n5722 0.152939
R13888 gnd.n5722 gnd.n5721 0.152939
R13889 gnd.n5721 gnd.n3085 0.152939
R13890 gnd.n4284 gnd.n4026 0.152939
R13891 gnd.n4285 gnd.n4284 0.152939
R13892 gnd.n4286 gnd.n4285 0.152939
R13893 gnd.n4286 gnd.n4014 0.152939
R13894 gnd.n4320 gnd.n4014 0.152939
R13895 gnd.n4321 gnd.n4320 0.152939
R13896 gnd.n4322 gnd.n4321 0.152939
R13897 gnd.n4322 gnd.n4008 0.152939
R13898 gnd.n4334 gnd.n4008 0.152939
R13899 gnd.n4335 gnd.n4334 0.152939
R13900 gnd.n4336 gnd.n4335 0.152939
R13901 gnd.n4336 gnd.n4002 0.152939
R13902 gnd.n4360 gnd.n4002 0.152939
R13903 gnd.n4360 gnd.n4359 0.152939
R13904 gnd.n4359 gnd.n4358 0.152939
R13905 gnd.n4358 gnd.n4003 0.152939
R13906 gnd.n4354 gnd.n4003 0.152939
R13907 gnd.n4354 gnd.n2643 0.152939
R13908 gnd.n6038 gnd.n2643 0.152939
R13909 gnd.n6038 gnd.n6037 0.152939
R13910 gnd.n6025 gnd.n2667 0.152939
R13911 gnd.n6025 gnd.n6024 0.152939
R13912 gnd.n6024 gnd.n6023 0.152939
R13913 gnd.n6023 gnd.n2669 0.152939
R13914 gnd.n6019 gnd.n2669 0.152939
R13915 gnd.n6019 gnd.n6018 0.152939
R13916 gnd.n3979 gnd.n3933 0.152939
R13917 gnd.n3979 gnd.n3978 0.152939
R13918 gnd.n3978 gnd.n3977 0.152939
R13919 gnd.n3977 gnd.n3934 0.152939
R13920 gnd.n3973 gnd.n3934 0.152939
R13921 gnd.n3973 gnd.n3972 0.152939
R13922 gnd.n3972 gnd.n3971 0.152939
R13923 gnd.n3971 gnd.n3938 0.152939
R13924 gnd.n3967 gnd.n3938 0.152939
R13925 gnd.n3967 gnd.n3966 0.152939
R13926 gnd.n3966 gnd.n3965 0.152939
R13927 gnd.n3965 gnd.n3942 0.152939
R13928 gnd.n3961 gnd.n3942 0.152939
R13929 gnd.n3961 gnd.n3960 0.152939
R13930 gnd.n3960 gnd.n3959 0.152939
R13931 gnd.n3959 gnd.n3946 0.152939
R13932 gnd.n3955 gnd.n3946 0.152939
R13933 gnd.n3955 gnd.n3954 0.152939
R13934 gnd.n3954 gnd.n3953 0.152939
R13935 gnd.n3953 gnd.n3950 0.152939
R13936 gnd.n3950 gnd.n3854 0.152939
R13937 gnd.n4496 gnd.n3854 0.152939
R13938 gnd.n4497 gnd.n4496 0.152939
R13939 gnd.n4498 gnd.n4497 0.152939
R13940 gnd.n4498 gnd.n3852 0.152939
R13941 gnd.n4504 gnd.n3852 0.152939
R13942 gnd.n4505 gnd.n4504 0.152939
R13943 gnd.n4512 gnd.n4505 0.152939
R13944 gnd.n4512 gnd.n4511 0.152939
R13945 gnd.n4511 gnd.n4510 0.152939
R13946 gnd.n4510 gnd.n4506 0.152939
R13947 gnd.n4506 gnd.n3736 0.152939
R13948 gnd.n4584 gnd.n3736 0.152939
R13949 gnd.n4585 gnd.n4584 0.152939
R13950 gnd.n4599 gnd.n4585 0.152939
R13951 gnd.n4599 gnd.n4598 0.152939
R13952 gnd.n4598 gnd.n4597 0.152939
R13953 gnd.n4597 gnd.n4586 0.152939
R13954 gnd.n4593 gnd.n4586 0.152939
R13955 gnd.n4593 gnd.n4592 0.152939
R13956 gnd.n4592 gnd.n3689 0.152939
R13957 gnd.n4668 gnd.n3689 0.152939
R13958 gnd.n4669 gnd.n4668 0.152939
R13959 gnd.n4696 gnd.n4669 0.152939
R13960 gnd.n4696 gnd.n4695 0.152939
R13961 gnd.n4695 gnd.n4694 0.152939
R13962 gnd.n4694 gnd.n4670 0.152939
R13963 gnd.n4690 gnd.n4670 0.152939
R13964 gnd.n4690 gnd.n4689 0.152939
R13965 gnd.n4689 gnd.n4688 0.152939
R13966 gnd.n4688 gnd.n4674 0.152939
R13967 gnd.n4684 gnd.n4674 0.152939
R13968 gnd.n4684 gnd.n4683 0.152939
R13969 gnd.n4683 gnd.n4682 0.152939
R13970 gnd.n4682 gnd.n3630 0.152939
R13971 gnd.n4815 gnd.n3630 0.152939
R13972 gnd.n4815 gnd.n4814 0.152939
R13973 gnd.n4814 gnd.n4813 0.152939
R13974 gnd.n4813 gnd.n3631 0.152939
R13975 gnd.n4809 gnd.n3631 0.152939
R13976 gnd.n4809 gnd.n4808 0.152939
R13977 gnd.n4808 gnd.n4807 0.152939
R13978 gnd.n4807 gnd.n4792 0.152939
R13979 gnd.n4803 gnd.n4792 0.152939
R13980 gnd.n4803 gnd.n4802 0.152939
R13981 gnd.n4802 gnd.n4801 0.152939
R13982 gnd.n4801 gnd.n4797 0.152939
R13983 gnd.n4797 gnd.n3565 0.152939
R13984 gnd.n4927 gnd.n3565 0.152939
R13985 gnd.n4927 gnd.n4926 0.152939
R13986 gnd.n4926 gnd.n4925 0.152939
R13987 gnd.n4925 gnd.n3566 0.152939
R13988 gnd.n4921 gnd.n3566 0.152939
R13989 gnd.n4921 gnd.n4920 0.152939
R13990 gnd.n4920 gnd.n4919 0.152939
R13991 gnd.n4919 gnd.n3513 0.152939
R13992 gnd.n5180 gnd.n3513 0.152939
R13993 gnd.n5181 gnd.n5180 0.152939
R13994 gnd.n5182 gnd.n5181 0.152939
R13995 gnd.n5182 gnd.n3503 0.152939
R13996 gnd.n5198 gnd.n3503 0.152939
R13997 gnd.n5199 gnd.n5198 0.152939
R13998 gnd.n5200 gnd.n5199 0.152939
R13999 gnd.n5200 gnd.n3491 0.152939
R14000 gnd.n5215 gnd.n3491 0.152939
R14001 gnd.n5216 gnd.n5215 0.152939
R14002 gnd.n5217 gnd.n5216 0.152939
R14003 gnd.n5217 gnd.n3479 0.152939
R14004 gnd.n5232 gnd.n3479 0.152939
R14005 gnd.n5233 gnd.n5232 0.152939
R14006 gnd.n5234 gnd.n5233 0.152939
R14007 gnd.n5234 gnd.n3466 0.152939
R14008 gnd.n5249 gnd.n3466 0.152939
R14009 gnd.n5250 gnd.n5249 0.152939
R14010 gnd.n5251 gnd.n5250 0.152939
R14011 gnd.n5251 gnd.n3455 0.152939
R14012 gnd.n5269 gnd.n3455 0.152939
R14013 gnd.n5270 gnd.n5269 0.152939
R14014 gnd.n5271 gnd.n5270 0.152939
R14015 gnd.n5271 gnd.n3094 0.152939
R14016 gnd.n5714 gnd.n3094 0.152939
R14017 gnd.n5713 gnd.n3095 0.152939
R14018 gnd.n5709 gnd.n3095 0.152939
R14019 gnd.n5709 gnd.n5708 0.152939
R14020 gnd.n5708 gnd.n5707 0.152939
R14021 gnd.n5707 gnd.n3099 0.152939
R14022 gnd.n5703 gnd.n3099 0.152939
R14023 gnd.n5342 gnd.n5304 0.152939
R14024 gnd.n5342 gnd.n5341 0.152939
R14025 gnd.n5341 gnd.n5340 0.152939
R14026 gnd.n5340 gnd.n5305 0.152939
R14027 gnd.n5336 gnd.n5305 0.152939
R14028 gnd.n5336 gnd.n5335 0.152939
R14029 gnd.n5335 gnd.n5334 0.152939
R14030 gnd.n5334 gnd.n5310 0.152939
R14031 gnd.n5330 gnd.n5310 0.152939
R14032 gnd.n5330 gnd.n3399 0.152939
R14033 gnd.n5391 gnd.n3399 0.152939
R14034 gnd.n5392 gnd.n5391 0.152939
R14035 gnd.n5393 gnd.n5392 0.152939
R14036 gnd.n5393 gnd.n3394 0.152939
R14037 gnd.n5406 gnd.n3394 0.152939
R14038 gnd.n5407 gnd.n5406 0.152939
R14039 gnd.n5412 gnd.n5407 0.152939
R14040 gnd.n5412 gnd.n5411 0.152939
R14041 gnd.n5411 gnd.n5410 0.152939
R14042 gnd.n5410 gnd.n67 0.152939
R14043 gnd.n7418 gnd.n7417 0.145814
R14044 gnd.n4256 gnd.n4255 0.145814
R14045 gnd.n4256 gnd.n4026 0.145814
R14046 gnd.n7418 gnd.n67 0.145814
R14047 gnd.n6018 gnd.n6017 0.128549
R14048 gnd.n5703 gnd.n5702 0.128549
R14049 gnd.n1643 gnd.n0 0.127478
R14050 gnd.n4295 gnd.n2544 0.0919634
R14051 gnd.n5373 gnd.n83 0.0919634
R14052 gnd.n1644 gnd.n1560 0.0767195
R14053 gnd.n1644 gnd.n1558 0.0767195
R14054 gnd.n6017 gnd.n2638 0.063
R14055 gnd.n5702 gnd.n3104 0.063
R14056 gnd.n401 gnd.n83 0.0614756
R14057 gnd.n4063 gnd.n2544 0.0614756
R14058 gnd.n3272 gnd.n3104 0.0538288
R14059 gnd.n7354 gnd.n386 0.0538288
R14060 gnd.n6157 gnd.n6156 0.0538288
R14061 gnd.n6045 gnd.n2638 0.0538288
R14062 gnd.n6335 gnd.n1048 0.0477147
R14063 gnd.n1500 gnd.n1396 0.0442063
R14064 gnd.n1514 gnd.n1396 0.0442063
R14065 gnd.n1515 gnd.n1514 0.0442063
R14066 gnd.n1516 gnd.n1515 0.0442063
R14067 gnd.n1516 gnd.n1384 0.0442063
R14068 gnd.n1530 gnd.n1384 0.0442063
R14069 gnd.n1531 gnd.n1530 0.0442063
R14070 gnd.n1532 gnd.n1531 0.0442063
R14071 gnd.n1532 gnd.n1371 0.0442063
R14072 gnd.n1741 gnd.n1371 0.0442063
R14073 gnd.n1744 gnd.n1743 0.0344674
R14074 gnd.n5524 gnd.n3272 0.0344674
R14075 gnd.n5524 gnd.n3274 0.0344674
R14076 gnd.n3298 gnd.n3274 0.0344674
R14077 gnd.n3299 gnd.n3298 0.0344674
R14078 gnd.n3300 gnd.n3299 0.0344674
R14079 gnd.n3301 gnd.n3300 0.0344674
R14080 gnd.n5317 gnd.n3301 0.0344674
R14081 gnd.n5317 gnd.n3319 0.0344674
R14082 gnd.n3320 gnd.n3319 0.0344674
R14083 gnd.n3321 gnd.n3320 0.0344674
R14084 gnd.n5323 gnd.n3321 0.0344674
R14085 gnd.n5323 gnd.n3339 0.0344674
R14086 gnd.n3340 gnd.n3339 0.0344674
R14087 gnd.n3341 gnd.n3340 0.0344674
R14088 gnd.n5400 gnd.n3341 0.0344674
R14089 gnd.n5400 gnd.n3356 0.0344674
R14090 gnd.n3357 gnd.n3356 0.0344674
R14091 gnd.n3358 gnd.n3357 0.0344674
R14092 gnd.n5420 gnd.n3358 0.0344674
R14093 gnd.n5421 gnd.n5420 0.0344674
R14094 gnd.n5421 gnd.n3387 0.0344674
R14095 gnd.n3387 gnd.n3382 0.0344674
R14096 gnd.n3383 gnd.n3382 0.0344674
R14097 gnd.n3384 gnd.n3383 0.0344674
R14098 gnd.n5431 gnd.n3384 0.0344674
R14099 gnd.n5431 gnd.n97 0.0344674
R14100 gnd.n98 gnd.n97 0.0344674
R14101 gnd.n99 gnd.n98 0.0344674
R14102 gnd.n7230 gnd.n99 0.0344674
R14103 gnd.n7230 gnd.n115 0.0344674
R14104 gnd.n116 gnd.n115 0.0344674
R14105 gnd.n117 gnd.n116 0.0344674
R14106 gnd.n7245 gnd.n117 0.0344674
R14107 gnd.n7245 gnd.n136 0.0344674
R14108 gnd.n137 gnd.n136 0.0344674
R14109 gnd.n138 gnd.n137 0.0344674
R14110 gnd.n7344 gnd.n138 0.0344674
R14111 gnd.n7344 gnd.n155 0.0344674
R14112 gnd.n156 gnd.n155 0.0344674
R14113 gnd.n157 gnd.n156 0.0344674
R14114 gnd.n173 gnd.n157 0.0344674
R14115 gnd.n7354 gnd.n173 0.0344674
R14116 gnd.n6156 gnd.n2450 0.0344674
R14117 gnd.n4080 gnd.n2450 0.0344674
R14118 gnd.n4080 gnd.n2472 0.0344674
R14119 gnd.n2473 gnd.n2472 0.0344674
R14120 gnd.n2474 gnd.n2473 0.0344674
R14121 gnd.n4086 gnd.n2474 0.0344674
R14122 gnd.n4086 gnd.n2491 0.0344674
R14123 gnd.n2492 gnd.n2491 0.0344674
R14124 gnd.n2493 gnd.n2492 0.0344674
R14125 gnd.n4176 gnd.n2493 0.0344674
R14126 gnd.n4176 gnd.n2511 0.0344674
R14127 gnd.n2512 gnd.n2511 0.0344674
R14128 gnd.n2513 gnd.n2512 0.0344674
R14129 gnd.n4179 gnd.n2513 0.0344674
R14130 gnd.n4179 gnd.n2532 0.0344674
R14131 gnd.n2533 gnd.n2532 0.0344674
R14132 gnd.n2534 gnd.n2533 0.0344674
R14133 gnd.n4058 gnd.n2534 0.0344674
R14134 gnd.n4244 gnd.n4058 0.0344674
R14135 gnd.n4245 gnd.n4244 0.0344674
R14136 gnd.n4245 gnd.n4044 0.0344674
R14137 gnd.n4044 gnd.n4040 0.0344674
R14138 gnd.n4041 gnd.n4040 0.0344674
R14139 gnd.n4269 gnd.n4041 0.0344674
R14140 gnd.n4269 gnd.n4042 0.0344674
R14141 gnd.n4042 gnd.n2559 0.0344674
R14142 gnd.n2560 gnd.n2559 0.0344674
R14143 gnd.n2561 gnd.n2560 0.0344674
R14144 gnd.n4012 gnd.n2561 0.0344674
R14145 gnd.n4012 gnd.n2577 0.0344674
R14146 gnd.n2578 gnd.n2577 0.0344674
R14147 gnd.n2579 gnd.n2578 0.0344674
R14148 gnd.n4006 gnd.n2579 0.0344674
R14149 gnd.n4006 gnd.n2598 0.0344674
R14150 gnd.n2599 gnd.n2598 0.0344674
R14151 gnd.n2600 gnd.n2599 0.0344674
R14152 gnd.n4345 gnd.n2600 0.0344674
R14153 gnd.n4345 gnd.n2618 0.0344674
R14154 gnd.n2619 gnd.n2618 0.0344674
R14155 gnd.n2620 gnd.n2619 0.0344674
R14156 gnd.n2637 gnd.n2620 0.0344674
R14157 gnd.n6045 gnd.n2637 0.0344674
R14158 gnd.n6016 gnd.n2674 0.0343753
R14159 gnd.n5701 gnd.n5700 0.0343753
R14160 gnd.n6036 gnd.n6035 0.0296328
R14161 gnd.n5303 gnd.n5302 0.0296328
R14162 gnd.n1364 gnd.n1363 0.0269946
R14163 gnd.n1754 gnd.n1752 0.0269946
R14164 gnd.n1753 gnd.n1346 0.0269946
R14165 gnd.n1773 gnd.n1772 0.0269946
R14166 gnd.n1775 gnd.n1774 0.0269946
R14167 gnd.n1340 gnd.n1338 0.0269946
R14168 gnd.n1785 gnd.n1783 0.0269946
R14169 gnd.n1784 gnd.n1319 0.0269946
R14170 gnd.n1804 gnd.n1803 0.0269946
R14171 gnd.n1806 gnd.n1805 0.0269946
R14172 gnd.n1314 gnd.n1312 0.0269946
R14173 gnd.n1816 gnd.n1814 0.0269946
R14174 gnd.n1815 gnd.n1293 0.0269946
R14175 gnd.n1835 gnd.n1834 0.0269946
R14176 gnd.n1837 gnd.n1836 0.0269946
R14177 gnd.n1288 gnd.n1286 0.0269946
R14178 gnd.n1847 gnd.n1845 0.0269946
R14179 gnd.n1846 gnd.n1268 0.0269946
R14180 gnd.n1866 gnd.n1865 0.0269946
R14181 gnd.n1868 gnd.n1867 0.0269946
R14182 gnd.n1262 gnd.n1260 0.0269946
R14183 gnd.n1878 gnd.n1876 0.0269946
R14184 gnd.n1877 gnd.n1243 0.0269946
R14185 gnd.n1897 gnd.n1896 0.0269946
R14186 gnd.n1899 gnd.n1898 0.0269946
R14187 gnd.n1237 gnd.n1235 0.0269946
R14188 gnd.n1909 gnd.n1907 0.0269946
R14189 gnd.n1908 gnd.n1218 0.0269946
R14190 gnd.n1928 gnd.n1927 0.0269946
R14191 gnd.n1930 gnd.n1929 0.0269946
R14192 gnd.n1212 gnd.n1211 0.0269946
R14193 gnd.n1940 gnd.n1207 0.0269946
R14194 gnd.n1939 gnd.n1209 0.0269946
R14195 gnd.n1208 gnd.n1190 0.0269946
R14196 gnd.n1962 gnd.n1191 0.0269946
R14197 gnd.n1961 gnd.n1192 0.0269946
R14198 gnd.n1956 gnd.n1166 0.0269946
R14199 gnd.n2030 gnd.n1164 0.0269946
R14200 gnd.n2032 gnd.n2031 0.0269946
R14201 gnd.n2034 gnd.n2033 0.0269946
R14202 gnd.n2044 gnd.n1157 0.0269946
R14203 gnd.n2046 gnd.n2045 0.0269946
R14204 gnd.n2047 gnd.n996 0.0269946
R14205 gnd.n2049 gnd.n997 0.0269946
R14206 gnd.n2051 gnd.n998 0.0269946
R14207 gnd.n2057 gnd.n2056 0.0269946
R14208 gnd.n2059 gnd.n2058 0.0269946
R14209 gnd.n2060 gnd.n1022 0.0269946
R14210 gnd.n2320 gnd.n1024 0.0269946
R14211 gnd.n2326 gnd.n2325 0.0269946
R14212 gnd.n2328 gnd.n2327 0.0269946
R14213 gnd.n6336 gnd.n1047 0.0269946
R14214 gnd.n6012 gnd.n2680 0.022519
R14215 gnd.n6011 gnd.n2681 0.022519
R14216 gnd.n6008 gnd.n6007 0.022519
R14217 gnd.n6004 gnd.n2686 0.022519
R14218 gnd.n6003 gnd.n2692 0.022519
R14219 gnd.n6000 gnd.n5999 0.022519
R14220 gnd.n5996 gnd.n2696 0.022519
R14221 gnd.n5995 gnd.n2700 0.022519
R14222 gnd.n5992 gnd.n5991 0.022519
R14223 gnd.n5988 gnd.n2704 0.022519
R14224 gnd.n5987 gnd.n2710 0.022519
R14225 gnd.n5984 gnd.n5983 0.022519
R14226 gnd.n5980 gnd.n2714 0.022519
R14227 gnd.n5979 gnd.n2718 0.022519
R14228 gnd.n5976 gnd.n5975 0.022519
R14229 gnd.n5972 gnd.n2722 0.022519
R14230 gnd.n5971 gnd.n2731 0.022519
R14231 gnd.n2736 gnd.n2735 0.022519
R14232 gnd.n6035 gnd.n2645 0.022519
R14233 gnd.n5697 gnd.n3105 0.022519
R14234 gnd.n5696 gnd.n3109 0.022519
R14235 gnd.n5693 gnd.n5692 0.022519
R14236 gnd.n5689 gnd.n3114 0.022519
R14237 gnd.n5688 gnd.n3118 0.022519
R14238 gnd.n5685 gnd.n5684 0.022519
R14239 gnd.n5681 gnd.n3122 0.022519
R14240 gnd.n5680 gnd.n3126 0.022519
R14241 gnd.n5677 gnd.n5676 0.022519
R14242 gnd.n5673 gnd.n3130 0.022519
R14243 gnd.n5672 gnd.n3134 0.022519
R14244 gnd.n5669 gnd.n5668 0.022519
R14245 gnd.n5665 gnd.n3138 0.022519
R14246 gnd.n5664 gnd.n3142 0.022519
R14247 gnd.n5661 gnd.n5660 0.022519
R14248 gnd.n5657 gnd.n3146 0.022519
R14249 gnd.n5656 gnd.n3152 0.022519
R14250 gnd.n3420 gnd.n3155 0.022519
R14251 gnd.n5302 gnd.n3419 0.022519
R14252 gnd.n5303 gnd.n3418 0.0218415
R14253 gnd.n6036 gnd.n2644 0.0218415
R14254 gnd.n1743 gnd.n1742 0.0202011
R14255 gnd.n1742 gnd.n1741 0.0148637
R14256 gnd.n2318 gnd.n2317 0.0144266
R14257 gnd.n2317 gnd.n1023 0.0130679
R14258 gnd.n2680 gnd.n2674 0.0123564
R14259 gnd.n6012 gnd.n6011 0.0123564
R14260 gnd.n6008 gnd.n2681 0.0123564
R14261 gnd.n6007 gnd.n2686 0.0123564
R14262 gnd.n6004 gnd.n6003 0.0123564
R14263 gnd.n6000 gnd.n2692 0.0123564
R14264 gnd.n5999 gnd.n2696 0.0123564
R14265 gnd.n5996 gnd.n5995 0.0123564
R14266 gnd.n5992 gnd.n2700 0.0123564
R14267 gnd.n5991 gnd.n2704 0.0123564
R14268 gnd.n5988 gnd.n5987 0.0123564
R14269 gnd.n5984 gnd.n2710 0.0123564
R14270 gnd.n5983 gnd.n2714 0.0123564
R14271 gnd.n5980 gnd.n5979 0.0123564
R14272 gnd.n5976 gnd.n2718 0.0123564
R14273 gnd.n5975 gnd.n2722 0.0123564
R14274 gnd.n5972 gnd.n5971 0.0123564
R14275 gnd.n2736 gnd.n2731 0.0123564
R14276 gnd.n2735 gnd.n2645 0.0123564
R14277 gnd.n5700 gnd.n3105 0.0123564
R14278 gnd.n5697 gnd.n5696 0.0123564
R14279 gnd.n5693 gnd.n3109 0.0123564
R14280 gnd.n5692 gnd.n3114 0.0123564
R14281 gnd.n5689 gnd.n5688 0.0123564
R14282 gnd.n5685 gnd.n3118 0.0123564
R14283 gnd.n5684 gnd.n3122 0.0123564
R14284 gnd.n5681 gnd.n5680 0.0123564
R14285 gnd.n5677 gnd.n3126 0.0123564
R14286 gnd.n5676 gnd.n3130 0.0123564
R14287 gnd.n5673 gnd.n5672 0.0123564
R14288 gnd.n5669 gnd.n3134 0.0123564
R14289 gnd.n5668 gnd.n3138 0.0123564
R14290 gnd.n5665 gnd.n5664 0.0123564
R14291 gnd.n5661 gnd.n3142 0.0123564
R14292 gnd.n5660 gnd.n3146 0.0123564
R14293 gnd.n5657 gnd.n5656 0.0123564
R14294 gnd.n3155 gnd.n3152 0.0123564
R14295 gnd.n3420 gnd.n3419 0.0123564
R14296 gnd.n1744 gnd.n1364 0.00797283
R14297 gnd.n1752 gnd.n1363 0.00797283
R14298 gnd.n1754 gnd.n1753 0.00797283
R14299 gnd.n1772 gnd.n1346 0.00797283
R14300 gnd.n1774 gnd.n1773 0.00797283
R14301 gnd.n1775 gnd.n1340 0.00797283
R14302 gnd.n1783 gnd.n1338 0.00797283
R14303 gnd.n1785 gnd.n1784 0.00797283
R14304 gnd.n1803 gnd.n1319 0.00797283
R14305 gnd.n1805 gnd.n1804 0.00797283
R14306 gnd.n1806 gnd.n1314 0.00797283
R14307 gnd.n1814 gnd.n1312 0.00797283
R14308 gnd.n1816 gnd.n1815 0.00797283
R14309 gnd.n1834 gnd.n1293 0.00797283
R14310 gnd.n1836 gnd.n1835 0.00797283
R14311 gnd.n1837 gnd.n1288 0.00797283
R14312 gnd.n1845 gnd.n1286 0.00797283
R14313 gnd.n1847 gnd.n1846 0.00797283
R14314 gnd.n1865 gnd.n1268 0.00797283
R14315 gnd.n1867 gnd.n1866 0.00797283
R14316 gnd.n1868 gnd.n1262 0.00797283
R14317 gnd.n1876 gnd.n1260 0.00797283
R14318 gnd.n1878 gnd.n1877 0.00797283
R14319 gnd.n1896 gnd.n1243 0.00797283
R14320 gnd.n1898 gnd.n1897 0.00797283
R14321 gnd.n1899 gnd.n1237 0.00797283
R14322 gnd.n1907 gnd.n1235 0.00797283
R14323 gnd.n1909 gnd.n1908 0.00797283
R14324 gnd.n1927 gnd.n1218 0.00797283
R14325 gnd.n1929 gnd.n1928 0.00797283
R14326 gnd.n1930 gnd.n1212 0.00797283
R14327 gnd.n1211 gnd.n1207 0.00797283
R14328 gnd.n1940 gnd.n1939 0.00797283
R14329 gnd.n1209 gnd.n1208 0.00797283
R14330 gnd.n1191 gnd.n1190 0.00797283
R14331 gnd.n1962 gnd.n1961 0.00797283
R14332 gnd.n1956 gnd.n1192 0.00797283
R14333 gnd.n1166 gnd.n1164 0.00797283
R14334 gnd.n2031 gnd.n2030 0.00797283
R14335 gnd.n2034 gnd.n2032 0.00797283
R14336 gnd.n2033 gnd.n1157 0.00797283
R14337 gnd.n2045 gnd.n2044 0.00797283
R14338 gnd.n2047 gnd.n2046 0.00797283
R14339 gnd.n2049 gnd.n996 0.00797283
R14340 gnd.n2051 gnd.n997 0.00797283
R14341 gnd.n2056 gnd.n998 0.00797283
R14342 gnd.n2058 gnd.n2057 0.00797283
R14343 gnd.n2060 gnd.n2059 0.00797283
R14344 gnd.n2318 gnd.n1022 0.00797283
R14345 gnd.n2320 gnd.n1023 0.00797283
R14346 gnd.n2325 gnd.n1024 0.00797283
R14347 gnd.n2328 gnd.n2326 0.00797283
R14348 gnd.n2327 gnd.n1047 0.00797283
R14349 gnd.n6336 gnd.n6335 0.00797283
R14350 gnd.n6017 gnd.n6016 0.00592005
R14351 gnd.n5702 gnd.n5701 0.00592005
R14352 a_n2982_13878.n136 a_n2982_13878.t94 512.366
R14353 a_n2982_13878.n135 a_n2982_13878.t83 512.366
R14354 a_n2982_13878.n134 a_n2982_13878.t72 512.366
R14355 a_n2982_13878.n138 a_n2982_13878.t102 512.366
R14356 a_n2982_13878.n137 a_n2982_13878.t91 512.366
R14357 a_n2982_13878.n133 a_n2982_13878.t90 512.366
R14358 a_n2982_13878.n140 a_n2982_13878.t98 512.366
R14359 a_n2982_13878.n139 a_n2982_13878.t81 512.366
R14360 a_n2982_13878.n132 a_n2982_13878.t82 512.366
R14361 a_n2982_13878.n142 a_n2982_13878.t85 512.366
R14362 a_n2982_13878.n141 a_n2982_13878.t95 512.366
R14363 a_n2982_13878.n131 a_n2982_13878.t111 512.366
R14364 a_n2982_13878.n31 a_n2982_13878.t110 538.698
R14365 a_n2982_13878.n117 a_n2982_13878.t87 512.366
R14366 a_n2982_13878.n116 a_n2982_13878.t92 512.366
R14367 a_n2982_13878.n108 a_n2982_13878.t80 512.366
R14368 a_n2982_13878.n115 a_n2982_13878.t97 512.366
R14369 a_n2982_13878.n114 a_n2982_13878.t106 512.366
R14370 a_n2982_13878.n109 a_n2982_13878.t107 512.366
R14371 a_n2982_13878.n113 a_n2982_13878.t74 512.366
R14372 a_n2982_13878.n112 a_n2982_13878.t89 512.366
R14373 a_n2982_13878.n110 a_n2982_13878.t77 512.366
R14374 a_n2982_13878.n111 a_n2982_13878.t84 512.366
R14375 a_n2982_13878.n25 a_n2982_13878.t40 538.698
R14376 a_n2982_13878.n124 a_n2982_13878.t52 512.366
R14377 a_n2982_13878.n123 a_n2982_13878.t30 512.366
R14378 a_n2982_13878.n93 a_n2982_13878.t64 512.366
R14379 a_n2982_13878.n122 a_n2982_13878.t38 512.366
R14380 a_n2982_13878.n121 a_n2982_13878.t54 512.366
R14381 a_n2982_13878.n94 a_n2982_13878.t32 512.366
R14382 a_n2982_13878.n120 a_n2982_13878.t48 512.366
R14383 a_n2982_13878.n119 a_n2982_13878.t56 512.366
R14384 a_n2982_13878.n95 a_n2982_13878.t50 512.366
R14385 a_n2982_13878.n118 a_n2982_13878.t66 512.366
R14386 a_n2982_13878.n13 a_n2982_13878.t34 538.698
R14387 a_n2982_13878.n150 a_n2982_13878.t62 512.366
R14388 a_n2982_13878.n88 a_n2982_13878.t24 512.366
R14389 a_n2982_13878.n151 a_n2982_13878.t44 512.366
R14390 a_n2982_13878.n87 a_n2982_13878.t22 512.366
R14391 a_n2982_13878.n152 a_n2982_13878.t58 512.366
R14392 a_n2982_13878.n153 a_n2982_13878.t36 512.366
R14393 a_n2982_13878.n86 a_n2982_13878.t46 512.366
R14394 a_n2982_13878.n154 a_n2982_13878.t28 512.366
R14395 a_n2982_13878.n85 a_n2982_13878.t26 512.366
R14396 a_n2982_13878.n155 a_n2982_13878.t60 512.366
R14397 a_n2982_13878.n19 a_n2982_13878.t109 538.698
R14398 a_n2982_13878.n144 a_n2982_13878.t78 512.366
R14399 a_n2982_13878.n92 a_n2982_13878.t79 512.366
R14400 a_n2982_13878.n145 a_n2982_13878.t104 512.366
R14401 a_n2982_13878.n91 a_n2982_13878.t105 512.366
R14402 a_n2982_13878.n146 a_n2982_13878.t76 512.366
R14403 a_n2982_13878.n147 a_n2982_13878.t100 512.366
R14404 a_n2982_13878.n90 a_n2982_13878.t101 512.366
R14405 a_n2982_13878.n148 a_n2982_13878.t73 512.366
R14406 a_n2982_13878.n89 a_n2982_13878.t86 512.366
R14407 a_n2982_13878.n149 a_n2982_13878.t96 512.366
R14408 a_n2982_13878.n0 a_n2982_13878.n82 70.1674
R14409 a_n2982_13878.n2 a_n2982_13878.n80 70.1674
R14410 a_n2982_13878.n4 a_n2982_13878.n78 70.1674
R14411 a_n2982_13878.n6 a_n2982_13878.n76 70.1674
R14412 a_n2982_13878.n51 a_n2982_13878.n26 70.5844
R14413 a_n2982_13878.n83 a_n2982_13878.n20 70.5844
R14414 a_n2982_13878.n26 a_n2982_13878.n49 70.1674
R14415 a_n2982_13878.n49 a_n2982_13878.n110 20.9683
R14416 a_n2982_13878.n48 a_n2982_13878.n27 74.73
R14417 a_n2982_13878.n112 a_n2982_13878.n48 11.843
R14418 a_n2982_13878.n47 a_n2982_13878.n27 80.4688
R14419 a_n2982_13878.n47 a_n2982_13878.n113 0.365327
R14420 a_n2982_13878.n28 a_n2982_13878.n46 75.0448
R14421 a_n2982_13878.n45 a_n2982_13878.n28 70.1674
R14422 a_n2982_13878.n115 a_n2982_13878.n45 20.9683
R14423 a_n2982_13878.n30 a_n2982_13878.n44 70.3058
R14424 a_n2982_13878.n44 a_n2982_13878.n108 20.6913
R14425 a_n2982_13878.n43 a_n2982_13878.n30 75.3623
R14426 a_n2982_13878.n116 a_n2982_13878.n43 10.5784
R14427 a_n2982_13878.n29 a_n2982_13878.n31 44.7878
R14428 a_n2982_13878.n20 a_n2982_13878.n58 70.1674
R14429 a_n2982_13878.n58 a_n2982_13878.n95 20.9683
R14430 a_n2982_13878.n57 a_n2982_13878.n21 74.73
R14431 a_n2982_13878.n119 a_n2982_13878.n57 11.843
R14432 a_n2982_13878.n56 a_n2982_13878.n21 80.4688
R14433 a_n2982_13878.n56 a_n2982_13878.n120 0.365327
R14434 a_n2982_13878.n22 a_n2982_13878.n55 75.0448
R14435 a_n2982_13878.n54 a_n2982_13878.n22 70.1674
R14436 a_n2982_13878.n122 a_n2982_13878.n54 20.9683
R14437 a_n2982_13878.n24 a_n2982_13878.n53 70.3058
R14438 a_n2982_13878.n53 a_n2982_13878.n93 20.6913
R14439 a_n2982_13878.n52 a_n2982_13878.n24 75.3623
R14440 a_n2982_13878.n123 a_n2982_13878.n52 10.5784
R14441 a_n2982_13878.n23 a_n2982_13878.n25 44.7878
R14442 a_n2982_13878.n9 a_n2982_13878.n74 70.5844
R14443 a_n2982_13878.n15 a_n2982_13878.n66 70.5844
R14444 a_n2982_13878.n65 a_n2982_13878.n15 70.1674
R14445 a_n2982_13878.n65 a_n2982_13878.n89 20.9683
R14446 a_n2982_13878.n14 a_n2982_13878.n64 74.73
R14447 a_n2982_13878.n148 a_n2982_13878.n64 11.843
R14448 a_n2982_13878.n63 a_n2982_13878.n14 80.4688
R14449 a_n2982_13878.n63 a_n2982_13878.n90 0.365327
R14450 a_n2982_13878.n16 a_n2982_13878.n62 75.0448
R14451 a_n2982_13878.n61 a_n2982_13878.n16 70.1674
R14452 a_n2982_13878.n61 a_n2982_13878.n91 20.9683
R14453 a_n2982_13878.n17 a_n2982_13878.n60 70.3058
R14454 a_n2982_13878.n145 a_n2982_13878.n60 20.6913
R14455 a_n2982_13878.n59 a_n2982_13878.n17 75.3623
R14456 a_n2982_13878.n59 a_n2982_13878.n92 10.5784
R14457 a_n2982_13878.n19 a_n2982_13878.n18 44.7878
R14458 a_n2982_13878.n73 a_n2982_13878.n9 70.1674
R14459 a_n2982_13878.n73 a_n2982_13878.n85 20.9683
R14460 a_n2982_13878.n8 a_n2982_13878.n72 74.73
R14461 a_n2982_13878.n154 a_n2982_13878.n72 11.843
R14462 a_n2982_13878.n71 a_n2982_13878.n8 80.4688
R14463 a_n2982_13878.n71 a_n2982_13878.n86 0.365327
R14464 a_n2982_13878.n10 a_n2982_13878.n70 75.0448
R14465 a_n2982_13878.n69 a_n2982_13878.n10 70.1674
R14466 a_n2982_13878.n69 a_n2982_13878.n87 20.9683
R14467 a_n2982_13878.n11 a_n2982_13878.n68 70.3058
R14468 a_n2982_13878.n151 a_n2982_13878.n68 20.6913
R14469 a_n2982_13878.n67 a_n2982_13878.n11 75.3623
R14470 a_n2982_13878.n67 a_n2982_13878.n88 10.5784
R14471 a_n2982_13878.n13 a_n2982_13878.n12 44.7878
R14472 a_n2982_13878.n76 a_n2982_13878.n131 20.9683
R14473 a_n2982_13878.n75 a_n2982_13878.n7 75.0448
R14474 a_n2982_13878.n141 a_n2982_13878.n75 11.2134
R14475 a_n2982_13878.n7 a_n2982_13878.n142 161.3
R14476 a_n2982_13878.n78 a_n2982_13878.n132 20.9683
R14477 a_n2982_13878.n77 a_n2982_13878.n5 75.0448
R14478 a_n2982_13878.n139 a_n2982_13878.n77 11.2134
R14479 a_n2982_13878.n5 a_n2982_13878.n140 161.3
R14480 a_n2982_13878.n80 a_n2982_13878.n133 20.9683
R14481 a_n2982_13878.n79 a_n2982_13878.n3 75.0448
R14482 a_n2982_13878.n137 a_n2982_13878.n79 11.2134
R14483 a_n2982_13878.n3 a_n2982_13878.n138 161.3
R14484 a_n2982_13878.n82 a_n2982_13878.n134 20.9683
R14485 a_n2982_13878.n81 a_n2982_13878.n1 75.0448
R14486 a_n2982_13878.n135 a_n2982_13878.n81 11.2134
R14487 a_n2982_13878.n1 a_n2982_13878.n136 161.3
R14488 a_n2982_13878.n41 a_n2982_13878.n105 81.2902
R14489 a_n2982_13878.n42 a_n2982_13878.n99 81.2902
R14490 a_n2982_13878.n32 a_n2982_13878.n96 81.2902
R14491 a_n2982_13878.n41 a_n2982_13878.n106 80.9324
R14492 a_n2982_13878.n34 a_n2982_13878.n107 80.9324
R14493 a_n2982_13878.n34 a_n2982_13878.n104 80.9324
R14494 a_n2982_13878.n34 a_n2982_13878.n103 80.9324
R14495 a_n2982_13878.n33 a_n2982_13878.n102 80.9324
R14496 a_n2982_13878.n42 a_n2982_13878.n100 80.9324
R14497 a_n2982_13878.n32 a_n2982_13878.n101 80.9324
R14498 a_n2982_13878.n32 a_n2982_13878.n98 80.9324
R14499 a_n2982_13878.n32 a_n2982_13878.n97 80.9324
R14500 a_n2982_13878.n39 a_n2982_13878.t35 74.6477
R14501 a_n2982_13878.n37 a_n2982_13878.t43 74.6477
R14502 a_n2982_13878.n36 a_n2982_13878.t41 74.2899
R14503 a_n2982_13878.n40 a_n2982_13878.t69 74.2897
R14504 a_n2982_13878.n40 a_n2982_13878.n157 70.6783
R14505 a_n2982_13878.n38 a_n2982_13878.n158 70.6783
R14506 a_n2982_13878.n38 a_n2982_13878.n159 70.6783
R14507 a_n2982_13878.n39 a_n2982_13878.n84 70.6783
R14508 a_n2982_13878.n37 a_n2982_13878.n125 70.6783
R14509 a_n2982_13878.n37 a_n2982_13878.n126 70.6783
R14510 a_n2982_13878.n35 a_n2982_13878.n127 70.6783
R14511 a_n2982_13878.n35 a_n2982_13878.n128 70.6783
R14512 a_n2982_13878.n36 a_n2982_13878.n129 70.6783
R14513 a_n2982_13878.n160 a_n2982_13878.n39 70.6782
R14514 a_n2982_13878.n136 a_n2982_13878.n135 48.2005
R14515 a_n2982_13878.t99 a_n2982_13878.n82 533.335
R14516 a_n2982_13878.n138 a_n2982_13878.n137 48.2005
R14517 a_n2982_13878.t108 a_n2982_13878.n80 533.335
R14518 a_n2982_13878.n140 a_n2982_13878.n139 48.2005
R14519 a_n2982_13878.t93 a_n2982_13878.n78 533.335
R14520 a_n2982_13878.n142 a_n2982_13878.n141 48.2005
R14521 a_n2982_13878.t88 a_n2982_13878.n76 533.335
R14522 a_n2982_13878.n117 a_n2982_13878.n116 48.2005
R14523 a_n2982_13878.n45 a_n2982_13878.n114 20.9683
R14524 a_n2982_13878.n113 a_n2982_13878.n109 48.2005
R14525 a_n2982_13878.n111 a_n2982_13878.n49 20.9683
R14526 a_n2982_13878.n124 a_n2982_13878.n123 48.2005
R14527 a_n2982_13878.n54 a_n2982_13878.n121 20.9683
R14528 a_n2982_13878.n120 a_n2982_13878.n94 48.2005
R14529 a_n2982_13878.n118 a_n2982_13878.n58 20.9683
R14530 a_n2982_13878.n150 a_n2982_13878.n88 48.2005
R14531 a_n2982_13878.n152 a_n2982_13878.n69 20.9683
R14532 a_n2982_13878.n153 a_n2982_13878.n86 48.2005
R14533 a_n2982_13878.n155 a_n2982_13878.n73 20.9683
R14534 a_n2982_13878.n144 a_n2982_13878.n92 48.2005
R14535 a_n2982_13878.n146 a_n2982_13878.n61 20.9683
R14536 a_n2982_13878.n147 a_n2982_13878.n90 48.2005
R14537 a_n2982_13878.n149 a_n2982_13878.n65 20.9683
R14538 a_n2982_13878.n115 a_n2982_13878.n44 21.4216
R14539 a_n2982_13878.n122 a_n2982_13878.n53 21.4216
R14540 a_n2982_13878.n87 a_n2982_13878.n68 21.4216
R14541 a_n2982_13878.n91 a_n2982_13878.n60 21.4216
R14542 a_n2982_13878.n51 a_n2982_13878.t103 532.5
R14543 a_n2982_13878.n83 a_n2982_13878.t42 532.5
R14544 a_n2982_13878.t68 a_n2982_13878.n74 532.5
R14545 a_n2982_13878.t75 a_n2982_13878.n66 532.5
R14546 a_n2982_13878.n33 a_n2982_13878.n32 31.7747
R14547 a_n2982_13878.n48 a_n2982_13878.n110 34.4824
R14548 a_n2982_13878.n57 a_n2982_13878.n95 34.4824
R14549 a_n2982_13878.n85 a_n2982_13878.n72 34.4824
R14550 a_n2982_13878.n89 a_n2982_13878.n64 34.4824
R14551 a_n2982_13878.n81 a_n2982_13878.n134 35.3134
R14552 a_n2982_13878.n79 a_n2982_13878.n133 35.3134
R14553 a_n2982_13878.n77 a_n2982_13878.n132 35.3134
R14554 a_n2982_13878.n75 a_n2982_13878.n131 35.3134
R14555 a_n2982_13878.n114 a_n2982_13878.n46 35.3134
R14556 a_n2982_13878.n46 a_n2982_13878.n109 11.2134
R14557 a_n2982_13878.n121 a_n2982_13878.n55 35.3134
R14558 a_n2982_13878.n55 a_n2982_13878.n94 11.2134
R14559 a_n2982_13878.n70 a_n2982_13878.n152 35.3134
R14560 a_n2982_13878.n153 a_n2982_13878.n70 11.2134
R14561 a_n2982_13878.n62 a_n2982_13878.n146 35.3134
R14562 a_n2982_13878.n147 a_n2982_13878.n62 11.2134
R14563 a_n2982_13878.n20 a_n2982_13878.n34 23.891
R14564 a_n2982_13878.n43 a_n2982_13878.n108 36.139
R14565 a_n2982_13878.n52 a_n2982_13878.n93 36.139
R14566 a_n2982_13878.n151 a_n2982_13878.n67 36.139
R14567 a_n2982_13878.n145 a_n2982_13878.n59 36.139
R14568 a_n2982_13878.n18 a_n2982_13878.n143 13.9285
R14569 a_n2982_13878.n26 a_n2982_13878.n50 13.724
R14570 a_n2982_13878.n130 a_n2982_13878.n23 12.4191
R14571 a_n2982_13878.n143 a_n2982_13878.n7 11.2486
R14572 a_n2982_13878.n0 a_n2982_13878.n50 11.2486
R14573 a_n2982_13878.n40 a_n2982_13878.n156 10.5745
R14574 a_n2982_13878.n156 a_n2982_13878.n9 8.58383
R14575 a_n2982_13878.n130 a_n2982_13878.n36 6.7311
R14576 a_n2982_13878.n156 a_n2982_13878.n50 5.3452
R14577 a_n2982_13878.n20 a_n2982_13878.n29 3.94368
R14578 a_n2982_13878.n12 a_n2982_13878.n15 3.94368
R14579 a_n2982_13878.n157 a_n2982_13878.t27 3.61217
R14580 a_n2982_13878.n157 a_n2982_13878.t61 3.61217
R14581 a_n2982_13878.n158 a_n2982_13878.t47 3.61217
R14582 a_n2982_13878.n158 a_n2982_13878.t29 3.61217
R14583 a_n2982_13878.n159 a_n2982_13878.t59 3.61217
R14584 a_n2982_13878.n159 a_n2982_13878.t37 3.61217
R14585 a_n2982_13878.n84 a_n2982_13878.t63 3.61217
R14586 a_n2982_13878.n84 a_n2982_13878.t25 3.61217
R14587 a_n2982_13878.n125 a_n2982_13878.t51 3.61217
R14588 a_n2982_13878.n125 a_n2982_13878.t67 3.61217
R14589 a_n2982_13878.n126 a_n2982_13878.t49 3.61217
R14590 a_n2982_13878.n126 a_n2982_13878.t57 3.61217
R14591 a_n2982_13878.n127 a_n2982_13878.t55 3.61217
R14592 a_n2982_13878.n127 a_n2982_13878.t33 3.61217
R14593 a_n2982_13878.n128 a_n2982_13878.t65 3.61217
R14594 a_n2982_13878.n128 a_n2982_13878.t39 3.61217
R14595 a_n2982_13878.n129 a_n2982_13878.t53 3.61217
R14596 a_n2982_13878.n129 a_n2982_13878.t31 3.61217
R14597 a_n2982_13878.n160 a_n2982_13878.t45 3.61217
R14598 a_n2982_13878.t23 a_n2982_13878.n160 3.61217
R14599 a_n2982_13878.n105 a_n2982_13878.t20 2.82907
R14600 a_n2982_13878.n105 a_n2982_13878.t10 2.82907
R14601 a_n2982_13878.n106 a_n2982_13878.t8 2.82907
R14602 a_n2982_13878.n106 a_n2982_13878.t14 2.82907
R14603 a_n2982_13878.n107 a_n2982_13878.t4 2.82907
R14604 a_n2982_13878.n107 a_n2982_13878.t71 2.82907
R14605 a_n2982_13878.n104 a_n2982_13878.t19 2.82907
R14606 a_n2982_13878.n104 a_n2982_13878.t7 2.82907
R14607 a_n2982_13878.n103 a_n2982_13878.t0 2.82907
R14608 a_n2982_13878.n103 a_n2982_13878.t21 2.82907
R14609 a_n2982_13878.n102 a_n2982_13878.t13 2.82907
R14610 a_n2982_13878.n102 a_n2982_13878.t70 2.82907
R14611 a_n2982_13878.n99 a_n2982_13878.t1 2.82907
R14612 a_n2982_13878.n99 a_n2982_13878.t18 2.82907
R14613 a_n2982_13878.n100 a_n2982_13878.t2 2.82907
R14614 a_n2982_13878.n100 a_n2982_13878.t12 2.82907
R14615 a_n2982_13878.n101 a_n2982_13878.t6 2.82907
R14616 a_n2982_13878.n101 a_n2982_13878.t5 2.82907
R14617 a_n2982_13878.n98 a_n2982_13878.t16 2.82907
R14618 a_n2982_13878.n98 a_n2982_13878.t15 2.82907
R14619 a_n2982_13878.n97 a_n2982_13878.t3 2.82907
R14620 a_n2982_13878.n97 a_n2982_13878.t11 2.82907
R14621 a_n2982_13878.n96 a_n2982_13878.t17 2.82907
R14622 a_n2982_13878.n96 a_n2982_13878.t9 2.82907
R14623 a_n2982_13878.n31 a_n2982_13878.n117 14.1668
R14624 a_n2982_13878.n111 a_n2982_13878.n51 22.3251
R14625 a_n2982_13878.n25 a_n2982_13878.n124 14.1668
R14626 a_n2982_13878.n118 a_n2982_13878.n83 22.3251
R14627 a_n2982_13878.n150 a_n2982_13878.n13 14.1668
R14628 a_n2982_13878.n74 a_n2982_13878.n155 22.3251
R14629 a_n2982_13878.n144 a_n2982_13878.n19 14.1668
R14630 a_n2982_13878.n66 a_n2982_13878.n149 22.3251
R14631 a_n2982_13878.n143 a_n2982_13878.n130 1.30542
R14632 a_n2982_13878.n4 a_n2982_13878.n3 1.04595
R14633 a_n2982_13878.n47 a_n2982_13878.n112 47.835
R14634 a_n2982_13878.n56 a_n2982_13878.n119 47.835
R14635 a_n2982_13878.n154 a_n2982_13878.n71 47.835
R14636 a_n2982_13878.n148 a_n2982_13878.n63 47.835
R14637 a_n2982_13878.n27 a_n2982_13878.n26 1.13686
R14638 a_n2982_13878.n15 a_n2982_13878.n14 1.13686
R14639 a_n2982_13878.n9 a_n2982_13878.n8 1.13686
R14640 a_n2982_13878.n21 a_n2982_13878.n20 1.09898
R14641 a_n2982_13878.n39 a_n2982_13878.n38 1.07378
R14642 a_n2982_13878.n36 a_n2982_13878.n35 1.07378
R14643 a_n2982_13878.n32 a_n2982_13878.n42 1.07378
R14644 a_n2982_13878.n30 a_n2982_13878.n29 0.758076
R14645 a_n2982_13878.n30 a_n2982_13878.n28 0.758076
R14646 a_n2982_13878.n28 a_n2982_13878.n27 0.758076
R14647 a_n2982_13878.n24 a_n2982_13878.n23 0.758076
R14648 a_n2982_13878.n24 a_n2982_13878.n22 0.758076
R14649 a_n2982_13878.n22 a_n2982_13878.n21 0.758076
R14650 a_n2982_13878.n17 a_n2982_13878.n18 0.758076
R14651 a_n2982_13878.n16 a_n2982_13878.n17 0.758076
R14652 a_n2982_13878.n14 a_n2982_13878.n16 0.758076
R14653 a_n2982_13878.n11 a_n2982_13878.n12 0.758076
R14654 a_n2982_13878.n10 a_n2982_13878.n11 0.758076
R14655 a_n2982_13878.n8 a_n2982_13878.n10 0.758076
R14656 a_n2982_13878.n7 a_n2982_13878.n6 0.758076
R14657 a_n2982_13878.n5 a_n2982_13878.n4 0.758076
R14658 a_n2982_13878.n3 a_n2982_13878.n2 0.758076
R14659 a_n2982_13878.n1 a_n2982_13878.n0 0.758076
R14660 a_n2982_13878.n34 a_n2982_13878.n41 0.716017
R14661 a_n2982_13878.n38 a_n2982_13878.n40 0.716017
R14662 a_n2982_13878.n35 a_n2982_13878.n37 0.716017
R14663 a_n2982_13878.n34 a_n2982_13878.n33 0.716017
R14664 a_n2982_13878.n6 a_n2982_13878.n5 0.67853
R14665 a_n2982_13878.n2 a_n2982_13878.n1 0.67853
R14666 vdd.n303 vdd.n267 756.745
R14667 vdd.n252 vdd.n216 756.745
R14668 vdd.n209 vdd.n173 756.745
R14669 vdd.n158 vdd.n122 756.745
R14670 vdd.n116 vdd.n80 756.745
R14671 vdd.n65 vdd.n29 756.745
R14672 vdd.n1953 vdd.n1917 756.745
R14673 vdd.n2004 vdd.n1968 756.745
R14674 vdd.n1859 vdd.n1823 756.745
R14675 vdd.n1910 vdd.n1874 756.745
R14676 vdd.n1766 vdd.n1730 756.745
R14677 vdd.n1817 vdd.n1781 756.745
R14678 vdd.n1143 vdd.t14 640.208
R14679 vdd.n838 vdd.t59 640.208
R14680 vdd.n1147 vdd.t56 640.208
R14681 vdd.n829 vdd.t83 640.208
R14682 vdd.n724 vdd.t36 640.208
R14683 vdd.n2535 vdd.t77 640.208
R14684 vdd.n661 vdd.t25 640.208
R14685 vdd.n2532 vdd.t66 640.208
R14686 vdd.n625 vdd.t10 640.208
R14687 vdd.n899 vdd.t73 640.208
R14688 vdd.n1565 vdd.t46 592.009
R14689 vdd.n1602 vdd.t70 592.009
R14690 vdd.n1476 vdd.t80 592.009
R14691 vdd.n2074 vdd.t40 592.009
R14692 vdd.n1076 vdd.t18 592.009
R14693 vdd.n1036 vdd.t22 592.009
R14694 vdd.n3293 vdd.t43 592.009
R14695 vdd.n427 vdd.t32 592.009
R14696 vdd.n387 vdd.t50 592.009
R14697 vdd.n580 vdd.t53 592.009
R14698 vdd.n543 vdd.t63 592.009
R14699 vdd.n3080 vdd.t28 592.009
R14700 vdd.n304 vdd.n303 585
R14701 vdd.n302 vdd.n269 585
R14702 vdd.n301 vdd.n300 585
R14703 vdd.n272 vdd.n270 585
R14704 vdd.n295 vdd.n294 585
R14705 vdd.n293 vdd.n292 585
R14706 vdd.n276 vdd.n275 585
R14707 vdd.n287 vdd.n286 585
R14708 vdd.n285 vdd.n284 585
R14709 vdd.n280 vdd.n279 585
R14710 vdd.n253 vdd.n252 585
R14711 vdd.n251 vdd.n218 585
R14712 vdd.n250 vdd.n249 585
R14713 vdd.n221 vdd.n219 585
R14714 vdd.n244 vdd.n243 585
R14715 vdd.n242 vdd.n241 585
R14716 vdd.n225 vdd.n224 585
R14717 vdd.n236 vdd.n235 585
R14718 vdd.n234 vdd.n233 585
R14719 vdd.n229 vdd.n228 585
R14720 vdd.n210 vdd.n209 585
R14721 vdd.n208 vdd.n175 585
R14722 vdd.n207 vdd.n206 585
R14723 vdd.n178 vdd.n176 585
R14724 vdd.n201 vdd.n200 585
R14725 vdd.n199 vdd.n198 585
R14726 vdd.n182 vdd.n181 585
R14727 vdd.n193 vdd.n192 585
R14728 vdd.n191 vdd.n190 585
R14729 vdd.n186 vdd.n185 585
R14730 vdd.n159 vdd.n158 585
R14731 vdd.n157 vdd.n124 585
R14732 vdd.n156 vdd.n155 585
R14733 vdd.n127 vdd.n125 585
R14734 vdd.n150 vdd.n149 585
R14735 vdd.n148 vdd.n147 585
R14736 vdd.n131 vdd.n130 585
R14737 vdd.n142 vdd.n141 585
R14738 vdd.n140 vdd.n139 585
R14739 vdd.n135 vdd.n134 585
R14740 vdd.n117 vdd.n116 585
R14741 vdd.n115 vdd.n82 585
R14742 vdd.n114 vdd.n113 585
R14743 vdd.n85 vdd.n83 585
R14744 vdd.n108 vdd.n107 585
R14745 vdd.n106 vdd.n105 585
R14746 vdd.n89 vdd.n88 585
R14747 vdd.n100 vdd.n99 585
R14748 vdd.n98 vdd.n97 585
R14749 vdd.n93 vdd.n92 585
R14750 vdd.n66 vdd.n65 585
R14751 vdd.n64 vdd.n31 585
R14752 vdd.n63 vdd.n62 585
R14753 vdd.n34 vdd.n32 585
R14754 vdd.n57 vdd.n56 585
R14755 vdd.n55 vdd.n54 585
R14756 vdd.n38 vdd.n37 585
R14757 vdd.n49 vdd.n48 585
R14758 vdd.n47 vdd.n46 585
R14759 vdd.n42 vdd.n41 585
R14760 vdd.n1954 vdd.n1953 585
R14761 vdd.n1952 vdd.n1919 585
R14762 vdd.n1951 vdd.n1950 585
R14763 vdd.n1922 vdd.n1920 585
R14764 vdd.n1945 vdd.n1944 585
R14765 vdd.n1943 vdd.n1942 585
R14766 vdd.n1926 vdd.n1925 585
R14767 vdd.n1937 vdd.n1936 585
R14768 vdd.n1935 vdd.n1934 585
R14769 vdd.n1930 vdd.n1929 585
R14770 vdd.n2005 vdd.n2004 585
R14771 vdd.n2003 vdd.n1970 585
R14772 vdd.n2002 vdd.n2001 585
R14773 vdd.n1973 vdd.n1971 585
R14774 vdd.n1996 vdd.n1995 585
R14775 vdd.n1994 vdd.n1993 585
R14776 vdd.n1977 vdd.n1976 585
R14777 vdd.n1988 vdd.n1987 585
R14778 vdd.n1986 vdd.n1985 585
R14779 vdd.n1981 vdd.n1980 585
R14780 vdd.n1860 vdd.n1859 585
R14781 vdd.n1858 vdd.n1825 585
R14782 vdd.n1857 vdd.n1856 585
R14783 vdd.n1828 vdd.n1826 585
R14784 vdd.n1851 vdd.n1850 585
R14785 vdd.n1849 vdd.n1848 585
R14786 vdd.n1832 vdd.n1831 585
R14787 vdd.n1843 vdd.n1842 585
R14788 vdd.n1841 vdd.n1840 585
R14789 vdd.n1836 vdd.n1835 585
R14790 vdd.n1911 vdd.n1910 585
R14791 vdd.n1909 vdd.n1876 585
R14792 vdd.n1908 vdd.n1907 585
R14793 vdd.n1879 vdd.n1877 585
R14794 vdd.n1902 vdd.n1901 585
R14795 vdd.n1900 vdd.n1899 585
R14796 vdd.n1883 vdd.n1882 585
R14797 vdd.n1894 vdd.n1893 585
R14798 vdd.n1892 vdd.n1891 585
R14799 vdd.n1887 vdd.n1886 585
R14800 vdd.n1767 vdd.n1766 585
R14801 vdd.n1765 vdd.n1732 585
R14802 vdd.n1764 vdd.n1763 585
R14803 vdd.n1735 vdd.n1733 585
R14804 vdd.n1758 vdd.n1757 585
R14805 vdd.n1756 vdd.n1755 585
R14806 vdd.n1739 vdd.n1738 585
R14807 vdd.n1750 vdd.n1749 585
R14808 vdd.n1748 vdd.n1747 585
R14809 vdd.n1743 vdd.n1742 585
R14810 vdd.n1818 vdd.n1817 585
R14811 vdd.n1816 vdd.n1783 585
R14812 vdd.n1815 vdd.n1814 585
R14813 vdd.n1786 vdd.n1784 585
R14814 vdd.n1809 vdd.n1808 585
R14815 vdd.n1807 vdd.n1806 585
R14816 vdd.n1790 vdd.n1789 585
R14817 vdd.n1801 vdd.n1800 585
R14818 vdd.n1799 vdd.n1798 585
R14819 vdd.n1794 vdd.n1793 585
R14820 vdd.n3409 vdd.n352 488.781
R14821 vdd.n3291 vdd.n350 488.781
R14822 vdd.n3213 vdd.n515 488.781
R14823 vdd.n3211 vdd.n517 488.781
R14824 vdd.n2069 vdd.n1358 488.781
R14825 vdd.n2072 vdd.n2071 488.781
R14826 vdd.n1671 vdd.n1436 488.781
R14827 vdd.n1669 vdd.n1439 488.781
R14828 vdd.n281 vdd.t156 329.043
R14829 vdd.n230 vdd.t238 329.043
R14830 vdd.n187 vdd.t145 329.043
R14831 vdd.n136 vdd.t114 329.043
R14832 vdd.n94 vdd.t118 329.043
R14833 vdd.n43 vdd.t5 329.043
R14834 vdd.n1931 vdd.t234 329.043
R14835 vdd.n1982 vdd.t147 329.043
R14836 vdd.n1837 vdd.t133 329.043
R14837 vdd.n1888 vdd.t116 329.043
R14838 vdd.n1744 vdd.t3 329.043
R14839 vdd.n1795 vdd.t123 329.043
R14840 vdd.n1565 vdd.t49 319.788
R14841 vdd.n1602 vdd.t72 319.788
R14842 vdd.n1476 vdd.t82 319.788
R14843 vdd.n2074 vdd.t41 319.788
R14844 vdd.n1076 vdd.t20 319.788
R14845 vdd.n1036 vdd.t23 319.788
R14846 vdd.n3293 vdd.t44 319.788
R14847 vdd.n427 vdd.t34 319.788
R14848 vdd.n387 vdd.t51 319.788
R14849 vdd.n580 vdd.t55 319.788
R14850 vdd.n543 vdd.t65 319.788
R14851 vdd.n3080 vdd.t31 319.788
R14852 vdd.n1566 vdd.t48 303.69
R14853 vdd.n1603 vdd.t71 303.69
R14854 vdd.n1477 vdd.t81 303.69
R14855 vdd.n2075 vdd.t42 303.69
R14856 vdd.n1077 vdd.t21 303.69
R14857 vdd.n1037 vdd.t24 303.69
R14858 vdd.n3294 vdd.t45 303.69
R14859 vdd.n428 vdd.t35 303.69
R14860 vdd.n388 vdd.t52 303.69
R14861 vdd.n581 vdd.t54 303.69
R14862 vdd.n544 vdd.t64 303.69
R14863 vdd.n3081 vdd.t30 303.69
R14864 vdd.n2802 vdd.n788 279.512
R14865 vdd.n3042 vdd.n635 279.512
R14866 vdd.n2979 vdd.n632 279.512
R14867 vdd.n2734 vdd.n2733 279.512
R14868 vdd.n2495 vdd.n826 279.512
R14869 vdd.n2426 vdd.n2425 279.512
R14870 vdd.n1183 vdd.n1182 279.512
R14871 vdd.n2220 vdd.n966 279.512
R14872 vdd.n2958 vdd.n633 279.512
R14873 vdd.n3045 vdd.n3044 279.512
R14874 vdd.n2607 vdd.n2530 279.512
R14875 vdd.n2538 vdd.n784 279.512
R14876 vdd.n2423 vdd.n836 279.512
R14877 vdd.n834 vdd.n808 279.512
R14878 vdd.n1308 vdd.n1003 279.512
R14879 vdd.n1108 vdd.n961 279.512
R14880 vdd.n2218 vdd.n969 254.619
R14881 vdd.n613 vdd.n516 254.619
R14882 vdd.n2960 vdd.n633 185
R14883 vdd.n3043 vdd.n633 185
R14884 vdd.n2962 vdd.n2961 185
R14885 vdd.n2961 vdd.n631 185
R14886 vdd.n2963 vdd.n667 185
R14887 vdd.n2973 vdd.n667 185
R14888 vdd.n2964 vdd.n676 185
R14889 vdd.n676 vdd.n674 185
R14890 vdd.n2966 vdd.n2965 185
R14891 vdd.n2967 vdd.n2966 185
R14892 vdd.n2919 vdd.n675 185
R14893 vdd.n675 vdd.n671 185
R14894 vdd.n2918 vdd.n2917 185
R14895 vdd.n2917 vdd.n2916 185
R14896 vdd.n678 vdd.n677 185
R14897 vdd.n679 vdd.n678 185
R14898 vdd.n2909 vdd.n2908 185
R14899 vdd.n2910 vdd.n2909 185
R14900 vdd.n2907 vdd.n687 185
R14901 vdd.n692 vdd.n687 185
R14902 vdd.n2906 vdd.n2905 185
R14903 vdd.n2905 vdd.n2904 185
R14904 vdd.n689 vdd.n688 185
R14905 vdd.n698 vdd.n689 185
R14906 vdd.n2897 vdd.n2896 185
R14907 vdd.n2898 vdd.n2897 185
R14908 vdd.n2895 vdd.n699 185
R14909 vdd.n705 vdd.n699 185
R14910 vdd.n2894 vdd.n2893 185
R14911 vdd.n2893 vdd.n2892 185
R14912 vdd.n701 vdd.n700 185
R14913 vdd.n702 vdd.n701 185
R14914 vdd.n2885 vdd.n2884 185
R14915 vdd.n2886 vdd.n2885 185
R14916 vdd.n2883 vdd.n712 185
R14917 vdd.n712 vdd.n709 185
R14918 vdd.n2882 vdd.n2881 185
R14919 vdd.n2881 vdd.n2880 185
R14920 vdd.n714 vdd.n713 185
R14921 vdd.n715 vdd.n714 185
R14922 vdd.n2873 vdd.n2872 185
R14923 vdd.n2874 vdd.n2873 185
R14924 vdd.n2871 vdd.n723 185
R14925 vdd.n729 vdd.n723 185
R14926 vdd.n2870 vdd.n2869 185
R14927 vdd.n2869 vdd.n2868 185
R14928 vdd.n2859 vdd.n726 185
R14929 vdd.n736 vdd.n726 185
R14930 vdd.n2861 vdd.n2860 185
R14931 vdd.n2862 vdd.n2861 185
R14932 vdd.n2858 vdd.n737 185
R14933 vdd.n737 vdd.n733 185
R14934 vdd.n2857 vdd.n2856 185
R14935 vdd.n2856 vdd.n2855 185
R14936 vdd.n739 vdd.n738 185
R14937 vdd.n740 vdd.n739 185
R14938 vdd.n2848 vdd.n2847 185
R14939 vdd.n2849 vdd.n2848 185
R14940 vdd.n2846 vdd.n748 185
R14941 vdd.n753 vdd.n748 185
R14942 vdd.n2845 vdd.n2844 185
R14943 vdd.n2844 vdd.n2843 185
R14944 vdd.n750 vdd.n749 185
R14945 vdd.n759 vdd.n750 185
R14946 vdd.n2836 vdd.n2835 185
R14947 vdd.n2837 vdd.n2836 185
R14948 vdd.n2834 vdd.n760 185
R14949 vdd.n2710 vdd.n760 185
R14950 vdd.n2833 vdd.n2832 185
R14951 vdd.n2832 vdd.n2831 185
R14952 vdd.n762 vdd.n761 185
R14953 vdd.n2716 vdd.n762 185
R14954 vdd.n2824 vdd.n2823 185
R14955 vdd.n2825 vdd.n2824 185
R14956 vdd.n2822 vdd.n771 185
R14957 vdd.n771 vdd.n768 185
R14958 vdd.n2821 vdd.n2820 185
R14959 vdd.n2820 vdd.n2819 185
R14960 vdd.n773 vdd.n772 185
R14961 vdd.n774 vdd.n773 185
R14962 vdd.n2812 vdd.n2811 185
R14963 vdd.n2813 vdd.n2812 185
R14964 vdd.n2810 vdd.n782 185
R14965 vdd.n2728 vdd.n782 185
R14966 vdd.n2809 vdd.n2808 185
R14967 vdd.n2808 vdd.n2807 185
R14968 vdd.n784 vdd.n783 185
R14969 vdd.n785 vdd.n784 185
R14970 vdd.n2539 vdd.n2538 185
R14971 vdd.n2541 vdd.n2540 185
R14972 vdd.n2543 vdd.n2542 185
R14973 vdd.n2545 vdd.n2544 185
R14974 vdd.n2547 vdd.n2546 185
R14975 vdd.n2549 vdd.n2548 185
R14976 vdd.n2551 vdd.n2550 185
R14977 vdd.n2553 vdd.n2552 185
R14978 vdd.n2555 vdd.n2554 185
R14979 vdd.n2557 vdd.n2556 185
R14980 vdd.n2559 vdd.n2558 185
R14981 vdd.n2561 vdd.n2560 185
R14982 vdd.n2563 vdd.n2562 185
R14983 vdd.n2565 vdd.n2564 185
R14984 vdd.n2567 vdd.n2566 185
R14985 vdd.n2569 vdd.n2568 185
R14986 vdd.n2571 vdd.n2570 185
R14987 vdd.n2573 vdd.n2572 185
R14988 vdd.n2575 vdd.n2574 185
R14989 vdd.n2577 vdd.n2576 185
R14990 vdd.n2579 vdd.n2578 185
R14991 vdd.n2581 vdd.n2580 185
R14992 vdd.n2583 vdd.n2582 185
R14993 vdd.n2585 vdd.n2584 185
R14994 vdd.n2587 vdd.n2586 185
R14995 vdd.n2589 vdd.n2588 185
R14996 vdd.n2591 vdd.n2590 185
R14997 vdd.n2593 vdd.n2592 185
R14998 vdd.n2595 vdd.n2594 185
R14999 vdd.n2597 vdd.n2596 185
R15000 vdd.n2599 vdd.n2598 185
R15001 vdd.n2601 vdd.n2600 185
R15002 vdd.n2603 vdd.n2602 185
R15003 vdd.n2605 vdd.n2604 185
R15004 vdd.n2606 vdd.n2530 185
R15005 vdd.n2800 vdd.n2530 185
R15006 vdd.n3046 vdd.n3045 185
R15007 vdd.n3047 vdd.n624 185
R15008 vdd.n3049 vdd.n3048 185
R15009 vdd.n3051 vdd.n622 185
R15010 vdd.n3053 vdd.n3052 185
R15011 vdd.n3054 vdd.n621 185
R15012 vdd.n3056 vdd.n3055 185
R15013 vdd.n3058 vdd.n619 185
R15014 vdd.n3060 vdd.n3059 185
R15015 vdd.n3061 vdd.n618 185
R15016 vdd.n3063 vdd.n3062 185
R15017 vdd.n3065 vdd.n616 185
R15018 vdd.n3067 vdd.n3066 185
R15019 vdd.n3068 vdd.n615 185
R15020 vdd.n3070 vdd.n3069 185
R15021 vdd.n3072 vdd.n614 185
R15022 vdd.n3073 vdd.n611 185
R15023 vdd.n3076 vdd.n3075 185
R15024 vdd.n612 vdd.n610 185
R15025 vdd.n2932 vdd.n2931 185
R15026 vdd.n2934 vdd.n2933 185
R15027 vdd.n2936 vdd.n2928 185
R15028 vdd.n2938 vdd.n2937 185
R15029 vdd.n2939 vdd.n2927 185
R15030 vdd.n2941 vdd.n2940 185
R15031 vdd.n2943 vdd.n2925 185
R15032 vdd.n2945 vdd.n2944 185
R15033 vdd.n2946 vdd.n2924 185
R15034 vdd.n2948 vdd.n2947 185
R15035 vdd.n2950 vdd.n2922 185
R15036 vdd.n2952 vdd.n2951 185
R15037 vdd.n2953 vdd.n2921 185
R15038 vdd.n2955 vdd.n2954 185
R15039 vdd.n2957 vdd.n2920 185
R15040 vdd.n2959 vdd.n2958 185
R15041 vdd.n2958 vdd.n613 185
R15042 vdd.n3044 vdd.n628 185
R15043 vdd.n3044 vdd.n3043 185
R15044 vdd.n2661 vdd.n630 185
R15045 vdd.n631 vdd.n630 185
R15046 vdd.n2662 vdd.n666 185
R15047 vdd.n2973 vdd.n666 185
R15048 vdd.n2664 vdd.n2663 185
R15049 vdd.n2663 vdd.n674 185
R15050 vdd.n2665 vdd.n673 185
R15051 vdd.n2967 vdd.n673 185
R15052 vdd.n2667 vdd.n2666 185
R15053 vdd.n2666 vdd.n671 185
R15054 vdd.n2668 vdd.n681 185
R15055 vdd.n2916 vdd.n681 185
R15056 vdd.n2670 vdd.n2669 185
R15057 vdd.n2669 vdd.n679 185
R15058 vdd.n2671 vdd.n686 185
R15059 vdd.n2910 vdd.n686 185
R15060 vdd.n2673 vdd.n2672 185
R15061 vdd.n2672 vdd.n692 185
R15062 vdd.n2674 vdd.n691 185
R15063 vdd.n2904 vdd.n691 185
R15064 vdd.n2676 vdd.n2675 185
R15065 vdd.n2675 vdd.n698 185
R15066 vdd.n2677 vdd.n697 185
R15067 vdd.n2898 vdd.n697 185
R15068 vdd.n2679 vdd.n2678 185
R15069 vdd.n2678 vdd.n705 185
R15070 vdd.n2680 vdd.n704 185
R15071 vdd.n2892 vdd.n704 185
R15072 vdd.n2682 vdd.n2681 185
R15073 vdd.n2681 vdd.n702 185
R15074 vdd.n2683 vdd.n711 185
R15075 vdd.n2886 vdd.n711 185
R15076 vdd.n2685 vdd.n2684 185
R15077 vdd.n2684 vdd.n709 185
R15078 vdd.n2686 vdd.n717 185
R15079 vdd.n2880 vdd.n717 185
R15080 vdd.n2688 vdd.n2687 185
R15081 vdd.n2687 vdd.n715 185
R15082 vdd.n2689 vdd.n722 185
R15083 vdd.n2874 vdd.n722 185
R15084 vdd.n2691 vdd.n2690 185
R15085 vdd.n2690 vdd.n729 185
R15086 vdd.n2692 vdd.n728 185
R15087 vdd.n2868 vdd.n728 185
R15088 vdd.n2694 vdd.n2693 185
R15089 vdd.n2693 vdd.n736 185
R15090 vdd.n2695 vdd.n735 185
R15091 vdd.n2862 vdd.n735 185
R15092 vdd.n2697 vdd.n2696 185
R15093 vdd.n2696 vdd.n733 185
R15094 vdd.n2698 vdd.n742 185
R15095 vdd.n2855 vdd.n742 185
R15096 vdd.n2700 vdd.n2699 185
R15097 vdd.n2699 vdd.n740 185
R15098 vdd.n2701 vdd.n747 185
R15099 vdd.n2849 vdd.n747 185
R15100 vdd.n2703 vdd.n2702 185
R15101 vdd.n2702 vdd.n753 185
R15102 vdd.n2704 vdd.n752 185
R15103 vdd.n2843 vdd.n752 185
R15104 vdd.n2706 vdd.n2705 185
R15105 vdd.n2705 vdd.n759 185
R15106 vdd.n2707 vdd.n758 185
R15107 vdd.n2837 vdd.n758 185
R15108 vdd.n2709 vdd.n2708 185
R15109 vdd.n2710 vdd.n2709 185
R15110 vdd.n2610 vdd.n764 185
R15111 vdd.n2831 vdd.n764 185
R15112 vdd.n2718 vdd.n2717 185
R15113 vdd.n2717 vdd.n2716 185
R15114 vdd.n2719 vdd.n770 185
R15115 vdd.n2825 vdd.n770 185
R15116 vdd.n2721 vdd.n2720 185
R15117 vdd.n2720 vdd.n768 185
R15118 vdd.n2722 vdd.n776 185
R15119 vdd.n2819 vdd.n776 185
R15120 vdd.n2724 vdd.n2723 185
R15121 vdd.n2723 vdd.n774 185
R15122 vdd.n2725 vdd.n781 185
R15123 vdd.n2813 vdd.n781 185
R15124 vdd.n2727 vdd.n2726 185
R15125 vdd.n2728 vdd.n2727 185
R15126 vdd.n2609 vdd.n787 185
R15127 vdd.n2807 vdd.n787 185
R15128 vdd.n2608 vdd.n2607 185
R15129 vdd.n2607 vdd.n785 185
R15130 vdd.n2069 vdd.n2068 185
R15131 vdd.n2070 vdd.n2069 185
R15132 vdd.n1359 vdd.n1357 185
R15133 vdd.n2061 vdd.n1357 185
R15134 vdd.n2064 vdd.n2063 185
R15135 vdd.n2063 vdd.n2062 185
R15136 vdd.n1362 vdd.n1361 185
R15137 vdd.n1363 vdd.n1362 185
R15138 vdd.n2050 vdd.n2049 185
R15139 vdd.n2051 vdd.n2050 185
R15140 vdd.n1371 vdd.n1370 185
R15141 vdd.n2042 vdd.n1370 185
R15142 vdd.n2045 vdd.n2044 185
R15143 vdd.n2044 vdd.n2043 185
R15144 vdd.n1374 vdd.n1373 185
R15145 vdd.n1380 vdd.n1374 185
R15146 vdd.n2033 vdd.n2032 185
R15147 vdd.n2034 vdd.n2033 185
R15148 vdd.n1382 vdd.n1381 185
R15149 vdd.n2025 vdd.n1381 185
R15150 vdd.n2028 vdd.n2027 185
R15151 vdd.n2027 vdd.n2026 185
R15152 vdd.n1385 vdd.n1384 185
R15153 vdd.n1386 vdd.n1385 185
R15154 vdd.n2016 vdd.n2015 185
R15155 vdd.n2017 vdd.n2016 185
R15156 vdd.n1394 vdd.n1393 185
R15157 vdd.n1393 vdd.n1392 185
R15158 vdd.n1729 vdd.n1728 185
R15159 vdd.n1728 vdd.n1727 185
R15160 vdd.n1397 vdd.n1396 185
R15161 vdd.n1403 vdd.n1397 185
R15162 vdd.n1718 vdd.n1717 185
R15163 vdd.n1719 vdd.n1718 185
R15164 vdd.n1405 vdd.n1404 185
R15165 vdd.n1710 vdd.n1404 185
R15166 vdd.n1713 vdd.n1712 185
R15167 vdd.n1712 vdd.n1711 185
R15168 vdd.n1408 vdd.n1407 185
R15169 vdd.n1415 vdd.n1408 185
R15170 vdd.n1701 vdd.n1700 185
R15171 vdd.n1702 vdd.n1701 185
R15172 vdd.n1417 vdd.n1416 185
R15173 vdd.n1416 vdd.n1414 185
R15174 vdd.n1696 vdd.n1695 185
R15175 vdd.n1695 vdd.n1694 185
R15176 vdd.n1420 vdd.n1419 185
R15177 vdd.n1421 vdd.n1420 185
R15178 vdd.n1685 vdd.n1684 185
R15179 vdd.n1686 vdd.n1685 185
R15180 vdd.n1429 vdd.n1428 185
R15181 vdd.n1428 vdd.n1427 185
R15182 vdd.n1680 vdd.n1679 185
R15183 vdd.n1679 vdd.n1678 185
R15184 vdd.n1432 vdd.n1431 185
R15185 vdd.n1438 vdd.n1432 185
R15186 vdd.n1669 vdd.n1668 185
R15187 vdd.n1670 vdd.n1669 185
R15188 vdd.n1665 vdd.n1439 185
R15189 vdd.n1664 vdd.n1442 185
R15190 vdd.n1663 vdd.n1443 185
R15191 vdd.n1443 vdd.n1437 185
R15192 vdd.n1446 vdd.n1444 185
R15193 vdd.n1659 vdd.n1448 185
R15194 vdd.n1658 vdd.n1449 185
R15195 vdd.n1657 vdd.n1451 185
R15196 vdd.n1454 vdd.n1452 185
R15197 vdd.n1653 vdd.n1456 185
R15198 vdd.n1652 vdd.n1457 185
R15199 vdd.n1651 vdd.n1459 185
R15200 vdd.n1462 vdd.n1460 185
R15201 vdd.n1647 vdd.n1464 185
R15202 vdd.n1646 vdd.n1465 185
R15203 vdd.n1645 vdd.n1467 185
R15204 vdd.n1470 vdd.n1468 185
R15205 vdd.n1641 vdd.n1472 185
R15206 vdd.n1640 vdd.n1473 185
R15207 vdd.n1639 vdd.n1475 185
R15208 vdd.n1480 vdd.n1478 185
R15209 vdd.n1635 vdd.n1482 185
R15210 vdd.n1634 vdd.n1483 185
R15211 vdd.n1633 vdd.n1485 185
R15212 vdd.n1488 vdd.n1486 185
R15213 vdd.n1629 vdd.n1490 185
R15214 vdd.n1628 vdd.n1491 185
R15215 vdd.n1627 vdd.n1493 185
R15216 vdd.n1496 vdd.n1494 185
R15217 vdd.n1623 vdd.n1498 185
R15218 vdd.n1622 vdd.n1499 185
R15219 vdd.n1621 vdd.n1501 185
R15220 vdd.n1504 vdd.n1502 185
R15221 vdd.n1617 vdd.n1506 185
R15222 vdd.n1616 vdd.n1507 185
R15223 vdd.n1615 vdd.n1509 185
R15224 vdd.n1512 vdd.n1510 185
R15225 vdd.n1611 vdd.n1514 185
R15226 vdd.n1610 vdd.n1515 185
R15227 vdd.n1609 vdd.n1517 185
R15228 vdd.n1520 vdd.n1518 185
R15229 vdd.n1605 vdd.n1522 185
R15230 vdd.n1604 vdd.n1601 185
R15231 vdd.n1599 vdd.n1523 185
R15232 vdd.n1598 vdd.n1597 185
R15233 vdd.n1528 vdd.n1525 185
R15234 vdd.n1593 vdd.n1529 185
R15235 vdd.n1592 vdd.n1531 185
R15236 vdd.n1591 vdd.n1532 185
R15237 vdd.n1536 vdd.n1533 185
R15238 vdd.n1587 vdd.n1537 185
R15239 vdd.n1586 vdd.n1539 185
R15240 vdd.n1585 vdd.n1540 185
R15241 vdd.n1544 vdd.n1541 185
R15242 vdd.n1581 vdd.n1545 185
R15243 vdd.n1580 vdd.n1547 185
R15244 vdd.n1579 vdd.n1548 185
R15245 vdd.n1552 vdd.n1549 185
R15246 vdd.n1575 vdd.n1553 185
R15247 vdd.n1574 vdd.n1555 185
R15248 vdd.n1573 vdd.n1556 185
R15249 vdd.n1560 vdd.n1557 185
R15250 vdd.n1569 vdd.n1561 185
R15251 vdd.n1568 vdd.n1563 185
R15252 vdd.n1564 vdd.n1436 185
R15253 vdd.n1437 vdd.n1436 185
R15254 vdd.n2073 vdd.n2072 185
R15255 vdd.n2077 vdd.n1353 185
R15256 vdd.n1352 vdd.n1346 185
R15257 vdd.n1350 vdd.n1349 185
R15258 vdd.n1348 vdd.n1107 185
R15259 vdd.n2081 vdd.n1104 185
R15260 vdd.n2083 vdd.n2082 185
R15261 vdd.n2085 vdd.n1102 185
R15262 vdd.n2087 vdd.n2086 185
R15263 vdd.n2088 vdd.n1097 185
R15264 vdd.n2090 vdd.n2089 185
R15265 vdd.n2092 vdd.n1095 185
R15266 vdd.n2094 vdd.n2093 185
R15267 vdd.n2095 vdd.n1090 185
R15268 vdd.n2097 vdd.n2096 185
R15269 vdd.n2099 vdd.n1088 185
R15270 vdd.n2101 vdd.n2100 185
R15271 vdd.n2102 vdd.n1084 185
R15272 vdd.n2104 vdd.n2103 185
R15273 vdd.n2106 vdd.n1081 185
R15274 vdd.n2108 vdd.n2107 185
R15275 vdd.n1082 vdd.n1075 185
R15276 vdd.n2112 vdd.n1079 185
R15277 vdd.n2113 vdd.n1071 185
R15278 vdd.n2115 vdd.n2114 185
R15279 vdd.n2117 vdd.n1069 185
R15280 vdd.n2119 vdd.n2118 185
R15281 vdd.n2120 vdd.n1064 185
R15282 vdd.n2122 vdd.n2121 185
R15283 vdd.n2124 vdd.n1062 185
R15284 vdd.n2126 vdd.n2125 185
R15285 vdd.n2127 vdd.n1057 185
R15286 vdd.n2129 vdd.n2128 185
R15287 vdd.n2131 vdd.n1055 185
R15288 vdd.n2133 vdd.n2132 185
R15289 vdd.n2134 vdd.n1050 185
R15290 vdd.n2136 vdd.n2135 185
R15291 vdd.n2138 vdd.n1048 185
R15292 vdd.n2140 vdd.n2139 185
R15293 vdd.n2141 vdd.n1044 185
R15294 vdd.n2143 vdd.n2142 185
R15295 vdd.n2145 vdd.n1041 185
R15296 vdd.n2147 vdd.n2146 185
R15297 vdd.n1042 vdd.n1035 185
R15298 vdd.n2151 vdd.n1039 185
R15299 vdd.n2152 vdd.n1031 185
R15300 vdd.n2154 vdd.n2153 185
R15301 vdd.n2156 vdd.n1029 185
R15302 vdd.n2158 vdd.n2157 185
R15303 vdd.n2159 vdd.n1024 185
R15304 vdd.n2161 vdd.n2160 185
R15305 vdd.n2163 vdd.n1022 185
R15306 vdd.n2165 vdd.n2164 185
R15307 vdd.n2166 vdd.n1017 185
R15308 vdd.n2168 vdd.n2167 185
R15309 vdd.n2170 vdd.n1015 185
R15310 vdd.n2172 vdd.n2171 185
R15311 vdd.n2173 vdd.n1013 185
R15312 vdd.n2175 vdd.n2174 185
R15313 vdd.n2178 vdd.n2177 185
R15314 vdd.n2180 vdd.n2179 185
R15315 vdd.n2182 vdd.n1011 185
R15316 vdd.n2184 vdd.n2183 185
R15317 vdd.n1358 vdd.n1010 185
R15318 vdd.n2071 vdd.n1356 185
R15319 vdd.n2071 vdd.n2070 185
R15320 vdd.n1366 vdd.n1355 185
R15321 vdd.n2061 vdd.n1355 185
R15322 vdd.n2060 vdd.n2059 185
R15323 vdd.n2062 vdd.n2060 185
R15324 vdd.n1365 vdd.n1364 185
R15325 vdd.n1364 vdd.n1363 185
R15326 vdd.n2053 vdd.n2052 185
R15327 vdd.n2052 vdd.n2051 185
R15328 vdd.n1369 vdd.n1368 185
R15329 vdd.n2042 vdd.n1369 185
R15330 vdd.n2041 vdd.n2040 185
R15331 vdd.n2043 vdd.n2041 185
R15332 vdd.n1376 vdd.n1375 185
R15333 vdd.n1380 vdd.n1375 185
R15334 vdd.n2036 vdd.n2035 185
R15335 vdd.n2035 vdd.n2034 185
R15336 vdd.n1379 vdd.n1378 185
R15337 vdd.n2025 vdd.n1379 185
R15338 vdd.n2024 vdd.n2023 185
R15339 vdd.n2026 vdd.n2024 185
R15340 vdd.n1388 vdd.n1387 185
R15341 vdd.n1387 vdd.n1386 185
R15342 vdd.n2019 vdd.n2018 185
R15343 vdd.n2018 vdd.n2017 185
R15344 vdd.n1391 vdd.n1390 185
R15345 vdd.n1392 vdd.n1391 185
R15346 vdd.n1726 vdd.n1725 185
R15347 vdd.n1727 vdd.n1726 185
R15348 vdd.n1399 vdd.n1398 185
R15349 vdd.n1403 vdd.n1398 185
R15350 vdd.n1721 vdd.n1720 185
R15351 vdd.n1720 vdd.n1719 185
R15352 vdd.n1402 vdd.n1401 185
R15353 vdd.n1710 vdd.n1402 185
R15354 vdd.n1709 vdd.n1708 185
R15355 vdd.n1711 vdd.n1709 185
R15356 vdd.n1410 vdd.n1409 185
R15357 vdd.n1415 vdd.n1409 185
R15358 vdd.n1704 vdd.n1703 185
R15359 vdd.n1703 vdd.n1702 185
R15360 vdd.n1413 vdd.n1412 185
R15361 vdd.n1414 vdd.n1413 185
R15362 vdd.n1693 vdd.n1692 185
R15363 vdd.n1694 vdd.n1693 185
R15364 vdd.n1423 vdd.n1422 185
R15365 vdd.n1422 vdd.n1421 185
R15366 vdd.n1688 vdd.n1687 185
R15367 vdd.n1687 vdd.n1686 185
R15368 vdd.n1426 vdd.n1425 185
R15369 vdd.n1427 vdd.n1426 185
R15370 vdd.n1677 vdd.n1676 185
R15371 vdd.n1678 vdd.n1677 185
R15372 vdd.n1434 vdd.n1433 185
R15373 vdd.n1438 vdd.n1433 185
R15374 vdd.n1672 vdd.n1671 185
R15375 vdd.n1671 vdd.n1670 185
R15376 vdd.n828 vdd.n826 185
R15377 vdd.n2424 vdd.n826 185
R15378 vdd.n2346 vdd.n846 185
R15379 vdd.n846 vdd.n833 185
R15380 vdd.n2348 vdd.n2347 185
R15381 vdd.n2349 vdd.n2348 185
R15382 vdd.n2345 vdd.n845 185
R15383 vdd.n1227 vdd.n845 185
R15384 vdd.n2344 vdd.n2343 185
R15385 vdd.n2343 vdd.n2342 185
R15386 vdd.n848 vdd.n847 185
R15387 vdd.n849 vdd.n848 185
R15388 vdd.n2333 vdd.n2332 185
R15389 vdd.n2334 vdd.n2333 185
R15390 vdd.n2331 vdd.n859 185
R15391 vdd.n859 vdd.n856 185
R15392 vdd.n2330 vdd.n2329 185
R15393 vdd.n2329 vdd.n2328 185
R15394 vdd.n861 vdd.n860 185
R15395 vdd.n1253 vdd.n861 185
R15396 vdd.n2321 vdd.n2320 185
R15397 vdd.n2322 vdd.n2321 185
R15398 vdd.n2319 vdd.n869 185
R15399 vdd.n874 vdd.n869 185
R15400 vdd.n2318 vdd.n2317 185
R15401 vdd.n2317 vdd.n2316 185
R15402 vdd.n871 vdd.n870 185
R15403 vdd.n880 vdd.n871 185
R15404 vdd.n2309 vdd.n2308 185
R15405 vdd.n2310 vdd.n2309 185
R15406 vdd.n2307 vdd.n881 185
R15407 vdd.n1265 vdd.n881 185
R15408 vdd.n2306 vdd.n2305 185
R15409 vdd.n2305 vdd.n2304 185
R15410 vdd.n883 vdd.n882 185
R15411 vdd.n884 vdd.n883 185
R15412 vdd.n2297 vdd.n2296 185
R15413 vdd.n2298 vdd.n2297 185
R15414 vdd.n2295 vdd.n893 185
R15415 vdd.n893 vdd.n890 185
R15416 vdd.n2294 vdd.n2293 185
R15417 vdd.n2293 vdd.n2292 185
R15418 vdd.n895 vdd.n894 185
R15419 vdd.n904 vdd.n895 185
R15420 vdd.n2284 vdd.n2283 185
R15421 vdd.n2285 vdd.n2284 185
R15422 vdd.n2282 vdd.n905 185
R15423 vdd.n911 vdd.n905 185
R15424 vdd.n2281 vdd.n2280 185
R15425 vdd.n2280 vdd.n2279 185
R15426 vdd.n907 vdd.n906 185
R15427 vdd.n908 vdd.n907 185
R15428 vdd.n2272 vdd.n2271 185
R15429 vdd.n2273 vdd.n2272 185
R15430 vdd.n2270 vdd.n918 185
R15431 vdd.n918 vdd.n915 185
R15432 vdd.n2269 vdd.n2268 185
R15433 vdd.n2268 vdd.n2267 185
R15434 vdd.n920 vdd.n919 185
R15435 vdd.n921 vdd.n920 185
R15436 vdd.n2260 vdd.n2259 185
R15437 vdd.n2261 vdd.n2260 185
R15438 vdd.n2258 vdd.n929 185
R15439 vdd.n934 vdd.n929 185
R15440 vdd.n2257 vdd.n2256 185
R15441 vdd.n2256 vdd.n2255 185
R15442 vdd.n931 vdd.n930 185
R15443 vdd.n940 vdd.n931 185
R15444 vdd.n2248 vdd.n2247 185
R15445 vdd.n2249 vdd.n2248 185
R15446 vdd.n2246 vdd.n941 185
R15447 vdd.n947 vdd.n941 185
R15448 vdd.n2245 vdd.n2244 185
R15449 vdd.n2244 vdd.n2243 185
R15450 vdd.n943 vdd.n942 185
R15451 vdd.n944 vdd.n943 185
R15452 vdd.n2236 vdd.n2235 185
R15453 vdd.n2237 vdd.n2236 185
R15454 vdd.n2234 vdd.n954 185
R15455 vdd.n954 vdd.n951 185
R15456 vdd.n2233 vdd.n2232 185
R15457 vdd.n2232 vdd.n2231 185
R15458 vdd.n956 vdd.n955 185
R15459 vdd.n965 vdd.n956 185
R15460 vdd.n2224 vdd.n2223 185
R15461 vdd.n2225 vdd.n2224 185
R15462 vdd.n2222 vdd.n966 185
R15463 vdd.n966 vdd.n962 185
R15464 vdd.n2221 vdd.n2220 185
R15465 vdd.n968 vdd.n967 185
R15466 vdd.n2217 vdd.n2216 185
R15467 vdd.n2218 vdd.n2217 185
R15468 vdd.n2215 vdd.n1004 185
R15469 vdd.n2214 vdd.n2213 185
R15470 vdd.n2212 vdd.n2211 185
R15471 vdd.n2210 vdd.n2209 185
R15472 vdd.n2208 vdd.n2207 185
R15473 vdd.n2206 vdd.n2205 185
R15474 vdd.n2204 vdd.n2203 185
R15475 vdd.n2202 vdd.n2201 185
R15476 vdd.n2200 vdd.n2199 185
R15477 vdd.n2198 vdd.n2197 185
R15478 vdd.n2196 vdd.n2195 185
R15479 vdd.n2194 vdd.n2193 185
R15480 vdd.n2192 vdd.n2191 185
R15481 vdd.n2190 vdd.n2189 185
R15482 vdd.n2188 vdd.n2187 185
R15483 vdd.n1149 vdd.n1005 185
R15484 vdd.n1151 vdd.n1150 185
R15485 vdd.n1153 vdd.n1152 185
R15486 vdd.n1155 vdd.n1154 185
R15487 vdd.n1157 vdd.n1156 185
R15488 vdd.n1159 vdd.n1158 185
R15489 vdd.n1161 vdd.n1160 185
R15490 vdd.n1163 vdd.n1162 185
R15491 vdd.n1165 vdd.n1164 185
R15492 vdd.n1167 vdd.n1166 185
R15493 vdd.n1169 vdd.n1168 185
R15494 vdd.n1171 vdd.n1170 185
R15495 vdd.n1173 vdd.n1172 185
R15496 vdd.n1175 vdd.n1174 185
R15497 vdd.n1178 vdd.n1177 185
R15498 vdd.n1180 vdd.n1179 185
R15499 vdd.n1182 vdd.n1181 185
R15500 vdd.n2427 vdd.n2426 185
R15501 vdd.n2429 vdd.n2428 185
R15502 vdd.n2431 vdd.n2430 185
R15503 vdd.n2434 vdd.n2433 185
R15504 vdd.n2436 vdd.n2435 185
R15505 vdd.n2438 vdd.n2437 185
R15506 vdd.n2440 vdd.n2439 185
R15507 vdd.n2442 vdd.n2441 185
R15508 vdd.n2444 vdd.n2443 185
R15509 vdd.n2446 vdd.n2445 185
R15510 vdd.n2448 vdd.n2447 185
R15511 vdd.n2450 vdd.n2449 185
R15512 vdd.n2452 vdd.n2451 185
R15513 vdd.n2454 vdd.n2453 185
R15514 vdd.n2456 vdd.n2455 185
R15515 vdd.n2458 vdd.n2457 185
R15516 vdd.n2460 vdd.n2459 185
R15517 vdd.n2462 vdd.n2461 185
R15518 vdd.n2464 vdd.n2463 185
R15519 vdd.n2466 vdd.n2465 185
R15520 vdd.n2468 vdd.n2467 185
R15521 vdd.n2470 vdd.n2469 185
R15522 vdd.n2472 vdd.n2471 185
R15523 vdd.n2474 vdd.n2473 185
R15524 vdd.n2476 vdd.n2475 185
R15525 vdd.n2478 vdd.n2477 185
R15526 vdd.n2480 vdd.n2479 185
R15527 vdd.n2482 vdd.n2481 185
R15528 vdd.n2484 vdd.n2483 185
R15529 vdd.n2486 vdd.n2485 185
R15530 vdd.n2488 vdd.n2487 185
R15531 vdd.n2490 vdd.n2489 185
R15532 vdd.n2492 vdd.n2491 185
R15533 vdd.n2493 vdd.n827 185
R15534 vdd.n2495 vdd.n2494 185
R15535 vdd.n2496 vdd.n2495 185
R15536 vdd.n2425 vdd.n831 185
R15537 vdd.n2425 vdd.n2424 185
R15538 vdd.n1225 vdd.n832 185
R15539 vdd.n833 vdd.n832 185
R15540 vdd.n1226 vdd.n843 185
R15541 vdd.n2349 vdd.n843 185
R15542 vdd.n1229 vdd.n1228 185
R15543 vdd.n1228 vdd.n1227 185
R15544 vdd.n1230 vdd.n850 185
R15545 vdd.n2342 vdd.n850 185
R15546 vdd.n1232 vdd.n1231 185
R15547 vdd.n1231 vdd.n849 185
R15548 vdd.n1233 vdd.n857 185
R15549 vdd.n2334 vdd.n857 185
R15550 vdd.n1235 vdd.n1234 185
R15551 vdd.n1234 vdd.n856 185
R15552 vdd.n1236 vdd.n862 185
R15553 vdd.n2328 vdd.n862 185
R15554 vdd.n1255 vdd.n1254 185
R15555 vdd.n1254 vdd.n1253 185
R15556 vdd.n1256 vdd.n867 185
R15557 vdd.n2322 vdd.n867 185
R15558 vdd.n1258 vdd.n1257 185
R15559 vdd.n1257 vdd.n874 185
R15560 vdd.n1259 vdd.n872 185
R15561 vdd.n2316 vdd.n872 185
R15562 vdd.n1261 vdd.n1260 185
R15563 vdd.n1260 vdd.n880 185
R15564 vdd.n1262 vdd.n878 185
R15565 vdd.n2310 vdd.n878 185
R15566 vdd.n1264 vdd.n1263 185
R15567 vdd.n1265 vdd.n1264 185
R15568 vdd.n1224 vdd.n885 185
R15569 vdd.n2304 vdd.n885 185
R15570 vdd.n1223 vdd.n1222 185
R15571 vdd.n1222 vdd.n884 185
R15572 vdd.n1221 vdd.n891 185
R15573 vdd.n2298 vdd.n891 185
R15574 vdd.n1220 vdd.n1219 185
R15575 vdd.n1219 vdd.n890 185
R15576 vdd.n1218 vdd.n896 185
R15577 vdd.n2292 vdd.n896 185
R15578 vdd.n1217 vdd.n1216 185
R15579 vdd.n1216 vdd.n904 185
R15580 vdd.n1215 vdd.n902 185
R15581 vdd.n2285 vdd.n902 185
R15582 vdd.n1214 vdd.n1213 185
R15583 vdd.n1213 vdd.n911 185
R15584 vdd.n1212 vdd.n909 185
R15585 vdd.n2279 vdd.n909 185
R15586 vdd.n1211 vdd.n1210 185
R15587 vdd.n1210 vdd.n908 185
R15588 vdd.n1209 vdd.n916 185
R15589 vdd.n2273 vdd.n916 185
R15590 vdd.n1208 vdd.n1207 185
R15591 vdd.n1207 vdd.n915 185
R15592 vdd.n1206 vdd.n922 185
R15593 vdd.n2267 vdd.n922 185
R15594 vdd.n1205 vdd.n1204 185
R15595 vdd.n1204 vdd.n921 185
R15596 vdd.n1203 vdd.n927 185
R15597 vdd.n2261 vdd.n927 185
R15598 vdd.n1202 vdd.n1201 185
R15599 vdd.n1201 vdd.n934 185
R15600 vdd.n1200 vdd.n932 185
R15601 vdd.n2255 vdd.n932 185
R15602 vdd.n1199 vdd.n1198 185
R15603 vdd.n1198 vdd.n940 185
R15604 vdd.n1197 vdd.n938 185
R15605 vdd.n2249 vdd.n938 185
R15606 vdd.n1196 vdd.n1195 185
R15607 vdd.n1195 vdd.n947 185
R15608 vdd.n1194 vdd.n945 185
R15609 vdd.n2243 vdd.n945 185
R15610 vdd.n1193 vdd.n1192 185
R15611 vdd.n1192 vdd.n944 185
R15612 vdd.n1191 vdd.n952 185
R15613 vdd.n2237 vdd.n952 185
R15614 vdd.n1190 vdd.n1189 185
R15615 vdd.n1189 vdd.n951 185
R15616 vdd.n1188 vdd.n957 185
R15617 vdd.n2231 vdd.n957 185
R15618 vdd.n1187 vdd.n1186 185
R15619 vdd.n1186 vdd.n965 185
R15620 vdd.n1185 vdd.n963 185
R15621 vdd.n2225 vdd.n963 185
R15622 vdd.n1184 vdd.n1183 185
R15623 vdd.n1183 vdd.n962 185
R15624 vdd.n3409 vdd.n3408 185
R15625 vdd.n3410 vdd.n3409 185
R15626 vdd.n347 vdd.n346 185
R15627 vdd.n3411 vdd.n347 185
R15628 vdd.n3414 vdd.n3413 185
R15629 vdd.n3413 vdd.n3412 185
R15630 vdd.n3415 vdd.n341 185
R15631 vdd.n341 vdd.n340 185
R15632 vdd.n3417 vdd.n3416 185
R15633 vdd.n3418 vdd.n3417 185
R15634 vdd.n336 vdd.n335 185
R15635 vdd.n3419 vdd.n336 185
R15636 vdd.n3422 vdd.n3421 185
R15637 vdd.n3421 vdd.n3420 185
R15638 vdd.n3423 vdd.n330 185
R15639 vdd.n330 vdd.n329 185
R15640 vdd.n3425 vdd.n3424 185
R15641 vdd.n3426 vdd.n3425 185
R15642 vdd.n324 vdd.n323 185
R15643 vdd.n3427 vdd.n324 185
R15644 vdd.n3430 vdd.n3429 185
R15645 vdd.n3429 vdd.n3428 185
R15646 vdd.n3431 vdd.n319 185
R15647 vdd.n325 vdd.n319 185
R15648 vdd.n3433 vdd.n3432 185
R15649 vdd.n3434 vdd.n3433 185
R15650 vdd.n315 vdd.n313 185
R15651 vdd.n3435 vdd.n315 185
R15652 vdd.n3438 vdd.n3437 185
R15653 vdd.n3437 vdd.n3436 185
R15654 vdd.n314 vdd.n312 185
R15655 vdd.n481 vdd.n314 185
R15656 vdd.n3260 vdd.n3259 185
R15657 vdd.n3261 vdd.n3260 185
R15658 vdd.n483 vdd.n482 185
R15659 vdd.n3252 vdd.n482 185
R15660 vdd.n3255 vdd.n3254 185
R15661 vdd.n3254 vdd.n3253 185
R15662 vdd.n486 vdd.n485 185
R15663 vdd.n493 vdd.n486 185
R15664 vdd.n3243 vdd.n3242 185
R15665 vdd.n3244 vdd.n3243 185
R15666 vdd.n495 vdd.n494 185
R15667 vdd.n494 vdd.n492 185
R15668 vdd.n3238 vdd.n3237 185
R15669 vdd.n3237 vdd.n3236 185
R15670 vdd.n498 vdd.n497 185
R15671 vdd.n499 vdd.n498 185
R15672 vdd.n3227 vdd.n3226 185
R15673 vdd.n3228 vdd.n3227 185
R15674 vdd.n507 vdd.n506 185
R15675 vdd.n506 vdd.n505 185
R15676 vdd.n3222 vdd.n3221 185
R15677 vdd.n3221 vdd.n3220 185
R15678 vdd.n510 vdd.n509 185
R15679 vdd.n511 vdd.n510 185
R15680 vdd.n3211 vdd.n3210 185
R15681 vdd.n3212 vdd.n3211 185
R15682 vdd.n3207 vdd.n517 185
R15683 vdd.n3206 vdd.n3205 185
R15684 vdd.n3203 vdd.n519 185
R15685 vdd.n3203 vdd.n516 185
R15686 vdd.n3202 vdd.n3201 185
R15687 vdd.n3200 vdd.n3199 185
R15688 vdd.n3198 vdd.n3197 185
R15689 vdd.n3196 vdd.n3195 185
R15690 vdd.n3194 vdd.n525 185
R15691 vdd.n3192 vdd.n3191 185
R15692 vdd.n3190 vdd.n526 185
R15693 vdd.n3189 vdd.n3188 185
R15694 vdd.n3186 vdd.n531 185
R15695 vdd.n3184 vdd.n3183 185
R15696 vdd.n3182 vdd.n532 185
R15697 vdd.n3181 vdd.n3180 185
R15698 vdd.n3178 vdd.n537 185
R15699 vdd.n3176 vdd.n3175 185
R15700 vdd.n3174 vdd.n538 185
R15701 vdd.n3173 vdd.n3172 185
R15702 vdd.n3170 vdd.n545 185
R15703 vdd.n3168 vdd.n3167 185
R15704 vdd.n3166 vdd.n546 185
R15705 vdd.n3165 vdd.n3164 185
R15706 vdd.n3162 vdd.n551 185
R15707 vdd.n3160 vdd.n3159 185
R15708 vdd.n3158 vdd.n552 185
R15709 vdd.n3157 vdd.n3156 185
R15710 vdd.n3154 vdd.n557 185
R15711 vdd.n3152 vdd.n3151 185
R15712 vdd.n3150 vdd.n558 185
R15713 vdd.n3149 vdd.n3148 185
R15714 vdd.n3146 vdd.n563 185
R15715 vdd.n3144 vdd.n3143 185
R15716 vdd.n3142 vdd.n564 185
R15717 vdd.n3141 vdd.n3140 185
R15718 vdd.n3138 vdd.n569 185
R15719 vdd.n3136 vdd.n3135 185
R15720 vdd.n3134 vdd.n570 185
R15721 vdd.n3133 vdd.n3132 185
R15722 vdd.n3130 vdd.n575 185
R15723 vdd.n3128 vdd.n3127 185
R15724 vdd.n3126 vdd.n576 185
R15725 vdd.n585 vdd.n579 185
R15726 vdd.n3122 vdd.n3121 185
R15727 vdd.n3119 vdd.n583 185
R15728 vdd.n3118 vdd.n3117 185
R15729 vdd.n3116 vdd.n3115 185
R15730 vdd.n3114 vdd.n589 185
R15731 vdd.n3112 vdd.n3111 185
R15732 vdd.n3110 vdd.n590 185
R15733 vdd.n3109 vdd.n3108 185
R15734 vdd.n3106 vdd.n595 185
R15735 vdd.n3104 vdd.n3103 185
R15736 vdd.n3102 vdd.n596 185
R15737 vdd.n3101 vdd.n3100 185
R15738 vdd.n3098 vdd.n601 185
R15739 vdd.n3096 vdd.n3095 185
R15740 vdd.n3094 vdd.n602 185
R15741 vdd.n3093 vdd.n3092 185
R15742 vdd.n3090 vdd.n3089 185
R15743 vdd.n3088 vdd.n3087 185
R15744 vdd.n3086 vdd.n3085 185
R15745 vdd.n3084 vdd.n3083 185
R15746 vdd.n3079 vdd.n515 185
R15747 vdd.n516 vdd.n515 185
R15748 vdd.n3292 vdd.n3291 185
R15749 vdd.n3296 vdd.n462 185
R15750 vdd.n3298 vdd.n3297 185
R15751 vdd.n3300 vdd.n460 185
R15752 vdd.n3302 vdd.n3301 185
R15753 vdd.n3303 vdd.n455 185
R15754 vdd.n3305 vdd.n3304 185
R15755 vdd.n3307 vdd.n453 185
R15756 vdd.n3309 vdd.n3308 185
R15757 vdd.n3310 vdd.n448 185
R15758 vdd.n3312 vdd.n3311 185
R15759 vdd.n3314 vdd.n446 185
R15760 vdd.n3316 vdd.n3315 185
R15761 vdd.n3317 vdd.n441 185
R15762 vdd.n3319 vdd.n3318 185
R15763 vdd.n3321 vdd.n439 185
R15764 vdd.n3323 vdd.n3322 185
R15765 vdd.n3324 vdd.n435 185
R15766 vdd.n3326 vdd.n3325 185
R15767 vdd.n3328 vdd.n432 185
R15768 vdd.n3330 vdd.n3329 185
R15769 vdd.n433 vdd.n426 185
R15770 vdd.n3334 vdd.n430 185
R15771 vdd.n3335 vdd.n422 185
R15772 vdd.n3337 vdd.n3336 185
R15773 vdd.n3339 vdd.n420 185
R15774 vdd.n3341 vdd.n3340 185
R15775 vdd.n3342 vdd.n415 185
R15776 vdd.n3344 vdd.n3343 185
R15777 vdd.n3346 vdd.n413 185
R15778 vdd.n3348 vdd.n3347 185
R15779 vdd.n3349 vdd.n408 185
R15780 vdd.n3351 vdd.n3350 185
R15781 vdd.n3353 vdd.n406 185
R15782 vdd.n3355 vdd.n3354 185
R15783 vdd.n3356 vdd.n401 185
R15784 vdd.n3358 vdd.n3357 185
R15785 vdd.n3360 vdd.n399 185
R15786 vdd.n3362 vdd.n3361 185
R15787 vdd.n3363 vdd.n395 185
R15788 vdd.n3365 vdd.n3364 185
R15789 vdd.n3367 vdd.n392 185
R15790 vdd.n3369 vdd.n3368 185
R15791 vdd.n393 vdd.n386 185
R15792 vdd.n3373 vdd.n390 185
R15793 vdd.n3374 vdd.n382 185
R15794 vdd.n3376 vdd.n3375 185
R15795 vdd.n3378 vdd.n380 185
R15796 vdd.n3380 vdd.n3379 185
R15797 vdd.n3381 vdd.n375 185
R15798 vdd.n3383 vdd.n3382 185
R15799 vdd.n3385 vdd.n373 185
R15800 vdd.n3387 vdd.n3386 185
R15801 vdd.n3388 vdd.n368 185
R15802 vdd.n3390 vdd.n3389 185
R15803 vdd.n3392 vdd.n366 185
R15804 vdd.n3394 vdd.n3393 185
R15805 vdd.n3395 vdd.n360 185
R15806 vdd.n3397 vdd.n3396 185
R15807 vdd.n3399 vdd.n359 185
R15808 vdd.n3400 vdd.n358 185
R15809 vdd.n3403 vdd.n3402 185
R15810 vdd.n3404 vdd.n356 185
R15811 vdd.n3405 vdd.n352 185
R15812 vdd.n3287 vdd.n350 185
R15813 vdd.n3410 vdd.n350 185
R15814 vdd.n3286 vdd.n349 185
R15815 vdd.n3411 vdd.n349 185
R15816 vdd.n3285 vdd.n348 185
R15817 vdd.n3412 vdd.n348 185
R15818 vdd.n468 vdd.n467 185
R15819 vdd.n467 vdd.n340 185
R15820 vdd.n3281 vdd.n339 185
R15821 vdd.n3418 vdd.n339 185
R15822 vdd.n3280 vdd.n338 185
R15823 vdd.n3419 vdd.n338 185
R15824 vdd.n3279 vdd.n337 185
R15825 vdd.n3420 vdd.n337 185
R15826 vdd.n471 vdd.n470 185
R15827 vdd.n470 vdd.n329 185
R15828 vdd.n3275 vdd.n328 185
R15829 vdd.n3426 vdd.n328 185
R15830 vdd.n3274 vdd.n327 185
R15831 vdd.n3427 vdd.n327 185
R15832 vdd.n3273 vdd.n326 185
R15833 vdd.n3428 vdd.n326 185
R15834 vdd.n474 vdd.n473 185
R15835 vdd.n473 vdd.n325 185
R15836 vdd.n3269 vdd.n318 185
R15837 vdd.n3434 vdd.n318 185
R15838 vdd.n3268 vdd.n317 185
R15839 vdd.n3435 vdd.n317 185
R15840 vdd.n3267 vdd.n316 185
R15841 vdd.n3436 vdd.n316 185
R15842 vdd.n480 vdd.n476 185
R15843 vdd.n481 vdd.n480 185
R15844 vdd.n3263 vdd.n3262 185
R15845 vdd.n3262 vdd.n3261 185
R15846 vdd.n479 vdd.n478 185
R15847 vdd.n3252 vdd.n479 185
R15848 vdd.n3251 vdd.n3250 185
R15849 vdd.n3253 vdd.n3251 185
R15850 vdd.n488 vdd.n487 185
R15851 vdd.n493 vdd.n487 185
R15852 vdd.n3246 vdd.n3245 185
R15853 vdd.n3245 vdd.n3244 185
R15854 vdd.n491 vdd.n490 185
R15855 vdd.n492 vdd.n491 185
R15856 vdd.n3235 vdd.n3234 185
R15857 vdd.n3236 vdd.n3235 185
R15858 vdd.n501 vdd.n500 185
R15859 vdd.n500 vdd.n499 185
R15860 vdd.n3230 vdd.n3229 185
R15861 vdd.n3229 vdd.n3228 185
R15862 vdd.n504 vdd.n503 185
R15863 vdd.n505 vdd.n504 185
R15864 vdd.n3219 vdd.n3218 185
R15865 vdd.n3220 vdd.n3219 185
R15866 vdd.n513 vdd.n512 185
R15867 vdd.n512 vdd.n511 185
R15868 vdd.n3214 vdd.n3213 185
R15869 vdd.n3213 vdd.n3212 185
R15870 vdd.n2803 vdd.n2802 185
R15871 vdd.n790 vdd.n789 185
R15872 vdd.n2799 vdd.n2798 185
R15873 vdd.n2800 vdd.n2799 185
R15874 vdd.n2797 vdd.n2531 185
R15875 vdd.n2796 vdd.n2795 185
R15876 vdd.n2794 vdd.n2793 185
R15877 vdd.n2792 vdd.n2791 185
R15878 vdd.n2790 vdd.n2789 185
R15879 vdd.n2788 vdd.n2787 185
R15880 vdd.n2786 vdd.n2785 185
R15881 vdd.n2784 vdd.n2783 185
R15882 vdd.n2782 vdd.n2781 185
R15883 vdd.n2780 vdd.n2779 185
R15884 vdd.n2778 vdd.n2777 185
R15885 vdd.n2776 vdd.n2775 185
R15886 vdd.n2774 vdd.n2773 185
R15887 vdd.n2772 vdd.n2771 185
R15888 vdd.n2770 vdd.n2769 185
R15889 vdd.n2768 vdd.n2767 185
R15890 vdd.n2766 vdd.n2765 185
R15891 vdd.n2764 vdd.n2763 185
R15892 vdd.n2762 vdd.n2761 185
R15893 vdd.n2760 vdd.n2759 185
R15894 vdd.n2758 vdd.n2757 185
R15895 vdd.n2756 vdd.n2755 185
R15896 vdd.n2754 vdd.n2753 185
R15897 vdd.n2752 vdd.n2751 185
R15898 vdd.n2750 vdd.n2749 185
R15899 vdd.n2748 vdd.n2747 185
R15900 vdd.n2746 vdd.n2745 185
R15901 vdd.n2744 vdd.n2743 185
R15902 vdd.n2742 vdd.n2741 185
R15903 vdd.n2739 vdd.n2738 185
R15904 vdd.n2737 vdd.n2736 185
R15905 vdd.n2735 vdd.n2734 185
R15906 vdd.n2980 vdd.n2979 185
R15907 vdd.n2981 vdd.n660 185
R15908 vdd.n2983 vdd.n2982 185
R15909 vdd.n2985 vdd.n658 185
R15910 vdd.n2987 vdd.n2986 185
R15911 vdd.n2988 vdd.n657 185
R15912 vdd.n2990 vdd.n2989 185
R15913 vdd.n2992 vdd.n655 185
R15914 vdd.n2994 vdd.n2993 185
R15915 vdd.n2995 vdd.n654 185
R15916 vdd.n2997 vdd.n2996 185
R15917 vdd.n2999 vdd.n652 185
R15918 vdd.n3001 vdd.n3000 185
R15919 vdd.n3002 vdd.n651 185
R15920 vdd.n3004 vdd.n3003 185
R15921 vdd.n3006 vdd.n649 185
R15922 vdd.n3008 vdd.n3007 185
R15923 vdd.n3010 vdd.n648 185
R15924 vdd.n3012 vdd.n3011 185
R15925 vdd.n3014 vdd.n646 185
R15926 vdd.n3016 vdd.n3015 185
R15927 vdd.n3017 vdd.n645 185
R15928 vdd.n3019 vdd.n3018 185
R15929 vdd.n3021 vdd.n643 185
R15930 vdd.n3023 vdd.n3022 185
R15931 vdd.n3024 vdd.n642 185
R15932 vdd.n3026 vdd.n3025 185
R15933 vdd.n3028 vdd.n640 185
R15934 vdd.n3030 vdd.n3029 185
R15935 vdd.n3031 vdd.n639 185
R15936 vdd.n3033 vdd.n3032 185
R15937 vdd.n3035 vdd.n638 185
R15938 vdd.n3036 vdd.n637 185
R15939 vdd.n3039 vdd.n3038 185
R15940 vdd.n3040 vdd.n635 185
R15941 vdd.n635 vdd.n613 185
R15942 vdd.n2977 vdd.n632 185
R15943 vdd.n3043 vdd.n632 185
R15944 vdd.n2976 vdd.n2975 185
R15945 vdd.n2975 vdd.n631 185
R15946 vdd.n2974 vdd.n664 185
R15947 vdd.n2974 vdd.n2973 185
R15948 vdd.n2617 vdd.n665 185
R15949 vdd.n674 vdd.n665 185
R15950 vdd.n2618 vdd.n672 185
R15951 vdd.n2967 vdd.n672 185
R15952 vdd.n2620 vdd.n2619 185
R15953 vdd.n2619 vdd.n671 185
R15954 vdd.n2621 vdd.n680 185
R15955 vdd.n2916 vdd.n680 185
R15956 vdd.n2623 vdd.n2622 185
R15957 vdd.n2622 vdd.n679 185
R15958 vdd.n2624 vdd.n685 185
R15959 vdd.n2910 vdd.n685 185
R15960 vdd.n2626 vdd.n2625 185
R15961 vdd.n2625 vdd.n692 185
R15962 vdd.n2627 vdd.n690 185
R15963 vdd.n2904 vdd.n690 185
R15964 vdd.n2629 vdd.n2628 185
R15965 vdd.n2628 vdd.n698 185
R15966 vdd.n2630 vdd.n696 185
R15967 vdd.n2898 vdd.n696 185
R15968 vdd.n2632 vdd.n2631 185
R15969 vdd.n2631 vdd.n705 185
R15970 vdd.n2633 vdd.n703 185
R15971 vdd.n2892 vdd.n703 185
R15972 vdd.n2635 vdd.n2634 185
R15973 vdd.n2634 vdd.n702 185
R15974 vdd.n2636 vdd.n710 185
R15975 vdd.n2886 vdd.n710 185
R15976 vdd.n2638 vdd.n2637 185
R15977 vdd.n2637 vdd.n709 185
R15978 vdd.n2639 vdd.n716 185
R15979 vdd.n2880 vdd.n716 185
R15980 vdd.n2641 vdd.n2640 185
R15981 vdd.n2640 vdd.n715 185
R15982 vdd.n2642 vdd.n721 185
R15983 vdd.n2874 vdd.n721 185
R15984 vdd.n2644 vdd.n2643 185
R15985 vdd.n2643 vdd.n729 185
R15986 vdd.n2645 vdd.n727 185
R15987 vdd.n2868 vdd.n727 185
R15988 vdd.n2647 vdd.n2646 185
R15989 vdd.n2646 vdd.n736 185
R15990 vdd.n2648 vdd.n734 185
R15991 vdd.n2862 vdd.n734 185
R15992 vdd.n2650 vdd.n2649 185
R15993 vdd.n2649 vdd.n733 185
R15994 vdd.n2651 vdd.n741 185
R15995 vdd.n2855 vdd.n741 185
R15996 vdd.n2653 vdd.n2652 185
R15997 vdd.n2652 vdd.n740 185
R15998 vdd.n2654 vdd.n746 185
R15999 vdd.n2849 vdd.n746 185
R16000 vdd.n2656 vdd.n2655 185
R16001 vdd.n2655 vdd.n753 185
R16002 vdd.n2657 vdd.n751 185
R16003 vdd.n2843 vdd.n751 185
R16004 vdd.n2659 vdd.n2658 185
R16005 vdd.n2658 vdd.n759 185
R16006 vdd.n2660 vdd.n757 185
R16007 vdd.n2837 vdd.n757 185
R16008 vdd.n2712 vdd.n2711 185
R16009 vdd.n2711 vdd.n2710 185
R16010 vdd.n2713 vdd.n763 185
R16011 vdd.n2831 vdd.n763 185
R16012 vdd.n2715 vdd.n2714 185
R16013 vdd.n2716 vdd.n2715 185
R16014 vdd.n2616 vdd.n769 185
R16015 vdd.n2825 vdd.n769 185
R16016 vdd.n2615 vdd.n2614 185
R16017 vdd.n2614 vdd.n768 185
R16018 vdd.n2613 vdd.n775 185
R16019 vdd.n2819 vdd.n775 185
R16020 vdd.n2612 vdd.n2611 185
R16021 vdd.n2611 vdd.n774 185
R16022 vdd.n2534 vdd.n780 185
R16023 vdd.n2813 vdd.n780 185
R16024 vdd.n2730 vdd.n2729 185
R16025 vdd.n2729 vdd.n2728 185
R16026 vdd.n2731 vdd.n786 185
R16027 vdd.n2807 vdd.n786 185
R16028 vdd.n2733 vdd.n2732 185
R16029 vdd.n2733 vdd.n785 185
R16030 vdd.n2804 vdd.n788 185
R16031 vdd.n788 vdd.n785 185
R16032 vdd.n2806 vdd.n2805 185
R16033 vdd.n2807 vdd.n2806 185
R16034 vdd.n779 vdd.n778 185
R16035 vdd.n2728 vdd.n779 185
R16036 vdd.n2815 vdd.n2814 185
R16037 vdd.n2814 vdd.n2813 185
R16038 vdd.n2816 vdd.n777 185
R16039 vdd.n777 vdd.n774 185
R16040 vdd.n2818 vdd.n2817 185
R16041 vdd.n2819 vdd.n2818 185
R16042 vdd.n767 vdd.n766 185
R16043 vdd.n768 vdd.n767 185
R16044 vdd.n2827 vdd.n2826 185
R16045 vdd.n2826 vdd.n2825 185
R16046 vdd.n2828 vdd.n765 185
R16047 vdd.n2716 vdd.n765 185
R16048 vdd.n2830 vdd.n2829 185
R16049 vdd.n2831 vdd.n2830 185
R16050 vdd.n756 vdd.n755 185
R16051 vdd.n2710 vdd.n756 185
R16052 vdd.n2839 vdd.n2838 185
R16053 vdd.n2838 vdd.n2837 185
R16054 vdd.n2840 vdd.n754 185
R16055 vdd.n759 vdd.n754 185
R16056 vdd.n2842 vdd.n2841 185
R16057 vdd.n2843 vdd.n2842 185
R16058 vdd.n745 vdd.n744 185
R16059 vdd.n753 vdd.n745 185
R16060 vdd.n2851 vdd.n2850 185
R16061 vdd.n2850 vdd.n2849 185
R16062 vdd.n2852 vdd.n743 185
R16063 vdd.n743 vdd.n740 185
R16064 vdd.n2854 vdd.n2853 185
R16065 vdd.n2855 vdd.n2854 185
R16066 vdd.n732 vdd.n731 185
R16067 vdd.n733 vdd.n732 185
R16068 vdd.n2864 vdd.n2863 185
R16069 vdd.n2863 vdd.n2862 185
R16070 vdd.n2865 vdd.n730 185
R16071 vdd.n736 vdd.n730 185
R16072 vdd.n2867 vdd.n2866 185
R16073 vdd.n2868 vdd.n2867 185
R16074 vdd.n720 vdd.n719 185
R16075 vdd.n729 vdd.n720 185
R16076 vdd.n2876 vdd.n2875 185
R16077 vdd.n2875 vdd.n2874 185
R16078 vdd.n2877 vdd.n718 185
R16079 vdd.n718 vdd.n715 185
R16080 vdd.n2879 vdd.n2878 185
R16081 vdd.n2880 vdd.n2879 185
R16082 vdd.n708 vdd.n707 185
R16083 vdd.n709 vdd.n708 185
R16084 vdd.n2888 vdd.n2887 185
R16085 vdd.n2887 vdd.n2886 185
R16086 vdd.n2889 vdd.n706 185
R16087 vdd.n706 vdd.n702 185
R16088 vdd.n2891 vdd.n2890 185
R16089 vdd.n2892 vdd.n2891 185
R16090 vdd.n695 vdd.n694 185
R16091 vdd.n705 vdd.n695 185
R16092 vdd.n2900 vdd.n2899 185
R16093 vdd.n2899 vdd.n2898 185
R16094 vdd.n2901 vdd.n693 185
R16095 vdd.n698 vdd.n693 185
R16096 vdd.n2903 vdd.n2902 185
R16097 vdd.n2904 vdd.n2903 185
R16098 vdd.n684 vdd.n683 185
R16099 vdd.n692 vdd.n684 185
R16100 vdd.n2912 vdd.n2911 185
R16101 vdd.n2911 vdd.n2910 185
R16102 vdd.n2913 vdd.n682 185
R16103 vdd.n682 vdd.n679 185
R16104 vdd.n2915 vdd.n2914 185
R16105 vdd.n2916 vdd.n2915 185
R16106 vdd.n670 vdd.n669 185
R16107 vdd.n671 vdd.n670 185
R16108 vdd.n2969 vdd.n2968 185
R16109 vdd.n2968 vdd.n2967 185
R16110 vdd.n2970 vdd.n668 185
R16111 vdd.n674 vdd.n668 185
R16112 vdd.n2972 vdd.n2971 185
R16113 vdd.n2973 vdd.n2972 185
R16114 vdd.n636 vdd.n634 185
R16115 vdd.n634 vdd.n631 185
R16116 vdd.n3042 vdd.n3041 185
R16117 vdd.n3043 vdd.n3042 185
R16118 vdd.n2423 vdd.n2422 185
R16119 vdd.n2424 vdd.n2423 185
R16120 vdd.n837 vdd.n835 185
R16121 vdd.n835 vdd.n833 185
R16122 vdd.n2338 vdd.n844 185
R16123 vdd.n2349 vdd.n844 185
R16124 vdd.n2339 vdd.n853 185
R16125 vdd.n1227 vdd.n853 185
R16126 vdd.n2341 vdd.n2340 185
R16127 vdd.n2342 vdd.n2341 185
R16128 vdd.n2337 vdd.n852 185
R16129 vdd.n852 vdd.n849 185
R16130 vdd.n2336 vdd.n2335 185
R16131 vdd.n2335 vdd.n2334 185
R16132 vdd.n855 vdd.n854 185
R16133 vdd.n856 vdd.n855 185
R16134 vdd.n2327 vdd.n2326 185
R16135 vdd.n2328 vdd.n2327 185
R16136 vdd.n2325 vdd.n864 185
R16137 vdd.n1253 vdd.n864 185
R16138 vdd.n2324 vdd.n2323 185
R16139 vdd.n2323 vdd.n2322 185
R16140 vdd.n866 vdd.n865 185
R16141 vdd.n874 vdd.n866 185
R16142 vdd.n2315 vdd.n2314 185
R16143 vdd.n2316 vdd.n2315 185
R16144 vdd.n2313 vdd.n875 185
R16145 vdd.n880 vdd.n875 185
R16146 vdd.n2312 vdd.n2311 185
R16147 vdd.n2311 vdd.n2310 185
R16148 vdd.n877 vdd.n876 185
R16149 vdd.n1265 vdd.n877 185
R16150 vdd.n2303 vdd.n2302 185
R16151 vdd.n2304 vdd.n2303 185
R16152 vdd.n2301 vdd.n887 185
R16153 vdd.n887 vdd.n884 185
R16154 vdd.n2300 vdd.n2299 185
R16155 vdd.n2299 vdd.n2298 185
R16156 vdd.n889 vdd.n888 185
R16157 vdd.n890 vdd.n889 185
R16158 vdd.n2291 vdd.n2290 185
R16159 vdd.n2292 vdd.n2291 185
R16160 vdd.n2288 vdd.n898 185
R16161 vdd.n904 vdd.n898 185
R16162 vdd.n2287 vdd.n2286 185
R16163 vdd.n2286 vdd.n2285 185
R16164 vdd.n901 vdd.n900 185
R16165 vdd.n911 vdd.n901 185
R16166 vdd.n2278 vdd.n2277 185
R16167 vdd.n2279 vdd.n2278 185
R16168 vdd.n2276 vdd.n912 185
R16169 vdd.n912 vdd.n908 185
R16170 vdd.n2275 vdd.n2274 185
R16171 vdd.n2274 vdd.n2273 185
R16172 vdd.n914 vdd.n913 185
R16173 vdd.n915 vdd.n914 185
R16174 vdd.n2266 vdd.n2265 185
R16175 vdd.n2267 vdd.n2266 185
R16176 vdd.n2264 vdd.n924 185
R16177 vdd.n924 vdd.n921 185
R16178 vdd.n2263 vdd.n2262 185
R16179 vdd.n2262 vdd.n2261 185
R16180 vdd.n926 vdd.n925 185
R16181 vdd.n934 vdd.n926 185
R16182 vdd.n2254 vdd.n2253 185
R16183 vdd.n2255 vdd.n2254 185
R16184 vdd.n2252 vdd.n935 185
R16185 vdd.n940 vdd.n935 185
R16186 vdd.n2251 vdd.n2250 185
R16187 vdd.n2250 vdd.n2249 185
R16188 vdd.n937 vdd.n936 185
R16189 vdd.n947 vdd.n937 185
R16190 vdd.n2242 vdd.n2241 185
R16191 vdd.n2243 vdd.n2242 185
R16192 vdd.n2240 vdd.n948 185
R16193 vdd.n948 vdd.n944 185
R16194 vdd.n2239 vdd.n2238 185
R16195 vdd.n2238 vdd.n2237 185
R16196 vdd.n950 vdd.n949 185
R16197 vdd.n951 vdd.n950 185
R16198 vdd.n2230 vdd.n2229 185
R16199 vdd.n2231 vdd.n2230 185
R16200 vdd.n2228 vdd.n959 185
R16201 vdd.n965 vdd.n959 185
R16202 vdd.n2227 vdd.n2226 185
R16203 vdd.n2226 vdd.n2225 185
R16204 vdd.n961 vdd.n960 185
R16205 vdd.n962 vdd.n961 185
R16206 vdd.n2354 vdd.n808 185
R16207 vdd.n2496 vdd.n808 185
R16208 vdd.n2356 vdd.n2355 185
R16209 vdd.n2358 vdd.n2357 185
R16210 vdd.n2360 vdd.n2359 185
R16211 vdd.n2362 vdd.n2361 185
R16212 vdd.n2364 vdd.n2363 185
R16213 vdd.n2366 vdd.n2365 185
R16214 vdd.n2368 vdd.n2367 185
R16215 vdd.n2370 vdd.n2369 185
R16216 vdd.n2372 vdd.n2371 185
R16217 vdd.n2374 vdd.n2373 185
R16218 vdd.n2376 vdd.n2375 185
R16219 vdd.n2378 vdd.n2377 185
R16220 vdd.n2380 vdd.n2379 185
R16221 vdd.n2382 vdd.n2381 185
R16222 vdd.n2384 vdd.n2383 185
R16223 vdd.n2386 vdd.n2385 185
R16224 vdd.n2388 vdd.n2387 185
R16225 vdd.n2390 vdd.n2389 185
R16226 vdd.n2392 vdd.n2391 185
R16227 vdd.n2394 vdd.n2393 185
R16228 vdd.n2396 vdd.n2395 185
R16229 vdd.n2398 vdd.n2397 185
R16230 vdd.n2400 vdd.n2399 185
R16231 vdd.n2402 vdd.n2401 185
R16232 vdd.n2404 vdd.n2403 185
R16233 vdd.n2406 vdd.n2405 185
R16234 vdd.n2408 vdd.n2407 185
R16235 vdd.n2410 vdd.n2409 185
R16236 vdd.n2412 vdd.n2411 185
R16237 vdd.n2414 vdd.n2413 185
R16238 vdd.n2416 vdd.n2415 185
R16239 vdd.n2418 vdd.n2417 185
R16240 vdd.n2420 vdd.n2419 185
R16241 vdd.n2421 vdd.n836 185
R16242 vdd.n2353 vdd.n834 185
R16243 vdd.n2424 vdd.n834 185
R16244 vdd.n2352 vdd.n2351 185
R16245 vdd.n2351 vdd.n833 185
R16246 vdd.n2350 vdd.n841 185
R16247 vdd.n2350 vdd.n2349 185
R16248 vdd.n1243 vdd.n842 185
R16249 vdd.n1227 vdd.n842 185
R16250 vdd.n1244 vdd.n851 185
R16251 vdd.n2342 vdd.n851 185
R16252 vdd.n1246 vdd.n1245 185
R16253 vdd.n1245 vdd.n849 185
R16254 vdd.n1247 vdd.n858 185
R16255 vdd.n2334 vdd.n858 185
R16256 vdd.n1249 vdd.n1248 185
R16257 vdd.n1248 vdd.n856 185
R16258 vdd.n1250 vdd.n863 185
R16259 vdd.n2328 vdd.n863 185
R16260 vdd.n1252 vdd.n1251 185
R16261 vdd.n1253 vdd.n1252 185
R16262 vdd.n1242 vdd.n868 185
R16263 vdd.n2322 vdd.n868 185
R16264 vdd.n1241 vdd.n1240 185
R16265 vdd.n1240 vdd.n874 185
R16266 vdd.n1239 vdd.n873 185
R16267 vdd.n2316 vdd.n873 185
R16268 vdd.n1238 vdd.n1237 185
R16269 vdd.n1237 vdd.n880 185
R16270 vdd.n1146 vdd.n879 185
R16271 vdd.n2310 vdd.n879 185
R16272 vdd.n1267 vdd.n1266 185
R16273 vdd.n1266 vdd.n1265 185
R16274 vdd.n1268 vdd.n886 185
R16275 vdd.n2304 vdd.n886 185
R16276 vdd.n1270 vdd.n1269 185
R16277 vdd.n1269 vdd.n884 185
R16278 vdd.n1271 vdd.n892 185
R16279 vdd.n2298 vdd.n892 185
R16280 vdd.n1273 vdd.n1272 185
R16281 vdd.n1272 vdd.n890 185
R16282 vdd.n1274 vdd.n897 185
R16283 vdd.n2292 vdd.n897 185
R16284 vdd.n1276 vdd.n1275 185
R16285 vdd.n1275 vdd.n904 185
R16286 vdd.n1277 vdd.n903 185
R16287 vdd.n2285 vdd.n903 185
R16288 vdd.n1279 vdd.n1278 185
R16289 vdd.n1278 vdd.n911 185
R16290 vdd.n1280 vdd.n910 185
R16291 vdd.n2279 vdd.n910 185
R16292 vdd.n1282 vdd.n1281 185
R16293 vdd.n1281 vdd.n908 185
R16294 vdd.n1283 vdd.n917 185
R16295 vdd.n2273 vdd.n917 185
R16296 vdd.n1285 vdd.n1284 185
R16297 vdd.n1284 vdd.n915 185
R16298 vdd.n1286 vdd.n923 185
R16299 vdd.n2267 vdd.n923 185
R16300 vdd.n1288 vdd.n1287 185
R16301 vdd.n1287 vdd.n921 185
R16302 vdd.n1289 vdd.n928 185
R16303 vdd.n2261 vdd.n928 185
R16304 vdd.n1291 vdd.n1290 185
R16305 vdd.n1290 vdd.n934 185
R16306 vdd.n1292 vdd.n933 185
R16307 vdd.n2255 vdd.n933 185
R16308 vdd.n1294 vdd.n1293 185
R16309 vdd.n1293 vdd.n940 185
R16310 vdd.n1295 vdd.n939 185
R16311 vdd.n2249 vdd.n939 185
R16312 vdd.n1297 vdd.n1296 185
R16313 vdd.n1296 vdd.n947 185
R16314 vdd.n1298 vdd.n946 185
R16315 vdd.n2243 vdd.n946 185
R16316 vdd.n1300 vdd.n1299 185
R16317 vdd.n1299 vdd.n944 185
R16318 vdd.n1301 vdd.n953 185
R16319 vdd.n2237 vdd.n953 185
R16320 vdd.n1303 vdd.n1302 185
R16321 vdd.n1302 vdd.n951 185
R16322 vdd.n1304 vdd.n958 185
R16323 vdd.n2231 vdd.n958 185
R16324 vdd.n1306 vdd.n1305 185
R16325 vdd.n1305 vdd.n965 185
R16326 vdd.n1307 vdd.n964 185
R16327 vdd.n2225 vdd.n964 185
R16328 vdd.n1309 vdd.n1308 185
R16329 vdd.n1308 vdd.n962 185
R16330 vdd.n1109 vdd.n1108 185
R16331 vdd.n1111 vdd.n1110 185
R16332 vdd.n1113 vdd.n1112 185
R16333 vdd.n1115 vdd.n1114 185
R16334 vdd.n1117 vdd.n1116 185
R16335 vdd.n1119 vdd.n1118 185
R16336 vdd.n1121 vdd.n1120 185
R16337 vdd.n1123 vdd.n1122 185
R16338 vdd.n1125 vdd.n1124 185
R16339 vdd.n1127 vdd.n1126 185
R16340 vdd.n1129 vdd.n1128 185
R16341 vdd.n1131 vdd.n1130 185
R16342 vdd.n1133 vdd.n1132 185
R16343 vdd.n1135 vdd.n1134 185
R16344 vdd.n1137 vdd.n1136 185
R16345 vdd.n1139 vdd.n1138 185
R16346 vdd.n1141 vdd.n1140 185
R16347 vdd.n1343 vdd.n1142 185
R16348 vdd.n1342 vdd.n1341 185
R16349 vdd.n1340 vdd.n1339 185
R16350 vdd.n1338 vdd.n1337 185
R16351 vdd.n1336 vdd.n1335 185
R16352 vdd.n1334 vdd.n1333 185
R16353 vdd.n1332 vdd.n1331 185
R16354 vdd.n1330 vdd.n1329 185
R16355 vdd.n1328 vdd.n1327 185
R16356 vdd.n1326 vdd.n1325 185
R16357 vdd.n1324 vdd.n1323 185
R16358 vdd.n1322 vdd.n1321 185
R16359 vdd.n1320 vdd.n1319 185
R16360 vdd.n1318 vdd.n1317 185
R16361 vdd.n1316 vdd.n1315 185
R16362 vdd.n1314 vdd.n1313 185
R16363 vdd.n1312 vdd.n1311 185
R16364 vdd.n1310 vdd.n1003 185
R16365 vdd.n2218 vdd.n1003 185
R16366 vdd.n303 vdd.n302 171.744
R16367 vdd.n302 vdd.n301 171.744
R16368 vdd.n301 vdd.n270 171.744
R16369 vdd.n294 vdd.n270 171.744
R16370 vdd.n294 vdd.n293 171.744
R16371 vdd.n293 vdd.n275 171.744
R16372 vdd.n286 vdd.n275 171.744
R16373 vdd.n286 vdd.n285 171.744
R16374 vdd.n285 vdd.n279 171.744
R16375 vdd.n252 vdd.n251 171.744
R16376 vdd.n251 vdd.n250 171.744
R16377 vdd.n250 vdd.n219 171.744
R16378 vdd.n243 vdd.n219 171.744
R16379 vdd.n243 vdd.n242 171.744
R16380 vdd.n242 vdd.n224 171.744
R16381 vdd.n235 vdd.n224 171.744
R16382 vdd.n235 vdd.n234 171.744
R16383 vdd.n234 vdd.n228 171.744
R16384 vdd.n209 vdd.n208 171.744
R16385 vdd.n208 vdd.n207 171.744
R16386 vdd.n207 vdd.n176 171.744
R16387 vdd.n200 vdd.n176 171.744
R16388 vdd.n200 vdd.n199 171.744
R16389 vdd.n199 vdd.n181 171.744
R16390 vdd.n192 vdd.n181 171.744
R16391 vdd.n192 vdd.n191 171.744
R16392 vdd.n191 vdd.n185 171.744
R16393 vdd.n158 vdd.n157 171.744
R16394 vdd.n157 vdd.n156 171.744
R16395 vdd.n156 vdd.n125 171.744
R16396 vdd.n149 vdd.n125 171.744
R16397 vdd.n149 vdd.n148 171.744
R16398 vdd.n148 vdd.n130 171.744
R16399 vdd.n141 vdd.n130 171.744
R16400 vdd.n141 vdd.n140 171.744
R16401 vdd.n140 vdd.n134 171.744
R16402 vdd.n116 vdd.n115 171.744
R16403 vdd.n115 vdd.n114 171.744
R16404 vdd.n114 vdd.n83 171.744
R16405 vdd.n107 vdd.n83 171.744
R16406 vdd.n107 vdd.n106 171.744
R16407 vdd.n106 vdd.n88 171.744
R16408 vdd.n99 vdd.n88 171.744
R16409 vdd.n99 vdd.n98 171.744
R16410 vdd.n98 vdd.n92 171.744
R16411 vdd.n65 vdd.n64 171.744
R16412 vdd.n64 vdd.n63 171.744
R16413 vdd.n63 vdd.n32 171.744
R16414 vdd.n56 vdd.n32 171.744
R16415 vdd.n56 vdd.n55 171.744
R16416 vdd.n55 vdd.n37 171.744
R16417 vdd.n48 vdd.n37 171.744
R16418 vdd.n48 vdd.n47 171.744
R16419 vdd.n47 vdd.n41 171.744
R16420 vdd.n1953 vdd.n1952 171.744
R16421 vdd.n1952 vdd.n1951 171.744
R16422 vdd.n1951 vdd.n1920 171.744
R16423 vdd.n1944 vdd.n1920 171.744
R16424 vdd.n1944 vdd.n1943 171.744
R16425 vdd.n1943 vdd.n1925 171.744
R16426 vdd.n1936 vdd.n1925 171.744
R16427 vdd.n1936 vdd.n1935 171.744
R16428 vdd.n1935 vdd.n1929 171.744
R16429 vdd.n2004 vdd.n2003 171.744
R16430 vdd.n2003 vdd.n2002 171.744
R16431 vdd.n2002 vdd.n1971 171.744
R16432 vdd.n1995 vdd.n1971 171.744
R16433 vdd.n1995 vdd.n1994 171.744
R16434 vdd.n1994 vdd.n1976 171.744
R16435 vdd.n1987 vdd.n1976 171.744
R16436 vdd.n1987 vdd.n1986 171.744
R16437 vdd.n1986 vdd.n1980 171.744
R16438 vdd.n1859 vdd.n1858 171.744
R16439 vdd.n1858 vdd.n1857 171.744
R16440 vdd.n1857 vdd.n1826 171.744
R16441 vdd.n1850 vdd.n1826 171.744
R16442 vdd.n1850 vdd.n1849 171.744
R16443 vdd.n1849 vdd.n1831 171.744
R16444 vdd.n1842 vdd.n1831 171.744
R16445 vdd.n1842 vdd.n1841 171.744
R16446 vdd.n1841 vdd.n1835 171.744
R16447 vdd.n1910 vdd.n1909 171.744
R16448 vdd.n1909 vdd.n1908 171.744
R16449 vdd.n1908 vdd.n1877 171.744
R16450 vdd.n1901 vdd.n1877 171.744
R16451 vdd.n1901 vdd.n1900 171.744
R16452 vdd.n1900 vdd.n1882 171.744
R16453 vdd.n1893 vdd.n1882 171.744
R16454 vdd.n1893 vdd.n1892 171.744
R16455 vdd.n1892 vdd.n1886 171.744
R16456 vdd.n1766 vdd.n1765 171.744
R16457 vdd.n1765 vdd.n1764 171.744
R16458 vdd.n1764 vdd.n1733 171.744
R16459 vdd.n1757 vdd.n1733 171.744
R16460 vdd.n1757 vdd.n1756 171.744
R16461 vdd.n1756 vdd.n1738 171.744
R16462 vdd.n1749 vdd.n1738 171.744
R16463 vdd.n1749 vdd.n1748 171.744
R16464 vdd.n1748 vdd.n1742 171.744
R16465 vdd.n1817 vdd.n1816 171.744
R16466 vdd.n1816 vdd.n1815 171.744
R16467 vdd.n1815 vdd.n1784 171.744
R16468 vdd.n1808 vdd.n1784 171.744
R16469 vdd.n1808 vdd.n1807 171.744
R16470 vdd.n1807 vdd.n1789 171.744
R16471 vdd.n1800 vdd.n1789 171.744
R16472 vdd.n1800 vdd.n1799 171.744
R16473 vdd.n1799 vdd.n1793 171.744
R16474 vdd.n3402 vdd.n356 146.341
R16475 vdd.n3400 vdd.n3399 146.341
R16476 vdd.n3397 vdd.n360 146.341
R16477 vdd.n3393 vdd.n3392 146.341
R16478 vdd.n3390 vdd.n368 146.341
R16479 vdd.n3386 vdd.n3385 146.341
R16480 vdd.n3383 vdd.n375 146.341
R16481 vdd.n3379 vdd.n3378 146.341
R16482 vdd.n3376 vdd.n382 146.341
R16483 vdd.n393 vdd.n390 146.341
R16484 vdd.n3368 vdd.n3367 146.341
R16485 vdd.n3365 vdd.n395 146.341
R16486 vdd.n3361 vdd.n3360 146.341
R16487 vdd.n3358 vdd.n401 146.341
R16488 vdd.n3354 vdd.n3353 146.341
R16489 vdd.n3351 vdd.n408 146.341
R16490 vdd.n3347 vdd.n3346 146.341
R16491 vdd.n3344 vdd.n415 146.341
R16492 vdd.n3340 vdd.n3339 146.341
R16493 vdd.n3337 vdd.n422 146.341
R16494 vdd.n433 vdd.n430 146.341
R16495 vdd.n3329 vdd.n3328 146.341
R16496 vdd.n3326 vdd.n435 146.341
R16497 vdd.n3322 vdd.n3321 146.341
R16498 vdd.n3319 vdd.n441 146.341
R16499 vdd.n3315 vdd.n3314 146.341
R16500 vdd.n3312 vdd.n448 146.341
R16501 vdd.n3308 vdd.n3307 146.341
R16502 vdd.n3305 vdd.n455 146.341
R16503 vdd.n3301 vdd.n3300 146.341
R16504 vdd.n3298 vdd.n462 146.341
R16505 vdd.n3213 vdd.n512 146.341
R16506 vdd.n3219 vdd.n512 146.341
R16507 vdd.n3219 vdd.n504 146.341
R16508 vdd.n3229 vdd.n504 146.341
R16509 vdd.n3229 vdd.n500 146.341
R16510 vdd.n3235 vdd.n500 146.341
R16511 vdd.n3235 vdd.n491 146.341
R16512 vdd.n3245 vdd.n491 146.341
R16513 vdd.n3245 vdd.n487 146.341
R16514 vdd.n3251 vdd.n487 146.341
R16515 vdd.n3251 vdd.n479 146.341
R16516 vdd.n3262 vdd.n479 146.341
R16517 vdd.n3262 vdd.n480 146.341
R16518 vdd.n480 vdd.n316 146.341
R16519 vdd.n317 vdd.n316 146.341
R16520 vdd.n318 vdd.n317 146.341
R16521 vdd.n473 vdd.n318 146.341
R16522 vdd.n473 vdd.n326 146.341
R16523 vdd.n327 vdd.n326 146.341
R16524 vdd.n328 vdd.n327 146.341
R16525 vdd.n470 vdd.n328 146.341
R16526 vdd.n470 vdd.n337 146.341
R16527 vdd.n338 vdd.n337 146.341
R16528 vdd.n339 vdd.n338 146.341
R16529 vdd.n467 vdd.n339 146.341
R16530 vdd.n467 vdd.n348 146.341
R16531 vdd.n349 vdd.n348 146.341
R16532 vdd.n350 vdd.n349 146.341
R16533 vdd.n3205 vdd.n3203 146.341
R16534 vdd.n3203 vdd.n3202 146.341
R16535 vdd.n3199 vdd.n3198 146.341
R16536 vdd.n3195 vdd.n3194 146.341
R16537 vdd.n3192 vdd.n526 146.341
R16538 vdd.n3188 vdd.n3186 146.341
R16539 vdd.n3184 vdd.n532 146.341
R16540 vdd.n3180 vdd.n3178 146.341
R16541 vdd.n3176 vdd.n538 146.341
R16542 vdd.n3172 vdd.n3170 146.341
R16543 vdd.n3168 vdd.n546 146.341
R16544 vdd.n3164 vdd.n3162 146.341
R16545 vdd.n3160 vdd.n552 146.341
R16546 vdd.n3156 vdd.n3154 146.341
R16547 vdd.n3152 vdd.n558 146.341
R16548 vdd.n3148 vdd.n3146 146.341
R16549 vdd.n3144 vdd.n564 146.341
R16550 vdd.n3140 vdd.n3138 146.341
R16551 vdd.n3136 vdd.n570 146.341
R16552 vdd.n3132 vdd.n3130 146.341
R16553 vdd.n3128 vdd.n576 146.341
R16554 vdd.n3121 vdd.n585 146.341
R16555 vdd.n3119 vdd.n3118 146.341
R16556 vdd.n3115 vdd.n3114 146.341
R16557 vdd.n3112 vdd.n590 146.341
R16558 vdd.n3108 vdd.n3106 146.341
R16559 vdd.n3104 vdd.n596 146.341
R16560 vdd.n3100 vdd.n3098 146.341
R16561 vdd.n3096 vdd.n602 146.341
R16562 vdd.n3092 vdd.n3090 146.341
R16563 vdd.n3087 vdd.n3086 146.341
R16564 vdd.n3083 vdd.n515 146.341
R16565 vdd.n3211 vdd.n510 146.341
R16566 vdd.n3221 vdd.n510 146.341
R16567 vdd.n3221 vdd.n506 146.341
R16568 vdd.n3227 vdd.n506 146.341
R16569 vdd.n3227 vdd.n498 146.341
R16570 vdd.n3237 vdd.n498 146.341
R16571 vdd.n3237 vdd.n494 146.341
R16572 vdd.n3243 vdd.n494 146.341
R16573 vdd.n3243 vdd.n486 146.341
R16574 vdd.n3254 vdd.n486 146.341
R16575 vdd.n3254 vdd.n482 146.341
R16576 vdd.n3260 vdd.n482 146.341
R16577 vdd.n3260 vdd.n314 146.341
R16578 vdd.n3437 vdd.n314 146.341
R16579 vdd.n3437 vdd.n315 146.341
R16580 vdd.n3433 vdd.n315 146.341
R16581 vdd.n3433 vdd.n319 146.341
R16582 vdd.n3429 vdd.n319 146.341
R16583 vdd.n3429 vdd.n324 146.341
R16584 vdd.n3425 vdd.n324 146.341
R16585 vdd.n3425 vdd.n330 146.341
R16586 vdd.n3421 vdd.n330 146.341
R16587 vdd.n3421 vdd.n336 146.341
R16588 vdd.n3417 vdd.n336 146.341
R16589 vdd.n3417 vdd.n341 146.341
R16590 vdd.n3413 vdd.n341 146.341
R16591 vdd.n3413 vdd.n347 146.341
R16592 vdd.n3409 vdd.n347 146.341
R16593 vdd.n2183 vdd.n2182 146.341
R16594 vdd.n2180 vdd.n2177 146.341
R16595 vdd.n2175 vdd.n1013 146.341
R16596 vdd.n2171 vdd.n2170 146.341
R16597 vdd.n2168 vdd.n1017 146.341
R16598 vdd.n2164 vdd.n2163 146.341
R16599 vdd.n2161 vdd.n1024 146.341
R16600 vdd.n2157 vdd.n2156 146.341
R16601 vdd.n2154 vdd.n1031 146.341
R16602 vdd.n1042 vdd.n1039 146.341
R16603 vdd.n2146 vdd.n2145 146.341
R16604 vdd.n2143 vdd.n1044 146.341
R16605 vdd.n2139 vdd.n2138 146.341
R16606 vdd.n2136 vdd.n1050 146.341
R16607 vdd.n2132 vdd.n2131 146.341
R16608 vdd.n2129 vdd.n1057 146.341
R16609 vdd.n2125 vdd.n2124 146.341
R16610 vdd.n2122 vdd.n1064 146.341
R16611 vdd.n2118 vdd.n2117 146.341
R16612 vdd.n2115 vdd.n1071 146.341
R16613 vdd.n1082 vdd.n1079 146.341
R16614 vdd.n2107 vdd.n2106 146.341
R16615 vdd.n2104 vdd.n1084 146.341
R16616 vdd.n2100 vdd.n2099 146.341
R16617 vdd.n2097 vdd.n1090 146.341
R16618 vdd.n2093 vdd.n2092 146.341
R16619 vdd.n2090 vdd.n1097 146.341
R16620 vdd.n2086 vdd.n2085 146.341
R16621 vdd.n2083 vdd.n1104 146.341
R16622 vdd.n1350 vdd.n1348 146.341
R16623 vdd.n1353 vdd.n1352 146.341
R16624 vdd.n1671 vdd.n1433 146.341
R16625 vdd.n1677 vdd.n1433 146.341
R16626 vdd.n1677 vdd.n1426 146.341
R16627 vdd.n1687 vdd.n1426 146.341
R16628 vdd.n1687 vdd.n1422 146.341
R16629 vdd.n1693 vdd.n1422 146.341
R16630 vdd.n1693 vdd.n1413 146.341
R16631 vdd.n1703 vdd.n1413 146.341
R16632 vdd.n1703 vdd.n1409 146.341
R16633 vdd.n1709 vdd.n1409 146.341
R16634 vdd.n1709 vdd.n1402 146.341
R16635 vdd.n1720 vdd.n1402 146.341
R16636 vdd.n1720 vdd.n1398 146.341
R16637 vdd.n1726 vdd.n1398 146.341
R16638 vdd.n1726 vdd.n1391 146.341
R16639 vdd.n2018 vdd.n1391 146.341
R16640 vdd.n2018 vdd.n1387 146.341
R16641 vdd.n2024 vdd.n1387 146.341
R16642 vdd.n2024 vdd.n1379 146.341
R16643 vdd.n2035 vdd.n1379 146.341
R16644 vdd.n2035 vdd.n1375 146.341
R16645 vdd.n2041 vdd.n1375 146.341
R16646 vdd.n2041 vdd.n1369 146.341
R16647 vdd.n2052 vdd.n1369 146.341
R16648 vdd.n2052 vdd.n1364 146.341
R16649 vdd.n2060 vdd.n1364 146.341
R16650 vdd.n2060 vdd.n1355 146.341
R16651 vdd.n2071 vdd.n1355 146.341
R16652 vdd.n1443 vdd.n1442 146.341
R16653 vdd.n1446 vdd.n1443 146.341
R16654 vdd.n1449 vdd.n1448 146.341
R16655 vdd.n1454 vdd.n1451 146.341
R16656 vdd.n1457 vdd.n1456 146.341
R16657 vdd.n1462 vdd.n1459 146.341
R16658 vdd.n1465 vdd.n1464 146.341
R16659 vdd.n1470 vdd.n1467 146.341
R16660 vdd.n1473 vdd.n1472 146.341
R16661 vdd.n1480 vdd.n1475 146.341
R16662 vdd.n1483 vdd.n1482 146.341
R16663 vdd.n1488 vdd.n1485 146.341
R16664 vdd.n1491 vdd.n1490 146.341
R16665 vdd.n1496 vdd.n1493 146.341
R16666 vdd.n1499 vdd.n1498 146.341
R16667 vdd.n1504 vdd.n1501 146.341
R16668 vdd.n1507 vdd.n1506 146.341
R16669 vdd.n1512 vdd.n1509 146.341
R16670 vdd.n1515 vdd.n1514 146.341
R16671 vdd.n1520 vdd.n1517 146.341
R16672 vdd.n1601 vdd.n1522 146.341
R16673 vdd.n1599 vdd.n1598 146.341
R16674 vdd.n1529 vdd.n1528 146.341
R16675 vdd.n1532 vdd.n1531 146.341
R16676 vdd.n1537 vdd.n1536 146.341
R16677 vdd.n1540 vdd.n1539 146.341
R16678 vdd.n1545 vdd.n1544 146.341
R16679 vdd.n1548 vdd.n1547 146.341
R16680 vdd.n1553 vdd.n1552 146.341
R16681 vdd.n1556 vdd.n1555 146.341
R16682 vdd.n1561 vdd.n1560 146.341
R16683 vdd.n1563 vdd.n1436 146.341
R16684 vdd.n1669 vdd.n1432 146.341
R16685 vdd.n1679 vdd.n1432 146.341
R16686 vdd.n1679 vdd.n1428 146.341
R16687 vdd.n1685 vdd.n1428 146.341
R16688 vdd.n1685 vdd.n1420 146.341
R16689 vdd.n1695 vdd.n1420 146.341
R16690 vdd.n1695 vdd.n1416 146.341
R16691 vdd.n1701 vdd.n1416 146.341
R16692 vdd.n1701 vdd.n1408 146.341
R16693 vdd.n1712 vdd.n1408 146.341
R16694 vdd.n1712 vdd.n1404 146.341
R16695 vdd.n1718 vdd.n1404 146.341
R16696 vdd.n1718 vdd.n1397 146.341
R16697 vdd.n1728 vdd.n1397 146.341
R16698 vdd.n1728 vdd.n1393 146.341
R16699 vdd.n2016 vdd.n1393 146.341
R16700 vdd.n2016 vdd.n1385 146.341
R16701 vdd.n2027 vdd.n1385 146.341
R16702 vdd.n2027 vdd.n1381 146.341
R16703 vdd.n2033 vdd.n1381 146.341
R16704 vdd.n2033 vdd.n1374 146.341
R16705 vdd.n2044 vdd.n1374 146.341
R16706 vdd.n2044 vdd.n1370 146.341
R16707 vdd.n2050 vdd.n1370 146.341
R16708 vdd.n2050 vdd.n1362 146.341
R16709 vdd.n2063 vdd.n1362 146.341
R16710 vdd.n2063 vdd.n1357 146.341
R16711 vdd.n2069 vdd.n1357 146.341
R16712 vdd.n1143 vdd.t17 127.284
R16713 vdd.n838 vdd.t61 127.284
R16714 vdd.n1147 vdd.t58 127.284
R16715 vdd.n829 vdd.t84 127.284
R16716 vdd.n724 vdd.t38 127.284
R16717 vdd.n724 vdd.t39 127.284
R16718 vdd.n2535 vdd.t79 127.284
R16719 vdd.n661 vdd.t26 127.284
R16720 vdd.n2532 vdd.t69 127.284
R16721 vdd.n625 vdd.t12 127.284
R16722 vdd.n899 vdd.t75 127.284
R16723 vdd.n899 vdd.t76 127.284
R16724 vdd.n22 vdd.n20 117.314
R16725 vdd.n17 vdd.n15 117.314
R16726 vdd.n27 vdd.n26 116.927
R16727 vdd.n24 vdd.n23 116.927
R16728 vdd.n22 vdd.n21 116.927
R16729 vdd.n17 vdd.n16 116.927
R16730 vdd.n19 vdd.n18 116.927
R16731 vdd.n27 vdd.n25 116.927
R16732 vdd.n1144 vdd.t16 111.188
R16733 vdd.n839 vdd.t62 111.188
R16734 vdd.n1148 vdd.t57 111.188
R16735 vdd.n830 vdd.t85 111.188
R16736 vdd.n2536 vdd.t78 111.188
R16737 vdd.n662 vdd.t27 111.188
R16738 vdd.n2533 vdd.t68 111.188
R16739 vdd.n626 vdd.t13 111.188
R16740 vdd.n2806 vdd.n788 99.5127
R16741 vdd.n2806 vdd.n779 99.5127
R16742 vdd.n2814 vdd.n779 99.5127
R16743 vdd.n2814 vdd.n777 99.5127
R16744 vdd.n2818 vdd.n777 99.5127
R16745 vdd.n2818 vdd.n767 99.5127
R16746 vdd.n2826 vdd.n767 99.5127
R16747 vdd.n2826 vdd.n765 99.5127
R16748 vdd.n2830 vdd.n765 99.5127
R16749 vdd.n2830 vdd.n756 99.5127
R16750 vdd.n2838 vdd.n756 99.5127
R16751 vdd.n2838 vdd.n754 99.5127
R16752 vdd.n2842 vdd.n754 99.5127
R16753 vdd.n2842 vdd.n745 99.5127
R16754 vdd.n2850 vdd.n745 99.5127
R16755 vdd.n2850 vdd.n743 99.5127
R16756 vdd.n2854 vdd.n743 99.5127
R16757 vdd.n2854 vdd.n732 99.5127
R16758 vdd.n2863 vdd.n732 99.5127
R16759 vdd.n2863 vdd.n730 99.5127
R16760 vdd.n2867 vdd.n730 99.5127
R16761 vdd.n2867 vdd.n720 99.5127
R16762 vdd.n2875 vdd.n720 99.5127
R16763 vdd.n2875 vdd.n718 99.5127
R16764 vdd.n2879 vdd.n718 99.5127
R16765 vdd.n2879 vdd.n708 99.5127
R16766 vdd.n2887 vdd.n708 99.5127
R16767 vdd.n2887 vdd.n706 99.5127
R16768 vdd.n2891 vdd.n706 99.5127
R16769 vdd.n2891 vdd.n695 99.5127
R16770 vdd.n2899 vdd.n695 99.5127
R16771 vdd.n2899 vdd.n693 99.5127
R16772 vdd.n2903 vdd.n693 99.5127
R16773 vdd.n2903 vdd.n684 99.5127
R16774 vdd.n2911 vdd.n684 99.5127
R16775 vdd.n2911 vdd.n682 99.5127
R16776 vdd.n2915 vdd.n682 99.5127
R16777 vdd.n2915 vdd.n670 99.5127
R16778 vdd.n2968 vdd.n670 99.5127
R16779 vdd.n2968 vdd.n668 99.5127
R16780 vdd.n2972 vdd.n668 99.5127
R16781 vdd.n2972 vdd.n634 99.5127
R16782 vdd.n3042 vdd.n634 99.5127
R16783 vdd.n3038 vdd.n635 99.5127
R16784 vdd.n3036 vdd.n3035 99.5127
R16785 vdd.n3033 vdd.n639 99.5127
R16786 vdd.n3029 vdd.n3028 99.5127
R16787 vdd.n3026 vdd.n642 99.5127
R16788 vdd.n3022 vdd.n3021 99.5127
R16789 vdd.n3019 vdd.n645 99.5127
R16790 vdd.n3015 vdd.n3014 99.5127
R16791 vdd.n3012 vdd.n648 99.5127
R16792 vdd.n3007 vdd.n3006 99.5127
R16793 vdd.n3004 vdd.n651 99.5127
R16794 vdd.n3000 vdd.n2999 99.5127
R16795 vdd.n2997 vdd.n654 99.5127
R16796 vdd.n2993 vdd.n2992 99.5127
R16797 vdd.n2990 vdd.n657 99.5127
R16798 vdd.n2986 vdd.n2985 99.5127
R16799 vdd.n2983 vdd.n660 99.5127
R16800 vdd.n2733 vdd.n786 99.5127
R16801 vdd.n2729 vdd.n786 99.5127
R16802 vdd.n2729 vdd.n780 99.5127
R16803 vdd.n2611 vdd.n780 99.5127
R16804 vdd.n2611 vdd.n775 99.5127
R16805 vdd.n2614 vdd.n775 99.5127
R16806 vdd.n2614 vdd.n769 99.5127
R16807 vdd.n2715 vdd.n769 99.5127
R16808 vdd.n2715 vdd.n763 99.5127
R16809 vdd.n2711 vdd.n763 99.5127
R16810 vdd.n2711 vdd.n757 99.5127
R16811 vdd.n2658 vdd.n757 99.5127
R16812 vdd.n2658 vdd.n751 99.5127
R16813 vdd.n2655 vdd.n751 99.5127
R16814 vdd.n2655 vdd.n746 99.5127
R16815 vdd.n2652 vdd.n746 99.5127
R16816 vdd.n2652 vdd.n741 99.5127
R16817 vdd.n2649 vdd.n741 99.5127
R16818 vdd.n2649 vdd.n734 99.5127
R16819 vdd.n2646 vdd.n734 99.5127
R16820 vdd.n2646 vdd.n727 99.5127
R16821 vdd.n2643 vdd.n727 99.5127
R16822 vdd.n2643 vdd.n721 99.5127
R16823 vdd.n2640 vdd.n721 99.5127
R16824 vdd.n2640 vdd.n716 99.5127
R16825 vdd.n2637 vdd.n716 99.5127
R16826 vdd.n2637 vdd.n710 99.5127
R16827 vdd.n2634 vdd.n710 99.5127
R16828 vdd.n2634 vdd.n703 99.5127
R16829 vdd.n2631 vdd.n703 99.5127
R16830 vdd.n2631 vdd.n696 99.5127
R16831 vdd.n2628 vdd.n696 99.5127
R16832 vdd.n2628 vdd.n690 99.5127
R16833 vdd.n2625 vdd.n690 99.5127
R16834 vdd.n2625 vdd.n685 99.5127
R16835 vdd.n2622 vdd.n685 99.5127
R16836 vdd.n2622 vdd.n680 99.5127
R16837 vdd.n2619 vdd.n680 99.5127
R16838 vdd.n2619 vdd.n672 99.5127
R16839 vdd.n672 vdd.n665 99.5127
R16840 vdd.n2974 vdd.n665 99.5127
R16841 vdd.n2975 vdd.n2974 99.5127
R16842 vdd.n2975 vdd.n632 99.5127
R16843 vdd.n2799 vdd.n790 99.5127
R16844 vdd.n2799 vdd.n2531 99.5127
R16845 vdd.n2795 vdd.n2794 99.5127
R16846 vdd.n2791 vdd.n2790 99.5127
R16847 vdd.n2787 vdd.n2786 99.5127
R16848 vdd.n2783 vdd.n2782 99.5127
R16849 vdd.n2779 vdd.n2778 99.5127
R16850 vdd.n2775 vdd.n2774 99.5127
R16851 vdd.n2771 vdd.n2770 99.5127
R16852 vdd.n2767 vdd.n2766 99.5127
R16853 vdd.n2763 vdd.n2762 99.5127
R16854 vdd.n2759 vdd.n2758 99.5127
R16855 vdd.n2755 vdd.n2754 99.5127
R16856 vdd.n2751 vdd.n2750 99.5127
R16857 vdd.n2747 vdd.n2746 99.5127
R16858 vdd.n2743 vdd.n2742 99.5127
R16859 vdd.n2738 vdd.n2737 99.5127
R16860 vdd.n2495 vdd.n827 99.5127
R16861 vdd.n2491 vdd.n2490 99.5127
R16862 vdd.n2487 vdd.n2486 99.5127
R16863 vdd.n2483 vdd.n2482 99.5127
R16864 vdd.n2479 vdd.n2478 99.5127
R16865 vdd.n2475 vdd.n2474 99.5127
R16866 vdd.n2471 vdd.n2470 99.5127
R16867 vdd.n2467 vdd.n2466 99.5127
R16868 vdd.n2463 vdd.n2462 99.5127
R16869 vdd.n2459 vdd.n2458 99.5127
R16870 vdd.n2455 vdd.n2454 99.5127
R16871 vdd.n2451 vdd.n2450 99.5127
R16872 vdd.n2447 vdd.n2446 99.5127
R16873 vdd.n2443 vdd.n2442 99.5127
R16874 vdd.n2439 vdd.n2438 99.5127
R16875 vdd.n2435 vdd.n2434 99.5127
R16876 vdd.n2430 vdd.n2429 99.5127
R16877 vdd.n1183 vdd.n963 99.5127
R16878 vdd.n1186 vdd.n963 99.5127
R16879 vdd.n1186 vdd.n957 99.5127
R16880 vdd.n1189 vdd.n957 99.5127
R16881 vdd.n1189 vdd.n952 99.5127
R16882 vdd.n1192 vdd.n952 99.5127
R16883 vdd.n1192 vdd.n945 99.5127
R16884 vdd.n1195 vdd.n945 99.5127
R16885 vdd.n1195 vdd.n938 99.5127
R16886 vdd.n1198 vdd.n938 99.5127
R16887 vdd.n1198 vdd.n932 99.5127
R16888 vdd.n1201 vdd.n932 99.5127
R16889 vdd.n1201 vdd.n927 99.5127
R16890 vdd.n1204 vdd.n927 99.5127
R16891 vdd.n1204 vdd.n922 99.5127
R16892 vdd.n1207 vdd.n922 99.5127
R16893 vdd.n1207 vdd.n916 99.5127
R16894 vdd.n1210 vdd.n916 99.5127
R16895 vdd.n1210 vdd.n909 99.5127
R16896 vdd.n1213 vdd.n909 99.5127
R16897 vdd.n1213 vdd.n902 99.5127
R16898 vdd.n1216 vdd.n902 99.5127
R16899 vdd.n1216 vdd.n896 99.5127
R16900 vdd.n1219 vdd.n896 99.5127
R16901 vdd.n1219 vdd.n891 99.5127
R16902 vdd.n1222 vdd.n891 99.5127
R16903 vdd.n1222 vdd.n885 99.5127
R16904 vdd.n1264 vdd.n885 99.5127
R16905 vdd.n1264 vdd.n878 99.5127
R16906 vdd.n1260 vdd.n878 99.5127
R16907 vdd.n1260 vdd.n872 99.5127
R16908 vdd.n1257 vdd.n872 99.5127
R16909 vdd.n1257 vdd.n867 99.5127
R16910 vdd.n1254 vdd.n867 99.5127
R16911 vdd.n1254 vdd.n862 99.5127
R16912 vdd.n1234 vdd.n862 99.5127
R16913 vdd.n1234 vdd.n857 99.5127
R16914 vdd.n1231 vdd.n857 99.5127
R16915 vdd.n1231 vdd.n850 99.5127
R16916 vdd.n1228 vdd.n850 99.5127
R16917 vdd.n1228 vdd.n843 99.5127
R16918 vdd.n843 vdd.n832 99.5127
R16919 vdd.n2425 vdd.n832 99.5127
R16920 vdd.n2217 vdd.n968 99.5127
R16921 vdd.n2217 vdd.n1004 99.5127
R16922 vdd.n2213 vdd.n2212 99.5127
R16923 vdd.n2209 vdd.n2208 99.5127
R16924 vdd.n2205 vdd.n2204 99.5127
R16925 vdd.n2201 vdd.n2200 99.5127
R16926 vdd.n2197 vdd.n2196 99.5127
R16927 vdd.n2193 vdd.n2192 99.5127
R16928 vdd.n2189 vdd.n2188 99.5127
R16929 vdd.n1150 vdd.n1149 99.5127
R16930 vdd.n1154 vdd.n1153 99.5127
R16931 vdd.n1158 vdd.n1157 99.5127
R16932 vdd.n1162 vdd.n1161 99.5127
R16933 vdd.n1166 vdd.n1165 99.5127
R16934 vdd.n1170 vdd.n1169 99.5127
R16935 vdd.n1174 vdd.n1173 99.5127
R16936 vdd.n1179 vdd.n1178 99.5127
R16937 vdd.n2224 vdd.n966 99.5127
R16938 vdd.n2224 vdd.n956 99.5127
R16939 vdd.n2232 vdd.n956 99.5127
R16940 vdd.n2232 vdd.n954 99.5127
R16941 vdd.n2236 vdd.n954 99.5127
R16942 vdd.n2236 vdd.n943 99.5127
R16943 vdd.n2244 vdd.n943 99.5127
R16944 vdd.n2244 vdd.n941 99.5127
R16945 vdd.n2248 vdd.n941 99.5127
R16946 vdd.n2248 vdd.n931 99.5127
R16947 vdd.n2256 vdd.n931 99.5127
R16948 vdd.n2256 vdd.n929 99.5127
R16949 vdd.n2260 vdd.n929 99.5127
R16950 vdd.n2260 vdd.n920 99.5127
R16951 vdd.n2268 vdd.n920 99.5127
R16952 vdd.n2268 vdd.n918 99.5127
R16953 vdd.n2272 vdd.n918 99.5127
R16954 vdd.n2272 vdd.n907 99.5127
R16955 vdd.n2280 vdd.n907 99.5127
R16956 vdd.n2280 vdd.n905 99.5127
R16957 vdd.n2284 vdd.n905 99.5127
R16958 vdd.n2284 vdd.n895 99.5127
R16959 vdd.n2293 vdd.n895 99.5127
R16960 vdd.n2293 vdd.n893 99.5127
R16961 vdd.n2297 vdd.n893 99.5127
R16962 vdd.n2297 vdd.n883 99.5127
R16963 vdd.n2305 vdd.n883 99.5127
R16964 vdd.n2305 vdd.n881 99.5127
R16965 vdd.n2309 vdd.n881 99.5127
R16966 vdd.n2309 vdd.n871 99.5127
R16967 vdd.n2317 vdd.n871 99.5127
R16968 vdd.n2317 vdd.n869 99.5127
R16969 vdd.n2321 vdd.n869 99.5127
R16970 vdd.n2321 vdd.n861 99.5127
R16971 vdd.n2329 vdd.n861 99.5127
R16972 vdd.n2329 vdd.n859 99.5127
R16973 vdd.n2333 vdd.n859 99.5127
R16974 vdd.n2333 vdd.n848 99.5127
R16975 vdd.n2343 vdd.n848 99.5127
R16976 vdd.n2343 vdd.n845 99.5127
R16977 vdd.n2348 vdd.n845 99.5127
R16978 vdd.n2348 vdd.n846 99.5127
R16979 vdd.n846 vdd.n826 99.5127
R16980 vdd.n2958 vdd.n2957 99.5127
R16981 vdd.n2955 vdd.n2921 99.5127
R16982 vdd.n2951 vdd.n2950 99.5127
R16983 vdd.n2948 vdd.n2924 99.5127
R16984 vdd.n2944 vdd.n2943 99.5127
R16985 vdd.n2941 vdd.n2927 99.5127
R16986 vdd.n2937 vdd.n2936 99.5127
R16987 vdd.n2934 vdd.n2931 99.5127
R16988 vdd.n3075 vdd.n612 99.5127
R16989 vdd.n3073 vdd.n3072 99.5127
R16990 vdd.n3070 vdd.n615 99.5127
R16991 vdd.n3066 vdd.n3065 99.5127
R16992 vdd.n3063 vdd.n618 99.5127
R16993 vdd.n3059 vdd.n3058 99.5127
R16994 vdd.n3056 vdd.n621 99.5127
R16995 vdd.n3052 vdd.n3051 99.5127
R16996 vdd.n3049 vdd.n624 99.5127
R16997 vdd.n2607 vdd.n787 99.5127
R16998 vdd.n2727 vdd.n787 99.5127
R16999 vdd.n2727 vdd.n781 99.5127
R17000 vdd.n2723 vdd.n781 99.5127
R17001 vdd.n2723 vdd.n776 99.5127
R17002 vdd.n2720 vdd.n776 99.5127
R17003 vdd.n2720 vdd.n770 99.5127
R17004 vdd.n2717 vdd.n770 99.5127
R17005 vdd.n2717 vdd.n764 99.5127
R17006 vdd.n2709 vdd.n764 99.5127
R17007 vdd.n2709 vdd.n758 99.5127
R17008 vdd.n2705 vdd.n758 99.5127
R17009 vdd.n2705 vdd.n752 99.5127
R17010 vdd.n2702 vdd.n752 99.5127
R17011 vdd.n2702 vdd.n747 99.5127
R17012 vdd.n2699 vdd.n747 99.5127
R17013 vdd.n2699 vdd.n742 99.5127
R17014 vdd.n2696 vdd.n742 99.5127
R17015 vdd.n2696 vdd.n735 99.5127
R17016 vdd.n2693 vdd.n735 99.5127
R17017 vdd.n2693 vdd.n728 99.5127
R17018 vdd.n2690 vdd.n728 99.5127
R17019 vdd.n2690 vdd.n722 99.5127
R17020 vdd.n2687 vdd.n722 99.5127
R17021 vdd.n2687 vdd.n717 99.5127
R17022 vdd.n2684 vdd.n717 99.5127
R17023 vdd.n2684 vdd.n711 99.5127
R17024 vdd.n2681 vdd.n711 99.5127
R17025 vdd.n2681 vdd.n704 99.5127
R17026 vdd.n2678 vdd.n704 99.5127
R17027 vdd.n2678 vdd.n697 99.5127
R17028 vdd.n2675 vdd.n697 99.5127
R17029 vdd.n2675 vdd.n691 99.5127
R17030 vdd.n2672 vdd.n691 99.5127
R17031 vdd.n2672 vdd.n686 99.5127
R17032 vdd.n2669 vdd.n686 99.5127
R17033 vdd.n2669 vdd.n681 99.5127
R17034 vdd.n2666 vdd.n681 99.5127
R17035 vdd.n2666 vdd.n673 99.5127
R17036 vdd.n2663 vdd.n673 99.5127
R17037 vdd.n2663 vdd.n666 99.5127
R17038 vdd.n666 vdd.n630 99.5127
R17039 vdd.n3044 vdd.n630 99.5127
R17040 vdd.n2542 vdd.n2541 99.5127
R17041 vdd.n2546 vdd.n2545 99.5127
R17042 vdd.n2550 vdd.n2549 99.5127
R17043 vdd.n2554 vdd.n2553 99.5127
R17044 vdd.n2558 vdd.n2557 99.5127
R17045 vdd.n2562 vdd.n2561 99.5127
R17046 vdd.n2566 vdd.n2565 99.5127
R17047 vdd.n2570 vdd.n2569 99.5127
R17048 vdd.n2574 vdd.n2573 99.5127
R17049 vdd.n2578 vdd.n2577 99.5127
R17050 vdd.n2582 vdd.n2581 99.5127
R17051 vdd.n2586 vdd.n2585 99.5127
R17052 vdd.n2590 vdd.n2589 99.5127
R17053 vdd.n2594 vdd.n2593 99.5127
R17054 vdd.n2598 vdd.n2597 99.5127
R17055 vdd.n2602 vdd.n2601 99.5127
R17056 vdd.n2604 vdd.n2530 99.5127
R17057 vdd.n2808 vdd.n784 99.5127
R17058 vdd.n2808 vdd.n782 99.5127
R17059 vdd.n2812 vdd.n782 99.5127
R17060 vdd.n2812 vdd.n773 99.5127
R17061 vdd.n2820 vdd.n773 99.5127
R17062 vdd.n2820 vdd.n771 99.5127
R17063 vdd.n2824 vdd.n771 99.5127
R17064 vdd.n2824 vdd.n762 99.5127
R17065 vdd.n2832 vdd.n762 99.5127
R17066 vdd.n2832 vdd.n760 99.5127
R17067 vdd.n2836 vdd.n760 99.5127
R17068 vdd.n2836 vdd.n750 99.5127
R17069 vdd.n2844 vdd.n750 99.5127
R17070 vdd.n2844 vdd.n748 99.5127
R17071 vdd.n2848 vdd.n748 99.5127
R17072 vdd.n2848 vdd.n739 99.5127
R17073 vdd.n2856 vdd.n739 99.5127
R17074 vdd.n2856 vdd.n737 99.5127
R17075 vdd.n2861 vdd.n737 99.5127
R17076 vdd.n2861 vdd.n726 99.5127
R17077 vdd.n2869 vdd.n726 99.5127
R17078 vdd.n2869 vdd.n723 99.5127
R17079 vdd.n2873 vdd.n723 99.5127
R17080 vdd.n2873 vdd.n714 99.5127
R17081 vdd.n2881 vdd.n714 99.5127
R17082 vdd.n2881 vdd.n712 99.5127
R17083 vdd.n2885 vdd.n712 99.5127
R17084 vdd.n2885 vdd.n701 99.5127
R17085 vdd.n2893 vdd.n701 99.5127
R17086 vdd.n2893 vdd.n699 99.5127
R17087 vdd.n2897 vdd.n699 99.5127
R17088 vdd.n2897 vdd.n689 99.5127
R17089 vdd.n2905 vdd.n689 99.5127
R17090 vdd.n2905 vdd.n687 99.5127
R17091 vdd.n2909 vdd.n687 99.5127
R17092 vdd.n2909 vdd.n678 99.5127
R17093 vdd.n2917 vdd.n678 99.5127
R17094 vdd.n2917 vdd.n675 99.5127
R17095 vdd.n2966 vdd.n675 99.5127
R17096 vdd.n2966 vdd.n676 99.5127
R17097 vdd.n676 vdd.n667 99.5127
R17098 vdd.n2961 vdd.n667 99.5127
R17099 vdd.n2961 vdd.n633 99.5127
R17100 vdd.n2419 vdd.n2418 99.5127
R17101 vdd.n2415 vdd.n2414 99.5127
R17102 vdd.n2411 vdd.n2410 99.5127
R17103 vdd.n2407 vdd.n2406 99.5127
R17104 vdd.n2403 vdd.n2402 99.5127
R17105 vdd.n2399 vdd.n2398 99.5127
R17106 vdd.n2395 vdd.n2394 99.5127
R17107 vdd.n2391 vdd.n2390 99.5127
R17108 vdd.n2387 vdd.n2386 99.5127
R17109 vdd.n2383 vdd.n2382 99.5127
R17110 vdd.n2379 vdd.n2378 99.5127
R17111 vdd.n2375 vdd.n2374 99.5127
R17112 vdd.n2371 vdd.n2370 99.5127
R17113 vdd.n2367 vdd.n2366 99.5127
R17114 vdd.n2363 vdd.n2362 99.5127
R17115 vdd.n2359 vdd.n2358 99.5127
R17116 vdd.n2355 vdd.n808 99.5127
R17117 vdd.n1308 vdd.n964 99.5127
R17118 vdd.n1305 vdd.n964 99.5127
R17119 vdd.n1305 vdd.n958 99.5127
R17120 vdd.n1302 vdd.n958 99.5127
R17121 vdd.n1302 vdd.n953 99.5127
R17122 vdd.n1299 vdd.n953 99.5127
R17123 vdd.n1299 vdd.n946 99.5127
R17124 vdd.n1296 vdd.n946 99.5127
R17125 vdd.n1296 vdd.n939 99.5127
R17126 vdd.n1293 vdd.n939 99.5127
R17127 vdd.n1293 vdd.n933 99.5127
R17128 vdd.n1290 vdd.n933 99.5127
R17129 vdd.n1290 vdd.n928 99.5127
R17130 vdd.n1287 vdd.n928 99.5127
R17131 vdd.n1287 vdd.n923 99.5127
R17132 vdd.n1284 vdd.n923 99.5127
R17133 vdd.n1284 vdd.n917 99.5127
R17134 vdd.n1281 vdd.n917 99.5127
R17135 vdd.n1281 vdd.n910 99.5127
R17136 vdd.n1278 vdd.n910 99.5127
R17137 vdd.n1278 vdd.n903 99.5127
R17138 vdd.n1275 vdd.n903 99.5127
R17139 vdd.n1275 vdd.n897 99.5127
R17140 vdd.n1272 vdd.n897 99.5127
R17141 vdd.n1272 vdd.n892 99.5127
R17142 vdd.n1269 vdd.n892 99.5127
R17143 vdd.n1269 vdd.n886 99.5127
R17144 vdd.n1266 vdd.n886 99.5127
R17145 vdd.n1266 vdd.n879 99.5127
R17146 vdd.n1237 vdd.n879 99.5127
R17147 vdd.n1237 vdd.n873 99.5127
R17148 vdd.n1240 vdd.n873 99.5127
R17149 vdd.n1240 vdd.n868 99.5127
R17150 vdd.n1252 vdd.n868 99.5127
R17151 vdd.n1252 vdd.n863 99.5127
R17152 vdd.n1248 vdd.n863 99.5127
R17153 vdd.n1248 vdd.n858 99.5127
R17154 vdd.n1245 vdd.n858 99.5127
R17155 vdd.n1245 vdd.n851 99.5127
R17156 vdd.n851 vdd.n842 99.5127
R17157 vdd.n2350 vdd.n842 99.5127
R17158 vdd.n2351 vdd.n2350 99.5127
R17159 vdd.n2351 vdd.n834 99.5127
R17160 vdd.n1112 vdd.n1111 99.5127
R17161 vdd.n1116 vdd.n1115 99.5127
R17162 vdd.n1120 vdd.n1119 99.5127
R17163 vdd.n1124 vdd.n1123 99.5127
R17164 vdd.n1128 vdd.n1127 99.5127
R17165 vdd.n1132 vdd.n1131 99.5127
R17166 vdd.n1136 vdd.n1135 99.5127
R17167 vdd.n1140 vdd.n1139 99.5127
R17168 vdd.n1341 vdd.n1142 99.5127
R17169 vdd.n1339 vdd.n1338 99.5127
R17170 vdd.n1335 vdd.n1334 99.5127
R17171 vdd.n1331 vdd.n1330 99.5127
R17172 vdd.n1327 vdd.n1326 99.5127
R17173 vdd.n1323 vdd.n1322 99.5127
R17174 vdd.n1319 vdd.n1318 99.5127
R17175 vdd.n1315 vdd.n1314 99.5127
R17176 vdd.n1311 vdd.n1003 99.5127
R17177 vdd.n2226 vdd.n961 99.5127
R17178 vdd.n2226 vdd.n959 99.5127
R17179 vdd.n2230 vdd.n959 99.5127
R17180 vdd.n2230 vdd.n950 99.5127
R17181 vdd.n2238 vdd.n950 99.5127
R17182 vdd.n2238 vdd.n948 99.5127
R17183 vdd.n2242 vdd.n948 99.5127
R17184 vdd.n2242 vdd.n937 99.5127
R17185 vdd.n2250 vdd.n937 99.5127
R17186 vdd.n2250 vdd.n935 99.5127
R17187 vdd.n2254 vdd.n935 99.5127
R17188 vdd.n2254 vdd.n926 99.5127
R17189 vdd.n2262 vdd.n926 99.5127
R17190 vdd.n2262 vdd.n924 99.5127
R17191 vdd.n2266 vdd.n924 99.5127
R17192 vdd.n2266 vdd.n914 99.5127
R17193 vdd.n2274 vdd.n914 99.5127
R17194 vdd.n2274 vdd.n912 99.5127
R17195 vdd.n2278 vdd.n912 99.5127
R17196 vdd.n2278 vdd.n901 99.5127
R17197 vdd.n2286 vdd.n901 99.5127
R17198 vdd.n2286 vdd.n898 99.5127
R17199 vdd.n2291 vdd.n898 99.5127
R17200 vdd.n2291 vdd.n889 99.5127
R17201 vdd.n2299 vdd.n889 99.5127
R17202 vdd.n2299 vdd.n887 99.5127
R17203 vdd.n2303 vdd.n887 99.5127
R17204 vdd.n2303 vdd.n877 99.5127
R17205 vdd.n2311 vdd.n877 99.5127
R17206 vdd.n2311 vdd.n875 99.5127
R17207 vdd.n2315 vdd.n875 99.5127
R17208 vdd.n2315 vdd.n866 99.5127
R17209 vdd.n2323 vdd.n866 99.5127
R17210 vdd.n2323 vdd.n864 99.5127
R17211 vdd.n2327 vdd.n864 99.5127
R17212 vdd.n2327 vdd.n855 99.5127
R17213 vdd.n2335 vdd.n855 99.5127
R17214 vdd.n2335 vdd.n852 99.5127
R17215 vdd.n2341 vdd.n852 99.5127
R17216 vdd.n2341 vdd.n853 99.5127
R17217 vdd.n853 vdd.n844 99.5127
R17218 vdd.n844 vdd.n835 99.5127
R17219 vdd.n2423 vdd.n835 99.5127
R17220 vdd.n9 vdd.n7 98.9633
R17221 vdd.n2 vdd.n0 98.9633
R17222 vdd.n9 vdd.n8 98.6055
R17223 vdd.n11 vdd.n10 98.6055
R17224 vdd.n13 vdd.n12 98.6055
R17225 vdd.n6 vdd.n5 98.6055
R17226 vdd.n4 vdd.n3 98.6055
R17227 vdd.n2 vdd.n1 98.6055
R17228 vdd.t156 vdd.n279 85.8723
R17229 vdd.t238 vdd.n228 85.8723
R17230 vdd.t145 vdd.n185 85.8723
R17231 vdd.t114 vdd.n134 85.8723
R17232 vdd.t118 vdd.n92 85.8723
R17233 vdd.t5 vdd.n41 85.8723
R17234 vdd.t234 vdd.n1929 85.8723
R17235 vdd.t147 vdd.n1980 85.8723
R17236 vdd.t133 vdd.n1835 85.8723
R17237 vdd.t116 vdd.n1886 85.8723
R17238 vdd.t3 vdd.n1742 85.8723
R17239 vdd.t123 vdd.n1793 85.8723
R17240 vdd.n725 vdd.n724 78.546
R17241 vdd.n2289 vdd.n899 78.546
R17242 vdd.n266 vdd.n265 75.1835
R17243 vdd.n264 vdd.n263 75.1835
R17244 vdd.n262 vdd.n261 75.1835
R17245 vdd.n260 vdd.n259 75.1835
R17246 vdd.n258 vdd.n257 75.1835
R17247 vdd.n172 vdd.n171 75.1835
R17248 vdd.n170 vdd.n169 75.1835
R17249 vdd.n168 vdd.n167 75.1835
R17250 vdd.n166 vdd.n165 75.1835
R17251 vdd.n164 vdd.n163 75.1835
R17252 vdd.n79 vdd.n78 75.1835
R17253 vdd.n77 vdd.n76 75.1835
R17254 vdd.n75 vdd.n74 75.1835
R17255 vdd.n73 vdd.n72 75.1835
R17256 vdd.n71 vdd.n70 75.1835
R17257 vdd.n1959 vdd.n1958 75.1835
R17258 vdd.n1961 vdd.n1960 75.1835
R17259 vdd.n1963 vdd.n1962 75.1835
R17260 vdd.n1965 vdd.n1964 75.1835
R17261 vdd.n1967 vdd.n1966 75.1835
R17262 vdd.n1865 vdd.n1864 75.1835
R17263 vdd.n1867 vdd.n1866 75.1835
R17264 vdd.n1869 vdd.n1868 75.1835
R17265 vdd.n1871 vdd.n1870 75.1835
R17266 vdd.n1873 vdd.n1872 75.1835
R17267 vdd.n1772 vdd.n1771 75.1835
R17268 vdd.n1774 vdd.n1773 75.1835
R17269 vdd.n1776 vdd.n1775 75.1835
R17270 vdd.n1778 vdd.n1777 75.1835
R17271 vdd.n1780 vdd.n1779 75.1835
R17272 vdd.n2800 vdd.n2513 72.8958
R17273 vdd.n2800 vdd.n2514 72.8958
R17274 vdd.n2800 vdd.n2515 72.8958
R17275 vdd.n2800 vdd.n2516 72.8958
R17276 vdd.n2800 vdd.n2517 72.8958
R17277 vdd.n2800 vdd.n2518 72.8958
R17278 vdd.n2800 vdd.n2519 72.8958
R17279 vdd.n2800 vdd.n2520 72.8958
R17280 vdd.n2800 vdd.n2521 72.8958
R17281 vdd.n2800 vdd.n2522 72.8958
R17282 vdd.n2800 vdd.n2523 72.8958
R17283 vdd.n2800 vdd.n2524 72.8958
R17284 vdd.n2800 vdd.n2525 72.8958
R17285 vdd.n2800 vdd.n2526 72.8958
R17286 vdd.n2800 vdd.n2527 72.8958
R17287 vdd.n2800 vdd.n2528 72.8958
R17288 vdd.n2800 vdd.n2529 72.8958
R17289 vdd.n629 vdd.n613 72.8958
R17290 vdd.n3050 vdd.n613 72.8958
R17291 vdd.n623 vdd.n613 72.8958
R17292 vdd.n3057 vdd.n613 72.8958
R17293 vdd.n620 vdd.n613 72.8958
R17294 vdd.n3064 vdd.n613 72.8958
R17295 vdd.n617 vdd.n613 72.8958
R17296 vdd.n3071 vdd.n613 72.8958
R17297 vdd.n3074 vdd.n613 72.8958
R17298 vdd.n2930 vdd.n613 72.8958
R17299 vdd.n2935 vdd.n613 72.8958
R17300 vdd.n2929 vdd.n613 72.8958
R17301 vdd.n2942 vdd.n613 72.8958
R17302 vdd.n2926 vdd.n613 72.8958
R17303 vdd.n2949 vdd.n613 72.8958
R17304 vdd.n2923 vdd.n613 72.8958
R17305 vdd.n2956 vdd.n613 72.8958
R17306 vdd.n2219 vdd.n2218 72.8958
R17307 vdd.n2218 vdd.n970 72.8958
R17308 vdd.n2218 vdd.n971 72.8958
R17309 vdd.n2218 vdd.n972 72.8958
R17310 vdd.n2218 vdd.n973 72.8958
R17311 vdd.n2218 vdd.n974 72.8958
R17312 vdd.n2218 vdd.n975 72.8958
R17313 vdd.n2218 vdd.n976 72.8958
R17314 vdd.n2218 vdd.n977 72.8958
R17315 vdd.n2218 vdd.n978 72.8958
R17316 vdd.n2218 vdd.n979 72.8958
R17317 vdd.n2218 vdd.n980 72.8958
R17318 vdd.n2218 vdd.n981 72.8958
R17319 vdd.n2218 vdd.n982 72.8958
R17320 vdd.n2218 vdd.n983 72.8958
R17321 vdd.n2218 vdd.n984 72.8958
R17322 vdd.n2218 vdd.n985 72.8958
R17323 vdd.n2496 vdd.n809 72.8958
R17324 vdd.n2496 vdd.n810 72.8958
R17325 vdd.n2496 vdd.n811 72.8958
R17326 vdd.n2496 vdd.n812 72.8958
R17327 vdd.n2496 vdd.n813 72.8958
R17328 vdd.n2496 vdd.n814 72.8958
R17329 vdd.n2496 vdd.n815 72.8958
R17330 vdd.n2496 vdd.n816 72.8958
R17331 vdd.n2496 vdd.n817 72.8958
R17332 vdd.n2496 vdd.n818 72.8958
R17333 vdd.n2496 vdd.n819 72.8958
R17334 vdd.n2496 vdd.n820 72.8958
R17335 vdd.n2496 vdd.n821 72.8958
R17336 vdd.n2496 vdd.n822 72.8958
R17337 vdd.n2496 vdd.n823 72.8958
R17338 vdd.n2496 vdd.n824 72.8958
R17339 vdd.n2496 vdd.n825 72.8958
R17340 vdd.n2801 vdd.n2800 72.8958
R17341 vdd.n2800 vdd.n2497 72.8958
R17342 vdd.n2800 vdd.n2498 72.8958
R17343 vdd.n2800 vdd.n2499 72.8958
R17344 vdd.n2800 vdd.n2500 72.8958
R17345 vdd.n2800 vdd.n2501 72.8958
R17346 vdd.n2800 vdd.n2502 72.8958
R17347 vdd.n2800 vdd.n2503 72.8958
R17348 vdd.n2800 vdd.n2504 72.8958
R17349 vdd.n2800 vdd.n2505 72.8958
R17350 vdd.n2800 vdd.n2506 72.8958
R17351 vdd.n2800 vdd.n2507 72.8958
R17352 vdd.n2800 vdd.n2508 72.8958
R17353 vdd.n2800 vdd.n2509 72.8958
R17354 vdd.n2800 vdd.n2510 72.8958
R17355 vdd.n2800 vdd.n2511 72.8958
R17356 vdd.n2800 vdd.n2512 72.8958
R17357 vdd.n2978 vdd.n613 72.8958
R17358 vdd.n2984 vdd.n613 72.8958
R17359 vdd.n659 vdd.n613 72.8958
R17360 vdd.n2991 vdd.n613 72.8958
R17361 vdd.n656 vdd.n613 72.8958
R17362 vdd.n2998 vdd.n613 72.8958
R17363 vdd.n653 vdd.n613 72.8958
R17364 vdd.n3005 vdd.n613 72.8958
R17365 vdd.n650 vdd.n613 72.8958
R17366 vdd.n3013 vdd.n613 72.8958
R17367 vdd.n647 vdd.n613 72.8958
R17368 vdd.n3020 vdd.n613 72.8958
R17369 vdd.n644 vdd.n613 72.8958
R17370 vdd.n3027 vdd.n613 72.8958
R17371 vdd.n641 vdd.n613 72.8958
R17372 vdd.n3034 vdd.n613 72.8958
R17373 vdd.n3037 vdd.n613 72.8958
R17374 vdd.n2496 vdd.n807 72.8958
R17375 vdd.n2496 vdd.n806 72.8958
R17376 vdd.n2496 vdd.n805 72.8958
R17377 vdd.n2496 vdd.n804 72.8958
R17378 vdd.n2496 vdd.n803 72.8958
R17379 vdd.n2496 vdd.n802 72.8958
R17380 vdd.n2496 vdd.n801 72.8958
R17381 vdd.n2496 vdd.n800 72.8958
R17382 vdd.n2496 vdd.n799 72.8958
R17383 vdd.n2496 vdd.n798 72.8958
R17384 vdd.n2496 vdd.n797 72.8958
R17385 vdd.n2496 vdd.n796 72.8958
R17386 vdd.n2496 vdd.n795 72.8958
R17387 vdd.n2496 vdd.n794 72.8958
R17388 vdd.n2496 vdd.n793 72.8958
R17389 vdd.n2496 vdd.n792 72.8958
R17390 vdd.n2496 vdd.n791 72.8958
R17391 vdd.n2218 vdd.n986 72.8958
R17392 vdd.n2218 vdd.n987 72.8958
R17393 vdd.n2218 vdd.n988 72.8958
R17394 vdd.n2218 vdd.n989 72.8958
R17395 vdd.n2218 vdd.n990 72.8958
R17396 vdd.n2218 vdd.n991 72.8958
R17397 vdd.n2218 vdd.n992 72.8958
R17398 vdd.n2218 vdd.n993 72.8958
R17399 vdd.n2218 vdd.n994 72.8958
R17400 vdd.n2218 vdd.n995 72.8958
R17401 vdd.n2218 vdd.n996 72.8958
R17402 vdd.n2218 vdd.n997 72.8958
R17403 vdd.n2218 vdd.n998 72.8958
R17404 vdd.n2218 vdd.n999 72.8958
R17405 vdd.n2218 vdd.n1000 72.8958
R17406 vdd.n2218 vdd.n1001 72.8958
R17407 vdd.n2218 vdd.n1002 72.8958
R17408 vdd.n1441 vdd.n1437 66.2847
R17409 vdd.n1447 vdd.n1437 66.2847
R17410 vdd.n1450 vdd.n1437 66.2847
R17411 vdd.n1455 vdd.n1437 66.2847
R17412 vdd.n1458 vdd.n1437 66.2847
R17413 vdd.n1463 vdd.n1437 66.2847
R17414 vdd.n1466 vdd.n1437 66.2847
R17415 vdd.n1471 vdd.n1437 66.2847
R17416 vdd.n1474 vdd.n1437 66.2847
R17417 vdd.n1481 vdd.n1437 66.2847
R17418 vdd.n1484 vdd.n1437 66.2847
R17419 vdd.n1489 vdd.n1437 66.2847
R17420 vdd.n1492 vdd.n1437 66.2847
R17421 vdd.n1497 vdd.n1437 66.2847
R17422 vdd.n1500 vdd.n1437 66.2847
R17423 vdd.n1505 vdd.n1437 66.2847
R17424 vdd.n1508 vdd.n1437 66.2847
R17425 vdd.n1513 vdd.n1437 66.2847
R17426 vdd.n1516 vdd.n1437 66.2847
R17427 vdd.n1521 vdd.n1437 66.2847
R17428 vdd.n1600 vdd.n1437 66.2847
R17429 vdd.n1524 vdd.n1437 66.2847
R17430 vdd.n1530 vdd.n1437 66.2847
R17431 vdd.n1535 vdd.n1437 66.2847
R17432 vdd.n1538 vdd.n1437 66.2847
R17433 vdd.n1543 vdd.n1437 66.2847
R17434 vdd.n1546 vdd.n1437 66.2847
R17435 vdd.n1551 vdd.n1437 66.2847
R17436 vdd.n1554 vdd.n1437 66.2847
R17437 vdd.n1559 vdd.n1437 66.2847
R17438 vdd.n1562 vdd.n1437 66.2847
R17439 vdd.n1354 vdd.n969 66.2847
R17440 vdd.n1351 vdd.n969 66.2847
R17441 vdd.n1347 vdd.n969 66.2847
R17442 vdd.n2084 vdd.n969 66.2847
R17443 vdd.n1103 vdd.n969 66.2847
R17444 vdd.n2091 vdd.n969 66.2847
R17445 vdd.n1096 vdd.n969 66.2847
R17446 vdd.n2098 vdd.n969 66.2847
R17447 vdd.n1089 vdd.n969 66.2847
R17448 vdd.n2105 vdd.n969 66.2847
R17449 vdd.n1083 vdd.n969 66.2847
R17450 vdd.n1078 vdd.n969 66.2847
R17451 vdd.n2116 vdd.n969 66.2847
R17452 vdd.n1070 vdd.n969 66.2847
R17453 vdd.n2123 vdd.n969 66.2847
R17454 vdd.n1063 vdd.n969 66.2847
R17455 vdd.n2130 vdd.n969 66.2847
R17456 vdd.n1056 vdd.n969 66.2847
R17457 vdd.n2137 vdd.n969 66.2847
R17458 vdd.n1049 vdd.n969 66.2847
R17459 vdd.n2144 vdd.n969 66.2847
R17460 vdd.n1043 vdd.n969 66.2847
R17461 vdd.n1038 vdd.n969 66.2847
R17462 vdd.n2155 vdd.n969 66.2847
R17463 vdd.n1030 vdd.n969 66.2847
R17464 vdd.n2162 vdd.n969 66.2847
R17465 vdd.n1023 vdd.n969 66.2847
R17466 vdd.n2169 vdd.n969 66.2847
R17467 vdd.n1016 vdd.n969 66.2847
R17468 vdd.n2176 vdd.n969 66.2847
R17469 vdd.n2181 vdd.n969 66.2847
R17470 vdd.n1012 vdd.n969 66.2847
R17471 vdd.n3204 vdd.n516 66.2847
R17472 vdd.n520 vdd.n516 66.2847
R17473 vdd.n523 vdd.n516 66.2847
R17474 vdd.n3193 vdd.n516 66.2847
R17475 vdd.n3187 vdd.n516 66.2847
R17476 vdd.n3185 vdd.n516 66.2847
R17477 vdd.n3179 vdd.n516 66.2847
R17478 vdd.n3177 vdd.n516 66.2847
R17479 vdd.n3171 vdd.n516 66.2847
R17480 vdd.n3169 vdd.n516 66.2847
R17481 vdd.n3163 vdd.n516 66.2847
R17482 vdd.n3161 vdd.n516 66.2847
R17483 vdd.n3155 vdd.n516 66.2847
R17484 vdd.n3153 vdd.n516 66.2847
R17485 vdd.n3147 vdd.n516 66.2847
R17486 vdd.n3145 vdd.n516 66.2847
R17487 vdd.n3139 vdd.n516 66.2847
R17488 vdd.n3137 vdd.n516 66.2847
R17489 vdd.n3131 vdd.n516 66.2847
R17490 vdd.n3129 vdd.n516 66.2847
R17491 vdd.n584 vdd.n516 66.2847
R17492 vdd.n3120 vdd.n516 66.2847
R17493 vdd.n586 vdd.n516 66.2847
R17494 vdd.n3113 vdd.n516 66.2847
R17495 vdd.n3107 vdd.n516 66.2847
R17496 vdd.n3105 vdd.n516 66.2847
R17497 vdd.n3099 vdd.n516 66.2847
R17498 vdd.n3097 vdd.n516 66.2847
R17499 vdd.n3091 vdd.n516 66.2847
R17500 vdd.n607 vdd.n516 66.2847
R17501 vdd.n609 vdd.n516 66.2847
R17502 vdd.n3290 vdd.n351 66.2847
R17503 vdd.n3299 vdd.n351 66.2847
R17504 vdd.n461 vdd.n351 66.2847
R17505 vdd.n3306 vdd.n351 66.2847
R17506 vdd.n454 vdd.n351 66.2847
R17507 vdd.n3313 vdd.n351 66.2847
R17508 vdd.n447 vdd.n351 66.2847
R17509 vdd.n3320 vdd.n351 66.2847
R17510 vdd.n440 vdd.n351 66.2847
R17511 vdd.n3327 vdd.n351 66.2847
R17512 vdd.n434 vdd.n351 66.2847
R17513 vdd.n429 vdd.n351 66.2847
R17514 vdd.n3338 vdd.n351 66.2847
R17515 vdd.n421 vdd.n351 66.2847
R17516 vdd.n3345 vdd.n351 66.2847
R17517 vdd.n414 vdd.n351 66.2847
R17518 vdd.n3352 vdd.n351 66.2847
R17519 vdd.n407 vdd.n351 66.2847
R17520 vdd.n3359 vdd.n351 66.2847
R17521 vdd.n400 vdd.n351 66.2847
R17522 vdd.n3366 vdd.n351 66.2847
R17523 vdd.n394 vdd.n351 66.2847
R17524 vdd.n389 vdd.n351 66.2847
R17525 vdd.n3377 vdd.n351 66.2847
R17526 vdd.n381 vdd.n351 66.2847
R17527 vdd.n3384 vdd.n351 66.2847
R17528 vdd.n374 vdd.n351 66.2847
R17529 vdd.n3391 vdd.n351 66.2847
R17530 vdd.n367 vdd.n351 66.2847
R17531 vdd.n3398 vdd.n351 66.2847
R17532 vdd.n3401 vdd.n351 66.2847
R17533 vdd.n355 vdd.n351 66.2847
R17534 vdd.n356 vdd.n355 52.4337
R17535 vdd.n3401 vdd.n3400 52.4337
R17536 vdd.n3398 vdd.n3397 52.4337
R17537 vdd.n3393 vdd.n367 52.4337
R17538 vdd.n3391 vdd.n3390 52.4337
R17539 vdd.n3386 vdd.n374 52.4337
R17540 vdd.n3384 vdd.n3383 52.4337
R17541 vdd.n3379 vdd.n381 52.4337
R17542 vdd.n3377 vdd.n3376 52.4337
R17543 vdd.n390 vdd.n389 52.4337
R17544 vdd.n3368 vdd.n394 52.4337
R17545 vdd.n3366 vdd.n3365 52.4337
R17546 vdd.n3361 vdd.n400 52.4337
R17547 vdd.n3359 vdd.n3358 52.4337
R17548 vdd.n3354 vdd.n407 52.4337
R17549 vdd.n3352 vdd.n3351 52.4337
R17550 vdd.n3347 vdd.n414 52.4337
R17551 vdd.n3345 vdd.n3344 52.4337
R17552 vdd.n3340 vdd.n421 52.4337
R17553 vdd.n3338 vdd.n3337 52.4337
R17554 vdd.n430 vdd.n429 52.4337
R17555 vdd.n3329 vdd.n434 52.4337
R17556 vdd.n3327 vdd.n3326 52.4337
R17557 vdd.n3322 vdd.n440 52.4337
R17558 vdd.n3320 vdd.n3319 52.4337
R17559 vdd.n3315 vdd.n447 52.4337
R17560 vdd.n3313 vdd.n3312 52.4337
R17561 vdd.n3308 vdd.n454 52.4337
R17562 vdd.n3306 vdd.n3305 52.4337
R17563 vdd.n3301 vdd.n461 52.4337
R17564 vdd.n3299 vdd.n3298 52.4337
R17565 vdd.n3291 vdd.n3290 52.4337
R17566 vdd.n3204 vdd.n517 52.4337
R17567 vdd.n3202 vdd.n520 52.4337
R17568 vdd.n3198 vdd.n523 52.4337
R17569 vdd.n3194 vdd.n3193 52.4337
R17570 vdd.n3187 vdd.n526 52.4337
R17571 vdd.n3186 vdd.n3185 52.4337
R17572 vdd.n3179 vdd.n532 52.4337
R17573 vdd.n3178 vdd.n3177 52.4337
R17574 vdd.n3171 vdd.n538 52.4337
R17575 vdd.n3170 vdd.n3169 52.4337
R17576 vdd.n3163 vdd.n546 52.4337
R17577 vdd.n3162 vdd.n3161 52.4337
R17578 vdd.n3155 vdd.n552 52.4337
R17579 vdd.n3154 vdd.n3153 52.4337
R17580 vdd.n3147 vdd.n558 52.4337
R17581 vdd.n3146 vdd.n3145 52.4337
R17582 vdd.n3139 vdd.n564 52.4337
R17583 vdd.n3138 vdd.n3137 52.4337
R17584 vdd.n3131 vdd.n570 52.4337
R17585 vdd.n3130 vdd.n3129 52.4337
R17586 vdd.n584 vdd.n576 52.4337
R17587 vdd.n3121 vdd.n3120 52.4337
R17588 vdd.n3118 vdd.n586 52.4337
R17589 vdd.n3114 vdd.n3113 52.4337
R17590 vdd.n3107 vdd.n590 52.4337
R17591 vdd.n3106 vdd.n3105 52.4337
R17592 vdd.n3099 vdd.n596 52.4337
R17593 vdd.n3098 vdd.n3097 52.4337
R17594 vdd.n3091 vdd.n602 52.4337
R17595 vdd.n3090 vdd.n607 52.4337
R17596 vdd.n3086 vdd.n609 52.4337
R17597 vdd.n2183 vdd.n1012 52.4337
R17598 vdd.n2181 vdd.n2180 52.4337
R17599 vdd.n2176 vdd.n2175 52.4337
R17600 vdd.n2171 vdd.n1016 52.4337
R17601 vdd.n2169 vdd.n2168 52.4337
R17602 vdd.n2164 vdd.n1023 52.4337
R17603 vdd.n2162 vdd.n2161 52.4337
R17604 vdd.n2157 vdd.n1030 52.4337
R17605 vdd.n2155 vdd.n2154 52.4337
R17606 vdd.n1039 vdd.n1038 52.4337
R17607 vdd.n2146 vdd.n1043 52.4337
R17608 vdd.n2144 vdd.n2143 52.4337
R17609 vdd.n2139 vdd.n1049 52.4337
R17610 vdd.n2137 vdd.n2136 52.4337
R17611 vdd.n2132 vdd.n1056 52.4337
R17612 vdd.n2130 vdd.n2129 52.4337
R17613 vdd.n2125 vdd.n1063 52.4337
R17614 vdd.n2123 vdd.n2122 52.4337
R17615 vdd.n2118 vdd.n1070 52.4337
R17616 vdd.n2116 vdd.n2115 52.4337
R17617 vdd.n1079 vdd.n1078 52.4337
R17618 vdd.n2107 vdd.n1083 52.4337
R17619 vdd.n2105 vdd.n2104 52.4337
R17620 vdd.n2100 vdd.n1089 52.4337
R17621 vdd.n2098 vdd.n2097 52.4337
R17622 vdd.n2093 vdd.n1096 52.4337
R17623 vdd.n2091 vdd.n2090 52.4337
R17624 vdd.n2086 vdd.n1103 52.4337
R17625 vdd.n2084 vdd.n2083 52.4337
R17626 vdd.n1348 vdd.n1347 52.4337
R17627 vdd.n1352 vdd.n1351 52.4337
R17628 vdd.n2072 vdd.n1354 52.4337
R17629 vdd.n1441 vdd.n1439 52.4337
R17630 vdd.n1447 vdd.n1446 52.4337
R17631 vdd.n1450 vdd.n1449 52.4337
R17632 vdd.n1455 vdd.n1454 52.4337
R17633 vdd.n1458 vdd.n1457 52.4337
R17634 vdd.n1463 vdd.n1462 52.4337
R17635 vdd.n1466 vdd.n1465 52.4337
R17636 vdd.n1471 vdd.n1470 52.4337
R17637 vdd.n1474 vdd.n1473 52.4337
R17638 vdd.n1481 vdd.n1480 52.4337
R17639 vdd.n1484 vdd.n1483 52.4337
R17640 vdd.n1489 vdd.n1488 52.4337
R17641 vdd.n1492 vdd.n1491 52.4337
R17642 vdd.n1497 vdd.n1496 52.4337
R17643 vdd.n1500 vdd.n1499 52.4337
R17644 vdd.n1505 vdd.n1504 52.4337
R17645 vdd.n1508 vdd.n1507 52.4337
R17646 vdd.n1513 vdd.n1512 52.4337
R17647 vdd.n1516 vdd.n1515 52.4337
R17648 vdd.n1521 vdd.n1520 52.4337
R17649 vdd.n1601 vdd.n1600 52.4337
R17650 vdd.n1598 vdd.n1524 52.4337
R17651 vdd.n1530 vdd.n1529 52.4337
R17652 vdd.n1535 vdd.n1532 52.4337
R17653 vdd.n1538 vdd.n1537 52.4337
R17654 vdd.n1543 vdd.n1540 52.4337
R17655 vdd.n1546 vdd.n1545 52.4337
R17656 vdd.n1551 vdd.n1548 52.4337
R17657 vdd.n1554 vdd.n1553 52.4337
R17658 vdd.n1559 vdd.n1556 52.4337
R17659 vdd.n1562 vdd.n1561 52.4337
R17660 vdd.n1442 vdd.n1441 52.4337
R17661 vdd.n1448 vdd.n1447 52.4337
R17662 vdd.n1451 vdd.n1450 52.4337
R17663 vdd.n1456 vdd.n1455 52.4337
R17664 vdd.n1459 vdd.n1458 52.4337
R17665 vdd.n1464 vdd.n1463 52.4337
R17666 vdd.n1467 vdd.n1466 52.4337
R17667 vdd.n1472 vdd.n1471 52.4337
R17668 vdd.n1475 vdd.n1474 52.4337
R17669 vdd.n1482 vdd.n1481 52.4337
R17670 vdd.n1485 vdd.n1484 52.4337
R17671 vdd.n1490 vdd.n1489 52.4337
R17672 vdd.n1493 vdd.n1492 52.4337
R17673 vdd.n1498 vdd.n1497 52.4337
R17674 vdd.n1501 vdd.n1500 52.4337
R17675 vdd.n1506 vdd.n1505 52.4337
R17676 vdd.n1509 vdd.n1508 52.4337
R17677 vdd.n1514 vdd.n1513 52.4337
R17678 vdd.n1517 vdd.n1516 52.4337
R17679 vdd.n1522 vdd.n1521 52.4337
R17680 vdd.n1600 vdd.n1599 52.4337
R17681 vdd.n1528 vdd.n1524 52.4337
R17682 vdd.n1531 vdd.n1530 52.4337
R17683 vdd.n1536 vdd.n1535 52.4337
R17684 vdd.n1539 vdd.n1538 52.4337
R17685 vdd.n1544 vdd.n1543 52.4337
R17686 vdd.n1547 vdd.n1546 52.4337
R17687 vdd.n1552 vdd.n1551 52.4337
R17688 vdd.n1555 vdd.n1554 52.4337
R17689 vdd.n1560 vdd.n1559 52.4337
R17690 vdd.n1563 vdd.n1562 52.4337
R17691 vdd.n1354 vdd.n1353 52.4337
R17692 vdd.n1351 vdd.n1350 52.4337
R17693 vdd.n1347 vdd.n1104 52.4337
R17694 vdd.n2085 vdd.n2084 52.4337
R17695 vdd.n1103 vdd.n1097 52.4337
R17696 vdd.n2092 vdd.n2091 52.4337
R17697 vdd.n1096 vdd.n1090 52.4337
R17698 vdd.n2099 vdd.n2098 52.4337
R17699 vdd.n1089 vdd.n1084 52.4337
R17700 vdd.n2106 vdd.n2105 52.4337
R17701 vdd.n1083 vdd.n1082 52.4337
R17702 vdd.n1078 vdd.n1071 52.4337
R17703 vdd.n2117 vdd.n2116 52.4337
R17704 vdd.n1070 vdd.n1064 52.4337
R17705 vdd.n2124 vdd.n2123 52.4337
R17706 vdd.n1063 vdd.n1057 52.4337
R17707 vdd.n2131 vdd.n2130 52.4337
R17708 vdd.n1056 vdd.n1050 52.4337
R17709 vdd.n2138 vdd.n2137 52.4337
R17710 vdd.n1049 vdd.n1044 52.4337
R17711 vdd.n2145 vdd.n2144 52.4337
R17712 vdd.n1043 vdd.n1042 52.4337
R17713 vdd.n1038 vdd.n1031 52.4337
R17714 vdd.n2156 vdd.n2155 52.4337
R17715 vdd.n1030 vdd.n1024 52.4337
R17716 vdd.n2163 vdd.n2162 52.4337
R17717 vdd.n1023 vdd.n1017 52.4337
R17718 vdd.n2170 vdd.n2169 52.4337
R17719 vdd.n1016 vdd.n1013 52.4337
R17720 vdd.n2177 vdd.n2176 52.4337
R17721 vdd.n2182 vdd.n2181 52.4337
R17722 vdd.n1358 vdd.n1012 52.4337
R17723 vdd.n3205 vdd.n3204 52.4337
R17724 vdd.n3199 vdd.n520 52.4337
R17725 vdd.n3195 vdd.n523 52.4337
R17726 vdd.n3193 vdd.n3192 52.4337
R17727 vdd.n3188 vdd.n3187 52.4337
R17728 vdd.n3185 vdd.n3184 52.4337
R17729 vdd.n3180 vdd.n3179 52.4337
R17730 vdd.n3177 vdd.n3176 52.4337
R17731 vdd.n3172 vdd.n3171 52.4337
R17732 vdd.n3169 vdd.n3168 52.4337
R17733 vdd.n3164 vdd.n3163 52.4337
R17734 vdd.n3161 vdd.n3160 52.4337
R17735 vdd.n3156 vdd.n3155 52.4337
R17736 vdd.n3153 vdd.n3152 52.4337
R17737 vdd.n3148 vdd.n3147 52.4337
R17738 vdd.n3145 vdd.n3144 52.4337
R17739 vdd.n3140 vdd.n3139 52.4337
R17740 vdd.n3137 vdd.n3136 52.4337
R17741 vdd.n3132 vdd.n3131 52.4337
R17742 vdd.n3129 vdd.n3128 52.4337
R17743 vdd.n585 vdd.n584 52.4337
R17744 vdd.n3120 vdd.n3119 52.4337
R17745 vdd.n3115 vdd.n586 52.4337
R17746 vdd.n3113 vdd.n3112 52.4337
R17747 vdd.n3108 vdd.n3107 52.4337
R17748 vdd.n3105 vdd.n3104 52.4337
R17749 vdd.n3100 vdd.n3099 52.4337
R17750 vdd.n3097 vdd.n3096 52.4337
R17751 vdd.n3092 vdd.n3091 52.4337
R17752 vdd.n3087 vdd.n607 52.4337
R17753 vdd.n3083 vdd.n609 52.4337
R17754 vdd.n3290 vdd.n462 52.4337
R17755 vdd.n3300 vdd.n3299 52.4337
R17756 vdd.n461 vdd.n455 52.4337
R17757 vdd.n3307 vdd.n3306 52.4337
R17758 vdd.n454 vdd.n448 52.4337
R17759 vdd.n3314 vdd.n3313 52.4337
R17760 vdd.n447 vdd.n441 52.4337
R17761 vdd.n3321 vdd.n3320 52.4337
R17762 vdd.n440 vdd.n435 52.4337
R17763 vdd.n3328 vdd.n3327 52.4337
R17764 vdd.n434 vdd.n433 52.4337
R17765 vdd.n429 vdd.n422 52.4337
R17766 vdd.n3339 vdd.n3338 52.4337
R17767 vdd.n421 vdd.n415 52.4337
R17768 vdd.n3346 vdd.n3345 52.4337
R17769 vdd.n414 vdd.n408 52.4337
R17770 vdd.n3353 vdd.n3352 52.4337
R17771 vdd.n407 vdd.n401 52.4337
R17772 vdd.n3360 vdd.n3359 52.4337
R17773 vdd.n400 vdd.n395 52.4337
R17774 vdd.n3367 vdd.n3366 52.4337
R17775 vdd.n394 vdd.n393 52.4337
R17776 vdd.n389 vdd.n382 52.4337
R17777 vdd.n3378 vdd.n3377 52.4337
R17778 vdd.n381 vdd.n375 52.4337
R17779 vdd.n3385 vdd.n3384 52.4337
R17780 vdd.n374 vdd.n368 52.4337
R17781 vdd.n3392 vdd.n3391 52.4337
R17782 vdd.n367 vdd.n360 52.4337
R17783 vdd.n3399 vdd.n3398 52.4337
R17784 vdd.n3402 vdd.n3401 52.4337
R17785 vdd.n355 vdd.n352 52.4337
R17786 vdd.t187 vdd.t200 51.4683
R17787 vdd.n258 vdd.n256 42.0461
R17788 vdd.n164 vdd.n162 42.0461
R17789 vdd.n71 vdd.n69 42.0461
R17790 vdd.n1959 vdd.n1957 42.0461
R17791 vdd.n1865 vdd.n1863 42.0461
R17792 vdd.n1772 vdd.n1770 42.0461
R17793 vdd.n308 vdd.n307 41.6884
R17794 vdd.n214 vdd.n213 41.6884
R17795 vdd.n121 vdd.n120 41.6884
R17796 vdd.n2009 vdd.n2008 41.6884
R17797 vdd.n1915 vdd.n1914 41.6884
R17798 vdd.n1822 vdd.n1821 41.6884
R17799 vdd.n1567 vdd.n1566 41.1157
R17800 vdd.n1604 vdd.n1603 41.1157
R17801 vdd.n1478 vdd.n1477 41.1157
R17802 vdd.n3295 vdd.n3294 41.1157
R17803 vdd.n3334 vdd.n428 41.1157
R17804 vdd.n3373 vdd.n388 41.1157
R17805 vdd.n3037 vdd.n3036 39.2114
R17806 vdd.n3034 vdd.n3033 39.2114
R17807 vdd.n3029 vdd.n641 39.2114
R17808 vdd.n3027 vdd.n3026 39.2114
R17809 vdd.n3022 vdd.n644 39.2114
R17810 vdd.n3020 vdd.n3019 39.2114
R17811 vdd.n3015 vdd.n647 39.2114
R17812 vdd.n3013 vdd.n3012 39.2114
R17813 vdd.n3007 vdd.n650 39.2114
R17814 vdd.n3005 vdd.n3004 39.2114
R17815 vdd.n3000 vdd.n653 39.2114
R17816 vdd.n2998 vdd.n2997 39.2114
R17817 vdd.n2993 vdd.n656 39.2114
R17818 vdd.n2991 vdd.n2990 39.2114
R17819 vdd.n2986 vdd.n659 39.2114
R17820 vdd.n2984 vdd.n2983 39.2114
R17821 vdd.n2979 vdd.n2978 39.2114
R17822 vdd.n2802 vdd.n2801 39.2114
R17823 vdd.n2531 vdd.n2497 39.2114
R17824 vdd.n2794 vdd.n2498 39.2114
R17825 vdd.n2790 vdd.n2499 39.2114
R17826 vdd.n2786 vdd.n2500 39.2114
R17827 vdd.n2782 vdd.n2501 39.2114
R17828 vdd.n2778 vdd.n2502 39.2114
R17829 vdd.n2774 vdd.n2503 39.2114
R17830 vdd.n2770 vdd.n2504 39.2114
R17831 vdd.n2766 vdd.n2505 39.2114
R17832 vdd.n2762 vdd.n2506 39.2114
R17833 vdd.n2758 vdd.n2507 39.2114
R17834 vdd.n2754 vdd.n2508 39.2114
R17835 vdd.n2750 vdd.n2509 39.2114
R17836 vdd.n2746 vdd.n2510 39.2114
R17837 vdd.n2742 vdd.n2511 39.2114
R17838 vdd.n2737 vdd.n2512 39.2114
R17839 vdd.n2491 vdd.n825 39.2114
R17840 vdd.n2487 vdd.n824 39.2114
R17841 vdd.n2483 vdd.n823 39.2114
R17842 vdd.n2479 vdd.n822 39.2114
R17843 vdd.n2475 vdd.n821 39.2114
R17844 vdd.n2471 vdd.n820 39.2114
R17845 vdd.n2467 vdd.n819 39.2114
R17846 vdd.n2463 vdd.n818 39.2114
R17847 vdd.n2459 vdd.n817 39.2114
R17848 vdd.n2455 vdd.n816 39.2114
R17849 vdd.n2451 vdd.n815 39.2114
R17850 vdd.n2447 vdd.n814 39.2114
R17851 vdd.n2443 vdd.n813 39.2114
R17852 vdd.n2439 vdd.n812 39.2114
R17853 vdd.n2435 vdd.n811 39.2114
R17854 vdd.n2430 vdd.n810 39.2114
R17855 vdd.n2426 vdd.n809 39.2114
R17856 vdd.n2220 vdd.n2219 39.2114
R17857 vdd.n1004 vdd.n970 39.2114
R17858 vdd.n2212 vdd.n971 39.2114
R17859 vdd.n2208 vdd.n972 39.2114
R17860 vdd.n2204 vdd.n973 39.2114
R17861 vdd.n2200 vdd.n974 39.2114
R17862 vdd.n2196 vdd.n975 39.2114
R17863 vdd.n2192 vdd.n976 39.2114
R17864 vdd.n2188 vdd.n977 39.2114
R17865 vdd.n1150 vdd.n978 39.2114
R17866 vdd.n1154 vdd.n979 39.2114
R17867 vdd.n1158 vdd.n980 39.2114
R17868 vdd.n1162 vdd.n981 39.2114
R17869 vdd.n1166 vdd.n982 39.2114
R17870 vdd.n1170 vdd.n983 39.2114
R17871 vdd.n1174 vdd.n984 39.2114
R17872 vdd.n1179 vdd.n985 39.2114
R17873 vdd.n2956 vdd.n2955 39.2114
R17874 vdd.n2951 vdd.n2923 39.2114
R17875 vdd.n2949 vdd.n2948 39.2114
R17876 vdd.n2944 vdd.n2926 39.2114
R17877 vdd.n2942 vdd.n2941 39.2114
R17878 vdd.n2937 vdd.n2929 39.2114
R17879 vdd.n2935 vdd.n2934 39.2114
R17880 vdd.n2930 vdd.n612 39.2114
R17881 vdd.n3074 vdd.n3073 39.2114
R17882 vdd.n3071 vdd.n3070 39.2114
R17883 vdd.n3066 vdd.n617 39.2114
R17884 vdd.n3064 vdd.n3063 39.2114
R17885 vdd.n3059 vdd.n620 39.2114
R17886 vdd.n3057 vdd.n3056 39.2114
R17887 vdd.n3052 vdd.n623 39.2114
R17888 vdd.n3050 vdd.n3049 39.2114
R17889 vdd.n3045 vdd.n629 39.2114
R17890 vdd.n2538 vdd.n2513 39.2114
R17891 vdd.n2542 vdd.n2514 39.2114
R17892 vdd.n2546 vdd.n2515 39.2114
R17893 vdd.n2550 vdd.n2516 39.2114
R17894 vdd.n2554 vdd.n2517 39.2114
R17895 vdd.n2558 vdd.n2518 39.2114
R17896 vdd.n2562 vdd.n2519 39.2114
R17897 vdd.n2566 vdd.n2520 39.2114
R17898 vdd.n2570 vdd.n2521 39.2114
R17899 vdd.n2574 vdd.n2522 39.2114
R17900 vdd.n2578 vdd.n2523 39.2114
R17901 vdd.n2582 vdd.n2524 39.2114
R17902 vdd.n2586 vdd.n2525 39.2114
R17903 vdd.n2590 vdd.n2526 39.2114
R17904 vdd.n2594 vdd.n2527 39.2114
R17905 vdd.n2598 vdd.n2528 39.2114
R17906 vdd.n2602 vdd.n2529 39.2114
R17907 vdd.n2541 vdd.n2513 39.2114
R17908 vdd.n2545 vdd.n2514 39.2114
R17909 vdd.n2549 vdd.n2515 39.2114
R17910 vdd.n2553 vdd.n2516 39.2114
R17911 vdd.n2557 vdd.n2517 39.2114
R17912 vdd.n2561 vdd.n2518 39.2114
R17913 vdd.n2565 vdd.n2519 39.2114
R17914 vdd.n2569 vdd.n2520 39.2114
R17915 vdd.n2573 vdd.n2521 39.2114
R17916 vdd.n2577 vdd.n2522 39.2114
R17917 vdd.n2581 vdd.n2523 39.2114
R17918 vdd.n2585 vdd.n2524 39.2114
R17919 vdd.n2589 vdd.n2525 39.2114
R17920 vdd.n2593 vdd.n2526 39.2114
R17921 vdd.n2597 vdd.n2527 39.2114
R17922 vdd.n2601 vdd.n2528 39.2114
R17923 vdd.n2604 vdd.n2529 39.2114
R17924 vdd.n629 vdd.n624 39.2114
R17925 vdd.n3051 vdd.n3050 39.2114
R17926 vdd.n623 vdd.n621 39.2114
R17927 vdd.n3058 vdd.n3057 39.2114
R17928 vdd.n620 vdd.n618 39.2114
R17929 vdd.n3065 vdd.n3064 39.2114
R17930 vdd.n617 vdd.n615 39.2114
R17931 vdd.n3072 vdd.n3071 39.2114
R17932 vdd.n3075 vdd.n3074 39.2114
R17933 vdd.n2931 vdd.n2930 39.2114
R17934 vdd.n2936 vdd.n2935 39.2114
R17935 vdd.n2929 vdd.n2927 39.2114
R17936 vdd.n2943 vdd.n2942 39.2114
R17937 vdd.n2926 vdd.n2924 39.2114
R17938 vdd.n2950 vdd.n2949 39.2114
R17939 vdd.n2923 vdd.n2921 39.2114
R17940 vdd.n2957 vdd.n2956 39.2114
R17941 vdd.n2219 vdd.n968 39.2114
R17942 vdd.n2213 vdd.n970 39.2114
R17943 vdd.n2209 vdd.n971 39.2114
R17944 vdd.n2205 vdd.n972 39.2114
R17945 vdd.n2201 vdd.n973 39.2114
R17946 vdd.n2197 vdd.n974 39.2114
R17947 vdd.n2193 vdd.n975 39.2114
R17948 vdd.n2189 vdd.n976 39.2114
R17949 vdd.n1149 vdd.n977 39.2114
R17950 vdd.n1153 vdd.n978 39.2114
R17951 vdd.n1157 vdd.n979 39.2114
R17952 vdd.n1161 vdd.n980 39.2114
R17953 vdd.n1165 vdd.n981 39.2114
R17954 vdd.n1169 vdd.n982 39.2114
R17955 vdd.n1173 vdd.n983 39.2114
R17956 vdd.n1178 vdd.n984 39.2114
R17957 vdd.n1182 vdd.n985 39.2114
R17958 vdd.n2429 vdd.n809 39.2114
R17959 vdd.n2434 vdd.n810 39.2114
R17960 vdd.n2438 vdd.n811 39.2114
R17961 vdd.n2442 vdd.n812 39.2114
R17962 vdd.n2446 vdd.n813 39.2114
R17963 vdd.n2450 vdd.n814 39.2114
R17964 vdd.n2454 vdd.n815 39.2114
R17965 vdd.n2458 vdd.n816 39.2114
R17966 vdd.n2462 vdd.n817 39.2114
R17967 vdd.n2466 vdd.n818 39.2114
R17968 vdd.n2470 vdd.n819 39.2114
R17969 vdd.n2474 vdd.n820 39.2114
R17970 vdd.n2478 vdd.n821 39.2114
R17971 vdd.n2482 vdd.n822 39.2114
R17972 vdd.n2486 vdd.n823 39.2114
R17973 vdd.n2490 vdd.n824 39.2114
R17974 vdd.n827 vdd.n825 39.2114
R17975 vdd.n2801 vdd.n790 39.2114
R17976 vdd.n2795 vdd.n2497 39.2114
R17977 vdd.n2791 vdd.n2498 39.2114
R17978 vdd.n2787 vdd.n2499 39.2114
R17979 vdd.n2783 vdd.n2500 39.2114
R17980 vdd.n2779 vdd.n2501 39.2114
R17981 vdd.n2775 vdd.n2502 39.2114
R17982 vdd.n2771 vdd.n2503 39.2114
R17983 vdd.n2767 vdd.n2504 39.2114
R17984 vdd.n2763 vdd.n2505 39.2114
R17985 vdd.n2759 vdd.n2506 39.2114
R17986 vdd.n2755 vdd.n2507 39.2114
R17987 vdd.n2751 vdd.n2508 39.2114
R17988 vdd.n2747 vdd.n2509 39.2114
R17989 vdd.n2743 vdd.n2510 39.2114
R17990 vdd.n2738 vdd.n2511 39.2114
R17991 vdd.n2734 vdd.n2512 39.2114
R17992 vdd.n2978 vdd.n660 39.2114
R17993 vdd.n2985 vdd.n2984 39.2114
R17994 vdd.n659 vdd.n657 39.2114
R17995 vdd.n2992 vdd.n2991 39.2114
R17996 vdd.n656 vdd.n654 39.2114
R17997 vdd.n2999 vdd.n2998 39.2114
R17998 vdd.n653 vdd.n651 39.2114
R17999 vdd.n3006 vdd.n3005 39.2114
R18000 vdd.n650 vdd.n648 39.2114
R18001 vdd.n3014 vdd.n3013 39.2114
R18002 vdd.n647 vdd.n645 39.2114
R18003 vdd.n3021 vdd.n3020 39.2114
R18004 vdd.n644 vdd.n642 39.2114
R18005 vdd.n3028 vdd.n3027 39.2114
R18006 vdd.n641 vdd.n639 39.2114
R18007 vdd.n3035 vdd.n3034 39.2114
R18008 vdd.n3038 vdd.n3037 39.2114
R18009 vdd.n836 vdd.n791 39.2114
R18010 vdd.n2418 vdd.n792 39.2114
R18011 vdd.n2414 vdd.n793 39.2114
R18012 vdd.n2410 vdd.n794 39.2114
R18013 vdd.n2406 vdd.n795 39.2114
R18014 vdd.n2402 vdd.n796 39.2114
R18015 vdd.n2398 vdd.n797 39.2114
R18016 vdd.n2394 vdd.n798 39.2114
R18017 vdd.n2390 vdd.n799 39.2114
R18018 vdd.n2386 vdd.n800 39.2114
R18019 vdd.n2382 vdd.n801 39.2114
R18020 vdd.n2378 vdd.n802 39.2114
R18021 vdd.n2374 vdd.n803 39.2114
R18022 vdd.n2370 vdd.n804 39.2114
R18023 vdd.n2366 vdd.n805 39.2114
R18024 vdd.n2362 vdd.n806 39.2114
R18025 vdd.n2358 vdd.n807 39.2114
R18026 vdd.n1108 vdd.n986 39.2114
R18027 vdd.n1112 vdd.n987 39.2114
R18028 vdd.n1116 vdd.n988 39.2114
R18029 vdd.n1120 vdd.n989 39.2114
R18030 vdd.n1124 vdd.n990 39.2114
R18031 vdd.n1128 vdd.n991 39.2114
R18032 vdd.n1132 vdd.n992 39.2114
R18033 vdd.n1136 vdd.n993 39.2114
R18034 vdd.n1140 vdd.n994 39.2114
R18035 vdd.n1341 vdd.n995 39.2114
R18036 vdd.n1338 vdd.n996 39.2114
R18037 vdd.n1334 vdd.n997 39.2114
R18038 vdd.n1330 vdd.n998 39.2114
R18039 vdd.n1326 vdd.n999 39.2114
R18040 vdd.n1322 vdd.n1000 39.2114
R18041 vdd.n1318 vdd.n1001 39.2114
R18042 vdd.n1314 vdd.n1002 39.2114
R18043 vdd.n2355 vdd.n807 39.2114
R18044 vdd.n2359 vdd.n806 39.2114
R18045 vdd.n2363 vdd.n805 39.2114
R18046 vdd.n2367 vdd.n804 39.2114
R18047 vdd.n2371 vdd.n803 39.2114
R18048 vdd.n2375 vdd.n802 39.2114
R18049 vdd.n2379 vdd.n801 39.2114
R18050 vdd.n2383 vdd.n800 39.2114
R18051 vdd.n2387 vdd.n799 39.2114
R18052 vdd.n2391 vdd.n798 39.2114
R18053 vdd.n2395 vdd.n797 39.2114
R18054 vdd.n2399 vdd.n796 39.2114
R18055 vdd.n2403 vdd.n795 39.2114
R18056 vdd.n2407 vdd.n794 39.2114
R18057 vdd.n2411 vdd.n793 39.2114
R18058 vdd.n2415 vdd.n792 39.2114
R18059 vdd.n2419 vdd.n791 39.2114
R18060 vdd.n1111 vdd.n986 39.2114
R18061 vdd.n1115 vdd.n987 39.2114
R18062 vdd.n1119 vdd.n988 39.2114
R18063 vdd.n1123 vdd.n989 39.2114
R18064 vdd.n1127 vdd.n990 39.2114
R18065 vdd.n1131 vdd.n991 39.2114
R18066 vdd.n1135 vdd.n992 39.2114
R18067 vdd.n1139 vdd.n993 39.2114
R18068 vdd.n1142 vdd.n994 39.2114
R18069 vdd.n1339 vdd.n995 39.2114
R18070 vdd.n1335 vdd.n996 39.2114
R18071 vdd.n1331 vdd.n997 39.2114
R18072 vdd.n1327 vdd.n998 39.2114
R18073 vdd.n1323 vdd.n999 39.2114
R18074 vdd.n1319 vdd.n1000 39.2114
R18075 vdd.n1315 vdd.n1001 39.2114
R18076 vdd.n1311 vdd.n1002 39.2114
R18077 vdd.n2076 vdd.n2075 37.2369
R18078 vdd.n2112 vdd.n1077 37.2369
R18079 vdd.n2151 vdd.n1037 37.2369
R18080 vdd.n3126 vdd.n581 37.2369
R18081 vdd.n545 vdd.n544 37.2369
R18082 vdd.n3082 vdd.n3081 37.2369
R18083 vdd.n1145 vdd.n1144 30.449
R18084 vdd.n840 vdd.n839 30.449
R18085 vdd.n1176 vdd.n1148 30.449
R18086 vdd.n2432 vdd.n830 30.449
R18087 vdd.n2537 vdd.n2536 30.449
R18088 vdd.n663 vdd.n662 30.449
R18089 vdd.n2740 vdd.n2533 30.449
R18090 vdd.n627 vdd.n626 30.449
R18091 vdd.n2222 vdd.n2221 29.8151
R18092 vdd.n2494 vdd.n828 29.8151
R18093 vdd.n2427 vdd.n831 29.8151
R18094 vdd.n1184 vdd.n1181 29.8151
R18095 vdd.n2735 vdd.n2732 29.8151
R18096 vdd.n2980 vdd.n2977 29.8151
R18097 vdd.n2804 vdd.n2803 29.8151
R18098 vdd.n3041 vdd.n3040 29.8151
R18099 vdd.n2960 vdd.n2959 29.8151
R18100 vdd.n3046 vdd.n628 29.8151
R18101 vdd.n2608 vdd.n2606 29.8151
R18102 vdd.n2539 vdd.n783 29.8151
R18103 vdd.n1109 vdd.n960 29.8151
R18104 vdd.n2422 vdd.n2421 29.8151
R18105 vdd.n2354 vdd.n2353 29.8151
R18106 vdd.n1310 vdd.n1309 29.8151
R18107 vdd.n1670 vdd.n1437 20.633
R18108 vdd.n2070 vdd.n969 20.633
R18109 vdd.n3212 vdd.n516 20.633
R18110 vdd.n3410 vdd.n351 20.633
R18111 vdd.n1672 vdd.n1434 19.3944
R18112 vdd.n1676 vdd.n1434 19.3944
R18113 vdd.n1676 vdd.n1425 19.3944
R18114 vdd.n1688 vdd.n1425 19.3944
R18115 vdd.n1688 vdd.n1423 19.3944
R18116 vdd.n1692 vdd.n1423 19.3944
R18117 vdd.n1692 vdd.n1412 19.3944
R18118 vdd.n1704 vdd.n1412 19.3944
R18119 vdd.n1704 vdd.n1410 19.3944
R18120 vdd.n1708 vdd.n1410 19.3944
R18121 vdd.n1708 vdd.n1401 19.3944
R18122 vdd.n1721 vdd.n1401 19.3944
R18123 vdd.n1721 vdd.n1399 19.3944
R18124 vdd.n1725 vdd.n1399 19.3944
R18125 vdd.n1725 vdd.n1390 19.3944
R18126 vdd.n2019 vdd.n1390 19.3944
R18127 vdd.n2019 vdd.n1388 19.3944
R18128 vdd.n2023 vdd.n1388 19.3944
R18129 vdd.n2023 vdd.n1378 19.3944
R18130 vdd.n2036 vdd.n1378 19.3944
R18131 vdd.n2036 vdd.n1376 19.3944
R18132 vdd.n2040 vdd.n1376 19.3944
R18133 vdd.n2040 vdd.n1368 19.3944
R18134 vdd.n2053 vdd.n1368 19.3944
R18135 vdd.n2053 vdd.n1365 19.3944
R18136 vdd.n2059 vdd.n1365 19.3944
R18137 vdd.n2059 vdd.n1366 19.3944
R18138 vdd.n1366 vdd.n1356 19.3944
R18139 vdd.n1597 vdd.n1523 19.3944
R18140 vdd.n1597 vdd.n1525 19.3944
R18141 vdd.n1593 vdd.n1525 19.3944
R18142 vdd.n1593 vdd.n1592 19.3944
R18143 vdd.n1592 vdd.n1591 19.3944
R18144 vdd.n1591 vdd.n1533 19.3944
R18145 vdd.n1587 vdd.n1533 19.3944
R18146 vdd.n1587 vdd.n1586 19.3944
R18147 vdd.n1586 vdd.n1585 19.3944
R18148 vdd.n1585 vdd.n1541 19.3944
R18149 vdd.n1581 vdd.n1541 19.3944
R18150 vdd.n1581 vdd.n1580 19.3944
R18151 vdd.n1580 vdd.n1579 19.3944
R18152 vdd.n1579 vdd.n1549 19.3944
R18153 vdd.n1575 vdd.n1549 19.3944
R18154 vdd.n1575 vdd.n1574 19.3944
R18155 vdd.n1574 vdd.n1573 19.3944
R18156 vdd.n1573 vdd.n1557 19.3944
R18157 vdd.n1569 vdd.n1557 19.3944
R18158 vdd.n1569 vdd.n1568 19.3944
R18159 vdd.n1635 vdd.n1634 19.3944
R18160 vdd.n1634 vdd.n1633 19.3944
R18161 vdd.n1633 vdd.n1486 19.3944
R18162 vdd.n1629 vdd.n1486 19.3944
R18163 vdd.n1629 vdd.n1628 19.3944
R18164 vdd.n1628 vdd.n1627 19.3944
R18165 vdd.n1627 vdd.n1494 19.3944
R18166 vdd.n1623 vdd.n1494 19.3944
R18167 vdd.n1623 vdd.n1622 19.3944
R18168 vdd.n1622 vdd.n1621 19.3944
R18169 vdd.n1621 vdd.n1502 19.3944
R18170 vdd.n1617 vdd.n1502 19.3944
R18171 vdd.n1617 vdd.n1616 19.3944
R18172 vdd.n1616 vdd.n1615 19.3944
R18173 vdd.n1615 vdd.n1510 19.3944
R18174 vdd.n1611 vdd.n1510 19.3944
R18175 vdd.n1611 vdd.n1610 19.3944
R18176 vdd.n1610 vdd.n1609 19.3944
R18177 vdd.n1609 vdd.n1518 19.3944
R18178 vdd.n1605 vdd.n1518 19.3944
R18179 vdd.n1665 vdd.n1664 19.3944
R18180 vdd.n1664 vdd.n1663 19.3944
R18181 vdd.n1663 vdd.n1444 19.3944
R18182 vdd.n1659 vdd.n1444 19.3944
R18183 vdd.n1659 vdd.n1658 19.3944
R18184 vdd.n1658 vdd.n1657 19.3944
R18185 vdd.n1657 vdd.n1452 19.3944
R18186 vdd.n1653 vdd.n1452 19.3944
R18187 vdd.n1653 vdd.n1652 19.3944
R18188 vdd.n1652 vdd.n1651 19.3944
R18189 vdd.n1651 vdd.n1460 19.3944
R18190 vdd.n1647 vdd.n1460 19.3944
R18191 vdd.n1647 vdd.n1646 19.3944
R18192 vdd.n1646 vdd.n1645 19.3944
R18193 vdd.n1645 vdd.n1468 19.3944
R18194 vdd.n1641 vdd.n1468 19.3944
R18195 vdd.n1641 vdd.n1640 19.3944
R18196 vdd.n1640 vdd.n1639 19.3944
R18197 vdd.n2108 vdd.n1075 19.3944
R18198 vdd.n2108 vdd.n1081 19.3944
R18199 vdd.n2103 vdd.n1081 19.3944
R18200 vdd.n2103 vdd.n2102 19.3944
R18201 vdd.n2102 vdd.n2101 19.3944
R18202 vdd.n2101 vdd.n1088 19.3944
R18203 vdd.n2096 vdd.n1088 19.3944
R18204 vdd.n2096 vdd.n2095 19.3944
R18205 vdd.n2095 vdd.n2094 19.3944
R18206 vdd.n2094 vdd.n1095 19.3944
R18207 vdd.n2089 vdd.n1095 19.3944
R18208 vdd.n2089 vdd.n2088 19.3944
R18209 vdd.n2088 vdd.n2087 19.3944
R18210 vdd.n2087 vdd.n1102 19.3944
R18211 vdd.n2082 vdd.n1102 19.3944
R18212 vdd.n2082 vdd.n2081 19.3944
R18213 vdd.n1349 vdd.n1107 19.3944
R18214 vdd.n2077 vdd.n1346 19.3944
R18215 vdd.n2147 vdd.n1035 19.3944
R18216 vdd.n2147 vdd.n1041 19.3944
R18217 vdd.n2142 vdd.n1041 19.3944
R18218 vdd.n2142 vdd.n2141 19.3944
R18219 vdd.n2141 vdd.n2140 19.3944
R18220 vdd.n2140 vdd.n1048 19.3944
R18221 vdd.n2135 vdd.n1048 19.3944
R18222 vdd.n2135 vdd.n2134 19.3944
R18223 vdd.n2134 vdd.n2133 19.3944
R18224 vdd.n2133 vdd.n1055 19.3944
R18225 vdd.n2128 vdd.n1055 19.3944
R18226 vdd.n2128 vdd.n2127 19.3944
R18227 vdd.n2127 vdd.n2126 19.3944
R18228 vdd.n2126 vdd.n1062 19.3944
R18229 vdd.n2121 vdd.n1062 19.3944
R18230 vdd.n2121 vdd.n2120 19.3944
R18231 vdd.n2120 vdd.n2119 19.3944
R18232 vdd.n2119 vdd.n1069 19.3944
R18233 vdd.n2114 vdd.n1069 19.3944
R18234 vdd.n2114 vdd.n2113 19.3944
R18235 vdd.n2184 vdd.n1010 19.3944
R18236 vdd.n2184 vdd.n1011 19.3944
R18237 vdd.n2179 vdd.n2178 19.3944
R18238 vdd.n2174 vdd.n2173 19.3944
R18239 vdd.n2173 vdd.n2172 19.3944
R18240 vdd.n2172 vdd.n1015 19.3944
R18241 vdd.n2167 vdd.n1015 19.3944
R18242 vdd.n2167 vdd.n2166 19.3944
R18243 vdd.n2166 vdd.n2165 19.3944
R18244 vdd.n2165 vdd.n1022 19.3944
R18245 vdd.n2160 vdd.n1022 19.3944
R18246 vdd.n2160 vdd.n2159 19.3944
R18247 vdd.n2159 vdd.n2158 19.3944
R18248 vdd.n2158 vdd.n1029 19.3944
R18249 vdd.n2153 vdd.n1029 19.3944
R18250 vdd.n2153 vdd.n2152 19.3944
R18251 vdd.n1668 vdd.n1431 19.3944
R18252 vdd.n1680 vdd.n1431 19.3944
R18253 vdd.n1680 vdd.n1429 19.3944
R18254 vdd.n1684 vdd.n1429 19.3944
R18255 vdd.n1684 vdd.n1419 19.3944
R18256 vdd.n1696 vdd.n1419 19.3944
R18257 vdd.n1696 vdd.n1417 19.3944
R18258 vdd.n1700 vdd.n1417 19.3944
R18259 vdd.n1700 vdd.n1407 19.3944
R18260 vdd.n1713 vdd.n1407 19.3944
R18261 vdd.n1713 vdd.n1405 19.3944
R18262 vdd.n1717 vdd.n1405 19.3944
R18263 vdd.n1717 vdd.n1396 19.3944
R18264 vdd.n1729 vdd.n1396 19.3944
R18265 vdd.n1729 vdd.n1394 19.3944
R18266 vdd.n2015 vdd.n1394 19.3944
R18267 vdd.n2015 vdd.n1384 19.3944
R18268 vdd.n2028 vdd.n1384 19.3944
R18269 vdd.n2028 vdd.n1382 19.3944
R18270 vdd.n2032 vdd.n1382 19.3944
R18271 vdd.n2032 vdd.n1373 19.3944
R18272 vdd.n2045 vdd.n1373 19.3944
R18273 vdd.n2045 vdd.n1371 19.3944
R18274 vdd.n2049 vdd.n1371 19.3944
R18275 vdd.n2049 vdd.n1361 19.3944
R18276 vdd.n2064 vdd.n1361 19.3944
R18277 vdd.n2064 vdd.n1359 19.3944
R18278 vdd.n2068 vdd.n1359 19.3944
R18279 vdd.n3214 vdd.n513 19.3944
R18280 vdd.n3218 vdd.n513 19.3944
R18281 vdd.n3218 vdd.n503 19.3944
R18282 vdd.n3230 vdd.n503 19.3944
R18283 vdd.n3230 vdd.n501 19.3944
R18284 vdd.n3234 vdd.n501 19.3944
R18285 vdd.n3234 vdd.n490 19.3944
R18286 vdd.n3246 vdd.n490 19.3944
R18287 vdd.n3246 vdd.n488 19.3944
R18288 vdd.n3250 vdd.n488 19.3944
R18289 vdd.n3250 vdd.n478 19.3944
R18290 vdd.n3263 vdd.n478 19.3944
R18291 vdd.n3263 vdd.n476 19.3944
R18292 vdd.n3267 vdd.n476 19.3944
R18293 vdd.n3268 vdd.n3267 19.3944
R18294 vdd.n3269 vdd.n3268 19.3944
R18295 vdd.n3269 vdd.n474 19.3944
R18296 vdd.n3273 vdd.n474 19.3944
R18297 vdd.n3274 vdd.n3273 19.3944
R18298 vdd.n3275 vdd.n3274 19.3944
R18299 vdd.n3275 vdd.n471 19.3944
R18300 vdd.n3279 vdd.n471 19.3944
R18301 vdd.n3280 vdd.n3279 19.3944
R18302 vdd.n3281 vdd.n3280 19.3944
R18303 vdd.n3281 vdd.n468 19.3944
R18304 vdd.n3285 vdd.n468 19.3944
R18305 vdd.n3286 vdd.n3285 19.3944
R18306 vdd.n3287 vdd.n3286 19.3944
R18307 vdd.n3330 vdd.n426 19.3944
R18308 vdd.n3330 vdd.n432 19.3944
R18309 vdd.n3325 vdd.n432 19.3944
R18310 vdd.n3325 vdd.n3324 19.3944
R18311 vdd.n3324 vdd.n3323 19.3944
R18312 vdd.n3323 vdd.n439 19.3944
R18313 vdd.n3318 vdd.n439 19.3944
R18314 vdd.n3318 vdd.n3317 19.3944
R18315 vdd.n3317 vdd.n3316 19.3944
R18316 vdd.n3316 vdd.n446 19.3944
R18317 vdd.n3311 vdd.n446 19.3944
R18318 vdd.n3311 vdd.n3310 19.3944
R18319 vdd.n3310 vdd.n3309 19.3944
R18320 vdd.n3309 vdd.n453 19.3944
R18321 vdd.n3304 vdd.n453 19.3944
R18322 vdd.n3304 vdd.n3303 19.3944
R18323 vdd.n3303 vdd.n3302 19.3944
R18324 vdd.n3302 vdd.n460 19.3944
R18325 vdd.n3297 vdd.n460 19.3944
R18326 vdd.n3297 vdd.n3296 19.3944
R18327 vdd.n3369 vdd.n386 19.3944
R18328 vdd.n3369 vdd.n392 19.3944
R18329 vdd.n3364 vdd.n392 19.3944
R18330 vdd.n3364 vdd.n3363 19.3944
R18331 vdd.n3363 vdd.n3362 19.3944
R18332 vdd.n3362 vdd.n399 19.3944
R18333 vdd.n3357 vdd.n399 19.3944
R18334 vdd.n3357 vdd.n3356 19.3944
R18335 vdd.n3356 vdd.n3355 19.3944
R18336 vdd.n3355 vdd.n406 19.3944
R18337 vdd.n3350 vdd.n406 19.3944
R18338 vdd.n3350 vdd.n3349 19.3944
R18339 vdd.n3349 vdd.n3348 19.3944
R18340 vdd.n3348 vdd.n413 19.3944
R18341 vdd.n3343 vdd.n413 19.3944
R18342 vdd.n3343 vdd.n3342 19.3944
R18343 vdd.n3342 vdd.n3341 19.3944
R18344 vdd.n3341 vdd.n420 19.3944
R18345 vdd.n3336 vdd.n420 19.3944
R18346 vdd.n3336 vdd.n3335 19.3944
R18347 vdd.n3405 vdd.n3404 19.3944
R18348 vdd.n3404 vdd.n3403 19.3944
R18349 vdd.n3403 vdd.n358 19.3944
R18350 vdd.n359 vdd.n358 19.3944
R18351 vdd.n3396 vdd.n359 19.3944
R18352 vdd.n3396 vdd.n3395 19.3944
R18353 vdd.n3395 vdd.n3394 19.3944
R18354 vdd.n3394 vdd.n366 19.3944
R18355 vdd.n3389 vdd.n366 19.3944
R18356 vdd.n3389 vdd.n3388 19.3944
R18357 vdd.n3388 vdd.n3387 19.3944
R18358 vdd.n3387 vdd.n373 19.3944
R18359 vdd.n3382 vdd.n373 19.3944
R18360 vdd.n3382 vdd.n3381 19.3944
R18361 vdd.n3381 vdd.n3380 19.3944
R18362 vdd.n3380 vdd.n380 19.3944
R18363 vdd.n3375 vdd.n380 19.3944
R18364 vdd.n3375 vdd.n3374 19.3944
R18365 vdd.n3210 vdd.n509 19.3944
R18366 vdd.n3222 vdd.n509 19.3944
R18367 vdd.n3222 vdd.n507 19.3944
R18368 vdd.n3226 vdd.n507 19.3944
R18369 vdd.n3226 vdd.n497 19.3944
R18370 vdd.n3238 vdd.n497 19.3944
R18371 vdd.n3238 vdd.n495 19.3944
R18372 vdd.n3242 vdd.n495 19.3944
R18373 vdd.n3242 vdd.n485 19.3944
R18374 vdd.n3255 vdd.n485 19.3944
R18375 vdd.n3255 vdd.n483 19.3944
R18376 vdd.n3259 vdd.n483 19.3944
R18377 vdd.n3259 vdd.n312 19.3944
R18378 vdd.n3438 vdd.n312 19.3944
R18379 vdd.n3438 vdd.n313 19.3944
R18380 vdd.n3432 vdd.n313 19.3944
R18381 vdd.n3432 vdd.n3431 19.3944
R18382 vdd.n3431 vdd.n3430 19.3944
R18383 vdd.n3430 vdd.n323 19.3944
R18384 vdd.n3424 vdd.n323 19.3944
R18385 vdd.n3424 vdd.n3423 19.3944
R18386 vdd.n3423 vdd.n3422 19.3944
R18387 vdd.n3422 vdd.n335 19.3944
R18388 vdd.n3416 vdd.n335 19.3944
R18389 vdd.n3416 vdd.n3415 19.3944
R18390 vdd.n3415 vdd.n3414 19.3944
R18391 vdd.n3414 vdd.n346 19.3944
R18392 vdd.n3408 vdd.n346 19.3944
R18393 vdd.n3167 vdd.n3166 19.3944
R18394 vdd.n3166 vdd.n3165 19.3944
R18395 vdd.n3165 vdd.n551 19.3944
R18396 vdd.n3159 vdd.n551 19.3944
R18397 vdd.n3159 vdd.n3158 19.3944
R18398 vdd.n3158 vdd.n3157 19.3944
R18399 vdd.n3157 vdd.n557 19.3944
R18400 vdd.n3151 vdd.n557 19.3944
R18401 vdd.n3151 vdd.n3150 19.3944
R18402 vdd.n3150 vdd.n3149 19.3944
R18403 vdd.n3149 vdd.n563 19.3944
R18404 vdd.n3143 vdd.n563 19.3944
R18405 vdd.n3143 vdd.n3142 19.3944
R18406 vdd.n3142 vdd.n3141 19.3944
R18407 vdd.n3141 vdd.n569 19.3944
R18408 vdd.n3135 vdd.n569 19.3944
R18409 vdd.n3135 vdd.n3134 19.3944
R18410 vdd.n3134 vdd.n3133 19.3944
R18411 vdd.n3133 vdd.n575 19.3944
R18412 vdd.n3127 vdd.n575 19.3944
R18413 vdd.n3207 vdd.n3206 19.3944
R18414 vdd.n3206 vdd.n519 19.3944
R18415 vdd.n3201 vdd.n3200 19.3944
R18416 vdd.n3197 vdd.n3196 19.3944
R18417 vdd.n3196 vdd.n525 19.3944
R18418 vdd.n3191 vdd.n525 19.3944
R18419 vdd.n3191 vdd.n3190 19.3944
R18420 vdd.n3190 vdd.n3189 19.3944
R18421 vdd.n3189 vdd.n531 19.3944
R18422 vdd.n3183 vdd.n531 19.3944
R18423 vdd.n3183 vdd.n3182 19.3944
R18424 vdd.n3182 vdd.n3181 19.3944
R18425 vdd.n3181 vdd.n537 19.3944
R18426 vdd.n3175 vdd.n537 19.3944
R18427 vdd.n3175 vdd.n3174 19.3944
R18428 vdd.n3174 vdd.n3173 19.3944
R18429 vdd.n3122 vdd.n579 19.3944
R18430 vdd.n3122 vdd.n583 19.3944
R18431 vdd.n3117 vdd.n583 19.3944
R18432 vdd.n3117 vdd.n3116 19.3944
R18433 vdd.n3116 vdd.n589 19.3944
R18434 vdd.n3111 vdd.n589 19.3944
R18435 vdd.n3111 vdd.n3110 19.3944
R18436 vdd.n3110 vdd.n3109 19.3944
R18437 vdd.n3109 vdd.n595 19.3944
R18438 vdd.n3103 vdd.n595 19.3944
R18439 vdd.n3103 vdd.n3102 19.3944
R18440 vdd.n3102 vdd.n3101 19.3944
R18441 vdd.n3101 vdd.n601 19.3944
R18442 vdd.n3095 vdd.n601 19.3944
R18443 vdd.n3095 vdd.n3094 19.3944
R18444 vdd.n3094 vdd.n3093 19.3944
R18445 vdd.n3089 vdd.n3088 19.3944
R18446 vdd.n3085 vdd.n3084 19.3944
R18447 vdd.n1604 vdd.n1523 19.0066
R18448 vdd.n2112 vdd.n1075 19.0066
R18449 vdd.n3334 vdd.n426 19.0066
R18450 vdd.n3126 vdd.n579 19.0066
R18451 vdd.n1144 vdd.n1143 16.0975
R18452 vdd.n839 vdd.n838 16.0975
R18453 vdd.n1566 vdd.n1565 16.0975
R18454 vdd.n1603 vdd.n1602 16.0975
R18455 vdd.n1477 vdd.n1476 16.0975
R18456 vdd.n2075 vdd.n2074 16.0975
R18457 vdd.n1077 vdd.n1076 16.0975
R18458 vdd.n1037 vdd.n1036 16.0975
R18459 vdd.n1148 vdd.n1147 16.0975
R18460 vdd.n830 vdd.n829 16.0975
R18461 vdd.n2536 vdd.n2535 16.0975
R18462 vdd.n3294 vdd.n3293 16.0975
R18463 vdd.n428 vdd.n427 16.0975
R18464 vdd.n388 vdd.n387 16.0975
R18465 vdd.n581 vdd.n580 16.0975
R18466 vdd.n544 vdd.n543 16.0975
R18467 vdd.n662 vdd.n661 16.0975
R18468 vdd.n2533 vdd.n2532 16.0975
R18469 vdd.n3081 vdd.n3080 16.0975
R18470 vdd.n626 vdd.n625 16.0975
R18471 vdd.t200 vdd.n2496 15.4182
R18472 vdd.n2800 vdd.t187 15.4182
R18473 vdd.n28 vdd.n27 14.5458
R18474 vdd.n304 vdd.n269 13.1884
R18475 vdd.n253 vdd.n218 13.1884
R18476 vdd.n210 vdd.n175 13.1884
R18477 vdd.n159 vdd.n124 13.1884
R18478 vdd.n117 vdd.n82 13.1884
R18479 vdd.n66 vdd.n31 13.1884
R18480 vdd.n1954 vdd.n1919 13.1884
R18481 vdd.n2005 vdd.n1970 13.1884
R18482 vdd.n1860 vdd.n1825 13.1884
R18483 vdd.n1911 vdd.n1876 13.1884
R18484 vdd.n1767 vdd.n1732 13.1884
R18485 vdd.n1818 vdd.n1783 13.1884
R18486 vdd.n2218 vdd.n962 13.1509
R18487 vdd.n3043 vdd.n613 13.1509
R18488 vdd.n1635 vdd.n1478 12.9944
R18489 vdd.n1639 vdd.n1478 12.9944
R18490 vdd.n2151 vdd.n1035 12.9944
R18491 vdd.n2152 vdd.n2151 12.9944
R18492 vdd.n3373 vdd.n386 12.9944
R18493 vdd.n3374 vdd.n3373 12.9944
R18494 vdd.n3167 vdd.n545 12.9944
R18495 vdd.n3173 vdd.n545 12.9944
R18496 vdd.n305 vdd.n267 12.8005
R18497 vdd.n300 vdd.n271 12.8005
R18498 vdd.n254 vdd.n216 12.8005
R18499 vdd.n249 vdd.n220 12.8005
R18500 vdd.n211 vdd.n173 12.8005
R18501 vdd.n206 vdd.n177 12.8005
R18502 vdd.n160 vdd.n122 12.8005
R18503 vdd.n155 vdd.n126 12.8005
R18504 vdd.n118 vdd.n80 12.8005
R18505 vdd.n113 vdd.n84 12.8005
R18506 vdd.n67 vdd.n29 12.8005
R18507 vdd.n62 vdd.n33 12.8005
R18508 vdd.n1955 vdd.n1917 12.8005
R18509 vdd.n1950 vdd.n1921 12.8005
R18510 vdd.n2006 vdd.n1968 12.8005
R18511 vdd.n2001 vdd.n1972 12.8005
R18512 vdd.n1861 vdd.n1823 12.8005
R18513 vdd.n1856 vdd.n1827 12.8005
R18514 vdd.n1912 vdd.n1874 12.8005
R18515 vdd.n1907 vdd.n1878 12.8005
R18516 vdd.n1768 vdd.n1730 12.8005
R18517 vdd.n1763 vdd.n1734 12.8005
R18518 vdd.n1819 vdd.n1781 12.8005
R18519 vdd.n1814 vdd.n1785 12.8005
R18520 vdd.n299 vdd.n272 12.0247
R18521 vdd.n248 vdd.n221 12.0247
R18522 vdd.n205 vdd.n178 12.0247
R18523 vdd.n154 vdd.n127 12.0247
R18524 vdd.n112 vdd.n85 12.0247
R18525 vdd.n61 vdd.n34 12.0247
R18526 vdd.n1949 vdd.n1922 12.0247
R18527 vdd.n2000 vdd.n1973 12.0247
R18528 vdd.n1855 vdd.n1828 12.0247
R18529 vdd.n1906 vdd.n1879 12.0247
R18530 vdd.n1762 vdd.n1735 12.0247
R18531 vdd.n1813 vdd.n1786 12.0247
R18532 vdd.n1670 vdd.n1438 11.337
R18533 vdd.n1678 vdd.n1427 11.337
R18534 vdd.n1686 vdd.n1427 11.337
R18535 vdd.n1694 vdd.n1421 11.337
R18536 vdd.n1702 vdd.n1414 11.337
R18537 vdd.n1711 vdd.n1710 11.337
R18538 vdd.n1719 vdd.n1403 11.337
R18539 vdd.n2017 vdd.n1392 11.337
R18540 vdd.n2026 vdd.n1386 11.337
R18541 vdd.n2034 vdd.n1380 11.337
R18542 vdd.n2043 vdd.n2042 11.337
R18543 vdd.n2051 vdd.n1363 11.337
R18544 vdd.n2062 vdd.n1363 11.337
R18545 vdd.n2062 vdd.n2061 11.337
R18546 vdd.n3220 vdd.n511 11.337
R18547 vdd.n3220 vdd.n505 11.337
R18548 vdd.n3228 vdd.n505 11.337
R18549 vdd.n3236 vdd.n499 11.337
R18550 vdd.n3244 vdd.n492 11.337
R18551 vdd.n3253 vdd.n3252 11.337
R18552 vdd.n3261 vdd.n481 11.337
R18553 vdd.n3435 vdd.n3434 11.337
R18554 vdd.n3428 vdd.n325 11.337
R18555 vdd.n3426 vdd.n329 11.337
R18556 vdd.n3420 vdd.n3419 11.337
R18557 vdd.n3418 vdd.n340 11.337
R18558 vdd.n3412 vdd.n340 11.337
R18559 vdd.n3411 vdd.n3410 11.337
R18560 vdd.n296 vdd.n295 11.249
R18561 vdd.n245 vdd.n244 11.249
R18562 vdd.n202 vdd.n201 11.249
R18563 vdd.n151 vdd.n150 11.249
R18564 vdd.n109 vdd.n108 11.249
R18565 vdd.n58 vdd.n57 11.249
R18566 vdd.n1946 vdd.n1945 11.249
R18567 vdd.n1997 vdd.n1996 11.249
R18568 vdd.n1852 vdd.n1851 11.249
R18569 vdd.n1903 vdd.n1902 11.249
R18570 vdd.n1759 vdd.n1758 11.249
R18571 vdd.n1810 vdd.n1809 11.249
R18572 vdd.n1686 vdd.t115 10.9969
R18573 vdd.t117 vdd.n3418 10.9969
R18574 vdd.n1415 vdd.t134 10.7702
R18575 vdd.t6 vdd.n3427 10.7702
R18576 vdd.n281 vdd.n280 10.7238
R18577 vdd.n230 vdd.n229 10.7238
R18578 vdd.n187 vdd.n186 10.7238
R18579 vdd.n136 vdd.n135 10.7238
R18580 vdd.n94 vdd.n93 10.7238
R18581 vdd.n43 vdd.n42 10.7238
R18582 vdd.n1931 vdd.n1930 10.7238
R18583 vdd.n1982 vdd.n1981 10.7238
R18584 vdd.n1837 vdd.n1836 10.7238
R18585 vdd.n1888 vdd.n1887 10.7238
R18586 vdd.n1744 vdd.n1743 10.7238
R18587 vdd.n1795 vdd.n1794 10.7238
R18588 vdd.n2223 vdd.n2222 10.6151
R18589 vdd.n2223 vdd.n955 10.6151
R18590 vdd.n2233 vdd.n955 10.6151
R18591 vdd.n2234 vdd.n2233 10.6151
R18592 vdd.n2235 vdd.n2234 10.6151
R18593 vdd.n2235 vdd.n942 10.6151
R18594 vdd.n2245 vdd.n942 10.6151
R18595 vdd.n2246 vdd.n2245 10.6151
R18596 vdd.n2247 vdd.n2246 10.6151
R18597 vdd.n2247 vdd.n930 10.6151
R18598 vdd.n2257 vdd.n930 10.6151
R18599 vdd.n2258 vdd.n2257 10.6151
R18600 vdd.n2259 vdd.n2258 10.6151
R18601 vdd.n2259 vdd.n919 10.6151
R18602 vdd.n2269 vdd.n919 10.6151
R18603 vdd.n2270 vdd.n2269 10.6151
R18604 vdd.n2271 vdd.n2270 10.6151
R18605 vdd.n2271 vdd.n906 10.6151
R18606 vdd.n2281 vdd.n906 10.6151
R18607 vdd.n2282 vdd.n2281 10.6151
R18608 vdd.n2283 vdd.n2282 10.6151
R18609 vdd.n2283 vdd.n894 10.6151
R18610 vdd.n2294 vdd.n894 10.6151
R18611 vdd.n2295 vdd.n2294 10.6151
R18612 vdd.n2296 vdd.n2295 10.6151
R18613 vdd.n2296 vdd.n882 10.6151
R18614 vdd.n2306 vdd.n882 10.6151
R18615 vdd.n2307 vdd.n2306 10.6151
R18616 vdd.n2308 vdd.n2307 10.6151
R18617 vdd.n2308 vdd.n870 10.6151
R18618 vdd.n2318 vdd.n870 10.6151
R18619 vdd.n2319 vdd.n2318 10.6151
R18620 vdd.n2320 vdd.n2319 10.6151
R18621 vdd.n2320 vdd.n860 10.6151
R18622 vdd.n2330 vdd.n860 10.6151
R18623 vdd.n2331 vdd.n2330 10.6151
R18624 vdd.n2332 vdd.n2331 10.6151
R18625 vdd.n2332 vdd.n847 10.6151
R18626 vdd.n2344 vdd.n847 10.6151
R18627 vdd.n2345 vdd.n2344 10.6151
R18628 vdd.n2347 vdd.n2345 10.6151
R18629 vdd.n2347 vdd.n2346 10.6151
R18630 vdd.n2346 vdd.n828 10.6151
R18631 vdd.n2494 vdd.n2493 10.6151
R18632 vdd.n2493 vdd.n2492 10.6151
R18633 vdd.n2492 vdd.n2489 10.6151
R18634 vdd.n2489 vdd.n2488 10.6151
R18635 vdd.n2488 vdd.n2485 10.6151
R18636 vdd.n2485 vdd.n2484 10.6151
R18637 vdd.n2484 vdd.n2481 10.6151
R18638 vdd.n2481 vdd.n2480 10.6151
R18639 vdd.n2480 vdd.n2477 10.6151
R18640 vdd.n2477 vdd.n2476 10.6151
R18641 vdd.n2476 vdd.n2473 10.6151
R18642 vdd.n2473 vdd.n2472 10.6151
R18643 vdd.n2472 vdd.n2469 10.6151
R18644 vdd.n2469 vdd.n2468 10.6151
R18645 vdd.n2468 vdd.n2465 10.6151
R18646 vdd.n2465 vdd.n2464 10.6151
R18647 vdd.n2464 vdd.n2461 10.6151
R18648 vdd.n2461 vdd.n2460 10.6151
R18649 vdd.n2460 vdd.n2457 10.6151
R18650 vdd.n2457 vdd.n2456 10.6151
R18651 vdd.n2456 vdd.n2453 10.6151
R18652 vdd.n2453 vdd.n2452 10.6151
R18653 vdd.n2452 vdd.n2449 10.6151
R18654 vdd.n2449 vdd.n2448 10.6151
R18655 vdd.n2448 vdd.n2445 10.6151
R18656 vdd.n2445 vdd.n2444 10.6151
R18657 vdd.n2444 vdd.n2441 10.6151
R18658 vdd.n2441 vdd.n2440 10.6151
R18659 vdd.n2440 vdd.n2437 10.6151
R18660 vdd.n2437 vdd.n2436 10.6151
R18661 vdd.n2436 vdd.n2433 10.6151
R18662 vdd.n2431 vdd.n2428 10.6151
R18663 vdd.n2428 vdd.n2427 10.6151
R18664 vdd.n1185 vdd.n1184 10.6151
R18665 vdd.n1187 vdd.n1185 10.6151
R18666 vdd.n1188 vdd.n1187 10.6151
R18667 vdd.n1190 vdd.n1188 10.6151
R18668 vdd.n1191 vdd.n1190 10.6151
R18669 vdd.n1193 vdd.n1191 10.6151
R18670 vdd.n1194 vdd.n1193 10.6151
R18671 vdd.n1196 vdd.n1194 10.6151
R18672 vdd.n1197 vdd.n1196 10.6151
R18673 vdd.n1199 vdd.n1197 10.6151
R18674 vdd.n1200 vdd.n1199 10.6151
R18675 vdd.n1202 vdd.n1200 10.6151
R18676 vdd.n1203 vdd.n1202 10.6151
R18677 vdd.n1205 vdd.n1203 10.6151
R18678 vdd.n1206 vdd.n1205 10.6151
R18679 vdd.n1208 vdd.n1206 10.6151
R18680 vdd.n1209 vdd.n1208 10.6151
R18681 vdd.n1211 vdd.n1209 10.6151
R18682 vdd.n1212 vdd.n1211 10.6151
R18683 vdd.n1214 vdd.n1212 10.6151
R18684 vdd.n1215 vdd.n1214 10.6151
R18685 vdd.n1217 vdd.n1215 10.6151
R18686 vdd.n1218 vdd.n1217 10.6151
R18687 vdd.n1220 vdd.n1218 10.6151
R18688 vdd.n1221 vdd.n1220 10.6151
R18689 vdd.n1223 vdd.n1221 10.6151
R18690 vdd.n1224 vdd.n1223 10.6151
R18691 vdd.n1263 vdd.n1224 10.6151
R18692 vdd.n1263 vdd.n1262 10.6151
R18693 vdd.n1262 vdd.n1261 10.6151
R18694 vdd.n1261 vdd.n1259 10.6151
R18695 vdd.n1259 vdd.n1258 10.6151
R18696 vdd.n1258 vdd.n1256 10.6151
R18697 vdd.n1256 vdd.n1255 10.6151
R18698 vdd.n1255 vdd.n1236 10.6151
R18699 vdd.n1236 vdd.n1235 10.6151
R18700 vdd.n1235 vdd.n1233 10.6151
R18701 vdd.n1233 vdd.n1232 10.6151
R18702 vdd.n1232 vdd.n1230 10.6151
R18703 vdd.n1230 vdd.n1229 10.6151
R18704 vdd.n1229 vdd.n1226 10.6151
R18705 vdd.n1226 vdd.n1225 10.6151
R18706 vdd.n1225 vdd.n831 10.6151
R18707 vdd.n2221 vdd.n967 10.6151
R18708 vdd.n2216 vdd.n967 10.6151
R18709 vdd.n2216 vdd.n2215 10.6151
R18710 vdd.n2215 vdd.n2214 10.6151
R18711 vdd.n2214 vdd.n2211 10.6151
R18712 vdd.n2211 vdd.n2210 10.6151
R18713 vdd.n2210 vdd.n2207 10.6151
R18714 vdd.n2207 vdd.n2206 10.6151
R18715 vdd.n2206 vdd.n2203 10.6151
R18716 vdd.n2203 vdd.n2202 10.6151
R18717 vdd.n2202 vdd.n2199 10.6151
R18718 vdd.n2199 vdd.n2198 10.6151
R18719 vdd.n2198 vdd.n2195 10.6151
R18720 vdd.n2195 vdd.n2194 10.6151
R18721 vdd.n2194 vdd.n2191 10.6151
R18722 vdd.n2191 vdd.n2190 10.6151
R18723 vdd.n2190 vdd.n2187 10.6151
R18724 vdd.n2187 vdd.n1005 10.6151
R18725 vdd.n1151 vdd.n1005 10.6151
R18726 vdd.n1152 vdd.n1151 10.6151
R18727 vdd.n1155 vdd.n1152 10.6151
R18728 vdd.n1156 vdd.n1155 10.6151
R18729 vdd.n1159 vdd.n1156 10.6151
R18730 vdd.n1160 vdd.n1159 10.6151
R18731 vdd.n1163 vdd.n1160 10.6151
R18732 vdd.n1164 vdd.n1163 10.6151
R18733 vdd.n1167 vdd.n1164 10.6151
R18734 vdd.n1168 vdd.n1167 10.6151
R18735 vdd.n1171 vdd.n1168 10.6151
R18736 vdd.n1172 vdd.n1171 10.6151
R18737 vdd.n1175 vdd.n1172 10.6151
R18738 vdd.n1180 vdd.n1177 10.6151
R18739 vdd.n1181 vdd.n1180 10.6151
R18740 vdd.n2732 vdd.n2731 10.6151
R18741 vdd.n2731 vdd.n2730 10.6151
R18742 vdd.n2730 vdd.n2534 10.6151
R18743 vdd.n2612 vdd.n2534 10.6151
R18744 vdd.n2613 vdd.n2612 10.6151
R18745 vdd.n2615 vdd.n2613 10.6151
R18746 vdd.n2616 vdd.n2615 10.6151
R18747 vdd.n2714 vdd.n2616 10.6151
R18748 vdd.n2714 vdd.n2713 10.6151
R18749 vdd.n2713 vdd.n2712 10.6151
R18750 vdd.n2712 vdd.n2660 10.6151
R18751 vdd.n2660 vdd.n2659 10.6151
R18752 vdd.n2659 vdd.n2657 10.6151
R18753 vdd.n2657 vdd.n2656 10.6151
R18754 vdd.n2656 vdd.n2654 10.6151
R18755 vdd.n2654 vdd.n2653 10.6151
R18756 vdd.n2653 vdd.n2651 10.6151
R18757 vdd.n2651 vdd.n2650 10.6151
R18758 vdd.n2650 vdd.n2648 10.6151
R18759 vdd.n2648 vdd.n2647 10.6151
R18760 vdd.n2647 vdd.n2645 10.6151
R18761 vdd.n2645 vdd.n2644 10.6151
R18762 vdd.n2644 vdd.n2642 10.6151
R18763 vdd.n2642 vdd.n2641 10.6151
R18764 vdd.n2641 vdd.n2639 10.6151
R18765 vdd.n2639 vdd.n2638 10.6151
R18766 vdd.n2638 vdd.n2636 10.6151
R18767 vdd.n2636 vdd.n2635 10.6151
R18768 vdd.n2635 vdd.n2633 10.6151
R18769 vdd.n2633 vdd.n2632 10.6151
R18770 vdd.n2632 vdd.n2630 10.6151
R18771 vdd.n2630 vdd.n2629 10.6151
R18772 vdd.n2629 vdd.n2627 10.6151
R18773 vdd.n2627 vdd.n2626 10.6151
R18774 vdd.n2626 vdd.n2624 10.6151
R18775 vdd.n2624 vdd.n2623 10.6151
R18776 vdd.n2623 vdd.n2621 10.6151
R18777 vdd.n2621 vdd.n2620 10.6151
R18778 vdd.n2620 vdd.n2618 10.6151
R18779 vdd.n2618 vdd.n2617 10.6151
R18780 vdd.n2617 vdd.n664 10.6151
R18781 vdd.n2976 vdd.n664 10.6151
R18782 vdd.n2977 vdd.n2976 10.6151
R18783 vdd.n2803 vdd.n789 10.6151
R18784 vdd.n2798 vdd.n789 10.6151
R18785 vdd.n2798 vdd.n2797 10.6151
R18786 vdd.n2797 vdd.n2796 10.6151
R18787 vdd.n2796 vdd.n2793 10.6151
R18788 vdd.n2793 vdd.n2792 10.6151
R18789 vdd.n2792 vdd.n2789 10.6151
R18790 vdd.n2789 vdd.n2788 10.6151
R18791 vdd.n2788 vdd.n2785 10.6151
R18792 vdd.n2785 vdd.n2784 10.6151
R18793 vdd.n2784 vdd.n2781 10.6151
R18794 vdd.n2781 vdd.n2780 10.6151
R18795 vdd.n2780 vdd.n2777 10.6151
R18796 vdd.n2777 vdd.n2776 10.6151
R18797 vdd.n2776 vdd.n2773 10.6151
R18798 vdd.n2773 vdd.n2772 10.6151
R18799 vdd.n2772 vdd.n2769 10.6151
R18800 vdd.n2769 vdd.n2768 10.6151
R18801 vdd.n2768 vdd.n2765 10.6151
R18802 vdd.n2765 vdd.n2764 10.6151
R18803 vdd.n2764 vdd.n2761 10.6151
R18804 vdd.n2761 vdd.n2760 10.6151
R18805 vdd.n2760 vdd.n2757 10.6151
R18806 vdd.n2757 vdd.n2756 10.6151
R18807 vdd.n2756 vdd.n2753 10.6151
R18808 vdd.n2753 vdd.n2752 10.6151
R18809 vdd.n2752 vdd.n2749 10.6151
R18810 vdd.n2749 vdd.n2748 10.6151
R18811 vdd.n2748 vdd.n2745 10.6151
R18812 vdd.n2745 vdd.n2744 10.6151
R18813 vdd.n2744 vdd.n2741 10.6151
R18814 vdd.n2739 vdd.n2736 10.6151
R18815 vdd.n2736 vdd.n2735 10.6151
R18816 vdd.n2805 vdd.n2804 10.6151
R18817 vdd.n2805 vdd.n778 10.6151
R18818 vdd.n2815 vdd.n778 10.6151
R18819 vdd.n2816 vdd.n2815 10.6151
R18820 vdd.n2817 vdd.n2816 10.6151
R18821 vdd.n2817 vdd.n766 10.6151
R18822 vdd.n2827 vdd.n766 10.6151
R18823 vdd.n2828 vdd.n2827 10.6151
R18824 vdd.n2829 vdd.n2828 10.6151
R18825 vdd.n2829 vdd.n755 10.6151
R18826 vdd.n2839 vdd.n755 10.6151
R18827 vdd.n2840 vdd.n2839 10.6151
R18828 vdd.n2841 vdd.n2840 10.6151
R18829 vdd.n2841 vdd.n744 10.6151
R18830 vdd.n2851 vdd.n744 10.6151
R18831 vdd.n2852 vdd.n2851 10.6151
R18832 vdd.n2853 vdd.n2852 10.6151
R18833 vdd.n2853 vdd.n731 10.6151
R18834 vdd.n2864 vdd.n731 10.6151
R18835 vdd.n2865 vdd.n2864 10.6151
R18836 vdd.n2866 vdd.n2865 10.6151
R18837 vdd.n2866 vdd.n719 10.6151
R18838 vdd.n2876 vdd.n719 10.6151
R18839 vdd.n2877 vdd.n2876 10.6151
R18840 vdd.n2878 vdd.n2877 10.6151
R18841 vdd.n2878 vdd.n707 10.6151
R18842 vdd.n2888 vdd.n707 10.6151
R18843 vdd.n2889 vdd.n2888 10.6151
R18844 vdd.n2890 vdd.n2889 10.6151
R18845 vdd.n2890 vdd.n694 10.6151
R18846 vdd.n2900 vdd.n694 10.6151
R18847 vdd.n2901 vdd.n2900 10.6151
R18848 vdd.n2902 vdd.n2901 10.6151
R18849 vdd.n2902 vdd.n683 10.6151
R18850 vdd.n2912 vdd.n683 10.6151
R18851 vdd.n2913 vdd.n2912 10.6151
R18852 vdd.n2914 vdd.n2913 10.6151
R18853 vdd.n2914 vdd.n669 10.6151
R18854 vdd.n2969 vdd.n669 10.6151
R18855 vdd.n2970 vdd.n2969 10.6151
R18856 vdd.n2971 vdd.n2970 10.6151
R18857 vdd.n2971 vdd.n636 10.6151
R18858 vdd.n3041 vdd.n636 10.6151
R18859 vdd.n3040 vdd.n3039 10.6151
R18860 vdd.n3039 vdd.n637 10.6151
R18861 vdd.n638 vdd.n637 10.6151
R18862 vdd.n3032 vdd.n638 10.6151
R18863 vdd.n3032 vdd.n3031 10.6151
R18864 vdd.n3031 vdd.n3030 10.6151
R18865 vdd.n3030 vdd.n640 10.6151
R18866 vdd.n3025 vdd.n640 10.6151
R18867 vdd.n3025 vdd.n3024 10.6151
R18868 vdd.n3024 vdd.n3023 10.6151
R18869 vdd.n3023 vdd.n643 10.6151
R18870 vdd.n3018 vdd.n643 10.6151
R18871 vdd.n3018 vdd.n3017 10.6151
R18872 vdd.n3017 vdd.n3016 10.6151
R18873 vdd.n3016 vdd.n646 10.6151
R18874 vdd.n3011 vdd.n646 10.6151
R18875 vdd.n3011 vdd.n3010 10.6151
R18876 vdd.n3010 vdd.n3008 10.6151
R18877 vdd.n3008 vdd.n649 10.6151
R18878 vdd.n3003 vdd.n649 10.6151
R18879 vdd.n3003 vdd.n3002 10.6151
R18880 vdd.n3002 vdd.n3001 10.6151
R18881 vdd.n3001 vdd.n652 10.6151
R18882 vdd.n2996 vdd.n652 10.6151
R18883 vdd.n2996 vdd.n2995 10.6151
R18884 vdd.n2995 vdd.n2994 10.6151
R18885 vdd.n2994 vdd.n655 10.6151
R18886 vdd.n2989 vdd.n655 10.6151
R18887 vdd.n2989 vdd.n2988 10.6151
R18888 vdd.n2988 vdd.n2987 10.6151
R18889 vdd.n2987 vdd.n658 10.6151
R18890 vdd.n2982 vdd.n2981 10.6151
R18891 vdd.n2981 vdd.n2980 10.6151
R18892 vdd.n2959 vdd.n2920 10.6151
R18893 vdd.n2954 vdd.n2920 10.6151
R18894 vdd.n2954 vdd.n2953 10.6151
R18895 vdd.n2953 vdd.n2952 10.6151
R18896 vdd.n2952 vdd.n2922 10.6151
R18897 vdd.n2947 vdd.n2922 10.6151
R18898 vdd.n2947 vdd.n2946 10.6151
R18899 vdd.n2946 vdd.n2945 10.6151
R18900 vdd.n2945 vdd.n2925 10.6151
R18901 vdd.n2940 vdd.n2925 10.6151
R18902 vdd.n2940 vdd.n2939 10.6151
R18903 vdd.n2939 vdd.n2938 10.6151
R18904 vdd.n2938 vdd.n2928 10.6151
R18905 vdd.n2933 vdd.n2928 10.6151
R18906 vdd.n2933 vdd.n2932 10.6151
R18907 vdd.n2932 vdd.n610 10.6151
R18908 vdd.n3076 vdd.n610 10.6151
R18909 vdd.n3076 vdd.n611 10.6151
R18910 vdd.n614 vdd.n611 10.6151
R18911 vdd.n3069 vdd.n614 10.6151
R18912 vdd.n3069 vdd.n3068 10.6151
R18913 vdd.n3068 vdd.n3067 10.6151
R18914 vdd.n3067 vdd.n616 10.6151
R18915 vdd.n3062 vdd.n616 10.6151
R18916 vdd.n3062 vdd.n3061 10.6151
R18917 vdd.n3061 vdd.n3060 10.6151
R18918 vdd.n3060 vdd.n619 10.6151
R18919 vdd.n3055 vdd.n619 10.6151
R18920 vdd.n3055 vdd.n3054 10.6151
R18921 vdd.n3054 vdd.n3053 10.6151
R18922 vdd.n3053 vdd.n622 10.6151
R18923 vdd.n3048 vdd.n3047 10.6151
R18924 vdd.n3047 vdd.n3046 10.6151
R18925 vdd.n2609 vdd.n2608 10.6151
R18926 vdd.n2726 vdd.n2609 10.6151
R18927 vdd.n2726 vdd.n2725 10.6151
R18928 vdd.n2725 vdd.n2724 10.6151
R18929 vdd.n2724 vdd.n2722 10.6151
R18930 vdd.n2722 vdd.n2721 10.6151
R18931 vdd.n2721 vdd.n2719 10.6151
R18932 vdd.n2719 vdd.n2718 10.6151
R18933 vdd.n2718 vdd.n2610 10.6151
R18934 vdd.n2708 vdd.n2610 10.6151
R18935 vdd.n2708 vdd.n2707 10.6151
R18936 vdd.n2707 vdd.n2706 10.6151
R18937 vdd.n2706 vdd.n2704 10.6151
R18938 vdd.n2704 vdd.n2703 10.6151
R18939 vdd.n2703 vdd.n2701 10.6151
R18940 vdd.n2701 vdd.n2700 10.6151
R18941 vdd.n2700 vdd.n2698 10.6151
R18942 vdd.n2698 vdd.n2697 10.6151
R18943 vdd.n2697 vdd.n2695 10.6151
R18944 vdd.n2695 vdd.n2694 10.6151
R18945 vdd.n2694 vdd.n2692 10.6151
R18946 vdd.n2692 vdd.n2691 10.6151
R18947 vdd.n2691 vdd.n2689 10.6151
R18948 vdd.n2689 vdd.n2688 10.6151
R18949 vdd.n2688 vdd.n2686 10.6151
R18950 vdd.n2686 vdd.n2685 10.6151
R18951 vdd.n2685 vdd.n2683 10.6151
R18952 vdd.n2683 vdd.n2682 10.6151
R18953 vdd.n2682 vdd.n2680 10.6151
R18954 vdd.n2680 vdd.n2679 10.6151
R18955 vdd.n2679 vdd.n2677 10.6151
R18956 vdd.n2677 vdd.n2676 10.6151
R18957 vdd.n2676 vdd.n2674 10.6151
R18958 vdd.n2674 vdd.n2673 10.6151
R18959 vdd.n2673 vdd.n2671 10.6151
R18960 vdd.n2671 vdd.n2670 10.6151
R18961 vdd.n2670 vdd.n2668 10.6151
R18962 vdd.n2668 vdd.n2667 10.6151
R18963 vdd.n2667 vdd.n2665 10.6151
R18964 vdd.n2665 vdd.n2664 10.6151
R18965 vdd.n2664 vdd.n2662 10.6151
R18966 vdd.n2662 vdd.n2661 10.6151
R18967 vdd.n2661 vdd.n628 10.6151
R18968 vdd.n2540 vdd.n2539 10.6151
R18969 vdd.n2543 vdd.n2540 10.6151
R18970 vdd.n2544 vdd.n2543 10.6151
R18971 vdd.n2547 vdd.n2544 10.6151
R18972 vdd.n2548 vdd.n2547 10.6151
R18973 vdd.n2551 vdd.n2548 10.6151
R18974 vdd.n2552 vdd.n2551 10.6151
R18975 vdd.n2555 vdd.n2552 10.6151
R18976 vdd.n2556 vdd.n2555 10.6151
R18977 vdd.n2559 vdd.n2556 10.6151
R18978 vdd.n2560 vdd.n2559 10.6151
R18979 vdd.n2563 vdd.n2560 10.6151
R18980 vdd.n2564 vdd.n2563 10.6151
R18981 vdd.n2567 vdd.n2564 10.6151
R18982 vdd.n2568 vdd.n2567 10.6151
R18983 vdd.n2571 vdd.n2568 10.6151
R18984 vdd.n2572 vdd.n2571 10.6151
R18985 vdd.n2575 vdd.n2572 10.6151
R18986 vdd.n2576 vdd.n2575 10.6151
R18987 vdd.n2579 vdd.n2576 10.6151
R18988 vdd.n2580 vdd.n2579 10.6151
R18989 vdd.n2583 vdd.n2580 10.6151
R18990 vdd.n2584 vdd.n2583 10.6151
R18991 vdd.n2587 vdd.n2584 10.6151
R18992 vdd.n2588 vdd.n2587 10.6151
R18993 vdd.n2591 vdd.n2588 10.6151
R18994 vdd.n2592 vdd.n2591 10.6151
R18995 vdd.n2595 vdd.n2592 10.6151
R18996 vdd.n2596 vdd.n2595 10.6151
R18997 vdd.n2599 vdd.n2596 10.6151
R18998 vdd.n2600 vdd.n2599 10.6151
R18999 vdd.n2605 vdd.n2603 10.6151
R19000 vdd.n2606 vdd.n2605 10.6151
R19001 vdd.n2809 vdd.n783 10.6151
R19002 vdd.n2810 vdd.n2809 10.6151
R19003 vdd.n2811 vdd.n2810 10.6151
R19004 vdd.n2811 vdd.n772 10.6151
R19005 vdd.n2821 vdd.n772 10.6151
R19006 vdd.n2822 vdd.n2821 10.6151
R19007 vdd.n2823 vdd.n2822 10.6151
R19008 vdd.n2823 vdd.n761 10.6151
R19009 vdd.n2833 vdd.n761 10.6151
R19010 vdd.n2834 vdd.n2833 10.6151
R19011 vdd.n2835 vdd.n2834 10.6151
R19012 vdd.n2835 vdd.n749 10.6151
R19013 vdd.n2845 vdd.n749 10.6151
R19014 vdd.n2846 vdd.n2845 10.6151
R19015 vdd.n2847 vdd.n2846 10.6151
R19016 vdd.n2847 vdd.n738 10.6151
R19017 vdd.n2857 vdd.n738 10.6151
R19018 vdd.n2858 vdd.n2857 10.6151
R19019 vdd.n2860 vdd.n2858 10.6151
R19020 vdd.n2860 vdd.n2859 10.6151
R19021 vdd.n2871 vdd.n2870 10.6151
R19022 vdd.n2872 vdd.n2871 10.6151
R19023 vdd.n2872 vdd.n713 10.6151
R19024 vdd.n2882 vdd.n713 10.6151
R19025 vdd.n2883 vdd.n2882 10.6151
R19026 vdd.n2884 vdd.n2883 10.6151
R19027 vdd.n2884 vdd.n700 10.6151
R19028 vdd.n2894 vdd.n700 10.6151
R19029 vdd.n2895 vdd.n2894 10.6151
R19030 vdd.n2896 vdd.n2895 10.6151
R19031 vdd.n2896 vdd.n688 10.6151
R19032 vdd.n2906 vdd.n688 10.6151
R19033 vdd.n2907 vdd.n2906 10.6151
R19034 vdd.n2908 vdd.n2907 10.6151
R19035 vdd.n2908 vdd.n677 10.6151
R19036 vdd.n2918 vdd.n677 10.6151
R19037 vdd.n2919 vdd.n2918 10.6151
R19038 vdd.n2965 vdd.n2919 10.6151
R19039 vdd.n2965 vdd.n2964 10.6151
R19040 vdd.n2964 vdd.n2963 10.6151
R19041 vdd.n2963 vdd.n2962 10.6151
R19042 vdd.n2962 vdd.n2960 10.6151
R19043 vdd.n2227 vdd.n960 10.6151
R19044 vdd.n2228 vdd.n2227 10.6151
R19045 vdd.n2229 vdd.n2228 10.6151
R19046 vdd.n2229 vdd.n949 10.6151
R19047 vdd.n2239 vdd.n949 10.6151
R19048 vdd.n2240 vdd.n2239 10.6151
R19049 vdd.n2241 vdd.n2240 10.6151
R19050 vdd.n2241 vdd.n936 10.6151
R19051 vdd.n2251 vdd.n936 10.6151
R19052 vdd.n2252 vdd.n2251 10.6151
R19053 vdd.n2253 vdd.n2252 10.6151
R19054 vdd.n2253 vdd.n925 10.6151
R19055 vdd.n2263 vdd.n925 10.6151
R19056 vdd.n2264 vdd.n2263 10.6151
R19057 vdd.n2265 vdd.n2264 10.6151
R19058 vdd.n2265 vdd.n913 10.6151
R19059 vdd.n2275 vdd.n913 10.6151
R19060 vdd.n2276 vdd.n2275 10.6151
R19061 vdd.n2277 vdd.n2276 10.6151
R19062 vdd.n2277 vdd.n900 10.6151
R19063 vdd.n2287 vdd.n900 10.6151
R19064 vdd.n2288 vdd.n2287 10.6151
R19065 vdd.n2290 vdd.n888 10.6151
R19066 vdd.n2300 vdd.n888 10.6151
R19067 vdd.n2301 vdd.n2300 10.6151
R19068 vdd.n2302 vdd.n2301 10.6151
R19069 vdd.n2302 vdd.n876 10.6151
R19070 vdd.n2312 vdd.n876 10.6151
R19071 vdd.n2313 vdd.n2312 10.6151
R19072 vdd.n2314 vdd.n2313 10.6151
R19073 vdd.n2314 vdd.n865 10.6151
R19074 vdd.n2324 vdd.n865 10.6151
R19075 vdd.n2325 vdd.n2324 10.6151
R19076 vdd.n2326 vdd.n2325 10.6151
R19077 vdd.n2326 vdd.n854 10.6151
R19078 vdd.n2336 vdd.n854 10.6151
R19079 vdd.n2337 vdd.n2336 10.6151
R19080 vdd.n2340 vdd.n2337 10.6151
R19081 vdd.n2340 vdd.n2339 10.6151
R19082 vdd.n2339 vdd.n2338 10.6151
R19083 vdd.n2338 vdd.n837 10.6151
R19084 vdd.n2422 vdd.n837 10.6151
R19085 vdd.n2421 vdd.n2420 10.6151
R19086 vdd.n2420 vdd.n2417 10.6151
R19087 vdd.n2417 vdd.n2416 10.6151
R19088 vdd.n2416 vdd.n2413 10.6151
R19089 vdd.n2413 vdd.n2412 10.6151
R19090 vdd.n2412 vdd.n2409 10.6151
R19091 vdd.n2409 vdd.n2408 10.6151
R19092 vdd.n2408 vdd.n2405 10.6151
R19093 vdd.n2405 vdd.n2404 10.6151
R19094 vdd.n2404 vdd.n2401 10.6151
R19095 vdd.n2401 vdd.n2400 10.6151
R19096 vdd.n2400 vdd.n2397 10.6151
R19097 vdd.n2397 vdd.n2396 10.6151
R19098 vdd.n2396 vdd.n2393 10.6151
R19099 vdd.n2393 vdd.n2392 10.6151
R19100 vdd.n2392 vdd.n2389 10.6151
R19101 vdd.n2389 vdd.n2388 10.6151
R19102 vdd.n2388 vdd.n2385 10.6151
R19103 vdd.n2385 vdd.n2384 10.6151
R19104 vdd.n2384 vdd.n2381 10.6151
R19105 vdd.n2381 vdd.n2380 10.6151
R19106 vdd.n2380 vdd.n2377 10.6151
R19107 vdd.n2377 vdd.n2376 10.6151
R19108 vdd.n2376 vdd.n2373 10.6151
R19109 vdd.n2373 vdd.n2372 10.6151
R19110 vdd.n2372 vdd.n2369 10.6151
R19111 vdd.n2369 vdd.n2368 10.6151
R19112 vdd.n2368 vdd.n2365 10.6151
R19113 vdd.n2365 vdd.n2364 10.6151
R19114 vdd.n2364 vdd.n2361 10.6151
R19115 vdd.n2361 vdd.n2360 10.6151
R19116 vdd.n2357 vdd.n2356 10.6151
R19117 vdd.n2356 vdd.n2354 10.6151
R19118 vdd.n1309 vdd.n1307 10.6151
R19119 vdd.n1307 vdd.n1306 10.6151
R19120 vdd.n1306 vdd.n1304 10.6151
R19121 vdd.n1304 vdd.n1303 10.6151
R19122 vdd.n1303 vdd.n1301 10.6151
R19123 vdd.n1301 vdd.n1300 10.6151
R19124 vdd.n1300 vdd.n1298 10.6151
R19125 vdd.n1298 vdd.n1297 10.6151
R19126 vdd.n1297 vdd.n1295 10.6151
R19127 vdd.n1295 vdd.n1294 10.6151
R19128 vdd.n1294 vdd.n1292 10.6151
R19129 vdd.n1292 vdd.n1291 10.6151
R19130 vdd.n1291 vdd.n1289 10.6151
R19131 vdd.n1289 vdd.n1288 10.6151
R19132 vdd.n1288 vdd.n1286 10.6151
R19133 vdd.n1286 vdd.n1285 10.6151
R19134 vdd.n1285 vdd.n1283 10.6151
R19135 vdd.n1283 vdd.n1282 10.6151
R19136 vdd.n1282 vdd.n1280 10.6151
R19137 vdd.n1280 vdd.n1279 10.6151
R19138 vdd.n1279 vdd.n1277 10.6151
R19139 vdd.n1277 vdd.n1276 10.6151
R19140 vdd.n1276 vdd.n1274 10.6151
R19141 vdd.n1274 vdd.n1273 10.6151
R19142 vdd.n1273 vdd.n1271 10.6151
R19143 vdd.n1271 vdd.n1270 10.6151
R19144 vdd.n1270 vdd.n1268 10.6151
R19145 vdd.n1268 vdd.n1267 10.6151
R19146 vdd.n1267 vdd.n1146 10.6151
R19147 vdd.n1238 vdd.n1146 10.6151
R19148 vdd.n1239 vdd.n1238 10.6151
R19149 vdd.n1241 vdd.n1239 10.6151
R19150 vdd.n1242 vdd.n1241 10.6151
R19151 vdd.n1251 vdd.n1242 10.6151
R19152 vdd.n1251 vdd.n1250 10.6151
R19153 vdd.n1250 vdd.n1249 10.6151
R19154 vdd.n1249 vdd.n1247 10.6151
R19155 vdd.n1247 vdd.n1246 10.6151
R19156 vdd.n1246 vdd.n1244 10.6151
R19157 vdd.n1244 vdd.n1243 10.6151
R19158 vdd.n1243 vdd.n841 10.6151
R19159 vdd.n2352 vdd.n841 10.6151
R19160 vdd.n2353 vdd.n2352 10.6151
R19161 vdd.n1110 vdd.n1109 10.6151
R19162 vdd.n1113 vdd.n1110 10.6151
R19163 vdd.n1114 vdd.n1113 10.6151
R19164 vdd.n1117 vdd.n1114 10.6151
R19165 vdd.n1118 vdd.n1117 10.6151
R19166 vdd.n1121 vdd.n1118 10.6151
R19167 vdd.n1122 vdd.n1121 10.6151
R19168 vdd.n1125 vdd.n1122 10.6151
R19169 vdd.n1126 vdd.n1125 10.6151
R19170 vdd.n1129 vdd.n1126 10.6151
R19171 vdd.n1130 vdd.n1129 10.6151
R19172 vdd.n1133 vdd.n1130 10.6151
R19173 vdd.n1134 vdd.n1133 10.6151
R19174 vdd.n1137 vdd.n1134 10.6151
R19175 vdd.n1138 vdd.n1137 10.6151
R19176 vdd.n1141 vdd.n1138 10.6151
R19177 vdd.n1343 vdd.n1141 10.6151
R19178 vdd.n1343 vdd.n1342 10.6151
R19179 vdd.n1342 vdd.n1340 10.6151
R19180 vdd.n1340 vdd.n1337 10.6151
R19181 vdd.n1337 vdd.n1336 10.6151
R19182 vdd.n1336 vdd.n1333 10.6151
R19183 vdd.n1333 vdd.n1332 10.6151
R19184 vdd.n1332 vdd.n1329 10.6151
R19185 vdd.n1329 vdd.n1328 10.6151
R19186 vdd.n1328 vdd.n1325 10.6151
R19187 vdd.n1325 vdd.n1324 10.6151
R19188 vdd.n1324 vdd.n1321 10.6151
R19189 vdd.n1321 vdd.n1320 10.6151
R19190 vdd.n1320 vdd.n1317 10.6151
R19191 vdd.n1317 vdd.n1316 10.6151
R19192 vdd.n1313 vdd.n1312 10.6151
R19193 vdd.n1312 vdd.n1310 10.6151
R19194 vdd.n1727 vdd.t90 10.5435
R19195 vdd.n2070 vdd.t19 10.5435
R19196 vdd.n3212 vdd.t29 10.5435
R19197 vdd.n3436 vdd.t101 10.5435
R19198 vdd.n292 vdd.n274 10.4732
R19199 vdd.n241 vdd.n223 10.4732
R19200 vdd.n198 vdd.n180 10.4732
R19201 vdd.n147 vdd.n129 10.4732
R19202 vdd.n105 vdd.n87 10.4732
R19203 vdd.n54 vdd.n36 10.4732
R19204 vdd.n1942 vdd.n1924 10.4732
R19205 vdd.n1993 vdd.n1975 10.4732
R19206 vdd.n1848 vdd.n1830 10.4732
R19207 vdd.n1899 vdd.n1881 10.4732
R19208 vdd.n1755 vdd.n1737 10.4732
R19209 vdd.n1806 vdd.n1788 10.4732
R19210 vdd.n2025 vdd.t119 10.3167
R19211 vdd.t121 vdd.n493 10.3167
R19212 vdd.n2187 vdd.n2186 9.98956
R19213 vdd.n3010 vdd.n3009 9.98956
R19214 vdd.n3077 vdd.n3076 9.98956
R19215 vdd.n2079 vdd.n1343 9.98956
R19216 vdd.n1678 vdd.t47 9.86327
R19217 vdd.n3412 vdd.t33 9.86327
R19218 vdd.n2424 vdd.t220 9.7499
R19219 vdd.t205 vdd.n785 9.7499
R19220 vdd.n291 vdd.n276 9.69747
R19221 vdd.n240 vdd.n225 9.69747
R19222 vdd.n197 vdd.n182 9.69747
R19223 vdd.n146 vdd.n131 9.69747
R19224 vdd.n104 vdd.n89 9.69747
R19225 vdd.n53 vdd.n38 9.69747
R19226 vdd.n1941 vdd.n1926 9.69747
R19227 vdd.n1992 vdd.n1977 9.69747
R19228 vdd.n1847 vdd.n1832 9.69747
R19229 vdd.n1898 vdd.n1883 9.69747
R19230 vdd.n1754 vdd.n1739 9.69747
R19231 vdd.n1805 vdd.n1790 9.69747
R19232 vdd.n307 vdd.n306 9.45567
R19233 vdd.n256 vdd.n255 9.45567
R19234 vdd.n213 vdd.n212 9.45567
R19235 vdd.n162 vdd.n161 9.45567
R19236 vdd.n120 vdd.n119 9.45567
R19237 vdd.n69 vdd.n68 9.45567
R19238 vdd.n1957 vdd.n1956 9.45567
R19239 vdd.n2008 vdd.n2007 9.45567
R19240 vdd.n1863 vdd.n1862 9.45567
R19241 vdd.n1914 vdd.n1913 9.45567
R19242 vdd.n1770 vdd.n1769 9.45567
R19243 vdd.n1821 vdd.n1820 9.45567
R19244 vdd.n2149 vdd.n1035 9.3005
R19245 vdd.n2148 vdd.n2147 9.3005
R19246 vdd.n1041 vdd.n1040 9.3005
R19247 vdd.n2142 vdd.n1045 9.3005
R19248 vdd.n2141 vdd.n1046 9.3005
R19249 vdd.n2140 vdd.n1047 9.3005
R19250 vdd.n1051 vdd.n1048 9.3005
R19251 vdd.n2135 vdd.n1052 9.3005
R19252 vdd.n2134 vdd.n1053 9.3005
R19253 vdd.n2133 vdd.n1054 9.3005
R19254 vdd.n1058 vdd.n1055 9.3005
R19255 vdd.n2128 vdd.n1059 9.3005
R19256 vdd.n2127 vdd.n1060 9.3005
R19257 vdd.n2126 vdd.n1061 9.3005
R19258 vdd.n1065 vdd.n1062 9.3005
R19259 vdd.n2121 vdd.n1066 9.3005
R19260 vdd.n2120 vdd.n1067 9.3005
R19261 vdd.n2119 vdd.n1068 9.3005
R19262 vdd.n1072 vdd.n1069 9.3005
R19263 vdd.n2114 vdd.n1073 9.3005
R19264 vdd.n2113 vdd.n1074 9.3005
R19265 vdd.n2112 vdd.n2111 9.3005
R19266 vdd.n2110 vdd.n1075 9.3005
R19267 vdd.n2109 vdd.n2108 9.3005
R19268 vdd.n1081 vdd.n1080 9.3005
R19269 vdd.n2103 vdd.n1085 9.3005
R19270 vdd.n2102 vdd.n1086 9.3005
R19271 vdd.n2101 vdd.n1087 9.3005
R19272 vdd.n1091 vdd.n1088 9.3005
R19273 vdd.n2096 vdd.n1092 9.3005
R19274 vdd.n2095 vdd.n1093 9.3005
R19275 vdd.n2094 vdd.n1094 9.3005
R19276 vdd.n1098 vdd.n1095 9.3005
R19277 vdd.n2089 vdd.n1099 9.3005
R19278 vdd.n2088 vdd.n1100 9.3005
R19279 vdd.n2087 vdd.n1101 9.3005
R19280 vdd.n1105 vdd.n1102 9.3005
R19281 vdd.n2082 vdd.n1106 9.3005
R19282 vdd.n2151 vdd.n2150 9.3005
R19283 vdd.n2173 vdd.n1006 9.3005
R19284 vdd.n2172 vdd.n1014 9.3005
R19285 vdd.n1018 vdd.n1015 9.3005
R19286 vdd.n2167 vdd.n1019 9.3005
R19287 vdd.n2166 vdd.n1020 9.3005
R19288 vdd.n2165 vdd.n1021 9.3005
R19289 vdd.n1025 vdd.n1022 9.3005
R19290 vdd.n2160 vdd.n1026 9.3005
R19291 vdd.n2159 vdd.n1027 9.3005
R19292 vdd.n2158 vdd.n1028 9.3005
R19293 vdd.n1032 vdd.n1029 9.3005
R19294 vdd.n2153 vdd.n1033 9.3005
R19295 vdd.n2152 vdd.n1034 9.3005
R19296 vdd.n2185 vdd.n2184 9.3005
R19297 vdd.n1010 vdd.n1009 9.3005
R19298 vdd.n2013 vdd.n1394 9.3005
R19299 vdd.n2015 vdd.n2014 9.3005
R19300 vdd.n1384 vdd.n1383 9.3005
R19301 vdd.n2029 vdd.n2028 9.3005
R19302 vdd.n2030 vdd.n1382 9.3005
R19303 vdd.n2032 vdd.n2031 9.3005
R19304 vdd.n1373 vdd.n1372 9.3005
R19305 vdd.n2046 vdd.n2045 9.3005
R19306 vdd.n2047 vdd.n1371 9.3005
R19307 vdd.n2049 vdd.n2048 9.3005
R19308 vdd.n1361 vdd.n1360 9.3005
R19309 vdd.n2065 vdd.n2064 9.3005
R19310 vdd.n2066 vdd.n1359 9.3005
R19311 vdd.n2068 vdd.n2067 9.3005
R19312 vdd.n283 vdd.n282 9.3005
R19313 vdd.n278 vdd.n277 9.3005
R19314 vdd.n289 vdd.n288 9.3005
R19315 vdd.n291 vdd.n290 9.3005
R19316 vdd.n274 vdd.n273 9.3005
R19317 vdd.n297 vdd.n296 9.3005
R19318 vdd.n299 vdd.n298 9.3005
R19319 vdd.n271 vdd.n268 9.3005
R19320 vdd.n306 vdd.n305 9.3005
R19321 vdd.n232 vdd.n231 9.3005
R19322 vdd.n227 vdd.n226 9.3005
R19323 vdd.n238 vdd.n237 9.3005
R19324 vdd.n240 vdd.n239 9.3005
R19325 vdd.n223 vdd.n222 9.3005
R19326 vdd.n246 vdd.n245 9.3005
R19327 vdd.n248 vdd.n247 9.3005
R19328 vdd.n220 vdd.n217 9.3005
R19329 vdd.n255 vdd.n254 9.3005
R19330 vdd.n189 vdd.n188 9.3005
R19331 vdd.n184 vdd.n183 9.3005
R19332 vdd.n195 vdd.n194 9.3005
R19333 vdd.n197 vdd.n196 9.3005
R19334 vdd.n180 vdd.n179 9.3005
R19335 vdd.n203 vdd.n202 9.3005
R19336 vdd.n205 vdd.n204 9.3005
R19337 vdd.n177 vdd.n174 9.3005
R19338 vdd.n212 vdd.n211 9.3005
R19339 vdd.n138 vdd.n137 9.3005
R19340 vdd.n133 vdd.n132 9.3005
R19341 vdd.n144 vdd.n143 9.3005
R19342 vdd.n146 vdd.n145 9.3005
R19343 vdd.n129 vdd.n128 9.3005
R19344 vdd.n152 vdd.n151 9.3005
R19345 vdd.n154 vdd.n153 9.3005
R19346 vdd.n126 vdd.n123 9.3005
R19347 vdd.n161 vdd.n160 9.3005
R19348 vdd.n96 vdd.n95 9.3005
R19349 vdd.n91 vdd.n90 9.3005
R19350 vdd.n102 vdd.n101 9.3005
R19351 vdd.n104 vdd.n103 9.3005
R19352 vdd.n87 vdd.n86 9.3005
R19353 vdd.n110 vdd.n109 9.3005
R19354 vdd.n112 vdd.n111 9.3005
R19355 vdd.n84 vdd.n81 9.3005
R19356 vdd.n119 vdd.n118 9.3005
R19357 vdd.n45 vdd.n44 9.3005
R19358 vdd.n40 vdd.n39 9.3005
R19359 vdd.n51 vdd.n50 9.3005
R19360 vdd.n53 vdd.n52 9.3005
R19361 vdd.n36 vdd.n35 9.3005
R19362 vdd.n59 vdd.n58 9.3005
R19363 vdd.n61 vdd.n60 9.3005
R19364 vdd.n33 vdd.n30 9.3005
R19365 vdd.n68 vdd.n67 9.3005
R19366 vdd.n3126 vdd.n3125 9.3005
R19367 vdd.n3127 vdd.n578 9.3005
R19368 vdd.n577 vdd.n575 9.3005
R19369 vdd.n3133 vdd.n574 9.3005
R19370 vdd.n3134 vdd.n573 9.3005
R19371 vdd.n3135 vdd.n572 9.3005
R19372 vdd.n571 vdd.n569 9.3005
R19373 vdd.n3141 vdd.n568 9.3005
R19374 vdd.n3142 vdd.n567 9.3005
R19375 vdd.n3143 vdd.n566 9.3005
R19376 vdd.n565 vdd.n563 9.3005
R19377 vdd.n3149 vdd.n562 9.3005
R19378 vdd.n3150 vdd.n561 9.3005
R19379 vdd.n3151 vdd.n560 9.3005
R19380 vdd.n559 vdd.n557 9.3005
R19381 vdd.n3157 vdd.n556 9.3005
R19382 vdd.n3158 vdd.n555 9.3005
R19383 vdd.n3159 vdd.n554 9.3005
R19384 vdd.n553 vdd.n551 9.3005
R19385 vdd.n3165 vdd.n550 9.3005
R19386 vdd.n3166 vdd.n549 9.3005
R19387 vdd.n3167 vdd.n548 9.3005
R19388 vdd.n547 vdd.n545 9.3005
R19389 vdd.n3173 vdd.n542 9.3005
R19390 vdd.n3174 vdd.n541 9.3005
R19391 vdd.n3175 vdd.n540 9.3005
R19392 vdd.n539 vdd.n537 9.3005
R19393 vdd.n3181 vdd.n536 9.3005
R19394 vdd.n3182 vdd.n535 9.3005
R19395 vdd.n3183 vdd.n534 9.3005
R19396 vdd.n533 vdd.n531 9.3005
R19397 vdd.n3189 vdd.n530 9.3005
R19398 vdd.n3190 vdd.n529 9.3005
R19399 vdd.n3191 vdd.n528 9.3005
R19400 vdd.n527 vdd.n525 9.3005
R19401 vdd.n3196 vdd.n524 9.3005
R19402 vdd.n3206 vdd.n518 9.3005
R19403 vdd.n3208 vdd.n3207 9.3005
R19404 vdd.n509 vdd.n508 9.3005
R19405 vdd.n3223 vdd.n3222 9.3005
R19406 vdd.n3224 vdd.n507 9.3005
R19407 vdd.n3226 vdd.n3225 9.3005
R19408 vdd.n497 vdd.n496 9.3005
R19409 vdd.n3239 vdd.n3238 9.3005
R19410 vdd.n3240 vdd.n495 9.3005
R19411 vdd.n3242 vdd.n3241 9.3005
R19412 vdd.n485 vdd.n484 9.3005
R19413 vdd.n3256 vdd.n3255 9.3005
R19414 vdd.n3257 vdd.n483 9.3005
R19415 vdd.n3259 vdd.n3258 9.3005
R19416 vdd.n312 vdd.n310 9.3005
R19417 vdd.n3210 vdd.n3209 9.3005
R19418 vdd.n3439 vdd.n3438 9.3005
R19419 vdd.n313 vdd.n311 9.3005
R19420 vdd.n3432 vdd.n320 9.3005
R19421 vdd.n3431 vdd.n321 9.3005
R19422 vdd.n3430 vdd.n322 9.3005
R19423 vdd.n331 vdd.n323 9.3005
R19424 vdd.n3424 vdd.n332 9.3005
R19425 vdd.n3423 vdd.n333 9.3005
R19426 vdd.n3422 vdd.n334 9.3005
R19427 vdd.n342 vdd.n335 9.3005
R19428 vdd.n3416 vdd.n343 9.3005
R19429 vdd.n3415 vdd.n344 9.3005
R19430 vdd.n3414 vdd.n345 9.3005
R19431 vdd.n353 vdd.n346 9.3005
R19432 vdd.n3408 vdd.n3407 9.3005
R19433 vdd.n3404 vdd.n354 9.3005
R19434 vdd.n3403 vdd.n357 9.3005
R19435 vdd.n361 vdd.n358 9.3005
R19436 vdd.n362 vdd.n359 9.3005
R19437 vdd.n3396 vdd.n363 9.3005
R19438 vdd.n3395 vdd.n364 9.3005
R19439 vdd.n3394 vdd.n365 9.3005
R19440 vdd.n369 vdd.n366 9.3005
R19441 vdd.n3389 vdd.n370 9.3005
R19442 vdd.n3388 vdd.n371 9.3005
R19443 vdd.n3387 vdd.n372 9.3005
R19444 vdd.n376 vdd.n373 9.3005
R19445 vdd.n3382 vdd.n377 9.3005
R19446 vdd.n3381 vdd.n378 9.3005
R19447 vdd.n3380 vdd.n379 9.3005
R19448 vdd.n383 vdd.n380 9.3005
R19449 vdd.n3375 vdd.n384 9.3005
R19450 vdd.n3374 vdd.n385 9.3005
R19451 vdd.n3373 vdd.n3372 9.3005
R19452 vdd.n3371 vdd.n386 9.3005
R19453 vdd.n3370 vdd.n3369 9.3005
R19454 vdd.n392 vdd.n391 9.3005
R19455 vdd.n3364 vdd.n396 9.3005
R19456 vdd.n3363 vdd.n397 9.3005
R19457 vdd.n3362 vdd.n398 9.3005
R19458 vdd.n402 vdd.n399 9.3005
R19459 vdd.n3357 vdd.n403 9.3005
R19460 vdd.n3356 vdd.n404 9.3005
R19461 vdd.n3355 vdd.n405 9.3005
R19462 vdd.n409 vdd.n406 9.3005
R19463 vdd.n3350 vdd.n410 9.3005
R19464 vdd.n3349 vdd.n411 9.3005
R19465 vdd.n3348 vdd.n412 9.3005
R19466 vdd.n416 vdd.n413 9.3005
R19467 vdd.n3343 vdd.n417 9.3005
R19468 vdd.n3342 vdd.n418 9.3005
R19469 vdd.n3341 vdd.n419 9.3005
R19470 vdd.n423 vdd.n420 9.3005
R19471 vdd.n3336 vdd.n424 9.3005
R19472 vdd.n3335 vdd.n425 9.3005
R19473 vdd.n3334 vdd.n3333 9.3005
R19474 vdd.n3332 vdd.n426 9.3005
R19475 vdd.n3331 vdd.n3330 9.3005
R19476 vdd.n432 vdd.n431 9.3005
R19477 vdd.n3325 vdd.n436 9.3005
R19478 vdd.n3324 vdd.n437 9.3005
R19479 vdd.n3323 vdd.n438 9.3005
R19480 vdd.n442 vdd.n439 9.3005
R19481 vdd.n3318 vdd.n443 9.3005
R19482 vdd.n3317 vdd.n444 9.3005
R19483 vdd.n3316 vdd.n445 9.3005
R19484 vdd.n449 vdd.n446 9.3005
R19485 vdd.n3311 vdd.n450 9.3005
R19486 vdd.n3310 vdd.n451 9.3005
R19487 vdd.n3309 vdd.n452 9.3005
R19488 vdd.n456 vdd.n453 9.3005
R19489 vdd.n3304 vdd.n457 9.3005
R19490 vdd.n3303 vdd.n458 9.3005
R19491 vdd.n3302 vdd.n459 9.3005
R19492 vdd.n463 vdd.n460 9.3005
R19493 vdd.n3297 vdd.n464 9.3005
R19494 vdd.n3296 vdd.n465 9.3005
R19495 vdd.n3292 vdd.n3289 9.3005
R19496 vdd.n3406 vdd.n3405 9.3005
R19497 vdd.n3216 vdd.n513 9.3005
R19498 vdd.n3218 vdd.n3217 9.3005
R19499 vdd.n503 vdd.n502 9.3005
R19500 vdd.n3231 vdd.n3230 9.3005
R19501 vdd.n3232 vdd.n501 9.3005
R19502 vdd.n3234 vdd.n3233 9.3005
R19503 vdd.n490 vdd.n489 9.3005
R19504 vdd.n3247 vdd.n3246 9.3005
R19505 vdd.n3248 vdd.n488 9.3005
R19506 vdd.n3250 vdd.n3249 9.3005
R19507 vdd.n478 vdd.n477 9.3005
R19508 vdd.n3264 vdd.n3263 9.3005
R19509 vdd.n3265 vdd.n476 9.3005
R19510 vdd.n3267 vdd.n3266 9.3005
R19511 vdd.n3268 vdd.n475 9.3005
R19512 vdd.n3270 vdd.n3269 9.3005
R19513 vdd.n3271 vdd.n474 9.3005
R19514 vdd.n3273 vdd.n3272 9.3005
R19515 vdd.n3274 vdd.n472 9.3005
R19516 vdd.n3276 vdd.n3275 9.3005
R19517 vdd.n3277 vdd.n471 9.3005
R19518 vdd.n3279 vdd.n3278 9.3005
R19519 vdd.n3280 vdd.n469 9.3005
R19520 vdd.n3282 vdd.n3281 9.3005
R19521 vdd.n3283 vdd.n468 9.3005
R19522 vdd.n3285 vdd.n3284 9.3005
R19523 vdd.n3286 vdd.n466 9.3005
R19524 vdd.n3288 vdd.n3287 9.3005
R19525 vdd.n3215 vdd.n3214 9.3005
R19526 vdd.n3079 vdd.n514 9.3005
R19527 vdd.n3084 vdd.n3078 9.3005
R19528 vdd.n3094 vdd.n605 9.3005
R19529 vdd.n3095 vdd.n604 9.3005
R19530 vdd.n603 vdd.n601 9.3005
R19531 vdd.n3101 vdd.n600 9.3005
R19532 vdd.n3102 vdd.n599 9.3005
R19533 vdd.n3103 vdd.n598 9.3005
R19534 vdd.n597 vdd.n595 9.3005
R19535 vdd.n3109 vdd.n594 9.3005
R19536 vdd.n3110 vdd.n593 9.3005
R19537 vdd.n3111 vdd.n592 9.3005
R19538 vdd.n591 vdd.n589 9.3005
R19539 vdd.n3116 vdd.n588 9.3005
R19540 vdd.n3117 vdd.n587 9.3005
R19541 vdd.n583 vdd.n582 9.3005
R19542 vdd.n3123 vdd.n3122 9.3005
R19543 vdd.n3124 vdd.n579 9.3005
R19544 vdd.n2078 vdd.n2077 9.3005
R19545 vdd.n2073 vdd.n1345 9.3005
R19546 vdd.n1674 vdd.n1434 9.3005
R19547 vdd.n1676 vdd.n1675 9.3005
R19548 vdd.n1425 vdd.n1424 9.3005
R19549 vdd.n1689 vdd.n1688 9.3005
R19550 vdd.n1690 vdd.n1423 9.3005
R19551 vdd.n1692 vdd.n1691 9.3005
R19552 vdd.n1412 vdd.n1411 9.3005
R19553 vdd.n1705 vdd.n1704 9.3005
R19554 vdd.n1706 vdd.n1410 9.3005
R19555 vdd.n1708 vdd.n1707 9.3005
R19556 vdd.n1401 vdd.n1400 9.3005
R19557 vdd.n1722 vdd.n1721 9.3005
R19558 vdd.n1723 vdd.n1399 9.3005
R19559 vdd.n1725 vdd.n1724 9.3005
R19560 vdd.n1390 vdd.n1389 9.3005
R19561 vdd.n2020 vdd.n2019 9.3005
R19562 vdd.n2021 vdd.n1388 9.3005
R19563 vdd.n2023 vdd.n2022 9.3005
R19564 vdd.n1378 vdd.n1377 9.3005
R19565 vdd.n2037 vdd.n2036 9.3005
R19566 vdd.n2038 vdd.n1376 9.3005
R19567 vdd.n2040 vdd.n2039 9.3005
R19568 vdd.n1368 vdd.n1367 9.3005
R19569 vdd.n2054 vdd.n2053 9.3005
R19570 vdd.n2055 vdd.n1365 9.3005
R19571 vdd.n2059 vdd.n2058 9.3005
R19572 vdd.n2057 vdd.n1366 9.3005
R19573 vdd.n2056 vdd.n1356 9.3005
R19574 vdd.n1673 vdd.n1672 9.3005
R19575 vdd.n1568 vdd.n1558 9.3005
R19576 vdd.n1570 vdd.n1569 9.3005
R19577 vdd.n1571 vdd.n1557 9.3005
R19578 vdd.n1573 vdd.n1572 9.3005
R19579 vdd.n1574 vdd.n1550 9.3005
R19580 vdd.n1576 vdd.n1575 9.3005
R19581 vdd.n1577 vdd.n1549 9.3005
R19582 vdd.n1579 vdd.n1578 9.3005
R19583 vdd.n1580 vdd.n1542 9.3005
R19584 vdd.n1582 vdd.n1581 9.3005
R19585 vdd.n1583 vdd.n1541 9.3005
R19586 vdd.n1585 vdd.n1584 9.3005
R19587 vdd.n1586 vdd.n1534 9.3005
R19588 vdd.n1588 vdd.n1587 9.3005
R19589 vdd.n1589 vdd.n1533 9.3005
R19590 vdd.n1591 vdd.n1590 9.3005
R19591 vdd.n1592 vdd.n1527 9.3005
R19592 vdd.n1594 vdd.n1593 9.3005
R19593 vdd.n1595 vdd.n1525 9.3005
R19594 vdd.n1597 vdd.n1596 9.3005
R19595 vdd.n1526 vdd.n1523 9.3005
R19596 vdd.n1604 vdd.n1519 9.3005
R19597 vdd.n1606 vdd.n1605 9.3005
R19598 vdd.n1607 vdd.n1518 9.3005
R19599 vdd.n1609 vdd.n1608 9.3005
R19600 vdd.n1610 vdd.n1511 9.3005
R19601 vdd.n1612 vdd.n1611 9.3005
R19602 vdd.n1613 vdd.n1510 9.3005
R19603 vdd.n1615 vdd.n1614 9.3005
R19604 vdd.n1616 vdd.n1503 9.3005
R19605 vdd.n1618 vdd.n1617 9.3005
R19606 vdd.n1619 vdd.n1502 9.3005
R19607 vdd.n1621 vdd.n1620 9.3005
R19608 vdd.n1622 vdd.n1495 9.3005
R19609 vdd.n1624 vdd.n1623 9.3005
R19610 vdd.n1625 vdd.n1494 9.3005
R19611 vdd.n1627 vdd.n1626 9.3005
R19612 vdd.n1628 vdd.n1487 9.3005
R19613 vdd.n1630 vdd.n1629 9.3005
R19614 vdd.n1631 vdd.n1486 9.3005
R19615 vdd.n1633 vdd.n1632 9.3005
R19616 vdd.n1634 vdd.n1479 9.3005
R19617 vdd.n1636 vdd.n1635 9.3005
R19618 vdd.n1637 vdd.n1478 9.3005
R19619 vdd.n1639 vdd.n1638 9.3005
R19620 vdd.n1640 vdd.n1469 9.3005
R19621 vdd.n1642 vdd.n1641 9.3005
R19622 vdd.n1643 vdd.n1468 9.3005
R19623 vdd.n1645 vdd.n1644 9.3005
R19624 vdd.n1646 vdd.n1461 9.3005
R19625 vdd.n1648 vdd.n1647 9.3005
R19626 vdd.n1649 vdd.n1460 9.3005
R19627 vdd.n1651 vdd.n1650 9.3005
R19628 vdd.n1652 vdd.n1453 9.3005
R19629 vdd.n1654 vdd.n1653 9.3005
R19630 vdd.n1655 vdd.n1452 9.3005
R19631 vdd.n1657 vdd.n1656 9.3005
R19632 vdd.n1658 vdd.n1445 9.3005
R19633 vdd.n1660 vdd.n1659 9.3005
R19634 vdd.n1661 vdd.n1444 9.3005
R19635 vdd.n1663 vdd.n1662 9.3005
R19636 vdd.n1664 vdd.n1440 9.3005
R19637 vdd.n1666 vdd.n1665 9.3005
R19638 vdd.n1564 vdd.n1435 9.3005
R19639 vdd.n1431 vdd.n1430 9.3005
R19640 vdd.n1681 vdd.n1680 9.3005
R19641 vdd.n1682 vdd.n1429 9.3005
R19642 vdd.n1684 vdd.n1683 9.3005
R19643 vdd.n1419 vdd.n1418 9.3005
R19644 vdd.n1697 vdd.n1696 9.3005
R19645 vdd.n1698 vdd.n1417 9.3005
R19646 vdd.n1700 vdd.n1699 9.3005
R19647 vdd.n1407 vdd.n1406 9.3005
R19648 vdd.n1714 vdd.n1713 9.3005
R19649 vdd.n1715 vdd.n1405 9.3005
R19650 vdd.n1717 vdd.n1716 9.3005
R19651 vdd.n1396 vdd.n1395 9.3005
R19652 vdd.n1668 vdd.n1667 9.3005
R19653 vdd.n2012 vdd.n1729 9.3005
R19654 vdd.n1933 vdd.n1932 9.3005
R19655 vdd.n1928 vdd.n1927 9.3005
R19656 vdd.n1939 vdd.n1938 9.3005
R19657 vdd.n1941 vdd.n1940 9.3005
R19658 vdd.n1924 vdd.n1923 9.3005
R19659 vdd.n1947 vdd.n1946 9.3005
R19660 vdd.n1949 vdd.n1948 9.3005
R19661 vdd.n1921 vdd.n1918 9.3005
R19662 vdd.n1956 vdd.n1955 9.3005
R19663 vdd.n1984 vdd.n1983 9.3005
R19664 vdd.n1979 vdd.n1978 9.3005
R19665 vdd.n1990 vdd.n1989 9.3005
R19666 vdd.n1992 vdd.n1991 9.3005
R19667 vdd.n1975 vdd.n1974 9.3005
R19668 vdd.n1998 vdd.n1997 9.3005
R19669 vdd.n2000 vdd.n1999 9.3005
R19670 vdd.n1972 vdd.n1969 9.3005
R19671 vdd.n2007 vdd.n2006 9.3005
R19672 vdd.n1839 vdd.n1838 9.3005
R19673 vdd.n1834 vdd.n1833 9.3005
R19674 vdd.n1845 vdd.n1844 9.3005
R19675 vdd.n1847 vdd.n1846 9.3005
R19676 vdd.n1830 vdd.n1829 9.3005
R19677 vdd.n1853 vdd.n1852 9.3005
R19678 vdd.n1855 vdd.n1854 9.3005
R19679 vdd.n1827 vdd.n1824 9.3005
R19680 vdd.n1862 vdd.n1861 9.3005
R19681 vdd.n1890 vdd.n1889 9.3005
R19682 vdd.n1885 vdd.n1884 9.3005
R19683 vdd.n1896 vdd.n1895 9.3005
R19684 vdd.n1898 vdd.n1897 9.3005
R19685 vdd.n1881 vdd.n1880 9.3005
R19686 vdd.n1904 vdd.n1903 9.3005
R19687 vdd.n1906 vdd.n1905 9.3005
R19688 vdd.n1878 vdd.n1875 9.3005
R19689 vdd.n1913 vdd.n1912 9.3005
R19690 vdd.n1746 vdd.n1745 9.3005
R19691 vdd.n1741 vdd.n1740 9.3005
R19692 vdd.n1752 vdd.n1751 9.3005
R19693 vdd.n1754 vdd.n1753 9.3005
R19694 vdd.n1737 vdd.n1736 9.3005
R19695 vdd.n1760 vdd.n1759 9.3005
R19696 vdd.n1762 vdd.n1761 9.3005
R19697 vdd.n1734 vdd.n1731 9.3005
R19698 vdd.n1769 vdd.n1768 9.3005
R19699 vdd.n1797 vdd.n1796 9.3005
R19700 vdd.n1792 vdd.n1791 9.3005
R19701 vdd.n1803 vdd.n1802 9.3005
R19702 vdd.n1805 vdd.n1804 9.3005
R19703 vdd.n1788 vdd.n1787 9.3005
R19704 vdd.n1811 vdd.n1810 9.3005
R19705 vdd.n1813 vdd.n1812 9.3005
R19706 vdd.n1785 vdd.n1782 9.3005
R19707 vdd.n1820 vdd.n1819 9.3005
R19708 vdd.n288 vdd.n287 8.92171
R19709 vdd.n237 vdd.n236 8.92171
R19710 vdd.n194 vdd.n193 8.92171
R19711 vdd.n143 vdd.n142 8.92171
R19712 vdd.n101 vdd.n100 8.92171
R19713 vdd.n50 vdd.n49 8.92171
R19714 vdd.n1938 vdd.n1937 8.92171
R19715 vdd.n1989 vdd.n1988 8.92171
R19716 vdd.n1844 vdd.n1843 8.92171
R19717 vdd.n1895 vdd.n1894 8.92171
R19718 vdd.n1751 vdd.n1750 8.92171
R19719 vdd.n1802 vdd.n1801 8.92171
R19720 vdd.n215 vdd.n121 8.81535
R19721 vdd.n1916 vdd.n1822 8.81535
R19722 vdd.n2051 vdd.t2 8.72962
R19723 vdd.n3228 vdd.t4 8.72962
R19724 vdd.t0 vdd.n2025 8.50289
R19725 vdd.n493 vdd.t130 8.50289
R19726 vdd.n28 vdd.n14 8.42249
R19727 vdd.n1727 vdd.t153 8.27616
R19728 vdd.n3436 vdd.t88 8.27616
R19729 vdd.n3440 vdd.n3439 8.16225
R19730 vdd.n2012 vdd.n2011 8.16225
R19731 vdd.n284 vdd.n278 8.14595
R19732 vdd.n233 vdd.n227 8.14595
R19733 vdd.n190 vdd.n184 8.14595
R19734 vdd.n139 vdd.n133 8.14595
R19735 vdd.n97 vdd.n91 8.14595
R19736 vdd.n46 vdd.n40 8.14595
R19737 vdd.n1934 vdd.n1928 8.14595
R19738 vdd.n1985 vdd.n1979 8.14595
R19739 vdd.n1840 vdd.n1834 8.14595
R19740 vdd.n1891 vdd.n1885 8.14595
R19741 vdd.n1747 vdd.n1741 8.14595
R19742 vdd.n1798 vdd.n1792 8.14595
R19743 vdd.t96 vdd.n1415 8.04943
R19744 vdd.n3427 vdd.t98 8.04943
R19745 vdd.n2225 vdd.n962 7.70933
R19746 vdd.n2225 vdd.n965 7.70933
R19747 vdd.n2231 vdd.n951 7.70933
R19748 vdd.n2237 vdd.n951 7.70933
R19749 vdd.n2237 vdd.n944 7.70933
R19750 vdd.n2243 vdd.n944 7.70933
R19751 vdd.n2243 vdd.n947 7.70933
R19752 vdd.n2249 vdd.n940 7.70933
R19753 vdd.n2255 vdd.n934 7.70933
R19754 vdd.n2261 vdd.n921 7.70933
R19755 vdd.n2267 vdd.n921 7.70933
R19756 vdd.n2273 vdd.n915 7.70933
R19757 vdd.n2279 vdd.n908 7.70933
R19758 vdd.n2279 vdd.n911 7.70933
R19759 vdd.n2285 vdd.n904 7.70933
R19760 vdd.n2292 vdd.n890 7.70933
R19761 vdd.n2298 vdd.n890 7.70933
R19762 vdd.n2304 vdd.n884 7.70933
R19763 vdd.n2310 vdd.n880 7.70933
R19764 vdd.n2316 vdd.n874 7.70933
R19765 vdd.n2334 vdd.n856 7.70933
R19766 vdd.n2334 vdd.n849 7.70933
R19767 vdd.n2342 vdd.n849 7.70933
R19768 vdd.n2424 vdd.n833 7.70933
R19769 vdd.n2807 vdd.n785 7.70933
R19770 vdd.n2819 vdd.n774 7.70933
R19771 vdd.n2819 vdd.n768 7.70933
R19772 vdd.n2825 vdd.n768 7.70933
R19773 vdd.n2837 vdd.n759 7.70933
R19774 vdd.n2843 vdd.n753 7.70933
R19775 vdd.n2855 vdd.n740 7.70933
R19776 vdd.n2862 vdd.n733 7.70933
R19777 vdd.n2862 vdd.n736 7.70933
R19778 vdd.n2868 vdd.n729 7.70933
R19779 vdd.n2874 vdd.n715 7.70933
R19780 vdd.n2880 vdd.n715 7.70933
R19781 vdd.n2886 vdd.n709 7.70933
R19782 vdd.n2892 vdd.n702 7.70933
R19783 vdd.n2892 vdd.n705 7.70933
R19784 vdd.n2898 vdd.n698 7.70933
R19785 vdd.n2904 vdd.n692 7.70933
R19786 vdd.n2910 vdd.n679 7.70933
R19787 vdd.n2916 vdd.n679 7.70933
R19788 vdd.n2916 vdd.n671 7.70933
R19789 vdd.n2967 vdd.n671 7.70933
R19790 vdd.n2967 vdd.n674 7.70933
R19791 vdd.n2973 vdd.n631 7.70933
R19792 vdd.n3043 vdd.n631 7.70933
R19793 vdd.n283 vdd.n280 7.3702
R19794 vdd.n232 vdd.n229 7.3702
R19795 vdd.n189 vdd.n186 7.3702
R19796 vdd.n138 vdd.n135 7.3702
R19797 vdd.n96 vdd.n93 7.3702
R19798 vdd.n45 vdd.n42 7.3702
R19799 vdd.n1933 vdd.n1930 7.3702
R19800 vdd.n1984 vdd.n1981 7.3702
R19801 vdd.n1839 vdd.n1836 7.3702
R19802 vdd.n1890 vdd.n1887 7.3702
R19803 vdd.n1746 vdd.n1743 7.3702
R19804 vdd.n1797 vdd.n1794 7.3702
R19805 vdd.n934 vdd.t225 7.36923
R19806 vdd.n2898 vdd.t202 7.36923
R19807 vdd.n1694 vdd.t149 7.1425
R19808 vdd.n2249 vdd.t177 7.1425
R19809 vdd.n1253 vdd.t173 7.1425
R19810 vdd.n2831 vdd.t176 7.1425
R19811 vdd.n692 vdd.t186 7.1425
R19812 vdd.n3420 vdd.t94 7.1425
R19813 vdd.n1605 vdd.n1604 6.98232
R19814 vdd.n2113 vdd.n2112 6.98232
R19815 vdd.n3335 vdd.n3334 6.98232
R19816 vdd.n3127 vdd.n3126 6.98232
R19817 vdd.n1710 vdd.t140 6.91577
R19818 vdd.n325 vdd.t86 6.91577
R19819 vdd.n1253 vdd.t174 6.80241
R19820 vdd.n2831 vdd.t218 6.80241
R19821 vdd.n2017 vdd.t92 6.68904
R19822 vdd.n3261 vdd.t128 6.68904
R19823 vdd.n1380 vdd.t143 6.46231
R19824 vdd.n2273 vdd.t184 6.46231
R19825 vdd.t189 vdd.n884 6.46231
R19826 vdd.n2855 vdd.t194 6.46231
R19827 vdd.t210 vdd.n709 6.46231
R19828 vdd.t112 vdd.n492 6.46231
R19829 vdd.n2349 vdd.t222 6.34895
R19830 vdd.n2728 vdd.t207 6.34895
R19831 vdd.n3440 vdd.n309 6.27748
R19832 vdd.n2011 vdd.n2010 6.27748
R19833 vdd.n2870 vdd.n725 6.2444
R19834 vdd.n2289 vdd.n2288 6.2444
R19835 vdd.n2310 vdd.t215 5.89549
R19836 vdd.n753 vdd.t190 5.89549
R19837 vdd.n284 vdd.n283 5.81868
R19838 vdd.n233 vdd.n232 5.81868
R19839 vdd.n190 vdd.n189 5.81868
R19840 vdd.n139 vdd.n138 5.81868
R19841 vdd.n97 vdd.n96 5.81868
R19842 vdd.n46 vdd.n45 5.81868
R19843 vdd.n1934 vdd.n1933 5.81868
R19844 vdd.n1985 vdd.n1984 5.81868
R19845 vdd.n1840 vdd.n1839 5.81868
R19846 vdd.n1891 vdd.n1890 5.81868
R19847 vdd.n1747 vdd.n1746 5.81868
R19848 vdd.n1798 vdd.n1797 5.81868
R19849 vdd.n2432 vdd.n2431 5.77611
R19850 vdd.n1177 vdd.n1176 5.77611
R19851 vdd.n2740 vdd.n2739 5.77611
R19852 vdd.n2982 vdd.n663 5.77611
R19853 vdd.n3048 vdd.n627 5.77611
R19854 vdd.n2603 vdd.n2537 5.77611
R19855 vdd.n2357 vdd.n840 5.77611
R19856 vdd.n1313 vdd.n1145 5.77611
R19857 vdd.n1567 vdd.n1564 5.62474
R19858 vdd.n2076 vdd.n2073 5.62474
R19859 vdd.n3295 vdd.n3292 5.62474
R19860 vdd.n3082 vdd.n3079 5.62474
R19861 vdd.n2285 vdd.t204 5.55539
R19862 vdd.n729 vdd.t180 5.55539
R19863 vdd.n287 vdd.n278 5.04292
R19864 vdd.n236 vdd.n227 5.04292
R19865 vdd.n193 vdd.n184 5.04292
R19866 vdd.n142 vdd.n133 5.04292
R19867 vdd.n100 vdd.n91 5.04292
R19868 vdd.n49 vdd.n40 5.04292
R19869 vdd.n1937 vdd.n1928 5.04292
R19870 vdd.n1988 vdd.n1979 5.04292
R19871 vdd.n1843 vdd.n1834 5.04292
R19872 vdd.n1894 vdd.n1885 5.04292
R19873 vdd.n1750 vdd.n1741 5.04292
R19874 vdd.n1801 vdd.n1792 5.04292
R19875 vdd.n2043 vdd.t143 4.8752
R19876 vdd.t183 vdd.t196 4.8752
R19877 vdd.t226 vdd.t172 4.8752
R19878 vdd.n3236 vdd.t112 4.8752
R19879 vdd.n2433 vdd.n2432 4.83952
R19880 vdd.n1176 vdd.n1175 4.83952
R19881 vdd.n2741 vdd.n2740 4.83952
R19882 vdd.n663 vdd.n658 4.83952
R19883 vdd.n627 vdd.n622 4.83952
R19884 vdd.n2600 vdd.n2537 4.83952
R19885 vdd.n2360 vdd.n840 4.83952
R19886 vdd.n1316 vdd.n1145 4.83952
R19887 vdd.n1227 vdd.t192 4.76184
R19888 vdd.n2813 vdd.t178 4.76184
R19889 vdd.n2081 vdd.n2080 4.74817
R19890 vdd.n1349 vdd.n1344 4.74817
R19891 vdd.n1011 vdd.n1008 4.74817
R19892 vdd.n2174 vdd.n1007 4.74817
R19893 vdd.n2179 vdd.n1008 4.74817
R19894 vdd.n2178 vdd.n1007 4.74817
R19895 vdd.n521 vdd.n519 4.74817
R19896 vdd.n3197 vdd.n522 4.74817
R19897 vdd.n3200 vdd.n522 4.74817
R19898 vdd.n3201 vdd.n521 4.74817
R19899 vdd.n3089 vdd.n606 4.74817
R19900 vdd.n3085 vdd.n608 4.74817
R19901 vdd.n3088 vdd.n608 4.74817
R19902 vdd.n3093 vdd.n606 4.74817
R19903 vdd.n2080 vdd.n1107 4.74817
R19904 vdd.n1346 vdd.n1344 4.74817
R19905 vdd.n309 vdd.n308 4.7074
R19906 vdd.n215 vdd.n214 4.7074
R19907 vdd.n2010 vdd.n2009 4.7074
R19908 vdd.n1916 vdd.n1915 4.7074
R19909 vdd.t92 vdd.n1386 4.64847
R19910 vdd.t185 vdd.n915 4.64847
R19911 vdd.n2304 vdd.t224 4.64847
R19912 vdd.t213 vdd.n740 4.64847
R19913 vdd.n2886 vdd.t209 4.64847
R19914 vdd.n3252 vdd.t128 4.64847
R19915 vdd.n904 vdd.t74 4.53511
R19916 vdd.n2868 vdd.t37 4.53511
R19917 vdd.n1719 vdd.t140 4.42174
R19918 vdd.n2231 vdd.t15 4.42174
R19919 vdd.n1227 vdd.t60 4.42174
R19920 vdd.n2813 vdd.t67 4.42174
R19921 vdd.n674 vdd.t11 4.42174
R19922 vdd.n3434 vdd.t86 4.42174
R19923 vdd.n2859 vdd.n725 4.37123
R19924 vdd.n2290 vdd.n2289 4.37123
R19925 vdd.n2328 vdd.t211 4.30838
R19926 vdd.n2716 vdd.t198 4.30838
R19927 vdd.n288 vdd.n276 4.26717
R19928 vdd.n237 vdd.n225 4.26717
R19929 vdd.n194 vdd.n182 4.26717
R19930 vdd.n143 vdd.n131 4.26717
R19931 vdd.n101 vdd.n89 4.26717
R19932 vdd.n50 vdd.n38 4.26717
R19933 vdd.n1938 vdd.n1926 4.26717
R19934 vdd.n1989 vdd.n1977 4.26717
R19935 vdd.n1844 vdd.n1832 4.26717
R19936 vdd.n1895 vdd.n1883 4.26717
R19937 vdd.n1751 vdd.n1739 4.26717
R19938 vdd.n1802 vdd.n1790 4.26717
R19939 vdd.t149 vdd.n1414 4.19501
R19940 vdd.t94 vdd.n329 4.19501
R19941 vdd.n309 vdd.n215 4.10845
R19942 vdd.n2010 vdd.n1916 4.10845
R19943 vdd.n265 vdd.t146 4.06363
R19944 vdd.n265 vdd.t95 4.06363
R19945 vdd.n263 vdd.t87 4.06363
R19946 vdd.n263 vdd.t7 4.06363
R19947 vdd.n261 vdd.t103 4.06363
R19948 vdd.n261 vdd.t162 4.06363
R19949 vdd.n259 vdd.t131 4.06363
R19950 vdd.n259 vdd.t231 4.06363
R19951 vdd.n257 vdd.t237 4.06363
R19952 vdd.n257 vdd.t132 4.06363
R19953 vdd.n171 vdd.t138 4.06363
R19954 vdd.n171 vdd.t232 4.06363
R19955 vdd.n169 vdd.t242 4.06363
R19956 vdd.n169 vdd.t230 4.06363
R19957 vdd.n167 vdd.t108 4.06363
R19958 vdd.n167 vdd.t228 4.06363
R19959 vdd.n165 vdd.t148 4.06363
R19960 vdd.n165 vdd.t129 4.06363
R19961 vdd.n163 vdd.t113 4.06363
R19962 vdd.n163 vdd.t168 4.06363
R19963 vdd.n78 vdd.t99 4.06363
R19964 vdd.n78 vdd.t241 4.06363
R19965 vdd.n76 vdd.t240 4.06363
R19966 vdd.n76 vdd.t136 4.06363
R19967 vdd.n74 vdd.t102 4.06363
R19968 vdd.n74 vdd.t89 4.06363
R19969 vdd.n72 vdd.t243 4.06363
R19970 vdd.n72 vdd.t160 4.06363
R19971 vdd.n70 vdd.t124 4.06363
R19972 vdd.n70 vdd.t122 4.06363
R19973 vdd.n1958 vdd.t164 4.06363
R19974 vdd.n1958 vdd.t165 4.06363
R19975 vdd.n1960 vdd.t137 4.06363
R19976 vdd.n1960 vdd.t139 4.06363
R19977 vdd.n1962 vdd.t154 4.06363
R19978 vdd.n1962 vdd.t161 4.06363
R19979 vdd.n1964 vdd.t229 4.06363
R19980 vdd.n1964 vdd.t141 4.06363
R19981 vdd.n1966 vdd.t236 4.06363
R19982 vdd.n1966 vdd.t97 4.06363
R19983 vdd.n1864 vdd.t167 4.06363
R19984 vdd.n1864 vdd.t151 4.06363
R19985 vdd.n1866 vdd.t93 4.06363
R19986 vdd.n1866 vdd.t1 4.06363
R19987 vdd.n1868 vdd.t158 4.06363
R19988 vdd.n1868 vdd.t100 4.06363
R19989 vdd.n1870 vdd.t235 4.06363
R19990 vdd.n1870 vdd.t157 4.06363
R19991 vdd.n1872 vdd.t169 4.06363
R19992 vdd.n1872 vdd.t233 4.06363
R19993 vdd.n1771 vdd.t120 4.06363
R19994 vdd.n1771 vdd.t144 4.06363
R19995 vdd.n1773 vdd.t159 4.06363
R19996 vdd.n1773 vdd.t155 4.06363
R19997 vdd.n1775 vdd.t166 4.06363
R19998 vdd.n1775 vdd.t91 4.06363
R19999 vdd.n1777 vdd.t135 4.06363
R20000 vdd.n1777 vdd.t239 4.06363
R20001 vdd.n1779 vdd.t150 4.06363
R20002 vdd.n1779 vdd.t152 4.06363
R20003 vdd.n940 vdd.t217 3.96828
R20004 vdd.n2322 vdd.t195 3.96828
R20005 vdd.n2710 vdd.t214 3.96828
R20006 vdd.n2904 vdd.t203 3.96828
R20007 vdd.n26 vdd.t9 3.9605
R20008 vdd.n26 vdd.t111 3.9605
R20009 vdd.n23 vdd.t171 3.9605
R20010 vdd.n23 vdd.t8 3.9605
R20011 vdd.n21 vdd.t170 3.9605
R20012 vdd.n21 vdd.t105 3.9605
R20013 vdd.n20 vdd.t127 3.9605
R20014 vdd.n20 vdd.t110 3.9605
R20015 vdd.n15 vdd.t163 3.9605
R20016 vdd.n15 vdd.t104 3.9605
R20017 vdd.n16 vdd.t126 3.9605
R20018 vdd.n16 vdd.t109 3.9605
R20019 vdd.n18 vdd.t106 3.9605
R20020 vdd.n18 vdd.t125 3.9605
R20021 vdd.n25 vdd.t107 3.9605
R20022 vdd.n25 vdd.t142 3.9605
R20023 vdd.n2255 vdd.t217 3.74155
R20024 vdd.n874 vdd.t195 3.74155
R20025 vdd.n2837 vdd.t214 3.74155
R20026 vdd.n698 vdd.t203 3.74155
R20027 vdd.n7 vdd.t227 3.61217
R20028 vdd.n7 vdd.t191 3.61217
R20029 vdd.n8 vdd.t199 3.61217
R20030 vdd.n8 vdd.t219 3.61217
R20031 vdd.n10 vdd.t208 3.61217
R20032 vdd.n10 vdd.t179 3.61217
R20033 vdd.n12 vdd.t188 3.61217
R20034 vdd.n12 vdd.t206 3.61217
R20035 vdd.n5 vdd.t221 3.61217
R20036 vdd.n5 vdd.t201 3.61217
R20037 vdd.n3 vdd.t193 3.61217
R20038 vdd.n3 vdd.t223 3.61217
R20039 vdd.n1 vdd.t175 3.61217
R20040 vdd.n1 vdd.t212 3.61217
R20041 vdd.n0 vdd.t216 3.61217
R20042 vdd.n0 vdd.t197 3.61217
R20043 vdd.n292 vdd.n291 3.49141
R20044 vdd.n241 vdd.n240 3.49141
R20045 vdd.n198 vdd.n197 3.49141
R20046 vdd.n147 vdd.n146 3.49141
R20047 vdd.n105 vdd.n104 3.49141
R20048 vdd.n54 vdd.n53 3.49141
R20049 vdd.n1942 vdd.n1941 3.49141
R20050 vdd.n1993 vdd.n1992 3.49141
R20051 vdd.n1848 vdd.n1847 3.49141
R20052 vdd.n1899 vdd.n1898 3.49141
R20053 vdd.n1755 vdd.n1754 3.49141
R20054 vdd.n1806 vdd.n1805 3.49141
R20055 vdd.t211 vdd.n856 3.40145
R20056 vdd.n2496 vdd.t220 3.40145
R20057 vdd.n2800 vdd.t205 3.40145
R20058 vdd.n2825 vdd.t198 3.40145
R20059 vdd.n1702 vdd.t96 3.28809
R20060 vdd.n965 vdd.t15 3.28809
R20061 vdd.n2349 vdd.t60 3.28809
R20062 vdd.n2728 vdd.t67 3.28809
R20063 vdd.n2973 vdd.t11 3.28809
R20064 vdd.t98 vdd.n3426 3.28809
R20065 vdd.n1403 vdd.t153 3.06136
R20066 vdd.n2267 vdd.t185 3.06136
R20067 vdd.n1265 vdd.t224 3.06136
R20068 vdd.n2849 vdd.t213 3.06136
R20069 vdd.t209 vdd.n702 3.06136
R20070 vdd.t88 vdd.n3435 3.06136
R20071 vdd.n2342 vdd.t192 2.94799
R20072 vdd.t178 vdd.n774 2.94799
R20073 vdd.n2026 vdd.t0 2.83463
R20074 vdd.n3253 vdd.t130 2.83463
R20075 vdd.n295 vdd.n274 2.71565
R20076 vdd.n244 vdd.n223 2.71565
R20077 vdd.n201 vdd.n180 2.71565
R20078 vdd.n150 vdd.n129 2.71565
R20079 vdd.n108 vdd.n87 2.71565
R20080 vdd.n57 vdd.n36 2.71565
R20081 vdd.n1945 vdd.n1924 2.71565
R20082 vdd.n1996 vdd.n1975 2.71565
R20083 vdd.n1851 vdd.n1830 2.71565
R20084 vdd.n1902 vdd.n1881 2.71565
R20085 vdd.n1758 vdd.n1737 2.71565
R20086 vdd.n1809 vdd.n1788 2.71565
R20087 vdd.n2042 vdd.t2 2.6079
R20088 vdd.t4 vdd.n499 2.6079
R20089 vdd.n2316 vdd.t196 2.49453
R20090 vdd.n759 vdd.t226 2.49453
R20091 vdd.n282 vdd.n281 2.4129
R20092 vdd.n231 vdd.n230 2.4129
R20093 vdd.n188 vdd.n187 2.4129
R20094 vdd.n137 vdd.n136 2.4129
R20095 vdd.n95 vdd.n94 2.4129
R20096 vdd.n44 vdd.n43 2.4129
R20097 vdd.n1932 vdd.n1931 2.4129
R20098 vdd.n1983 vdd.n1982 2.4129
R20099 vdd.n1838 vdd.n1837 2.4129
R20100 vdd.n1889 vdd.n1888 2.4129
R20101 vdd.n1745 vdd.n1744 2.4129
R20102 vdd.n1796 vdd.n1795 2.4129
R20103 vdd.n2186 vdd.n1008 2.27742
R20104 vdd.n2186 vdd.n1007 2.27742
R20105 vdd.n3009 vdd.n522 2.27742
R20106 vdd.n3009 vdd.n521 2.27742
R20107 vdd.n3077 vdd.n608 2.27742
R20108 vdd.n3077 vdd.n606 2.27742
R20109 vdd.n2080 vdd.n2079 2.27742
R20110 vdd.n2079 vdd.n1344 2.27742
R20111 vdd.n911 vdd.t204 2.15444
R20112 vdd.n2292 vdd.t182 2.15444
R20113 vdd.n736 vdd.t181 2.15444
R20114 vdd.n2874 vdd.t180 2.15444
R20115 vdd.n296 vdd.n272 1.93989
R20116 vdd.n245 vdd.n221 1.93989
R20117 vdd.n202 vdd.n178 1.93989
R20118 vdd.n151 vdd.n127 1.93989
R20119 vdd.n109 vdd.n85 1.93989
R20120 vdd.n58 vdd.n34 1.93989
R20121 vdd.n1946 vdd.n1922 1.93989
R20122 vdd.n1997 vdd.n1973 1.93989
R20123 vdd.n1852 vdd.n1828 1.93989
R20124 vdd.n1903 vdd.n1879 1.93989
R20125 vdd.n1759 vdd.n1735 1.93989
R20126 vdd.n1810 vdd.n1786 1.93989
R20127 vdd.n1265 vdd.t215 1.81434
R20128 vdd.n2849 vdd.t190 1.81434
R20129 vdd.n1438 vdd.t47 1.47425
R20130 vdd.t33 vdd.n3411 1.47425
R20131 vdd.t222 vdd.n833 1.36088
R20132 vdd.n2807 vdd.t207 1.36088
R20133 vdd.t184 vdd.n908 1.24752
R20134 vdd.n2298 vdd.t189 1.24752
R20135 vdd.t194 vdd.n733 1.24752
R20136 vdd.n2880 vdd.t210 1.24752
R20137 vdd.n307 vdd.n267 1.16414
R20138 vdd.n300 vdd.n299 1.16414
R20139 vdd.n256 vdd.n216 1.16414
R20140 vdd.n249 vdd.n248 1.16414
R20141 vdd.n213 vdd.n173 1.16414
R20142 vdd.n206 vdd.n205 1.16414
R20143 vdd.n162 vdd.n122 1.16414
R20144 vdd.n155 vdd.n154 1.16414
R20145 vdd.n120 vdd.n80 1.16414
R20146 vdd.n113 vdd.n112 1.16414
R20147 vdd.n69 vdd.n29 1.16414
R20148 vdd.n62 vdd.n61 1.16414
R20149 vdd.n1957 vdd.n1917 1.16414
R20150 vdd.n1950 vdd.n1949 1.16414
R20151 vdd.n2008 vdd.n1968 1.16414
R20152 vdd.n2001 vdd.n2000 1.16414
R20153 vdd.n1863 vdd.n1823 1.16414
R20154 vdd.n1856 vdd.n1855 1.16414
R20155 vdd.n1914 vdd.n1874 1.16414
R20156 vdd.n1907 vdd.n1906 1.16414
R20157 vdd.n1770 vdd.n1730 1.16414
R20158 vdd.n1763 vdd.n1762 1.16414
R20159 vdd.n1821 vdd.n1781 1.16414
R20160 vdd.n1814 vdd.n1813 1.16414
R20161 vdd.n2011 vdd.n28 1.11236
R20162 vdd vdd.n3440 1.10453
R20163 vdd.n2034 vdd.t119 1.02079
R20164 vdd.t74 vdd.t182 1.02079
R20165 vdd.t181 vdd.t37 1.02079
R20166 vdd.n3244 vdd.t121 1.02079
R20167 vdd.n1568 vdd.n1567 0.970197
R20168 vdd.n2077 vdd.n2076 0.970197
R20169 vdd.n3296 vdd.n3295 0.970197
R20170 vdd.n3084 vdd.n3082 0.970197
R20171 vdd.n2322 vdd.t174 0.907421
R20172 vdd.n2710 vdd.t218 0.907421
R20173 vdd.t90 vdd.n1392 0.794056
R20174 vdd.n2061 vdd.t19 0.794056
R20175 vdd.t29 vdd.n511 0.794056
R20176 vdd.n481 vdd.t101 0.794056
R20177 vdd.n1711 vdd.t134 0.567326
R20178 vdd.n947 vdd.t177 0.567326
R20179 vdd.n2328 vdd.t173 0.567326
R20180 vdd.n2716 vdd.t176 0.567326
R20181 vdd.n2910 vdd.t186 0.567326
R20182 vdd.n3428 vdd.t6 0.567326
R20183 vdd.n2067 vdd.n1009 0.509646
R20184 vdd.n3209 vdd.n3208 0.509646
R20185 vdd.n3407 vdd.n3406 0.509646
R20186 vdd.n3289 vdd.n3288 0.509646
R20187 vdd.n3215 vdd.n514 0.509646
R20188 vdd.n2056 vdd.n1345 0.509646
R20189 vdd.n1673 vdd.n1435 0.509646
R20190 vdd.n1667 vdd.n1666 0.509646
R20191 vdd.n4 vdd.n2 0.459552
R20192 vdd.n11 vdd.n9 0.459552
R20193 vdd.n305 vdd.n304 0.388379
R20194 vdd.n271 vdd.n269 0.388379
R20195 vdd.n254 vdd.n253 0.388379
R20196 vdd.n220 vdd.n218 0.388379
R20197 vdd.n211 vdd.n210 0.388379
R20198 vdd.n177 vdd.n175 0.388379
R20199 vdd.n160 vdd.n159 0.388379
R20200 vdd.n126 vdd.n124 0.388379
R20201 vdd.n118 vdd.n117 0.388379
R20202 vdd.n84 vdd.n82 0.388379
R20203 vdd.n67 vdd.n66 0.388379
R20204 vdd.n33 vdd.n31 0.388379
R20205 vdd.n1955 vdd.n1954 0.388379
R20206 vdd.n1921 vdd.n1919 0.388379
R20207 vdd.n2006 vdd.n2005 0.388379
R20208 vdd.n1972 vdd.n1970 0.388379
R20209 vdd.n1861 vdd.n1860 0.388379
R20210 vdd.n1827 vdd.n1825 0.388379
R20211 vdd.n1912 vdd.n1911 0.388379
R20212 vdd.n1878 vdd.n1876 0.388379
R20213 vdd.n1768 vdd.n1767 0.388379
R20214 vdd.n1734 vdd.n1732 0.388379
R20215 vdd.n1819 vdd.n1818 0.388379
R20216 vdd.n1785 vdd.n1783 0.388379
R20217 vdd.n19 vdd.n17 0.387128
R20218 vdd.n24 vdd.n22 0.387128
R20219 vdd.n6 vdd.n4 0.358259
R20220 vdd.n13 vdd.n11 0.358259
R20221 vdd.n260 vdd.n258 0.358259
R20222 vdd.n262 vdd.n260 0.358259
R20223 vdd.n264 vdd.n262 0.358259
R20224 vdd.n266 vdd.n264 0.358259
R20225 vdd.n308 vdd.n266 0.358259
R20226 vdd.n166 vdd.n164 0.358259
R20227 vdd.n168 vdd.n166 0.358259
R20228 vdd.n170 vdd.n168 0.358259
R20229 vdd.n172 vdd.n170 0.358259
R20230 vdd.n214 vdd.n172 0.358259
R20231 vdd.n73 vdd.n71 0.358259
R20232 vdd.n75 vdd.n73 0.358259
R20233 vdd.n77 vdd.n75 0.358259
R20234 vdd.n79 vdd.n77 0.358259
R20235 vdd.n121 vdd.n79 0.358259
R20236 vdd.n2009 vdd.n1967 0.358259
R20237 vdd.n1967 vdd.n1965 0.358259
R20238 vdd.n1965 vdd.n1963 0.358259
R20239 vdd.n1963 vdd.n1961 0.358259
R20240 vdd.n1961 vdd.n1959 0.358259
R20241 vdd.n1915 vdd.n1873 0.358259
R20242 vdd.n1873 vdd.n1871 0.358259
R20243 vdd.n1871 vdd.n1869 0.358259
R20244 vdd.n1869 vdd.n1867 0.358259
R20245 vdd.n1867 vdd.n1865 0.358259
R20246 vdd.n1822 vdd.n1780 0.358259
R20247 vdd.n1780 vdd.n1778 0.358259
R20248 vdd.n1778 vdd.n1776 0.358259
R20249 vdd.n1776 vdd.n1774 0.358259
R20250 vdd.n1774 vdd.n1772 0.358259
R20251 vdd.t115 vdd.n1421 0.340595
R20252 vdd.n2261 vdd.t225 0.340595
R20253 vdd.n880 vdd.t183 0.340595
R20254 vdd.n2843 vdd.t172 0.340595
R20255 vdd.n705 vdd.t202 0.340595
R20256 vdd.n3419 vdd.t117 0.340595
R20257 vdd.n14 vdd.n6 0.334552
R20258 vdd.n14 vdd.n13 0.334552
R20259 vdd.n27 vdd.n19 0.21707
R20260 vdd.n27 vdd.n24 0.21707
R20261 vdd.n306 vdd.n268 0.155672
R20262 vdd.n298 vdd.n268 0.155672
R20263 vdd.n298 vdd.n297 0.155672
R20264 vdd.n297 vdd.n273 0.155672
R20265 vdd.n290 vdd.n273 0.155672
R20266 vdd.n290 vdd.n289 0.155672
R20267 vdd.n289 vdd.n277 0.155672
R20268 vdd.n282 vdd.n277 0.155672
R20269 vdd.n255 vdd.n217 0.155672
R20270 vdd.n247 vdd.n217 0.155672
R20271 vdd.n247 vdd.n246 0.155672
R20272 vdd.n246 vdd.n222 0.155672
R20273 vdd.n239 vdd.n222 0.155672
R20274 vdd.n239 vdd.n238 0.155672
R20275 vdd.n238 vdd.n226 0.155672
R20276 vdd.n231 vdd.n226 0.155672
R20277 vdd.n212 vdd.n174 0.155672
R20278 vdd.n204 vdd.n174 0.155672
R20279 vdd.n204 vdd.n203 0.155672
R20280 vdd.n203 vdd.n179 0.155672
R20281 vdd.n196 vdd.n179 0.155672
R20282 vdd.n196 vdd.n195 0.155672
R20283 vdd.n195 vdd.n183 0.155672
R20284 vdd.n188 vdd.n183 0.155672
R20285 vdd.n161 vdd.n123 0.155672
R20286 vdd.n153 vdd.n123 0.155672
R20287 vdd.n153 vdd.n152 0.155672
R20288 vdd.n152 vdd.n128 0.155672
R20289 vdd.n145 vdd.n128 0.155672
R20290 vdd.n145 vdd.n144 0.155672
R20291 vdd.n144 vdd.n132 0.155672
R20292 vdd.n137 vdd.n132 0.155672
R20293 vdd.n119 vdd.n81 0.155672
R20294 vdd.n111 vdd.n81 0.155672
R20295 vdd.n111 vdd.n110 0.155672
R20296 vdd.n110 vdd.n86 0.155672
R20297 vdd.n103 vdd.n86 0.155672
R20298 vdd.n103 vdd.n102 0.155672
R20299 vdd.n102 vdd.n90 0.155672
R20300 vdd.n95 vdd.n90 0.155672
R20301 vdd.n68 vdd.n30 0.155672
R20302 vdd.n60 vdd.n30 0.155672
R20303 vdd.n60 vdd.n59 0.155672
R20304 vdd.n59 vdd.n35 0.155672
R20305 vdd.n52 vdd.n35 0.155672
R20306 vdd.n52 vdd.n51 0.155672
R20307 vdd.n51 vdd.n39 0.155672
R20308 vdd.n44 vdd.n39 0.155672
R20309 vdd.n1956 vdd.n1918 0.155672
R20310 vdd.n1948 vdd.n1918 0.155672
R20311 vdd.n1948 vdd.n1947 0.155672
R20312 vdd.n1947 vdd.n1923 0.155672
R20313 vdd.n1940 vdd.n1923 0.155672
R20314 vdd.n1940 vdd.n1939 0.155672
R20315 vdd.n1939 vdd.n1927 0.155672
R20316 vdd.n1932 vdd.n1927 0.155672
R20317 vdd.n2007 vdd.n1969 0.155672
R20318 vdd.n1999 vdd.n1969 0.155672
R20319 vdd.n1999 vdd.n1998 0.155672
R20320 vdd.n1998 vdd.n1974 0.155672
R20321 vdd.n1991 vdd.n1974 0.155672
R20322 vdd.n1991 vdd.n1990 0.155672
R20323 vdd.n1990 vdd.n1978 0.155672
R20324 vdd.n1983 vdd.n1978 0.155672
R20325 vdd.n1862 vdd.n1824 0.155672
R20326 vdd.n1854 vdd.n1824 0.155672
R20327 vdd.n1854 vdd.n1853 0.155672
R20328 vdd.n1853 vdd.n1829 0.155672
R20329 vdd.n1846 vdd.n1829 0.155672
R20330 vdd.n1846 vdd.n1845 0.155672
R20331 vdd.n1845 vdd.n1833 0.155672
R20332 vdd.n1838 vdd.n1833 0.155672
R20333 vdd.n1913 vdd.n1875 0.155672
R20334 vdd.n1905 vdd.n1875 0.155672
R20335 vdd.n1905 vdd.n1904 0.155672
R20336 vdd.n1904 vdd.n1880 0.155672
R20337 vdd.n1897 vdd.n1880 0.155672
R20338 vdd.n1897 vdd.n1896 0.155672
R20339 vdd.n1896 vdd.n1884 0.155672
R20340 vdd.n1889 vdd.n1884 0.155672
R20341 vdd.n1769 vdd.n1731 0.155672
R20342 vdd.n1761 vdd.n1731 0.155672
R20343 vdd.n1761 vdd.n1760 0.155672
R20344 vdd.n1760 vdd.n1736 0.155672
R20345 vdd.n1753 vdd.n1736 0.155672
R20346 vdd.n1753 vdd.n1752 0.155672
R20347 vdd.n1752 vdd.n1740 0.155672
R20348 vdd.n1745 vdd.n1740 0.155672
R20349 vdd.n1820 vdd.n1782 0.155672
R20350 vdd.n1812 vdd.n1782 0.155672
R20351 vdd.n1812 vdd.n1811 0.155672
R20352 vdd.n1811 vdd.n1787 0.155672
R20353 vdd.n1804 vdd.n1787 0.155672
R20354 vdd.n1804 vdd.n1803 0.155672
R20355 vdd.n1803 vdd.n1791 0.155672
R20356 vdd.n1796 vdd.n1791 0.155672
R20357 vdd.n1014 vdd.n1006 0.152939
R20358 vdd.n1018 vdd.n1014 0.152939
R20359 vdd.n1019 vdd.n1018 0.152939
R20360 vdd.n1020 vdd.n1019 0.152939
R20361 vdd.n1021 vdd.n1020 0.152939
R20362 vdd.n1025 vdd.n1021 0.152939
R20363 vdd.n1026 vdd.n1025 0.152939
R20364 vdd.n1027 vdd.n1026 0.152939
R20365 vdd.n1028 vdd.n1027 0.152939
R20366 vdd.n1032 vdd.n1028 0.152939
R20367 vdd.n1033 vdd.n1032 0.152939
R20368 vdd.n1034 vdd.n1033 0.152939
R20369 vdd.n2150 vdd.n1034 0.152939
R20370 vdd.n2150 vdd.n2149 0.152939
R20371 vdd.n2149 vdd.n2148 0.152939
R20372 vdd.n2148 vdd.n1040 0.152939
R20373 vdd.n1045 vdd.n1040 0.152939
R20374 vdd.n1046 vdd.n1045 0.152939
R20375 vdd.n1047 vdd.n1046 0.152939
R20376 vdd.n1051 vdd.n1047 0.152939
R20377 vdd.n1052 vdd.n1051 0.152939
R20378 vdd.n1053 vdd.n1052 0.152939
R20379 vdd.n1054 vdd.n1053 0.152939
R20380 vdd.n1058 vdd.n1054 0.152939
R20381 vdd.n1059 vdd.n1058 0.152939
R20382 vdd.n1060 vdd.n1059 0.152939
R20383 vdd.n1061 vdd.n1060 0.152939
R20384 vdd.n1065 vdd.n1061 0.152939
R20385 vdd.n1066 vdd.n1065 0.152939
R20386 vdd.n1067 vdd.n1066 0.152939
R20387 vdd.n1068 vdd.n1067 0.152939
R20388 vdd.n1072 vdd.n1068 0.152939
R20389 vdd.n1073 vdd.n1072 0.152939
R20390 vdd.n1074 vdd.n1073 0.152939
R20391 vdd.n2111 vdd.n1074 0.152939
R20392 vdd.n2111 vdd.n2110 0.152939
R20393 vdd.n2110 vdd.n2109 0.152939
R20394 vdd.n2109 vdd.n1080 0.152939
R20395 vdd.n1085 vdd.n1080 0.152939
R20396 vdd.n1086 vdd.n1085 0.152939
R20397 vdd.n1087 vdd.n1086 0.152939
R20398 vdd.n1091 vdd.n1087 0.152939
R20399 vdd.n1092 vdd.n1091 0.152939
R20400 vdd.n1093 vdd.n1092 0.152939
R20401 vdd.n1094 vdd.n1093 0.152939
R20402 vdd.n1098 vdd.n1094 0.152939
R20403 vdd.n1099 vdd.n1098 0.152939
R20404 vdd.n1100 vdd.n1099 0.152939
R20405 vdd.n1101 vdd.n1100 0.152939
R20406 vdd.n1105 vdd.n1101 0.152939
R20407 vdd.n1106 vdd.n1105 0.152939
R20408 vdd.n2185 vdd.n1009 0.152939
R20409 vdd.n2014 vdd.n2013 0.152939
R20410 vdd.n2014 vdd.n1383 0.152939
R20411 vdd.n2029 vdd.n1383 0.152939
R20412 vdd.n2030 vdd.n2029 0.152939
R20413 vdd.n2031 vdd.n2030 0.152939
R20414 vdd.n2031 vdd.n1372 0.152939
R20415 vdd.n2046 vdd.n1372 0.152939
R20416 vdd.n2047 vdd.n2046 0.152939
R20417 vdd.n2048 vdd.n2047 0.152939
R20418 vdd.n2048 vdd.n1360 0.152939
R20419 vdd.n2065 vdd.n1360 0.152939
R20420 vdd.n2066 vdd.n2065 0.152939
R20421 vdd.n2067 vdd.n2066 0.152939
R20422 vdd.n527 vdd.n524 0.152939
R20423 vdd.n528 vdd.n527 0.152939
R20424 vdd.n529 vdd.n528 0.152939
R20425 vdd.n530 vdd.n529 0.152939
R20426 vdd.n533 vdd.n530 0.152939
R20427 vdd.n534 vdd.n533 0.152939
R20428 vdd.n535 vdd.n534 0.152939
R20429 vdd.n536 vdd.n535 0.152939
R20430 vdd.n539 vdd.n536 0.152939
R20431 vdd.n540 vdd.n539 0.152939
R20432 vdd.n541 vdd.n540 0.152939
R20433 vdd.n542 vdd.n541 0.152939
R20434 vdd.n547 vdd.n542 0.152939
R20435 vdd.n548 vdd.n547 0.152939
R20436 vdd.n549 vdd.n548 0.152939
R20437 vdd.n550 vdd.n549 0.152939
R20438 vdd.n553 vdd.n550 0.152939
R20439 vdd.n554 vdd.n553 0.152939
R20440 vdd.n555 vdd.n554 0.152939
R20441 vdd.n556 vdd.n555 0.152939
R20442 vdd.n559 vdd.n556 0.152939
R20443 vdd.n560 vdd.n559 0.152939
R20444 vdd.n561 vdd.n560 0.152939
R20445 vdd.n562 vdd.n561 0.152939
R20446 vdd.n565 vdd.n562 0.152939
R20447 vdd.n566 vdd.n565 0.152939
R20448 vdd.n567 vdd.n566 0.152939
R20449 vdd.n568 vdd.n567 0.152939
R20450 vdd.n571 vdd.n568 0.152939
R20451 vdd.n572 vdd.n571 0.152939
R20452 vdd.n573 vdd.n572 0.152939
R20453 vdd.n574 vdd.n573 0.152939
R20454 vdd.n577 vdd.n574 0.152939
R20455 vdd.n578 vdd.n577 0.152939
R20456 vdd.n3125 vdd.n578 0.152939
R20457 vdd.n3125 vdd.n3124 0.152939
R20458 vdd.n3124 vdd.n3123 0.152939
R20459 vdd.n3123 vdd.n582 0.152939
R20460 vdd.n587 vdd.n582 0.152939
R20461 vdd.n588 vdd.n587 0.152939
R20462 vdd.n591 vdd.n588 0.152939
R20463 vdd.n592 vdd.n591 0.152939
R20464 vdd.n593 vdd.n592 0.152939
R20465 vdd.n594 vdd.n593 0.152939
R20466 vdd.n597 vdd.n594 0.152939
R20467 vdd.n598 vdd.n597 0.152939
R20468 vdd.n599 vdd.n598 0.152939
R20469 vdd.n600 vdd.n599 0.152939
R20470 vdd.n603 vdd.n600 0.152939
R20471 vdd.n604 vdd.n603 0.152939
R20472 vdd.n605 vdd.n604 0.152939
R20473 vdd.n3208 vdd.n518 0.152939
R20474 vdd.n3209 vdd.n508 0.152939
R20475 vdd.n3223 vdd.n508 0.152939
R20476 vdd.n3224 vdd.n3223 0.152939
R20477 vdd.n3225 vdd.n3224 0.152939
R20478 vdd.n3225 vdd.n496 0.152939
R20479 vdd.n3239 vdd.n496 0.152939
R20480 vdd.n3240 vdd.n3239 0.152939
R20481 vdd.n3241 vdd.n3240 0.152939
R20482 vdd.n3241 vdd.n484 0.152939
R20483 vdd.n3256 vdd.n484 0.152939
R20484 vdd.n3257 vdd.n3256 0.152939
R20485 vdd.n3258 vdd.n3257 0.152939
R20486 vdd.n3258 vdd.n310 0.152939
R20487 vdd.n320 vdd.n311 0.152939
R20488 vdd.n321 vdd.n320 0.152939
R20489 vdd.n322 vdd.n321 0.152939
R20490 vdd.n331 vdd.n322 0.152939
R20491 vdd.n332 vdd.n331 0.152939
R20492 vdd.n333 vdd.n332 0.152939
R20493 vdd.n334 vdd.n333 0.152939
R20494 vdd.n342 vdd.n334 0.152939
R20495 vdd.n343 vdd.n342 0.152939
R20496 vdd.n344 vdd.n343 0.152939
R20497 vdd.n345 vdd.n344 0.152939
R20498 vdd.n353 vdd.n345 0.152939
R20499 vdd.n3407 vdd.n353 0.152939
R20500 vdd.n3406 vdd.n354 0.152939
R20501 vdd.n357 vdd.n354 0.152939
R20502 vdd.n361 vdd.n357 0.152939
R20503 vdd.n362 vdd.n361 0.152939
R20504 vdd.n363 vdd.n362 0.152939
R20505 vdd.n364 vdd.n363 0.152939
R20506 vdd.n365 vdd.n364 0.152939
R20507 vdd.n369 vdd.n365 0.152939
R20508 vdd.n370 vdd.n369 0.152939
R20509 vdd.n371 vdd.n370 0.152939
R20510 vdd.n372 vdd.n371 0.152939
R20511 vdd.n376 vdd.n372 0.152939
R20512 vdd.n377 vdd.n376 0.152939
R20513 vdd.n378 vdd.n377 0.152939
R20514 vdd.n379 vdd.n378 0.152939
R20515 vdd.n383 vdd.n379 0.152939
R20516 vdd.n384 vdd.n383 0.152939
R20517 vdd.n385 vdd.n384 0.152939
R20518 vdd.n3372 vdd.n385 0.152939
R20519 vdd.n3372 vdd.n3371 0.152939
R20520 vdd.n3371 vdd.n3370 0.152939
R20521 vdd.n3370 vdd.n391 0.152939
R20522 vdd.n396 vdd.n391 0.152939
R20523 vdd.n397 vdd.n396 0.152939
R20524 vdd.n398 vdd.n397 0.152939
R20525 vdd.n402 vdd.n398 0.152939
R20526 vdd.n403 vdd.n402 0.152939
R20527 vdd.n404 vdd.n403 0.152939
R20528 vdd.n405 vdd.n404 0.152939
R20529 vdd.n409 vdd.n405 0.152939
R20530 vdd.n410 vdd.n409 0.152939
R20531 vdd.n411 vdd.n410 0.152939
R20532 vdd.n412 vdd.n411 0.152939
R20533 vdd.n416 vdd.n412 0.152939
R20534 vdd.n417 vdd.n416 0.152939
R20535 vdd.n418 vdd.n417 0.152939
R20536 vdd.n419 vdd.n418 0.152939
R20537 vdd.n423 vdd.n419 0.152939
R20538 vdd.n424 vdd.n423 0.152939
R20539 vdd.n425 vdd.n424 0.152939
R20540 vdd.n3333 vdd.n425 0.152939
R20541 vdd.n3333 vdd.n3332 0.152939
R20542 vdd.n3332 vdd.n3331 0.152939
R20543 vdd.n3331 vdd.n431 0.152939
R20544 vdd.n436 vdd.n431 0.152939
R20545 vdd.n437 vdd.n436 0.152939
R20546 vdd.n438 vdd.n437 0.152939
R20547 vdd.n442 vdd.n438 0.152939
R20548 vdd.n443 vdd.n442 0.152939
R20549 vdd.n444 vdd.n443 0.152939
R20550 vdd.n445 vdd.n444 0.152939
R20551 vdd.n449 vdd.n445 0.152939
R20552 vdd.n450 vdd.n449 0.152939
R20553 vdd.n451 vdd.n450 0.152939
R20554 vdd.n452 vdd.n451 0.152939
R20555 vdd.n456 vdd.n452 0.152939
R20556 vdd.n457 vdd.n456 0.152939
R20557 vdd.n458 vdd.n457 0.152939
R20558 vdd.n459 vdd.n458 0.152939
R20559 vdd.n463 vdd.n459 0.152939
R20560 vdd.n464 vdd.n463 0.152939
R20561 vdd.n465 vdd.n464 0.152939
R20562 vdd.n3289 vdd.n465 0.152939
R20563 vdd.n3216 vdd.n3215 0.152939
R20564 vdd.n3217 vdd.n3216 0.152939
R20565 vdd.n3217 vdd.n502 0.152939
R20566 vdd.n3231 vdd.n502 0.152939
R20567 vdd.n3232 vdd.n3231 0.152939
R20568 vdd.n3233 vdd.n3232 0.152939
R20569 vdd.n3233 vdd.n489 0.152939
R20570 vdd.n3247 vdd.n489 0.152939
R20571 vdd.n3248 vdd.n3247 0.152939
R20572 vdd.n3249 vdd.n3248 0.152939
R20573 vdd.n3249 vdd.n477 0.152939
R20574 vdd.n3264 vdd.n477 0.152939
R20575 vdd.n3265 vdd.n3264 0.152939
R20576 vdd.n3266 vdd.n3265 0.152939
R20577 vdd.n3266 vdd.n475 0.152939
R20578 vdd.n3270 vdd.n475 0.152939
R20579 vdd.n3271 vdd.n3270 0.152939
R20580 vdd.n3272 vdd.n3271 0.152939
R20581 vdd.n3272 vdd.n472 0.152939
R20582 vdd.n3276 vdd.n472 0.152939
R20583 vdd.n3277 vdd.n3276 0.152939
R20584 vdd.n3278 vdd.n3277 0.152939
R20585 vdd.n3278 vdd.n469 0.152939
R20586 vdd.n3282 vdd.n469 0.152939
R20587 vdd.n3283 vdd.n3282 0.152939
R20588 vdd.n3284 vdd.n3283 0.152939
R20589 vdd.n3284 vdd.n466 0.152939
R20590 vdd.n3288 vdd.n466 0.152939
R20591 vdd.n3078 vdd.n514 0.152939
R20592 vdd.n2078 vdd.n1345 0.152939
R20593 vdd.n1674 vdd.n1673 0.152939
R20594 vdd.n1675 vdd.n1674 0.152939
R20595 vdd.n1675 vdd.n1424 0.152939
R20596 vdd.n1689 vdd.n1424 0.152939
R20597 vdd.n1690 vdd.n1689 0.152939
R20598 vdd.n1691 vdd.n1690 0.152939
R20599 vdd.n1691 vdd.n1411 0.152939
R20600 vdd.n1705 vdd.n1411 0.152939
R20601 vdd.n1706 vdd.n1705 0.152939
R20602 vdd.n1707 vdd.n1706 0.152939
R20603 vdd.n1707 vdd.n1400 0.152939
R20604 vdd.n1722 vdd.n1400 0.152939
R20605 vdd.n1723 vdd.n1722 0.152939
R20606 vdd.n1724 vdd.n1723 0.152939
R20607 vdd.n1724 vdd.n1389 0.152939
R20608 vdd.n2020 vdd.n1389 0.152939
R20609 vdd.n2021 vdd.n2020 0.152939
R20610 vdd.n2022 vdd.n2021 0.152939
R20611 vdd.n2022 vdd.n1377 0.152939
R20612 vdd.n2037 vdd.n1377 0.152939
R20613 vdd.n2038 vdd.n2037 0.152939
R20614 vdd.n2039 vdd.n2038 0.152939
R20615 vdd.n2039 vdd.n1367 0.152939
R20616 vdd.n2054 vdd.n1367 0.152939
R20617 vdd.n2055 vdd.n2054 0.152939
R20618 vdd.n2058 vdd.n2055 0.152939
R20619 vdd.n2058 vdd.n2057 0.152939
R20620 vdd.n2057 vdd.n2056 0.152939
R20621 vdd.n1666 vdd.n1440 0.152939
R20622 vdd.n1662 vdd.n1440 0.152939
R20623 vdd.n1662 vdd.n1661 0.152939
R20624 vdd.n1661 vdd.n1660 0.152939
R20625 vdd.n1660 vdd.n1445 0.152939
R20626 vdd.n1656 vdd.n1445 0.152939
R20627 vdd.n1656 vdd.n1655 0.152939
R20628 vdd.n1655 vdd.n1654 0.152939
R20629 vdd.n1654 vdd.n1453 0.152939
R20630 vdd.n1650 vdd.n1453 0.152939
R20631 vdd.n1650 vdd.n1649 0.152939
R20632 vdd.n1649 vdd.n1648 0.152939
R20633 vdd.n1648 vdd.n1461 0.152939
R20634 vdd.n1644 vdd.n1461 0.152939
R20635 vdd.n1644 vdd.n1643 0.152939
R20636 vdd.n1643 vdd.n1642 0.152939
R20637 vdd.n1642 vdd.n1469 0.152939
R20638 vdd.n1638 vdd.n1469 0.152939
R20639 vdd.n1638 vdd.n1637 0.152939
R20640 vdd.n1637 vdd.n1636 0.152939
R20641 vdd.n1636 vdd.n1479 0.152939
R20642 vdd.n1632 vdd.n1479 0.152939
R20643 vdd.n1632 vdd.n1631 0.152939
R20644 vdd.n1631 vdd.n1630 0.152939
R20645 vdd.n1630 vdd.n1487 0.152939
R20646 vdd.n1626 vdd.n1487 0.152939
R20647 vdd.n1626 vdd.n1625 0.152939
R20648 vdd.n1625 vdd.n1624 0.152939
R20649 vdd.n1624 vdd.n1495 0.152939
R20650 vdd.n1620 vdd.n1495 0.152939
R20651 vdd.n1620 vdd.n1619 0.152939
R20652 vdd.n1619 vdd.n1618 0.152939
R20653 vdd.n1618 vdd.n1503 0.152939
R20654 vdd.n1614 vdd.n1503 0.152939
R20655 vdd.n1614 vdd.n1613 0.152939
R20656 vdd.n1613 vdd.n1612 0.152939
R20657 vdd.n1612 vdd.n1511 0.152939
R20658 vdd.n1608 vdd.n1511 0.152939
R20659 vdd.n1608 vdd.n1607 0.152939
R20660 vdd.n1607 vdd.n1606 0.152939
R20661 vdd.n1606 vdd.n1519 0.152939
R20662 vdd.n1526 vdd.n1519 0.152939
R20663 vdd.n1596 vdd.n1526 0.152939
R20664 vdd.n1596 vdd.n1595 0.152939
R20665 vdd.n1595 vdd.n1594 0.152939
R20666 vdd.n1594 vdd.n1527 0.152939
R20667 vdd.n1590 vdd.n1527 0.152939
R20668 vdd.n1590 vdd.n1589 0.152939
R20669 vdd.n1589 vdd.n1588 0.152939
R20670 vdd.n1588 vdd.n1534 0.152939
R20671 vdd.n1584 vdd.n1534 0.152939
R20672 vdd.n1584 vdd.n1583 0.152939
R20673 vdd.n1583 vdd.n1582 0.152939
R20674 vdd.n1582 vdd.n1542 0.152939
R20675 vdd.n1578 vdd.n1542 0.152939
R20676 vdd.n1578 vdd.n1577 0.152939
R20677 vdd.n1577 vdd.n1576 0.152939
R20678 vdd.n1576 vdd.n1550 0.152939
R20679 vdd.n1572 vdd.n1550 0.152939
R20680 vdd.n1572 vdd.n1571 0.152939
R20681 vdd.n1571 vdd.n1570 0.152939
R20682 vdd.n1570 vdd.n1558 0.152939
R20683 vdd.n1558 vdd.n1435 0.152939
R20684 vdd.n1667 vdd.n1430 0.152939
R20685 vdd.n1681 vdd.n1430 0.152939
R20686 vdd.n1682 vdd.n1681 0.152939
R20687 vdd.n1683 vdd.n1682 0.152939
R20688 vdd.n1683 vdd.n1418 0.152939
R20689 vdd.n1697 vdd.n1418 0.152939
R20690 vdd.n1698 vdd.n1697 0.152939
R20691 vdd.n1699 vdd.n1698 0.152939
R20692 vdd.n1699 vdd.n1406 0.152939
R20693 vdd.n1714 vdd.n1406 0.152939
R20694 vdd.n1715 vdd.n1714 0.152939
R20695 vdd.n1716 vdd.n1715 0.152939
R20696 vdd.n1716 vdd.n1395 0.152939
R20697 vdd.n2013 vdd.n2012 0.145814
R20698 vdd.n3439 vdd.n310 0.145814
R20699 vdd.n3439 vdd.n311 0.145814
R20700 vdd.n2012 vdd.n1395 0.145814
R20701 vdd.n2186 vdd.n2185 0.110256
R20702 vdd.n3009 vdd.n518 0.110256
R20703 vdd.n3078 vdd.n3077 0.110256
R20704 vdd.n2079 vdd.n2078 0.110256
R20705 vdd.n2186 vdd.n1006 0.0431829
R20706 vdd.n2079 vdd.n1106 0.0431829
R20707 vdd.n3009 vdd.n524 0.0431829
R20708 vdd.n3077 vdd.n605 0.0431829
R20709 vdd vdd.n28 0.00833333
R20710 a_n2804_13878.n2 a_n2804_13878.n0 98.9633
R20711 a_n2804_13878.n5 a_n2804_13878.n3 98.7517
R20712 a_n2804_13878.n25 a_n2804_13878.n24 98.6055
R20713 a_n2804_13878.n27 a_n2804_13878.n26 98.6055
R20714 a_n2804_13878.n2 a_n2804_13878.n1 98.6055
R20715 a_n2804_13878.n13 a_n2804_13878.n12 98.6055
R20716 a_n2804_13878.n11 a_n2804_13878.n10 98.6055
R20717 a_n2804_13878.n9 a_n2804_13878.n8 98.6055
R20718 a_n2804_13878.n7 a_n2804_13878.n6 98.6055
R20719 a_n2804_13878.n5 a_n2804_13878.n4 98.6055
R20720 a_n2804_13878.n29 a_n2804_13878.n28 98.6054
R20721 a_n2804_13878.n23 a_n2804_13878.n22 98.6054
R20722 a_n2804_13878.n15 a_n2804_13878.t1 74.6477
R20723 a_n2804_13878.n20 a_n2804_13878.t2 74.2899
R20724 a_n2804_13878.n17 a_n2804_13878.t3 74.2899
R20725 a_n2804_13878.n16 a_n2804_13878.t0 74.2899
R20726 a_n2804_13878.n19 a_n2804_13878.n18 70.6783
R20727 a_n2804_13878.n15 a_n2804_13878.n14 70.6783
R20728 a_n2804_13878.n21 a_n2804_13878.n13 15.7159
R20729 a_n2804_13878.n23 a_n2804_13878.n21 12.6495
R20730 a_n2804_13878.n21 a_n2804_13878.n20 8.38735
R20731 a_n2804_13878.n22 a_n2804_13878.t15 3.61217
R20732 a_n2804_13878.n22 a_n2804_13878.t24 3.61217
R20733 a_n2804_13878.n24 a_n2804_13878.t28 3.61217
R20734 a_n2804_13878.n24 a_n2804_13878.t14 3.61217
R20735 a_n2804_13878.n26 a_n2804_13878.t18 3.61217
R20736 a_n2804_13878.n26 a_n2804_13878.t19 3.61217
R20737 a_n2804_13878.n1 a_n2804_13878.t8 3.61217
R20738 a_n2804_13878.n1 a_n2804_13878.t20 3.61217
R20739 a_n2804_13878.n0 a_n2804_13878.t25 3.61217
R20740 a_n2804_13878.n0 a_n2804_13878.t31 3.61217
R20741 a_n2804_13878.n18 a_n2804_13878.t6 3.61217
R20742 a_n2804_13878.n18 a_n2804_13878.t7 3.61217
R20743 a_n2804_13878.n14 a_n2804_13878.t4 3.61217
R20744 a_n2804_13878.n14 a_n2804_13878.t5 3.61217
R20745 a_n2804_13878.n12 a_n2804_13878.t21 3.61217
R20746 a_n2804_13878.n12 a_n2804_13878.t9 3.61217
R20747 a_n2804_13878.n10 a_n2804_13878.t26 3.61217
R20748 a_n2804_13878.n10 a_n2804_13878.t11 3.61217
R20749 a_n2804_13878.n8 a_n2804_13878.t10 3.61217
R20750 a_n2804_13878.n8 a_n2804_13878.t13 3.61217
R20751 a_n2804_13878.n6 a_n2804_13878.t23 3.61217
R20752 a_n2804_13878.n6 a_n2804_13878.t16 3.61217
R20753 a_n2804_13878.n4 a_n2804_13878.t27 3.61217
R20754 a_n2804_13878.n4 a_n2804_13878.t17 3.61217
R20755 a_n2804_13878.n3 a_n2804_13878.t12 3.61217
R20756 a_n2804_13878.n3 a_n2804_13878.t22 3.61217
R20757 a_n2804_13878.n29 a_n2804_13878.t29 3.61217
R20758 a_n2804_13878.t30 a_n2804_13878.n29 3.61217
R20759 a_n2804_13878.n16 a_n2804_13878.n15 0.358259
R20760 a_n2804_13878.n19 a_n2804_13878.n17 0.358259
R20761 a_n2804_13878.n20 a_n2804_13878.n19 0.358259
R20762 a_n2804_13878.n28 a_n2804_13878.n2 0.358259
R20763 a_n2804_13878.n28 a_n2804_13878.n27 0.358259
R20764 a_n2804_13878.n27 a_n2804_13878.n25 0.358259
R20765 a_n2804_13878.n25 a_n2804_13878.n23 0.358259
R20766 a_n2804_13878.n7 a_n2804_13878.n5 0.146627
R20767 a_n2804_13878.n9 a_n2804_13878.n7 0.146627
R20768 a_n2804_13878.n11 a_n2804_13878.n9 0.146627
R20769 a_n2804_13878.n13 a_n2804_13878.n11 0.146627
R20770 a_n2804_13878.n17 a_n2804_13878.n16 0.101793
R20771 a_n8300_8799.n145 a_n8300_8799.t113 490.524
R20772 a_n8300_8799.n156 a_n8300_8799.t49 490.524
R20773 a_n8300_8799.n168 a_n8300_8799.t97 490.524
R20774 a_n8300_8799.n111 a_n8300_8799.t89 490.524
R20775 a_n8300_8799.n122 a_n8300_8799.t96 490.524
R20776 a_n8300_8799.n134 a_n8300_8799.t98 490.524
R20777 a_n8300_8799.n34 a_n8300_8799.t51 484.3
R20778 a_n8300_8799.n151 a_n8300_8799.t50 464.166
R20779 a_n8300_8799.n150 a_n8300_8799.t100 464.166
R20780 a_n8300_8799.n141 a_n8300_8799.t61 464.166
R20781 a_n8300_8799.n149 a_n8300_8799.t53 464.166
R20782 a_n8300_8799.n148 a_n8300_8799.t105 464.166
R20783 a_n8300_8799.n142 a_n8300_8799.t77 464.166
R20784 a_n8300_8799.n147 a_n8300_8799.t62 464.166
R20785 a_n8300_8799.n146 a_n8300_8799.t117 464.166
R20786 a_n8300_8799.n143 a_n8300_8799.t88 464.166
R20787 a_n8300_8799.n144 a_n8300_8799.t64 464.166
R20788 a_n8300_8799.n43 a_n8300_8799.t57 484.3
R20789 a_n8300_8799.n162 a_n8300_8799.t56 464.166
R20790 a_n8300_8799.n161 a_n8300_8799.t112 464.166
R20791 a_n8300_8799.n152 a_n8300_8799.t66 464.166
R20792 a_n8300_8799.n160 a_n8300_8799.t60 464.166
R20793 a_n8300_8799.n159 a_n8300_8799.t114 464.166
R20794 a_n8300_8799.n153 a_n8300_8799.t86 464.166
R20795 a_n8300_8799.n158 a_n8300_8799.t69 464.166
R20796 a_n8300_8799.n157 a_n8300_8799.t52 464.166
R20797 a_n8300_8799.n154 a_n8300_8799.t95 464.166
R20798 a_n8300_8799.n155 a_n8300_8799.t70 464.166
R20799 a_n8300_8799.n52 a_n8300_8799.t85 484.3
R20800 a_n8300_8799.n174 a_n8300_8799.t99 464.166
R20801 a_n8300_8799.n173 a_n8300_8799.t59 464.166
R20802 a_n8300_8799.n164 a_n8300_8799.t110 464.166
R20803 a_n8300_8799.n172 a_n8300_8799.t73 464.166
R20804 a_n8300_8799.n171 a_n8300_8799.t104 464.166
R20805 a_n8300_8799.n165 a_n8300_8799.t63 464.166
R20806 a_n8300_8799.n170 a_n8300_8799.t91 464.166
R20807 a_n8300_8799.n169 a_n8300_8799.t55 464.166
R20808 a_n8300_8799.n166 a_n8300_8799.t82 464.166
R20809 a_n8300_8799.n167 a_n8300_8799.t68 464.166
R20810 a_n8300_8799.n110 a_n8300_8799.t111 464.166
R20811 a_n8300_8799.n109 a_n8300_8799.t65 464.166
R20812 a_n8300_8799.n112 a_n8300_8799.t87 464.166
R20813 a_n8300_8799.n108 a_n8300_8799.t107 464.166
R20814 a_n8300_8799.n113 a_n8300_8799.t108 464.166
R20815 a_n8300_8799.n114 a_n8300_8799.t76 464.166
R20816 a_n8300_8799.n107 a_n8300_8799.t94 464.166
R20817 a_n8300_8799.n115 a_n8300_8799.t106 464.166
R20818 a_n8300_8799.n106 a_n8300_8799.t74 464.166
R20819 a_n8300_8799.n116 a_n8300_8799.t75 464.166
R20820 a_n8300_8799.n121 a_n8300_8799.t119 464.166
R20821 a_n8300_8799.n120 a_n8300_8799.t71 464.166
R20822 a_n8300_8799.n123 a_n8300_8799.t93 464.166
R20823 a_n8300_8799.n119 a_n8300_8799.t116 464.166
R20824 a_n8300_8799.n124 a_n8300_8799.t118 464.166
R20825 a_n8300_8799.n125 a_n8300_8799.t83 464.166
R20826 a_n8300_8799.n118 a_n8300_8799.t103 464.166
R20827 a_n8300_8799.n126 a_n8300_8799.t115 464.166
R20828 a_n8300_8799.n117 a_n8300_8799.t79 464.166
R20829 a_n8300_8799.n127 a_n8300_8799.t80 464.166
R20830 a_n8300_8799.n133 a_n8300_8799.t67 464.166
R20831 a_n8300_8799.n132 a_n8300_8799.t81 464.166
R20832 a_n8300_8799.n135 a_n8300_8799.t54 464.166
R20833 a_n8300_8799.n131 a_n8300_8799.t90 464.166
R20834 a_n8300_8799.n136 a_n8300_8799.t78 464.166
R20835 a_n8300_8799.n137 a_n8300_8799.t102 464.166
R20836 a_n8300_8799.n130 a_n8300_8799.t72 464.166
R20837 a_n8300_8799.n138 a_n8300_8799.t109 464.166
R20838 a_n8300_8799.n129 a_n8300_8799.t58 464.166
R20839 a_n8300_8799.n139 a_n8300_8799.t48 464.166
R20840 a_n8300_8799.n42 a_n8300_8799.n41 75.3623
R20841 a_n8300_8799.n40 a_n8300_8799.n20 70.3058
R20842 a_n8300_8799.n20 a_n8300_8799.n39 70.1674
R20843 a_n8300_8799.n39 a_n8300_8799.n142 20.9683
R20844 a_n8300_8799.n38 a_n8300_8799.n21 75.0448
R20845 a_n8300_8799.n148 a_n8300_8799.n38 11.2134
R20846 a_n8300_8799.n37 a_n8300_8799.n21 80.4688
R20847 a_n8300_8799.n23 a_n8300_8799.n36 74.73
R20848 a_n8300_8799.n35 a_n8300_8799.n23 70.1674
R20849 a_n8300_8799.n151 a_n8300_8799.n35 20.9683
R20850 a_n8300_8799.n22 a_n8300_8799.n34 70.5844
R20851 a_n8300_8799.n51 a_n8300_8799.n50 75.3623
R20852 a_n8300_8799.n49 a_n8300_8799.n16 70.3058
R20853 a_n8300_8799.n16 a_n8300_8799.n48 70.1674
R20854 a_n8300_8799.n48 a_n8300_8799.n153 20.9683
R20855 a_n8300_8799.n47 a_n8300_8799.n17 75.0448
R20856 a_n8300_8799.n159 a_n8300_8799.n47 11.2134
R20857 a_n8300_8799.n46 a_n8300_8799.n17 80.4688
R20858 a_n8300_8799.n19 a_n8300_8799.n45 74.73
R20859 a_n8300_8799.n44 a_n8300_8799.n19 70.1674
R20860 a_n8300_8799.n162 a_n8300_8799.n44 20.9683
R20861 a_n8300_8799.n18 a_n8300_8799.n43 70.5844
R20862 a_n8300_8799.n60 a_n8300_8799.n59 75.3623
R20863 a_n8300_8799.n58 a_n8300_8799.n12 70.3058
R20864 a_n8300_8799.n12 a_n8300_8799.n57 70.1674
R20865 a_n8300_8799.n57 a_n8300_8799.n165 20.9683
R20866 a_n8300_8799.n56 a_n8300_8799.n13 75.0448
R20867 a_n8300_8799.n171 a_n8300_8799.n56 11.2134
R20868 a_n8300_8799.n55 a_n8300_8799.n13 80.4688
R20869 a_n8300_8799.n15 a_n8300_8799.n54 74.73
R20870 a_n8300_8799.n53 a_n8300_8799.n15 70.1674
R20871 a_n8300_8799.n174 a_n8300_8799.n53 20.9683
R20872 a_n8300_8799.n14 a_n8300_8799.n52 70.5844
R20873 a_n8300_8799.n8 a_n8300_8799.n69 70.5844
R20874 a_n8300_8799.n68 a_n8300_8799.n9 70.1674
R20875 a_n8300_8799.n68 a_n8300_8799.n106 20.9683
R20876 a_n8300_8799.n9 a_n8300_8799.n67 74.73
R20877 a_n8300_8799.n115 a_n8300_8799.n67 11.843
R20878 a_n8300_8799.n66 a_n8300_8799.n10 80.4688
R20879 a_n8300_8799.n66 a_n8300_8799.n107 0.365327
R20880 a_n8300_8799.n10 a_n8300_8799.n65 75.0448
R20881 a_n8300_8799.n64 a_n8300_8799.n11 70.1674
R20882 a_n8300_8799.n64 a_n8300_8799.n108 20.9683
R20883 a_n8300_8799.n11 a_n8300_8799.n63 70.3058
R20884 a_n8300_8799.n112 a_n8300_8799.n63 20.6913
R20885 a_n8300_8799.n62 a_n8300_8799.n61 75.3623
R20886 a_n8300_8799.n4 a_n8300_8799.n78 70.5844
R20887 a_n8300_8799.n77 a_n8300_8799.n5 70.1674
R20888 a_n8300_8799.n77 a_n8300_8799.n117 20.9683
R20889 a_n8300_8799.n5 a_n8300_8799.n76 74.73
R20890 a_n8300_8799.n126 a_n8300_8799.n76 11.843
R20891 a_n8300_8799.n75 a_n8300_8799.n6 80.4688
R20892 a_n8300_8799.n75 a_n8300_8799.n118 0.365327
R20893 a_n8300_8799.n6 a_n8300_8799.n74 75.0448
R20894 a_n8300_8799.n73 a_n8300_8799.n7 70.1674
R20895 a_n8300_8799.n73 a_n8300_8799.n119 20.9683
R20896 a_n8300_8799.n7 a_n8300_8799.n72 70.3058
R20897 a_n8300_8799.n123 a_n8300_8799.n72 20.6913
R20898 a_n8300_8799.n71 a_n8300_8799.n70 75.3623
R20899 a_n8300_8799.n0 a_n8300_8799.n87 70.5844
R20900 a_n8300_8799.n86 a_n8300_8799.n1 70.1674
R20901 a_n8300_8799.n86 a_n8300_8799.n129 20.9683
R20902 a_n8300_8799.n1 a_n8300_8799.n85 74.73
R20903 a_n8300_8799.n138 a_n8300_8799.n85 11.843
R20904 a_n8300_8799.n84 a_n8300_8799.n2 80.4688
R20905 a_n8300_8799.n84 a_n8300_8799.n130 0.365327
R20906 a_n8300_8799.n2 a_n8300_8799.n83 75.0448
R20907 a_n8300_8799.n82 a_n8300_8799.n3 70.1674
R20908 a_n8300_8799.n82 a_n8300_8799.n131 20.9683
R20909 a_n8300_8799.n3 a_n8300_8799.n81 70.3058
R20910 a_n8300_8799.n135 a_n8300_8799.n81 20.6913
R20911 a_n8300_8799.n80 a_n8300_8799.n79 75.3623
R20912 a_n8300_8799.n27 a_n8300_8799.n88 98.9633
R20913 a_n8300_8799.n184 a_n8300_8799.n32 98.9632
R20914 a_n8300_8799.n32 a_n8300_8799.n183 98.6055
R20915 a_n8300_8799.n32 a_n8300_8799.n182 98.6055
R20916 a_n8300_8799.n31 a_n8300_8799.n181 98.6055
R20917 a_n8300_8799.n31 a_n8300_8799.n180 98.6055
R20918 a_n8300_8799.n30 a_n8300_8799.n179 98.6055
R20919 a_n8300_8799.n29 a_n8300_8799.n93 98.6055
R20920 a_n8300_8799.n29 a_n8300_8799.n92 98.6055
R20921 a_n8300_8799.n28 a_n8300_8799.n91 98.6055
R20922 a_n8300_8799.n28 a_n8300_8799.n90 98.6055
R20923 a_n8300_8799.n27 a_n8300_8799.n89 98.6055
R20924 a_n8300_8799.n25 a_n8300_8799.n94 81.2902
R20925 a_n8300_8799.n33 a_n8300_8799.n100 81.2902
R20926 a_n8300_8799.n24 a_n8300_8799.n97 81.2902
R20927 a_n8300_8799.n26 a_n8300_8799.n103 80.9324
R20928 a_n8300_8799.n26 a_n8300_8799.n104 80.9324
R20929 a_n8300_8799.n25 a_n8300_8799.n105 80.9324
R20930 a_n8300_8799.n25 a_n8300_8799.n96 80.9324
R20931 a_n8300_8799.n25 a_n8300_8799.n95 80.9324
R20932 a_n8300_8799.n33 a_n8300_8799.n101 80.9324
R20933 a_n8300_8799.n24 a_n8300_8799.n102 80.9324
R20934 a_n8300_8799.n24 a_n8300_8799.n99 80.9324
R20935 a_n8300_8799.n24 a_n8300_8799.n98 80.9324
R20936 a_n8300_8799.n35 a_n8300_8799.n150 20.9683
R20937 a_n8300_8799.n149 a_n8300_8799.n148 48.2005
R20938 a_n8300_8799.n147 a_n8300_8799.n39 20.9683
R20939 a_n8300_8799.n144 a_n8300_8799.n143 48.2005
R20940 a_n8300_8799.n44 a_n8300_8799.n161 20.9683
R20941 a_n8300_8799.n160 a_n8300_8799.n159 48.2005
R20942 a_n8300_8799.n158 a_n8300_8799.n48 20.9683
R20943 a_n8300_8799.n155 a_n8300_8799.n154 48.2005
R20944 a_n8300_8799.n53 a_n8300_8799.n173 20.9683
R20945 a_n8300_8799.n172 a_n8300_8799.n171 48.2005
R20946 a_n8300_8799.n170 a_n8300_8799.n57 20.9683
R20947 a_n8300_8799.n167 a_n8300_8799.n166 48.2005
R20948 a_n8300_8799.n110 a_n8300_8799.n109 48.2005
R20949 a_n8300_8799.n113 a_n8300_8799.n64 20.9683
R20950 a_n8300_8799.n114 a_n8300_8799.n107 48.2005
R20951 a_n8300_8799.n116 a_n8300_8799.n68 20.9683
R20952 a_n8300_8799.n121 a_n8300_8799.n120 48.2005
R20953 a_n8300_8799.n124 a_n8300_8799.n73 20.9683
R20954 a_n8300_8799.n125 a_n8300_8799.n118 48.2005
R20955 a_n8300_8799.n127 a_n8300_8799.n77 20.9683
R20956 a_n8300_8799.n133 a_n8300_8799.n132 48.2005
R20957 a_n8300_8799.n136 a_n8300_8799.n82 20.9683
R20958 a_n8300_8799.n137 a_n8300_8799.n130 48.2005
R20959 a_n8300_8799.n139 a_n8300_8799.n86 20.9683
R20960 a_n8300_8799.n37 a_n8300_8799.n141 47.835
R20961 a_n8300_8799.n40 a_n8300_8799.n146 20.6913
R20962 a_n8300_8799.n46 a_n8300_8799.n152 47.835
R20963 a_n8300_8799.n49 a_n8300_8799.n157 20.6913
R20964 a_n8300_8799.n55 a_n8300_8799.n164 47.835
R20965 a_n8300_8799.n58 a_n8300_8799.n169 20.6913
R20966 a_n8300_8799.n108 a_n8300_8799.n63 21.4216
R20967 a_n8300_8799.n119 a_n8300_8799.n72 21.4216
R20968 a_n8300_8799.n131 a_n8300_8799.n81 21.4216
R20969 a_n8300_8799.t92 a_n8300_8799.n69 484.3
R20970 a_n8300_8799.t101 a_n8300_8799.n78 484.3
R20971 a_n8300_8799.t84 a_n8300_8799.n87 484.3
R20972 a_n8300_8799.n62 a_n8300_8799.n111 45.0871
R20973 a_n8300_8799.n71 a_n8300_8799.n122 45.0871
R20974 a_n8300_8799.n80 a_n8300_8799.n134 45.0871
R20975 a_n8300_8799.n42 a_n8300_8799.n145 45.0871
R20976 a_n8300_8799.n51 a_n8300_8799.n156 45.0871
R20977 a_n8300_8799.n60 a_n8300_8799.n168 45.0871
R20978 a_n8300_8799.n30 a_n8300_8799.n178 33.8967
R20979 a_n8300_8799.n26 a_n8300_8799.n24 32.5134
R20980 a_n8300_8799.n36 a_n8300_8799.n141 11.843
R20981 a_n8300_8799.n146 a_n8300_8799.n41 36.139
R20982 a_n8300_8799.n45 a_n8300_8799.n152 11.843
R20983 a_n8300_8799.n157 a_n8300_8799.n50 36.139
R20984 a_n8300_8799.n54 a_n8300_8799.n164 11.843
R20985 a_n8300_8799.n169 a_n8300_8799.n59 36.139
R20986 a_n8300_8799.n112 a_n8300_8799.n61 36.139
R20987 a_n8300_8799.n106 a_n8300_8799.n67 34.4824
R20988 a_n8300_8799.n123 a_n8300_8799.n70 36.139
R20989 a_n8300_8799.n117 a_n8300_8799.n76 34.4824
R20990 a_n8300_8799.n135 a_n8300_8799.n79 36.139
R20991 a_n8300_8799.n129 a_n8300_8799.n85 34.4824
R20992 a_n8300_8799.n38 a_n8300_8799.n142 35.3134
R20993 a_n8300_8799.n47 a_n8300_8799.n153 35.3134
R20994 a_n8300_8799.n56 a_n8300_8799.n165 35.3134
R20995 a_n8300_8799.n65 a_n8300_8799.n113 35.3134
R20996 a_n8300_8799.n114 a_n8300_8799.n65 11.2134
R20997 a_n8300_8799.n74 a_n8300_8799.n124 35.3134
R20998 a_n8300_8799.n125 a_n8300_8799.n74 11.2134
R20999 a_n8300_8799.n83 a_n8300_8799.n136 35.3134
R21000 a_n8300_8799.n137 a_n8300_8799.n83 11.2134
R21001 a_n8300_8799.n150 a_n8300_8799.n36 34.4824
R21002 a_n8300_8799.n41 a_n8300_8799.n143 10.5784
R21003 a_n8300_8799.n161 a_n8300_8799.n45 34.4824
R21004 a_n8300_8799.n50 a_n8300_8799.n154 10.5784
R21005 a_n8300_8799.n173 a_n8300_8799.n54 34.4824
R21006 a_n8300_8799.n59 a_n8300_8799.n166 10.5784
R21007 a_n8300_8799.n61 a_n8300_8799.n109 10.5784
R21008 a_n8300_8799.n70 a_n8300_8799.n120 10.5784
R21009 a_n8300_8799.n79 a_n8300_8799.n132 10.5784
R21010 a_n8300_8799.n178 a_n8300_8799.n29 20.9925
R21011 a_n8300_8799.n145 a_n8300_8799.n144 14.1472
R21012 a_n8300_8799.n156 a_n8300_8799.n155 14.1472
R21013 a_n8300_8799.n168 a_n8300_8799.n167 14.1472
R21014 a_n8300_8799.n111 a_n8300_8799.n110 14.1472
R21015 a_n8300_8799.n122 a_n8300_8799.n121 14.1472
R21016 a_n8300_8799.n134 a_n8300_8799.n133 14.1472
R21017 a_n8300_8799.n177 a_n8300_8799.n25 12.3339
R21018 a_n8300_8799.n178 a_n8300_8799.n177 11.4887
R21019 a_n8300_8799.n163 a_n8300_8799.n22 9.01755
R21020 a_n8300_8799.n128 a_n8300_8799.n8 9.01755
R21021 a_n8300_8799.n176 a_n8300_8799.n140 7.1766
R21022 a_n8300_8799.n176 a_n8300_8799.n175 6.83037
R21023 a_n8300_8799.n163 a_n8300_8799.n18 4.90959
R21024 a_n8300_8799.n175 a_n8300_8799.n14 4.90959
R21025 a_n8300_8799.n128 a_n8300_8799.n4 4.90959
R21026 a_n8300_8799.n140 a_n8300_8799.n0 4.90959
R21027 a_n8300_8799.n175 a_n8300_8799.n163 4.10845
R21028 a_n8300_8799.n140 a_n8300_8799.n128 4.10845
R21029 a_n8300_8799.n183 a_n8300_8799.t26 3.61217
R21030 a_n8300_8799.n183 a_n8300_8799.t40 3.61217
R21031 a_n8300_8799.n182 a_n8300_8799.t31 3.61217
R21032 a_n8300_8799.n182 a_n8300_8799.t36 3.61217
R21033 a_n8300_8799.n181 a_n8300_8799.t23 3.61217
R21034 a_n8300_8799.n181 a_n8300_8799.t35 3.61217
R21035 a_n8300_8799.n180 a_n8300_8799.t34 3.61217
R21036 a_n8300_8799.n180 a_n8300_8799.t30 3.61217
R21037 a_n8300_8799.n179 a_n8300_8799.t42 3.61217
R21038 a_n8300_8799.n179 a_n8300_8799.t22 3.61217
R21039 a_n8300_8799.n93 a_n8300_8799.t37 3.61217
R21040 a_n8300_8799.n93 a_n8300_8799.t39 3.61217
R21041 a_n8300_8799.n92 a_n8300_8799.t38 3.61217
R21042 a_n8300_8799.n92 a_n8300_8799.t25 3.61217
R21043 a_n8300_8799.n91 a_n8300_8799.t33 3.61217
R21044 a_n8300_8799.n91 a_n8300_8799.t29 3.61217
R21045 a_n8300_8799.n90 a_n8300_8799.t32 3.61217
R21046 a_n8300_8799.n90 a_n8300_8799.t27 3.61217
R21047 a_n8300_8799.n89 a_n8300_8799.t24 3.61217
R21048 a_n8300_8799.n89 a_n8300_8799.t41 3.61217
R21049 a_n8300_8799.n88 a_n8300_8799.t20 3.61217
R21050 a_n8300_8799.n88 a_n8300_8799.t28 3.61217
R21051 a_n8300_8799.t19 a_n8300_8799.n184 3.61217
R21052 a_n8300_8799.n184 a_n8300_8799.t21 3.61217
R21053 a_n8300_8799.n177 a_n8300_8799.n176 3.4105
R21054 a_n8300_8799.n103 a_n8300_8799.t15 2.82907
R21055 a_n8300_8799.n103 a_n8300_8799.t1 2.82907
R21056 a_n8300_8799.n104 a_n8300_8799.t0 2.82907
R21057 a_n8300_8799.n104 a_n8300_8799.t47 2.82907
R21058 a_n8300_8799.n105 a_n8300_8799.t8 2.82907
R21059 a_n8300_8799.n105 a_n8300_8799.t44 2.82907
R21060 a_n8300_8799.n96 a_n8300_8799.t16 2.82907
R21061 a_n8300_8799.n96 a_n8300_8799.t10 2.82907
R21062 a_n8300_8799.n95 a_n8300_8799.t5 2.82907
R21063 a_n8300_8799.n95 a_n8300_8799.t18 2.82907
R21064 a_n8300_8799.n94 a_n8300_8799.t13 2.82907
R21065 a_n8300_8799.n94 a_n8300_8799.t2 2.82907
R21066 a_n8300_8799.n100 a_n8300_8799.t46 2.82907
R21067 a_n8300_8799.n100 a_n8300_8799.t9 2.82907
R21068 a_n8300_8799.n101 a_n8300_8799.t11 2.82907
R21069 a_n8300_8799.n101 a_n8300_8799.t17 2.82907
R21070 a_n8300_8799.n102 a_n8300_8799.t45 2.82907
R21071 a_n8300_8799.n102 a_n8300_8799.t14 2.82907
R21072 a_n8300_8799.n99 a_n8300_8799.t4 2.82907
R21073 a_n8300_8799.n99 a_n8300_8799.t12 2.82907
R21074 a_n8300_8799.n98 a_n8300_8799.t43 2.82907
R21075 a_n8300_8799.n98 a_n8300_8799.t3 2.82907
R21076 a_n8300_8799.n97 a_n8300_8799.t7 2.82907
R21077 a_n8300_8799.n97 a_n8300_8799.t6 2.82907
R21078 a_n8300_8799.n34 a_n8300_8799.n151 22.3251
R21079 a_n8300_8799.n43 a_n8300_8799.n162 22.3251
R21080 a_n8300_8799.n52 a_n8300_8799.n174 22.3251
R21081 a_n8300_8799.n69 a_n8300_8799.n116 22.3251
R21082 a_n8300_8799.n78 a_n8300_8799.n127 22.3251
R21083 a_n8300_8799.n87 a_n8300_8799.n139 22.3251
R21084 a_n8300_8799.n37 a_n8300_8799.n149 0.365327
R21085 a_n8300_8799.n147 a_n8300_8799.n40 21.4216
R21086 a_n8300_8799.n46 a_n8300_8799.n160 0.365327
R21087 a_n8300_8799.n158 a_n8300_8799.n49 21.4216
R21088 a_n8300_8799.n55 a_n8300_8799.n172 0.365327
R21089 a_n8300_8799.n170 a_n8300_8799.n58 21.4216
R21090 a_n8300_8799.n115 a_n8300_8799.n66 47.835
R21091 a_n8300_8799.n126 a_n8300_8799.n75 47.835
R21092 a_n8300_8799.n138 a_n8300_8799.n84 47.835
R21093 a_n8300_8799.n25 a_n8300_8799.n26 1.43153
R21094 a_n8300_8799.n24 a_n8300_8799.n33 1.07378
R21095 a_n8300_8799.n23 a_n8300_8799.n21 0.758076
R21096 a_n8300_8799.n21 a_n8300_8799.n20 0.758076
R21097 a_n8300_8799.n42 a_n8300_8799.n20 0.758076
R21098 a_n8300_8799.n19 a_n8300_8799.n17 0.758076
R21099 a_n8300_8799.n17 a_n8300_8799.n16 0.758076
R21100 a_n8300_8799.n51 a_n8300_8799.n16 0.758076
R21101 a_n8300_8799.n15 a_n8300_8799.n13 0.758076
R21102 a_n8300_8799.n13 a_n8300_8799.n12 0.758076
R21103 a_n8300_8799.n60 a_n8300_8799.n12 0.758076
R21104 a_n8300_8799.n11 a_n8300_8799.n10 0.758076
R21105 a_n8300_8799.n10 a_n8300_8799.n9 0.758076
R21106 a_n8300_8799.n9 a_n8300_8799.n8 0.758076
R21107 a_n8300_8799.n7 a_n8300_8799.n6 0.758076
R21108 a_n8300_8799.n6 a_n8300_8799.n5 0.758076
R21109 a_n8300_8799.n5 a_n8300_8799.n4 0.758076
R21110 a_n8300_8799.n3 a_n8300_8799.n2 0.758076
R21111 a_n8300_8799.n2 a_n8300_8799.n1 0.758076
R21112 a_n8300_8799.n1 a_n8300_8799.n0 0.758076
R21113 a_n8300_8799.n32 a_n8300_8799.n31 0.716017
R21114 a_n8300_8799.n31 a_n8300_8799.n30 0.716017
R21115 a_n8300_8799.n29 a_n8300_8799.n28 0.716017
R21116 a_n8300_8799.n28 a_n8300_8799.n27 0.716017
R21117 a_n8300_8799.n80 a_n8300_8799.n3 0.568682
R21118 a_n8300_8799.n71 a_n8300_8799.n7 0.568682
R21119 a_n8300_8799.n62 a_n8300_8799.n11 0.568682
R21120 a_n8300_8799.n15 a_n8300_8799.n14 0.568682
R21121 a_n8300_8799.n19 a_n8300_8799.n18 0.568682
R21122 a_n8300_8799.n23 a_n8300_8799.n22 0.568682
R21123 CSoutput.n19 CSoutput.t160 184.661
R21124 CSoutput.n78 CSoutput.n77 165.8
R21125 CSoutput.n76 CSoutput.n0 165.8
R21126 CSoutput.n75 CSoutput.n74 165.8
R21127 CSoutput.n73 CSoutput.n72 165.8
R21128 CSoutput.n71 CSoutput.n2 165.8
R21129 CSoutput.n69 CSoutput.n68 165.8
R21130 CSoutput.n67 CSoutput.n3 165.8
R21131 CSoutput.n66 CSoutput.n65 165.8
R21132 CSoutput.n63 CSoutput.n4 165.8
R21133 CSoutput.n61 CSoutput.n60 165.8
R21134 CSoutput.n59 CSoutput.n5 165.8
R21135 CSoutput.n58 CSoutput.n57 165.8
R21136 CSoutput.n55 CSoutput.n6 165.8
R21137 CSoutput.n54 CSoutput.n53 165.8
R21138 CSoutput.n52 CSoutput.n51 165.8
R21139 CSoutput.n50 CSoutput.n8 165.8
R21140 CSoutput.n48 CSoutput.n47 165.8
R21141 CSoutput.n46 CSoutput.n9 165.8
R21142 CSoutput.n45 CSoutput.n44 165.8
R21143 CSoutput.n42 CSoutput.n10 165.8
R21144 CSoutput.n41 CSoutput.n40 165.8
R21145 CSoutput.n39 CSoutput.n38 165.8
R21146 CSoutput.n37 CSoutput.n12 165.8
R21147 CSoutput.n35 CSoutput.n34 165.8
R21148 CSoutput.n33 CSoutput.n13 165.8
R21149 CSoutput.n32 CSoutput.n31 165.8
R21150 CSoutput.n29 CSoutput.n14 165.8
R21151 CSoutput.n28 CSoutput.n27 165.8
R21152 CSoutput.n26 CSoutput.n25 165.8
R21153 CSoutput.n24 CSoutput.n16 165.8
R21154 CSoutput.n22 CSoutput.n21 165.8
R21155 CSoutput.n20 CSoutput.n17 165.8
R21156 CSoutput.n77 CSoutput.t164 162.194
R21157 CSoutput.n18 CSoutput.t150 120.501
R21158 CSoutput.n23 CSoutput.t152 120.501
R21159 CSoutput.n15 CSoutput.t165 120.501
R21160 CSoutput.n30 CSoutput.t153 120.501
R21161 CSoutput.n36 CSoutput.t156 120.501
R21162 CSoutput.n11 CSoutput.t148 120.501
R21163 CSoutput.n43 CSoutput.t161 120.501
R21164 CSoutput.n49 CSoutput.t157 120.501
R21165 CSoutput.n7 CSoutput.t151 120.501
R21166 CSoutput.n56 CSoutput.t147 120.501
R21167 CSoutput.n62 CSoutput.t158 120.501
R21168 CSoutput.n64 CSoutput.t159 120.501
R21169 CSoutput.n70 CSoutput.t149 120.501
R21170 CSoutput.n1 CSoutput.t145 120.501
R21171 CSoutput.n290 CSoutput.n288 103.469
R21172 CSoutput.n278 CSoutput.n276 103.469
R21173 CSoutput.n267 CSoutput.n265 103.469
R21174 CSoutput.n104 CSoutput.n102 103.469
R21175 CSoutput.n92 CSoutput.n90 103.469
R21176 CSoutput.n81 CSoutput.n79 103.469
R21177 CSoutput.n296 CSoutput.n295 103.111
R21178 CSoutput.n294 CSoutput.n293 103.111
R21179 CSoutput.n292 CSoutput.n291 103.111
R21180 CSoutput.n290 CSoutput.n289 103.111
R21181 CSoutput.n286 CSoutput.n285 103.111
R21182 CSoutput.n284 CSoutput.n283 103.111
R21183 CSoutput.n282 CSoutput.n281 103.111
R21184 CSoutput.n280 CSoutput.n279 103.111
R21185 CSoutput.n278 CSoutput.n277 103.111
R21186 CSoutput.n275 CSoutput.n274 103.111
R21187 CSoutput.n273 CSoutput.n272 103.111
R21188 CSoutput.n271 CSoutput.n270 103.111
R21189 CSoutput.n269 CSoutput.n268 103.111
R21190 CSoutput.n267 CSoutput.n266 103.111
R21191 CSoutput.n104 CSoutput.n103 103.111
R21192 CSoutput.n106 CSoutput.n105 103.111
R21193 CSoutput.n108 CSoutput.n107 103.111
R21194 CSoutput.n110 CSoutput.n109 103.111
R21195 CSoutput.n112 CSoutput.n111 103.111
R21196 CSoutput.n92 CSoutput.n91 103.111
R21197 CSoutput.n94 CSoutput.n93 103.111
R21198 CSoutput.n96 CSoutput.n95 103.111
R21199 CSoutput.n98 CSoutput.n97 103.111
R21200 CSoutput.n100 CSoutput.n99 103.111
R21201 CSoutput.n81 CSoutput.n80 103.111
R21202 CSoutput.n83 CSoutput.n82 103.111
R21203 CSoutput.n85 CSoutput.n84 103.111
R21204 CSoutput.n87 CSoutput.n86 103.111
R21205 CSoutput.n89 CSoutput.n88 103.111
R21206 CSoutput.n298 CSoutput.n297 103.111
R21207 CSoutput.n326 CSoutput.n324 81.5057
R21208 CSoutput.n314 CSoutput.n312 81.5057
R21209 CSoutput.n303 CSoutput.n301 81.5057
R21210 CSoutput.n362 CSoutput.n360 81.5057
R21211 CSoutput.n350 CSoutput.n348 81.5057
R21212 CSoutput.n339 CSoutput.n337 81.5057
R21213 CSoutput.n334 CSoutput.n333 80.9324
R21214 CSoutput.n332 CSoutput.n331 80.9324
R21215 CSoutput.n330 CSoutput.n329 80.9324
R21216 CSoutput.n328 CSoutput.n327 80.9324
R21217 CSoutput.n326 CSoutput.n325 80.9324
R21218 CSoutput.n322 CSoutput.n321 80.9324
R21219 CSoutput.n320 CSoutput.n319 80.9324
R21220 CSoutput.n318 CSoutput.n317 80.9324
R21221 CSoutput.n316 CSoutput.n315 80.9324
R21222 CSoutput.n314 CSoutput.n313 80.9324
R21223 CSoutput.n311 CSoutput.n310 80.9324
R21224 CSoutput.n309 CSoutput.n308 80.9324
R21225 CSoutput.n307 CSoutput.n306 80.9324
R21226 CSoutput.n305 CSoutput.n304 80.9324
R21227 CSoutput.n303 CSoutput.n302 80.9324
R21228 CSoutput.n362 CSoutput.n361 80.9324
R21229 CSoutput.n364 CSoutput.n363 80.9324
R21230 CSoutput.n366 CSoutput.n365 80.9324
R21231 CSoutput.n368 CSoutput.n367 80.9324
R21232 CSoutput.n370 CSoutput.n369 80.9324
R21233 CSoutput.n350 CSoutput.n349 80.9324
R21234 CSoutput.n352 CSoutput.n351 80.9324
R21235 CSoutput.n354 CSoutput.n353 80.9324
R21236 CSoutput.n356 CSoutput.n355 80.9324
R21237 CSoutput.n358 CSoutput.n357 80.9324
R21238 CSoutput.n339 CSoutput.n338 80.9324
R21239 CSoutput.n341 CSoutput.n340 80.9324
R21240 CSoutput.n343 CSoutput.n342 80.9324
R21241 CSoutput.n345 CSoutput.n344 80.9324
R21242 CSoutput.n347 CSoutput.n346 80.9324
R21243 CSoutput.n25 CSoutput.n24 48.1486
R21244 CSoutput.n69 CSoutput.n3 48.1486
R21245 CSoutput.n38 CSoutput.n37 48.1486
R21246 CSoutput.n42 CSoutput.n41 48.1486
R21247 CSoutput.n51 CSoutput.n50 48.1486
R21248 CSoutput.n55 CSoutput.n54 48.1486
R21249 CSoutput.n22 CSoutput.n17 46.462
R21250 CSoutput.n72 CSoutput.n71 46.462
R21251 CSoutput.n20 CSoutput.n19 44.9055
R21252 CSoutput.n29 CSoutput.n28 43.7635
R21253 CSoutput.n65 CSoutput.n63 43.7635
R21254 CSoutput.n35 CSoutput.n13 41.7396
R21255 CSoutput.n57 CSoutput.n5 41.7396
R21256 CSoutput.n44 CSoutput.n9 37.0171
R21257 CSoutput.n48 CSoutput.n9 37.0171
R21258 CSoutput.n76 CSoutput.n75 34.9932
R21259 CSoutput.n31 CSoutput.n13 32.2947
R21260 CSoutput.n61 CSoutput.n5 32.2947
R21261 CSoutput.n30 CSoutput.n29 29.6014
R21262 CSoutput.n63 CSoutput.n62 29.6014
R21263 CSoutput.n19 CSoutput.n18 28.4085
R21264 CSoutput.n18 CSoutput.n17 25.1176
R21265 CSoutput.n72 CSoutput.n1 25.1176
R21266 CSoutput.n43 CSoutput.n42 22.0922
R21267 CSoutput.n50 CSoutput.n49 22.0922
R21268 CSoutput.n77 CSoutput.n76 21.8586
R21269 CSoutput.n37 CSoutput.n36 18.9681
R21270 CSoutput.n56 CSoutput.n55 18.9681
R21271 CSoutput.n25 CSoutput.n15 17.6292
R21272 CSoutput.n64 CSoutput.n3 17.6292
R21273 CSoutput.n24 CSoutput.n23 15.844
R21274 CSoutput.n70 CSoutput.n69 15.844
R21275 CSoutput.n38 CSoutput.n11 14.5051
R21276 CSoutput.n54 CSoutput.n7 14.5051
R21277 CSoutput.n373 CSoutput.n78 11.4982
R21278 CSoutput.n41 CSoutput.n11 11.3811
R21279 CSoutput.n51 CSoutput.n7 11.3811
R21280 CSoutput.n23 CSoutput.n22 10.0422
R21281 CSoutput.n71 CSoutput.n70 10.0422
R21282 CSoutput.n287 CSoutput.n275 9.25285
R21283 CSoutput.n101 CSoutput.n89 9.25285
R21284 CSoutput.n323 CSoutput.n311 8.98182
R21285 CSoutput.n359 CSoutput.n347 8.98182
R21286 CSoutput.n336 CSoutput.n300 8.65726
R21287 CSoutput.n28 CSoutput.n15 8.25698
R21288 CSoutput.n65 CSoutput.n64 8.25698
R21289 CSoutput.n300 CSoutput.n299 7.12641
R21290 CSoutput.n114 CSoutput.n113 7.12641
R21291 CSoutput.n36 CSoutput.n35 6.91809
R21292 CSoutput.n57 CSoutput.n56 6.91809
R21293 CSoutput.n336 CSoutput.n335 6.02792
R21294 CSoutput.n372 CSoutput.n371 6.02792
R21295 CSoutput.n335 CSoutput.n334 5.25266
R21296 CSoutput.n323 CSoutput.n322 5.25266
R21297 CSoutput.n371 CSoutput.n370 5.25266
R21298 CSoutput.n359 CSoutput.n358 5.25266
R21299 CSoutput.n299 CSoutput.n298 5.1449
R21300 CSoutput.n287 CSoutput.n286 5.1449
R21301 CSoutput.n113 CSoutput.n112 5.1449
R21302 CSoutput.n101 CSoutput.n100 5.1449
R21303 CSoutput.n373 CSoutput.n114 5.06482
R21304 CSoutput.n205 CSoutput.n158 4.5005
R21305 CSoutput.n174 CSoutput.n158 4.5005
R21306 CSoutput.n169 CSoutput.n153 4.5005
R21307 CSoutput.n169 CSoutput.n155 4.5005
R21308 CSoutput.n169 CSoutput.n152 4.5005
R21309 CSoutput.n169 CSoutput.n156 4.5005
R21310 CSoutput.n169 CSoutput.n151 4.5005
R21311 CSoutput.n169 CSoutput.t162 4.5005
R21312 CSoutput.n169 CSoutput.n150 4.5005
R21313 CSoutput.n169 CSoutput.n157 4.5005
R21314 CSoutput.n169 CSoutput.n158 4.5005
R21315 CSoutput.n167 CSoutput.n153 4.5005
R21316 CSoutput.n167 CSoutput.n155 4.5005
R21317 CSoutput.n167 CSoutput.n152 4.5005
R21318 CSoutput.n167 CSoutput.n156 4.5005
R21319 CSoutput.n167 CSoutput.n151 4.5005
R21320 CSoutput.n167 CSoutput.t162 4.5005
R21321 CSoutput.n167 CSoutput.n150 4.5005
R21322 CSoutput.n167 CSoutput.n157 4.5005
R21323 CSoutput.n167 CSoutput.n158 4.5005
R21324 CSoutput.n166 CSoutput.n153 4.5005
R21325 CSoutput.n166 CSoutput.n155 4.5005
R21326 CSoutput.n166 CSoutput.n152 4.5005
R21327 CSoutput.n166 CSoutput.n156 4.5005
R21328 CSoutput.n166 CSoutput.n151 4.5005
R21329 CSoutput.n166 CSoutput.t162 4.5005
R21330 CSoutput.n166 CSoutput.n150 4.5005
R21331 CSoutput.n166 CSoutput.n157 4.5005
R21332 CSoutput.n166 CSoutput.n158 4.5005
R21333 CSoutput.n251 CSoutput.n153 4.5005
R21334 CSoutput.n251 CSoutput.n155 4.5005
R21335 CSoutput.n251 CSoutput.n152 4.5005
R21336 CSoutput.n251 CSoutput.n156 4.5005
R21337 CSoutput.n251 CSoutput.n151 4.5005
R21338 CSoutput.n251 CSoutput.t162 4.5005
R21339 CSoutput.n251 CSoutput.n150 4.5005
R21340 CSoutput.n251 CSoutput.n157 4.5005
R21341 CSoutput.n251 CSoutput.n158 4.5005
R21342 CSoutput.n249 CSoutput.n153 4.5005
R21343 CSoutput.n249 CSoutput.n155 4.5005
R21344 CSoutput.n249 CSoutput.n152 4.5005
R21345 CSoutput.n249 CSoutput.n156 4.5005
R21346 CSoutput.n249 CSoutput.n151 4.5005
R21347 CSoutput.n249 CSoutput.t162 4.5005
R21348 CSoutput.n249 CSoutput.n150 4.5005
R21349 CSoutput.n249 CSoutput.n157 4.5005
R21350 CSoutput.n247 CSoutput.n153 4.5005
R21351 CSoutput.n247 CSoutput.n155 4.5005
R21352 CSoutput.n247 CSoutput.n152 4.5005
R21353 CSoutput.n247 CSoutput.n156 4.5005
R21354 CSoutput.n247 CSoutput.n151 4.5005
R21355 CSoutput.n247 CSoutput.t162 4.5005
R21356 CSoutput.n247 CSoutput.n150 4.5005
R21357 CSoutput.n247 CSoutput.n157 4.5005
R21358 CSoutput.n177 CSoutput.n153 4.5005
R21359 CSoutput.n177 CSoutput.n155 4.5005
R21360 CSoutput.n177 CSoutput.n152 4.5005
R21361 CSoutput.n177 CSoutput.n156 4.5005
R21362 CSoutput.n177 CSoutput.n151 4.5005
R21363 CSoutput.n177 CSoutput.t162 4.5005
R21364 CSoutput.n177 CSoutput.n150 4.5005
R21365 CSoutput.n177 CSoutput.n157 4.5005
R21366 CSoutput.n177 CSoutput.n158 4.5005
R21367 CSoutput.n176 CSoutput.n153 4.5005
R21368 CSoutput.n176 CSoutput.n155 4.5005
R21369 CSoutput.n176 CSoutput.n152 4.5005
R21370 CSoutput.n176 CSoutput.n156 4.5005
R21371 CSoutput.n176 CSoutput.n151 4.5005
R21372 CSoutput.n176 CSoutput.t162 4.5005
R21373 CSoutput.n176 CSoutput.n150 4.5005
R21374 CSoutput.n176 CSoutput.n157 4.5005
R21375 CSoutput.n176 CSoutput.n158 4.5005
R21376 CSoutput.n180 CSoutput.n153 4.5005
R21377 CSoutput.n180 CSoutput.n155 4.5005
R21378 CSoutput.n180 CSoutput.n152 4.5005
R21379 CSoutput.n180 CSoutput.n156 4.5005
R21380 CSoutput.n180 CSoutput.n151 4.5005
R21381 CSoutput.n180 CSoutput.t162 4.5005
R21382 CSoutput.n180 CSoutput.n150 4.5005
R21383 CSoutput.n180 CSoutput.n157 4.5005
R21384 CSoutput.n180 CSoutput.n158 4.5005
R21385 CSoutput.n179 CSoutput.n153 4.5005
R21386 CSoutput.n179 CSoutput.n155 4.5005
R21387 CSoutput.n179 CSoutput.n152 4.5005
R21388 CSoutput.n179 CSoutput.n156 4.5005
R21389 CSoutput.n179 CSoutput.n151 4.5005
R21390 CSoutput.n179 CSoutput.t162 4.5005
R21391 CSoutput.n179 CSoutput.n150 4.5005
R21392 CSoutput.n179 CSoutput.n157 4.5005
R21393 CSoutput.n179 CSoutput.n158 4.5005
R21394 CSoutput.n162 CSoutput.n153 4.5005
R21395 CSoutput.n162 CSoutput.n155 4.5005
R21396 CSoutput.n162 CSoutput.n152 4.5005
R21397 CSoutput.n162 CSoutput.n156 4.5005
R21398 CSoutput.n162 CSoutput.n151 4.5005
R21399 CSoutput.n162 CSoutput.t162 4.5005
R21400 CSoutput.n162 CSoutput.n150 4.5005
R21401 CSoutput.n162 CSoutput.n157 4.5005
R21402 CSoutput.n162 CSoutput.n158 4.5005
R21403 CSoutput.n254 CSoutput.n153 4.5005
R21404 CSoutput.n254 CSoutput.n155 4.5005
R21405 CSoutput.n254 CSoutput.n152 4.5005
R21406 CSoutput.n254 CSoutput.n156 4.5005
R21407 CSoutput.n254 CSoutput.n151 4.5005
R21408 CSoutput.n254 CSoutput.t162 4.5005
R21409 CSoutput.n254 CSoutput.n150 4.5005
R21410 CSoutput.n254 CSoutput.n157 4.5005
R21411 CSoutput.n254 CSoutput.n158 4.5005
R21412 CSoutput.n241 CSoutput.n212 4.5005
R21413 CSoutput.n241 CSoutput.n218 4.5005
R21414 CSoutput.n199 CSoutput.n188 4.5005
R21415 CSoutput.n199 CSoutput.n190 4.5005
R21416 CSoutput.n199 CSoutput.n187 4.5005
R21417 CSoutput.n199 CSoutput.n191 4.5005
R21418 CSoutput.n199 CSoutput.n186 4.5005
R21419 CSoutput.n199 CSoutput.t155 4.5005
R21420 CSoutput.n199 CSoutput.n185 4.5005
R21421 CSoutput.n199 CSoutput.n192 4.5005
R21422 CSoutput.n241 CSoutput.n199 4.5005
R21423 CSoutput.n220 CSoutput.n188 4.5005
R21424 CSoutput.n220 CSoutput.n190 4.5005
R21425 CSoutput.n220 CSoutput.n187 4.5005
R21426 CSoutput.n220 CSoutput.n191 4.5005
R21427 CSoutput.n220 CSoutput.n186 4.5005
R21428 CSoutput.n220 CSoutput.t155 4.5005
R21429 CSoutput.n220 CSoutput.n185 4.5005
R21430 CSoutput.n220 CSoutput.n192 4.5005
R21431 CSoutput.n241 CSoutput.n220 4.5005
R21432 CSoutput.n198 CSoutput.n188 4.5005
R21433 CSoutput.n198 CSoutput.n190 4.5005
R21434 CSoutput.n198 CSoutput.n187 4.5005
R21435 CSoutput.n198 CSoutput.n191 4.5005
R21436 CSoutput.n198 CSoutput.n186 4.5005
R21437 CSoutput.n198 CSoutput.t155 4.5005
R21438 CSoutput.n198 CSoutput.n185 4.5005
R21439 CSoutput.n198 CSoutput.n192 4.5005
R21440 CSoutput.n241 CSoutput.n198 4.5005
R21441 CSoutput.n222 CSoutput.n188 4.5005
R21442 CSoutput.n222 CSoutput.n190 4.5005
R21443 CSoutput.n222 CSoutput.n187 4.5005
R21444 CSoutput.n222 CSoutput.n191 4.5005
R21445 CSoutput.n222 CSoutput.n186 4.5005
R21446 CSoutput.n222 CSoutput.t155 4.5005
R21447 CSoutput.n222 CSoutput.n185 4.5005
R21448 CSoutput.n222 CSoutput.n192 4.5005
R21449 CSoutput.n241 CSoutput.n222 4.5005
R21450 CSoutput.n188 CSoutput.n183 4.5005
R21451 CSoutput.n190 CSoutput.n183 4.5005
R21452 CSoutput.n187 CSoutput.n183 4.5005
R21453 CSoutput.n191 CSoutput.n183 4.5005
R21454 CSoutput.n186 CSoutput.n183 4.5005
R21455 CSoutput.t155 CSoutput.n183 4.5005
R21456 CSoutput.n185 CSoutput.n183 4.5005
R21457 CSoutput.n192 CSoutput.n183 4.5005
R21458 CSoutput.n244 CSoutput.n188 4.5005
R21459 CSoutput.n244 CSoutput.n190 4.5005
R21460 CSoutput.n244 CSoutput.n187 4.5005
R21461 CSoutput.n244 CSoutput.n191 4.5005
R21462 CSoutput.n244 CSoutput.n186 4.5005
R21463 CSoutput.n244 CSoutput.t155 4.5005
R21464 CSoutput.n244 CSoutput.n185 4.5005
R21465 CSoutput.n244 CSoutput.n192 4.5005
R21466 CSoutput.n242 CSoutput.n188 4.5005
R21467 CSoutput.n242 CSoutput.n190 4.5005
R21468 CSoutput.n242 CSoutput.n187 4.5005
R21469 CSoutput.n242 CSoutput.n191 4.5005
R21470 CSoutput.n242 CSoutput.n186 4.5005
R21471 CSoutput.n242 CSoutput.t155 4.5005
R21472 CSoutput.n242 CSoutput.n185 4.5005
R21473 CSoutput.n242 CSoutput.n192 4.5005
R21474 CSoutput.n242 CSoutput.n241 4.5005
R21475 CSoutput.n224 CSoutput.n188 4.5005
R21476 CSoutput.n224 CSoutput.n190 4.5005
R21477 CSoutput.n224 CSoutput.n187 4.5005
R21478 CSoutput.n224 CSoutput.n191 4.5005
R21479 CSoutput.n224 CSoutput.n186 4.5005
R21480 CSoutput.n224 CSoutput.t155 4.5005
R21481 CSoutput.n224 CSoutput.n185 4.5005
R21482 CSoutput.n224 CSoutput.n192 4.5005
R21483 CSoutput.n241 CSoutput.n224 4.5005
R21484 CSoutput.n196 CSoutput.n188 4.5005
R21485 CSoutput.n196 CSoutput.n190 4.5005
R21486 CSoutput.n196 CSoutput.n187 4.5005
R21487 CSoutput.n196 CSoutput.n191 4.5005
R21488 CSoutput.n196 CSoutput.n186 4.5005
R21489 CSoutput.n196 CSoutput.t155 4.5005
R21490 CSoutput.n196 CSoutput.n185 4.5005
R21491 CSoutput.n196 CSoutput.n192 4.5005
R21492 CSoutput.n241 CSoutput.n196 4.5005
R21493 CSoutput.n226 CSoutput.n188 4.5005
R21494 CSoutput.n226 CSoutput.n190 4.5005
R21495 CSoutput.n226 CSoutput.n187 4.5005
R21496 CSoutput.n226 CSoutput.n191 4.5005
R21497 CSoutput.n226 CSoutput.n186 4.5005
R21498 CSoutput.n226 CSoutput.t155 4.5005
R21499 CSoutput.n226 CSoutput.n185 4.5005
R21500 CSoutput.n226 CSoutput.n192 4.5005
R21501 CSoutput.n241 CSoutput.n226 4.5005
R21502 CSoutput.n195 CSoutput.n188 4.5005
R21503 CSoutput.n195 CSoutput.n190 4.5005
R21504 CSoutput.n195 CSoutput.n187 4.5005
R21505 CSoutput.n195 CSoutput.n191 4.5005
R21506 CSoutput.n195 CSoutput.n186 4.5005
R21507 CSoutput.n195 CSoutput.t155 4.5005
R21508 CSoutput.n195 CSoutput.n185 4.5005
R21509 CSoutput.n195 CSoutput.n192 4.5005
R21510 CSoutput.n241 CSoutput.n195 4.5005
R21511 CSoutput.n240 CSoutput.n188 4.5005
R21512 CSoutput.n240 CSoutput.n190 4.5005
R21513 CSoutput.n240 CSoutput.n187 4.5005
R21514 CSoutput.n240 CSoutput.n191 4.5005
R21515 CSoutput.n240 CSoutput.n186 4.5005
R21516 CSoutput.n240 CSoutput.t155 4.5005
R21517 CSoutput.n240 CSoutput.n185 4.5005
R21518 CSoutput.n240 CSoutput.n192 4.5005
R21519 CSoutput.n241 CSoutput.n240 4.5005
R21520 CSoutput.n239 CSoutput.n124 4.5005
R21521 CSoutput.n140 CSoutput.n124 4.5005
R21522 CSoutput.n135 CSoutput.n119 4.5005
R21523 CSoutput.n135 CSoutput.n121 4.5005
R21524 CSoutput.n135 CSoutput.n118 4.5005
R21525 CSoutput.n135 CSoutput.n122 4.5005
R21526 CSoutput.n135 CSoutput.n117 4.5005
R21527 CSoutput.n135 CSoutput.t154 4.5005
R21528 CSoutput.n135 CSoutput.n116 4.5005
R21529 CSoutput.n135 CSoutput.n123 4.5005
R21530 CSoutput.n135 CSoutput.n124 4.5005
R21531 CSoutput.n133 CSoutput.n119 4.5005
R21532 CSoutput.n133 CSoutput.n121 4.5005
R21533 CSoutput.n133 CSoutput.n118 4.5005
R21534 CSoutput.n133 CSoutput.n122 4.5005
R21535 CSoutput.n133 CSoutput.n117 4.5005
R21536 CSoutput.n133 CSoutput.t154 4.5005
R21537 CSoutput.n133 CSoutput.n116 4.5005
R21538 CSoutput.n133 CSoutput.n123 4.5005
R21539 CSoutput.n133 CSoutput.n124 4.5005
R21540 CSoutput.n132 CSoutput.n119 4.5005
R21541 CSoutput.n132 CSoutput.n121 4.5005
R21542 CSoutput.n132 CSoutput.n118 4.5005
R21543 CSoutput.n132 CSoutput.n122 4.5005
R21544 CSoutput.n132 CSoutput.n117 4.5005
R21545 CSoutput.n132 CSoutput.t154 4.5005
R21546 CSoutput.n132 CSoutput.n116 4.5005
R21547 CSoutput.n132 CSoutput.n123 4.5005
R21548 CSoutput.n132 CSoutput.n124 4.5005
R21549 CSoutput.n261 CSoutput.n119 4.5005
R21550 CSoutput.n261 CSoutput.n121 4.5005
R21551 CSoutput.n261 CSoutput.n118 4.5005
R21552 CSoutput.n261 CSoutput.n122 4.5005
R21553 CSoutput.n261 CSoutput.n117 4.5005
R21554 CSoutput.n261 CSoutput.t154 4.5005
R21555 CSoutput.n261 CSoutput.n116 4.5005
R21556 CSoutput.n261 CSoutput.n123 4.5005
R21557 CSoutput.n261 CSoutput.n124 4.5005
R21558 CSoutput.n259 CSoutput.n119 4.5005
R21559 CSoutput.n259 CSoutput.n121 4.5005
R21560 CSoutput.n259 CSoutput.n118 4.5005
R21561 CSoutput.n259 CSoutput.n122 4.5005
R21562 CSoutput.n259 CSoutput.n117 4.5005
R21563 CSoutput.n259 CSoutput.t154 4.5005
R21564 CSoutput.n259 CSoutput.n116 4.5005
R21565 CSoutput.n259 CSoutput.n123 4.5005
R21566 CSoutput.n257 CSoutput.n119 4.5005
R21567 CSoutput.n257 CSoutput.n121 4.5005
R21568 CSoutput.n257 CSoutput.n118 4.5005
R21569 CSoutput.n257 CSoutput.n122 4.5005
R21570 CSoutput.n257 CSoutput.n117 4.5005
R21571 CSoutput.n257 CSoutput.t154 4.5005
R21572 CSoutput.n257 CSoutput.n116 4.5005
R21573 CSoutput.n257 CSoutput.n123 4.5005
R21574 CSoutput.n143 CSoutput.n119 4.5005
R21575 CSoutput.n143 CSoutput.n121 4.5005
R21576 CSoutput.n143 CSoutput.n118 4.5005
R21577 CSoutput.n143 CSoutput.n122 4.5005
R21578 CSoutput.n143 CSoutput.n117 4.5005
R21579 CSoutput.n143 CSoutput.t154 4.5005
R21580 CSoutput.n143 CSoutput.n116 4.5005
R21581 CSoutput.n143 CSoutput.n123 4.5005
R21582 CSoutput.n143 CSoutput.n124 4.5005
R21583 CSoutput.n142 CSoutput.n119 4.5005
R21584 CSoutput.n142 CSoutput.n121 4.5005
R21585 CSoutput.n142 CSoutput.n118 4.5005
R21586 CSoutput.n142 CSoutput.n122 4.5005
R21587 CSoutput.n142 CSoutput.n117 4.5005
R21588 CSoutput.n142 CSoutput.t154 4.5005
R21589 CSoutput.n142 CSoutput.n116 4.5005
R21590 CSoutput.n142 CSoutput.n123 4.5005
R21591 CSoutput.n142 CSoutput.n124 4.5005
R21592 CSoutput.n146 CSoutput.n119 4.5005
R21593 CSoutput.n146 CSoutput.n121 4.5005
R21594 CSoutput.n146 CSoutput.n118 4.5005
R21595 CSoutput.n146 CSoutput.n122 4.5005
R21596 CSoutput.n146 CSoutput.n117 4.5005
R21597 CSoutput.n146 CSoutput.t154 4.5005
R21598 CSoutput.n146 CSoutput.n116 4.5005
R21599 CSoutput.n146 CSoutput.n123 4.5005
R21600 CSoutput.n146 CSoutput.n124 4.5005
R21601 CSoutput.n145 CSoutput.n119 4.5005
R21602 CSoutput.n145 CSoutput.n121 4.5005
R21603 CSoutput.n145 CSoutput.n118 4.5005
R21604 CSoutput.n145 CSoutput.n122 4.5005
R21605 CSoutput.n145 CSoutput.n117 4.5005
R21606 CSoutput.n145 CSoutput.t154 4.5005
R21607 CSoutput.n145 CSoutput.n116 4.5005
R21608 CSoutput.n145 CSoutput.n123 4.5005
R21609 CSoutput.n145 CSoutput.n124 4.5005
R21610 CSoutput.n128 CSoutput.n119 4.5005
R21611 CSoutput.n128 CSoutput.n121 4.5005
R21612 CSoutput.n128 CSoutput.n118 4.5005
R21613 CSoutput.n128 CSoutput.n122 4.5005
R21614 CSoutput.n128 CSoutput.n117 4.5005
R21615 CSoutput.n128 CSoutput.t154 4.5005
R21616 CSoutput.n128 CSoutput.n116 4.5005
R21617 CSoutput.n128 CSoutput.n123 4.5005
R21618 CSoutput.n128 CSoutput.n124 4.5005
R21619 CSoutput.n264 CSoutput.n119 4.5005
R21620 CSoutput.n264 CSoutput.n121 4.5005
R21621 CSoutput.n264 CSoutput.n118 4.5005
R21622 CSoutput.n264 CSoutput.n122 4.5005
R21623 CSoutput.n264 CSoutput.n117 4.5005
R21624 CSoutput.n264 CSoutput.t154 4.5005
R21625 CSoutput.n264 CSoutput.n116 4.5005
R21626 CSoutput.n264 CSoutput.n123 4.5005
R21627 CSoutput.n264 CSoutput.n124 4.5005
R21628 CSoutput.n299 CSoutput.n287 4.10845
R21629 CSoutput.n113 CSoutput.n101 4.10845
R21630 CSoutput.n297 CSoutput.t55 4.06363
R21631 CSoutput.n297 CSoutput.t6 4.06363
R21632 CSoutput.n295 CSoutput.t2 4.06363
R21633 CSoutput.n295 CSoutput.t31 4.06363
R21634 CSoutput.n293 CSoutput.t42 4.06363
R21635 CSoutput.n293 CSoutput.t57 4.06363
R21636 CSoutput.n291 CSoutput.t66 4.06363
R21637 CSoutput.n291 CSoutput.t14 4.06363
R21638 CSoutput.n289 CSoutput.t19 4.06363
R21639 CSoutput.n289 CSoutput.t58 4.06363
R21640 CSoutput.n288 CSoutput.t68 4.06363
R21641 CSoutput.n288 CSoutput.t69 4.06363
R21642 CSoutput.n285 CSoutput.t49 4.06363
R21643 CSoutput.n285 CSoutput.t70 4.06363
R21644 CSoutput.n283 CSoutput.t67 4.06363
R21645 CSoutput.n283 CSoutput.t24 4.06363
R21646 CSoutput.n281 CSoutput.t33 4.06363
R21647 CSoutput.n281 CSoutput.t50 4.06363
R21648 CSoutput.n279 CSoutput.t59 4.06363
R21649 CSoutput.n279 CSoutput.t5 4.06363
R21650 CSoutput.n277 CSoutput.t7 4.06363
R21651 CSoutput.n277 CSoutput.t53 4.06363
R21652 CSoutput.n276 CSoutput.t62 4.06363
R21653 CSoutput.n276 CSoutput.t63 4.06363
R21654 CSoutput.n274 CSoutput.t51 4.06363
R21655 CSoutput.n274 CSoutput.t22 4.06363
R21656 CSoutput.n272 CSoutput.t64 4.06363
R21657 CSoutput.n272 CSoutput.t37 4.06363
R21658 CSoutput.n270 CSoutput.t56 4.06363
R21659 CSoutput.n270 CSoutput.t28 4.06363
R21660 CSoutput.n268 CSoutput.t46 4.06363
R21661 CSoutput.n268 CSoutput.t15 4.06363
R21662 CSoutput.n266 CSoutput.t60 4.06363
R21663 CSoutput.n266 CSoutput.t9 4.06363
R21664 CSoutput.n265 CSoutput.t34 4.06363
R21665 CSoutput.n265 CSoutput.t20 4.06363
R21666 CSoutput.n102 CSoutput.t44 4.06363
R21667 CSoutput.n102 CSoutput.t27 4.06363
R21668 CSoutput.n103 CSoutput.t13 4.06363
R21669 CSoutput.n103 CSoutput.t45 4.06363
R21670 CSoutput.n105 CSoutput.t43 4.06363
R21671 CSoutput.n105 CSoutput.t25 4.06363
R21672 CSoutput.n107 CSoutput.t12 4.06363
R21673 CSoutput.n107 CSoutput.t11 4.06363
R21674 CSoutput.n109 CSoutput.t54 4.06363
R21675 CSoutput.n109 CSoutput.t32 4.06363
R21676 CSoutput.n111 CSoutput.t30 4.06363
R21677 CSoutput.n111 CSoutput.t8 4.06363
R21678 CSoutput.n90 CSoutput.t39 4.06363
R21679 CSoutput.n90 CSoutput.t18 4.06363
R21680 CSoutput.n91 CSoutput.t4 4.06363
R21681 CSoutput.n91 CSoutput.t40 4.06363
R21682 CSoutput.n93 CSoutput.t36 4.06363
R21683 CSoutput.n93 CSoutput.t16 4.06363
R21684 CSoutput.n95 CSoutput.t3 4.06363
R21685 CSoutput.n95 CSoutput.t1 4.06363
R21686 CSoutput.n97 CSoutput.t48 4.06363
R21687 CSoutput.n97 CSoutput.t26 4.06363
R21688 CSoutput.n99 CSoutput.t23 4.06363
R21689 CSoutput.n99 CSoutput.t0 4.06363
R21690 CSoutput.n79 CSoutput.t71 4.06363
R21691 CSoutput.n79 CSoutput.t35 4.06363
R21692 CSoutput.n80 CSoutput.t10 4.06363
R21693 CSoutput.n80 CSoutput.t61 4.06363
R21694 CSoutput.n82 CSoutput.t17 4.06363
R21695 CSoutput.n82 CSoutput.t47 4.06363
R21696 CSoutput.n84 CSoutput.t29 4.06363
R21697 CSoutput.n84 CSoutput.t41 4.06363
R21698 CSoutput.n86 CSoutput.t38 4.06363
R21699 CSoutput.n86 CSoutput.t65 4.06363
R21700 CSoutput.n88 CSoutput.t21 4.06363
R21701 CSoutput.n88 CSoutput.t52 4.06363
R21702 CSoutput.n44 CSoutput.n43 3.79402
R21703 CSoutput.n49 CSoutput.n48 3.79402
R21704 CSoutput.n335 CSoutput.n323 3.72967
R21705 CSoutput.n371 CSoutput.n359 3.72967
R21706 CSoutput.n373 CSoutput.n372 3.57343
R21707 CSoutput.n372 CSoutput.n336 3.04641
R21708 CSoutput.n333 CSoutput.t116 2.82907
R21709 CSoutput.n333 CSoutput.t73 2.82907
R21710 CSoutput.n331 CSoutput.t142 2.82907
R21711 CSoutput.n331 CSoutput.t131 2.82907
R21712 CSoutput.n329 CSoutput.t98 2.82907
R21713 CSoutput.n329 CSoutput.t107 2.82907
R21714 CSoutput.n327 CSoutput.t72 2.82907
R21715 CSoutput.n327 CSoutput.t138 2.82907
R21716 CSoutput.n325 CSoutput.t132 2.82907
R21717 CSoutput.n325 CSoutput.t87 2.82907
R21718 CSoutput.n324 CSoutput.t80 2.82907
R21719 CSoutput.n324 CSoutput.t141 2.82907
R21720 CSoutput.n321 CSoutput.t83 2.82907
R21721 CSoutput.n321 CSoutput.t93 2.82907
R21722 CSoutput.n319 CSoutput.t91 2.82907
R21723 CSoutput.n319 CSoutput.t79 2.82907
R21724 CSoutput.n317 CSoutput.t104 2.82907
R21725 CSoutput.n317 CSoutput.t84 2.82907
R21726 CSoutput.n315 CSoutput.t85 2.82907
R21727 CSoutput.n315 CSoutput.t92 2.82907
R21728 CSoutput.n313 CSoutput.t90 2.82907
R21729 CSoutput.n313 CSoutput.t102 2.82907
R21730 CSoutput.n312 CSoutput.t103 2.82907
R21731 CSoutput.n312 CSoutput.t86 2.82907
R21732 CSoutput.n310 CSoutput.t125 2.82907
R21733 CSoutput.n310 CSoutput.t95 2.82907
R21734 CSoutput.n308 CSoutput.t76 2.82907
R21735 CSoutput.n308 CSoutput.t111 2.82907
R21736 CSoutput.n306 CSoutput.t94 2.82907
R21737 CSoutput.n306 CSoutput.t105 2.82907
R21738 CSoutput.n304 CSoutput.t106 2.82907
R21739 CSoutput.n304 CSoutput.t137 2.82907
R21740 CSoutput.n302 CSoutput.t121 2.82907
R21741 CSoutput.n302 CSoutput.t74 2.82907
R21742 CSoutput.n301 CSoutput.t134 2.82907
R21743 CSoutput.n301 CSoutput.t81 2.82907
R21744 CSoutput.n360 CSoutput.t129 2.82907
R21745 CSoutput.n360 CSoutput.t140 2.82907
R21746 CSoutput.n361 CSoutput.t143 2.82907
R21747 CSoutput.n361 CSoutput.t120 2.82907
R21748 CSoutput.n363 CSoutput.t124 2.82907
R21749 CSoutput.n363 CSoutput.t135 2.82907
R21750 CSoutput.n365 CSoutput.t82 2.82907
R21751 CSoutput.n365 CSoutput.t114 2.82907
R21752 CSoutput.n367 CSoutput.t119 2.82907
R21753 CSoutput.n367 CSoutput.t130 2.82907
R21754 CSoutput.n369 CSoutput.t136 2.82907
R21755 CSoutput.n369 CSoutput.t123 2.82907
R21756 CSoutput.n348 CSoutput.t100 2.82907
R21757 CSoutput.n348 CSoutput.t117 2.82907
R21758 CSoutput.n349 CSoutput.t118 2.82907
R21759 CSoutput.n349 CSoutput.t109 2.82907
R21760 CSoutput.n351 CSoutput.t108 2.82907
R21761 CSoutput.n351 CSoutput.t101 2.82907
R21762 CSoutput.n353 CSoutput.t96 2.82907
R21763 CSoutput.n353 CSoutput.t88 2.82907
R21764 CSoutput.n355 CSoutput.t89 2.82907
R21765 CSoutput.n355 CSoutput.t110 2.82907
R21766 CSoutput.n357 CSoutput.t112 2.82907
R21767 CSoutput.n357 CSoutput.t75 2.82907
R21768 CSoutput.n337 CSoutput.t113 2.82907
R21769 CSoutput.n337 CSoutput.t77 2.82907
R21770 CSoutput.n338 CSoutput.t97 2.82907
R21771 CSoutput.n338 CSoutput.t139 2.82907
R21772 CSoutput.n340 CSoutput.t78 2.82907
R21773 CSoutput.n340 CSoutput.t127 2.82907
R21774 CSoutput.n342 CSoutput.t126 2.82907
R21775 CSoutput.n342 CSoutput.t115 2.82907
R21776 CSoutput.n344 CSoutput.t128 2.82907
R21777 CSoutput.n344 CSoutput.t99 2.82907
R21778 CSoutput.n346 CSoutput.t122 2.82907
R21779 CSoutput.n346 CSoutput.t133 2.82907
R21780 CSoutput.n300 CSoutput.n114 2.78353
R21781 CSoutput.n75 CSoutput.n1 2.45513
R21782 CSoutput.n205 CSoutput.n203 2.251
R21783 CSoutput.n205 CSoutput.n202 2.251
R21784 CSoutput.n205 CSoutput.n201 2.251
R21785 CSoutput.n205 CSoutput.n200 2.251
R21786 CSoutput.n174 CSoutput.n173 2.251
R21787 CSoutput.n174 CSoutput.n172 2.251
R21788 CSoutput.n174 CSoutput.n171 2.251
R21789 CSoutput.n174 CSoutput.n170 2.251
R21790 CSoutput.n247 CSoutput.n246 2.251
R21791 CSoutput.n212 CSoutput.n210 2.251
R21792 CSoutput.n212 CSoutput.n209 2.251
R21793 CSoutput.n212 CSoutput.n208 2.251
R21794 CSoutput.n230 CSoutput.n212 2.251
R21795 CSoutput.n218 CSoutput.n217 2.251
R21796 CSoutput.n218 CSoutput.n216 2.251
R21797 CSoutput.n218 CSoutput.n215 2.251
R21798 CSoutput.n218 CSoutput.n214 2.251
R21799 CSoutput.n244 CSoutput.n184 2.251
R21800 CSoutput.n239 CSoutput.n237 2.251
R21801 CSoutput.n239 CSoutput.n236 2.251
R21802 CSoutput.n239 CSoutput.n235 2.251
R21803 CSoutput.n239 CSoutput.n234 2.251
R21804 CSoutput.n140 CSoutput.n139 2.251
R21805 CSoutput.n140 CSoutput.n138 2.251
R21806 CSoutput.n140 CSoutput.n137 2.251
R21807 CSoutput.n140 CSoutput.n136 2.251
R21808 CSoutput.n257 CSoutput.n256 2.251
R21809 CSoutput.n174 CSoutput.n154 2.2505
R21810 CSoutput.n169 CSoutput.n154 2.2505
R21811 CSoutput.n167 CSoutput.n154 2.2505
R21812 CSoutput.n166 CSoutput.n154 2.2505
R21813 CSoutput.n251 CSoutput.n154 2.2505
R21814 CSoutput.n249 CSoutput.n154 2.2505
R21815 CSoutput.n247 CSoutput.n154 2.2505
R21816 CSoutput.n177 CSoutput.n154 2.2505
R21817 CSoutput.n176 CSoutput.n154 2.2505
R21818 CSoutput.n180 CSoutput.n154 2.2505
R21819 CSoutput.n179 CSoutput.n154 2.2505
R21820 CSoutput.n162 CSoutput.n154 2.2505
R21821 CSoutput.n254 CSoutput.n154 2.2505
R21822 CSoutput.n254 CSoutput.n253 2.2505
R21823 CSoutput.n218 CSoutput.n189 2.2505
R21824 CSoutput.n199 CSoutput.n189 2.2505
R21825 CSoutput.n220 CSoutput.n189 2.2505
R21826 CSoutput.n198 CSoutput.n189 2.2505
R21827 CSoutput.n222 CSoutput.n189 2.2505
R21828 CSoutput.n189 CSoutput.n183 2.2505
R21829 CSoutput.n244 CSoutput.n189 2.2505
R21830 CSoutput.n242 CSoutput.n189 2.2505
R21831 CSoutput.n224 CSoutput.n189 2.2505
R21832 CSoutput.n196 CSoutput.n189 2.2505
R21833 CSoutput.n226 CSoutput.n189 2.2505
R21834 CSoutput.n195 CSoutput.n189 2.2505
R21835 CSoutput.n240 CSoutput.n189 2.2505
R21836 CSoutput.n240 CSoutput.n193 2.2505
R21837 CSoutput.n140 CSoutput.n120 2.2505
R21838 CSoutput.n135 CSoutput.n120 2.2505
R21839 CSoutput.n133 CSoutput.n120 2.2505
R21840 CSoutput.n132 CSoutput.n120 2.2505
R21841 CSoutput.n261 CSoutput.n120 2.2505
R21842 CSoutput.n259 CSoutput.n120 2.2505
R21843 CSoutput.n257 CSoutput.n120 2.2505
R21844 CSoutput.n143 CSoutput.n120 2.2505
R21845 CSoutput.n142 CSoutput.n120 2.2505
R21846 CSoutput.n146 CSoutput.n120 2.2505
R21847 CSoutput.n145 CSoutput.n120 2.2505
R21848 CSoutput.n128 CSoutput.n120 2.2505
R21849 CSoutput.n264 CSoutput.n120 2.2505
R21850 CSoutput.n264 CSoutput.n263 2.2505
R21851 CSoutput.n182 CSoutput.n175 2.25024
R21852 CSoutput.n182 CSoutput.n168 2.25024
R21853 CSoutput.n250 CSoutput.n182 2.25024
R21854 CSoutput.n182 CSoutput.n178 2.25024
R21855 CSoutput.n182 CSoutput.n181 2.25024
R21856 CSoutput.n182 CSoutput.n149 2.25024
R21857 CSoutput.n232 CSoutput.n229 2.25024
R21858 CSoutput.n232 CSoutput.n228 2.25024
R21859 CSoutput.n232 CSoutput.n227 2.25024
R21860 CSoutput.n232 CSoutput.n194 2.25024
R21861 CSoutput.n232 CSoutput.n231 2.25024
R21862 CSoutput.n233 CSoutput.n232 2.25024
R21863 CSoutput.n148 CSoutput.n141 2.25024
R21864 CSoutput.n148 CSoutput.n134 2.25024
R21865 CSoutput.n260 CSoutput.n148 2.25024
R21866 CSoutput.n148 CSoutput.n144 2.25024
R21867 CSoutput.n148 CSoutput.n147 2.25024
R21868 CSoutput.n148 CSoutput.n115 2.25024
R21869 CSoutput.n249 CSoutput.n159 1.50111
R21870 CSoutput.n197 CSoutput.n183 1.50111
R21871 CSoutput.n259 CSoutput.n125 1.50111
R21872 CSoutput.n205 CSoutput.n204 1.501
R21873 CSoutput.n212 CSoutput.n211 1.501
R21874 CSoutput.n239 CSoutput.n238 1.501
R21875 CSoutput.n253 CSoutput.n164 1.12536
R21876 CSoutput.n253 CSoutput.n165 1.12536
R21877 CSoutput.n253 CSoutput.n252 1.12536
R21878 CSoutput.n213 CSoutput.n193 1.12536
R21879 CSoutput.n219 CSoutput.n193 1.12536
R21880 CSoutput.n221 CSoutput.n193 1.12536
R21881 CSoutput.n263 CSoutput.n130 1.12536
R21882 CSoutput.n263 CSoutput.n131 1.12536
R21883 CSoutput.n263 CSoutput.n262 1.12536
R21884 CSoutput.n253 CSoutput.n160 1.12536
R21885 CSoutput.n253 CSoutput.n161 1.12536
R21886 CSoutput.n253 CSoutput.n163 1.12536
R21887 CSoutput.n243 CSoutput.n193 1.12536
R21888 CSoutput.n223 CSoutput.n193 1.12536
R21889 CSoutput.n225 CSoutput.n193 1.12536
R21890 CSoutput.n263 CSoutput.n126 1.12536
R21891 CSoutput.n263 CSoutput.n127 1.12536
R21892 CSoutput.n263 CSoutput.n129 1.12536
R21893 CSoutput.n31 CSoutput.n30 0.669944
R21894 CSoutput.n62 CSoutput.n61 0.669944
R21895 CSoutput.n328 CSoutput.n326 0.573776
R21896 CSoutput.n330 CSoutput.n328 0.573776
R21897 CSoutput.n332 CSoutput.n330 0.573776
R21898 CSoutput.n334 CSoutput.n332 0.573776
R21899 CSoutput.n316 CSoutput.n314 0.573776
R21900 CSoutput.n318 CSoutput.n316 0.573776
R21901 CSoutput.n320 CSoutput.n318 0.573776
R21902 CSoutput.n322 CSoutput.n320 0.573776
R21903 CSoutput.n305 CSoutput.n303 0.573776
R21904 CSoutput.n307 CSoutput.n305 0.573776
R21905 CSoutput.n309 CSoutput.n307 0.573776
R21906 CSoutput.n311 CSoutput.n309 0.573776
R21907 CSoutput.n370 CSoutput.n368 0.573776
R21908 CSoutput.n368 CSoutput.n366 0.573776
R21909 CSoutput.n366 CSoutput.n364 0.573776
R21910 CSoutput.n364 CSoutput.n362 0.573776
R21911 CSoutput.n358 CSoutput.n356 0.573776
R21912 CSoutput.n356 CSoutput.n354 0.573776
R21913 CSoutput.n354 CSoutput.n352 0.573776
R21914 CSoutput.n352 CSoutput.n350 0.573776
R21915 CSoutput.n347 CSoutput.n345 0.573776
R21916 CSoutput.n345 CSoutput.n343 0.573776
R21917 CSoutput.n343 CSoutput.n341 0.573776
R21918 CSoutput.n341 CSoutput.n339 0.573776
R21919 CSoutput.n373 CSoutput.n264 0.53442
R21920 CSoutput.n292 CSoutput.n290 0.358259
R21921 CSoutput.n294 CSoutput.n292 0.358259
R21922 CSoutput.n296 CSoutput.n294 0.358259
R21923 CSoutput.n298 CSoutput.n296 0.358259
R21924 CSoutput.n280 CSoutput.n278 0.358259
R21925 CSoutput.n282 CSoutput.n280 0.358259
R21926 CSoutput.n284 CSoutput.n282 0.358259
R21927 CSoutput.n286 CSoutput.n284 0.358259
R21928 CSoutput.n269 CSoutput.n267 0.358259
R21929 CSoutput.n271 CSoutput.n269 0.358259
R21930 CSoutput.n273 CSoutput.n271 0.358259
R21931 CSoutput.n275 CSoutput.n273 0.358259
R21932 CSoutput.n112 CSoutput.n110 0.358259
R21933 CSoutput.n110 CSoutput.n108 0.358259
R21934 CSoutput.n108 CSoutput.n106 0.358259
R21935 CSoutput.n106 CSoutput.n104 0.358259
R21936 CSoutput.n100 CSoutput.n98 0.358259
R21937 CSoutput.n98 CSoutput.n96 0.358259
R21938 CSoutput.n96 CSoutput.n94 0.358259
R21939 CSoutput.n94 CSoutput.n92 0.358259
R21940 CSoutput.n89 CSoutput.n87 0.358259
R21941 CSoutput.n87 CSoutput.n85 0.358259
R21942 CSoutput.n85 CSoutput.n83 0.358259
R21943 CSoutput.n83 CSoutput.n81 0.358259
R21944 CSoutput.n21 CSoutput.n20 0.169105
R21945 CSoutput.n21 CSoutput.n16 0.169105
R21946 CSoutput.n26 CSoutput.n16 0.169105
R21947 CSoutput.n27 CSoutput.n26 0.169105
R21948 CSoutput.n27 CSoutput.n14 0.169105
R21949 CSoutput.n32 CSoutput.n14 0.169105
R21950 CSoutput.n33 CSoutput.n32 0.169105
R21951 CSoutput.n34 CSoutput.n33 0.169105
R21952 CSoutput.n34 CSoutput.n12 0.169105
R21953 CSoutput.n39 CSoutput.n12 0.169105
R21954 CSoutput.n40 CSoutput.n39 0.169105
R21955 CSoutput.n40 CSoutput.n10 0.169105
R21956 CSoutput.n45 CSoutput.n10 0.169105
R21957 CSoutput.n46 CSoutput.n45 0.169105
R21958 CSoutput.n47 CSoutput.n46 0.169105
R21959 CSoutput.n47 CSoutput.n8 0.169105
R21960 CSoutput.n52 CSoutput.n8 0.169105
R21961 CSoutput.n53 CSoutput.n52 0.169105
R21962 CSoutput.n53 CSoutput.n6 0.169105
R21963 CSoutput.n58 CSoutput.n6 0.169105
R21964 CSoutput.n59 CSoutput.n58 0.169105
R21965 CSoutput.n60 CSoutput.n59 0.169105
R21966 CSoutput.n60 CSoutput.n4 0.169105
R21967 CSoutput.n66 CSoutput.n4 0.169105
R21968 CSoutput.n67 CSoutput.n66 0.169105
R21969 CSoutput.n68 CSoutput.n67 0.169105
R21970 CSoutput.n68 CSoutput.n2 0.169105
R21971 CSoutput.n73 CSoutput.n2 0.169105
R21972 CSoutput.n74 CSoutput.n73 0.169105
R21973 CSoutput.n74 CSoutput.n0 0.169105
R21974 CSoutput.n78 CSoutput.n0 0.169105
R21975 CSoutput.n207 CSoutput.n206 0.0910737
R21976 CSoutput.n258 CSoutput.n255 0.0723685
R21977 CSoutput.n212 CSoutput.n207 0.0522944
R21978 CSoutput.n255 CSoutput.n254 0.0499135
R21979 CSoutput.n206 CSoutput.n205 0.0499135
R21980 CSoutput.n240 CSoutput.n239 0.0464294
R21981 CSoutput.n248 CSoutput.n245 0.0391444
R21982 CSoutput.n207 CSoutput.t163 0.023435
R21983 CSoutput.n255 CSoutput.t144 0.02262
R21984 CSoutput.n206 CSoutput.t146 0.02262
R21985 CSoutput CSoutput.n373 0.0052
R21986 CSoutput.n177 CSoutput.n160 0.00365111
R21987 CSoutput.n180 CSoutput.n161 0.00365111
R21988 CSoutput.n163 CSoutput.n162 0.00365111
R21989 CSoutput.n205 CSoutput.n164 0.00365111
R21990 CSoutput.n169 CSoutput.n165 0.00365111
R21991 CSoutput.n252 CSoutput.n166 0.00365111
R21992 CSoutput.n243 CSoutput.n242 0.00365111
R21993 CSoutput.n223 CSoutput.n196 0.00365111
R21994 CSoutput.n225 CSoutput.n195 0.00365111
R21995 CSoutput.n213 CSoutput.n212 0.00365111
R21996 CSoutput.n219 CSoutput.n199 0.00365111
R21997 CSoutput.n221 CSoutput.n198 0.00365111
R21998 CSoutput.n143 CSoutput.n126 0.00365111
R21999 CSoutput.n146 CSoutput.n127 0.00365111
R22000 CSoutput.n129 CSoutput.n128 0.00365111
R22001 CSoutput.n239 CSoutput.n130 0.00365111
R22002 CSoutput.n135 CSoutput.n131 0.00365111
R22003 CSoutput.n262 CSoutput.n132 0.00365111
R22004 CSoutput.n174 CSoutput.n164 0.00340054
R22005 CSoutput.n167 CSoutput.n165 0.00340054
R22006 CSoutput.n252 CSoutput.n251 0.00340054
R22007 CSoutput.n247 CSoutput.n160 0.00340054
R22008 CSoutput.n176 CSoutput.n161 0.00340054
R22009 CSoutput.n179 CSoutput.n163 0.00340054
R22010 CSoutput.n218 CSoutput.n213 0.00340054
R22011 CSoutput.n220 CSoutput.n219 0.00340054
R22012 CSoutput.n222 CSoutput.n221 0.00340054
R22013 CSoutput.n244 CSoutput.n243 0.00340054
R22014 CSoutput.n224 CSoutput.n223 0.00340054
R22015 CSoutput.n226 CSoutput.n225 0.00340054
R22016 CSoutput.n140 CSoutput.n130 0.00340054
R22017 CSoutput.n133 CSoutput.n131 0.00340054
R22018 CSoutput.n262 CSoutput.n261 0.00340054
R22019 CSoutput.n257 CSoutput.n126 0.00340054
R22020 CSoutput.n142 CSoutput.n127 0.00340054
R22021 CSoutput.n145 CSoutput.n129 0.00340054
R22022 CSoutput.n175 CSoutput.n169 0.00252698
R22023 CSoutput.n168 CSoutput.n166 0.00252698
R22024 CSoutput.n250 CSoutput.n249 0.00252698
R22025 CSoutput.n178 CSoutput.n176 0.00252698
R22026 CSoutput.n181 CSoutput.n179 0.00252698
R22027 CSoutput.n254 CSoutput.n149 0.00252698
R22028 CSoutput.n175 CSoutput.n174 0.00252698
R22029 CSoutput.n168 CSoutput.n167 0.00252698
R22030 CSoutput.n251 CSoutput.n250 0.00252698
R22031 CSoutput.n178 CSoutput.n177 0.00252698
R22032 CSoutput.n181 CSoutput.n180 0.00252698
R22033 CSoutput.n162 CSoutput.n149 0.00252698
R22034 CSoutput.n229 CSoutput.n199 0.00252698
R22035 CSoutput.n228 CSoutput.n198 0.00252698
R22036 CSoutput.n227 CSoutput.n183 0.00252698
R22037 CSoutput.n224 CSoutput.n194 0.00252698
R22038 CSoutput.n231 CSoutput.n226 0.00252698
R22039 CSoutput.n240 CSoutput.n233 0.00252698
R22040 CSoutput.n229 CSoutput.n218 0.00252698
R22041 CSoutput.n228 CSoutput.n220 0.00252698
R22042 CSoutput.n227 CSoutput.n222 0.00252698
R22043 CSoutput.n242 CSoutput.n194 0.00252698
R22044 CSoutput.n231 CSoutput.n196 0.00252698
R22045 CSoutput.n233 CSoutput.n195 0.00252698
R22046 CSoutput.n141 CSoutput.n135 0.00252698
R22047 CSoutput.n134 CSoutput.n132 0.00252698
R22048 CSoutput.n260 CSoutput.n259 0.00252698
R22049 CSoutput.n144 CSoutput.n142 0.00252698
R22050 CSoutput.n147 CSoutput.n145 0.00252698
R22051 CSoutput.n264 CSoutput.n115 0.00252698
R22052 CSoutput.n141 CSoutput.n140 0.00252698
R22053 CSoutput.n134 CSoutput.n133 0.00252698
R22054 CSoutput.n261 CSoutput.n260 0.00252698
R22055 CSoutput.n144 CSoutput.n143 0.00252698
R22056 CSoutput.n147 CSoutput.n146 0.00252698
R22057 CSoutput.n128 CSoutput.n115 0.00252698
R22058 CSoutput.n249 CSoutput.n248 0.0020275
R22059 CSoutput.n248 CSoutput.n247 0.0020275
R22060 CSoutput.n245 CSoutput.n183 0.0020275
R22061 CSoutput.n245 CSoutput.n244 0.0020275
R22062 CSoutput.n259 CSoutput.n258 0.0020275
R22063 CSoutput.n258 CSoutput.n257 0.0020275
R22064 CSoutput.n159 CSoutput.n158 0.00166668
R22065 CSoutput.n241 CSoutput.n197 0.00166668
R22066 CSoutput.n125 CSoutput.n124 0.00166668
R22067 CSoutput.n263 CSoutput.n125 0.00133328
R22068 CSoutput.n197 CSoutput.n193 0.00133328
R22069 CSoutput.n253 CSoutput.n159 0.00133328
R22070 CSoutput.n256 CSoutput.n148 0.001
R22071 CSoutput.n234 CSoutput.n148 0.001
R22072 CSoutput.n136 CSoutput.n116 0.001
R22073 CSoutput.n235 CSoutput.n116 0.001
R22074 CSoutput.n137 CSoutput.n117 0.001
R22075 CSoutput.n236 CSoutput.n117 0.001
R22076 CSoutput.n138 CSoutput.n118 0.001
R22077 CSoutput.n237 CSoutput.n118 0.001
R22078 CSoutput.n139 CSoutput.n119 0.001
R22079 CSoutput.n238 CSoutput.n119 0.001
R22080 CSoutput.n232 CSoutput.n184 0.001
R22081 CSoutput.n232 CSoutput.n230 0.001
R22082 CSoutput.n214 CSoutput.n185 0.001
R22083 CSoutput.n208 CSoutput.n185 0.001
R22084 CSoutput.n215 CSoutput.n186 0.001
R22085 CSoutput.n209 CSoutput.n186 0.001
R22086 CSoutput.n216 CSoutput.n187 0.001
R22087 CSoutput.n210 CSoutput.n187 0.001
R22088 CSoutput.n217 CSoutput.n188 0.001
R22089 CSoutput.n211 CSoutput.n188 0.001
R22090 CSoutput.n246 CSoutput.n182 0.001
R22091 CSoutput.n200 CSoutput.n182 0.001
R22092 CSoutput.n170 CSoutput.n150 0.001
R22093 CSoutput.n201 CSoutput.n150 0.001
R22094 CSoutput.n171 CSoutput.n151 0.001
R22095 CSoutput.n202 CSoutput.n151 0.001
R22096 CSoutput.n172 CSoutput.n152 0.001
R22097 CSoutput.n203 CSoutput.n152 0.001
R22098 CSoutput.n173 CSoutput.n153 0.001
R22099 CSoutput.n204 CSoutput.n153 0.001
R22100 CSoutput.n204 CSoutput.n154 0.001
R22101 CSoutput.n203 CSoutput.n155 0.001
R22102 CSoutput.n202 CSoutput.n156 0.001
R22103 CSoutput.n201 CSoutput.t162 0.001
R22104 CSoutput.n200 CSoutput.n157 0.001
R22105 CSoutput.n173 CSoutput.n155 0.001
R22106 CSoutput.n172 CSoutput.n156 0.001
R22107 CSoutput.n171 CSoutput.t162 0.001
R22108 CSoutput.n170 CSoutput.n157 0.001
R22109 CSoutput.n246 CSoutput.n158 0.001
R22110 CSoutput.n211 CSoutput.n189 0.001
R22111 CSoutput.n210 CSoutput.n190 0.001
R22112 CSoutput.n209 CSoutput.n191 0.001
R22113 CSoutput.n208 CSoutput.t155 0.001
R22114 CSoutput.n230 CSoutput.n192 0.001
R22115 CSoutput.n217 CSoutput.n190 0.001
R22116 CSoutput.n216 CSoutput.n191 0.001
R22117 CSoutput.n215 CSoutput.t155 0.001
R22118 CSoutput.n214 CSoutput.n192 0.001
R22119 CSoutput.n241 CSoutput.n184 0.001
R22120 CSoutput.n238 CSoutput.n120 0.001
R22121 CSoutput.n237 CSoutput.n121 0.001
R22122 CSoutput.n236 CSoutput.n122 0.001
R22123 CSoutput.n235 CSoutput.t154 0.001
R22124 CSoutput.n234 CSoutput.n123 0.001
R22125 CSoutput.n139 CSoutput.n121 0.001
R22126 CSoutput.n138 CSoutput.n122 0.001
R22127 CSoutput.n137 CSoutput.t154 0.001
R22128 CSoutput.n136 CSoutput.n123 0.001
R22129 CSoutput.n256 CSoutput.n124 0.001
R22130 diffpairibias.n0 diffpairibias.t27 436.822
R22131 diffpairibias.n27 diffpairibias.t24 435.479
R22132 diffpairibias.n26 diffpairibias.t21 435.479
R22133 diffpairibias.n25 diffpairibias.t22 435.479
R22134 diffpairibias.n24 diffpairibias.t26 435.479
R22135 diffpairibias.n23 diffpairibias.t20 435.479
R22136 diffpairibias.n0 diffpairibias.t23 435.479
R22137 diffpairibias.n1 diffpairibias.t28 435.479
R22138 diffpairibias.n2 diffpairibias.t25 435.479
R22139 diffpairibias.n3 diffpairibias.t29 435.479
R22140 diffpairibias.n13 diffpairibias.t14 377.536
R22141 diffpairibias.n13 diffpairibias.t0 376.193
R22142 diffpairibias.n14 diffpairibias.t10 376.193
R22143 diffpairibias.n15 diffpairibias.t12 376.193
R22144 diffpairibias.n16 diffpairibias.t6 376.193
R22145 diffpairibias.n17 diffpairibias.t2 376.193
R22146 diffpairibias.n18 diffpairibias.t16 376.193
R22147 diffpairibias.n19 diffpairibias.t4 376.193
R22148 diffpairibias.n20 diffpairibias.t18 376.193
R22149 diffpairibias.n21 diffpairibias.t8 376.193
R22150 diffpairibias.n4 diffpairibias.t15 113.368
R22151 diffpairibias.n4 diffpairibias.t1 112.698
R22152 diffpairibias.n5 diffpairibias.t11 112.698
R22153 diffpairibias.n6 diffpairibias.t13 112.698
R22154 diffpairibias.n7 diffpairibias.t7 112.698
R22155 diffpairibias.n8 diffpairibias.t3 112.698
R22156 diffpairibias.n9 diffpairibias.t17 112.698
R22157 diffpairibias.n10 diffpairibias.t5 112.698
R22158 diffpairibias.n11 diffpairibias.t19 112.698
R22159 diffpairibias.n12 diffpairibias.t9 112.698
R22160 diffpairibias.n22 diffpairibias.n21 4.77242
R22161 diffpairibias.n22 diffpairibias.n12 4.30807
R22162 diffpairibias.n23 diffpairibias.n22 4.13945
R22163 diffpairibias.n21 diffpairibias.n20 1.34352
R22164 diffpairibias.n20 diffpairibias.n19 1.34352
R22165 diffpairibias.n19 diffpairibias.n18 1.34352
R22166 diffpairibias.n18 diffpairibias.n17 1.34352
R22167 diffpairibias.n17 diffpairibias.n16 1.34352
R22168 diffpairibias.n16 diffpairibias.n15 1.34352
R22169 diffpairibias.n15 diffpairibias.n14 1.34352
R22170 diffpairibias.n14 diffpairibias.n13 1.34352
R22171 diffpairibias.n3 diffpairibias.n2 1.34352
R22172 diffpairibias.n2 diffpairibias.n1 1.34352
R22173 diffpairibias.n1 diffpairibias.n0 1.34352
R22174 diffpairibias.n24 diffpairibias.n23 1.34352
R22175 diffpairibias.n25 diffpairibias.n24 1.34352
R22176 diffpairibias.n26 diffpairibias.n25 1.34352
R22177 diffpairibias.n27 diffpairibias.n26 1.34352
R22178 diffpairibias.n28 diffpairibias.n27 0.862419
R22179 diffpairibias diffpairibias.n28 0.684875
R22180 diffpairibias.n12 diffpairibias.n11 0.672012
R22181 diffpairibias.n11 diffpairibias.n10 0.672012
R22182 diffpairibias.n10 diffpairibias.n9 0.672012
R22183 diffpairibias.n9 diffpairibias.n8 0.672012
R22184 diffpairibias.n8 diffpairibias.n7 0.672012
R22185 diffpairibias.n7 diffpairibias.n6 0.672012
R22186 diffpairibias.n6 diffpairibias.n5 0.672012
R22187 diffpairibias.n5 diffpairibias.n4 0.672012
R22188 diffpairibias.n28 diffpairibias.n3 0.190907
R22189 a_n3827_n3924.n51 a_n3827_n3924.t43 214.994
R22190 a_n3827_n3924.t50 a_n3827_n3924.n58 214.994
R22191 a_n3827_n3924.n51 a_n3827_n3924.t47 214.321
R22192 a_n3827_n3924.n53 a_n3827_n3924.t42 214.321
R22193 a_n3827_n3924.n54 a_n3827_n3924.t45 214.321
R22194 a_n3827_n3924.n55 a_n3827_n3924.t41 214.321
R22195 a_n3827_n3924.n56 a_n3827_n3924.t46 214.321
R22196 a_n3827_n3924.n57 a_n3827_n3924.t49 214.321
R22197 a_n3827_n3924.n0 a_n3827_n3924.t48 214.321
R22198 a_n3827_n3924.n58 a_n3827_n3924.t44 214.321
R22199 a_n3827_n3924.n14 a_n3827_n3924.t27 55.8337
R22200 a_n3827_n3924.n13 a_n3827_n3924.t20 55.8337
R22201 a_n3827_n3924.n2 a_n3827_n3924.t26 55.8337
R22202 a_n3827_n3924.n25 a_n3827_n3924.t2 55.8335
R22203 a_n3827_n3924.n49 a_n3827_n3924.t36 55.8335
R22204 a_n3827_n3924.n38 a_n3827_n3924.t35 55.8335
R22205 a_n3827_n3924.n37 a_n3827_n3924.t19 55.8335
R22206 a_n3827_n3924.n26 a_n3827_n3924.t14 55.8335
R22207 a_n3827_n3924.n24 a_n3827_n3924.n23 53.0052
R22208 a_n3827_n3924.n22 a_n3827_n3924.n21 53.0052
R22209 a_n3827_n3924.n20 a_n3827_n3924.n19 53.0052
R22210 a_n3827_n3924.n18 a_n3827_n3924.n17 53.0052
R22211 a_n3827_n3924.n16 a_n3827_n3924.n15 53.0052
R22212 a_n3827_n3924.n12 a_n3827_n3924.n11 53.0052
R22213 a_n3827_n3924.n10 a_n3827_n3924.n9 53.0052
R22214 a_n3827_n3924.n8 a_n3827_n3924.n7 53.0052
R22215 a_n3827_n3924.n6 a_n3827_n3924.n5 53.0052
R22216 a_n3827_n3924.n4 a_n3827_n3924.n3 53.0052
R22217 a_n3827_n3924.n48 a_n3827_n3924.n47 53.0051
R22218 a_n3827_n3924.n46 a_n3827_n3924.n45 53.0051
R22219 a_n3827_n3924.n44 a_n3827_n3924.n43 53.0051
R22220 a_n3827_n3924.n42 a_n3827_n3924.n41 53.0051
R22221 a_n3827_n3924.n40 a_n3827_n3924.n39 53.0051
R22222 a_n3827_n3924.n36 a_n3827_n3924.n35 53.0051
R22223 a_n3827_n3924.n34 a_n3827_n3924.n33 53.0051
R22224 a_n3827_n3924.n32 a_n3827_n3924.n31 53.0051
R22225 a_n3827_n3924.n30 a_n3827_n3924.n29 53.0051
R22226 a_n3827_n3924.n28 a_n3827_n3924.n27 53.0051
R22227 a_n3827_n3924.n2 a_n3827_n3924.n1 12.1555
R22228 a_n3827_n3924.n50 a_n3827_n3924.n25 12.1555
R22229 a_n3827_n3924.n26 a_n3827_n3924.n1 5.07593
R22230 a_n3827_n3924.n50 a_n3827_n3924.n49 5.07593
R22231 a_n3827_n3924.n47 a_n3827_n3924.t25 2.82907
R22232 a_n3827_n3924.n47 a_n3827_n3924.t6 2.82907
R22233 a_n3827_n3924.n45 a_n3827_n3924.t12 2.82907
R22234 a_n3827_n3924.n45 a_n3827_n3924.t7 2.82907
R22235 a_n3827_n3924.n43 a_n3827_n3924.t31 2.82907
R22236 a_n3827_n3924.n43 a_n3827_n3924.t13 2.82907
R22237 a_n3827_n3924.n41 a_n3827_n3924.t21 2.82907
R22238 a_n3827_n3924.n41 a_n3827_n3924.t34 2.82907
R22239 a_n3827_n3924.n39 a_n3827_n3924.t18 2.82907
R22240 a_n3827_n3924.n39 a_n3827_n3924.t8 2.82907
R22241 a_n3827_n3924.n35 a_n3827_n3924.t33 2.82907
R22242 a_n3827_n3924.n35 a_n3827_n3924.t54 2.82907
R22243 a_n3827_n3924.n33 a_n3827_n3924.t29 2.82907
R22244 a_n3827_n3924.n33 a_n3827_n3924.t23 2.82907
R22245 a_n3827_n3924.n31 a_n3827_n3924.t24 2.82907
R22246 a_n3827_n3924.n31 a_n3827_n3924.t53 2.82907
R22247 a_n3827_n3924.n29 a_n3827_n3924.t4 2.82907
R22248 a_n3827_n3924.n29 a_n3827_n3924.t5 2.82907
R22249 a_n3827_n3924.n27 a_n3827_n3924.t11 2.82907
R22250 a_n3827_n3924.n27 a_n3827_n3924.t51 2.82907
R22251 a_n3827_n3924.n23 a_n3827_n3924.t56 2.82907
R22252 a_n3827_n3924.n23 a_n3827_n3924.t30 2.82907
R22253 a_n3827_n3924.n21 a_n3827_n3924.t52 2.82907
R22254 a_n3827_n3924.n21 a_n3827_n3924.t0 2.82907
R22255 a_n3827_n3924.n19 a_n3827_n3924.t22 2.82907
R22256 a_n3827_n3924.n19 a_n3827_n3924.t17 2.82907
R22257 a_n3827_n3924.n17 a_n3827_n3924.t39 2.82907
R22258 a_n3827_n3924.n17 a_n3827_n3924.t32 2.82907
R22259 a_n3827_n3924.n15 a_n3827_n3924.t3 2.82907
R22260 a_n3827_n3924.n15 a_n3827_n3924.t10 2.82907
R22261 a_n3827_n3924.n11 a_n3827_n3924.t28 2.82907
R22262 a_n3827_n3924.n11 a_n3827_n3924.t38 2.82907
R22263 a_n3827_n3924.n9 a_n3827_n3924.t57 2.82907
R22264 a_n3827_n3924.n9 a_n3827_n3924.t16 2.82907
R22265 a_n3827_n3924.n7 a_n3827_n3924.t15 2.82907
R22266 a_n3827_n3924.n7 a_n3827_n3924.t9 2.82907
R22267 a_n3827_n3924.n5 a_n3827_n3924.t40 2.82907
R22268 a_n3827_n3924.n5 a_n3827_n3924.t37 2.82907
R22269 a_n3827_n3924.n3 a_n3827_n3924.t55 2.82907
R22270 a_n3827_n3924.n3 a_n3827_n3924.t1 2.82907
R22271 a_n3827_n3924.n0 a_n3827_n3924.n1 1.95694
R22272 a_n3827_n3924.n52 a_n3827_n3924.n50 1.95694
R22273 a_n3827_n3924.n58 a_n3827_n3924.n0 0.672012
R22274 a_n3827_n3924.n57 a_n3827_n3924.n56 0.672012
R22275 a_n3827_n3924.n56 a_n3827_n3924.n55 0.672012
R22276 a_n3827_n3924.n55 a_n3827_n3924.n54 0.672012
R22277 a_n3827_n3924.n54 a_n3827_n3924.n53 0.672012
R22278 a_n3827_n3924.n0 a_n3827_n3924.n57 0.672012
R22279 a_n3827_n3924.n53 a_n3827_n3924.n52 0.501227
R22280 a_n3827_n3924.n4 a_n3827_n3924.n2 0.358259
R22281 a_n3827_n3924.n6 a_n3827_n3924.n4 0.358259
R22282 a_n3827_n3924.n8 a_n3827_n3924.n6 0.358259
R22283 a_n3827_n3924.n10 a_n3827_n3924.n8 0.358259
R22284 a_n3827_n3924.n12 a_n3827_n3924.n10 0.358259
R22285 a_n3827_n3924.n13 a_n3827_n3924.n12 0.358259
R22286 a_n3827_n3924.n16 a_n3827_n3924.n14 0.358259
R22287 a_n3827_n3924.n18 a_n3827_n3924.n16 0.358259
R22288 a_n3827_n3924.n20 a_n3827_n3924.n18 0.358259
R22289 a_n3827_n3924.n22 a_n3827_n3924.n20 0.358259
R22290 a_n3827_n3924.n24 a_n3827_n3924.n22 0.358259
R22291 a_n3827_n3924.n25 a_n3827_n3924.n24 0.358259
R22292 a_n3827_n3924.n28 a_n3827_n3924.n26 0.358259
R22293 a_n3827_n3924.n30 a_n3827_n3924.n28 0.358259
R22294 a_n3827_n3924.n32 a_n3827_n3924.n30 0.358259
R22295 a_n3827_n3924.n34 a_n3827_n3924.n32 0.358259
R22296 a_n3827_n3924.n36 a_n3827_n3924.n34 0.358259
R22297 a_n3827_n3924.n37 a_n3827_n3924.n36 0.358259
R22298 a_n3827_n3924.n40 a_n3827_n3924.n38 0.358259
R22299 a_n3827_n3924.n42 a_n3827_n3924.n40 0.358259
R22300 a_n3827_n3924.n44 a_n3827_n3924.n42 0.358259
R22301 a_n3827_n3924.n46 a_n3827_n3924.n44 0.358259
R22302 a_n3827_n3924.n48 a_n3827_n3924.n46 0.358259
R22303 a_n3827_n3924.n49 a_n3827_n3924.n48 0.358259
R22304 a_n3827_n3924.n14 a_n3827_n3924.n13 0.235414
R22305 a_n3827_n3924.n38 a_n3827_n3924.n37 0.235414
R22306 a_n3827_n3924.n52 a_n3827_n3924.n51 0.171285
R22307 a_n2982_8322.n28 a_n2982_8322.t20 74.6477
R22308 a_n2982_8322.n13 a_n2982_8322.t9 74.6477
R22309 a_n2982_8322.n1 a_n2982_8322.t35 74.6474
R22310 a_n2982_8322.n20 a_n2982_8322.t14 74.2899
R22311 a_n2982_8322.n10 a_n2982_8322.t15 74.2899
R22312 a_n2982_8322.n14 a_n2982_8322.t7 74.2899
R22313 a_n2982_8322.n15 a_n2982_8322.t10 74.2899
R22314 a_n2982_8322.n18 a_n2982_8322.t11 74.2899
R22315 a_n2982_8322.n28 a_n2982_8322.n27 70.6783
R22316 a_n2982_8322.n26 a_n2982_8322.n25 70.6783
R22317 a_n2982_8322.n24 a_n2982_8322.n23 70.6783
R22318 a_n2982_8322.n22 a_n2982_8322.n21 70.6783
R22319 a_n2982_8322.n1 a_n2982_8322.n0 70.6783
R22320 a_n2982_8322.n3 a_n2982_8322.n2 70.6783
R22321 a_n2982_8322.n5 a_n2982_8322.n4 70.6783
R22322 a_n2982_8322.n7 a_n2982_8322.n6 70.6783
R22323 a_n2982_8322.n9 a_n2982_8322.n8 70.6783
R22324 a_n2982_8322.n13 a_n2982_8322.n12 70.6783
R22325 a_n2982_8322.n17 a_n2982_8322.n16 70.6783
R22326 a_n2982_8322.n30 a_n2982_8322.n29 70.6782
R22327 a_n2982_8322.n20 a_n2982_8322.n19 24.9022
R22328 a_n2982_8322.n11 a_n2982_8322.t0 9.63019
R22329 a_n2982_8322.n19 a_n2982_8322.n18 8.38735
R22330 a_n2982_8322.n11 a_n2982_8322.n10 6.90998
R22331 a_n2982_8322.n19 a_n2982_8322.n11 5.3452
R22332 a_n2982_8322.n27 a_n2982_8322.t33 3.61217
R22333 a_n2982_8322.n27 a_n2982_8322.t29 3.61217
R22334 a_n2982_8322.n25 a_n2982_8322.t17 3.61217
R22335 a_n2982_8322.n25 a_n2982_8322.t16 3.61217
R22336 a_n2982_8322.n23 a_n2982_8322.t30 3.61217
R22337 a_n2982_8322.n23 a_n2982_8322.t23 3.61217
R22338 a_n2982_8322.n21 a_n2982_8322.t27 3.61217
R22339 a_n2982_8322.n21 a_n2982_8322.t25 3.61217
R22340 a_n2982_8322.n0 a_n2982_8322.t28 3.61217
R22341 a_n2982_8322.n0 a_n2982_8322.t24 3.61217
R22342 a_n2982_8322.n2 a_n2982_8322.t21 3.61217
R22343 a_n2982_8322.n2 a_n2982_8322.t37 3.61217
R22344 a_n2982_8322.n4 a_n2982_8322.t34 3.61217
R22345 a_n2982_8322.n4 a_n2982_8322.t22 3.61217
R22346 a_n2982_8322.n6 a_n2982_8322.t19 3.61217
R22347 a_n2982_8322.n6 a_n2982_8322.t18 3.61217
R22348 a_n2982_8322.n8 a_n2982_8322.t32 3.61217
R22349 a_n2982_8322.n8 a_n2982_8322.t31 3.61217
R22350 a_n2982_8322.n12 a_n2982_8322.t13 3.61217
R22351 a_n2982_8322.n12 a_n2982_8322.t12 3.61217
R22352 a_n2982_8322.n16 a_n2982_8322.t8 3.61217
R22353 a_n2982_8322.n16 a_n2982_8322.t6 3.61217
R22354 a_n2982_8322.t36 a_n2982_8322.n30 3.61217
R22355 a_n2982_8322.n30 a_n2982_8322.t26 3.61217
R22356 a_n2982_8322.n10 a_n2982_8322.n9 0.358259
R22357 a_n2982_8322.n9 a_n2982_8322.n7 0.358259
R22358 a_n2982_8322.n7 a_n2982_8322.n5 0.358259
R22359 a_n2982_8322.n5 a_n2982_8322.n3 0.358259
R22360 a_n2982_8322.n3 a_n2982_8322.n1 0.358259
R22361 a_n2982_8322.n18 a_n2982_8322.n17 0.358259
R22362 a_n2982_8322.n17 a_n2982_8322.n15 0.358259
R22363 a_n2982_8322.n14 a_n2982_8322.n13 0.358259
R22364 a_n2982_8322.n22 a_n2982_8322.n20 0.358259
R22365 a_n2982_8322.n24 a_n2982_8322.n22 0.358259
R22366 a_n2982_8322.n26 a_n2982_8322.n24 0.358259
R22367 a_n2982_8322.n29 a_n2982_8322.n26 0.358259
R22368 a_n2982_8322.n29 a_n2982_8322.n28 0.358259
R22369 a_n2982_8322.n15 a_n2982_8322.n14 0.101793
R22370 a_n2982_8322.t5 a_n2982_8322.t3 0.0788333
R22371 a_n2982_8322.t1 a_n2982_8322.t2 0.0788333
R22372 a_n2982_8322.t0 a_n2982_8322.t4 0.0788333
R22373 a_n2982_8322.t1 a_n2982_8322.t5 0.0318333
R22374 a_n2982_8322.t0 a_n2982_8322.t2 0.0318333
R22375 a_n2982_8322.t3 a_n2982_8322.t2 0.0318333
R22376 a_n2982_8322.t4 a_n2982_8322.t1 0.0318333
R22377 plus.n43 plus.t25 442.325
R22378 plus.n11 plus.t12 442.325
R22379 plus.n42 plus.t5 415.966
R22380 plus.n41 plus.t20 415.966
R22381 plus.n47 plus.t26 415.966
R22382 plus.n39 plus.t11 415.966
R22383 plus.n52 plus.t6 415.966
R22384 plus.n54 plus.t10 415.966
R22385 plus.n37 plus.t19 415.966
R22386 plus.n59 plus.t8 415.966
R22387 plus.n35 plus.t16 415.966
R22388 plus.n64 plus.t28 415.966
R22389 plus.n66 plus.t21 415.966
R22390 plus.n32 plus.t23 415.966
R22391 plus.n30 plus.t13 415.966
R22392 plus.n29 plus.t27 415.966
R22393 plus.n3 plus.t22 415.966
R22394 plus.n23 plus.t7 415.966
R22395 plus.n22 plus.t18 415.966
R22396 plus.n6 plus.t14 415.966
R22397 plus.n17 plus.t24 415.966
R22398 plus.n15 plus.t17 415.966
R22399 plus.n9 plus.t9 415.966
R22400 plus.n10 plus.t15 415.966
R22401 plus.n70 plus.t3 243.97
R22402 plus.n70 plus.n69 223.454
R22403 plus.n72 plus.n71 223.454
R22404 plus.n67 plus.n66 161.3
R22405 plus.n65 plus.n34 161.3
R22406 plus.n64 plus.n63 161.3
R22407 plus.n62 plus.n35 161.3
R22408 plus.n61 plus.n60 161.3
R22409 plus.n59 plus.n36 161.3
R22410 plus.n58 plus.n57 161.3
R22411 plus.n56 plus.n37 161.3
R22412 plus.n55 plus.n54 161.3
R22413 plus.n53 plus.n38 161.3
R22414 plus.n52 plus.n51 161.3
R22415 plus.n50 plus.n39 161.3
R22416 plus.n49 plus.n48 161.3
R22417 plus.n47 plus.n40 161.3
R22418 plus.n46 plus.n45 161.3
R22419 plus.n44 plus.n41 161.3
R22420 plus.n12 plus.n9 161.3
R22421 plus.n14 plus.n13 161.3
R22422 plus.n15 plus.n8 161.3
R22423 plus.n16 plus.n7 161.3
R22424 plus.n18 plus.n17 161.3
R22425 plus.n19 plus.n6 161.3
R22426 plus.n21 plus.n20 161.3
R22427 plus.n22 plus.n5 161.3
R22428 plus.n23 plus.n4 161.3
R22429 plus.n25 plus.n24 161.3
R22430 plus.n26 plus.n3 161.3
R22431 plus.n28 plus.n27 161.3
R22432 plus.n29 plus.n2 161.3
R22433 plus.n30 plus.n1 161.3
R22434 plus.n31 plus.n0 161.3
R22435 plus.n33 plus.n32 161.3
R22436 plus.n42 plus.n41 48.2005
R22437 plus.n52 plus.n39 48.2005
R22438 plus.n54 plus.n37 48.2005
R22439 plus.n64 plus.n35 48.2005
R22440 plus.n30 plus.n29 48.2005
R22441 plus.n23 plus.n22 48.2005
R22442 plus.n17 plus.n6 48.2005
R22443 plus.n10 plus.n9 48.2005
R22444 plus.n48 plus.n47 47.4702
R22445 plus.n59 plus.n58 47.4702
R22446 plus.n24 plus.n3 47.4702
R22447 plus.n16 plus.n15 47.4702
R22448 plus.n66 plus.n65 46.0096
R22449 plus.n32 plus.n31 46.0096
R22450 plus.n44 plus.n43 45.0871
R22451 plus.n12 plus.n11 45.0871
R22452 plus.n68 plus.n67 31.0554
R22453 plus.n47 plus.n46 25.5611
R22454 plus.n60 plus.n59 25.5611
R22455 plus.n28 plus.n3 25.5611
R22456 plus.n15 plus.n14 25.5611
R22457 plus.n53 plus.n52 24.1005
R22458 plus.n54 plus.n53 24.1005
R22459 plus.n22 plus.n21 24.1005
R22460 plus.n21 plus.n6 24.1005
R22461 plus.n46 plus.n41 22.6399
R22462 plus.n60 plus.n35 22.6399
R22463 plus.n29 plus.n28 22.6399
R22464 plus.n14 plus.n9 22.6399
R22465 plus.n69 plus.t4 19.8005
R22466 plus.n69 plus.t1 19.8005
R22467 plus.n71 plus.t0 19.8005
R22468 plus.n71 plus.t2 19.8005
R22469 plus plus.n73 14.3678
R22470 plus.n43 plus.n42 14.1472
R22471 plus.n11 plus.n10 14.1472
R22472 plus.n68 plus.n33 11.7259
R22473 plus.n73 plus.n72 5.40567
R22474 plus.n65 plus.n64 2.19141
R22475 plus.n31 plus.n30 2.19141
R22476 plus.n73 plus.n68 1.188
R22477 plus.n48 plus.n39 0.730803
R22478 plus.n58 plus.n37 0.730803
R22479 plus.n24 plus.n23 0.730803
R22480 plus.n17 plus.n16 0.730803
R22481 plus.n72 plus.n70 0.716017
R22482 plus.n45 plus.n44 0.189894
R22483 plus.n45 plus.n40 0.189894
R22484 plus.n49 plus.n40 0.189894
R22485 plus.n50 plus.n49 0.189894
R22486 plus.n51 plus.n50 0.189894
R22487 plus.n51 plus.n38 0.189894
R22488 plus.n55 plus.n38 0.189894
R22489 plus.n56 plus.n55 0.189894
R22490 plus.n57 plus.n56 0.189894
R22491 plus.n57 plus.n36 0.189894
R22492 plus.n61 plus.n36 0.189894
R22493 plus.n62 plus.n61 0.189894
R22494 plus.n63 plus.n62 0.189894
R22495 plus.n63 plus.n34 0.189894
R22496 plus.n67 plus.n34 0.189894
R22497 plus.n33 plus.n0 0.189894
R22498 plus.n1 plus.n0 0.189894
R22499 plus.n2 plus.n1 0.189894
R22500 plus.n27 plus.n2 0.189894
R22501 plus.n27 plus.n26 0.189894
R22502 plus.n26 plus.n25 0.189894
R22503 plus.n25 plus.n4 0.189894
R22504 plus.n5 plus.n4 0.189894
R22505 plus.n20 plus.n5 0.189894
R22506 plus.n20 plus.n19 0.189894
R22507 plus.n19 plus.n18 0.189894
R22508 plus.n18 plus.n7 0.189894
R22509 plus.n8 plus.n7 0.189894
R22510 plus.n13 plus.n8 0.189894
R22511 plus.n13 plus.n12 0.189894
R22512 minus.n45 minus.t26 442.325
R22513 minus.n9 minus.t12 442.325
R22514 minus.n66 minus.t16 415.966
R22515 minus.n64 minus.t28 415.966
R22516 minus.n63 minus.t21 415.966
R22517 minus.n37 minus.t14 415.966
R22518 minus.n57 minus.t23 415.966
R22519 minus.n56 minus.t11 415.966
R22520 minus.n40 minus.t5 415.966
R22521 minus.n51 minus.t17 415.966
R22522 minus.n49 minus.t10 415.966
R22523 minus.n43 minus.t25 415.966
R22524 minus.n44 minus.t7 415.966
R22525 minus.n8 minus.t18 415.966
R22526 minus.n7 minus.t8 415.966
R22527 minus.n13 minus.t13 415.966
R22528 minus.n5 minus.t24 415.966
R22529 minus.n18 minus.t19 415.966
R22530 minus.n20 minus.t22 415.966
R22531 minus.n3 minus.t6 415.966
R22532 minus.n25 minus.t20 415.966
R22533 minus.n1 minus.t27 415.966
R22534 minus.n30 minus.t15 415.966
R22535 minus.n32 minus.t9 415.966
R22536 minus.n72 minus.t3 243.255
R22537 minus.n71 minus.n69 224.169
R22538 minus.n71 minus.n70 223.454
R22539 minus.n46 minus.n43 161.3
R22540 minus.n48 minus.n47 161.3
R22541 minus.n49 minus.n42 161.3
R22542 minus.n50 minus.n41 161.3
R22543 minus.n52 minus.n51 161.3
R22544 minus.n53 minus.n40 161.3
R22545 minus.n55 minus.n54 161.3
R22546 minus.n56 minus.n39 161.3
R22547 minus.n57 minus.n38 161.3
R22548 minus.n59 minus.n58 161.3
R22549 minus.n60 minus.n37 161.3
R22550 minus.n62 minus.n61 161.3
R22551 minus.n63 minus.n36 161.3
R22552 minus.n64 minus.n35 161.3
R22553 minus.n65 minus.n34 161.3
R22554 minus.n67 minus.n66 161.3
R22555 minus.n33 minus.n32 161.3
R22556 minus.n31 minus.n0 161.3
R22557 minus.n30 minus.n29 161.3
R22558 minus.n28 minus.n1 161.3
R22559 minus.n27 minus.n26 161.3
R22560 minus.n25 minus.n2 161.3
R22561 minus.n24 minus.n23 161.3
R22562 minus.n22 minus.n3 161.3
R22563 minus.n21 minus.n20 161.3
R22564 minus.n19 minus.n4 161.3
R22565 minus.n18 minus.n17 161.3
R22566 minus.n16 minus.n5 161.3
R22567 minus.n15 minus.n14 161.3
R22568 minus.n13 minus.n6 161.3
R22569 minus.n12 minus.n11 161.3
R22570 minus.n10 minus.n7 161.3
R22571 minus.n64 minus.n63 48.2005
R22572 minus.n57 minus.n56 48.2005
R22573 minus.n51 minus.n40 48.2005
R22574 minus.n44 minus.n43 48.2005
R22575 minus.n8 minus.n7 48.2005
R22576 minus.n18 minus.n5 48.2005
R22577 minus.n20 minus.n3 48.2005
R22578 minus.n30 minus.n1 48.2005
R22579 minus.n58 minus.n37 47.4702
R22580 minus.n50 minus.n49 47.4702
R22581 minus.n14 minus.n13 47.4702
R22582 minus.n25 minus.n24 47.4702
R22583 minus.n66 minus.n65 46.0096
R22584 minus.n32 minus.n31 46.0096
R22585 minus.n10 minus.n9 45.0871
R22586 minus.n46 minus.n45 45.0871
R22587 minus.n68 minus.n67 31.2713
R22588 minus.n62 minus.n37 25.5611
R22589 minus.n49 minus.n48 25.5611
R22590 minus.n13 minus.n12 25.5611
R22591 minus.n26 minus.n25 25.5611
R22592 minus.n56 minus.n55 24.1005
R22593 minus.n55 minus.n40 24.1005
R22594 minus.n19 minus.n18 24.1005
R22595 minus.n20 minus.n19 24.1005
R22596 minus.n63 minus.n62 22.6399
R22597 minus.n48 minus.n43 22.6399
R22598 minus.n12 minus.n7 22.6399
R22599 minus.n26 minus.n1 22.6399
R22600 minus.n70 minus.t2 19.8005
R22601 minus.n70 minus.t0 19.8005
R22602 minus.n69 minus.t1 19.8005
R22603 minus.n69 minus.t4 19.8005
R22604 minus.n45 minus.n44 14.1472
R22605 minus.n9 minus.n8 14.1472
R22606 minus.n68 minus.n33 11.9418
R22607 minus minus.n73 11.5306
R22608 minus.n73 minus.n72 4.80222
R22609 minus.n65 minus.n64 2.19141
R22610 minus.n31 minus.n30 2.19141
R22611 minus.n73 minus.n68 0.972091
R22612 minus.n58 minus.n57 0.730803
R22613 minus.n51 minus.n50 0.730803
R22614 minus.n14 minus.n5 0.730803
R22615 minus.n24 minus.n3 0.730803
R22616 minus.n72 minus.n71 0.716017
R22617 minus.n67 minus.n34 0.189894
R22618 minus.n35 minus.n34 0.189894
R22619 minus.n36 minus.n35 0.189894
R22620 minus.n61 minus.n36 0.189894
R22621 minus.n61 minus.n60 0.189894
R22622 minus.n60 minus.n59 0.189894
R22623 minus.n59 minus.n38 0.189894
R22624 minus.n39 minus.n38 0.189894
R22625 minus.n54 minus.n39 0.189894
R22626 minus.n54 minus.n53 0.189894
R22627 minus.n53 minus.n52 0.189894
R22628 minus.n52 minus.n41 0.189894
R22629 minus.n42 minus.n41 0.189894
R22630 minus.n47 minus.n42 0.189894
R22631 minus.n47 minus.n46 0.189894
R22632 minus.n11 minus.n10 0.189894
R22633 minus.n11 minus.n6 0.189894
R22634 minus.n15 minus.n6 0.189894
R22635 minus.n16 minus.n15 0.189894
R22636 minus.n17 minus.n16 0.189894
R22637 minus.n17 minus.n4 0.189894
R22638 minus.n21 minus.n4 0.189894
R22639 minus.n22 minus.n21 0.189894
R22640 minus.n23 minus.n22 0.189894
R22641 minus.n23 minus.n2 0.189894
R22642 minus.n27 minus.n2 0.189894
R22643 minus.n28 minus.n27 0.189894
R22644 minus.n29 minus.n28 0.189894
R22645 minus.n29 minus.n0 0.189894
R22646 minus.n33 minus.n0 0.189894
R22647 outputibias.n27 outputibias.n1 289.615
R22648 outputibias.n58 outputibias.n32 289.615
R22649 outputibias.n90 outputibias.n64 289.615
R22650 outputibias.n122 outputibias.n96 289.615
R22651 outputibias.n28 outputibias.n27 185
R22652 outputibias.n26 outputibias.n25 185
R22653 outputibias.n5 outputibias.n4 185
R22654 outputibias.n20 outputibias.n19 185
R22655 outputibias.n18 outputibias.n17 185
R22656 outputibias.n9 outputibias.n8 185
R22657 outputibias.n12 outputibias.n11 185
R22658 outputibias.n59 outputibias.n58 185
R22659 outputibias.n57 outputibias.n56 185
R22660 outputibias.n36 outputibias.n35 185
R22661 outputibias.n51 outputibias.n50 185
R22662 outputibias.n49 outputibias.n48 185
R22663 outputibias.n40 outputibias.n39 185
R22664 outputibias.n43 outputibias.n42 185
R22665 outputibias.n91 outputibias.n90 185
R22666 outputibias.n89 outputibias.n88 185
R22667 outputibias.n68 outputibias.n67 185
R22668 outputibias.n83 outputibias.n82 185
R22669 outputibias.n81 outputibias.n80 185
R22670 outputibias.n72 outputibias.n71 185
R22671 outputibias.n75 outputibias.n74 185
R22672 outputibias.n123 outputibias.n122 185
R22673 outputibias.n121 outputibias.n120 185
R22674 outputibias.n100 outputibias.n99 185
R22675 outputibias.n115 outputibias.n114 185
R22676 outputibias.n113 outputibias.n112 185
R22677 outputibias.n104 outputibias.n103 185
R22678 outputibias.n107 outputibias.n106 185
R22679 outputibias.n0 outputibias.t10 178.945
R22680 outputibias.n133 outputibias.t8 177.018
R22681 outputibias.n132 outputibias.t11 177.018
R22682 outputibias.n0 outputibias.t9 177.018
R22683 outputibias.t7 outputibias.n10 147.661
R22684 outputibias.t1 outputibias.n41 147.661
R22685 outputibias.t3 outputibias.n73 147.661
R22686 outputibias.t5 outputibias.n105 147.661
R22687 outputibias.n128 outputibias.t6 132.363
R22688 outputibias.n128 outputibias.t0 130.436
R22689 outputibias.n129 outputibias.t2 130.436
R22690 outputibias.n130 outputibias.t4 130.436
R22691 outputibias.n27 outputibias.n26 104.615
R22692 outputibias.n26 outputibias.n4 104.615
R22693 outputibias.n19 outputibias.n4 104.615
R22694 outputibias.n19 outputibias.n18 104.615
R22695 outputibias.n18 outputibias.n8 104.615
R22696 outputibias.n11 outputibias.n8 104.615
R22697 outputibias.n58 outputibias.n57 104.615
R22698 outputibias.n57 outputibias.n35 104.615
R22699 outputibias.n50 outputibias.n35 104.615
R22700 outputibias.n50 outputibias.n49 104.615
R22701 outputibias.n49 outputibias.n39 104.615
R22702 outputibias.n42 outputibias.n39 104.615
R22703 outputibias.n90 outputibias.n89 104.615
R22704 outputibias.n89 outputibias.n67 104.615
R22705 outputibias.n82 outputibias.n67 104.615
R22706 outputibias.n82 outputibias.n81 104.615
R22707 outputibias.n81 outputibias.n71 104.615
R22708 outputibias.n74 outputibias.n71 104.615
R22709 outputibias.n122 outputibias.n121 104.615
R22710 outputibias.n121 outputibias.n99 104.615
R22711 outputibias.n114 outputibias.n99 104.615
R22712 outputibias.n114 outputibias.n113 104.615
R22713 outputibias.n113 outputibias.n103 104.615
R22714 outputibias.n106 outputibias.n103 104.615
R22715 outputibias.n63 outputibias.n31 95.6354
R22716 outputibias.n63 outputibias.n62 94.6732
R22717 outputibias.n95 outputibias.n94 94.6732
R22718 outputibias.n127 outputibias.n126 94.6732
R22719 outputibias.n11 outputibias.t7 52.3082
R22720 outputibias.n42 outputibias.t1 52.3082
R22721 outputibias.n74 outputibias.t3 52.3082
R22722 outputibias.n106 outputibias.t5 52.3082
R22723 outputibias.n12 outputibias.n10 15.6674
R22724 outputibias.n43 outputibias.n41 15.6674
R22725 outputibias.n75 outputibias.n73 15.6674
R22726 outputibias.n107 outputibias.n105 15.6674
R22727 outputibias.n13 outputibias.n9 12.8005
R22728 outputibias.n44 outputibias.n40 12.8005
R22729 outputibias.n76 outputibias.n72 12.8005
R22730 outputibias.n108 outputibias.n104 12.8005
R22731 outputibias.n17 outputibias.n16 12.0247
R22732 outputibias.n48 outputibias.n47 12.0247
R22733 outputibias.n80 outputibias.n79 12.0247
R22734 outputibias.n112 outputibias.n111 12.0247
R22735 outputibias.n20 outputibias.n7 11.249
R22736 outputibias.n51 outputibias.n38 11.249
R22737 outputibias.n83 outputibias.n70 11.249
R22738 outputibias.n115 outputibias.n102 11.249
R22739 outputibias.n21 outputibias.n5 10.4732
R22740 outputibias.n52 outputibias.n36 10.4732
R22741 outputibias.n84 outputibias.n68 10.4732
R22742 outputibias.n116 outputibias.n100 10.4732
R22743 outputibias.n25 outputibias.n24 9.69747
R22744 outputibias.n56 outputibias.n55 9.69747
R22745 outputibias.n88 outputibias.n87 9.69747
R22746 outputibias.n120 outputibias.n119 9.69747
R22747 outputibias.n31 outputibias.n30 9.45567
R22748 outputibias.n62 outputibias.n61 9.45567
R22749 outputibias.n94 outputibias.n93 9.45567
R22750 outputibias.n126 outputibias.n125 9.45567
R22751 outputibias.n30 outputibias.n29 9.3005
R22752 outputibias.n3 outputibias.n2 9.3005
R22753 outputibias.n24 outputibias.n23 9.3005
R22754 outputibias.n22 outputibias.n21 9.3005
R22755 outputibias.n7 outputibias.n6 9.3005
R22756 outputibias.n16 outputibias.n15 9.3005
R22757 outputibias.n14 outputibias.n13 9.3005
R22758 outputibias.n61 outputibias.n60 9.3005
R22759 outputibias.n34 outputibias.n33 9.3005
R22760 outputibias.n55 outputibias.n54 9.3005
R22761 outputibias.n53 outputibias.n52 9.3005
R22762 outputibias.n38 outputibias.n37 9.3005
R22763 outputibias.n47 outputibias.n46 9.3005
R22764 outputibias.n45 outputibias.n44 9.3005
R22765 outputibias.n93 outputibias.n92 9.3005
R22766 outputibias.n66 outputibias.n65 9.3005
R22767 outputibias.n87 outputibias.n86 9.3005
R22768 outputibias.n85 outputibias.n84 9.3005
R22769 outputibias.n70 outputibias.n69 9.3005
R22770 outputibias.n79 outputibias.n78 9.3005
R22771 outputibias.n77 outputibias.n76 9.3005
R22772 outputibias.n125 outputibias.n124 9.3005
R22773 outputibias.n98 outputibias.n97 9.3005
R22774 outputibias.n119 outputibias.n118 9.3005
R22775 outputibias.n117 outputibias.n116 9.3005
R22776 outputibias.n102 outputibias.n101 9.3005
R22777 outputibias.n111 outputibias.n110 9.3005
R22778 outputibias.n109 outputibias.n108 9.3005
R22779 outputibias.n28 outputibias.n3 8.92171
R22780 outputibias.n59 outputibias.n34 8.92171
R22781 outputibias.n91 outputibias.n66 8.92171
R22782 outputibias.n123 outputibias.n98 8.92171
R22783 outputibias.n29 outputibias.n1 8.14595
R22784 outputibias.n60 outputibias.n32 8.14595
R22785 outputibias.n92 outputibias.n64 8.14595
R22786 outputibias.n124 outputibias.n96 8.14595
R22787 outputibias.n31 outputibias.n1 5.81868
R22788 outputibias.n62 outputibias.n32 5.81868
R22789 outputibias.n94 outputibias.n64 5.81868
R22790 outputibias.n126 outputibias.n96 5.81868
R22791 outputibias.n131 outputibias.n130 5.20947
R22792 outputibias.n29 outputibias.n28 5.04292
R22793 outputibias.n60 outputibias.n59 5.04292
R22794 outputibias.n92 outputibias.n91 5.04292
R22795 outputibias.n124 outputibias.n123 5.04292
R22796 outputibias.n131 outputibias.n127 4.42209
R22797 outputibias.n14 outputibias.n10 4.38594
R22798 outputibias.n45 outputibias.n41 4.38594
R22799 outputibias.n77 outputibias.n73 4.38594
R22800 outputibias.n109 outputibias.n105 4.38594
R22801 outputibias.n132 outputibias.n131 4.28454
R22802 outputibias.n25 outputibias.n3 4.26717
R22803 outputibias.n56 outputibias.n34 4.26717
R22804 outputibias.n88 outputibias.n66 4.26717
R22805 outputibias.n120 outputibias.n98 4.26717
R22806 outputibias.n24 outputibias.n5 3.49141
R22807 outputibias.n55 outputibias.n36 3.49141
R22808 outputibias.n87 outputibias.n68 3.49141
R22809 outputibias.n119 outputibias.n100 3.49141
R22810 outputibias.n21 outputibias.n20 2.71565
R22811 outputibias.n52 outputibias.n51 2.71565
R22812 outputibias.n84 outputibias.n83 2.71565
R22813 outputibias.n116 outputibias.n115 2.71565
R22814 outputibias.n17 outputibias.n7 1.93989
R22815 outputibias.n48 outputibias.n38 1.93989
R22816 outputibias.n80 outputibias.n70 1.93989
R22817 outputibias.n112 outputibias.n102 1.93989
R22818 outputibias.n130 outputibias.n129 1.9266
R22819 outputibias.n129 outputibias.n128 1.9266
R22820 outputibias.n133 outputibias.n132 1.92658
R22821 outputibias.n134 outputibias.n133 1.29913
R22822 outputibias.n16 outputibias.n9 1.16414
R22823 outputibias.n47 outputibias.n40 1.16414
R22824 outputibias.n79 outputibias.n72 1.16414
R22825 outputibias.n111 outputibias.n104 1.16414
R22826 outputibias.n127 outputibias.n95 0.962709
R22827 outputibias.n95 outputibias.n63 0.962709
R22828 outputibias.n13 outputibias.n12 0.388379
R22829 outputibias.n44 outputibias.n43 0.388379
R22830 outputibias.n76 outputibias.n75 0.388379
R22831 outputibias.n108 outputibias.n107 0.388379
R22832 outputibias.n134 outputibias.n0 0.337251
R22833 outputibias outputibias.n134 0.302375
R22834 outputibias.n30 outputibias.n2 0.155672
R22835 outputibias.n23 outputibias.n2 0.155672
R22836 outputibias.n23 outputibias.n22 0.155672
R22837 outputibias.n22 outputibias.n6 0.155672
R22838 outputibias.n15 outputibias.n6 0.155672
R22839 outputibias.n15 outputibias.n14 0.155672
R22840 outputibias.n61 outputibias.n33 0.155672
R22841 outputibias.n54 outputibias.n33 0.155672
R22842 outputibias.n54 outputibias.n53 0.155672
R22843 outputibias.n53 outputibias.n37 0.155672
R22844 outputibias.n46 outputibias.n37 0.155672
R22845 outputibias.n46 outputibias.n45 0.155672
R22846 outputibias.n93 outputibias.n65 0.155672
R22847 outputibias.n86 outputibias.n65 0.155672
R22848 outputibias.n86 outputibias.n85 0.155672
R22849 outputibias.n85 outputibias.n69 0.155672
R22850 outputibias.n78 outputibias.n69 0.155672
R22851 outputibias.n78 outputibias.n77 0.155672
R22852 outputibias.n125 outputibias.n97 0.155672
R22853 outputibias.n118 outputibias.n97 0.155672
R22854 outputibias.n118 outputibias.n117 0.155672
R22855 outputibias.n117 outputibias.n101 0.155672
R22856 outputibias.n110 outputibias.n101 0.155672
R22857 outputibias.n110 outputibias.n109 0.155672
R22858 output.n41 output.n15 289.615
R22859 output.n72 output.n46 289.615
R22860 output.n104 output.n78 289.615
R22861 output.n136 output.n110 289.615
R22862 output.n77 output.n45 197.26
R22863 output.n77 output.n76 196.298
R22864 output.n109 output.n108 196.298
R22865 output.n141 output.n140 196.298
R22866 output.n42 output.n41 185
R22867 output.n40 output.n39 185
R22868 output.n19 output.n18 185
R22869 output.n34 output.n33 185
R22870 output.n32 output.n31 185
R22871 output.n23 output.n22 185
R22872 output.n26 output.n25 185
R22873 output.n73 output.n72 185
R22874 output.n71 output.n70 185
R22875 output.n50 output.n49 185
R22876 output.n65 output.n64 185
R22877 output.n63 output.n62 185
R22878 output.n54 output.n53 185
R22879 output.n57 output.n56 185
R22880 output.n105 output.n104 185
R22881 output.n103 output.n102 185
R22882 output.n82 output.n81 185
R22883 output.n97 output.n96 185
R22884 output.n95 output.n94 185
R22885 output.n86 output.n85 185
R22886 output.n89 output.n88 185
R22887 output.n137 output.n136 185
R22888 output.n135 output.n134 185
R22889 output.n114 output.n113 185
R22890 output.n129 output.n128 185
R22891 output.n127 output.n126 185
R22892 output.n118 output.n117 185
R22893 output.n121 output.n120 185
R22894 output.t17 output.n24 147.661
R22895 output.t18 output.n55 147.661
R22896 output.t19 output.n87 147.661
R22897 output.t16 output.n119 147.661
R22898 output.n41 output.n40 104.615
R22899 output.n40 output.n18 104.615
R22900 output.n33 output.n18 104.615
R22901 output.n33 output.n32 104.615
R22902 output.n32 output.n22 104.615
R22903 output.n25 output.n22 104.615
R22904 output.n72 output.n71 104.615
R22905 output.n71 output.n49 104.615
R22906 output.n64 output.n49 104.615
R22907 output.n64 output.n63 104.615
R22908 output.n63 output.n53 104.615
R22909 output.n56 output.n53 104.615
R22910 output.n104 output.n103 104.615
R22911 output.n103 output.n81 104.615
R22912 output.n96 output.n81 104.615
R22913 output.n96 output.n95 104.615
R22914 output.n95 output.n85 104.615
R22915 output.n88 output.n85 104.615
R22916 output.n136 output.n135 104.615
R22917 output.n135 output.n113 104.615
R22918 output.n128 output.n113 104.615
R22919 output.n128 output.n127 104.615
R22920 output.n127 output.n117 104.615
R22921 output.n120 output.n117 104.615
R22922 output.n1 output.t1 77.056
R22923 output.n14 output.t3 76.6694
R22924 output.n1 output.n0 72.7095
R22925 output.n3 output.n2 72.7095
R22926 output.n5 output.n4 72.7095
R22927 output.n7 output.n6 72.7095
R22928 output.n9 output.n8 72.7095
R22929 output.n11 output.n10 72.7095
R22930 output.n13 output.n12 72.7095
R22931 output.n25 output.t17 52.3082
R22932 output.n56 output.t18 52.3082
R22933 output.n88 output.t19 52.3082
R22934 output.n120 output.t16 52.3082
R22935 output.n26 output.n24 15.6674
R22936 output.n57 output.n55 15.6674
R22937 output.n89 output.n87 15.6674
R22938 output.n121 output.n119 15.6674
R22939 output.n27 output.n23 12.8005
R22940 output.n58 output.n54 12.8005
R22941 output.n90 output.n86 12.8005
R22942 output.n122 output.n118 12.8005
R22943 output.n31 output.n30 12.0247
R22944 output.n62 output.n61 12.0247
R22945 output.n94 output.n93 12.0247
R22946 output.n126 output.n125 12.0247
R22947 output.n34 output.n21 11.249
R22948 output.n65 output.n52 11.249
R22949 output.n97 output.n84 11.249
R22950 output.n129 output.n116 11.249
R22951 output.n35 output.n19 10.4732
R22952 output.n66 output.n50 10.4732
R22953 output.n98 output.n82 10.4732
R22954 output.n130 output.n114 10.4732
R22955 output.n39 output.n38 9.69747
R22956 output.n70 output.n69 9.69747
R22957 output.n102 output.n101 9.69747
R22958 output.n134 output.n133 9.69747
R22959 output.n45 output.n44 9.45567
R22960 output.n76 output.n75 9.45567
R22961 output.n108 output.n107 9.45567
R22962 output.n140 output.n139 9.45567
R22963 output.n44 output.n43 9.3005
R22964 output.n17 output.n16 9.3005
R22965 output.n38 output.n37 9.3005
R22966 output.n36 output.n35 9.3005
R22967 output.n21 output.n20 9.3005
R22968 output.n30 output.n29 9.3005
R22969 output.n28 output.n27 9.3005
R22970 output.n75 output.n74 9.3005
R22971 output.n48 output.n47 9.3005
R22972 output.n69 output.n68 9.3005
R22973 output.n67 output.n66 9.3005
R22974 output.n52 output.n51 9.3005
R22975 output.n61 output.n60 9.3005
R22976 output.n59 output.n58 9.3005
R22977 output.n107 output.n106 9.3005
R22978 output.n80 output.n79 9.3005
R22979 output.n101 output.n100 9.3005
R22980 output.n99 output.n98 9.3005
R22981 output.n84 output.n83 9.3005
R22982 output.n93 output.n92 9.3005
R22983 output.n91 output.n90 9.3005
R22984 output.n139 output.n138 9.3005
R22985 output.n112 output.n111 9.3005
R22986 output.n133 output.n132 9.3005
R22987 output.n131 output.n130 9.3005
R22988 output.n116 output.n115 9.3005
R22989 output.n125 output.n124 9.3005
R22990 output.n123 output.n122 9.3005
R22991 output.n42 output.n17 8.92171
R22992 output.n73 output.n48 8.92171
R22993 output.n105 output.n80 8.92171
R22994 output.n137 output.n112 8.92171
R22995 output output.n141 8.15037
R22996 output.n43 output.n15 8.14595
R22997 output.n74 output.n46 8.14595
R22998 output.n106 output.n78 8.14595
R22999 output.n138 output.n110 8.14595
R23000 output.n45 output.n15 5.81868
R23001 output.n76 output.n46 5.81868
R23002 output.n108 output.n78 5.81868
R23003 output.n140 output.n110 5.81868
R23004 output.n43 output.n42 5.04292
R23005 output.n74 output.n73 5.04292
R23006 output.n106 output.n105 5.04292
R23007 output.n138 output.n137 5.04292
R23008 output.n28 output.n24 4.38594
R23009 output.n59 output.n55 4.38594
R23010 output.n91 output.n87 4.38594
R23011 output.n123 output.n119 4.38594
R23012 output.n39 output.n17 4.26717
R23013 output.n70 output.n48 4.26717
R23014 output.n102 output.n80 4.26717
R23015 output.n134 output.n112 4.26717
R23016 output.n0 output.t12 3.9605
R23017 output.n0 output.t15 3.9605
R23018 output.n2 output.t5 3.9605
R23019 output.n2 output.t4 3.9605
R23020 output.n4 output.t10 3.9605
R23021 output.n4 output.t14 3.9605
R23022 output.n6 output.t2 3.9605
R23023 output.n6 output.t6 3.9605
R23024 output.n8 output.t7 3.9605
R23025 output.n8 output.t13 3.9605
R23026 output.n10 output.t0 3.9605
R23027 output.n10 output.t8 3.9605
R23028 output.n12 output.t11 3.9605
R23029 output.n12 output.t9 3.9605
R23030 output.n38 output.n19 3.49141
R23031 output.n69 output.n50 3.49141
R23032 output.n101 output.n82 3.49141
R23033 output.n133 output.n114 3.49141
R23034 output.n35 output.n34 2.71565
R23035 output.n66 output.n65 2.71565
R23036 output.n98 output.n97 2.71565
R23037 output.n130 output.n129 2.71565
R23038 output.n31 output.n21 1.93989
R23039 output.n62 output.n52 1.93989
R23040 output.n94 output.n84 1.93989
R23041 output.n126 output.n116 1.93989
R23042 output.n30 output.n23 1.16414
R23043 output.n61 output.n54 1.16414
R23044 output.n93 output.n86 1.16414
R23045 output.n125 output.n118 1.16414
R23046 output.n141 output.n109 0.962709
R23047 output.n109 output.n77 0.962709
R23048 output.n27 output.n26 0.388379
R23049 output.n58 output.n57 0.388379
R23050 output.n90 output.n89 0.388379
R23051 output.n122 output.n121 0.388379
R23052 output.n14 output.n13 0.387128
R23053 output.n13 output.n11 0.387128
R23054 output.n11 output.n9 0.387128
R23055 output.n9 output.n7 0.387128
R23056 output.n7 output.n5 0.387128
R23057 output.n5 output.n3 0.387128
R23058 output.n3 output.n1 0.387128
R23059 output.n44 output.n16 0.155672
R23060 output.n37 output.n16 0.155672
R23061 output.n37 output.n36 0.155672
R23062 output.n36 output.n20 0.155672
R23063 output.n29 output.n20 0.155672
R23064 output.n29 output.n28 0.155672
R23065 output.n75 output.n47 0.155672
R23066 output.n68 output.n47 0.155672
R23067 output.n68 output.n67 0.155672
R23068 output.n67 output.n51 0.155672
R23069 output.n60 output.n51 0.155672
R23070 output.n60 output.n59 0.155672
R23071 output.n107 output.n79 0.155672
R23072 output.n100 output.n79 0.155672
R23073 output.n100 output.n99 0.155672
R23074 output.n99 output.n83 0.155672
R23075 output.n92 output.n83 0.155672
R23076 output.n92 output.n91 0.155672
R23077 output.n139 output.n111 0.155672
R23078 output.n132 output.n111 0.155672
R23079 output.n132 output.n131 0.155672
R23080 output.n131 output.n115 0.155672
R23081 output.n124 output.n115 0.155672
R23082 output.n124 output.n123 0.155672
R23083 output output.n14 0.126227
C0 minus commonsourceibias 0.331305f
C1 plus commonsourceibias 0.276969f
C2 output outputibias 2.34152f
C3 vdd output 7.23429f
C4 CSoutput output 6.13881f
C5 CSoutput outputibias 0.032386f
C6 vdd CSoutput 92.9691f
C7 minus diffpairibias 2.98e-19
C8 commonsourceibias output 0.006808f
C9 CSoutput minus 2.75386f
C10 vdd plus 0.084873f
C11 commonsourceibias outputibias 0.003832f
C12 plus diffpairibias 2.75e-19
C13 vdd commonsourceibias 0.004218f
C14 CSoutput plus 0.852171f
C15 commonsourceibias diffpairibias 0.064336f
C16 CSoutput commonsourceibias 42.3358f
C17 minus plus 9.09051f
C18 diffpairibias gnd 60.00273f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.14503p
C22 plus gnd 33.1377f
C23 minus gnd 27.462212f
C24 CSoutput gnd 0.1075p
C25 vdd gnd 0.479853p
C26 output.t1 gnd 0.464308f
C27 output.t12 gnd 0.044422f
C28 output.t15 gnd 0.044422f
C29 output.n0 gnd 0.364624f
C30 output.n1 gnd 0.614102f
C31 output.t5 gnd 0.044422f
C32 output.t4 gnd 0.044422f
C33 output.n2 gnd 0.364624f
C34 output.n3 gnd 0.350265f
C35 output.t10 gnd 0.044422f
C36 output.t14 gnd 0.044422f
C37 output.n4 gnd 0.364624f
C38 output.n5 gnd 0.350265f
C39 output.t2 gnd 0.044422f
C40 output.t6 gnd 0.044422f
C41 output.n6 gnd 0.364624f
C42 output.n7 gnd 0.350265f
C43 output.t7 gnd 0.044422f
C44 output.t13 gnd 0.044422f
C45 output.n8 gnd 0.364624f
C46 output.n9 gnd 0.350265f
C47 output.t0 gnd 0.044422f
C48 output.t8 gnd 0.044422f
C49 output.n10 gnd 0.364624f
C50 output.n11 gnd 0.350265f
C51 output.t11 gnd 0.044422f
C52 output.t9 gnd 0.044422f
C53 output.n12 gnd 0.364624f
C54 output.n13 gnd 0.350265f
C55 output.t3 gnd 0.462979f
C56 output.n14 gnd 0.28994f
C57 output.n15 gnd 0.015803f
C58 output.n16 gnd 0.011243f
C59 output.n17 gnd 0.006041f
C60 output.n18 gnd 0.01428f
C61 output.n19 gnd 0.006397f
C62 output.n20 gnd 0.011243f
C63 output.n21 gnd 0.006041f
C64 output.n22 gnd 0.01428f
C65 output.n23 gnd 0.006397f
C66 output.n24 gnd 0.048111f
C67 output.t17 gnd 0.023274f
C68 output.n25 gnd 0.01071f
C69 output.n26 gnd 0.008435f
C70 output.n27 gnd 0.006041f
C71 output.n28 gnd 0.267512f
C72 output.n29 gnd 0.011243f
C73 output.n30 gnd 0.006041f
C74 output.n31 gnd 0.006397f
C75 output.n32 gnd 0.01428f
C76 output.n33 gnd 0.01428f
C77 output.n34 gnd 0.006397f
C78 output.n35 gnd 0.006041f
C79 output.n36 gnd 0.011243f
C80 output.n37 gnd 0.011243f
C81 output.n38 gnd 0.006041f
C82 output.n39 gnd 0.006397f
C83 output.n40 gnd 0.01428f
C84 output.n41 gnd 0.030913f
C85 output.n42 gnd 0.006397f
C86 output.n43 gnd 0.006041f
C87 output.n44 gnd 0.025987f
C88 output.n45 gnd 0.097665f
C89 output.n46 gnd 0.015803f
C90 output.n47 gnd 0.011243f
C91 output.n48 gnd 0.006041f
C92 output.n49 gnd 0.01428f
C93 output.n50 gnd 0.006397f
C94 output.n51 gnd 0.011243f
C95 output.n52 gnd 0.006041f
C96 output.n53 gnd 0.01428f
C97 output.n54 gnd 0.006397f
C98 output.n55 gnd 0.048111f
C99 output.t18 gnd 0.023274f
C100 output.n56 gnd 0.01071f
C101 output.n57 gnd 0.008435f
C102 output.n58 gnd 0.006041f
C103 output.n59 gnd 0.267512f
C104 output.n60 gnd 0.011243f
C105 output.n61 gnd 0.006041f
C106 output.n62 gnd 0.006397f
C107 output.n63 gnd 0.01428f
C108 output.n64 gnd 0.01428f
C109 output.n65 gnd 0.006397f
C110 output.n66 gnd 0.006041f
C111 output.n67 gnd 0.011243f
C112 output.n68 gnd 0.011243f
C113 output.n69 gnd 0.006041f
C114 output.n70 gnd 0.006397f
C115 output.n71 gnd 0.01428f
C116 output.n72 gnd 0.030913f
C117 output.n73 gnd 0.006397f
C118 output.n74 gnd 0.006041f
C119 output.n75 gnd 0.025987f
C120 output.n76 gnd 0.09306f
C121 output.n77 gnd 1.65264f
C122 output.n78 gnd 0.015803f
C123 output.n79 gnd 0.011243f
C124 output.n80 gnd 0.006041f
C125 output.n81 gnd 0.01428f
C126 output.n82 gnd 0.006397f
C127 output.n83 gnd 0.011243f
C128 output.n84 gnd 0.006041f
C129 output.n85 gnd 0.01428f
C130 output.n86 gnd 0.006397f
C131 output.n87 gnd 0.048111f
C132 output.t19 gnd 0.023274f
C133 output.n88 gnd 0.01071f
C134 output.n89 gnd 0.008435f
C135 output.n90 gnd 0.006041f
C136 output.n91 gnd 0.267512f
C137 output.n92 gnd 0.011243f
C138 output.n93 gnd 0.006041f
C139 output.n94 gnd 0.006397f
C140 output.n95 gnd 0.01428f
C141 output.n96 gnd 0.01428f
C142 output.n97 gnd 0.006397f
C143 output.n98 gnd 0.006041f
C144 output.n99 gnd 0.011243f
C145 output.n100 gnd 0.011243f
C146 output.n101 gnd 0.006041f
C147 output.n102 gnd 0.006397f
C148 output.n103 gnd 0.01428f
C149 output.n104 gnd 0.030913f
C150 output.n105 gnd 0.006397f
C151 output.n106 gnd 0.006041f
C152 output.n107 gnd 0.025987f
C153 output.n108 gnd 0.09306f
C154 output.n109 gnd 0.713089f
C155 output.n110 gnd 0.015803f
C156 output.n111 gnd 0.011243f
C157 output.n112 gnd 0.006041f
C158 output.n113 gnd 0.01428f
C159 output.n114 gnd 0.006397f
C160 output.n115 gnd 0.011243f
C161 output.n116 gnd 0.006041f
C162 output.n117 gnd 0.01428f
C163 output.n118 gnd 0.006397f
C164 output.n119 gnd 0.048111f
C165 output.t16 gnd 0.023274f
C166 output.n120 gnd 0.01071f
C167 output.n121 gnd 0.008435f
C168 output.n122 gnd 0.006041f
C169 output.n123 gnd 0.267512f
C170 output.n124 gnd 0.011243f
C171 output.n125 gnd 0.006041f
C172 output.n126 gnd 0.006397f
C173 output.n127 gnd 0.01428f
C174 output.n128 gnd 0.01428f
C175 output.n129 gnd 0.006397f
C176 output.n130 gnd 0.006041f
C177 output.n131 gnd 0.011243f
C178 output.n132 gnd 0.011243f
C179 output.n133 gnd 0.006041f
C180 output.n134 gnd 0.006397f
C181 output.n135 gnd 0.01428f
C182 output.n136 gnd 0.030913f
C183 output.n137 gnd 0.006397f
C184 output.n138 gnd 0.006041f
C185 output.n139 gnd 0.025987f
C186 output.n140 gnd 0.09306f
C187 output.n141 gnd 1.67353f
C188 outputibias.t9 gnd 0.11477f
C189 outputibias.t10 gnd 0.115567f
C190 outputibias.n0 gnd 0.130108f
C191 outputibias.n1 gnd 0.001372f
C192 outputibias.n2 gnd 9.76e-19
C193 outputibias.n3 gnd 5.24e-19
C194 outputibias.n4 gnd 0.001239f
C195 outputibias.n5 gnd 5.55e-19
C196 outputibias.n6 gnd 9.76e-19
C197 outputibias.n7 gnd 5.24e-19
C198 outputibias.n8 gnd 0.001239f
C199 outputibias.n9 gnd 5.55e-19
C200 outputibias.n10 gnd 0.004176f
C201 outputibias.t7 gnd 0.00202f
C202 outputibias.n11 gnd 9.3e-19
C203 outputibias.n12 gnd 7.32e-19
C204 outputibias.n13 gnd 5.24e-19
C205 outputibias.n14 gnd 0.02322f
C206 outputibias.n15 gnd 9.76e-19
C207 outputibias.n16 gnd 5.24e-19
C208 outputibias.n17 gnd 5.55e-19
C209 outputibias.n18 gnd 0.001239f
C210 outputibias.n19 gnd 0.001239f
C211 outputibias.n20 gnd 5.55e-19
C212 outputibias.n21 gnd 5.24e-19
C213 outputibias.n22 gnd 9.76e-19
C214 outputibias.n23 gnd 9.76e-19
C215 outputibias.n24 gnd 5.24e-19
C216 outputibias.n25 gnd 5.55e-19
C217 outputibias.n26 gnd 0.001239f
C218 outputibias.n27 gnd 0.002683f
C219 outputibias.n28 gnd 5.55e-19
C220 outputibias.n29 gnd 5.24e-19
C221 outputibias.n30 gnd 0.002256f
C222 outputibias.n31 gnd 0.005781f
C223 outputibias.n32 gnd 0.001372f
C224 outputibias.n33 gnd 9.76e-19
C225 outputibias.n34 gnd 5.24e-19
C226 outputibias.n35 gnd 0.001239f
C227 outputibias.n36 gnd 5.55e-19
C228 outputibias.n37 gnd 9.76e-19
C229 outputibias.n38 gnd 5.24e-19
C230 outputibias.n39 gnd 0.001239f
C231 outputibias.n40 gnd 5.55e-19
C232 outputibias.n41 gnd 0.004176f
C233 outputibias.t1 gnd 0.00202f
C234 outputibias.n42 gnd 9.3e-19
C235 outputibias.n43 gnd 7.32e-19
C236 outputibias.n44 gnd 5.24e-19
C237 outputibias.n45 gnd 0.02322f
C238 outputibias.n46 gnd 9.76e-19
C239 outputibias.n47 gnd 5.24e-19
C240 outputibias.n48 gnd 5.55e-19
C241 outputibias.n49 gnd 0.001239f
C242 outputibias.n50 gnd 0.001239f
C243 outputibias.n51 gnd 5.55e-19
C244 outputibias.n52 gnd 5.24e-19
C245 outputibias.n53 gnd 9.76e-19
C246 outputibias.n54 gnd 9.76e-19
C247 outputibias.n55 gnd 5.24e-19
C248 outputibias.n56 gnd 5.55e-19
C249 outputibias.n57 gnd 0.001239f
C250 outputibias.n58 gnd 0.002683f
C251 outputibias.n59 gnd 5.55e-19
C252 outputibias.n60 gnd 5.24e-19
C253 outputibias.n61 gnd 0.002256f
C254 outputibias.n62 gnd 0.005197f
C255 outputibias.n63 gnd 0.121892f
C256 outputibias.n64 gnd 0.001372f
C257 outputibias.n65 gnd 9.76e-19
C258 outputibias.n66 gnd 5.24e-19
C259 outputibias.n67 gnd 0.001239f
C260 outputibias.n68 gnd 5.55e-19
C261 outputibias.n69 gnd 9.76e-19
C262 outputibias.n70 gnd 5.24e-19
C263 outputibias.n71 gnd 0.001239f
C264 outputibias.n72 gnd 5.55e-19
C265 outputibias.n73 gnd 0.004176f
C266 outputibias.t3 gnd 0.00202f
C267 outputibias.n74 gnd 9.3e-19
C268 outputibias.n75 gnd 7.32e-19
C269 outputibias.n76 gnd 5.24e-19
C270 outputibias.n77 gnd 0.02322f
C271 outputibias.n78 gnd 9.76e-19
C272 outputibias.n79 gnd 5.24e-19
C273 outputibias.n80 gnd 5.55e-19
C274 outputibias.n81 gnd 0.001239f
C275 outputibias.n82 gnd 0.001239f
C276 outputibias.n83 gnd 5.55e-19
C277 outputibias.n84 gnd 5.24e-19
C278 outputibias.n85 gnd 9.76e-19
C279 outputibias.n86 gnd 9.76e-19
C280 outputibias.n87 gnd 5.24e-19
C281 outputibias.n88 gnd 5.55e-19
C282 outputibias.n89 gnd 0.001239f
C283 outputibias.n90 gnd 0.002683f
C284 outputibias.n91 gnd 5.55e-19
C285 outputibias.n92 gnd 5.24e-19
C286 outputibias.n93 gnd 0.002256f
C287 outputibias.n94 gnd 0.005197f
C288 outputibias.n95 gnd 0.064513f
C289 outputibias.n96 gnd 0.001372f
C290 outputibias.n97 gnd 9.76e-19
C291 outputibias.n98 gnd 5.24e-19
C292 outputibias.n99 gnd 0.001239f
C293 outputibias.n100 gnd 5.55e-19
C294 outputibias.n101 gnd 9.76e-19
C295 outputibias.n102 gnd 5.24e-19
C296 outputibias.n103 gnd 0.001239f
C297 outputibias.n104 gnd 5.55e-19
C298 outputibias.n105 gnd 0.004176f
C299 outputibias.t5 gnd 0.00202f
C300 outputibias.n106 gnd 9.3e-19
C301 outputibias.n107 gnd 7.32e-19
C302 outputibias.n108 gnd 5.24e-19
C303 outputibias.n109 gnd 0.02322f
C304 outputibias.n110 gnd 9.76e-19
C305 outputibias.n111 gnd 5.24e-19
C306 outputibias.n112 gnd 5.55e-19
C307 outputibias.n113 gnd 0.001239f
C308 outputibias.n114 gnd 0.001239f
C309 outputibias.n115 gnd 5.55e-19
C310 outputibias.n116 gnd 5.24e-19
C311 outputibias.n117 gnd 9.76e-19
C312 outputibias.n118 gnd 9.76e-19
C313 outputibias.n119 gnd 5.24e-19
C314 outputibias.n120 gnd 5.55e-19
C315 outputibias.n121 gnd 0.001239f
C316 outputibias.n122 gnd 0.002683f
C317 outputibias.n123 gnd 5.55e-19
C318 outputibias.n124 gnd 5.24e-19
C319 outputibias.n125 gnd 0.002256f
C320 outputibias.n126 gnd 0.005197f
C321 outputibias.n127 gnd 0.084814f
C322 outputibias.t4 gnd 0.108319f
C323 outputibias.t2 gnd 0.108319f
C324 outputibias.t0 gnd 0.108319f
C325 outputibias.t6 gnd 0.109238f
C326 outputibias.n128 gnd 0.134674f
C327 outputibias.n129 gnd 0.07244f
C328 outputibias.n130 gnd 0.079818f
C329 outputibias.n131 gnd 0.164901f
C330 outputibias.t11 gnd 0.11477f
C331 outputibias.n132 gnd 0.067481f
C332 outputibias.t8 gnd 0.11477f
C333 outputibias.n133 gnd 0.065115f
C334 outputibias.n134 gnd 0.029159f
C335 minus.n0 gnd 0.033094f
C336 minus.t27 gnd 0.33435f
C337 minus.n1 gnd 0.154274f
C338 minus.n2 gnd 0.033094f
C339 minus.t6 gnd 0.33435f
C340 minus.n3 gnd 0.151214f
C341 minus.n4 gnd 0.033094f
C342 minus.t24 gnd 0.33435f
C343 minus.n5 gnd 0.151214f
C344 minus.n6 gnd 0.033094f
C345 minus.t8 gnd 0.33435f
C346 minus.n7 gnd 0.154274f
C347 minus.t12 gnd 0.343352f
C348 minus.t18 gnd 0.33435f
C349 minus.n8 gnd 0.15819f
C350 minus.n9 gnd 0.143194f
C351 minus.n10 gnd 0.134377f
C352 minus.n11 gnd 0.033094f
C353 minus.n12 gnd 0.00751f
C354 minus.t13 gnd 0.33435f
C355 minus.n13 gnd 0.154581f
C356 minus.n14 gnd 0.00751f
C357 minus.n15 gnd 0.033094f
C358 minus.n16 gnd 0.033094f
C359 minus.n17 gnd 0.033094f
C360 minus.t19 gnd 0.33435f
C361 minus.n18 gnd 0.154479f
C362 minus.n19 gnd 0.00751f
C363 minus.t22 gnd 0.33435f
C364 minus.n20 gnd 0.154479f
C365 minus.n21 gnd 0.033094f
C366 minus.n22 gnd 0.033094f
C367 minus.n23 gnd 0.033094f
C368 minus.n24 gnd 0.00751f
C369 minus.t20 gnd 0.33435f
C370 minus.n25 gnd 0.154581f
C371 minus.n26 gnd 0.00751f
C372 minus.n27 gnd 0.033094f
C373 minus.n28 gnd 0.033094f
C374 minus.n29 gnd 0.033094f
C375 minus.t15 gnd 0.33435f
C376 minus.n30 gnd 0.151418f
C377 minus.n31 gnd 0.00751f
C378 minus.t9 gnd 0.33435f
C379 minus.n32 gnd 0.150806f
C380 minus.n33 gnd 0.371412f
C381 minus.n34 gnd 0.033094f
C382 minus.t16 gnd 0.33435f
C383 minus.t28 gnd 0.33435f
C384 minus.n35 gnd 0.033094f
C385 minus.t21 gnd 0.33435f
C386 minus.n36 gnd 0.033094f
C387 minus.t14 gnd 0.33435f
C388 minus.n37 gnd 0.154581f
C389 minus.n38 gnd 0.033094f
C390 minus.t23 gnd 0.33435f
C391 minus.t11 gnd 0.33435f
C392 minus.n39 gnd 0.033094f
C393 minus.t5 gnd 0.33435f
C394 minus.n40 gnd 0.154479f
C395 minus.n41 gnd 0.033094f
C396 minus.t17 gnd 0.33435f
C397 minus.t10 gnd 0.33435f
C398 minus.n42 gnd 0.033094f
C399 minus.t25 gnd 0.33435f
C400 minus.n43 gnd 0.154274f
C401 minus.t26 gnd 0.343352f
C402 minus.t7 gnd 0.33435f
C403 minus.n44 gnd 0.15819f
C404 minus.n45 gnd 0.143194f
C405 minus.n46 gnd 0.134377f
C406 minus.n47 gnd 0.033094f
C407 minus.n48 gnd 0.00751f
C408 minus.n49 gnd 0.154581f
C409 minus.n50 gnd 0.00751f
C410 minus.n51 gnd 0.151214f
C411 minus.n52 gnd 0.033094f
C412 minus.n53 gnd 0.033094f
C413 minus.n54 gnd 0.033094f
C414 minus.n55 gnd 0.00751f
C415 minus.n56 gnd 0.154479f
C416 minus.n57 gnd 0.151214f
C417 minus.n58 gnd 0.00751f
C418 minus.n59 gnd 0.033094f
C419 minus.n60 gnd 0.033094f
C420 minus.n61 gnd 0.033094f
C421 minus.n62 gnd 0.00751f
C422 minus.n63 gnd 0.154274f
C423 minus.n64 gnd 0.151418f
C424 minus.n65 gnd 0.00751f
C425 minus.n66 gnd 0.150806f
C426 minus.n67 gnd 1.00426f
C427 minus.n68 gnd 1.52338f
C428 minus.t1 gnd 0.010202f
C429 minus.t4 gnd 0.010202f
C430 minus.n69 gnd 0.033547f
C431 minus.t2 gnd 0.010202f
C432 minus.t0 gnd 0.010202f
C433 minus.n70 gnd 0.033087f
C434 minus.n71 gnd 0.282383f
C435 minus.t3 gnd 0.056783f
C436 minus.n72 gnd 0.154094f
C437 minus.n73 gnd 2.07222f
C438 plus.n0 gnd 0.023974f
C439 plus.t23 gnd 0.242206f
C440 plus.n1 gnd 0.023974f
C441 plus.t13 gnd 0.242206f
C442 plus.n2 gnd 0.023974f
C443 plus.t27 gnd 0.242206f
C444 plus.t22 gnd 0.242206f
C445 plus.n3 gnd 0.111979f
C446 plus.n4 gnd 0.023974f
C447 plus.t7 gnd 0.242206f
C448 plus.n5 gnd 0.023974f
C449 plus.t18 gnd 0.242206f
C450 plus.t14 gnd 0.242206f
C451 plus.n6 gnd 0.111906f
C452 plus.n7 gnd 0.023974f
C453 plus.t24 gnd 0.242206f
C454 plus.n8 gnd 0.023974f
C455 plus.t17 gnd 0.242206f
C456 plus.t9 gnd 0.242206f
C457 plus.n9 gnd 0.111758f
C458 plus.t12 gnd 0.248727f
C459 plus.t15 gnd 0.242206f
C460 plus.n10 gnd 0.114594f
C461 plus.n11 gnd 0.103731f
C462 plus.n12 gnd 0.097344f
C463 plus.n13 gnd 0.023974f
C464 plus.n14 gnd 0.00544f
C465 plus.n15 gnd 0.111979f
C466 plus.n16 gnd 0.00544f
C467 plus.n17 gnd 0.109541f
C468 plus.n18 gnd 0.023974f
C469 plus.n19 gnd 0.023974f
C470 plus.n20 gnd 0.023974f
C471 plus.n21 gnd 0.00544f
C472 plus.n22 gnd 0.111906f
C473 plus.n23 gnd 0.109541f
C474 plus.n24 gnd 0.00544f
C475 plus.n25 gnd 0.023974f
C476 plus.n26 gnd 0.023974f
C477 plus.n27 gnd 0.023974f
C478 plus.n28 gnd 0.00544f
C479 plus.n29 gnd 0.111758f
C480 plus.n30 gnd 0.109688f
C481 plus.n31 gnd 0.00544f
C482 plus.n32 gnd 0.109245f
C483 plus.n33 gnd 0.262859f
C484 plus.n34 gnd 0.023974f
C485 plus.t16 gnd 0.242206f
C486 plus.n35 gnd 0.111758f
C487 plus.t28 gnd 0.242206f
C488 plus.n36 gnd 0.023974f
C489 plus.t19 gnd 0.242206f
C490 plus.n37 gnd 0.109541f
C491 plus.n38 gnd 0.023974f
C492 plus.t11 gnd 0.242206f
C493 plus.n39 gnd 0.109541f
C494 plus.t6 gnd 0.242206f
C495 plus.n40 gnd 0.023974f
C496 plus.t20 gnd 0.242206f
C497 plus.n41 gnd 0.111758f
C498 plus.t25 gnd 0.248727f
C499 plus.t5 gnd 0.242206f
C500 plus.n42 gnd 0.114594f
C501 plus.n43 gnd 0.103731f
C502 plus.n44 gnd 0.097344f
C503 plus.n45 gnd 0.023974f
C504 plus.n46 gnd 0.00544f
C505 plus.t26 gnd 0.242206f
C506 plus.n47 gnd 0.111979f
C507 plus.n48 gnd 0.00544f
C508 plus.n49 gnd 0.023974f
C509 plus.n50 gnd 0.023974f
C510 plus.n51 gnd 0.023974f
C511 plus.n52 gnd 0.111906f
C512 plus.n53 gnd 0.00544f
C513 plus.t10 gnd 0.242206f
C514 plus.n54 gnd 0.111906f
C515 plus.n55 gnd 0.023974f
C516 plus.n56 gnd 0.023974f
C517 plus.n57 gnd 0.023974f
C518 plus.n58 gnd 0.00544f
C519 plus.t8 gnd 0.242206f
C520 plus.n59 gnd 0.111979f
C521 plus.n60 gnd 0.00544f
C522 plus.n61 gnd 0.023974f
C523 plus.n62 gnd 0.023974f
C524 plus.n63 gnd 0.023974f
C525 plus.n64 gnd 0.109688f
C526 plus.n65 gnd 0.00544f
C527 plus.t21 gnd 0.242206f
C528 plus.n66 gnd 0.109245f
C529 plus.n67 gnd 0.717857f
C530 plus.n68 gnd 1.0941f
C531 plus.t3 gnd 0.041386f
C532 plus.t4 gnd 0.00739f
C533 plus.t1 gnd 0.00739f
C534 plus.n69 gnd 0.023968f
C535 plus.n70 gnd 0.18607f
C536 plus.t0 gnd 0.00739f
C537 plus.t2 gnd 0.00739f
C538 plus.n71 gnd 0.023968f
C539 plus.n72 gnd 0.139668f
C540 plus.n73 gnd 2.65334f
C541 a_n2982_8322.t26 gnd 0.100219f
C542 a_n2982_8322.t2 gnd 20.791302f
C543 a_n2982_8322.t3 gnd 20.6455f
C544 a_n2982_8322.t5 gnd 20.6455f
C545 a_n2982_8322.t1 gnd 20.791302f
C546 a_n2982_8322.t4 gnd 20.6455f
C547 a_n2982_8322.t0 gnd 28.6983f
C548 a_n2982_8322.t35 gnd 0.938395f
C549 a_n2982_8322.t28 gnd 0.100219f
C550 a_n2982_8322.t24 gnd 0.100219f
C551 a_n2982_8322.n0 gnd 0.705941f
C552 a_n2982_8322.n1 gnd 0.788787f
C553 a_n2982_8322.t21 gnd 0.100219f
C554 a_n2982_8322.t37 gnd 0.100219f
C555 a_n2982_8322.n2 gnd 0.705941f
C556 a_n2982_8322.n3 gnd 0.400772f
C557 a_n2982_8322.t34 gnd 0.100219f
C558 a_n2982_8322.t22 gnd 0.100219f
C559 a_n2982_8322.n4 gnd 0.705941f
C560 a_n2982_8322.n5 gnd 0.400772f
C561 a_n2982_8322.t19 gnd 0.100219f
C562 a_n2982_8322.t18 gnd 0.100219f
C563 a_n2982_8322.n6 gnd 0.705941f
C564 a_n2982_8322.n7 gnd 0.400772f
C565 a_n2982_8322.t32 gnd 0.100219f
C566 a_n2982_8322.t31 gnd 0.100219f
C567 a_n2982_8322.n8 gnd 0.705941f
C568 a_n2982_8322.n9 gnd 0.400772f
C569 a_n2982_8322.t15 gnd 0.936529f
C570 a_n2982_8322.n10 gnd 1.11212f
C571 a_n2982_8322.n11 gnd 3.23133f
C572 a_n2982_8322.t9 gnd 0.938398f
C573 a_n2982_8322.t13 gnd 0.100219f
C574 a_n2982_8322.t12 gnd 0.100219f
C575 a_n2982_8322.n12 gnd 0.705941f
C576 a_n2982_8322.n13 gnd 0.788785f
C577 a_n2982_8322.t7 gnd 0.936529f
C578 a_n2982_8322.n14 gnd 0.396928f
C579 a_n2982_8322.t10 gnd 0.936529f
C580 a_n2982_8322.n15 gnd 0.396928f
C581 a_n2982_8322.t8 gnd 0.100219f
C582 a_n2982_8322.t6 gnd 0.100219f
C583 a_n2982_8322.n16 gnd 0.705941f
C584 a_n2982_8322.n17 gnd 0.400772f
C585 a_n2982_8322.t11 gnd 0.936529f
C586 a_n2982_8322.n18 gnd 1.47227f
C587 a_n2982_8322.n19 gnd 2.35273f
C588 a_n2982_8322.t14 gnd 0.936529f
C589 a_n2982_8322.n20 gnd 1.8725f
C590 a_n2982_8322.t27 gnd 0.100219f
C591 a_n2982_8322.t25 gnd 0.100219f
C592 a_n2982_8322.n21 gnd 0.705941f
C593 a_n2982_8322.n22 gnd 0.400772f
C594 a_n2982_8322.t30 gnd 0.100219f
C595 a_n2982_8322.t23 gnd 0.100219f
C596 a_n2982_8322.n23 gnd 0.705941f
C597 a_n2982_8322.n24 gnd 0.400772f
C598 a_n2982_8322.t17 gnd 0.100219f
C599 a_n2982_8322.t16 gnd 0.100219f
C600 a_n2982_8322.n25 gnd 0.705941f
C601 a_n2982_8322.n26 gnd 0.400772f
C602 a_n2982_8322.t20 gnd 0.938398f
C603 a_n2982_8322.t33 gnd 0.100219f
C604 a_n2982_8322.t29 gnd 0.100219f
C605 a_n2982_8322.n27 gnd 0.705941f
C606 a_n2982_8322.n28 gnd 0.788785f
C607 a_n2982_8322.n29 gnd 0.40077f
C608 a_n2982_8322.n30 gnd 0.705943f
C609 a_n2982_8322.t36 gnd 0.100219f
C610 a_n3827_n3924.n0 gnd 1.10033f
C611 a_n3827_n3924.n1 gnd 0.958536f
C612 a_n3827_n3924.t26 gnd 1.06719f
C613 a_n3827_n3924.n2 gnd 0.920943f
C614 a_n3827_n3924.t55 gnd 0.102682f
C615 a_n3827_n3924.t1 gnd 0.102682f
C616 a_n3827_n3924.n3 gnd 0.838616f
C617 a_n3827_n3924.n4 gnd 0.340114f
C618 a_n3827_n3924.t40 gnd 0.102682f
C619 a_n3827_n3924.t37 gnd 0.102682f
C620 a_n3827_n3924.n5 gnd 0.838616f
C621 a_n3827_n3924.n6 gnd 0.340114f
C622 a_n3827_n3924.t15 gnd 0.102682f
C623 a_n3827_n3924.t9 gnd 0.102682f
C624 a_n3827_n3924.n7 gnd 0.838616f
C625 a_n3827_n3924.n8 gnd 0.340114f
C626 a_n3827_n3924.t57 gnd 0.102682f
C627 a_n3827_n3924.t16 gnd 0.102682f
C628 a_n3827_n3924.n9 gnd 0.838616f
C629 a_n3827_n3924.n10 gnd 0.340114f
C630 a_n3827_n3924.t28 gnd 0.102682f
C631 a_n3827_n3924.t38 gnd 0.102682f
C632 a_n3827_n3924.n11 gnd 0.838616f
C633 a_n3827_n3924.n12 gnd 0.340114f
C634 a_n3827_n3924.t20 gnd 1.06719f
C635 a_n3827_n3924.n13 gnd 0.362194f
C636 a_n3827_n3924.t27 gnd 1.06719f
C637 a_n3827_n3924.n14 gnd 0.362194f
C638 a_n3827_n3924.t3 gnd 0.102682f
C639 a_n3827_n3924.t10 gnd 0.102682f
C640 a_n3827_n3924.n15 gnd 0.838616f
C641 a_n3827_n3924.n16 gnd 0.340114f
C642 a_n3827_n3924.t39 gnd 0.102682f
C643 a_n3827_n3924.t32 gnd 0.102682f
C644 a_n3827_n3924.n17 gnd 0.838616f
C645 a_n3827_n3924.n18 gnd 0.340114f
C646 a_n3827_n3924.t22 gnd 0.102682f
C647 a_n3827_n3924.t17 gnd 0.102682f
C648 a_n3827_n3924.n19 gnd 0.838616f
C649 a_n3827_n3924.n20 gnd 0.340114f
C650 a_n3827_n3924.t52 gnd 0.102682f
C651 a_n3827_n3924.t0 gnd 0.102682f
C652 a_n3827_n3924.n21 gnd 0.838616f
C653 a_n3827_n3924.n22 gnd 0.340114f
C654 a_n3827_n3924.t56 gnd 0.102682f
C655 a_n3827_n3924.t30 gnd 0.102682f
C656 a_n3827_n3924.n23 gnd 0.838616f
C657 a_n3827_n3924.n24 gnd 0.340114f
C658 a_n3827_n3924.t2 gnd 1.06718f
C659 a_n3827_n3924.n25 gnd 0.920947f
C660 a_n3827_n3924.t14 gnd 1.06718f
C661 a_n3827_n3924.n26 gnd 0.58539f
C662 a_n3827_n3924.t11 gnd 0.102682f
C663 a_n3827_n3924.t51 gnd 0.102682f
C664 a_n3827_n3924.n27 gnd 0.838615f
C665 a_n3827_n3924.n28 gnd 0.340116f
C666 a_n3827_n3924.t4 gnd 0.102682f
C667 a_n3827_n3924.t5 gnd 0.102682f
C668 a_n3827_n3924.n29 gnd 0.838615f
C669 a_n3827_n3924.n30 gnd 0.340116f
C670 a_n3827_n3924.t24 gnd 0.102682f
C671 a_n3827_n3924.t53 gnd 0.102682f
C672 a_n3827_n3924.n31 gnd 0.838615f
C673 a_n3827_n3924.n32 gnd 0.340116f
C674 a_n3827_n3924.t29 gnd 0.102682f
C675 a_n3827_n3924.t23 gnd 0.102682f
C676 a_n3827_n3924.n33 gnd 0.838615f
C677 a_n3827_n3924.n34 gnd 0.340116f
C678 a_n3827_n3924.t33 gnd 0.102682f
C679 a_n3827_n3924.t54 gnd 0.102682f
C680 a_n3827_n3924.n35 gnd 0.838615f
C681 a_n3827_n3924.n36 gnd 0.340116f
C682 a_n3827_n3924.t19 gnd 1.06718f
C683 a_n3827_n3924.n37 gnd 0.362198f
C684 a_n3827_n3924.t35 gnd 1.06718f
C685 a_n3827_n3924.n38 gnd 0.362198f
C686 a_n3827_n3924.t18 gnd 0.102682f
C687 a_n3827_n3924.t8 gnd 0.102682f
C688 a_n3827_n3924.n39 gnd 0.838615f
C689 a_n3827_n3924.n40 gnd 0.340116f
C690 a_n3827_n3924.t21 gnd 0.102682f
C691 a_n3827_n3924.t34 gnd 0.102682f
C692 a_n3827_n3924.n41 gnd 0.838615f
C693 a_n3827_n3924.n42 gnd 0.340116f
C694 a_n3827_n3924.t31 gnd 0.102682f
C695 a_n3827_n3924.t13 gnd 0.102682f
C696 a_n3827_n3924.n43 gnd 0.838615f
C697 a_n3827_n3924.n44 gnd 0.340116f
C698 a_n3827_n3924.t12 gnd 0.102682f
C699 a_n3827_n3924.t7 gnd 0.102682f
C700 a_n3827_n3924.n45 gnd 0.838615f
C701 a_n3827_n3924.n46 gnd 0.340116f
C702 a_n3827_n3924.t25 gnd 0.102682f
C703 a_n3827_n3924.t6 gnd 0.102682f
C704 a_n3827_n3924.n47 gnd 0.838615f
C705 a_n3827_n3924.n48 gnd 0.340116f
C706 a_n3827_n3924.t36 gnd 1.06718f
C707 a_n3827_n3924.n49 gnd 0.58539f
C708 a_n3827_n3924.n50 gnd 0.958536f
C709 a_n3827_n3924.t43 gnd 1.32959f
C710 a_n3827_n3924.t47 gnd 1.32595f
C711 a_n3827_n3924.n51 gnd 1.82937f
C712 a_n3827_n3924.n52 gnd 0.504753f
C713 a_n3827_n3924.t42 gnd 1.32595f
C714 a_n3827_n3924.n53 gnd 0.844057f
C715 a_n3827_n3924.t45 gnd 1.32595f
C716 a_n3827_n3924.n54 gnd 0.933892f
C717 a_n3827_n3924.t41 gnd 1.32595f
C718 a_n3827_n3924.n55 gnd 0.933892f
C719 a_n3827_n3924.t46 gnd 1.32595f
C720 a_n3827_n3924.n56 gnd 0.933892f
C721 a_n3827_n3924.t49 gnd 1.32595f
C722 a_n3827_n3924.n57 gnd 0.918983f
C723 a_n3827_n3924.t48 gnd 1.32595f
C724 a_n3827_n3924.t44 gnd 1.32595f
C725 a_n3827_n3924.n58 gnd 1.5379f
C726 a_n3827_n3924.t50 gnd 1.32785f
C727 diffpairibias.t27 gnd 0.090128f
C728 diffpairibias.t23 gnd 0.08996f
C729 diffpairibias.n0 gnd 0.105991f
C730 diffpairibias.t28 gnd 0.08996f
C731 diffpairibias.n1 gnd 0.051736f
C732 diffpairibias.t25 gnd 0.08996f
C733 diffpairibias.n2 gnd 0.051736f
C734 diffpairibias.t29 gnd 0.08996f
C735 diffpairibias.n3 gnd 0.041084f
C736 diffpairibias.t15 gnd 0.086371f
C737 diffpairibias.t1 gnd 0.085993f
C738 diffpairibias.n4 gnd 0.13579f
C739 diffpairibias.t11 gnd 0.085993f
C740 diffpairibias.n5 gnd 0.072463f
C741 diffpairibias.t13 gnd 0.085993f
C742 diffpairibias.n6 gnd 0.072463f
C743 diffpairibias.t7 gnd 0.085993f
C744 diffpairibias.n7 gnd 0.072463f
C745 diffpairibias.t3 gnd 0.085993f
C746 diffpairibias.n8 gnd 0.072463f
C747 diffpairibias.t17 gnd 0.085993f
C748 diffpairibias.n9 gnd 0.072463f
C749 diffpairibias.t5 gnd 0.085993f
C750 diffpairibias.n10 gnd 0.072463f
C751 diffpairibias.t19 gnd 0.085993f
C752 diffpairibias.n11 gnd 0.072463f
C753 diffpairibias.t9 gnd 0.085993f
C754 diffpairibias.n12 gnd 0.102883f
C755 diffpairibias.t14 gnd 0.086899f
C756 diffpairibias.t0 gnd 0.086748f
C757 diffpairibias.n13 gnd 0.094648f
C758 diffpairibias.t10 gnd 0.086748f
C759 diffpairibias.n14 gnd 0.052262f
C760 diffpairibias.t12 gnd 0.086748f
C761 diffpairibias.n15 gnd 0.052262f
C762 diffpairibias.t6 gnd 0.086748f
C763 diffpairibias.n16 gnd 0.052262f
C764 diffpairibias.t2 gnd 0.086748f
C765 diffpairibias.n17 gnd 0.052262f
C766 diffpairibias.t16 gnd 0.086748f
C767 diffpairibias.n18 gnd 0.052262f
C768 diffpairibias.t4 gnd 0.086748f
C769 diffpairibias.n19 gnd 0.052262f
C770 diffpairibias.t18 gnd 0.086748f
C771 diffpairibias.n20 gnd 0.052262f
C772 diffpairibias.t8 gnd 0.086748f
C773 diffpairibias.n21 gnd 0.061849f
C774 diffpairibias.n22 gnd 0.233513f
C775 diffpairibias.t20 gnd 0.08996f
C776 diffpairibias.n23 gnd 0.051747f
C777 diffpairibias.t26 gnd 0.08996f
C778 diffpairibias.n24 gnd 0.051736f
C779 diffpairibias.t22 gnd 0.08996f
C780 diffpairibias.n25 gnd 0.051736f
C781 diffpairibias.t21 gnd 0.08996f
C782 diffpairibias.n26 gnd 0.051736f
C783 diffpairibias.t24 gnd 0.08996f
C784 diffpairibias.n27 gnd 0.04729f
C785 diffpairibias.n28 gnd 0.047711f
C786 CSoutput.n0 gnd 0.041367f
C787 CSoutput.t145 gnd 0.273631f
C788 CSoutput.n1 gnd 0.123558f
C789 CSoutput.n2 gnd 0.041367f
C790 CSoutput.t149 gnd 0.273631f
C791 CSoutput.n3 gnd 0.032786f
C792 CSoutput.n4 gnd 0.041367f
C793 CSoutput.t158 gnd 0.273631f
C794 CSoutput.n5 gnd 0.028272f
C795 CSoutput.n6 gnd 0.041367f
C796 CSoutput.t147 gnd 0.273631f
C797 CSoutput.t151 gnd 0.273631f
C798 CSoutput.n7 gnd 0.122211f
C799 CSoutput.n8 gnd 0.041367f
C800 CSoutput.t157 gnd 0.273631f
C801 CSoutput.n9 gnd 0.026956f
C802 CSoutput.n10 gnd 0.041367f
C803 CSoutput.t161 gnd 0.273631f
C804 CSoutput.t148 gnd 0.273631f
C805 CSoutput.n11 gnd 0.122211f
C806 CSoutput.n12 gnd 0.041367f
C807 CSoutput.t156 gnd 0.273631f
C808 CSoutput.n13 gnd 0.028272f
C809 CSoutput.n14 gnd 0.041367f
C810 CSoutput.t153 gnd 0.273631f
C811 CSoutput.t165 gnd 0.273631f
C812 CSoutput.n15 gnd 0.122211f
C813 CSoutput.n16 gnd 0.041367f
C814 CSoutput.t152 gnd 0.273631f
C815 CSoutput.n17 gnd 0.030196f
C816 CSoutput.t160 gnd 0.326996f
C817 CSoutput.t150 gnd 0.273631f
C818 CSoutput.n18 gnd 0.156016f
C819 CSoutput.n19 gnd 0.15139f
C820 CSoutput.n20 gnd 0.17563f
C821 CSoutput.n21 gnd 0.041367f
C822 CSoutput.n22 gnd 0.034525f
C823 CSoutput.n23 gnd 0.122211f
C824 CSoutput.n24 gnd 0.033281f
C825 CSoutput.n25 gnd 0.032786f
C826 CSoutput.n26 gnd 0.041367f
C827 CSoutput.n27 gnd 0.041367f
C828 CSoutput.n28 gnd 0.034259f
C829 CSoutput.n29 gnd 0.029087f
C830 CSoutput.n30 gnd 0.124932f
C831 CSoutput.n31 gnd 0.029488f
C832 CSoutput.n32 gnd 0.041367f
C833 CSoutput.n33 gnd 0.041367f
C834 CSoutput.n34 gnd 0.041367f
C835 CSoutput.n35 gnd 0.033895f
C836 CSoutput.n36 gnd 0.122211f
C837 CSoutput.n37 gnd 0.032415f
C838 CSoutput.n38 gnd 0.033652f
C839 CSoutput.n39 gnd 0.041367f
C840 CSoutput.n40 gnd 0.041367f
C841 CSoutput.n41 gnd 0.034518f
C842 CSoutput.n42 gnd 0.031549f
C843 CSoutput.n43 gnd 0.122211f
C844 CSoutput.n44 gnd 0.032349f
C845 CSoutput.n45 gnd 0.041367f
C846 CSoutput.n46 gnd 0.041367f
C847 CSoutput.n47 gnd 0.041367f
C848 CSoutput.n48 gnd 0.032349f
C849 CSoutput.n49 gnd 0.122211f
C850 CSoutput.n50 gnd 0.031549f
C851 CSoutput.n51 gnd 0.034518f
C852 CSoutput.n52 gnd 0.041367f
C853 CSoutput.n53 gnd 0.041367f
C854 CSoutput.n54 gnd 0.033652f
C855 CSoutput.n55 gnd 0.032415f
C856 CSoutput.n56 gnd 0.122211f
C857 CSoutput.n57 gnd 0.033895f
C858 CSoutput.n58 gnd 0.041367f
C859 CSoutput.n59 gnd 0.041367f
C860 CSoutput.n60 gnd 0.041367f
C861 CSoutput.n61 gnd 0.029488f
C862 CSoutput.n62 gnd 0.124932f
C863 CSoutput.n63 gnd 0.029087f
C864 CSoutput.t159 gnd 0.273631f
C865 CSoutput.n64 gnd 0.122211f
C866 CSoutput.n65 gnd 0.034259f
C867 CSoutput.n66 gnd 0.041367f
C868 CSoutput.n67 gnd 0.041367f
C869 CSoutput.n68 gnd 0.041367f
C870 CSoutput.n69 gnd 0.033281f
C871 CSoutput.n70 gnd 0.122211f
C872 CSoutput.n71 gnd 0.034525f
C873 CSoutput.n72 gnd 0.030196f
C874 CSoutput.n73 gnd 0.041367f
C875 CSoutput.n74 gnd 0.041367f
C876 CSoutput.n75 gnd 0.031315f
C877 CSoutput.n76 gnd 0.018598f
C878 CSoutput.t164 gnd 0.307444f
C879 CSoutput.n77 gnd 0.152726f
C880 CSoutput.n78 gnd 0.624793f
C881 CSoutput.t71 gnd 0.051599f
C882 CSoutput.t35 gnd 0.051599f
C883 CSoutput.n79 gnd 0.399496f
C884 CSoutput.t10 gnd 0.051599f
C885 CSoutput.t61 gnd 0.051599f
C886 CSoutput.n80 gnd 0.398784f
C887 CSoutput.n81 gnd 0.404765f
C888 CSoutput.t17 gnd 0.051599f
C889 CSoutput.t47 gnd 0.051599f
C890 CSoutput.n82 gnd 0.398784f
C891 CSoutput.n83 gnd 0.199451f
C892 CSoutput.t29 gnd 0.051599f
C893 CSoutput.t41 gnd 0.051599f
C894 CSoutput.n84 gnd 0.398784f
C895 CSoutput.n85 gnd 0.199451f
C896 CSoutput.t38 gnd 0.051599f
C897 CSoutput.t65 gnd 0.051599f
C898 CSoutput.n86 gnd 0.398784f
C899 CSoutput.n87 gnd 0.199451f
C900 CSoutput.t21 gnd 0.051599f
C901 CSoutput.t52 gnd 0.051599f
C902 CSoutput.n88 gnd 0.398784f
C903 CSoutput.n89 gnd 0.365747f
C904 CSoutput.t39 gnd 0.051599f
C905 CSoutput.t18 gnd 0.051599f
C906 CSoutput.n90 gnd 0.399496f
C907 CSoutput.t4 gnd 0.051599f
C908 CSoutput.t40 gnd 0.051599f
C909 CSoutput.n91 gnd 0.398784f
C910 CSoutput.n92 gnd 0.404765f
C911 CSoutput.t36 gnd 0.051599f
C912 CSoutput.t16 gnd 0.051599f
C913 CSoutput.n93 gnd 0.398784f
C914 CSoutput.n94 gnd 0.199451f
C915 CSoutput.t3 gnd 0.051599f
C916 CSoutput.t1 gnd 0.051599f
C917 CSoutput.n95 gnd 0.398784f
C918 CSoutput.n96 gnd 0.199451f
C919 CSoutput.t48 gnd 0.051599f
C920 CSoutput.t26 gnd 0.051599f
C921 CSoutput.n97 gnd 0.398784f
C922 CSoutput.n98 gnd 0.199451f
C923 CSoutput.t23 gnd 0.051599f
C924 CSoutput.t0 gnd 0.051599f
C925 CSoutput.n99 gnd 0.398784f
C926 CSoutput.n100 gnd 0.297432f
C927 CSoutput.n101 gnd 0.37506f
C928 CSoutput.t44 gnd 0.051599f
C929 CSoutput.t27 gnd 0.051599f
C930 CSoutput.n102 gnd 0.399496f
C931 CSoutput.t13 gnd 0.051599f
C932 CSoutput.t45 gnd 0.051599f
C933 CSoutput.n103 gnd 0.398784f
C934 CSoutput.n104 gnd 0.404765f
C935 CSoutput.t43 gnd 0.051599f
C936 CSoutput.t25 gnd 0.051599f
C937 CSoutput.n105 gnd 0.398784f
C938 CSoutput.n106 gnd 0.199451f
C939 CSoutput.t12 gnd 0.051599f
C940 CSoutput.t11 gnd 0.051599f
C941 CSoutput.n107 gnd 0.398784f
C942 CSoutput.n108 gnd 0.199451f
C943 CSoutput.t54 gnd 0.051599f
C944 CSoutput.t32 gnd 0.051599f
C945 CSoutput.n109 gnd 0.398784f
C946 CSoutput.n110 gnd 0.199451f
C947 CSoutput.t30 gnd 0.051599f
C948 CSoutput.t8 gnd 0.051599f
C949 CSoutput.n111 gnd 0.398784f
C950 CSoutput.n112 gnd 0.297432f
C951 CSoutput.n113 gnd 0.419221f
C952 CSoutput.n114 gnd 7.73775f
C953 CSoutput.n116 gnd 0.731767f
C954 CSoutput.n117 gnd 0.548825f
C955 CSoutput.n118 gnd 0.731767f
C956 CSoutput.n119 gnd 0.731767f
C957 CSoutput.n120 gnd 1.97014f
C958 CSoutput.n121 gnd 0.731767f
C959 CSoutput.n122 gnd 0.731767f
C960 CSoutput.t154 gnd 0.914709f
C961 CSoutput.n123 gnd 0.731767f
C962 CSoutput.n124 gnd 0.731767f
C963 CSoutput.n128 gnd 0.731767f
C964 CSoutput.n132 gnd 0.731767f
C965 CSoutput.n133 gnd 0.731767f
C966 CSoutput.n135 gnd 0.731767f
C967 CSoutput.n140 gnd 0.731767f
C968 CSoutput.n142 gnd 0.731767f
C969 CSoutput.n143 gnd 0.731767f
C970 CSoutput.n145 gnd 0.731767f
C971 CSoutput.n146 gnd 0.731767f
C972 CSoutput.n148 gnd 0.731767f
C973 CSoutput.t144 gnd 12.2277f
C974 CSoutput.n150 gnd 0.731767f
C975 CSoutput.n151 gnd 0.548825f
C976 CSoutput.n152 gnd 0.731767f
C977 CSoutput.n153 gnd 0.731767f
C978 CSoutput.n154 gnd 1.97014f
C979 CSoutput.n155 gnd 0.731767f
C980 CSoutput.n156 gnd 0.731767f
C981 CSoutput.t162 gnd 0.914709f
C982 CSoutput.n157 gnd 0.731767f
C983 CSoutput.n158 gnd 0.731767f
C984 CSoutput.n162 gnd 0.731767f
C985 CSoutput.n166 gnd 0.731767f
C986 CSoutput.n167 gnd 0.731767f
C987 CSoutput.n169 gnd 0.731767f
C988 CSoutput.n174 gnd 0.731767f
C989 CSoutput.n176 gnd 0.731767f
C990 CSoutput.n177 gnd 0.731767f
C991 CSoutput.n179 gnd 0.731767f
C992 CSoutput.n180 gnd 0.731767f
C993 CSoutput.n182 gnd 0.731767f
C994 CSoutput.n183 gnd 0.548825f
C995 CSoutput.n185 gnd 0.731767f
C996 CSoutput.n186 gnd 0.548825f
C997 CSoutput.n187 gnd 0.731767f
C998 CSoutput.n188 gnd 0.731767f
C999 CSoutput.n189 gnd 1.97014f
C1000 CSoutput.n190 gnd 0.731767f
C1001 CSoutput.n191 gnd 0.731767f
C1002 CSoutput.t155 gnd 0.914709f
C1003 CSoutput.n192 gnd 0.731767f
C1004 CSoutput.n193 gnd 1.97014f
C1005 CSoutput.n195 gnd 0.731767f
C1006 CSoutput.n196 gnd 0.731767f
C1007 CSoutput.n198 gnd 0.731767f
C1008 CSoutput.n199 gnd 0.731767f
C1009 CSoutput.t163 gnd 12.0285f
C1010 CSoutput.t146 gnd 12.2277f
C1011 CSoutput.n205 gnd 2.29566f
C1012 CSoutput.n206 gnd 9.35169f
C1013 CSoutput.n207 gnd 9.743f
C1014 CSoutput.n212 gnd 2.48682f
C1015 CSoutput.n218 gnd 0.731767f
C1016 CSoutput.n220 gnd 0.731767f
C1017 CSoutput.n222 gnd 0.731767f
C1018 CSoutput.n224 gnd 0.731767f
C1019 CSoutput.n226 gnd 0.731767f
C1020 CSoutput.n232 gnd 0.731767f
C1021 CSoutput.n239 gnd 1.34251f
C1022 CSoutput.n240 gnd 1.34251f
C1023 CSoutput.n241 gnd 0.731767f
C1024 CSoutput.n242 gnd 0.731767f
C1025 CSoutput.n244 gnd 0.548825f
C1026 CSoutput.n245 gnd 0.47002f
C1027 CSoutput.n247 gnd 0.548825f
C1028 CSoutput.n248 gnd 0.47002f
C1029 CSoutput.n249 gnd 0.548825f
C1030 CSoutput.n251 gnd 0.731767f
C1031 CSoutput.n253 gnd 1.97014f
C1032 CSoutput.n254 gnd 2.29566f
C1033 CSoutput.n255 gnd 8.601151f
C1034 CSoutput.n257 gnd 0.548825f
C1035 CSoutput.n258 gnd 1.41216f
C1036 CSoutput.n259 gnd 0.548825f
C1037 CSoutput.n261 gnd 0.731767f
C1038 CSoutput.n263 gnd 1.97014f
C1039 CSoutput.n264 gnd 4.29129f
C1040 CSoutput.t34 gnd 0.051599f
C1041 CSoutput.t20 gnd 0.051599f
C1042 CSoutput.n265 gnd 0.399496f
C1043 CSoutput.t60 gnd 0.051599f
C1044 CSoutput.t9 gnd 0.051599f
C1045 CSoutput.n266 gnd 0.398784f
C1046 CSoutput.n267 gnd 0.404765f
C1047 CSoutput.t46 gnd 0.051599f
C1048 CSoutput.t15 gnd 0.051599f
C1049 CSoutput.n268 gnd 0.398784f
C1050 CSoutput.n269 gnd 0.199451f
C1051 CSoutput.t56 gnd 0.051599f
C1052 CSoutput.t28 gnd 0.051599f
C1053 CSoutput.n270 gnd 0.398784f
C1054 CSoutput.n271 gnd 0.199451f
C1055 CSoutput.t64 gnd 0.051599f
C1056 CSoutput.t37 gnd 0.051599f
C1057 CSoutput.n272 gnd 0.398784f
C1058 CSoutput.n273 gnd 0.199451f
C1059 CSoutput.t51 gnd 0.051599f
C1060 CSoutput.t22 gnd 0.051599f
C1061 CSoutput.n274 gnd 0.398784f
C1062 CSoutput.n275 gnd 0.365747f
C1063 CSoutput.t62 gnd 0.051599f
C1064 CSoutput.t63 gnd 0.051599f
C1065 CSoutput.n276 gnd 0.399496f
C1066 CSoutput.t7 gnd 0.051599f
C1067 CSoutput.t53 gnd 0.051599f
C1068 CSoutput.n277 gnd 0.398784f
C1069 CSoutput.n278 gnd 0.404765f
C1070 CSoutput.t59 gnd 0.051599f
C1071 CSoutput.t5 gnd 0.051599f
C1072 CSoutput.n279 gnd 0.398784f
C1073 CSoutput.n280 gnd 0.199451f
C1074 CSoutput.t33 gnd 0.051599f
C1075 CSoutput.t50 gnd 0.051599f
C1076 CSoutput.n281 gnd 0.398784f
C1077 CSoutput.n282 gnd 0.199451f
C1078 CSoutput.t67 gnd 0.051599f
C1079 CSoutput.t24 gnd 0.051599f
C1080 CSoutput.n283 gnd 0.398784f
C1081 CSoutput.n284 gnd 0.199451f
C1082 CSoutput.t49 gnd 0.051599f
C1083 CSoutput.t70 gnd 0.051599f
C1084 CSoutput.n285 gnd 0.398784f
C1085 CSoutput.n286 gnd 0.297432f
C1086 CSoutput.n287 gnd 0.37506f
C1087 CSoutput.t68 gnd 0.051599f
C1088 CSoutput.t69 gnd 0.051599f
C1089 CSoutput.n288 gnd 0.399496f
C1090 CSoutput.t19 gnd 0.051599f
C1091 CSoutput.t58 gnd 0.051599f
C1092 CSoutput.n289 gnd 0.398784f
C1093 CSoutput.n290 gnd 0.404765f
C1094 CSoutput.t66 gnd 0.051599f
C1095 CSoutput.t14 gnd 0.051599f
C1096 CSoutput.n291 gnd 0.398784f
C1097 CSoutput.n292 gnd 0.199451f
C1098 CSoutput.t42 gnd 0.051599f
C1099 CSoutput.t57 gnd 0.051599f
C1100 CSoutput.n293 gnd 0.398784f
C1101 CSoutput.n294 gnd 0.199451f
C1102 CSoutput.t2 gnd 0.051599f
C1103 CSoutput.t31 gnd 0.051599f
C1104 CSoutput.n295 gnd 0.398784f
C1105 CSoutput.n296 gnd 0.199451f
C1106 CSoutput.t55 gnd 0.051599f
C1107 CSoutput.t6 gnd 0.051599f
C1108 CSoutput.n297 gnd 0.398783f
C1109 CSoutput.n298 gnd 0.297433f
C1110 CSoutput.n299 gnd 0.419221f
C1111 CSoutput.n300 gnd 11.0842f
C1112 CSoutput.t134 gnd 0.045149f
C1113 CSoutput.t81 gnd 0.045149f
C1114 CSoutput.n301 gnd 0.400288f
C1115 CSoutput.t121 gnd 0.045149f
C1116 CSoutput.t74 gnd 0.045149f
C1117 CSoutput.n302 gnd 0.398953f
C1118 CSoutput.n303 gnd 0.37175f
C1119 CSoutput.t106 gnd 0.045149f
C1120 CSoutput.t137 gnd 0.045149f
C1121 CSoutput.n304 gnd 0.398953f
C1122 CSoutput.n305 gnd 0.183255f
C1123 CSoutput.t94 gnd 0.045149f
C1124 CSoutput.t105 gnd 0.045149f
C1125 CSoutput.n306 gnd 0.398953f
C1126 CSoutput.n307 gnd 0.183255f
C1127 CSoutput.t76 gnd 0.045149f
C1128 CSoutput.t111 gnd 0.045149f
C1129 CSoutput.n308 gnd 0.398953f
C1130 CSoutput.n309 gnd 0.183255f
C1131 CSoutput.t125 gnd 0.045149f
C1132 CSoutput.t95 gnd 0.045149f
C1133 CSoutput.n310 gnd 0.398953f
C1134 CSoutput.n311 gnd 0.338004f
C1135 CSoutput.t103 gnd 0.045149f
C1136 CSoutput.t86 gnd 0.045149f
C1137 CSoutput.n312 gnd 0.400288f
C1138 CSoutput.t90 gnd 0.045149f
C1139 CSoutput.t102 gnd 0.045149f
C1140 CSoutput.n313 gnd 0.398953f
C1141 CSoutput.n314 gnd 0.37175f
C1142 CSoutput.t85 gnd 0.045149f
C1143 CSoutput.t92 gnd 0.045149f
C1144 CSoutput.n315 gnd 0.398953f
C1145 CSoutput.n316 gnd 0.183255f
C1146 CSoutput.t104 gnd 0.045149f
C1147 CSoutput.t84 gnd 0.045149f
C1148 CSoutput.n317 gnd 0.398953f
C1149 CSoutput.n318 gnd 0.183255f
C1150 CSoutput.t91 gnd 0.045149f
C1151 CSoutput.t79 gnd 0.045149f
C1152 CSoutput.n319 gnd 0.398953f
C1153 CSoutput.n320 gnd 0.183255f
C1154 CSoutput.t83 gnd 0.045149f
C1155 CSoutput.t93 gnd 0.045149f
C1156 CSoutput.n321 gnd 0.398953f
C1157 CSoutput.n322 gnd 0.278221f
C1158 CSoutput.n323 gnd 0.350923f
C1159 CSoutput.t80 gnd 0.045149f
C1160 CSoutput.t141 gnd 0.045149f
C1161 CSoutput.n324 gnd 0.400288f
C1162 CSoutput.t132 gnd 0.045149f
C1163 CSoutput.t87 gnd 0.045149f
C1164 CSoutput.n325 gnd 0.398953f
C1165 CSoutput.n326 gnd 0.37175f
C1166 CSoutput.t72 gnd 0.045149f
C1167 CSoutput.t138 gnd 0.045149f
C1168 CSoutput.n327 gnd 0.398953f
C1169 CSoutput.n328 gnd 0.183255f
C1170 CSoutput.t98 gnd 0.045149f
C1171 CSoutput.t107 gnd 0.045149f
C1172 CSoutput.n329 gnd 0.398953f
C1173 CSoutput.n330 gnd 0.183255f
C1174 CSoutput.t142 gnd 0.045149f
C1175 CSoutput.t131 gnd 0.045149f
C1176 CSoutput.n331 gnd 0.398953f
C1177 CSoutput.n332 gnd 0.183255f
C1178 CSoutput.t116 gnd 0.045149f
C1179 CSoutput.t73 gnd 0.045149f
C1180 CSoutput.n333 gnd 0.398953f
C1181 CSoutput.n334 gnd 0.278221f
C1182 CSoutput.n335 gnd 0.376836f
C1183 CSoutput.n336 gnd 11.2107f
C1184 CSoutput.t113 gnd 0.045149f
C1185 CSoutput.t77 gnd 0.045149f
C1186 CSoutput.n337 gnd 0.400288f
C1187 CSoutput.t97 gnd 0.045149f
C1188 CSoutput.t139 gnd 0.045149f
C1189 CSoutput.n338 gnd 0.398953f
C1190 CSoutput.n339 gnd 0.37175f
C1191 CSoutput.t78 gnd 0.045149f
C1192 CSoutput.t127 gnd 0.045149f
C1193 CSoutput.n340 gnd 0.398953f
C1194 CSoutput.n341 gnd 0.183255f
C1195 CSoutput.t126 gnd 0.045149f
C1196 CSoutput.t115 gnd 0.045149f
C1197 CSoutput.n342 gnd 0.398953f
C1198 CSoutput.n343 gnd 0.183255f
C1199 CSoutput.t128 gnd 0.045149f
C1200 CSoutput.t99 gnd 0.045149f
C1201 CSoutput.n344 gnd 0.398953f
C1202 CSoutput.n345 gnd 0.183255f
C1203 CSoutput.t122 gnd 0.045149f
C1204 CSoutput.t133 gnd 0.045149f
C1205 CSoutput.n346 gnd 0.398953f
C1206 CSoutput.n347 gnd 0.338004f
C1207 CSoutput.t100 gnd 0.045149f
C1208 CSoutput.t117 gnd 0.045149f
C1209 CSoutput.n348 gnd 0.400288f
C1210 CSoutput.t118 gnd 0.045149f
C1211 CSoutput.t109 gnd 0.045149f
C1212 CSoutput.n349 gnd 0.398953f
C1213 CSoutput.n350 gnd 0.37175f
C1214 CSoutput.t108 gnd 0.045149f
C1215 CSoutput.t101 gnd 0.045149f
C1216 CSoutput.n351 gnd 0.398953f
C1217 CSoutput.n352 gnd 0.183255f
C1218 CSoutput.t96 gnd 0.045149f
C1219 CSoutput.t88 gnd 0.045149f
C1220 CSoutput.n353 gnd 0.398953f
C1221 CSoutput.n354 gnd 0.183255f
C1222 CSoutput.t89 gnd 0.045149f
C1223 CSoutput.t110 gnd 0.045149f
C1224 CSoutput.n355 gnd 0.398953f
C1225 CSoutput.n356 gnd 0.183255f
C1226 CSoutput.t112 gnd 0.045149f
C1227 CSoutput.t75 gnd 0.045149f
C1228 CSoutput.n357 gnd 0.398953f
C1229 CSoutput.n358 gnd 0.278221f
C1230 CSoutput.n359 gnd 0.350923f
C1231 CSoutput.t129 gnd 0.045149f
C1232 CSoutput.t140 gnd 0.045149f
C1233 CSoutput.n360 gnd 0.400288f
C1234 CSoutput.t143 gnd 0.045149f
C1235 CSoutput.t120 gnd 0.045149f
C1236 CSoutput.n361 gnd 0.398953f
C1237 CSoutput.n362 gnd 0.37175f
C1238 CSoutput.t124 gnd 0.045149f
C1239 CSoutput.t135 gnd 0.045149f
C1240 CSoutput.n363 gnd 0.398953f
C1241 CSoutput.n364 gnd 0.183255f
C1242 CSoutput.t82 gnd 0.045149f
C1243 CSoutput.t114 gnd 0.045149f
C1244 CSoutput.n365 gnd 0.398953f
C1245 CSoutput.n366 gnd 0.183255f
C1246 CSoutput.t119 gnd 0.045149f
C1247 CSoutput.t130 gnd 0.045149f
C1248 CSoutput.n367 gnd 0.398953f
C1249 CSoutput.n368 gnd 0.183255f
C1250 CSoutput.t136 gnd 0.045149f
C1251 CSoutput.t123 gnd 0.045149f
C1252 CSoutput.n369 gnd 0.398953f
C1253 CSoutput.n370 gnd 0.278221f
C1254 CSoutput.n371 gnd 0.376836f
C1255 CSoutput.n372 gnd 6.49258f
C1256 CSoutput.n373 gnd 12.4894f
C1257 a_n8300_8799.n0 gnd 0.183261f
C1258 a_n8300_8799.n1 gnd 0.21461f
C1259 a_n8300_8799.n2 gnd 0.21461f
C1260 a_n8300_8799.n3 gnd 0.21461f
C1261 a_n8300_8799.n4 gnd 0.183261f
C1262 a_n8300_8799.n5 gnd 0.21461f
C1263 a_n8300_8799.n6 gnd 0.21461f
C1264 a_n8300_8799.n7 gnd 0.21461f
C1265 a_n8300_8799.n8 gnd 0.353995f
C1266 a_n8300_8799.n9 gnd 0.21461f
C1267 a_n8300_8799.n10 gnd 0.21461f
C1268 a_n8300_8799.n11 gnd 0.21461f
C1269 a_n8300_8799.n12 gnd 0.21461f
C1270 a_n8300_8799.n13 gnd 0.21461f
C1271 a_n8300_8799.n14 gnd 0.183261f
C1272 a_n8300_8799.n15 gnd 0.21461f
C1273 a_n8300_8799.n16 gnd 0.21461f
C1274 a_n8300_8799.n17 gnd 0.21461f
C1275 a_n8300_8799.n18 gnd 0.183261f
C1276 a_n8300_8799.n19 gnd 0.21461f
C1277 a_n8300_8799.n20 gnd 0.21461f
C1278 a_n8300_8799.n21 gnd 0.21461f
C1279 a_n8300_8799.n22 gnd 0.353995f
C1280 a_n8300_8799.n23 gnd 0.21461f
C1281 a_n8300_8799.n24 gnd 3.52204f
C1282 a_n8300_8799.n25 gnd 1.79585f
C1283 a_n8300_8799.n26 gnd 3.05554f
C1284 a_n8300_8799.n27 gnd 1.05358f
C1285 a_n8300_8799.n28 gnd 1.03866f
C1286 a_n8300_8799.n29 gnd 3.11527f
C1287 a_n8300_8799.n30 gnd 3.79872f
C1288 a_n8300_8799.n31 gnd 1.03866f
C1289 a_n8300_8799.n32 gnd 1.57291f
C1290 a_n8300_8799.n33 gnd 0.722524f
C1291 a_n8300_8799.n34 gnd 0.259534f
C1292 a_n8300_8799.n36 gnd 0.007994f
C1293 a_n8300_8799.n37 gnd 0.012082f
C1294 a_n8300_8799.n38 gnd 0.008309f
C1295 a_n8300_8799.n40 gnd 4.15e-19
C1296 a_n8300_8799.n41 gnd 0.008611f
C1297 a_n8300_8799.n42 gnd 0.271503f
C1298 a_n8300_8799.n43 gnd 0.259534f
C1299 a_n8300_8799.n45 gnd 0.007994f
C1300 a_n8300_8799.n46 gnd 0.012082f
C1301 a_n8300_8799.n47 gnd 0.008309f
C1302 a_n8300_8799.n49 gnd 4.15e-19
C1303 a_n8300_8799.n50 gnd 0.008611f
C1304 a_n8300_8799.n51 gnd 0.271503f
C1305 a_n8300_8799.n52 gnd 0.259534f
C1306 a_n8300_8799.n54 gnd 0.007994f
C1307 a_n8300_8799.n55 gnd 0.012082f
C1308 a_n8300_8799.n56 gnd 0.008309f
C1309 a_n8300_8799.n58 gnd 4.15e-19
C1310 a_n8300_8799.n59 gnd 0.008611f
C1311 a_n8300_8799.n60 gnd 0.271503f
C1312 a_n8300_8799.n61 gnd 0.008611f
C1313 a_n8300_8799.n62 gnd 0.271503f
C1314 a_n8300_8799.n63 gnd 4.15e-19
C1315 a_n8300_8799.n65 gnd 0.008309f
C1316 a_n8300_8799.n66 gnd 0.012082f
C1317 a_n8300_8799.n67 gnd 0.007994f
C1318 a_n8300_8799.n69 gnd 0.259534f
C1319 a_n8300_8799.n70 gnd 0.008611f
C1320 a_n8300_8799.n71 gnd 0.271503f
C1321 a_n8300_8799.n72 gnd 4.15e-19
C1322 a_n8300_8799.n74 gnd 0.008309f
C1323 a_n8300_8799.n75 gnd 0.012082f
C1324 a_n8300_8799.n76 gnd 0.007994f
C1325 a_n8300_8799.n78 gnd 0.259534f
C1326 a_n8300_8799.n79 gnd 0.008611f
C1327 a_n8300_8799.n80 gnd 0.271503f
C1328 a_n8300_8799.n81 gnd 4.15e-19
C1329 a_n8300_8799.n83 gnd 0.008309f
C1330 a_n8300_8799.n84 gnd 0.012082f
C1331 a_n8300_8799.n85 gnd 0.007994f
C1332 a_n8300_8799.n87 gnd 0.259534f
C1333 a_n8300_8799.t21 gnd 0.148856f
C1334 a_n8300_8799.t20 gnd 0.148856f
C1335 a_n8300_8799.t28 gnd 0.148856f
C1336 a_n8300_8799.n88 gnd 1.17405f
C1337 a_n8300_8799.t24 gnd 0.148856f
C1338 a_n8300_8799.t41 gnd 0.148856f
C1339 a_n8300_8799.n89 gnd 1.17211f
C1340 a_n8300_8799.t32 gnd 0.148856f
C1341 a_n8300_8799.t27 gnd 0.148856f
C1342 a_n8300_8799.n90 gnd 1.17211f
C1343 a_n8300_8799.t33 gnd 0.148856f
C1344 a_n8300_8799.t29 gnd 0.148856f
C1345 a_n8300_8799.n91 gnd 1.17211f
C1346 a_n8300_8799.t38 gnd 0.148856f
C1347 a_n8300_8799.t25 gnd 0.148856f
C1348 a_n8300_8799.n92 gnd 1.17211f
C1349 a_n8300_8799.t37 gnd 0.148856f
C1350 a_n8300_8799.t39 gnd 0.148856f
C1351 a_n8300_8799.n93 gnd 1.17211f
C1352 a_n8300_8799.t13 gnd 0.115777f
C1353 a_n8300_8799.t2 gnd 0.115777f
C1354 a_n8300_8799.n94 gnd 1.02467f
C1355 a_n8300_8799.t5 gnd 0.115777f
C1356 a_n8300_8799.t18 gnd 0.115777f
C1357 a_n8300_8799.n95 gnd 1.02304f
C1358 a_n8300_8799.t16 gnd 0.115777f
C1359 a_n8300_8799.t10 gnd 0.115777f
C1360 a_n8300_8799.n96 gnd 1.02304f
C1361 a_n8300_8799.t7 gnd 0.115777f
C1362 a_n8300_8799.t6 gnd 0.115777f
C1363 a_n8300_8799.n97 gnd 1.02467f
C1364 a_n8300_8799.t43 gnd 0.115777f
C1365 a_n8300_8799.t3 gnd 0.115777f
C1366 a_n8300_8799.n98 gnd 1.02304f
C1367 a_n8300_8799.t4 gnd 0.115777f
C1368 a_n8300_8799.t12 gnd 0.115777f
C1369 a_n8300_8799.n99 gnd 1.02304f
C1370 a_n8300_8799.t46 gnd 0.115777f
C1371 a_n8300_8799.t9 gnd 0.115777f
C1372 a_n8300_8799.n100 gnd 1.02467f
C1373 a_n8300_8799.t11 gnd 0.115777f
C1374 a_n8300_8799.t17 gnd 0.115777f
C1375 a_n8300_8799.n101 gnd 1.02304f
C1376 a_n8300_8799.t45 gnd 0.115777f
C1377 a_n8300_8799.t14 gnd 0.115777f
C1378 a_n8300_8799.n102 gnd 1.02304f
C1379 a_n8300_8799.t15 gnd 0.115777f
C1380 a_n8300_8799.t1 gnd 0.115777f
C1381 a_n8300_8799.n103 gnd 1.02304f
C1382 a_n8300_8799.t0 gnd 0.115777f
C1383 a_n8300_8799.t47 gnd 0.115777f
C1384 a_n8300_8799.n104 gnd 1.02304f
C1385 a_n8300_8799.t8 gnd 0.115777f
C1386 a_n8300_8799.t44 gnd 0.115777f
C1387 a_n8300_8799.n105 gnd 1.02304f
C1388 a_n8300_8799.t74 gnd 0.617225f
C1389 a_n8300_8799.n106 gnd 0.27935f
C1390 a_n8300_8799.t75 gnd 0.617225f
C1391 a_n8300_8799.t94 gnd 0.617225f
C1392 a_n8300_8799.n107 gnd 0.270206f
C1393 a_n8300_8799.t107 gnd 0.617225f
C1394 a_n8300_8799.n108 gnd 0.281966f
C1395 a_n8300_8799.t108 gnd 0.617225f
C1396 a_n8300_8799.t65 gnd 0.617225f
C1397 a_n8300_8799.n109 gnd 0.275168f
C1398 a_n8300_8799.t89 gnd 0.631731f
C1399 a_n8300_8799.t111 gnd 0.617225f
C1400 a_n8300_8799.n110 gnd 0.281517f
C1401 a_n8300_8799.n111 gnd 0.257292f
C1402 a_n8300_8799.t87 gnd 0.617225f
C1403 a_n8300_8799.n112 gnd 0.279228f
C1404 a_n8300_8799.n113 gnd 0.279365f
C1405 a_n8300_8799.t76 gnd 0.617225f
C1406 a_n8300_8799.n114 gnd 0.275499f
C1407 a_n8300_8799.t106 gnd 0.617225f
C1408 a_n8300_8799.n115 gnd 0.275757f
C1409 a_n8300_8799.n116 gnd 0.281517f
C1410 a_n8300_8799.t92 gnd 0.62843f
C1411 a_n8300_8799.t79 gnd 0.617225f
C1412 a_n8300_8799.n117 gnd 0.27935f
C1413 a_n8300_8799.t80 gnd 0.617225f
C1414 a_n8300_8799.t103 gnd 0.617225f
C1415 a_n8300_8799.n118 gnd 0.270206f
C1416 a_n8300_8799.t116 gnd 0.617225f
C1417 a_n8300_8799.n119 gnd 0.281966f
C1418 a_n8300_8799.t118 gnd 0.617225f
C1419 a_n8300_8799.t71 gnd 0.617225f
C1420 a_n8300_8799.n120 gnd 0.275168f
C1421 a_n8300_8799.t96 gnd 0.631731f
C1422 a_n8300_8799.t119 gnd 0.617225f
C1423 a_n8300_8799.n121 gnd 0.281517f
C1424 a_n8300_8799.n122 gnd 0.257292f
C1425 a_n8300_8799.t93 gnd 0.617225f
C1426 a_n8300_8799.n123 gnd 0.279228f
C1427 a_n8300_8799.n124 gnd 0.279365f
C1428 a_n8300_8799.t83 gnd 0.617225f
C1429 a_n8300_8799.n125 gnd 0.275499f
C1430 a_n8300_8799.t115 gnd 0.617225f
C1431 a_n8300_8799.n126 gnd 0.275757f
C1432 a_n8300_8799.n127 gnd 0.281517f
C1433 a_n8300_8799.t101 gnd 0.62843f
C1434 a_n8300_8799.n128 gnd 0.926624f
C1435 a_n8300_8799.t58 gnd 0.617225f
C1436 a_n8300_8799.n129 gnd 0.27935f
C1437 a_n8300_8799.t48 gnd 0.617225f
C1438 a_n8300_8799.t72 gnd 0.617225f
C1439 a_n8300_8799.n130 gnd 0.270206f
C1440 a_n8300_8799.t90 gnd 0.617225f
C1441 a_n8300_8799.n131 gnd 0.281966f
C1442 a_n8300_8799.t78 gnd 0.617225f
C1443 a_n8300_8799.t81 gnd 0.617225f
C1444 a_n8300_8799.n132 gnd 0.275168f
C1445 a_n8300_8799.t98 gnd 0.631731f
C1446 a_n8300_8799.t67 gnd 0.617225f
C1447 a_n8300_8799.n133 gnd 0.281517f
C1448 a_n8300_8799.n134 gnd 0.257292f
C1449 a_n8300_8799.t54 gnd 0.617225f
C1450 a_n8300_8799.n135 gnd 0.279228f
C1451 a_n8300_8799.n136 gnd 0.279365f
C1452 a_n8300_8799.t102 gnd 0.617225f
C1453 a_n8300_8799.n137 gnd 0.275499f
C1454 a_n8300_8799.t109 gnd 0.617225f
C1455 a_n8300_8799.n138 gnd 0.275757f
C1456 a_n8300_8799.n139 gnd 0.281517f
C1457 a_n8300_8799.t84 gnd 0.62843f
C1458 a_n8300_8799.n140 gnd 1.90527f
C1459 a_n8300_8799.t51 gnd 0.62843f
C1460 a_n8300_8799.t50 gnd 0.617225f
C1461 a_n8300_8799.t100 gnd 0.617225f
C1462 a_n8300_8799.t61 gnd 0.617225f
C1463 a_n8300_8799.n141 gnd 0.275757f
C1464 a_n8300_8799.t53 gnd 0.617225f
C1465 a_n8300_8799.t105 gnd 0.617225f
C1466 a_n8300_8799.t77 gnd 0.617225f
C1467 a_n8300_8799.n142 gnd 0.279365f
C1468 a_n8300_8799.t62 gnd 0.617225f
C1469 a_n8300_8799.t117 gnd 0.617225f
C1470 a_n8300_8799.t88 gnd 0.617225f
C1471 a_n8300_8799.n143 gnd 0.275168f
C1472 a_n8300_8799.t113 gnd 0.631731f
C1473 a_n8300_8799.t64 gnd 0.617225f
C1474 a_n8300_8799.n144 gnd 0.281517f
C1475 a_n8300_8799.n145 gnd 0.257292f
C1476 a_n8300_8799.n146 gnd 0.279228f
C1477 a_n8300_8799.n147 gnd 0.281966f
C1478 a_n8300_8799.n148 gnd 0.275499f
C1479 a_n8300_8799.n149 gnd 0.270206f
C1480 a_n8300_8799.n150 gnd 0.27935f
C1481 a_n8300_8799.n151 gnd 0.281517f
C1482 a_n8300_8799.t57 gnd 0.62843f
C1483 a_n8300_8799.t56 gnd 0.617225f
C1484 a_n8300_8799.t112 gnd 0.617225f
C1485 a_n8300_8799.t66 gnd 0.617225f
C1486 a_n8300_8799.n152 gnd 0.275757f
C1487 a_n8300_8799.t60 gnd 0.617225f
C1488 a_n8300_8799.t114 gnd 0.617225f
C1489 a_n8300_8799.t86 gnd 0.617225f
C1490 a_n8300_8799.n153 gnd 0.279365f
C1491 a_n8300_8799.t69 gnd 0.617225f
C1492 a_n8300_8799.t52 gnd 0.617225f
C1493 a_n8300_8799.t95 gnd 0.617225f
C1494 a_n8300_8799.n154 gnd 0.275168f
C1495 a_n8300_8799.t49 gnd 0.631731f
C1496 a_n8300_8799.t70 gnd 0.617225f
C1497 a_n8300_8799.n155 gnd 0.281517f
C1498 a_n8300_8799.n156 gnd 0.257292f
C1499 a_n8300_8799.n157 gnd 0.279228f
C1500 a_n8300_8799.n158 gnd 0.281966f
C1501 a_n8300_8799.n159 gnd 0.275499f
C1502 a_n8300_8799.n160 gnd 0.270206f
C1503 a_n8300_8799.n161 gnd 0.27935f
C1504 a_n8300_8799.n162 gnd 0.281517f
C1505 a_n8300_8799.n163 gnd 0.926624f
C1506 a_n8300_8799.t85 gnd 0.62843f
C1507 a_n8300_8799.t99 gnd 0.617225f
C1508 a_n8300_8799.t59 gnd 0.617225f
C1509 a_n8300_8799.t110 gnd 0.617225f
C1510 a_n8300_8799.n164 gnd 0.275757f
C1511 a_n8300_8799.t73 gnd 0.617225f
C1512 a_n8300_8799.t104 gnd 0.617225f
C1513 a_n8300_8799.t63 gnd 0.617225f
C1514 a_n8300_8799.n165 gnd 0.279365f
C1515 a_n8300_8799.t91 gnd 0.617225f
C1516 a_n8300_8799.t55 gnd 0.617225f
C1517 a_n8300_8799.t82 gnd 0.617225f
C1518 a_n8300_8799.n166 gnd 0.275168f
C1519 a_n8300_8799.t97 gnd 0.631731f
C1520 a_n8300_8799.t68 gnd 0.617225f
C1521 a_n8300_8799.n167 gnd 0.281517f
C1522 a_n8300_8799.n168 gnd 0.257292f
C1523 a_n8300_8799.n169 gnd 0.279228f
C1524 a_n8300_8799.n170 gnd 0.281966f
C1525 a_n8300_8799.n171 gnd 0.275499f
C1526 a_n8300_8799.n172 gnd 0.270206f
C1527 a_n8300_8799.n173 gnd 0.27935f
C1528 a_n8300_8799.n174 gnd 0.281517f
C1529 a_n8300_8799.n175 gnd 1.4618f
C1530 a_n8300_8799.n176 gnd 17.9394f
C1531 a_n8300_8799.n177 gnd 4.51719f
C1532 a_n8300_8799.n178 gnd 7.87732f
C1533 a_n8300_8799.t42 gnd 0.148856f
C1534 a_n8300_8799.t22 gnd 0.148856f
C1535 a_n8300_8799.n179 gnd 1.17211f
C1536 a_n8300_8799.t34 gnd 0.148856f
C1537 a_n8300_8799.t30 gnd 0.148856f
C1538 a_n8300_8799.n180 gnd 1.17211f
C1539 a_n8300_8799.t23 gnd 0.148856f
C1540 a_n8300_8799.t35 gnd 0.148856f
C1541 a_n8300_8799.n181 gnd 1.17211f
C1542 a_n8300_8799.t31 gnd 0.148856f
C1543 a_n8300_8799.t36 gnd 0.148856f
C1544 a_n8300_8799.n182 gnd 1.17211f
C1545 a_n8300_8799.t26 gnd 0.148856f
C1546 a_n8300_8799.t40 gnd 0.148856f
C1547 a_n8300_8799.n183 gnd 1.17211f
C1548 a_n8300_8799.n184 gnd 1.17405f
C1549 a_n8300_8799.t19 gnd 0.148856f
C1550 a_n2804_13878.t29 gnd 0.194878f
C1551 a_n2804_13878.t25 gnd 0.194878f
C1552 a_n2804_13878.t31 gnd 0.194878f
C1553 a_n2804_13878.n0 gnd 1.53703f
C1554 a_n2804_13878.t8 gnd 0.194878f
C1555 a_n2804_13878.t20 gnd 0.194878f
C1556 a_n2804_13878.n1 gnd 1.5345f
C1557 a_n2804_13878.n2 gnd 1.37932f
C1558 a_n2804_13878.t12 gnd 0.194878f
C1559 a_n2804_13878.t22 gnd 0.194878f
C1560 a_n2804_13878.n3 gnd 1.53612f
C1561 a_n2804_13878.t27 gnd 0.194878f
C1562 a_n2804_13878.t17 gnd 0.194878f
C1563 a_n2804_13878.n4 gnd 1.5345f
C1564 a_n2804_13878.n5 gnd 2.14416f
C1565 a_n2804_13878.t23 gnd 0.194878f
C1566 a_n2804_13878.t16 gnd 0.194878f
C1567 a_n2804_13878.n6 gnd 1.5345f
C1568 a_n2804_13878.n7 gnd 1.04587f
C1569 a_n2804_13878.t10 gnd 0.194878f
C1570 a_n2804_13878.t13 gnd 0.194878f
C1571 a_n2804_13878.n8 gnd 1.5345f
C1572 a_n2804_13878.n9 gnd 1.04587f
C1573 a_n2804_13878.t26 gnd 0.194878f
C1574 a_n2804_13878.t11 gnd 0.194878f
C1575 a_n2804_13878.n10 gnd 1.5345f
C1576 a_n2804_13878.n11 gnd 1.04587f
C1577 a_n2804_13878.t21 gnd 0.194878f
C1578 a_n2804_13878.t9 gnd 0.194878f
C1579 a_n2804_13878.n12 gnd 1.5345f
C1580 a_n2804_13878.n13 gnd 4.90989f
C1581 a_n2804_13878.t1 gnd 1.82474f
C1582 a_n2804_13878.t4 gnd 0.194878f
C1583 a_n2804_13878.t5 gnd 0.194878f
C1584 a_n2804_13878.n14 gnd 1.37272f
C1585 a_n2804_13878.n15 gnd 1.53381f
C1586 a_n2804_13878.t0 gnd 1.8211f
C1587 a_n2804_13878.n16 gnd 0.771835f
C1588 a_n2804_13878.t3 gnd 1.8211f
C1589 a_n2804_13878.n17 gnd 0.771835f
C1590 a_n2804_13878.t6 gnd 0.194878f
C1591 a_n2804_13878.t7 gnd 0.194878f
C1592 a_n2804_13878.n18 gnd 1.37272f
C1593 a_n2804_13878.n19 gnd 0.77931f
C1594 a_n2804_13878.t2 gnd 1.8211f
C1595 a_n2804_13878.n20 gnd 2.86287f
C1596 a_n2804_13878.n21 gnd 3.75497f
C1597 a_n2804_13878.t15 gnd 0.194878f
C1598 a_n2804_13878.t24 gnd 0.194878f
C1599 a_n2804_13878.n22 gnd 1.53449f
C1600 a_n2804_13878.n23 gnd 2.50654f
C1601 a_n2804_13878.t28 gnd 0.194878f
C1602 a_n2804_13878.t14 gnd 0.194878f
C1603 a_n2804_13878.n24 gnd 1.5345f
C1604 a_n2804_13878.n25 gnd 0.679894f
C1605 a_n2804_13878.t18 gnd 0.194878f
C1606 a_n2804_13878.t19 gnd 0.194878f
C1607 a_n2804_13878.n26 gnd 1.5345f
C1608 a_n2804_13878.n27 gnd 0.679894f
C1609 a_n2804_13878.n28 gnd 0.679892f
C1610 a_n2804_13878.n29 gnd 1.5345f
C1611 a_n2804_13878.t30 gnd 0.194878f
C1612 vdd.t216 gnd 0.032423f
C1613 vdd.t197 gnd 0.032423f
C1614 vdd.n0 gnd 0.255722f
C1615 vdd.t175 gnd 0.032423f
C1616 vdd.t212 gnd 0.032423f
C1617 vdd.n1 gnd 0.2553f
C1618 vdd.n2 gnd 0.235436f
C1619 vdd.t193 gnd 0.032423f
C1620 vdd.t223 gnd 0.032423f
C1621 vdd.n3 gnd 0.2553f
C1622 vdd.n4 gnd 0.119069f
C1623 vdd.t221 gnd 0.032423f
C1624 vdd.t201 gnd 0.032423f
C1625 vdd.n5 gnd 0.2553f
C1626 vdd.n6 gnd 0.111724f
C1627 vdd.t227 gnd 0.032423f
C1628 vdd.t191 gnd 0.032423f
C1629 vdd.n7 gnd 0.255722f
C1630 vdd.t199 gnd 0.032423f
C1631 vdd.t219 gnd 0.032423f
C1632 vdd.n8 gnd 0.2553f
C1633 vdd.n9 gnd 0.235436f
C1634 vdd.t208 gnd 0.032423f
C1635 vdd.t179 gnd 0.032423f
C1636 vdd.n10 gnd 0.2553f
C1637 vdd.n11 gnd 0.119069f
C1638 vdd.t188 gnd 0.032423f
C1639 vdd.t206 gnd 0.032423f
C1640 vdd.n12 gnd 0.2553f
C1641 vdd.n13 gnd 0.111724f
C1642 vdd.n14 gnd 0.078987f
C1643 vdd.t163 gnd 0.018013f
C1644 vdd.t104 gnd 0.018013f
C1645 vdd.n15 gnd 0.165798f
C1646 vdd.t126 gnd 0.018013f
C1647 vdd.t109 gnd 0.018013f
C1648 vdd.n16 gnd 0.165313f
C1649 vdd.n17 gnd 0.287696f
C1650 vdd.t106 gnd 0.018013f
C1651 vdd.t125 gnd 0.018013f
C1652 vdd.n18 gnd 0.165313f
C1653 vdd.n19 gnd 0.119024f
C1654 vdd.t127 gnd 0.018013f
C1655 vdd.t110 gnd 0.018013f
C1656 vdd.n20 gnd 0.165798f
C1657 vdd.t170 gnd 0.018013f
C1658 vdd.t105 gnd 0.018013f
C1659 vdd.n21 gnd 0.165313f
C1660 vdd.n22 gnd 0.287696f
C1661 vdd.t171 gnd 0.018013f
C1662 vdd.t8 gnd 0.018013f
C1663 vdd.n23 gnd 0.165313f
C1664 vdd.n24 gnd 0.119024f
C1665 vdd.t107 gnd 0.018013f
C1666 vdd.t142 gnd 0.018013f
C1667 vdd.n25 gnd 0.165313f
C1668 vdd.t9 gnd 0.018013f
C1669 vdd.t111 gnd 0.018013f
C1670 vdd.n26 gnd 0.165313f
C1671 vdd.n27 gnd 18.0989f
C1672 vdd.n28 gnd 7.13208f
C1673 vdd.n29 gnd 0.004913f
C1674 vdd.n30 gnd 0.004559f
C1675 vdd.n31 gnd 0.002522f
C1676 vdd.n32 gnd 0.00579f
C1677 vdd.n33 gnd 0.00245f
C1678 vdd.n34 gnd 0.002594f
C1679 vdd.n35 gnd 0.004559f
C1680 vdd.n36 gnd 0.00245f
C1681 vdd.n37 gnd 0.00579f
C1682 vdd.n38 gnd 0.002594f
C1683 vdd.n39 gnd 0.004559f
C1684 vdd.n40 gnd 0.00245f
C1685 vdd.n41 gnd 0.004343f
C1686 vdd.n42 gnd 0.004356f
C1687 vdd.t5 gnd 0.01244f
C1688 vdd.n43 gnd 0.027678f
C1689 vdd.n44 gnd 0.144045f
C1690 vdd.n45 gnd 0.00245f
C1691 vdd.n46 gnd 0.002594f
C1692 vdd.n47 gnd 0.00579f
C1693 vdd.n48 gnd 0.00579f
C1694 vdd.n49 gnd 0.002594f
C1695 vdd.n50 gnd 0.00245f
C1696 vdd.n51 gnd 0.004559f
C1697 vdd.n52 gnd 0.004559f
C1698 vdd.n53 gnd 0.00245f
C1699 vdd.n54 gnd 0.002594f
C1700 vdd.n55 gnd 0.00579f
C1701 vdd.n56 gnd 0.00579f
C1702 vdd.n57 gnd 0.002594f
C1703 vdd.n58 gnd 0.00245f
C1704 vdd.n59 gnd 0.004559f
C1705 vdd.n60 gnd 0.004559f
C1706 vdd.n61 gnd 0.00245f
C1707 vdd.n62 gnd 0.002594f
C1708 vdd.n63 gnd 0.00579f
C1709 vdd.n64 gnd 0.00579f
C1710 vdd.n65 gnd 0.013689f
C1711 vdd.n66 gnd 0.002522f
C1712 vdd.n67 gnd 0.00245f
C1713 vdd.n68 gnd 0.011783f
C1714 vdd.n69 gnd 0.008226f
C1715 vdd.t124 gnd 0.02882f
C1716 vdd.t122 gnd 0.02882f
C1717 vdd.n70 gnd 0.198072f
C1718 vdd.n71 gnd 0.155753f
C1719 vdd.t243 gnd 0.02882f
C1720 vdd.t160 gnd 0.02882f
C1721 vdd.n72 gnd 0.198072f
C1722 vdd.n73 gnd 0.125692f
C1723 vdd.t102 gnd 0.02882f
C1724 vdd.t89 gnd 0.02882f
C1725 vdd.n74 gnd 0.198072f
C1726 vdd.n75 gnd 0.125692f
C1727 vdd.t240 gnd 0.02882f
C1728 vdd.t136 gnd 0.02882f
C1729 vdd.n76 gnd 0.198072f
C1730 vdd.n77 gnd 0.125692f
C1731 vdd.t99 gnd 0.02882f
C1732 vdd.t241 gnd 0.02882f
C1733 vdd.n78 gnd 0.198072f
C1734 vdd.n79 gnd 0.125692f
C1735 vdd.n80 gnd 0.004913f
C1736 vdd.n81 gnd 0.004559f
C1737 vdd.n82 gnd 0.002522f
C1738 vdd.n83 gnd 0.00579f
C1739 vdd.n84 gnd 0.00245f
C1740 vdd.n85 gnd 0.002594f
C1741 vdd.n86 gnd 0.004559f
C1742 vdd.n87 gnd 0.00245f
C1743 vdd.n88 gnd 0.00579f
C1744 vdd.n89 gnd 0.002594f
C1745 vdd.n90 gnd 0.004559f
C1746 vdd.n91 gnd 0.00245f
C1747 vdd.n92 gnd 0.004343f
C1748 vdd.n93 gnd 0.004356f
C1749 vdd.t118 gnd 0.01244f
C1750 vdd.n94 gnd 0.027678f
C1751 vdd.n95 gnd 0.144045f
C1752 vdd.n96 gnd 0.00245f
C1753 vdd.n97 gnd 0.002594f
C1754 vdd.n98 gnd 0.00579f
C1755 vdd.n99 gnd 0.00579f
C1756 vdd.n100 gnd 0.002594f
C1757 vdd.n101 gnd 0.00245f
C1758 vdd.n102 gnd 0.004559f
C1759 vdd.n103 gnd 0.004559f
C1760 vdd.n104 gnd 0.00245f
C1761 vdd.n105 gnd 0.002594f
C1762 vdd.n106 gnd 0.00579f
C1763 vdd.n107 gnd 0.00579f
C1764 vdd.n108 gnd 0.002594f
C1765 vdd.n109 gnd 0.00245f
C1766 vdd.n110 gnd 0.004559f
C1767 vdd.n111 gnd 0.004559f
C1768 vdd.n112 gnd 0.00245f
C1769 vdd.n113 gnd 0.002594f
C1770 vdd.n114 gnd 0.00579f
C1771 vdd.n115 gnd 0.00579f
C1772 vdd.n116 gnd 0.013689f
C1773 vdd.n117 gnd 0.002522f
C1774 vdd.n118 gnd 0.00245f
C1775 vdd.n119 gnd 0.011783f
C1776 vdd.n120 gnd 0.007968f
C1777 vdd.n121 gnd 0.093515f
C1778 vdd.n122 gnd 0.004913f
C1779 vdd.n123 gnd 0.004559f
C1780 vdd.n124 gnd 0.002522f
C1781 vdd.n125 gnd 0.00579f
C1782 vdd.n126 gnd 0.00245f
C1783 vdd.n127 gnd 0.002594f
C1784 vdd.n128 gnd 0.004559f
C1785 vdd.n129 gnd 0.00245f
C1786 vdd.n130 gnd 0.00579f
C1787 vdd.n131 gnd 0.002594f
C1788 vdd.n132 gnd 0.004559f
C1789 vdd.n133 gnd 0.00245f
C1790 vdd.n134 gnd 0.004343f
C1791 vdd.n135 gnd 0.004356f
C1792 vdd.t114 gnd 0.01244f
C1793 vdd.n136 gnd 0.027678f
C1794 vdd.n137 gnd 0.144045f
C1795 vdd.n138 gnd 0.00245f
C1796 vdd.n139 gnd 0.002594f
C1797 vdd.n140 gnd 0.00579f
C1798 vdd.n141 gnd 0.00579f
C1799 vdd.n142 gnd 0.002594f
C1800 vdd.n143 gnd 0.00245f
C1801 vdd.n144 gnd 0.004559f
C1802 vdd.n145 gnd 0.004559f
C1803 vdd.n146 gnd 0.00245f
C1804 vdd.n147 gnd 0.002594f
C1805 vdd.n148 gnd 0.00579f
C1806 vdd.n149 gnd 0.00579f
C1807 vdd.n150 gnd 0.002594f
C1808 vdd.n151 gnd 0.00245f
C1809 vdd.n152 gnd 0.004559f
C1810 vdd.n153 gnd 0.004559f
C1811 vdd.n154 gnd 0.00245f
C1812 vdd.n155 gnd 0.002594f
C1813 vdd.n156 gnd 0.00579f
C1814 vdd.n157 gnd 0.00579f
C1815 vdd.n158 gnd 0.013689f
C1816 vdd.n159 gnd 0.002522f
C1817 vdd.n160 gnd 0.00245f
C1818 vdd.n161 gnd 0.011783f
C1819 vdd.n162 gnd 0.008226f
C1820 vdd.t113 gnd 0.02882f
C1821 vdd.t168 gnd 0.02882f
C1822 vdd.n163 gnd 0.198072f
C1823 vdd.n164 gnd 0.155753f
C1824 vdd.t148 gnd 0.02882f
C1825 vdd.t129 gnd 0.02882f
C1826 vdd.n165 gnd 0.198072f
C1827 vdd.n166 gnd 0.125692f
C1828 vdd.t108 gnd 0.02882f
C1829 vdd.t228 gnd 0.02882f
C1830 vdd.n167 gnd 0.198072f
C1831 vdd.n168 gnd 0.125692f
C1832 vdd.t242 gnd 0.02882f
C1833 vdd.t230 gnd 0.02882f
C1834 vdd.n169 gnd 0.198072f
C1835 vdd.n170 gnd 0.125692f
C1836 vdd.t138 gnd 0.02882f
C1837 vdd.t232 gnd 0.02882f
C1838 vdd.n171 gnd 0.198072f
C1839 vdd.n172 gnd 0.125692f
C1840 vdd.n173 gnd 0.004913f
C1841 vdd.n174 gnd 0.004559f
C1842 vdd.n175 gnd 0.002522f
C1843 vdd.n176 gnd 0.00579f
C1844 vdd.n177 gnd 0.00245f
C1845 vdd.n178 gnd 0.002594f
C1846 vdd.n179 gnd 0.004559f
C1847 vdd.n180 gnd 0.00245f
C1848 vdd.n181 gnd 0.00579f
C1849 vdd.n182 gnd 0.002594f
C1850 vdd.n183 gnd 0.004559f
C1851 vdd.n184 gnd 0.00245f
C1852 vdd.n185 gnd 0.004343f
C1853 vdd.n186 gnd 0.004356f
C1854 vdd.t145 gnd 0.01244f
C1855 vdd.n187 gnd 0.027678f
C1856 vdd.n188 gnd 0.144045f
C1857 vdd.n189 gnd 0.00245f
C1858 vdd.n190 gnd 0.002594f
C1859 vdd.n191 gnd 0.00579f
C1860 vdd.n192 gnd 0.00579f
C1861 vdd.n193 gnd 0.002594f
C1862 vdd.n194 gnd 0.00245f
C1863 vdd.n195 gnd 0.004559f
C1864 vdd.n196 gnd 0.004559f
C1865 vdd.n197 gnd 0.00245f
C1866 vdd.n198 gnd 0.002594f
C1867 vdd.n199 gnd 0.00579f
C1868 vdd.n200 gnd 0.00579f
C1869 vdd.n201 gnd 0.002594f
C1870 vdd.n202 gnd 0.00245f
C1871 vdd.n203 gnd 0.004559f
C1872 vdd.n204 gnd 0.004559f
C1873 vdd.n205 gnd 0.00245f
C1874 vdd.n206 gnd 0.002594f
C1875 vdd.n207 gnd 0.00579f
C1876 vdd.n208 gnd 0.00579f
C1877 vdd.n209 gnd 0.013689f
C1878 vdd.n210 gnd 0.002522f
C1879 vdd.n211 gnd 0.00245f
C1880 vdd.n212 gnd 0.011783f
C1881 vdd.n213 gnd 0.007968f
C1882 vdd.n214 gnd 0.055632f
C1883 vdd.n215 gnd 0.200457f
C1884 vdd.n216 gnd 0.004913f
C1885 vdd.n217 gnd 0.004559f
C1886 vdd.n218 gnd 0.002522f
C1887 vdd.n219 gnd 0.00579f
C1888 vdd.n220 gnd 0.00245f
C1889 vdd.n221 gnd 0.002594f
C1890 vdd.n222 gnd 0.004559f
C1891 vdd.n223 gnd 0.00245f
C1892 vdd.n224 gnd 0.00579f
C1893 vdd.n225 gnd 0.002594f
C1894 vdd.n226 gnd 0.004559f
C1895 vdd.n227 gnd 0.00245f
C1896 vdd.n228 gnd 0.004343f
C1897 vdd.n229 gnd 0.004356f
C1898 vdd.t238 gnd 0.01244f
C1899 vdd.n230 gnd 0.027678f
C1900 vdd.n231 gnd 0.144045f
C1901 vdd.n232 gnd 0.00245f
C1902 vdd.n233 gnd 0.002594f
C1903 vdd.n234 gnd 0.00579f
C1904 vdd.n235 gnd 0.00579f
C1905 vdd.n236 gnd 0.002594f
C1906 vdd.n237 gnd 0.00245f
C1907 vdd.n238 gnd 0.004559f
C1908 vdd.n239 gnd 0.004559f
C1909 vdd.n240 gnd 0.00245f
C1910 vdd.n241 gnd 0.002594f
C1911 vdd.n242 gnd 0.00579f
C1912 vdd.n243 gnd 0.00579f
C1913 vdd.n244 gnd 0.002594f
C1914 vdd.n245 gnd 0.00245f
C1915 vdd.n246 gnd 0.004559f
C1916 vdd.n247 gnd 0.004559f
C1917 vdd.n248 gnd 0.00245f
C1918 vdd.n249 gnd 0.002594f
C1919 vdd.n250 gnd 0.00579f
C1920 vdd.n251 gnd 0.00579f
C1921 vdd.n252 gnd 0.013689f
C1922 vdd.n253 gnd 0.002522f
C1923 vdd.n254 gnd 0.00245f
C1924 vdd.n255 gnd 0.011783f
C1925 vdd.n256 gnd 0.008226f
C1926 vdd.t237 gnd 0.02882f
C1927 vdd.t132 gnd 0.02882f
C1928 vdd.n257 gnd 0.198072f
C1929 vdd.n258 gnd 0.155753f
C1930 vdd.t131 gnd 0.02882f
C1931 vdd.t231 gnd 0.02882f
C1932 vdd.n259 gnd 0.198072f
C1933 vdd.n260 gnd 0.125692f
C1934 vdd.t103 gnd 0.02882f
C1935 vdd.t162 gnd 0.02882f
C1936 vdd.n261 gnd 0.198072f
C1937 vdd.n262 gnd 0.125692f
C1938 vdd.t87 gnd 0.02882f
C1939 vdd.t7 gnd 0.02882f
C1940 vdd.n263 gnd 0.198072f
C1941 vdd.n264 gnd 0.125692f
C1942 vdd.t146 gnd 0.02882f
C1943 vdd.t95 gnd 0.02882f
C1944 vdd.n265 gnd 0.198072f
C1945 vdd.n266 gnd 0.125692f
C1946 vdd.n267 gnd 0.004913f
C1947 vdd.n268 gnd 0.004559f
C1948 vdd.n269 gnd 0.002522f
C1949 vdd.n270 gnd 0.00579f
C1950 vdd.n271 gnd 0.00245f
C1951 vdd.n272 gnd 0.002594f
C1952 vdd.n273 gnd 0.004559f
C1953 vdd.n274 gnd 0.00245f
C1954 vdd.n275 gnd 0.00579f
C1955 vdd.n276 gnd 0.002594f
C1956 vdd.n277 gnd 0.004559f
C1957 vdd.n278 gnd 0.00245f
C1958 vdd.n279 gnd 0.004343f
C1959 vdd.n280 gnd 0.004356f
C1960 vdd.t156 gnd 0.01244f
C1961 vdd.n281 gnd 0.027678f
C1962 vdd.n282 gnd 0.144045f
C1963 vdd.n283 gnd 0.00245f
C1964 vdd.n284 gnd 0.002594f
C1965 vdd.n285 gnd 0.00579f
C1966 vdd.n286 gnd 0.00579f
C1967 vdd.n287 gnd 0.002594f
C1968 vdd.n288 gnd 0.00245f
C1969 vdd.n289 gnd 0.004559f
C1970 vdd.n290 gnd 0.004559f
C1971 vdd.n291 gnd 0.00245f
C1972 vdd.n292 gnd 0.002594f
C1973 vdd.n293 gnd 0.00579f
C1974 vdd.n294 gnd 0.00579f
C1975 vdd.n295 gnd 0.002594f
C1976 vdd.n296 gnd 0.00245f
C1977 vdd.n297 gnd 0.004559f
C1978 vdd.n298 gnd 0.004559f
C1979 vdd.n299 gnd 0.00245f
C1980 vdd.n300 gnd 0.002594f
C1981 vdd.n301 gnd 0.00579f
C1982 vdd.n302 gnd 0.00579f
C1983 vdd.n303 gnd 0.013689f
C1984 vdd.n304 gnd 0.002522f
C1985 vdd.n305 gnd 0.00245f
C1986 vdd.n306 gnd 0.011783f
C1987 vdd.n307 gnd 0.007968f
C1988 vdd.n308 gnd 0.055632f
C1989 vdd.n309 gnd 0.220309f
C1990 vdd.n310 gnd 0.008921f
C1991 vdd.n311 gnd 0.008921f
C1992 vdd.n312 gnd 0.007205f
C1993 vdd.n313 gnd 0.007205f
C1994 vdd.n314 gnd 0.008952f
C1995 vdd.n315 gnd 0.008952f
C1996 vdd.t101 gnd 0.45741f
C1997 vdd.n316 gnd 0.008952f
C1998 vdd.n317 gnd 0.008952f
C1999 vdd.n318 gnd 0.008952f
C2000 vdd.t86 gnd 0.45741f
C2001 vdd.n319 gnd 0.008952f
C2002 vdd.n320 gnd 0.008952f
C2003 vdd.n321 gnd 0.008952f
C2004 vdd.n322 gnd 0.008952f
C2005 vdd.n323 gnd 0.007205f
C2006 vdd.n324 gnd 0.008952f
C2007 vdd.n325 gnd 0.73643f
C2008 vdd.n326 gnd 0.008952f
C2009 vdd.n327 gnd 0.008952f
C2010 vdd.n328 gnd 0.008952f
C2011 vdd.n329 gnd 0.626652f
C2012 vdd.n330 gnd 0.008952f
C2013 vdd.n331 gnd 0.008952f
C2014 vdd.n332 gnd 0.008952f
C2015 vdd.n333 gnd 0.008952f
C2016 vdd.n334 gnd 0.008952f
C2017 vdd.n335 gnd 0.007205f
C2018 vdd.n336 gnd 0.008952f
C2019 vdd.t94 gnd 0.45741f
C2020 vdd.n337 gnd 0.008952f
C2021 vdd.n338 gnd 0.008952f
C2022 vdd.n339 gnd 0.008952f
C2023 vdd.n340 gnd 0.91482f
C2024 vdd.n341 gnd 0.008952f
C2025 vdd.n342 gnd 0.008952f
C2026 vdd.n343 gnd 0.008952f
C2027 vdd.n344 gnd 0.008952f
C2028 vdd.n345 gnd 0.008952f
C2029 vdd.n346 gnd 0.007205f
C2030 vdd.n347 gnd 0.008952f
C2031 vdd.n348 gnd 0.008952f
C2032 vdd.n349 gnd 0.008952f
C2033 vdd.n350 gnd 0.021096f
C2034 vdd.n351 gnd 2.10409f
C2035 vdd.n352 gnd 0.021425f
C2036 vdd.n353 gnd 0.008952f
C2037 vdd.n354 gnd 0.008952f
C2038 vdd.n356 gnd 0.008952f
C2039 vdd.n357 gnd 0.008952f
C2040 vdd.n358 gnd 0.007205f
C2041 vdd.n359 gnd 0.007205f
C2042 vdd.n360 gnd 0.008952f
C2043 vdd.n361 gnd 0.008952f
C2044 vdd.n362 gnd 0.008952f
C2045 vdd.n363 gnd 0.008952f
C2046 vdd.n364 gnd 0.008952f
C2047 vdd.n365 gnd 0.008952f
C2048 vdd.n366 gnd 0.007205f
C2049 vdd.n368 gnd 0.008952f
C2050 vdd.n369 gnd 0.008952f
C2051 vdd.n370 gnd 0.008952f
C2052 vdd.n371 gnd 0.008952f
C2053 vdd.n372 gnd 0.008952f
C2054 vdd.n373 gnd 0.007205f
C2055 vdd.n375 gnd 0.008952f
C2056 vdd.n376 gnd 0.008952f
C2057 vdd.n377 gnd 0.008952f
C2058 vdd.n378 gnd 0.008952f
C2059 vdd.n379 gnd 0.008952f
C2060 vdd.n380 gnd 0.007205f
C2061 vdd.n382 gnd 0.008952f
C2062 vdd.n383 gnd 0.008952f
C2063 vdd.n384 gnd 0.008952f
C2064 vdd.n385 gnd 0.008952f
C2065 vdd.n386 gnd 0.006016f
C2066 vdd.t52 gnd 0.110129f
C2067 vdd.t51 gnd 0.117698f
C2068 vdd.t50 gnd 0.143827f
C2069 vdd.n387 gnd 0.184366f
C2070 vdd.n388 gnd 0.155622f
C2071 vdd.n390 gnd 0.008952f
C2072 vdd.n391 gnd 0.008952f
C2073 vdd.n392 gnd 0.007205f
C2074 vdd.n393 gnd 0.008952f
C2075 vdd.n395 gnd 0.008952f
C2076 vdd.n396 gnd 0.008952f
C2077 vdd.n397 gnd 0.008952f
C2078 vdd.n398 gnd 0.008952f
C2079 vdd.n399 gnd 0.007205f
C2080 vdd.n401 gnd 0.008952f
C2081 vdd.n402 gnd 0.008952f
C2082 vdd.n403 gnd 0.008952f
C2083 vdd.n404 gnd 0.008952f
C2084 vdd.n405 gnd 0.008952f
C2085 vdd.n406 gnd 0.007205f
C2086 vdd.n408 gnd 0.008952f
C2087 vdd.n409 gnd 0.008952f
C2088 vdd.n410 gnd 0.008952f
C2089 vdd.n411 gnd 0.008952f
C2090 vdd.n412 gnd 0.008952f
C2091 vdd.n413 gnd 0.007205f
C2092 vdd.n415 gnd 0.008952f
C2093 vdd.n416 gnd 0.008952f
C2094 vdd.n417 gnd 0.008952f
C2095 vdd.n418 gnd 0.008952f
C2096 vdd.n419 gnd 0.008952f
C2097 vdd.n420 gnd 0.007205f
C2098 vdd.n422 gnd 0.008952f
C2099 vdd.n423 gnd 0.008952f
C2100 vdd.n424 gnd 0.008952f
C2101 vdd.n425 gnd 0.008952f
C2102 vdd.n426 gnd 0.007133f
C2103 vdd.t35 gnd 0.110129f
C2104 vdd.t34 gnd 0.117698f
C2105 vdd.t32 gnd 0.143827f
C2106 vdd.n427 gnd 0.184366f
C2107 vdd.n428 gnd 0.155622f
C2108 vdd.n430 gnd 0.008952f
C2109 vdd.n431 gnd 0.008952f
C2110 vdd.n432 gnd 0.007205f
C2111 vdd.n433 gnd 0.008952f
C2112 vdd.n435 gnd 0.008952f
C2113 vdd.n436 gnd 0.008952f
C2114 vdd.n437 gnd 0.008952f
C2115 vdd.n438 gnd 0.008952f
C2116 vdd.n439 gnd 0.007205f
C2117 vdd.n441 gnd 0.008952f
C2118 vdd.n442 gnd 0.008952f
C2119 vdd.n443 gnd 0.008952f
C2120 vdd.n444 gnd 0.008952f
C2121 vdd.n445 gnd 0.008952f
C2122 vdd.n446 gnd 0.007205f
C2123 vdd.n448 gnd 0.008952f
C2124 vdd.n449 gnd 0.008952f
C2125 vdd.n450 gnd 0.008952f
C2126 vdd.n451 gnd 0.008952f
C2127 vdd.n452 gnd 0.008952f
C2128 vdd.n453 gnd 0.007205f
C2129 vdd.n455 gnd 0.008952f
C2130 vdd.n456 gnd 0.008952f
C2131 vdd.n457 gnd 0.008952f
C2132 vdd.n458 gnd 0.008952f
C2133 vdd.n459 gnd 0.008952f
C2134 vdd.n460 gnd 0.007205f
C2135 vdd.n462 gnd 0.008952f
C2136 vdd.n463 gnd 0.008952f
C2137 vdd.n464 gnd 0.008952f
C2138 vdd.n465 gnd 0.008952f
C2139 vdd.n466 gnd 0.008952f
C2140 vdd.n467 gnd 0.008952f
C2141 vdd.n468 gnd 0.007205f
C2142 vdd.n469 gnd 0.008952f
C2143 vdd.n470 gnd 0.008952f
C2144 vdd.n471 gnd 0.007205f
C2145 vdd.n472 gnd 0.008952f
C2146 vdd.n473 gnd 0.008952f
C2147 vdd.n474 gnd 0.007205f
C2148 vdd.n475 gnd 0.008952f
C2149 vdd.n476 gnd 0.007205f
C2150 vdd.n477 gnd 0.008952f
C2151 vdd.n478 gnd 0.007205f
C2152 vdd.n479 gnd 0.008952f
C2153 vdd.n480 gnd 0.008952f
C2154 vdd.t128 gnd 0.45741f
C2155 vdd.n481 gnd 0.489429f
C2156 vdd.n482 gnd 0.008952f
C2157 vdd.n483 gnd 0.007205f
C2158 vdd.n484 gnd 0.008952f
C2159 vdd.n485 gnd 0.007205f
C2160 vdd.n486 gnd 0.008952f
C2161 vdd.t130 gnd 0.45741f
C2162 vdd.n487 gnd 0.008952f
C2163 vdd.n488 gnd 0.007205f
C2164 vdd.n489 gnd 0.008952f
C2165 vdd.n490 gnd 0.007205f
C2166 vdd.n491 gnd 0.008952f
C2167 vdd.n492 gnd 0.718134f
C2168 vdd.n493 gnd 0.759301f
C2169 vdd.t121 gnd 0.45741f
C2170 vdd.n494 gnd 0.008952f
C2171 vdd.n495 gnd 0.007205f
C2172 vdd.n496 gnd 0.008952f
C2173 vdd.n497 gnd 0.007205f
C2174 vdd.n498 gnd 0.008952f
C2175 vdd.n499 gnd 0.562614f
C2176 vdd.n500 gnd 0.008952f
C2177 vdd.n501 gnd 0.007205f
C2178 vdd.n502 gnd 0.008952f
C2179 vdd.n503 gnd 0.007205f
C2180 vdd.n504 gnd 0.008952f
C2181 vdd.n505 gnd 0.91482f
C2182 vdd.t4 gnd 0.45741f
C2183 vdd.n506 gnd 0.008952f
C2184 vdd.n507 gnd 0.007205f
C2185 vdd.n508 gnd 0.008952f
C2186 vdd.n509 gnd 0.007205f
C2187 vdd.n510 gnd 0.008952f
C2188 vdd.n511 gnd 0.489429f
C2189 vdd.n512 gnd 0.008952f
C2190 vdd.n513 gnd 0.007205f
C2191 vdd.n514 gnd 0.021425f
C2192 vdd.n515 gnd 0.021425f
C2193 vdd.n516 gnd 11.105901f
C2194 vdd.t29 gnd 0.45741f
C2195 vdd.n517 gnd 0.021425f
C2196 vdd.n518 gnd 0.007698f
C2197 vdd.n519 gnd 0.007205f
C2198 vdd.n524 gnd 0.005729f
C2199 vdd.n525 gnd 0.007205f
C2200 vdd.n526 gnd 0.008952f
C2201 vdd.n527 gnd 0.008952f
C2202 vdd.n528 gnd 0.008952f
C2203 vdd.n529 gnd 0.008952f
C2204 vdd.n530 gnd 0.008952f
C2205 vdd.n531 gnd 0.007205f
C2206 vdd.n532 gnd 0.008952f
C2207 vdd.n533 gnd 0.008952f
C2208 vdd.n534 gnd 0.008952f
C2209 vdd.n535 gnd 0.008952f
C2210 vdd.n536 gnd 0.008952f
C2211 vdd.n537 gnd 0.007205f
C2212 vdd.n538 gnd 0.008952f
C2213 vdd.n539 gnd 0.008952f
C2214 vdd.n540 gnd 0.008952f
C2215 vdd.n541 gnd 0.008952f
C2216 vdd.n542 gnd 0.008952f
C2217 vdd.t64 gnd 0.110129f
C2218 vdd.t65 gnd 0.117698f
C2219 vdd.t63 gnd 0.143827f
C2220 vdd.n543 gnd 0.184366f
C2221 vdd.n544 gnd 0.154901f
C2222 vdd.n545 gnd 0.014698f
C2223 vdd.n546 gnd 0.008952f
C2224 vdd.n547 gnd 0.008952f
C2225 vdd.n548 gnd 0.008952f
C2226 vdd.n549 gnd 0.008952f
C2227 vdd.n550 gnd 0.008952f
C2228 vdd.n551 gnd 0.007205f
C2229 vdd.n552 gnd 0.008952f
C2230 vdd.n553 gnd 0.008952f
C2231 vdd.n554 gnd 0.008952f
C2232 vdd.n555 gnd 0.008952f
C2233 vdd.n556 gnd 0.008952f
C2234 vdd.n557 gnd 0.007205f
C2235 vdd.n558 gnd 0.008952f
C2236 vdd.n559 gnd 0.008952f
C2237 vdd.n560 gnd 0.008952f
C2238 vdd.n561 gnd 0.008952f
C2239 vdd.n562 gnd 0.008952f
C2240 vdd.n563 gnd 0.007205f
C2241 vdd.n564 gnd 0.008952f
C2242 vdd.n565 gnd 0.008952f
C2243 vdd.n566 gnd 0.008952f
C2244 vdd.n567 gnd 0.008952f
C2245 vdd.n568 gnd 0.008952f
C2246 vdd.n569 gnd 0.007205f
C2247 vdd.n570 gnd 0.008952f
C2248 vdd.n571 gnd 0.008952f
C2249 vdd.n572 gnd 0.008952f
C2250 vdd.n573 gnd 0.008952f
C2251 vdd.n574 gnd 0.008952f
C2252 vdd.n575 gnd 0.007205f
C2253 vdd.n576 gnd 0.008952f
C2254 vdd.n577 gnd 0.008952f
C2255 vdd.n578 gnd 0.008952f
C2256 vdd.n579 gnd 0.007133f
C2257 vdd.t54 gnd 0.110129f
C2258 vdd.t55 gnd 0.117698f
C2259 vdd.t53 gnd 0.143827f
C2260 vdd.n580 gnd 0.184366f
C2261 vdd.n581 gnd 0.154901f
C2262 vdd.n582 gnd 0.008952f
C2263 vdd.n583 gnd 0.007205f
C2264 vdd.n585 gnd 0.008952f
C2265 vdd.n587 gnd 0.008952f
C2266 vdd.n588 gnd 0.008952f
C2267 vdd.n589 gnd 0.007205f
C2268 vdd.n590 gnd 0.008952f
C2269 vdd.n591 gnd 0.008952f
C2270 vdd.n592 gnd 0.008952f
C2271 vdd.n593 gnd 0.008952f
C2272 vdd.n594 gnd 0.008952f
C2273 vdd.n595 gnd 0.007205f
C2274 vdd.n596 gnd 0.008952f
C2275 vdd.n597 gnd 0.008952f
C2276 vdd.n598 gnd 0.008952f
C2277 vdd.n599 gnd 0.008952f
C2278 vdd.n600 gnd 0.008952f
C2279 vdd.n601 gnd 0.007205f
C2280 vdd.n602 gnd 0.008952f
C2281 vdd.n603 gnd 0.008952f
C2282 vdd.n604 gnd 0.008952f
C2283 vdd.n605 gnd 0.005729f
C2284 vdd.n610 gnd 0.006087f
C2285 vdd.n611 gnd 0.006087f
C2286 vdd.n612 gnd 0.006087f
C2287 vdd.n613 gnd 10.804f
C2288 vdd.n614 gnd 0.006087f
C2289 vdd.n615 gnd 0.006087f
C2290 vdd.n616 gnd 0.006087f
C2291 vdd.n618 gnd 0.006087f
C2292 vdd.n619 gnd 0.006087f
C2293 vdd.n621 gnd 0.006087f
C2294 vdd.n622 gnd 0.004431f
C2295 vdd.n624 gnd 0.006087f
C2296 vdd.t13 gnd 0.245981f
C2297 vdd.t12 gnd 0.251792f
C2298 vdd.t10 gnd 0.160586f
C2299 vdd.n625 gnd 0.086788f
C2300 vdd.n626 gnd 0.049229f
C2301 vdd.n627 gnd 0.0087f
C2302 vdd.n628 gnd 0.013821f
C2303 vdd.n630 gnd 0.006087f
C2304 vdd.n631 gnd 0.622078f
C2305 vdd.n632 gnd 0.013034f
C2306 vdd.n633 gnd 0.013034f
C2307 vdd.n634 gnd 0.006087f
C2308 vdd.n635 gnd 0.013821f
C2309 vdd.n636 gnd 0.006087f
C2310 vdd.n637 gnd 0.006087f
C2311 vdd.n638 gnd 0.006087f
C2312 vdd.n639 gnd 0.006087f
C2313 vdd.n640 gnd 0.006087f
C2314 vdd.n642 gnd 0.006087f
C2315 vdd.n643 gnd 0.006087f
C2316 vdd.n645 gnd 0.006087f
C2317 vdd.n646 gnd 0.006087f
C2318 vdd.n648 gnd 0.006087f
C2319 vdd.n649 gnd 0.006087f
C2320 vdd.n651 gnd 0.006087f
C2321 vdd.n652 gnd 0.006087f
C2322 vdd.n654 gnd 0.006087f
C2323 vdd.n655 gnd 0.006087f
C2324 vdd.n657 gnd 0.006087f
C2325 vdd.n658 gnd 0.004431f
C2326 vdd.n660 gnd 0.006087f
C2327 vdd.t27 gnd 0.245981f
C2328 vdd.t26 gnd 0.251792f
C2329 vdd.t25 gnd 0.160586f
C2330 vdd.n661 gnd 0.086788f
C2331 vdd.n662 gnd 0.049229f
C2332 vdd.n663 gnd 0.0087f
C2333 vdd.n664 gnd 0.006087f
C2334 vdd.n665 gnd 0.006087f
C2335 vdd.t11 gnd 0.311039f
C2336 vdd.n666 gnd 0.006087f
C2337 vdd.n667 gnd 0.006087f
C2338 vdd.n668 gnd 0.006087f
C2339 vdd.n669 gnd 0.006087f
C2340 vdd.n670 gnd 0.006087f
C2341 vdd.n671 gnd 0.622078f
C2342 vdd.n672 gnd 0.006087f
C2343 vdd.n673 gnd 0.006087f
C2344 vdd.n674 gnd 0.489429f
C2345 vdd.n675 gnd 0.006087f
C2346 vdd.n676 gnd 0.006087f
C2347 vdd.n677 gnd 0.006087f
C2348 vdd.n678 gnd 0.006087f
C2349 vdd.n679 gnd 0.622078f
C2350 vdd.n680 gnd 0.006087f
C2351 vdd.n681 gnd 0.006087f
C2352 vdd.n682 gnd 0.006087f
C2353 vdd.n683 gnd 0.006087f
C2354 vdd.n684 gnd 0.006087f
C2355 vdd.t186 gnd 0.311039f
C2356 vdd.n685 gnd 0.006087f
C2357 vdd.n686 gnd 0.006087f
C2358 vdd.n687 gnd 0.006087f
C2359 vdd.n688 gnd 0.006087f
C2360 vdd.n689 gnd 0.006087f
C2361 vdd.t203 gnd 0.311039f
C2362 vdd.n690 gnd 0.006087f
C2363 vdd.n691 gnd 0.006087f
C2364 vdd.n692 gnd 0.599207f
C2365 vdd.n693 gnd 0.006087f
C2366 vdd.n694 gnd 0.006087f
C2367 vdd.n695 gnd 0.006087f
C2368 vdd.t202 gnd 0.311039f
C2369 vdd.n696 gnd 0.006087f
C2370 vdd.n697 gnd 0.006087f
C2371 vdd.n698 gnd 0.461984f
C2372 vdd.n699 gnd 0.006087f
C2373 vdd.n700 gnd 0.006087f
C2374 vdd.n701 gnd 0.006087f
C2375 vdd.n702 gnd 0.43454f
C2376 vdd.n703 gnd 0.006087f
C2377 vdd.n704 gnd 0.006087f
C2378 vdd.n705 gnd 0.324761f
C2379 vdd.n706 gnd 0.006087f
C2380 vdd.n707 gnd 0.006087f
C2381 vdd.n708 gnd 0.006087f
C2382 vdd.n709 gnd 0.571763f
C2383 vdd.n710 gnd 0.006087f
C2384 vdd.n711 gnd 0.006087f
C2385 vdd.t209 gnd 0.311039f
C2386 vdd.n712 gnd 0.006087f
C2387 vdd.n713 gnd 0.006087f
C2388 vdd.n714 gnd 0.006087f
C2389 vdd.n715 gnd 0.622078f
C2390 vdd.n716 gnd 0.006087f
C2391 vdd.n717 gnd 0.006087f
C2392 vdd.t210 gnd 0.311039f
C2393 vdd.n718 gnd 0.006087f
C2394 vdd.n719 gnd 0.006087f
C2395 vdd.n720 gnd 0.006087f
C2396 vdd.t180 gnd 0.311039f
C2397 vdd.n721 gnd 0.006087f
C2398 vdd.n722 gnd 0.006087f
C2399 vdd.n723 gnd 0.006087f
C2400 vdd.t38 gnd 0.251792f
C2401 vdd.t36 gnd 0.160586f
C2402 vdd.t39 gnd 0.251792f
C2403 vdd.n724 gnd 0.141517f
C2404 vdd.n725 gnd 0.017634f
C2405 vdd.n726 gnd 0.006087f
C2406 vdd.t37 gnd 0.224131f
C2407 vdd.n727 gnd 0.006087f
C2408 vdd.n728 gnd 0.006087f
C2409 vdd.n729 gnd 0.53517f
C2410 vdd.n730 gnd 0.006087f
C2411 vdd.n731 gnd 0.006087f
C2412 vdd.n732 gnd 0.006087f
C2413 vdd.n733 gnd 0.361354f
C2414 vdd.n734 gnd 0.006087f
C2415 vdd.n735 gnd 0.006087f
C2416 vdd.t181 gnd 0.128075f
C2417 vdd.n736 gnd 0.397947f
C2418 vdd.n737 gnd 0.006087f
C2419 vdd.n738 gnd 0.006087f
C2420 vdd.n739 gnd 0.006087f
C2421 vdd.n740 gnd 0.498577f
C2422 vdd.n741 gnd 0.006087f
C2423 vdd.n742 gnd 0.006087f
C2424 vdd.t194 gnd 0.311039f
C2425 vdd.n743 gnd 0.006087f
C2426 vdd.n744 gnd 0.006087f
C2427 vdd.n745 gnd 0.006087f
C2428 vdd.t190 gnd 0.311039f
C2429 vdd.n746 gnd 0.006087f
C2430 vdd.n747 gnd 0.006087f
C2431 vdd.t213 gnd 0.311039f
C2432 vdd.n748 gnd 0.006087f
C2433 vdd.n749 gnd 0.006087f
C2434 vdd.n750 gnd 0.006087f
C2435 vdd.t172 gnd 0.210409f
C2436 vdd.n751 gnd 0.006087f
C2437 vdd.n752 gnd 0.006087f
C2438 vdd.n753 gnd 0.548892f
C2439 vdd.n754 gnd 0.006087f
C2440 vdd.n755 gnd 0.006087f
C2441 vdd.n756 gnd 0.006087f
C2442 vdd.t214 gnd 0.311039f
C2443 vdd.n757 gnd 0.006087f
C2444 vdd.n758 gnd 0.006087f
C2445 vdd.t226 gnd 0.297317f
C2446 vdd.n759 gnd 0.411669f
C2447 vdd.n760 gnd 0.006087f
C2448 vdd.n761 gnd 0.006087f
C2449 vdd.n762 gnd 0.006087f
C2450 vdd.t176 gnd 0.311039f
C2451 vdd.n763 gnd 0.006087f
C2452 vdd.n764 gnd 0.006087f
C2453 vdd.t218 gnd 0.311039f
C2454 vdd.n765 gnd 0.006087f
C2455 vdd.n766 gnd 0.006087f
C2456 vdd.n767 gnd 0.006087f
C2457 vdd.n768 gnd 0.622078f
C2458 vdd.n769 gnd 0.006087f
C2459 vdd.n770 gnd 0.006087f
C2460 vdd.t198 gnd 0.311039f
C2461 vdd.n771 gnd 0.006087f
C2462 vdd.n772 gnd 0.006087f
C2463 vdd.n773 gnd 0.006087f
C2464 vdd.n774 gnd 0.429965f
C2465 vdd.n775 gnd 0.006087f
C2466 vdd.n776 gnd 0.006087f
C2467 vdd.n777 gnd 0.006087f
C2468 vdd.n778 gnd 0.006087f
C2469 vdd.n779 gnd 0.006087f
C2470 vdd.t67 gnd 0.311039f
C2471 vdd.n780 gnd 0.006087f
C2472 vdd.n781 gnd 0.006087f
C2473 vdd.t178 gnd 0.311039f
C2474 vdd.n782 gnd 0.006087f
C2475 vdd.n783 gnd 0.013034f
C2476 vdd.n784 gnd 0.013034f
C2477 vdd.n785 gnd 0.704411f
C2478 vdd.n786 gnd 0.006087f
C2479 vdd.n787 gnd 0.006087f
C2480 vdd.t207 gnd 0.311039f
C2481 vdd.n788 gnd 0.013034f
C2482 vdd.n789 gnd 0.006087f
C2483 vdd.n790 gnd 0.006087f
C2484 vdd.t220 gnd 0.530596f
C2485 vdd.n808 gnd 0.013821f
C2486 vdd.n826 gnd 0.013034f
C2487 vdd.n827 gnd 0.006087f
C2488 vdd.n828 gnd 0.013034f
C2489 vdd.t85 gnd 0.245981f
C2490 vdd.t84 gnd 0.251792f
C2491 vdd.t83 gnd 0.160586f
C2492 vdd.n829 gnd 0.086788f
C2493 vdd.n830 gnd 0.049229f
C2494 vdd.n831 gnd 0.013821f
C2495 vdd.n832 gnd 0.006087f
C2496 vdd.n833 gnd 0.365928f
C2497 vdd.n834 gnd 0.013034f
C2498 vdd.n835 gnd 0.006087f
C2499 vdd.n836 gnd 0.013821f
C2500 vdd.n837 gnd 0.006087f
C2501 vdd.t62 gnd 0.245981f
C2502 vdd.t61 gnd 0.251792f
C2503 vdd.t59 gnd 0.160586f
C2504 vdd.n838 gnd 0.086788f
C2505 vdd.n839 gnd 0.049229f
C2506 vdd.n840 gnd 0.0087f
C2507 vdd.n841 gnd 0.006087f
C2508 vdd.n842 gnd 0.006087f
C2509 vdd.t60 gnd 0.311039f
C2510 vdd.n843 gnd 0.006087f
C2511 vdd.t222 gnd 0.311039f
C2512 vdd.n844 gnd 0.006087f
C2513 vdd.n845 gnd 0.006087f
C2514 vdd.n846 gnd 0.006087f
C2515 vdd.n847 gnd 0.006087f
C2516 vdd.n848 gnd 0.006087f
C2517 vdd.n849 gnd 0.622078f
C2518 vdd.n850 gnd 0.006087f
C2519 vdd.n851 gnd 0.006087f
C2520 vdd.t192 gnd 0.311039f
C2521 vdd.n852 gnd 0.006087f
C2522 vdd.n853 gnd 0.006087f
C2523 vdd.n854 gnd 0.006087f
C2524 vdd.n855 gnd 0.006087f
C2525 vdd.n856 gnd 0.448262f
C2526 vdd.n857 gnd 0.006087f
C2527 vdd.n858 gnd 0.006087f
C2528 vdd.n859 gnd 0.006087f
C2529 vdd.n860 gnd 0.006087f
C2530 vdd.n861 gnd 0.006087f
C2531 vdd.t173 gnd 0.311039f
C2532 vdd.n862 gnd 0.006087f
C2533 vdd.n863 gnd 0.006087f
C2534 vdd.t211 gnd 0.311039f
C2535 vdd.n864 gnd 0.006087f
C2536 vdd.n865 gnd 0.006087f
C2537 vdd.n866 gnd 0.006087f
C2538 vdd.t195 gnd 0.311039f
C2539 vdd.n867 gnd 0.006087f
C2540 vdd.n868 gnd 0.006087f
C2541 vdd.t174 gnd 0.311039f
C2542 vdd.n869 gnd 0.006087f
C2543 vdd.n870 gnd 0.006087f
C2544 vdd.n871 gnd 0.006087f
C2545 vdd.t196 gnd 0.297317f
C2546 vdd.n872 gnd 0.006087f
C2547 vdd.n873 gnd 0.006087f
C2548 vdd.n874 gnd 0.461984f
C2549 vdd.n875 gnd 0.006087f
C2550 vdd.n876 gnd 0.006087f
C2551 vdd.n877 gnd 0.006087f
C2552 vdd.t215 gnd 0.311039f
C2553 vdd.n878 gnd 0.006087f
C2554 vdd.n879 gnd 0.006087f
C2555 vdd.t183 gnd 0.210409f
C2556 vdd.n880 gnd 0.324761f
C2557 vdd.n881 gnd 0.006087f
C2558 vdd.n882 gnd 0.006087f
C2559 vdd.n883 gnd 0.006087f
C2560 vdd.n884 gnd 0.571763f
C2561 vdd.n885 gnd 0.006087f
C2562 vdd.n886 gnd 0.006087f
C2563 vdd.t224 gnd 0.311039f
C2564 vdd.n887 gnd 0.006087f
C2565 vdd.n888 gnd 0.006087f
C2566 vdd.n889 gnd 0.006087f
C2567 vdd.n890 gnd 0.622078f
C2568 vdd.n891 gnd 0.006087f
C2569 vdd.n892 gnd 0.006087f
C2570 vdd.t189 gnd 0.311039f
C2571 vdd.n893 gnd 0.006087f
C2572 vdd.n894 gnd 0.006087f
C2573 vdd.n895 gnd 0.006087f
C2574 vdd.t182 gnd 0.128075f
C2575 vdd.n896 gnd 0.006087f
C2576 vdd.n897 gnd 0.006087f
C2577 vdd.n898 gnd 0.006087f
C2578 vdd.t75 gnd 0.251792f
C2579 vdd.t73 gnd 0.160586f
C2580 vdd.t76 gnd 0.251792f
C2581 vdd.n899 gnd 0.141517f
C2582 vdd.n900 gnd 0.006087f
C2583 vdd.n901 gnd 0.006087f
C2584 vdd.t204 gnd 0.311039f
C2585 vdd.n902 gnd 0.006087f
C2586 vdd.n903 gnd 0.006087f
C2587 vdd.t74 gnd 0.224131f
C2588 vdd.n904 gnd 0.494003f
C2589 vdd.n905 gnd 0.006087f
C2590 vdd.n906 gnd 0.006087f
C2591 vdd.n907 gnd 0.006087f
C2592 vdd.n908 gnd 0.361354f
C2593 vdd.n909 gnd 0.006087f
C2594 vdd.n910 gnd 0.006087f
C2595 vdd.n911 gnd 0.397947f
C2596 vdd.n912 gnd 0.006087f
C2597 vdd.n913 gnd 0.006087f
C2598 vdd.n914 gnd 0.006087f
C2599 vdd.n915 gnd 0.498577f
C2600 vdd.n916 gnd 0.006087f
C2601 vdd.n917 gnd 0.006087f
C2602 vdd.t184 gnd 0.311039f
C2603 vdd.n918 gnd 0.006087f
C2604 vdd.n919 gnd 0.006087f
C2605 vdd.n920 gnd 0.006087f
C2606 vdd.n921 gnd 0.622078f
C2607 vdd.n922 gnd 0.006087f
C2608 vdd.n923 gnd 0.006087f
C2609 vdd.t185 gnd 0.311039f
C2610 vdd.n924 gnd 0.006087f
C2611 vdd.n925 gnd 0.006087f
C2612 vdd.n926 gnd 0.006087f
C2613 vdd.t225 gnd 0.311039f
C2614 vdd.n927 gnd 0.006087f
C2615 vdd.n928 gnd 0.006087f
C2616 vdd.n929 gnd 0.006087f
C2617 vdd.n930 gnd 0.006087f
C2618 vdd.n931 gnd 0.006087f
C2619 vdd.t217 gnd 0.311039f
C2620 vdd.n932 gnd 0.006087f
C2621 vdd.n933 gnd 0.006087f
C2622 vdd.n934 gnd 0.608355f
C2623 vdd.n935 gnd 0.006087f
C2624 vdd.n936 gnd 0.006087f
C2625 vdd.n937 gnd 0.006087f
C2626 vdd.t177 gnd 0.311039f
C2627 vdd.n938 gnd 0.006087f
C2628 vdd.n939 gnd 0.006087f
C2629 vdd.n940 gnd 0.471132f
C2630 vdd.n941 gnd 0.006087f
C2631 vdd.n942 gnd 0.006087f
C2632 vdd.n943 gnd 0.006087f
C2633 vdd.n944 gnd 0.622078f
C2634 vdd.n945 gnd 0.006087f
C2635 vdd.n946 gnd 0.006087f
C2636 vdd.n947 gnd 0.333909f
C2637 vdd.n948 gnd 0.006087f
C2638 vdd.n949 gnd 0.006087f
C2639 vdd.n950 gnd 0.006087f
C2640 vdd.n951 gnd 0.622078f
C2641 vdd.n952 gnd 0.006087f
C2642 vdd.n953 gnd 0.006087f
C2643 vdd.n954 gnd 0.006087f
C2644 vdd.n955 gnd 0.006087f
C2645 vdd.n956 gnd 0.006087f
C2646 vdd.t15 gnd 0.311039f
C2647 vdd.n957 gnd 0.006087f
C2648 vdd.n958 gnd 0.006087f
C2649 vdd.n959 gnd 0.006087f
C2650 vdd.n960 gnd 0.013034f
C2651 vdd.n961 gnd 0.013034f
C2652 vdd.n962 gnd 0.841635f
C2653 vdd.n963 gnd 0.006087f
C2654 vdd.n964 gnd 0.006087f
C2655 vdd.n965 gnd 0.443688f
C2656 vdd.n966 gnd 0.013034f
C2657 vdd.n967 gnd 0.006087f
C2658 vdd.n968 gnd 0.006087f
C2659 vdd.n969 gnd 11.105901f
C2660 vdd.n1003 gnd 0.013821f
C2661 vdd.n1004 gnd 0.006087f
C2662 vdd.n1005 gnd 0.006087f
C2663 vdd.n1006 gnd 0.005729f
C2664 vdd.n1009 gnd 0.021425f
C2665 vdd.n1010 gnd 0.00598f
C2666 vdd.n1011 gnd 0.007205f
C2667 vdd.n1013 gnd 0.008952f
C2668 vdd.n1014 gnd 0.008952f
C2669 vdd.n1015 gnd 0.007205f
C2670 vdd.n1017 gnd 0.008952f
C2671 vdd.n1018 gnd 0.008952f
C2672 vdd.n1019 gnd 0.008952f
C2673 vdd.n1020 gnd 0.008952f
C2674 vdd.n1021 gnd 0.008952f
C2675 vdd.n1022 gnd 0.007205f
C2676 vdd.n1024 gnd 0.008952f
C2677 vdd.n1025 gnd 0.008952f
C2678 vdd.n1026 gnd 0.008952f
C2679 vdd.n1027 gnd 0.008952f
C2680 vdd.n1028 gnd 0.008952f
C2681 vdd.n1029 gnd 0.007205f
C2682 vdd.n1031 gnd 0.008952f
C2683 vdd.n1032 gnd 0.008952f
C2684 vdd.n1033 gnd 0.008952f
C2685 vdd.n1034 gnd 0.008952f
C2686 vdd.n1035 gnd 0.006016f
C2687 vdd.t24 gnd 0.110129f
C2688 vdd.t23 gnd 0.117698f
C2689 vdd.t22 gnd 0.143827f
C2690 vdd.n1036 gnd 0.184366f
C2691 vdd.n1037 gnd 0.154901f
C2692 vdd.n1039 gnd 0.008952f
C2693 vdd.n1040 gnd 0.008952f
C2694 vdd.n1041 gnd 0.007205f
C2695 vdd.n1042 gnd 0.008952f
C2696 vdd.n1044 gnd 0.008952f
C2697 vdd.n1045 gnd 0.008952f
C2698 vdd.n1046 gnd 0.008952f
C2699 vdd.n1047 gnd 0.008952f
C2700 vdd.n1048 gnd 0.007205f
C2701 vdd.n1050 gnd 0.008952f
C2702 vdd.n1051 gnd 0.008952f
C2703 vdd.n1052 gnd 0.008952f
C2704 vdd.n1053 gnd 0.008952f
C2705 vdd.n1054 gnd 0.008952f
C2706 vdd.n1055 gnd 0.007205f
C2707 vdd.n1057 gnd 0.008952f
C2708 vdd.n1058 gnd 0.008952f
C2709 vdd.n1059 gnd 0.008952f
C2710 vdd.n1060 gnd 0.008952f
C2711 vdd.n1061 gnd 0.008952f
C2712 vdd.n1062 gnd 0.007205f
C2713 vdd.n1064 gnd 0.008952f
C2714 vdd.n1065 gnd 0.008952f
C2715 vdd.n1066 gnd 0.008952f
C2716 vdd.n1067 gnd 0.008952f
C2717 vdd.n1068 gnd 0.008952f
C2718 vdd.n1069 gnd 0.007205f
C2719 vdd.n1071 gnd 0.008952f
C2720 vdd.n1072 gnd 0.008952f
C2721 vdd.n1073 gnd 0.008952f
C2722 vdd.n1074 gnd 0.008952f
C2723 vdd.n1075 gnd 0.007133f
C2724 vdd.t21 gnd 0.110129f
C2725 vdd.t20 gnd 0.117698f
C2726 vdd.t18 gnd 0.143827f
C2727 vdd.n1076 gnd 0.184366f
C2728 vdd.n1077 gnd 0.154901f
C2729 vdd.n1079 gnd 0.008952f
C2730 vdd.n1080 gnd 0.008952f
C2731 vdd.n1081 gnd 0.007205f
C2732 vdd.n1082 gnd 0.008952f
C2733 vdd.n1084 gnd 0.008952f
C2734 vdd.n1085 gnd 0.008952f
C2735 vdd.n1086 gnd 0.008952f
C2736 vdd.n1087 gnd 0.008952f
C2737 vdd.n1088 gnd 0.007205f
C2738 vdd.n1090 gnd 0.008952f
C2739 vdd.n1091 gnd 0.008952f
C2740 vdd.n1092 gnd 0.008952f
C2741 vdd.n1093 gnd 0.008952f
C2742 vdd.n1094 gnd 0.008952f
C2743 vdd.n1095 gnd 0.007205f
C2744 vdd.n1097 gnd 0.008952f
C2745 vdd.n1098 gnd 0.008952f
C2746 vdd.n1099 gnd 0.008952f
C2747 vdd.n1100 gnd 0.008952f
C2748 vdd.n1101 gnd 0.008952f
C2749 vdd.n1102 gnd 0.007205f
C2750 vdd.n1104 gnd 0.008952f
C2751 vdd.n1105 gnd 0.008952f
C2752 vdd.n1106 gnd 0.005729f
C2753 vdd.n1107 gnd 0.007205f
C2754 vdd.n1108 gnd 0.013821f
C2755 vdd.n1109 gnd 0.013821f
C2756 vdd.n1110 gnd 0.006087f
C2757 vdd.n1111 gnd 0.006087f
C2758 vdd.n1112 gnd 0.006087f
C2759 vdd.n1113 gnd 0.006087f
C2760 vdd.n1114 gnd 0.006087f
C2761 vdd.n1115 gnd 0.006087f
C2762 vdd.n1116 gnd 0.006087f
C2763 vdd.n1117 gnd 0.006087f
C2764 vdd.n1118 gnd 0.006087f
C2765 vdd.n1119 gnd 0.006087f
C2766 vdd.n1120 gnd 0.006087f
C2767 vdd.n1121 gnd 0.006087f
C2768 vdd.n1122 gnd 0.006087f
C2769 vdd.n1123 gnd 0.006087f
C2770 vdd.n1124 gnd 0.006087f
C2771 vdd.n1125 gnd 0.006087f
C2772 vdd.n1126 gnd 0.006087f
C2773 vdd.n1127 gnd 0.006087f
C2774 vdd.n1128 gnd 0.006087f
C2775 vdd.n1129 gnd 0.006087f
C2776 vdd.n1130 gnd 0.006087f
C2777 vdd.n1131 gnd 0.006087f
C2778 vdd.n1132 gnd 0.006087f
C2779 vdd.n1133 gnd 0.006087f
C2780 vdd.n1134 gnd 0.006087f
C2781 vdd.n1135 gnd 0.006087f
C2782 vdd.n1136 gnd 0.006087f
C2783 vdd.n1137 gnd 0.006087f
C2784 vdd.n1138 gnd 0.006087f
C2785 vdd.n1139 gnd 0.006087f
C2786 vdd.n1140 gnd 0.006087f
C2787 vdd.n1141 gnd 0.006087f
C2788 vdd.n1142 gnd 0.006087f
C2789 vdd.t16 gnd 0.245981f
C2790 vdd.t17 gnd 0.251792f
C2791 vdd.t14 gnd 0.160586f
C2792 vdd.n1143 gnd 0.086788f
C2793 vdd.n1144 gnd 0.049229f
C2794 vdd.n1145 gnd 0.0087f
C2795 vdd.n1146 gnd 0.006087f
C2796 vdd.t57 gnd 0.245981f
C2797 vdd.t58 gnd 0.251792f
C2798 vdd.t56 gnd 0.160586f
C2799 vdd.n1147 gnd 0.086788f
C2800 vdd.n1148 gnd 0.049229f
C2801 vdd.n1149 gnd 0.006087f
C2802 vdd.n1150 gnd 0.006087f
C2803 vdd.n1151 gnd 0.006087f
C2804 vdd.n1152 gnd 0.006087f
C2805 vdd.n1153 gnd 0.006087f
C2806 vdd.n1154 gnd 0.006087f
C2807 vdd.n1155 gnd 0.006087f
C2808 vdd.n1156 gnd 0.006087f
C2809 vdd.n1157 gnd 0.006087f
C2810 vdd.n1158 gnd 0.006087f
C2811 vdd.n1159 gnd 0.006087f
C2812 vdd.n1160 gnd 0.006087f
C2813 vdd.n1161 gnd 0.006087f
C2814 vdd.n1162 gnd 0.006087f
C2815 vdd.n1163 gnd 0.006087f
C2816 vdd.n1164 gnd 0.006087f
C2817 vdd.n1165 gnd 0.006087f
C2818 vdd.n1166 gnd 0.006087f
C2819 vdd.n1167 gnd 0.006087f
C2820 vdd.n1168 gnd 0.006087f
C2821 vdd.n1169 gnd 0.006087f
C2822 vdd.n1170 gnd 0.006087f
C2823 vdd.n1171 gnd 0.006087f
C2824 vdd.n1172 gnd 0.006087f
C2825 vdd.n1173 gnd 0.006087f
C2826 vdd.n1174 gnd 0.006087f
C2827 vdd.n1175 gnd 0.004431f
C2828 vdd.n1176 gnd 0.0087f
C2829 vdd.n1177 gnd 0.0047f
C2830 vdd.n1178 gnd 0.006087f
C2831 vdd.n1179 gnd 0.006087f
C2832 vdd.n1180 gnd 0.006087f
C2833 vdd.n1181 gnd 0.013821f
C2834 vdd.n1182 gnd 0.013821f
C2835 vdd.n1183 gnd 0.013034f
C2836 vdd.n1184 gnd 0.013034f
C2837 vdd.n1185 gnd 0.006087f
C2838 vdd.n1186 gnd 0.006087f
C2839 vdd.n1187 gnd 0.006087f
C2840 vdd.n1188 gnd 0.006087f
C2841 vdd.n1189 gnd 0.006087f
C2842 vdd.n1190 gnd 0.006087f
C2843 vdd.n1191 gnd 0.006087f
C2844 vdd.n1192 gnd 0.006087f
C2845 vdd.n1193 gnd 0.006087f
C2846 vdd.n1194 gnd 0.006087f
C2847 vdd.n1195 gnd 0.006087f
C2848 vdd.n1196 gnd 0.006087f
C2849 vdd.n1197 gnd 0.006087f
C2850 vdd.n1198 gnd 0.006087f
C2851 vdd.n1199 gnd 0.006087f
C2852 vdd.n1200 gnd 0.006087f
C2853 vdd.n1201 gnd 0.006087f
C2854 vdd.n1202 gnd 0.006087f
C2855 vdd.n1203 gnd 0.006087f
C2856 vdd.n1204 gnd 0.006087f
C2857 vdd.n1205 gnd 0.006087f
C2858 vdd.n1206 gnd 0.006087f
C2859 vdd.n1207 gnd 0.006087f
C2860 vdd.n1208 gnd 0.006087f
C2861 vdd.n1209 gnd 0.006087f
C2862 vdd.n1210 gnd 0.006087f
C2863 vdd.n1211 gnd 0.006087f
C2864 vdd.n1212 gnd 0.006087f
C2865 vdd.n1213 gnd 0.006087f
C2866 vdd.n1214 gnd 0.006087f
C2867 vdd.n1215 gnd 0.006087f
C2868 vdd.n1216 gnd 0.006087f
C2869 vdd.n1217 gnd 0.006087f
C2870 vdd.n1218 gnd 0.006087f
C2871 vdd.n1219 gnd 0.006087f
C2872 vdd.n1220 gnd 0.006087f
C2873 vdd.n1221 gnd 0.006087f
C2874 vdd.n1222 gnd 0.006087f
C2875 vdd.n1223 gnd 0.006087f
C2876 vdd.n1224 gnd 0.006087f
C2877 vdd.n1225 gnd 0.006087f
C2878 vdd.n1226 gnd 0.006087f
C2879 vdd.n1227 gnd 0.370502f
C2880 vdd.n1228 gnd 0.006087f
C2881 vdd.n1229 gnd 0.006087f
C2882 vdd.n1230 gnd 0.006087f
C2883 vdd.n1231 gnd 0.006087f
C2884 vdd.n1232 gnd 0.006087f
C2885 vdd.n1233 gnd 0.006087f
C2886 vdd.n1234 gnd 0.006087f
C2887 vdd.n1235 gnd 0.006087f
C2888 vdd.n1236 gnd 0.006087f
C2889 vdd.n1237 gnd 0.006087f
C2890 vdd.n1238 gnd 0.006087f
C2891 vdd.n1239 gnd 0.006087f
C2892 vdd.n1240 gnd 0.006087f
C2893 vdd.n1241 gnd 0.006087f
C2894 vdd.n1242 gnd 0.006087f
C2895 vdd.n1243 gnd 0.006087f
C2896 vdd.n1244 gnd 0.006087f
C2897 vdd.n1245 gnd 0.006087f
C2898 vdd.n1246 gnd 0.006087f
C2899 vdd.n1247 gnd 0.006087f
C2900 vdd.n1248 gnd 0.006087f
C2901 vdd.n1249 gnd 0.006087f
C2902 vdd.n1250 gnd 0.006087f
C2903 vdd.n1251 gnd 0.006087f
C2904 vdd.n1252 gnd 0.006087f
C2905 vdd.n1253 gnd 0.562614f
C2906 vdd.n1254 gnd 0.006087f
C2907 vdd.n1255 gnd 0.006087f
C2908 vdd.n1256 gnd 0.006087f
C2909 vdd.n1257 gnd 0.006087f
C2910 vdd.n1258 gnd 0.006087f
C2911 vdd.n1259 gnd 0.006087f
C2912 vdd.n1260 gnd 0.006087f
C2913 vdd.n1261 gnd 0.006087f
C2914 vdd.n1262 gnd 0.006087f
C2915 vdd.n1263 gnd 0.006087f
C2916 vdd.n1264 gnd 0.006087f
C2917 vdd.n1265 gnd 0.196686f
C2918 vdd.n1266 gnd 0.006087f
C2919 vdd.n1267 gnd 0.006087f
C2920 vdd.n1268 gnd 0.006087f
C2921 vdd.n1269 gnd 0.006087f
C2922 vdd.n1270 gnd 0.006087f
C2923 vdd.n1271 gnd 0.006087f
C2924 vdd.n1272 gnd 0.006087f
C2925 vdd.n1273 gnd 0.006087f
C2926 vdd.n1274 gnd 0.006087f
C2927 vdd.n1275 gnd 0.006087f
C2928 vdd.n1276 gnd 0.006087f
C2929 vdd.n1277 gnd 0.006087f
C2930 vdd.n1278 gnd 0.006087f
C2931 vdd.n1279 gnd 0.006087f
C2932 vdd.n1280 gnd 0.006087f
C2933 vdd.n1281 gnd 0.006087f
C2934 vdd.n1282 gnd 0.006087f
C2935 vdd.n1283 gnd 0.006087f
C2936 vdd.n1284 gnd 0.006087f
C2937 vdd.n1285 gnd 0.006087f
C2938 vdd.n1286 gnd 0.006087f
C2939 vdd.n1287 gnd 0.006087f
C2940 vdd.n1288 gnd 0.006087f
C2941 vdd.n1289 gnd 0.006087f
C2942 vdd.n1290 gnd 0.006087f
C2943 vdd.n1291 gnd 0.006087f
C2944 vdd.n1292 gnd 0.006087f
C2945 vdd.n1293 gnd 0.006087f
C2946 vdd.n1294 gnd 0.006087f
C2947 vdd.n1295 gnd 0.006087f
C2948 vdd.n1296 gnd 0.006087f
C2949 vdd.n1297 gnd 0.006087f
C2950 vdd.n1298 gnd 0.006087f
C2951 vdd.n1299 gnd 0.006087f
C2952 vdd.n1300 gnd 0.006087f
C2953 vdd.n1301 gnd 0.006087f
C2954 vdd.n1302 gnd 0.006087f
C2955 vdd.n1303 gnd 0.006087f
C2956 vdd.n1304 gnd 0.006087f
C2957 vdd.n1305 gnd 0.006087f
C2958 vdd.n1306 gnd 0.006087f
C2959 vdd.n1307 gnd 0.006087f
C2960 vdd.n1308 gnd 0.013034f
C2961 vdd.n1309 gnd 0.013034f
C2962 vdd.n1310 gnd 0.013821f
C2963 vdd.n1311 gnd 0.006087f
C2964 vdd.n1312 gnd 0.006087f
C2965 vdd.n1313 gnd 0.0047f
C2966 vdd.n1314 gnd 0.006087f
C2967 vdd.n1315 gnd 0.006087f
C2968 vdd.n1316 gnd 0.004431f
C2969 vdd.n1317 gnd 0.006087f
C2970 vdd.n1318 gnd 0.006087f
C2971 vdd.n1319 gnd 0.006087f
C2972 vdd.n1320 gnd 0.006087f
C2973 vdd.n1321 gnd 0.006087f
C2974 vdd.n1322 gnd 0.006087f
C2975 vdd.n1323 gnd 0.006087f
C2976 vdd.n1324 gnd 0.006087f
C2977 vdd.n1325 gnd 0.006087f
C2978 vdd.n1326 gnd 0.006087f
C2979 vdd.n1327 gnd 0.006087f
C2980 vdd.n1328 gnd 0.006087f
C2981 vdd.n1329 gnd 0.006087f
C2982 vdd.n1330 gnd 0.006087f
C2983 vdd.n1331 gnd 0.006087f
C2984 vdd.n1332 gnd 0.006087f
C2985 vdd.n1333 gnd 0.006087f
C2986 vdd.n1334 gnd 0.006087f
C2987 vdd.n1335 gnd 0.006087f
C2988 vdd.n1336 gnd 0.006087f
C2989 vdd.n1337 gnd 0.006087f
C2990 vdd.n1338 gnd 0.006087f
C2991 vdd.n1339 gnd 0.006087f
C2992 vdd.n1340 gnd 0.006087f
C2993 vdd.n1341 gnd 0.006087f
C2994 vdd.n1342 gnd 0.006087f
C2995 vdd.n1343 gnd 0.041006f
C2996 vdd.n1345 gnd 0.021425f
C2997 vdd.n1346 gnd 0.007205f
C2998 vdd.n1348 gnd 0.008952f
C2999 vdd.n1349 gnd 0.007205f
C3000 vdd.n1350 gnd 0.008952f
C3001 vdd.n1352 gnd 0.008952f
C3002 vdd.n1353 gnd 0.008952f
C3003 vdd.n1355 gnd 0.008952f
C3004 vdd.n1356 gnd 0.00598f
C3005 vdd.t19 gnd 0.45741f
C3006 vdd.n1357 gnd 0.008952f
C3007 vdd.n1358 gnd 0.021425f
C3008 vdd.n1359 gnd 0.007205f
C3009 vdd.n1360 gnd 0.008952f
C3010 vdd.n1361 gnd 0.007205f
C3011 vdd.n1362 gnd 0.008952f
C3012 vdd.n1363 gnd 0.91482f
C3013 vdd.n1364 gnd 0.008952f
C3014 vdd.n1365 gnd 0.007205f
C3015 vdd.n1366 gnd 0.007205f
C3016 vdd.n1367 gnd 0.008952f
C3017 vdd.n1368 gnd 0.007205f
C3018 vdd.n1369 gnd 0.008952f
C3019 vdd.t2 gnd 0.45741f
C3020 vdd.n1370 gnd 0.008952f
C3021 vdd.n1371 gnd 0.007205f
C3022 vdd.n1372 gnd 0.008952f
C3023 vdd.n1373 gnd 0.007205f
C3024 vdd.n1374 gnd 0.008952f
C3025 vdd.t143 gnd 0.45741f
C3026 vdd.n1375 gnd 0.008952f
C3027 vdd.n1376 gnd 0.007205f
C3028 vdd.n1377 gnd 0.008952f
C3029 vdd.n1378 gnd 0.007205f
C3030 vdd.n1379 gnd 0.008952f
C3031 vdd.t119 gnd 0.45741f
C3032 vdd.n1380 gnd 0.718134f
C3033 vdd.n1381 gnd 0.008952f
C3034 vdd.n1382 gnd 0.007205f
C3035 vdd.n1383 gnd 0.008952f
C3036 vdd.n1384 gnd 0.007205f
C3037 vdd.n1385 gnd 0.008952f
C3038 vdd.n1386 gnd 0.644948f
C3039 vdd.n1387 gnd 0.008952f
C3040 vdd.n1388 gnd 0.007205f
C3041 vdd.n1389 gnd 0.008952f
C3042 vdd.n1390 gnd 0.007205f
C3043 vdd.n1391 gnd 0.008952f
C3044 vdd.n1392 gnd 0.489429f
C3045 vdd.t92 gnd 0.45741f
C3046 vdd.n1393 gnd 0.008952f
C3047 vdd.n1394 gnd 0.007205f
C3048 vdd.n1395 gnd 0.008921f
C3049 vdd.n1396 gnd 0.007205f
C3050 vdd.n1397 gnd 0.008952f
C3051 vdd.t153 gnd 0.45741f
C3052 vdd.n1398 gnd 0.008952f
C3053 vdd.n1399 gnd 0.007205f
C3054 vdd.n1400 gnd 0.008952f
C3055 vdd.n1401 gnd 0.007205f
C3056 vdd.n1402 gnd 0.008952f
C3057 vdd.t140 gnd 0.45741f
C3058 vdd.n1403 gnd 0.580911f
C3059 vdd.n1404 gnd 0.008952f
C3060 vdd.n1405 gnd 0.007205f
C3061 vdd.n1406 gnd 0.008952f
C3062 vdd.n1407 gnd 0.007205f
C3063 vdd.n1408 gnd 0.008952f
C3064 vdd.t134 gnd 0.45741f
C3065 vdd.n1409 gnd 0.008952f
C3066 vdd.n1410 gnd 0.007205f
C3067 vdd.n1411 gnd 0.008952f
C3068 vdd.n1412 gnd 0.007205f
C3069 vdd.n1413 gnd 0.008952f
C3070 vdd.n1414 gnd 0.626652f
C3071 vdd.n1415 gnd 0.759301f
C3072 vdd.t96 gnd 0.45741f
C3073 vdd.n1416 gnd 0.008952f
C3074 vdd.n1417 gnd 0.007205f
C3075 vdd.n1418 gnd 0.008952f
C3076 vdd.n1419 gnd 0.007205f
C3077 vdd.n1420 gnd 0.008952f
C3078 vdd.n1421 gnd 0.471132f
C3079 vdd.n1422 gnd 0.008952f
C3080 vdd.n1423 gnd 0.007205f
C3081 vdd.n1424 gnd 0.008952f
C3082 vdd.n1425 gnd 0.007205f
C3083 vdd.n1426 gnd 0.008952f
C3084 vdd.n1427 gnd 0.91482f
C3085 vdd.t115 gnd 0.45741f
C3086 vdd.n1428 gnd 0.008952f
C3087 vdd.n1429 gnd 0.007205f
C3088 vdd.n1430 gnd 0.008952f
C3089 vdd.n1431 gnd 0.007205f
C3090 vdd.n1432 gnd 0.008952f
C3091 vdd.t47 gnd 0.45741f
C3092 vdd.n1433 gnd 0.008952f
C3093 vdd.n1434 gnd 0.007205f
C3094 vdd.n1435 gnd 0.021425f
C3095 vdd.n1436 gnd 0.021425f
C3096 vdd.n1437 gnd 2.10409f
C3097 vdd.n1438 gnd 0.516873f
C3098 vdd.n1439 gnd 0.021425f
C3099 vdd.n1440 gnd 0.008952f
C3100 vdd.n1442 gnd 0.008952f
C3101 vdd.n1443 gnd 0.008952f
C3102 vdd.n1444 gnd 0.007205f
C3103 vdd.n1445 gnd 0.008952f
C3104 vdd.n1446 gnd 0.008952f
C3105 vdd.n1448 gnd 0.008952f
C3106 vdd.n1449 gnd 0.008952f
C3107 vdd.n1451 gnd 0.008952f
C3108 vdd.n1452 gnd 0.007205f
C3109 vdd.n1453 gnd 0.008952f
C3110 vdd.n1454 gnd 0.008952f
C3111 vdd.n1456 gnd 0.008952f
C3112 vdd.n1457 gnd 0.008952f
C3113 vdd.n1459 gnd 0.008952f
C3114 vdd.n1460 gnd 0.007205f
C3115 vdd.n1461 gnd 0.008952f
C3116 vdd.n1462 gnd 0.008952f
C3117 vdd.n1464 gnd 0.008952f
C3118 vdd.n1465 gnd 0.008952f
C3119 vdd.n1467 gnd 0.008952f
C3120 vdd.n1468 gnd 0.007205f
C3121 vdd.n1469 gnd 0.008952f
C3122 vdd.n1470 gnd 0.008952f
C3123 vdd.n1472 gnd 0.008952f
C3124 vdd.n1473 gnd 0.008952f
C3125 vdd.n1475 gnd 0.008952f
C3126 vdd.t81 gnd 0.110129f
C3127 vdd.t82 gnd 0.117698f
C3128 vdd.t80 gnd 0.143827f
C3129 vdd.n1476 gnd 0.184366f
C3130 vdd.n1477 gnd 0.155622f
C3131 vdd.n1478 gnd 0.015419f
C3132 vdd.n1479 gnd 0.008952f
C3133 vdd.n1480 gnd 0.008952f
C3134 vdd.n1482 gnd 0.008952f
C3135 vdd.n1483 gnd 0.008952f
C3136 vdd.n1485 gnd 0.008952f
C3137 vdd.n1486 gnd 0.007205f
C3138 vdd.n1487 gnd 0.008952f
C3139 vdd.n1488 gnd 0.008952f
C3140 vdd.n1490 gnd 0.008952f
C3141 vdd.n1491 gnd 0.008952f
C3142 vdd.n1493 gnd 0.008952f
C3143 vdd.n1494 gnd 0.007205f
C3144 vdd.n1495 gnd 0.008952f
C3145 vdd.n1496 gnd 0.008952f
C3146 vdd.n1498 gnd 0.008952f
C3147 vdd.n1499 gnd 0.008952f
C3148 vdd.n1501 gnd 0.008952f
C3149 vdd.n1502 gnd 0.007205f
C3150 vdd.n1503 gnd 0.008952f
C3151 vdd.n1504 gnd 0.008952f
C3152 vdd.n1506 gnd 0.008952f
C3153 vdd.n1507 gnd 0.008952f
C3154 vdd.n1509 gnd 0.008952f
C3155 vdd.n1510 gnd 0.007205f
C3156 vdd.n1511 gnd 0.008952f
C3157 vdd.n1512 gnd 0.008952f
C3158 vdd.n1514 gnd 0.008952f
C3159 vdd.n1515 gnd 0.008952f
C3160 vdd.n1517 gnd 0.008952f
C3161 vdd.n1518 gnd 0.007205f
C3162 vdd.n1519 gnd 0.008952f
C3163 vdd.n1520 gnd 0.008952f
C3164 vdd.n1522 gnd 0.008952f
C3165 vdd.n1523 gnd 0.007133f
C3166 vdd.n1525 gnd 0.007205f
C3167 vdd.n1526 gnd 0.008952f
C3168 vdd.n1527 gnd 0.008952f
C3169 vdd.n1528 gnd 0.008952f
C3170 vdd.n1529 gnd 0.008952f
C3171 vdd.n1531 gnd 0.008952f
C3172 vdd.n1532 gnd 0.008952f
C3173 vdd.n1533 gnd 0.007205f
C3174 vdd.n1534 gnd 0.008952f
C3175 vdd.n1536 gnd 0.008952f
C3176 vdd.n1537 gnd 0.008952f
C3177 vdd.n1539 gnd 0.008952f
C3178 vdd.n1540 gnd 0.008952f
C3179 vdd.n1541 gnd 0.007205f
C3180 vdd.n1542 gnd 0.008952f
C3181 vdd.n1544 gnd 0.008952f
C3182 vdd.n1545 gnd 0.008952f
C3183 vdd.n1547 gnd 0.008952f
C3184 vdd.n1548 gnd 0.008952f
C3185 vdd.n1549 gnd 0.007205f
C3186 vdd.n1550 gnd 0.008952f
C3187 vdd.n1552 gnd 0.008952f
C3188 vdd.n1553 gnd 0.008952f
C3189 vdd.n1555 gnd 0.008952f
C3190 vdd.n1556 gnd 0.008952f
C3191 vdd.n1557 gnd 0.007205f
C3192 vdd.n1558 gnd 0.008952f
C3193 vdd.n1560 gnd 0.008952f
C3194 vdd.n1561 gnd 0.008952f
C3195 vdd.n1563 gnd 0.008952f
C3196 vdd.n1564 gnd 0.003422f
C3197 vdd.t48 gnd 0.110129f
C3198 vdd.t49 gnd 0.117698f
C3199 vdd.t46 gnd 0.143827f
C3200 vdd.n1565 gnd 0.184366f
C3201 vdd.n1566 gnd 0.155622f
C3202 vdd.n1567 gnd 0.011816f
C3203 vdd.n1568 gnd 0.003783f
C3204 vdd.n1569 gnd 0.007205f
C3205 vdd.n1570 gnd 0.008952f
C3206 vdd.n1571 gnd 0.008952f
C3207 vdd.n1572 gnd 0.008952f
C3208 vdd.n1573 gnd 0.007205f
C3209 vdd.n1574 gnd 0.007205f
C3210 vdd.n1575 gnd 0.007205f
C3211 vdd.n1576 gnd 0.008952f
C3212 vdd.n1577 gnd 0.008952f
C3213 vdd.n1578 gnd 0.008952f
C3214 vdd.n1579 gnd 0.007205f
C3215 vdd.n1580 gnd 0.007205f
C3216 vdd.n1581 gnd 0.007205f
C3217 vdd.n1582 gnd 0.008952f
C3218 vdd.n1583 gnd 0.008952f
C3219 vdd.n1584 gnd 0.008952f
C3220 vdd.n1585 gnd 0.007205f
C3221 vdd.n1586 gnd 0.007205f
C3222 vdd.n1587 gnd 0.007205f
C3223 vdd.n1588 gnd 0.008952f
C3224 vdd.n1589 gnd 0.008952f
C3225 vdd.n1590 gnd 0.008952f
C3226 vdd.n1591 gnd 0.007205f
C3227 vdd.n1592 gnd 0.007205f
C3228 vdd.n1593 gnd 0.007205f
C3229 vdd.n1594 gnd 0.008952f
C3230 vdd.n1595 gnd 0.008952f
C3231 vdd.n1596 gnd 0.008952f
C3232 vdd.n1597 gnd 0.007205f
C3233 vdd.n1598 gnd 0.008952f
C3234 vdd.n1599 gnd 0.008952f
C3235 vdd.n1601 gnd 0.008952f
C3236 vdd.t71 gnd 0.110129f
C3237 vdd.t72 gnd 0.117698f
C3238 vdd.t70 gnd 0.143827f
C3239 vdd.n1602 gnd 0.184366f
C3240 vdd.n1603 gnd 0.155622f
C3241 vdd.n1604 gnd 0.015419f
C3242 vdd.n1605 gnd 0.004899f
C3243 vdd.n1606 gnd 0.008952f
C3244 vdd.n1607 gnd 0.008952f
C3245 vdd.n1608 gnd 0.008952f
C3246 vdd.n1609 gnd 0.007205f
C3247 vdd.n1610 gnd 0.007205f
C3248 vdd.n1611 gnd 0.007205f
C3249 vdd.n1612 gnd 0.008952f
C3250 vdd.n1613 gnd 0.008952f
C3251 vdd.n1614 gnd 0.008952f
C3252 vdd.n1615 gnd 0.007205f
C3253 vdd.n1616 gnd 0.007205f
C3254 vdd.n1617 gnd 0.007205f
C3255 vdd.n1618 gnd 0.008952f
C3256 vdd.n1619 gnd 0.008952f
C3257 vdd.n1620 gnd 0.008952f
C3258 vdd.n1621 gnd 0.007205f
C3259 vdd.n1622 gnd 0.007205f
C3260 vdd.n1623 gnd 0.007205f
C3261 vdd.n1624 gnd 0.008952f
C3262 vdd.n1625 gnd 0.008952f
C3263 vdd.n1626 gnd 0.008952f
C3264 vdd.n1627 gnd 0.007205f
C3265 vdd.n1628 gnd 0.007205f
C3266 vdd.n1629 gnd 0.007205f
C3267 vdd.n1630 gnd 0.008952f
C3268 vdd.n1631 gnd 0.008952f
C3269 vdd.n1632 gnd 0.008952f
C3270 vdd.n1633 gnd 0.007205f
C3271 vdd.n1634 gnd 0.007205f
C3272 vdd.n1635 gnd 0.006016f
C3273 vdd.n1636 gnd 0.008952f
C3274 vdd.n1637 gnd 0.008952f
C3275 vdd.n1638 gnd 0.008952f
C3276 vdd.n1639 gnd 0.006016f
C3277 vdd.n1640 gnd 0.007205f
C3278 vdd.n1641 gnd 0.007205f
C3279 vdd.n1642 gnd 0.008952f
C3280 vdd.n1643 gnd 0.008952f
C3281 vdd.n1644 gnd 0.008952f
C3282 vdd.n1645 gnd 0.007205f
C3283 vdd.n1646 gnd 0.007205f
C3284 vdd.n1647 gnd 0.007205f
C3285 vdd.n1648 gnd 0.008952f
C3286 vdd.n1649 gnd 0.008952f
C3287 vdd.n1650 gnd 0.008952f
C3288 vdd.n1651 gnd 0.007205f
C3289 vdd.n1652 gnd 0.007205f
C3290 vdd.n1653 gnd 0.007205f
C3291 vdd.n1654 gnd 0.008952f
C3292 vdd.n1655 gnd 0.008952f
C3293 vdd.n1656 gnd 0.008952f
C3294 vdd.n1657 gnd 0.007205f
C3295 vdd.n1658 gnd 0.007205f
C3296 vdd.n1659 gnd 0.007205f
C3297 vdd.n1660 gnd 0.008952f
C3298 vdd.n1661 gnd 0.008952f
C3299 vdd.n1662 gnd 0.008952f
C3300 vdd.n1663 gnd 0.007205f
C3301 vdd.n1664 gnd 0.007205f
C3302 vdd.n1665 gnd 0.00598f
C3303 vdd.n1666 gnd 0.021425f
C3304 vdd.n1667 gnd 0.021096f
C3305 vdd.n1668 gnd 0.00598f
C3306 vdd.n1669 gnd 0.021096f
C3307 vdd.n1670 gnd 1.2899f
C3308 vdd.n1671 gnd 0.021096f
C3309 vdd.n1672 gnd 0.00598f
C3310 vdd.n1673 gnd 0.021096f
C3311 vdd.n1674 gnd 0.008952f
C3312 vdd.n1675 gnd 0.008952f
C3313 vdd.n1676 gnd 0.007205f
C3314 vdd.n1677 gnd 0.008952f
C3315 vdd.n1678 gnd 0.855357f
C3316 vdd.n1679 gnd 0.008952f
C3317 vdd.n1680 gnd 0.007205f
C3318 vdd.n1681 gnd 0.008952f
C3319 vdd.n1682 gnd 0.008952f
C3320 vdd.n1683 gnd 0.008952f
C3321 vdd.n1684 gnd 0.007205f
C3322 vdd.n1685 gnd 0.008952f
C3323 vdd.n1686 gnd 0.901098f
C3324 vdd.n1687 gnd 0.008952f
C3325 vdd.n1688 gnd 0.007205f
C3326 vdd.n1689 gnd 0.008952f
C3327 vdd.n1690 gnd 0.008952f
C3328 vdd.n1691 gnd 0.008952f
C3329 vdd.n1692 gnd 0.007205f
C3330 vdd.n1693 gnd 0.008952f
C3331 vdd.t149 gnd 0.45741f
C3332 vdd.n1694 gnd 0.745578f
C3333 vdd.n1695 gnd 0.008952f
C3334 vdd.n1696 gnd 0.007205f
C3335 vdd.n1697 gnd 0.008952f
C3336 vdd.n1698 gnd 0.008952f
C3337 vdd.n1699 gnd 0.008952f
C3338 vdd.n1700 gnd 0.007205f
C3339 vdd.n1701 gnd 0.008952f
C3340 vdd.n1702 gnd 0.590059f
C3341 vdd.n1703 gnd 0.008952f
C3342 vdd.n1704 gnd 0.007205f
C3343 vdd.n1705 gnd 0.008952f
C3344 vdd.n1706 gnd 0.008952f
C3345 vdd.n1707 gnd 0.008952f
C3346 vdd.n1708 gnd 0.007205f
C3347 vdd.n1709 gnd 0.008952f
C3348 vdd.n1710 gnd 0.73643f
C3349 vdd.n1711 gnd 0.480281f
C3350 vdd.n1712 gnd 0.008952f
C3351 vdd.n1713 gnd 0.007205f
C3352 vdd.n1714 gnd 0.008952f
C3353 vdd.n1715 gnd 0.008952f
C3354 vdd.n1716 gnd 0.008952f
C3355 vdd.n1717 gnd 0.007205f
C3356 vdd.n1718 gnd 0.008952f
C3357 vdd.n1719 gnd 0.6358f
C3358 vdd.n1720 gnd 0.008952f
C3359 vdd.n1721 gnd 0.007205f
C3360 vdd.n1722 gnd 0.008952f
C3361 vdd.n1723 gnd 0.008952f
C3362 vdd.n1724 gnd 0.008952f
C3363 vdd.n1725 gnd 0.007205f
C3364 vdd.n1726 gnd 0.008952f
C3365 vdd.t90 gnd 0.45741f
C3366 vdd.n1727 gnd 0.759301f
C3367 vdd.n1728 gnd 0.008952f
C3368 vdd.n1729 gnd 0.007205f
C3369 vdd.n1730 gnd 0.004913f
C3370 vdd.n1731 gnd 0.004559f
C3371 vdd.n1732 gnd 0.002522f
C3372 vdd.n1733 gnd 0.00579f
C3373 vdd.n1734 gnd 0.00245f
C3374 vdd.n1735 gnd 0.002594f
C3375 vdd.n1736 gnd 0.004559f
C3376 vdd.n1737 gnd 0.00245f
C3377 vdd.n1738 gnd 0.00579f
C3378 vdd.n1739 gnd 0.002594f
C3379 vdd.n1740 gnd 0.004559f
C3380 vdd.n1741 gnd 0.00245f
C3381 vdd.n1742 gnd 0.004343f
C3382 vdd.n1743 gnd 0.004356f
C3383 vdd.t3 gnd 0.01244f
C3384 vdd.n1744 gnd 0.027678f
C3385 vdd.n1745 gnd 0.144045f
C3386 vdd.n1746 gnd 0.00245f
C3387 vdd.n1747 gnd 0.002594f
C3388 vdd.n1748 gnd 0.00579f
C3389 vdd.n1749 gnd 0.00579f
C3390 vdd.n1750 gnd 0.002594f
C3391 vdd.n1751 gnd 0.00245f
C3392 vdd.n1752 gnd 0.004559f
C3393 vdd.n1753 gnd 0.004559f
C3394 vdd.n1754 gnd 0.00245f
C3395 vdd.n1755 gnd 0.002594f
C3396 vdd.n1756 gnd 0.00579f
C3397 vdd.n1757 gnd 0.00579f
C3398 vdd.n1758 gnd 0.002594f
C3399 vdd.n1759 gnd 0.00245f
C3400 vdd.n1760 gnd 0.004559f
C3401 vdd.n1761 gnd 0.004559f
C3402 vdd.n1762 gnd 0.00245f
C3403 vdd.n1763 gnd 0.002594f
C3404 vdd.n1764 gnd 0.00579f
C3405 vdd.n1765 gnd 0.00579f
C3406 vdd.n1766 gnd 0.013689f
C3407 vdd.n1767 gnd 0.002522f
C3408 vdd.n1768 gnd 0.00245f
C3409 vdd.n1769 gnd 0.011783f
C3410 vdd.n1770 gnd 0.008226f
C3411 vdd.t120 gnd 0.02882f
C3412 vdd.t144 gnd 0.02882f
C3413 vdd.n1771 gnd 0.198072f
C3414 vdd.n1772 gnd 0.155753f
C3415 vdd.t159 gnd 0.02882f
C3416 vdd.t155 gnd 0.02882f
C3417 vdd.n1773 gnd 0.198072f
C3418 vdd.n1774 gnd 0.125692f
C3419 vdd.t166 gnd 0.02882f
C3420 vdd.t91 gnd 0.02882f
C3421 vdd.n1775 gnd 0.198072f
C3422 vdd.n1776 gnd 0.125692f
C3423 vdd.t135 gnd 0.02882f
C3424 vdd.t239 gnd 0.02882f
C3425 vdd.n1777 gnd 0.198072f
C3426 vdd.n1778 gnd 0.125692f
C3427 vdd.t150 gnd 0.02882f
C3428 vdd.t152 gnd 0.02882f
C3429 vdd.n1779 gnd 0.198072f
C3430 vdd.n1780 gnd 0.125692f
C3431 vdd.n1781 gnd 0.004913f
C3432 vdd.n1782 gnd 0.004559f
C3433 vdd.n1783 gnd 0.002522f
C3434 vdd.n1784 gnd 0.00579f
C3435 vdd.n1785 gnd 0.00245f
C3436 vdd.n1786 gnd 0.002594f
C3437 vdd.n1787 gnd 0.004559f
C3438 vdd.n1788 gnd 0.00245f
C3439 vdd.n1789 gnd 0.00579f
C3440 vdd.n1790 gnd 0.002594f
C3441 vdd.n1791 gnd 0.004559f
C3442 vdd.n1792 gnd 0.00245f
C3443 vdd.n1793 gnd 0.004343f
C3444 vdd.n1794 gnd 0.004356f
C3445 vdd.t123 gnd 0.01244f
C3446 vdd.n1795 gnd 0.027678f
C3447 vdd.n1796 gnd 0.144045f
C3448 vdd.n1797 gnd 0.00245f
C3449 vdd.n1798 gnd 0.002594f
C3450 vdd.n1799 gnd 0.00579f
C3451 vdd.n1800 gnd 0.00579f
C3452 vdd.n1801 gnd 0.002594f
C3453 vdd.n1802 gnd 0.00245f
C3454 vdd.n1803 gnd 0.004559f
C3455 vdd.n1804 gnd 0.004559f
C3456 vdd.n1805 gnd 0.00245f
C3457 vdd.n1806 gnd 0.002594f
C3458 vdd.n1807 gnd 0.00579f
C3459 vdd.n1808 gnd 0.00579f
C3460 vdd.n1809 gnd 0.002594f
C3461 vdd.n1810 gnd 0.00245f
C3462 vdd.n1811 gnd 0.004559f
C3463 vdd.n1812 gnd 0.004559f
C3464 vdd.n1813 gnd 0.00245f
C3465 vdd.n1814 gnd 0.002594f
C3466 vdd.n1815 gnd 0.00579f
C3467 vdd.n1816 gnd 0.00579f
C3468 vdd.n1817 gnd 0.013689f
C3469 vdd.n1818 gnd 0.002522f
C3470 vdd.n1819 gnd 0.00245f
C3471 vdd.n1820 gnd 0.011783f
C3472 vdd.n1821 gnd 0.007968f
C3473 vdd.n1822 gnd 0.093515f
C3474 vdd.n1823 gnd 0.004913f
C3475 vdd.n1824 gnd 0.004559f
C3476 vdd.n1825 gnd 0.002522f
C3477 vdd.n1826 gnd 0.00579f
C3478 vdd.n1827 gnd 0.00245f
C3479 vdd.n1828 gnd 0.002594f
C3480 vdd.n1829 gnd 0.004559f
C3481 vdd.n1830 gnd 0.00245f
C3482 vdd.n1831 gnd 0.00579f
C3483 vdd.n1832 gnd 0.002594f
C3484 vdd.n1833 gnd 0.004559f
C3485 vdd.n1834 gnd 0.00245f
C3486 vdd.n1835 gnd 0.004343f
C3487 vdd.n1836 gnd 0.004356f
C3488 vdd.t133 gnd 0.01244f
C3489 vdd.n1837 gnd 0.027678f
C3490 vdd.n1838 gnd 0.144045f
C3491 vdd.n1839 gnd 0.00245f
C3492 vdd.n1840 gnd 0.002594f
C3493 vdd.n1841 gnd 0.00579f
C3494 vdd.n1842 gnd 0.00579f
C3495 vdd.n1843 gnd 0.002594f
C3496 vdd.n1844 gnd 0.00245f
C3497 vdd.n1845 gnd 0.004559f
C3498 vdd.n1846 gnd 0.004559f
C3499 vdd.n1847 gnd 0.00245f
C3500 vdd.n1848 gnd 0.002594f
C3501 vdd.n1849 gnd 0.00579f
C3502 vdd.n1850 gnd 0.00579f
C3503 vdd.n1851 gnd 0.002594f
C3504 vdd.n1852 gnd 0.00245f
C3505 vdd.n1853 gnd 0.004559f
C3506 vdd.n1854 gnd 0.004559f
C3507 vdd.n1855 gnd 0.00245f
C3508 vdd.n1856 gnd 0.002594f
C3509 vdd.n1857 gnd 0.00579f
C3510 vdd.n1858 gnd 0.00579f
C3511 vdd.n1859 gnd 0.013689f
C3512 vdd.n1860 gnd 0.002522f
C3513 vdd.n1861 gnd 0.00245f
C3514 vdd.n1862 gnd 0.011783f
C3515 vdd.n1863 gnd 0.008226f
C3516 vdd.t167 gnd 0.02882f
C3517 vdd.t151 gnd 0.02882f
C3518 vdd.n1864 gnd 0.198072f
C3519 vdd.n1865 gnd 0.155753f
C3520 vdd.t93 gnd 0.02882f
C3521 vdd.t1 gnd 0.02882f
C3522 vdd.n1866 gnd 0.198072f
C3523 vdd.n1867 gnd 0.125692f
C3524 vdd.t158 gnd 0.02882f
C3525 vdd.t100 gnd 0.02882f
C3526 vdd.n1868 gnd 0.198072f
C3527 vdd.n1869 gnd 0.125692f
C3528 vdd.t235 gnd 0.02882f
C3529 vdd.t157 gnd 0.02882f
C3530 vdd.n1870 gnd 0.198072f
C3531 vdd.n1871 gnd 0.125692f
C3532 vdd.t169 gnd 0.02882f
C3533 vdd.t233 gnd 0.02882f
C3534 vdd.n1872 gnd 0.198072f
C3535 vdd.n1873 gnd 0.125692f
C3536 vdd.n1874 gnd 0.004913f
C3537 vdd.n1875 gnd 0.004559f
C3538 vdd.n1876 gnd 0.002522f
C3539 vdd.n1877 gnd 0.00579f
C3540 vdd.n1878 gnd 0.00245f
C3541 vdd.n1879 gnd 0.002594f
C3542 vdd.n1880 gnd 0.004559f
C3543 vdd.n1881 gnd 0.00245f
C3544 vdd.n1882 gnd 0.00579f
C3545 vdd.n1883 gnd 0.002594f
C3546 vdd.n1884 gnd 0.004559f
C3547 vdd.n1885 gnd 0.00245f
C3548 vdd.n1886 gnd 0.004343f
C3549 vdd.n1887 gnd 0.004356f
C3550 vdd.t116 gnd 0.01244f
C3551 vdd.n1888 gnd 0.027678f
C3552 vdd.n1889 gnd 0.144045f
C3553 vdd.n1890 gnd 0.00245f
C3554 vdd.n1891 gnd 0.002594f
C3555 vdd.n1892 gnd 0.00579f
C3556 vdd.n1893 gnd 0.00579f
C3557 vdd.n1894 gnd 0.002594f
C3558 vdd.n1895 gnd 0.00245f
C3559 vdd.n1896 gnd 0.004559f
C3560 vdd.n1897 gnd 0.004559f
C3561 vdd.n1898 gnd 0.00245f
C3562 vdd.n1899 gnd 0.002594f
C3563 vdd.n1900 gnd 0.00579f
C3564 vdd.n1901 gnd 0.00579f
C3565 vdd.n1902 gnd 0.002594f
C3566 vdd.n1903 gnd 0.00245f
C3567 vdd.n1904 gnd 0.004559f
C3568 vdd.n1905 gnd 0.004559f
C3569 vdd.n1906 gnd 0.00245f
C3570 vdd.n1907 gnd 0.002594f
C3571 vdd.n1908 gnd 0.00579f
C3572 vdd.n1909 gnd 0.00579f
C3573 vdd.n1910 gnd 0.013689f
C3574 vdd.n1911 gnd 0.002522f
C3575 vdd.n1912 gnd 0.00245f
C3576 vdd.n1913 gnd 0.011783f
C3577 vdd.n1914 gnd 0.007968f
C3578 vdd.n1915 gnd 0.055632f
C3579 vdd.n1916 gnd 0.200457f
C3580 vdd.n1917 gnd 0.004913f
C3581 vdd.n1918 gnd 0.004559f
C3582 vdd.n1919 gnd 0.002522f
C3583 vdd.n1920 gnd 0.00579f
C3584 vdd.n1921 gnd 0.00245f
C3585 vdd.n1922 gnd 0.002594f
C3586 vdd.n1923 gnd 0.004559f
C3587 vdd.n1924 gnd 0.00245f
C3588 vdd.n1925 gnd 0.00579f
C3589 vdd.n1926 gnd 0.002594f
C3590 vdd.n1927 gnd 0.004559f
C3591 vdd.n1928 gnd 0.00245f
C3592 vdd.n1929 gnd 0.004343f
C3593 vdd.n1930 gnd 0.004356f
C3594 vdd.t234 gnd 0.01244f
C3595 vdd.n1931 gnd 0.027678f
C3596 vdd.n1932 gnd 0.144045f
C3597 vdd.n1933 gnd 0.00245f
C3598 vdd.n1934 gnd 0.002594f
C3599 vdd.n1935 gnd 0.00579f
C3600 vdd.n1936 gnd 0.00579f
C3601 vdd.n1937 gnd 0.002594f
C3602 vdd.n1938 gnd 0.00245f
C3603 vdd.n1939 gnd 0.004559f
C3604 vdd.n1940 gnd 0.004559f
C3605 vdd.n1941 gnd 0.00245f
C3606 vdd.n1942 gnd 0.002594f
C3607 vdd.n1943 gnd 0.00579f
C3608 vdd.n1944 gnd 0.00579f
C3609 vdd.n1945 gnd 0.002594f
C3610 vdd.n1946 gnd 0.00245f
C3611 vdd.n1947 gnd 0.004559f
C3612 vdd.n1948 gnd 0.004559f
C3613 vdd.n1949 gnd 0.00245f
C3614 vdd.n1950 gnd 0.002594f
C3615 vdd.n1951 gnd 0.00579f
C3616 vdd.n1952 gnd 0.00579f
C3617 vdd.n1953 gnd 0.013689f
C3618 vdd.n1954 gnd 0.002522f
C3619 vdd.n1955 gnd 0.00245f
C3620 vdd.n1956 gnd 0.011783f
C3621 vdd.n1957 gnd 0.008226f
C3622 vdd.t164 gnd 0.02882f
C3623 vdd.t165 gnd 0.02882f
C3624 vdd.n1958 gnd 0.198072f
C3625 vdd.n1959 gnd 0.155753f
C3626 vdd.t137 gnd 0.02882f
C3627 vdd.t139 gnd 0.02882f
C3628 vdd.n1960 gnd 0.198072f
C3629 vdd.n1961 gnd 0.125692f
C3630 vdd.t154 gnd 0.02882f
C3631 vdd.t161 gnd 0.02882f
C3632 vdd.n1962 gnd 0.198072f
C3633 vdd.n1963 gnd 0.125692f
C3634 vdd.t229 gnd 0.02882f
C3635 vdd.t141 gnd 0.02882f
C3636 vdd.n1964 gnd 0.198072f
C3637 vdd.n1965 gnd 0.125692f
C3638 vdd.t236 gnd 0.02882f
C3639 vdd.t97 gnd 0.02882f
C3640 vdd.n1966 gnd 0.198072f
C3641 vdd.n1967 gnd 0.125692f
C3642 vdd.n1968 gnd 0.004913f
C3643 vdd.n1969 gnd 0.004559f
C3644 vdd.n1970 gnd 0.002522f
C3645 vdd.n1971 gnd 0.00579f
C3646 vdd.n1972 gnd 0.00245f
C3647 vdd.n1973 gnd 0.002594f
C3648 vdd.n1974 gnd 0.004559f
C3649 vdd.n1975 gnd 0.00245f
C3650 vdd.n1976 gnd 0.00579f
C3651 vdd.n1977 gnd 0.002594f
C3652 vdd.n1978 gnd 0.004559f
C3653 vdd.n1979 gnd 0.00245f
C3654 vdd.n1980 gnd 0.004343f
C3655 vdd.n1981 gnd 0.004356f
C3656 vdd.t147 gnd 0.01244f
C3657 vdd.n1982 gnd 0.027678f
C3658 vdd.n1983 gnd 0.144045f
C3659 vdd.n1984 gnd 0.00245f
C3660 vdd.n1985 gnd 0.002594f
C3661 vdd.n1986 gnd 0.00579f
C3662 vdd.n1987 gnd 0.00579f
C3663 vdd.n1988 gnd 0.002594f
C3664 vdd.n1989 gnd 0.00245f
C3665 vdd.n1990 gnd 0.004559f
C3666 vdd.n1991 gnd 0.004559f
C3667 vdd.n1992 gnd 0.00245f
C3668 vdd.n1993 gnd 0.002594f
C3669 vdd.n1994 gnd 0.00579f
C3670 vdd.n1995 gnd 0.00579f
C3671 vdd.n1996 gnd 0.002594f
C3672 vdd.n1997 gnd 0.00245f
C3673 vdd.n1998 gnd 0.004559f
C3674 vdd.n1999 gnd 0.004559f
C3675 vdd.n2000 gnd 0.00245f
C3676 vdd.n2001 gnd 0.002594f
C3677 vdd.n2002 gnd 0.00579f
C3678 vdd.n2003 gnd 0.00579f
C3679 vdd.n2004 gnd 0.013689f
C3680 vdd.n2005 gnd 0.002522f
C3681 vdd.n2006 gnd 0.00245f
C3682 vdd.n2007 gnd 0.011783f
C3683 vdd.n2008 gnd 0.007968f
C3684 vdd.n2009 gnd 0.055632f
C3685 vdd.n2010 gnd 0.220309f
C3686 vdd.n2011 gnd 2.30733f
C3687 vdd.n2012 gnd 0.532874f
C3688 vdd.n2013 gnd 0.008921f
C3689 vdd.n2014 gnd 0.008952f
C3690 vdd.n2015 gnd 0.007205f
C3691 vdd.n2016 gnd 0.008952f
C3692 vdd.n2017 gnd 0.727282f
C3693 vdd.n2018 gnd 0.008952f
C3694 vdd.n2019 gnd 0.007205f
C3695 vdd.n2020 gnd 0.008952f
C3696 vdd.n2021 gnd 0.008952f
C3697 vdd.n2022 gnd 0.008952f
C3698 vdd.n2023 gnd 0.007205f
C3699 vdd.n2024 gnd 0.008952f
C3700 vdd.n2025 gnd 0.759301f
C3701 vdd.t0 gnd 0.45741f
C3702 vdd.n2026 gnd 0.571763f
C3703 vdd.n2027 gnd 0.008952f
C3704 vdd.n2028 gnd 0.007205f
C3705 vdd.n2029 gnd 0.008952f
C3706 vdd.n2030 gnd 0.008952f
C3707 vdd.n2031 gnd 0.008952f
C3708 vdd.n2032 gnd 0.007205f
C3709 vdd.n2033 gnd 0.008952f
C3710 vdd.n2034 gnd 0.498577f
C3711 vdd.n2035 gnd 0.008952f
C3712 vdd.n2036 gnd 0.007205f
C3713 vdd.n2037 gnd 0.008952f
C3714 vdd.n2038 gnd 0.008952f
C3715 vdd.n2039 gnd 0.008952f
C3716 vdd.n2040 gnd 0.007205f
C3717 vdd.n2041 gnd 0.008952f
C3718 vdd.n2042 gnd 0.562614f
C3719 vdd.n2043 gnd 0.654096f
C3720 vdd.n2044 gnd 0.008952f
C3721 vdd.n2045 gnd 0.007205f
C3722 vdd.n2046 gnd 0.008952f
C3723 vdd.n2047 gnd 0.008952f
C3724 vdd.n2048 gnd 0.008952f
C3725 vdd.n2049 gnd 0.007205f
C3726 vdd.n2050 gnd 0.008952f
C3727 vdd.n2051 gnd 0.809616f
C3728 vdd.n2052 gnd 0.008952f
C3729 vdd.n2053 gnd 0.007205f
C3730 vdd.n2054 gnd 0.008952f
C3731 vdd.n2055 gnd 0.008952f
C3732 vdd.n2056 gnd 0.021096f
C3733 vdd.n2057 gnd 0.008952f
C3734 vdd.n2058 gnd 0.008952f
C3735 vdd.n2059 gnd 0.007205f
C3736 vdd.n2060 gnd 0.008952f
C3737 vdd.n2061 gnd 0.489429f
C3738 vdd.n2062 gnd 0.91482f
C3739 vdd.n2063 gnd 0.008952f
C3740 vdd.n2064 gnd 0.007205f
C3741 vdd.n2065 gnd 0.008952f
C3742 vdd.n2066 gnd 0.008952f
C3743 vdd.n2067 gnd 0.021096f
C3744 vdd.n2068 gnd 0.00598f
C3745 vdd.n2069 gnd 0.021096f
C3746 vdd.n2070 gnd 1.25788f
C3747 vdd.n2071 gnd 0.021096f
C3748 vdd.n2072 gnd 0.021425f
C3749 vdd.n2073 gnd 0.003422f
C3750 vdd.t42 gnd 0.110129f
C3751 vdd.t41 gnd 0.117698f
C3752 vdd.t40 gnd 0.143827f
C3753 vdd.n2074 gnd 0.184366f
C3754 vdd.n2075 gnd 0.154901f
C3755 vdd.n2076 gnd 0.011096f
C3756 vdd.n2077 gnd 0.003783f
C3757 vdd.n2078 gnd 0.007698f
C3758 vdd.n2079 gnd 0.950314f
C3759 vdd.n2081 gnd 0.007205f
C3760 vdd.n2082 gnd 0.007205f
C3761 vdd.n2083 gnd 0.008952f
C3762 vdd.n2085 gnd 0.008952f
C3763 vdd.n2086 gnd 0.008952f
C3764 vdd.n2087 gnd 0.007205f
C3765 vdd.n2088 gnd 0.007205f
C3766 vdd.n2089 gnd 0.007205f
C3767 vdd.n2090 gnd 0.008952f
C3768 vdd.n2092 gnd 0.008952f
C3769 vdd.n2093 gnd 0.008952f
C3770 vdd.n2094 gnd 0.007205f
C3771 vdd.n2095 gnd 0.007205f
C3772 vdd.n2096 gnd 0.007205f
C3773 vdd.n2097 gnd 0.008952f
C3774 vdd.n2099 gnd 0.008952f
C3775 vdd.n2100 gnd 0.008952f
C3776 vdd.n2101 gnd 0.007205f
C3777 vdd.n2102 gnd 0.007205f
C3778 vdd.n2103 gnd 0.007205f
C3779 vdd.n2104 gnd 0.008952f
C3780 vdd.n2106 gnd 0.008952f
C3781 vdd.n2107 gnd 0.008952f
C3782 vdd.n2108 gnd 0.007205f
C3783 vdd.n2109 gnd 0.008952f
C3784 vdd.n2110 gnd 0.008952f
C3785 vdd.n2111 gnd 0.008952f
C3786 vdd.n2112 gnd 0.014698f
C3787 vdd.n2113 gnd 0.004899f
C3788 vdd.n2114 gnd 0.007205f
C3789 vdd.n2115 gnd 0.008952f
C3790 vdd.n2117 gnd 0.008952f
C3791 vdd.n2118 gnd 0.008952f
C3792 vdd.n2119 gnd 0.007205f
C3793 vdd.n2120 gnd 0.007205f
C3794 vdd.n2121 gnd 0.007205f
C3795 vdd.n2122 gnd 0.008952f
C3796 vdd.n2124 gnd 0.008952f
C3797 vdd.n2125 gnd 0.008952f
C3798 vdd.n2126 gnd 0.007205f
C3799 vdd.n2127 gnd 0.007205f
C3800 vdd.n2128 gnd 0.007205f
C3801 vdd.n2129 gnd 0.008952f
C3802 vdd.n2131 gnd 0.008952f
C3803 vdd.n2132 gnd 0.008952f
C3804 vdd.n2133 gnd 0.007205f
C3805 vdd.n2134 gnd 0.007205f
C3806 vdd.n2135 gnd 0.007205f
C3807 vdd.n2136 gnd 0.008952f
C3808 vdd.n2138 gnd 0.008952f
C3809 vdd.n2139 gnd 0.008952f
C3810 vdd.n2140 gnd 0.007205f
C3811 vdd.n2141 gnd 0.007205f
C3812 vdd.n2142 gnd 0.007205f
C3813 vdd.n2143 gnd 0.008952f
C3814 vdd.n2145 gnd 0.008952f
C3815 vdd.n2146 gnd 0.008952f
C3816 vdd.n2147 gnd 0.007205f
C3817 vdd.n2148 gnd 0.008952f
C3818 vdd.n2149 gnd 0.008952f
C3819 vdd.n2150 gnd 0.008952f
C3820 vdd.n2151 gnd 0.014698f
C3821 vdd.n2152 gnd 0.006016f
C3822 vdd.n2153 gnd 0.007205f
C3823 vdd.n2154 gnd 0.008952f
C3824 vdd.n2156 gnd 0.008952f
C3825 vdd.n2157 gnd 0.008952f
C3826 vdd.n2158 gnd 0.007205f
C3827 vdd.n2159 gnd 0.007205f
C3828 vdd.n2160 gnd 0.007205f
C3829 vdd.n2161 gnd 0.008952f
C3830 vdd.n2163 gnd 0.008952f
C3831 vdd.n2164 gnd 0.008952f
C3832 vdd.n2165 gnd 0.007205f
C3833 vdd.n2166 gnd 0.007205f
C3834 vdd.n2167 gnd 0.007205f
C3835 vdd.n2168 gnd 0.008952f
C3836 vdd.n2170 gnd 0.008952f
C3837 vdd.n2171 gnd 0.008952f
C3838 vdd.n2172 gnd 0.007205f
C3839 vdd.n2173 gnd 0.007205f
C3840 vdd.n2174 gnd 0.007205f
C3841 vdd.n2175 gnd 0.008952f
C3842 vdd.n2177 gnd 0.008952f
C3843 vdd.n2178 gnd 0.007205f
C3844 vdd.n2179 gnd 0.007205f
C3845 vdd.n2180 gnd 0.008952f
C3846 vdd.n2182 gnd 0.008952f
C3847 vdd.n2183 gnd 0.008952f
C3848 vdd.n2184 gnd 0.007205f
C3849 vdd.n2185 gnd 0.007698f
C3850 vdd.n2186 gnd 0.950314f
C3851 vdd.n2187 gnd 0.041006f
C3852 vdd.n2188 gnd 0.006087f
C3853 vdd.n2189 gnd 0.006087f
C3854 vdd.n2190 gnd 0.006087f
C3855 vdd.n2191 gnd 0.006087f
C3856 vdd.n2192 gnd 0.006087f
C3857 vdd.n2193 gnd 0.006087f
C3858 vdd.n2194 gnd 0.006087f
C3859 vdd.n2195 gnd 0.006087f
C3860 vdd.n2196 gnd 0.006087f
C3861 vdd.n2197 gnd 0.006087f
C3862 vdd.n2198 gnd 0.006087f
C3863 vdd.n2199 gnd 0.006087f
C3864 vdd.n2200 gnd 0.006087f
C3865 vdd.n2201 gnd 0.006087f
C3866 vdd.n2202 gnd 0.006087f
C3867 vdd.n2203 gnd 0.006087f
C3868 vdd.n2204 gnd 0.006087f
C3869 vdd.n2205 gnd 0.006087f
C3870 vdd.n2206 gnd 0.006087f
C3871 vdd.n2207 gnd 0.006087f
C3872 vdd.n2208 gnd 0.006087f
C3873 vdd.n2209 gnd 0.006087f
C3874 vdd.n2210 gnd 0.006087f
C3875 vdd.n2211 gnd 0.006087f
C3876 vdd.n2212 gnd 0.006087f
C3877 vdd.n2213 gnd 0.006087f
C3878 vdd.n2214 gnd 0.006087f
C3879 vdd.n2215 gnd 0.006087f
C3880 vdd.n2216 gnd 0.006087f
C3881 vdd.n2217 gnd 0.006087f
C3882 vdd.n2218 gnd 10.804f
C3883 vdd.n2220 gnd 0.013821f
C3884 vdd.n2221 gnd 0.013821f
C3885 vdd.n2222 gnd 0.013034f
C3886 vdd.n2223 gnd 0.006087f
C3887 vdd.n2224 gnd 0.006087f
C3888 vdd.n2225 gnd 0.622078f
C3889 vdd.n2226 gnd 0.006087f
C3890 vdd.n2227 gnd 0.006087f
C3891 vdd.n2228 gnd 0.006087f
C3892 vdd.n2229 gnd 0.006087f
C3893 vdd.n2230 gnd 0.006087f
C3894 vdd.n2231 gnd 0.489429f
C3895 vdd.n2232 gnd 0.006087f
C3896 vdd.n2233 gnd 0.006087f
C3897 vdd.n2234 gnd 0.006087f
C3898 vdd.n2235 gnd 0.006087f
C3899 vdd.n2236 gnd 0.006087f
C3900 vdd.n2237 gnd 0.622078f
C3901 vdd.n2238 gnd 0.006087f
C3902 vdd.n2239 gnd 0.006087f
C3903 vdd.n2240 gnd 0.006087f
C3904 vdd.n2241 gnd 0.006087f
C3905 vdd.n2242 gnd 0.006087f
C3906 vdd.n2243 gnd 0.622078f
C3907 vdd.n2244 gnd 0.006087f
C3908 vdd.n2245 gnd 0.006087f
C3909 vdd.n2246 gnd 0.006087f
C3910 vdd.n2247 gnd 0.006087f
C3911 vdd.n2248 gnd 0.006087f
C3912 vdd.n2249 gnd 0.599207f
C3913 vdd.n2250 gnd 0.006087f
C3914 vdd.n2251 gnd 0.006087f
C3915 vdd.n2252 gnd 0.006087f
C3916 vdd.n2253 gnd 0.006087f
C3917 vdd.n2254 gnd 0.006087f
C3918 vdd.n2255 gnd 0.461984f
C3919 vdd.n2256 gnd 0.006087f
C3920 vdd.n2257 gnd 0.006087f
C3921 vdd.n2258 gnd 0.006087f
C3922 vdd.n2259 gnd 0.006087f
C3923 vdd.n2260 gnd 0.006087f
C3924 vdd.n2261 gnd 0.324761f
C3925 vdd.n2262 gnd 0.006087f
C3926 vdd.n2263 gnd 0.006087f
C3927 vdd.n2264 gnd 0.006087f
C3928 vdd.n2265 gnd 0.006087f
C3929 vdd.n2266 gnd 0.006087f
C3930 vdd.n2267 gnd 0.43454f
C3931 vdd.n2268 gnd 0.006087f
C3932 vdd.n2269 gnd 0.006087f
C3933 vdd.n2270 gnd 0.006087f
C3934 vdd.n2271 gnd 0.006087f
C3935 vdd.n2272 gnd 0.006087f
C3936 vdd.n2273 gnd 0.571763f
C3937 vdd.n2274 gnd 0.006087f
C3938 vdd.n2275 gnd 0.006087f
C3939 vdd.n2276 gnd 0.006087f
C3940 vdd.n2277 gnd 0.006087f
C3941 vdd.n2278 gnd 0.006087f
C3942 vdd.n2279 gnd 0.622078f
C3943 vdd.n2280 gnd 0.006087f
C3944 vdd.n2281 gnd 0.006087f
C3945 vdd.n2282 gnd 0.006087f
C3946 vdd.n2283 gnd 0.006087f
C3947 vdd.n2284 gnd 0.006087f
C3948 vdd.n2285 gnd 0.53517f
C3949 vdd.n2286 gnd 0.006087f
C3950 vdd.n2287 gnd 0.006087f
C3951 vdd.n2288 gnd 0.004834f
C3952 vdd.n2289 gnd 0.017634f
C3953 vdd.n2290 gnd 0.004297f
C3954 vdd.n2291 gnd 0.006087f
C3955 vdd.n2292 gnd 0.397947f
C3956 vdd.n2293 gnd 0.006087f
C3957 vdd.n2294 gnd 0.006087f
C3958 vdd.n2295 gnd 0.006087f
C3959 vdd.n2296 gnd 0.006087f
C3960 vdd.n2297 gnd 0.006087f
C3961 vdd.n2298 gnd 0.361354f
C3962 vdd.n2299 gnd 0.006087f
C3963 vdd.n2300 gnd 0.006087f
C3964 vdd.n2301 gnd 0.006087f
C3965 vdd.n2302 gnd 0.006087f
C3966 vdd.n2303 gnd 0.006087f
C3967 vdd.n2304 gnd 0.498577f
C3968 vdd.n2305 gnd 0.006087f
C3969 vdd.n2306 gnd 0.006087f
C3970 vdd.n2307 gnd 0.006087f
C3971 vdd.n2308 gnd 0.006087f
C3972 vdd.n2309 gnd 0.006087f
C3973 vdd.n2310 gnd 0.548892f
C3974 vdd.n2311 gnd 0.006087f
C3975 vdd.n2312 gnd 0.006087f
C3976 vdd.n2313 gnd 0.006087f
C3977 vdd.n2314 gnd 0.006087f
C3978 vdd.n2315 gnd 0.006087f
C3979 vdd.n2316 gnd 0.411669f
C3980 vdd.n2317 gnd 0.006087f
C3981 vdd.n2318 gnd 0.006087f
C3982 vdd.n2319 gnd 0.006087f
C3983 vdd.n2320 gnd 0.006087f
C3984 vdd.n2321 gnd 0.006087f
C3985 vdd.n2322 gnd 0.196686f
C3986 vdd.n2323 gnd 0.006087f
C3987 vdd.n2324 gnd 0.006087f
C3988 vdd.n2325 gnd 0.006087f
C3989 vdd.n2326 gnd 0.006087f
C3990 vdd.n2327 gnd 0.006087f
C3991 vdd.n2328 gnd 0.196686f
C3992 vdd.n2329 gnd 0.006087f
C3993 vdd.n2330 gnd 0.006087f
C3994 vdd.n2331 gnd 0.006087f
C3995 vdd.n2332 gnd 0.006087f
C3996 vdd.n2333 gnd 0.006087f
C3997 vdd.n2334 gnd 0.622078f
C3998 vdd.n2335 gnd 0.006087f
C3999 vdd.n2336 gnd 0.006087f
C4000 vdd.n2337 gnd 0.006087f
C4001 vdd.n2338 gnd 0.006087f
C4002 vdd.n2339 gnd 0.006087f
C4003 vdd.n2340 gnd 0.006087f
C4004 vdd.n2341 gnd 0.006087f
C4005 vdd.n2342 gnd 0.429965f
C4006 vdd.n2343 gnd 0.006087f
C4007 vdd.n2344 gnd 0.006087f
C4008 vdd.n2345 gnd 0.006087f
C4009 vdd.n2346 gnd 0.006087f
C4010 vdd.n2347 gnd 0.006087f
C4011 vdd.n2348 gnd 0.006087f
C4012 vdd.n2349 gnd 0.388799f
C4013 vdd.n2350 gnd 0.006087f
C4014 vdd.n2351 gnd 0.006087f
C4015 vdd.n2352 gnd 0.006087f
C4016 vdd.n2353 gnd 0.013821f
C4017 vdd.n2354 gnd 0.013034f
C4018 vdd.n2355 gnd 0.006087f
C4019 vdd.n2356 gnd 0.006087f
C4020 vdd.n2357 gnd 0.0047f
C4021 vdd.n2358 gnd 0.006087f
C4022 vdd.n2359 gnd 0.006087f
C4023 vdd.n2360 gnd 0.004431f
C4024 vdd.n2361 gnd 0.006087f
C4025 vdd.n2362 gnd 0.006087f
C4026 vdd.n2363 gnd 0.006087f
C4027 vdd.n2364 gnd 0.006087f
C4028 vdd.n2365 gnd 0.006087f
C4029 vdd.n2366 gnd 0.006087f
C4030 vdd.n2367 gnd 0.006087f
C4031 vdd.n2368 gnd 0.006087f
C4032 vdd.n2369 gnd 0.006087f
C4033 vdd.n2370 gnd 0.006087f
C4034 vdd.n2371 gnd 0.006087f
C4035 vdd.n2372 gnd 0.006087f
C4036 vdd.n2373 gnd 0.006087f
C4037 vdd.n2374 gnd 0.006087f
C4038 vdd.n2375 gnd 0.006087f
C4039 vdd.n2376 gnd 0.006087f
C4040 vdd.n2377 gnd 0.006087f
C4041 vdd.n2378 gnd 0.006087f
C4042 vdd.n2379 gnd 0.006087f
C4043 vdd.n2380 gnd 0.006087f
C4044 vdd.n2381 gnd 0.006087f
C4045 vdd.n2382 gnd 0.006087f
C4046 vdd.n2383 gnd 0.006087f
C4047 vdd.n2384 gnd 0.006087f
C4048 vdd.n2385 gnd 0.006087f
C4049 vdd.n2386 gnd 0.006087f
C4050 vdd.n2387 gnd 0.006087f
C4051 vdd.n2388 gnd 0.006087f
C4052 vdd.n2389 gnd 0.006087f
C4053 vdd.n2390 gnd 0.006087f
C4054 vdd.n2391 gnd 0.006087f
C4055 vdd.n2392 gnd 0.006087f
C4056 vdd.n2393 gnd 0.006087f
C4057 vdd.n2394 gnd 0.006087f
C4058 vdd.n2395 gnd 0.006087f
C4059 vdd.n2396 gnd 0.006087f
C4060 vdd.n2397 gnd 0.006087f
C4061 vdd.n2398 gnd 0.006087f
C4062 vdd.n2399 gnd 0.006087f
C4063 vdd.n2400 gnd 0.006087f
C4064 vdd.n2401 gnd 0.006087f
C4065 vdd.n2402 gnd 0.006087f
C4066 vdd.n2403 gnd 0.006087f
C4067 vdd.n2404 gnd 0.006087f
C4068 vdd.n2405 gnd 0.006087f
C4069 vdd.n2406 gnd 0.006087f
C4070 vdd.n2407 gnd 0.006087f
C4071 vdd.n2408 gnd 0.006087f
C4072 vdd.n2409 gnd 0.006087f
C4073 vdd.n2410 gnd 0.006087f
C4074 vdd.n2411 gnd 0.006087f
C4075 vdd.n2412 gnd 0.006087f
C4076 vdd.n2413 gnd 0.006087f
C4077 vdd.n2414 gnd 0.006087f
C4078 vdd.n2415 gnd 0.006087f
C4079 vdd.n2416 gnd 0.006087f
C4080 vdd.n2417 gnd 0.006087f
C4081 vdd.n2418 gnd 0.006087f
C4082 vdd.n2419 gnd 0.006087f
C4083 vdd.n2420 gnd 0.006087f
C4084 vdd.n2421 gnd 0.013821f
C4085 vdd.n2422 gnd 0.013034f
C4086 vdd.n2423 gnd 0.013034f
C4087 vdd.n2424 gnd 0.704411f
C4088 vdd.n2425 gnd 0.013034f
C4089 vdd.n2426 gnd 0.013821f
C4090 vdd.n2427 gnd 0.013034f
C4091 vdd.n2428 gnd 0.006087f
C4092 vdd.n2429 gnd 0.006087f
C4093 vdd.n2430 gnd 0.006087f
C4094 vdd.n2431 gnd 0.0047f
C4095 vdd.n2432 gnd 0.0087f
C4096 vdd.n2433 gnd 0.004431f
C4097 vdd.n2434 gnd 0.006087f
C4098 vdd.n2435 gnd 0.006087f
C4099 vdd.n2436 gnd 0.006087f
C4100 vdd.n2437 gnd 0.006087f
C4101 vdd.n2438 gnd 0.006087f
C4102 vdd.n2439 gnd 0.006087f
C4103 vdd.n2440 gnd 0.006087f
C4104 vdd.n2441 gnd 0.006087f
C4105 vdd.n2442 gnd 0.006087f
C4106 vdd.n2443 gnd 0.006087f
C4107 vdd.n2444 gnd 0.006087f
C4108 vdd.n2445 gnd 0.006087f
C4109 vdd.n2446 gnd 0.006087f
C4110 vdd.n2447 gnd 0.006087f
C4111 vdd.n2448 gnd 0.006087f
C4112 vdd.n2449 gnd 0.006087f
C4113 vdd.n2450 gnd 0.006087f
C4114 vdd.n2451 gnd 0.006087f
C4115 vdd.n2452 gnd 0.006087f
C4116 vdd.n2453 gnd 0.006087f
C4117 vdd.n2454 gnd 0.006087f
C4118 vdd.n2455 gnd 0.006087f
C4119 vdd.n2456 gnd 0.006087f
C4120 vdd.n2457 gnd 0.006087f
C4121 vdd.n2458 gnd 0.006087f
C4122 vdd.n2459 gnd 0.006087f
C4123 vdd.n2460 gnd 0.006087f
C4124 vdd.n2461 gnd 0.006087f
C4125 vdd.n2462 gnd 0.006087f
C4126 vdd.n2463 gnd 0.006087f
C4127 vdd.n2464 gnd 0.006087f
C4128 vdd.n2465 gnd 0.006087f
C4129 vdd.n2466 gnd 0.006087f
C4130 vdd.n2467 gnd 0.006087f
C4131 vdd.n2468 gnd 0.006087f
C4132 vdd.n2469 gnd 0.006087f
C4133 vdd.n2470 gnd 0.006087f
C4134 vdd.n2471 gnd 0.006087f
C4135 vdd.n2472 gnd 0.006087f
C4136 vdd.n2473 gnd 0.006087f
C4137 vdd.n2474 gnd 0.006087f
C4138 vdd.n2475 gnd 0.006087f
C4139 vdd.n2476 gnd 0.006087f
C4140 vdd.n2477 gnd 0.006087f
C4141 vdd.n2478 gnd 0.006087f
C4142 vdd.n2479 gnd 0.006087f
C4143 vdd.n2480 gnd 0.006087f
C4144 vdd.n2481 gnd 0.006087f
C4145 vdd.n2482 gnd 0.006087f
C4146 vdd.n2483 gnd 0.006087f
C4147 vdd.n2484 gnd 0.006087f
C4148 vdd.n2485 gnd 0.006087f
C4149 vdd.n2486 gnd 0.006087f
C4150 vdd.n2487 gnd 0.006087f
C4151 vdd.n2488 gnd 0.006087f
C4152 vdd.n2489 gnd 0.006087f
C4153 vdd.n2490 gnd 0.006087f
C4154 vdd.n2491 gnd 0.006087f
C4155 vdd.n2492 gnd 0.006087f
C4156 vdd.n2493 gnd 0.006087f
C4157 vdd.n2494 gnd 0.013821f
C4158 vdd.n2495 gnd 0.013821f
C4159 vdd.n2496 gnd 0.759301f
C4160 vdd.t200 gnd 2.69872f
C4161 vdd.t187 gnd 2.69872f
C4162 vdd.n2530 gnd 0.013821f
C4163 vdd.t205 gnd 0.530596f
C4164 vdd.n2531 gnd 0.006087f
C4165 vdd.t68 gnd 0.245981f
C4166 vdd.t69 gnd 0.251792f
C4167 vdd.t66 gnd 0.160586f
C4168 vdd.n2532 gnd 0.086788f
C4169 vdd.n2533 gnd 0.049229f
C4170 vdd.n2534 gnd 0.006087f
C4171 vdd.t78 gnd 0.245981f
C4172 vdd.t79 gnd 0.251792f
C4173 vdd.t77 gnd 0.160586f
C4174 vdd.n2535 gnd 0.086788f
C4175 vdd.n2536 gnd 0.049229f
C4176 vdd.n2537 gnd 0.0087f
C4177 vdd.n2538 gnd 0.013821f
C4178 vdd.n2539 gnd 0.013821f
C4179 vdd.n2540 gnd 0.006087f
C4180 vdd.n2541 gnd 0.006087f
C4181 vdd.n2542 gnd 0.006087f
C4182 vdd.n2543 gnd 0.006087f
C4183 vdd.n2544 gnd 0.006087f
C4184 vdd.n2545 gnd 0.006087f
C4185 vdd.n2546 gnd 0.006087f
C4186 vdd.n2547 gnd 0.006087f
C4187 vdd.n2548 gnd 0.006087f
C4188 vdd.n2549 gnd 0.006087f
C4189 vdd.n2550 gnd 0.006087f
C4190 vdd.n2551 gnd 0.006087f
C4191 vdd.n2552 gnd 0.006087f
C4192 vdd.n2553 gnd 0.006087f
C4193 vdd.n2554 gnd 0.006087f
C4194 vdd.n2555 gnd 0.006087f
C4195 vdd.n2556 gnd 0.006087f
C4196 vdd.n2557 gnd 0.006087f
C4197 vdd.n2558 gnd 0.006087f
C4198 vdd.n2559 gnd 0.006087f
C4199 vdd.n2560 gnd 0.006087f
C4200 vdd.n2561 gnd 0.006087f
C4201 vdd.n2562 gnd 0.006087f
C4202 vdd.n2563 gnd 0.006087f
C4203 vdd.n2564 gnd 0.006087f
C4204 vdd.n2565 gnd 0.006087f
C4205 vdd.n2566 gnd 0.006087f
C4206 vdd.n2567 gnd 0.006087f
C4207 vdd.n2568 gnd 0.006087f
C4208 vdd.n2569 gnd 0.006087f
C4209 vdd.n2570 gnd 0.006087f
C4210 vdd.n2571 gnd 0.006087f
C4211 vdd.n2572 gnd 0.006087f
C4212 vdd.n2573 gnd 0.006087f
C4213 vdd.n2574 gnd 0.006087f
C4214 vdd.n2575 gnd 0.006087f
C4215 vdd.n2576 gnd 0.006087f
C4216 vdd.n2577 gnd 0.006087f
C4217 vdd.n2578 gnd 0.006087f
C4218 vdd.n2579 gnd 0.006087f
C4219 vdd.n2580 gnd 0.006087f
C4220 vdd.n2581 gnd 0.006087f
C4221 vdd.n2582 gnd 0.006087f
C4222 vdd.n2583 gnd 0.006087f
C4223 vdd.n2584 gnd 0.006087f
C4224 vdd.n2585 gnd 0.006087f
C4225 vdd.n2586 gnd 0.006087f
C4226 vdd.n2587 gnd 0.006087f
C4227 vdd.n2588 gnd 0.006087f
C4228 vdd.n2589 gnd 0.006087f
C4229 vdd.n2590 gnd 0.006087f
C4230 vdd.n2591 gnd 0.006087f
C4231 vdd.n2592 gnd 0.006087f
C4232 vdd.n2593 gnd 0.006087f
C4233 vdd.n2594 gnd 0.006087f
C4234 vdd.n2595 gnd 0.006087f
C4235 vdd.n2596 gnd 0.006087f
C4236 vdd.n2597 gnd 0.006087f
C4237 vdd.n2598 gnd 0.006087f
C4238 vdd.n2599 gnd 0.006087f
C4239 vdd.n2600 gnd 0.004431f
C4240 vdd.n2601 gnd 0.006087f
C4241 vdd.n2602 gnd 0.006087f
C4242 vdd.n2603 gnd 0.0047f
C4243 vdd.n2604 gnd 0.006087f
C4244 vdd.n2605 gnd 0.006087f
C4245 vdd.n2606 gnd 0.013821f
C4246 vdd.n2607 gnd 0.013034f
C4247 vdd.n2608 gnd 0.013034f
C4248 vdd.n2609 gnd 0.006087f
C4249 vdd.n2610 gnd 0.006087f
C4250 vdd.n2611 gnd 0.006087f
C4251 vdd.n2612 gnd 0.006087f
C4252 vdd.n2613 gnd 0.006087f
C4253 vdd.n2614 gnd 0.006087f
C4254 vdd.n2615 gnd 0.006087f
C4255 vdd.n2616 gnd 0.006087f
C4256 vdd.n2617 gnd 0.006087f
C4257 vdd.n2618 gnd 0.006087f
C4258 vdd.n2619 gnd 0.006087f
C4259 vdd.n2620 gnd 0.006087f
C4260 vdd.n2621 gnd 0.006087f
C4261 vdd.n2622 gnd 0.006087f
C4262 vdd.n2623 gnd 0.006087f
C4263 vdd.n2624 gnd 0.006087f
C4264 vdd.n2625 gnd 0.006087f
C4265 vdd.n2626 gnd 0.006087f
C4266 vdd.n2627 gnd 0.006087f
C4267 vdd.n2628 gnd 0.006087f
C4268 vdd.n2629 gnd 0.006087f
C4269 vdd.n2630 gnd 0.006087f
C4270 vdd.n2631 gnd 0.006087f
C4271 vdd.n2632 gnd 0.006087f
C4272 vdd.n2633 gnd 0.006087f
C4273 vdd.n2634 gnd 0.006087f
C4274 vdd.n2635 gnd 0.006087f
C4275 vdd.n2636 gnd 0.006087f
C4276 vdd.n2637 gnd 0.006087f
C4277 vdd.n2638 gnd 0.006087f
C4278 vdd.n2639 gnd 0.006087f
C4279 vdd.n2640 gnd 0.006087f
C4280 vdd.n2641 gnd 0.006087f
C4281 vdd.n2642 gnd 0.006087f
C4282 vdd.n2643 gnd 0.006087f
C4283 vdd.n2644 gnd 0.006087f
C4284 vdd.n2645 gnd 0.006087f
C4285 vdd.n2646 gnd 0.006087f
C4286 vdd.n2647 gnd 0.006087f
C4287 vdd.n2648 gnd 0.006087f
C4288 vdd.n2649 gnd 0.006087f
C4289 vdd.n2650 gnd 0.006087f
C4290 vdd.n2651 gnd 0.006087f
C4291 vdd.n2652 gnd 0.006087f
C4292 vdd.n2653 gnd 0.006087f
C4293 vdd.n2654 gnd 0.006087f
C4294 vdd.n2655 gnd 0.006087f
C4295 vdd.n2656 gnd 0.006087f
C4296 vdd.n2657 gnd 0.006087f
C4297 vdd.n2658 gnd 0.006087f
C4298 vdd.n2659 gnd 0.006087f
C4299 vdd.n2660 gnd 0.006087f
C4300 vdd.n2661 gnd 0.006087f
C4301 vdd.n2662 gnd 0.006087f
C4302 vdd.n2663 gnd 0.006087f
C4303 vdd.n2664 gnd 0.006087f
C4304 vdd.n2665 gnd 0.006087f
C4305 vdd.n2666 gnd 0.006087f
C4306 vdd.n2667 gnd 0.006087f
C4307 vdd.n2668 gnd 0.006087f
C4308 vdd.n2669 gnd 0.006087f
C4309 vdd.n2670 gnd 0.006087f
C4310 vdd.n2671 gnd 0.006087f
C4311 vdd.n2672 gnd 0.006087f
C4312 vdd.n2673 gnd 0.006087f
C4313 vdd.n2674 gnd 0.006087f
C4314 vdd.n2675 gnd 0.006087f
C4315 vdd.n2676 gnd 0.006087f
C4316 vdd.n2677 gnd 0.006087f
C4317 vdd.n2678 gnd 0.006087f
C4318 vdd.n2679 gnd 0.006087f
C4319 vdd.n2680 gnd 0.006087f
C4320 vdd.n2681 gnd 0.006087f
C4321 vdd.n2682 gnd 0.006087f
C4322 vdd.n2683 gnd 0.006087f
C4323 vdd.n2684 gnd 0.006087f
C4324 vdd.n2685 gnd 0.006087f
C4325 vdd.n2686 gnd 0.006087f
C4326 vdd.n2687 gnd 0.006087f
C4327 vdd.n2688 gnd 0.006087f
C4328 vdd.n2689 gnd 0.006087f
C4329 vdd.n2690 gnd 0.006087f
C4330 vdd.n2691 gnd 0.006087f
C4331 vdd.n2692 gnd 0.006087f
C4332 vdd.n2693 gnd 0.006087f
C4333 vdd.n2694 gnd 0.006087f
C4334 vdd.n2695 gnd 0.006087f
C4335 vdd.n2696 gnd 0.006087f
C4336 vdd.n2697 gnd 0.006087f
C4337 vdd.n2698 gnd 0.006087f
C4338 vdd.n2699 gnd 0.006087f
C4339 vdd.n2700 gnd 0.006087f
C4340 vdd.n2701 gnd 0.006087f
C4341 vdd.n2702 gnd 0.006087f
C4342 vdd.n2703 gnd 0.006087f
C4343 vdd.n2704 gnd 0.006087f
C4344 vdd.n2705 gnd 0.006087f
C4345 vdd.n2706 gnd 0.006087f
C4346 vdd.n2707 gnd 0.006087f
C4347 vdd.n2708 gnd 0.006087f
C4348 vdd.n2709 gnd 0.006087f
C4349 vdd.n2710 gnd 0.196686f
C4350 vdd.n2711 gnd 0.006087f
C4351 vdd.n2712 gnd 0.006087f
C4352 vdd.n2713 gnd 0.006087f
C4353 vdd.n2714 gnd 0.006087f
C4354 vdd.n2715 gnd 0.006087f
C4355 vdd.n2716 gnd 0.196686f
C4356 vdd.n2717 gnd 0.006087f
C4357 vdd.n2718 gnd 0.006087f
C4358 vdd.n2719 gnd 0.006087f
C4359 vdd.n2720 gnd 0.006087f
C4360 vdd.n2721 gnd 0.006087f
C4361 vdd.n2722 gnd 0.006087f
C4362 vdd.n2723 gnd 0.006087f
C4363 vdd.n2724 gnd 0.006087f
C4364 vdd.n2725 gnd 0.006087f
C4365 vdd.n2726 gnd 0.006087f
C4366 vdd.n2727 gnd 0.006087f
C4367 vdd.n2728 gnd 0.388799f
C4368 vdd.n2729 gnd 0.006087f
C4369 vdd.n2730 gnd 0.006087f
C4370 vdd.n2731 gnd 0.006087f
C4371 vdd.n2732 gnd 0.013034f
C4372 vdd.n2733 gnd 0.013034f
C4373 vdd.n2734 gnd 0.013821f
C4374 vdd.n2735 gnd 0.013821f
C4375 vdd.n2736 gnd 0.006087f
C4376 vdd.n2737 gnd 0.006087f
C4377 vdd.n2738 gnd 0.006087f
C4378 vdd.n2739 gnd 0.0047f
C4379 vdd.n2740 gnd 0.0087f
C4380 vdd.n2741 gnd 0.004431f
C4381 vdd.n2742 gnd 0.006087f
C4382 vdd.n2743 gnd 0.006087f
C4383 vdd.n2744 gnd 0.006087f
C4384 vdd.n2745 gnd 0.006087f
C4385 vdd.n2746 gnd 0.006087f
C4386 vdd.n2747 gnd 0.006087f
C4387 vdd.n2748 gnd 0.006087f
C4388 vdd.n2749 gnd 0.006087f
C4389 vdd.n2750 gnd 0.006087f
C4390 vdd.n2751 gnd 0.006087f
C4391 vdd.n2752 gnd 0.006087f
C4392 vdd.n2753 gnd 0.006087f
C4393 vdd.n2754 gnd 0.006087f
C4394 vdd.n2755 gnd 0.006087f
C4395 vdd.n2756 gnd 0.006087f
C4396 vdd.n2757 gnd 0.006087f
C4397 vdd.n2758 gnd 0.006087f
C4398 vdd.n2759 gnd 0.006087f
C4399 vdd.n2760 gnd 0.006087f
C4400 vdd.n2761 gnd 0.006087f
C4401 vdd.n2762 gnd 0.006087f
C4402 vdd.n2763 gnd 0.006087f
C4403 vdd.n2764 gnd 0.006087f
C4404 vdd.n2765 gnd 0.006087f
C4405 vdd.n2766 gnd 0.006087f
C4406 vdd.n2767 gnd 0.006087f
C4407 vdd.n2768 gnd 0.006087f
C4408 vdd.n2769 gnd 0.006087f
C4409 vdd.n2770 gnd 0.006087f
C4410 vdd.n2771 gnd 0.006087f
C4411 vdd.n2772 gnd 0.006087f
C4412 vdd.n2773 gnd 0.006087f
C4413 vdd.n2774 gnd 0.006087f
C4414 vdd.n2775 gnd 0.006087f
C4415 vdd.n2776 gnd 0.006087f
C4416 vdd.n2777 gnd 0.006087f
C4417 vdd.n2778 gnd 0.006087f
C4418 vdd.n2779 gnd 0.006087f
C4419 vdd.n2780 gnd 0.006087f
C4420 vdd.n2781 gnd 0.006087f
C4421 vdd.n2782 gnd 0.006087f
C4422 vdd.n2783 gnd 0.006087f
C4423 vdd.n2784 gnd 0.006087f
C4424 vdd.n2785 gnd 0.006087f
C4425 vdd.n2786 gnd 0.006087f
C4426 vdd.n2787 gnd 0.006087f
C4427 vdd.n2788 gnd 0.006087f
C4428 vdd.n2789 gnd 0.006087f
C4429 vdd.n2790 gnd 0.006087f
C4430 vdd.n2791 gnd 0.006087f
C4431 vdd.n2792 gnd 0.006087f
C4432 vdd.n2793 gnd 0.006087f
C4433 vdd.n2794 gnd 0.006087f
C4434 vdd.n2795 gnd 0.006087f
C4435 vdd.n2796 gnd 0.006087f
C4436 vdd.n2797 gnd 0.006087f
C4437 vdd.n2798 gnd 0.006087f
C4438 vdd.n2799 gnd 0.006087f
C4439 vdd.n2800 gnd 0.759301f
C4440 vdd.n2802 gnd 0.013821f
C4441 vdd.n2803 gnd 0.013821f
C4442 vdd.n2804 gnd 0.013034f
C4443 vdd.n2805 gnd 0.006087f
C4444 vdd.n2806 gnd 0.006087f
C4445 vdd.n2807 gnd 0.365928f
C4446 vdd.n2808 gnd 0.006087f
C4447 vdd.n2809 gnd 0.006087f
C4448 vdd.n2810 gnd 0.006087f
C4449 vdd.n2811 gnd 0.006087f
C4450 vdd.n2812 gnd 0.006087f
C4451 vdd.n2813 gnd 0.370502f
C4452 vdd.n2814 gnd 0.006087f
C4453 vdd.n2815 gnd 0.006087f
C4454 vdd.n2816 gnd 0.006087f
C4455 vdd.n2817 gnd 0.006087f
C4456 vdd.n2818 gnd 0.006087f
C4457 vdd.n2819 gnd 0.622078f
C4458 vdd.n2820 gnd 0.006087f
C4459 vdd.n2821 gnd 0.006087f
C4460 vdd.n2822 gnd 0.006087f
C4461 vdd.n2823 gnd 0.006087f
C4462 vdd.n2824 gnd 0.006087f
C4463 vdd.n2825 gnd 0.448262f
C4464 vdd.n2826 gnd 0.006087f
C4465 vdd.n2827 gnd 0.006087f
C4466 vdd.n2828 gnd 0.006087f
C4467 vdd.n2829 gnd 0.006087f
C4468 vdd.n2830 gnd 0.006087f
C4469 vdd.n2831 gnd 0.562614f
C4470 vdd.n2832 gnd 0.006087f
C4471 vdd.n2833 gnd 0.006087f
C4472 vdd.n2834 gnd 0.006087f
C4473 vdd.n2835 gnd 0.006087f
C4474 vdd.n2836 gnd 0.006087f
C4475 vdd.n2837 gnd 0.461984f
C4476 vdd.n2838 gnd 0.006087f
C4477 vdd.n2839 gnd 0.006087f
C4478 vdd.n2840 gnd 0.006087f
C4479 vdd.n2841 gnd 0.006087f
C4480 vdd.n2842 gnd 0.006087f
C4481 vdd.n2843 gnd 0.324761f
C4482 vdd.n2844 gnd 0.006087f
C4483 vdd.n2845 gnd 0.006087f
C4484 vdd.n2846 gnd 0.006087f
C4485 vdd.n2847 gnd 0.006087f
C4486 vdd.n2848 gnd 0.006087f
C4487 vdd.n2849 gnd 0.196686f
C4488 vdd.n2850 gnd 0.006087f
C4489 vdd.n2851 gnd 0.006087f
C4490 vdd.n2852 gnd 0.006087f
C4491 vdd.n2853 gnd 0.006087f
C4492 vdd.n2854 gnd 0.006087f
C4493 vdd.n2855 gnd 0.571763f
C4494 vdd.n2856 gnd 0.006087f
C4495 vdd.n2857 gnd 0.006087f
C4496 vdd.n2858 gnd 0.006087f
C4497 vdd.n2859 gnd 0.004297f
C4498 vdd.n2860 gnd 0.006087f
C4499 vdd.n2861 gnd 0.006087f
C4500 vdd.n2862 gnd 0.622078f
C4501 vdd.n2863 gnd 0.006087f
C4502 vdd.n2864 gnd 0.006087f
C4503 vdd.n2865 gnd 0.006087f
C4504 vdd.n2866 gnd 0.006087f
C4505 vdd.n2867 gnd 0.006087f
C4506 vdd.n2868 gnd 0.494003f
C4507 vdd.n2869 gnd 0.006087f
C4508 vdd.n2870 gnd 0.004834f
C4509 vdd.n2871 gnd 0.006087f
C4510 vdd.n2872 gnd 0.006087f
C4511 vdd.n2873 gnd 0.006087f
C4512 vdd.n2874 gnd 0.397947f
C4513 vdd.n2875 gnd 0.006087f
C4514 vdd.n2876 gnd 0.006087f
C4515 vdd.n2877 gnd 0.006087f
C4516 vdd.n2878 gnd 0.006087f
C4517 vdd.n2879 gnd 0.006087f
C4518 vdd.n2880 gnd 0.361354f
C4519 vdd.n2881 gnd 0.006087f
C4520 vdd.n2882 gnd 0.006087f
C4521 vdd.n2883 gnd 0.006087f
C4522 vdd.n2884 gnd 0.006087f
C4523 vdd.n2885 gnd 0.006087f
C4524 vdd.n2886 gnd 0.498577f
C4525 vdd.n2887 gnd 0.006087f
C4526 vdd.n2888 gnd 0.006087f
C4527 vdd.n2889 gnd 0.006087f
C4528 vdd.n2890 gnd 0.006087f
C4529 vdd.n2891 gnd 0.006087f
C4530 vdd.n2892 gnd 0.622078f
C4531 vdd.n2893 gnd 0.006087f
C4532 vdd.n2894 gnd 0.006087f
C4533 vdd.n2895 gnd 0.006087f
C4534 vdd.n2896 gnd 0.006087f
C4535 vdd.n2897 gnd 0.006087f
C4536 vdd.n2898 gnd 0.608355f
C4537 vdd.n2899 gnd 0.006087f
C4538 vdd.n2900 gnd 0.006087f
C4539 vdd.n2901 gnd 0.006087f
C4540 vdd.n2902 gnd 0.006087f
C4541 vdd.n2903 gnd 0.006087f
C4542 vdd.n2904 gnd 0.471132f
C4543 vdd.n2905 gnd 0.006087f
C4544 vdd.n2906 gnd 0.006087f
C4545 vdd.n2907 gnd 0.006087f
C4546 vdd.n2908 gnd 0.006087f
C4547 vdd.n2909 gnd 0.006087f
C4548 vdd.n2910 gnd 0.333909f
C4549 vdd.n2911 gnd 0.006087f
C4550 vdd.n2912 gnd 0.006087f
C4551 vdd.n2913 gnd 0.006087f
C4552 vdd.n2914 gnd 0.006087f
C4553 vdd.n2915 gnd 0.006087f
C4554 vdd.n2916 gnd 0.622078f
C4555 vdd.n2917 gnd 0.006087f
C4556 vdd.n2918 gnd 0.006087f
C4557 vdd.n2919 gnd 0.006087f
C4558 vdd.n2920 gnd 0.006087f
C4559 vdd.n2921 gnd 0.006087f
C4560 vdd.n2922 gnd 0.006087f
C4561 vdd.n2924 gnd 0.006087f
C4562 vdd.n2925 gnd 0.006087f
C4563 vdd.n2927 gnd 0.006087f
C4564 vdd.n2928 gnd 0.006087f
C4565 vdd.n2931 gnd 0.006087f
C4566 vdd.n2932 gnd 0.006087f
C4567 vdd.n2933 gnd 0.006087f
C4568 vdd.n2934 gnd 0.006087f
C4569 vdd.n2936 gnd 0.006087f
C4570 vdd.n2937 gnd 0.006087f
C4571 vdd.n2938 gnd 0.006087f
C4572 vdd.n2939 gnd 0.006087f
C4573 vdd.n2940 gnd 0.006087f
C4574 vdd.n2941 gnd 0.006087f
C4575 vdd.n2943 gnd 0.006087f
C4576 vdd.n2944 gnd 0.006087f
C4577 vdd.n2945 gnd 0.006087f
C4578 vdd.n2946 gnd 0.006087f
C4579 vdd.n2947 gnd 0.006087f
C4580 vdd.n2948 gnd 0.006087f
C4581 vdd.n2950 gnd 0.006087f
C4582 vdd.n2951 gnd 0.006087f
C4583 vdd.n2952 gnd 0.006087f
C4584 vdd.n2953 gnd 0.006087f
C4585 vdd.n2954 gnd 0.006087f
C4586 vdd.n2955 gnd 0.006087f
C4587 vdd.n2957 gnd 0.006087f
C4588 vdd.n2958 gnd 0.013821f
C4589 vdd.n2959 gnd 0.013821f
C4590 vdd.n2960 gnd 0.013034f
C4591 vdd.n2961 gnd 0.006087f
C4592 vdd.n2962 gnd 0.006087f
C4593 vdd.n2963 gnd 0.006087f
C4594 vdd.n2964 gnd 0.006087f
C4595 vdd.n2965 gnd 0.006087f
C4596 vdd.n2966 gnd 0.006087f
C4597 vdd.n2967 gnd 0.622078f
C4598 vdd.n2968 gnd 0.006087f
C4599 vdd.n2969 gnd 0.006087f
C4600 vdd.n2970 gnd 0.006087f
C4601 vdd.n2971 gnd 0.006087f
C4602 vdd.n2972 gnd 0.006087f
C4603 vdd.n2973 gnd 0.443688f
C4604 vdd.n2974 gnd 0.006087f
C4605 vdd.n2975 gnd 0.006087f
C4606 vdd.n2976 gnd 0.006087f
C4607 vdd.n2977 gnd 0.013821f
C4608 vdd.n2979 gnd 0.013821f
C4609 vdd.n2980 gnd 0.013034f
C4610 vdd.n2981 gnd 0.006087f
C4611 vdd.n2982 gnd 0.0047f
C4612 vdd.n2983 gnd 0.006087f
C4613 vdd.n2985 gnd 0.006087f
C4614 vdd.n2986 gnd 0.006087f
C4615 vdd.n2987 gnd 0.006087f
C4616 vdd.n2988 gnd 0.006087f
C4617 vdd.n2989 gnd 0.006087f
C4618 vdd.n2990 gnd 0.006087f
C4619 vdd.n2992 gnd 0.006087f
C4620 vdd.n2993 gnd 0.006087f
C4621 vdd.n2994 gnd 0.006087f
C4622 vdd.n2995 gnd 0.006087f
C4623 vdd.n2996 gnd 0.006087f
C4624 vdd.n2997 gnd 0.006087f
C4625 vdd.n2999 gnd 0.006087f
C4626 vdd.n3000 gnd 0.006087f
C4627 vdd.n3001 gnd 0.006087f
C4628 vdd.n3002 gnd 0.006087f
C4629 vdd.n3003 gnd 0.006087f
C4630 vdd.n3004 gnd 0.006087f
C4631 vdd.n3006 gnd 0.006087f
C4632 vdd.n3007 gnd 0.006087f
C4633 vdd.n3008 gnd 0.006087f
C4634 vdd.n3009 gnd 0.953733f
C4635 vdd.n3010 gnd 0.037587f
C4636 vdd.n3011 gnd 0.006087f
C4637 vdd.n3012 gnd 0.006087f
C4638 vdd.n3014 gnd 0.006087f
C4639 vdd.n3015 gnd 0.006087f
C4640 vdd.n3016 gnd 0.006087f
C4641 vdd.n3017 gnd 0.006087f
C4642 vdd.n3018 gnd 0.006087f
C4643 vdd.n3019 gnd 0.006087f
C4644 vdd.n3021 gnd 0.006087f
C4645 vdd.n3022 gnd 0.006087f
C4646 vdd.n3023 gnd 0.006087f
C4647 vdd.n3024 gnd 0.006087f
C4648 vdd.n3025 gnd 0.006087f
C4649 vdd.n3026 gnd 0.006087f
C4650 vdd.n3028 gnd 0.006087f
C4651 vdd.n3029 gnd 0.006087f
C4652 vdd.n3030 gnd 0.006087f
C4653 vdd.n3031 gnd 0.006087f
C4654 vdd.n3032 gnd 0.006087f
C4655 vdd.n3033 gnd 0.006087f
C4656 vdd.n3035 gnd 0.006087f
C4657 vdd.n3036 gnd 0.006087f
C4658 vdd.n3038 gnd 0.006087f
C4659 vdd.n3039 gnd 0.006087f
C4660 vdd.n3040 gnd 0.013821f
C4661 vdd.n3041 gnd 0.013034f
C4662 vdd.n3042 gnd 0.013034f
C4663 vdd.n3043 gnd 0.841635f
C4664 vdd.n3044 gnd 0.013034f
C4665 vdd.n3045 gnd 0.013821f
C4666 vdd.n3046 gnd 0.013034f
C4667 vdd.n3047 gnd 0.006087f
C4668 vdd.n3048 gnd 0.0047f
C4669 vdd.n3049 gnd 0.006087f
C4670 vdd.n3051 gnd 0.006087f
C4671 vdd.n3052 gnd 0.006087f
C4672 vdd.n3053 gnd 0.006087f
C4673 vdd.n3054 gnd 0.006087f
C4674 vdd.n3055 gnd 0.006087f
C4675 vdd.n3056 gnd 0.006087f
C4676 vdd.n3058 gnd 0.006087f
C4677 vdd.n3059 gnd 0.006087f
C4678 vdd.n3060 gnd 0.006087f
C4679 vdd.n3061 gnd 0.006087f
C4680 vdd.n3062 gnd 0.006087f
C4681 vdd.n3063 gnd 0.006087f
C4682 vdd.n3065 gnd 0.006087f
C4683 vdd.n3066 gnd 0.006087f
C4684 vdd.n3067 gnd 0.006087f
C4685 vdd.n3068 gnd 0.006087f
C4686 vdd.n3069 gnd 0.006087f
C4687 vdd.n3070 gnd 0.006087f
C4688 vdd.n3072 gnd 0.006087f
C4689 vdd.n3073 gnd 0.006087f
C4690 vdd.n3075 gnd 0.006087f
C4691 vdd.n3076 gnd 0.037587f
C4692 vdd.n3077 gnd 0.953733f
C4693 vdd.n3078 gnd 0.007698f
C4694 vdd.n3079 gnd 0.003422f
C4695 vdd.t30 gnd 0.110129f
C4696 vdd.t31 gnd 0.117698f
C4697 vdd.t28 gnd 0.143827f
C4698 vdd.n3080 gnd 0.184366f
C4699 vdd.n3081 gnd 0.154901f
C4700 vdd.n3082 gnd 0.011096f
C4701 vdd.n3083 gnd 0.008952f
C4702 vdd.n3084 gnd 0.003783f
C4703 vdd.n3085 gnd 0.007205f
C4704 vdd.n3086 gnd 0.008952f
C4705 vdd.n3087 gnd 0.008952f
C4706 vdd.n3088 gnd 0.007205f
C4707 vdd.n3089 gnd 0.007205f
C4708 vdd.n3090 gnd 0.008952f
C4709 vdd.n3092 gnd 0.008952f
C4710 vdd.n3093 gnd 0.007205f
C4711 vdd.n3094 gnd 0.007205f
C4712 vdd.n3095 gnd 0.007205f
C4713 vdd.n3096 gnd 0.008952f
C4714 vdd.n3098 gnd 0.008952f
C4715 vdd.n3100 gnd 0.008952f
C4716 vdd.n3101 gnd 0.007205f
C4717 vdd.n3102 gnd 0.007205f
C4718 vdd.n3103 gnd 0.007205f
C4719 vdd.n3104 gnd 0.008952f
C4720 vdd.n3106 gnd 0.008952f
C4721 vdd.n3108 gnd 0.008952f
C4722 vdd.n3109 gnd 0.007205f
C4723 vdd.n3110 gnd 0.007205f
C4724 vdd.n3111 gnd 0.007205f
C4725 vdd.n3112 gnd 0.008952f
C4726 vdd.n3114 gnd 0.008952f
C4727 vdd.n3115 gnd 0.008952f
C4728 vdd.n3116 gnd 0.007205f
C4729 vdd.n3117 gnd 0.007205f
C4730 vdd.n3118 gnd 0.008952f
C4731 vdd.n3119 gnd 0.008952f
C4732 vdd.n3121 gnd 0.008952f
C4733 vdd.n3122 gnd 0.007205f
C4734 vdd.n3123 gnd 0.008952f
C4735 vdd.n3124 gnd 0.008952f
C4736 vdd.n3125 gnd 0.008952f
C4737 vdd.n3126 gnd 0.014698f
C4738 vdd.n3127 gnd 0.004899f
C4739 vdd.n3128 gnd 0.008952f
C4740 vdd.n3130 gnd 0.008952f
C4741 vdd.n3132 gnd 0.008952f
C4742 vdd.n3133 gnd 0.007205f
C4743 vdd.n3134 gnd 0.007205f
C4744 vdd.n3135 gnd 0.007205f
C4745 vdd.n3136 gnd 0.008952f
C4746 vdd.n3138 gnd 0.008952f
C4747 vdd.n3140 gnd 0.008952f
C4748 vdd.n3141 gnd 0.007205f
C4749 vdd.n3142 gnd 0.007205f
C4750 vdd.n3143 gnd 0.007205f
C4751 vdd.n3144 gnd 0.008952f
C4752 vdd.n3146 gnd 0.008952f
C4753 vdd.n3148 gnd 0.008952f
C4754 vdd.n3149 gnd 0.007205f
C4755 vdd.n3150 gnd 0.007205f
C4756 vdd.n3151 gnd 0.007205f
C4757 vdd.n3152 gnd 0.008952f
C4758 vdd.n3154 gnd 0.008952f
C4759 vdd.n3156 gnd 0.008952f
C4760 vdd.n3157 gnd 0.007205f
C4761 vdd.n3158 gnd 0.007205f
C4762 vdd.n3159 gnd 0.007205f
C4763 vdd.n3160 gnd 0.008952f
C4764 vdd.n3162 gnd 0.008952f
C4765 vdd.n3164 gnd 0.008952f
C4766 vdd.n3165 gnd 0.007205f
C4767 vdd.n3166 gnd 0.007205f
C4768 vdd.n3167 gnd 0.006016f
C4769 vdd.n3168 gnd 0.008952f
C4770 vdd.n3170 gnd 0.008952f
C4771 vdd.n3172 gnd 0.008952f
C4772 vdd.n3173 gnd 0.006016f
C4773 vdd.n3174 gnd 0.007205f
C4774 vdd.n3175 gnd 0.007205f
C4775 vdd.n3176 gnd 0.008952f
C4776 vdd.n3178 gnd 0.008952f
C4777 vdd.n3180 gnd 0.008952f
C4778 vdd.n3181 gnd 0.007205f
C4779 vdd.n3182 gnd 0.007205f
C4780 vdd.n3183 gnd 0.007205f
C4781 vdd.n3184 gnd 0.008952f
C4782 vdd.n3186 gnd 0.008952f
C4783 vdd.n3188 gnd 0.008952f
C4784 vdd.n3189 gnd 0.007205f
C4785 vdd.n3190 gnd 0.007205f
C4786 vdd.n3191 gnd 0.007205f
C4787 vdd.n3192 gnd 0.008952f
C4788 vdd.n3194 gnd 0.008952f
C4789 vdd.n3195 gnd 0.008952f
C4790 vdd.n3196 gnd 0.007205f
C4791 vdd.n3197 gnd 0.007205f
C4792 vdd.n3198 gnd 0.008952f
C4793 vdd.n3199 gnd 0.008952f
C4794 vdd.n3200 gnd 0.007205f
C4795 vdd.n3201 gnd 0.007205f
C4796 vdd.n3202 gnd 0.008952f
C4797 vdd.n3203 gnd 0.008952f
C4798 vdd.n3205 gnd 0.008952f
C4799 vdd.n3206 gnd 0.007205f
C4800 vdd.n3207 gnd 0.00598f
C4801 vdd.n3208 gnd 0.021425f
C4802 vdd.n3209 gnd 0.021096f
C4803 vdd.n3210 gnd 0.00598f
C4804 vdd.n3211 gnd 0.021096f
C4805 vdd.n3212 gnd 1.25788f
C4806 vdd.n3213 gnd 0.021096f
C4807 vdd.n3214 gnd 0.00598f
C4808 vdd.n3215 gnd 0.021096f
C4809 vdd.n3216 gnd 0.008952f
C4810 vdd.n3217 gnd 0.008952f
C4811 vdd.n3218 gnd 0.007205f
C4812 vdd.n3219 gnd 0.008952f
C4813 vdd.n3220 gnd 0.91482f
C4814 vdd.n3221 gnd 0.008952f
C4815 vdd.n3222 gnd 0.007205f
C4816 vdd.n3223 gnd 0.008952f
C4817 vdd.n3224 gnd 0.008952f
C4818 vdd.n3225 gnd 0.008952f
C4819 vdd.n3226 gnd 0.007205f
C4820 vdd.n3227 gnd 0.008952f
C4821 vdd.n3228 gnd 0.809616f
C4822 vdd.n3229 gnd 0.008952f
C4823 vdd.n3230 gnd 0.007205f
C4824 vdd.n3231 gnd 0.008952f
C4825 vdd.n3232 gnd 0.008952f
C4826 vdd.n3233 gnd 0.008952f
C4827 vdd.n3234 gnd 0.007205f
C4828 vdd.n3235 gnd 0.008952f
C4829 vdd.t112 gnd 0.45741f
C4830 vdd.n3236 gnd 0.654096f
C4831 vdd.n3237 gnd 0.008952f
C4832 vdd.n3238 gnd 0.007205f
C4833 vdd.n3239 gnd 0.008952f
C4834 vdd.n3240 gnd 0.008952f
C4835 vdd.n3241 gnd 0.008952f
C4836 vdd.n3242 gnd 0.007205f
C4837 vdd.n3243 gnd 0.008952f
C4838 vdd.n3244 gnd 0.498577f
C4839 vdd.n3245 gnd 0.008952f
C4840 vdd.n3246 gnd 0.007205f
C4841 vdd.n3247 gnd 0.008952f
C4842 vdd.n3248 gnd 0.008952f
C4843 vdd.n3249 gnd 0.008952f
C4844 vdd.n3250 gnd 0.007205f
C4845 vdd.n3251 gnd 0.008952f
C4846 vdd.n3252 gnd 0.644948f
C4847 vdd.n3253 gnd 0.571763f
C4848 vdd.n3254 gnd 0.008952f
C4849 vdd.n3255 gnd 0.007205f
C4850 vdd.n3256 gnd 0.008952f
C4851 vdd.n3257 gnd 0.008952f
C4852 vdd.n3258 gnd 0.008952f
C4853 vdd.n3259 gnd 0.007205f
C4854 vdd.n3260 gnd 0.008952f
C4855 vdd.n3261 gnd 0.727282f
C4856 vdd.n3262 gnd 0.008952f
C4857 vdd.n3263 gnd 0.007205f
C4858 vdd.n3264 gnd 0.008952f
C4859 vdd.n3265 gnd 0.008952f
C4860 vdd.n3266 gnd 0.008952f
C4861 vdd.n3267 gnd 0.007205f
C4862 vdd.n3268 gnd 0.007205f
C4863 vdd.n3269 gnd 0.007205f
C4864 vdd.n3270 gnd 0.008952f
C4865 vdd.n3271 gnd 0.008952f
C4866 vdd.n3272 gnd 0.008952f
C4867 vdd.n3273 gnd 0.007205f
C4868 vdd.n3274 gnd 0.007205f
C4869 vdd.n3275 gnd 0.007205f
C4870 vdd.n3276 gnd 0.008952f
C4871 vdd.n3277 gnd 0.008952f
C4872 vdd.n3278 gnd 0.008952f
C4873 vdd.n3279 gnd 0.007205f
C4874 vdd.n3280 gnd 0.007205f
C4875 vdd.n3281 gnd 0.007205f
C4876 vdd.n3282 gnd 0.008952f
C4877 vdd.n3283 gnd 0.008952f
C4878 vdd.n3284 gnd 0.008952f
C4879 vdd.n3285 gnd 0.007205f
C4880 vdd.n3286 gnd 0.007205f
C4881 vdd.n3287 gnd 0.00598f
C4882 vdd.n3288 gnd 0.021096f
C4883 vdd.n3289 gnd 0.021425f
C4884 vdd.n3291 gnd 0.021425f
C4885 vdd.n3292 gnd 0.003422f
C4886 vdd.t45 gnd 0.110129f
C4887 vdd.t44 gnd 0.117698f
C4888 vdd.t43 gnd 0.143827f
C4889 vdd.n3293 gnd 0.184366f
C4890 vdd.n3294 gnd 0.155622f
C4891 vdd.n3295 gnd 0.011816f
C4892 vdd.n3296 gnd 0.003783f
C4893 vdd.n3297 gnd 0.007205f
C4894 vdd.n3298 gnd 0.008952f
C4895 vdd.n3300 gnd 0.008952f
C4896 vdd.n3301 gnd 0.008952f
C4897 vdd.n3302 gnd 0.007205f
C4898 vdd.n3303 gnd 0.007205f
C4899 vdd.n3304 gnd 0.007205f
C4900 vdd.n3305 gnd 0.008952f
C4901 vdd.n3307 gnd 0.008952f
C4902 vdd.n3308 gnd 0.008952f
C4903 vdd.n3309 gnd 0.007205f
C4904 vdd.n3310 gnd 0.007205f
C4905 vdd.n3311 gnd 0.007205f
C4906 vdd.n3312 gnd 0.008952f
C4907 vdd.n3314 gnd 0.008952f
C4908 vdd.n3315 gnd 0.008952f
C4909 vdd.n3316 gnd 0.007205f
C4910 vdd.n3317 gnd 0.007205f
C4911 vdd.n3318 gnd 0.007205f
C4912 vdd.n3319 gnd 0.008952f
C4913 vdd.n3321 gnd 0.008952f
C4914 vdd.n3322 gnd 0.008952f
C4915 vdd.n3323 gnd 0.007205f
C4916 vdd.n3324 gnd 0.007205f
C4917 vdd.n3325 gnd 0.007205f
C4918 vdd.n3326 gnd 0.008952f
C4919 vdd.n3328 gnd 0.008952f
C4920 vdd.n3329 gnd 0.008952f
C4921 vdd.n3330 gnd 0.007205f
C4922 vdd.n3331 gnd 0.008952f
C4923 vdd.n3332 gnd 0.008952f
C4924 vdd.n3333 gnd 0.008952f
C4925 vdd.n3334 gnd 0.015419f
C4926 vdd.n3335 gnd 0.004899f
C4927 vdd.n3336 gnd 0.007205f
C4928 vdd.n3337 gnd 0.008952f
C4929 vdd.n3339 gnd 0.008952f
C4930 vdd.n3340 gnd 0.008952f
C4931 vdd.n3341 gnd 0.007205f
C4932 vdd.n3342 gnd 0.007205f
C4933 vdd.n3343 gnd 0.007205f
C4934 vdd.n3344 gnd 0.008952f
C4935 vdd.n3346 gnd 0.008952f
C4936 vdd.n3347 gnd 0.008952f
C4937 vdd.n3348 gnd 0.007205f
C4938 vdd.n3349 gnd 0.007205f
C4939 vdd.n3350 gnd 0.007205f
C4940 vdd.n3351 gnd 0.008952f
C4941 vdd.n3353 gnd 0.008952f
C4942 vdd.n3354 gnd 0.008952f
C4943 vdd.n3355 gnd 0.007205f
C4944 vdd.n3356 gnd 0.007205f
C4945 vdd.n3357 gnd 0.007205f
C4946 vdd.n3358 gnd 0.008952f
C4947 vdd.n3360 gnd 0.008952f
C4948 vdd.n3361 gnd 0.008952f
C4949 vdd.n3362 gnd 0.007205f
C4950 vdd.n3363 gnd 0.007205f
C4951 vdd.n3364 gnd 0.007205f
C4952 vdd.n3365 gnd 0.008952f
C4953 vdd.n3367 gnd 0.008952f
C4954 vdd.n3368 gnd 0.008952f
C4955 vdd.n3369 gnd 0.007205f
C4956 vdd.n3370 gnd 0.008952f
C4957 vdd.n3371 gnd 0.008952f
C4958 vdd.n3372 gnd 0.008952f
C4959 vdd.n3373 gnd 0.015419f
C4960 vdd.n3374 gnd 0.006016f
C4961 vdd.n3375 gnd 0.007205f
C4962 vdd.n3376 gnd 0.008952f
C4963 vdd.n3378 gnd 0.008952f
C4964 vdd.n3379 gnd 0.008952f
C4965 vdd.n3380 gnd 0.007205f
C4966 vdd.n3381 gnd 0.007205f
C4967 vdd.n3382 gnd 0.007205f
C4968 vdd.n3383 gnd 0.008952f
C4969 vdd.n3385 gnd 0.008952f
C4970 vdd.n3386 gnd 0.008952f
C4971 vdd.n3387 gnd 0.007205f
C4972 vdd.n3388 gnd 0.007205f
C4973 vdd.n3389 gnd 0.007205f
C4974 vdd.n3390 gnd 0.008952f
C4975 vdd.n3392 gnd 0.008952f
C4976 vdd.n3393 gnd 0.008952f
C4977 vdd.n3394 gnd 0.007205f
C4978 vdd.n3395 gnd 0.007205f
C4979 vdd.n3396 gnd 0.007205f
C4980 vdd.n3397 gnd 0.008952f
C4981 vdd.n3399 gnd 0.008952f
C4982 vdd.n3400 gnd 0.008952f
C4983 vdd.n3402 gnd 0.008952f
C4984 vdd.n3403 gnd 0.007205f
C4985 vdd.n3404 gnd 0.007205f
C4986 vdd.n3405 gnd 0.00598f
C4987 vdd.n3406 gnd 0.021425f
C4988 vdd.n3407 gnd 0.021096f
C4989 vdd.n3408 gnd 0.00598f
C4990 vdd.n3409 gnd 0.021096f
C4991 vdd.n3410 gnd 1.2899f
C4992 vdd.n3411 gnd 0.516873f
C4993 vdd.t33 gnd 0.45741f
C4994 vdd.n3412 gnd 0.855357f
C4995 vdd.n3413 gnd 0.008952f
C4996 vdd.n3414 gnd 0.007205f
C4997 vdd.n3415 gnd 0.007205f
C4998 vdd.n3416 gnd 0.007205f
C4999 vdd.n3417 gnd 0.008952f
C5000 vdd.n3418 gnd 0.901098f
C5001 vdd.t117 gnd 0.45741f
C5002 vdd.n3419 gnd 0.471132f
C5003 vdd.n3420 gnd 0.745578f
C5004 vdd.n3421 gnd 0.008952f
C5005 vdd.n3422 gnd 0.007205f
C5006 vdd.n3423 gnd 0.007205f
C5007 vdd.n3424 gnd 0.007205f
C5008 vdd.n3425 gnd 0.008952f
C5009 vdd.n3426 gnd 0.590059f
C5010 vdd.t98 gnd 0.45741f
C5011 vdd.n3427 gnd 0.759301f
C5012 vdd.t6 gnd 0.45741f
C5013 vdd.n3428 gnd 0.480281f
C5014 vdd.n3429 gnd 0.008952f
C5015 vdd.n3430 gnd 0.007205f
C5016 vdd.n3431 gnd 0.007205f
C5017 vdd.n3432 gnd 0.007205f
C5018 vdd.n3433 gnd 0.008952f
C5019 vdd.n3434 gnd 0.6358f
C5020 vdd.n3435 gnd 0.580911f
C5021 vdd.t88 gnd 0.45741f
C5022 vdd.n3436 gnd 0.759301f
C5023 vdd.n3437 gnd 0.008952f
C5024 vdd.n3438 gnd 0.007205f
C5025 vdd.n3439 gnd 0.532874f
C5026 vdd.n3440 gnd 2.2976f
C5027 a_n2982_13878.n0 gnd 0.930299f
C5028 a_n2982_13878.n1 gnd 0.204505f
C5029 a_n2982_13878.n2 gnd 0.150622f
C5030 a_n2982_13878.n3 gnd 0.23673f
C5031 a_n2982_13878.n4 gnd 0.182847f
C5032 a_n2982_13878.n5 gnd 0.204505f
C5033 a_n2982_13878.n6 gnd 0.150622f
C5034 a_n2982_13878.n7 gnd 0.984182f
C5035 a_n2982_13878.n8 gnd 0.215533f
C5036 a_n2982_13878.n9 gnd 0.758602f
C5037 a_n2982_13878.n10 gnd 0.215533f
C5038 a_n2982_13878.n11 gnd 0.215533f
C5039 a_n2982_13878.n12 gnd 0.490874f
C5040 a_n2982_13878.n13 gnd 0.282596f
C5041 a_n2982_13878.n14 gnd 0.215533f
C5042 a_n2982_13878.n15 gnd 0.544757f
C5043 a_n2982_13878.n16 gnd 0.215533f
C5044 a_n2982_13878.n17 gnd 0.215533f
C5045 a_n2982_13878.n18 gnd 0.958966f
C5046 a_n2982_13878.n19 gnd 0.282596f
C5047 a_n2982_13878.n20 gnd 3.20753f
C5048 a_n2982_13878.n21 gnd 0.215533f
C5049 a_n2982_13878.n22 gnd 0.215533f
C5050 a_n2982_13878.n23 gnd 0.868451f
C5051 a_n2982_13878.n24 gnd 0.215533f
C5052 a_n2982_13878.n25 gnd 0.282596f
C5053 a_n2982_13878.n26 gnd 1.00004f
C5054 a_n2982_13878.n27 gnd 0.215533f
C5055 a_n2982_13878.n28 gnd 0.215533f
C5056 a_n2982_13878.n29 gnd 0.490874f
C5057 a_n2982_13878.n30 gnd 0.215533f
C5058 a_n2982_13878.n31 gnd 0.282596f
C5059 a_n2982_13878.n32 gnd 3.4865f
C5060 a_n2982_13878.n33 gnd 2.65557f
C5061 a_n2982_13878.n34 gnd 3.74061f
C5062 a_n2982_13878.n35 gnd 1.19566f
C5063 a_n2982_13878.n36 gnd 2.1833f
C5064 a_n2982_13878.n37 gnd 1.77446f
C5065 a_n2982_13878.n38 gnd 1.19566f
C5066 a_n2982_13878.n39 gnd 1.77446f
C5067 a_n2982_13878.n40 gnd 2.38801f
C5068 a_n2982_13878.n41 gnd 0.725631f
C5069 a_n2982_13878.n42 gnd 0.725634f
C5070 a_n2982_13878.n43 gnd 0.008648f
C5071 a_n2982_13878.n44 gnd 4.17e-19
C5072 a_n2982_13878.n46 gnd 0.008345f
C5073 a_n2982_13878.n47 gnd 0.012134f
C5074 a_n2982_13878.n48 gnd 0.008028f
C5075 a_n2982_13878.n50 gnd 1.69354f
C5076 a_n2982_13878.n51 gnd 0.285885f
C5077 a_n2982_13878.n52 gnd 0.008648f
C5078 a_n2982_13878.n53 gnd 4.17e-19
C5079 a_n2982_13878.n55 gnd 0.008345f
C5080 a_n2982_13878.n56 gnd 0.012134f
C5081 a_n2982_13878.n57 gnd 0.008028f
C5082 a_n2982_13878.n59 gnd 0.008648f
C5083 a_n2982_13878.n60 gnd 4.17e-19
C5084 a_n2982_13878.n62 gnd 0.008345f
C5085 a_n2982_13878.n63 gnd 0.012134f
C5086 a_n2982_13878.n64 gnd 0.008028f
C5087 a_n2982_13878.n66 gnd 0.285885f
C5088 a_n2982_13878.n67 gnd 0.008648f
C5089 a_n2982_13878.n68 gnd 4.17e-19
C5090 a_n2982_13878.n70 gnd 0.008345f
C5091 a_n2982_13878.n71 gnd 0.012134f
C5092 a_n2982_13878.n72 gnd 0.008028f
C5093 a_n2982_13878.n74 gnd 0.285885f
C5094 a_n2982_13878.n75 gnd 0.008345f
C5095 a_n2982_13878.n76 gnd 0.284719f
C5096 a_n2982_13878.n77 gnd 0.008345f
C5097 a_n2982_13878.n78 gnd 0.284719f
C5098 a_n2982_13878.n79 gnd 0.008345f
C5099 a_n2982_13878.n80 gnd 0.284719f
C5100 a_n2982_13878.n81 gnd 0.008345f
C5101 a_n2982_13878.n82 gnd 0.284719f
C5102 a_n2982_13878.n83 gnd 0.285885f
C5103 a_n2982_13878.t45 gnd 0.149496f
C5104 a_n2982_13878.t35 gnd 1.39981f
C5105 a_n2982_13878.t63 gnd 0.149496f
C5106 a_n2982_13878.t25 gnd 0.149496f
C5107 a_n2982_13878.n84 gnd 1.05305f
C5108 a_n2982_13878.t26 gnd 0.695384f
C5109 a_n2982_13878.n85 gnd 0.305719f
C5110 a_n2982_13878.t60 gnd 0.695384f
C5111 a_n2982_13878.t46 gnd 0.695384f
C5112 a_n2982_13878.n86 gnd 0.296537f
C5113 a_n2982_13878.t22 gnd 0.695384f
C5114 a_n2982_13878.n87 gnd 0.308347f
C5115 a_n2982_13878.t58 gnd 0.695384f
C5116 a_n2982_13878.t24 gnd 0.695384f
C5117 a_n2982_13878.n88 gnd 0.30152f
C5118 a_n2982_13878.t34 gnd 0.70986f
C5119 a_n2982_13878.t86 gnd 0.695384f
C5120 a_n2982_13878.n89 gnd 0.305719f
C5121 a_n2982_13878.t96 gnd 0.695384f
C5122 a_n2982_13878.t101 gnd 0.695384f
C5123 a_n2982_13878.n90 gnd 0.296537f
C5124 a_n2982_13878.t105 gnd 0.695384f
C5125 a_n2982_13878.n91 gnd 0.308347f
C5126 a_n2982_13878.t76 gnd 0.695384f
C5127 a_n2982_13878.t79 gnd 0.695384f
C5128 a_n2982_13878.n92 gnd 0.30152f
C5129 a_n2982_13878.t109 gnd 0.70986f
C5130 a_n2982_13878.t40 gnd 0.70986f
C5131 a_n2982_13878.t52 gnd 0.695384f
C5132 a_n2982_13878.t30 gnd 0.695384f
C5133 a_n2982_13878.t64 gnd 0.695384f
C5134 a_n2982_13878.n93 gnd 0.305597f
C5135 a_n2982_13878.t38 gnd 0.695384f
C5136 a_n2982_13878.t54 gnd 0.695384f
C5137 a_n2982_13878.t32 gnd 0.695384f
C5138 a_n2982_13878.n94 gnd 0.301852f
C5139 a_n2982_13878.t48 gnd 0.695384f
C5140 a_n2982_13878.t56 gnd 0.695384f
C5141 a_n2982_13878.t50 gnd 0.695384f
C5142 a_n2982_13878.n95 gnd 0.305719f
C5143 a_n2982_13878.t66 gnd 0.695384f
C5144 a_n2982_13878.t42 gnd 0.70657f
C5145 a_n2982_13878.t17 gnd 0.116275f
C5146 a_n2982_13878.t9 gnd 0.116275f
C5147 a_n2982_13878.n96 gnd 1.02908f
C5148 a_n2982_13878.t3 gnd 0.116275f
C5149 a_n2982_13878.t11 gnd 0.116275f
C5150 a_n2982_13878.n97 gnd 1.02744f
C5151 a_n2982_13878.t16 gnd 0.116275f
C5152 a_n2982_13878.t15 gnd 0.116275f
C5153 a_n2982_13878.n98 gnd 1.02744f
C5154 a_n2982_13878.t1 gnd 0.116275f
C5155 a_n2982_13878.t18 gnd 0.116275f
C5156 a_n2982_13878.n99 gnd 1.02908f
C5157 a_n2982_13878.t2 gnd 0.116275f
C5158 a_n2982_13878.t12 gnd 0.116275f
C5159 a_n2982_13878.n100 gnd 1.02744f
C5160 a_n2982_13878.t6 gnd 0.116275f
C5161 a_n2982_13878.t5 gnd 0.116275f
C5162 a_n2982_13878.n101 gnd 1.02744f
C5163 a_n2982_13878.t13 gnd 0.116275f
C5164 a_n2982_13878.t70 gnd 0.116275f
C5165 a_n2982_13878.n102 gnd 1.02744f
C5166 a_n2982_13878.t0 gnd 0.116275f
C5167 a_n2982_13878.t21 gnd 0.116275f
C5168 a_n2982_13878.n103 gnd 1.02744f
C5169 a_n2982_13878.t19 gnd 0.116275f
C5170 a_n2982_13878.t7 gnd 0.116275f
C5171 a_n2982_13878.n104 gnd 1.02744f
C5172 a_n2982_13878.t20 gnd 0.116275f
C5173 a_n2982_13878.t10 gnd 0.116275f
C5174 a_n2982_13878.n105 gnd 1.02908f
C5175 a_n2982_13878.t8 gnd 0.116275f
C5176 a_n2982_13878.t14 gnd 0.116275f
C5177 a_n2982_13878.n106 gnd 1.02744f
C5178 a_n2982_13878.t4 gnd 0.116275f
C5179 a_n2982_13878.t71 gnd 0.116275f
C5180 a_n2982_13878.n107 gnd 1.02744f
C5181 a_n2982_13878.t110 gnd 0.70986f
C5182 a_n2982_13878.t87 gnd 0.695384f
C5183 a_n2982_13878.t92 gnd 0.695384f
C5184 a_n2982_13878.t80 gnd 0.695384f
C5185 a_n2982_13878.n108 gnd 0.305597f
C5186 a_n2982_13878.t97 gnd 0.695384f
C5187 a_n2982_13878.t106 gnd 0.695384f
C5188 a_n2982_13878.t107 gnd 0.695384f
C5189 a_n2982_13878.n109 gnd 0.301852f
C5190 a_n2982_13878.t74 gnd 0.695384f
C5191 a_n2982_13878.t89 gnd 0.695384f
C5192 a_n2982_13878.t77 gnd 0.695384f
C5193 a_n2982_13878.n110 gnd 0.305719f
C5194 a_n2982_13878.t84 gnd 0.695384f
C5195 a_n2982_13878.t103 gnd 0.70657f
C5196 a_n2982_13878.n111 gnd 0.307896f
C5197 a_n2982_13878.n112 gnd 0.302112f
C5198 a_n2982_13878.n113 gnd 0.296537f
C5199 a_n2982_13878.n114 gnd 0.305735f
C5200 a_n2982_13878.n115 gnd 0.308347f
C5201 a_n2982_13878.n116 gnd 0.30152f
C5202 a_n2982_13878.n117 gnd 0.307896f
C5203 a_n2982_13878.n118 gnd 0.307896f
C5204 a_n2982_13878.n119 gnd 0.302112f
C5205 a_n2982_13878.n120 gnd 0.296537f
C5206 a_n2982_13878.n121 gnd 0.305735f
C5207 a_n2982_13878.n122 gnd 0.308347f
C5208 a_n2982_13878.n123 gnd 0.30152f
C5209 a_n2982_13878.n124 gnd 0.307896f
C5210 a_n2982_13878.t43 gnd 1.39981f
C5211 a_n2982_13878.t51 gnd 0.149496f
C5212 a_n2982_13878.t67 gnd 0.149496f
C5213 a_n2982_13878.n125 gnd 1.05305f
C5214 a_n2982_13878.t49 gnd 0.149496f
C5215 a_n2982_13878.t57 gnd 0.149496f
C5216 a_n2982_13878.n126 gnd 1.05305f
C5217 a_n2982_13878.t55 gnd 0.149496f
C5218 a_n2982_13878.t33 gnd 0.149496f
C5219 a_n2982_13878.n127 gnd 1.05305f
C5220 a_n2982_13878.t65 gnd 0.149496f
C5221 a_n2982_13878.t39 gnd 0.149496f
C5222 a_n2982_13878.n128 gnd 1.05305f
C5223 a_n2982_13878.t53 gnd 0.149496f
C5224 a_n2982_13878.t31 gnd 0.149496f
C5225 a_n2982_13878.n129 gnd 1.05305f
C5226 a_n2982_13878.t41 gnd 1.39702f
C5227 a_n2982_13878.n130 gnd 1.0237f
C5228 a_n2982_13878.t85 gnd 0.695384f
C5229 a_n2982_13878.t95 gnd 0.695384f
C5230 a_n2982_13878.t111 gnd 0.695384f
C5231 a_n2982_13878.n131 gnd 0.305735f
C5232 a_n2982_13878.t98 gnd 0.695384f
C5233 a_n2982_13878.t81 gnd 0.695384f
C5234 a_n2982_13878.t82 gnd 0.695384f
C5235 a_n2982_13878.n132 gnd 0.305735f
C5236 a_n2982_13878.t102 gnd 0.695384f
C5237 a_n2982_13878.t91 gnd 0.695384f
C5238 a_n2982_13878.t90 gnd 0.695384f
C5239 a_n2982_13878.n133 gnd 0.305735f
C5240 a_n2982_13878.t94 gnd 0.695384f
C5241 a_n2982_13878.t83 gnd 0.695384f
C5242 a_n2982_13878.t72 gnd 0.695384f
C5243 a_n2982_13878.n134 gnd 0.305735f
C5244 a_n2982_13878.t99 gnd 0.707035f
C5245 a_n2982_13878.n135 gnd 0.301852f
C5246 a_n2982_13878.n136 gnd 0.296371f
C5247 a_n2982_13878.t108 gnd 0.707035f
C5248 a_n2982_13878.n137 gnd 0.301852f
C5249 a_n2982_13878.n138 gnd 0.296371f
C5250 a_n2982_13878.t93 gnd 0.707035f
C5251 a_n2982_13878.n139 gnd 0.301852f
C5252 a_n2982_13878.n140 gnd 0.296371f
C5253 a_n2982_13878.t88 gnd 0.707035f
C5254 a_n2982_13878.n141 gnd 0.301852f
C5255 a_n2982_13878.n142 gnd 0.296371f
C5256 a_n2982_13878.n143 gnd 1.36231f
C5257 a_n2982_13878.t78 gnd 0.695384f
C5258 a_n2982_13878.n144 gnd 0.307896f
C5259 a_n2982_13878.t104 gnd 0.695384f
C5260 a_n2982_13878.n145 gnd 0.305597f
C5261 a_n2982_13878.n146 gnd 0.305735f
C5262 a_n2982_13878.t100 gnd 0.695384f
C5263 a_n2982_13878.n147 gnd 0.301852f
C5264 a_n2982_13878.t73 gnd 0.695384f
C5265 a_n2982_13878.n148 gnd 0.302112f
C5266 a_n2982_13878.n149 gnd 0.307896f
C5267 a_n2982_13878.t75 gnd 0.70657f
C5268 a_n2982_13878.t62 gnd 0.695384f
C5269 a_n2982_13878.n150 gnd 0.307896f
C5270 a_n2982_13878.t44 gnd 0.695384f
C5271 a_n2982_13878.n151 gnd 0.305597f
C5272 a_n2982_13878.n152 gnd 0.305735f
C5273 a_n2982_13878.t36 gnd 0.695384f
C5274 a_n2982_13878.n153 gnd 0.301852f
C5275 a_n2982_13878.t28 gnd 0.695384f
C5276 a_n2982_13878.n154 gnd 0.302112f
C5277 a_n2982_13878.n155 gnd 0.307896f
C5278 a_n2982_13878.t68 gnd 0.70657f
C5279 a_n2982_13878.n156 gnd 1.34634f
C5280 a_n2982_13878.t69 gnd 1.39701f
C5281 a_n2982_13878.t27 gnd 0.149496f
C5282 a_n2982_13878.t61 gnd 0.149496f
C5283 a_n2982_13878.n157 gnd 1.05305f
C5284 a_n2982_13878.t47 gnd 0.149496f
C5285 a_n2982_13878.t29 gnd 0.149496f
C5286 a_n2982_13878.n158 gnd 1.05305f
C5287 a_n2982_13878.t59 gnd 0.149496f
C5288 a_n2982_13878.t37 gnd 0.149496f
C5289 a_n2982_13878.n159 gnd 1.05305f
C5290 a_n2982_13878.n160 gnd 1.05305f
C5291 a_n2982_13878.t23 gnd 0.149496f
C5292 commonsourceibias.n0 gnd 0.012299f
C5293 commonsourceibias.t57 gnd 0.18623f
C5294 commonsourceibias.t110 gnd 0.172196f
C5295 commonsourceibias.n1 gnd 0.068706f
C5296 commonsourceibias.n2 gnd 0.009217f
C5297 commonsourceibias.t70 gnd 0.172196f
C5298 commonsourceibias.n3 gnd 0.007456f
C5299 commonsourceibias.n4 gnd 0.009217f
C5300 commonsourceibias.t117 gnd 0.172196f
C5301 commonsourceibias.n5 gnd 0.008898f
C5302 commonsourceibias.n6 gnd 0.009217f
C5303 commonsourceibias.t85 gnd 0.172196f
C5304 commonsourceibias.n7 gnd 0.068706f
C5305 commonsourceibias.t54 gnd 0.172196f
C5306 commonsourceibias.n8 gnd 0.007444f
C5307 commonsourceibias.n9 gnd 0.012299f
C5308 commonsourceibias.t2 gnd 0.18623f
C5309 commonsourceibias.t42 gnd 0.172196f
C5310 commonsourceibias.n10 gnd 0.068706f
C5311 commonsourceibias.n11 gnd 0.009217f
C5312 commonsourceibias.t44 gnd 0.172196f
C5313 commonsourceibias.n12 gnd 0.007456f
C5314 commonsourceibias.n13 gnd 0.009217f
C5315 commonsourceibias.t32 gnd 0.172196f
C5316 commonsourceibias.n14 gnd 0.008898f
C5317 commonsourceibias.n15 gnd 0.009217f
C5318 commonsourceibias.t24 gnd 0.172196f
C5319 commonsourceibias.n16 gnd 0.068706f
C5320 commonsourceibias.t4 gnd 0.172196f
C5321 commonsourceibias.n17 gnd 0.007444f
C5322 commonsourceibias.n18 gnd 0.009217f
C5323 commonsourceibias.t14 gnd 0.172196f
C5324 commonsourceibias.t22 gnd 0.172196f
C5325 commonsourceibias.n19 gnd 0.068706f
C5326 commonsourceibias.n20 gnd 0.009217f
C5327 commonsourceibias.t36 gnd 0.172196f
C5328 commonsourceibias.n21 gnd 0.068706f
C5329 commonsourceibias.n22 gnd 0.009217f
C5330 commonsourceibias.t26 gnd 0.172196f
C5331 commonsourceibias.n23 gnd 0.068706f
C5332 commonsourceibias.n24 gnd 0.046399f
C5333 commonsourceibias.t8 gnd 0.172196f
C5334 commonsourceibias.t16 gnd 0.194303f
C5335 commonsourceibias.n25 gnd 0.079733f
C5336 commonsourceibias.n26 gnd 0.082545f
C5337 commonsourceibias.n27 gnd 0.01136f
C5338 commonsourceibias.n28 gnd 0.012567f
C5339 commonsourceibias.n29 gnd 0.009217f
C5340 commonsourceibias.n30 gnd 0.009217f
C5341 commonsourceibias.n31 gnd 0.012485f
C5342 commonsourceibias.n32 gnd 0.007456f
C5343 commonsourceibias.n33 gnd 0.01264f
C5344 commonsourceibias.n34 gnd 0.009217f
C5345 commonsourceibias.n35 gnd 0.009217f
C5346 commonsourceibias.n36 gnd 0.012717f
C5347 commonsourceibias.n37 gnd 0.010966f
C5348 commonsourceibias.n38 gnd 0.008898f
C5349 commonsourceibias.n39 gnd 0.009217f
C5350 commonsourceibias.n40 gnd 0.009217f
C5351 commonsourceibias.n41 gnd 0.011274f
C5352 commonsourceibias.n42 gnd 0.012653f
C5353 commonsourceibias.n43 gnd 0.068706f
C5354 commonsourceibias.n44 gnd 0.012568f
C5355 commonsourceibias.n45 gnd 0.009217f
C5356 commonsourceibias.n46 gnd 0.009217f
C5357 commonsourceibias.n47 gnd 0.009217f
C5358 commonsourceibias.n48 gnd 0.012568f
C5359 commonsourceibias.n49 gnd 0.068706f
C5360 commonsourceibias.n50 gnd 0.012653f
C5361 commonsourceibias.n51 gnd 0.011274f
C5362 commonsourceibias.n52 gnd 0.009217f
C5363 commonsourceibias.n53 gnd 0.009217f
C5364 commonsourceibias.n54 gnd 0.009217f
C5365 commonsourceibias.n55 gnd 0.010966f
C5366 commonsourceibias.n56 gnd 0.012717f
C5367 commonsourceibias.n57 gnd 0.068706f
C5368 commonsourceibias.n58 gnd 0.01264f
C5369 commonsourceibias.n59 gnd 0.009217f
C5370 commonsourceibias.n60 gnd 0.009217f
C5371 commonsourceibias.n61 gnd 0.009217f
C5372 commonsourceibias.n62 gnd 0.012485f
C5373 commonsourceibias.n63 gnd 0.068706f
C5374 commonsourceibias.n64 gnd 0.012567f
C5375 commonsourceibias.n65 gnd 0.01136f
C5376 commonsourceibias.n66 gnd 0.009217f
C5377 commonsourceibias.n67 gnd 0.009217f
C5378 commonsourceibias.n68 gnd 0.009349f
C5379 commonsourceibias.n69 gnd 0.009666f
C5380 commonsourceibias.n70 gnd 0.082208f
C5381 commonsourceibias.n71 gnd 0.091197f
C5382 commonsourceibias.t3 gnd 0.019889f
C5383 commonsourceibias.t43 gnd 0.019889f
C5384 commonsourceibias.n72 gnd 0.175743f
C5385 commonsourceibias.n73 gnd 0.151855f
C5386 commonsourceibias.t45 gnd 0.019889f
C5387 commonsourceibias.t33 gnd 0.019889f
C5388 commonsourceibias.n74 gnd 0.175743f
C5389 commonsourceibias.n75 gnd 0.080726f
C5390 commonsourceibias.t25 gnd 0.019889f
C5391 commonsourceibias.t5 gnd 0.019889f
C5392 commonsourceibias.n76 gnd 0.175743f
C5393 commonsourceibias.n77 gnd 0.067443f
C5394 commonsourceibias.t9 gnd 0.019889f
C5395 commonsourceibias.t17 gnd 0.019889f
C5396 commonsourceibias.n78 gnd 0.176331f
C5397 commonsourceibias.t37 gnd 0.019889f
C5398 commonsourceibias.t27 gnd 0.019889f
C5399 commonsourceibias.n79 gnd 0.175743f
C5400 commonsourceibias.n80 gnd 0.16376f
C5401 commonsourceibias.t15 gnd 0.019889f
C5402 commonsourceibias.t23 gnd 0.019889f
C5403 commonsourceibias.n81 gnd 0.175743f
C5404 commonsourceibias.n82 gnd 0.067443f
C5405 commonsourceibias.n83 gnd 0.081666f
C5406 commonsourceibias.n84 gnd 0.009217f
C5407 commonsourceibias.t97 gnd 0.172196f
C5408 commonsourceibias.t86 gnd 0.172196f
C5409 commonsourceibias.n85 gnd 0.068706f
C5410 commonsourceibias.n86 gnd 0.009217f
C5411 commonsourceibias.t115 gnd 0.172196f
C5412 commonsourceibias.n87 gnd 0.068706f
C5413 commonsourceibias.n88 gnd 0.009217f
C5414 commonsourceibias.t80 gnd 0.172196f
C5415 commonsourceibias.n89 gnd 0.068706f
C5416 commonsourceibias.n90 gnd 0.046399f
C5417 commonsourceibias.t66 gnd 0.172196f
C5418 commonsourceibias.t96 gnd 0.194303f
C5419 commonsourceibias.n91 gnd 0.079733f
C5420 commonsourceibias.n92 gnd 0.082545f
C5421 commonsourceibias.n93 gnd 0.01136f
C5422 commonsourceibias.n94 gnd 0.012567f
C5423 commonsourceibias.n95 gnd 0.009217f
C5424 commonsourceibias.n96 gnd 0.009217f
C5425 commonsourceibias.n97 gnd 0.012485f
C5426 commonsourceibias.n98 gnd 0.007456f
C5427 commonsourceibias.n99 gnd 0.01264f
C5428 commonsourceibias.n100 gnd 0.009217f
C5429 commonsourceibias.n101 gnd 0.009217f
C5430 commonsourceibias.n102 gnd 0.012717f
C5431 commonsourceibias.n103 gnd 0.010966f
C5432 commonsourceibias.n104 gnd 0.008898f
C5433 commonsourceibias.n105 gnd 0.009217f
C5434 commonsourceibias.n106 gnd 0.009217f
C5435 commonsourceibias.n107 gnd 0.011274f
C5436 commonsourceibias.n108 gnd 0.012653f
C5437 commonsourceibias.n109 gnd 0.068706f
C5438 commonsourceibias.n110 gnd 0.012568f
C5439 commonsourceibias.n111 gnd 0.009172f
C5440 commonsourceibias.n112 gnd 0.066626f
C5441 commonsourceibias.n113 gnd 0.009172f
C5442 commonsourceibias.n114 gnd 0.012568f
C5443 commonsourceibias.n115 gnd 0.068706f
C5444 commonsourceibias.n116 gnd 0.012653f
C5445 commonsourceibias.n117 gnd 0.011274f
C5446 commonsourceibias.n118 gnd 0.009217f
C5447 commonsourceibias.n119 gnd 0.009217f
C5448 commonsourceibias.n120 gnd 0.009217f
C5449 commonsourceibias.n121 gnd 0.010966f
C5450 commonsourceibias.n122 gnd 0.012717f
C5451 commonsourceibias.n123 gnd 0.068706f
C5452 commonsourceibias.n124 gnd 0.01264f
C5453 commonsourceibias.n125 gnd 0.009217f
C5454 commonsourceibias.n126 gnd 0.009217f
C5455 commonsourceibias.n127 gnd 0.009217f
C5456 commonsourceibias.n128 gnd 0.012485f
C5457 commonsourceibias.n129 gnd 0.068706f
C5458 commonsourceibias.n130 gnd 0.012567f
C5459 commonsourceibias.n131 gnd 0.01136f
C5460 commonsourceibias.n132 gnd 0.009217f
C5461 commonsourceibias.n133 gnd 0.009217f
C5462 commonsourceibias.n134 gnd 0.009349f
C5463 commonsourceibias.n135 gnd 0.009666f
C5464 commonsourceibias.n136 gnd 0.082208f
C5465 commonsourceibias.n137 gnd 0.05322f
C5466 commonsourceibias.n138 gnd 0.012299f
C5467 commonsourceibias.t88 gnd 0.18623f
C5468 commonsourceibias.t105 gnd 0.172196f
C5469 commonsourceibias.n139 gnd 0.068706f
C5470 commonsourceibias.n140 gnd 0.009217f
C5471 commonsourceibias.t101 gnd 0.172196f
C5472 commonsourceibias.n141 gnd 0.007456f
C5473 commonsourceibias.n142 gnd 0.009217f
C5474 commonsourceibias.t89 gnd 0.172196f
C5475 commonsourceibias.n143 gnd 0.008898f
C5476 commonsourceibias.n144 gnd 0.009217f
C5477 commonsourceibias.t106 gnd 0.172196f
C5478 commonsourceibias.n145 gnd 0.068706f
C5479 commonsourceibias.t99 gnd 0.172196f
C5480 commonsourceibias.n146 gnd 0.007444f
C5481 commonsourceibias.n147 gnd 0.009217f
C5482 commonsourceibias.t87 gnd 0.172196f
C5483 commonsourceibias.t107 gnd 0.172196f
C5484 commonsourceibias.n148 gnd 0.068706f
C5485 commonsourceibias.n149 gnd 0.009217f
C5486 commonsourceibias.t100 gnd 0.172196f
C5487 commonsourceibias.n150 gnd 0.068706f
C5488 commonsourceibias.n151 gnd 0.009217f
C5489 commonsourceibias.t112 gnd 0.172196f
C5490 commonsourceibias.n152 gnd 0.068706f
C5491 commonsourceibias.n153 gnd 0.046399f
C5492 commonsourceibias.t108 gnd 0.172196f
C5493 commonsourceibias.t98 gnd 0.194303f
C5494 commonsourceibias.n154 gnd 0.079733f
C5495 commonsourceibias.n155 gnd 0.082545f
C5496 commonsourceibias.n156 gnd 0.01136f
C5497 commonsourceibias.n157 gnd 0.012567f
C5498 commonsourceibias.n158 gnd 0.009217f
C5499 commonsourceibias.n159 gnd 0.009217f
C5500 commonsourceibias.n160 gnd 0.012485f
C5501 commonsourceibias.n161 gnd 0.007456f
C5502 commonsourceibias.n162 gnd 0.01264f
C5503 commonsourceibias.n163 gnd 0.009217f
C5504 commonsourceibias.n164 gnd 0.009217f
C5505 commonsourceibias.n165 gnd 0.012717f
C5506 commonsourceibias.n166 gnd 0.010966f
C5507 commonsourceibias.n167 gnd 0.008898f
C5508 commonsourceibias.n168 gnd 0.009217f
C5509 commonsourceibias.n169 gnd 0.009217f
C5510 commonsourceibias.n170 gnd 0.011274f
C5511 commonsourceibias.n171 gnd 0.012653f
C5512 commonsourceibias.n172 gnd 0.068706f
C5513 commonsourceibias.n173 gnd 0.012568f
C5514 commonsourceibias.n174 gnd 0.009217f
C5515 commonsourceibias.n175 gnd 0.009217f
C5516 commonsourceibias.n176 gnd 0.009217f
C5517 commonsourceibias.n177 gnd 0.012568f
C5518 commonsourceibias.n178 gnd 0.068706f
C5519 commonsourceibias.n179 gnd 0.012653f
C5520 commonsourceibias.n180 gnd 0.011274f
C5521 commonsourceibias.n181 gnd 0.009217f
C5522 commonsourceibias.n182 gnd 0.009217f
C5523 commonsourceibias.n183 gnd 0.009217f
C5524 commonsourceibias.n184 gnd 0.010966f
C5525 commonsourceibias.n185 gnd 0.012717f
C5526 commonsourceibias.n186 gnd 0.068706f
C5527 commonsourceibias.n187 gnd 0.01264f
C5528 commonsourceibias.n188 gnd 0.009217f
C5529 commonsourceibias.n189 gnd 0.009217f
C5530 commonsourceibias.n190 gnd 0.009217f
C5531 commonsourceibias.n191 gnd 0.012485f
C5532 commonsourceibias.n192 gnd 0.068706f
C5533 commonsourceibias.n193 gnd 0.012567f
C5534 commonsourceibias.n194 gnd 0.01136f
C5535 commonsourceibias.n195 gnd 0.009217f
C5536 commonsourceibias.n196 gnd 0.009217f
C5537 commonsourceibias.n197 gnd 0.009349f
C5538 commonsourceibias.n198 gnd 0.009666f
C5539 commonsourceibias.n199 gnd 0.082208f
C5540 commonsourceibias.n200 gnd 0.027976f
C5541 commonsourceibias.n201 gnd 0.147064f
C5542 commonsourceibias.n202 gnd 0.012299f
C5543 commonsourceibias.t50 gnd 0.172196f
C5544 commonsourceibias.n203 gnd 0.068706f
C5545 commonsourceibias.n204 gnd 0.009217f
C5546 commonsourceibias.t59 gnd 0.172196f
C5547 commonsourceibias.n205 gnd 0.007456f
C5548 commonsourceibias.n206 gnd 0.009217f
C5549 commonsourceibias.t104 gnd 0.172196f
C5550 commonsourceibias.n207 gnd 0.008898f
C5551 commonsourceibias.n208 gnd 0.009217f
C5552 commonsourceibias.t119 gnd 0.172196f
C5553 commonsourceibias.n209 gnd 0.068706f
C5554 commonsourceibias.t53 gnd 0.172196f
C5555 commonsourceibias.n210 gnd 0.007444f
C5556 commonsourceibias.n211 gnd 0.009217f
C5557 commonsourceibias.t93 gnd 0.172196f
C5558 commonsourceibias.t84 gnd 0.172196f
C5559 commonsourceibias.n212 gnd 0.068706f
C5560 commonsourceibias.n213 gnd 0.009217f
C5561 commonsourceibias.t49 gnd 0.172196f
C5562 commonsourceibias.n214 gnd 0.068706f
C5563 commonsourceibias.n215 gnd 0.009217f
C5564 commonsourceibias.t60 gnd 0.172196f
C5565 commonsourceibias.n216 gnd 0.068706f
C5566 commonsourceibias.n217 gnd 0.046399f
C5567 commonsourceibias.t75 gnd 0.172196f
C5568 commonsourceibias.t118 gnd 0.194303f
C5569 commonsourceibias.n218 gnd 0.079733f
C5570 commonsourceibias.n219 gnd 0.082545f
C5571 commonsourceibias.n220 gnd 0.01136f
C5572 commonsourceibias.n221 gnd 0.012567f
C5573 commonsourceibias.n222 gnd 0.009217f
C5574 commonsourceibias.n223 gnd 0.009217f
C5575 commonsourceibias.n224 gnd 0.012485f
C5576 commonsourceibias.n225 gnd 0.007456f
C5577 commonsourceibias.n226 gnd 0.01264f
C5578 commonsourceibias.n227 gnd 0.009217f
C5579 commonsourceibias.n228 gnd 0.009217f
C5580 commonsourceibias.n229 gnd 0.012717f
C5581 commonsourceibias.n230 gnd 0.010966f
C5582 commonsourceibias.n231 gnd 0.008898f
C5583 commonsourceibias.n232 gnd 0.009217f
C5584 commonsourceibias.n233 gnd 0.009217f
C5585 commonsourceibias.n234 gnd 0.011274f
C5586 commonsourceibias.n235 gnd 0.012653f
C5587 commonsourceibias.n236 gnd 0.068706f
C5588 commonsourceibias.n237 gnd 0.012568f
C5589 commonsourceibias.n238 gnd 0.009217f
C5590 commonsourceibias.n239 gnd 0.009217f
C5591 commonsourceibias.n240 gnd 0.009217f
C5592 commonsourceibias.n241 gnd 0.012568f
C5593 commonsourceibias.n242 gnd 0.068706f
C5594 commonsourceibias.n243 gnd 0.012653f
C5595 commonsourceibias.n244 gnd 0.011274f
C5596 commonsourceibias.n245 gnd 0.009217f
C5597 commonsourceibias.n246 gnd 0.009217f
C5598 commonsourceibias.n247 gnd 0.009217f
C5599 commonsourceibias.n248 gnd 0.010966f
C5600 commonsourceibias.n249 gnd 0.012717f
C5601 commonsourceibias.n250 gnd 0.068706f
C5602 commonsourceibias.n251 gnd 0.01264f
C5603 commonsourceibias.n252 gnd 0.009217f
C5604 commonsourceibias.n253 gnd 0.009217f
C5605 commonsourceibias.n254 gnd 0.009217f
C5606 commonsourceibias.n255 gnd 0.012485f
C5607 commonsourceibias.n256 gnd 0.068706f
C5608 commonsourceibias.n257 gnd 0.012567f
C5609 commonsourceibias.n258 gnd 0.01136f
C5610 commonsourceibias.n259 gnd 0.009217f
C5611 commonsourceibias.n260 gnd 0.009217f
C5612 commonsourceibias.n261 gnd 0.009349f
C5613 commonsourceibias.n262 gnd 0.009666f
C5614 commonsourceibias.t111 gnd 0.18623f
C5615 commonsourceibias.n263 gnd 0.082208f
C5616 commonsourceibias.n264 gnd 0.027976f
C5617 commonsourceibias.n265 gnd 0.517265f
C5618 commonsourceibias.n266 gnd 0.012299f
C5619 commonsourceibias.t114 gnd 0.18623f
C5620 commonsourceibias.t78 gnd 0.172196f
C5621 commonsourceibias.n267 gnd 0.068706f
C5622 commonsourceibias.n268 gnd 0.009217f
C5623 commonsourceibias.t52 gnd 0.172196f
C5624 commonsourceibias.n269 gnd 0.007456f
C5625 commonsourceibias.n270 gnd 0.009217f
C5626 commonsourceibias.t94 gnd 0.172196f
C5627 commonsourceibias.n271 gnd 0.008898f
C5628 commonsourceibias.n272 gnd 0.009217f
C5629 commonsourceibias.t113 gnd 0.172196f
C5630 commonsourceibias.n273 gnd 0.007444f
C5631 commonsourceibias.n274 gnd 0.009217f
C5632 commonsourceibias.t76 gnd 0.172196f
C5633 commonsourceibias.t65 gnd 0.172196f
C5634 commonsourceibias.n275 gnd 0.068706f
C5635 commonsourceibias.n276 gnd 0.009217f
C5636 commonsourceibias.t92 gnd 0.172196f
C5637 commonsourceibias.n277 gnd 0.068706f
C5638 commonsourceibias.n278 gnd 0.009217f
C5639 commonsourceibias.t63 gnd 0.172196f
C5640 commonsourceibias.n279 gnd 0.068706f
C5641 commonsourceibias.n280 gnd 0.046399f
C5642 commonsourceibias.t58 gnd 0.172196f
C5643 commonsourceibias.t69 gnd 0.194303f
C5644 commonsourceibias.n281 gnd 0.079733f
C5645 commonsourceibias.n282 gnd 0.082545f
C5646 commonsourceibias.n283 gnd 0.01136f
C5647 commonsourceibias.n284 gnd 0.012567f
C5648 commonsourceibias.n285 gnd 0.009217f
C5649 commonsourceibias.n286 gnd 0.009217f
C5650 commonsourceibias.n287 gnd 0.012485f
C5651 commonsourceibias.n288 gnd 0.007456f
C5652 commonsourceibias.n289 gnd 0.01264f
C5653 commonsourceibias.n290 gnd 0.009217f
C5654 commonsourceibias.n291 gnd 0.009217f
C5655 commonsourceibias.n292 gnd 0.012717f
C5656 commonsourceibias.n293 gnd 0.010966f
C5657 commonsourceibias.n294 gnd 0.008898f
C5658 commonsourceibias.n295 gnd 0.009217f
C5659 commonsourceibias.n296 gnd 0.009217f
C5660 commonsourceibias.n297 gnd 0.011274f
C5661 commonsourceibias.n298 gnd 0.012653f
C5662 commonsourceibias.n299 gnd 0.068706f
C5663 commonsourceibias.n300 gnd 0.012568f
C5664 commonsourceibias.n301 gnd 0.009172f
C5665 commonsourceibias.t47 gnd 0.019889f
C5666 commonsourceibias.t1 gnd 0.019889f
C5667 commonsourceibias.n302 gnd 0.176331f
C5668 commonsourceibias.t7 gnd 0.019889f
C5669 commonsourceibias.t21 gnd 0.019889f
C5670 commonsourceibias.n303 gnd 0.175743f
C5671 commonsourceibias.n304 gnd 0.16376f
C5672 commonsourceibias.t11 gnd 0.019889f
C5673 commonsourceibias.t35 gnd 0.019889f
C5674 commonsourceibias.n305 gnd 0.175743f
C5675 commonsourceibias.n306 gnd 0.067443f
C5676 commonsourceibias.n307 gnd 0.012299f
C5677 commonsourceibias.t28 gnd 0.172196f
C5678 commonsourceibias.n308 gnd 0.068706f
C5679 commonsourceibias.n309 gnd 0.009217f
C5680 commonsourceibias.t30 gnd 0.172196f
C5681 commonsourceibias.n310 gnd 0.007456f
C5682 commonsourceibias.n311 gnd 0.009217f
C5683 commonsourceibias.t18 gnd 0.172196f
C5684 commonsourceibias.n312 gnd 0.008898f
C5685 commonsourceibias.n313 gnd 0.009217f
C5686 commonsourceibias.t40 gnd 0.172196f
C5687 commonsourceibias.n314 gnd 0.007444f
C5688 commonsourceibias.n315 gnd 0.009217f
C5689 commonsourceibias.t34 gnd 0.172196f
C5690 commonsourceibias.t10 gnd 0.172196f
C5691 commonsourceibias.n316 gnd 0.068706f
C5692 commonsourceibias.n317 gnd 0.009217f
C5693 commonsourceibias.t20 gnd 0.172196f
C5694 commonsourceibias.n318 gnd 0.068706f
C5695 commonsourceibias.n319 gnd 0.009217f
C5696 commonsourceibias.t6 gnd 0.172196f
C5697 commonsourceibias.n320 gnd 0.068706f
C5698 commonsourceibias.n321 gnd 0.046399f
C5699 commonsourceibias.t0 gnd 0.172196f
C5700 commonsourceibias.t46 gnd 0.194303f
C5701 commonsourceibias.n322 gnd 0.079733f
C5702 commonsourceibias.n323 gnd 0.082545f
C5703 commonsourceibias.n324 gnd 0.01136f
C5704 commonsourceibias.n325 gnd 0.012567f
C5705 commonsourceibias.n326 gnd 0.009217f
C5706 commonsourceibias.n327 gnd 0.009217f
C5707 commonsourceibias.n328 gnd 0.012485f
C5708 commonsourceibias.n329 gnd 0.007456f
C5709 commonsourceibias.n330 gnd 0.01264f
C5710 commonsourceibias.n331 gnd 0.009217f
C5711 commonsourceibias.n332 gnd 0.009217f
C5712 commonsourceibias.n333 gnd 0.012717f
C5713 commonsourceibias.n334 gnd 0.010966f
C5714 commonsourceibias.n335 gnd 0.008898f
C5715 commonsourceibias.n336 gnd 0.009217f
C5716 commonsourceibias.n337 gnd 0.009217f
C5717 commonsourceibias.n338 gnd 0.011274f
C5718 commonsourceibias.n339 gnd 0.012653f
C5719 commonsourceibias.n340 gnd 0.068706f
C5720 commonsourceibias.n341 gnd 0.012568f
C5721 commonsourceibias.n342 gnd 0.009217f
C5722 commonsourceibias.n343 gnd 0.009217f
C5723 commonsourceibias.n344 gnd 0.009217f
C5724 commonsourceibias.n345 gnd 0.012568f
C5725 commonsourceibias.n346 gnd 0.068706f
C5726 commonsourceibias.n347 gnd 0.012653f
C5727 commonsourceibias.t12 gnd 0.172196f
C5728 commonsourceibias.n348 gnd 0.068706f
C5729 commonsourceibias.n349 gnd 0.011274f
C5730 commonsourceibias.n350 gnd 0.009217f
C5731 commonsourceibias.n351 gnd 0.009217f
C5732 commonsourceibias.n352 gnd 0.009217f
C5733 commonsourceibias.n353 gnd 0.010966f
C5734 commonsourceibias.n354 gnd 0.012717f
C5735 commonsourceibias.n355 gnd 0.068706f
C5736 commonsourceibias.n356 gnd 0.01264f
C5737 commonsourceibias.n357 gnd 0.009217f
C5738 commonsourceibias.n358 gnd 0.009217f
C5739 commonsourceibias.n359 gnd 0.009217f
C5740 commonsourceibias.n360 gnd 0.012485f
C5741 commonsourceibias.n361 gnd 0.068706f
C5742 commonsourceibias.n362 gnd 0.012567f
C5743 commonsourceibias.n363 gnd 0.01136f
C5744 commonsourceibias.n364 gnd 0.009217f
C5745 commonsourceibias.n365 gnd 0.009217f
C5746 commonsourceibias.n366 gnd 0.009349f
C5747 commonsourceibias.n367 gnd 0.009666f
C5748 commonsourceibias.t38 gnd 0.18623f
C5749 commonsourceibias.n368 gnd 0.082208f
C5750 commonsourceibias.n369 gnd 0.091197f
C5751 commonsourceibias.t29 gnd 0.019889f
C5752 commonsourceibias.t39 gnd 0.019889f
C5753 commonsourceibias.n370 gnd 0.175743f
C5754 commonsourceibias.n371 gnd 0.151855f
C5755 commonsourceibias.t19 gnd 0.019889f
C5756 commonsourceibias.t31 gnd 0.019889f
C5757 commonsourceibias.n372 gnd 0.175743f
C5758 commonsourceibias.n373 gnd 0.080726f
C5759 commonsourceibias.t41 gnd 0.019889f
C5760 commonsourceibias.t13 gnd 0.019889f
C5761 commonsourceibias.n374 gnd 0.175743f
C5762 commonsourceibias.n375 gnd 0.067443f
C5763 commonsourceibias.n376 gnd 0.081666f
C5764 commonsourceibias.n377 gnd 0.066626f
C5765 commonsourceibias.n378 gnd 0.009172f
C5766 commonsourceibias.n379 gnd 0.012568f
C5767 commonsourceibias.n380 gnd 0.068706f
C5768 commonsourceibias.n381 gnd 0.012653f
C5769 commonsourceibias.t64 gnd 0.172196f
C5770 commonsourceibias.n382 gnd 0.068706f
C5771 commonsourceibias.n383 gnd 0.011274f
C5772 commonsourceibias.n384 gnd 0.009217f
C5773 commonsourceibias.n385 gnd 0.009217f
C5774 commonsourceibias.n386 gnd 0.009217f
C5775 commonsourceibias.n387 gnd 0.010966f
C5776 commonsourceibias.n388 gnd 0.012717f
C5777 commonsourceibias.n389 gnd 0.068706f
C5778 commonsourceibias.n390 gnd 0.01264f
C5779 commonsourceibias.n391 gnd 0.009217f
C5780 commonsourceibias.n392 gnd 0.009217f
C5781 commonsourceibias.n393 gnd 0.009217f
C5782 commonsourceibias.n394 gnd 0.012485f
C5783 commonsourceibias.n395 gnd 0.068706f
C5784 commonsourceibias.n396 gnd 0.012567f
C5785 commonsourceibias.n397 gnd 0.01136f
C5786 commonsourceibias.n398 gnd 0.009217f
C5787 commonsourceibias.n399 gnd 0.009217f
C5788 commonsourceibias.n400 gnd 0.009349f
C5789 commonsourceibias.n401 gnd 0.009666f
C5790 commonsourceibias.n402 gnd 0.082208f
C5791 commonsourceibias.n403 gnd 0.05322f
C5792 commonsourceibias.n404 gnd 0.012299f
C5793 commonsourceibias.t91 gnd 0.172196f
C5794 commonsourceibias.n405 gnd 0.068706f
C5795 commonsourceibias.n406 gnd 0.009217f
C5796 commonsourceibias.t82 gnd 0.172196f
C5797 commonsourceibias.n407 gnd 0.007456f
C5798 commonsourceibias.n408 gnd 0.009217f
C5799 commonsourceibias.t73 gnd 0.172196f
C5800 commonsourceibias.n409 gnd 0.008898f
C5801 commonsourceibias.n410 gnd 0.009217f
C5802 commonsourceibias.t83 gnd 0.172196f
C5803 commonsourceibias.n411 gnd 0.007444f
C5804 commonsourceibias.n412 gnd 0.009217f
C5805 commonsourceibias.t103 gnd 0.172196f
C5806 commonsourceibias.t95 gnd 0.172196f
C5807 commonsourceibias.n413 gnd 0.068706f
C5808 commonsourceibias.n414 gnd 0.009217f
C5809 commonsourceibias.t81 gnd 0.172196f
C5810 commonsourceibias.n415 gnd 0.068706f
C5811 commonsourceibias.n416 gnd 0.009217f
C5812 commonsourceibias.t102 gnd 0.172196f
C5813 commonsourceibias.n417 gnd 0.068706f
C5814 commonsourceibias.n418 gnd 0.046399f
C5815 commonsourceibias.t116 gnd 0.172196f
C5816 commonsourceibias.t79 gnd 0.194303f
C5817 commonsourceibias.n419 gnd 0.079733f
C5818 commonsourceibias.n420 gnd 0.082545f
C5819 commonsourceibias.n421 gnd 0.01136f
C5820 commonsourceibias.n422 gnd 0.012567f
C5821 commonsourceibias.n423 gnd 0.009217f
C5822 commonsourceibias.n424 gnd 0.009217f
C5823 commonsourceibias.n425 gnd 0.012485f
C5824 commonsourceibias.n426 gnd 0.007456f
C5825 commonsourceibias.n427 gnd 0.01264f
C5826 commonsourceibias.n428 gnd 0.009217f
C5827 commonsourceibias.n429 gnd 0.009217f
C5828 commonsourceibias.n430 gnd 0.012717f
C5829 commonsourceibias.n431 gnd 0.010966f
C5830 commonsourceibias.n432 gnd 0.008898f
C5831 commonsourceibias.n433 gnd 0.009217f
C5832 commonsourceibias.n434 gnd 0.009217f
C5833 commonsourceibias.n435 gnd 0.011274f
C5834 commonsourceibias.n436 gnd 0.012653f
C5835 commonsourceibias.n437 gnd 0.068706f
C5836 commonsourceibias.n438 gnd 0.012568f
C5837 commonsourceibias.n439 gnd 0.009217f
C5838 commonsourceibias.n440 gnd 0.009217f
C5839 commonsourceibias.n441 gnd 0.009217f
C5840 commonsourceibias.n442 gnd 0.012568f
C5841 commonsourceibias.n443 gnd 0.068706f
C5842 commonsourceibias.n444 gnd 0.012653f
C5843 commonsourceibias.t90 gnd 0.172196f
C5844 commonsourceibias.n445 gnd 0.068706f
C5845 commonsourceibias.n446 gnd 0.011274f
C5846 commonsourceibias.n447 gnd 0.009217f
C5847 commonsourceibias.n448 gnd 0.009217f
C5848 commonsourceibias.n449 gnd 0.009217f
C5849 commonsourceibias.n450 gnd 0.010966f
C5850 commonsourceibias.n451 gnd 0.012717f
C5851 commonsourceibias.n452 gnd 0.068706f
C5852 commonsourceibias.n453 gnd 0.01264f
C5853 commonsourceibias.n454 gnd 0.009217f
C5854 commonsourceibias.n455 gnd 0.009217f
C5855 commonsourceibias.n456 gnd 0.009217f
C5856 commonsourceibias.n457 gnd 0.012485f
C5857 commonsourceibias.n458 gnd 0.068706f
C5858 commonsourceibias.n459 gnd 0.012567f
C5859 commonsourceibias.n460 gnd 0.01136f
C5860 commonsourceibias.n461 gnd 0.009217f
C5861 commonsourceibias.n462 gnd 0.009217f
C5862 commonsourceibias.n463 gnd 0.009349f
C5863 commonsourceibias.n464 gnd 0.009666f
C5864 commonsourceibias.t74 gnd 0.18623f
C5865 commonsourceibias.n465 gnd 0.082208f
C5866 commonsourceibias.n466 gnd 0.027976f
C5867 commonsourceibias.n467 gnd 0.147064f
C5868 commonsourceibias.n468 gnd 0.012299f
C5869 commonsourceibias.t62 gnd 0.172196f
C5870 commonsourceibias.n469 gnd 0.068706f
C5871 commonsourceibias.n470 gnd 0.009217f
C5872 commonsourceibias.t71 gnd 0.172196f
C5873 commonsourceibias.n471 gnd 0.007456f
C5874 commonsourceibias.n472 gnd 0.009217f
C5875 commonsourceibias.t48 gnd 0.172196f
C5876 commonsourceibias.n473 gnd 0.008898f
C5877 commonsourceibias.n474 gnd 0.009217f
C5878 commonsourceibias.t67 gnd 0.172196f
C5879 commonsourceibias.n475 gnd 0.007444f
C5880 commonsourceibias.n476 gnd 0.009217f
C5881 commonsourceibias.t77 gnd 0.172196f
C5882 commonsourceibias.t109 gnd 0.172196f
C5883 commonsourceibias.n477 gnd 0.068706f
C5884 commonsourceibias.n478 gnd 0.009217f
C5885 commonsourceibias.t61 gnd 0.172196f
C5886 commonsourceibias.n479 gnd 0.068706f
C5887 commonsourceibias.n480 gnd 0.009217f
C5888 commonsourceibias.t72 gnd 0.172196f
C5889 commonsourceibias.n481 gnd 0.068706f
C5890 commonsourceibias.n482 gnd 0.046399f
C5891 commonsourceibias.t68 gnd 0.172196f
C5892 commonsourceibias.t55 gnd 0.194303f
C5893 commonsourceibias.n483 gnd 0.079733f
C5894 commonsourceibias.n484 gnd 0.082545f
C5895 commonsourceibias.n485 gnd 0.01136f
C5896 commonsourceibias.n486 gnd 0.012567f
C5897 commonsourceibias.n487 gnd 0.009217f
C5898 commonsourceibias.n488 gnd 0.009217f
C5899 commonsourceibias.n489 gnd 0.012485f
C5900 commonsourceibias.n490 gnd 0.007456f
C5901 commonsourceibias.n491 gnd 0.01264f
C5902 commonsourceibias.n492 gnd 0.009217f
C5903 commonsourceibias.n493 gnd 0.009217f
C5904 commonsourceibias.n494 gnd 0.012717f
C5905 commonsourceibias.n495 gnd 0.010966f
C5906 commonsourceibias.n496 gnd 0.008898f
C5907 commonsourceibias.n497 gnd 0.009217f
C5908 commonsourceibias.n498 gnd 0.009217f
C5909 commonsourceibias.n499 gnd 0.011274f
C5910 commonsourceibias.n500 gnd 0.012653f
C5911 commonsourceibias.n501 gnd 0.068706f
C5912 commonsourceibias.n502 gnd 0.012568f
C5913 commonsourceibias.n503 gnd 0.009217f
C5914 commonsourceibias.n504 gnd 0.009217f
C5915 commonsourceibias.n505 gnd 0.009217f
C5916 commonsourceibias.n506 gnd 0.012568f
C5917 commonsourceibias.n507 gnd 0.068706f
C5918 commonsourceibias.n508 gnd 0.012653f
C5919 commonsourceibias.t56 gnd 0.172196f
C5920 commonsourceibias.n509 gnd 0.068706f
C5921 commonsourceibias.n510 gnd 0.011274f
C5922 commonsourceibias.n511 gnd 0.009217f
C5923 commonsourceibias.n512 gnd 0.009217f
C5924 commonsourceibias.n513 gnd 0.009217f
C5925 commonsourceibias.n514 gnd 0.010966f
C5926 commonsourceibias.n515 gnd 0.012717f
C5927 commonsourceibias.n516 gnd 0.068706f
C5928 commonsourceibias.n517 gnd 0.01264f
C5929 commonsourceibias.n518 gnd 0.009217f
C5930 commonsourceibias.n519 gnd 0.009217f
C5931 commonsourceibias.n520 gnd 0.009217f
C5932 commonsourceibias.n521 gnd 0.012485f
C5933 commonsourceibias.n522 gnd 0.068706f
C5934 commonsourceibias.n523 gnd 0.012567f
C5935 commonsourceibias.n524 gnd 0.01136f
C5936 commonsourceibias.n525 gnd 0.009217f
C5937 commonsourceibias.n526 gnd 0.009217f
C5938 commonsourceibias.n527 gnd 0.009349f
C5939 commonsourceibias.n528 gnd 0.009666f
C5940 commonsourceibias.t51 gnd 0.18623f
C5941 commonsourceibias.n529 gnd 0.082208f
C5942 commonsourceibias.n530 gnd 0.027976f
C5943 commonsourceibias.n531 gnd 0.194274f
C5944 commonsourceibias.n532 gnd 5.09694f
.ends

