* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t46 plus.t0 drain_left.t10 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X1 source.t22 minus.t0 drain_right.t23 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X2 drain_right.t22 minus.t1 source.t20 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X3 source.t45 plus.t1 drain_left.t5 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X4 drain_left.t16 plus.t2 source.t44 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X5 source.t7 minus.t2 drain_right.t21 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=1
X6 drain_left.t23 plus.t3 source.t43 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X7 a_n4174_n1488# a_n4174_n1488# a_n4174_n1488# a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=1
X8 drain_left.t14 plus.t4 source.t42 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X9 drain_left.t6 plus.t5 source.t41 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X10 drain_right.t20 minus.t3 source.t21 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X11 source.t19 minus.t4 drain_right.t19 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X12 drain_left.t20 plus.t6 source.t40 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X13 drain_left.t17 plus.t7 source.t39 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=1
X14 source.t38 plus.t8 drain_left.t12 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X15 source.t37 plus.t9 drain_left.t0 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X16 source.t36 plus.t10 drain_left.t13 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X17 drain_right.t18 minus.t5 source.t1 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X18 source.t6 minus.t6 drain_right.t17 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X19 drain_left.t15 plus.t11 source.t35 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X20 source.t34 plus.t12 drain_left.t8 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X21 drain_left.t1 plus.t13 source.t33 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X22 source.t32 plus.t14 drain_left.t11 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X23 drain_left.t2 plus.t15 source.t31 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=1
X24 source.t4 minus.t7 drain_right.t16 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X25 drain_right.t15 minus.t8 source.t5 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X26 source.t13 minus.t9 drain_right.t14 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X27 drain_left.t7 plus.t16 source.t30 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X28 source.t29 plus.t17 drain_left.t21 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X29 a_n4174_n1488# a_n4174_n1488# a_n4174_n1488# a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=1
X30 drain_right.t13 minus.t10 source.t10 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X31 drain_right.t12 minus.t11 source.t2 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X32 drain_right.t11 minus.t12 source.t12 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=1
X33 source.t16 minus.t13 drain_right.t10 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X34 drain_right.t9 minus.t14 source.t9 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=1
X35 source.t14 minus.t15 drain_right.t8 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X36 drain_left.t18 plus.t18 source.t28 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X37 source.t27 plus.t19 drain_left.t22 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X38 drain_right.t7 minus.t16 source.t18 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X39 drain_left.t19 plus.t20 source.t26 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X40 source.t25 plus.t21 drain_left.t4 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=1
X41 a_n4174_n1488# a_n4174_n1488# a_n4174_n1488# a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=1
X42 source.t11 minus.t17 drain_right.t6 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X43 drain_right.t5 minus.t18 source.t17 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X44 source.t24 plus.t22 drain_left.t9 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X45 source.t15 minus.t19 drain_right.t4 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X46 a_n4174_n1488# a_n4174_n1488# a_n4174_n1488# a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=1
X47 source.t23 plus.t23 drain_left.t3 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=1
X48 source.t47 minus.t20 drain_right.t3 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X49 drain_right.t2 minus.t21 source.t8 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X50 drain_right.t1 minus.t22 source.t3 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X51 source.t0 minus.t23 drain_right.t0 a_n4174_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=1
R0 plus.n17 plus.n14 161.3
R1 plus.n19 plus.n18 161.3
R2 plus.n21 plus.n20 161.3
R3 plus.n22 plus.n12 161.3
R4 plus.n24 plus.n23 161.3
R5 plus.n26 plus.n25 161.3
R6 plus.n27 plus.n10 161.3
R7 plus.n29 plus.n28 161.3
R8 plus.n31 plus.n30 161.3
R9 plus.n32 plus.n8 161.3
R10 plus.n35 plus.n34 161.3
R11 plus.n36 plus.n7 161.3
R12 plus.n38 plus.n37 161.3
R13 plus.n40 plus.n6 161.3
R14 plus.n43 plus.n42 161.3
R15 plus.n44 plus.n5 161.3
R16 plus.n46 plus.n45 161.3
R17 plus.n47 plus.n4 161.3
R18 plus.n50 plus.n49 161.3
R19 plus.n51 plus.n3 161.3
R20 plus.n53 plus.n52 161.3
R21 plus.n55 plus.n2 161.3
R22 plus.n57 plus.n56 161.3
R23 plus.n59 plus.n58 161.3
R24 plus.n60 plus.n0 161.3
R25 plus.n81 plus.n78 161.3
R26 plus.n83 plus.n82 161.3
R27 plus.n85 plus.n84 161.3
R28 plus.n86 plus.n76 161.3
R29 plus.n88 plus.n87 161.3
R30 plus.n90 plus.n89 161.3
R31 plus.n91 plus.n74 161.3
R32 plus.n93 plus.n92 161.3
R33 plus.n95 plus.n94 161.3
R34 plus.n96 plus.n72 161.3
R35 plus.n99 plus.n98 161.3
R36 plus.n100 plus.n71 161.3
R37 plus.n102 plus.n101 161.3
R38 plus.n104 plus.n69 161.3
R39 plus.n106 plus.n105 161.3
R40 plus.n107 plus.n68 161.3
R41 plus.n109 plus.n108 161.3
R42 plus.n110 plus.n67 161.3
R43 plus.n113 plus.n112 161.3
R44 plus.n114 plus.n66 161.3
R45 plus.n116 plus.n115 161.3
R46 plus.n118 plus.n65 161.3
R47 plus.n120 plus.n119 161.3
R48 plus.n122 plus.n121 161.3
R49 plus.n123 plus.n63 161.3
R50 plus.n15 plus.t23 133.606
R51 plus.n79 plus.t15 133.606
R52 plus.n61 plus.t7 111.584
R53 plus.n124 plus.t21 111.584
R54 plus.n62 plus.n61 80.6037
R55 plus.n125 plus.n124 80.6037
R56 plus.n1 plus.t12 72.3005
R57 plus.n54 plus.t16 72.3005
R58 plus.n48 plus.t8 72.3005
R59 plus.n41 plus.t13 72.3005
R60 plus.n39 plus.t17 72.3005
R61 plus.n33 plus.t6 72.3005
R62 plus.n9 plus.t14 72.3005
R63 plus.n11 plus.t3 72.3005
R64 plus.n13 plus.t0 72.3005
R65 plus.n16 plus.t2 72.3005
R66 plus.n64 plus.t11 72.3005
R67 plus.n117 plus.t1 72.3005
R68 plus.n111 plus.t5 72.3005
R69 plus.n70 plus.t19 72.3005
R70 plus.n103 plus.t4 72.3005
R71 plus.n97 plus.t10 72.3005
R72 plus.n73 plus.t20 72.3005
R73 plus.n75 plus.t22 72.3005
R74 plus.n77 plus.t18 72.3005
R75 plus.n80 plus.t9 72.3005
R76 plus.n56 plus.n55 56.5617
R77 plus.n42 plus.n40 56.5617
R78 plus.n32 plus.n31 56.5617
R79 plus.n18 plus.n17 56.5617
R80 plus.n119 plus.n118 56.5617
R81 plus.n105 plus.n104 56.5617
R82 plus.n96 plus.n95 56.5617
R83 plus.n82 plus.n81 56.5617
R84 plus.n47 plus.n46 56.0773
R85 plus.n27 plus.n26 56.0773
R86 plus.n110 plus.n109 56.0773
R87 plus.n91 plus.n90 56.0773
R88 plus.n61 plus.n60 46.0096
R89 plus.n124 plus.n123 46.0096
R90 plus.n49 plus.n3 41.5458
R91 plus.n23 plus.n22 41.5458
R92 plus.n112 plus.n66 41.5458
R93 plus.n87 plus.n86 41.5458
R94 plus.n38 plus.n7 40.577
R95 plus.n34 plus.n7 40.577
R96 plus.n102 plus.n71 40.577
R97 plus.n98 plus.n71 40.577
R98 plus.n53 plus.n3 39.6083
R99 plus.n22 plus.n21 39.6083
R100 plus.n116 plus.n66 39.6083
R101 plus.n86 plus.n85 39.6083
R102 plus plus.n125 35.7154
R103 plus.n16 plus.n15 33.0515
R104 plus.n80 plus.n79 33.0515
R105 plus.n15 plus.n14 28.5514
R106 plus.n79 plus.n78 28.5514
R107 plus.n60 plus.n59 26.0455
R108 plus.n123 plus.n122 26.0455
R109 plus.n46 plus.n5 25.0767
R110 plus.n28 plus.n27 25.0767
R111 plus.n109 plus.n68 25.0767
R112 plus.n92 plus.n91 25.0767
R113 plus.n42 plus.n41 24.3464
R114 plus.n31 plus.n9 24.3464
R115 plus.n105 plus.n70 24.3464
R116 plus.n95 plus.n73 24.3464
R117 plus.n56 plus.n1 23.8546
R118 plus.n17 plus.n16 23.8546
R119 plus.n119 plus.n64 23.8546
R120 plus.n81 plus.n80 23.8546
R121 plus.n55 plus.n54 16.9689
R122 plus.n18 plus.n13 16.9689
R123 plus.n118 plus.n117 16.9689
R124 plus.n82 plus.n77 16.9689
R125 plus.n40 plus.n39 16.477
R126 plus.n33 plus.n32 16.477
R127 plus.n104 plus.n103 16.477
R128 plus.n97 plus.n96 16.477
R129 plus.n48 plus.n47 15.9852
R130 plus.n26 plus.n11 15.9852
R131 plus.n111 plus.n110 15.9852
R132 plus.n90 plus.n75 15.9852
R133 plus plus.n62 9.0464
R134 plus.n49 plus.n48 8.60764
R135 plus.n23 plus.n11 8.60764
R136 plus.n112 plus.n111 8.60764
R137 plus.n87 plus.n75 8.60764
R138 plus.n39 plus.n38 8.11581
R139 plus.n34 plus.n33 8.11581
R140 plus.n103 plus.n102 8.11581
R141 plus.n98 plus.n97 8.11581
R142 plus.n54 plus.n53 7.62397
R143 plus.n21 plus.n13 7.62397
R144 plus.n117 plus.n116 7.62397
R145 plus.n85 plus.n77 7.62397
R146 plus.n59 plus.n1 0.738255
R147 plus.n122 plus.n64 0.738255
R148 plus.n62 plus.n0 0.285035
R149 plus.n125 plus.n63 0.285035
R150 plus.n41 plus.n5 0.246418
R151 plus.n28 plus.n9 0.246418
R152 plus.n70 plus.n68 0.246418
R153 plus.n92 plus.n73 0.246418
R154 plus.n19 plus.n14 0.189894
R155 plus.n20 plus.n19 0.189894
R156 plus.n20 plus.n12 0.189894
R157 plus.n24 plus.n12 0.189894
R158 plus.n25 plus.n24 0.189894
R159 plus.n25 plus.n10 0.189894
R160 plus.n29 plus.n10 0.189894
R161 plus.n30 plus.n29 0.189894
R162 plus.n30 plus.n8 0.189894
R163 plus.n35 plus.n8 0.189894
R164 plus.n36 plus.n35 0.189894
R165 plus.n37 plus.n36 0.189894
R166 plus.n37 plus.n6 0.189894
R167 plus.n43 plus.n6 0.189894
R168 plus.n44 plus.n43 0.189894
R169 plus.n45 plus.n44 0.189894
R170 plus.n45 plus.n4 0.189894
R171 plus.n50 plus.n4 0.189894
R172 plus.n51 plus.n50 0.189894
R173 plus.n52 plus.n51 0.189894
R174 plus.n52 plus.n2 0.189894
R175 plus.n57 plus.n2 0.189894
R176 plus.n58 plus.n57 0.189894
R177 plus.n58 plus.n0 0.189894
R178 plus.n121 plus.n63 0.189894
R179 plus.n121 plus.n120 0.189894
R180 plus.n120 plus.n65 0.189894
R181 plus.n115 plus.n65 0.189894
R182 plus.n115 plus.n114 0.189894
R183 plus.n114 plus.n113 0.189894
R184 plus.n113 plus.n67 0.189894
R185 plus.n108 plus.n67 0.189894
R186 plus.n108 plus.n107 0.189894
R187 plus.n107 plus.n106 0.189894
R188 plus.n106 plus.n69 0.189894
R189 plus.n101 plus.n69 0.189894
R190 plus.n101 plus.n100 0.189894
R191 plus.n100 plus.n99 0.189894
R192 plus.n99 plus.n72 0.189894
R193 plus.n94 plus.n72 0.189894
R194 plus.n94 plus.n93 0.189894
R195 plus.n93 plus.n74 0.189894
R196 plus.n89 plus.n74 0.189894
R197 plus.n89 plus.n88 0.189894
R198 plus.n88 plus.n76 0.189894
R199 plus.n84 plus.n76 0.189894
R200 plus.n84 plus.n83 0.189894
R201 plus.n83 plus.n78 0.189894
R202 drain_left.n13 drain_left.n11 80.9197
R203 drain_left.n7 drain_left.n5 80.9196
R204 drain_left.n2 drain_left.n0 80.9196
R205 drain_left.n21 drain_left.n20 79.7731
R206 drain_left.n19 drain_left.n18 79.7731
R207 drain_left.n17 drain_left.n16 79.7731
R208 drain_left.n15 drain_left.n14 79.7731
R209 drain_left.n13 drain_left.n12 79.7731
R210 drain_left.n7 drain_left.n6 79.773
R211 drain_left.n9 drain_left.n8 79.773
R212 drain_left.n4 drain_left.n3 79.773
R213 drain_left.n2 drain_left.n1 79.773
R214 drain_left drain_left.n10 31.4411
R215 drain_left drain_left.n21 6.79977
R216 drain_left.n5 drain_left.t0 6.6005
R217 drain_left.n5 drain_left.t2 6.6005
R218 drain_left.n6 drain_left.t9 6.6005
R219 drain_left.n6 drain_left.t18 6.6005
R220 drain_left.n8 drain_left.t13 6.6005
R221 drain_left.n8 drain_left.t19 6.6005
R222 drain_left.n3 drain_left.t22 6.6005
R223 drain_left.n3 drain_left.t14 6.6005
R224 drain_left.n1 drain_left.t5 6.6005
R225 drain_left.n1 drain_left.t6 6.6005
R226 drain_left.n0 drain_left.t4 6.6005
R227 drain_left.n0 drain_left.t15 6.6005
R228 drain_left.n20 drain_left.t8 6.6005
R229 drain_left.n20 drain_left.t17 6.6005
R230 drain_left.n18 drain_left.t12 6.6005
R231 drain_left.n18 drain_left.t7 6.6005
R232 drain_left.n16 drain_left.t21 6.6005
R233 drain_left.n16 drain_left.t1 6.6005
R234 drain_left.n14 drain_left.t11 6.6005
R235 drain_left.n14 drain_left.t20 6.6005
R236 drain_left.n12 drain_left.t10 6.6005
R237 drain_left.n12 drain_left.t23 6.6005
R238 drain_left.n11 drain_left.t3 6.6005
R239 drain_left.n11 drain_left.t16 6.6005
R240 drain_left.n9 drain_left.n7 1.14705
R241 drain_left.n4 drain_left.n2 1.14705
R242 drain_left.n15 drain_left.n13 1.14705
R243 drain_left.n17 drain_left.n15 1.14705
R244 drain_left.n19 drain_left.n17 1.14705
R245 drain_left.n21 drain_left.n19 1.14705
R246 drain_left.n10 drain_left.n9 0.51843
R247 drain_left.n10 drain_left.n4 0.51843
R248 source.n0 source.t39 69.6943
R249 source.n11 source.t23 69.6943
R250 source.n12 source.t9 69.6943
R251 source.n23 source.t7 69.6943
R252 source.n47 source.t12 69.6942
R253 source.n36 source.t0 69.6942
R254 source.n35 source.t31 69.6942
R255 source.n24 source.t25 69.6942
R256 source.n2 source.n1 63.0943
R257 source.n4 source.n3 63.0943
R258 source.n6 source.n5 63.0943
R259 source.n8 source.n7 63.0943
R260 source.n10 source.n9 63.0943
R261 source.n14 source.n13 63.0943
R262 source.n16 source.n15 63.0943
R263 source.n18 source.n17 63.0943
R264 source.n20 source.n19 63.0943
R265 source.n22 source.n21 63.0943
R266 source.n46 source.n45 63.0942
R267 source.n44 source.n43 63.0942
R268 source.n42 source.n41 63.0942
R269 source.n40 source.n39 63.0942
R270 source.n38 source.n37 63.0942
R271 source.n34 source.n33 63.0942
R272 source.n32 source.n31 63.0942
R273 source.n30 source.n29 63.0942
R274 source.n28 source.n27 63.0942
R275 source.n26 source.n25 63.0942
R276 source.n24 source.n23 15.6161
R277 source.n48 source.n0 9.77989
R278 source.n45 source.t17 6.6005
R279 source.n45 source.t4 6.6005
R280 source.n43 source.t2 6.6005
R281 source.n43 source.t14 6.6005
R282 source.n41 source.t3 6.6005
R283 source.n41 source.t47 6.6005
R284 source.n39 source.t5 6.6005
R285 source.n39 source.t16 6.6005
R286 source.n37 source.t8 6.6005
R287 source.n37 source.t13 6.6005
R288 source.n33 source.t28 6.6005
R289 source.n33 source.t37 6.6005
R290 source.n31 source.t26 6.6005
R291 source.n31 source.t24 6.6005
R292 source.n29 source.t42 6.6005
R293 source.n29 source.t36 6.6005
R294 source.n27 source.t41 6.6005
R295 source.n27 source.t27 6.6005
R296 source.n25 source.t35 6.6005
R297 source.n25 source.t45 6.6005
R298 source.n1 source.t30 6.6005
R299 source.n1 source.t34 6.6005
R300 source.n3 source.t33 6.6005
R301 source.n3 source.t38 6.6005
R302 source.n5 source.t40 6.6005
R303 source.n5 source.t29 6.6005
R304 source.n7 source.t43 6.6005
R305 source.n7 source.t32 6.6005
R306 source.n9 source.t44 6.6005
R307 source.n9 source.t46 6.6005
R308 source.n13 source.t18 6.6005
R309 source.n13 source.t11 6.6005
R310 source.n15 source.t21 6.6005
R311 source.n15 source.t15 6.6005
R312 source.n17 source.t1 6.6005
R313 source.n17 source.t22 6.6005
R314 source.n19 source.t20 6.6005
R315 source.n19 source.t19 6.6005
R316 source.n21 source.t10 6.6005
R317 source.n21 source.t6 6.6005
R318 source.n48 source.n47 5.83671
R319 source.n23 source.n22 1.14705
R320 source.n22 source.n20 1.14705
R321 source.n20 source.n18 1.14705
R322 source.n18 source.n16 1.14705
R323 source.n16 source.n14 1.14705
R324 source.n14 source.n12 1.14705
R325 source.n11 source.n10 1.14705
R326 source.n10 source.n8 1.14705
R327 source.n8 source.n6 1.14705
R328 source.n6 source.n4 1.14705
R329 source.n4 source.n2 1.14705
R330 source.n2 source.n0 1.14705
R331 source.n26 source.n24 1.14705
R332 source.n28 source.n26 1.14705
R333 source.n30 source.n28 1.14705
R334 source.n32 source.n30 1.14705
R335 source.n34 source.n32 1.14705
R336 source.n35 source.n34 1.14705
R337 source.n38 source.n36 1.14705
R338 source.n40 source.n38 1.14705
R339 source.n42 source.n40 1.14705
R340 source.n44 source.n42 1.14705
R341 source.n46 source.n44 1.14705
R342 source.n47 source.n46 1.14705
R343 source.n12 source.n11 0.470328
R344 source.n36 source.n35 0.470328
R345 source source.n48 0.188
R346 minus.n60 minus.n0 161.3
R347 minus.n59 minus.n58 161.3
R348 minus.n57 minus.n56 161.3
R349 minus.n55 minus.n2 161.3
R350 minus.n53 minus.n52 161.3
R351 minus.n51 minus.n3 161.3
R352 minus.n50 minus.n49 161.3
R353 minus.n47 minus.n4 161.3
R354 minus.n46 minus.n45 161.3
R355 minus.n44 minus.n5 161.3
R356 minus.n43 minus.n42 161.3
R357 minus.n41 minus.n6 161.3
R358 minus.n39 minus.n38 161.3
R359 minus.n37 minus.n8 161.3
R360 minus.n36 minus.n35 161.3
R361 minus.n33 minus.n9 161.3
R362 minus.n32 minus.n31 161.3
R363 minus.n30 minus.n29 161.3
R364 minus.n28 minus.n11 161.3
R365 minus.n27 minus.n26 161.3
R366 minus.n25 minus.n24 161.3
R367 minus.n23 minus.n13 161.3
R368 minus.n22 minus.n21 161.3
R369 minus.n20 minus.n19 161.3
R370 minus.n18 minus.n15 161.3
R371 minus.n123 minus.n63 161.3
R372 minus.n122 minus.n121 161.3
R373 minus.n120 minus.n119 161.3
R374 minus.n118 minus.n65 161.3
R375 minus.n116 minus.n115 161.3
R376 minus.n114 minus.n66 161.3
R377 minus.n113 minus.n112 161.3
R378 minus.n110 minus.n67 161.3
R379 minus.n109 minus.n108 161.3
R380 minus.n107 minus.n68 161.3
R381 minus.n106 minus.n105 161.3
R382 minus.n103 minus.n69 161.3
R383 minus.n101 minus.n100 161.3
R384 minus.n99 minus.n70 161.3
R385 minus.n98 minus.n97 161.3
R386 minus.n95 minus.n71 161.3
R387 minus.n94 minus.n93 161.3
R388 minus.n92 minus.n91 161.3
R389 minus.n90 minus.n73 161.3
R390 minus.n89 minus.n88 161.3
R391 minus.n87 minus.n86 161.3
R392 minus.n85 minus.n75 161.3
R393 minus.n84 minus.n83 161.3
R394 minus.n82 minus.n81 161.3
R395 minus.n80 minus.n77 161.3
R396 minus.n16 minus.t14 133.606
R397 minus.n78 minus.t23 133.606
R398 minus.n61 minus.t2 111.584
R399 minus.n124 minus.t12 111.584
R400 minus.n62 minus.n61 80.6037
R401 minus.n125 minus.n124 80.6037
R402 minus.n17 minus.t17 72.3005
R403 minus.n14 minus.t16 72.3005
R404 minus.n12 minus.t19 72.3005
R405 minus.n10 minus.t3 72.3005
R406 minus.n34 minus.t0 72.3005
R407 minus.n40 minus.t5 72.3005
R408 minus.n7 minus.t4 72.3005
R409 minus.n48 minus.t1 72.3005
R410 minus.n54 minus.t6 72.3005
R411 minus.n1 minus.t10 72.3005
R412 minus.n79 minus.t21 72.3005
R413 minus.n76 minus.t9 72.3005
R414 minus.n74 minus.t8 72.3005
R415 minus.n72 minus.t13 72.3005
R416 minus.n96 minus.t22 72.3005
R417 minus.n102 minus.t20 72.3005
R418 minus.n104 minus.t11 72.3005
R419 minus.n111 minus.t15 72.3005
R420 minus.n117 minus.t18 72.3005
R421 minus.n64 minus.t7 72.3005
R422 minus.n19 minus.n18 56.5617
R423 minus.n33 minus.n32 56.5617
R424 minus.n42 minus.n41 56.5617
R425 minus.n56 minus.n55 56.5617
R426 minus.n81 minus.n80 56.5617
R427 minus.n95 minus.n94 56.5617
R428 minus.n105 minus.n103 56.5617
R429 minus.n119 minus.n118 56.5617
R430 minus.n28 minus.n27 56.0773
R431 minus.n47 minus.n46 56.0773
R432 minus.n90 minus.n89 56.0773
R433 minus.n110 minus.n109 56.0773
R434 minus.n61 minus.n60 46.0096
R435 minus.n124 minus.n123 46.0096
R436 minus.n24 minus.n23 41.5458
R437 minus.n49 minus.n3 41.5458
R438 minus.n86 minus.n85 41.5458
R439 minus.n112 minus.n66 41.5458
R440 minus.n35 minus.n8 40.577
R441 minus.n39 minus.n8 40.577
R442 minus.n97 minus.n70 40.577
R443 minus.n101 minus.n70 40.577
R444 minus.n23 minus.n22 39.6083
R445 minus.n53 minus.n3 39.6083
R446 minus.n85 minus.n84 39.6083
R447 minus.n116 minus.n66 39.6083
R448 minus.n126 minus.n62 38.4252
R449 minus.n17 minus.n16 33.0515
R450 minus.n79 minus.n78 33.0515
R451 minus.n16 minus.n15 28.5514
R452 minus.n78 minus.n77 28.5514
R453 minus.n60 minus.n59 26.0455
R454 minus.n123 minus.n122 26.0455
R455 minus.n29 minus.n28 25.0767
R456 minus.n46 minus.n5 25.0767
R457 minus.n91 minus.n90 25.0767
R458 minus.n109 minus.n68 25.0767
R459 minus.n32 minus.n10 24.3464
R460 minus.n42 minus.n7 24.3464
R461 minus.n94 minus.n72 24.3464
R462 minus.n105 minus.n104 24.3464
R463 minus.n18 minus.n17 23.8546
R464 minus.n56 minus.n1 23.8546
R465 minus.n80 minus.n79 23.8546
R466 minus.n119 minus.n64 23.8546
R467 minus.n19 minus.n14 16.9689
R468 minus.n55 minus.n54 16.9689
R469 minus.n81 minus.n76 16.9689
R470 minus.n118 minus.n117 16.9689
R471 minus.n34 minus.n33 16.477
R472 minus.n41 minus.n40 16.477
R473 minus.n96 minus.n95 16.477
R474 minus.n103 minus.n102 16.477
R475 minus.n27 minus.n12 15.9852
R476 minus.n48 minus.n47 15.9852
R477 minus.n89 minus.n74 15.9852
R478 minus.n111 minus.n110 15.9852
R479 minus.n24 minus.n12 8.60764
R480 minus.n49 minus.n48 8.60764
R481 minus.n86 minus.n74 8.60764
R482 minus.n112 minus.n111 8.60764
R483 minus.n35 minus.n34 8.11581
R484 minus.n40 minus.n39 8.11581
R485 minus.n97 minus.n96 8.11581
R486 minus.n102 minus.n101 8.11581
R487 minus.n22 minus.n14 7.62397
R488 minus.n54 minus.n53 7.62397
R489 minus.n84 minus.n76 7.62397
R490 minus.n117 minus.n116 7.62397
R491 minus.n126 minus.n125 6.81155
R492 minus.n59 minus.n1 0.738255
R493 minus.n122 minus.n64 0.738255
R494 minus.n62 minus.n0 0.285035
R495 minus.n125 minus.n63 0.285035
R496 minus.n29 minus.n10 0.246418
R497 minus.n7 minus.n5 0.246418
R498 minus.n91 minus.n72 0.246418
R499 minus.n104 minus.n68 0.246418
R500 minus.n58 minus.n0 0.189894
R501 minus.n58 minus.n57 0.189894
R502 minus.n57 minus.n2 0.189894
R503 minus.n52 minus.n2 0.189894
R504 minus.n52 minus.n51 0.189894
R505 minus.n51 minus.n50 0.189894
R506 minus.n50 minus.n4 0.189894
R507 minus.n45 minus.n4 0.189894
R508 minus.n45 minus.n44 0.189894
R509 minus.n44 minus.n43 0.189894
R510 minus.n43 minus.n6 0.189894
R511 minus.n38 minus.n6 0.189894
R512 minus.n38 minus.n37 0.189894
R513 minus.n37 minus.n36 0.189894
R514 minus.n36 minus.n9 0.189894
R515 minus.n31 minus.n9 0.189894
R516 minus.n31 minus.n30 0.189894
R517 minus.n30 minus.n11 0.189894
R518 minus.n26 minus.n11 0.189894
R519 minus.n26 minus.n25 0.189894
R520 minus.n25 minus.n13 0.189894
R521 minus.n21 minus.n13 0.189894
R522 minus.n21 minus.n20 0.189894
R523 minus.n20 minus.n15 0.189894
R524 minus.n82 minus.n77 0.189894
R525 minus.n83 minus.n82 0.189894
R526 minus.n83 minus.n75 0.189894
R527 minus.n87 minus.n75 0.189894
R528 minus.n88 minus.n87 0.189894
R529 minus.n88 minus.n73 0.189894
R530 minus.n92 minus.n73 0.189894
R531 minus.n93 minus.n92 0.189894
R532 minus.n93 minus.n71 0.189894
R533 minus.n98 minus.n71 0.189894
R534 minus.n99 minus.n98 0.189894
R535 minus.n100 minus.n99 0.189894
R536 minus.n100 minus.n69 0.189894
R537 minus.n106 minus.n69 0.189894
R538 minus.n107 minus.n106 0.189894
R539 minus.n108 minus.n107 0.189894
R540 minus.n108 minus.n67 0.189894
R541 minus.n113 minus.n67 0.189894
R542 minus.n114 minus.n113 0.189894
R543 minus.n115 minus.n114 0.189894
R544 minus.n115 minus.n65 0.189894
R545 minus.n120 minus.n65 0.189894
R546 minus.n121 minus.n120 0.189894
R547 minus.n121 minus.n63 0.189894
R548 minus minus.n126 0.188
R549 drain_right.n13 drain_right.n11 80.9197
R550 drain_right.n7 drain_right.n5 80.9196
R551 drain_right.n2 drain_right.n0 80.9196
R552 drain_right.n13 drain_right.n12 79.7731
R553 drain_right.n15 drain_right.n14 79.7731
R554 drain_right.n17 drain_right.n16 79.7731
R555 drain_right.n19 drain_right.n18 79.7731
R556 drain_right.n21 drain_right.n20 79.7731
R557 drain_right.n7 drain_right.n6 79.773
R558 drain_right.n9 drain_right.n8 79.773
R559 drain_right.n4 drain_right.n3 79.773
R560 drain_right.n2 drain_right.n1 79.773
R561 drain_right drain_right.n10 30.8879
R562 drain_right drain_right.n21 6.79977
R563 drain_right.n5 drain_right.t16 6.6005
R564 drain_right.n5 drain_right.t11 6.6005
R565 drain_right.n6 drain_right.t8 6.6005
R566 drain_right.n6 drain_right.t5 6.6005
R567 drain_right.n8 drain_right.t3 6.6005
R568 drain_right.n8 drain_right.t12 6.6005
R569 drain_right.n3 drain_right.t10 6.6005
R570 drain_right.n3 drain_right.t1 6.6005
R571 drain_right.n1 drain_right.t14 6.6005
R572 drain_right.n1 drain_right.t15 6.6005
R573 drain_right.n0 drain_right.t0 6.6005
R574 drain_right.n0 drain_right.t2 6.6005
R575 drain_right.n11 drain_right.t6 6.6005
R576 drain_right.n11 drain_right.t9 6.6005
R577 drain_right.n12 drain_right.t4 6.6005
R578 drain_right.n12 drain_right.t7 6.6005
R579 drain_right.n14 drain_right.t23 6.6005
R580 drain_right.n14 drain_right.t20 6.6005
R581 drain_right.n16 drain_right.t19 6.6005
R582 drain_right.n16 drain_right.t18 6.6005
R583 drain_right.n18 drain_right.t17 6.6005
R584 drain_right.n18 drain_right.t22 6.6005
R585 drain_right.n20 drain_right.t21 6.6005
R586 drain_right.n20 drain_right.t13 6.6005
R587 drain_right.n9 drain_right.n7 1.14705
R588 drain_right.n4 drain_right.n2 1.14705
R589 drain_right.n21 drain_right.n19 1.14705
R590 drain_right.n19 drain_right.n17 1.14705
R591 drain_right.n17 drain_right.n15 1.14705
R592 drain_right.n15 drain_right.n13 1.14705
R593 drain_right.n10 drain_right.n9 0.51843
R594 drain_right.n10 drain_right.n4 0.51843
C0 plus drain_left 5.53495f
C1 drain_right source 10.1116f
C2 drain_right minus 5.11354f
C3 plus drain_right 0.588209f
C4 minus source 6.30846f
C5 plus source 6.32246f
C6 plus minus 6.696569f
C7 drain_right drain_left 2.34071f
C8 drain_left source 10.1074f
C9 drain_left minus 0.181512f
C10 drain_right a_n4174_n1488# 7.30295f
C11 drain_left a_n4174_n1488# 7.89609f
C12 source a_n4174_n1488# 4.50549f
C13 minus a_n4174_n1488# 16.292759f
C14 plus a_n4174_n1488# 17.774471f
C15 drain_right.t0 a_n4174_n1488# 0.07024f
C16 drain_right.t2 a_n4174_n1488# 0.07024f
C17 drain_right.n0 a_n4174_n1488# 0.513195f
C18 drain_right.t14 a_n4174_n1488# 0.07024f
C19 drain_right.t15 a_n4174_n1488# 0.07024f
C20 drain_right.n1 a_n4174_n1488# 0.506563f
C21 drain_right.n2 a_n4174_n1488# 0.917488f
C22 drain_right.t10 a_n4174_n1488# 0.07024f
C23 drain_right.t1 a_n4174_n1488# 0.07024f
C24 drain_right.n3 a_n4174_n1488# 0.506563f
C25 drain_right.n4 a_n4174_n1488# 0.397405f
C26 drain_right.t16 a_n4174_n1488# 0.07024f
C27 drain_right.t11 a_n4174_n1488# 0.07024f
C28 drain_right.n5 a_n4174_n1488# 0.513195f
C29 drain_right.t8 a_n4174_n1488# 0.07024f
C30 drain_right.t5 a_n4174_n1488# 0.07024f
C31 drain_right.n6 a_n4174_n1488# 0.506563f
C32 drain_right.n7 a_n4174_n1488# 0.917489f
C33 drain_right.t3 a_n4174_n1488# 0.07024f
C34 drain_right.t12 a_n4174_n1488# 0.07024f
C35 drain_right.n8 a_n4174_n1488# 0.506563f
C36 drain_right.n9 a_n4174_n1488# 0.397405f
C37 drain_right.n10 a_n4174_n1488# 1.58022f
C38 drain_right.t6 a_n4174_n1488# 0.07024f
C39 drain_right.t9 a_n4174_n1488# 0.07024f
C40 drain_right.n11 a_n4174_n1488# 0.513197f
C41 drain_right.t4 a_n4174_n1488# 0.07024f
C42 drain_right.t7 a_n4174_n1488# 0.07024f
C43 drain_right.n12 a_n4174_n1488# 0.506566f
C44 drain_right.n13 a_n4174_n1488# 0.917484f
C45 drain_right.t23 a_n4174_n1488# 0.07024f
C46 drain_right.t20 a_n4174_n1488# 0.07024f
C47 drain_right.n14 a_n4174_n1488# 0.506566f
C48 drain_right.n15 a_n4174_n1488# 0.456091f
C49 drain_right.t19 a_n4174_n1488# 0.07024f
C50 drain_right.t18 a_n4174_n1488# 0.07024f
C51 drain_right.n16 a_n4174_n1488# 0.506566f
C52 drain_right.n17 a_n4174_n1488# 0.456091f
C53 drain_right.t17 a_n4174_n1488# 0.07024f
C54 drain_right.t22 a_n4174_n1488# 0.07024f
C55 drain_right.n18 a_n4174_n1488# 0.506566f
C56 drain_right.n19 a_n4174_n1488# 0.456091f
C57 drain_right.t21 a_n4174_n1488# 0.07024f
C58 drain_right.t13 a_n4174_n1488# 0.07024f
C59 drain_right.n20 a_n4174_n1488# 0.506566f
C60 drain_right.n21 a_n4174_n1488# 0.728715f
C61 minus.n0 a_n4174_n1488# 0.04848f
C62 minus.t10 a_n4174_n1488# 0.271513f
C63 minus.n1 a_n4174_n1488# 0.135078f
C64 minus.n2 a_n4174_n1488# 0.036331f
C65 minus.t6 a_n4174_n1488# 0.271513f
C66 minus.n3 a_n4174_n1488# 0.02939f
C67 minus.n4 a_n4174_n1488# 0.036331f
C68 minus.t1 a_n4174_n1488# 0.271513f
C69 minus.n5 a_n4174_n1488# 0.035075f
C70 minus.n6 a_n4174_n1488# 0.036331f
C71 minus.t4 a_n4174_n1488# 0.271513f
C72 minus.n7 a_n4174_n1488# 0.135078f
C73 minus.t5 a_n4174_n1488# 0.271513f
C74 minus.n8 a_n4174_n1488# 0.029344f
C75 minus.n9 a_n4174_n1488# 0.036331f
C76 minus.t0 a_n4174_n1488# 0.271513f
C77 minus.t3 a_n4174_n1488# 0.271513f
C78 minus.n10 a_n4174_n1488# 0.135078f
C79 minus.n11 a_n4174_n1488# 0.036331f
C80 minus.t19 a_n4174_n1488# 0.271513f
C81 minus.n12 a_n4174_n1488# 0.135078f
C82 minus.n13 a_n4174_n1488# 0.036331f
C83 minus.t16 a_n4174_n1488# 0.271513f
C84 minus.n14 a_n4174_n1488# 0.135078f
C85 minus.n15 a_n4174_n1488# 0.182901f
C86 minus.t17 a_n4174_n1488# 0.271513f
C87 minus.t14 a_n4174_n1488# 0.359245f
C88 minus.n16 a_n4174_n1488# 0.177959f
C89 minus.n17 a_n4174_n1488# 0.189629f
C90 minus.n18 a_n4174_n1488# 0.044779f
C91 minus.n19 a_n4174_n1488# 0.049539f
C92 minus.n20 a_n4174_n1488# 0.036331f
C93 minus.n21 a_n4174_n1488# 0.036331f
C94 minus.n22 a_n4174_n1488# 0.049215f
C95 minus.n23 a_n4174_n1488# 0.02939f
C96 minus.n24 a_n4174_n1488# 0.049826f
C97 minus.n25 a_n4174_n1488# 0.036331f
C98 minus.n26 a_n4174_n1488# 0.036331f
C99 minus.n27 a_n4174_n1488# 0.05013f
C100 minus.n28 a_n4174_n1488# 0.043226f
C101 minus.n29 a_n4174_n1488# 0.035075f
C102 minus.n30 a_n4174_n1488# 0.036331f
C103 minus.n31 a_n4174_n1488# 0.036331f
C104 minus.n32 a_n4174_n1488# 0.044439f
C105 minus.n33 a_n4174_n1488# 0.049879f
C106 minus.n34 a_n4174_n1488# 0.135078f
C107 minus.n35 a_n4174_n1488# 0.049543f
C108 minus.n36 a_n4174_n1488# 0.036331f
C109 minus.n37 a_n4174_n1488# 0.036331f
C110 minus.n38 a_n4174_n1488# 0.036331f
C111 minus.n39 a_n4174_n1488# 0.049543f
C112 minus.n40 a_n4174_n1488# 0.135078f
C113 minus.n41 a_n4174_n1488# 0.049879f
C114 minus.n42 a_n4174_n1488# 0.044439f
C115 minus.n43 a_n4174_n1488# 0.036331f
C116 minus.n44 a_n4174_n1488# 0.036331f
C117 minus.n45 a_n4174_n1488# 0.036331f
C118 minus.n46 a_n4174_n1488# 0.043226f
C119 minus.n47 a_n4174_n1488# 0.05013f
C120 minus.n48 a_n4174_n1488# 0.135078f
C121 minus.n49 a_n4174_n1488# 0.049826f
C122 minus.n50 a_n4174_n1488# 0.036331f
C123 minus.n51 a_n4174_n1488# 0.036331f
C124 minus.n52 a_n4174_n1488# 0.036331f
C125 minus.n53 a_n4174_n1488# 0.049215f
C126 minus.n54 a_n4174_n1488# 0.135078f
C127 minus.n55 a_n4174_n1488# 0.049539f
C128 minus.n56 a_n4174_n1488# 0.044779f
C129 minus.n57 a_n4174_n1488# 0.036331f
C130 minus.n58 a_n4174_n1488# 0.036331f
C131 minus.n59 a_n4174_n1488# 0.036855f
C132 minus.n60 a_n4174_n1488# 0.038101f
C133 minus.t2 a_n4174_n1488# 0.326833f
C134 minus.n61 a_n4174_n1488# 0.188299f
C135 minus.n62 a_n4174_n1488# 1.42934f
C136 minus.n63 a_n4174_n1488# 0.04848f
C137 minus.t7 a_n4174_n1488# 0.271513f
C138 minus.n64 a_n4174_n1488# 0.135078f
C139 minus.n65 a_n4174_n1488# 0.036331f
C140 minus.t18 a_n4174_n1488# 0.271513f
C141 minus.n66 a_n4174_n1488# 0.02939f
C142 minus.n67 a_n4174_n1488# 0.036331f
C143 minus.t15 a_n4174_n1488# 0.271513f
C144 minus.n68 a_n4174_n1488# 0.035075f
C145 minus.n69 a_n4174_n1488# 0.036331f
C146 minus.t20 a_n4174_n1488# 0.271513f
C147 minus.n70 a_n4174_n1488# 0.029344f
C148 minus.n71 a_n4174_n1488# 0.036331f
C149 minus.t22 a_n4174_n1488# 0.271513f
C150 minus.t13 a_n4174_n1488# 0.271513f
C151 minus.n72 a_n4174_n1488# 0.135078f
C152 minus.n73 a_n4174_n1488# 0.036331f
C153 minus.t8 a_n4174_n1488# 0.271513f
C154 minus.n74 a_n4174_n1488# 0.135078f
C155 minus.n75 a_n4174_n1488# 0.036331f
C156 minus.t9 a_n4174_n1488# 0.271513f
C157 minus.n76 a_n4174_n1488# 0.135078f
C158 minus.n77 a_n4174_n1488# 0.182901f
C159 minus.t21 a_n4174_n1488# 0.271513f
C160 minus.t23 a_n4174_n1488# 0.359245f
C161 minus.n78 a_n4174_n1488# 0.177959f
C162 minus.n79 a_n4174_n1488# 0.189629f
C163 minus.n80 a_n4174_n1488# 0.044779f
C164 minus.n81 a_n4174_n1488# 0.049539f
C165 minus.n82 a_n4174_n1488# 0.036331f
C166 minus.n83 a_n4174_n1488# 0.036331f
C167 minus.n84 a_n4174_n1488# 0.049215f
C168 minus.n85 a_n4174_n1488# 0.02939f
C169 minus.n86 a_n4174_n1488# 0.049826f
C170 minus.n87 a_n4174_n1488# 0.036331f
C171 minus.n88 a_n4174_n1488# 0.036331f
C172 minus.n89 a_n4174_n1488# 0.05013f
C173 minus.n90 a_n4174_n1488# 0.043226f
C174 minus.n91 a_n4174_n1488# 0.035075f
C175 minus.n92 a_n4174_n1488# 0.036331f
C176 minus.n93 a_n4174_n1488# 0.036331f
C177 minus.n94 a_n4174_n1488# 0.044439f
C178 minus.n95 a_n4174_n1488# 0.049879f
C179 minus.n96 a_n4174_n1488# 0.135078f
C180 minus.n97 a_n4174_n1488# 0.049543f
C181 minus.n98 a_n4174_n1488# 0.036331f
C182 minus.n99 a_n4174_n1488# 0.036331f
C183 minus.n100 a_n4174_n1488# 0.036331f
C184 minus.n101 a_n4174_n1488# 0.049543f
C185 minus.n102 a_n4174_n1488# 0.135078f
C186 minus.n103 a_n4174_n1488# 0.049879f
C187 minus.t11 a_n4174_n1488# 0.271513f
C188 minus.n104 a_n4174_n1488# 0.135078f
C189 minus.n105 a_n4174_n1488# 0.044439f
C190 minus.n106 a_n4174_n1488# 0.036331f
C191 minus.n107 a_n4174_n1488# 0.036331f
C192 minus.n108 a_n4174_n1488# 0.036331f
C193 minus.n109 a_n4174_n1488# 0.043226f
C194 minus.n110 a_n4174_n1488# 0.05013f
C195 minus.n111 a_n4174_n1488# 0.135078f
C196 minus.n112 a_n4174_n1488# 0.049826f
C197 minus.n113 a_n4174_n1488# 0.036331f
C198 minus.n114 a_n4174_n1488# 0.036331f
C199 minus.n115 a_n4174_n1488# 0.036331f
C200 minus.n116 a_n4174_n1488# 0.049215f
C201 minus.n117 a_n4174_n1488# 0.135078f
C202 minus.n118 a_n4174_n1488# 0.049539f
C203 minus.n119 a_n4174_n1488# 0.044779f
C204 minus.n120 a_n4174_n1488# 0.036331f
C205 minus.n121 a_n4174_n1488# 0.036331f
C206 minus.n122 a_n4174_n1488# 0.036855f
C207 minus.n123 a_n4174_n1488# 0.038101f
C208 minus.t12 a_n4174_n1488# 0.326833f
C209 minus.n124 a_n4174_n1488# 0.188299f
C210 minus.n125 a_n4174_n1488# 0.276472f
C211 minus.n126 a_n4174_n1488# 1.702f
C212 source.t39 a_n4174_n1488# 0.584366f
C213 source.n0 a_n4174_n1488# 0.898462f
C214 source.t30 a_n4174_n1488# 0.070373f
C215 source.t34 a_n4174_n1488# 0.070373f
C216 source.n1 a_n4174_n1488# 0.446206f
C217 source.n2 a_n4174_n1488# 0.477928f
C218 source.t33 a_n4174_n1488# 0.070373f
C219 source.t38 a_n4174_n1488# 0.070373f
C220 source.n3 a_n4174_n1488# 0.446206f
C221 source.n4 a_n4174_n1488# 0.477928f
C222 source.t40 a_n4174_n1488# 0.070373f
C223 source.t29 a_n4174_n1488# 0.070373f
C224 source.n5 a_n4174_n1488# 0.446206f
C225 source.n6 a_n4174_n1488# 0.477928f
C226 source.t43 a_n4174_n1488# 0.070373f
C227 source.t32 a_n4174_n1488# 0.070373f
C228 source.n7 a_n4174_n1488# 0.446206f
C229 source.n8 a_n4174_n1488# 0.477928f
C230 source.t44 a_n4174_n1488# 0.070373f
C231 source.t46 a_n4174_n1488# 0.070373f
C232 source.n9 a_n4174_n1488# 0.446206f
C233 source.n10 a_n4174_n1488# 0.477928f
C234 source.t23 a_n4174_n1488# 0.584366f
C235 source.n11 a_n4174_n1488# 0.466966f
C236 source.t9 a_n4174_n1488# 0.584366f
C237 source.n12 a_n4174_n1488# 0.466966f
C238 source.t18 a_n4174_n1488# 0.070373f
C239 source.t11 a_n4174_n1488# 0.070373f
C240 source.n13 a_n4174_n1488# 0.446206f
C241 source.n14 a_n4174_n1488# 0.477928f
C242 source.t21 a_n4174_n1488# 0.070373f
C243 source.t15 a_n4174_n1488# 0.070373f
C244 source.n15 a_n4174_n1488# 0.446206f
C245 source.n16 a_n4174_n1488# 0.477928f
C246 source.t1 a_n4174_n1488# 0.070373f
C247 source.t22 a_n4174_n1488# 0.070373f
C248 source.n17 a_n4174_n1488# 0.446206f
C249 source.n18 a_n4174_n1488# 0.477928f
C250 source.t20 a_n4174_n1488# 0.070373f
C251 source.t19 a_n4174_n1488# 0.070373f
C252 source.n19 a_n4174_n1488# 0.446206f
C253 source.n20 a_n4174_n1488# 0.477928f
C254 source.t10 a_n4174_n1488# 0.070373f
C255 source.t6 a_n4174_n1488# 0.070373f
C256 source.n21 a_n4174_n1488# 0.446206f
C257 source.n22 a_n4174_n1488# 0.477928f
C258 source.t7 a_n4174_n1488# 0.584366f
C259 source.n23 a_n4174_n1488# 1.22213f
C260 source.t25 a_n4174_n1488# 0.584363f
C261 source.n24 a_n4174_n1488# 1.22214f
C262 source.t35 a_n4174_n1488# 0.070373f
C263 source.t45 a_n4174_n1488# 0.070373f
C264 source.n25 a_n4174_n1488# 0.446203f
C265 source.n26 a_n4174_n1488# 0.477931f
C266 source.t41 a_n4174_n1488# 0.070373f
C267 source.t27 a_n4174_n1488# 0.070373f
C268 source.n27 a_n4174_n1488# 0.446203f
C269 source.n28 a_n4174_n1488# 0.477931f
C270 source.t42 a_n4174_n1488# 0.070373f
C271 source.t36 a_n4174_n1488# 0.070373f
C272 source.n29 a_n4174_n1488# 0.446203f
C273 source.n30 a_n4174_n1488# 0.477931f
C274 source.t26 a_n4174_n1488# 0.070373f
C275 source.t24 a_n4174_n1488# 0.070373f
C276 source.n31 a_n4174_n1488# 0.446203f
C277 source.n32 a_n4174_n1488# 0.477931f
C278 source.t28 a_n4174_n1488# 0.070373f
C279 source.t37 a_n4174_n1488# 0.070373f
C280 source.n33 a_n4174_n1488# 0.446203f
C281 source.n34 a_n4174_n1488# 0.477931f
C282 source.t31 a_n4174_n1488# 0.584363f
C283 source.n35 a_n4174_n1488# 0.466969f
C284 source.t0 a_n4174_n1488# 0.584363f
C285 source.n36 a_n4174_n1488# 0.466969f
C286 source.t8 a_n4174_n1488# 0.070373f
C287 source.t13 a_n4174_n1488# 0.070373f
C288 source.n37 a_n4174_n1488# 0.446203f
C289 source.n38 a_n4174_n1488# 0.477931f
C290 source.t5 a_n4174_n1488# 0.070373f
C291 source.t16 a_n4174_n1488# 0.070373f
C292 source.n39 a_n4174_n1488# 0.446203f
C293 source.n40 a_n4174_n1488# 0.477931f
C294 source.t3 a_n4174_n1488# 0.070373f
C295 source.t47 a_n4174_n1488# 0.070373f
C296 source.n41 a_n4174_n1488# 0.446203f
C297 source.n42 a_n4174_n1488# 0.477931f
C298 source.t2 a_n4174_n1488# 0.070373f
C299 source.t14 a_n4174_n1488# 0.070373f
C300 source.n43 a_n4174_n1488# 0.446203f
C301 source.n44 a_n4174_n1488# 0.477931f
C302 source.t17 a_n4174_n1488# 0.070373f
C303 source.t4 a_n4174_n1488# 0.070373f
C304 source.n45 a_n4174_n1488# 0.446203f
C305 source.n46 a_n4174_n1488# 0.477931f
C306 source.t12 a_n4174_n1488# 0.584363f
C307 source.n47 a_n4174_n1488# 0.67978f
C308 source.n48 a_n4174_n1488# 0.887141f
C309 drain_left.t4 a_n4174_n1488# 0.071373f
C310 drain_left.t15 a_n4174_n1488# 0.071373f
C311 drain_left.n0 a_n4174_n1488# 0.521471f
C312 drain_left.t5 a_n4174_n1488# 0.071373f
C313 drain_left.t6 a_n4174_n1488# 0.071373f
C314 drain_left.n1 a_n4174_n1488# 0.514733f
C315 drain_left.n2 a_n4174_n1488# 0.932285f
C316 drain_left.t22 a_n4174_n1488# 0.071373f
C317 drain_left.t14 a_n4174_n1488# 0.071373f
C318 drain_left.n3 a_n4174_n1488# 0.514733f
C319 drain_left.n4 a_n4174_n1488# 0.403814f
C320 drain_left.t0 a_n4174_n1488# 0.071373f
C321 drain_left.t2 a_n4174_n1488# 0.071373f
C322 drain_left.n5 a_n4174_n1488# 0.521471f
C323 drain_left.t9 a_n4174_n1488# 0.071373f
C324 drain_left.t18 a_n4174_n1488# 0.071373f
C325 drain_left.n6 a_n4174_n1488# 0.514733f
C326 drain_left.n7 a_n4174_n1488# 0.932285f
C327 drain_left.t13 a_n4174_n1488# 0.071373f
C328 drain_left.t19 a_n4174_n1488# 0.071373f
C329 drain_left.n8 a_n4174_n1488# 0.514733f
C330 drain_left.n9 a_n4174_n1488# 0.403814f
C331 drain_left.n10 a_n4174_n1488# 1.66391f
C332 drain_left.t3 a_n4174_n1488# 0.071373f
C333 drain_left.t16 a_n4174_n1488# 0.071373f
C334 drain_left.n11 a_n4174_n1488# 0.521474f
C335 drain_left.t10 a_n4174_n1488# 0.071373f
C336 drain_left.t23 a_n4174_n1488# 0.071373f
C337 drain_left.n12 a_n4174_n1488# 0.514736f
C338 drain_left.n13 a_n4174_n1488# 0.93228f
C339 drain_left.t11 a_n4174_n1488# 0.071373f
C340 drain_left.t20 a_n4174_n1488# 0.071373f
C341 drain_left.n14 a_n4174_n1488# 0.514736f
C342 drain_left.n15 a_n4174_n1488# 0.463446f
C343 drain_left.t21 a_n4174_n1488# 0.071373f
C344 drain_left.t1 a_n4174_n1488# 0.071373f
C345 drain_left.n16 a_n4174_n1488# 0.514736f
C346 drain_left.n17 a_n4174_n1488# 0.463446f
C347 drain_left.t12 a_n4174_n1488# 0.071373f
C348 drain_left.t7 a_n4174_n1488# 0.071373f
C349 drain_left.n18 a_n4174_n1488# 0.514736f
C350 drain_left.n19 a_n4174_n1488# 0.463446f
C351 drain_left.t8 a_n4174_n1488# 0.071373f
C352 drain_left.t17 a_n4174_n1488# 0.071373f
C353 drain_left.n20 a_n4174_n1488# 0.514736f
C354 drain_left.n21 a_n4174_n1488# 0.740467f
C355 plus.n0 a_n4174_n1488# 0.049753f
C356 plus.t7 a_n4174_n1488# 0.335418f
C357 plus.t12 a_n4174_n1488# 0.278644f
C358 plus.n1 a_n4174_n1488# 0.138625f
C359 plus.n2 a_n4174_n1488# 0.037285f
C360 plus.t16 a_n4174_n1488# 0.278644f
C361 plus.n3 a_n4174_n1488# 0.030162f
C362 plus.n4 a_n4174_n1488# 0.037285f
C363 plus.t8 a_n4174_n1488# 0.278644f
C364 plus.n5 a_n4174_n1488# 0.035996f
C365 plus.n6 a_n4174_n1488# 0.037285f
C366 plus.t17 a_n4174_n1488# 0.278644f
C367 plus.n7 a_n4174_n1488# 0.030114f
C368 plus.n8 a_n4174_n1488# 0.037285f
C369 plus.t6 a_n4174_n1488# 0.278644f
C370 plus.t14 a_n4174_n1488# 0.278644f
C371 plus.n9 a_n4174_n1488# 0.138625f
C372 plus.n10 a_n4174_n1488# 0.037285f
C373 plus.t3 a_n4174_n1488# 0.278644f
C374 plus.n11 a_n4174_n1488# 0.138625f
C375 plus.n12 a_n4174_n1488# 0.037285f
C376 plus.t0 a_n4174_n1488# 0.278644f
C377 plus.n13 a_n4174_n1488# 0.138625f
C378 plus.n14 a_n4174_n1488# 0.187705f
C379 plus.t2 a_n4174_n1488# 0.278644f
C380 plus.t23 a_n4174_n1488# 0.36868f
C381 plus.n15 a_n4174_n1488# 0.182633f
C382 plus.n16 a_n4174_n1488# 0.19461f
C383 plus.n17 a_n4174_n1488# 0.045955f
C384 plus.n18 a_n4174_n1488# 0.05084f
C385 plus.n19 a_n4174_n1488# 0.037285f
C386 plus.n20 a_n4174_n1488# 0.037285f
C387 plus.n21 a_n4174_n1488# 0.050508f
C388 plus.n22 a_n4174_n1488# 0.030162f
C389 plus.n23 a_n4174_n1488# 0.051134f
C390 plus.n24 a_n4174_n1488# 0.037285f
C391 plus.n25 a_n4174_n1488# 0.037285f
C392 plus.n26 a_n4174_n1488# 0.051446f
C393 plus.n27 a_n4174_n1488# 0.044361f
C394 plus.n28 a_n4174_n1488# 0.035996f
C395 plus.n29 a_n4174_n1488# 0.037285f
C396 plus.n30 a_n4174_n1488# 0.037285f
C397 plus.n31 a_n4174_n1488# 0.045606f
C398 plus.n32 a_n4174_n1488# 0.051189f
C399 plus.n33 a_n4174_n1488# 0.138625f
C400 plus.n34 a_n4174_n1488# 0.050845f
C401 plus.n35 a_n4174_n1488# 0.037285f
C402 plus.n36 a_n4174_n1488# 0.037285f
C403 plus.n37 a_n4174_n1488# 0.037285f
C404 plus.n38 a_n4174_n1488# 0.050845f
C405 plus.n39 a_n4174_n1488# 0.138625f
C406 plus.n40 a_n4174_n1488# 0.051189f
C407 plus.t13 a_n4174_n1488# 0.278644f
C408 plus.n41 a_n4174_n1488# 0.138625f
C409 plus.n42 a_n4174_n1488# 0.045606f
C410 plus.n43 a_n4174_n1488# 0.037285f
C411 plus.n44 a_n4174_n1488# 0.037285f
C412 plus.n45 a_n4174_n1488# 0.037285f
C413 plus.n46 a_n4174_n1488# 0.044361f
C414 plus.n47 a_n4174_n1488# 0.051446f
C415 plus.n48 a_n4174_n1488# 0.138625f
C416 plus.n49 a_n4174_n1488# 0.051134f
C417 plus.n50 a_n4174_n1488# 0.037285f
C418 plus.n51 a_n4174_n1488# 0.037285f
C419 plus.n52 a_n4174_n1488# 0.037285f
C420 plus.n53 a_n4174_n1488# 0.050508f
C421 plus.n54 a_n4174_n1488# 0.138625f
C422 plus.n55 a_n4174_n1488# 0.05084f
C423 plus.n56 a_n4174_n1488# 0.045955f
C424 plus.n57 a_n4174_n1488# 0.037285f
C425 plus.n58 a_n4174_n1488# 0.037285f
C426 plus.n59 a_n4174_n1488# 0.037823f
C427 plus.n60 a_n4174_n1488# 0.039101f
C428 plus.n61 a_n4174_n1488# 0.193244f
C429 plus.n62 a_n4174_n1488# 0.320038f
C430 plus.n63 a_n4174_n1488# 0.049753f
C431 plus.t21 a_n4174_n1488# 0.335418f
C432 plus.t11 a_n4174_n1488# 0.278644f
C433 plus.n64 a_n4174_n1488# 0.138625f
C434 plus.n65 a_n4174_n1488# 0.037285f
C435 plus.t1 a_n4174_n1488# 0.278644f
C436 plus.n66 a_n4174_n1488# 0.030162f
C437 plus.n67 a_n4174_n1488# 0.037285f
C438 plus.t5 a_n4174_n1488# 0.278644f
C439 plus.n68 a_n4174_n1488# 0.035996f
C440 plus.n69 a_n4174_n1488# 0.037285f
C441 plus.t19 a_n4174_n1488# 0.278644f
C442 plus.n70 a_n4174_n1488# 0.138625f
C443 plus.t4 a_n4174_n1488# 0.278644f
C444 plus.n71 a_n4174_n1488# 0.030114f
C445 plus.n72 a_n4174_n1488# 0.037285f
C446 plus.t10 a_n4174_n1488# 0.278644f
C447 plus.t20 a_n4174_n1488# 0.278644f
C448 plus.n73 a_n4174_n1488# 0.138625f
C449 plus.n74 a_n4174_n1488# 0.037285f
C450 plus.t22 a_n4174_n1488# 0.278644f
C451 plus.n75 a_n4174_n1488# 0.138625f
C452 plus.n76 a_n4174_n1488# 0.037285f
C453 plus.t18 a_n4174_n1488# 0.278644f
C454 plus.n77 a_n4174_n1488# 0.138625f
C455 plus.n78 a_n4174_n1488# 0.187705f
C456 plus.t9 a_n4174_n1488# 0.278644f
C457 plus.t15 a_n4174_n1488# 0.36868f
C458 plus.n79 a_n4174_n1488# 0.182633f
C459 plus.n80 a_n4174_n1488# 0.19461f
C460 plus.n81 a_n4174_n1488# 0.045955f
C461 plus.n82 a_n4174_n1488# 0.05084f
C462 plus.n83 a_n4174_n1488# 0.037285f
C463 plus.n84 a_n4174_n1488# 0.037285f
C464 plus.n85 a_n4174_n1488# 0.050508f
C465 plus.n86 a_n4174_n1488# 0.030162f
C466 plus.n87 a_n4174_n1488# 0.051134f
C467 plus.n88 a_n4174_n1488# 0.037285f
C468 plus.n89 a_n4174_n1488# 0.037285f
C469 plus.n90 a_n4174_n1488# 0.051446f
C470 plus.n91 a_n4174_n1488# 0.044361f
C471 plus.n92 a_n4174_n1488# 0.035996f
C472 plus.n93 a_n4174_n1488# 0.037285f
C473 plus.n94 a_n4174_n1488# 0.037285f
C474 plus.n95 a_n4174_n1488# 0.045606f
C475 plus.n96 a_n4174_n1488# 0.051189f
C476 plus.n97 a_n4174_n1488# 0.138625f
C477 plus.n98 a_n4174_n1488# 0.050845f
C478 plus.n99 a_n4174_n1488# 0.037285f
C479 plus.n100 a_n4174_n1488# 0.037285f
C480 plus.n101 a_n4174_n1488# 0.037285f
C481 plus.n102 a_n4174_n1488# 0.050845f
C482 plus.n103 a_n4174_n1488# 0.138625f
C483 plus.n104 a_n4174_n1488# 0.051189f
C484 plus.n105 a_n4174_n1488# 0.045606f
C485 plus.n106 a_n4174_n1488# 0.037285f
C486 plus.n107 a_n4174_n1488# 0.037285f
C487 plus.n108 a_n4174_n1488# 0.037285f
C488 plus.n109 a_n4174_n1488# 0.044361f
C489 plus.n110 a_n4174_n1488# 0.051446f
C490 plus.n111 a_n4174_n1488# 0.138625f
C491 plus.n112 a_n4174_n1488# 0.051134f
C492 plus.n113 a_n4174_n1488# 0.037285f
C493 plus.n114 a_n4174_n1488# 0.037285f
C494 plus.n115 a_n4174_n1488# 0.037285f
C495 plus.n116 a_n4174_n1488# 0.050508f
C496 plus.n117 a_n4174_n1488# 0.138625f
C497 plus.n118 a_n4174_n1488# 0.05084f
C498 plus.n119 a_n4174_n1488# 0.045955f
C499 plus.n120 a_n4174_n1488# 0.037285f
C500 plus.n121 a_n4174_n1488# 0.037285f
C501 plus.n122 a_n4174_n1488# 0.037823f
C502 plus.n123 a_n4174_n1488# 0.039101f
C503 plus.n124 a_n4174_n1488# 0.193244f
C504 plus.n125 a_n4174_n1488# 1.38129f
.ends

