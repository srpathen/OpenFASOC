* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t15 plus.t0 drain_left.t3 a_n2046_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X1 drain_left.t6 plus.t1 source.t14 a_n2046_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X2 drain_left.t5 plus.t2 source.t13 a_n2046_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=1
X3 a_n2046_n1488# a_n2046_n1488# a_n2046_n1488# a_n2046_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=9.36 ps=54.24 w=3 l=1
X4 source.t12 plus.t3 drain_left.t0 a_n2046_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X5 drain_left.t7 plus.t4 source.t11 a_n2046_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=1
X6 drain_right.t7 minus.t0 source.t4 a_n2046_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=1
X7 source.t1 minus.t1 drain_right.t6 a_n2046_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X8 drain_right.t5 minus.t2 source.t0 a_n2046_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=1.17 ps=6.78 w=3 l=1
X9 drain_left.t2 plus.t5 source.t10 a_n2046_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X10 a_n2046_n1488# a_n2046_n1488# a_n2046_n1488# a_n2046_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=1
X11 drain_right.t4 minus.t3 source.t3 a_n2046_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X12 a_n2046_n1488# a_n2046_n1488# a_n2046_n1488# a_n2046_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=1
X13 source.t6 minus.t4 drain_right.t3 a_n2046_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X14 source.t9 plus.t6 drain_left.t1 a_n2046_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=1
X15 source.t5 minus.t5 drain_right.t2 a_n2046_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=1
X16 source.t8 plus.t7 drain_left.t4 a_n2046_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=1
X17 drain_right.t1 minus.t6 source.t7 a_n2046_n1488# sky130_fd_pr__nfet_01v8 ad=0.495 pd=3.33 as=0.495 ps=3.33 w=3 l=1
X18 a_n2046_n1488# a_n2046_n1488# a_n2046_n1488# a_n2046_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0 ps=0 w=3 l=1
X19 source.t2 minus.t7 drain_right.t0 a_n2046_n1488# sky130_fd_pr__nfet_01v8 ad=1.17 pd=6.78 as=0.495 ps=3.33 w=3 l=1
R0 plus.n5 plus.n4 161.3
R1 plus.n6 plus.n1 161.3
R2 plus.n8 plus.n7 161.3
R3 plus.n10 plus.n0 161.3
R4 plus.n18 plus.n17 161.3
R5 plus.n19 plus.n14 161.3
R6 plus.n21 plus.n20 161.3
R7 plus.n23 plus.n13 161.3
R8 plus.n2 plus.t7 126.844
R9 plus.n15 plus.t4 126.844
R10 plus.n11 plus.t2 111.584
R11 plus.n24 plus.t6 111.584
R12 plus.n12 plus.n11 80.6037
R13 plus.n25 plus.n24 80.6037
R14 plus.n9 plus.t0 72.3005
R15 plus.n3 plus.t1 72.3005
R16 plus.n22 plus.t5 72.3005
R17 plus.n16 plus.t3 72.3005
R18 plus.n11 plus.n10 56.3158
R19 plus.n24 plus.n23 56.3158
R20 plus.n3 plus.n2 46.9082
R21 plus.n16 plus.n15 46.9082
R22 plus.n5 plus.n2 43.8991
R23 plus.n18 plus.n15 43.8991
R24 plus.n8 plus.n1 40.577
R25 plus.n4 plus.n1 40.577
R26 plus.n21 plus.n14 40.577
R27 plus.n17 plus.n14 40.577
R28 plus plus.n25 27.723
R29 plus.n10 plus.n9 16.477
R30 plus.n23 plus.n22 16.477
R31 plus plus.n12 9.11458
R32 plus.n9 plus.n8 8.11581
R33 plus.n4 plus.n3 8.11581
R34 plus.n22 plus.n21 8.11581
R35 plus.n17 plus.n16 8.11581
R36 plus.n12 plus.n0 0.285035
R37 plus.n25 plus.n13 0.285035
R38 plus.n6 plus.n5 0.189894
R39 plus.n7 plus.n6 0.189894
R40 plus.n7 plus.n0 0.189894
R41 plus.n20 plus.n13 0.189894
R42 plus.n20 plus.n19 0.189894
R43 plus.n19 plus.n18 0.189894
R44 drain_left.n5 drain_left.n3 80.9197
R45 drain_left.n2 drain_left.n1 80.2909
R46 drain_left.n2 drain_left.n0 80.2909
R47 drain_left.n5 drain_left.n4 79.7731
R48 drain_left drain_left.n2 24.5618
R49 drain_left drain_left.n5 6.79977
R50 drain_left.n1 drain_left.t0 6.6005
R51 drain_left.n1 drain_left.t7 6.6005
R52 drain_left.n0 drain_left.t1 6.6005
R53 drain_left.n0 drain_left.t2 6.6005
R54 drain_left.n4 drain_left.t3 6.6005
R55 drain_left.n4 drain_left.t5 6.6005
R56 drain_left.n3 drain_left.t4 6.6005
R57 drain_left.n3 drain_left.t6 6.6005
R58 source.n0 source.t13 69.6943
R59 source.n3 source.t8 69.6943
R60 source.n4 source.t0 69.6943
R61 source.n7 source.t5 69.6943
R62 source.n15 source.t4 69.6942
R63 source.n12 source.t2 69.6942
R64 source.n11 source.t11 69.6942
R65 source.n8 source.t9 69.6942
R66 source.n2 source.n1 63.0943
R67 source.n6 source.n5 63.0943
R68 source.n14 source.n13 63.0942
R69 source.n10 source.n9 63.0942
R70 source.n8 source.n7 15.6161
R71 source.n16 source.n0 9.77989
R72 source.n13 source.t7 6.6005
R73 source.n13 source.t1 6.6005
R74 source.n9 source.t10 6.6005
R75 source.n9 source.t12 6.6005
R76 source.n1 source.t14 6.6005
R77 source.n1 source.t15 6.6005
R78 source.n5 source.t3 6.6005
R79 source.n5 source.t6 6.6005
R80 source.n16 source.n15 5.83671
R81 source.n7 source.n6 1.14705
R82 source.n6 source.n4 1.14705
R83 source.n3 source.n2 1.14705
R84 source.n2 source.n0 1.14705
R85 source.n10 source.n8 1.14705
R86 source.n11 source.n10 1.14705
R87 source.n14 source.n12 1.14705
R88 source.n15 source.n14 1.14705
R89 source.n4 source.n3 0.470328
R90 source.n12 source.n11 0.470328
R91 source source.n16 0.188
R92 minus.n10 minus.n0 161.3
R93 minus.n8 minus.n7 161.3
R94 minus.n6 minus.n1 161.3
R95 minus.n5 minus.n4 161.3
R96 minus.n23 minus.n13 161.3
R97 minus.n21 minus.n20 161.3
R98 minus.n19 minus.n14 161.3
R99 minus.n18 minus.n17 161.3
R100 minus.n2 minus.t2 126.844
R101 minus.n15 minus.t7 126.844
R102 minus.n11 minus.t5 111.584
R103 minus.n24 minus.t0 111.584
R104 minus.n12 minus.n11 80.6037
R105 minus.n25 minus.n24 80.6037
R106 minus.n3 minus.t4 72.3005
R107 minus.n9 minus.t3 72.3005
R108 minus.n16 minus.t6 72.3005
R109 minus.n22 minus.t1 72.3005
R110 minus.n11 minus.n10 56.3158
R111 minus.n24 minus.n23 56.3158
R112 minus.n3 minus.n2 46.9082
R113 minus.n16 minus.n15 46.9082
R114 minus.n5 minus.n2 43.8991
R115 minus.n18 minus.n15 43.8991
R116 minus.n4 minus.n1 40.577
R117 minus.n8 minus.n1 40.577
R118 minus.n17 minus.n14 40.577
R119 minus.n21 minus.n14 40.577
R120 minus.n26 minus.n12 30.4328
R121 minus.n10 minus.n9 16.477
R122 minus.n23 minus.n22 16.477
R123 minus.n4 minus.n3 8.11581
R124 minus.n9 minus.n8 8.11581
R125 minus.n17 minus.n16 8.11581
R126 minus.n22 minus.n21 8.11581
R127 minus.n26 minus.n25 6.87973
R128 minus.n12 minus.n0 0.285035
R129 minus.n25 minus.n13 0.285035
R130 minus.n7 minus.n0 0.189894
R131 minus.n7 minus.n6 0.189894
R132 minus.n6 minus.n5 0.189894
R133 minus.n19 minus.n18 0.189894
R134 minus.n20 minus.n19 0.189894
R135 minus.n20 minus.n13 0.189894
R136 minus minus.n26 0.188
R137 drain_right.n5 drain_right.n3 80.9197
R138 drain_right.n2 drain_right.n1 80.2909
R139 drain_right.n2 drain_right.n0 80.2909
R140 drain_right.n5 drain_right.n4 79.7731
R141 drain_right drain_right.n2 24.0086
R142 drain_right drain_right.n5 6.79977
R143 drain_right.n1 drain_right.t6 6.6005
R144 drain_right.n1 drain_right.t7 6.6005
R145 drain_right.n0 drain_right.t0 6.6005
R146 drain_right.n0 drain_right.t1 6.6005
R147 drain_right.n3 drain_right.t3 6.6005
R148 drain_right.n3 drain_right.t5 6.6005
R149 drain_right.n4 drain_right.t2 6.6005
R150 drain_right.n4 drain_right.t4 6.6005
C0 minus source 2.28559f
C1 minus drain_left 0.177055f
C2 minus drain_right 1.93186f
C3 plus source 2.29958f
C4 plus drain_left 2.13188f
C5 source drain_left 4.27854f
C6 drain_right plus 0.360895f
C7 drain_right source 4.28211f
C8 drain_right drain_left 0.975109f
C9 minus plus 4.02258f
C10 drain_right a_n2046_n1488# 3.67876f
C11 drain_left a_n2046_n1488# 4.4497f
C12 source a_n2046_n1488# 3.814498f
C13 minus a_n2046_n1488# 7.187183f
C14 plus a_n2046_n1488# 8.3693f
C15 drain_right.t0 a_n2046_n1488# 0.041029f
C16 drain_right.t1 a_n2046_n1488# 0.041029f
C17 drain_right.n0 a_n2046_n1488# 0.297441f
C18 drain_right.t6 a_n2046_n1488# 0.041029f
C19 drain_right.t7 a_n2046_n1488# 0.041029f
C20 drain_right.n1 a_n2046_n1488# 0.297441f
C21 drain_right.n2 a_n2046_n1488# 1.02683f
C22 drain_right.t3 a_n2046_n1488# 0.041029f
C23 drain_right.t5 a_n2046_n1488# 0.041029f
C24 drain_right.n3 a_n2046_n1488# 0.299774f
C25 drain_right.t2 a_n2046_n1488# 0.041029f
C26 drain_right.t4 a_n2046_n1488# 0.041029f
C27 drain_right.n4 a_n2046_n1488# 0.2959f
C28 drain_right.n5 a_n2046_n1488# 0.695178f
C29 minus.n0 a_n2046_n1488# 0.042394f
C30 minus.t3 a_n2046_n1488# 0.23743f
C31 minus.n1 a_n2046_n1488# 0.02566f
C32 minus.t2 a_n2046_n1488# 0.305957f
C33 minus.n2 a_n2046_n1488# 0.163098f
C34 minus.t4 a_n2046_n1488# 0.23743f
C35 minus.n3 a_n2046_n1488# 0.146392f
C36 minus.n4 a_n2046_n1488# 0.043324f
C37 minus.n5 a_n2046_n1488# 0.136009f
C38 minus.n6 a_n2046_n1488# 0.031771f
C39 minus.n7 a_n2046_n1488# 0.031771f
C40 minus.n8 a_n2046_n1488# 0.043324f
C41 minus.n9 a_n2046_n1488# 0.118121f
C42 minus.n10 a_n2046_n1488# 0.043578f
C43 minus.t5 a_n2046_n1488# 0.285806f
C44 minus.n11 a_n2046_n1488# 0.16727f
C45 minus.n12 a_n2046_n1488# 0.869196f
C46 minus.n13 a_n2046_n1488# 0.042394f
C47 minus.t1 a_n2046_n1488# 0.23743f
C48 minus.n14 a_n2046_n1488# 0.02566f
C49 minus.t7 a_n2046_n1488# 0.305957f
C50 minus.n15 a_n2046_n1488# 0.163098f
C51 minus.t6 a_n2046_n1488# 0.23743f
C52 minus.n16 a_n2046_n1488# 0.146392f
C53 minus.n17 a_n2046_n1488# 0.043324f
C54 minus.n18 a_n2046_n1488# 0.136009f
C55 minus.n19 a_n2046_n1488# 0.031771f
C56 minus.n20 a_n2046_n1488# 0.031771f
C57 minus.n21 a_n2046_n1488# 0.043324f
C58 minus.n22 a_n2046_n1488# 0.118121f
C59 minus.n23 a_n2046_n1488# 0.043578f
C60 minus.t0 a_n2046_n1488# 0.285806f
C61 minus.n24 a_n2046_n1488# 0.16727f
C62 minus.n25 a_n2046_n1488# 0.246717f
C63 minus.n26 a_n2046_n1488# 1.04455f
C64 source.t13 a_n2046_n1488# 0.489384f
C65 source.n0 a_n2046_n1488# 0.752427f
C66 source.t14 a_n2046_n1488# 0.058935f
C67 source.t15 a_n2046_n1488# 0.058935f
C68 source.n1 a_n2046_n1488# 0.37368f
C69 source.n2 a_n2046_n1488# 0.400246f
C70 source.t8 a_n2046_n1488# 0.489384f
C71 source.n3 a_n2046_n1488# 0.391066f
C72 source.t0 a_n2046_n1488# 0.489384f
C73 source.n4 a_n2046_n1488# 0.391066f
C74 source.t3 a_n2046_n1488# 0.058935f
C75 source.t6 a_n2046_n1488# 0.058935f
C76 source.n5 a_n2046_n1488# 0.37368f
C77 source.n6 a_n2046_n1488# 0.400246f
C78 source.t5 a_n2046_n1488# 0.489384f
C79 source.n7 a_n2046_n1488# 1.02349f
C80 source.t9 a_n2046_n1488# 0.489381f
C81 source.n8 a_n2046_n1488# 1.02349f
C82 source.t10 a_n2046_n1488# 0.058935f
C83 source.t12 a_n2046_n1488# 0.058935f
C84 source.n9 a_n2046_n1488# 0.373677f
C85 source.n10 a_n2046_n1488# 0.400249f
C86 source.t11 a_n2046_n1488# 0.489381f
C87 source.n11 a_n2046_n1488# 0.391068f
C88 source.t2 a_n2046_n1488# 0.489381f
C89 source.n12 a_n2046_n1488# 0.391068f
C90 source.t7 a_n2046_n1488# 0.058935f
C91 source.t1 a_n2046_n1488# 0.058935f
C92 source.n13 a_n2046_n1488# 0.373677f
C93 source.n14 a_n2046_n1488# 0.400249f
C94 source.t4 a_n2046_n1488# 0.489381f
C95 source.n15 a_n2046_n1488# 0.569289f
C96 source.n16 a_n2046_n1488# 0.742946f
C97 drain_left.t1 a_n2046_n1488# 0.06012f
C98 drain_left.t2 a_n2046_n1488# 0.06012f
C99 drain_left.n0 a_n2046_n1488# 0.435841f
C100 drain_left.t0 a_n2046_n1488# 0.06012f
C101 drain_left.t7 a_n2046_n1488# 0.06012f
C102 drain_left.n1 a_n2046_n1488# 0.435841f
C103 drain_left.n2 a_n2046_n1488# 1.55477f
C104 drain_left.t4 a_n2046_n1488# 0.06012f
C105 drain_left.t6 a_n2046_n1488# 0.06012f
C106 drain_left.n3 a_n2046_n1488# 0.439259f
C107 drain_left.t3 a_n2046_n1488# 0.06012f
C108 drain_left.t5 a_n2046_n1488# 0.06012f
C109 drain_left.n4 a_n2046_n1488# 0.433583f
C110 drain_left.n5 a_n2046_n1488# 1.01864f
C111 plus.n0 a_n2046_n1488# 0.057108f
C112 plus.t2 a_n2046_n1488# 0.385001f
C113 plus.t0 a_n2046_n1488# 0.319835f
C114 plus.n1 a_n2046_n1488# 0.034566f
C115 plus.t7 a_n2046_n1488# 0.412146f
C116 plus.n2 a_n2046_n1488# 0.219704f
C117 plus.t1 a_n2046_n1488# 0.319835f
C118 plus.n3 a_n2046_n1488# 0.197201f
C119 plus.n4 a_n2046_n1488# 0.058361f
C120 plus.n5 a_n2046_n1488# 0.183214f
C121 plus.n6 a_n2046_n1488# 0.042797f
C122 plus.n7 a_n2046_n1488# 0.042797f
C123 plus.n8 a_n2046_n1488# 0.058361f
C124 plus.n9 a_n2046_n1488# 0.159118f
C125 plus.n10 a_n2046_n1488# 0.058703f
C126 plus.n11 a_n2046_n1488# 0.225324f
C127 plus.n12 a_n2046_n1488# 0.374399f
C128 plus.n13 a_n2046_n1488# 0.057108f
C129 plus.t6 a_n2046_n1488# 0.385001f
C130 plus.t5 a_n2046_n1488# 0.319835f
C131 plus.n14 a_n2046_n1488# 0.034566f
C132 plus.t4 a_n2046_n1488# 0.412146f
C133 plus.n15 a_n2046_n1488# 0.219704f
C134 plus.t3 a_n2046_n1488# 0.319835f
C135 plus.n16 a_n2046_n1488# 0.197201f
C136 plus.n17 a_n2046_n1488# 0.058361f
C137 plus.n18 a_n2046_n1488# 0.183214f
C138 plus.n19 a_n2046_n1488# 0.042797f
C139 plus.n20 a_n2046_n1488# 0.042797f
C140 plus.n21 a_n2046_n1488# 0.058361f
C141 plus.n22 a_n2046_n1488# 0.159118f
C142 plus.n23 a_n2046_n1488# 0.058703f
C143 plus.n24 a_n2046_n1488# 0.225324f
C144 plus.n25 a_n2046_n1488# 1.10302f
.ends

