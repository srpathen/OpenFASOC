* NGSPICE file created from opamp92.ext - technology: sky130A

.subckt opamp92 gnd CSoutput output vdd plus minus commonsourceibias outputibias diffpairibias
X0 CSoutput.t143 a_n8300_8799.t44 vdd.t257 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X1 a_n2472_13878.t27 a_n2650_13878.t64 vdd.t22 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X2 a_n2472_13878.t19 a_n2650_13878.t10 a_n2650_13878.t11 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 vdd.t256 a_n8300_8799.t45 CSoutput.t142 vdd.t210 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X4 CSoutput.t141 a_n8300_8799.t46 vdd.t255 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X5 gnd.t302 commonsourceibias.t64 CSoutput.t149 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X6 a_n3827_n3924.t20 diffpairibias.t20 gnd.t15 gnd.t14 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X7 CSoutput.t140 a_n8300_8799.t47 vdd.t254 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X8 commonsourceibias.t63 commonsourceibias.t62 gnd.t301 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X9 gnd.t174 gnd.t172 gnd.t173 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X10 vdd.t126 CSoutput.t160 output.t18 gnd.t321 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X11 a_n2650_8322.t27 a_n2650_13878.t65 a_n8300_8799.t13 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X12 gnd.t171 gnd.t169 gnd.t170 gnd.t87 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X13 CSoutput.t4 commonsourceibias.t65 gnd.t300 gnd.t267 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X14 gnd.t168 gnd.t166 gnd.t167 gnd.t120 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X15 CSoutput.t139 a_n8300_8799.t48 vdd.t253 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X16 gnd.t299 commonsourceibias.t60 commonsourceibias.t61 gnd.t249 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X17 gnd.t165 gnd.t163 gnd.t164 gnd.t113 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X18 gnd.t162 gnd.t161 plus.t4 gnd.t120 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X19 CSoutput.t5 commonsourceibias.t66 gnd.t298 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X20 a_n8300_8799.t33 plus.t5 a_n3827_n3924.t38 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X21 vdd.t252 a_n8300_8799.t49 CSoutput.t138 vdd.t203 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X22 gnd.t160 gnd.t158 gnd.t159 gnd.t87 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X23 minus.t4 gnd.t155 gnd.t157 gnd.t156 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X24 commonsourceibias.t33 commonsourceibias.t32 gnd.t295 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X25 a_n8300_8799.t1 a_n2650_13878.t66 a_n2650_8322.t26 vdd.t3 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X26 CSoutput.t18 commonsourceibias.t67 gnd.t297 gnd.t257 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X27 vdd.t251 a_n8300_8799.t50 CSoutput.t137 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X28 vdd.t250 a_n8300_8799.t51 CSoutput.t136 vdd.t223 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X29 a_n8300_8799.t2 a_n2650_13878.t67 a_n2650_8322.t25 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X30 a_n8300_8799.t25 plus.t6 a_n3827_n3924.t35 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X31 commonsourceibias.t35 commonsourceibias.t34 gnd.t296 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 gnd.t154 gnd.t152 gnd.t153 gnd.t73 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X33 CSoutput.t161 a_n2650_8322.t33 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X34 CSoutput.t135 a_n8300_8799.t52 vdd.t249 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X35 CSoutput.t19 commonsourceibias.t68 gnd.t294 gnd.t175 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X36 a_n3827_n3924.t19 diffpairibias.t21 gnd.t53 gnd.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X37 a_n3827_n3924.t42 minus.t5 a_n2650_13878.t55 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X38 CSoutput.t134 a_n8300_8799.t53 vdd.t248 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X39 gnd.t151 gnd.t148 gnd.t150 gnd.t149 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X40 gnd.t293 commonsourceibias.t69 CSoutput.t158 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X41 a_n3827_n3924.t57 plus.t7 a_n8300_8799.t43 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X42 vdd.t247 a_n8300_8799.t54 CSoutput.t133 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X43 gnd.t292 commonsourceibias.t30 commonsourceibias.t31 gnd.t251 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X44 a_n2650_13878.t62 minus.t6 a_n3827_n3924.t50 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X45 a_n3827_n3924.t53 plus.t8 a_n8300_8799.t39 gnd.t324 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X46 output.t17 CSoutput.t162 vdd.t128 gnd.t320 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X47 a_n3827_n3924.t8 minus.t7 a_n2650_13878.t4 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X48 CSoutput.t132 a_n8300_8799.t55 vdd.t246 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X49 commonsourceibias.t47 commonsourceibias.t46 gnd.t290 gnd.t269 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X50 vdd.t110 vdd.t108 vdd.t109 vdd.t44 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X51 gnd.t291 commonsourceibias.t70 CSoutput.t159 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 a_n2472_13878.t18 a_n2650_13878.t24 a_n2650_13878.t25 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X53 a_n2650_13878.t17 a_n2650_13878.t16 a_n2472_13878.t17 vdd.t113 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X54 CSoutput.t163 a_n2650_8322.t32 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X55 gnd.t289 commonsourceibias.t71 CSoutput.t153 gnd.t177 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X56 CSoutput.t131 a_n8300_8799.t56 vdd.t245 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X57 output.t16 CSoutput.t164 vdd.t129 gnd.t319 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X58 a_n3827_n3924.t5 minus.t8 a_n2650_13878.t1 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X59 vdd.t107 vdd.t105 vdd.t106 vdd.t82 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X60 vdd.t234 a_n8300_8799.t57 CSoutput.t130 vdd.t203 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X61 gnd.t288 commonsourceibias.t44 commonsourceibias.t45 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X62 diffpairibias.t19 diffpairibias.t18 gnd.t62 gnd.t61 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X63 commonsourceibias.t43 commonsourceibias.t42 gnd.t287 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X64 a_n2650_13878.t9 a_n2650_13878.t8 a_n2472_13878.t16 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X65 a_n8300_8799.t15 a_n2650_13878.t68 a_n2650_8322.t24 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X66 CSoutput.t129 a_n8300_8799.t58 vdd.t244 vdd.t212 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X67 commonsourceibias.t41 commonsourceibias.t40 gnd.t286 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X68 a_n2650_13878.t48 minus.t9 a_n3827_n3924.t24 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X69 a_n2650_13878.t7 a_n2650_13878.t6 a_n2472_13878.t15 vdd.t20 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X70 gnd.t147 gnd.t145 plus.t3 gnd.t146 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X71 vdd.t243 a_n8300_8799.t59 CSoutput.t128 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X72 vdd.t242 a_n8300_8799.t60 CSoutput.t127 vdd.t223 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X73 a_n8300_8799.t16 a_n2650_13878.t69 a_n2650_8322.t23 vdd.t28 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X74 gnd.t144 gnd.t142 gnd.t143 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X75 diffpairibias.t17 diffpairibias.t16 gnd.t39 gnd.t38 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X76 gnd.t285 commonsourceibias.t38 commonsourceibias.t39 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X77 CSoutput.t126 a_n8300_8799.t61 vdd.t233 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X78 CSoutput.t154 commonsourceibias.t72 gnd.t284 gnd.t267 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X79 output.t2 outputibias.t8 gnd.t58 gnd.t57 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X80 a_n2650_8322.t22 a_n2650_13878.t70 a_n8300_8799.t28 vdd.t20 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X81 vdd.t104 vdd.t102 vdd.t103 vdd.t69 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X82 CSoutput.t125 a_n8300_8799.t62 vdd.t241 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X83 vdd.t121 CSoutput.t165 output.t15 gnd.t318 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X84 plus.t2 gnd.t139 gnd.t141 gnd.t140 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X85 vdd.t122 CSoutput.t166 output.t14 gnd.t317 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X86 gnd.t283 commonsourceibias.t36 commonsourceibias.t37 gnd.t177 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X87 CSoutput.t12 commonsourceibias.t73 gnd.t282 gnd.t269 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 CSoutput.t13 commonsourceibias.t74 gnd.t281 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 a_n8300_8799.t40 plus.t9 a_n3827_n3924.t54 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X90 CSoutput.t42 commonsourceibias.t75 gnd.t280 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X91 outputibias.t7 outputibias.t6 gnd.t42 gnd.t41 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X92 CSoutput.t43 commonsourceibias.t76 gnd.t279 gnd.t257 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X93 a_n3827_n3924.t18 diffpairibias.t22 gnd.t50 gnd.t49 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X94 vdd.t235 a_n8300_8799.t63 CSoutput.t124 vdd.t201 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X95 a_n3827_n3924.t7 minus.t10 a_n2650_13878.t3 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X96 vdd.t240 a_n8300_8799.t64 CSoutput.t123 vdd.t227 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X97 a_n2650_13878.t23 a_n2650_13878.t22 a_n2472_13878.t14 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X98 vdd.t239 a_n8300_8799.t65 CSoutput.t122 vdd.t182 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X99 vdd.t238 a_n8300_8799.t66 CSoutput.t121 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X100 a_n8300_8799.t29 a_n2650_13878.t71 a_n2650_8322.t21 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X101 a_n2650_13878.t21 a_n2650_13878.t20 a_n2472_13878.t13 vdd.t18 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X102 a_n2650_13878.t60 minus.t11 a_n3827_n3924.t48 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X103 gnd.t278 commonsourceibias.t2 commonsourceibias.t3 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X104 a_n3827_n3924.t56 plus.t10 a_n8300_8799.t42 gnd.t305 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X105 gnd.t277 commonsourceibias.t0 commonsourceibias.t1 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X106 vdd.t237 a_n8300_8799.t67 CSoutput.t120 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X107 CSoutput.t119 a_n8300_8799.t68 vdd.t236 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X108 diffpairibias.t15 diffpairibias.t14 gnd.t17 gnd.t16 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X109 a_n3827_n3924.t51 minus.t12 a_n2650_13878.t63 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X110 vdd.t101 vdd.t99 vdd.t100 vdd.t86 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X111 CSoutput.t118 a_n8300_8799.t69 vdd.t232 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X112 gnd.t276 commonsourceibias.t77 CSoutput.t29 gnd.t214 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X113 vdd.t98 vdd.t95 vdd.t97 vdd.t96 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X114 gnd.t275 commonsourceibias.t78 CSoutput.t30 gnd.t251 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X115 gnd.t274 commonsourceibias.t79 CSoutput.t14 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X116 gnd.t273 commonsourceibias.t80 CSoutput.t15 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X117 CSoutput.t117 a_n8300_8799.t70 vdd.t231 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X118 output.t13 CSoutput.t167 vdd.t123 gnd.t316 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X119 vdd.t230 a_n8300_8799.t71 CSoutput.t116 vdd.t227 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X120 vdd.t10 CSoutput.t168 output.t12 gnd.t315 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X121 vdd.t259 a_n2650_13878.t72 a_n2650_8322.t7 vdd.t258 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X122 a_n2650_13878.t39 a_n2650_13878.t38 a_n2472_13878.t12 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X123 gnd.t272 commonsourceibias.t81 CSoutput.t144 gnd.t249 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X124 vdd.t94 vdd.t92 vdd.t93 vdd.t69 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X125 vdd.t91 vdd.t89 vdd.t90 vdd.t62 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X126 gnd.t138 gnd.t136 gnd.t137 gnd.t99 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X127 a_n2650_8322.t6 a_n2650_13878.t73 vdd.t261 vdd.t260 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X128 a_n3827_n3924.t17 diffpairibias.t23 gnd.t29 gnd.t28 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X129 CSoutput.t115 a_n8300_8799.t72 vdd.t229 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X130 a_n2650_13878.t59 minus.t13 a_n3827_n3924.t47 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X131 a_n3827_n3924.t27 plus.t11 a_n8300_8799.t18 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X132 vdd.t265 a_n2650_13878.t74 a_n2472_13878.t26 vdd.t264 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X133 gnd.t135 gnd.t133 minus.t3 gnd.t134 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X134 gnd.t271 commonsourceibias.t82 CSoutput.t145 gnd.t244 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X135 vdd.t88 vdd.t85 vdd.t87 vdd.t86 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X136 vdd.t228 a_n8300_8799.t73 CSoutput.t114 vdd.t227 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X137 vdd.t226 a_n8300_8799.t74 CSoutput.t113 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X138 a_n8300_8799.t19 plus.t12 a_n3827_n3924.t28 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X139 vdd.t84 vdd.t81 vdd.t83 vdd.t82 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X140 a_n2650_8322.t5 a_n2650_13878.t75 vdd.t267 vdd.t266 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X141 a_n2650_13878.t2 minus.t14 a_n3827_n3924.t6 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X142 a_n8300_8799.t5 a_n2650_13878.t76 a_n2650_8322.t20 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X143 CSoutput.t112 a_n8300_8799.t75 vdd.t225 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X144 diffpairibias.t13 diffpairibias.t12 gnd.t304 gnd.t303 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X145 vdd.t224 a_n8300_8799.t76 CSoutput.t111 vdd.t223 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X146 a_n2650_13878.t13 a_n2650_13878.t12 a_n2472_13878.t11 vdd.t26 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X147 vdd.t222 a_n8300_8799.t77 CSoutput.t110 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X148 a_n8300_8799.t6 a_n2650_13878.t77 a_n2650_8322.t19 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X149 CSoutput.t109 a_n8300_8799.t78 vdd.t221 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X150 CSoutput.t146 commonsourceibias.t83 gnd.t270 gnd.t269 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X151 commonsourceibias.t5 commonsourceibias.t4 gnd.t268 gnd.t267 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X152 CSoutput.t147 commonsourceibias.t84 gnd.t266 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X153 a_n2472_13878.t10 a_n2650_13878.t32 a_n2650_13878.t33 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X154 CSoutput.t20 commonsourceibias.t85 gnd.t265 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X155 vdd.t11 CSoutput.t169 output.t11 gnd.t314 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X156 a_n8300_8799.t36 plus.t13 a_n3827_n3924.t44 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X157 a_n3827_n3924.t4 minus.t15 a_n2650_13878.t0 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X158 a_n3827_n3924.t9 minus.t16 a_n2650_13878.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X159 CSoutput.t21 commonsourceibias.t86 gnd.t264 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X160 gnd.t263 commonsourceibias.t87 CSoutput.t33 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X161 CSoutput.t108 a_n8300_8799.t79 vdd.t220 vdd.t212 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X162 gnd.t262 commonsourceibias.t56 commonsourceibias.t57 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X163 a_n2650_13878.t58 minus.t17 a_n3827_n3924.t46 gnd.t55 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X164 vdd.t6 a_n2650_13878.t78 a_n2650_8322.t4 vdd.t5 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X165 a_n2472_13878.t9 a_n2650_13878.t34 a_n2650_13878.t35 vdd.t3 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X166 vdd.t219 a_n8300_8799.t80 CSoutput.t107 vdd.t210 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X167 vdd.t80 vdd.t78 vdd.t79 vdd.t62 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X168 commonsourceibias.t55 commonsourceibias.t54 gnd.t261 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X169 a_n2650_13878.t37 a_n2650_13878.t36 a_n2472_13878.t8 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X170 gnd.t260 commonsourceibias.t52 commonsourceibias.t53 gnd.t244 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X171 vdd.t218 a_n8300_8799.t81 CSoutput.t106 vdd.t165 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X172 gnd.t259 commonsourceibias.t50 commonsourceibias.t51 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X173 a_n3827_n3924.t16 diffpairibias.t24 gnd.t25 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X174 commonsourceibias.t49 commonsourceibias.t48 gnd.t258 gnd.t257 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X175 a_n3827_n3924.t15 diffpairibias.t25 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X176 outputibias.t5 outputibias.t4 gnd.t37 gnd.t36 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X177 gnd.t256 commonsourceibias.t88 CSoutput.t34 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X178 a_n2650_13878.t61 minus.t18 a_n3827_n3924.t49 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X179 vdd.t217 a_n8300_8799.t82 CSoutput.t105 vdd.t201 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X180 gnd.t255 commonsourceibias.t89 CSoutput.t0 gnd.t214 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X181 gnd.t254 commonsourceibias.t90 CSoutput.t1 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X182 gnd.t252 commonsourceibias.t91 CSoutput.t6 gnd.t251 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X183 gnd.t132 gnd.t130 minus.t2 gnd.t131 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X184 gnd.t250 commonsourceibias.t92 CSoutput.t7 gnd.t249 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X185 a_n2472_13878.t7 a_n2650_13878.t40 a_n2650_13878.t41 vdd.t34 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X186 a_n2650_8322.t18 a_n2650_13878.t79 a_n8300_8799.t4 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X187 vdd.t77 vdd.t75 vdd.t76 vdd.t40 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X188 CSoutput.t104 a_n8300_8799.t83 vdd.t216 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X189 commonsourceibias.t7 commonsourceibias.t6 gnd.t248 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X190 CSoutput.t103 a_n8300_8799.t84 vdd.t215 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X191 a_n2650_13878.t56 minus.t19 a_n3827_n3924.t43 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X192 outputibias.t3 outputibias.t2 gnd.t326 gnd.t325 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X193 gnd.t247 commonsourceibias.t93 CSoutput.t35 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X194 CSoutput.t36 commonsourceibias.t94 gnd.t246 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X195 diffpairibias.t11 diffpairibias.t10 gnd.t60 gnd.t59 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X196 a_n2472_13878.t25 a_n2650_13878.t80 vdd.t115 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X197 gnd.t245 commonsourceibias.t95 CSoutput.t44 gnd.t244 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X198 vdd.t117 a_n2650_13878.t81 a_n2472_13878.t24 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X199 gnd.t243 commonsourceibias.t12 commonsourceibias.t13 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X200 CSoutput.t102 a_n8300_8799.t85 vdd.t213 vdd.t212 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X201 a_n3827_n3924.t1 plus.t14 a_n8300_8799.t7 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X202 vdd.t211 a_n8300_8799.t86 CSoutput.t101 vdd.t210 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X203 commonsourceibias.t11 commonsourceibias.t10 gnd.t242 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X204 vdd.t209 a_n8300_8799.t87 CSoutput.t100 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X205 CSoutput.t45 commonsourceibias.t96 gnd.t241 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X206 CSoutput.t99 a_n8300_8799.t88 vdd.t207 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X207 a_n3827_n3924.t45 minus.t20 a_n2650_13878.t57 gnd.t324 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X208 a_n2472_13878.t6 a_n2650_13878.t42 a_n2650_13878.t43 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X209 diffpairibias.t9 diffpairibias.t8 gnd.t323 gnd.t322 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X210 a_n3827_n3924.t3 plus.t15 a_n8300_8799.t9 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X211 a_n3827_n3924.t25 minus.t21 a_n2650_13878.t49 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X212 a_n8300_8799.t14 plus.t16 a_n3827_n3924.t23 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X213 vdd.t206 a_n8300_8799.t89 CSoutput.t98 vdd.t165 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X214 gnd.t240 commonsourceibias.t8 commonsourceibias.t9 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X215 CSoutput.t24 commonsourceibias.t97 gnd.t238 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X216 a_n2650_8322.t17 a_n2650_13878.t82 a_n8300_8799.t20 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X217 CSoutput.t97 a_n8300_8799.t90 vdd.t205 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X218 diffpairibias.t7 diffpairibias.t6 gnd.t31 gnd.t30 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X219 vdd.t204 a_n8300_8799.t91 CSoutput.t96 vdd.t203 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X220 a_n2472_13878.t5 a_n2650_13878.t44 a_n2650_13878.t45 vdd.t28 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X221 vdd.t74 vdd.t72 vdd.t73 vdd.t51 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X222 vdd.t112 a_n2650_13878.t83 a_n2650_8322.t3 vdd.t111 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X223 vdd.t202 a_n8300_8799.t92 CSoutput.t95 vdd.t201 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X224 vdd.t12 CSoutput.t170 output.t10 gnd.t313 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X225 CSoutput.t171 a_n2650_8322.t31 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X226 CSoutput.t31 commonsourceibias.t98 gnd.t237 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X227 CSoutput.t16 commonsourceibias.t99 gnd.t236 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X228 gnd.t234 commonsourceibias.t100 CSoutput.t8 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X229 CSoutput.t94 a_n8300_8799.t93 vdd.t200 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X230 gnd.t129 gnd.t126 gnd.t128 gnd.t127 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X231 a_n2472_13878.t23 a_n2650_13878.t84 vdd.t269 vdd.t268 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X232 outputibias.t1 outputibias.t0 gnd.t64 gnd.t63 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X233 vdd.t71 vdd.t68 vdd.t70 vdd.t69 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X234 CSoutput.t37 commonsourceibias.t101 gnd.t232 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 vdd.t67 vdd.t65 vdd.t66 vdd.t51 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X236 commonsourceibias.t59 commonsourceibias.t58 gnd.t231 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X237 plus.t1 gnd.t123 gnd.t125 gnd.t124 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X238 vdd.t199 a_n8300_8799.t94 CSoutput.t93 vdd.t182 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X239 CSoutput.t172 a_n2650_8322.t30 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X240 CSoutput.t92 a_n8300_8799.t95 vdd.t198 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X241 gnd.t122 gnd.t119 gnd.t121 gnd.t120 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X242 gnd.t118 gnd.t116 minus.t1 gnd.t117 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X243 gnd.t115 gnd.t112 gnd.t114 gnd.t113 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X244 gnd.t111 gnd.t109 gnd.t110 gnd.t99 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X245 gnd.t108 gnd.t105 gnd.t107 gnd.t106 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X246 vdd.t197 a_n8300_8799.t96 CSoutput.t91 vdd.t176 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X247 a_n3827_n3924.t14 diffpairibias.t26 gnd.t13 gnd.t12 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X248 vdd.t271 a_n2650_13878.t85 a_n2650_8322.t2 vdd.t270 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X249 a_n2650_8322.t16 a_n2650_13878.t86 a_n8300_8799.t26 vdd.t26 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X250 gnd.t229 commonsourceibias.t102 CSoutput.t2 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X251 CSoutput.t90 a_n8300_8799.t97 vdd.t196 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X252 vdd.t64 vdd.t61 vdd.t63 vdd.t62 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X253 vdd.t60 vdd.t58 vdd.t59 vdd.t36 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X254 vdd.t195 a_n8300_8799.t98 CSoutput.t89 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X255 vdd.t194 a_n8300_8799.t99 CSoutput.t88 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X256 output.t1 outputibias.t9 gnd.t27 gnd.t26 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X257 gnd.t227 commonsourceibias.t103 CSoutput.t9 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X258 CSoutput.t38 commonsourceibias.t104 gnd.t226 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X259 a_n3827_n3924.t30 plus.t17 a_n8300_8799.t22 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X260 vdd.t57 vdd.t54 vdd.t56 vdd.t55 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X261 vdd.t193 a_n8300_8799.t100 CSoutput.t87 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X262 a_n8300_8799.t21 plus.t18 a_n3827_n3924.t29 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X263 CSoutput.t86 a_n8300_8799.t101 vdd.t192 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X264 a_n3827_n3924.t41 minus.t22 a_n2650_13878.t54 gnd.t305 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X265 gnd.t225 commonsourceibias.t105 CSoutput.t46 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X266 a_n2472_13878.t4 a_n2650_13878.t30 a_n2650_13878.t31 vdd.t30 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X267 CSoutput.t85 a_n8300_8799.t102 vdd.t190 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X268 CSoutput.t25 commonsourceibias.t106 gnd.t224 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X269 a_n2650_8322.t15 a_n2650_13878.t87 a_n8300_8799.t27 vdd.t113 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X270 vdd.t53 vdd.t50 vdd.t52 vdd.t51 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X271 diffpairibias.t5 diffpairibias.t4 gnd.t328 gnd.t327 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X272 vdd.t49 vdd.t47 vdd.t48 vdd.t36 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X273 a_n3827_n3924.t22 minus.t23 a_n2650_13878.t47 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X274 a_n8300_8799.t32 plus.t19 a_n3827_n3924.t37 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X275 commonsourceibias.t29 commonsourceibias.t28 gnd.t223 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X276 gnd.t221 commonsourceibias.t107 CSoutput.t32 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X277 gnd.t104 gnd.t102 gnd.t103 gnd.t73 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X278 CSoutput.t17 commonsourceibias.t108 gnd.t220 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X279 gnd.t215 commonsourceibias.t14 commonsourceibias.t15 gnd.t214 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X280 CSoutput.t84 a_n8300_8799.t103 vdd.t189 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X281 CSoutput.t83 a_n8300_8799.t104 vdd.t187 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X282 CSoutput.t82 a_n8300_8799.t105 vdd.t185 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X283 a_n3827_n3924.t13 diffpairibias.t27 gnd.t34 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X284 vdd.t184 a_n8300_8799.t106 CSoutput.t81 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X285 CSoutput.t10 commonsourceibias.t109 gnd.t219 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X286 vdd.t183 a_n8300_8799.t107 CSoutput.t80 vdd.t182 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X287 a_n2650_8322.t1 a_n2650_13878.t88 vdd.t15 vdd.t14 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X288 CSoutput.t79 a_n8300_8799.t108 vdd.t181 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X289 CSoutput.t148 commonsourceibias.t110 gnd.t217 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X290 a_n3827_n3924.t34 plus.t20 a_n8300_8799.t24 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X291 vdd.t179 a_n8300_8799.t109 CSoutput.t78 vdd.t176 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X292 CSoutput.t77 a_n8300_8799.t110 vdd.t178 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X293 vdd.t17 a_n2650_13878.t89 a_n2472_13878.t22 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X294 gnd.t216 commonsourceibias.t16 commonsourceibias.t17 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X295 vdd.t177 a_n8300_8799.t111 CSoutput.t76 vdd.t176 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X296 CSoutput.t75 a_n8300_8799.t112 vdd.t175 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X297 output.t9 CSoutput.t173 vdd.t127 gnd.t312 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X298 CSoutput.t23 commonsourceibias.t111 gnd.t213 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X299 CSoutput.t74 a_n8300_8799.t113 vdd.t173 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X300 gnd.t212 commonsourceibias.t112 CSoutput.t22 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X301 vdd.t172 a_n8300_8799.t114 CSoutput.t73 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X302 a_n8300_8799.t31 plus.t21 a_n3827_n3924.t36 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X303 vdd.t170 a_n8300_8799.t115 CSoutput.t72 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X304 CSoutput.t155 commonsourceibias.t113 gnd.t211 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X305 a_n3827_n3924.t32 minus.t24 a_n2650_13878.t51 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X306 commonsourceibias.t21 commonsourceibias.t20 gnd.t204 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X307 a_n2650_8322.t14 a_n2650_13878.t90 a_n8300_8799.t34 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X308 CSoutput.t150 commonsourceibias.t114 gnd.t209 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X309 a_n8300_8799.t35 a_n2650_13878.t91 a_n2650_8322.t13 vdd.t30 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X310 output.t8 CSoutput.t174 vdd.t32 gnd.t311 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X311 gnd.t207 commonsourceibias.t22 commonsourceibias.t23 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X312 a_n2472_13878.t21 a_n2650_13878.t92 vdd.t120 vdd.t119 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X313 gnd.t205 commonsourceibias.t115 CSoutput.t26 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X314 vdd.t46 vdd.t43 vdd.t45 vdd.t44 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X315 vdd.t169 a_n8300_8799.t116 CSoutput.t71 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X316 vdd.t42 vdd.t39 vdd.t41 vdd.t40 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X317 CSoutput.t70 a_n8300_8799.t117 vdd.t168 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X318 gnd.t101 gnd.t98 gnd.t100 gnd.t99 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X319 vdd.t38 vdd.t35 vdd.t37 vdd.t36 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X320 a_n8300_8799.t10 plus.t22 a_n3827_n3924.t10 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X321 commonsourceibias.t19 commonsourceibias.t18 gnd.t202 gnd.t201 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X322 a_n8300_8799.t30 a_n2650_13878.t93 a_n2650_8322.t12 vdd.t34 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X323 a_n2650_8322.t11 a_n2650_13878.t94 a_n8300_8799.t11 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X324 CSoutput.t175 a_n2650_8322.t29 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X325 a_n2650_13878.t53 minus.t25 a_n3827_n3924.t40 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X326 vdd.t166 a_n8300_8799.t118 CSoutput.t69 vdd.t165 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X327 CSoutput.t68 a_n8300_8799.t119 vdd.t161 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X328 CSoutput.t67 a_n8300_8799.t120 vdd.t164 vdd.t145 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X329 gnd.t200 commonsourceibias.t24 commonsourceibias.t25 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X330 CSoutput.t66 a_n8300_8799.t121 vdd.t163 vdd.t145 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X331 a_n2472_13878.t3 a_n2650_13878.t28 a_n2650_13878.t29 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X332 vdd.t162 a_n8300_8799.t122 CSoutput.t65 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X333 gnd.t199 commonsourceibias.t116 CSoutput.t156 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X334 CSoutput.t151 commonsourceibias.t117 gnd.t197 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X335 a_n3827_n3924.t2 plus.t23 a_n8300_8799.t8 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X336 output.t7 CSoutput.t176 vdd.t33 gnd.t310 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X337 gnd.t195 commonsourceibias.t118 CSoutput.t39 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X338 a_n8300_8799.t23 plus.t24 a_n3827_n3924.t33 gnd.t55 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X339 a_n3827_n3924.t12 diffpairibias.t28 gnd.t44 gnd.t43 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X340 vdd.t159 a_n8300_8799.t123 CSoutput.t64 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X341 gnd.t97 gnd.t94 gnd.t96 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X342 CSoutput.t63 a_n8300_8799.t124 vdd.t158 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X343 gnd.t93 gnd.t90 gnd.t92 gnd.t91 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X344 a_n2650_13878.t19 a_n2650_13878.t18 a_n2472_13878.t2 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X345 gnd.t89 gnd.t86 gnd.t88 gnd.t87 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X346 a_n8300_8799.t12 a_n2650_13878.t95 a_n2650_8322.t10 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X347 output.t19 outputibias.t10 gnd.t330 gnd.t329 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X348 vdd.t157 a_n8300_8799.t125 CSoutput.t62 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X349 gnd.t193 commonsourceibias.t119 CSoutput.t27 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X350 CSoutput.t61 a_n8300_8799.t126 vdd.t156 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X351 a_n3827_n3924.t0 plus.t25 a_n8300_8799.t3 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X352 vdd.t124 CSoutput.t177 output.t6 gnd.t309 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X353 gnd.t85 gnd.t82 gnd.t84 gnd.t83 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X354 CSoutput.t157 commonsourceibias.t120 gnd.t191 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X355 CSoutput.t152 commonsourceibias.t121 gnd.t189 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X356 diffpairibias.t3 diffpairibias.t2 gnd.t11 gnd.t10 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X357 vdd.t154 a_n8300_8799.t127 CSoutput.t60 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X358 CSoutput.t59 a_n8300_8799.t128 vdd.t144 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X359 output.t0 outputibias.t11 gnd.t22 gnd.t21 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X360 CSoutput.t58 a_n8300_8799.t129 vdd.t152 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X361 a_n2650_8322.t9 a_n2650_13878.t96 a_n8300_8799.t0 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X362 vdd.t150 a_n8300_8799.t130 CSoutput.t57 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X363 CSoutput.t56 a_n8300_8799.t131 vdd.t148 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X364 diffpairibias.t1 diffpairibias.t0 gnd.t46 gnd.t45 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X365 gnd.t81 gnd.t79 plus.t0 gnd.t80 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X366 a_n8300_8799.t17 plus.t26 a_n3827_n3924.t26 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X367 minus.t0 gnd.t76 gnd.t78 gnd.t77 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X368 CSoutput.t40 commonsourceibias.t122 gnd.t187 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X369 CSoutput.t178 a_n2650_8322.t28 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X370 vdd.t2 a_n2650_13878.t97 a_n2472_13878.t20 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X371 gnd.t185 commonsourceibias.t123 CSoutput.t3 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X372 CSoutput.t55 a_n8300_8799.t132 vdd.t146 vdd.t145 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X373 gnd.t75 gnd.t72 gnd.t74 gnd.t73 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X374 gnd.t71 gnd.t68 gnd.t70 gnd.t69 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X375 vdd.t125 CSoutput.t179 output.t5 gnd.t308 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X376 vdd.t143 a_n8300_8799.t133 CSoutput.t54 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X377 vdd.t141 a_n8300_8799.t134 CSoutput.t53 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X378 CSoutput.t11 commonsourceibias.t124 gnd.t183 gnd.t175 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X379 CSoutput.t52 a_n8300_8799.t135 vdd.t139 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X380 output.t4 CSoutput.t180 vdd.t24 gnd.t307 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X381 gnd.t182 commonsourceibias.t125 CSoutput.t41 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X382 a_n2650_13878.t52 minus.t26 a_n3827_n3924.t39 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X383 gnd.t180 commonsourceibias.t126 CSoutput.t47 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X384 a_n2650_8322.t8 a_n2650_13878.t98 a_n8300_8799.t37 vdd.t18 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X385 vdd.t137 a_n8300_8799.t136 CSoutput.t51 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X386 vdd.t135 a_n8300_8799.t137 CSoutput.t50 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X387 CSoutput.t49 a_n8300_8799.t138 vdd.t133 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X388 output.t3 CSoutput.t181 vdd.t25 gnd.t306 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X389 gnd.t178 commonsourceibias.t127 CSoutput.t28 gnd.t177 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X390 a_n3827_n3924.t52 plus.t27 a_n8300_8799.t38 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X391 a_n2650_8322.t0 a_n2650_13878.t99 vdd.t263 vdd.t262 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X392 a_n2650_13878.t46 minus.t27 a_n3827_n3924.t21 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X393 a_n2472_13878.t1 a_n2650_13878.t14 a_n2650_13878.t15 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X394 commonsourceibias.t27 commonsourceibias.t26 gnd.t176 gnd.t175 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X395 a_n3827_n3924.t11 diffpairibias.t29 gnd.t48 gnd.t47 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X396 a_n2650_13878.t50 minus.t28 a_n3827_n3924.t31 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X397 CSoutput.t48 a_n8300_8799.t139 vdd.t131 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X398 a_n3827_n3924.t55 plus.t28 a_n8300_8799.t41 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X399 a_n2650_13878.t27 a_n2650_13878.t26 a_n2472_13878.t0 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 a_n8300_8799.n185 a_n8300_8799.t131 485.149
R1 a_n8300_8799.n201 a_n8300_8799.t46 485.149
R2 a_n8300_8799.n218 a_n8300_8799.t110 485.149
R3 a_n8300_8799.n134 a_n8300_8799.t96 485.149
R4 a_n8300_8799.n150 a_n8300_8799.t109 485.149
R5 a_n8300_8799.n167 a_n8300_8799.t111 485.149
R6 a_n8300_8799.n195 a_n8300_8799.t94 464.166
R7 a_n8300_8799.n194 a_n8300_8799.t47 464.166
R8 a_n8300_8799.n180 a_n8300_8799.t98 464.166
R9 a_n8300_8799.n193 a_n8300_8799.t97 464.166
R10 a_n8300_8799.n192 a_n8300_8799.t49 464.166
R11 a_n8300_8799.n181 a_n8300_8799.t48 464.166
R12 a_n8300_8799.n191 a_n8300_8799.t116 464.166
R13 a_n8300_8799.n190 a_n8300_8799.t61 464.166
R14 a_n8300_8799.n182 a_n8300_8799.t51 464.166
R15 a_n8300_8799.n189 a_n8300_8799.t120 464.166
R16 a_n8300_8799.n188 a_n8300_8799.t82 464.166
R17 a_n8300_8799.n183 a_n8300_8799.t62 464.166
R18 a_n8300_8799.n187 a_n8300_8799.t137 464.166
R19 a_n8300_8799.n186 a_n8300_8799.t95 464.166
R20 a_n8300_8799.n184 a_n8300_8799.t64 464.166
R21 a_n8300_8799.n211 a_n8300_8799.t107 464.166
R22 a_n8300_8799.n210 a_n8300_8799.t55 464.166
R23 a_n8300_8799.n196 a_n8300_8799.t114 464.166
R24 a_n8300_8799.n209 a_n8300_8799.t113 464.166
R25 a_n8300_8799.n208 a_n8300_8799.t57 464.166
R26 a_n8300_8799.n197 a_n8300_8799.t56 464.166
R27 a_n8300_8799.n207 a_n8300_8799.t130 464.166
R28 a_n8300_8799.n206 a_n8300_8799.t69 464.166
R29 a_n8300_8799.n198 a_n8300_8799.t60 464.166
R30 a_n8300_8799.n205 a_n8300_8799.t132 464.166
R31 a_n8300_8799.n204 a_n8300_8799.t92 464.166
R32 a_n8300_8799.n199 a_n8300_8799.t72 464.166
R33 a_n8300_8799.n203 a_n8300_8799.t50 464.166
R34 a_n8300_8799.n202 a_n8300_8799.t108 464.166
R35 a_n8300_8799.n200 a_n8300_8799.t73 464.166
R36 a_n8300_8799.n228 a_n8300_8799.t65 464.166
R37 a_n8300_8799.n227 a_n8300_8799.t135 464.166
R38 a_n8300_8799.n213 a_n8300_8799.t106 464.166
R39 a_n8300_8799.n226 a_n8300_8799.t129 464.166
R40 a_n8300_8799.n225 a_n8300_8799.t91 464.166
R41 a_n8300_8799.n214 a_n8300_8799.t112 464.166
R42 a_n8300_8799.n224 a_n8300_8799.t59 464.166
R43 a_n8300_8799.n223 a_n8300_8799.t126 464.166
R44 a_n8300_8799.n215 a_n8300_8799.t76 464.166
R45 a_n8300_8799.n222 a_n8300_8799.t121 464.166
R46 a_n8300_8799.n221 a_n8300_8799.t63 464.166
R47 a_n8300_8799.n216 a_n8300_8799.t101 464.166
R48 a_n8300_8799.n220 a_n8300_8799.t54 464.166
R49 a_n8300_8799.n219 a_n8300_8799.t88 464.166
R50 a_n8300_8799.n217 a_n8300_8799.t71 464.166
R51 a_n8300_8799.n133 a_n8300_8799.t128 464.166
R52 a_n8300_8799.n136 a_n8300_8799.t66 464.166
R53 a_n8300_8799.n132 a_n8300_8799.t93 464.166
R54 a_n8300_8799.n137 a_n8300_8799.t123 464.166
R55 a_n8300_8799.n138 a_n8300_8799.t124 464.166
R56 a_n8300_8799.n139 a_n8300_8799.t81 464.166
R57 a_n8300_8799.n140 a_n8300_8799.t105 464.166
R58 a_n8300_8799.n131 a_n8300_8799.t122 464.166
R59 a_n8300_8799.n141 a_n8300_8799.t79 464.166
R60 a_n8300_8799.n142 a_n8300_8799.t80 464.166
R61 a_n8300_8799.n143 a_n8300_8799.t102 464.166
R62 a_n8300_8799.n144 a_n8300_8799.t67 464.166
R63 a_n8300_8799.n130 a_n8300_8799.t68 464.166
R64 a_n8300_8799.n145 a_n8300_8799.t99 464.166
R65 a_n8300_8799.n149 a_n8300_8799.t139 464.166
R66 a_n8300_8799.n152 a_n8300_8799.t74 464.166
R67 a_n8300_8799.n148 a_n8300_8799.t103 464.166
R68 a_n8300_8799.n153 a_n8300_8799.t136 464.166
R69 a_n8300_8799.n154 a_n8300_8799.t138 464.166
R70 a_n8300_8799.n155 a_n8300_8799.t89 464.166
R71 a_n8300_8799.n156 a_n8300_8799.t119 464.166
R72 a_n8300_8799.n147 a_n8300_8799.t134 464.166
R73 a_n8300_8799.n157 a_n8300_8799.t85 464.166
R74 a_n8300_8799.n158 a_n8300_8799.t86 464.166
R75 a_n8300_8799.n159 a_n8300_8799.t117 464.166
R76 a_n8300_8799.n160 a_n8300_8799.t77 464.166
R77 a_n8300_8799.n146 a_n8300_8799.t78 464.166
R78 a_n8300_8799.n161 a_n8300_8799.t115 464.166
R79 a_n8300_8799.n166 a_n8300_8799.t70 464.166
R80 a_n8300_8799.n169 a_n8300_8799.t87 464.166
R81 a_n8300_8799.n165 a_n8300_8799.t53 464.166
R82 a_n8300_8799.n170 a_n8300_8799.t100 464.166
R83 a_n8300_8799.n171 a_n8300_8799.t83 464.166
R84 a_n8300_8799.n172 a_n8300_8799.t118 464.166
R85 a_n8300_8799.n173 a_n8300_8799.t75 464.166
R86 a_n8300_8799.n164 a_n8300_8799.t125 464.166
R87 a_n8300_8799.n174 a_n8300_8799.t58 464.166
R88 a_n8300_8799.n175 a_n8300_8799.t45 464.166
R89 a_n8300_8799.n176 a_n8300_8799.t90 464.166
R90 a_n8300_8799.n177 a_n8300_8799.t127 464.166
R91 a_n8300_8799.n163 a_n8300_8799.t104 464.166
R92 a_n8300_8799.n178 a_n8300_8799.t133 464.166
R93 a_n8300_8799.n54 a_n8300_8799.n30 74.4178
R94 a_n8300_8799.n186 a_n8300_8799.n54 12.4674
R95 a_n8300_8799.n53 a_n8300_8799.n30 80.107
R96 a_n8300_8799.n53 a_n8300_8799.n187 1.08907
R97 a_n8300_8799.n31 a_n8300_8799.n52 75.3623
R98 a_n8300_8799.n51 a_n8300_8799.n31 70.3058
R99 a_n8300_8799.n33 a_n8300_8799.n50 70.1674
R100 a_n8300_8799.n50 a_n8300_8799.n182 20.9683
R101 a_n8300_8799.n49 a_n8300_8799.n33 75.0448
R102 a_n8300_8799.n190 a_n8300_8799.n49 11.2134
R103 a_n8300_8799.n48 a_n8300_8799.n32 80.4688
R104 a_n8300_8799.n32 a_n8300_8799.n47 74.73
R105 a_n8300_8799.n46 a_n8300_8799.n34 70.1674
R106 a_n8300_8799.n193 a_n8300_8799.n46 20.9683
R107 a_n8300_8799.n34 a_n8300_8799.n45 70.5844
R108 a_n8300_8799.n45 a_n8300_8799.n180 20.1342
R109 a_n8300_8799.n44 a_n8300_8799.n35 75.6825
R110 a_n8300_8799.n194 a_n8300_8799.n44 9.93802
R111 a_n8300_8799.n35 a_n8300_8799.n195 161.3
R112 a_n8300_8799.n65 a_n8300_8799.n24 74.4178
R113 a_n8300_8799.n202 a_n8300_8799.n65 12.4674
R114 a_n8300_8799.n64 a_n8300_8799.n24 80.107
R115 a_n8300_8799.n64 a_n8300_8799.n203 1.08907
R116 a_n8300_8799.n25 a_n8300_8799.n63 75.3623
R117 a_n8300_8799.n62 a_n8300_8799.n25 70.3058
R118 a_n8300_8799.n27 a_n8300_8799.n61 70.1674
R119 a_n8300_8799.n61 a_n8300_8799.n198 20.9683
R120 a_n8300_8799.n60 a_n8300_8799.n27 75.0448
R121 a_n8300_8799.n206 a_n8300_8799.n60 11.2134
R122 a_n8300_8799.n59 a_n8300_8799.n26 80.4688
R123 a_n8300_8799.n26 a_n8300_8799.n58 74.73
R124 a_n8300_8799.n57 a_n8300_8799.n28 70.1674
R125 a_n8300_8799.n209 a_n8300_8799.n57 20.9683
R126 a_n8300_8799.n28 a_n8300_8799.n56 70.5844
R127 a_n8300_8799.n56 a_n8300_8799.n196 20.1342
R128 a_n8300_8799.n55 a_n8300_8799.n29 75.6825
R129 a_n8300_8799.n210 a_n8300_8799.n55 9.93802
R130 a_n8300_8799.n29 a_n8300_8799.n211 161.3
R131 a_n8300_8799.n76 a_n8300_8799.n18 74.4178
R132 a_n8300_8799.n219 a_n8300_8799.n76 12.4674
R133 a_n8300_8799.n75 a_n8300_8799.n18 80.107
R134 a_n8300_8799.n75 a_n8300_8799.n220 1.08907
R135 a_n8300_8799.n19 a_n8300_8799.n74 75.3623
R136 a_n8300_8799.n73 a_n8300_8799.n19 70.3058
R137 a_n8300_8799.n21 a_n8300_8799.n72 70.1674
R138 a_n8300_8799.n72 a_n8300_8799.n215 20.9683
R139 a_n8300_8799.n71 a_n8300_8799.n21 75.0448
R140 a_n8300_8799.n223 a_n8300_8799.n71 11.2134
R141 a_n8300_8799.n70 a_n8300_8799.n20 80.4688
R142 a_n8300_8799.n20 a_n8300_8799.n69 74.73
R143 a_n8300_8799.n68 a_n8300_8799.n22 70.1674
R144 a_n8300_8799.n226 a_n8300_8799.n68 20.9683
R145 a_n8300_8799.n22 a_n8300_8799.n67 70.5844
R146 a_n8300_8799.n67 a_n8300_8799.n213 20.1342
R147 a_n8300_8799.n66 a_n8300_8799.n23 75.6825
R148 a_n8300_8799.n227 a_n8300_8799.n66 9.93802
R149 a_n8300_8799.n23 a_n8300_8799.n228 161.3
R150 a_n8300_8799.n13 a_n8300_8799.n87 70.1674
R151 a_n8300_8799.n145 a_n8300_8799.n87 20.9683
R152 a_n8300_8799.n86 a_n8300_8799.n13 74.4178
R153 a_n8300_8799.n86 a_n8300_8799.n130 12.4674
R154 a_n8300_8799.n12 a_n8300_8799.n85 80.107
R155 a_n8300_8799.n144 a_n8300_8799.n85 1.08907
R156 a_n8300_8799.n84 a_n8300_8799.n12 75.3623
R157 a_n8300_8799.n14 a_n8300_8799.n83 70.3058
R158 a_n8300_8799.n82 a_n8300_8799.n14 70.1674
R159 a_n8300_8799.n82 a_n8300_8799.n131 20.9683
R160 a_n8300_8799.n15 a_n8300_8799.n81 75.0448
R161 a_n8300_8799.n140 a_n8300_8799.n81 11.2134
R162 a_n8300_8799.n80 a_n8300_8799.n15 80.4688
R163 a_n8300_8799.n16 a_n8300_8799.n79 74.73
R164 a_n8300_8799.n78 a_n8300_8799.n16 70.1674
R165 a_n8300_8799.n78 a_n8300_8799.n132 20.9683
R166 a_n8300_8799.n17 a_n8300_8799.n77 70.5844
R167 a_n8300_8799.n136 a_n8300_8799.n77 20.1342
R168 a_n8300_8799.n135 a_n8300_8799.n17 161.3
R169 a_n8300_8799.n7 a_n8300_8799.n98 70.1674
R170 a_n8300_8799.n161 a_n8300_8799.n98 20.9683
R171 a_n8300_8799.n97 a_n8300_8799.n7 74.4178
R172 a_n8300_8799.n97 a_n8300_8799.n146 12.4674
R173 a_n8300_8799.n6 a_n8300_8799.n96 80.107
R174 a_n8300_8799.n160 a_n8300_8799.n96 1.08907
R175 a_n8300_8799.n95 a_n8300_8799.n6 75.3623
R176 a_n8300_8799.n8 a_n8300_8799.n94 70.3058
R177 a_n8300_8799.n93 a_n8300_8799.n8 70.1674
R178 a_n8300_8799.n93 a_n8300_8799.n147 20.9683
R179 a_n8300_8799.n9 a_n8300_8799.n92 75.0448
R180 a_n8300_8799.n156 a_n8300_8799.n92 11.2134
R181 a_n8300_8799.n91 a_n8300_8799.n9 80.4688
R182 a_n8300_8799.n10 a_n8300_8799.n90 74.73
R183 a_n8300_8799.n89 a_n8300_8799.n10 70.1674
R184 a_n8300_8799.n89 a_n8300_8799.n148 20.9683
R185 a_n8300_8799.n11 a_n8300_8799.n88 70.5844
R186 a_n8300_8799.n152 a_n8300_8799.n88 20.1342
R187 a_n8300_8799.n151 a_n8300_8799.n11 161.3
R188 a_n8300_8799.n1 a_n8300_8799.n109 70.1674
R189 a_n8300_8799.n178 a_n8300_8799.n109 20.9683
R190 a_n8300_8799.n108 a_n8300_8799.n1 74.4178
R191 a_n8300_8799.n108 a_n8300_8799.n163 12.4674
R192 a_n8300_8799.n0 a_n8300_8799.n107 80.107
R193 a_n8300_8799.n177 a_n8300_8799.n107 1.08907
R194 a_n8300_8799.n106 a_n8300_8799.n0 75.3623
R195 a_n8300_8799.n2 a_n8300_8799.n105 70.3058
R196 a_n8300_8799.n104 a_n8300_8799.n2 70.1674
R197 a_n8300_8799.n104 a_n8300_8799.n164 20.9683
R198 a_n8300_8799.n3 a_n8300_8799.n103 75.0448
R199 a_n8300_8799.n173 a_n8300_8799.n103 11.2134
R200 a_n8300_8799.n102 a_n8300_8799.n3 80.4688
R201 a_n8300_8799.n4 a_n8300_8799.n101 74.73
R202 a_n8300_8799.n100 a_n8300_8799.n4 70.1674
R203 a_n8300_8799.n100 a_n8300_8799.n165 20.9683
R204 a_n8300_8799.n5 a_n8300_8799.n99 70.5844
R205 a_n8300_8799.n169 a_n8300_8799.n99 20.1342
R206 a_n8300_8799.n168 a_n8300_8799.n5 161.3
R207 a_n8300_8799.n41 a_n8300_8799.n110 98.9633
R208 a_n8300_8799.n39 a_n8300_8799.n113 98.9631
R209 a_n8300_8799.n42 a_n8300_8799.n233 98.6055
R210 a_n8300_8799.n41 a_n8300_8799.n112 98.6055
R211 a_n8300_8799.n41 a_n8300_8799.n111 98.6055
R212 a_n8300_8799.n39 a_n8300_8799.n114 98.6055
R213 a_n8300_8799.n39 a_n8300_8799.n115 98.6055
R214 a_n8300_8799.n40 a_n8300_8799.n116 98.6055
R215 a_n8300_8799.n40 a_n8300_8799.n117 98.6055
R216 a_n8300_8799.n234 a_n8300_8799.n42 98.6054
R217 a_n8300_8799.n37 a_n8300_8799.n118 81.2902
R218 a_n8300_8799.n43 a_n8300_8799.n124 81.2902
R219 a_n8300_8799.n36 a_n8300_8799.n121 81.2902
R220 a_n8300_8799.n38 a_n8300_8799.n127 80.9324
R221 a_n8300_8799.n38 a_n8300_8799.n128 80.9324
R222 a_n8300_8799.n37 a_n8300_8799.n129 80.9324
R223 a_n8300_8799.n37 a_n8300_8799.n120 80.9324
R224 a_n8300_8799.n37 a_n8300_8799.n119 80.9324
R225 a_n8300_8799.n43 a_n8300_8799.n125 80.9324
R226 a_n8300_8799.n36 a_n8300_8799.n126 80.9324
R227 a_n8300_8799.n36 a_n8300_8799.n123 80.9324
R228 a_n8300_8799.n36 a_n8300_8799.n122 80.9324
R229 a_n8300_8799.n30 a_n8300_8799.n185 70.4033
R230 a_n8300_8799.n24 a_n8300_8799.n201 70.4033
R231 a_n8300_8799.n18 a_n8300_8799.n218 70.4033
R232 a_n8300_8799.n17 a_n8300_8799.n134 70.4033
R233 a_n8300_8799.n11 a_n8300_8799.n150 70.4033
R234 a_n8300_8799.n5 a_n8300_8799.n167 70.4033
R235 a_n8300_8799.n195 a_n8300_8799.n194 48.2005
R236 a_n8300_8799.n46 a_n8300_8799.n192 20.9683
R237 a_n8300_8799.n191 a_n8300_8799.n190 48.2005
R238 a_n8300_8799.n189 a_n8300_8799.n50 20.9683
R239 a_n8300_8799.n187 a_n8300_8799.n183 48.2005
R240 a_n8300_8799.n211 a_n8300_8799.n210 48.2005
R241 a_n8300_8799.n57 a_n8300_8799.n208 20.9683
R242 a_n8300_8799.n207 a_n8300_8799.n206 48.2005
R243 a_n8300_8799.n205 a_n8300_8799.n61 20.9683
R244 a_n8300_8799.n203 a_n8300_8799.n199 48.2005
R245 a_n8300_8799.n228 a_n8300_8799.n227 48.2005
R246 a_n8300_8799.n68 a_n8300_8799.n225 20.9683
R247 a_n8300_8799.n224 a_n8300_8799.n223 48.2005
R248 a_n8300_8799.n222 a_n8300_8799.n72 20.9683
R249 a_n8300_8799.n220 a_n8300_8799.n216 48.2005
R250 a_n8300_8799.n137 a_n8300_8799.n78 20.9683
R251 a_n8300_8799.n140 a_n8300_8799.n139 48.2005
R252 a_n8300_8799.n141 a_n8300_8799.n82 20.9683
R253 a_n8300_8799.n144 a_n8300_8799.n143 48.2005
R254 a_n8300_8799.t44 a_n8300_8799.n87 485.135
R255 a_n8300_8799.n153 a_n8300_8799.n89 20.9683
R256 a_n8300_8799.n156 a_n8300_8799.n155 48.2005
R257 a_n8300_8799.n157 a_n8300_8799.n93 20.9683
R258 a_n8300_8799.n160 a_n8300_8799.n159 48.2005
R259 a_n8300_8799.t52 a_n8300_8799.n98 485.135
R260 a_n8300_8799.n170 a_n8300_8799.n100 20.9683
R261 a_n8300_8799.n173 a_n8300_8799.n172 48.2005
R262 a_n8300_8799.n174 a_n8300_8799.n104 20.9683
R263 a_n8300_8799.n177 a_n8300_8799.n176 48.2005
R264 a_n8300_8799.t84 a_n8300_8799.n109 485.135
R265 a_n8300_8799.n48 a_n8300_8799.n181 47.835
R266 a_n8300_8799.n51 a_n8300_8799.n188 20.6913
R267 a_n8300_8799.n59 a_n8300_8799.n197 47.835
R268 a_n8300_8799.n62 a_n8300_8799.n204 20.6913
R269 a_n8300_8799.n70 a_n8300_8799.n214 47.835
R270 a_n8300_8799.n73 a_n8300_8799.n221 20.6913
R271 a_n8300_8799.n138 a_n8300_8799.n80 47.835
R272 a_n8300_8799.n142 a_n8300_8799.n83 20.6913
R273 a_n8300_8799.n154 a_n8300_8799.n91 47.835
R274 a_n8300_8799.n158 a_n8300_8799.n94 20.6913
R275 a_n8300_8799.n171 a_n8300_8799.n102 47.835
R276 a_n8300_8799.n175 a_n8300_8799.n105 20.6913
R277 a_n8300_8799.n193 a_n8300_8799.n45 22.3251
R278 a_n8300_8799.n209 a_n8300_8799.n56 22.3251
R279 a_n8300_8799.n226 a_n8300_8799.n67 22.3251
R280 a_n8300_8799.n132 a_n8300_8799.n77 22.3251
R281 a_n8300_8799.n148 a_n8300_8799.n88 22.3251
R282 a_n8300_8799.n165 a_n8300_8799.n99 22.3251
R283 a_n8300_8799.n232 a_n8300_8799.n40 32.8234
R284 a_n8300_8799.n38 a_n8300_8799.n36 32.5134
R285 a_n8300_8799.n54 a_n8300_8799.n184 33.6462
R286 a_n8300_8799.n65 a_n8300_8799.n200 33.6462
R287 a_n8300_8799.n76 a_n8300_8799.n217 33.6462
R288 a_n8300_8799.n136 a_n8300_8799.n135 27.0217
R289 a_n8300_8799.n145 a_n8300_8799.n86 33.6462
R290 a_n8300_8799.n152 a_n8300_8799.n151 27.0217
R291 a_n8300_8799.n161 a_n8300_8799.n97 33.6462
R292 a_n8300_8799.n169 a_n8300_8799.n168 27.0217
R293 a_n8300_8799.n178 a_n8300_8799.n108 33.6462
R294 a_n8300_8799.n47 a_n8300_8799.n181 11.843
R295 a_n8300_8799.n188 a_n8300_8799.n52 36.139
R296 a_n8300_8799.n58 a_n8300_8799.n197 11.843
R297 a_n8300_8799.n204 a_n8300_8799.n63 36.139
R298 a_n8300_8799.n69 a_n8300_8799.n214 11.843
R299 a_n8300_8799.n221 a_n8300_8799.n74 36.139
R300 a_n8300_8799.n138 a_n8300_8799.n79 11.843
R301 a_n8300_8799.n142 a_n8300_8799.n84 36.139
R302 a_n8300_8799.n154 a_n8300_8799.n90 11.843
R303 a_n8300_8799.n158 a_n8300_8799.n95 36.139
R304 a_n8300_8799.n171 a_n8300_8799.n101 11.843
R305 a_n8300_8799.n175 a_n8300_8799.n106 36.139
R306 a_n8300_8799.n49 a_n8300_8799.n182 35.3134
R307 a_n8300_8799.n60 a_n8300_8799.n198 35.3134
R308 a_n8300_8799.n71 a_n8300_8799.n215 35.3134
R309 a_n8300_8799.n131 a_n8300_8799.n81 35.3134
R310 a_n8300_8799.n147 a_n8300_8799.n92 35.3134
R311 a_n8300_8799.n164 a_n8300_8799.n103 35.3134
R312 a_n8300_8799.n192 a_n8300_8799.n47 34.4824
R313 a_n8300_8799.n52 a_n8300_8799.n183 10.5784
R314 a_n8300_8799.n208 a_n8300_8799.n58 34.4824
R315 a_n8300_8799.n63 a_n8300_8799.n199 10.5784
R316 a_n8300_8799.n225 a_n8300_8799.n69 34.4824
R317 a_n8300_8799.n74 a_n8300_8799.n216 10.5784
R318 a_n8300_8799.n79 a_n8300_8799.n137 34.4824
R319 a_n8300_8799.n143 a_n8300_8799.n84 10.5784
R320 a_n8300_8799.n90 a_n8300_8799.n153 34.4824
R321 a_n8300_8799.n159 a_n8300_8799.n95 10.5784
R322 a_n8300_8799.n101 a_n8300_8799.n170 34.4824
R323 a_n8300_8799.n176 a_n8300_8799.n106 10.5784
R324 a_n8300_8799.n44 a_n8300_8799.n180 36.9592
R325 a_n8300_8799.n55 a_n8300_8799.n196 36.9592
R326 a_n8300_8799.n66 a_n8300_8799.n213 36.9592
R327 a_n8300_8799.n135 a_n8300_8799.n133 21.1793
R328 a_n8300_8799.n151 a_n8300_8799.n149 21.1793
R329 a_n8300_8799.n168 a_n8300_8799.n166 21.1793
R330 a_n8300_8799.n185 a_n8300_8799.n184 20.9576
R331 a_n8300_8799.n201 a_n8300_8799.n200 20.9576
R332 a_n8300_8799.n218 a_n8300_8799.n217 20.9576
R333 a_n8300_8799.n134 a_n8300_8799.n133 20.9576
R334 a_n8300_8799.n150 a_n8300_8799.n149 20.9576
R335 a_n8300_8799.n167 a_n8300_8799.n166 20.9576
R336 a_n8300_8799.n42 a_n8300_8799.n232 19.9193
R337 a_n8300_8799.n231 a_n8300_8799.n37 12.3339
R338 a_n8300_8799.n232 a_n8300_8799.n231 11.4887
R339 a_n8300_8799.n212 a_n8300_8799.n35 9.07815
R340 a_n8300_8799.n162 a_n8300_8799.n13 9.07815
R341 a_n8300_8799.n230 a_n8300_8799.n179 7.07257
R342 a_n8300_8799.n230 a_n8300_8799.n229 6.72634
R343 a_n8300_8799.n212 a_n8300_8799.n29 4.9702
R344 a_n8300_8799.n229 a_n8300_8799.n23 4.9702
R345 a_n8300_8799.n162 a_n8300_8799.n7 4.9702
R346 a_n8300_8799.n179 a_n8300_8799.n1 4.9702
R347 a_n8300_8799.n229 a_n8300_8799.n212 4.10845
R348 a_n8300_8799.n179 a_n8300_8799.n162 4.10845
R349 a_n8300_8799.n233 a_n8300_8799.t4 3.61217
R350 a_n8300_8799.n233 a_n8300_8799.t16 3.61217
R351 a_n8300_8799.n112 a_n8300_8799.t27 3.61217
R352 a_n8300_8799.n112 a_n8300_8799.t12 3.61217
R353 a_n8300_8799.n111 a_n8300_8799.t20 3.61217
R354 a_n8300_8799.n111 a_n8300_8799.t29 3.61217
R355 a_n8300_8799.n110 a_n8300_8799.t37 3.61217
R356 a_n8300_8799.n110 a_n8300_8799.t6 3.61217
R357 a_n8300_8799.n113 a_n8300_8799.t26 3.61217
R358 a_n8300_8799.n113 a_n8300_8799.t2 3.61217
R359 a_n8300_8799.n114 a_n8300_8799.t13 3.61217
R360 a_n8300_8799.n114 a_n8300_8799.t5 3.61217
R361 a_n8300_8799.n115 a_n8300_8799.t34 3.61217
R362 a_n8300_8799.n115 a_n8300_8799.t35 3.61217
R363 a_n8300_8799.n116 a_n8300_8799.t11 3.61217
R364 a_n8300_8799.n116 a_n8300_8799.t15 3.61217
R365 a_n8300_8799.n117 a_n8300_8799.t28 3.61217
R366 a_n8300_8799.n117 a_n8300_8799.t30 3.61217
R367 a_n8300_8799.t0 a_n8300_8799.n234 3.61217
R368 a_n8300_8799.n234 a_n8300_8799.t1 3.61217
R369 a_n8300_8799.n231 a_n8300_8799.n230 3.4105
R370 a_n8300_8799.n127 a_n8300_8799.t41 2.82907
R371 a_n8300_8799.n127 a_n8300_8799.t31 2.82907
R372 a_n8300_8799.n128 a_n8300_8799.t39 2.82907
R373 a_n8300_8799.n128 a_n8300_8799.t14 2.82907
R374 a_n8300_8799.n129 a_n8300_8799.t42 2.82907
R375 a_n8300_8799.n129 a_n8300_8799.t32 2.82907
R376 a_n8300_8799.n120 a_n8300_8799.t18 2.82907
R377 a_n8300_8799.n120 a_n8300_8799.t25 2.82907
R378 a_n8300_8799.n119 a_n8300_8799.t24 2.82907
R379 a_n8300_8799.n119 a_n8300_8799.t17 2.82907
R380 a_n8300_8799.n118 a_n8300_8799.t3 2.82907
R381 a_n8300_8799.n118 a_n8300_8799.t33 2.82907
R382 a_n8300_8799.n124 a_n8300_8799.t9 2.82907
R383 a_n8300_8799.n124 a_n8300_8799.t19 2.82907
R384 a_n8300_8799.n125 a_n8300_8799.t22 2.82907
R385 a_n8300_8799.n125 a_n8300_8799.t40 2.82907
R386 a_n8300_8799.n126 a_n8300_8799.t7 2.82907
R387 a_n8300_8799.n126 a_n8300_8799.t23 2.82907
R388 a_n8300_8799.n123 a_n8300_8799.t43 2.82907
R389 a_n8300_8799.n123 a_n8300_8799.t21 2.82907
R390 a_n8300_8799.n122 a_n8300_8799.t38 2.82907
R391 a_n8300_8799.n122 a_n8300_8799.t10 2.82907
R392 a_n8300_8799.n121 a_n8300_8799.t8 2.82907
R393 a_n8300_8799.n121 a_n8300_8799.t36 2.82907
R394 a_n8300_8799.n53 a_n8300_8799.n186 47.0982
R395 a_n8300_8799.n64 a_n8300_8799.n202 47.0982
R396 a_n8300_8799.n75 a_n8300_8799.n219 47.0982
R397 a_n8300_8799.n130 a_n8300_8799.n85 47.0982
R398 a_n8300_8799.n146 a_n8300_8799.n96 47.0982
R399 a_n8300_8799.n163 a_n8300_8799.n107 47.0982
R400 a_n8300_8799.n48 a_n8300_8799.n191 0.365327
R401 a_n8300_8799.n189 a_n8300_8799.n51 21.4216
R402 a_n8300_8799.n59 a_n8300_8799.n207 0.365327
R403 a_n8300_8799.n205 a_n8300_8799.n62 21.4216
R404 a_n8300_8799.n70 a_n8300_8799.n224 0.365327
R405 a_n8300_8799.n222 a_n8300_8799.n73 21.4216
R406 a_n8300_8799.n139 a_n8300_8799.n80 0.365327
R407 a_n8300_8799.n83 a_n8300_8799.n141 21.4216
R408 a_n8300_8799.n155 a_n8300_8799.n91 0.365327
R409 a_n8300_8799.n94 a_n8300_8799.n157 21.4216
R410 a_n8300_8799.n172 a_n8300_8799.n102 0.365327
R411 a_n8300_8799.n105 a_n8300_8799.n174 21.4216
R412 a_n8300_8799.n37 a_n8300_8799.n38 1.43153
R413 a_n8300_8799.n31 a_n8300_8799.n30 1.13686
R414 a_n8300_8799.n25 a_n8300_8799.n24 1.13686
R415 a_n8300_8799.n19 a_n8300_8799.n18 1.13686
R416 a_n8300_8799.n13 a_n8300_8799.n12 1.13686
R417 a_n8300_8799.n7 a_n8300_8799.n6 1.13686
R418 a_n8300_8799.n1 a_n8300_8799.n0 1.13686
R419 a_n8300_8799.n42 a_n8300_8799.n41 1.07378
R420 a_n8300_8799.n40 a_n8300_8799.n39 1.07378
R421 a_n8300_8799.n36 a_n8300_8799.n43 1.07378
R422 a_n8300_8799.n35 a_n8300_8799.n34 0.758076
R423 a_n8300_8799.n32 a_n8300_8799.n34 0.758076
R424 a_n8300_8799.n33 a_n8300_8799.n32 0.758076
R425 a_n8300_8799.n33 a_n8300_8799.n31 0.758076
R426 a_n8300_8799.n29 a_n8300_8799.n28 0.758076
R427 a_n8300_8799.n26 a_n8300_8799.n28 0.758076
R428 a_n8300_8799.n27 a_n8300_8799.n26 0.758076
R429 a_n8300_8799.n27 a_n8300_8799.n25 0.758076
R430 a_n8300_8799.n23 a_n8300_8799.n22 0.758076
R431 a_n8300_8799.n20 a_n8300_8799.n22 0.758076
R432 a_n8300_8799.n21 a_n8300_8799.n20 0.758076
R433 a_n8300_8799.n21 a_n8300_8799.n19 0.758076
R434 a_n8300_8799.n16 a_n8300_8799.n17 0.758076
R435 a_n8300_8799.n15 a_n8300_8799.n16 0.758076
R436 a_n8300_8799.n14 a_n8300_8799.n15 0.758076
R437 a_n8300_8799.n12 a_n8300_8799.n14 0.758076
R438 a_n8300_8799.n10 a_n8300_8799.n11 0.758076
R439 a_n8300_8799.n9 a_n8300_8799.n10 0.758076
R440 a_n8300_8799.n8 a_n8300_8799.n9 0.758076
R441 a_n8300_8799.n6 a_n8300_8799.n8 0.758076
R442 a_n8300_8799.n4 a_n8300_8799.n5 0.758076
R443 a_n8300_8799.n3 a_n8300_8799.n4 0.758076
R444 a_n8300_8799.n2 a_n8300_8799.n3 0.758076
R445 a_n8300_8799.n0 a_n8300_8799.n2 0.758076
R446 vdd.n315 vdd.n279 756.745
R447 vdd.n260 vdd.n224 756.745
R448 vdd.n217 vdd.n181 756.745
R449 vdd.n162 vdd.n126 756.745
R450 vdd.n120 vdd.n84 756.745
R451 vdd.n65 vdd.n29 756.745
R452 vdd.n1764 vdd.n1728 756.745
R453 vdd.n1819 vdd.n1783 756.745
R454 vdd.n1666 vdd.n1630 756.745
R455 vdd.n1721 vdd.n1685 756.745
R456 vdd.n1569 vdd.n1533 756.745
R457 vdd.n1624 vdd.n1588 756.745
R458 vdd.n1107 vdd.t43 640.208
R459 vdd.n968 vdd.t81 640.208
R460 vdd.n1101 vdd.t108 640.208
R461 vdd.n959 vdd.t105 640.208
R462 vdd.n856 vdd.t54 640.208
R463 vdd.n2678 vdd.t99 640.208
R464 vdd.n804 vdd.t75 640.208
R465 vdd.n2747 vdd.t85 640.208
R466 vdd.n768 vdd.t39 640.208
R467 vdd.n1029 vdd.t95 640.208
R468 vdd.n1228 vdd.t68 592.009
R469 vdd.n1384 vdd.t92 592.009
R470 vdd.n1420 vdd.t102 592.009
R471 vdd.n2117 vdd.t61 592.009
R472 vdd.n1967 vdd.t78 592.009
R473 vdd.n1927 vdd.t89 592.009
R474 vdd.n405 vdd.t65 592.009
R475 vdd.n419 vdd.t50 592.009
R476 vdd.n431 vdd.t72 592.009
R477 vdd.n723 vdd.t35 592.009
R478 vdd.n686 vdd.t47 592.009
R479 vdd.n3195 vdd.t58 592.009
R480 vdd.n316 vdd.n315 585
R481 vdd.n314 vdd.n281 585
R482 vdd.n313 vdd.n312 585
R483 vdd.n284 vdd.n282 585
R484 vdd.n307 vdd.n306 585
R485 vdd.n305 vdd.n304 585
R486 vdd.n288 vdd.n287 585
R487 vdd.n299 vdd.n298 585
R488 vdd.n297 vdd.n296 585
R489 vdd.n292 vdd.n291 585
R490 vdd.n261 vdd.n260 585
R491 vdd.n259 vdd.n226 585
R492 vdd.n258 vdd.n257 585
R493 vdd.n229 vdd.n227 585
R494 vdd.n252 vdd.n251 585
R495 vdd.n250 vdd.n249 585
R496 vdd.n233 vdd.n232 585
R497 vdd.n244 vdd.n243 585
R498 vdd.n242 vdd.n241 585
R499 vdd.n237 vdd.n236 585
R500 vdd.n218 vdd.n217 585
R501 vdd.n216 vdd.n183 585
R502 vdd.n215 vdd.n214 585
R503 vdd.n186 vdd.n184 585
R504 vdd.n209 vdd.n208 585
R505 vdd.n207 vdd.n206 585
R506 vdd.n190 vdd.n189 585
R507 vdd.n201 vdd.n200 585
R508 vdd.n199 vdd.n198 585
R509 vdd.n194 vdd.n193 585
R510 vdd.n163 vdd.n162 585
R511 vdd.n161 vdd.n128 585
R512 vdd.n160 vdd.n159 585
R513 vdd.n131 vdd.n129 585
R514 vdd.n154 vdd.n153 585
R515 vdd.n152 vdd.n151 585
R516 vdd.n135 vdd.n134 585
R517 vdd.n146 vdd.n145 585
R518 vdd.n144 vdd.n143 585
R519 vdd.n139 vdd.n138 585
R520 vdd.n121 vdd.n120 585
R521 vdd.n119 vdd.n86 585
R522 vdd.n118 vdd.n117 585
R523 vdd.n89 vdd.n87 585
R524 vdd.n112 vdd.n111 585
R525 vdd.n110 vdd.n109 585
R526 vdd.n93 vdd.n92 585
R527 vdd.n104 vdd.n103 585
R528 vdd.n102 vdd.n101 585
R529 vdd.n97 vdd.n96 585
R530 vdd.n66 vdd.n65 585
R531 vdd.n64 vdd.n31 585
R532 vdd.n63 vdd.n62 585
R533 vdd.n34 vdd.n32 585
R534 vdd.n57 vdd.n56 585
R535 vdd.n55 vdd.n54 585
R536 vdd.n38 vdd.n37 585
R537 vdd.n49 vdd.n48 585
R538 vdd.n47 vdd.n46 585
R539 vdd.n42 vdd.n41 585
R540 vdd.n1765 vdd.n1764 585
R541 vdd.n1763 vdd.n1730 585
R542 vdd.n1762 vdd.n1761 585
R543 vdd.n1733 vdd.n1731 585
R544 vdd.n1756 vdd.n1755 585
R545 vdd.n1754 vdd.n1753 585
R546 vdd.n1737 vdd.n1736 585
R547 vdd.n1748 vdd.n1747 585
R548 vdd.n1746 vdd.n1745 585
R549 vdd.n1741 vdd.n1740 585
R550 vdd.n1820 vdd.n1819 585
R551 vdd.n1818 vdd.n1785 585
R552 vdd.n1817 vdd.n1816 585
R553 vdd.n1788 vdd.n1786 585
R554 vdd.n1811 vdd.n1810 585
R555 vdd.n1809 vdd.n1808 585
R556 vdd.n1792 vdd.n1791 585
R557 vdd.n1803 vdd.n1802 585
R558 vdd.n1801 vdd.n1800 585
R559 vdd.n1796 vdd.n1795 585
R560 vdd.n1667 vdd.n1666 585
R561 vdd.n1665 vdd.n1632 585
R562 vdd.n1664 vdd.n1663 585
R563 vdd.n1635 vdd.n1633 585
R564 vdd.n1658 vdd.n1657 585
R565 vdd.n1656 vdd.n1655 585
R566 vdd.n1639 vdd.n1638 585
R567 vdd.n1650 vdd.n1649 585
R568 vdd.n1648 vdd.n1647 585
R569 vdd.n1643 vdd.n1642 585
R570 vdd.n1722 vdd.n1721 585
R571 vdd.n1720 vdd.n1687 585
R572 vdd.n1719 vdd.n1718 585
R573 vdd.n1690 vdd.n1688 585
R574 vdd.n1713 vdd.n1712 585
R575 vdd.n1711 vdd.n1710 585
R576 vdd.n1694 vdd.n1693 585
R577 vdd.n1705 vdd.n1704 585
R578 vdd.n1703 vdd.n1702 585
R579 vdd.n1698 vdd.n1697 585
R580 vdd.n1570 vdd.n1569 585
R581 vdd.n1568 vdd.n1535 585
R582 vdd.n1567 vdd.n1566 585
R583 vdd.n1538 vdd.n1536 585
R584 vdd.n1561 vdd.n1560 585
R585 vdd.n1559 vdd.n1558 585
R586 vdd.n1542 vdd.n1541 585
R587 vdd.n1553 vdd.n1552 585
R588 vdd.n1551 vdd.n1550 585
R589 vdd.n1546 vdd.n1545 585
R590 vdd.n1625 vdd.n1624 585
R591 vdd.n1623 vdd.n1590 585
R592 vdd.n1622 vdd.n1621 585
R593 vdd.n1593 vdd.n1591 585
R594 vdd.n1616 vdd.n1615 585
R595 vdd.n1614 vdd.n1613 585
R596 vdd.n1597 vdd.n1596 585
R597 vdd.n1608 vdd.n1607 585
R598 vdd.n1606 vdd.n1605 585
R599 vdd.n1601 vdd.n1600 585
R600 vdd.n445 vdd.n370 462.44
R601 vdd.n3433 vdd.n372 462.44
R602 vdd.n3328 vdd.n657 462.44
R603 vdd.n3326 vdd.n660 462.44
R604 vdd.n2112 vdd.n1127 462.44
R605 vdd.n2115 vdd.n2114 462.44
R606 vdd.n1455 vdd.n1225 462.44
R607 vdd.n1452 vdd.n1223 462.44
R608 vdd.n293 vdd.t148 329.043
R609 vdd.n238 vdd.t199 329.043
R610 vdd.n195 vdd.t255 329.043
R611 vdd.n140 vdd.t183 329.043
R612 vdd.n98 vdd.t178 329.043
R613 vdd.n43 vdd.t239 329.043
R614 vdd.n1742 vdd.t257 329.043
R615 vdd.n1797 vdd.t197 329.043
R616 vdd.n1644 vdd.t249 329.043
R617 vdd.n1699 vdd.t179 329.043
R618 vdd.n1547 vdd.t215 329.043
R619 vdd.n1602 vdd.t177 329.043
R620 vdd.n1228 vdd.t71 319.788
R621 vdd.n1384 vdd.t94 319.788
R622 vdd.n1420 vdd.t104 319.788
R623 vdd.n2117 vdd.t63 319.788
R624 vdd.n1967 vdd.t79 319.788
R625 vdd.n1927 vdd.t90 319.788
R626 vdd.n405 vdd.t66 319.788
R627 vdd.n419 vdd.t52 319.788
R628 vdd.n431 vdd.t73 319.788
R629 vdd.n723 vdd.t38 319.788
R630 vdd.n686 vdd.t49 319.788
R631 vdd.n3195 vdd.t60 319.788
R632 vdd.n1229 vdd.t70 303.69
R633 vdd.n1385 vdd.t93 303.69
R634 vdd.n1421 vdd.t103 303.69
R635 vdd.n2118 vdd.t64 303.69
R636 vdd.n1968 vdd.t80 303.69
R637 vdd.n1928 vdd.t91 303.69
R638 vdd.n406 vdd.t67 303.69
R639 vdd.n420 vdd.t53 303.69
R640 vdd.n432 vdd.t74 303.69
R641 vdd.n724 vdd.t37 303.69
R642 vdd.n687 vdd.t48 303.69
R643 vdd.n3196 vdd.t59 303.69
R644 vdd.n2933 vdd.n918 285.366
R645 vdd.n3157 vdd.n778 285.366
R646 vdd.n3094 vdd.n775 285.366
R647 vdd.n2812 vdd.n915 285.366
R648 vdd.n2642 vdd.n956 285.366
R649 vdd.n2573 vdd.n2572 285.366
R650 vdd.n2313 vdd.n1082 285.366
R651 vdd.n2383 vdd.n1084 285.366
R652 vdd.n3073 vdd.n776 285.366
R653 vdd.n3160 vdd.n3159 285.366
R654 vdd.n2926 vdd.n916 285.366
R655 vdd.n2935 vdd.n914 285.366
R656 vdd.n2570 vdd.n966 285.366
R657 vdd.n964 vdd.n938 285.366
R658 vdd.n2199 vdd.n1083 285.366
R659 vdd.n2385 vdd.n1080 285.366
R660 vdd.n1125 vdd.n1081 216.982
R661 vdd.n756 vdd.n658 216.982
R662 vdd.n3075 vdd.n776 185
R663 vdd.n3158 vdd.n776 185
R664 vdd.n3077 vdd.n3076 185
R665 vdd.n3076 vdd.n774 185
R666 vdd.n3078 vdd.n810 185
R667 vdd.n3088 vdd.n810 185
R668 vdd.n3079 vdd.n819 185
R669 vdd.n819 vdd.n817 185
R670 vdd.n3081 vdd.n3080 185
R671 vdd.n3082 vdd.n3081 185
R672 vdd.n3034 vdd.n818 185
R673 vdd.n818 vdd.n814 185
R674 vdd.n3033 vdd.n3032 185
R675 vdd.n3032 vdd.n3031 185
R676 vdd.n821 vdd.n820 185
R677 vdd.n822 vdd.n821 185
R678 vdd.n3024 vdd.n3023 185
R679 vdd.n3025 vdd.n3024 185
R680 vdd.n3022 vdd.n830 185
R681 vdd.n835 vdd.n830 185
R682 vdd.n3021 vdd.n3020 185
R683 vdd.n3020 vdd.n3019 185
R684 vdd.n832 vdd.n831 185
R685 vdd.n841 vdd.n832 185
R686 vdd.n3012 vdd.n3011 185
R687 vdd.n3013 vdd.n3012 185
R688 vdd.n3010 vdd.n842 185
R689 vdd.n848 vdd.n842 185
R690 vdd.n3009 vdd.n3008 185
R691 vdd.n3008 vdd.n3007 185
R692 vdd.n844 vdd.n843 185
R693 vdd.n845 vdd.n844 185
R694 vdd.n3000 vdd.n2999 185
R695 vdd.n3001 vdd.n3000 185
R696 vdd.n2998 vdd.n855 185
R697 vdd.n855 vdd.n852 185
R698 vdd.n2996 vdd.n2995 185
R699 vdd.n2995 vdd.n2994 185
R700 vdd.n858 vdd.n857 185
R701 vdd.n859 vdd.n858 185
R702 vdd.n2987 vdd.n2986 185
R703 vdd.n2988 vdd.n2987 185
R704 vdd.n2985 vdd.n867 185
R705 vdd.n872 vdd.n867 185
R706 vdd.n2984 vdd.n2983 185
R707 vdd.n2983 vdd.n2982 185
R708 vdd.n869 vdd.n868 185
R709 vdd.n2894 vdd.n869 185
R710 vdd.n2975 vdd.n2974 185
R711 vdd.n2976 vdd.n2975 185
R712 vdd.n2973 vdd.n879 185
R713 vdd.n879 vdd.n876 185
R714 vdd.n2972 vdd.n2971 185
R715 vdd.n2971 vdd.n2970 185
R716 vdd.n881 vdd.n880 185
R717 vdd.n882 vdd.n881 185
R718 vdd.n2963 vdd.n2962 185
R719 vdd.n2964 vdd.n2963 185
R720 vdd.n2961 vdd.n890 185
R721 vdd.n2906 vdd.n890 185
R722 vdd.n2960 vdd.n2959 185
R723 vdd.n2959 vdd.n2958 185
R724 vdd.n892 vdd.n891 185
R725 vdd.n901 vdd.n892 185
R726 vdd.n2951 vdd.n2950 185
R727 vdd.n2952 vdd.n2951 185
R728 vdd.n2949 vdd.n902 185
R729 vdd.n902 vdd.n898 185
R730 vdd.n2948 vdd.n2947 185
R731 vdd.n2947 vdd.n2946 185
R732 vdd.n904 vdd.n903 185
R733 vdd.n2918 vdd.n904 185
R734 vdd.n2939 vdd.n2938 185
R735 vdd.n2940 vdd.n2939 185
R736 vdd.n2937 vdd.n912 185
R737 vdd.n917 vdd.n912 185
R738 vdd.n2936 vdd.n2935 185
R739 vdd.n2935 vdd.n2934 185
R740 vdd.n914 vdd.n913 185
R741 vdd.n2682 vdd.n2681 185
R742 vdd.n2684 vdd.n2683 185
R743 vdd.n2686 vdd.n2685 185
R744 vdd.n2688 vdd.n2687 185
R745 vdd.n2690 vdd.n2689 185
R746 vdd.n2692 vdd.n2691 185
R747 vdd.n2694 vdd.n2693 185
R748 vdd.n2696 vdd.n2695 185
R749 vdd.n2698 vdd.n2697 185
R750 vdd.n2700 vdd.n2699 185
R751 vdd.n2702 vdd.n2701 185
R752 vdd.n2704 vdd.n2703 185
R753 vdd.n2706 vdd.n2705 185
R754 vdd.n2708 vdd.n2707 185
R755 vdd.n2710 vdd.n2709 185
R756 vdd.n2712 vdd.n2711 185
R757 vdd.n2714 vdd.n2713 185
R758 vdd.n2716 vdd.n2715 185
R759 vdd.n2718 vdd.n2717 185
R760 vdd.n2720 vdd.n2719 185
R761 vdd.n2722 vdd.n2721 185
R762 vdd.n2724 vdd.n2723 185
R763 vdd.n2726 vdd.n2725 185
R764 vdd.n2728 vdd.n2727 185
R765 vdd.n2730 vdd.n2729 185
R766 vdd.n2732 vdd.n2731 185
R767 vdd.n2734 vdd.n2733 185
R768 vdd.n2736 vdd.n2735 185
R769 vdd.n2738 vdd.n2737 185
R770 vdd.n2740 vdd.n2739 185
R771 vdd.n2742 vdd.n2741 185
R772 vdd.n2744 vdd.n2743 185
R773 vdd.n2745 vdd.n2677 185
R774 vdd.n2926 vdd.n2925 185
R775 vdd.n2927 vdd.n2926 185
R776 vdd.n3161 vdd.n3160 185
R777 vdd.n3162 vdd.n767 185
R778 vdd.n3164 vdd.n3163 185
R779 vdd.n3166 vdd.n765 185
R780 vdd.n3168 vdd.n3167 185
R781 vdd.n3169 vdd.n764 185
R782 vdd.n3171 vdd.n3170 185
R783 vdd.n3173 vdd.n762 185
R784 vdd.n3175 vdd.n3174 185
R785 vdd.n3176 vdd.n761 185
R786 vdd.n3178 vdd.n3177 185
R787 vdd.n3180 vdd.n759 185
R788 vdd.n3182 vdd.n3181 185
R789 vdd.n3183 vdd.n758 185
R790 vdd.n3185 vdd.n3184 185
R791 vdd.n3187 vdd.n757 185
R792 vdd.n3188 vdd.n754 185
R793 vdd.n3191 vdd.n3190 185
R794 vdd.n755 vdd.n753 185
R795 vdd.n3047 vdd.n3046 185
R796 vdd.n3049 vdd.n3048 185
R797 vdd.n3051 vdd.n3043 185
R798 vdd.n3053 vdd.n3052 185
R799 vdd.n3054 vdd.n3042 185
R800 vdd.n3056 vdd.n3055 185
R801 vdd.n3058 vdd.n3040 185
R802 vdd.n3060 vdd.n3059 185
R803 vdd.n3061 vdd.n3039 185
R804 vdd.n3063 vdd.n3062 185
R805 vdd.n3065 vdd.n3037 185
R806 vdd.n3067 vdd.n3066 185
R807 vdd.n3068 vdd.n3036 185
R808 vdd.n3070 vdd.n3069 185
R809 vdd.n3072 vdd.n3035 185
R810 vdd.n3074 vdd.n3073 185
R811 vdd.n3073 vdd.n756 185
R812 vdd.n3159 vdd.n771 185
R813 vdd.n3159 vdd.n3158 185
R814 vdd.n2825 vdd.n773 185
R815 vdd.n774 vdd.n773 185
R816 vdd.n2826 vdd.n809 185
R817 vdd.n3088 vdd.n809 185
R818 vdd.n2828 vdd.n2827 185
R819 vdd.n2827 vdd.n817 185
R820 vdd.n2829 vdd.n816 185
R821 vdd.n3082 vdd.n816 185
R822 vdd.n2831 vdd.n2830 185
R823 vdd.n2830 vdd.n814 185
R824 vdd.n2832 vdd.n824 185
R825 vdd.n3031 vdd.n824 185
R826 vdd.n2834 vdd.n2833 185
R827 vdd.n2833 vdd.n822 185
R828 vdd.n2835 vdd.n829 185
R829 vdd.n3025 vdd.n829 185
R830 vdd.n2837 vdd.n2836 185
R831 vdd.n2836 vdd.n835 185
R832 vdd.n2838 vdd.n834 185
R833 vdd.n3019 vdd.n834 185
R834 vdd.n2840 vdd.n2839 185
R835 vdd.n2839 vdd.n841 185
R836 vdd.n2841 vdd.n840 185
R837 vdd.n3013 vdd.n840 185
R838 vdd.n2843 vdd.n2842 185
R839 vdd.n2842 vdd.n848 185
R840 vdd.n2844 vdd.n847 185
R841 vdd.n3007 vdd.n847 185
R842 vdd.n2846 vdd.n2845 185
R843 vdd.n2845 vdd.n845 185
R844 vdd.n2847 vdd.n854 185
R845 vdd.n3001 vdd.n854 185
R846 vdd.n2849 vdd.n2848 185
R847 vdd.n2848 vdd.n852 185
R848 vdd.n2850 vdd.n861 185
R849 vdd.n2994 vdd.n861 185
R850 vdd.n2852 vdd.n2851 185
R851 vdd.n2851 vdd.n859 185
R852 vdd.n2853 vdd.n866 185
R853 vdd.n2988 vdd.n866 185
R854 vdd.n2855 vdd.n2854 185
R855 vdd.n2854 vdd.n872 185
R856 vdd.n2856 vdd.n871 185
R857 vdd.n2982 vdd.n871 185
R858 vdd.n2896 vdd.n2895 185
R859 vdd.n2895 vdd.n2894 185
R860 vdd.n2897 vdd.n878 185
R861 vdd.n2976 vdd.n878 185
R862 vdd.n2899 vdd.n2898 185
R863 vdd.n2898 vdd.n876 185
R864 vdd.n2900 vdd.n884 185
R865 vdd.n2970 vdd.n884 185
R866 vdd.n2902 vdd.n2901 185
R867 vdd.n2901 vdd.n882 185
R868 vdd.n2903 vdd.n889 185
R869 vdd.n2964 vdd.n889 185
R870 vdd.n2905 vdd.n2904 185
R871 vdd.n2906 vdd.n2905 185
R872 vdd.n2824 vdd.n894 185
R873 vdd.n2958 vdd.n894 185
R874 vdd.n2823 vdd.n2822 185
R875 vdd.n2822 vdd.n901 185
R876 vdd.n2821 vdd.n900 185
R877 vdd.n2952 vdd.n900 185
R878 vdd.n2820 vdd.n2819 185
R879 vdd.n2819 vdd.n898 185
R880 vdd.n2746 vdd.n906 185
R881 vdd.n2946 vdd.n906 185
R882 vdd.n2920 vdd.n2919 185
R883 vdd.n2919 vdd.n2918 185
R884 vdd.n2921 vdd.n911 185
R885 vdd.n2940 vdd.n911 185
R886 vdd.n2923 vdd.n2922 185
R887 vdd.n2922 vdd.n917 185
R888 vdd.n2924 vdd.n916 185
R889 vdd.n2934 vdd.n916 185
R890 vdd.n2112 vdd.n2111 185
R891 vdd.n2113 vdd.n2112 185
R892 vdd.n1128 vdd.n1126 185
R893 vdd.n1126 vdd.n1124 185
R894 vdd.n1894 vdd.n1893 185
R895 vdd.n1893 vdd.n1892 185
R896 vdd.n1131 vdd.n1130 185
R897 vdd.n1132 vdd.n1131 185
R898 vdd.n1881 vdd.n1880 185
R899 vdd.n1882 vdd.n1881 185
R900 vdd.n1140 vdd.n1139 185
R901 vdd.n1873 vdd.n1139 185
R902 vdd.n1876 vdd.n1875 185
R903 vdd.n1875 vdd.n1874 185
R904 vdd.n1143 vdd.n1142 185
R905 vdd.n1149 vdd.n1143 185
R906 vdd.n1864 vdd.n1863 185
R907 vdd.n1865 vdd.n1864 185
R908 vdd.n1151 vdd.n1150 185
R909 vdd.n1856 vdd.n1150 185
R910 vdd.n1859 vdd.n1858 185
R911 vdd.n1858 vdd.n1857 185
R912 vdd.n1154 vdd.n1153 185
R913 vdd.n1155 vdd.n1154 185
R914 vdd.n1847 vdd.n1846 185
R915 vdd.n1848 vdd.n1847 185
R916 vdd.n1163 vdd.n1162 185
R917 vdd.n1162 vdd.n1161 185
R918 vdd.n1842 vdd.n1841 185
R919 vdd.n1841 vdd.n1840 185
R920 vdd.n1166 vdd.n1165 185
R921 vdd.n1172 vdd.n1166 185
R922 vdd.n1831 vdd.n1830 185
R923 vdd.n1832 vdd.n1831 185
R924 vdd.n1174 vdd.n1173 185
R925 vdd.n1528 vdd.n1173 185
R926 vdd.n1531 vdd.n1530 185
R927 vdd.n1530 vdd.n1529 185
R928 vdd.n1177 vdd.n1176 185
R929 vdd.n1184 vdd.n1177 185
R930 vdd.n1519 vdd.n1518 185
R931 vdd.n1520 vdd.n1519 185
R932 vdd.n1186 vdd.n1185 185
R933 vdd.n1185 vdd.n1183 185
R934 vdd.n1514 vdd.n1513 185
R935 vdd.n1513 vdd.n1512 185
R936 vdd.n1189 vdd.n1188 185
R937 vdd.n1190 vdd.n1189 185
R938 vdd.n1503 vdd.n1502 185
R939 vdd.n1504 vdd.n1503 185
R940 vdd.n1197 vdd.n1196 185
R941 vdd.n1495 vdd.n1196 185
R942 vdd.n1498 vdd.n1497 185
R943 vdd.n1497 vdd.n1496 185
R944 vdd.n1200 vdd.n1199 185
R945 vdd.n1206 vdd.n1200 185
R946 vdd.n1486 vdd.n1485 185
R947 vdd.n1487 vdd.n1486 185
R948 vdd.n1208 vdd.n1207 185
R949 vdd.n1478 vdd.n1207 185
R950 vdd.n1481 vdd.n1480 185
R951 vdd.n1480 vdd.n1479 185
R952 vdd.n1211 vdd.n1210 185
R953 vdd.n1212 vdd.n1211 185
R954 vdd.n1469 vdd.n1468 185
R955 vdd.n1470 vdd.n1469 185
R956 vdd.n1220 vdd.n1219 185
R957 vdd.n1219 vdd.n1218 185
R958 vdd.n1464 vdd.n1463 185
R959 vdd.n1463 vdd.n1462 185
R960 vdd.n1223 vdd.n1222 185
R961 vdd.n1224 vdd.n1223 185
R962 vdd.n1452 vdd.n1451 185
R963 vdd.n1450 vdd.n1263 185
R964 vdd.n1265 vdd.n1262 185
R965 vdd.n1454 vdd.n1262 185
R966 vdd.n1446 vdd.n1267 185
R967 vdd.n1445 vdd.n1268 185
R968 vdd.n1444 vdd.n1269 185
R969 vdd.n1272 vdd.n1270 185
R970 vdd.n1440 vdd.n1273 185
R971 vdd.n1439 vdd.n1274 185
R972 vdd.n1438 vdd.n1275 185
R973 vdd.n1278 vdd.n1276 185
R974 vdd.n1434 vdd.n1279 185
R975 vdd.n1433 vdd.n1280 185
R976 vdd.n1432 vdd.n1281 185
R977 vdd.n1284 vdd.n1282 185
R978 vdd.n1428 vdd.n1285 185
R979 vdd.n1427 vdd.n1286 185
R980 vdd.n1426 vdd.n1287 185
R981 vdd.n1418 vdd.n1288 185
R982 vdd.n1422 vdd.n1419 185
R983 vdd.n1417 vdd.n1290 185
R984 vdd.n1416 vdd.n1291 185
R985 vdd.n1294 vdd.n1292 185
R986 vdd.n1412 vdd.n1295 185
R987 vdd.n1411 vdd.n1296 185
R988 vdd.n1410 vdd.n1297 185
R989 vdd.n1300 vdd.n1298 185
R990 vdd.n1406 vdd.n1301 185
R991 vdd.n1405 vdd.n1302 185
R992 vdd.n1404 vdd.n1303 185
R993 vdd.n1306 vdd.n1304 185
R994 vdd.n1400 vdd.n1307 185
R995 vdd.n1399 vdd.n1308 185
R996 vdd.n1398 vdd.n1309 185
R997 vdd.n1312 vdd.n1310 185
R998 vdd.n1394 vdd.n1313 185
R999 vdd.n1393 vdd.n1314 185
R1000 vdd.n1392 vdd.n1315 185
R1001 vdd.n1318 vdd.n1316 185
R1002 vdd.n1388 vdd.n1319 185
R1003 vdd.n1387 vdd.n1320 185
R1004 vdd.n1386 vdd.n1383 185
R1005 vdd.n1323 vdd.n1321 185
R1006 vdd.n1379 vdd.n1324 185
R1007 vdd.n1378 vdd.n1325 185
R1008 vdd.n1377 vdd.n1326 185
R1009 vdd.n1329 vdd.n1327 185
R1010 vdd.n1373 vdd.n1330 185
R1011 vdd.n1372 vdd.n1331 185
R1012 vdd.n1371 vdd.n1332 185
R1013 vdd.n1335 vdd.n1333 185
R1014 vdd.n1367 vdd.n1336 185
R1015 vdd.n1366 vdd.n1337 185
R1016 vdd.n1365 vdd.n1338 185
R1017 vdd.n1341 vdd.n1339 185
R1018 vdd.n1361 vdd.n1342 185
R1019 vdd.n1360 vdd.n1343 185
R1020 vdd.n1359 vdd.n1344 185
R1021 vdd.n1347 vdd.n1345 185
R1022 vdd.n1355 vdd.n1348 185
R1023 vdd.n1354 vdd.n1349 185
R1024 vdd.n1353 vdd.n1350 185
R1025 vdd.n1351 vdd.n1231 185
R1026 vdd.n1456 vdd.n1455 185
R1027 vdd.n1455 vdd.n1454 185
R1028 vdd.n2116 vdd.n2115 185
R1029 vdd.n2120 vdd.n1120 185
R1030 vdd.n1996 vdd.n1119 185
R1031 vdd.n1999 vdd.n1998 185
R1032 vdd.n2001 vdd.n2000 185
R1033 vdd.n2004 vdd.n2003 185
R1034 vdd.n2006 vdd.n2005 185
R1035 vdd.n2008 vdd.n1994 185
R1036 vdd.n2010 vdd.n2009 185
R1037 vdd.n2011 vdd.n1988 185
R1038 vdd.n2013 vdd.n2012 185
R1039 vdd.n2015 vdd.n1986 185
R1040 vdd.n2017 vdd.n2016 185
R1041 vdd.n2018 vdd.n1981 185
R1042 vdd.n2020 vdd.n2019 185
R1043 vdd.n2022 vdd.n1979 185
R1044 vdd.n2024 vdd.n2023 185
R1045 vdd.n2025 vdd.n1975 185
R1046 vdd.n2027 vdd.n2026 185
R1047 vdd.n2029 vdd.n1972 185
R1048 vdd.n2031 vdd.n2030 185
R1049 vdd.n1973 vdd.n1966 185
R1050 vdd.n2035 vdd.n1970 185
R1051 vdd.n2036 vdd.n1962 185
R1052 vdd.n2038 vdd.n2037 185
R1053 vdd.n2040 vdd.n1960 185
R1054 vdd.n2042 vdd.n2041 185
R1055 vdd.n2043 vdd.n1955 185
R1056 vdd.n2045 vdd.n2044 185
R1057 vdd.n2047 vdd.n1953 185
R1058 vdd.n2049 vdd.n2048 185
R1059 vdd.n2050 vdd.n1948 185
R1060 vdd.n2052 vdd.n2051 185
R1061 vdd.n2054 vdd.n1946 185
R1062 vdd.n2056 vdd.n2055 185
R1063 vdd.n2057 vdd.n1941 185
R1064 vdd.n2059 vdd.n2058 185
R1065 vdd.n2061 vdd.n1939 185
R1066 vdd.n2063 vdd.n2062 185
R1067 vdd.n2064 vdd.n1935 185
R1068 vdd.n2066 vdd.n2065 185
R1069 vdd.n2068 vdd.n1932 185
R1070 vdd.n2070 vdd.n2069 185
R1071 vdd.n1933 vdd.n1926 185
R1072 vdd.n2074 vdd.n1930 185
R1073 vdd.n2075 vdd.n1922 185
R1074 vdd.n2077 vdd.n2076 185
R1075 vdd.n2079 vdd.n1920 185
R1076 vdd.n2081 vdd.n2080 185
R1077 vdd.n2082 vdd.n1915 185
R1078 vdd.n2084 vdd.n2083 185
R1079 vdd.n2086 vdd.n1913 185
R1080 vdd.n2088 vdd.n2087 185
R1081 vdd.n2089 vdd.n1908 185
R1082 vdd.n2091 vdd.n2090 185
R1083 vdd.n2093 vdd.n1907 185
R1084 vdd.n2094 vdd.n1904 185
R1085 vdd.n2097 vdd.n2096 185
R1086 vdd.n1906 vdd.n1902 185
R1087 vdd.n2101 vdd.n1900 185
R1088 vdd.n2103 vdd.n2102 185
R1089 vdd.n2105 vdd.n1898 185
R1090 vdd.n2107 vdd.n2106 185
R1091 vdd.n2108 vdd.n1127 185
R1092 vdd.n2114 vdd.n1123 185
R1093 vdd.n2114 vdd.n2113 185
R1094 vdd.n1135 vdd.n1122 185
R1095 vdd.n1124 vdd.n1122 185
R1096 vdd.n1891 vdd.n1890 185
R1097 vdd.n1892 vdd.n1891 185
R1098 vdd.n1134 vdd.n1133 185
R1099 vdd.n1133 vdd.n1132 185
R1100 vdd.n1884 vdd.n1883 185
R1101 vdd.n1883 vdd.n1882 185
R1102 vdd.n1138 vdd.n1137 185
R1103 vdd.n1873 vdd.n1138 185
R1104 vdd.n1872 vdd.n1871 185
R1105 vdd.n1874 vdd.n1872 185
R1106 vdd.n1145 vdd.n1144 185
R1107 vdd.n1149 vdd.n1144 185
R1108 vdd.n1867 vdd.n1866 185
R1109 vdd.n1866 vdd.n1865 185
R1110 vdd.n1148 vdd.n1147 185
R1111 vdd.n1856 vdd.n1148 185
R1112 vdd.n1855 vdd.n1854 185
R1113 vdd.n1857 vdd.n1855 185
R1114 vdd.n1157 vdd.n1156 185
R1115 vdd.n1156 vdd.n1155 185
R1116 vdd.n1850 vdd.n1849 185
R1117 vdd.n1849 vdd.n1848 185
R1118 vdd.n1160 vdd.n1159 185
R1119 vdd.n1161 vdd.n1160 185
R1120 vdd.n1839 vdd.n1838 185
R1121 vdd.n1840 vdd.n1839 185
R1122 vdd.n1168 vdd.n1167 185
R1123 vdd.n1172 vdd.n1167 185
R1124 vdd.n1834 vdd.n1833 185
R1125 vdd.n1833 vdd.n1832 185
R1126 vdd.n1171 vdd.n1170 185
R1127 vdd.n1528 vdd.n1171 185
R1128 vdd.n1527 vdd.n1526 185
R1129 vdd.n1529 vdd.n1527 185
R1130 vdd.n1179 vdd.n1178 185
R1131 vdd.n1184 vdd.n1178 185
R1132 vdd.n1522 vdd.n1521 185
R1133 vdd.n1521 vdd.n1520 185
R1134 vdd.n1182 vdd.n1181 185
R1135 vdd.n1183 vdd.n1182 185
R1136 vdd.n1511 vdd.n1510 185
R1137 vdd.n1512 vdd.n1511 185
R1138 vdd.n1192 vdd.n1191 185
R1139 vdd.n1191 vdd.n1190 185
R1140 vdd.n1506 vdd.n1505 185
R1141 vdd.n1505 vdd.n1504 185
R1142 vdd.n1195 vdd.n1194 185
R1143 vdd.n1495 vdd.n1195 185
R1144 vdd.n1494 vdd.n1493 185
R1145 vdd.n1496 vdd.n1494 185
R1146 vdd.n1202 vdd.n1201 185
R1147 vdd.n1206 vdd.n1201 185
R1148 vdd.n1489 vdd.n1488 185
R1149 vdd.n1488 vdd.n1487 185
R1150 vdd.n1205 vdd.n1204 185
R1151 vdd.n1478 vdd.n1205 185
R1152 vdd.n1477 vdd.n1476 185
R1153 vdd.n1479 vdd.n1477 185
R1154 vdd.n1214 vdd.n1213 185
R1155 vdd.n1213 vdd.n1212 185
R1156 vdd.n1472 vdd.n1471 185
R1157 vdd.n1471 vdd.n1470 185
R1158 vdd.n1217 vdd.n1216 185
R1159 vdd.n1218 vdd.n1217 185
R1160 vdd.n1461 vdd.n1460 185
R1161 vdd.n1462 vdd.n1461 185
R1162 vdd.n1226 vdd.n1225 185
R1163 vdd.n1225 vdd.n1224 185
R1164 vdd.n958 vdd.n956 185
R1165 vdd.n2571 vdd.n956 185
R1166 vdd.n2493 vdd.n976 185
R1167 vdd.n976 vdd.n963 185
R1168 vdd.n2495 vdd.n2494 185
R1169 vdd.n2496 vdd.n2495 185
R1170 vdd.n2492 vdd.n975 185
R1171 vdd.n2251 vdd.n975 185
R1172 vdd.n2491 vdd.n2490 185
R1173 vdd.n2490 vdd.n2489 185
R1174 vdd.n978 vdd.n977 185
R1175 vdd.n979 vdd.n978 185
R1176 vdd.n2480 vdd.n2479 185
R1177 vdd.n2481 vdd.n2480 185
R1178 vdd.n2478 vdd.n989 185
R1179 vdd.n989 vdd.n986 185
R1180 vdd.n2477 vdd.n2476 185
R1181 vdd.n2476 vdd.n2475 185
R1182 vdd.n991 vdd.n990 185
R1183 vdd.n2263 vdd.n991 185
R1184 vdd.n2468 vdd.n2467 185
R1185 vdd.n2469 vdd.n2468 185
R1186 vdd.n2466 vdd.n999 185
R1187 vdd.n1004 vdd.n999 185
R1188 vdd.n2465 vdd.n2464 185
R1189 vdd.n2464 vdd.n2463 185
R1190 vdd.n1001 vdd.n1000 185
R1191 vdd.n1010 vdd.n1001 185
R1192 vdd.n2456 vdd.n2455 185
R1193 vdd.n2457 vdd.n2456 185
R1194 vdd.n2454 vdd.n1011 185
R1195 vdd.n2275 vdd.n1011 185
R1196 vdd.n2453 vdd.n2452 185
R1197 vdd.n2452 vdd.n2451 185
R1198 vdd.n1013 vdd.n1012 185
R1199 vdd.n1014 vdd.n1013 185
R1200 vdd.n2444 vdd.n2443 185
R1201 vdd.n2445 vdd.n2444 185
R1202 vdd.n2442 vdd.n1023 185
R1203 vdd.n1023 vdd.n1020 185
R1204 vdd.n2441 vdd.n2440 185
R1205 vdd.n2440 vdd.n2439 185
R1206 vdd.n1025 vdd.n1024 185
R1207 vdd.n1034 vdd.n1025 185
R1208 vdd.n2431 vdd.n2430 185
R1209 vdd.n2432 vdd.n2431 185
R1210 vdd.n2429 vdd.n1035 185
R1211 vdd.n1041 vdd.n1035 185
R1212 vdd.n2428 vdd.n2427 185
R1213 vdd.n2427 vdd.n2426 185
R1214 vdd.n1037 vdd.n1036 185
R1215 vdd.n1038 vdd.n1037 185
R1216 vdd.n2419 vdd.n2418 185
R1217 vdd.n2420 vdd.n2419 185
R1218 vdd.n2417 vdd.n1048 185
R1219 vdd.n1048 vdd.n1045 185
R1220 vdd.n2416 vdd.n2415 185
R1221 vdd.n2415 vdd.n2414 185
R1222 vdd.n1050 vdd.n1049 185
R1223 vdd.n1051 vdd.n1050 185
R1224 vdd.n2407 vdd.n2406 185
R1225 vdd.n2408 vdd.n2407 185
R1226 vdd.n2405 vdd.n1060 185
R1227 vdd.n1060 vdd.n1057 185
R1228 vdd.n2404 vdd.n2403 185
R1229 vdd.n2403 vdd.n2402 185
R1230 vdd.n1062 vdd.n1061 185
R1231 vdd.n1063 vdd.n1062 185
R1232 vdd.n2395 vdd.n2394 185
R1233 vdd.n2396 vdd.n2395 185
R1234 vdd.n2393 vdd.n1072 185
R1235 vdd.n1072 vdd.n1069 185
R1236 vdd.n2392 vdd.n2391 185
R1237 vdd.n2391 vdd.n2390 185
R1238 vdd.n1074 vdd.n1073 185
R1239 vdd.n1075 vdd.n1074 185
R1240 vdd.n2383 vdd.n2382 185
R1241 vdd.n2384 vdd.n2383 185
R1242 vdd.n2381 vdd.n1084 185
R1243 vdd.n2380 vdd.n2379 185
R1244 vdd.n2377 vdd.n1085 185
R1245 vdd.n2377 vdd.n1081 185
R1246 vdd.n2376 vdd.n2375 185
R1247 vdd.n2374 vdd.n2373 185
R1248 vdd.n2372 vdd.n1087 185
R1249 vdd.n2370 vdd.n2369 185
R1250 vdd.n2368 vdd.n1088 185
R1251 vdd.n2367 vdd.n2366 185
R1252 vdd.n2364 vdd.n1089 185
R1253 vdd.n2362 vdd.n2361 185
R1254 vdd.n2360 vdd.n1090 185
R1255 vdd.n2359 vdd.n2358 185
R1256 vdd.n2356 vdd.n1091 185
R1257 vdd.n2354 vdd.n2353 185
R1258 vdd.n2352 vdd.n1092 185
R1259 vdd.n2351 vdd.n2350 185
R1260 vdd.n2348 vdd.n1093 185
R1261 vdd.n2346 vdd.n2345 185
R1262 vdd.n2344 vdd.n1094 185
R1263 vdd.n2343 vdd.n2342 185
R1264 vdd.n2340 vdd.n1095 185
R1265 vdd.n2338 vdd.n2337 185
R1266 vdd.n2336 vdd.n1096 185
R1267 vdd.n2335 vdd.n2334 185
R1268 vdd.n2332 vdd.n1097 185
R1269 vdd.n2330 vdd.n2329 185
R1270 vdd.n2328 vdd.n1098 185
R1271 vdd.n2327 vdd.n2326 185
R1272 vdd.n2324 vdd.n1099 185
R1273 vdd.n2322 vdd.n2321 185
R1274 vdd.n2320 vdd.n1100 185
R1275 vdd.n2318 vdd.n2317 185
R1276 vdd.n2315 vdd.n1103 185
R1277 vdd.n2313 vdd.n2312 185
R1278 vdd.n2574 vdd.n2573 185
R1279 vdd.n2576 vdd.n2575 185
R1280 vdd.n2578 vdd.n2577 185
R1281 vdd.n2581 vdd.n2580 185
R1282 vdd.n2583 vdd.n2582 185
R1283 vdd.n2585 vdd.n2584 185
R1284 vdd.n2587 vdd.n2586 185
R1285 vdd.n2589 vdd.n2588 185
R1286 vdd.n2591 vdd.n2590 185
R1287 vdd.n2593 vdd.n2592 185
R1288 vdd.n2595 vdd.n2594 185
R1289 vdd.n2597 vdd.n2596 185
R1290 vdd.n2599 vdd.n2598 185
R1291 vdd.n2601 vdd.n2600 185
R1292 vdd.n2603 vdd.n2602 185
R1293 vdd.n2605 vdd.n2604 185
R1294 vdd.n2607 vdd.n2606 185
R1295 vdd.n2609 vdd.n2608 185
R1296 vdd.n2611 vdd.n2610 185
R1297 vdd.n2613 vdd.n2612 185
R1298 vdd.n2615 vdd.n2614 185
R1299 vdd.n2617 vdd.n2616 185
R1300 vdd.n2619 vdd.n2618 185
R1301 vdd.n2621 vdd.n2620 185
R1302 vdd.n2623 vdd.n2622 185
R1303 vdd.n2625 vdd.n2624 185
R1304 vdd.n2627 vdd.n2626 185
R1305 vdd.n2629 vdd.n2628 185
R1306 vdd.n2631 vdd.n2630 185
R1307 vdd.n2633 vdd.n2632 185
R1308 vdd.n2635 vdd.n2634 185
R1309 vdd.n2637 vdd.n2636 185
R1310 vdd.n2639 vdd.n2638 185
R1311 vdd.n2640 vdd.n957 185
R1312 vdd.n2642 vdd.n2641 185
R1313 vdd.n2643 vdd.n2642 185
R1314 vdd.n2572 vdd.n961 185
R1315 vdd.n2572 vdd.n2571 185
R1316 vdd.n2249 vdd.n962 185
R1317 vdd.n963 vdd.n962 185
R1318 vdd.n2250 vdd.n973 185
R1319 vdd.n2496 vdd.n973 185
R1320 vdd.n2253 vdd.n2252 185
R1321 vdd.n2252 vdd.n2251 185
R1322 vdd.n2254 vdd.n980 185
R1323 vdd.n2489 vdd.n980 185
R1324 vdd.n2256 vdd.n2255 185
R1325 vdd.n2255 vdd.n979 185
R1326 vdd.n2257 vdd.n987 185
R1327 vdd.n2481 vdd.n987 185
R1328 vdd.n2259 vdd.n2258 185
R1329 vdd.n2258 vdd.n986 185
R1330 vdd.n2260 vdd.n992 185
R1331 vdd.n2475 vdd.n992 185
R1332 vdd.n2262 vdd.n2261 185
R1333 vdd.n2263 vdd.n2262 185
R1334 vdd.n2248 vdd.n997 185
R1335 vdd.n2469 vdd.n997 185
R1336 vdd.n2247 vdd.n2246 185
R1337 vdd.n2246 vdd.n1004 185
R1338 vdd.n2245 vdd.n1002 185
R1339 vdd.n2463 vdd.n1002 185
R1340 vdd.n2244 vdd.n2243 185
R1341 vdd.n2243 vdd.n1010 185
R1342 vdd.n1104 vdd.n1008 185
R1343 vdd.n2457 vdd.n1008 185
R1344 vdd.n2277 vdd.n2276 185
R1345 vdd.n2276 vdd.n2275 185
R1346 vdd.n2278 vdd.n1015 185
R1347 vdd.n2451 vdd.n1015 185
R1348 vdd.n2280 vdd.n2279 185
R1349 vdd.n2279 vdd.n1014 185
R1350 vdd.n2281 vdd.n1021 185
R1351 vdd.n2445 vdd.n1021 185
R1352 vdd.n2283 vdd.n2282 185
R1353 vdd.n2282 vdd.n1020 185
R1354 vdd.n2284 vdd.n1026 185
R1355 vdd.n2439 vdd.n1026 185
R1356 vdd.n2286 vdd.n2285 185
R1357 vdd.n2285 vdd.n1034 185
R1358 vdd.n2287 vdd.n1032 185
R1359 vdd.n2432 vdd.n1032 185
R1360 vdd.n2289 vdd.n2288 185
R1361 vdd.n2288 vdd.n1041 185
R1362 vdd.n2290 vdd.n1039 185
R1363 vdd.n2426 vdd.n1039 185
R1364 vdd.n2292 vdd.n2291 185
R1365 vdd.n2291 vdd.n1038 185
R1366 vdd.n2293 vdd.n1046 185
R1367 vdd.n2420 vdd.n1046 185
R1368 vdd.n2295 vdd.n2294 185
R1369 vdd.n2294 vdd.n1045 185
R1370 vdd.n2296 vdd.n1052 185
R1371 vdd.n2414 vdd.n1052 185
R1372 vdd.n2298 vdd.n2297 185
R1373 vdd.n2297 vdd.n1051 185
R1374 vdd.n2299 vdd.n1058 185
R1375 vdd.n2408 vdd.n1058 185
R1376 vdd.n2301 vdd.n2300 185
R1377 vdd.n2300 vdd.n1057 185
R1378 vdd.n2302 vdd.n1064 185
R1379 vdd.n2402 vdd.n1064 185
R1380 vdd.n2304 vdd.n2303 185
R1381 vdd.n2303 vdd.n1063 185
R1382 vdd.n2305 vdd.n1070 185
R1383 vdd.n2396 vdd.n1070 185
R1384 vdd.n2307 vdd.n2306 185
R1385 vdd.n2306 vdd.n1069 185
R1386 vdd.n2308 vdd.n1076 185
R1387 vdd.n2390 vdd.n1076 185
R1388 vdd.n2310 vdd.n2309 185
R1389 vdd.n2309 vdd.n1075 185
R1390 vdd.n2311 vdd.n1082 185
R1391 vdd.n2384 vdd.n1082 185
R1392 vdd.n370 vdd.n369 185
R1393 vdd.n3436 vdd.n370 185
R1394 vdd.n3439 vdd.n3438 185
R1395 vdd.n3438 vdd.n3437 185
R1396 vdd.n3440 vdd.n364 185
R1397 vdd.n364 vdd.n363 185
R1398 vdd.n3442 vdd.n3441 185
R1399 vdd.n3443 vdd.n3442 185
R1400 vdd.n359 vdd.n358 185
R1401 vdd.n3444 vdd.n359 185
R1402 vdd.n3447 vdd.n3446 185
R1403 vdd.n3446 vdd.n3445 185
R1404 vdd.n3448 vdd.n353 185
R1405 vdd.n3418 vdd.n353 185
R1406 vdd.n3450 vdd.n3449 185
R1407 vdd.n3451 vdd.n3450 185
R1408 vdd.n348 vdd.n347 185
R1409 vdd.n3452 vdd.n348 185
R1410 vdd.n3455 vdd.n3454 185
R1411 vdd.n3454 vdd.n3453 185
R1412 vdd.n3456 vdd.n342 185
R1413 vdd.n349 vdd.n342 185
R1414 vdd.n3458 vdd.n3457 185
R1415 vdd.n3459 vdd.n3458 185
R1416 vdd.n338 vdd.n337 185
R1417 vdd.n3460 vdd.n338 185
R1418 vdd.n3463 vdd.n3462 185
R1419 vdd.n3462 vdd.n3461 185
R1420 vdd.n3464 vdd.n333 185
R1421 vdd.n333 vdd.n332 185
R1422 vdd.n3466 vdd.n3465 185
R1423 vdd.n3467 vdd.n3466 185
R1424 vdd.n327 vdd.n325 185
R1425 vdd.n3468 vdd.n327 185
R1426 vdd.n3471 vdd.n3470 185
R1427 vdd.n3470 vdd.n3469 185
R1428 vdd.n326 vdd.n324 185
R1429 vdd.n328 vdd.n326 185
R1430 vdd.n3394 vdd.n3393 185
R1431 vdd.n3395 vdd.n3394 185
R1432 vdd.n615 vdd.n614 185
R1433 vdd.n614 vdd.n613 185
R1434 vdd.n3389 vdd.n3388 185
R1435 vdd.n3388 vdd.n3387 185
R1436 vdd.n618 vdd.n617 185
R1437 vdd.n624 vdd.n618 185
R1438 vdd.n3375 vdd.n3374 185
R1439 vdd.n3376 vdd.n3375 185
R1440 vdd.n626 vdd.n625 185
R1441 vdd.n3367 vdd.n625 185
R1442 vdd.n3370 vdd.n3369 185
R1443 vdd.n3369 vdd.n3368 185
R1444 vdd.n629 vdd.n628 185
R1445 vdd.n636 vdd.n629 185
R1446 vdd.n3358 vdd.n3357 185
R1447 vdd.n3359 vdd.n3358 185
R1448 vdd.n638 vdd.n637 185
R1449 vdd.n637 vdd.n635 185
R1450 vdd.n3353 vdd.n3352 185
R1451 vdd.n3352 vdd.n3351 185
R1452 vdd.n641 vdd.n640 185
R1453 vdd.n642 vdd.n641 185
R1454 vdd.n3342 vdd.n3341 185
R1455 vdd.n3343 vdd.n3342 185
R1456 vdd.n650 vdd.n649 185
R1457 vdd.n649 vdd.n648 185
R1458 vdd.n3337 vdd.n3336 185
R1459 vdd.n3336 vdd.n3335 185
R1460 vdd.n653 vdd.n652 185
R1461 vdd.n659 vdd.n653 185
R1462 vdd.n3326 vdd.n3325 185
R1463 vdd.n3327 vdd.n3326 185
R1464 vdd.n3322 vdd.n660 185
R1465 vdd.n3321 vdd.n3320 185
R1466 vdd.n3318 vdd.n662 185
R1467 vdd.n3318 vdd.n658 185
R1468 vdd.n3317 vdd.n3316 185
R1469 vdd.n3315 vdd.n3314 185
R1470 vdd.n3313 vdd.n3312 185
R1471 vdd.n3311 vdd.n3310 185
R1472 vdd.n3309 vdd.n668 185
R1473 vdd.n3307 vdd.n3306 185
R1474 vdd.n3305 vdd.n669 185
R1475 vdd.n3304 vdd.n3303 185
R1476 vdd.n3301 vdd.n674 185
R1477 vdd.n3299 vdd.n3298 185
R1478 vdd.n3297 vdd.n675 185
R1479 vdd.n3296 vdd.n3295 185
R1480 vdd.n3293 vdd.n680 185
R1481 vdd.n3291 vdd.n3290 185
R1482 vdd.n3289 vdd.n681 185
R1483 vdd.n3288 vdd.n3287 185
R1484 vdd.n3285 vdd.n688 185
R1485 vdd.n3283 vdd.n3282 185
R1486 vdd.n3281 vdd.n689 185
R1487 vdd.n3280 vdd.n3279 185
R1488 vdd.n3277 vdd.n694 185
R1489 vdd.n3275 vdd.n3274 185
R1490 vdd.n3273 vdd.n695 185
R1491 vdd.n3272 vdd.n3271 185
R1492 vdd.n3269 vdd.n700 185
R1493 vdd.n3267 vdd.n3266 185
R1494 vdd.n3265 vdd.n701 185
R1495 vdd.n3264 vdd.n3263 185
R1496 vdd.n3261 vdd.n706 185
R1497 vdd.n3259 vdd.n3258 185
R1498 vdd.n3257 vdd.n707 185
R1499 vdd.n3256 vdd.n3255 185
R1500 vdd.n3253 vdd.n712 185
R1501 vdd.n3251 vdd.n3250 185
R1502 vdd.n3249 vdd.n713 185
R1503 vdd.n3248 vdd.n3247 185
R1504 vdd.n3245 vdd.n718 185
R1505 vdd.n3243 vdd.n3242 185
R1506 vdd.n3241 vdd.n719 185
R1507 vdd.n728 vdd.n722 185
R1508 vdd.n3237 vdd.n3236 185
R1509 vdd.n3234 vdd.n726 185
R1510 vdd.n3233 vdd.n3232 185
R1511 vdd.n3231 vdd.n3230 185
R1512 vdd.n3229 vdd.n732 185
R1513 vdd.n3227 vdd.n3226 185
R1514 vdd.n3225 vdd.n733 185
R1515 vdd.n3224 vdd.n3223 185
R1516 vdd.n3221 vdd.n738 185
R1517 vdd.n3219 vdd.n3218 185
R1518 vdd.n3217 vdd.n739 185
R1519 vdd.n3216 vdd.n3215 185
R1520 vdd.n3213 vdd.n744 185
R1521 vdd.n3211 vdd.n3210 185
R1522 vdd.n3209 vdd.n745 185
R1523 vdd.n3208 vdd.n3207 185
R1524 vdd.n3205 vdd.n3204 185
R1525 vdd.n3203 vdd.n3202 185
R1526 vdd.n3201 vdd.n3200 185
R1527 vdd.n3199 vdd.n3198 185
R1528 vdd.n3194 vdd.n657 185
R1529 vdd.n658 vdd.n657 185
R1530 vdd.n3433 vdd.n3432 185
R1531 vdd.n599 vdd.n404 185
R1532 vdd.n598 vdd.n597 185
R1533 vdd.n596 vdd.n595 185
R1534 vdd.n594 vdd.n409 185
R1535 vdd.n590 vdd.n589 185
R1536 vdd.n588 vdd.n587 185
R1537 vdd.n586 vdd.n585 185
R1538 vdd.n584 vdd.n411 185
R1539 vdd.n580 vdd.n579 185
R1540 vdd.n578 vdd.n577 185
R1541 vdd.n576 vdd.n575 185
R1542 vdd.n574 vdd.n413 185
R1543 vdd.n570 vdd.n569 185
R1544 vdd.n568 vdd.n567 185
R1545 vdd.n566 vdd.n565 185
R1546 vdd.n564 vdd.n415 185
R1547 vdd.n560 vdd.n559 185
R1548 vdd.n558 vdd.n557 185
R1549 vdd.n556 vdd.n555 185
R1550 vdd.n554 vdd.n417 185
R1551 vdd.n550 vdd.n549 185
R1552 vdd.n548 vdd.n547 185
R1553 vdd.n546 vdd.n545 185
R1554 vdd.n544 vdd.n421 185
R1555 vdd.n540 vdd.n539 185
R1556 vdd.n538 vdd.n537 185
R1557 vdd.n536 vdd.n535 185
R1558 vdd.n534 vdd.n423 185
R1559 vdd.n530 vdd.n529 185
R1560 vdd.n528 vdd.n527 185
R1561 vdd.n526 vdd.n525 185
R1562 vdd.n524 vdd.n425 185
R1563 vdd.n520 vdd.n519 185
R1564 vdd.n518 vdd.n517 185
R1565 vdd.n516 vdd.n515 185
R1566 vdd.n514 vdd.n427 185
R1567 vdd.n510 vdd.n509 185
R1568 vdd.n508 vdd.n507 185
R1569 vdd.n506 vdd.n505 185
R1570 vdd.n504 vdd.n429 185
R1571 vdd.n500 vdd.n499 185
R1572 vdd.n498 vdd.n497 185
R1573 vdd.n496 vdd.n495 185
R1574 vdd.n494 vdd.n433 185
R1575 vdd.n490 vdd.n489 185
R1576 vdd.n488 vdd.n487 185
R1577 vdd.n486 vdd.n485 185
R1578 vdd.n484 vdd.n435 185
R1579 vdd.n480 vdd.n479 185
R1580 vdd.n478 vdd.n477 185
R1581 vdd.n476 vdd.n475 185
R1582 vdd.n474 vdd.n437 185
R1583 vdd.n470 vdd.n469 185
R1584 vdd.n468 vdd.n467 185
R1585 vdd.n466 vdd.n465 185
R1586 vdd.n464 vdd.n439 185
R1587 vdd.n460 vdd.n459 185
R1588 vdd.n458 vdd.n457 185
R1589 vdd.n456 vdd.n455 185
R1590 vdd.n454 vdd.n441 185
R1591 vdd.n450 vdd.n449 185
R1592 vdd.n448 vdd.n447 185
R1593 vdd.n446 vdd.n445 185
R1594 vdd.n3429 vdd.n372 185
R1595 vdd.n3436 vdd.n372 185
R1596 vdd.n3428 vdd.n371 185
R1597 vdd.n3437 vdd.n371 185
R1598 vdd.n3427 vdd.n3426 185
R1599 vdd.n3426 vdd.n363 185
R1600 vdd.n602 vdd.n362 185
R1601 vdd.n3443 vdd.n362 185
R1602 vdd.n3422 vdd.n361 185
R1603 vdd.n3444 vdd.n361 185
R1604 vdd.n3421 vdd.n360 185
R1605 vdd.n3445 vdd.n360 185
R1606 vdd.n3420 vdd.n3419 185
R1607 vdd.n3419 vdd.n3418 185
R1608 vdd.n604 vdd.n352 185
R1609 vdd.n3451 vdd.n352 185
R1610 vdd.n3414 vdd.n351 185
R1611 vdd.n3452 vdd.n351 185
R1612 vdd.n3413 vdd.n350 185
R1613 vdd.n3453 vdd.n350 185
R1614 vdd.n3412 vdd.n3411 185
R1615 vdd.n3411 vdd.n349 185
R1616 vdd.n606 vdd.n341 185
R1617 vdd.n3459 vdd.n341 185
R1618 vdd.n3407 vdd.n340 185
R1619 vdd.n3460 vdd.n340 185
R1620 vdd.n3406 vdd.n339 185
R1621 vdd.n3461 vdd.n339 185
R1622 vdd.n3405 vdd.n3404 185
R1623 vdd.n3404 vdd.n332 185
R1624 vdd.n608 vdd.n331 185
R1625 vdd.n3467 vdd.n331 185
R1626 vdd.n3400 vdd.n330 185
R1627 vdd.n3468 vdd.n330 185
R1628 vdd.n3399 vdd.n329 185
R1629 vdd.n3469 vdd.n329 185
R1630 vdd.n3398 vdd.n3397 185
R1631 vdd.n3397 vdd.n328 185
R1632 vdd.n3396 vdd.n610 185
R1633 vdd.n3396 vdd.n3395 185
R1634 vdd.n3384 vdd.n612 185
R1635 vdd.n613 vdd.n612 185
R1636 vdd.n3386 vdd.n3385 185
R1637 vdd.n3387 vdd.n3386 185
R1638 vdd.n620 vdd.n619 185
R1639 vdd.n624 vdd.n619 185
R1640 vdd.n3378 vdd.n3377 185
R1641 vdd.n3377 vdd.n3376 185
R1642 vdd.n623 vdd.n622 185
R1643 vdd.n3367 vdd.n623 185
R1644 vdd.n3366 vdd.n3365 185
R1645 vdd.n3368 vdd.n3366 185
R1646 vdd.n631 vdd.n630 185
R1647 vdd.n636 vdd.n630 185
R1648 vdd.n3361 vdd.n3360 185
R1649 vdd.n3360 vdd.n3359 185
R1650 vdd.n634 vdd.n633 185
R1651 vdd.n635 vdd.n634 185
R1652 vdd.n3350 vdd.n3349 185
R1653 vdd.n3351 vdd.n3350 185
R1654 vdd.n644 vdd.n643 185
R1655 vdd.n643 vdd.n642 185
R1656 vdd.n3345 vdd.n3344 185
R1657 vdd.n3344 vdd.n3343 185
R1658 vdd.n647 vdd.n646 185
R1659 vdd.n648 vdd.n647 185
R1660 vdd.n3334 vdd.n3333 185
R1661 vdd.n3335 vdd.n3334 185
R1662 vdd.n655 vdd.n654 185
R1663 vdd.n659 vdd.n654 185
R1664 vdd.n3329 vdd.n3328 185
R1665 vdd.n3328 vdd.n3327 185
R1666 vdd.n2931 vdd.n918 185
R1667 vdd.n2930 vdd.n2929 185
R1668 vdd.n920 vdd.n919 185
R1669 vdd.n2927 vdd.n920 185
R1670 vdd.n2750 vdd.n2749 185
R1671 vdd.n2752 vdd.n2751 185
R1672 vdd.n2754 vdd.n2753 185
R1673 vdd.n2756 vdd.n2755 185
R1674 vdd.n2758 vdd.n2757 185
R1675 vdd.n2760 vdd.n2759 185
R1676 vdd.n2762 vdd.n2761 185
R1677 vdd.n2764 vdd.n2763 185
R1678 vdd.n2766 vdd.n2765 185
R1679 vdd.n2768 vdd.n2767 185
R1680 vdd.n2770 vdd.n2769 185
R1681 vdd.n2772 vdd.n2771 185
R1682 vdd.n2774 vdd.n2773 185
R1683 vdd.n2776 vdd.n2775 185
R1684 vdd.n2778 vdd.n2777 185
R1685 vdd.n2780 vdd.n2779 185
R1686 vdd.n2782 vdd.n2781 185
R1687 vdd.n2784 vdd.n2783 185
R1688 vdd.n2786 vdd.n2785 185
R1689 vdd.n2788 vdd.n2787 185
R1690 vdd.n2790 vdd.n2789 185
R1691 vdd.n2792 vdd.n2791 185
R1692 vdd.n2794 vdd.n2793 185
R1693 vdd.n2796 vdd.n2795 185
R1694 vdd.n2798 vdd.n2797 185
R1695 vdd.n2800 vdd.n2799 185
R1696 vdd.n2802 vdd.n2801 185
R1697 vdd.n2804 vdd.n2803 185
R1698 vdd.n2806 vdd.n2805 185
R1699 vdd.n2809 vdd.n2808 185
R1700 vdd.n2811 vdd.n2810 185
R1701 vdd.n2813 vdd.n2812 185
R1702 vdd.n3095 vdd.n3094 185
R1703 vdd.n3096 vdd.n803 185
R1704 vdd.n3098 vdd.n3097 185
R1705 vdd.n3100 vdd.n801 185
R1706 vdd.n3102 vdd.n3101 185
R1707 vdd.n3103 vdd.n800 185
R1708 vdd.n3105 vdd.n3104 185
R1709 vdd.n3107 vdd.n798 185
R1710 vdd.n3109 vdd.n3108 185
R1711 vdd.n3110 vdd.n797 185
R1712 vdd.n3112 vdd.n3111 185
R1713 vdd.n3114 vdd.n795 185
R1714 vdd.n3116 vdd.n3115 185
R1715 vdd.n3117 vdd.n794 185
R1716 vdd.n3119 vdd.n3118 185
R1717 vdd.n3121 vdd.n792 185
R1718 vdd.n3123 vdd.n3122 185
R1719 vdd.n3125 vdd.n791 185
R1720 vdd.n3127 vdd.n3126 185
R1721 vdd.n3129 vdd.n789 185
R1722 vdd.n3131 vdd.n3130 185
R1723 vdd.n3132 vdd.n788 185
R1724 vdd.n3134 vdd.n3133 185
R1725 vdd.n3136 vdd.n786 185
R1726 vdd.n3138 vdd.n3137 185
R1727 vdd.n3139 vdd.n785 185
R1728 vdd.n3141 vdd.n3140 185
R1729 vdd.n3143 vdd.n783 185
R1730 vdd.n3145 vdd.n3144 185
R1731 vdd.n3146 vdd.n782 185
R1732 vdd.n3148 vdd.n3147 185
R1733 vdd.n3150 vdd.n781 185
R1734 vdd.n3151 vdd.n780 185
R1735 vdd.n3154 vdd.n3153 185
R1736 vdd.n3155 vdd.n778 185
R1737 vdd.n778 vdd.n756 185
R1738 vdd.n3092 vdd.n775 185
R1739 vdd.n3158 vdd.n775 185
R1740 vdd.n3091 vdd.n3090 185
R1741 vdd.n3090 vdd.n774 185
R1742 vdd.n3089 vdd.n807 185
R1743 vdd.n3089 vdd.n3088 185
R1744 vdd.n2863 vdd.n808 185
R1745 vdd.n817 vdd.n808 185
R1746 vdd.n2864 vdd.n815 185
R1747 vdd.n3082 vdd.n815 185
R1748 vdd.n2866 vdd.n2865 185
R1749 vdd.n2865 vdd.n814 185
R1750 vdd.n2867 vdd.n823 185
R1751 vdd.n3031 vdd.n823 185
R1752 vdd.n2869 vdd.n2868 185
R1753 vdd.n2868 vdd.n822 185
R1754 vdd.n2870 vdd.n828 185
R1755 vdd.n3025 vdd.n828 185
R1756 vdd.n2872 vdd.n2871 185
R1757 vdd.n2871 vdd.n835 185
R1758 vdd.n2873 vdd.n833 185
R1759 vdd.n3019 vdd.n833 185
R1760 vdd.n2875 vdd.n2874 185
R1761 vdd.n2874 vdd.n841 185
R1762 vdd.n2876 vdd.n839 185
R1763 vdd.n3013 vdd.n839 185
R1764 vdd.n2878 vdd.n2877 185
R1765 vdd.n2877 vdd.n848 185
R1766 vdd.n2879 vdd.n846 185
R1767 vdd.n3007 vdd.n846 185
R1768 vdd.n2881 vdd.n2880 185
R1769 vdd.n2880 vdd.n845 185
R1770 vdd.n2882 vdd.n853 185
R1771 vdd.n3001 vdd.n853 185
R1772 vdd.n2884 vdd.n2883 185
R1773 vdd.n2883 vdd.n852 185
R1774 vdd.n2885 vdd.n860 185
R1775 vdd.n2994 vdd.n860 185
R1776 vdd.n2887 vdd.n2886 185
R1777 vdd.n2886 vdd.n859 185
R1778 vdd.n2888 vdd.n865 185
R1779 vdd.n2988 vdd.n865 185
R1780 vdd.n2890 vdd.n2889 185
R1781 vdd.n2889 vdd.n872 185
R1782 vdd.n2891 vdd.n870 185
R1783 vdd.n2982 vdd.n870 185
R1784 vdd.n2893 vdd.n2892 185
R1785 vdd.n2894 vdd.n2893 185
R1786 vdd.n2862 vdd.n877 185
R1787 vdd.n2976 vdd.n877 185
R1788 vdd.n2861 vdd.n2860 185
R1789 vdd.n2860 vdd.n876 185
R1790 vdd.n2859 vdd.n883 185
R1791 vdd.n2970 vdd.n883 185
R1792 vdd.n2858 vdd.n2857 185
R1793 vdd.n2857 vdd.n882 185
R1794 vdd.n2818 vdd.n888 185
R1795 vdd.n2964 vdd.n888 185
R1796 vdd.n2908 vdd.n2907 185
R1797 vdd.n2907 vdd.n2906 185
R1798 vdd.n2909 vdd.n893 185
R1799 vdd.n2958 vdd.n893 185
R1800 vdd.n2911 vdd.n2910 185
R1801 vdd.n2910 vdd.n901 185
R1802 vdd.n2912 vdd.n899 185
R1803 vdd.n2952 vdd.n899 185
R1804 vdd.n2914 vdd.n2913 185
R1805 vdd.n2913 vdd.n898 185
R1806 vdd.n2915 vdd.n905 185
R1807 vdd.n2946 vdd.n905 185
R1808 vdd.n2917 vdd.n2916 185
R1809 vdd.n2918 vdd.n2917 185
R1810 vdd.n2817 vdd.n910 185
R1811 vdd.n2940 vdd.n910 185
R1812 vdd.n2816 vdd.n2815 185
R1813 vdd.n2815 vdd.n917 185
R1814 vdd.n2814 vdd.n915 185
R1815 vdd.n2934 vdd.n915 185
R1816 vdd.n2933 vdd.n2932 185
R1817 vdd.n2934 vdd.n2933 185
R1818 vdd.n909 vdd.n908 185
R1819 vdd.n917 vdd.n909 185
R1820 vdd.n2942 vdd.n2941 185
R1821 vdd.n2941 vdd.n2940 185
R1822 vdd.n2943 vdd.n907 185
R1823 vdd.n2918 vdd.n907 185
R1824 vdd.n2945 vdd.n2944 185
R1825 vdd.n2946 vdd.n2945 185
R1826 vdd.n897 vdd.n896 185
R1827 vdd.n898 vdd.n897 185
R1828 vdd.n2954 vdd.n2953 185
R1829 vdd.n2953 vdd.n2952 185
R1830 vdd.n2955 vdd.n895 185
R1831 vdd.n901 vdd.n895 185
R1832 vdd.n2957 vdd.n2956 185
R1833 vdd.n2958 vdd.n2957 185
R1834 vdd.n887 vdd.n886 185
R1835 vdd.n2906 vdd.n887 185
R1836 vdd.n2966 vdd.n2965 185
R1837 vdd.n2965 vdd.n2964 185
R1838 vdd.n2967 vdd.n885 185
R1839 vdd.n885 vdd.n882 185
R1840 vdd.n2969 vdd.n2968 185
R1841 vdd.n2970 vdd.n2969 185
R1842 vdd.n875 vdd.n874 185
R1843 vdd.n876 vdd.n875 185
R1844 vdd.n2978 vdd.n2977 185
R1845 vdd.n2977 vdd.n2976 185
R1846 vdd.n2979 vdd.n873 185
R1847 vdd.n2894 vdd.n873 185
R1848 vdd.n2981 vdd.n2980 185
R1849 vdd.n2982 vdd.n2981 185
R1850 vdd.n864 vdd.n863 185
R1851 vdd.n872 vdd.n864 185
R1852 vdd.n2990 vdd.n2989 185
R1853 vdd.n2989 vdd.n2988 185
R1854 vdd.n2991 vdd.n862 185
R1855 vdd.n862 vdd.n859 185
R1856 vdd.n2993 vdd.n2992 185
R1857 vdd.n2994 vdd.n2993 185
R1858 vdd.n851 vdd.n850 185
R1859 vdd.n852 vdd.n851 185
R1860 vdd.n3003 vdd.n3002 185
R1861 vdd.n3002 vdd.n3001 185
R1862 vdd.n3004 vdd.n849 185
R1863 vdd.n849 vdd.n845 185
R1864 vdd.n3006 vdd.n3005 185
R1865 vdd.n3007 vdd.n3006 185
R1866 vdd.n838 vdd.n837 185
R1867 vdd.n848 vdd.n838 185
R1868 vdd.n3015 vdd.n3014 185
R1869 vdd.n3014 vdd.n3013 185
R1870 vdd.n3016 vdd.n836 185
R1871 vdd.n841 vdd.n836 185
R1872 vdd.n3018 vdd.n3017 185
R1873 vdd.n3019 vdd.n3018 185
R1874 vdd.n827 vdd.n826 185
R1875 vdd.n835 vdd.n827 185
R1876 vdd.n3027 vdd.n3026 185
R1877 vdd.n3026 vdd.n3025 185
R1878 vdd.n3028 vdd.n825 185
R1879 vdd.n825 vdd.n822 185
R1880 vdd.n3030 vdd.n3029 185
R1881 vdd.n3031 vdd.n3030 185
R1882 vdd.n813 vdd.n812 185
R1883 vdd.n814 vdd.n813 185
R1884 vdd.n3084 vdd.n3083 185
R1885 vdd.n3083 vdd.n3082 185
R1886 vdd.n3085 vdd.n811 185
R1887 vdd.n817 vdd.n811 185
R1888 vdd.n3087 vdd.n3086 185
R1889 vdd.n3088 vdd.n3087 185
R1890 vdd.n779 vdd.n777 185
R1891 vdd.n777 vdd.n774 185
R1892 vdd.n3157 vdd.n3156 185
R1893 vdd.n3158 vdd.n3157 185
R1894 vdd.n2570 vdd.n2569 185
R1895 vdd.n2571 vdd.n2570 185
R1896 vdd.n967 vdd.n965 185
R1897 vdd.n965 vdd.n963 185
R1898 vdd.n2485 vdd.n974 185
R1899 vdd.n2496 vdd.n974 185
R1900 vdd.n2486 vdd.n983 185
R1901 vdd.n2251 vdd.n983 185
R1902 vdd.n2488 vdd.n2487 185
R1903 vdd.n2489 vdd.n2488 185
R1904 vdd.n2484 vdd.n982 185
R1905 vdd.n982 vdd.n979 185
R1906 vdd.n2483 vdd.n2482 185
R1907 vdd.n2482 vdd.n2481 185
R1908 vdd.n985 vdd.n984 185
R1909 vdd.n986 vdd.n985 185
R1910 vdd.n2474 vdd.n2473 185
R1911 vdd.n2475 vdd.n2474 185
R1912 vdd.n2472 vdd.n994 185
R1913 vdd.n2263 vdd.n994 185
R1914 vdd.n2471 vdd.n2470 185
R1915 vdd.n2470 vdd.n2469 185
R1916 vdd.n996 vdd.n995 185
R1917 vdd.n1004 vdd.n996 185
R1918 vdd.n2462 vdd.n2461 185
R1919 vdd.n2463 vdd.n2462 185
R1920 vdd.n2460 vdd.n1005 185
R1921 vdd.n1010 vdd.n1005 185
R1922 vdd.n2459 vdd.n2458 185
R1923 vdd.n2458 vdd.n2457 185
R1924 vdd.n1007 vdd.n1006 185
R1925 vdd.n2275 vdd.n1007 185
R1926 vdd.n2450 vdd.n2449 185
R1927 vdd.n2451 vdd.n2450 185
R1928 vdd.n2448 vdd.n1017 185
R1929 vdd.n1017 vdd.n1014 185
R1930 vdd.n2447 vdd.n2446 185
R1931 vdd.n2446 vdd.n2445 185
R1932 vdd.n1019 vdd.n1018 185
R1933 vdd.n1020 vdd.n1019 185
R1934 vdd.n2438 vdd.n2437 185
R1935 vdd.n2439 vdd.n2438 185
R1936 vdd.n2435 vdd.n1028 185
R1937 vdd.n1034 vdd.n1028 185
R1938 vdd.n2434 vdd.n2433 185
R1939 vdd.n2433 vdd.n2432 185
R1940 vdd.n1031 vdd.n1030 185
R1941 vdd.n1041 vdd.n1031 185
R1942 vdd.n2425 vdd.n2424 185
R1943 vdd.n2426 vdd.n2425 185
R1944 vdd.n2423 vdd.n1042 185
R1945 vdd.n1042 vdd.n1038 185
R1946 vdd.n2422 vdd.n2421 185
R1947 vdd.n2421 vdd.n2420 185
R1948 vdd.n1044 vdd.n1043 185
R1949 vdd.n1045 vdd.n1044 185
R1950 vdd.n2413 vdd.n2412 185
R1951 vdd.n2414 vdd.n2413 185
R1952 vdd.n2411 vdd.n1054 185
R1953 vdd.n1054 vdd.n1051 185
R1954 vdd.n2410 vdd.n2409 185
R1955 vdd.n2409 vdd.n2408 185
R1956 vdd.n1056 vdd.n1055 185
R1957 vdd.n1057 vdd.n1056 185
R1958 vdd.n2401 vdd.n2400 185
R1959 vdd.n2402 vdd.n2401 185
R1960 vdd.n2399 vdd.n1066 185
R1961 vdd.n1066 vdd.n1063 185
R1962 vdd.n2398 vdd.n2397 185
R1963 vdd.n2397 vdd.n2396 185
R1964 vdd.n1068 vdd.n1067 185
R1965 vdd.n1069 vdd.n1068 185
R1966 vdd.n2389 vdd.n2388 185
R1967 vdd.n2390 vdd.n2389 185
R1968 vdd.n2387 vdd.n1078 185
R1969 vdd.n1078 vdd.n1075 185
R1970 vdd.n2386 vdd.n2385 185
R1971 vdd.n2385 vdd.n2384 185
R1972 vdd.n2501 vdd.n938 185
R1973 vdd.n2643 vdd.n938 185
R1974 vdd.n2503 vdd.n2502 185
R1975 vdd.n2505 vdd.n2504 185
R1976 vdd.n2507 vdd.n2506 185
R1977 vdd.n2509 vdd.n2508 185
R1978 vdd.n2511 vdd.n2510 185
R1979 vdd.n2513 vdd.n2512 185
R1980 vdd.n2515 vdd.n2514 185
R1981 vdd.n2517 vdd.n2516 185
R1982 vdd.n2519 vdd.n2518 185
R1983 vdd.n2521 vdd.n2520 185
R1984 vdd.n2523 vdd.n2522 185
R1985 vdd.n2525 vdd.n2524 185
R1986 vdd.n2527 vdd.n2526 185
R1987 vdd.n2529 vdd.n2528 185
R1988 vdd.n2531 vdd.n2530 185
R1989 vdd.n2533 vdd.n2532 185
R1990 vdd.n2535 vdd.n2534 185
R1991 vdd.n2537 vdd.n2536 185
R1992 vdd.n2539 vdd.n2538 185
R1993 vdd.n2541 vdd.n2540 185
R1994 vdd.n2543 vdd.n2542 185
R1995 vdd.n2545 vdd.n2544 185
R1996 vdd.n2547 vdd.n2546 185
R1997 vdd.n2549 vdd.n2548 185
R1998 vdd.n2551 vdd.n2550 185
R1999 vdd.n2553 vdd.n2552 185
R2000 vdd.n2555 vdd.n2554 185
R2001 vdd.n2557 vdd.n2556 185
R2002 vdd.n2559 vdd.n2558 185
R2003 vdd.n2561 vdd.n2560 185
R2004 vdd.n2563 vdd.n2562 185
R2005 vdd.n2565 vdd.n2564 185
R2006 vdd.n2567 vdd.n2566 185
R2007 vdd.n2568 vdd.n966 185
R2008 vdd.n2500 vdd.n964 185
R2009 vdd.n2571 vdd.n964 185
R2010 vdd.n2499 vdd.n2498 185
R2011 vdd.n2498 vdd.n963 185
R2012 vdd.n2497 vdd.n971 185
R2013 vdd.n2497 vdd.n2496 185
R2014 vdd.n2235 vdd.n972 185
R2015 vdd.n2251 vdd.n972 185
R2016 vdd.n2236 vdd.n981 185
R2017 vdd.n2489 vdd.n981 185
R2018 vdd.n2238 vdd.n2237 185
R2019 vdd.n2237 vdd.n979 185
R2020 vdd.n2239 vdd.n988 185
R2021 vdd.n2481 vdd.n988 185
R2022 vdd.n2241 vdd.n2240 185
R2023 vdd.n2240 vdd.n986 185
R2024 vdd.n2242 vdd.n993 185
R2025 vdd.n2475 vdd.n993 185
R2026 vdd.n2265 vdd.n2264 185
R2027 vdd.n2264 vdd.n2263 185
R2028 vdd.n2266 vdd.n998 185
R2029 vdd.n2469 vdd.n998 185
R2030 vdd.n2268 vdd.n2267 185
R2031 vdd.n2267 vdd.n1004 185
R2032 vdd.n2269 vdd.n1003 185
R2033 vdd.n2463 vdd.n1003 185
R2034 vdd.n2271 vdd.n2270 185
R2035 vdd.n2270 vdd.n1010 185
R2036 vdd.n2272 vdd.n1009 185
R2037 vdd.n2457 vdd.n1009 185
R2038 vdd.n2274 vdd.n2273 185
R2039 vdd.n2275 vdd.n2274 185
R2040 vdd.n2234 vdd.n1016 185
R2041 vdd.n2451 vdd.n1016 185
R2042 vdd.n2233 vdd.n2232 185
R2043 vdd.n2232 vdd.n1014 185
R2044 vdd.n2231 vdd.n1022 185
R2045 vdd.n2445 vdd.n1022 185
R2046 vdd.n2230 vdd.n2229 185
R2047 vdd.n2229 vdd.n1020 185
R2048 vdd.n2228 vdd.n1027 185
R2049 vdd.n2439 vdd.n1027 185
R2050 vdd.n2227 vdd.n2226 185
R2051 vdd.n2226 vdd.n1034 185
R2052 vdd.n2225 vdd.n1033 185
R2053 vdd.n2432 vdd.n1033 185
R2054 vdd.n2224 vdd.n2223 185
R2055 vdd.n2223 vdd.n1041 185
R2056 vdd.n2222 vdd.n1040 185
R2057 vdd.n2426 vdd.n1040 185
R2058 vdd.n2221 vdd.n2220 185
R2059 vdd.n2220 vdd.n1038 185
R2060 vdd.n2219 vdd.n1047 185
R2061 vdd.n2420 vdd.n1047 185
R2062 vdd.n2218 vdd.n2217 185
R2063 vdd.n2217 vdd.n1045 185
R2064 vdd.n2216 vdd.n1053 185
R2065 vdd.n2414 vdd.n1053 185
R2066 vdd.n2215 vdd.n2214 185
R2067 vdd.n2214 vdd.n1051 185
R2068 vdd.n2213 vdd.n1059 185
R2069 vdd.n2408 vdd.n1059 185
R2070 vdd.n2212 vdd.n2211 185
R2071 vdd.n2211 vdd.n1057 185
R2072 vdd.n2210 vdd.n1065 185
R2073 vdd.n2402 vdd.n1065 185
R2074 vdd.n2209 vdd.n2208 185
R2075 vdd.n2208 vdd.n1063 185
R2076 vdd.n2207 vdd.n1071 185
R2077 vdd.n2396 vdd.n1071 185
R2078 vdd.n2206 vdd.n2205 185
R2079 vdd.n2205 vdd.n1069 185
R2080 vdd.n2204 vdd.n1077 185
R2081 vdd.n2390 vdd.n1077 185
R2082 vdd.n2203 vdd.n2202 185
R2083 vdd.n2202 vdd.n1075 185
R2084 vdd.n2201 vdd.n1083 185
R2085 vdd.n2384 vdd.n1083 185
R2086 vdd.n1080 vdd.n1079 185
R2087 vdd.n2133 vdd.n2131 185
R2088 vdd.n2136 vdd.n2135 185
R2089 vdd.n2137 vdd.n2130 185
R2090 vdd.n2139 vdd.n2138 185
R2091 vdd.n2141 vdd.n2129 185
R2092 vdd.n2144 vdd.n2143 185
R2093 vdd.n2145 vdd.n2128 185
R2094 vdd.n2147 vdd.n2146 185
R2095 vdd.n2149 vdd.n2127 185
R2096 vdd.n2152 vdd.n2151 185
R2097 vdd.n2153 vdd.n2126 185
R2098 vdd.n2155 vdd.n2154 185
R2099 vdd.n2157 vdd.n2125 185
R2100 vdd.n2160 vdd.n2159 185
R2101 vdd.n2161 vdd.n2124 185
R2102 vdd.n2163 vdd.n2162 185
R2103 vdd.n2165 vdd.n2123 185
R2104 vdd.n2168 vdd.n2167 185
R2105 vdd.n2169 vdd.n1114 185
R2106 vdd.n2171 vdd.n2170 185
R2107 vdd.n2173 vdd.n1113 185
R2108 vdd.n2176 vdd.n2175 185
R2109 vdd.n2177 vdd.n1112 185
R2110 vdd.n2179 vdd.n2178 185
R2111 vdd.n2181 vdd.n1111 185
R2112 vdd.n2184 vdd.n2183 185
R2113 vdd.n2185 vdd.n1110 185
R2114 vdd.n2187 vdd.n2186 185
R2115 vdd.n2189 vdd.n1109 185
R2116 vdd.n2192 vdd.n2191 185
R2117 vdd.n2193 vdd.n1106 185
R2118 vdd.n2196 vdd.n2195 185
R2119 vdd.n2198 vdd.n1105 185
R2120 vdd.n2200 vdd.n2199 185
R2121 vdd.n2199 vdd.n1081 185
R2122 vdd.n315 vdd.n314 171.744
R2123 vdd.n314 vdd.n313 171.744
R2124 vdd.n313 vdd.n282 171.744
R2125 vdd.n306 vdd.n282 171.744
R2126 vdd.n306 vdd.n305 171.744
R2127 vdd.n305 vdd.n287 171.744
R2128 vdd.n298 vdd.n287 171.744
R2129 vdd.n298 vdd.n297 171.744
R2130 vdd.n297 vdd.n291 171.744
R2131 vdd.n260 vdd.n259 171.744
R2132 vdd.n259 vdd.n258 171.744
R2133 vdd.n258 vdd.n227 171.744
R2134 vdd.n251 vdd.n227 171.744
R2135 vdd.n251 vdd.n250 171.744
R2136 vdd.n250 vdd.n232 171.744
R2137 vdd.n243 vdd.n232 171.744
R2138 vdd.n243 vdd.n242 171.744
R2139 vdd.n242 vdd.n236 171.744
R2140 vdd.n217 vdd.n216 171.744
R2141 vdd.n216 vdd.n215 171.744
R2142 vdd.n215 vdd.n184 171.744
R2143 vdd.n208 vdd.n184 171.744
R2144 vdd.n208 vdd.n207 171.744
R2145 vdd.n207 vdd.n189 171.744
R2146 vdd.n200 vdd.n189 171.744
R2147 vdd.n200 vdd.n199 171.744
R2148 vdd.n199 vdd.n193 171.744
R2149 vdd.n162 vdd.n161 171.744
R2150 vdd.n161 vdd.n160 171.744
R2151 vdd.n160 vdd.n129 171.744
R2152 vdd.n153 vdd.n129 171.744
R2153 vdd.n153 vdd.n152 171.744
R2154 vdd.n152 vdd.n134 171.744
R2155 vdd.n145 vdd.n134 171.744
R2156 vdd.n145 vdd.n144 171.744
R2157 vdd.n144 vdd.n138 171.744
R2158 vdd.n120 vdd.n119 171.744
R2159 vdd.n119 vdd.n118 171.744
R2160 vdd.n118 vdd.n87 171.744
R2161 vdd.n111 vdd.n87 171.744
R2162 vdd.n111 vdd.n110 171.744
R2163 vdd.n110 vdd.n92 171.744
R2164 vdd.n103 vdd.n92 171.744
R2165 vdd.n103 vdd.n102 171.744
R2166 vdd.n102 vdd.n96 171.744
R2167 vdd.n65 vdd.n64 171.744
R2168 vdd.n64 vdd.n63 171.744
R2169 vdd.n63 vdd.n32 171.744
R2170 vdd.n56 vdd.n32 171.744
R2171 vdd.n56 vdd.n55 171.744
R2172 vdd.n55 vdd.n37 171.744
R2173 vdd.n48 vdd.n37 171.744
R2174 vdd.n48 vdd.n47 171.744
R2175 vdd.n47 vdd.n41 171.744
R2176 vdd.n1764 vdd.n1763 171.744
R2177 vdd.n1763 vdd.n1762 171.744
R2178 vdd.n1762 vdd.n1731 171.744
R2179 vdd.n1755 vdd.n1731 171.744
R2180 vdd.n1755 vdd.n1754 171.744
R2181 vdd.n1754 vdd.n1736 171.744
R2182 vdd.n1747 vdd.n1736 171.744
R2183 vdd.n1747 vdd.n1746 171.744
R2184 vdd.n1746 vdd.n1740 171.744
R2185 vdd.n1819 vdd.n1818 171.744
R2186 vdd.n1818 vdd.n1817 171.744
R2187 vdd.n1817 vdd.n1786 171.744
R2188 vdd.n1810 vdd.n1786 171.744
R2189 vdd.n1810 vdd.n1809 171.744
R2190 vdd.n1809 vdd.n1791 171.744
R2191 vdd.n1802 vdd.n1791 171.744
R2192 vdd.n1802 vdd.n1801 171.744
R2193 vdd.n1801 vdd.n1795 171.744
R2194 vdd.n1666 vdd.n1665 171.744
R2195 vdd.n1665 vdd.n1664 171.744
R2196 vdd.n1664 vdd.n1633 171.744
R2197 vdd.n1657 vdd.n1633 171.744
R2198 vdd.n1657 vdd.n1656 171.744
R2199 vdd.n1656 vdd.n1638 171.744
R2200 vdd.n1649 vdd.n1638 171.744
R2201 vdd.n1649 vdd.n1648 171.744
R2202 vdd.n1648 vdd.n1642 171.744
R2203 vdd.n1721 vdd.n1720 171.744
R2204 vdd.n1720 vdd.n1719 171.744
R2205 vdd.n1719 vdd.n1688 171.744
R2206 vdd.n1712 vdd.n1688 171.744
R2207 vdd.n1712 vdd.n1711 171.744
R2208 vdd.n1711 vdd.n1693 171.744
R2209 vdd.n1704 vdd.n1693 171.744
R2210 vdd.n1704 vdd.n1703 171.744
R2211 vdd.n1703 vdd.n1697 171.744
R2212 vdd.n1569 vdd.n1568 171.744
R2213 vdd.n1568 vdd.n1567 171.744
R2214 vdd.n1567 vdd.n1536 171.744
R2215 vdd.n1560 vdd.n1536 171.744
R2216 vdd.n1560 vdd.n1559 171.744
R2217 vdd.n1559 vdd.n1541 171.744
R2218 vdd.n1552 vdd.n1541 171.744
R2219 vdd.n1552 vdd.n1551 171.744
R2220 vdd.n1551 vdd.n1545 171.744
R2221 vdd.n1624 vdd.n1623 171.744
R2222 vdd.n1623 vdd.n1622 171.744
R2223 vdd.n1622 vdd.n1591 171.744
R2224 vdd.n1615 vdd.n1591 171.744
R2225 vdd.n1615 vdd.n1614 171.744
R2226 vdd.n1614 vdd.n1596 171.744
R2227 vdd.n1607 vdd.n1596 171.744
R2228 vdd.n1607 vdd.n1606 171.744
R2229 vdd.n1606 vdd.n1600 171.744
R2230 vdd.n449 vdd.n448 146.341
R2231 vdd.n455 vdd.n454 146.341
R2232 vdd.n459 vdd.n458 146.341
R2233 vdd.n465 vdd.n464 146.341
R2234 vdd.n469 vdd.n468 146.341
R2235 vdd.n475 vdd.n474 146.341
R2236 vdd.n479 vdd.n478 146.341
R2237 vdd.n485 vdd.n484 146.341
R2238 vdd.n489 vdd.n488 146.341
R2239 vdd.n495 vdd.n494 146.341
R2240 vdd.n499 vdd.n498 146.341
R2241 vdd.n505 vdd.n504 146.341
R2242 vdd.n509 vdd.n508 146.341
R2243 vdd.n515 vdd.n514 146.341
R2244 vdd.n519 vdd.n518 146.341
R2245 vdd.n525 vdd.n524 146.341
R2246 vdd.n529 vdd.n528 146.341
R2247 vdd.n535 vdd.n534 146.341
R2248 vdd.n539 vdd.n538 146.341
R2249 vdd.n545 vdd.n544 146.341
R2250 vdd.n549 vdd.n548 146.341
R2251 vdd.n555 vdd.n554 146.341
R2252 vdd.n559 vdd.n558 146.341
R2253 vdd.n565 vdd.n564 146.341
R2254 vdd.n569 vdd.n568 146.341
R2255 vdd.n575 vdd.n574 146.341
R2256 vdd.n579 vdd.n578 146.341
R2257 vdd.n585 vdd.n584 146.341
R2258 vdd.n589 vdd.n588 146.341
R2259 vdd.n595 vdd.n594 146.341
R2260 vdd.n597 vdd.n404 146.341
R2261 vdd.n3328 vdd.n654 146.341
R2262 vdd.n3334 vdd.n654 146.341
R2263 vdd.n3334 vdd.n647 146.341
R2264 vdd.n3344 vdd.n647 146.341
R2265 vdd.n3344 vdd.n643 146.341
R2266 vdd.n3350 vdd.n643 146.341
R2267 vdd.n3350 vdd.n634 146.341
R2268 vdd.n3360 vdd.n634 146.341
R2269 vdd.n3360 vdd.n630 146.341
R2270 vdd.n3366 vdd.n630 146.341
R2271 vdd.n3366 vdd.n623 146.341
R2272 vdd.n3377 vdd.n623 146.341
R2273 vdd.n3377 vdd.n619 146.341
R2274 vdd.n3386 vdd.n619 146.341
R2275 vdd.n3386 vdd.n612 146.341
R2276 vdd.n3396 vdd.n612 146.341
R2277 vdd.n3397 vdd.n3396 146.341
R2278 vdd.n3397 vdd.n329 146.341
R2279 vdd.n330 vdd.n329 146.341
R2280 vdd.n331 vdd.n330 146.341
R2281 vdd.n3404 vdd.n331 146.341
R2282 vdd.n3404 vdd.n339 146.341
R2283 vdd.n340 vdd.n339 146.341
R2284 vdd.n341 vdd.n340 146.341
R2285 vdd.n3411 vdd.n341 146.341
R2286 vdd.n3411 vdd.n350 146.341
R2287 vdd.n351 vdd.n350 146.341
R2288 vdd.n352 vdd.n351 146.341
R2289 vdd.n3419 vdd.n352 146.341
R2290 vdd.n3419 vdd.n360 146.341
R2291 vdd.n361 vdd.n360 146.341
R2292 vdd.n362 vdd.n361 146.341
R2293 vdd.n3426 vdd.n362 146.341
R2294 vdd.n3426 vdd.n371 146.341
R2295 vdd.n372 vdd.n371 146.341
R2296 vdd.n3320 vdd.n3318 146.341
R2297 vdd.n3318 vdd.n3317 146.341
R2298 vdd.n3314 vdd.n3313 146.341
R2299 vdd.n3310 vdd.n3309 146.341
R2300 vdd.n3307 vdd.n669 146.341
R2301 vdd.n3303 vdd.n3301 146.341
R2302 vdd.n3299 vdd.n675 146.341
R2303 vdd.n3295 vdd.n3293 146.341
R2304 vdd.n3291 vdd.n681 146.341
R2305 vdd.n3287 vdd.n3285 146.341
R2306 vdd.n3283 vdd.n689 146.341
R2307 vdd.n3279 vdd.n3277 146.341
R2308 vdd.n3275 vdd.n695 146.341
R2309 vdd.n3271 vdd.n3269 146.341
R2310 vdd.n3267 vdd.n701 146.341
R2311 vdd.n3263 vdd.n3261 146.341
R2312 vdd.n3259 vdd.n707 146.341
R2313 vdd.n3255 vdd.n3253 146.341
R2314 vdd.n3251 vdd.n713 146.341
R2315 vdd.n3247 vdd.n3245 146.341
R2316 vdd.n3243 vdd.n719 146.341
R2317 vdd.n3236 vdd.n728 146.341
R2318 vdd.n3234 vdd.n3233 146.341
R2319 vdd.n3230 vdd.n3229 146.341
R2320 vdd.n3227 vdd.n733 146.341
R2321 vdd.n3223 vdd.n3221 146.341
R2322 vdd.n3219 vdd.n739 146.341
R2323 vdd.n3215 vdd.n3213 146.341
R2324 vdd.n3211 vdd.n745 146.341
R2325 vdd.n3207 vdd.n3205 146.341
R2326 vdd.n3202 vdd.n3201 146.341
R2327 vdd.n3198 vdd.n657 146.341
R2328 vdd.n3326 vdd.n653 146.341
R2329 vdd.n3336 vdd.n653 146.341
R2330 vdd.n3336 vdd.n649 146.341
R2331 vdd.n3342 vdd.n649 146.341
R2332 vdd.n3342 vdd.n641 146.341
R2333 vdd.n3352 vdd.n641 146.341
R2334 vdd.n3352 vdd.n637 146.341
R2335 vdd.n3358 vdd.n637 146.341
R2336 vdd.n3358 vdd.n629 146.341
R2337 vdd.n3369 vdd.n629 146.341
R2338 vdd.n3369 vdd.n625 146.341
R2339 vdd.n3375 vdd.n625 146.341
R2340 vdd.n3375 vdd.n618 146.341
R2341 vdd.n3388 vdd.n618 146.341
R2342 vdd.n3388 vdd.n614 146.341
R2343 vdd.n3394 vdd.n614 146.341
R2344 vdd.n3394 vdd.n326 146.341
R2345 vdd.n3470 vdd.n326 146.341
R2346 vdd.n3470 vdd.n327 146.341
R2347 vdd.n3466 vdd.n327 146.341
R2348 vdd.n3466 vdd.n333 146.341
R2349 vdd.n3462 vdd.n333 146.341
R2350 vdd.n3462 vdd.n338 146.341
R2351 vdd.n3458 vdd.n338 146.341
R2352 vdd.n3458 vdd.n342 146.341
R2353 vdd.n3454 vdd.n342 146.341
R2354 vdd.n3454 vdd.n348 146.341
R2355 vdd.n3450 vdd.n348 146.341
R2356 vdd.n3450 vdd.n353 146.341
R2357 vdd.n3446 vdd.n353 146.341
R2358 vdd.n3446 vdd.n359 146.341
R2359 vdd.n3442 vdd.n359 146.341
R2360 vdd.n3442 vdd.n364 146.341
R2361 vdd.n3438 vdd.n364 146.341
R2362 vdd.n3438 vdd.n370 146.341
R2363 vdd.n2106 vdd.n2105 146.341
R2364 vdd.n2103 vdd.n1900 146.341
R2365 vdd.n2096 vdd.n1906 146.341
R2366 vdd.n2094 vdd.n2093 146.341
R2367 vdd.n2091 vdd.n1908 146.341
R2368 vdd.n2087 vdd.n2086 146.341
R2369 vdd.n2084 vdd.n1915 146.341
R2370 vdd.n2080 vdd.n2079 146.341
R2371 vdd.n2077 vdd.n1922 146.341
R2372 vdd.n1933 vdd.n1930 146.341
R2373 vdd.n2069 vdd.n2068 146.341
R2374 vdd.n2066 vdd.n1935 146.341
R2375 vdd.n2062 vdd.n2061 146.341
R2376 vdd.n2059 vdd.n1941 146.341
R2377 vdd.n2055 vdd.n2054 146.341
R2378 vdd.n2052 vdd.n1948 146.341
R2379 vdd.n2048 vdd.n2047 146.341
R2380 vdd.n2045 vdd.n1955 146.341
R2381 vdd.n2041 vdd.n2040 146.341
R2382 vdd.n2038 vdd.n1962 146.341
R2383 vdd.n1973 vdd.n1970 146.341
R2384 vdd.n2030 vdd.n2029 146.341
R2385 vdd.n2027 vdd.n1975 146.341
R2386 vdd.n2023 vdd.n2022 146.341
R2387 vdd.n2020 vdd.n1981 146.341
R2388 vdd.n2016 vdd.n2015 146.341
R2389 vdd.n2013 vdd.n1988 146.341
R2390 vdd.n2009 vdd.n2008 146.341
R2391 vdd.n2006 vdd.n2003 146.341
R2392 vdd.n2001 vdd.n1998 146.341
R2393 vdd.n1996 vdd.n1120 146.341
R2394 vdd.n1461 vdd.n1225 146.341
R2395 vdd.n1461 vdd.n1217 146.341
R2396 vdd.n1471 vdd.n1217 146.341
R2397 vdd.n1471 vdd.n1213 146.341
R2398 vdd.n1477 vdd.n1213 146.341
R2399 vdd.n1477 vdd.n1205 146.341
R2400 vdd.n1488 vdd.n1205 146.341
R2401 vdd.n1488 vdd.n1201 146.341
R2402 vdd.n1494 vdd.n1201 146.341
R2403 vdd.n1494 vdd.n1195 146.341
R2404 vdd.n1505 vdd.n1195 146.341
R2405 vdd.n1505 vdd.n1191 146.341
R2406 vdd.n1511 vdd.n1191 146.341
R2407 vdd.n1511 vdd.n1182 146.341
R2408 vdd.n1521 vdd.n1182 146.341
R2409 vdd.n1521 vdd.n1178 146.341
R2410 vdd.n1527 vdd.n1178 146.341
R2411 vdd.n1527 vdd.n1171 146.341
R2412 vdd.n1833 vdd.n1171 146.341
R2413 vdd.n1833 vdd.n1167 146.341
R2414 vdd.n1839 vdd.n1167 146.341
R2415 vdd.n1839 vdd.n1160 146.341
R2416 vdd.n1849 vdd.n1160 146.341
R2417 vdd.n1849 vdd.n1156 146.341
R2418 vdd.n1855 vdd.n1156 146.341
R2419 vdd.n1855 vdd.n1148 146.341
R2420 vdd.n1866 vdd.n1148 146.341
R2421 vdd.n1866 vdd.n1144 146.341
R2422 vdd.n1872 vdd.n1144 146.341
R2423 vdd.n1872 vdd.n1138 146.341
R2424 vdd.n1883 vdd.n1138 146.341
R2425 vdd.n1883 vdd.n1133 146.341
R2426 vdd.n1891 vdd.n1133 146.341
R2427 vdd.n1891 vdd.n1122 146.341
R2428 vdd.n2114 vdd.n1122 146.341
R2429 vdd.n1263 vdd.n1262 146.341
R2430 vdd.n1267 vdd.n1262 146.341
R2431 vdd.n1269 vdd.n1268 146.341
R2432 vdd.n1273 vdd.n1272 146.341
R2433 vdd.n1275 vdd.n1274 146.341
R2434 vdd.n1279 vdd.n1278 146.341
R2435 vdd.n1281 vdd.n1280 146.341
R2436 vdd.n1285 vdd.n1284 146.341
R2437 vdd.n1287 vdd.n1286 146.341
R2438 vdd.n1419 vdd.n1418 146.341
R2439 vdd.n1291 vdd.n1290 146.341
R2440 vdd.n1295 vdd.n1294 146.341
R2441 vdd.n1297 vdd.n1296 146.341
R2442 vdd.n1301 vdd.n1300 146.341
R2443 vdd.n1303 vdd.n1302 146.341
R2444 vdd.n1307 vdd.n1306 146.341
R2445 vdd.n1309 vdd.n1308 146.341
R2446 vdd.n1313 vdd.n1312 146.341
R2447 vdd.n1315 vdd.n1314 146.341
R2448 vdd.n1319 vdd.n1318 146.341
R2449 vdd.n1383 vdd.n1320 146.341
R2450 vdd.n1324 vdd.n1323 146.341
R2451 vdd.n1326 vdd.n1325 146.341
R2452 vdd.n1330 vdd.n1329 146.341
R2453 vdd.n1332 vdd.n1331 146.341
R2454 vdd.n1336 vdd.n1335 146.341
R2455 vdd.n1338 vdd.n1337 146.341
R2456 vdd.n1342 vdd.n1341 146.341
R2457 vdd.n1344 vdd.n1343 146.341
R2458 vdd.n1348 vdd.n1347 146.341
R2459 vdd.n1350 vdd.n1349 146.341
R2460 vdd.n1455 vdd.n1231 146.341
R2461 vdd.n1463 vdd.n1223 146.341
R2462 vdd.n1463 vdd.n1219 146.341
R2463 vdd.n1469 vdd.n1219 146.341
R2464 vdd.n1469 vdd.n1211 146.341
R2465 vdd.n1480 vdd.n1211 146.341
R2466 vdd.n1480 vdd.n1207 146.341
R2467 vdd.n1486 vdd.n1207 146.341
R2468 vdd.n1486 vdd.n1200 146.341
R2469 vdd.n1497 vdd.n1200 146.341
R2470 vdd.n1497 vdd.n1196 146.341
R2471 vdd.n1503 vdd.n1196 146.341
R2472 vdd.n1503 vdd.n1189 146.341
R2473 vdd.n1513 vdd.n1189 146.341
R2474 vdd.n1513 vdd.n1185 146.341
R2475 vdd.n1519 vdd.n1185 146.341
R2476 vdd.n1519 vdd.n1177 146.341
R2477 vdd.n1530 vdd.n1177 146.341
R2478 vdd.n1530 vdd.n1173 146.341
R2479 vdd.n1831 vdd.n1173 146.341
R2480 vdd.n1831 vdd.n1166 146.341
R2481 vdd.n1841 vdd.n1166 146.341
R2482 vdd.n1841 vdd.n1162 146.341
R2483 vdd.n1847 vdd.n1162 146.341
R2484 vdd.n1847 vdd.n1154 146.341
R2485 vdd.n1858 vdd.n1154 146.341
R2486 vdd.n1858 vdd.n1150 146.341
R2487 vdd.n1864 vdd.n1150 146.341
R2488 vdd.n1864 vdd.n1143 146.341
R2489 vdd.n1875 vdd.n1143 146.341
R2490 vdd.n1875 vdd.n1139 146.341
R2491 vdd.n1881 vdd.n1139 146.341
R2492 vdd.n1881 vdd.n1131 146.341
R2493 vdd.n1893 vdd.n1131 146.341
R2494 vdd.n1893 vdd.n1126 146.341
R2495 vdd.n2112 vdd.n1126 146.341
R2496 vdd.n1107 vdd.t46 127.284
R2497 vdd.n968 vdd.t83 127.284
R2498 vdd.n1101 vdd.t110 127.284
R2499 vdd.n959 vdd.t106 127.284
R2500 vdd.n856 vdd.t56 127.284
R2501 vdd.n856 vdd.t57 127.284
R2502 vdd.n2678 vdd.t101 127.284
R2503 vdd.n804 vdd.t76 127.284
R2504 vdd.n2747 vdd.t88 127.284
R2505 vdd.n768 vdd.t41 127.284
R2506 vdd.n1029 vdd.t97 127.284
R2507 vdd.n1029 vdd.t98 127.284
R2508 vdd.n22 vdd.n20 117.314
R2509 vdd.n17 vdd.n15 117.314
R2510 vdd.n27 vdd.n26 116.927
R2511 vdd.n24 vdd.n23 116.927
R2512 vdd.n22 vdd.n21 116.927
R2513 vdd.n17 vdd.n16 116.927
R2514 vdd.n19 vdd.n18 116.927
R2515 vdd.n27 vdd.n25 116.927
R2516 vdd.n1108 vdd.t45 111.188
R2517 vdd.n969 vdd.t84 111.188
R2518 vdd.n1102 vdd.t109 111.188
R2519 vdd.n960 vdd.t107 111.188
R2520 vdd.n2679 vdd.t100 111.188
R2521 vdd.n805 vdd.t77 111.188
R2522 vdd.n2748 vdd.t87 111.188
R2523 vdd.n769 vdd.t42 111.188
R2524 vdd.n2933 vdd.n909 99.5127
R2525 vdd.n2941 vdd.n909 99.5127
R2526 vdd.n2941 vdd.n907 99.5127
R2527 vdd.n2945 vdd.n907 99.5127
R2528 vdd.n2945 vdd.n897 99.5127
R2529 vdd.n2953 vdd.n897 99.5127
R2530 vdd.n2953 vdd.n895 99.5127
R2531 vdd.n2957 vdd.n895 99.5127
R2532 vdd.n2957 vdd.n887 99.5127
R2533 vdd.n2965 vdd.n887 99.5127
R2534 vdd.n2965 vdd.n885 99.5127
R2535 vdd.n2969 vdd.n885 99.5127
R2536 vdd.n2969 vdd.n875 99.5127
R2537 vdd.n2977 vdd.n875 99.5127
R2538 vdd.n2977 vdd.n873 99.5127
R2539 vdd.n2981 vdd.n873 99.5127
R2540 vdd.n2981 vdd.n864 99.5127
R2541 vdd.n2989 vdd.n864 99.5127
R2542 vdd.n2989 vdd.n862 99.5127
R2543 vdd.n2993 vdd.n862 99.5127
R2544 vdd.n2993 vdd.n851 99.5127
R2545 vdd.n3002 vdd.n851 99.5127
R2546 vdd.n3002 vdd.n849 99.5127
R2547 vdd.n3006 vdd.n849 99.5127
R2548 vdd.n3006 vdd.n838 99.5127
R2549 vdd.n3014 vdd.n838 99.5127
R2550 vdd.n3014 vdd.n836 99.5127
R2551 vdd.n3018 vdd.n836 99.5127
R2552 vdd.n3018 vdd.n827 99.5127
R2553 vdd.n3026 vdd.n827 99.5127
R2554 vdd.n3026 vdd.n825 99.5127
R2555 vdd.n3030 vdd.n825 99.5127
R2556 vdd.n3030 vdd.n813 99.5127
R2557 vdd.n3083 vdd.n813 99.5127
R2558 vdd.n3083 vdd.n811 99.5127
R2559 vdd.n3087 vdd.n811 99.5127
R2560 vdd.n3087 vdd.n777 99.5127
R2561 vdd.n3157 vdd.n777 99.5127
R2562 vdd.n3153 vdd.n778 99.5127
R2563 vdd.n3151 vdd.n3150 99.5127
R2564 vdd.n3148 vdd.n782 99.5127
R2565 vdd.n3144 vdd.n3143 99.5127
R2566 vdd.n3141 vdd.n785 99.5127
R2567 vdd.n3137 vdd.n3136 99.5127
R2568 vdd.n3134 vdd.n788 99.5127
R2569 vdd.n3130 vdd.n3129 99.5127
R2570 vdd.n3127 vdd.n791 99.5127
R2571 vdd.n3122 vdd.n3121 99.5127
R2572 vdd.n3119 vdd.n794 99.5127
R2573 vdd.n3115 vdd.n3114 99.5127
R2574 vdd.n3112 vdd.n797 99.5127
R2575 vdd.n3108 vdd.n3107 99.5127
R2576 vdd.n3105 vdd.n800 99.5127
R2577 vdd.n3101 vdd.n3100 99.5127
R2578 vdd.n3098 vdd.n803 99.5127
R2579 vdd.n2815 vdd.n915 99.5127
R2580 vdd.n2815 vdd.n910 99.5127
R2581 vdd.n2917 vdd.n910 99.5127
R2582 vdd.n2917 vdd.n905 99.5127
R2583 vdd.n2913 vdd.n905 99.5127
R2584 vdd.n2913 vdd.n899 99.5127
R2585 vdd.n2910 vdd.n899 99.5127
R2586 vdd.n2910 vdd.n893 99.5127
R2587 vdd.n2907 vdd.n893 99.5127
R2588 vdd.n2907 vdd.n888 99.5127
R2589 vdd.n2857 vdd.n888 99.5127
R2590 vdd.n2857 vdd.n883 99.5127
R2591 vdd.n2860 vdd.n883 99.5127
R2592 vdd.n2860 vdd.n877 99.5127
R2593 vdd.n2893 vdd.n877 99.5127
R2594 vdd.n2893 vdd.n870 99.5127
R2595 vdd.n2889 vdd.n870 99.5127
R2596 vdd.n2889 vdd.n865 99.5127
R2597 vdd.n2886 vdd.n865 99.5127
R2598 vdd.n2886 vdd.n860 99.5127
R2599 vdd.n2883 vdd.n860 99.5127
R2600 vdd.n2883 vdd.n853 99.5127
R2601 vdd.n2880 vdd.n853 99.5127
R2602 vdd.n2880 vdd.n846 99.5127
R2603 vdd.n2877 vdd.n846 99.5127
R2604 vdd.n2877 vdd.n839 99.5127
R2605 vdd.n2874 vdd.n839 99.5127
R2606 vdd.n2874 vdd.n833 99.5127
R2607 vdd.n2871 vdd.n833 99.5127
R2608 vdd.n2871 vdd.n828 99.5127
R2609 vdd.n2868 vdd.n828 99.5127
R2610 vdd.n2868 vdd.n823 99.5127
R2611 vdd.n2865 vdd.n823 99.5127
R2612 vdd.n2865 vdd.n815 99.5127
R2613 vdd.n815 vdd.n808 99.5127
R2614 vdd.n3089 vdd.n808 99.5127
R2615 vdd.n3090 vdd.n3089 99.5127
R2616 vdd.n3090 vdd.n775 99.5127
R2617 vdd.n2929 vdd.n920 99.5127
R2618 vdd.n2749 vdd.n920 99.5127
R2619 vdd.n2753 vdd.n2752 99.5127
R2620 vdd.n2757 vdd.n2756 99.5127
R2621 vdd.n2761 vdd.n2760 99.5127
R2622 vdd.n2765 vdd.n2764 99.5127
R2623 vdd.n2769 vdd.n2768 99.5127
R2624 vdd.n2773 vdd.n2772 99.5127
R2625 vdd.n2777 vdd.n2776 99.5127
R2626 vdd.n2781 vdd.n2780 99.5127
R2627 vdd.n2785 vdd.n2784 99.5127
R2628 vdd.n2789 vdd.n2788 99.5127
R2629 vdd.n2793 vdd.n2792 99.5127
R2630 vdd.n2797 vdd.n2796 99.5127
R2631 vdd.n2801 vdd.n2800 99.5127
R2632 vdd.n2805 vdd.n2804 99.5127
R2633 vdd.n2810 vdd.n2809 99.5127
R2634 vdd.n2642 vdd.n957 99.5127
R2635 vdd.n2638 vdd.n2637 99.5127
R2636 vdd.n2634 vdd.n2633 99.5127
R2637 vdd.n2630 vdd.n2629 99.5127
R2638 vdd.n2626 vdd.n2625 99.5127
R2639 vdd.n2622 vdd.n2621 99.5127
R2640 vdd.n2618 vdd.n2617 99.5127
R2641 vdd.n2614 vdd.n2613 99.5127
R2642 vdd.n2610 vdd.n2609 99.5127
R2643 vdd.n2606 vdd.n2605 99.5127
R2644 vdd.n2602 vdd.n2601 99.5127
R2645 vdd.n2598 vdd.n2597 99.5127
R2646 vdd.n2594 vdd.n2593 99.5127
R2647 vdd.n2590 vdd.n2589 99.5127
R2648 vdd.n2586 vdd.n2585 99.5127
R2649 vdd.n2582 vdd.n2581 99.5127
R2650 vdd.n2577 vdd.n2576 99.5127
R2651 vdd.n2309 vdd.n1082 99.5127
R2652 vdd.n2309 vdd.n1076 99.5127
R2653 vdd.n2306 vdd.n1076 99.5127
R2654 vdd.n2306 vdd.n1070 99.5127
R2655 vdd.n2303 vdd.n1070 99.5127
R2656 vdd.n2303 vdd.n1064 99.5127
R2657 vdd.n2300 vdd.n1064 99.5127
R2658 vdd.n2300 vdd.n1058 99.5127
R2659 vdd.n2297 vdd.n1058 99.5127
R2660 vdd.n2297 vdd.n1052 99.5127
R2661 vdd.n2294 vdd.n1052 99.5127
R2662 vdd.n2294 vdd.n1046 99.5127
R2663 vdd.n2291 vdd.n1046 99.5127
R2664 vdd.n2291 vdd.n1039 99.5127
R2665 vdd.n2288 vdd.n1039 99.5127
R2666 vdd.n2288 vdd.n1032 99.5127
R2667 vdd.n2285 vdd.n1032 99.5127
R2668 vdd.n2285 vdd.n1026 99.5127
R2669 vdd.n2282 vdd.n1026 99.5127
R2670 vdd.n2282 vdd.n1021 99.5127
R2671 vdd.n2279 vdd.n1021 99.5127
R2672 vdd.n2279 vdd.n1015 99.5127
R2673 vdd.n2276 vdd.n1015 99.5127
R2674 vdd.n2276 vdd.n1008 99.5127
R2675 vdd.n2243 vdd.n1008 99.5127
R2676 vdd.n2243 vdd.n1002 99.5127
R2677 vdd.n2246 vdd.n1002 99.5127
R2678 vdd.n2246 vdd.n997 99.5127
R2679 vdd.n2262 vdd.n997 99.5127
R2680 vdd.n2262 vdd.n992 99.5127
R2681 vdd.n2258 vdd.n992 99.5127
R2682 vdd.n2258 vdd.n987 99.5127
R2683 vdd.n2255 vdd.n987 99.5127
R2684 vdd.n2255 vdd.n980 99.5127
R2685 vdd.n2252 vdd.n980 99.5127
R2686 vdd.n2252 vdd.n973 99.5127
R2687 vdd.n973 vdd.n962 99.5127
R2688 vdd.n2572 vdd.n962 99.5127
R2689 vdd.n2379 vdd.n2377 99.5127
R2690 vdd.n2377 vdd.n2376 99.5127
R2691 vdd.n2373 vdd.n2372 99.5127
R2692 vdd.n2370 vdd.n1088 99.5127
R2693 vdd.n2366 vdd.n2364 99.5127
R2694 vdd.n2362 vdd.n1090 99.5127
R2695 vdd.n2358 vdd.n2356 99.5127
R2696 vdd.n2354 vdd.n1092 99.5127
R2697 vdd.n2350 vdd.n2348 99.5127
R2698 vdd.n2346 vdd.n1094 99.5127
R2699 vdd.n2342 vdd.n2340 99.5127
R2700 vdd.n2338 vdd.n1096 99.5127
R2701 vdd.n2334 vdd.n2332 99.5127
R2702 vdd.n2330 vdd.n1098 99.5127
R2703 vdd.n2326 vdd.n2324 99.5127
R2704 vdd.n2322 vdd.n1100 99.5127
R2705 vdd.n2317 vdd.n2315 99.5127
R2706 vdd.n2383 vdd.n1074 99.5127
R2707 vdd.n2391 vdd.n1074 99.5127
R2708 vdd.n2391 vdd.n1072 99.5127
R2709 vdd.n2395 vdd.n1072 99.5127
R2710 vdd.n2395 vdd.n1062 99.5127
R2711 vdd.n2403 vdd.n1062 99.5127
R2712 vdd.n2403 vdd.n1060 99.5127
R2713 vdd.n2407 vdd.n1060 99.5127
R2714 vdd.n2407 vdd.n1050 99.5127
R2715 vdd.n2415 vdd.n1050 99.5127
R2716 vdd.n2415 vdd.n1048 99.5127
R2717 vdd.n2419 vdd.n1048 99.5127
R2718 vdd.n2419 vdd.n1037 99.5127
R2719 vdd.n2427 vdd.n1037 99.5127
R2720 vdd.n2427 vdd.n1035 99.5127
R2721 vdd.n2431 vdd.n1035 99.5127
R2722 vdd.n2431 vdd.n1025 99.5127
R2723 vdd.n2440 vdd.n1025 99.5127
R2724 vdd.n2440 vdd.n1023 99.5127
R2725 vdd.n2444 vdd.n1023 99.5127
R2726 vdd.n2444 vdd.n1013 99.5127
R2727 vdd.n2452 vdd.n1013 99.5127
R2728 vdd.n2452 vdd.n1011 99.5127
R2729 vdd.n2456 vdd.n1011 99.5127
R2730 vdd.n2456 vdd.n1001 99.5127
R2731 vdd.n2464 vdd.n1001 99.5127
R2732 vdd.n2464 vdd.n999 99.5127
R2733 vdd.n2468 vdd.n999 99.5127
R2734 vdd.n2468 vdd.n991 99.5127
R2735 vdd.n2476 vdd.n991 99.5127
R2736 vdd.n2476 vdd.n989 99.5127
R2737 vdd.n2480 vdd.n989 99.5127
R2738 vdd.n2480 vdd.n978 99.5127
R2739 vdd.n2490 vdd.n978 99.5127
R2740 vdd.n2490 vdd.n975 99.5127
R2741 vdd.n2495 vdd.n975 99.5127
R2742 vdd.n2495 vdd.n976 99.5127
R2743 vdd.n976 vdd.n956 99.5127
R2744 vdd.n3073 vdd.n3072 99.5127
R2745 vdd.n3070 vdd.n3036 99.5127
R2746 vdd.n3066 vdd.n3065 99.5127
R2747 vdd.n3063 vdd.n3039 99.5127
R2748 vdd.n3059 vdd.n3058 99.5127
R2749 vdd.n3056 vdd.n3042 99.5127
R2750 vdd.n3052 vdd.n3051 99.5127
R2751 vdd.n3049 vdd.n3046 99.5127
R2752 vdd.n3190 vdd.n755 99.5127
R2753 vdd.n3188 vdd.n3187 99.5127
R2754 vdd.n3185 vdd.n758 99.5127
R2755 vdd.n3181 vdd.n3180 99.5127
R2756 vdd.n3178 vdd.n761 99.5127
R2757 vdd.n3174 vdd.n3173 99.5127
R2758 vdd.n3171 vdd.n764 99.5127
R2759 vdd.n3167 vdd.n3166 99.5127
R2760 vdd.n3164 vdd.n767 99.5127
R2761 vdd.n2922 vdd.n916 99.5127
R2762 vdd.n2922 vdd.n911 99.5127
R2763 vdd.n2919 vdd.n911 99.5127
R2764 vdd.n2919 vdd.n906 99.5127
R2765 vdd.n2819 vdd.n906 99.5127
R2766 vdd.n2819 vdd.n900 99.5127
R2767 vdd.n2822 vdd.n900 99.5127
R2768 vdd.n2822 vdd.n894 99.5127
R2769 vdd.n2905 vdd.n894 99.5127
R2770 vdd.n2905 vdd.n889 99.5127
R2771 vdd.n2901 vdd.n889 99.5127
R2772 vdd.n2901 vdd.n884 99.5127
R2773 vdd.n2898 vdd.n884 99.5127
R2774 vdd.n2898 vdd.n878 99.5127
R2775 vdd.n2895 vdd.n878 99.5127
R2776 vdd.n2895 vdd.n871 99.5127
R2777 vdd.n2854 vdd.n871 99.5127
R2778 vdd.n2854 vdd.n866 99.5127
R2779 vdd.n2851 vdd.n866 99.5127
R2780 vdd.n2851 vdd.n861 99.5127
R2781 vdd.n2848 vdd.n861 99.5127
R2782 vdd.n2848 vdd.n854 99.5127
R2783 vdd.n2845 vdd.n854 99.5127
R2784 vdd.n2845 vdd.n847 99.5127
R2785 vdd.n2842 vdd.n847 99.5127
R2786 vdd.n2842 vdd.n840 99.5127
R2787 vdd.n2839 vdd.n840 99.5127
R2788 vdd.n2839 vdd.n834 99.5127
R2789 vdd.n2836 vdd.n834 99.5127
R2790 vdd.n2836 vdd.n829 99.5127
R2791 vdd.n2833 vdd.n829 99.5127
R2792 vdd.n2833 vdd.n824 99.5127
R2793 vdd.n2830 vdd.n824 99.5127
R2794 vdd.n2830 vdd.n816 99.5127
R2795 vdd.n2827 vdd.n816 99.5127
R2796 vdd.n2827 vdd.n809 99.5127
R2797 vdd.n809 vdd.n773 99.5127
R2798 vdd.n3159 vdd.n773 99.5127
R2799 vdd.n2683 vdd.n2682 99.5127
R2800 vdd.n2687 vdd.n2686 99.5127
R2801 vdd.n2691 vdd.n2690 99.5127
R2802 vdd.n2695 vdd.n2694 99.5127
R2803 vdd.n2699 vdd.n2698 99.5127
R2804 vdd.n2703 vdd.n2702 99.5127
R2805 vdd.n2707 vdd.n2706 99.5127
R2806 vdd.n2711 vdd.n2710 99.5127
R2807 vdd.n2715 vdd.n2714 99.5127
R2808 vdd.n2719 vdd.n2718 99.5127
R2809 vdd.n2723 vdd.n2722 99.5127
R2810 vdd.n2727 vdd.n2726 99.5127
R2811 vdd.n2731 vdd.n2730 99.5127
R2812 vdd.n2735 vdd.n2734 99.5127
R2813 vdd.n2739 vdd.n2738 99.5127
R2814 vdd.n2743 vdd.n2742 99.5127
R2815 vdd.n2926 vdd.n2677 99.5127
R2816 vdd.n2935 vdd.n912 99.5127
R2817 vdd.n2939 vdd.n912 99.5127
R2818 vdd.n2939 vdd.n904 99.5127
R2819 vdd.n2947 vdd.n904 99.5127
R2820 vdd.n2947 vdd.n902 99.5127
R2821 vdd.n2951 vdd.n902 99.5127
R2822 vdd.n2951 vdd.n892 99.5127
R2823 vdd.n2959 vdd.n892 99.5127
R2824 vdd.n2959 vdd.n890 99.5127
R2825 vdd.n2963 vdd.n890 99.5127
R2826 vdd.n2963 vdd.n881 99.5127
R2827 vdd.n2971 vdd.n881 99.5127
R2828 vdd.n2971 vdd.n879 99.5127
R2829 vdd.n2975 vdd.n879 99.5127
R2830 vdd.n2975 vdd.n869 99.5127
R2831 vdd.n2983 vdd.n869 99.5127
R2832 vdd.n2983 vdd.n867 99.5127
R2833 vdd.n2987 vdd.n867 99.5127
R2834 vdd.n2987 vdd.n858 99.5127
R2835 vdd.n2995 vdd.n858 99.5127
R2836 vdd.n2995 vdd.n855 99.5127
R2837 vdd.n3000 vdd.n855 99.5127
R2838 vdd.n3000 vdd.n844 99.5127
R2839 vdd.n3008 vdd.n844 99.5127
R2840 vdd.n3008 vdd.n842 99.5127
R2841 vdd.n3012 vdd.n842 99.5127
R2842 vdd.n3012 vdd.n832 99.5127
R2843 vdd.n3020 vdd.n832 99.5127
R2844 vdd.n3020 vdd.n830 99.5127
R2845 vdd.n3024 vdd.n830 99.5127
R2846 vdd.n3024 vdd.n821 99.5127
R2847 vdd.n3032 vdd.n821 99.5127
R2848 vdd.n3032 vdd.n818 99.5127
R2849 vdd.n3081 vdd.n818 99.5127
R2850 vdd.n3081 vdd.n819 99.5127
R2851 vdd.n819 vdd.n810 99.5127
R2852 vdd.n3076 vdd.n810 99.5127
R2853 vdd.n3076 vdd.n776 99.5127
R2854 vdd.n2566 vdd.n2565 99.5127
R2855 vdd.n2562 vdd.n2561 99.5127
R2856 vdd.n2558 vdd.n2557 99.5127
R2857 vdd.n2554 vdd.n2553 99.5127
R2858 vdd.n2550 vdd.n2549 99.5127
R2859 vdd.n2546 vdd.n2545 99.5127
R2860 vdd.n2542 vdd.n2541 99.5127
R2861 vdd.n2538 vdd.n2537 99.5127
R2862 vdd.n2534 vdd.n2533 99.5127
R2863 vdd.n2530 vdd.n2529 99.5127
R2864 vdd.n2526 vdd.n2525 99.5127
R2865 vdd.n2522 vdd.n2521 99.5127
R2866 vdd.n2518 vdd.n2517 99.5127
R2867 vdd.n2514 vdd.n2513 99.5127
R2868 vdd.n2510 vdd.n2509 99.5127
R2869 vdd.n2506 vdd.n2505 99.5127
R2870 vdd.n2502 vdd.n938 99.5127
R2871 vdd.n2202 vdd.n1083 99.5127
R2872 vdd.n2202 vdd.n1077 99.5127
R2873 vdd.n2205 vdd.n1077 99.5127
R2874 vdd.n2205 vdd.n1071 99.5127
R2875 vdd.n2208 vdd.n1071 99.5127
R2876 vdd.n2208 vdd.n1065 99.5127
R2877 vdd.n2211 vdd.n1065 99.5127
R2878 vdd.n2211 vdd.n1059 99.5127
R2879 vdd.n2214 vdd.n1059 99.5127
R2880 vdd.n2214 vdd.n1053 99.5127
R2881 vdd.n2217 vdd.n1053 99.5127
R2882 vdd.n2217 vdd.n1047 99.5127
R2883 vdd.n2220 vdd.n1047 99.5127
R2884 vdd.n2220 vdd.n1040 99.5127
R2885 vdd.n2223 vdd.n1040 99.5127
R2886 vdd.n2223 vdd.n1033 99.5127
R2887 vdd.n2226 vdd.n1033 99.5127
R2888 vdd.n2226 vdd.n1027 99.5127
R2889 vdd.n2229 vdd.n1027 99.5127
R2890 vdd.n2229 vdd.n1022 99.5127
R2891 vdd.n2232 vdd.n1022 99.5127
R2892 vdd.n2232 vdd.n1016 99.5127
R2893 vdd.n2274 vdd.n1016 99.5127
R2894 vdd.n2274 vdd.n1009 99.5127
R2895 vdd.n2270 vdd.n1009 99.5127
R2896 vdd.n2270 vdd.n1003 99.5127
R2897 vdd.n2267 vdd.n1003 99.5127
R2898 vdd.n2267 vdd.n998 99.5127
R2899 vdd.n2264 vdd.n998 99.5127
R2900 vdd.n2264 vdd.n993 99.5127
R2901 vdd.n2240 vdd.n993 99.5127
R2902 vdd.n2240 vdd.n988 99.5127
R2903 vdd.n2237 vdd.n988 99.5127
R2904 vdd.n2237 vdd.n981 99.5127
R2905 vdd.n981 vdd.n972 99.5127
R2906 vdd.n2497 vdd.n972 99.5127
R2907 vdd.n2498 vdd.n2497 99.5127
R2908 vdd.n2498 vdd.n964 99.5127
R2909 vdd.n2135 vdd.n2133 99.5127
R2910 vdd.n2139 vdd.n2130 99.5127
R2911 vdd.n2143 vdd.n2141 99.5127
R2912 vdd.n2147 vdd.n2128 99.5127
R2913 vdd.n2151 vdd.n2149 99.5127
R2914 vdd.n2155 vdd.n2126 99.5127
R2915 vdd.n2159 vdd.n2157 99.5127
R2916 vdd.n2163 vdd.n2124 99.5127
R2917 vdd.n2167 vdd.n2165 99.5127
R2918 vdd.n2171 vdd.n1114 99.5127
R2919 vdd.n2175 vdd.n2173 99.5127
R2920 vdd.n2179 vdd.n1112 99.5127
R2921 vdd.n2183 vdd.n2181 99.5127
R2922 vdd.n2187 vdd.n1110 99.5127
R2923 vdd.n2191 vdd.n2189 99.5127
R2924 vdd.n2196 vdd.n1106 99.5127
R2925 vdd.n2199 vdd.n2198 99.5127
R2926 vdd.n2385 vdd.n1078 99.5127
R2927 vdd.n2389 vdd.n1078 99.5127
R2928 vdd.n2389 vdd.n1068 99.5127
R2929 vdd.n2397 vdd.n1068 99.5127
R2930 vdd.n2397 vdd.n1066 99.5127
R2931 vdd.n2401 vdd.n1066 99.5127
R2932 vdd.n2401 vdd.n1056 99.5127
R2933 vdd.n2409 vdd.n1056 99.5127
R2934 vdd.n2409 vdd.n1054 99.5127
R2935 vdd.n2413 vdd.n1054 99.5127
R2936 vdd.n2413 vdd.n1044 99.5127
R2937 vdd.n2421 vdd.n1044 99.5127
R2938 vdd.n2421 vdd.n1042 99.5127
R2939 vdd.n2425 vdd.n1042 99.5127
R2940 vdd.n2425 vdd.n1031 99.5127
R2941 vdd.n2433 vdd.n1031 99.5127
R2942 vdd.n2433 vdd.n1028 99.5127
R2943 vdd.n2438 vdd.n1028 99.5127
R2944 vdd.n2438 vdd.n1019 99.5127
R2945 vdd.n2446 vdd.n1019 99.5127
R2946 vdd.n2446 vdd.n1017 99.5127
R2947 vdd.n2450 vdd.n1017 99.5127
R2948 vdd.n2450 vdd.n1007 99.5127
R2949 vdd.n2458 vdd.n1007 99.5127
R2950 vdd.n2458 vdd.n1005 99.5127
R2951 vdd.n2462 vdd.n1005 99.5127
R2952 vdd.n2462 vdd.n996 99.5127
R2953 vdd.n2470 vdd.n996 99.5127
R2954 vdd.n2470 vdd.n994 99.5127
R2955 vdd.n2474 vdd.n994 99.5127
R2956 vdd.n2474 vdd.n985 99.5127
R2957 vdd.n2482 vdd.n985 99.5127
R2958 vdd.n2482 vdd.n982 99.5127
R2959 vdd.n2488 vdd.n982 99.5127
R2960 vdd.n2488 vdd.n983 99.5127
R2961 vdd.n983 vdd.n974 99.5127
R2962 vdd.n974 vdd.n965 99.5127
R2963 vdd.n2570 vdd.n965 99.5127
R2964 vdd.n9 vdd.n7 98.9633
R2965 vdd.n2 vdd.n0 98.9633
R2966 vdd.n9 vdd.n8 98.6055
R2967 vdd.n11 vdd.n10 98.6055
R2968 vdd.n13 vdd.n12 98.6055
R2969 vdd.n6 vdd.n5 98.6055
R2970 vdd.n4 vdd.n3 98.6055
R2971 vdd.n2 vdd.n1 98.6055
R2972 vdd.t148 vdd.n291 85.8723
R2973 vdd.t199 vdd.n236 85.8723
R2974 vdd.t255 vdd.n193 85.8723
R2975 vdd.t183 vdd.n138 85.8723
R2976 vdd.t178 vdd.n96 85.8723
R2977 vdd.t239 vdd.n41 85.8723
R2978 vdd.t257 vdd.n1740 85.8723
R2979 vdd.t197 vdd.n1795 85.8723
R2980 vdd.t249 vdd.n1642 85.8723
R2981 vdd.t179 vdd.n1697 85.8723
R2982 vdd.t215 vdd.n1545 85.8723
R2983 vdd.t177 vdd.n1600 85.8723
R2984 vdd.n2997 vdd.n856 78.546
R2985 vdd.n2436 vdd.n1029 78.546
R2986 vdd.n278 vdd.n277 75.1835
R2987 vdd.n276 vdd.n275 75.1835
R2988 vdd.n274 vdd.n273 75.1835
R2989 vdd.n272 vdd.n271 75.1835
R2990 vdd.n270 vdd.n269 75.1835
R2991 vdd.n268 vdd.n267 75.1835
R2992 vdd.n266 vdd.n265 75.1835
R2993 vdd.n180 vdd.n179 75.1835
R2994 vdd.n178 vdd.n177 75.1835
R2995 vdd.n176 vdd.n175 75.1835
R2996 vdd.n174 vdd.n173 75.1835
R2997 vdd.n172 vdd.n171 75.1835
R2998 vdd.n170 vdd.n169 75.1835
R2999 vdd.n168 vdd.n167 75.1835
R3000 vdd.n83 vdd.n82 75.1835
R3001 vdd.n81 vdd.n80 75.1835
R3002 vdd.n79 vdd.n78 75.1835
R3003 vdd.n77 vdd.n76 75.1835
R3004 vdd.n75 vdd.n74 75.1835
R3005 vdd.n73 vdd.n72 75.1835
R3006 vdd.n71 vdd.n70 75.1835
R3007 vdd.n1770 vdd.n1769 75.1835
R3008 vdd.n1772 vdd.n1771 75.1835
R3009 vdd.n1774 vdd.n1773 75.1835
R3010 vdd.n1776 vdd.n1775 75.1835
R3011 vdd.n1778 vdd.n1777 75.1835
R3012 vdd.n1780 vdd.n1779 75.1835
R3013 vdd.n1782 vdd.n1781 75.1835
R3014 vdd.n1672 vdd.n1671 75.1835
R3015 vdd.n1674 vdd.n1673 75.1835
R3016 vdd.n1676 vdd.n1675 75.1835
R3017 vdd.n1678 vdd.n1677 75.1835
R3018 vdd.n1680 vdd.n1679 75.1835
R3019 vdd.n1682 vdd.n1681 75.1835
R3020 vdd.n1684 vdd.n1683 75.1835
R3021 vdd.n1575 vdd.n1574 75.1835
R3022 vdd.n1577 vdd.n1576 75.1835
R3023 vdd.n1579 vdd.n1578 75.1835
R3024 vdd.n1581 vdd.n1580 75.1835
R3025 vdd.n1583 vdd.n1582 75.1835
R3026 vdd.n1585 vdd.n1584 75.1835
R3027 vdd.n1587 vdd.n1586 75.1835
R3028 vdd.n2927 vdd.n2660 72.8958
R3029 vdd.n2927 vdd.n2661 72.8958
R3030 vdd.n2927 vdd.n2662 72.8958
R3031 vdd.n2927 vdd.n2663 72.8958
R3032 vdd.n2927 vdd.n2664 72.8958
R3033 vdd.n2927 vdd.n2665 72.8958
R3034 vdd.n2927 vdd.n2666 72.8958
R3035 vdd.n2927 vdd.n2667 72.8958
R3036 vdd.n2927 vdd.n2668 72.8958
R3037 vdd.n2927 vdd.n2669 72.8958
R3038 vdd.n2927 vdd.n2670 72.8958
R3039 vdd.n2927 vdd.n2671 72.8958
R3040 vdd.n2927 vdd.n2672 72.8958
R3041 vdd.n2927 vdd.n2673 72.8958
R3042 vdd.n2927 vdd.n2674 72.8958
R3043 vdd.n2927 vdd.n2675 72.8958
R3044 vdd.n2927 vdd.n2676 72.8958
R3045 vdd.n772 vdd.n756 72.8958
R3046 vdd.n3165 vdd.n756 72.8958
R3047 vdd.n766 vdd.n756 72.8958
R3048 vdd.n3172 vdd.n756 72.8958
R3049 vdd.n763 vdd.n756 72.8958
R3050 vdd.n3179 vdd.n756 72.8958
R3051 vdd.n760 vdd.n756 72.8958
R3052 vdd.n3186 vdd.n756 72.8958
R3053 vdd.n3189 vdd.n756 72.8958
R3054 vdd.n3045 vdd.n756 72.8958
R3055 vdd.n3050 vdd.n756 72.8958
R3056 vdd.n3044 vdd.n756 72.8958
R3057 vdd.n3057 vdd.n756 72.8958
R3058 vdd.n3041 vdd.n756 72.8958
R3059 vdd.n3064 vdd.n756 72.8958
R3060 vdd.n3038 vdd.n756 72.8958
R3061 vdd.n3071 vdd.n756 72.8958
R3062 vdd.n2378 vdd.n1081 72.8958
R3063 vdd.n1086 vdd.n1081 72.8958
R3064 vdd.n2371 vdd.n1081 72.8958
R3065 vdd.n2365 vdd.n1081 72.8958
R3066 vdd.n2363 vdd.n1081 72.8958
R3067 vdd.n2357 vdd.n1081 72.8958
R3068 vdd.n2355 vdd.n1081 72.8958
R3069 vdd.n2349 vdd.n1081 72.8958
R3070 vdd.n2347 vdd.n1081 72.8958
R3071 vdd.n2341 vdd.n1081 72.8958
R3072 vdd.n2339 vdd.n1081 72.8958
R3073 vdd.n2333 vdd.n1081 72.8958
R3074 vdd.n2331 vdd.n1081 72.8958
R3075 vdd.n2325 vdd.n1081 72.8958
R3076 vdd.n2323 vdd.n1081 72.8958
R3077 vdd.n2316 vdd.n1081 72.8958
R3078 vdd.n2314 vdd.n1081 72.8958
R3079 vdd.n2643 vdd.n939 72.8958
R3080 vdd.n2643 vdd.n940 72.8958
R3081 vdd.n2643 vdd.n941 72.8958
R3082 vdd.n2643 vdd.n942 72.8958
R3083 vdd.n2643 vdd.n943 72.8958
R3084 vdd.n2643 vdd.n944 72.8958
R3085 vdd.n2643 vdd.n945 72.8958
R3086 vdd.n2643 vdd.n946 72.8958
R3087 vdd.n2643 vdd.n947 72.8958
R3088 vdd.n2643 vdd.n948 72.8958
R3089 vdd.n2643 vdd.n949 72.8958
R3090 vdd.n2643 vdd.n950 72.8958
R3091 vdd.n2643 vdd.n951 72.8958
R3092 vdd.n2643 vdd.n952 72.8958
R3093 vdd.n2643 vdd.n953 72.8958
R3094 vdd.n2643 vdd.n954 72.8958
R3095 vdd.n2643 vdd.n955 72.8958
R3096 vdd.n2928 vdd.n2927 72.8958
R3097 vdd.n2927 vdd.n2644 72.8958
R3098 vdd.n2927 vdd.n2645 72.8958
R3099 vdd.n2927 vdd.n2646 72.8958
R3100 vdd.n2927 vdd.n2647 72.8958
R3101 vdd.n2927 vdd.n2648 72.8958
R3102 vdd.n2927 vdd.n2649 72.8958
R3103 vdd.n2927 vdd.n2650 72.8958
R3104 vdd.n2927 vdd.n2651 72.8958
R3105 vdd.n2927 vdd.n2652 72.8958
R3106 vdd.n2927 vdd.n2653 72.8958
R3107 vdd.n2927 vdd.n2654 72.8958
R3108 vdd.n2927 vdd.n2655 72.8958
R3109 vdd.n2927 vdd.n2656 72.8958
R3110 vdd.n2927 vdd.n2657 72.8958
R3111 vdd.n2927 vdd.n2658 72.8958
R3112 vdd.n2927 vdd.n2659 72.8958
R3113 vdd.n3093 vdd.n756 72.8958
R3114 vdd.n3099 vdd.n756 72.8958
R3115 vdd.n802 vdd.n756 72.8958
R3116 vdd.n3106 vdd.n756 72.8958
R3117 vdd.n799 vdd.n756 72.8958
R3118 vdd.n3113 vdd.n756 72.8958
R3119 vdd.n796 vdd.n756 72.8958
R3120 vdd.n3120 vdd.n756 72.8958
R3121 vdd.n793 vdd.n756 72.8958
R3122 vdd.n3128 vdd.n756 72.8958
R3123 vdd.n790 vdd.n756 72.8958
R3124 vdd.n3135 vdd.n756 72.8958
R3125 vdd.n787 vdd.n756 72.8958
R3126 vdd.n3142 vdd.n756 72.8958
R3127 vdd.n784 vdd.n756 72.8958
R3128 vdd.n3149 vdd.n756 72.8958
R3129 vdd.n3152 vdd.n756 72.8958
R3130 vdd.n2643 vdd.n937 72.8958
R3131 vdd.n2643 vdd.n936 72.8958
R3132 vdd.n2643 vdd.n935 72.8958
R3133 vdd.n2643 vdd.n934 72.8958
R3134 vdd.n2643 vdd.n933 72.8958
R3135 vdd.n2643 vdd.n932 72.8958
R3136 vdd.n2643 vdd.n931 72.8958
R3137 vdd.n2643 vdd.n930 72.8958
R3138 vdd.n2643 vdd.n929 72.8958
R3139 vdd.n2643 vdd.n928 72.8958
R3140 vdd.n2643 vdd.n927 72.8958
R3141 vdd.n2643 vdd.n926 72.8958
R3142 vdd.n2643 vdd.n925 72.8958
R3143 vdd.n2643 vdd.n924 72.8958
R3144 vdd.n2643 vdd.n923 72.8958
R3145 vdd.n2643 vdd.n922 72.8958
R3146 vdd.n2643 vdd.n921 72.8958
R3147 vdd.n2132 vdd.n1081 72.8958
R3148 vdd.n2134 vdd.n1081 72.8958
R3149 vdd.n2140 vdd.n1081 72.8958
R3150 vdd.n2142 vdd.n1081 72.8958
R3151 vdd.n2148 vdd.n1081 72.8958
R3152 vdd.n2150 vdd.n1081 72.8958
R3153 vdd.n2156 vdd.n1081 72.8958
R3154 vdd.n2158 vdd.n1081 72.8958
R3155 vdd.n2164 vdd.n1081 72.8958
R3156 vdd.n2166 vdd.n1081 72.8958
R3157 vdd.n2172 vdd.n1081 72.8958
R3158 vdd.n2174 vdd.n1081 72.8958
R3159 vdd.n2180 vdd.n1081 72.8958
R3160 vdd.n2182 vdd.n1081 72.8958
R3161 vdd.n2188 vdd.n1081 72.8958
R3162 vdd.n2190 vdd.n1081 72.8958
R3163 vdd.n2197 vdd.n1081 72.8958
R3164 vdd.n1454 vdd.n1453 66.2847
R3165 vdd.n1454 vdd.n1232 66.2847
R3166 vdd.n1454 vdd.n1233 66.2847
R3167 vdd.n1454 vdd.n1234 66.2847
R3168 vdd.n1454 vdd.n1235 66.2847
R3169 vdd.n1454 vdd.n1236 66.2847
R3170 vdd.n1454 vdd.n1237 66.2847
R3171 vdd.n1454 vdd.n1238 66.2847
R3172 vdd.n1454 vdd.n1239 66.2847
R3173 vdd.n1454 vdd.n1240 66.2847
R3174 vdd.n1454 vdd.n1241 66.2847
R3175 vdd.n1454 vdd.n1242 66.2847
R3176 vdd.n1454 vdd.n1243 66.2847
R3177 vdd.n1454 vdd.n1244 66.2847
R3178 vdd.n1454 vdd.n1245 66.2847
R3179 vdd.n1454 vdd.n1246 66.2847
R3180 vdd.n1454 vdd.n1247 66.2847
R3181 vdd.n1454 vdd.n1248 66.2847
R3182 vdd.n1454 vdd.n1249 66.2847
R3183 vdd.n1454 vdd.n1250 66.2847
R3184 vdd.n1454 vdd.n1251 66.2847
R3185 vdd.n1454 vdd.n1252 66.2847
R3186 vdd.n1454 vdd.n1253 66.2847
R3187 vdd.n1454 vdd.n1254 66.2847
R3188 vdd.n1454 vdd.n1255 66.2847
R3189 vdd.n1454 vdd.n1256 66.2847
R3190 vdd.n1454 vdd.n1257 66.2847
R3191 vdd.n1454 vdd.n1258 66.2847
R3192 vdd.n1454 vdd.n1259 66.2847
R3193 vdd.n1454 vdd.n1260 66.2847
R3194 vdd.n1454 vdd.n1261 66.2847
R3195 vdd.n1125 vdd.n1121 66.2847
R3196 vdd.n1997 vdd.n1125 66.2847
R3197 vdd.n2002 vdd.n1125 66.2847
R3198 vdd.n2007 vdd.n1125 66.2847
R3199 vdd.n1995 vdd.n1125 66.2847
R3200 vdd.n2014 vdd.n1125 66.2847
R3201 vdd.n1987 vdd.n1125 66.2847
R3202 vdd.n2021 vdd.n1125 66.2847
R3203 vdd.n1980 vdd.n1125 66.2847
R3204 vdd.n2028 vdd.n1125 66.2847
R3205 vdd.n1974 vdd.n1125 66.2847
R3206 vdd.n1969 vdd.n1125 66.2847
R3207 vdd.n2039 vdd.n1125 66.2847
R3208 vdd.n1961 vdd.n1125 66.2847
R3209 vdd.n2046 vdd.n1125 66.2847
R3210 vdd.n1954 vdd.n1125 66.2847
R3211 vdd.n2053 vdd.n1125 66.2847
R3212 vdd.n1947 vdd.n1125 66.2847
R3213 vdd.n2060 vdd.n1125 66.2847
R3214 vdd.n1940 vdd.n1125 66.2847
R3215 vdd.n2067 vdd.n1125 66.2847
R3216 vdd.n1934 vdd.n1125 66.2847
R3217 vdd.n1929 vdd.n1125 66.2847
R3218 vdd.n2078 vdd.n1125 66.2847
R3219 vdd.n1921 vdd.n1125 66.2847
R3220 vdd.n2085 vdd.n1125 66.2847
R3221 vdd.n1914 vdd.n1125 66.2847
R3222 vdd.n2092 vdd.n1125 66.2847
R3223 vdd.n2095 vdd.n1125 66.2847
R3224 vdd.n1905 vdd.n1125 66.2847
R3225 vdd.n2104 vdd.n1125 66.2847
R3226 vdd.n1899 vdd.n1125 66.2847
R3227 vdd.n3319 vdd.n658 66.2847
R3228 vdd.n663 vdd.n658 66.2847
R3229 vdd.n666 vdd.n658 66.2847
R3230 vdd.n3308 vdd.n658 66.2847
R3231 vdd.n3302 vdd.n658 66.2847
R3232 vdd.n3300 vdd.n658 66.2847
R3233 vdd.n3294 vdd.n658 66.2847
R3234 vdd.n3292 vdd.n658 66.2847
R3235 vdd.n3286 vdd.n658 66.2847
R3236 vdd.n3284 vdd.n658 66.2847
R3237 vdd.n3278 vdd.n658 66.2847
R3238 vdd.n3276 vdd.n658 66.2847
R3239 vdd.n3270 vdd.n658 66.2847
R3240 vdd.n3268 vdd.n658 66.2847
R3241 vdd.n3262 vdd.n658 66.2847
R3242 vdd.n3260 vdd.n658 66.2847
R3243 vdd.n3254 vdd.n658 66.2847
R3244 vdd.n3252 vdd.n658 66.2847
R3245 vdd.n3246 vdd.n658 66.2847
R3246 vdd.n3244 vdd.n658 66.2847
R3247 vdd.n727 vdd.n658 66.2847
R3248 vdd.n3235 vdd.n658 66.2847
R3249 vdd.n729 vdd.n658 66.2847
R3250 vdd.n3228 vdd.n658 66.2847
R3251 vdd.n3222 vdd.n658 66.2847
R3252 vdd.n3220 vdd.n658 66.2847
R3253 vdd.n3214 vdd.n658 66.2847
R3254 vdd.n3212 vdd.n658 66.2847
R3255 vdd.n3206 vdd.n658 66.2847
R3256 vdd.n750 vdd.n658 66.2847
R3257 vdd.n752 vdd.n658 66.2847
R3258 vdd.n3435 vdd.n3434 66.2847
R3259 vdd.n3435 vdd.n403 66.2847
R3260 vdd.n3435 vdd.n402 66.2847
R3261 vdd.n3435 vdd.n401 66.2847
R3262 vdd.n3435 vdd.n400 66.2847
R3263 vdd.n3435 vdd.n399 66.2847
R3264 vdd.n3435 vdd.n398 66.2847
R3265 vdd.n3435 vdd.n397 66.2847
R3266 vdd.n3435 vdd.n396 66.2847
R3267 vdd.n3435 vdd.n395 66.2847
R3268 vdd.n3435 vdd.n394 66.2847
R3269 vdd.n3435 vdd.n393 66.2847
R3270 vdd.n3435 vdd.n392 66.2847
R3271 vdd.n3435 vdd.n391 66.2847
R3272 vdd.n3435 vdd.n390 66.2847
R3273 vdd.n3435 vdd.n389 66.2847
R3274 vdd.n3435 vdd.n388 66.2847
R3275 vdd.n3435 vdd.n387 66.2847
R3276 vdd.n3435 vdd.n386 66.2847
R3277 vdd.n3435 vdd.n385 66.2847
R3278 vdd.n3435 vdd.n384 66.2847
R3279 vdd.n3435 vdd.n383 66.2847
R3280 vdd.n3435 vdd.n382 66.2847
R3281 vdd.n3435 vdd.n381 66.2847
R3282 vdd.n3435 vdd.n380 66.2847
R3283 vdd.n3435 vdd.n379 66.2847
R3284 vdd.n3435 vdd.n378 66.2847
R3285 vdd.n3435 vdd.n377 66.2847
R3286 vdd.n3435 vdd.n376 66.2847
R3287 vdd.n3435 vdd.n375 66.2847
R3288 vdd.n3435 vdd.n374 66.2847
R3289 vdd.n3435 vdd.n373 66.2847
R3290 vdd.n448 vdd.n373 52.4337
R3291 vdd.n454 vdd.n374 52.4337
R3292 vdd.n458 vdd.n375 52.4337
R3293 vdd.n464 vdd.n376 52.4337
R3294 vdd.n468 vdd.n377 52.4337
R3295 vdd.n474 vdd.n378 52.4337
R3296 vdd.n478 vdd.n379 52.4337
R3297 vdd.n484 vdd.n380 52.4337
R3298 vdd.n488 vdd.n381 52.4337
R3299 vdd.n494 vdd.n382 52.4337
R3300 vdd.n498 vdd.n383 52.4337
R3301 vdd.n504 vdd.n384 52.4337
R3302 vdd.n508 vdd.n385 52.4337
R3303 vdd.n514 vdd.n386 52.4337
R3304 vdd.n518 vdd.n387 52.4337
R3305 vdd.n524 vdd.n388 52.4337
R3306 vdd.n528 vdd.n389 52.4337
R3307 vdd.n534 vdd.n390 52.4337
R3308 vdd.n538 vdd.n391 52.4337
R3309 vdd.n544 vdd.n392 52.4337
R3310 vdd.n548 vdd.n393 52.4337
R3311 vdd.n554 vdd.n394 52.4337
R3312 vdd.n558 vdd.n395 52.4337
R3313 vdd.n564 vdd.n396 52.4337
R3314 vdd.n568 vdd.n397 52.4337
R3315 vdd.n574 vdd.n398 52.4337
R3316 vdd.n578 vdd.n399 52.4337
R3317 vdd.n584 vdd.n400 52.4337
R3318 vdd.n588 vdd.n401 52.4337
R3319 vdd.n594 vdd.n402 52.4337
R3320 vdd.n597 vdd.n403 52.4337
R3321 vdd.n3434 vdd.n3433 52.4337
R3322 vdd.n3319 vdd.n660 52.4337
R3323 vdd.n3317 vdd.n663 52.4337
R3324 vdd.n3313 vdd.n666 52.4337
R3325 vdd.n3309 vdd.n3308 52.4337
R3326 vdd.n3302 vdd.n669 52.4337
R3327 vdd.n3301 vdd.n3300 52.4337
R3328 vdd.n3294 vdd.n675 52.4337
R3329 vdd.n3293 vdd.n3292 52.4337
R3330 vdd.n3286 vdd.n681 52.4337
R3331 vdd.n3285 vdd.n3284 52.4337
R3332 vdd.n3278 vdd.n689 52.4337
R3333 vdd.n3277 vdd.n3276 52.4337
R3334 vdd.n3270 vdd.n695 52.4337
R3335 vdd.n3269 vdd.n3268 52.4337
R3336 vdd.n3262 vdd.n701 52.4337
R3337 vdd.n3261 vdd.n3260 52.4337
R3338 vdd.n3254 vdd.n707 52.4337
R3339 vdd.n3253 vdd.n3252 52.4337
R3340 vdd.n3246 vdd.n713 52.4337
R3341 vdd.n3245 vdd.n3244 52.4337
R3342 vdd.n727 vdd.n719 52.4337
R3343 vdd.n3236 vdd.n3235 52.4337
R3344 vdd.n3233 vdd.n729 52.4337
R3345 vdd.n3229 vdd.n3228 52.4337
R3346 vdd.n3222 vdd.n733 52.4337
R3347 vdd.n3221 vdd.n3220 52.4337
R3348 vdd.n3214 vdd.n739 52.4337
R3349 vdd.n3213 vdd.n3212 52.4337
R3350 vdd.n3206 vdd.n745 52.4337
R3351 vdd.n3205 vdd.n750 52.4337
R3352 vdd.n3201 vdd.n752 52.4337
R3353 vdd.n2106 vdd.n1899 52.4337
R3354 vdd.n2104 vdd.n2103 52.4337
R3355 vdd.n1906 vdd.n1905 52.4337
R3356 vdd.n2095 vdd.n2094 52.4337
R3357 vdd.n2092 vdd.n2091 52.4337
R3358 vdd.n2087 vdd.n1914 52.4337
R3359 vdd.n2085 vdd.n2084 52.4337
R3360 vdd.n2080 vdd.n1921 52.4337
R3361 vdd.n2078 vdd.n2077 52.4337
R3362 vdd.n1930 vdd.n1929 52.4337
R3363 vdd.n2069 vdd.n1934 52.4337
R3364 vdd.n2067 vdd.n2066 52.4337
R3365 vdd.n2062 vdd.n1940 52.4337
R3366 vdd.n2060 vdd.n2059 52.4337
R3367 vdd.n2055 vdd.n1947 52.4337
R3368 vdd.n2053 vdd.n2052 52.4337
R3369 vdd.n2048 vdd.n1954 52.4337
R3370 vdd.n2046 vdd.n2045 52.4337
R3371 vdd.n2041 vdd.n1961 52.4337
R3372 vdd.n2039 vdd.n2038 52.4337
R3373 vdd.n1970 vdd.n1969 52.4337
R3374 vdd.n2030 vdd.n1974 52.4337
R3375 vdd.n2028 vdd.n2027 52.4337
R3376 vdd.n2023 vdd.n1980 52.4337
R3377 vdd.n2021 vdd.n2020 52.4337
R3378 vdd.n2016 vdd.n1987 52.4337
R3379 vdd.n2014 vdd.n2013 52.4337
R3380 vdd.n2009 vdd.n1995 52.4337
R3381 vdd.n2007 vdd.n2006 52.4337
R3382 vdd.n2002 vdd.n2001 52.4337
R3383 vdd.n1997 vdd.n1996 52.4337
R3384 vdd.n2115 vdd.n1121 52.4337
R3385 vdd.n1453 vdd.n1452 52.4337
R3386 vdd.n1267 vdd.n1232 52.4337
R3387 vdd.n1269 vdd.n1233 52.4337
R3388 vdd.n1273 vdd.n1234 52.4337
R3389 vdd.n1275 vdd.n1235 52.4337
R3390 vdd.n1279 vdd.n1236 52.4337
R3391 vdd.n1281 vdd.n1237 52.4337
R3392 vdd.n1285 vdd.n1238 52.4337
R3393 vdd.n1287 vdd.n1239 52.4337
R3394 vdd.n1419 vdd.n1240 52.4337
R3395 vdd.n1291 vdd.n1241 52.4337
R3396 vdd.n1295 vdd.n1242 52.4337
R3397 vdd.n1297 vdd.n1243 52.4337
R3398 vdd.n1301 vdd.n1244 52.4337
R3399 vdd.n1303 vdd.n1245 52.4337
R3400 vdd.n1307 vdd.n1246 52.4337
R3401 vdd.n1309 vdd.n1247 52.4337
R3402 vdd.n1313 vdd.n1248 52.4337
R3403 vdd.n1315 vdd.n1249 52.4337
R3404 vdd.n1319 vdd.n1250 52.4337
R3405 vdd.n1383 vdd.n1251 52.4337
R3406 vdd.n1324 vdd.n1252 52.4337
R3407 vdd.n1326 vdd.n1253 52.4337
R3408 vdd.n1330 vdd.n1254 52.4337
R3409 vdd.n1332 vdd.n1255 52.4337
R3410 vdd.n1336 vdd.n1256 52.4337
R3411 vdd.n1338 vdd.n1257 52.4337
R3412 vdd.n1342 vdd.n1258 52.4337
R3413 vdd.n1344 vdd.n1259 52.4337
R3414 vdd.n1348 vdd.n1260 52.4337
R3415 vdd.n1350 vdd.n1261 52.4337
R3416 vdd.n1453 vdd.n1263 52.4337
R3417 vdd.n1268 vdd.n1232 52.4337
R3418 vdd.n1272 vdd.n1233 52.4337
R3419 vdd.n1274 vdd.n1234 52.4337
R3420 vdd.n1278 vdd.n1235 52.4337
R3421 vdd.n1280 vdd.n1236 52.4337
R3422 vdd.n1284 vdd.n1237 52.4337
R3423 vdd.n1286 vdd.n1238 52.4337
R3424 vdd.n1418 vdd.n1239 52.4337
R3425 vdd.n1290 vdd.n1240 52.4337
R3426 vdd.n1294 vdd.n1241 52.4337
R3427 vdd.n1296 vdd.n1242 52.4337
R3428 vdd.n1300 vdd.n1243 52.4337
R3429 vdd.n1302 vdd.n1244 52.4337
R3430 vdd.n1306 vdd.n1245 52.4337
R3431 vdd.n1308 vdd.n1246 52.4337
R3432 vdd.n1312 vdd.n1247 52.4337
R3433 vdd.n1314 vdd.n1248 52.4337
R3434 vdd.n1318 vdd.n1249 52.4337
R3435 vdd.n1320 vdd.n1250 52.4337
R3436 vdd.n1323 vdd.n1251 52.4337
R3437 vdd.n1325 vdd.n1252 52.4337
R3438 vdd.n1329 vdd.n1253 52.4337
R3439 vdd.n1331 vdd.n1254 52.4337
R3440 vdd.n1335 vdd.n1255 52.4337
R3441 vdd.n1337 vdd.n1256 52.4337
R3442 vdd.n1341 vdd.n1257 52.4337
R3443 vdd.n1343 vdd.n1258 52.4337
R3444 vdd.n1347 vdd.n1259 52.4337
R3445 vdd.n1349 vdd.n1260 52.4337
R3446 vdd.n1261 vdd.n1231 52.4337
R3447 vdd.n1121 vdd.n1120 52.4337
R3448 vdd.n1998 vdd.n1997 52.4337
R3449 vdd.n2003 vdd.n2002 52.4337
R3450 vdd.n2008 vdd.n2007 52.4337
R3451 vdd.n1995 vdd.n1988 52.4337
R3452 vdd.n2015 vdd.n2014 52.4337
R3453 vdd.n1987 vdd.n1981 52.4337
R3454 vdd.n2022 vdd.n2021 52.4337
R3455 vdd.n1980 vdd.n1975 52.4337
R3456 vdd.n2029 vdd.n2028 52.4337
R3457 vdd.n1974 vdd.n1973 52.4337
R3458 vdd.n1969 vdd.n1962 52.4337
R3459 vdd.n2040 vdd.n2039 52.4337
R3460 vdd.n1961 vdd.n1955 52.4337
R3461 vdd.n2047 vdd.n2046 52.4337
R3462 vdd.n1954 vdd.n1948 52.4337
R3463 vdd.n2054 vdd.n2053 52.4337
R3464 vdd.n1947 vdd.n1941 52.4337
R3465 vdd.n2061 vdd.n2060 52.4337
R3466 vdd.n1940 vdd.n1935 52.4337
R3467 vdd.n2068 vdd.n2067 52.4337
R3468 vdd.n1934 vdd.n1933 52.4337
R3469 vdd.n1929 vdd.n1922 52.4337
R3470 vdd.n2079 vdd.n2078 52.4337
R3471 vdd.n1921 vdd.n1915 52.4337
R3472 vdd.n2086 vdd.n2085 52.4337
R3473 vdd.n1914 vdd.n1908 52.4337
R3474 vdd.n2093 vdd.n2092 52.4337
R3475 vdd.n2096 vdd.n2095 52.4337
R3476 vdd.n1905 vdd.n1900 52.4337
R3477 vdd.n2105 vdd.n2104 52.4337
R3478 vdd.n1899 vdd.n1127 52.4337
R3479 vdd.n3320 vdd.n3319 52.4337
R3480 vdd.n3314 vdd.n663 52.4337
R3481 vdd.n3310 vdd.n666 52.4337
R3482 vdd.n3308 vdd.n3307 52.4337
R3483 vdd.n3303 vdd.n3302 52.4337
R3484 vdd.n3300 vdd.n3299 52.4337
R3485 vdd.n3295 vdd.n3294 52.4337
R3486 vdd.n3292 vdd.n3291 52.4337
R3487 vdd.n3287 vdd.n3286 52.4337
R3488 vdd.n3284 vdd.n3283 52.4337
R3489 vdd.n3279 vdd.n3278 52.4337
R3490 vdd.n3276 vdd.n3275 52.4337
R3491 vdd.n3271 vdd.n3270 52.4337
R3492 vdd.n3268 vdd.n3267 52.4337
R3493 vdd.n3263 vdd.n3262 52.4337
R3494 vdd.n3260 vdd.n3259 52.4337
R3495 vdd.n3255 vdd.n3254 52.4337
R3496 vdd.n3252 vdd.n3251 52.4337
R3497 vdd.n3247 vdd.n3246 52.4337
R3498 vdd.n3244 vdd.n3243 52.4337
R3499 vdd.n728 vdd.n727 52.4337
R3500 vdd.n3235 vdd.n3234 52.4337
R3501 vdd.n3230 vdd.n729 52.4337
R3502 vdd.n3228 vdd.n3227 52.4337
R3503 vdd.n3223 vdd.n3222 52.4337
R3504 vdd.n3220 vdd.n3219 52.4337
R3505 vdd.n3215 vdd.n3214 52.4337
R3506 vdd.n3212 vdd.n3211 52.4337
R3507 vdd.n3207 vdd.n3206 52.4337
R3508 vdd.n3202 vdd.n750 52.4337
R3509 vdd.n3198 vdd.n752 52.4337
R3510 vdd.n3434 vdd.n404 52.4337
R3511 vdd.n595 vdd.n403 52.4337
R3512 vdd.n589 vdd.n402 52.4337
R3513 vdd.n585 vdd.n401 52.4337
R3514 vdd.n579 vdd.n400 52.4337
R3515 vdd.n575 vdd.n399 52.4337
R3516 vdd.n569 vdd.n398 52.4337
R3517 vdd.n565 vdd.n397 52.4337
R3518 vdd.n559 vdd.n396 52.4337
R3519 vdd.n555 vdd.n395 52.4337
R3520 vdd.n549 vdd.n394 52.4337
R3521 vdd.n545 vdd.n393 52.4337
R3522 vdd.n539 vdd.n392 52.4337
R3523 vdd.n535 vdd.n391 52.4337
R3524 vdd.n529 vdd.n390 52.4337
R3525 vdd.n525 vdd.n389 52.4337
R3526 vdd.n519 vdd.n388 52.4337
R3527 vdd.n515 vdd.n387 52.4337
R3528 vdd.n509 vdd.n386 52.4337
R3529 vdd.n505 vdd.n385 52.4337
R3530 vdd.n499 vdd.n384 52.4337
R3531 vdd.n495 vdd.n383 52.4337
R3532 vdd.n489 vdd.n382 52.4337
R3533 vdd.n485 vdd.n381 52.4337
R3534 vdd.n479 vdd.n380 52.4337
R3535 vdd.n475 vdd.n379 52.4337
R3536 vdd.n469 vdd.n378 52.4337
R3537 vdd.n465 vdd.n377 52.4337
R3538 vdd.n459 vdd.n376 52.4337
R3539 vdd.n455 vdd.n375 52.4337
R3540 vdd.n449 vdd.n374 52.4337
R3541 vdd.n445 vdd.n373 52.4337
R3542 vdd.t119 vdd.t111 51.4683
R3543 vdd.n266 vdd.n264 42.0461
R3544 vdd.n168 vdd.n166 42.0461
R3545 vdd.n71 vdd.n69 42.0461
R3546 vdd.n1770 vdd.n1768 42.0461
R3547 vdd.n1672 vdd.n1670 42.0461
R3548 vdd.n1575 vdd.n1573 42.0461
R3549 vdd.n320 vdd.n319 41.6884
R3550 vdd.n222 vdd.n221 41.6884
R3551 vdd.n125 vdd.n124 41.6884
R3552 vdd.n1824 vdd.n1823 41.6884
R3553 vdd.n1726 vdd.n1725 41.6884
R3554 vdd.n1629 vdd.n1628 41.6884
R3555 vdd.n1230 vdd.n1229 41.1157
R3556 vdd.n1386 vdd.n1385 41.1157
R3557 vdd.n1422 vdd.n1421 41.1157
R3558 vdd.n407 vdd.n406 41.1157
R3559 vdd.n547 vdd.n420 41.1157
R3560 vdd.n433 vdd.n432 41.1157
R3561 vdd.n3152 vdd.n3151 39.2114
R3562 vdd.n3149 vdd.n3148 39.2114
R3563 vdd.n3144 vdd.n784 39.2114
R3564 vdd.n3142 vdd.n3141 39.2114
R3565 vdd.n3137 vdd.n787 39.2114
R3566 vdd.n3135 vdd.n3134 39.2114
R3567 vdd.n3130 vdd.n790 39.2114
R3568 vdd.n3128 vdd.n3127 39.2114
R3569 vdd.n3122 vdd.n793 39.2114
R3570 vdd.n3120 vdd.n3119 39.2114
R3571 vdd.n3115 vdd.n796 39.2114
R3572 vdd.n3113 vdd.n3112 39.2114
R3573 vdd.n3108 vdd.n799 39.2114
R3574 vdd.n3106 vdd.n3105 39.2114
R3575 vdd.n3101 vdd.n802 39.2114
R3576 vdd.n3099 vdd.n3098 39.2114
R3577 vdd.n3094 vdd.n3093 39.2114
R3578 vdd.n2928 vdd.n918 39.2114
R3579 vdd.n2749 vdd.n2644 39.2114
R3580 vdd.n2753 vdd.n2645 39.2114
R3581 vdd.n2757 vdd.n2646 39.2114
R3582 vdd.n2761 vdd.n2647 39.2114
R3583 vdd.n2765 vdd.n2648 39.2114
R3584 vdd.n2769 vdd.n2649 39.2114
R3585 vdd.n2773 vdd.n2650 39.2114
R3586 vdd.n2777 vdd.n2651 39.2114
R3587 vdd.n2781 vdd.n2652 39.2114
R3588 vdd.n2785 vdd.n2653 39.2114
R3589 vdd.n2789 vdd.n2654 39.2114
R3590 vdd.n2793 vdd.n2655 39.2114
R3591 vdd.n2797 vdd.n2656 39.2114
R3592 vdd.n2801 vdd.n2657 39.2114
R3593 vdd.n2805 vdd.n2658 39.2114
R3594 vdd.n2810 vdd.n2659 39.2114
R3595 vdd.n2638 vdd.n955 39.2114
R3596 vdd.n2634 vdd.n954 39.2114
R3597 vdd.n2630 vdd.n953 39.2114
R3598 vdd.n2626 vdd.n952 39.2114
R3599 vdd.n2622 vdd.n951 39.2114
R3600 vdd.n2618 vdd.n950 39.2114
R3601 vdd.n2614 vdd.n949 39.2114
R3602 vdd.n2610 vdd.n948 39.2114
R3603 vdd.n2606 vdd.n947 39.2114
R3604 vdd.n2602 vdd.n946 39.2114
R3605 vdd.n2598 vdd.n945 39.2114
R3606 vdd.n2594 vdd.n944 39.2114
R3607 vdd.n2590 vdd.n943 39.2114
R3608 vdd.n2586 vdd.n942 39.2114
R3609 vdd.n2582 vdd.n941 39.2114
R3610 vdd.n2577 vdd.n940 39.2114
R3611 vdd.n2573 vdd.n939 39.2114
R3612 vdd.n2378 vdd.n1084 39.2114
R3613 vdd.n2376 vdd.n1086 39.2114
R3614 vdd.n2372 vdd.n2371 39.2114
R3615 vdd.n2365 vdd.n1088 39.2114
R3616 vdd.n2364 vdd.n2363 39.2114
R3617 vdd.n2357 vdd.n1090 39.2114
R3618 vdd.n2356 vdd.n2355 39.2114
R3619 vdd.n2349 vdd.n1092 39.2114
R3620 vdd.n2348 vdd.n2347 39.2114
R3621 vdd.n2341 vdd.n1094 39.2114
R3622 vdd.n2340 vdd.n2339 39.2114
R3623 vdd.n2333 vdd.n1096 39.2114
R3624 vdd.n2332 vdd.n2331 39.2114
R3625 vdd.n2325 vdd.n1098 39.2114
R3626 vdd.n2324 vdd.n2323 39.2114
R3627 vdd.n2316 vdd.n1100 39.2114
R3628 vdd.n2315 vdd.n2314 39.2114
R3629 vdd.n3071 vdd.n3070 39.2114
R3630 vdd.n3066 vdd.n3038 39.2114
R3631 vdd.n3064 vdd.n3063 39.2114
R3632 vdd.n3059 vdd.n3041 39.2114
R3633 vdd.n3057 vdd.n3056 39.2114
R3634 vdd.n3052 vdd.n3044 39.2114
R3635 vdd.n3050 vdd.n3049 39.2114
R3636 vdd.n3045 vdd.n755 39.2114
R3637 vdd.n3189 vdd.n3188 39.2114
R3638 vdd.n3186 vdd.n3185 39.2114
R3639 vdd.n3181 vdd.n760 39.2114
R3640 vdd.n3179 vdd.n3178 39.2114
R3641 vdd.n3174 vdd.n763 39.2114
R3642 vdd.n3172 vdd.n3171 39.2114
R3643 vdd.n3167 vdd.n766 39.2114
R3644 vdd.n3165 vdd.n3164 39.2114
R3645 vdd.n3160 vdd.n772 39.2114
R3646 vdd.n2660 vdd.n914 39.2114
R3647 vdd.n2683 vdd.n2661 39.2114
R3648 vdd.n2687 vdd.n2662 39.2114
R3649 vdd.n2691 vdd.n2663 39.2114
R3650 vdd.n2695 vdd.n2664 39.2114
R3651 vdd.n2699 vdd.n2665 39.2114
R3652 vdd.n2703 vdd.n2666 39.2114
R3653 vdd.n2707 vdd.n2667 39.2114
R3654 vdd.n2711 vdd.n2668 39.2114
R3655 vdd.n2715 vdd.n2669 39.2114
R3656 vdd.n2719 vdd.n2670 39.2114
R3657 vdd.n2723 vdd.n2671 39.2114
R3658 vdd.n2727 vdd.n2672 39.2114
R3659 vdd.n2731 vdd.n2673 39.2114
R3660 vdd.n2735 vdd.n2674 39.2114
R3661 vdd.n2739 vdd.n2675 39.2114
R3662 vdd.n2743 vdd.n2676 39.2114
R3663 vdd.n2682 vdd.n2660 39.2114
R3664 vdd.n2686 vdd.n2661 39.2114
R3665 vdd.n2690 vdd.n2662 39.2114
R3666 vdd.n2694 vdd.n2663 39.2114
R3667 vdd.n2698 vdd.n2664 39.2114
R3668 vdd.n2702 vdd.n2665 39.2114
R3669 vdd.n2706 vdd.n2666 39.2114
R3670 vdd.n2710 vdd.n2667 39.2114
R3671 vdd.n2714 vdd.n2668 39.2114
R3672 vdd.n2718 vdd.n2669 39.2114
R3673 vdd.n2722 vdd.n2670 39.2114
R3674 vdd.n2726 vdd.n2671 39.2114
R3675 vdd.n2730 vdd.n2672 39.2114
R3676 vdd.n2734 vdd.n2673 39.2114
R3677 vdd.n2738 vdd.n2674 39.2114
R3678 vdd.n2742 vdd.n2675 39.2114
R3679 vdd.n2677 vdd.n2676 39.2114
R3680 vdd.n772 vdd.n767 39.2114
R3681 vdd.n3166 vdd.n3165 39.2114
R3682 vdd.n766 vdd.n764 39.2114
R3683 vdd.n3173 vdd.n3172 39.2114
R3684 vdd.n763 vdd.n761 39.2114
R3685 vdd.n3180 vdd.n3179 39.2114
R3686 vdd.n760 vdd.n758 39.2114
R3687 vdd.n3187 vdd.n3186 39.2114
R3688 vdd.n3190 vdd.n3189 39.2114
R3689 vdd.n3046 vdd.n3045 39.2114
R3690 vdd.n3051 vdd.n3050 39.2114
R3691 vdd.n3044 vdd.n3042 39.2114
R3692 vdd.n3058 vdd.n3057 39.2114
R3693 vdd.n3041 vdd.n3039 39.2114
R3694 vdd.n3065 vdd.n3064 39.2114
R3695 vdd.n3038 vdd.n3036 39.2114
R3696 vdd.n3072 vdd.n3071 39.2114
R3697 vdd.n2379 vdd.n2378 39.2114
R3698 vdd.n2373 vdd.n1086 39.2114
R3699 vdd.n2371 vdd.n2370 39.2114
R3700 vdd.n2366 vdd.n2365 39.2114
R3701 vdd.n2363 vdd.n2362 39.2114
R3702 vdd.n2358 vdd.n2357 39.2114
R3703 vdd.n2355 vdd.n2354 39.2114
R3704 vdd.n2350 vdd.n2349 39.2114
R3705 vdd.n2347 vdd.n2346 39.2114
R3706 vdd.n2342 vdd.n2341 39.2114
R3707 vdd.n2339 vdd.n2338 39.2114
R3708 vdd.n2334 vdd.n2333 39.2114
R3709 vdd.n2331 vdd.n2330 39.2114
R3710 vdd.n2326 vdd.n2325 39.2114
R3711 vdd.n2323 vdd.n2322 39.2114
R3712 vdd.n2317 vdd.n2316 39.2114
R3713 vdd.n2314 vdd.n2313 39.2114
R3714 vdd.n2576 vdd.n939 39.2114
R3715 vdd.n2581 vdd.n940 39.2114
R3716 vdd.n2585 vdd.n941 39.2114
R3717 vdd.n2589 vdd.n942 39.2114
R3718 vdd.n2593 vdd.n943 39.2114
R3719 vdd.n2597 vdd.n944 39.2114
R3720 vdd.n2601 vdd.n945 39.2114
R3721 vdd.n2605 vdd.n946 39.2114
R3722 vdd.n2609 vdd.n947 39.2114
R3723 vdd.n2613 vdd.n948 39.2114
R3724 vdd.n2617 vdd.n949 39.2114
R3725 vdd.n2621 vdd.n950 39.2114
R3726 vdd.n2625 vdd.n951 39.2114
R3727 vdd.n2629 vdd.n952 39.2114
R3728 vdd.n2633 vdd.n953 39.2114
R3729 vdd.n2637 vdd.n954 39.2114
R3730 vdd.n957 vdd.n955 39.2114
R3731 vdd.n2929 vdd.n2928 39.2114
R3732 vdd.n2752 vdd.n2644 39.2114
R3733 vdd.n2756 vdd.n2645 39.2114
R3734 vdd.n2760 vdd.n2646 39.2114
R3735 vdd.n2764 vdd.n2647 39.2114
R3736 vdd.n2768 vdd.n2648 39.2114
R3737 vdd.n2772 vdd.n2649 39.2114
R3738 vdd.n2776 vdd.n2650 39.2114
R3739 vdd.n2780 vdd.n2651 39.2114
R3740 vdd.n2784 vdd.n2652 39.2114
R3741 vdd.n2788 vdd.n2653 39.2114
R3742 vdd.n2792 vdd.n2654 39.2114
R3743 vdd.n2796 vdd.n2655 39.2114
R3744 vdd.n2800 vdd.n2656 39.2114
R3745 vdd.n2804 vdd.n2657 39.2114
R3746 vdd.n2809 vdd.n2658 39.2114
R3747 vdd.n2812 vdd.n2659 39.2114
R3748 vdd.n3093 vdd.n803 39.2114
R3749 vdd.n3100 vdd.n3099 39.2114
R3750 vdd.n802 vdd.n800 39.2114
R3751 vdd.n3107 vdd.n3106 39.2114
R3752 vdd.n799 vdd.n797 39.2114
R3753 vdd.n3114 vdd.n3113 39.2114
R3754 vdd.n796 vdd.n794 39.2114
R3755 vdd.n3121 vdd.n3120 39.2114
R3756 vdd.n793 vdd.n791 39.2114
R3757 vdd.n3129 vdd.n3128 39.2114
R3758 vdd.n790 vdd.n788 39.2114
R3759 vdd.n3136 vdd.n3135 39.2114
R3760 vdd.n787 vdd.n785 39.2114
R3761 vdd.n3143 vdd.n3142 39.2114
R3762 vdd.n784 vdd.n782 39.2114
R3763 vdd.n3150 vdd.n3149 39.2114
R3764 vdd.n3153 vdd.n3152 39.2114
R3765 vdd.n966 vdd.n921 39.2114
R3766 vdd.n2565 vdd.n922 39.2114
R3767 vdd.n2561 vdd.n923 39.2114
R3768 vdd.n2557 vdd.n924 39.2114
R3769 vdd.n2553 vdd.n925 39.2114
R3770 vdd.n2549 vdd.n926 39.2114
R3771 vdd.n2545 vdd.n927 39.2114
R3772 vdd.n2541 vdd.n928 39.2114
R3773 vdd.n2537 vdd.n929 39.2114
R3774 vdd.n2533 vdd.n930 39.2114
R3775 vdd.n2529 vdd.n931 39.2114
R3776 vdd.n2525 vdd.n932 39.2114
R3777 vdd.n2521 vdd.n933 39.2114
R3778 vdd.n2517 vdd.n934 39.2114
R3779 vdd.n2513 vdd.n935 39.2114
R3780 vdd.n2509 vdd.n936 39.2114
R3781 vdd.n2505 vdd.n937 39.2114
R3782 vdd.n2132 vdd.n1080 39.2114
R3783 vdd.n2135 vdd.n2134 39.2114
R3784 vdd.n2140 vdd.n2139 39.2114
R3785 vdd.n2143 vdd.n2142 39.2114
R3786 vdd.n2148 vdd.n2147 39.2114
R3787 vdd.n2151 vdd.n2150 39.2114
R3788 vdd.n2156 vdd.n2155 39.2114
R3789 vdd.n2159 vdd.n2158 39.2114
R3790 vdd.n2164 vdd.n2163 39.2114
R3791 vdd.n2167 vdd.n2166 39.2114
R3792 vdd.n2172 vdd.n2171 39.2114
R3793 vdd.n2175 vdd.n2174 39.2114
R3794 vdd.n2180 vdd.n2179 39.2114
R3795 vdd.n2183 vdd.n2182 39.2114
R3796 vdd.n2188 vdd.n2187 39.2114
R3797 vdd.n2191 vdd.n2190 39.2114
R3798 vdd.n2197 vdd.n2196 39.2114
R3799 vdd.n2502 vdd.n937 39.2114
R3800 vdd.n2506 vdd.n936 39.2114
R3801 vdd.n2510 vdd.n935 39.2114
R3802 vdd.n2514 vdd.n934 39.2114
R3803 vdd.n2518 vdd.n933 39.2114
R3804 vdd.n2522 vdd.n932 39.2114
R3805 vdd.n2526 vdd.n931 39.2114
R3806 vdd.n2530 vdd.n930 39.2114
R3807 vdd.n2534 vdd.n929 39.2114
R3808 vdd.n2538 vdd.n928 39.2114
R3809 vdd.n2542 vdd.n927 39.2114
R3810 vdd.n2546 vdd.n926 39.2114
R3811 vdd.n2550 vdd.n925 39.2114
R3812 vdd.n2554 vdd.n924 39.2114
R3813 vdd.n2558 vdd.n923 39.2114
R3814 vdd.n2562 vdd.n922 39.2114
R3815 vdd.n2566 vdd.n921 39.2114
R3816 vdd.n2133 vdd.n2132 39.2114
R3817 vdd.n2134 vdd.n2130 39.2114
R3818 vdd.n2141 vdd.n2140 39.2114
R3819 vdd.n2142 vdd.n2128 39.2114
R3820 vdd.n2149 vdd.n2148 39.2114
R3821 vdd.n2150 vdd.n2126 39.2114
R3822 vdd.n2157 vdd.n2156 39.2114
R3823 vdd.n2158 vdd.n2124 39.2114
R3824 vdd.n2165 vdd.n2164 39.2114
R3825 vdd.n2166 vdd.n1114 39.2114
R3826 vdd.n2173 vdd.n2172 39.2114
R3827 vdd.n2174 vdd.n1112 39.2114
R3828 vdd.n2181 vdd.n2180 39.2114
R3829 vdd.n2182 vdd.n1110 39.2114
R3830 vdd.n2189 vdd.n2188 39.2114
R3831 vdd.n2190 vdd.n1106 39.2114
R3832 vdd.n2198 vdd.n2197 39.2114
R3833 vdd.n2119 vdd.n2118 37.2369
R3834 vdd.n2035 vdd.n1968 37.2369
R3835 vdd.n2074 vdd.n1928 37.2369
R3836 vdd.n3241 vdd.n724 37.2369
R3837 vdd.n688 vdd.n687 37.2369
R3838 vdd.n3197 vdd.n3196 37.2369
R3839 vdd.n2194 vdd.n1108 30.449
R3840 vdd.n970 vdd.n969 30.449
R3841 vdd.n2319 vdd.n1102 30.449
R3842 vdd.n2579 vdd.n960 30.449
R3843 vdd.n2680 vdd.n2679 30.449
R3844 vdd.n806 vdd.n805 30.449
R3845 vdd.n2807 vdd.n2748 30.449
R3846 vdd.n770 vdd.n769 30.449
R3847 vdd.n2382 vdd.n2381 30.4395
R3848 vdd.n2641 vdd.n958 30.4395
R3849 vdd.n2574 vdd.n961 30.4395
R3850 vdd.n2312 vdd.n2311 30.4395
R3851 vdd.n2814 vdd.n2813 30.4395
R3852 vdd.n3095 vdd.n3092 30.4395
R3853 vdd.n2932 vdd.n2931 30.4395
R3854 vdd.n3156 vdd.n3155 30.4395
R3855 vdd.n3075 vdd.n3074 30.4395
R3856 vdd.n3161 vdd.n771 30.4395
R3857 vdd.n2925 vdd.n2924 30.4395
R3858 vdd.n2936 vdd.n913 30.4395
R3859 vdd.n2386 vdd.n1079 30.4395
R3860 vdd.n2569 vdd.n2568 30.4395
R3861 vdd.n2501 vdd.n2500 30.4395
R3862 vdd.n2201 vdd.n2200 30.4395
R3863 vdd.n1460 vdd.n1226 19.3944
R3864 vdd.n1460 vdd.n1216 19.3944
R3865 vdd.n1472 vdd.n1216 19.3944
R3866 vdd.n1472 vdd.n1214 19.3944
R3867 vdd.n1476 vdd.n1214 19.3944
R3868 vdd.n1476 vdd.n1204 19.3944
R3869 vdd.n1489 vdd.n1204 19.3944
R3870 vdd.n1489 vdd.n1202 19.3944
R3871 vdd.n1493 vdd.n1202 19.3944
R3872 vdd.n1493 vdd.n1194 19.3944
R3873 vdd.n1506 vdd.n1194 19.3944
R3874 vdd.n1506 vdd.n1192 19.3944
R3875 vdd.n1510 vdd.n1192 19.3944
R3876 vdd.n1510 vdd.n1181 19.3944
R3877 vdd.n1522 vdd.n1181 19.3944
R3878 vdd.n1522 vdd.n1179 19.3944
R3879 vdd.n1526 vdd.n1179 19.3944
R3880 vdd.n1526 vdd.n1170 19.3944
R3881 vdd.n1834 vdd.n1170 19.3944
R3882 vdd.n1834 vdd.n1168 19.3944
R3883 vdd.n1838 vdd.n1168 19.3944
R3884 vdd.n1838 vdd.n1159 19.3944
R3885 vdd.n1850 vdd.n1159 19.3944
R3886 vdd.n1850 vdd.n1157 19.3944
R3887 vdd.n1854 vdd.n1157 19.3944
R3888 vdd.n1854 vdd.n1147 19.3944
R3889 vdd.n1867 vdd.n1147 19.3944
R3890 vdd.n1867 vdd.n1145 19.3944
R3891 vdd.n1871 vdd.n1145 19.3944
R3892 vdd.n1871 vdd.n1137 19.3944
R3893 vdd.n1884 vdd.n1137 19.3944
R3894 vdd.n1884 vdd.n1134 19.3944
R3895 vdd.n1890 vdd.n1134 19.3944
R3896 vdd.n1890 vdd.n1135 19.3944
R3897 vdd.n1135 vdd.n1123 19.3944
R3898 vdd.n1379 vdd.n1321 19.3944
R3899 vdd.n1379 vdd.n1378 19.3944
R3900 vdd.n1378 vdd.n1377 19.3944
R3901 vdd.n1377 vdd.n1327 19.3944
R3902 vdd.n1373 vdd.n1327 19.3944
R3903 vdd.n1373 vdd.n1372 19.3944
R3904 vdd.n1372 vdd.n1371 19.3944
R3905 vdd.n1371 vdd.n1333 19.3944
R3906 vdd.n1367 vdd.n1333 19.3944
R3907 vdd.n1367 vdd.n1366 19.3944
R3908 vdd.n1366 vdd.n1365 19.3944
R3909 vdd.n1365 vdd.n1339 19.3944
R3910 vdd.n1361 vdd.n1339 19.3944
R3911 vdd.n1361 vdd.n1360 19.3944
R3912 vdd.n1360 vdd.n1359 19.3944
R3913 vdd.n1359 vdd.n1345 19.3944
R3914 vdd.n1355 vdd.n1345 19.3944
R3915 vdd.n1355 vdd.n1354 19.3944
R3916 vdd.n1354 vdd.n1353 19.3944
R3917 vdd.n1353 vdd.n1351 19.3944
R3918 vdd.n1417 vdd.n1416 19.3944
R3919 vdd.n1416 vdd.n1292 19.3944
R3920 vdd.n1412 vdd.n1292 19.3944
R3921 vdd.n1412 vdd.n1411 19.3944
R3922 vdd.n1411 vdd.n1410 19.3944
R3923 vdd.n1410 vdd.n1298 19.3944
R3924 vdd.n1406 vdd.n1298 19.3944
R3925 vdd.n1406 vdd.n1405 19.3944
R3926 vdd.n1405 vdd.n1404 19.3944
R3927 vdd.n1404 vdd.n1304 19.3944
R3928 vdd.n1400 vdd.n1304 19.3944
R3929 vdd.n1400 vdd.n1399 19.3944
R3930 vdd.n1399 vdd.n1398 19.3944
R3931 vdd.n1398 vdd.n1310 19.3944
R3932 vdd.n1394 vdd.n1310 19.3944
R3933 vdd.n1394 vdd.n1393 19.3944
R3934 vdd.n1393 vdd.n1392 19.3944
R3935 vdd.n1392 vdd.n1316 19.3944
R3936 vdd.n1388 vdd.n1316 19.3944
R3937 vdd.n1388 vdd.n1387 19.3944
R3938 vdd.n1451 vdd.n1450 19.3944
R3939 vdd.n1450 vdd.n1265 19.3944
R3940 vdd.n1446 vdd.n1265 19.3944
R3941 vdd.n1446 vdd.n1445 19.3944
R3942 vdd.n1445 vdd.n1444 19.3944
R3943 vdd.n1444 vdd.n1270 19.3944
R3944 vdd.n1440 vdd.n1270 19.3944
R3945 vdd.n1440 vdd.n1439 19.3944
R3946 vdd.n1439 vdd.n1438 19.3944
R3947 vdd.n1438 vdd.n1276 19.3944
R3948 vdd.n1434 vdd.n1276 19.3944
R3949 vdd.n1434 vdd.n1433 19.3944
R3950 vdd.n1433 vdd.n1432 19.3944
R3951 vdd.n1432 vdd.n1282 19.3944
R3952 vdd.n1428 vdd.n1282 19.3944
R3953 vdd.n1428 vdd.n1427 19.3944
R3954 vdd.n1427 vdd.n1426 19.3944
R3955 vdd.n1426 vdd.n1288 19.3944
R3956 vdd.n2031 vdd.n1966 19.3944
R3957 vdd.n2031 vdd.n1972 19.3944
R3958 vdd.n2026 vdd.n1972 19.3944
R3959 vdd.n2026 vdd.n2025 19.3944
R3960 vdd.n2025 vdd.n2024 19.3944
R3961 vdd.n2024 vdd.n1979 19.3944
R3962 vdd.n2019 vdd.n1979 19.3944
R3963 vdd.n2019 vdd.n2018 19.3944
R3964 vdd.n2018 vdd.n2017 19.3944
R3965 vdd.n2017 vdd.n1986 19.3944
R3966 vdd.n2012 vdd.n1986 19.3944
R3967 vdd.n2012 vdd.n2011 19.3944
R3968 vdd.n2011 vdd.n2010 19.3944
R3969 vdd.n2010 vdd.n1994 19.3944
R3970 vdd.n2005 vdd.n1994 19.3944
R3971 vdd.n2005 vdd.n2004 19.3944
R3972 vdd.n2000 vdd.n1999 19.3944
R3973 vdd.n2120 vdd.n1119 19.3944
R3974 vdd.n2070 vdd.n1926 19.3944
R3975 vdd.n2070 vdd.n1932 19.3944
R3976 vdd.n2065 vdd.n1932 19.3944
R3977 vdd.n2065 vdd.n2064 19.3944
R3978 vdd.n2064 vdd.n2063 19.3944
R3979 vdd.n2063 vdd.n1939 19.3944
R3980 vdd.n2058 vdd.n1939 19.3944
R3981 vdd.n2058 vdd.n2057 19.3944
R3982 vdd.n2057 vdd.n2056 19.3944
R3983 vdd.n2056 vdd.n1946 19.3944
R3984 vdd.n2051 vdd.n1946 19.3944
R3985 vdd.n2051 vdd.n2050 19.3944
R3986 vdd.n2050 vdd.n2049 19.3944
R3987 vdd.n2049 vdd.n1953 19.3944
R3988 vdd.n2044 vdd.n1953 19.3944
R3989 vdd.n2044 vdd.n2043 19.3944
R3990 vdd.n2043 vdd.n2042 19.3944
R3991 vdd.n2042 vdd.n1960 19.3944
R3992 vdd.n2037 vdd.n1960 19.3944
R3993 vdd.n2037 vdd.n2036 19.3944
R3994 vdd.n2108 vdd.n2107 19.3944
R3995 vdd.n2107 vdd.n1898 19.3944
R3996 vdd.n2102 vdd.n2101 19.3944
R3997 vdd.n2097 vdd.n1902 19.3944
R3998 vdd.n2097 vdd.n1904 19.3944
R3999 vdd.n1907 vdd.n1904 19.3944
R4000 vdd.n2090 vdd.n1907 19.3944
R4001 vdd.n2090 vdd.n2089 19.3944
R4002 vdd.n2089 vdd.n2088 19.3944
R4003 vdd.n2088 vdd.n1913 19.3944
R4004 vdd.n2083 vdd.n1913 19.3944
R4005 vdd.n2083 vdd.n2082 19.3944
R4006 vdd.n2082 vdd.n2081 19.3944
R4007 vdd.n2081 vdd.n1920 19.3944
R4008 vdd.n2076 vdd.n1920 19.3944
R4009 vdd.n2076 vdd.n2075 19.3944
R4010 vdd.n1464 vdd.n1222 19.3944
R4011 vdd.n1464 vdd.n1220 19.3944
R4012 vdd.n1468 vdd.n1220 19.3944
R4013 vdd.n1468 vdd.n1210 19.3944
R4014 vdd.n1481 vdd.n1210 19.3944
R4015 vdd.n1481 vdd.n1208 19.3944
R4016 vdd.n1485 vdd.n1208 19.3944
R4017 vdd.n1485 vdd.n1199 19.3944
R4018 vdd.n1498 vdd.n1199 19.3944
R4019 vdd.n1498 vdd.n1197 19.3944
R4020 vdd.n1502 vdd.n1197 19.3944
R4021 vdd.n1502 vdd.n1188 19.3944
R4022 vdd.n1514 vdd.n1188 19.3944
R4023 vdd.n1514 vdd.n1186 19.3944
R4024 vdd.n1518 vdd.n1186 19.3944
R4025 vdd.n1518 vdd.n1176 19.3944
R4026 vdd.n1531 vdd.n1176 19.3944
R4027 vdd.n1531 vdd.n1174 19.3944
R4028 vdd.n1830 vdd.n1174 19.3944
R4029 vdd.n1830 vdd.n1165 19.3944
R4030 vdd.n1842 vdd.n1165 19.3944
R4031 vdd.n1842 vdd.n1163 19.3944
R4032 vdd.n1846 vdd.n1163 19.3944
R4033 vdd.n1846 vdd.n1153 19.3944
R4034 vdd.n1859 vdd.n1153 19.3944
R4035 vdd.n1859 vdd.n1151 19.3944
R4036 vdd.n1863 vdd.n1151 19.3944
R4037 vdd.n1863 vdd.n1142 19.3944
R4038 vdd.n1876 vdd.n1142 19.3944
R4039 vdd.n1876 vdd.n1140 19.3944
R4040 vdd.n1880 vdd.n1140 19.3944
R4041 vdd.n1880 vdd.n1130 19.3944
R4042 vdd.n1894 vdd.n1130 19.3944
R4043 vdd.n1894 vdd.n1128 19.3944
R4044 vdd.n2111 vdd.n1128 19.3944
R4045 vdd.n3329 vdd.n655 19.3944
R4046 vdd.n3333 vdd.n655 19.3944
R4047 vdd.n3333 vdd.n646 19.3944
R4048 vdd.n3345 vdd.n646 19.3944
R4049 vdd.n3345 vdd.n644 19.3944
R4050 vdd.n3349 vdd.n644 19.3944
R4051 vdd.n3349 vdd.n633 19.3944
R4052 vdd.n3361 vdd.n633 19.3944
R4053 vdd.n3361 vdd.n631 19.3944
R4054 vdd.n3365 vdd.n631 19.3944
R4055 vdd.n3365 vdd.n622 19.3944
R4056 vdd.n3378 vdd.n622 19.3944
R4057 vdd.n3378 vdd.n620 19.3944
R4058 vdd.n3385 vdd.n620 19.3944
R4059 vdd.n3385 vdd.n3384 19.3944
R4060 vdd.n3384 vdd.n610 19.3944
R4061 vdd.n3398 vdd.n610 19.3944
R4062 vdd.n3399 vdd.n3398 19.3944
R4063 vdd.n3400 vdd.n3399 19.3944
R4064 vdd.n3400 vdd.n608 19.3944
R4065 vdd.n3405 vdd.n608 19.3944
R4066 vdd.n3406 vdd.n3405 19.3944
R4067 vdd.n3407 vdd.n3406 19.3944
R4068 vdd.n3407 vdd.n606 19.3944
R4069 vdd.n3412 vdd.n606 19.3944
R4070 vdd.n3413 vdd.n3412 19.3944
R4071 vdd.n3414 vdd.n3413 19.3944
R4072 vdd.n3414 vdd.n604 19.3944
R4073 vdd.n3420 vdd.n604 19.3944
R4074 vdd.n3421 vdd.n3420 19.3944
R4075 vdd.n3422 vdd.n3421 19.3944
R4076 vdd.n3422 vdd.n602 19.3944
R4077 vdd.n3427 vdd.n602 19.3944
R4078 vdd.n3428 vdd.n3427 19.3944
R4079 vdd.n3429 vdd.n3428 19.3944
R4080 vdd.n550 vdd.n417 19.3944
R4081 vdd.n556 vdd.n417 19.3944
R4082 vdd.n557 vdd.n556 19.3944
R4083 vdd.n560 vdd.n557 19.3944
R4084 vdd.n560 vdd.n415 19.3944
R4085 vdd.n566 vdd.n415 19.3944
R4086 vdd.n567 vdd.n566 19.3944
R4087 vdd.n570 vdd.n567 19.3944
R4088 vdd.n570 vdd.n413 19.3944
R4089 vdd.n576 vdd.n413 19.3944
R4090 vdd.n577 vdd.n576 19.3944
R4091 vdd.n580 vdd.n577 19.3944
R4092 vdd.n580 vdd.n411 19.3944
R4093 vdd.n586 vdd.n411 19.3944
R4094 vdd.n587 vdd.n586 19.3944
R4095 vdd.n590 vdd.n587 19.3944
R4096 vdd.n590 vdd.n409 19.3944
R4097 vdd.n596 vdd.n409 19.3944
R4098 vdd.n598 vdd.n596 19.3944
R4099 vdd.n599 vdd.n598 19.3944
R4100 vdd.n497 vdd.n496 19.3944
R4101 vdd.n500 vdd.n497 19.3944
R4102 vdd.n500 vdd.n429 19.3944
R4103 vdd.n506 vdd.n429 19.3944
R4104 vdd.n507 vdd.n506 19.3944
R4105 vdd.n510 vdd.n507 19.3944
R4106 vdd.n510 vdd.n427 19.3944
R4107 vdd.n516 vdd.n427 19.3944
R4108 vdd.n517 vdd.n516 19.3944
R4109 vdd.n520 vdd.n517 19.3944
R4110 vdd.n520 vdd.n425 19.3944
R4111 vdd.n526 vdd.n425 19.3944
R4112 vdd.n527 vdd.n526 19.3944
R4113 vdd.n530 vdd.n527 19.3944
R4114 vdd.n530 vdd.n423 19.3944
R4115 vdd.n536 vdd.n423 19.3944
R4116 vdd.n537 vdd.n536 19.3944
R4117 vdd.n540 vdd.n537 19.3944
R4118 vdd.n540 vdd.n421 19.3944
R4119 vdd.n546 vdd.n421 19.3944
R4120 vdd.n447 vdd.n446 19.3944
R4121 vdd.n450 vdd.n447 19.3944
R4122 vdd.n450 vdd.n441 19.3944
R4123 vdd.n456 vdd.n441 19.3944
R4124 vdd.n457 vdd.n456 19.3944
R4125 vdd.n460 vdd.n457 19.3944
R4126 vdd.n460 vdd.n439 19.3944
R4127 vdd.n466 vdd.n439 19.3944
R4128 vdd.n467 vdd.n466 19.3944
R4129 vdd.n470 vdd.n467 19.3944
R4130 vdd.n470 vdd.n437 19.3944
R4131 vdd.n476 vdd.n437 19.3944
R4132 vdd.n477 vdd.n476 19.3944
R4133 vdd.n480 vdd.n477 19.3944
R4134 vdd.n480 vdd.n435 19.3944
R4135 vdd.n486 vdd.n435 19.3944
R4136 vdd.n487 vdd.n486 19.3944
R4137 vdd.n490 vdd.n487 19.3944
R4138 vdd.n3325 vdd.n652 19.3944
R4139 vdd.n3337 vdd.n652 19.3944
R4140 vdd.n3337 vdd.n650 19.3944
R4141 vdd.n3341 vdd.n650 19.3944
R4142 vdd.n3341 vdd.n640 19.3944
R4143 vdd.n3353 vdd.n640 19.3944
R4144 vdd.n3353 vdd.n638 19.3944
R4145 vdd.n3357 vdd.n638 19.3944
R4146 vdd.n3357 vdd.n628 19.3944
R4147 vdd.n3370 vdd.n628 19.3944
R4148 vdd.n3370 vdd.n626 19.3944
R4149 vdd.n3374 vdd.n626 19.3944
R4150 vdd.n3374 vdd.n617 19.3944
R4151 vdd.n3389 vdd.n617 19.3944
R4152 vdd.n3389 vdd.n615 19.3944
R4153 vdd.n3393 vdd.n615 19.3944
R4154 vdd.n3393 vdd.n324 19.3944
R4155 vdd.n3471 vdd.n324 19.3944
R4156 vdd.n3471 vdd.n325 19.3944
R4157 vdd.n3465 vdd.n325 19.3944
R4158 vdd.n3465 vdd.n3464 19.3944
R4159 vdd.n3464 vdd.n3463 19.3944
R4160 vdd.n3463 vdd.n337 19.3944
R4161 vdd.n3457 vdd.n337 19.3944
R4162 vdd.n3457 vdd.n3456 19.3944
R4163 vdd.n3456 vdd.n3455 19.3944
R4164 vdd.n3455 vdd.n347 19.3944
R4165 vdd.n3449 vdd.n347 19.3944
R4166 vdd.n3449 vdd.n3448 19.3944
R4167 vdd.n3448 vdd.n3447 19.3944
R4168 vdd.n3447 vdd.n358 19.3944
R4169 vdd.n3441 vdd.n358 19.3944
R4170 vdd.n3441 vdd.n3440 19.3944
R4171 vdd.n3440 vdd.n3439 19.3944
R4172 vdd.n3439 vdd.n369 19.3944
R4173 vdd.n3282 vdd.n3281 19.3944
R4174 vdd.n3281 vdd.n3280 19.3944
R4175 vdd.n3280 vdd.n694 19.3944
R4176 vdd.n3274 vdd.n694 19.3944
R4177 vdd.n3274 vdd.n3273 19.3944
R4178 vdd.n3273 vdd.n3272 19.3944
R4179 vdd.n3272 vdd.n700 19.3944
R4180 vdd.n3266 vdd.n700 19.3944
R4181 vdd.n3266 vdd.n3265 19.3944
R4182 vdd.n3265 vdd.n3264 19.3944
R4183 vdd.n3264 vdd.n706 19.3944
R4184 vdd.n3258 vdd.n706 19.3944
R4185 vdd.n3258 vdd.n3257 19.3944
R4186 vdd.n3257 vdd.n3256 19.3944
R4187 vdd.n3256 vdd.n712 19.3944
R4188 vdd.n3250 vdd.n712 19.3944
R4189 vdd.n3250 vdd.n3249 19.3944
R4190 vdd.n3249 vdd.n3248 19.3944
R4191 vdd.n3248 vdd.n718 19.3944
R4192 vdd.n3242 vdd.n718 19.3944
R4193 vdd.n3322 vdd.n3321 19.3944
R4194 vdd.n3321 vdd.n662 19.3944
R4195 vdd.n3316 vdd.n3315 19.3944
R4196 vdd.n3312 vdd.n3311 19.3944
R4197 vdd.n3311 vdd.n668 19.3944
R4198 vdd.n3306 vdd.n668 19.3944
R4199 vdd.n3306 vdd.n3305 19.3944
R4200 vdd.n3305 vdd.n3304 19.3944
R4201 vdd.n3304 vdd.n674 19.3944
R4202 vdd.n3298 vdd.n674 19.3944
R4203 vdd.n3298 vdd.n3297 19.3944
R4204 vdd.n3297 vdd.n3296 19.3944
R4205 vdd.n3296 vdd.n680 19.3944
R4206 vdd.n3290 vdd.n680 19.3944
R4207 vdd.n3290 vdd.n3289 19.3944
R4208 vdd.n3289 vdd.n3288 19.3944
R4209 vdd.n3237 vdd.n722 19.3944
R4210 vdd.n3237 vdd.n726 19.3944
R4211 vdd.n3232 vdd.n726 19.3944
R4212 vdd.n3232 vdd.n3231 19.3944
R4213 vdd.n3231 vdd.n732 19.3944
R4214 vdd.n3226 vdd.n732 19.3944
R4215 vdd.n3226 vdd.n3225 19.3944
R4216 vdd.n3225 vdd.n3224 19.3944
R4217 vdd.n3224 vdd.n738 19.3944
R4218 vdd.n3218 vdd.n738 19.3944
R4219 vdd.n3218 vdd.n3217 19.3944
R4220 vdd.n3217 vdd.n3216 19.3944
R4221 vdd.n3216 vdd.n744 19.3944
R4222 vdd.n3210 vdd.n744 19.3944
R4223 vdd.n3210 vdd.n3209 19.3944
R4224 vdd.n3209 vdd.n3208 19.3944
R4225 vdd.n3204 vdd.n3203 19.3944
R4226 vdd.n3200 vdd.n3199 19.3944
R4227 vdd.n1386 vdd.n1321 19.0066
R4228 vdd.n2035 vdd.n1966 19.0066
R4229 vdd.n550 vdd.n547 19.0066
R4230 vdd.n3241 vdd.n722 19.0066
R4231 vdd.n1454 vdd.n1224 18.5924
R4232 vdd.n2113 vdd.n1125 18.5924
R4233 vdd.n3327 vdd.n658 18.5924
R4234 vdd.n3436 vdd.n3435 18.5924
R4235 vdd.n1108 vdd.n1107 16.0975
R4236 vdd.n969 vdd.n968 16.0975
R4237 vdd.n1229 vdd.n1228 16.0975
R4238 vdd.n1385 vdd.n1384 16.0975
R4239 vdd.n1421 vdd.n1420 16.0975
R4240 vdd.n2118 vdd.n2117 16.0975
R4241 vdd.n1968 vdd.n1967 16.0975
R4242 vdd.n1928 vdd.n1927 16.0975
R4243 vdd.n1102 vdd.n1101 16.0975
R4244 vdd.n960 vdd.n959 16.0975
R4245 vdd.n2679 vdd.n2678 16.0975
R4246 vdd.n406 vdd.n405 16.0975
R4247 vdd.n420 vdd.n419 16.0975
R4248 vdd.n432 vdd.n431 16.0975
R4249 vdd.n724 vdd.n723 16.0975
R4250 vdd.n687 vdd.n686 16.0975
R4251 vdd.n805 vdd.n804 16.0975
R4252 vdd.n2748 vdd.n2747 16.0975
R4253 vdd.n3196 vdd.n3195 16.0975
R4254 vdd.n769 vdd.n768 16.0975
R4255 vdd.t111 vdd.n2643 15.4182
R4256 vdd.n2927 vdd.t119 15.4182
R4257 vdd.n28 vdd.n27 14.8356
R4258 vdd.n2384 vdd.n1081 13.6043
R4259 vdd.n3158 vdd.n756 13.6043
R4260 vdd.n316 vdd.n281 13.1884
R4261 vdd.n261 vdd.n226 13.1884
R4262 vdd.n218 vdd.n183 13.1884
R4263 vdd.n163 vdd.n128 13.1884
R4264 vdd.n121 vdd.n86 13.1884
R4265 vdd.n66 vdd.n31 13.1884
R4266 vdd.n1765 vdd.n1730 13.1884
R4267 vdd.n1820 vdd.n1785 13.1884
R4268 vdd.n1667 vdd.n1632 13.1884
R4269 vdd.n1722 vdd.n1687 13.1884
R4270 vdd.n1570 vdd.n1535 13.1884
R4271 vdd.n1625 vdd.n1590 13.1884
R4272 vdd.n1422 vdd.n1417 12.9944
R4273 vdd.n1422 vdd.n1288 12.9944
R4274 vdd.n2074 vdd.n1926 12.9944
R4275 vdd.n2075 vdd.n2074 12.9944
R4276 vdd.n496 vdd.n433 12.9944
R4277 vdd.n490 vdd.n433 12.9944
R4278 vdd.n3282 vdd.n688 12.9944
R4279 vdd.n3288 vdd.n688 12.9944
R4280 vdd.n317 vdd.n279 12.8005
R4281 vdd.n312 vdd.n283 12.8005
R4282 vdd.n262 vdd.n224 12.8005
R4283 vdd.n257 vdd.n228 12.8005
R4284 vdd.n219 vdd.n181 12.8005
R4285 vdd.n214 vdd.n185 12.8005
R4286 vdd.n164 vdd.n126 12.8005
R4287 vdd.n159 vdd.n130 12.8005
R4288 vdd.n122 vdd.n84 12.8005
R4289 vdd.n117 vdd.n88 12.8005
R4290 vdd.n67 vdd.n29 12.8005
R4291 vdd.n62 vdd.n33 12.8005
R4292 vdd.n1766 vdd.n1728 12.8005
R4293 vdd.n1761 vdd.n1732 12.8005
R4294 vdd.n1821 vdd.n1783 12.8005
R4295 vdd.n1816 vdd.n1787 12.8005
R4296 vdd.n1668 vdd.n1630 12.8005
R4297 vdd.n1663 vdd.n1634 12.8005
R4298 vdd.n1723 vdd.n1685 12.8005
R4299 vdd.n1718 vdd.n1689 12.8005
R4300 vdd.n1571 vdd.n1533 12.8005
R4301 vdd.n1566 vdd.n1537 12.8005
R4302 vdd.n1626 vdd.n1588 12.8005
R4303 vdd.n1621 vdd.n1592 12.8005
R4304 vdd.n311 vdd.n284 12.0247
R4305 vdd.n256 vdd.n229 12.0247
R4306 vdd.n213 vdd.n186 12.0247
R4307 vdd.n158 vdd.n131 12.0247
R4308 vdd.n116 vdd.n89 12.0247
R4309 vdd.n61 vdd.n34 12.0247
R4310 vdd.n1760 vdd.n1733 12.0247
R4311 vdd.n1815 vdd.n1788 12.0247
R4312 vdd.n1662 vdd.n1635 12.0247
R4313 vdd.n1717 vdd.n1690 12.0247
R4314 vdd.n1565 vdd.n1538 12.0247
R4315 vdd.n1620 vdd.n1593 12.0247
R4316 vdd.n1462 vdd.n1224 11.337
R4317 vdd.n1470 vdd.n1218 11.337
R4318 vdd.n1470 vdd.n1212 11.337
R4319 vdd.n1479 vdd.n1212 11.337
R4320 vdd.n1487 vdd.n1206 11.337
R4321 vdd.n1496 vdd.n1495 11.337
R4322 vdd.n1512 vdd.n1190 11.337
R4323 vdd.n1520 vdd.n1183 11.337
R4324 vdd.n1529 vdd.n1528 11.337
R4325 vdd.n1832 vdd.n1172 11.337
R4326 vdd.n1848 vdd.n1161 11.337
R4327 vdd.n1857 vdd.n1155 11.337
R4328 vdd.n1865 vdd.n1149 11.337
R4329 vdd.n1874 vdd.n1873 11.337
R4330 vdd.n1882 vdd.n1132 11.337
R4331 vdd.n1892 vdd.n1132 11.337
R4332 vdd.n2113 vdd.n1124 11.337
R4333 vdd.n3327 vdd.n659 11.337
R4334 vdd.n3335 vdd.n648 11.337
R4335 vdd.n3343 vdd.n648 11.337
R4336 vdd.n3351 vdd.n642 11.337
R4337 vdd.n3359 vdd.n635 11.337
R4338 vdd.n3368 vdd.n3367 11.337
R4339 vdd.n3376 vdd.n624 11.337
R4340 vdd.n3395 vdd.n613 11.337
R4341 vdd.n3469 vdd.n328 11.337
R4342 vdd.n3467 vdd.n332 11.337
R4343 vdd.n3461 vdd.n3460 11.337
R4344 vdd.n3453 vdd.n349 11.337
R4345 vdd.n3452 vdd.n3451 11.337
R4346 vdd.n3445 vdd.n3444 11.337
R4347 vdd.n3444 vdd.n3443 11.337
R4348 vdd.n3443 vdd.n363 11.337
R4349 vdd.n3437 vdd.n3436 11.337
R4350 vdd.n308 vdd.n307 11.249
R4351 vdd.n253 vdd.n252 11.249
R4352 vdd.n210 vdd.n209 11.249
R4353 vdd.n155 vdd.n154 11.249
R4354 vdd.n113 vdd.n112 11.249
R4355 vdd.n58 vdd.n57 11.249
R4356 vdd.n1757 vdd.n1756 11.249
R4357 vdd.n1812 vdd.n1811 11.249
R4358 vdd.n1659 vdd.n1658 11.249
R4359 vdd.n1714 vdd.n1713 11.249
R4360 vdd.n1562 vdd.n1561 11.249
R4361 vdd.n1617 vdd.n1616 11.249
R4362 vdd.n1882 vdd.t214 10.7702
R4363 vdd.n3343 vdd.t182 10.7702
R4364 vdd.n293 vdd.n292 10.7238
R4365 vdd.n238 vdd.n237 10.7238
R4366 vdd.n195 vdd.n194 10.7238
R4367 vdd.n140 vdd.n139 10.7238
R4368 vdd.n98 vdd.n97 10.7238
R4369 vdd.n43 vdd.n42 10.7238
R4370 vdd.n1742 vdd.n1741 10.7238
R4371 vdd.n1797 vdd.n1796 10.7238
R4372 vdd.n1644 vdd.n1643 10.7238
R4373 vdd.n1699 vdd.n1698 10.7238
R4374 vdd.n1547 vdd.n1546 10.7238
R4375 vdd.n1602 vdd.n1601 10.7238
R4376 vdd.n2382 vdd.n1073 10.6151
R4377 vdd.n2392 vdd.n1073 10.6151
R4378 vdd.n2393 vdd.n2392 10.6151
R4379 vdd.n2394 vdd.n2393 10.6151
R4380 vdd.n2394 vdd.n1061 10.6151
R4381 vdd.n2404 vdd.n1061 10.6151
R4382 vdd.n2405 vdd.n2404 10.6151
R4383 vdd.n2406 vdd.n2405 10.6151
R4384 vdd.n2406 vdd.n1049 10.6151
R4385 vdd.n2416 vdd.n1049 10.6151
R4386 vdd.n2417 vdd.n2416 10.6151
R4387 vdd.n2418 vdd.n2417 10.6151
R4388 vdd.n2418 vdd.n1036 10.6151
R4389 vdd.n2428 vdd.n1036 10.6151
R4390 vdd.n2429 vdd.n2428 10.6151
R4391 vdd.n2430 vdd.n2429 10.6151
R4392 vdd.n2430 vdd.n1024 10.6151
R4393 vdd.n2441 vdd.n1024 10.6151
R4394 vdd.n2442 vdd.n2441 10.6151
R4395 vdd.n2443 vdd.n2442 10.6151
R4396 vdd.n2443 vdd.n1012 10.6151
R4397 vdd.n2453 vdd.n1012 10.6151
R4398 vdd.n2454 vdd.n2453 10.6151
R4399 vdd.n2455 vdd.n2454 10.6151
R4400 vdd.n2455 vdd.n1000 10.6151
R4401 vdd.n2465 vdd.n1000 10.6151
R4402 vdd.n2466 vdd.n2465 10.6151
R4403 vdd.n2467 vdd.n2466 10.6151
R4404 vdd.n2467 vdd.n990 10.6151
R4405 vdd.n2477 vdd.n990 10.6151
R4406 vdd.n2478 vdd.n2477 10.6151
R4407 vdd.n2479 vdd.n2478 10.6151
R4408 vdd.n2479 vdd.n977 10.6151
R4409 vdd.n2491 vdd.n977 10.6151
R4410 vdd.n2492 vdd.n2491 10.6151
R4411 vdd.n2494 vdd.n2492 10.6151
R4412 vdd.n2494 vdd.n2493 10.6151
R4413 vdd.n2493 vdd.n958 10.6151
R4414 vdd.n2641 vdd.n2640 10.6151
R4415 vdd.n2640 vdd.n2639 10.6151
R4416 vdd.n2639 vdd.n2636 10.6151
R4417 vdd.n2636 vdd.n2635 10.6151
R4418 vdd.n2635 vdd.n2632 10.6151
R4419 vdd.n2632 vdd.n2631 10.6151
R4420 vdd.n2631 vdd.n2628 10.6151
R4421 vdd.n2628 vdd.n2627 10.6151
R4422 vdd.n2627 vdd.n2624 10.6151
R4423 vdd.n2624 vdd.n2623 10.6151
R4424 vdd.n2623 vdd.n2620 10.6151
R4425 vdd.n2620 vdd.n2619 10.6151
R4426 vdd.n2619 vdd.n2616 10.6151
R4427 vdd.n2616 vdd.n2615 10.6151
R4428 vdd.n2615 vdd.n2612 10.6151
R4429 vdd.n2612 vdd.n2611 10.6151
R4430 vdd.n2611 vdd.n2608 10.6151
R4431 vdd.n2608 vdd.n2607 10.6151
R4432 vdd.n2607 vdd.n2604 10.6151
R4433 vdd.n2604 vdd.n2603 10.6151
R4434 vdd.n2603 vdd.n2600 10.6151
R4435 vdd.n2600 vdd.n2599 10.6151
R4436 vdd.n2599 vdd.n2596 10.6151
R4437 vdd.n2596 vdd.n2595 10.6151
R4438 vdd.n2595 vdd.n2592 10.6151
R4439 vdd.n2592 vdd.n2591 10.6151
R4440 vdd.n2591 vdd.n2588 10.6151
R4441 vdd.n2588 vdd.n2587 10.6151
R4442 vdd.n2587 vdd.n2584 10.6151
R4443 vdd.n2584 vdd.n2583 10.6151
R4444 vdd.n2583 vdd.n2580 10.6151
R4445 vdd.n2578 vdd.n2575 10.6151
R4446 vdd.n2575 vdd.n2574 10.6151
R4447 vdd.n2311 vdd.n2310 10.6151
R4448 vdd.n2310 vdd.n2308 10.6151
R4449 vdd.n2308 vdd.n2307 10.6151
R4450 vdd.n2307 vdd.n2305 10.6151
R4451 vdd.n2305 vdd.n2304 10.6151
R4452 vdd.n2304 vdd.n2302 10.6151
R4453 vdd.n2302 vdd.n2301 10.6151
R4454 vdd.n2301 vdd.n2299 10.6151
R4455 vdd.n2299 vdd.n2298 10.6151
R4456 vdd.n2298 vdd.n2296 10.6151
R4457 vdd.n2296 vdd.n2295 10.6151
R4458 vdd.n2295 vdd.n2293 10.6151
R4459 vdd.n2293 vdd.n2292 10.6151
R4460 vdd.n2292 vdd.n2290 10.6151
R4461 vdd.n2290 vdd.n2289 10.6151
R4462 vdd.n2289 vdd.n2287 10.6151
R4463 vdd.n2287 vdd.n2286 10.6151
R4464 vdd.n2286 vdd.n2284 10.6151
R4465 vdd.n2284 vdd.n2283 10.6151
R4466 vdd.n2283 vdd.n2281 10.6151
R4467 vdd.n2281 vdd.n2280 10.6151
R4468 vdd.n2280 vdd.n2278 10.6151
R4469 vdd.n2278 vdd.n2277 10.6151
R4470 vdd.n2277 vdd.n1104 10.6151
R4471 vdd.n2244 vdd.n1104 10.6151
R4472 vdd.n2245 vdd.n2244 10.6151
R4473 vdd.n2247 vdd.n2245 10.6151
R4474 vdd.n2248 vdd.n2247 10.6151
R4475 vdd.n2261 vdd.n2248 10.6151
R4476 vdd.n2261 vdd.n2260 10.6151
R4477 vdd.n2260 vdd.n2259 10.6151
R4478 vdd.n2259 vdd.n2257 10.6151
R4479 vdd.n2257 vdd.n2256 10.6151
R4480 vdd.n2256 vdd.n2254 10.6151
R4481 vdd.n2254 vdd.n2253 10.6151
R4482 vdd.n2253 vdd.n2250 10.6151
R4483 vdd.n2250 vdd.n2249 10.6151
R4484 vdd.n2249 vdd.n961 10.6151
R4485 vdd.n2381 vdd.n2380 10.6151
R4486 vdd.n2380 vdd.n1085 10.6151
R4487 vdd.n2375 vdd.n1085 10.6151
R4488 vdd.n2375 vdd.n2374 10.6151
R4489 vdd.n2374 vdd.n1087 10.6151
R4490 vdd.n2369 vdd.n1087 10.6151
R4491 vdd.n2369 vdd.n2368 10.6151
R4492 vdd.n2368 vdd.n2367 10.6151
R4493 vdd.n2367 vdd.n1089 10.6151
R4494 vdd.n2361 vdd.n1089 10.6151
R4495 vdd.n2361 vdd.n2360 10.6151
R4496 vdd.n2360 vdd.n2359 10.6151
R4497 vdd.n2359 vdd.n1091 10.6151
R4498 vdd.n2353 vdd.n1091 10.6151
R4499 vdd.n2353 vdd.n2352 10.6151
R4500 vdd.n2352 vdd.n2351 10.6151
R4501 vdd.n2351 vdd.n1093 10.6151
R4502 vdd.n2345 vdd.n1093 10.6151
R4503 vdd.n2345 vdd.n2344 10.6151
R4504 vdd.n2344 vdd.n2343 10.6151
R4505 vdd.n2343 vdd.n1095 10.6151
R4506 vdd.n2337 vdd.n1095 10.6151
R4507 vdd.n2337 vdd.n2336 10.6151
R4508 vdd.n2336 vdd.n2335 10.6151
R4509 vdd.n2335 vdd.n1097 10.6151
R4510 vdd.n2329 vdd.n1097 10.6151
R4511 vdd.n2329 vdd.n2328 10.6151
R4512 vdd.n2328 vdd.n2327 10.6151
R4513 vdd.n2327 vdd.n1099 10.6151
R4514 vdd.n2321 vdd.n1099 10.6151
R4515 vdd.n2321 vdd.n2320 10.6151
R4516 vdd.n2318 vdd.n1103 10.6151
R4517 vdd.n2312 vdd.n1103 10.6151
R4518 vdd.n2816 vdd.n2814 10.6151
R4519 vdd.n2817 vdd.n2816 10.6151
R4520 vdd.n2916 vdd.n2817 10.6151
R4521 vdd.n2916 vdd.n2915 10.6151
R4522 vdd.n2915 vdd.n2914 10.6151
R4523 vdd.n2914 vdd.n2912 10.6151
R4524 vdd.n2912 vdd.n2911 10.6151
R4525 vdd.n2911 vdd.n2909 10.6151
R4526 vdd.n2909 vdd.n2908 10.6151
R4527 vdd.n2908 vdd.n2818 10.6151
R4528 vdd.n2858 vdd.n2818 10.6151
R4529 vdd.n2859 vdd.n2858 10.6151
R4530 vdd.n2861 vdd.n2859 10.6151
R4531 vdd.n2862 vdd.n2861 10.6151
R4532 vdd.n2892 vdd.n2862 10.6151
R4533 vdd.n2892 vdd.n2891 10.6151
R4534 vdd.n2891 vdd.n2890 10.6151
R4535 vdd.n2890 vdd.n2888 10.6151
R4536 vdd.n2888 vdd.n2887 10.6151
R4537 vdd.n2887 vdd.n2885 10.6151
R4538 vdd.n2885 vdd.n2884 10.6151
R4539 vdd.n2884 vdd.n2882 10.6151
R4540 vdd.n2882 vdd.n2881 10.6151
R4541 vdd.n2881 vdd.n2879 10.6151
R4542 vdd.n2879 vdd.n2878 10.6151
R4543 vdd.n2878 vdd.n2876 10.6151
R4544 vdd.n2876 vdd.n2875 10.6151
R4545 vdd.n2875 vdd.n2873 10.6151
R4546 vdd.n2873 vdd.n2872 10.6151
R4547 vdd.n2872 vdd.n2870 10.6151
R4548 vdd.n2870 vdd.n2869 10.6151
R4549 vdd.n2869 vdd.n2867 10.6151
R4550 vdd.n2867 vdd.n2866 10.6151
R4551 vdd.n2866 vdd.n2864 10.6151
R4552 vdd.n2864 vdd.n2863 10.6151
R4553 vdd.n2863 vdd.n807 10.6151
R4554 vdd.n3091 vdd.n807 10.6151
R4555 vdd.n3092 vdd.n3091 10.6151
R4556 vdd.n2931 vdd.n2930 10.6151
R4557 vdd.n2930 vdd.n919 10.6151
R4558 vdd.n2750 vdd.n919 10.6151
R4559 vdd.n2751 vdd.n2750 10.6151
R4560 vdd.n2754 vdd.n2751 10.6151
R4561 vdd.n2755 vdd.n2754 10.6151
R4562 vdd.n2758 vdd.n2755 10.6151
R4563 vdd.n2759 vdd.n2758 10.6151
R4564 vdd.n2762 vdd.n2759 10.6151
R4565 vdd.n2763 vdd.n2762 10.6151
R4566 vdd.n2766 vdd.n2763 10.6151
R4567 vdd.n2767 vdd.n2766 10.6151
R4568 vdd.n2770 vdd.n2767 10.6151
R4569 vdd.n2771 vdd.n2770 10.6151
R4570 vdd.n2774 vdd.n2771 10.6151
R4571 vdd.n2775 vdd.n2774 10.6151
R4572 vdd.n2778 vdd.n2775 10.6151
R4573 vdd.n2779 vdd.n2778 10.6151
R4574 vdd.n2782 vdd.n2779 10.6151
R4575 vdd.n2783 vdd.n2782 10.6151
R4576 vdd.n2786 vdd.n2783 10.6151
R4577 vdd.n2787 vdd.n2786 10.6151
R4578 vdd.n2790 vdd.n2787 10.6151
R4579 vdd.n2791 vdd.n2790 10.6151
R4580 vdd.n2794 vdd.n2791 10.6151
R4581 vdd.n2795 vdd.n2794 10.6151
R4582 vdd.n2798 vdd.n2795 10.6151
R4583 vdd.n2799 vdd.n2798 10.6151
R4584 vdd.n2802 vdd.n2799 10.6151
R4585 vdd.n2803 vdd.n2802 10.6151
R4586 vdd.n2806 vdd.n2803 10.6151
R4587 vdd.n2811 vdd.n2808 10.6151
R4588 vdd.n2813 vdd.n2811 10.6151
R4589 vdd.n2932 vdd.n908 10.6151
R4590 vdd.n2942 vdd.n908 10.6151
R4591 vdd.n2943 vdd.n2942 10.6151
R4592 vdd.n2944 vdd.n2943 10.6151
R4593 vdd.n2944 vdd.n896 10.6151
R4594 vdd.n2954 vdd.n896 10.6151
R4595 vdd.n2955 vdd.n2954 10.6151
R4596 vdd.n2956 vdd.n2955 10.6151
R4597 vdd.n2956 vdd.n886 10.6151
R4598 vdd.n2966 vdd.n886 10.6151
R4599 vdd.n2967 vdd.n2966 10.6151
R4600 vdd.n2968 vdd.n2967 10.6151
R4601 vdd.n2968 vdd.n874 10.6151
R4602 vdd.n2978 vdd.n874 10.6151
R4603 vdd.n2979 vdd.n2978 10.6151
R4604 vdd.n2980 vdd.n2979 10.6151
R4605 vdd.n2980 vdd.n863 10.6151
R4606 vdd.n2990 vdd.n863 10.6151
R4607 vdd.n2991 vdd.n2990 10.6151
R4608 vdd.n2992 vdd.n2991 10.6151
R4609 vdd.n2992 vdd.n850 10.6151
R4610 vdd.n3003 vdd.n850 10.6151
R4611 vdd.n3004 vdd.n3003 10.6151
R4612 vdd.n3005 vdd.n3004 10.6151
R4613 vdd.n3005 vdd.n837 10.6151
R4614 vdd.n3015 vdd.n837 10.6151
R4615 vdd.n3016 vdd.n3015 10.6151
R4616 vdd.n3017 vdd.n3016 10.6151
R4617 vdd.n3017 vdd.n826 10.6151
R4618 vdd.n3027 vdd.n826 10.6151
R4619 vdd.n3028 vdd.n3027 10.6151
R4620 vdd.n3029 vdd.n3028 10.6151
R4621 vdd.n3029 vdd.n812 10.6151
R4622 vdd.n3084 vdd.n812 10.6151
R4623 vdd.n3085 vdd.n3084 10.6151
R4624 vdd.n3086 vdd.n3085 10.6151
R4625 vdd.n3086 vdd.n779 10.6151
R4626 vdd.n3156 vdd.n779 10.6151
R4627 vdd.n3155 vdd.n3154 10.6151
R4628 vdd.n3154 vdd.n780 10.6151
R4629 vdd.n781 vdd.n780 10.6151
R4630 vdd.n3147 vdd.n781 10.6151
R4631 vdd.n3147 vdd.n3146 10.6151
R4632 vdd.n3146 vdd.n3145 10.6151
R4633 vdd.n3145 vdd.n783 10.6151
R4634 vdd.n3140 vdd.n783 10.6151
R4635 vdd.n3140 vdd.n3139 10.6151
R4636 vdd.n3139 vdd.n3138 10.6151
R4637 vdd.n3138 vdd.n786 10.6151
R4638 vdd.n3133 vdd.n786 10.6151
R4639 vdd.n3133 vdd.n3132 10.6151
R4640 vdd.n3132 vdd.n3131 10.6151
R4641 vdd.n3131 vdd.n789 10.6151
R4642 vdd.n3126 vdd.n789 10.6151
R4643 vdd.n3126 vdd.n3125 10.6151
R4644 vdd.n3125 vdd.n3123 10.6151
R4645 vdd.n3123 vdd.n792 10.6151
R4646 vdd.n3118 vdd.n792 10.6151
R4647 vdd.n3118 vdd.n3117 10.6151
R4648 vdd.n3117 vdd.n3116 10.6151
R4649 vdd.n3116 vdd.n795 10.6151
R4650 vdd.n3111 vdd.n795 10.6151
R4651 vdd.n3111 vdd.n3110 10.6151
R4652 vdd.n3110 vdd.n3109 10.6151
R4653 vdd.n3109 vdd.n798 10.6151
R4654 vdd.n3104 vdd.n798 10.6151
R4655 vdd.n3104 vdd.n3103 10.6151
R4656 vdd.n3103 vdd.n3102 10.6151
R4657 vdd.n3102 vdd.n801 10.6151
R4658 vdd.n3097 vdd.n3096 10.6151
R4659 vdd.n3096 vdd.n3095 10.6151
R4660 vdd.n3074 vdd.n3035 10.6151
R4661 vdd.n3069 vdd.n3035 10.6151
R4662 vdd.n3069 vdd.n3068 10.6151
R4663 vdd.n3068 vdd.n3067 10.6151
R4664 vdd.n3067 vdd.n3037 10.6151
R4665 vdd.n3062 vdd.n3037 10.6151
R4666 vdd.n3062 vdd.n3061 10.6151
R4667 vdd.n3061 vdd.n3060 10.6151
R4668 vdd.n3060 vdd.n3040 10.6151
R4669 vdd.n3055 vdd.n3040 10.6151
R4670 vdd.n3055 vdd.n3054 10.6151
R4671 vdd.n3054 vdd.n3053 10.6151
R4672 vdd.n3053 vdd.n3043 10.6151
R4673 vdd.n3048 vdd.n3043 10.6151
R4674 vdd.n3048 vdd.n3047 10.6151
R4675 vdd.n3047 vdd.n753 10.6151
R4676 vdd.n3191 vdd.n753 10.6151
R4677 vdd.n3191 vdd.n754 10.6151
R4678 vdd.n757 vdd.n754 10.6151
R4679 vdd.n3184 vdd.n757 10.6151
R4680 vdd.n3184 vdd.n3183 10.6151
R4681 vdd.n3183 vdd.n3182 10.6151
R4682 vdd.n3182 vdd.n759 10.6151
R4683 vdd.n3177 vdd.n759 10.6151
R4684 vdd.n3177 vdd.n3176 10.6151
R4685 vdd.n3176 vdd.n3175 10.6151
R4686 vdd.n3175 vdd.n762 10.6151
R4687 vdd.n3170 vdd.n762 10.6151
R4688 vdd.n3170 vdd.n3169 10.6151
R4689 vdd.n3169 vdd.n3168 10.6151
R4690 vdd.n3168 vdd.n765 10.6151
R4691 vdd.n3163 vdd.n3162 10.6151
R4692 vdd.n3162 vdd.n3161 10.6151
R4693 vdd.n2924 vdd.n2923 10.6151
R4694 vdd.n2923 vdd.n2921 10.6151
R4695 vdd.n2921 vdd.n2920 10.6151
R4696 vdd.n2920 vdd.n2746 10.6151
R4697 vdd.n2820 vdd.n2746 10.6151
R4698 vdd.n2821 vdd.n2820 10.6151
R4699 vdd.n2823 vdd.n2821 10.6151
R4700 vdd.n2824 vdd.n2823 10.6151
R4701 vdd.n2904 vdd.n2824 10.6151
R4702 vdd.n2904 vdd.n2903 10.6151
R4703 vdd.n2903 vdd.n2902 10.6151
R4704 vdd.n2902 vdd.n2900 10.6151
R4705 vdd.n2900 vdd.n2899 10.6151
R4706 vdd.n2899 vdd.n2897 10.6151
R4707 vdd.n2897 vdd.n2896 10.6151
R4708 vdd.n2896 vdd.n2856 10.6151
R4709 vdd.n2856 vdd.n2855 10.6151
R4710 vdd.n2855 vdd.n2853 10.6151
R4711 vdd.n2853 vdd.n2852 10.6151
R4712 vdd.n2852 vdd.n2850 10.6151
R4713 vdd.n2850 vdd.n2849 10.6151
R4714 vdd.n2849 vdd.n2847 10.6151
R4715 vdd.n2847 vdd.n2846 10.6151
R4716 vdd.n2846 vdd.n2844 10.6151
R4717 vdd.n2844 vdd.n2843 10.6151
R4718 vdd.n2843 vdd.n2841 10.6151
R4719 vdd.n2841 vdd.n2840 10.6151
R4720 vdd.n2840 vdd.n2838 10.6151
R4721 vdd.n2838 vdd.n2837 10.6151
R4722 vdd.n2837 vdd.n2835 10.6151
R4723 vdd.n2835 vdd.n2834 10.6151
R4724 vdd.n2834 vdd.n2832 10.6151
R4725 vdd.n2832 vdd.n2831 10.6151
R4726 vdd.n2831 vdd.n2829 10.6151
R4727 vdd.n2829 vdd.n2828 10.6151
R4728 vdd.n2828 vdd.n2826 10.6151
R4729 vdd.n2826 vdd.n2825 10.6151
R4730 vdd.n2825 vdd.n771 10.6151
R4731 vdd.n2681 vdd.n913 10.6151
R4732 vdd.n2684 vdd.n2681 10.6151
R4733 vdd.n2685 vdd.n2684 10.6151
R4734 vdd.n2688 vdd.n2685 10.6151
R4735 vdd.n2689 vdd.n2688 10.6151
R4736 vdd.n2692 vdd.n2689 10.6151
R4737 vdd.n2693 vdd.n2692 10.6151
R4738 vdd.n2696 vdd.n2693 10.6151
R4739 vdd.n2697 vdd.n2696 10.6151
R4740 vdd.n2700 vdd.n2697 10.6151
R4741 vdd.n2701 vdd.n2700 10.6151
R4742 vdd.n2704 vdd.n2701 10.6151
R4743 vdd.n2705 vdd.n2704 10.6151
R4744 vdd.n2708 vdd.n2705 10.6151
R4745 vdd.n2709 vdd.n2708 10.6151
R4746 vdd.n2712 vdd.n2709 10.6151
R4747 vdd.n2713 vdd.n2712 10.6151
R4748 vdd.n2716 vdd.n2713 10.6151
R4749 vdd.n2717 vdd.n2716 10.6151
R4750 vdd.n2720 vdd.n2717 10.6151
R4751 vdd.n2721 vdd.n2720 10.6151
R4752 vdd.n2724 vdd.n2721 10.6151
R4753 vdd.n2725 vdd.n2724 10.6151
R4754 vdd.n2728 vdd.n2725 10.6151
R4755 vdd.n2729 vdd.n2728 10.6151
R4756 vdd.n2732 vdd.n2729 10.6151
R4757 vdd.n2733 vdd.n2732 10.6151
R4758 vdd.n2736 vdd.n2733 10.6151
R4759 vdd.n2737 vdd.n2736 10.6151
R4760 vdd.n2740 vdd.n2737 10.6151
R4761 vdd.n2741 vdd.n2740 10.6151
R4762 vdd.n2745 vdd.n2744 10.6151
R4763 vdd.n2925 vdd.n2745 10.6151
R4764 vdd.n2937 vdd.n2936 10.6151
R4765 vdd.n2938 vdd.n2937 10.6151
R4766 vdd.n2938 vdd.n903 10.6151
R4767 vdd.n2948 vdd.n903 10.6151
R4768 vdd.n2949 vdd.n2948 10.6151
R4769 vdd.n2950 vdd.n2949 10.6151
R4770 vdd.n2950 vdd.n891 10.6151
R4771 vdd.n2960 vdd.n891 10.6151
R4772 vdd.n2961 vdd.n2960 10.6151
R4773 vdd.n2962 vdd.n2961 10.6151
R4774 vdd.n2962 vdd.n880 10.6151
R4775 vdd.n2972 vdd.n880 10.6151
R4776 vdd.n2973 vdd.n2972 10.6151
R4777 vdd.n2974 vdd.n2973 10.6151
R4778 vdd.n2974 vdd.n868 10.6151
R4779 vdd.n2984 vdd.n868 10.6151
R4780 vdd.n2985 vdd.n2984 10.6151
R4781 vdd.n2986 vdd.n2985 10.6151
R4782 vdd.n2986 vdd.n857 10.6151
R4783 vdd.n2996 vdd.n857 10.6151
R4784 vdd.n2999 vdd.n2998 10.6151
R4785 vdd.n2999 vdd.n843 10.6151
R4786 vdd.n3009 vdd.n843 10.6151
R4787 vdd.n3010 vdd.n3009 10.6151
R4788 vdd.n3011 vdd.n3010 10.6151
R4789 vdd.n3011 vdd.n831 10.6151
R4790 vdd.n3021 vdd.n831 10.6151
R4791 vdd.n3022 vdd.n3021 10.6151
R4792 vdd.n3023 vdd.n3022 10.6151
R4793 vdd.n3023 vdd.n820 10.6151
R4794 vdd.n3033 vdd.n820 10.6151
R4795 vdd.n3034 vdd.n3033 10.6151
R4796 vdd.n3080 vdd.n3034 10.6151
R4797 vdd.n3080 vdd.n3079 10.6151
R4798 vdd.n3079 vdd.n3078 10.6151
R4799 vdd.n3078 vdd.n3077 10.6151
R4800 vdd.n3077 vdd.n3075 10.6151
R4801 vdd.n2387 vdd.n2386 10.6151
R4802 vdd.n2388 vdd.n2387 10.6151
R4803 vdd.n2388 vdd.n1067 10.6151
R4804 vdd.n2398 vdd.n1067 10.6151
R4805 vdd.n2399 vdd.n2398 10.6151
R4806 vdd.n2400 vdd.n2399 10.6151
R4807 vdd.n2400 vdd.n1055 10.6151
R4808 vdd.n2410 vdd.n1055 10.6151
R4809 vdd.n2411 vdd.n2410 10.6151
R4810 vdd.n2412 vdd.n2411 10.6151
R4811 vdd.n2412 vdd.n1043 10.6151
R4812 vdd.n2422 vdd.n1043 10.6151
R4813 vdd.n2423 vdd.n2422 10.6151
R4814 vdd.n2424 vdd.n2423 10.6151
R4815 vdd.n2424 vdd.n1030 10.6151
R4816 vdd.n2434 vdd.n1030 10.6151
R4817 vdd.n2435 vdd.n2434 10.6151
R4818 vdd.n2437 vdd.n1018 10.6151
R4819 vdd.n2447 vdd.n1018 10.6151
R4820 vdd.n2448 vdd.n2447 10.6151
R4821 vdd.n2449 vdd.n2448 10.6151
R4822 vdd.n2449 vdd.n1006 10.6151
R4823 vdd.n2459 vdd.n1006 10.6151
R4824 vdd.n2460 vdd.n2459 10.6151
R4825 vdd.n2461 vdd.n2460 10.6151
R4826 vdd.n2461 vdd.n995 10.6151
R4827 vdd.n2471 vdd.n995 10.6151
R4828 vdd.n2472 vdd.n2471 10.6151
R4829 vdd.n2473 vdd.n2472 10.6151
R4830 vdd.n2473 vdd.n984 10.6151
R4831 vdd.n2483 vdd.n984 10.6151
R4832 vdd.n2484 vdd.n2483 10.6151
R4833 vdd.n2487 vdd.n2484 10.6151
R4834 vdd.n2487 vdd.n2486 10.6151
R4835 vdd.n2486 vdd.n2485 10.6151
R4836 vdd.n2485 vdd.n967 10.6151
R4837 vdd.n2569 vdd.n967 10.6151
R4838 vdd.n2568 vdd.n2567 10.6151
R4839 vdd.n2567 vdd.n2564 10.6151
R4840 vdd.n2564 vdd.n2563 10.6151
R4841 vdd.n2563 vdd.n2560 10.6151
R4842 vdd.n2560 vdd.n2559 10.6151
R4843 vdd.n2559 vdd.n2556 10.6151
R4844 vdd.n2556 vdd.n2555 10.6151
R4845 vdd.n2555 vdd.n2552 10.6151
R4846 vdd.n2552 vdd.n2551 10.6151
R4847 vdd.n2551 vdd.n2548 10.6151
R4848 vdd.n2548 vdd.n2547 10.6151
R4849 vdd.n2547 vdd.n2544 10.6151
R4850 vdd.n2544 vdd.n2543 10.6151
R4851 vdd.n2543 vdd.n2540 10.6151
R4852 vdd.n2540 vdd.n2539 10.6151
R4853 vdd.n2539 vdd.n2536 10.6151
R4854 vdd.n2536 vdd.n2535 10.6151
R4855 vdd.n2535 vdd.n2532 10.6151
R4856 vdd.n2532 vdd.n2531 10.6151
R4857 vdd.n2531 vdd.n2528 10.6151
R4858 vdd.n2528 vdd.n2527 10.6151
R4859 vdd.n2527 vdd.n2524 10.6151
R4860 vdd.n2524 vdd.n2523 10.6151
R4861 vdd.n2523 vdd.n2520 10.6151
R4862 vdd.n2520 vdd.n2519 10.6151
R4863 vdd.n2519 vdd.n2516 10.6151
R4864 vdd.n2516 vdd.n2515 10.6151
R4865 vdd.n2515 vdd.n2512 10.6151
R4866 vdd.n2512 vdd.n2511 10.6151
R4867 vdd.n2511 vdd.n2508 10.6151
R4868 vdd.n2508 vdd.n2507 10.6151
R4869 vdd.n2504 vdd.n2503 10.6151
R4870 vdd.n2503 vdd.n2501 10.6151
R4871 vdd.n2203 vdd.n2201 10.6151
R4872 vdd.n2204 vdd.n2203 10.6151
R4873 vdd.n2206 vdd.n2204 10.6151
R4874 vdd.n2207 vdd.n2206 10.6151
R4875 vdd.n2209 vdd.n2207 10.6151
R4876 vdd.n2210 vdd.n2209 10.6151
R4877 vdd.n2212 vdd.n2210 10.6151
R4878 vdd.n2213 vdd.n2212 10.6151
R4879 vdd.n2215 vdd.n2213 10.6151
R4880 vdd.n2216 vdd.n2215 10.6151
R4881 vdd.n2218 vdd.n2216 10.6151
R4882 vdd.n2219 vdd.n2218 10.6151
R4883 vdd.n2221 vdd.n2219 10.6151
R4884 vdd.n2222 vdd.n2221 10.6151
R4885 vdd.n2224 vdd.n2222 10.6151
R4886 vdd.n2225 vdd.n2224 10.6151
R4887 vdd.n2227 vdd.n2225 10.6151
R4888 vdd.n2228 vdd.n2227 10.6151
R4889 vdd.n2230 vdd.n2228 10.6151
R4890 vdd.n2231 vdd.n2230 10.6151
R4891 vdd.n2233 vdd.n2231 10.6151
R4892 vdd.n2234 vdd.n2233 10.6151
R4893 vdd.n2273 vdd.n2234 10.6151
R4894 vdd.n2273 vdd.n2272 10.6151
R4895 vdd.n2272 vdd.n2271 10.6151
R4896 vdd.n2271 vdd.n2269 10.6151
R4897 vdd.n2269 vdd.n2268 10.6151
R4898 vdd.n2268 vdd.n2266 10.6151
R4899 vdd.n2266 vdd.n2265 10.6151
R4900 vdd.n2265 vdd.n2242 10.6151
R4901 vdd.n2242 vdd.n2241 10.6151
R4902 vdd.n2241 vdd.n2239 10.6151
R4903 vdd.n2239 vdd.n2238 10.6151
R4904 vdd.n2238 vdd.n2236 10.6151
R4905 vdd.n2236 vdd.n2235 10.6151
R4906 vdd.n2235 vdd.n971 10.6151
R4907 vdd.n2499 vdd.n971 10.6151
R4908 vdd.n2500 vdd.n2499 10.6151
R4909 vdd.n2131 vdd.n1079 10.6151
R4910 vdd.n2136 vdd.n2131 10.6151
R4911 vdd.n2137 vdd.n2136 10.6151
R4912 vdd.n2138 vdd.n2137 10.6151
R4913 vdd.n2138 vdd.n2129 10.6151
R4914 vdd.n2144 vdd.n2129 10.6151
R4915 vdd.n2145 vdd.n2144 10.6151
R4916 vdd.n2146 vdd.n2145 10.6151
R4917 vdd.n2146 vdd.n2127 10.6151
R4918 vdd.n2152 vdd.n2127 10.6151
R4919 vdd.n2153 vdd.n2152 10.6151
R4920 vdd.n2154 vdd.n2153 10.6151
R4921 vdd.n2154 vdd.n2125 10.6151
R4922 vdd.n2160 vdd.n2125 10.6151
R4923 vdd.n2161 vdd.n2160 10.6151
R4924 vdd.n2162 vdd.n2161 10.6151
R4925 vdd.n2162 vdd.n2123 10.6151
R4926 vdd.n2168 vdd.n2123 10.6151
R4927 vdd.n2169 vdd.n2168 10.6151
R4928 vdd.n2170 vdd.n2169 10.6151
R4929 vdd.n2170 vdd.n1113 10.6151
R4930 vdd.n2176 vdd.n1113 10.6151
R4931 vdd.n2177 vdd.n2176 10.6151
R4932 vdd.n2178 vdd.n2177 10.6151
R4933 vdd.n2178 vdd.n1111 10.6151
R4934 vdd.n2184 vdd.n1111 10.6151
R4935 vdd.n2185 vdd.n2184 10.6151
R4936 vdd.n2186 vdd.n2185 10.6151
R4937 vdd.n2186 vdd.n1109 10.6151
R4938 vdd.n2192 vdd.n1109 10.6151
R4939 vdd.n2193 vdd.n2192 10.6151
R4940 vdd.n2195 vdd.n1105 10.6151
R4941 vdd.n2200 vdd.n1105 10.6151
R4942 vdd.t153 vdd.n1856 10.5435
R4943 vdd.n636 vdd.t151 10.5435
R4944 vdd.n304 vdd.n286 10.4732
R4945 vdd.n249 vdd.n231 10.4732
R4946 vdd.n206 vdd.n188 10.4732
R4947 vdd.n151 vdd.n133 10.4732
R4948 vdd.n109 vdd.n91 10.4732
R4949 vdd.n54 vdd.n36 10.4732
R4950 vdd.n1753 vdd.n1735 10.4732
R4951 vdd.n1808 vdd.n1790 10.4732
R4952 vdd.n1655 vdd.n1637 10.4732
R4953 vdd.n1710 vdd.n1692 10.4732
R4954 vdd.n1558 vdd.n1540 10.4732
R4955 vdd.n1613 vdd.n1595 10.4732
R4956 vdd.n1840 vdd.t212 10.3167
R4957 vdd.n3387 vdd.t149 10.3167
R4958 vdd.n2571 vdd.t260 10.2034
R4959 vdd.n2934 vdd.t116 10.2034
R4960 vdd.t165 vdd.n1184 10.09
R4961 vdd.n1892 vdd.t62 10.09
R4962 vdd.n3335 vdd.t36 10.09
R4963 vdd.n3468 vdd.t145 10.09
R4964 vdd.n2099 vdd.n1093 9.88581
R4965 vdd.n3125 vdd.n3124 9.88581
R4966 vdd.n3192 vdd.n3191 9.88581
R4967 vdd.n2123 vdd.n2122 9.88581
R4968 vdd.n1504 vdd.t188 9.86327
R4969 vdd.n3459 vdd.t134 9.86327
R4970 vdd.n303 vdd.n288 9.69747
R4971 vdd.n248 vdd.n233 9.69747
R4972 vdd.n205 vdd.n190 9.69747
R4973 vdd.n150 vdd.n135 9.69747
R4974 vdd.n108 vdd.n93 9.69747
R4975 vdd.n53 vdd.n38 9.69747
R4976 vdd.n1752 vdd.n1737 9.69747
R4977 vdd.n1807 vdd.n1792 9.69747
R4978 vdd.n1654 vdd.n1639 9.69747
R4979 vdd.n1709 vdd.n1694 9.69747
R4980 vdd.n1557 vdd.n1542 9.69747
R4981 vdd.n1612 vdd.n1597 9.69747
R4982 vdd.t176 vdd.n1478 9.63654
R4983 vdd.n3418 vdd.t147 9.63654
R4984 vdd.n319 vdd.n318 9.45567
R4985 vdd.n264 vdd.n263 9.45567
R4986 vdd.n221 vdd.n220 9.45567
R4987 vdd.n166 vdd.n165 9.45567
R4988 vdd.n124 vdd.n123 9.45567
R4989 vdd.n69 vdd.n68 9.45567
R4990 vdd.n1768 vdd.n1767 9.45567
R4991 vdd.n1823 vdd.n1822 9.45567
R4992 vdd.n1670 vdd.n1669 9.45567
R4993 vdd.n1725 vdd.n1724 9.45567
R4994 vdd.n1573 vdd.n1572 9.45567
R4995 vdd.n1628 vdd.n1627 9.45567
R4996 vdd.n2072 vdd.n1926 9.3005
R4997 vdd.n2071 vdd.n2070 9.3005
R4998 vdd.n1932 vdd.n1931 9.3005
R4999 vdd.n2065 vdd.n1936 9.3005
R5000 vdd.n2064 vdd.n1937 9.3005
R5001 vdd.n2063 vdd.n1938 9.3005
R5002 vdd.n1942 vdd.n1939 9.3005
R5003 vdd.n2058 vdd.n1943 9.3005
R5004 vdd.n2057 vdd.n1944 9.3005
R5005 vdd.n2056 vdd.n1945 9.3005
R5006 vdd.n1949 vdd.n1946 9.3005
R5007 vdd.n2051 vdd.n1950 9.3005
R5008 vdd.n2050 vdd.n1951 9.3005
R5009 vdd.n2049 vdd.n1952 9.3005
R5010 vdd.n1956 vdd.n1953 9.3005
R5011 vdd.n2044 vdd.n1957 9.3005
R5012 vdd.n2043 vdd.n1958 9.3005
R5013 vdd.n2042 vdd.n1959 9.3005
R5014 vdd.n1963 vdd.n1960 9.3005
R5015 vdd.n2037 vdd.n1964 9.3005
R5016 vdd.n2036 vdd.n1965 9.3005
R5017 vdd.n2035 vdd.n2034 9.3005
R5018 vdd.n2033 vdd.n1966 9.3005
R5019 vdd.n2032 vdd.n2031 9.3005
R5020 vdd.n1972 vdd.n1971 9.3005
R5021 vdd.n2026 vdd.n1976 9.3005
R5022 vdd.n2025 vdd.n1977 9.3005
R5023 vdd.n2024 vdd.n1978 9.3005
R5024 vdd.n1982 vdd.n1979 9.3005
R5025 vdd.n2019 vdd.n1983 9.3005
R5026 vdd.n2018 vdd.n1984 9.3005
R5027 vdd.n2017 vdd.n1985 9.3005
R5028 vdd.n1989 vdd.n1986 9.3005
R5029 vdd.n2012 vdd.n1990 9.3005
R5030 vdd.n2011 vdd.n1991 9.3005
R5031 vdd.n2010 vdd.n1992 9.3005
R5032 vdd.n1994 vdd.n1993 9.3005
R5033 vdd.n2005 vdd.n1115 9.3005
R5034 vdd.n2074 vdd.n2073 9.3005
R5035 vdd.n2098 vdd.n2097 9.3005
R5036 vdd.n1904 vdd.n1903 9.3005
R5037 vdd.n1909 vdd.n1907 9.3005
R5038 vdd.n2090 vdd.n1910 9.3005
R5039 vdd.n2089 vdd.n1911 9.3005
R5040 vdd.n2088 vdd.n1912 9.3005
R5041 vdd.n1916 vdd.n1913 9.3005
R5042 vdd.n2083 vdd.n1917 9.3005
R5043 vdd.n2082 vdd.n1918 9.3005
R5044 vdd.n2081 vdd.n1919 9.3005
R5045 vdd.n1923 vdd.n1920 9.3005
R5046 vdd.n2076 vdd.n1924 9.3005
R5047 vdd.n2075 vdd.n1925 9.3005
R5048 vdd.n2107 vdd.n1897 9.3005
R5049 vdd.n2109 vdd.n2108 9.3005
R5050 vdd.n1828 vdd.n1174 9.3005
R5051 vdd.n1830 vdd.n1829 9.3005
R5052 vdd.n1165 vdd.n1164 9.3005
R5053 vdd.n1843 vdd.n1842 9.3005
R5054 vdd.n1844 vdd.n1163 9.3005
R5055 vdd.n1846 vdd.n1845 9.3005
R5056 vdd.n1153 vdd.n1152 9.3005
R5057 vdd.n1860 vdd.n1859 9.3005
R5058 vdd.n1861 vdd.n1151 9.3005
R5059 vdd.n1863 vdd.n1862 9.3005
R5060 vdd.n1142 vdd.n1141 9.3005
R5061 vdd.n1877 vdd.n1876 9.3005
R5062 vdd.n1878 vdd.n1140 9.3005
R5063 vdd.n1880 vdd.n1879 9.3005
R5064 vdd.n1130 vdd.n1129 9.3005
R5065 vdd.n1895 vdd.n1894 9.3005
R5066 vdd.n1896 vdd.n1128 9.3005
R5067 vdd.n2111 vdd.n2110 9.3005
R5068 vdd.n295 vdd.n294 9.3005
R5069 vdd.n290 vdd.n289 9.3005
R5070 vdd.n301 vdd.n300 9.3005
R5071 vdd.n303 vdd.n302 9.3005
R5072 vdd.n286 vdd.n285 9.3005
R5073 vdd.n309 vdd.n308 9.3005
R5074 vdd.n311 vdd.n310 9.3005
R5075 vdd.n283 vdd.n280 9.3005
R5076 vdd.n318 vdd.n317 9.3005
R5077 vdd.n240 vdd.n239 9.3005
R5078 vdd.n235 vdd.n234 9.3005
R5079 vdd.n246 vdd.n245 9.3005
R5080 vdd.n248 vdd.n247 9.3005
R5081 vdd.n231 vdd.n230 9.3005
R5082 vdd.n254 vdd.n253 9.3005
R5083 vdd.n256 vdd.n255 9.3005
R5084 vdd.n228 vdd.n225 9.3005
R5085 vdd.n263 vdd.n262 9.3005
R5086 vdd.n197 vdd.n196 9.3005
R5087 vdd.n192 vdd.n191 9.3005
R5088 vdd.n203 vdd.n202 9.3005
R5089 vdd.n205 vdd.n204 9.3005
R5090 vdd.n188 vdd.n187 9.3005
R5091 vdd.n211 vdd.n210 9.3005
R5092 vdd.n213 vdd.n212 9.3005
R5093 vdd.n185 vdd.n182 9.3005
R5094 vdd.n220 vdd.n219 9.3005
R5095 vdd.n142 vdd.n141 9.3005
R5096 vdd.n137 vdd.n136 9.3005
R5097 vdd.n148 vdd.n147 9.3005
R5098 vdd.n150 vdd.n149 9.3005
R5099 vdd.n133 vdd.n132 9.3005
R5100 vdd.n156 vdd.n155 9.3005
R5101 vdd.n158 vdd.n157 9.3005
R5102 vdd.n130 vdd.n127 9.3005
R5103 vdd.n165 vdd.n164 9.3005
R5104 vdd.n100 vdd.n99 9.3005
R5105 vdd.n95 vdd.n94 9.3005
R5106 vdd.n106 vdd.n105 9.3005
R5107 vdd.n108 vdd.n107 9.3005
R5108 vdd.n91 vdd.n90 9.3005
R5109 vdd.n114 vdd.n113 9.3005
R5110 vdd.n116 vdd.n115 9.3005
R5111 vdd.n88 vdd.n85 9.3005
R5112 vdd.n123 vdd.n122 9.3005
R5113 vdd.n45 vdd.n44 9.3005
R5114 vdd.n40 vdd.n39 9.3005
R5115 vdd.n51 vdd.n50 9.3005
R5116 vdd.n53 vdd.n52 9.3005
R5117 vdd.n36 vdd.n35 9.3005
R5118 vdd.n59 vdd.n58 9.3005
R5119 vdd.n61 vdd.n60 9.3005
R5120 vdd.n33 vdd.n30 9.3005
R5121 vdd.n68 vdd.n67 9.3005
R5122 vdd.n3241 vdd.n3240 9.3005
R5123 vdd.n3242 vdd.n721 9.3005
R5124 vdd.n720 vdd.n718 9.3005
R5125 vdd.n3248 vdd.n717 9.3005
R5126 vdd.n3249 vdd.n716 9.3005
R5127 vdd.n3250 vdd.n715 9.3005
R5128 vdd.n714 vdd.n712 9.3005
R5129 vdd.n3256 vdd.n711 9.3005
R5130 vdd.n3257 vdd.n710 9.3005
R5131 vdd.n3258 vdd.n709 9.3005
R5132 vdd.n708 vdd.n706 9.3005
R5133 vdd.n3264 vdd.n705 9.3005
R5134 vdd.n3265 vdd.n704 9.3005
R5135 vdd.n3266 vdd.n703 9.3005
R5136 vdd.n702 vdd.n700 9.3005
R5137 vdd.n3272 vdd.n699 9.3005
R5138 vdd.n3273 vdd.n698 9.3005
R5139 vdd.n3274 vdd.n697 9.3005
R5140 vdd.n696 vdd.n694 9.3005
R5141 vdd.n3280 vdd.n693 9.3005
R5142 vdd.n3281 vdd.n692 9.3005
R5143 vdd.n3282 vdd.n691 9.3005
R5144 vdd.n690 vdd.n688 9.3005
R5145 vdd.n3288 vdd.n685 9.3005
R5146 vdd.n3289 vdd.n684 9.3005
R5147 vdd.n3290 vdd.n683 9.3005
R5148 vdd.n682 vdd.n680 9.3005
R5149 vdd.n3296 vdd.n679 9.3005
R5150 vdd.n3297 vdd.n678 9.3005
R5151 vdd.n3298 vdd.n677 9.3005
R5152 vdd.n676 vdd.n674 9.3005
R5153 vdd.n3304 vdd.n673 9.3005
R5154 vdd.n3305 vdd.n672 9.3005
R5155 vdd.n3306 vdd.n671 9.3005
R5156 vdd.n670 vdd.n668 9.3005
R5157 vdd.n3311 vdd.n667 9.3005
R5158 vdd.n3321 vdd.n661 9.3005
R5159 vdd.n3323 vdd.n3322 9.3005
R5160 vdd.n652 vdd.n651 9.3005
R5161 vdd.n3338 vdd.n3337 9.3005
R5162 vdd.n3339 vdd.n650 9.3005
R5163 vdd.n3341 vdd.n3340 9.3005
R5164 vdd.n640 vdd.n639 9.3005
R5165 vdd.n3354 vdd.n3353 9.3005
R5166 vdd.n3355 vdd.n638 9.3005
R5167 vdd.n3357 vdd.n3356 9.3005
R5168 vdd.n628 vdd.n627 9.3005
R5169 vdd.n3371 vdd.n3370 9.3005
R5170 vdd.n3372 vdd.n626 9.3005
R5171 vdd.n3374 vdd.n3373 9.3005
R5172 vdd.n617 vdd.n616 9.3005
R5173 vdd.n3390 vdd.n3389 9.3005
R5174 vdd.n3391 vdd.n615 9.3005
R5175 vdd.n3393 vdd.n3392 9.3005
R5176 vdd.n324 vdd.n322 9.3005
R5177 vdd.n3325 vdd.n3324 9.3005
R5178 vdd.n3472 vdd.n3471 9.3005
R5179 vdd.n325 vdd.n323 9.3005
R5180 vdd.n3465 vdd.n334 9.3005
R5181 vdd.n3464 vdd.n335 9.3005
R5182 vdd.n3463 vdd.n336 9.3005
R5183 vdd.n343 vdd.n337 9.3005
R5184 vdd.n3457 vdd.n344 9.3005
R5185 vdd.n3456 vdd.n345 9.3005
R5186 vdd.n3455 vdd.n346 9.3005
R5187 vdd.n354 vdd.n347 9.3005
R5188 vdd.n3449 vdd.n355 9.3005
R5189 vdd.n3448 vdd.n356 9.3005
R5190 vdd.n3447 vdd.n357 9.3005
R5191 vdd.n365 vdd.n358 9.3005
R5192 vdd.n3441 vdd.n366 9.3005
R5193 vdd.n3440 vdd.n367 9.3005
R5194 vdd.n3439 vdd.n368 9.3005
R5195 vdd.n443 vdd.n369 9.3005
R5196 vdd.n447 vdd.n442 9.3005
R5197 vdd.n451 vdd.n450 9.3005
R5198 vdd.n452 vdd.n441 9.3005
R5199 vdd.n456 vdd.n453 9.3005
R5200 vdd.n457 vdd.n440 9.3005
R5201 vdd.n461 vdd.n460 9.3005
R5202 vdd.n462 vdd.n439 9.3005
R5203 vdd.n466 vdd.n463 9.3005
R5204 vdd.n467 vdd.n438 9.3005
R5205 vdd.n471 vdd.n470 9.3005
R5206 vdd.n472 vdd.n437 9.3005
R5207 vdd.n476 vdd.n473 9.3005
R5208 vdd.n477 vdd.n436 9.3005
R5209 vdd.n481 vdd.n480 9.3005
R5210 vdd.n482 vdd.n435 9.3005
R5211 vdd.n486 vdd.n483 9.3005
R5212 vdd.n487 vdd.n434 9.3005
R5213 vdd.n491 vdd.n490 9.3005
R5214 vdd.n492 vdd.n433 9.3005
R5215 vdd.n496 vdd.n493 9.3005
R5216 vdd.n497 vdd.n430 9.3005
R5217 vdd.n501 vdd.n500 9.3005
R5218 vdd.n502 vdd.n429 9.3005
R5219 vdd.n506 vdd.n503 9.3005
R5220 vdd.n507 vdd.n428 9.3005
R5221 vdd.n511 vdd.n510 9.3005
R5222 vdd.n512 vdd.n427 9.3005
R5223 vdd.n516 vdd.n513 9.3005
R5224 vdd.n517 vdd.n426 9.3005
R5225 vdd.n521 vdd.n520 9.3005
R5226 vdd.n522 vdd.n425 9.3005
R5227 vdd.n526 vdd.n523 9.3005
R5228 vdd.n527 vdd.n424 9.3005
R5229 vdd.n531 vdd.n530 9.3005
R5230 vdd.n532 vdd.n423 9.3005
R5231 vdd.n536 vdd.n533 9.3005
R5232 vdd.n537 vdd.n422 9.3005
R5233 vdd.n541 vdd.n540 9.3005
R5234 vdd.n542 vdd.n421 9.3005
R5235 vdd.n546 vdd.n543 9.3005
R5236 vdd.n547 vdd.n418 9.3005
R5237 vdd.n551 vdd.n550 9.3005
R5238 vdd.n552 vdd.n417 9.3005
R5239 vdd.n556 vdd.n553 9.3005
R5240 vdd.n557 vdd.n416 9.3005
R5241 vdd.n561 vdd.n560 9.3005
R5242 vdd.n562 vdd.n415 9.3005
R5243 vdd.n566 vdd.n563 9.3005
R5244 vdd.n567 vdd.n414 9.3005
R5245 vdd.n571 vdd.n570 9.3005
R5246 vdd.n572 vdd.n413 9.3005
R5247 vdd.n576 vdd.n573 9.3005
R5248 vdd.n577 vdd.n412 9.3005
R5249 vdd.n581 vdd.n580 9.3005
R5250 vdd.n582 vdd.n411 9.3005
R5251 vdd.n586 vdd.n583 9.3005
R5252 vdd.n587 vdd.n410 9.3005
R5253 vdd.n591 vdd.n590 9.3005
R5254 vdd.n592 vdd.n409 9.3005
R5255 vdd.n596 vdd.n593 9.3005
R5256 vdd.n598 vdd.n408 9.3005
R5257 vdd.n600 vdd.n599 9.3005
R5258 vdd.n3432 vdd.n3431 9.3005
R5259 vdd.n446 vdd.n444 9.3005
R5260 vdd.n3331 vdd.n655 9.3005
R5261 vdd.n3333 vdd.n3332 9.3005
R5262 vdd.n646 vdd.n645 9.3005
R5263 vdd.n3346 vdd.n3345 9.3005
R5264 vdd.n3347 vdd.n644 9.3005
R5265 vdd.n3349 vdd.n3348 9.3005
R5266 vdd.n633 vdd.n632 9.3005
R5267 vdd.n3362 vdd.n3361 9.3005
R5268 vdd.n3363 vdd.n631 9.3005
R5269 vdd.n3365 vdd.n3364 9.3005
R5270 vdd.n622 vdd.n621 9.3005
R5271 vdd.n3379 vdd.n3378 9.3005
R5272 vdd.n3380 vdd.n620 9.3005
R5273 vdd.n3385 vdd.n3381 9.3005
R5274 vdd.n3384 vdd.n3383 9.3005
R5275 vdd.n3382 vdd.n610 9.3005
R5276 vdd.n3398 vdd.n611 9.3005
R5277 vdd.n3399 vdd.n609 9.3005
R5278 vdd.n3401 vdd.n3400 9.3005
R5279 vdd.n3402 vdd.n608 9.3005
R5280 vdd.n3405 vdd.n3403 9.3005
R5281 vdd.n3406 vdd.n607 9.3005
R5282 vdd.n3408 vdd.n3407 9.3005
R5283 vdd.n3409 vdd.n606 9.3005
R5284 vdd.n3412 vdd.n3410 9.3005
R5285 vdd.n3413 vdd.n605 9.3005
R5286 vdd.n3415 vdd.n3414 9.3005
R5287 vdd.n3416 vdd.n604 9.3005
R5288 vdd.n3420 vdd.n3417 9.3005
R5289 vdd.n3421 vdd.n603 9.3005
R5290 vdd.n3423 vdd.n3422 9.3005
R5291 vdd.n3424 vdd.n602 9.3005
R5292 vdd.n3427 vdd.n3425 9.3005
R5293 vdd.n3428 vdd.n601 9.3005
R5294 vdd.n3430 vdd.n3429 9.3005
R5295 vdd.n3330 vdd.n3329 9.3005
R5296 vdd.n3194 vdd.n656 9.3005
R5297 vdd.n3199 vdd.n3193 9.3005
R5298 vdd.n3209 vdd.n748 9.3005
R5299 vdd.n3210 vdd.n747 9.3005
R5300 vdd.n746 vdd.n744 9.3005
R5301 vdd.n3216 vdd.n743 9.3005
R5302 vdd.n3217 vdd.n742 9.3005
R5303 vdd.n3218 vdd.n741 9.3005
R5304 vdd.n740 vdd.n738 9.3005
R5305 vdd.n3224 vdd.n737 9.3005
R5306 vdd.n3225 vdd.n736 9.3005
R5307 vdd.n3226 vdd.n735 9.3005
R5308 vdd.n734 vdd.n732 9.3005
R5309 vdd.n3231 vdd.n731 9.3005
R5310 vdd.n3232 vdd.n730 9.3005
R5311 vdd.n726 vdd.n725 9.3005
R5312 vdd.n3238 vdd.n3237 9.3005
R5313 vdd.n3239 vdd.n722 9.3005
R5314 vdd.n2121 vdd.n2120 9.3005
R5315 vdd.n2116 vdd.n1118 9.3005
R5316 vdd.n1460 vdd.n1459 9.3005
R5317 vdd.n1216 vdd.n1215 9.3005
R5318 vdd.n1473 vdd.n1472 9.3005
R5319 vdd.n1474 vdd.n1214 9.3005
R5320 vdd.n1476 vdd.n1475 9.3005
R5321 vdd.n1204 vdd.n1203 9.3005
R5322 vdd.n1490 vdd.n1489 9.3005
R5323 vdd.n1491 vdd.n1202 9.3005
R5324 vdd.n1493 vdd.n1492 9.3005
R5325 vdd.n1194 vdd.n1193 9.3005
R5326 vdd.n1507 vdd.n1506 9.3005
R5327 vdd.n1508 vdd.n1192 9.3005
R5328 vdd.n1510 vdd.n1509 9.3005
R5329 vdd.n1181 vdd.n1180 9.3005
R5330 vdd.n1523 vdd.n1522 9.3005
R5331 vdd.n1524 vdd.n1179 9.3005
R5332 vdd.n1526 vdd.n1525 9.3005
R5333 vdd.n1170 vdd.n1169 9.3005
R5334 vdd.n1835 vdd.n1834 9.3005
R5335 vdd.n1836 vdd.n1168 9.3005
R5336 vdd.n1838 vdd.n1837 9.3005
R5337 vdd.n1159 vdd.n1158 9.3005
R5338 vdd.n1851 vdd.n1850 9.3005
R5339 vdd.n1852 vdd.n1157 9.3005
R5340 vdd.n1854 vdd.n1853 9.3005
R5341 vdd.n1147 vdd.n1146 9.3005
R5342 vdd.n1868 vdd.n1867 9.3005
R5343 vdd.n1869 vdd.n1145 9.3005
R5344 vdd.n1871 vdd.n1870 9.3005
R5345 vdd.n1137 vdd.n1136 9.3005
R5346 vdd.n1885 vdd.n1884 9.3005
R5347 vdd.n1886 vdd.n1134 9.3005
R5348 vdd.n1890 vdd.n1889 9.3005
R5349 vdd.n1888 vdd.n1135 9.3005
R5350 vdd.n1887 vdd.n1123 9.3005
R5351 vdd.n1458 vdd.n1226 9.3005
R5352 vdd.n1351 vdd.n1227 9.3005
R5353 vdd.n1353 vdd.n1352 9.3005
R5354 vdd.n1354 vdd.n1346 9.3005
R5355 vdd.n1356 vdd.n1355 9.3005
R5356 vdd.n1357 vdd.n1345 9.3005
R5357 vdd.n1359 vdd.n1358 9.3005
R5358 vdd.n1360 vdd.n1340 9.3005
R5359 vdd.n1362 vdd.n1361 9.3005
R5360 vdd.n1363 vdd.n1339 9.3005
R5361 vdd.n1365 vdd.n1364 9.3005
R5362 vdd.n1366 vdd.n1334 9.3005
R5363 vdd.n1368 vdd.n1367 9.3005
R5364 vdd.n1369 vdd.n1333 9.3005
R5365 vdd.n1371 vdd.n1370 9.3005
R5366 vdd.n1372 vdd.n1328 9.3005
R5367 vdd.n1374 vdd.n1373 9.3005
R5368 vdd.n1375 vdd.n1327 9.3005
R5369 vdd.n1377 vdd.n1376 9.3005
R5370 vdd.n1378 vdd.n1322 9.3005
R5371 vdd.n1380 vdd.n1379 9.3005
R5372 vdd.n1381 vdd.n1321 9.3005
R5373 vdd.n1386 vdd.n1382 9.3005
R5374 vdd.n1387 vdd.n1317 9.3005
R5375 vdd.n1389 vdd.n1388 9.3005
R5376 vdd.n1390 vdd.n1316 9.3005
R5377 vdd.n1392 vdd.n1391 9.3005
R5378 vdd.n1393 vdd.n1311 9.3005
R5379 vdd.n1395 vdd.n1394 9.3005
R5380 vdd.n1396 vdd.n1310 9.3005
R5381 vdd.n1398 vdd.n1397 9.3005
R5382 vdd.n1399 vdd.n1305 9.3005
R5383 vdd.n1401 vdd.n1400 9.3005
R5384 vdd.n1402 vdd.n1304 9.3005
R5385 vdd.n1404 vdd.n1403 9.3005
R5386 vdd.n1405 vdd.n1299 9.3005
R5387 vdd.n1407 vdd.n1406 9.3005
R5388 vdd.n1408 vdd.n1298 9.3005
R5389 vdd.n1410 vdd.n1409 9.3005
R5390 vdd.n1411 vdd.n1293 9.3005
R5391 vdd.n1413 vdd.n1412 9.3005
R5392 vdd.n1414 vdd.n1292 9.3005
R5393 vdd.n1416 vdd.n1415 9.3005
R5394 vdd.n1417 vdd.n1289 9.3005
R5395 vdd.n1423 vdd.n1422 9.3005
R5396 vdd.n1424 vdd.n1288 9.3005
R5397 vdd.n1426 vdd.n1425 9.3005
R5398 vdd.n1427 vdd.n1283 9.3005
R5399 vdd.n1429 vdd.n1428 9.3005
R5400 vdd.n1430 vdd.n1282 9.3005
R5401 vdd.n1432 vdd.n1431 9.3005
R5402 vdd.n1433 vdd.n1277 9.3005
R5403 vdd.n1435 vdd.n1434 9.3005
R5404 vdd.n1436 vdd.n1276 9.3005
R5405 vdd.n1438 vdd.n1437 9.3005
R5406 vdd.n1439 vdd.n1271 9.3005
R5407 vdd.n1441 vdd.n1440 9.3005
R5408 vdd.n1442 vdd.n1270 9.3005
R5409 vdd.n1444 vdd.n1443 9.3005
R5410 vdd.n1445 vdd.n1266 9.3005
R5411 vdd.n1447 vdd.n1446 9.3005
R5412 vdd.n1448 vdd.n1265 9.3005
R5413 vdd.n1450 vdd.n1449 9.3005
R5414 vdd.n1451 vdd.n1264 9.3005
R5415 vdd.n1457 vdd.n1456 9.3005
R5416 vdd.n1465 vdd.n1464 9.3005
R5417 vdd.n1466 vdd.n1220 9.3005
R5418 vdd.n1468 vdd.n1467 9.3005
R5419 vdd.n1210 vdd.n1209 9.3005
R5420 vdd.n1482 vdd.n1481 9.3005
R5421 vdd.n1483 vdd.n1208 9.3005
R5422 vdd.n1485 vdd.n1484 9.3005
R5423 vdd.n1199 vdd.n1198 9.3005
R5424 vdd.n1499 vdd.n1498 9.3005
R5425 vdd.n1500 vdd.n1197 9.3005
R5426 vdd.n1502 vdd.n1501 9.3005
R5427 vdd.n1188 vdd.n1187 9.3005
R5428 vdd.n1515 vdd.n1514 9.3005
R5429 vdd.n1516 vdd.n1186 9.3005
R5430 vdd.n1518 vdd.n1517 9.3005
R5431 vdd.n1176 vdd.n1175 9.3005
R5432 vdd.n1532 vdd.n1531 9.3005
R5433 vdd.n1222 vdd.n1221 9.3005
R5434 vdd.n1744 vdd.n1743 9.3005
R5435 vdd.n1739 vdd.n1738 9.3005
R5436 vdd.n1750 vdd.n1749 9.3005
R5437 vdd.n1752 vdd.n1751 9.3005
R5438 vdd.n1735 vdd.n1734 9.3005
R5439 vdd.n1758 vdd.n1757 9.3005
R5440 vdd.n1760 vdd.n1759 9.3005
R5441 vdd.n1732 vdd.n1729 9.3005
R5442 vdd.n1767 vdd.n1766 9.3005
R5443 vdd.n1799 vdd.n1798 9.3005
R5444 vdd.n1794 vdd.n1793 9.3005
R5445 vdd.n1805 vdd.n1804 9.3005
R5446 vdd.n1807 vdd.n1806 9.3005
R5447 vdd.n1790 vdd.n1789 9.3005
R5448 vdd.n1813 vdd.n1812 9.3005
R5449 vdd.n1815 vdd.n1814 9.3005
R5450 vdd.n1787 vdd.n1784 9.3005
R5451 vdd.n1822 vdd.n1821 9.3005
R5452 vdd.n1646 vdd.n1645 9.3005
R5453 vdd.n1641 vdd.n1640 9.3005
R5454 vdd.n1652 vdd.n1651 9.3005
R5455 vdd.n1654 vdd.n1653 9.3005
R5456 vdd.n1637 vdd.n1636 9.3005
R5457 vdd.n1660 vdd.n1659 9.3005
R5458 vdd.n1662 vdd.n1661 9.3005
R5459 vdd.n1634 vdd.n1631 9.3005
R5460 vdd.n1669 vdd.n1668 9.3005
R5461 vdd.n1701 vdd.n1700 9.3005
R5462 vdd.n1696 vdd.n1695 9.3005
R5463 vdd.n1707 vdd.n1706 9.3005
R5464 vdd.n1709 vdd.n1708 9.3005
R5465 vdd.n1692 vdd.n1691 9.3005
R5466 vdd.n1715 vdd.n1714 9.3005
R5467 vdd.n1717 vdd.n1716 9.3005
R5468 vdd.n1689 vdd.n1686 9.3005
R5469 vdd.n1724 vdd.n1723 9.3005
R5470 vdd.n1549 vdd.n1548 9.3005
R5471 vdd.n1544 vdd.n1543 9.3005
R5472 vdd.n1555 vdd.n1554 9.3005
R5473 vdd.n1557 vdd.n1556 9.3005
R5474 vdd.n1540 vdd.n1539 9.3005
R5475 vdd.n1563 vdd.n1562 9.3005
R5476 vdd.n1565 vdd.n1564 9.3005
R5477 vdd.n1537 vdd.n1534 9.3005
R5478 vdd.n1572 vdd.n1571 9.3005
R5479 vdd.n1604 vdd.n1603 9.3005
R5480 vdd.n1599 vdd.n1598 9.3005
R5481 vdd.n1610 vdd.n1609 9.3005
R5482 vdd.n1612 vdd.n1611 9.3005
R5483 vdd.n1595 vdd.n1594 9.3005
R5484 vdd.n1618 vdd.n1617 9.3005
R5485 vdd.n1620 vdd.n1619 9.3005
R5486 vdd.n1592 vdd.n1589 9.3005
R5487 vdd.n1627 vdd.n1626 9.3005
R5488 vdd.n1478 vdd.t130 9.18308
R5489 vdd.n3418 vdd.t227 9.18308
R5490 vdd.n1504 vdd.t136 8.95635
R5491 vdd.t191 vdd.n3459 8.95635
R5492 vdd.n300 vdd.n299 8.92171
R5493 vdd.n245 vdd.n244 8.92171
R5494 vdd.n202 vdd.n201 8.92171
R5495 vdd.n147 vdd.n146 8.92171
R5496 vdd.n105 vdd.n104 8.92171
R5497 vdd.n50 vdd.n49 8.92171
R5498 vdd.n1749 vdd.n1748 8.92171
R5499 vdd.n1804 vdd.n1803 8.92171
R5500 vdd.n1651 vdd.n1650 8.92171
R5501 vdd.n1706 vdd.n1705 8.92171
R5502 vdd.n1554 vdd.n1553 8.92171
R5503 vdd.n1609 vdd.n1608 8.92171
R5504 vdd.n223 vdd.n125 8.81535
R5505 vdd.n1727 vdd.n1629 8.81535
R5506 vdd.n1184 vdd.t160 8.72962
R5507 vdd.t223 vdd.n3468 8.72962
R5508 vdd.n1840 vdd.t210 8.50289
R5509 vdd.n3387 vdd.t174 8.50289
R5510 vdd.n28 vdd.n14 8.42249
R5511 vdd.n1856 vdd.t186 8.27616
R5512 vdd.t171 vdd.n636 8.27616
R5513 vdd.n3474 vdd.n3473 8.16225
R5514 vdd.n1827 vdd.n1826 8.16225
R5515 vdd.n296 vdd.n290 8.14595
R5516 vdd.n241 vdd.n235 8.14595
R5517 vdd.n198 vdd.n192 8.14595
R5518 vdd.n143 vdd.n137 8.14595
R5519 vdd.n101 vdd.n95 8.14595
R5520 vdd.n46 vdd.n40 8.14595
R5521 vdd.n1745 vdd.n1739 8.14595
R5522 vdd.n1800 vdd.n1794 8.14595
R5523 vdd.n1647 vdd.n1641 8.14595
R5524 vdd.n1702 vdd.n1696 8.14595
R5525 vdd.n1550 vdd.n1544 8.14595
R5526 vdd.n1605 vdd.n1599 8.14595
R5527 vdd.t69 vdd.n1218 7.8227
R5528 vdd.t51 vdd.n363 7.8227
R5529 vdd.n2384 vdd.n1075 7.70933
R5530 vdd.n2390 vdd.n1075 7.70933
R5531 vdd.n2396 vdd.n1069 7.70933
R5532 vdd.n2396 vdd.n1063 7.70933
R5533 vdd.n2402 vdd.n1063 7.70933
R5534 vdd.n2402 vdd.n1057 7.70933
R5535 vdd.n2408 vdd.n1057 7.70933
R5536 vdd.n2414 vdd.n1051 7.70933
R5537 vdd.n2420 vdd.n1045 7.70933
R5538 vdd.n2426 vdd.n1038 7.70933
R5539 vdd.n2426 vdd.n1041 7.70933
R5540 vdd.n2432 vdd.n1034 7.70933
R5541 vdd.n2439 vdd.n1020 7.70933
R5542 vdd.n2445 vdd.n1020 7.70933
R5543 vdd.n2451 vdd.n1014 7.70933
R5544 vdd.n2457 vdd.n1010 7.70933
R5545 vdd.n2463 vdd.n1004 7.70933
R5546 vdd.n2481 vdd.n986 7.70933
R5547 vdd.n2481 vdd.n979 7.70933
R5548 vdd.n2489 vdd.n979 7.70933
R5549 vdd.n2571 vdd.n963 7.70933
R5550 vdd.n2934 vdd.n917 7.70933
R5551 vdd.n2946 vdd.n898 7.70933
R5552 vdd.n2952 vdd.n898 7.70933
R5553 vdd.n2952 vdd.n901 7.70933
R5554 vdd.n2970 vdd.n882 7.70933
R5555 vdd.n2976 vdd.n876 7.70933
R5556 vdd.n2982 vdd.n872 7.70933
R5557 vdd.n2988 vdd.n859 7.70933
R5558 vdd.n2994 vdd.n859 7.70933
R5559 vdd.n3001 vdd.n852 7.70933
R5560 vdd.n3007 vdd.n845 7.70933
R5561 vdd.n3007 vdd.n848 7.70933
R5562 vdd.n3013 vdd.n841 7.70933
R5563 vdd.n3019 vdd.n835 7.70933
R5564 vdd.n3025 vdd.n822 7.70933
R5565 vdd.n3031 vdd.n822 7.70933
R5566 vdd.n3031 vdd.n814 7.70933
R5567 vdd.n3082 vdd.n814 7.70933
R5568 vdd.n3082 vdd.n817 7.70933
R5569 vdd.n3088 vdd.n774 7.70933
R5570 vdd.n3158 vdd.n774 7.70933
R5571 vdd.t20 vdd.n1051 7.59597
R5572 vdd.n2263 vdd.t4 7.59597
R5573 vdd.n2906 vdd.t18 7.59597
R5574 vdd.n835 vdd.t28 7.59597
R5575 vdd.n295 vdd.n292 7.3702
R5576 vdd.n240 vdd.n237 7.3702
R5577 vdd.n197 vdd.n194 7.3702
R5578 vdd.n142 vdd.n139 7.3702
R5579 vdd.n100 vdd.n97 7.3702
R5580 vdd.n45 vdd.n42 7.3702
R5581 vdd.n1744 vdd.n1741 7.3702
R5582 vdd.n1799 vdd.n1796 7.3702
R5583 vdd.n1646 vdd.n1643 7.3702
R5584 vdd.n1701 vdd.n1698 7.3702
R5585 vdd.n1549 vdd.n1546 7.3702
R5586 vdd.n1604 vdd.n1601 7.3702
R5587 vdd.n1387 vdd.n1386 6.98232
R5588 vdd.n2036 vdd.n2035 6.98232
R5589 vdd.n547 vdd.n546 6.98232
R5590 vdd.n3242 vdd.n3241 6.98232
R5591 vdd.n1874 vdd.t142 6.91577
R5592 vdd.n2420 vdd.t19 6.91577
R5593 vdd.n3013 vdd.t3 6.91577
R5594 vdd.n3351 vdd.t138 6.91577
R5595 vdd.n2998 vdd.n2997 6.86879
R5596 vdd.n2436 vdd.n2435 6.86879
R5597 vdd.n2496 vdd.t258 6.80241
R5598 vdd.n2940 vdd.t114 6.80241
R5599 vdd.t167 vdd.n1155 6.68904
R5600 vdd.n3367 vdd.t203 6.68904
R5601 vdd.n1832 vdd.t140 6.46231
R5602 vdd.n3395 vdd.t155 6.46231
R5603 vdd.n2263 vdd.t262 6.34895
R5604 vdd.n2906 vdd.t264 6.34895
R5605 vdd.n3474 vdd.n321 6.32949
R5606 vdd.n1826 vdd.n1825 6.32949
R5607 vdd.t132 vdd.n1183 6.23558
R5608 vdd.t201 vdd.n332 6.23558
R5609 vdd.n1496 vdd.t208 6.00885
R5610 vdd.t30 vdd.n1014 6.00885
R5611 vdd.n872 vdd.t113 6.00885
R5612 vdd.n3453 vdd.t180 6.00885
R5613 vdd.n296 vdd.n295 5.81868
R5614 vdd.n241 vdd.n240 5.81868
R5615 vdd.n198 vdd.n197 5.81868
R5616 vdd.n143 vdd.n142 5.81868
R5617 vdd.n101 vdd.n100 5.81868
R5618 vdd.n46 vdd.n45 5.81868
R5619 vdd.n1745 vdd.n1744 5.81868
R5620 vdd.n1800 vdd.n1799 5.81868
R5621 vdd.n1647 vdd.n1646 5.81868
R5622 vdd.n1702 vdd.n1701 5.81868
R5623 vdd.n1550 vdd.n1549 5.81868
R5624 vdd.n1605 vdd.n1604 5.81868
R5625 vdd.n2579 vdd.n2578 5.77611
R5626 vdd.n2319 vdd.n2318 5.77611
R5627 vdd.n2808 vdd.n2807 5.77611
R5628 vdd.n3097 vdd.n806 5.77611
R5629 vdd.n3163 vdd.n770 5.77611
R5630 vdd.n2744 vdd.n2680 5.77611
R5631 vdd.n2504 vdd.n970 5.77611
R5632 vdd.n2195 vdd.n2194 5.77611
R5633 vdd.n1456 vdd.n1230 5.62474
R5634 vdd.n2119 vdd.n2116 5.62474
R5635 vdd.n3432 vdd.n407 5.62474
R5636 vdd.n3197 vdd.n3194 5.62474
R5637 vdd.n2457 vdd.t266 5.44203
R5638 vdd.n2976 vdd.t16 5.44203
R5639 vdd.n1206 vdd.t208 5.32866
R5640 vdd.t180 vdd.n3452 5.32866
R5641 vdd.n1512 vdd.t132 5.10193
R5642 vdd.n2432 vdd.t27 5.10193
R5643 vdd.n2451 vdd.t23 5.10193
R5644 vdd.n2982 vdd.t118 5.10193
R5645 vdd.n3001 vdd.t0 5.10193
R5646 vdd.n3461 vdd.t201 5.10193
R5647 vdd.n299 vdd.n290 5.04292
R5648 vdd.n244 vdd.n235 5.04292
R5649 vdd.n201 vdd.n192 5.04292
R5650 vdd.n146 vdd.n137 5.04292
R5651 vdd.n104 vdd.n95 5.04292
R5652 vdd.n49 vdd.n40 5.04292
R5653 vdd.n1748 vdd.n1739 5.04292
R5654 vdd.n1803 vdd.n1794 5.04292
R5655 vdd.n1650 vdd.n1641 5.04292
R5656 vdd.n1705 vdd.n1696 5.04292
R5657 vdd.n1553 vdd.n1544 5.04292
R5658 vdd.n1608 vdd.n1599 5.04292
R5659 vdd.n1034 vdd.t96 4.98857
R5660 vdd.t55 vdd.n852 4.98857
R5661 vdd.n1528 vdd.t140 4.8752
R5662 vdd.t44 vdd.n1069 4.8752
R5663 vdd.t8 vdd.t270 4.8752
R5664 vdd.n2251 vdd.t82 4.8752
R5665 vdd.n2918 vdd.t86 4.8752
R5666 vdd.t21 vdd.t29 4.8752
R5667 vdd.n817 vdd.t40 4.8752
R5668 vdd.t155 vdd.n328 4.8752
R5669 vdd.n2580 vdd.n2579 4.83952
R5670 vdd.n2320 vdd.n2319 4.83952
R5671 vdd.n2807 vdd.n2806 4.83952
R5672 vdd.n806 vdd.n801 4.83952
R5673 vdd.n770 vdd.n765 4.83952
R5674 vdd.n2741 vdd.n2680 4.83952
R5675 vdd.n2507 vdd.n970 4.83952
R5676 vdd.n2194 vdd.n2193 4.83952
R5677 vdd.n2475 vdd.t5 4.76184
R5678 vdd.n2958 vdd.t268 4.76184
R5679 vdd.n2004 vdd.n1116 4.74817
R5680 vdd.n1999 vdd.n1117 4.74817
R5681 vdd.n1901 vdd.n1898 4.74817
R5682 vdd.n2100 vdd.n1902 4.74817
R5683 vdd.n2102 vdd.n1901 4.74817
R5684 vdd.n2101 vdd.n2100 4.74817
R5685 vdd.n664 vdd.n662 4.74817
R5686 vdd.n3312 vdd.n665 4.74817
R5687 vdd.n3315 vdd.n665 4.74817
R5688 vdd.n3316 vdd.n664 4.74817
R5689 vdd.n3204 vdd.n749 4.74817
R5690 vdd.n3200 vdd.n751 4.74817
R5691 vdd.n3203 vdd.n751 4.74817
R5692 vdd.n3208 vdd.n749 4.74817
R5693 vdd.n2000 vdd.n1116 4.74817
R5694 vdd.n1119 vdd.n1117 4.74817
R5695 vdd.n321 vdd.n320 4.7074
R5696 vdd.n223 vdd.n222 4.7074
R5697 vdd.n1825 vdd.n1824 4.7074
R5698 vdd.n1727 vdd.n1726 4.7074
R5699 vdd.n1848 vdd.t167 4.64847
R5700 vdd.n3376 vdd.t203 4.64847
R5701 vdd.n1149 vdd.t142 4.42174
R5702 vdd.t138 vdd.n635 4.42174
R5703 vdd.n2251 vdd.t14 4.30838
R5704 vdd.n2918 vdd.t1 4.30838
R5705 vdd.n300 vdd.n288 4.26717
R5706 vdd.n245 vdd.n233 4.26717
R5707 vdd.n202 vdd.n190 4.26717
R5708 vdd.n147 vdd.n135 4.26717
R5709 vdd.n105 vdd.n93 4.26717
R5710 vdd.n50 vdd.n38 4.26717
R5711 vdd.n1749 vdd.n1737 4.26717
R5712 vdd.n1804 vdd.n1792 4.26717
R5713 vdd.n1651 vdd.n1639 4.26717
R5714 vdd.n1706 vdd.n1694 4.26717
R5715 vdd.n1554 vdd.n1542 4.26717
R5716 vdd.n1609 vdd.n1597 4.26717
R5717 vdd.t34 vdd.n1045 4.19501
R5718 vdd.n1004 vdd.t26 4.19501
R5719 vdd.t9 vdd.n882 4.19501
R5720 vdd.n841 vdd.t7 4.19501
R5721 vdd.n321 vdd.n223 4.10845
R5722 vdd.n1825 vdd.n1727 4.10845
R5723 vdd.n277 vdd.t198 4.06363
R5724 vdd.n277 vdd.t240 4.06363
R5725 vdd.n275 vdd.t241 4.06363
R5726 vdd.n275 vdd.t135 4.06363
R5727 vdd.n273 vdd.t164 4.06363
R5728 vdd.n273 vdd.t217 4.06363
R5729 vdd.n271 vdd.t233 4.06363
R5730 vdd.n271 vdd.t250 4.06363
R5731 vdd.n269 vdd.t253 4.06363
R5732 vdd.n269 vdd.t169 4.06363
R5733 vdd.n267 vdd.t196 4.06363
R5734 vdd.n267 vdd.t252 4.06363
R5735 vdd.n265 vdd.t254 4.06363
R5736 vdd.n265 vdd.t195 4.06363
R5737 vdd.n179 vdd.t181 4.06363
R5738 vdd.n179 vdd.t228 4.06363
R5739 vdd.n177 vdd.t229 4.06363
R5740 vdd.n177 vdd.t251 4.06363
R5741 vdd.n175 vdd.t146 4.06363
R5742 vdd.n175 vdd.t202 4.06363
R5743 vdd.n173 vdd.t232 4.06363
R5744 vdd.n173 vdd.t242 4.06363
R5745 vdd.n171 vdd.t245 4.06363
R5746 vdd.n171 vdd.t150 4.06363
R5747 vdd.n169 vdd.t173 4.06363
R5748 vdd.n169 vdd.t234 4.06363
R5749 vdd.n167 vdd.t246 4.06363
R5750 vdd.n167 vdd.t172 4.06363
R5751 vdd.n82 vdd.t207 4.06363
R5752 vdd.n82 vdd.t230 4.06363
R5753 vdd.n80 vdd.t192 4.06363
R5754 vdd.n80 vdd.t247 4.06363
R5755 vdd.n78 vdd.t163 4.06363
R5756 vdd.n78 vdd.t235 4.06363
R5757 vdd.n76 vdd.t156 4.06363
R5758 vdd.n76 vdd.t224 4.06363
R5759 vdd.n74 vdd.t175 4.06363
R5760 vdd.n74 vdd.t243 4.06363
R5761 vdd.n72 vdd.t152 4.06363
R5762 vdd.n72 vdd.t204 4.06363
R5763 vdd.n70 vdd.t139 4.06363
R5764 vdd.n70 vdd.t184 4.06363
R5765 vdd.n1769 vdd.t236 4.06363
R5766 vdd.n1769 vdd.t194 4.06363
R5767 vdd.n1771 vdd.t190 4.06363
R5768 vdd.n1771 vdd.t237 4.06363
R5769 vdd.n1773 vdd.t220 4.06363
R5770 vdd.n1773 vdd.t219 4.06363
R5771 vdd.n1775 vdd.t185 4.06363
R5772 vdd.n1775 vdd.t162 4.06363
R5773 vdd.n1777 vdd.t158 4.06363
R5774 vdd.n1777 vdd.t218 4.06363
R5775 vdd.n1779 vdd.t200 4.06363
R5776 vdd.n1779 vdd.t159 4.06363
R5777 vdd.n1781 vdd.t144 4.06363
R5778 vdd.n1781 vdd.t238 4.06363
R5779 vdd.n1671 vdd.t221 4.06363
R5780 vdd.n1671 vdd.t170 4.06363
R5781 vdd.n1673 vdd.t168 4.06363
R5782 vdd.n1673 vdd.t222 4.06363
R5783 vdd.n1675 vdd.t213 4.06363
R5784 vdd.n1675 vdd.t211 4.06363
R5785 vdd.n1677 vdd.t161 4.06363
R5786 vdd.n1677 vdd.t141 4.06363
R5787 vdd.n1679 vdd.t133 4.06363
R5788 vdd.n1679 vdd.t206 4.06363
R5789 vdd.n1681 vdd.t189 4.06363
R5790 vdd.n1681 vdd.t137 4.06363
R5791 vdd.n1683 vdd.t131 4.06363
R5792 vdd.n1683 vdd.t226 4.06363
R5793 vdd.n1574 vdd.t187 4.06363
R5794 vdd.n1574 vdd.t143 4.06363
R5795 vdd.n1576 vdd.t205 4.06363
R5796 vdd.n1576 vdd.t154 4.06363
R5797 vdd.n1578 vdd.t244 4.06363
R5798 vdd.n1578 vdd.t256 4.06363
R5799 vdd.n1580 vdd.t225 4.06363
R5800 vdd.n1580 vdd.t157 4.06363
R5801 vdd.n1582 vdd.t216 4.06363
R5802 vdd.n1582 vdd.t166 4.06363
R5803 vdd.n1584 vdd.t248 4.06363
R5804 vdd.n1584 vdd.t193 4.06363
R5805 vdd.n1586 vdd.t231 4.06363
R5806 vdd.n1586 vdd.t209 4.06363
R5807 vdd.n26 vdd.t25 3.9605
R5808 vdd.n26 vdd.t126 3.9605
R5809 vdd.n23 vdd.t123 3.9605
R5810 vdd.n23 vdd.t124 3.9605
R5811 vdd.n21 vdd.t32 3.9605
R5812 vdd.n21 vdd.t12 3.9605
R5813 vdd.n20 vdd.t129 3.9605
R5814 vdd.n20 vdd.t122 3.9605
R5815 vdd.n15 vdd.t127 3.9605
R5816 vdd.n15 vdd.t121 3.9605
R5817 vdd.n16 vdd.t128 3.9605
R5818 vdd.n16 vdd.t125 3.9605
R5819 vdd.n18 vdd.t33 3.9605
R5820 vdd.n18 vdd.t10 3.9605
R5821 vdd.n25 vdd.t24 3.9605
R5822 vdd.n25 vdd.t11 3.9605
R5823 vdd.n2997 vdd.n2996 3.74684
R5824 vdd.n2437 vdd.n2436 3.74684
R5825 vdd.n7 vdd.t22 3.61217
R5826 vdd.n7 vdd.t17 3.61217
R5827 vdd.n8 vdd.t269 3.61217
R5828 vdd.n8 vdd.t265 3.61217
R5829 vdd.n10 vdd.t115 3.61217
R5830 vdd.n10 vdd.t2 3.61217
R5831 vdd.n12 vdd.t120 3.61217
R5832 vdd.n12 vdd.t117 3.61217
R5833 vdd.n5 vdd.t261 3.61217
R5834 vdd.n5 vdd.t112 3.61217
R5835 vdd.n3 vdd.t15 3.61217
R5836 vdd.n3 vdd.t259 3.61217
R5837 vdd.n1 vdd.t263 3.61217
R5838 vdd.n1 vdd.t6 3.61217
R5839 vdd.n0 vdd.t267 3.61217
R5840 vdd.n0 vdd.t271 3.61217
R5841 vdd.n1462 vdd.t69 3.51482
R5842 vdd.n2414 vdd.t34 3.51482
R5843 vdd.n2469 vdd.t26 3.51482
R5844 vdd.n2964 vdd.t9 3.51482
R5845 vdd.n3019 vdd.t7 3.51482
R5846 vdd.n3437 vdd.t51 3.51482
R5847 vdd.n304 vdd.n303 3.49141
R5848 vdd.n249 vdd.n248 3.49141
R5849 vdd.n206 vdd.n205 3.49141
R5850 vdd.n151 vdd.n150 3.49141
R5851 vdd.n109 vdd.n108 3.49141
R5852 vdd.n54 vdd.n53 3.49141
R5853 vdd.n1753 vdd.n1752 3.49141
R5854 vdd.n1808 vdd.n1807 3.49141
R5855 vdd.n1655 vdd.n1654 3.49141
R5856 vdd.n1710 vdd.n1709 3.49141
R5857 vdd.n1558 vdd.n1557 3.49141
R5858 vdd.n1613 vdd.n1612 3.49141
R5859 vdd.n2489 vdd.t14 3.40145
R5860 vdd.n2643 vdd.t260 3.40145
R5861 vdd.n2927 vdd.t116 3.40145
R5862 vdd.n2946 vdd.t1 3.40145
R5863 vdd.n1865 vdd.t186 3.06136
R5864 vdd.n3359 vdd.t171 3.06136
R5865 vdd.t5 vdd.n986 2.94799
R5866 vdd.n901 vdd.t268 2.94799
R5867 vdd.t210 vdd.n1161 2.83463
R5868 vdd.n2390 vdd.t44 2.83463
R5869 vdd.n2496 vdd.t82 2.83463
R5870 vdd.n2940 vdd.t86 2.83463
R5871 vdd.n3088 vdd.t40 2.83463
R5872 vdd.n624 vdd.t174 2.83463
R5873 vdd.n307 vdd.n286 2.71565
R5874 vdd.n252 vdd.n231 2.71565
R5875 vdd.n209 vdd.n188 2.71565
R5876 vdd.n154 vdd.n133 2.71565
R5877 vdd.n112 vdd.n91 2.71565
R5878 vdd.n57 vdd.n36 2.71565
R5879 vdd.n1756 vdd.n1735 2.71565
R5880 vdd.n1811 vdd.n1790 2.71565
R5881 vdd.n1658 vdd.n1637 2.71565
R5882 vdd.n1713 vdd.n1692 2.71565
R5883 vdd.n1561 vdd.n1540 2.71565
R5884 vdd.n1616 vdd.n1595 2.71565
R5885 vdd.n1529 vdd.t160 2.6079
R5886 vdd.n1041 vdd.t27 2.6079
R5887 vdd.n2275 vdd.t23 2.6079
R5888 vdd.n2894 vdd.t118 2.6079
R5889 vdd.t0 vdd.n845 2.6079
R5890 vdd.n3469 vdd.t223 2.6079
R5891 vdd.n294 vdd.n293 2.4129
R5892 vdd.n239 vdd.n238 2.4129
R5893 vdd.n196 vdd.n195 2.4129
R5894 vdd.n141 vdd.n140 2.4129
R5895 vdd.n99 vdd.n98 2.4129
R5896 vdd.n44 vdd.n43 2.4129
R5897 vdd.n1743 vdd.n1742 2.4129
R5898 vdd.n1798 vdd.n1797 2.4129
R5899 vdd.n1645 vdd.n1644 2.4129
R5900 vdd.n1700 vdd.n1699 2.4129
R5901 vdd.n1548 vdd.n1547 2.4129
R5902 vdd.n1603 vdd.n1602 2.4129
R5903 vdd.t136 vdd.n1190 2.38117
R5904 vdd.n3460 vdd.t191 2.38117
R5905 vdd.n2099 vdd.n1901 2.27742
R5906 vdd.n2100 vdd.n2099 2.27742
R5907 vdd.n3124 vdd.n665 2.27742
R5908 vdd.n3124 vdd.n664 2.27742
R5909 vdd.n3192 vdd.n751 2.27742
R5910 vdd.n3192 vdd.n749 2.27742
R5911 vdd.n2122 vdd.n1116 2.27742
R5912 vdd.n2122 vdd.n1117 2.27742
R5913 vdd.n2275 vdd.t266 2.2678
R5914 vdd.n2894 vdd.t16 2.2678
R5915 vdd.n1487 vdd.t130 2.15444
R5916 vdd.n3451 vdd.t227 2.15444
R5917 vdd.n2463 vdd.t270 2.04107
R5918 vdd.n2970 vdd.t21 2.04107
R5919 vdd.n308 vdd.n284 1.93989
R5920 vdd.n253 vdd.n229 1.93989
R5921 vdd.n210 vdd.n186 1.93989
R5922 vdd.n155 vdd.n131 1.93989
R5923 vdd.n113 vdd.n89 1.93989
R5924 vdd.n58 vdd.n34 1.93989
R5925 vdd.n1757 vdd.n1733 1.93989
R5926 vdd.n1812 vdd.n1788 1.93989
R5927 vdd.n1659 vdd.n1635 1.93989
R5928 vdd.n1714 vdd.n1690 1.93989
R5929 vdd.n1562 vdd.n1538 1.93989
R5930 vdd.n1617 vdd.n1593 1.93989
R5931 vdd.n1479 vdd.t176 1.70098
R5932 vdd.n2439 vdd.t31 1.70098
R5933 vdd.n2445 vdd.t30 1.70098
R5934 vdd.n2988 vdd.t113 1.70098
R5935 vdd.n2994 vdd.t13 1.70098
R5936 vdd.n3445 vdd.t147 1.70098
R5937 vdd.n1495 vdd.t188 1.47425
R5938 vdd.n349 vdd.t134 1.47425
R5939 vdd.n2469 vdd.t262 1.36088
R5940 vdd.n2964 vdd.t264 1.36088
R5941 vdd.n1520 vdd.t165 1.24752
R5942 vdd.t62 vdd.n1124 1.24752
R5943 vdd.n659 vdd.t36 1.24752
R5944 vdd.t145 vdd.n3467 1.24752
R5945 vdd.n319 vdd.n279 1.16414
R5946 vdd.n312 vdd.n311 1.16414
R5947 vdd.n264 vdd.n224 1.16414
R5948 vdd.n257 vdd.n256 1.16414
R5949 vdd.n221 vdd.n181 1.16414
R5950 vdd.n214 vdd.n213 1.16414
R5951 vdd.n166 vdd.n126 1.16414
R5952 vdd.n159 vdd.n158 1.16414
R5953 vdd.n124 vdd.n84 1.16414
R5954 vdd.n117 vdd.n116 1.16414
R5955 vdd.n69 vdd.n29 1.16414
R5956 vdd.n62 vdd.n61 1.16414
R5957 vdd.n1768 vdd.n1728 1.16414
R5958 vdd.n1761 vdd.n1760 1.16414
R5959 vdd.n1823 vdd.n1783 1.16414
R5960 vdd.n1816 vdd.n1815 1.16414
R5961 vdd.n1670 vdd.n1630 1.16414
R5962 vdd.n1663 vdd.n1662 1.16414
R5963 vdd.n1725 vdd.n1685 1.16414
R5964 vdd.n1718 vdd.n1717 1.16414
R5965 vdd.n1573 vdd.n1533 1.16414
R5966 vdd.n1566 vdd.n1565 1.16414
R5967 vdd.n1628 vdd.n1588 1.16414
R5968 vdd.n1621 vdd.n1620 1.16414
R5969 vdd.n1826 vdd.n28 1.06035
R5970 vdd vdd.n3474 1.05252
R5971 vdd.n1172 vdd.t212 1.02079
R5972 vdd.t96 vdd.t31 1.02079
R5973 vdd.t13 vdd.t55 1.02079
R5974 vdd.t149 vdd.n613 1.02079
R5975 vdd.n1351 vdd.n1230 0.970197
R5976 vdd.n2120 vdd.n2119 0.970197
R5977 vdd.n599 vdd.n407 0.970197
R5978 vdd.n3199 vdd.n3197 0.970197
R5979 vdd.t258 vdd.n963 0.907421
R5980 vdd.n917 vdd.t114 0.907421
R5981 vdd.n1857 vdd.t153 0.794056
R5982 vdd.t19 vdd.n1038 0.794056
R5983 vdd.n1010 vdd.t8 0.794056
R5984 vdd.t29 vdd.n876 0.794056
R5985 vdd.n848 vdd.t3 0.794056
R5986 vdd.n3368 vdd.t151 0.794056
R5987 vdd.n1873 vdd.t214 0.567326
R5988 vdd.t182 vdd.n642 0.567326
R5989 vdd.n2110 vdd.n2109 0.482207
R5990 vdd.n3324 vdd.n3323 0.482207
R5991 vdd.n444 vdd.n443 0.482207
R5992 vdd.n3431 vdd.n3430 0.482207
R5993 vdd.n3330 vdd.n656 0.482207
R5994 vdd.n1887 vdd.n1118 0.482207
R5995 vdd.n1458 vdd.n1457 0.482207
R5996 vdd.n1264 vdd.n1221 0.482207
R5997 vdd.n4 vdd.n2 0.459552
R5998 vdd.n11 vdd.n9 0.459552
R5999 vdd.n317 vdd.n316 0.388379
R6000 vdd.n283 vdd.n281 0.388379
R6001 vdd.n262 vdd.n261 0.388379
R6002 vdd.n228 vdd.n226 0.388379
R6003 vdd.n219 vdd.n218 0.388379
R6004 vdd.n185 vdd.n183 0.388379
R6005 vdd.n164 vdd.n163 0.388379
R6006 vdd.n130 vdd.n128 0.388379
R6007 vdd.n122 vdd.n121 0.388379
R6008 vdd.n88 vdd.n86 0.388379
R6009 vdd.n67 vdd.n66 0.388379
R6010 vdd.n33 vdd.n31 0.388379
R6011 vdd.n1766 vdd.n1765 0.388379
R6012 vdd.n1732 vdd.n1730 0.388379
R6013 vdd.n1821 vdd.n1820 0.388379
R6014 vdd.n1787 vdd.n1785 0.388379
R6015 vdd.n1668 vdd.n1667 0.388379
R6016 vdd.n1634 vdd.n1632 0.388379
R6017 vdd.n1723 vdd.n1722 0.388379
R6018 vdd.n1689 vdd.n1687 0.388379
R6019 vdd.n1571 vdd.n1570 0.388379
R6020 vdd.n1537 vdd.n1535 0.388379
R6021 vdd.n1626 vdd.n1625 0.388379
R6022 vdd.n1592 vdd.n1590 0.388379
R6023 vdd.n19 vdd.n17 0.387128
R6024 vdd.n24 vdd.n22 0.387128
R6025 vdd.n6 vdd.n4 0.358259
R6026 vdd.n13 vdd.n11 0.358259
R6027 vdd.n268 vdd.n266 0.358259
R6028 vdd.n270 vdd.n268 0.358259
R6029 vdd.n272 vdd.n270 0.358259
R6030 vdd.n274 vdd.n272 0.358259
R6031 vdd.n276 vdd.n274 0.358259
R6032 vdd.n278 vdd.n276 0.358259
R6033 vdd.n320 vdd.n278 0.358259
R6034 vdd.n170 vdd.n168 0.358259
R6035 vdd.n172 vdd.n170 0.358259
R6036 vdd.n174 vdd.n172 0.358259
R6037 vdd.n176 vdd.n174 0.358259
R6038 vdd.n178 vdd.n176 0.358259
R6039 vdd.n180 vdd.n178 0.358259
R6040 vdd.n222 vdd.n180 0.358259
R6041 vdd.n73 vdd.n71 0.358259
R6042 vdd.n75 vdd.n73 0.358259
R6043 vdd.n77 vdd.n75 0.358259
R6044 vdd.n79 vdd.n77 0.358259
R6045 vdd.n81 vdd.n79 0.358259
R6046 vdd.n83 vdd.n81 0.358259
R6047 vdd.n125 vdd.n83 0.358259
R6048 vdd.n1824 vdd.n1782 0.358259
R6049 vdd.n1782 vdd.n1780 0.358259
R6050 vdd.n1780 vdd.n1778 0.358259
R6051 vdd.n1778 vdd.n1776 0.358259
R6052 vdd.n1776 vdd.n1774 0.358259
R6053 vdd.n1774 vdd.n1772 0.358259
R6054 vdd.n1772 vdd.n1770 0.358259
R6055 vdd.n1726 vdd.n1684 0.358259
R6056 vdd.n1684 vdd.n1682 0.358259
R6057 vdd.n1682 vdd.n1680 0.358259
R6058 vdd.n1680 vdd.n1678 0.358259
R6059 vdd.n1678 vdd.n1676 0.358259
R6060 vdd.n1676 vdd.n1674 0.358259
R6061 vdd.n1674 vdd.n1672 0.358259
R6062 vdd.n1629 vdd.n1587 0.358259
R6063 vdd.n1587 vdd.n1585 0.358259
R6064 vdd.n1585 vdd.n1583 0.358259
R6065 vdd.n1583 vdd.n1581 0.358259
R6066 vdd.n1581 vdd.n1579 0.358259
R6067 vdd.n1579 vdd.n1577 0.358259
R6068 vdd.n1577 vdd.n1575 0.358259
R6069 vdd.n14 vdd.n6 0.334552
R6070 vdd.n14 vdd.n13 0.334552
R6071 vdd.n27 vdd.n19 0.21707
R6072 vdd.n27 vdd.n24 0.21707
R6073 vdd.n318 vdd.n280 0.155672
R6074 vdd.n310 vdd.n280 0.155672
R6075 vdd.n310 vdd.n309 0.155672
R6076 vdd.n309 vdd.n285 0.155672
R6077 vdd.n302 vdd.n285 0.155672
R6078 vdd.n302 vdd.n301 0.155672
R6079 vdd.n301 vdd.n289 0.155672
R6080 vdd.n294 vdd.n289 0.155672
R6081 vdd.n263 vdd.n225 0.155672
R6082 vdd.n255 vdd.n225 0.155672
R6083 vdd.n255 vdd.n254 0.155672
R6084 vdd.n254 vdd.n230 0.155672
R6085 vdd.n247 vdd.n230 0.155672
R6086 vdd.n247 vdd.n246 0.155672
R6087 vdd.n246 vdd.n234 0.155672
R6088 vdd.n239 vdd.n234 0.155672
R6089 vdd.n220 vdd.n182 0.155672
R6090 vdd.n212 vdd.n182 0.155672
R6091 vdd.n212 vdd.n211 0.155672
R6092 vdd.n211 vdd.n187 0.155672
R6093 vdd.n204 vdd.n187 0.155672
R6094 vdd.n204 vdd.n203 0.155672
R6095 vdd.n203 vdd.n191 0.155672
R6096 vdd.n196 vdd.n191 0.155672
R6097 vdd.n165 vdd.n127 0.155672
R6098 vdd.n157 vdd.n127 0.155672
R6099 vdd.n157 vdd.n156 0.155672
R6100 vdd.n156 vdd.n132 0.155672
R6101 vdd.n149 vdd.n132 0.155672
R6102 vdd.n149 vdd.n148 0.155672
R6103 vdd.n148 vdd.n136 0.155672
R6104 vdd.n141 vdd.n136 0.155672
R6105 vdd.n123 vdd.n85 0.155672
R6106 vdd.n115 vdd.n85 0.155672
R6107 vdd.n115 vdd.n114 0.155672
R6108 vdd.n114 vdd.n90 0.155672
R6109 vdd.n107 vdd.n90 0.155672
R6110 vdd.n107 vdd.n106 0.155672
R6111 vdd.n106 vdd.n94 0.155672
R6112 vdd.n99 vdd.n94 0.155672
R6113 vdd.n68 vdd.n30 0.155672
R6114 vdd.n60 vdd.n30 0.155672
R6115 vdd.n60 vdd.n59 0.155672
R6116 vdd.n59 vdd.n35 0.155672
R6117 vdd.n52 vdd.n35 0.155672
R6118 vdd.n52 vdd.n51 0.155672
R6119 vdd.n51 vdd.n39 0.155672
R6120 vdd.n44 vdd.n39 0.155672
R6121 vdd.n1767 vdd.n1729 0.155672
R6122 vdd.n1759 vdd.n1729 0.155672
R6123 vdd.n1759 vdd.n1758 0.155672
R6124 vdd.n1758 vdd.n1734 0.155672
R6125 vdd.n1751 vdd.n1734 0.155672
R6126 vdd.n1751 vdd.n1750 0.155672
R6127 vdd.n1750 vdd.n1738 0.155672
R6128 vdd.n1743 vdd.n1738 0.155672
R6129 vdd.n1822 vdd.n1784 0.155672
R6130 vdd.n1814 vdd.n1784 0.155672
R6131 vdd.n1814 vdd.n1813 0.155672
R6132 vdd.n1813 vdd.n1789 0.155672
R6133 vdd.n1806 vdd.n1789 0.155672
R6134 vdd.n1806 vdd.n1805 0.155672
R6135 vdd.n1805 vdd.n1793 0.155672
R6136 vdd.n1798 vdd.n1793 0.155672
R6137 vdd.n1669 vdd.n1631 0.155672
R6138 vdd.n1661 vdd.n1631 0.155672
R6139 vdd.n1661 vdd.n1660 0.155672
R6140 vdd.n1660 vdd.n1636 0.155672
R6141 vdd.n1653 vdd.n1636 0.155672
R6142 vdd.n1653 vdd.n1652 0.155672
R6143 vdd.n1652 vdd.n1640 0.155672
R6144 vdd.n1645 vdd.n1640 0.155672
R6145 vdd.n1724 vdd.n1686 0.155672
R6146 vdd.n1716 vdd.n1686 0.155672
R6147 vdd.n1716 vdd.n1715 0.155672
R6148 vdd.n1715 vdd.n1691 0.155672
R6149 vdd.n1708 vdd.n1691 0.155672
R6150 vdd.n1708 vdd.n1707 0.155672
R6151 vdd.n1707 vdd.n1695 0.155672
R6152 vdd.n1700 vdd.n1695 0.155672
R6153 vdd.n1572 vdd.n1534 0.155672
R6154 vdd.n1564 vdd.n1534 0.155672
R6155 vdd.n1564 vdd.n1563 0.155672
R6156 vdd.n1563 vdd.n1539 0.155672
R6157 vdd.n1556 vdd.n1539 0.155672
R6158 vdd.n1556 vdd.n1555 0.155672
R6159 vdd.n1555 vdd.n1543 0.155672
R6160 vdd.n1548 vdd.n1543 0.155672
R6161 vdd.n1627 vdd.n1589 0.155672
R6162 vdd.n1619 vdd.n1589 0.155672
R6163 vdd.n1619 vdd.n1618 0.155672
R6164 vdd.n1618 vdd.n1594 0.155672
R6165 vdd.n1611 vdd.n1594 0.155672
R6166 vdd.n1611 vdd.n1610 0.155672
R6167 vdd.n1610 vdd.n1598 0.155672
R6168 vdd.n1603 vdd.n1598 0.155672
R6169 vdd.n2098 vdd.n1903 0.152939
R6170 vdd.n1909 vdd.n1903 0.152939
R6171 vdd.n1910 vdd.n1909 0.152939
R6172 vdd.n1911 vdd.n1910 0.152939
R6173 vdd.n1912 vdd.n1911 0.152939
R6174 vdd.n1916 vdd.n1912 0.152939
R6175 vdd.n1917 vdd.n1916 0.152939
R6176 vdd.n1918 vdd.n1917 0.152939
R6177 vdd.n1919 vdd.n1918 0.152939
R6178 vdd.n1923 vdd.n1919 0.152939
R6179 vdd.n1924 vdd.n1923 0.152939
R6180 vdd.n1925 vdd.n1924 0.152939
R6181 vdd.n2073 vdd.n1925 0.152939
R6182 vdd.n2073 vdd.n2072 0.152939
R6183 vdd.n2072 vdd.n2071 0.152939
R6184 vdd.n2071 vdd.n1931 0.152939
R6185 vdd.n1936 vdd.n1931 0.152939
R6186 vdd.n1937 vdd.n1936 0.152939
R6187 vdd.n1938 vdd.n1937 0.152939
R6188 vdd.n1942 vdd.n1938 0.152939
R6189 vdd.n1943 vdd.n1942 0.152939
R6190 vdd.n1944 vdd.n1943 0.152939
R6191 vdd.n1945 vdd.n1944 0.152939
R6192 vdd.n1949 vdd.n1945 0.152939
R6193 vdd.n1950 vdd.n1949 0.152939
R6194 vdd.n1951 vdd.n1950 0.152939
R6195 vdd.n1952 vdd.n1951 0.152939
R6196 vdd.n1956 vdd.n1952 0.152939
R6197 vdd.n1957 vdd.n1956 0.152939
R6198 vdd.n1958 vdd.n1957 0.152939
R6199 vdd.n1959 vdd.n1958 0.152939
R6200 vdd.n1963 vdd.n1959 0.152939
R6201 vdd.n1964 vdd.n1963 0.152939
R6202 vdd.n1965 vdd.n1964 0.152939
R6203 vdd.n2034 vdd.n1965 0.152939
R6204 vdd.n2034 vdd.n2033 0.152939
R6205 vdd.n2033 vdd.n2032 0.152939
R6206 vdd.n2032 vdd.n1971 0.152939
R6207 vdd.n1976 vdd.n1971 0.152939
R6208 vdd.n1977 vdd.n1976 0.152939
R6209 vdd.n1978 vdd.n1977 0.152939
R6210 vdd.n1982 vdd.n1978 0.152939
R6211 vdd.n1983 vdd.n1982 0.152939
R6212 vdd.n1984 vdd.n1983 0.152939
R6213 vdd.n1985 vdd.n1984 0.152939
R6214 vdd.n1989 vdd.n1985 0.152939
R6215 vdd.n1990 vdd.n1989 0.152939
R6216 vdd.n1991 vdd.n1990 0.152939
R6217 vdd.n1992 vdd.n1991 0.152939
R6218 vdd.n1993 vdd.n1992 0.152939
R6219 vdd.n1993 vdd.n1115 0.152939
R6220 vdd.n2109 vdd.n1897 0.152939
R6221 vdd.n1829 vdd.n1828 0.152939
R6222 vdd.n1829 vdd.n1164 0.152939
R6223 vdd.n1843 vdd.n1164 0.152939
R6224 vdd.n1844 vdd.n1843 0.152939
R6225 vdd.n1845 vdd.n1844 0.152939
R6226 vdd.n1845 vdd.n1152 0.152939
R6227 vdd.n1860 vdd.n1152 0.152939
R6228 vdd.n1861 vdd.n1860 0.152939
R6229 vdd.n1862 vdd.n1861 0.152939
R6230 vdd.n1862 vdd.n1141 0.152939
R6231 vdd.n1877 vdd.n1141 0.152939
R6232 vdd.n1878 vdd.n1877 0.152939
R6233 vdd.n1879 vdd.n1878 0.152939
R6234 vdd.n1879 vdd.n1129 0.152939
R6235 vdd.n1895 vdd.n1129 0.152939
R6236 vdd.n1896 vdd.n1895 0.152939
R6237 vdd.n2110 vdd.n1896 0.152939
R6238 vdd.n670 vdd.n667 0.152939
R6239 vdd.n671 vdd.n670 0.152939
R6240 vdd.n672 vdd.n671 0.152939
R6241 vdd.n673 vdd.n672 0.152939
R6242 vdd.n676 vdd.n673 0.152939
R6243 vdd.n677 vdd.n676 0.152939
R6244 vdd.n678 vdd.n677 0.152939
R6245 vdd.n679 vdd.n678 0.152939
R6246 vdd.n682 vdd.n679 0.152939
R6247 vdd.n683 vdd.n682 0.152939
R6248 vdd.n684 vdd.n683 0.152939
R6249 vdd.n685 vdd.n684 0.152939
R6250 vdd.n690 vdd.n685 0.152939
R6251 vdd.n691 vdd.n690 0.152939
R6252 vdd.n692 vdd.n691 0.152939
R6253 vdd.n693 vdd.n692 0.152939
R6254 vdd.n696 vdd.n693 0.152939
R6255 vdd.n697 vdd.n696 0.152939
R6256 vdd.n698 vdd.n697 0.152939
R6257 vdd.n699 vdd.n698 0.152939
R6258 vdd.n702 vdd.n699 0.152939
R6259 vdd.n703 vdd.n702 0.152939
R6260 vdd.n704 vdd.n703 0.152939
R6261 vdd.n705 vdd.n704 0.152939
R6262 vdd.n708 vdd.n705 0.152939
R6263 vdd.n709 vdd.n708 0.152939
R6264 vdd.n710 vdd.n709 0.152939
R6265 vdd.n711 vdd.n710 0.152939
R6266 vdd.n714 vdd.n711 0.152939
R6267 vdd.n715 vdd.n714 0.152939
R6268 vdd.n716 vdd.n715 0.152939
R6269 vdd.n717 vdd.n716 0.152939
R6270 vdd.n720 vdd.n717 0.152939
R6271 vdd.n721 vdd.n720 0.152939
R6272 vdd.n3240 vdd.n721 0.152939
R6273 vdd.n3240 vdd.n3239 0.152939
R6274 vdd.n3239 vdd.n3238 0.152939
R6275 vdd.n3238 vdd.n725 0.152939
R6276 vdd.n730 vdd.n725 0.152939
R6277 vdd.n731 vdd.n730 0.152939
R6278 vdd.n734 vdd.n731 0.152939
R6279 vdd.n735 vdd.n734 0.152939
R6280 vdd.n736 vdd.n735 0.152939
R6281 vdd.n737 vdd.n736 0.152939
R6282 vdd.n740 vdd.n737 0.152939
R6283 vdd.n741 vdd.n740 0.152939
R6284 vdd.n742 vdd.n741 0.152939
R6285 vdd.n743 vdd.n742 0.152939
R6286 vdd.n746 vdd.n743 0.152939
R6287 vdd.n747 vdd.n746 0.152939
R6288 vdd.n748 vdd.n747 0.152939
R6289 vdd.n3323 vdd.n661 0.152939
R6290 vdd.n3324 vdd.n651 0.152939
R6291 vdd.n3338 vdd.n651 0.152939
R6292 vdd.n3339 vdd.n3338 0.152939
R6293 vdd.n3340 vdd.n3339 0.152939
R6294 vdd.n3340 vdd.n639 0.152939
R6295 vdd.n3354 vdd.n639 0.152939
R6296 vdd.n3355 vdd.n3354 0.152939
R6297 vdd.n3356 vdd.n3355 0.152939
R6298 vdd.n3356 vdd.n627 0.152939
R6299 vdd.n3371 vdd.n627 0.152939
R6300 vdd.n3372 vdd.n3371 0.152939
R6301 vdd.n3373 vdd.n3372 0.152939
R6302 vdd.n3373 vdd.n616 0.152939
R6303 vdd.n3390 vdd.n616 0.152939
R6304 vdd.n3391 vdd.n3390 0.152939
R6305 vdd.n3392 vdd.n3391 0.152939
R6306 vdd.n3392 vdd.n322 0.152939
R6307 vdd.n3472 vdd.n323 0.152939
R6308 vdd.n334 vdd.n323 0.152939
R6309 vdd.n335 vdd.n334 0.152939
R6310 vdd.n336 vdd.n335 0.152939
R6311 vdd.n343 vdd.n336 0.152939
R6312 vdd.n344 vdd.n343 0.152939
R6313 vdd.n345 vdd.n344 0.152939
R6314 vdd.n346 vdd.n345 0.152939
R6315 vdd.n354 vdd.n346 0.152939
R6316 vdd.n355 vdd.n354 0.152939
R6317 vdd.n356 vdd.n355 0.152939
R6318 vdd.n357 vdd.n356 0.152939
R6319 vdd.n365 vdd.n357 0.152939
R6320 vdd.n366 vdd.n365 0.152939
R6321 vdd.n367 vdd.n366 0.152939
R6322 vdd.n368 vdd.n367 0.152939
R6323 vdd.n443 vdd.n368 0.152939
R6324 vdd.n444 vdd.n442 0.152939
R6325 vdd.n451 vdd.n442 0.152939
R6326 vdd.n452 vdd.n451 0.152939
R6327 vdd.n453 vdd.n452 0.152939
R6328 vdd.n453 vdd.n440 0.152939
R6329 vdd.n461 vdd.n440 0.152939
R6330 vdd.n462 vdd.n461 0.152939
R6331 vdd.n463 vdd.n462 0.152939
R6332 vdd.n463 vdd.n438 0.152939
R6333 vdd.n471 vdd.n438 0.152939
R6334 vdd.n472 vdd.n471 0.152939
R6335 vdd.n473 vdd.n472 0.152939
R6336 vdd.n473 vdd.n436 0.152939
R6337 vdd.n481 vdd.n436 0.152939
R6338 vdd.n482 vdd.n481 0.152939
R6339 vdd.n483 vdd.n482 0.152939
R6340 vdd.n483 vdd.n434 0.152939
R6341 vdd.n491 vdd.n434 0.152939
R6342 vdd.n492 vdd.n491 0.152939
R6343 vdd.n493 vdd.n492 0.152939
R6344 vdd.n493 vdd.n430 0.152939
R6345 vdd.n501 vdd.n430 0.152939
R6346 vdd.n502 vdd.n501 0.152939
R6347 vdd.n503 vdd.n502 0.152939
R6348 vdd.n503 vdd.n428 0.152939
R6349 vdd.n511 vdd.n428 0.152939
R6350 vdd.n512 vdd.n511 0.152939
R6351 vdd.n513 vdd.n512 0.152939
R6352 vdd.n513 vdd.n426 0.152939
R6353 vdd.n521 vdd.n426 0.152939
R6354 vdd.n522 vdd.n521 0.152939
R6355 vdd.n523 vdd.n522 0.152939
R6356 vdd.n523 vdd.n424 0.152939
R6357 vdd.n531 vdd.n424 0.152939
R6358 vdd.n532 vdd.n531 0.152939
R6359 vdd.n533 vdd.n532 0.152939
R6360 vdd.n533 vdd.n422 0.152939
R6361 vdd.n541 vdd.n422 0.152939
R6362 vdd.n542 vdd.n541 0.152939
R6363 vdd.n543 vdd.n542 0.152939
R6364 vdd.n543 vdd.n418 0.152939
R6365 vdd.n551 vdd.n418 0.152939
R6366 vdd.n552 vdd.n551 0.152939
R6367 vdd.n553 vdd.n552 0.152939
R6368 vdd.n553 vdd.n416 0.152939
R6369 vdd.n561 vdd.n416 0.152939
R6370 vdd.n562 vdd.n561 0.152939
R6371 vdd.n563 vdd.n562 0.152939
R6372 vdd.n563 vdd.n414 0.152939
R6373 vdd.n571 vdd.n414 0.152939
R6374 vdd.n572 vdd.n571 0.152939
R6375 vdd.n573 vdd.n572 0.152939
R6376 vdd.n573 vdd.n412 0.152939
R6377 vdd.n581 vdd.n412 0.152939
R6378 vdd.n582 vdd.n581 0.152939
R6379 vdd.n583 vdd.n582 0.152939
R6380 vdd.n583 vdd.n410 0.152939
R6381 vdd.n591 vdd.n410 0.152939
R6382 vdd.n592 vdd.n591 0.152939
R6383 vdd.n593 vdd.n592 0.152939
R6384 vdd.n593 vdd.n408 0.152939
R6385 vdd.n600 vdd.n408 0.152939
R6386 vdd.n3431 vdd.n600 0.152939
R6387 vdd.n3331 vdd.n3330 0.152939
R6388 vdd.n3332 vdd.n3331 0.152939
R6389 vdd.n3332 vdd.n645 0.152939
R6390 vdd.n3346 vdd.n645 0.152939
R6391 vdd.n3347 vdd.n3346 0.152939
R6392 vdd.n3348 vdd.n3347 0.152939
R6393 vdd.n3348 vdd.n632 0.152939
R6394 vdd.n3362 vdd.n632 0.152939
R6395 vdd.n3363 vdd.n3362 0.152939
R6396 vdd.n3364 vdd.n3363 0.152939
R6397 vdd.n3364 vdd.n621 0.152939
R6398 vdd.n3379 vdd.n621 0.152939
R6399 vdd.n3380 vdd.n3379 0.152939
R6400 vdd.n3381 vdd.n3380 0.152939
R6401 vdd.n3383 vdd.n3381 0.152939
R6402 vdd.n3383 vdd.n3382 0.152939
R6403 vdd.n3382 vdd.n611 0.152939
R6404 vdd.n611 vdd.n609 0.152939
R6405 vdd.n3401 vdd.n609 0.152939
R6406 vdd.n3402 vdd.n3401 0.152939
R6407 vdd.n3403 vdd.n3402 0.152939
R6408 vdd.n3403 vdd.n607 0.152939
R6409 vdd.n3408 vdd.n607 0.152939
R6410 vdd.n3409 vdd.n3408 0.152939
R6411 vdd.n3410 vdd.n3409 0.152939
R6412 vdd.n3410 vdd.n605 0.152939
R6413 vdd.n3415 vdd.n605 0.152939
R6414 vdd.n3416 vdd.n3415 0.152939
R6415 vdd.n3417 vdd.n3416 0.152939
R6416 vdd.n3417 vdd.n603 0.152939
R6417 vdd.n3423 vdd.n603 0.152939
R6418 vdd.n3424 vdd.n3423 0.152939
R6419 vdd.n3425 vdd.n3424 0.152939
R6420 vdd.n3425 vdd.n601 0.152939
R6421 vdd.n3430 vdd.n601 0.152939
R6422 vdd.n3193 vdd.n656 0.152939
R6423 vdd.n2121 vdd.n1118 0.152939
R6424 vdd.n1459 vdd.n1458 0.152939
R6425 vdd.n1459 vdd.n1215 0.152939
R6426 vdd.n1473 vdd.n1215 0.152939
R6427 vdd.n1474 vdd.n1473 0.152939
R6428 vdd.n1475 vdd.n1474 0.152939
R6429 vdd.n1475 vdd.n1203 0.152939
R6430 vdd.n1490 vdd.n1203 0.152939
R6431 vdd.n1491 vdd.n1490 0.152939
R6432 vdd.n1492 vdd.n1491 0.152939
R6433 vdd.n1492 vdd.n1193 0.152939
R6434 vdd.n1507 vdd.n1193 0.152939
R6435 vdd.n1508 vdd.n1507 0.152939
R6436 vdd.n1509 vdd.n1508 0.152939
R6437 vdd.n1509 vdd.n1180 0.152939
R6438 vdd.n1523 vdd.n1180 0.152939
R6439 vdd.n1524 vdd.n1523 0.152939
R6440 vdd.n1525 vdd.n1524 0.152939
R6441 vdd.n1525 vdd.n1169 0.152939
R6442 vdd.n1835 vdd.n1169 0.152939
R6443 vdd.n1836 vdd.n1835 0.152939
R6444 vdd.n1837 vdd.n1836 0.152939
R6445 vdd.n1837 vdd.n1158 0.152939
R6446 vdd.n1851 vdd.n1158 0.152939
R6447 vdd.n1852 vdd.n1851 0.152939
R6448 vdd.n1853 vdd.n1852 0.152939
R6449 vdd.n1853 vdd.n1146 0.152939
R6450 vdd.n1868 vdd.n1146 0.152939
R6451 vdd.n1869 vdd.n1868 0.152939
R6452 vdd.n1870 vdd.n1869 0.152939
R6453 vdd.n1870 vdd.n1136 0.152939
R6454 vdd.n1885 vdd.n1136 0.152939
R6455 vdd.n1886 vdd.n1885 0.152939
R6456 vdd.n1889 vdd.n1886 0.152939
R6457 vdd.n1889 vdd.n1888 0.152939
R6458 vdd.n1888 vdd.n1887 0.152939
R6459 vdd.n1449 vdd.n1264 0.152939
R6460 vdd.n1449 vdd.n1448 0.152939
R6461 vdd.n1448 vdd.n1447 0.152939
R6462 vdd.n1447 vdd.n1266 0.152939
R6463 vdd.n1443 vdd.n1266 0.152939
R6464 vdd.n1443 vdd.n1442 0.152939
R6465 vdd.n1442 vdd.n1441 0.152939
R6466 vdd.n1441 vdd.n1271 0.152939
R6467 vdd.n1437 vdd.n1271 0.152939
R6468 vdd.n1437 vdd.n1436 0.152939
R6469 vdd.n1436 vdd.n1435 0.152939
R6470 vdd.n1435 vdd.n1277 0.152939
R6471 vdd.n1431 vdd.n1277 0.152939
R6472 vdd.n1431 vdd.n1430 0.152939
R6473 vdd.n1430 vdd.n1429 0.152939
R6474 vdd.n1429 vdd.n1283 0.152939
R6475 vdd.n1425 vdd.n1283 0.152939
R6476 vdd.n1425 vdd.n1424 0.152939
R6477 vdd.n1424 vdd.n1423 0.152939
R6478 vdd.n1423 vdd.n1289 0.152939
R6479 vdd.n1415 vdd.n1289 0.152939
R6480 vdd.n1415 vdd.n1414 0.152939
R6481 vdd.n1414 vdd.n1413 0.152939
R6482 vdd.n1413 vdd.n1293 0.152939
R6483 vdd.n1409 vdd.n1293 0.152939
R6484 vdd.n1409 vdd.n1408 0.152939
R6485 vdd.n1408 vdd.n1407 0.152939
R6486 vdd.n1407 vdd.n1299 0.152939
R6487 vdd.n1403 vdd.n1299 0.152939
R6488 vdd.n1403 vdd.n1402 0.152939
R6489 vdd.n1402 vdd.n1401 0.152939
R6490 vdd.n1401 vdd.n1305 0.152939
R6491 vdd.n1397 vdd.n1305 0.152939
R6492 vdd.n1397 vdd.n1396 0.152939
R6493 vdd.n1396 vdd.n1395 0.152939
R6494 vdd.n1395 vdd.n1311 0.152939
R6495 vdd.n1391 vdd.n1311 0.152939
R6496 vdd.n1391 vdd.n1390 0.152939
R6497 vdd.n1390 vdd.n1389 0.152939
R6498 vdd.n1389 vdd.n1317 0.152939
R6499 vdd.n1382 vdd.n1317 0.152939
R6500 vdd.n1382 vdd.n1381 0.152939
R6501 vdd.n1381 vdd.n1380 0.152939
R6502 vdd.n1380 vdd.n1322 0.152939
R6503 vdd.n1376 vdd.n1322 0.152939
R6504 vdd.n1376 vdd.n1375 0.152939
R6505 vdd.n1375 vdd.n1374 0.152939
R6506 vdd.n1374 vdd.n1328 0.152939
R6507 vdd.n1370 vdd.n1328 0.152939
R6508 vdd.n1370 vdd.n1369 0.152939
R6509 vdd.n1369 vdd.n1368 0.152939
R6510 vdd.n1368 vdd.n1334 0.152939
R6511 vdd.n1364 vdd.n1334 0.152939
R6512 vdd.n1364 vdd.n1363 0.152939
R6513 vdd.n1363 vdd.n1362 0.152939
R6514 vdd.n1362 vdd.n1340 0.152939
R6515 vdd.n1358 vdd.n1340 0.152939
R6516 vdd.n1358 vdd.n1357 0.152939
R6517 vdd.n1357 vdd.n1356 0.152939
R6518 vdd.n1356 vdd.n1346 0.152939
R6519 vdd.n1352 vdd.n1346 0.152939
R6520 vdd.n1352 vdd.n1227 0.152939
R6521 vdd.n1457 vdd.n1227 0.152939
R6522 vdd.n1465 vdd.n1221 0.152939
R6523 vdd.n1466 vdd.n1465 0.152939
R6524 vdd.n1467 vdd.n1466 0.152939
R6525 vdd.n1467 vdd.n1209 0.152939
R6526 vdd.n1482 vdd.n1209 0.152939
R6527 vdd.n1483 vdd.n1482 0.152939
R6528 vdd.n1484 vdd.n1483 0.152939
R6529 vdd.n1484 vdd.n1198 0.152939
R6530 vdd.n1499 vdd.n1198 0.152939
R6531 vdd.n1500 vdd.n1499 0.152939
R6532 vdd.n1501 vdd.n1500 0.152939
R6533 vdd.n1501 vdd.n1187 0.152939
R6534 vdd.n1515 vdd.n1187 0.152939
R6535 vdd.n1516 vdd.n1515 0.152939
R6536 vdd.n1517 vdd.n1516 0.152939
R6537 vdd.n1517 vdd.n1175 0.152939
R6538 vdd.n1532 vdd.n1175 0.152939
R6539 vdd.n2408 vdd.t20 0.113865
R6540 vdd.n2475 vdd.t4 0.113865
R6541 vdd.n2958 vdd.t18 0.113865
R6542 vdd.n3025 vdd.t28 0.113865
R6543 vdd.n2099 vdd.n1897 0.110256
R6544 vdd.n3124 vdd.n661 0.110256
R6545 vdd.n3193 vdd.n3192 0.110256
R6546 vdd.n2122 vdd.n2121 0.110256
R6547 vdd.n1828 vdd.n1827 0.0695946
R6548 vdd.n3473 vdd.n322 0.0695946
R6549 vdd.n3473 vdd.n3472 0.0695946
R6550 vdd.n1827 vdd.n1532 0.0695946
R6551 vdd.n2099 vdd.n2098 0.0431829
R6552 vdd.n2122 vdd.n1115 0.0431829
R6553 vdd.n3124 vdd.n667 0.0431829
R6554 vdd.n3192 vdd.n748 0.0431829
R6555 vdd vdd.n28 0.00833333
R6556 CSoutput.n19 CSoutput.t164 184.661
R6557 CSoutput.n78 CSoutput.n77 165.8
R6558 CSoutput.n76 CSoutput.n0 165.8
R6559 CSoutput.n75 CSoutput.n74 165.8
R6560 CSoutput.n73 CSoutput.n72 165.8
R6561 CSoutput.n71 CSoutput.n2 165.8
R6562 CSoutput.n69 CSoutput.n68 165.8
R6563 CSoutput.n67 CSoutput.n3 165.8
R6564 CSoutput.n66 CSoutput.n65 165.8
R6565 CSoutput.n63 CSoutput.n4 165.8
R6566 CSoutput.n61 CSoutput.n60 165.8
R6567 CSoutput.n59 CSoutput.n5 165.8
R6568 CSoutput.n58 CSoutput.n57 165.8
R6569 CSoutput.n55 CSoutput.n6 165.8
R6570 CSoutput.n54 CSoutput.n53 165.8
R6571 CSoutput.n52 CSoutput.n51 165.8
R6572 CSoutput.n50 CSoutput.n8 165.8
R6573 CSoutput.n48 CSoutput.n47 165.8
R6574 CSoutput.n46 CSoutput.n9 165.8
R6575 CSoutput.n45 CSoutput.n44 165.8
R6576 CSoutput.n42 CSoutput.n10 165.8
R6577 CSoutput.n41 CSoutput.n40 165.8
R6578 CSoutput.n39 CSoutput.n38 165.8
R6579 CSoutput.n37 CSoutput.n12 165.8
R6580 CSoutput.n35 CSoutput.n34 165.8
R6581 CSoutput.n33 CSoutput.n13 165.8
R6582 CSoutput.n32 CSoutput.n31 165.8
R6583 CSoutput.n29 CSoutput.n14 165.8
R6584 CSoutput.n28 CSoutput.n27 165.8
R6585 CSoutput.n26 CSoutput.n25 165.8
R6586 CSoutput.n24 CSoutput.n16 165.8
R6587 CSoutput.n22 CSoutput.n21 165.8
R6588 CSoutput.n20 CSoutput.n17 165.8
R6589 CSoutput.n77 CSoutput.t165 162.194
R6590 CSoutput.n18 CSoutput.t166 120.501
R6591 CSoutput.n23 CSoutput.t174 120.501
R6592 CSoutput.n15 CSoutput.t170 120.501
R6593 CSoutput.n30 CSoutput.t167 120.501
R6594 CSoutput.n36 CSoutput.t177 120.501
R6595 CSoutput.n11 CSoutput.t180 120.501
R6596 CSoutput.n43 CSoutput.t169 120.501
R6597 CSoutput.n49 CSoutput.t181 120.501
R6598 CSoutput.n7 CSoutput.t160 120.501
R6599 CSoutput.n56 CSoutput.t176 120.501
R6600 CSoutput.n62 CSoutput.t168 120.501
R6601 CSoutput.n64 CSoutput.t162 120.501
R6602 CSoutput.n70 CSoutput.t179 120.501
R6603 CSoutput.n1 CSoutput.t173 120.501
R6604 CSoutput.n310 CSoutput.n308 103.469
R6605 CSoutput.n294 CSoutput.n292 103.469
R6606 CSoutput.n279 CSoutput.n277 103.469
R6607 CSoutput.n112 CSoutput.n110 103.469
R6608 CSoutput.n96 CSoutput.n94 103.469
R6609 CSoutput.n81 CSoutput.n79 103.469
R6610 CSoutput.n320 CSoutput.n319 103.111
R6611 CSoutput.n318 CSoutput.n317 103.111
R6612 CSoutput.n316 CSoutput.n315 103.111
R6613 CSoutput.n314 CSoutput.n313 103.111
R6614 CSoutput.n312 CSoutput.n311 103.111
R6615 CSoutput.n310 CSoutput.n309 103.111
R6616 CSoutput.n306 CSoutput.n305 103.111
R6617 CSoutput.n304 CSoutput.n303 103.111
R6618 CSoutput.n302 CSoutput.n301 103.111
R6619 CSoutput.n300 CSoutput.n299 103.111
R6620 CSoutput.n298 CSoutput.n297 103.111
R6621 CSoutput.n296 CSoutput.n295 103.111
R6622 CSoutput.n294 CSoutput.n293 103.111
R6623 CSoutput.n291 CSoutput.n290 103.111
R6624 CSoutput.n289 CSoutput.n288 103.111
R6625 CSoutput.n287 CSoutput.n286 103.111
R6626 CSoutput.n285 CSoutput.n284 103.111
R6627 CSoutput.n283 CSoutput.n282 103.111
R6628 CSoutput.n281 CSoutput.n280 103.111
R6629 CSoutput.n279 CSoutput.n278 103.111
R6630 CSoutput.n112 CSoutput.n111 103.111
R6631 CSoutput.n114 CSoutput.n113 103.111
R6632 CSoutput.n116 CSoutput.n115 103.111
R6633 CSoutput.n118 CSoutput.n117 103.111
R6634 CSoutput.n120 CSoutput.n119 103.111
R6635 CSoutput.n122 CSoutput.n121 103.111
R6636 CSoutput.n124 CSoutput.n123 103.111
R6637 CSoutput.n96 CSoutput.n95 103.111
R6638 CSoutput.n98 CSoutput.n97 103.111
R6639 CSoutput.n100 CSoutput.n99 103.111
R6640 CSoutput.n102 CSoutput.n101 103.111
R6641 CSoutput.n104 CSoutput.n103 103.111
R6642 CSoutput.n106 CSoutput.n105 103.111
R6643 CSoutput.n108 CSoutput.n107 103.111
R6644 CSoutput.n81 CSoutput.n80 103.111
R6645 CSoutput.n83 CSoutput.n82 103.111
R6646 CSoutput.n85 CSoutput.n84 103.111
R6647 CSoutput.n87 CSoutput.n86 103.111
R6648 CSoutput.n89 CSoutput.n88 103.111
R6649 CSoutput.n91 CSoutput.n90 103.111
R6650 CSoutput.n93 CSoutput.n92 103.111
R6651 CSoutput.n322 CSoutput.n321 103.111
R6652 CSoutput.n342 CSoutput.n340 81.5057
R6653 CSoutput.n327 CSoutput.n325 81.5057
R6654 CSoutput.n374 CSoutput.n372 81.5057
R6655 CSoutput.n359 CSoutput.n357 81.5057
R6656 CSoutput.n354 CSoutput.n353 80.9324
R6657 CSoutput.n352 CSoutput.n351 80.9324
R6658 CSoutput.n350 CSoutput.n349 80.9324
R6659 CSoutput.n348 CSoutput.n347 80.9324
R6660 CSoutput.n346 CSoutput.n345 80.9324
R6661 CSoutput.n344 CSoutput.n343 80.9324
R6662 CSoutput.n342 CSoutput.n341 80.9324
R6663 CSoutput.n339 CSoutput.n338 80.9324
R6664 CSoutput.n337 CSoutput.n336 80.9324
R6665 CSoutput.n335 CSoutput.n334 80.9324
R6666 CSoutput.n333 CSoutput.n332 80.9324
R6667 CSoutput.n331 CSoutput.n330 80.9324
R6668 CSoutput.n329 CSoutput.n328 80.9324
R6669 CSoutput.n327 CSoutput.n326 80.9324
R6670 CSoutput.n374 CSoutput.n373 80.9324
R6671 CSoutput.n376 CSoutput.n375 80.9324
R6672 CSoutput.n378 CSoutput.n377 80.9324
R6673 CSoutput.n380 CSoutput.n379 80.9324
R6674 CSoutput.n382 CSoutput.n381 80.9324
R6675 CSoutput.n384 CSoutput.n383 80.9324
R6676 CSoutput.n386 CSoutput.n385 80.9324
R6677 CSoutput.n359 CSoutput.n358 80.9324
R6678 CSoutput.n361 CSoutput.n360 80.9324
R6679 CSoutput.n363 CSoutput.n362 80.9324
R6680 CSoutput.n365 CSoutput.n364 80.9324
R6681 CSoutput.n367 CSoutput.n366 80.9324
R6682 CSoutput.n369 CSoutput.n368 80.9324
R6683 CSoutput.n371 CSoutput.n370 80.9324
R6684 CSoutput.n25 CSoutput.n24 48.1486
R6685 CSoutput.n69 CSoutput.n3 48.1486
R6686 CSoutput.n38 CSoutput.n37 48.1486
R6687 CSoutput.n42 CSoutput.n41 48.1486
R6688 CSoutput.n51 CSoutput.n50 48.1486
R6689 CSoutput.n55 CSoutput.n54 48.1486
R6690 CSoutput.n22 CSoutput.n17 46.462
R6691 CSoutput.n72 CSoutput.n71 46.462
R6692 CSoutput.n20 CSoutput.n19 44.9055
R6693 CSoutput.n29 CSoutput.n28 43.7635
R6694 CSoutput.n65 CSoutput.n63 43.7635
R6695 CSoutput.n35 CSoutput.n13 41.7396
R6696 CSoutput.n57 CSoutput.n5 41.7396
R6697 CSoutput.n44 CSoutput.n9 37.0171
R6698 CSoutput.n48 CSoutput.n9 37.0171
R6699 CSoutput.n76 CSoutput.n75 34.9932
R6700 CSoutput.n31 CSoutput.n13 32.2947
R6701 CSoutput.n61 CSoutput.n5 32.2947
R6702 CSoutput.n30 CSoutput.n29 29.6014
R6703 CSoutput.n63 CSoutput.n62 29.6014
R6704 CSoutput.n19 CSoutput.n18 28.4085
R6705 CSoutput.n18 CSoutput.n17 25.1176
R6706 CSoutput.n72 CSoutput.n1 25.1176
R6707 CSoutput.n43 CSoutput.n42 22.0922
R6708 CSoutput.n50 CSoutput.n49 22.0922
R6709 CSoutput.n77 CSoutput.n76 21.8586
R6710 CSoutput.n37 CSoutput.n36 18.9681
R6711 CSoutput.n56 CSoutput.n55 18.9681
R6712 CSoutput.n25 CSoutput.n15 17.6292
R6713 CSoutput.n64 CSoutput.n3 17.6292
R6714 CSoutput.n24 CSoutput.n23 15.844
R6715 CSoutput.n70 CSoutput.n69 15.844
R6716 CSoutput.n38 CSoutput.n11 14.5051
R6717 CSoutput.n54 CSoutput.n7 14.5051
R6718 CSoutput.n389 CSoutput.n78 11.6139
R6719 CSoutput.n41 CSoutput.n11 11.3811
R6720 CSoutput.n51 CSoutput.n7 11.3811
R6721 CSoutput.n23 CSoutput.n22 10.0422
R6722 CSoutput.n71 CSoutput.n70 10.0422
R6723 CSoutput.n307 CSoutput.n291 9.25285
R6724 CSoutput.n109 CSoutput.n93 9.25285
R6725 CSoutput.n355 CSoutput.n339 8.97993
R6726 CSoutput.n387 CSoutput.n371 8.97993
R6727 CSoutput.n356 CSoutput.n324 8.82395
R6728 CSoutput.n28 CSoutput.n15 8.25698
R6729 CSoutput.n65 CSoutput.n64 8.25698
R6730 CSoutput.n356 CSoutput.n355 7.89345
R6731 CSoutput.n388 CSoutput.n387 7.89345
R6732 CSoutput.n324 CSoutput.n323 7.12641
R6733 CSoutput.n126 CSoutput.n125 7.12641
R6734 CSoutput.n36 CSoutput.n35 6.91809
R6735 CSoutput.n57 CSoutput.n56 6.91809
R6736 CSoutput.n355 CSoutput.n354 5.25266
R6737 CSoutput.n387 CSoutput.n386 5.25266
R6738 CSoutput.n389 CSoutput.n126 5.23151
R6739 CSoutput.n323 CSoutput.n322 5.1449
R6740 CSoutput.n307 CSoutput.n306 5.1449
R6741 CSoutput.n125 CSoutput.n124 5.1449
R6742 CSoutput.n109 CSoutput.n108 5.1449
R6743 CSoutput.n217 CSoutput.n170 4.5005
R6744 CSoutput.n186 CSoutput.n170 4.5005
R6745 CSoutput.n181 CSoutput.n165 4.5005
R6746 CSoutput.n181 CSoutput.n167 4.5005
R6747 CSoutput.n181 CSoutput.n164 4.5005
R6748 CSoutput.n181 CSoutput.n168 4.5005
R6749 CSoutput.n181 CSoutput.n163 4.5005
R6750 CSoutput.n181 CSoutput.t175 4.5005
R6751 CSoutput.n181 CSoutput.n162 4.5005
R6752 CSoutput.n181 CSoutput.n169 4.5005
R6753 CSoutput.n181 CSoutput.n170 4.5005
R6754 CSoutput.n179 CSoutput.n165 4.5005
R6755 CSoutput.n179 CSoutput.n167 4.5005
R6756 CSoutput.n179 CSoutput.n164 4.5005
R6757 CSoutput.n179 CSoutput.n168 4.5005
R6758 CSoutput.n179 CSoutput.n163 4.5005
R6759 CSoutput.n179 CSoutput.t175 4.5005
R6760 CSoutput.n179 CSoutput.n162 4.5005
R6761 CSoutput.n179 CSoutput.n169 4.5005
R6762 CSoutput.n179 CSoutput.n170 4.5005
R6763 CSoutput.n178 CSoutput.n165 4.5005
R6764 CSoutput.n178 CSoutput.n167 4.5005
R6765 CSoutput.n178 CSoutput.n164 4.5005
R6766 CSoutput.n178 CSoutput.n168 4.5005
R6767 CSoutput.n178 CSoutput.n163 4.5005
R6768 CSoutput.n178 CSoutput.t175 4.5005
R6769 CSoutput.n178 CSoutput.n162 4.5005
R6770 CSoutput.n178 CSoutput.n169 4.5005
R6771 CSoutput.n178 CSoutput.n170 4.5005
R6772 CSoutput.n263 CSoutput.n165 4.5005
R6773 CSoutput.n263 CSoutput.n167 4.5005
R6774 CSoutput.n263 CSoutput.n164 4.5005
R6775 CSoutput.n263 CSoutput.n168 4.5005
R6776 CSoutput.n263 CSoutput.n163 4.5005
R6777 CSoutput.n263 CSoutput.t175 4.5005
R6778 CSoutput.n263 CSoutput.n162 4.5005
R6779 CSoutput.n263 CSoutput.n169 4.5005
R6780 CSoutput.n263 CSoutput.n170 4.5005
R6781 CSoutput.n261 CSoutput.n165 4.5005
R6782 CSoutput.n261 CSoutput.n167 4.5005
R6783 CSoutput.n261 CSoutput.n164 4.5005
R6784 CSoutput.n261 CSoutput.n168 4.5005
R6785 CSoutput.n261 CSoutput.n163 4.5005
R6786 CSoutput.n261 CSoutput.t175 4.5005
R6787 CSoutput.n261 CSoutput.n162 4.5005
R6788 CSoutput.n261 CSoutput.n169 4.5005
R6789 CSoutput.n259 CSoutput.n165 4.5005
R6790 CSoutput.n259 CSoutput.n167 4.5005
R6791 CSoutput.n259 CSoutput.n164 4.5005
R6792 CSoutput.n259 CSoutput.n168 4.5005
R6793 CSoutput.n259 CSoutput.n163 4.5005
R6794 CSoutput.n259 CSoutput.t175 4.5005
R6795 CSoutput.n259 CSoutput.n162 4.5005
R6796 CSoutput.n259 CSoutput.n169 4.5005
R6797 CSoutput.n189 CSoutput.n165 4.5005
R6798 CSoutput.n189 CSoutput.n167 4.5005
R6799 CSoutput.n189 CSoutput.n164 4.5005
R6800 CSoutput.n189 CSoutput.n168 4.5005
R6801 CSoutput.n189 CSoutput.n163 4.5005
R6802 CSoutput.n189 CSoutput.t175 4.5005
R6803 CSoutput.n189 CSoutput.n162 4.5005
R6804 CSoutput.n189 CSoutput.n169 4.5005
R6805 CSoutput.n189 CSoutput.n170 4.5005
R6806 CSoutput.n188 CSoutput.n165 4.5005
R6807 CSoutput.n188 CSoutput.n167 4.5005
R6808 CSoutput.n188 CSoutput.n164 4.5005
R6809 CSoutput.n188 CSoutput.n168 4.5005
R6810 CSoutput.n188 CSoutput.n163 4.5005
R6811 CSoutput.n188 CSoutput.t175 4.5005
R6812 CSoutput.n188 CSoutput.n162 4.5005
R6813 CSoutput.n188 CSoutput.n169 4.5005
R6814 CSoutput.n188 CSoutput.n170 4.5005
R6815 CSoutput.n192 CSoutput.n165 4.5005
R6816 CSoutput.n192 CSoutput.n167 4.5005
R6817 CSoutput.n192 CSoutput.n164 4.5005
R6818 CSoutput.n192 CSoutput.n168 4.5005
R6819 CSoutput.n192 CSoutput.n163 4.5005
R6820 CSoutput.n192 CSoutput.t175 4.5005
R6821 CSoutput.n192 CSoutput.n162 4.5005
R6822 CSoutput.n192 CSoutput.n169 4.5005
R6823 CSoutput.n192 CSoutput.n170 4.5005
R6824 CSoutput.n191 CSoutput.n165 4.5005
R6825 CSoutput.n191 CSoutput.n167 4.5005
R6826 CSoutput.n191 CSoutput.n164 4.5005
R6827 CSoutput.n191 CSoutput.n168 4.5005
R6828 CSoutput.n191 CSoutput.n163 4.5005
R6829 CSoutput.n191 CSoutput.t175 4.5005
R6830 CSoutput.n191 CSoutput.n162 4.5005
R6831 CSoutput.n191 CSoutput.n169 4.5005
R6832 CSoutput.n191 CSoutput.n170 4.5005
R6833 CSoutput.n174 CSoutput.n165 4.5005
R6834 CSoutput.n174 CSoutput.n167 4.5005
R6835 CSoutput.n174 CSoutput.n164 4.5005
R6836 CSoutput.n174 CSoutput.n168 4.5005
R6837 CSoutput.n174 CSoutput.n163 4.5005
R6838 CSoutput.n174 CSoutput.t175 4.5005
R6839 CSoutput.n174 CSoutput.n162 4.5005
R6840 CSoutput.n174 CSoutput.n169 4.5005
R6841 CSoutput.n174 CSoutput.n170 4.5005
R6842 CSoutput.n266 CSoutput.n165 4.5005
R6843 CSoutput.n266 CSoutput.n167 4.5005
R6844 CSoutput.n266 CSoutput.n164 4.5005
R6845 CSoutput.n266 CSoutput.n168 4.5005
R6846 CSoutput.n266 CSoutput.n163 4.5005
R6847 CSoutput.n266 CSoutput.t175 4.5005
R6848 CSoutput.n266 CSoutput.n162 4.5005
R6849 CSoutput.n266 CSoutput.n169 4.5005
R6850 CSoutput.n266 CSoutput.n170 4.5005
R6851 CSoutput.n253 CSoutput.n224 4.5005
R6852 CSoutput.n253 CSoutput.n230 4.5005
R6853 CSoutput.n211 CSoutput.n200 4.5005
R6854 CSoutput.n211 CSoutput.n202 4.5005
R6855 CSoutput.n211 CSoutput.n199 4.5005
R6856 CSoutput.n211 CSoutput.n203 4.5005
R6857 CSoutput.n211 CSoutput.n198 4.5005
R6858 CSoutput.n211 CSoutput.t171 4.5005
R6859 CSoutput.n211 CSoutput.n197 4.5005
R6860 CSoutput.n211 CSoutput.n204 4.5005
R6861 CSoutput.n253 CSoutput.n211 4.5005
R6862 CSoutput.n232 CSoutput.n200 4.5005
R6863 CSoutput.n232 CSoutput.n202 4.5005
R6864 CSoutput.n232 CSoutput.n199 4.5005
R6865 CSoutput.n232 CSoutput.n203 4.5005
R6866 CSoutput.n232 CSoutput.n198 4.5005
R6867 CSoutput.n232 CSoutput.t171 4.5005
R6868 CSoutput.n232 CSoutput.n197 4.5005
R6869 CSoutput.n232 CSoutput.n204 4.5005
R6870 CSoutput.n253 CSoutput.n232 4.5005
R6871 CSoutput.n210 CSoutput.n200 4.5005
R6872 CSoutput.n210 CSoutput.n202 4.5005
R6873 CSoutput.n210 CSoutput.n199 4.5005
R6874 CSoutput.n210 CSoutput.n203 4.5005
R6875 CSoutput.n210 CSoutput.n198 4.5005
R6876 CSoutput.n210 CSoutput.t171 4.5005
R6877 CSoutput.n210 CSoutput.n197 4.5005
R6878 CSoutput.n210 CSoutput.n204 4.5005
R6879 CSoutput.n253 CSoutput.n210 4.5005
R6880 CSoutput.n234 CSoutput.n200 4.5005
R6881 CSoutput.n234 CSoutput.n202 4.5005
R6882 CSoutput.n234 CSoutput.n199 4.5005
R6883 CSoutput.n234 CSoutput.n203 4.5005
R6884 CSoutput.n234 CSoutput.n198 4.5005
R6885 CSoutput.n234 CSoutput.t171 4.5005
R6886 CSoutput.n234 CSoutput.n197 4.5005
R6887 CSoutput.n234 CSoutput.n204 4.5005
R6888 CSoutput.n253 CSoutput.n234 4.5005
R6889 CSoutput.n200 CSoutput.n195 4.5005
R6890 CSoutput.n202 CSoutput.n195 4.5005
R6891 CSoutput.n199 CSoutput.n195 4.5005
R6892 CSoutput.n203 CSoutput.n195 4.5005
R6893 CSoutput.n198 CSoutput.n195 4.5005
R6894 CSoutput.t171 CSoutput.n195 4.5005
R6895 CSoutput.n197 CSoutput.n195 4.5005
R6896 CSoutput.n204 CSoutput.n195 4.5005
R6897 CSoutput.n256 CSoutput.n200 4.5005
R6898 CSoutput.n256 CSoutput.n202 4.5005
R6899 CSoutput.n256 CSoutput.n199 4.5005
R6900 CSoutput.n256 CSoutput.n203 4.5005
R6901 CSoutput.n256 CSoutput.n198 4.5005
R6902 CSoutput.n256 CSoutput.t171 4.5005
R6903 CSoutput.n256 CSoutput.n197 4.5005
R6904 CSoutput.n256 CSoutput.n204 4.5005
R6905 CSoutput.n254 CSoutput.n200 4.5005
R6906 CSoutput.n254 CSoutput.n202 4.5005
R6907 CSoutput.n254 CSoutput.n199 4.5005
R6908 CSoutput.n254 CSoutput.n203 4.5005
R6909 CSoutput.n254 CSoutput.n198 4.5005
R6910 CSoutput.n254 CSoutput.t171 4.5005
R6911 CSoutput.n254 CSoutput.n197 4.5005
R6912 CSoutput.n254 CSoutput.n204 4.5005
R6913 CSoutput.n254 CSoutput.n253 4.5005
R6914 CSoutput.n236 CSoutput.n200 4.5005
R6915 CSoutput.n236 CSoutput.n202 4.5005
R6916 CSoutput.n236 CSoutput.n199 4.5005
R6917 CSoutput.n236 CSoutput.n203 4.5005
R6918 CSoutput.n236 CSoutput.n198 4.5005
R6919 CSoutput.n236 CSoutput.t171 4.5005
R6920 CSoutput.n236 CSoutput.n197 4.5005
R6921 CSoutput.n236 CSoutput.n204 4.5005
R6922 CSoutput.n253 CSoutput.n236 4.5005
R6923 CSoutput.n208 CSoutput.n200 4.5005
R6924 CSoutput.n208 CSoutput.n202 4.5005
R6925 CSoutput.n208 CSoutput.n199 4.5005
R6926 CSoutput.n208 CSoutput.n203 4.5005
R6927 CSoutput.n208 CSoutput.n198 4.5005
R6928 CSoutput.n208 CSoutput.t171 4.5005
R6929 CSoutput.n208 CSoutput.n197 4.5005
R6930 CSoutput.n208 CSoutput.n204 4.5005
R6931 CSoutput.n253 CSoutput.n208 4.5005
R6932 CSoutput.n238 CSoutput.n200 4.5005
R6933 CSoutput.n238 CSoutput.n202 4.5005
R6934 CSoutput.n238 CSoutput.n199 4.5005
R6935 CSoutput.n238 CSoutput.n203 4.5005
R6936 CSoutput.n238 CSoutput.n198 4.5005
R6937 CSoutput.n238 CSoutput.t171 4.5005
R6938 CSoutput.n238 CSoutput.n197 4.5005
R6939 CSoutput.n238 CSoutput.n204 4.5005
R6940 CSoutput.n253 CSoutput.n238 4.5005
R6941 CSoutput.n207 CSoutput.n200 4.5005
R6942 CSoutput.n207 CSoutput.n202 4.5005
R6943 CSoutput.n207 CSoutput.n199 4.5005
R6944 CSoutput.n207 CSoutput.n203 4.5005
R6945 CSoutput.n207 CSoutput.n198 4.5005
R6946 CSoutput.n207 CSoutput.t171 4.5005
R6947 CSoutput.n207 CSoutput.n197 4.5005
R6948 CSoutput.n207 CSoutput.n204 4.5005
R6949 CSoutput.n253 CSoutput.n207 4.5005
R6950 CSoutput.n252 CSoutput.n200 4.5005
R6951 CSoutput.n252 CSoutput.n202 4.5005
R6952 CSoutput.n252 CSoutput.n199 4.5005
R6953 CSoutput.n252 CSoutput.n203 4.5005
R6954 CSoutput.n252 CSoutput.n198 4.5005
R6955 CSoutput.n252 CSoutput.t171 4.5005
R6956 CSoutput.n252 CSoutput.n197 4.5005
R6957 CSoutput.n252 CSoutput.n204 4.5005
R6958 CSoutput.n253 CSoutput.n252 4.5005
R6959 CSoutput.n251 CSoutput.n136 4.5005
R6960 CSoutput.n152 CSoutput.n136 4.5005
R6961 CSoutput.n147 CSoutput.n131 4.5005
R6962 CSoutput.n147 CSoutput.n133 4.5005
R6963 CSoutput.n147 CSoutput.n130 4.5005
R6964 CSoutput.n147 CSoutput.n134 4.5005
R6965 CSoutput.n147 CSoutput.n129 4.5005
R6966 CSoutput.n147 CSoutput.t161 4.5005
R6967 CSoutput.n147 CSoutput.n128 4.5005
R6968 CSoutput.n147 CSoutput.n135 4.5005
R6969 CSoutput.n147 CSoutput.n136 4.5005
R6970 CSoutput.n145 CSoutput.n131 4.5005
R6971 CSoutput.n145 CSoutput.n133 4.5005
R6972 CSoutput.n145 CSoutput.n130 4.5005
R6973 CSoutput.n145 CSoutput.n134 4.5005
R6974 CSoutput.n145 CSoutput.n129 4.5005
R6975 CSoutput.n145 CSoutput.t161 4.5005
R6976 CSoutput.n145 CSoutput.n128 4.5005
R6977 CSoutput.n145 CSoutput.n135 4.5005
R6978 CSoutput.n145 CSoutput.n136 4.5005
R6979 CSoutput.n144 CSoutput.n131 4.5005
R6980 CSoutput.n144 CSoutput.n133 4.5005
R6981 CSoutput.n144 CSoutput.n130 4.5005
R6982 CSoutput.n144 CSoutput.n134 4.5005
R6983 CSoutput.n144 CSoutput.n129 4.5005
R6984 CSoutput.n144 CSoutput.t161 4.5005
R6985 CSoutput.n144 CSoutput.n128 4.5005
R6986 CSoutput.n144 CSoutput.n135 4.5005
R6987 CSoutput.n144 CSoutput.n136 4.5005
R6988 CSoutput.n273 CSoutput.n131 4.5005
R6989 CSoutput.n273 CSoutput.n133 4.5005
R6990 CSoutput.n273 CSoutput.n130 4.5005
R6991 CSoutput.n273 CSoutput.n134 4.5005
R6992 CSoutput.n273 CSoutput.n129 4.5005
R6993 CSoutput.n273 CSoutput.t161 4.5005
R6994 CSoutput.n273 CSoutput.n128 4.5005
R6995 CSoutput.n273 CSoutput.n135 4.5005
R6996 CSoutput.n273 CSoutput.n136 4.5005
R6997 CSoutput.n271 CSoutput.n131 4.5005
R6998 CSoutput.n271 CSoutput.n133 4.5005
R6999 CSoutput.n271 CSoutput.n130 4.5005
R7000 CSoutput.n271 CSoutput.n134 4.5005
R7001 CSoutput.n271 CSoutput.n129 4.5005
R7002 CSoutput.n271 CSoutput.t161 4.5005
R7003 CSoutput.n271 CSoutput.n128 4.5005
R7004 CSoutput.n271 CSoutput.n135 4.5005
R7005 CSoutput.n269 CSoutput.n131 4.5005
R7006 CSoutput.n269 CSoutput.n133 4.5005
R7007 CSoutput.n269 CSoutput.n130 4.5005
R7008 CSoutput.n269 CSoutput.n134 4.5005
R7009 CSoutput.n269 CSoutput.n129 4.5005
R7010 CSoutput.n269 CSoutput.t161 4.5005
R7011 CSoutput.n269 CSoutput.n128 4.5005
R7012 CSoutput.n269 CSoutput.n135 4.5005
R7013 CSoutput.n155 CSoutput.n131 4.5005
R7014 CSoutput.n155 CSoutput.n133 4.5005
R7015 CSoutput.n155 CSoutput.n130 4.5005
R7016 CSoutput.n155 CSoutput.n134 4.5005
R7017 CSoutput.n155 CSoutput.n129 4.5005
R7018 CSoutput.n155 CSoutput.t161 4.5005
R7019 CSoutput.n155 CSoutput.n128 4.5005
R7020 CSoutput.n155 CSoutput.n135 4.5005
R7021 CSoutput.n155 CSoutput.n136 4.5005
R7022 CSoutput.n154 CSoutput.n131 4.5005
R7023 CSoutput.n154 CSoutput.n133 4.5005
R7024 CSoutput.n154 CSoutput.n130 4.5005
R7025 CSoutput.n154 CSoutput.n134 4.5005
R7026 CSoutput.n154 CSoutput.n129 4.5005
R7027 CSoutput.n154 CSoutput.t161 4.5005
R7028 CSoutput.n154 CSoutput.n128 4.5005
R7029 CSoutput.n154 CSoutput.n135 4.5005
R7030 CSoutput.n154 CSoutput.n136 4.5005
R7031 CSoutput.n158 CSoutput.n131 4.5005
R7032 CSoutput.n158 CSoutput.n133 4.5005
R7033 CSoutput.n158 CSoutput.n130 4.5005
R7034 CSoutput.n158 CSoutput.n134 4.5005
R7035 CSoutput.n158 CSoutput.n129 4.5005
R7036 CSoutput.n158 CSoutput.t161 4.5005
R7037 CSoutput.n158 CSoutput.n128 4.5005
R7038 CSoutput.n158 CSoutput.n135 4.5005
R7039 CSoutput.n158 CSoutput.n136 4.5005
R7040 CSoutput.n157 CSoutput.n131 4.5005
R7041 CSoutput.n157 CSoutput.n133 4.5005
R7042 CSoutput.n157 CSoutput.n130 4.5005
R7043 CSoutput.n157 CSoutput.n134 4.5005
R7044 CSoutput.n157 CSoutput.n129 4.5005
R7045 CSoutput.n157 CSoutput.t161 4.5005
R7046 CSoutput.n157 CSoutput.n128 4.5005
R7047 CSoutput.n157 CSoutput.n135 4.5005
R7048 CSoutput.n157 CSoutput.n136 4.5005
R7049 CSoutput.n140 CSoutput.n131 4.5005
R7050 CSoutput.n140 CSoutput.n133 4.5005
R7051 CSoutput.n140 CSoutput.n130 4.5005
R7052 CSoutput.n140 CSoutput.n134 4.5005
R7053 CSoutput.n140 CSoutput.n129 4.5005
R7054 CSoutput.n140 CSoutput.t161 4.5005
R7055 CSoutput.n140 CSoutput.n128 4.5005
R7056 CSoutput.n140 CSoutput.n135 4.5005
R7057 CSoutput.n140 CSoutput.n136 4.5005
R7058 CSoutput.n276 CSoutput.n131 4.5005
R7059 CSoutput.n276 CSoutput.n133 4.5005
R7060 CSoutput.n276 CSoutput.n130 4.5005
R7061 CSoutput.n276 CSoutput.n134 4.5005
R7062 CSoutput.n276 CSoutput.n129 4.5005
R7063 CSoutput.n276 CSoutput.t161 4.5005
R7064 CSoutput.n276 CSoutput.n128 4.5005
R7065 CSoutput.n276 CSoutput.n135 4.5005
R7066 CSoutput.n276 CSoutput.n136 4.5005
R7067 CSoutput.n323 CSoutput.n307 4.10845
R7068 CSoutput.n125 CSoutput.n109 4.10845
R7069 CSoutput.n321 CSoutput.t123 4.06363
R7070 CSoutput.n321 CSoutput.t56 4.06363
R7071 CSoutput.n319 CSoutput.t50 4.06363
R7072 CSoutput.n319 CSoutput.t92 4.06363
R7073 CSoutput.n317 CSoutput.t105 4.06363
R7074 CSoutput.n317 CSoutput.t125 4.06363
R7075 CSoutput.n315 CSoutput.t136 4.06363
R7076 CSoutput.n315 CSoutput.t67 4.06363
R7077 CSoutput.n313 CSoutput.t71 4.06363
R7078 CSoutput.n313 CSoutput.t126 4.06363
R7079 CSoutput.n311 CSoutput.t138 4.06363
R7080 CSoutput.n311 CSoutput.t139 4.06363
R7081 CSoutput.n309 CSoutput.t89 4.06363
R7082 CSoutput.n309 CSoutput.t90 4.06363
R7083 CSoutput.n308 CSoutput.t93 4.06363
R7084 CSoutput.n308 CSoutput.t140 4.06363
R7085 CSoutput.n305 CSoutput.t114 4.06363
R7086 CSoutput.n305 CSoutput.t141 4.06363
R7087 CSoutput.n303 CSoutput.t137 4.06363
R7088 CSoutput.n303 CSoutput.t79 4.06363
R7089 CSoutput.n301 CSoutput.t95 4.06363
R7090 CSoutput.n301 CSoutput.t115 4.06363
R7091 CSoutput.n299 CSoutput.t127 4.06363
R7092 CSoutput.n299 CSoutput.t55 4.06363
R7093 CSoutput.n297 CSoutput.t57 4.06363
R7094 CSoutput.n297 CSoutput.t118 4.06363
R7095 CSoutput.n295 CSoutput.t130 4.06363
R7096 CSoutput.n295 CSoutput.t131 4.06363
R7097 CSoutput.n293 CSoutput.t73 4.06363
R7098 CSoutput.n293 CSoutput.t74 4.06363
R7099 CSoutput.n292 CSoutput.t80 4.06363
R7100 CSoutput.n292 CSoutput.t132 4.06363
R7101 CSoutput.n290 CSoutput.t116 4.06363
R7102 CSoutput.n290 CSoutput.t77 4.06363
R7103 CSoutput.n288 CSoutput.t133 4.06363
R7104 CSoutput.n288 CSoutput.t99 4.06363
R7105 CSoutput.n286 CSoutput.t124 4.06363
R7106 CSoutput.n286 CSoutput.t86 4.06363
R7107 CSoutput.n284 CSoutput.t111 4.06363
R7108 CSoutput.n284 CSoutput.t66 4.06363
R7109 CSoutput.n282 CSoutput.t128 4.06363
R7110 CSoutput.n282 CSoutput.t61 4.06363
R7111 CSoutput.n280 CSoutput.t96 4.06363
R7112 CSoutput.n280 CSoutput.t75 4.06363
R7113 CSoutput.n278 CSoutput.t81 4.06363
R7114 CSoutput.n278 CSoutput.t58 4.06363
R7115 CSoutput.n277 CSoutput.t122 4.06363
R7116 CSoutput.n277 CSoutput.t52 4.06363
R7117 CSoutput.n110 CSoutput.t88 4.06363
R7118 CSoutput.n110 CSoutput.t143 4.06363
R7119 CSoutput.n111 CSoutput.t120 4.06363
R7120 CSoutput.n111 CSoutput.t119 4.06363
R7121 CSoutput.n113 CSoutput.t107 4.06363
R7122 CSoutput.n113 CSoutput.t85 4.06363
R7123 CSoutput.n115 CSoutput.t65 4.06363
R7124 CSoutput.n115 CSoutput.t108 4.06363
R7125 CSoutput.n117 CSoutput.t106 4.06363
R7126 CSoutput.n117 CSoutput.t82 4.06363
R7127 CSoutput.n119 CSoutput.t64 4.06363
R7128 CSoutput.n119 CSoutput.t63 4.06363
R7129 CSoutput.n121 CSoutput.t121 4.06363
R7130 CSoutput.n121 CSoutput.t94 4.06363
R7131 CSoutput.n123 CSoutput.t91 4.06363
R7132 CSoutput.n123 CSoutput.t59 4.06363
R7133 CSoutput.n94 CSoutput.t72 4.06363
R7134 CSoutput.n94 CSoutput.t135 4.06363
R7135 CSoutput.n95 CSoutput.t110 4.06363
R7136 CSoutput.n95 CSoutput.t109 4.06363
R7137 CSoutput.n97 CSoutput.t101 4.06363
R7138 CSoutput.n97 CSoutput.t70 4.06363
R7139 CSoutput.n99 CSoutput.t53 4.06363
R7140 CSoutput.n99 CSoutput.t102 4.06363
R7141 CSoutput.n101 CSoutput.t98 4.06363
R7142 CSoutput.n101 CSoutput.t68 4.06363
R7143 CSoutput.n103 CSoutput.t51 4.06363
R7144 CSoutput.n103 CSoutput.t49 4.06363
R7145 CSoutput.n105 CSoutput.t113 4.06363
R7146 CSoutput.n105 CSoutput.t84 4.06363
R7147 CSoutput.n107 CSoutput.t78 4.06363
R7148 CSoutput.n107 CSoutput.t48 4.06363
R7149 CSoutput.n79 CSoutput.t54 4.06363
R7150 CSoutput.n79 CSoutput.t103 4.06363
R7151 CSoutput.n80 CSoutput.t60 4.06363
R7152 CSoutput.n80 CSoutput.t83 4.06363
R7153 CSoutput.n82 CSoutput.t142 4.06363
R7154 CSoutput.n82 CSoutput.t97 4.06363
R7155 CSoutput.n84 CSoutput.t62 4.06363
R7156 CSoutput.n84 CSoutput.t129 4.06363
R7157 CSoutput.n86 CSoutput.t69 4.06363
R7158 CSoutput.n86 CSoutput.t112 4.06363
R7159 CSoutput.n88 CSoutput.t87 4.06363
R7160 CSoutput.n88 CSoutput.t104 4.06363
R7161 CSoutput.n90 CSoutput.t100 4.06363
R7162 CSoutput.n90 CSoutput.t134 4.06363
R7163 CSoutput.n92 CSoutput.t76 4.06363
R7164 CSoutput.n92 CSoutput.t117 4.06363
R7165 CSoutput.n44 CSoutput.n43 3.79402
R7166 CSoutput.n49 CSoutput.n48 3.79402
R7167 CSoutput.n389 CSoutput.n388 3.57343
R7168 CSoutput.n388 CSoutput.n356 3.3798
R7169 CSoutput.n353 CSoutput.t29 2.82907
R7170 CSoutput.n353 CSoutput.t42 2.82907
R7171 CSoutput.n351 CSoutput.t145 2.82907
R7172 CSoutput.n351 CSoutput.t45 2.82907
R7173 CSoutput.n349 CSoutput.t28 2.82907
R7174 CSoutput.n349 CSoutput.t21 2.82907
R7175 CSoutput.n347 CSoutput.t35 2.82907
R7176 CSoutput.n347 CSoutput.t17 2.82907
R7177 CSoutput.n345 CSoutput.t159 2.82907
R7178 CSoutput.n345 CSoutput.t18 2.82907
R7179 CSoutput.n343 CSoutput.t33 2.82907
R7180 CSoutput.n343 CSoutput.t37 2.82907
R7181 CSoutput.n341 CSoutput.t32 2.82907
R7182 CSoutput.n341 CSoutput.t13 2.82907
R7183 CSoutput.n340 CSoutput.t144 2.82907
R7184 CSoutput.n340 CSoutput.t36 2.82907
R7185 CSoutput.n338 CSoutput.t0 2.82907
R7186 CSoutput.n338 CSoutput.t20 2.82907
R7187 CSoutput.n336 CSoutput.t44 2.82907
R7188 CSoutput.n336 CSoutput.t10 2.82907
R7189 CSoutput.n334 CSoutput.t153 2.82907
R7190 CSoutput.n334 CSoutput.t16 2.82907
R7191 CSoutput.n332 CSoutput.t46 2.82907
R7192 CSoutput.n332 CSoutput.t152 2.82907
R7193 CSoutput.n330 CSoutput.t15 2.82907
R7194 CSoutput.n330 CSoutput.t43 2.82907
R7195 CSoutput.n328 CSoutput.t8 2.82907
R7196 CSoutput.n328 CSoutput.t150 2.82907
R7197 CSoutput.n326 CSoutput.t27 2.82907
R7198 CSoutput.n326 CSoutput.t147 2.82907
R7199 CSoutput.n325 CSoutput.t7 2.82907
R7200 CSoutput.n325 CSoutput.t25 2.82907
R7201 CSoutput.n372 CSoutput.t22 2.82907
R7202 CSoutput.n372 CSoutput.t24 2.82907
R7203 CSoutput.n373 CSoutput.t34 2.82907
R7204 CSoutput.n373 CSoutput.t11 2.82907
R7205 CSoutput.n375 CSoutput.t39 2.82907
R7206 CSoutput.n375 CSoutput.t38 2.82907
R7207 CSoutput.n377 CSoutput.t14 2.82907
R7208 CSoutput.n377 CSoutput.t4 2.82907
R7209 CSoutput.n379 CSoutput.t41 2.82907
R7210 CSoutput.n379 CSoutput.t23 2.82907
R7211 CSoutput.n381 CSoutput.t9 2.82907
R7212 CSoutput.n381 CSoutput.t157 2.82907
R7213 CSoutput.n383 CSoutput.t26 2.82907
R7214 CSoutput.n383 CSoutput.t31 2.82907
R7215 CSoutput.n385 CSoutput.t30 2.82907
R7216 CSoutput.n385 CSoutput.t12 2.82907
R7217 CSoutput.n357 CSoutput.t3 2.82907
R7218 CSoutput.n357 CSoutput.t148 2.82907
R7219 CSoutput.n358 CSoutput.t2 2.82907
R7220 CSoutput.n358 CSoutput.t19 2.82907
R7221 CSoutput.n360 CSoutput.t149 2.82907
R7222 CSoutput.n360 CSoutput.t151 2.82907
R7223 CSoutput.n362 CSoutput.t1 2.82907
R7224 CSoutput.n362 CSoutput.t154 2.82907
R7225 CSoutput.n364 CSoutput.t158 2.82907
R7226 CSoutput.n364 CSoutput.t40 2.82907
R7227 CSoutput.n366 CSoutput.t156 2.82907
R7228 CSoutput.n366 CSoutput.t5 2.82907
R7229 CSoutput.n368 CSoutput.t47 2.82907
R7230 CSoutput.n368 CSoutput.t155 2.82907
R7231 CSoutput.n370 CSoutput.t6 2.82907
R7232 CSoutput.n370 CSoutput.t146 2.82907
R7233 CSoutput.n324 CSoutput.n126 2.78353
R7234 CSoutput.n75 CSoutput.n1 2.45513
R7235 CSoutput.n217 CSoutput.n215 2.251
R7236 CSoutput.n217 CSoutput.n214 2.251
R7237 CSoutput.n217 CSoutput.n213 2.251
R7238 CSoutput.n217 CSoutput.n212 2.251
R7239 CSoutput.n186 CSoutput.n185 2.251
R7240 CSoutput.n186 CSoutput.n184 2.251
R7241 CSoutput.n186 CSoutput.n183 2.251
R7242 CSoutput.n186 CSoutput.n182 2.251
R7243 CSoutput.n259 CSoutput.n258 2.251
R7244 CSoutput.n224 CSoutput.n222 2.251
R7245 CSoutput.n224 CSoutput.n221 2.251
R7246 CSoutput.n224 CSoutput.n220 2.251
R7247 CSoutput.n242 CSoutput.n224 2.251
R7248 CSoutput.n230 CSoutput.n229 2.251
R7249 CSoutput.n230 CSoutput.n228 2.251
R7250 CSoutput.n230 CSoutput.n227 2.251
R7251 CSoutput.n230 CSoutput.n226 2.251
R7252 CSoutput.n256 CSoutput.n196 2.251
R7253 CSoutput.n251 CSoutput.n249 2.251
R7254 CSoutput.n251 CSoutput.n248 2.251
R7255 CSoutput.n251 CSoutput.n247 2.251
R7256 CSoutput.n251 CSoutput.n246 2.251
R7257 CSoutput.n152 CSoutput.n151 2.251
R7258 CSoutput.n152 CSoutput.n150 2.251
R7259 CSoutput.n152 CSoutput.n149 2.251
R7260 CSoutput.n152 CSoutput.n148 2.251
R7261 CSoutput.n269 CSoutput.n268 2.251
R7262 CSoutput.n186 CSoutput.n166 2.2505
R7263 CSoutput.n181 CSoutput.n166 2.2505
R7264 CSoutput.n179 CSoutput.n166 2.2505
R7265 CSoutput.n178 CSoutput.n166 2.2505
R7266 CSoutput.n263 CSoutput.n166 2.2505
R7267 CSoutput.n261 CSoutput.n166 2.2505
R7268 CSoutput.n259 CSoutput.n166 2.2505
R7269 CSoutput.n189 CSoutput.n166 2.2505
R7270 CSoutput.n188 CSoutput.n166 2.2505
R7271 CSoutput.n192 CSoutput.n166 2.2505
R7272 CSoutput.n191 CSoutput.n166 2.2505
R7273 CSoutput.n174 CSoutput.n166 2.2505
R7274 CSoutput.n266 CSoutput.n166 2.2505
R7275 CSoutput.n266 CSoutput.n265 2.2505
R7276 CSoutput.n230 CSoutput.n201 2.2505
R7277 CSoutput.n211 CSoutput.n201 2.2505
R7278 CSoutput.n232 CSoutput.n201 2.2505
R7279 CSoutput.n210 CSoutput.n201 2.2505
R7280 CSoutput.n234 CSoutput.n201 2.2505
R7281 CSoutput.n201 CSoutput.n195 2.2505
R7282 CSoutput.n256 CSoutput.n201 2.2505
R7283 CSoutput.n254 CSoutput.n201 2.2505
R7284 CSoutput.n236 CSoutput.n201 2.2505
R7285 CSoutput.n208 CSoutput.n201 2.2505
R7286 CSoutput.n238 CSoutput.n201 2.2505
R7287 CSoutput.n207 CSoutput.n201 2.2505
R7288 CSoutput.n252 CSoutput.n201 2.2505
R7289 CSoutput.n252 CSoutput.n205 2.2505
R7290 CSoutput.n152 CSoutput.n132 2.2505
R7291 CSoutput.n147 CSoutput.n132 2.2505
R7292 CSoutput.n145 CSoutput.n132 2.2505
R7293 CSoutput.n144 CSoutput.n132 2.2505
R7294 CSoutput.n273 CSoutput.n132 2.2505
R7295 CSoutput.n271 CSoutput.n132 2.2505
R7296 CSoutput.n269 CSoutput.n132 2.2505
R7297 CSoutput.n155 CSoutput.n132 2.2505
R7298 CSoutput.n154 CSoutput.n132 2.2505
R7299 CSoutput.n158 CSoutput.n132 2.2505
R7300 CSoutput.n157 CSoutput.n132 2.2505
R7301 CSoutput.n140 CSoutput.n132 2.2505
R7302 CSoutput.n276 CSoutput.n132 2.2505
R7303 CSoutput.n276 CSoutput.n275 2.2505
R7304 CSoutput.n194 CSoutput.n187 2.25024
R7305 CSoutput.n194 CSoutput.n180 2.25024
R7306 CSoutput.n262 CSoutput.n194 2.25024
R7307 CSoutput.n194 CSoutput.n190 2.25024
R7308 CSoutput.n194 CSoutput.n193 2.25024
R7309 CSoutput.n194 CSoutput.n161 2.25024
R7310 CSoutput.n244 CSoutput.n241 2.25024
R7311 CSoutput.n244 CSoutput.n240 2.25024
R7312 CSoutput.n244 CSoutput.n239 2.25024
R7313 CSoutput.n244 CSoutput.n206 2.25024
R7314 CSoutput.n244 CSoutput.n243 2.25024
R7315 CSoutput.n245 CSoutput.n244 2.25024
R7316 CSoutput.n160 CSoutput.n153 2.25024
R7317 CSoutput.n160 CSoutput.n146 2.25024
R7318 CSoutput.n272 CSoutput.n160 2.25024
R7319 CSoutput.n160 CSoutput.n156 2.25024
R7320 CSoutput.n160 CSoutput.n159 2.25024
R7321 CSoutput.n160 CSoutput.n127 2.25024
R7322 CSoutput.n261 CSoutput.n171 1.50111
R7323 CSoutput.n209 CSoutput.n195 1.50111
R7324 CSoutput.n271 CSoutput.n137 1.50111
R7325 CSoutput.n217 CSoutput.n216 1.501
R7326 CSoutput.n224 CSoutput.n223 1.501
R7327 CSoutput.n251 CSoutput.n250 1.501
R7328 CSoutput.n265 CSoutput.n176 1.12536
R7329 CSoutput.n265 CSoutput.n177 1.12536
R7330 CSoutput.n265 CSoutput.n264 1.12536
R7331 CSoutput.n225 CSoutput.n205 1.12536
R7332 CSoutput.n231 CSoutput.n205 1.12536
R7333 CSoutput.n233 CSoutput.n205 1.12536
R7334 CSoutput.n275 CSoutput.n142 1.12536
R7335 CSoutput.n275 CSoutput.n143 1.12536
R7336 CSoutput.n275 CSoutput.n274 1.12536
R7337 CSoutput.n265 CSoutput.n172 1.12536
R7338 CSoutput.n265 CSoutput.n173 1.12536
R7339 CSoutput.n265 CSoutput.n175 1.12536
R7340 CSoutput.n255 CSoutput.n205 1.12536
R7341 CSoutput.n235 CSoutput.n205 1.12536
R7342 CSoutput.n237 CSoutput.n205 1.12536
R7343 CSoutput.n275 CSoutput.n138 1.12536
R7344 CSoutput.n275 CSoutput.n139 1.12536
R7345 CSoutput.n275 CSoutput.n141 1.12536
R7346 CSoutput.n31 CSoutput.n30 0.669944
R7347 CSoutput.n62 CSoutput.n61 0.669944
R7348 CSoutput.n344 CSoutput.n342 0.573776
R7349 CSoutput.n346 CSoutput.n344 0.573776
R7350 CSoutput.n348 CSoutput.n346 0.573776
R7351 CSoutput.n350 CSoutput.n348 0.573776
R7352 CSoutput.n352 CSoutput.n350 0.573776
R7353 CSoutput.n354 CSoutput.n352 0.573776
R7354 CSoutput.n329 CSoutput.n327 0.573776
R7355 CSoutput.n331 CSoutput.n329 0.573776
R7356 CSoutput.n333 CSoutput.n331 0.573776
R7357 CSoutput.n335 CSoutput.n333 0.573776
R7358 CSoutput.n337 CSoutput.n335 0.573776
R7359 CSoutput.n339 CSoutput.n337 0.573776
R7360 CSoutput.n386 CSoutput.n384 0.573776
R7361 CSoutput.n384 CSoutput.n382 0.573776
R7362 CSoutput.n382 CSoutput.n380 0.573776
R7363 CSoutput.n380 CSoutput.n378 0.573776
R7364 CSoutput.n378 CSoutput.n376 0.573776
R7365 CSoutput.n376 CSoutput.n374 0.573776
R7366 CSoutput.n371 CSoutput.n369 0.573776
R7367 CSoutput.n369 CSoutput.n367 0.573776
R7368 CSoutput.n367 CSoutput.n365 0.573776
R7369 CSoutput.n365 CSoutput.n363 0.573776
R7370 CSoutput.n363 CSoutput.n361 0.573776
R7371 CSoutput.n361 CSoutput.n359 0.573776
R7372 CSoutput.n389 CSoutput.n276 0.53442
R7373 CSoutput.n312 CSoutput.n310 0.358259
R7374 CSoutput.n314 CSoutput.n312 0.358259
R7375 CSoutput.n316 CSoutput.n314 0.358259
R7376 CSoutput.n318 CSoutput.n316 0.358259
R7377 CSoutput.n320 CSoutput.n318 0.358259
R7378 CSoutput.n322 CSoutput.n320 0.358259
R7379 CSoutput.n296 CSoutput.n294 0.358259
R7380 CSoutput.n298 CSoutput.n296 0.358259
R7381 CSoutput.n300 CSoutput.n298 0.358259
R7382 CSoutput.n302 CSoutput.n300 0.358259
R7383 CSoutput.n304 CSoutput.n302 0.358259
R7384 CSoutput.n306 CSoutput.n304 0.358259
R7385 CSoutput.n281 CSoutput.n279 0.358259
R7386 CSoutput.n283 CSoutput.n281 0.358259
R7387 CSoutput.n285 CSoutput.n283 0.358259
R7388 CSoutput.n287 CSoutput.n285 0.358259
R7389 CSoutput.n289 CSoutput.n287 0.358259
R7390 CSoutput.n291 CSoutput.n289 0.358259
R7391 CSoutput.n124 CSoutput.n122 0.358259
R7392 CSoutput.n122 CSoutput.n120 0.358259
R7393 CSoutput.n120 CSoutput.n118 0.358259
R7394 CSoutput.n118 CSoutput.n116 0.358259
R7395 CSoutput.n116 CSoutput.n114 0.358259
R7396 CSoutput.n114 CSoutput.n112 0.358259
R7397 CSoutput.n108 CSoutput.n106 0.358259
R7398 CSoutput.n106 CSoutput.n104 0.358259
R7399 CSoutput.n104 CSoutput.n102 0.358259
R7400 CSoutput.n102 CSoutput.n100 0.358259
R7401 CSoutput.n100 CSoutput.n98 0.358259
R7402 CSoutput.n98 CSoutput.n96 0.358259
R7403 CSoutput.n93 CSoutput.n91 0.358259
R7404 CSoutput.n91 CSoutput.n89 0.358259
R7405 CSoutput.n89 CSoutput.n87 0.358259
R7406 CSoutput.n87 CSoutput.n85 0.358259
R7407 CSoutput.n85 CSoutput.n83 0.358259
R7408 CSoutput.n83 CSoutput.n81 0.358259
R7409 CSoutput.n21 CSoutput.n20 0.169105
R7410 CSoutput.n21 CSoutput.n16 0.169105
R7411 CSoutput.n26 CSoutput.n16 0.169105
R7412 CSoutput.n27 CSoutput.n26 0.169105
R7413 CSoutput.n27 CSoutput.n14 0.169105
R7414 CSoutput.n32 CSoutput.n14 0.169105
R7415 CSoutput.n33 CSoutput.n32 0.169105
R7416 CSoutput.n34 CSoutput.n33 0.169105
R7417 CSoutput.n34 CSoutput.n12 0.169105
R7418 CSoutput.n39 CSoutput.n12 0.169105
R7419 CSoutput.n40 CSoutput.n39 0.169105
R7420 CSoutput.n40 CSoutput.n10 0.169105
R7421 CSoutput.n45 CSoutput.n10 0.169105
R7422 CSoutput.n46 CSoutput.n45 0.169105
R7423 CSoutput.n47 CSoutput.n46 0.169105
R7424 CSoutput.n47 CSoutput.n8 0.169105
R7425 CSoutput.n52 CSoutput.n8 0.169105
R7426 CSoutput.n53 CSoutput.n52 0.169105
R7427 CSoutput.n53 CSoutput.n6 0.169105
R7428 CSoutput.n58 CSoutput.n6 0.169105
R7429 CSoutput.n59 CSoutput.n58 0.169105
R7430 CSoutput.n60 CSoutput.n59 0.169105
R7431 CSoutput.n60 CSoutput.n4 0.169105
R7432 CSoutput.n66 CSoutput.n4 0.169105
R7433 CSoutput.n67 CSoutput.n66 0.169105
R7434 CSoutput.n68 CSoutput.n67 0.169105
R7435 CSoutput.n68 CSoutput.n2 0.169105
R7436 CSoutput.n73 CSoutput.n2 0.169105
R7437 CSoutput.n74 CSoutput.n73 0.169105
R7438 CSoutput.n74 CSoutput.n0 0.169105
R7439 CSoutput.n78 CSoutput.n0 0.169105
R7440 CSoutput.n219 CSoutput.n218 0.0910737
R7441 CSoutput.n270 CSoutput.n267 0.0723685
R7442 CSoutput.n224 CSoutput.n219 0.0522944
R7443 CSoutput.n267 CSoutput.n266 0.0499135
R7444 CSoutput.n218 CSoutput.n217 0.0499135
R7445 CSoutput.n252 CSoutput.n251 0.0464294
R7446 CSoutput.n260 CSoutput.n257 0.0391444
R7447 CSoutput.n219 CSoutput.t178 0.023435
R7448 CSoutput.n267 CSoutput.t172 0.02262
R7449 CSoutput.n218 CSoutput.t163 0.02262
R7450 CSoutput CSoutput.n389 0.0052
R7451 CSoutput.n189 CSoutput.n172 0.00365111
R7452 CSoutput.n192 CSoutput.n173 0.00365111
R7453 CSoutput.n175 CSoutput.n174 0.00365111
R7454 CSoutput.n217 CSoutput.n176 0.00365111
R7455 CSoutput.n181 CSoutput.n177 0.00365111
R7456 CSoutput.n264 CSoutput.n178 0.00365111
R7457 CSoutput.n255 CSoutput.n254 0.00365111
R7458 CSoutput.n235 CSoutput.n208 0.00365111
R7459 CSoutput.n237 CSoutput.n207 0.00365111
R7460 CSoutput.n225 CSoutput.n224 0.00365111
R7461 CSoutput.n231 CSoutput.n211 0.00365111
R7462 CSoutput.n233 CSoutput.n210 0.00365111
R7463 CSoutput.n155 CSoutput.n138 0.00365111
R7464 CSoutput.n158 CSoutput.n139 0.00365111
R7465 CSoutput.n141 CSoutput.n140 0.00365111
R7466 CSoutput.n251 CSoutput.n142 0.00365111
R7467 CSoutput.n147 CSoutput.n143 0.00365111
R7468 CSoutput.n274 CSoutput.n144 0.00365111
R7469 CSoutput.n186 CSoutput.n176 0.00340054
R7470 CSoutput.n179 CSoutput.n177 0.00340054
R7471 CSoutput.n264 CSoutput.n263 0.00340054
R7472 CSoutput.n259 CSoutput.n172 0.00340054
R7473 CSoutput.n188 CSoutput.n173 0.00340054
R7474 CSoutput.n191 CSoutput.n175 0.00340054
R7475 CSoutput.n230 CSoutput.n225 0.00340054
R7476 CSoutput.n232 CSoutput.n231 0.00340054
R7477 CSoutput.n234 CSoutput.n233 0.00340054
R7478 CSoutput.n256 CSoutput.n255 0.00340054
R7479 CSoutput.n236 CSoutput.n235 0.00340054
R7480 CSoutput.n238 CSoutput.n237 0.00340054
R7481 CSoutput.n152 CSoutput.n142 0.00340054
R7482 CSoutput.n145 CSoutput.n143 0.00340054
R7483 CSoutput.n274 CSoutput.n273 0.00340054
R7484 CSoutput.n269 CSoutput.n138 0.00340054
R7485 CSoutput.n154 CSoutput.n139 0.00340054
R7486 CSoutput.n157 CSoutput.n141 0.00340054
R7487 CSoutput.n187 CSoutput.n181 0.00252698
R7488 CSoutput.n180 CSoutput.n178 0.00252698
R7489 CSoutput.n262 CSoutput.n261 0.00252698
R7490 CSoutput.n190 CSoutput.n188 0.00252698
R7491 CSoutput.n193 CSoutput.n191 0.00252698
R7492 CSoutput.n266 CSoutput.n161 0.00252698
R7493 CSoutput.n187 CSoutput.n186 0.00252698
R7494 CSoutput.n180 CSoutput.n179 0.00252698
R7495 CSoutput.n263 CSoutput.n262 0.00252698
R7496 CSoutput.n190 CSoutput.n189 0.00252698
R7497 CSoutput.n193 CSoutput.n192 0.00252698
R7498 CSoutput.n174 CSoutput.n161 0.00252698
R7499 CSoutput.n241 CSoutput.n211 0.00252698
R7500 CSoutput.n240 CSoutput.n210 0.00252698
R7501 CSoutput.n239 CSoutput.n195 0.00252698
R7502 CSoutput.n236 CSoutput.n206 0.00252698
R7503 CSoutput.n243 CSoutput.n238 0.00252698
R7504 CSoutput.n252 CSoutput.n245 0.00252698
R7505 CSoutput.n241 CSoutput.n230 0.00252698
R7506 CSoutput.n240 CSoutput.n232 0.00252698
R7507 CSoutput.n239 CSoutput.n234 0.00252698
R7508 CSoutput.n254 CSoutput.n206 0.00252698
R7509 CSoutput.n243 CSoutput.n208 0.00252698
R7510 CSoutput.n245 CSoutput.n207 0.00252698
R7511 CSoutput.n153 CSoutput.n147 0.00252698
R7512 CSoutput.n146 CSoutput.n144 0.00252698
R7513 CSoutput.n272 CSoutput.n271 0.00252698
R7514 CSoutput.n156 CSoutput.n154 0.00252698
R7515 CSoutput.n159 CSoutput.n157 0.00252698
R7516 CSoutput.n276 CSoutput.n127 0.00252698
R7517 CSoutput.n153 CSoutput.n152 0.00252698
R7518 CSoutput.n146 CSoutput.n145 0.00252698
R7519 CSoutput.n273 CSoutput.n272 0.00252698
R7520 CSoutput.n156 CSoutput.n155 0.00252698
R7521 CSoutput.n159 CSoutput.n158 0.00252698
R7522 CSoutput.n140 CSoutput.n127 0.00252698
R7523 CSoutput.n261 CSoutput.n260 0.0020275
R7524 CSoutput.n260 CSoutput.n259 0.0020275
R7525 CSoutput.n257 CSoutput.n195 0.0020275
R7526 CSoutput.n257 CSoutput.n256 0.0020275
R7527 CSoutput.n271 CSoutput.n270 0.0020275
R7528 CSoutput.n270 CSoutput.n269 0.0020275
R7529 CSoutput.n171 CSoutput.n170 0.00166668
R7530 CSoutput.n253 CSoutput.n209 0.00166668
R7531 CSoutput.n137 CSoutput.n136 0.00166668
R7532 CSoutput.n275 CSoutput.n137 0.00133328
R7533 CSoutput.n209 CSoutput.n205 0.00133328
R7534 CSoutput.n265 CSoutput.n171 0.00133328
R7535 CSoutput.n268 CSoutput.n160 0.001
R7536 CSoutput.n246 CSoutput.n160 0.001
R7537 CSoutput.n148 CSoutput.n128 0.001
R7538 CSoutput.n247 CSoutput.n128 0.001
R7539 CSoutput.n149 CSoutput.n129 0.001
R7540 CSoutput.n248 CSoutput.n129 0.001
R7541 CSoutput.n150 CSoutput.n130 0.001
R7542 CSoutput.n249 CSoutput.n130 0.001
R7543 CSoutput.n151 CSoutput.n131 0.001
R7544 CSoutput.n250 CSoutput.n131 0.001
R7545 CSoutput.n244 CSoutput.n196 0.001
R7546 CSoutput.n244 CSoutput.n242 0.001
R7547 CSoutput.n226 CSoutput.n197 0.001
R7548 CSoutput.n220 CSoutput.n197 0.001
R7549 CSoutput.n227 CSoutput.n198 0.001
R7550 CSoutput.n221 CSoutput.n198 0.001
R7551 CSoutput.n228 CSoutput.n199 0.001
R7552 CSoutput.n222 CSoutput.n199 0.001
R7553 CSoutput.n229 CSoutput.n200 0.001
R7554 CSoutput.n223 CSoutput.n200 0.001
R7555 CSoutput.n258 CSoutput.n194 0.001
R7556 CSoutput.n212 CSoutput.n194 0.001
R7557 CSoutput.n182 CSoutput.n162 0.001
R7558 CSoutput.n213 CSoutput.n162 0.001
R7559 CSoutput.n183 CSoutput.n163 0.001
R7560 CSoutput.n214 CSoutput.n163 0.001
R7561 CSoutput.n184 CSoutput.n164 0.001
R7562 CSoutput.n215 CSoutput.n164 0.001
R7563 CSoutput.n185 CSoutput.n165 0.001
R7564 CSoutput.n216 CSoutput.n165 0.001
R7565 CSoutput.n216 CSoutput.n166 0.001
R7566 CSoutput.n215 CSoutput.n167 0.001
R7567 CSoutput.n214 CSoutput.n168 0.001
R7568 CSoutput.n213 CSoutput.t175 0.001
R7569 CSoutput.n212 CSoutput.n169 0.001
R7570 CSoutput.n185 CSoutput.n167 0.001
R7571 CSoutput.n184 CSoutput.n168 0.001
R7572 CSoutput.n183 CSoutput.t175 0.001
R7573 CSoutput.n182 CSoutput.n169 0.001
R7574 CSoutput.n258 CSoutput.n170 0.001
R7575 CSoutput.n223 CSoutput.n201 0.001
R7576 CSoutput.n222 CSoutput.n202 0.001
R7577 CSoutput.n221 CSoutput.n203 0.001
R7578 CSoutput.n220 CSoutput.t171 0.001
R7579 CSoutput.n242 CSoutput.n204 0.001
R7580 CSoutput.n229 CSoutput.n202 0.001
R7581 CSoutput.n228 CSoutput.n203 0.001
R7582 CSoutput.n227 CSoutput.t171 0.001
R7583 CSoutput.n226 CSoutput.n204 0.001
R7584 CSoutput.n253 CSoutput.n196 0.001
R7585 CSoutput.n250 CSoutput.n132 0.001
R7586 CSoutput.n249 CSoutput.n133 0.001
R7587 CSoutput.n248 CSoutput.n134 0.001
R7588 CSoutput.n247 CSoutput.t161 0.001
R7589 CSoutput.n246 CSoutput.n135 0.001
R7590 CSoutput.n151 CSoutput.n133 0.001
R7591 CSoutput.n150 CSoutput.n134 0.001
R7592 CSoutput.n149 CSoutput.t161 0.001
R7593 CSoutput.n148 CSoutput.n135 0.001
R7594 CSoutput.n268 CSoutput.n136 0.001
R7595 a_n2650_13878.n136 a_n2650_13878.t6 512.366
R7596 a_n2650_13878.n135 a_n2650_13878.t40 512.366
R7597 a_n2650_13878.n71 a_n2650_13878.t38 512.366
R7598 a_n2650_13878.n134 a_n2650_13878.t42 512.366
R7599 a_n2650_13878.n133 a_n2650_13878.t18 512.366
R7600 a_n2650_13878.n72 a_n2650_13878.t30 512.366
R7601 a_n2650_13878.n132 a_n2650_13878.t22 512.366
R7602 a_n2650_13878.n131 a_n2650_13878.t28 512.366
R7603 a_n2650_13878.n73 a_n2650_13878.t12 512.366
R7604 a_n2650_13878.n118 a_n2650_13878.t98 512.366
R7605 a_n2650_13878.n117 a_n2650_13878.t77 512.366
R7606 a_n2650_13878.n74 a_n2650_13878.t82 512.366
R7607 a_n2650_13878.n116 a_n2650_13878.t71 512.366
R7608 a_n2650_13878.n115 a_n2650_13878.t87 512.366
R7609 a_n2650_13878.n75 a_n2650_13878.t95 512.366
R7610 a_n2650_13878.n114 a_n2650_13878.t96 512.366
R7611 a_n2650_13878.n113 a_n2650_13878.t66 512.366
R7612 a_n2650_13878.n76 a_n2650_13878.t79 512.366
R7613 a_n2650_13878.n92 a_n2650_13878.t20 512.366
R7614 a_n2650_13878.n93 a_n2650_13878.t10 512.366
R7615 a_n2650_13878.n82 a_n2650_13878.t26 512.366
R7616 a_n2650_13878.n94 a_n2650_13878.t32 512.366
R7617 a_n2650_13878.n95 a_n2650_13878.t16 512.366
R7618 a_n2650_13878.n96 a_n2650_13878.t24 512.366
R7619 a_n2650_13878.n97 a_n2650_13878.t36 512.366
R7620 a_n2650_13878.n81 a_n2650_13878.t34 512.366
R7621 a_n2650_13878.n98 a_n2650_13878.t8 512.366
R7622 a_n2650_13878.n85 a_n2650_13878.t70 512.366
R7623 a_n2650_13878.n86 a_n2650_13878.t93 512.366
R7624 a_n2650_13878.n84 a_n2650_13878.t94 512.366
R7625 a_n2650_13878.n87 a_n2650_13878.t68 512.366
R7626 a_n2650_13878.n88 a_n2650_13878.t90 512.366
R7627 a_n2650_13878.n89 a_n2650_13878.t91 512.366
R7628 a_n2650_13878.n90 a_n2650_13878.t65 512.366
R7629 a_n2650_13878.n83 a_n2650_13878.t76 512.366
R7630 a_n2650_13878.n91 a_n2650_13878.t86 512.366
R7631 a_n2650_13878.n110 a_n2650_13878.t84 512.366
R7632 a_n2650_13878.n100 a_n2650_13878.t74 512.366
R7633 a_n2650_13878.n111 a_n2650_13878.t64 512.366
R7634 a_n2650_13878.n108 a_n2650_13878.t92 512.366
R7635 a_n2650_13878.n101 a_n2650_13878.t81 512.366
R7636 a_n2650_13878.n109 a_n2650_13878.t80 512.366
R7637 a_n2650_13878.n106 a_n2650_13878.t88 512.366
R7638 a_n2650_13878.n102 a_n2650_13878.t72 512.366
R7639 a_n2650_13878.n107 a_n2650_13878.t73 512.366
R7640 a_n2650_13878.n104 a_n2650_13878.t75 512.366
R7641 a_n2650_13878.n103 a_n2650_13878.t85 512.366
R7642 a_n2650_13878.n105 a_n2650_13878.t99 512.366
R7643 a_n2650_13878.n34 a_n2650_13878.n70 70.1674
R7644 a_n2650_13878.n4 a_n2650_13878.n63 70.1674
R7645 a_n2650_13878.n17 a_n2650_13878.n48 70.1674
R7646 a_n2650_13878.n21 a_n2650_13878.n41 70.1674
R7647 a_n2650_13878.n91 a_n2650_13878.n41 20.9683
R7648 a_n2650_13878.n40 a_n2650_13878.n21 74.73
R7649 a_n2650_13878.n40 a_n2650_13878.n83 11.843
R7650 a_n2650_13878.n20 a_n2650_13878.n39 80.4688
R7651 a_n2650_13878.n90 a_n2650_13878.n39 0.365327
R7652 a_n2650_13878.n38 a_n2650_13878.n20 75.0448
R7653 a_n2650_13878.n22 a_n2650_13878.n37 70.1674
R7654 a_n2650_13878.n87 a_n2650_13878.n37 20.9683
R7655 a_n2650_13878.n36 a_n2650_13878.n22 70.3058
R7656 a_n2650_13878.n36 a_n2650_13878.n84 20.6913
R7657 a_n2650_13878.n23 a_n2650_13878.n35 75.3623
R7658 a_n2650_13878.n86 a_n2650_13878.n35 10.5784
R7659 a_n2650_13878.n85 a_n2650_13878.n23 161.3
R7660 a_n2650_13878.n98 a_n2650_13878.n48 20.9683
R7661 a_n2650_13878.n47 a_n2650_13878.n17 74.73
R7662 a_n2650_13878.n47 a_n2650_13878.n81 11.843
R7663 a_n2650_13878.n16 a_n2650_13878.n46 80.4688
R7664 a_n2650_13878.n97 a_n2650_13878.n46 0.365327
R7665 a_n2650_13878.n45 a_n2650_13878.n16 75.0448
R7666 a_n2650_13878.n18 a_n2650_13878.n44 70.1674
R7667 a_n2650_13878.n94 a_n2650_13878.n44 20.9683
R7668 a_n2650_13878.n43 a_n2650_13878.n18 70.3058
R7669 a_n2650_13878.n43 a_n2650_13878.n82 20.6913
R7670 a_n2650_13878.n19 a_n2650_13878.n42 75.3623
R7671 a_n2650_13878.n93 a_n2650_13878.n42 10.5784
R7672 a_n2650_13878.n92 a_n2650_13878.n19 161.3
R7673 a_n2650_13878.n7 a_n2650_13878.n56 70.1674
R7674 a_n2650_13878.n9 a_n2650_13878.n54 70.1674
R7675 a_n2650_13878.n11 a_n2650_13878.n52 70.1674
R7676 a_n2650_13878.n14 a_n2650_13878.n50 70.1674
R7677 a_n2650_13878.n105 a_n2650_13878.n50 20.9683
R7678 a_n2650_13878.n49 a_n2650_13878.n15 75.0448
R7679 a_n2650_13878.n49 a_n2650_13878.n103 11.2134
R7680 a_n2650_13878.n15 a_n2650_13878.n104 161.3
R7681 a_n2650_13878.n107 a_n2650_13878.n52 20.9683
R7682 a_n2650_13878.n51 a_n2650_13878.n12 75.0448
R7683 a_n2650_13878.n51 a_n2650_13878.n102 11.2134
R7684 a_n2650_13878.n12 a_n2650_13878.n106 161.3
R7685 a_n2650_13878.n109 a_n2650_13878.n54 20.9683
R7686 a_n2650_13878.n53 a_n2650_13878.n10 75.0448
R7687 a_n2650_13878.n53 a_n2650_13878.n101 11.2134
R7688 a_n2650_13878.n10 a_n2650_13878.n108 161.3
R7689 a_n2650_13878.n111 a_n2650_13878.n56 20.9683
R7690 a_n2650_13878.n55 a_n2650_13878.n8 75.0448
R7691 a_n2650_13878.n55 a_n2650_13878.n100 11.2134
R7692 a_n2650_13878.n8 a_n2650_13878.n110 161.3
R7693 a_n2650_13878.n63 a_n2650_13878.n76 20.9683
R7694 a_n2650_13878.n62 a_n2650_13878.n4 74.73
R7695 a_n2650_13878.n113 a_n2650_13878.n62 11.843
R7696 a_n2650_13878.n61 a_n2650_13878.n3 80.4688
R7697 a_n2650_13878.n61 a_n2650_13878.n114 0.365327
R7698 a_n2650_13878.n3 a_n2650_13878.n60 75.0448
R7699 a_n2650_13878.n59 a_n2650_13878.n5 70.1674
R7700 a_n2650_13878.n116 a_n2650_13878.n59 20.9683
R7701 a_n2650_13878.n5 a_n2650_13878.n58 70.3058
R7702 a_n2650_13878.n58 a_n2650_13878.n74 20.6913
R7703 a_n2650_13878.n57 a_n2650_13878.n6 75.3623
R7704 a_n2650_13878.n117 a_n2650_13878.n57 10.5784
R7705 a_n2650_13878.n6 a_n2650_13878.n118 161.3
R7706 a_n2650_13878.n70 a_n2650_13878.n73 20.9683
R7707 a_n2650_13878.n69 a_n2650_13878.n34 74.73
R7708 a_n2650_13878.n131 a_n2650_13878.n69 11.843
R7709 a_n2650_13878.n68 a_n2650_13878.n1 80.4688
R7710 a_n2650_13878.n68 a_n2650_13878.n132 0.365327
R7711 a_n2650_13878.n1 a_n2650_13878.n67 75.0448
R7712 a_n2650_13878.n66 a_n2650_13878.n0 70.1674
R7713 a_n2650_13878.n134 a_n2650_13878.n66 20.9683
R7714 a_n2650_13878.n0 a_n2650_13878.n65 70.3058
R7715 a_n2650_13878.n65 a_n2650_13878.n71 20.6913
R7716 a_n2650_13878.n64 a_n2650_13878.n2 75.3623
R7717 a_n2650_13878.n135 a_n2650_13878.n64 10.5784
R7718 a_n2650_13878.n2 a_n2650_13878.n136 161.3
R7719 a_n2650_13878.n32 a_n2650_13878.n128 81.2902
R7720 a_n2650_13878.n33 a_n2650_13878.n122 81.2902
R7721 a_n2650_13878.n24 a_n2650_13878.n119 81.2902
R7722 a_n2650_13878.n32 a_n2650_13878.n129 80.9324
R7723 a_n2650_13878.n26 a_n2650_13878.n130 80.9324
R7724 a_n2650_13878.n26 a_n2650_13878.n127 80.9324
R7725 a_n2650_13878.n26 a_n2650_13878.n126 80.9324
R7726 a_n2650_13878.n25 a_n2650_13878.n125 80.9324
R7727 a_n2650_13878.n33 a_n2650_13878.n123 80.9324
R7728 a_n2650_13878.n24 a_n2650_13878.n124 80.9324
R7729 a_n2650_13878.n24 a_n2650_13878.n121 80.9324
R7730 a_n2650_13878.n24 a_n2650_13878.n120 80.9324
R7731 a_n2650_13878.n30 a_n2650_13878.t15 74.6477
R7732 a_n2650_13878.n27 a_n2650_13878.t21 74.6477
R7733 a_n2650_13878.t7 a_n2650_13878.n142 74.2899
R7734 a_n2650_13878.n29 a_n2650_13878.t45 74.2897
R7735 a_n2650_13878.n30 a_n2650_13878.n138 70.6783
R7736 a_n2650_13878.n30 a_n2650_13878.n139 70.6783
R7737 a_n2650_13878.n31 a_n2650_13878.n140 70.6783
R7738 a_n2650_13878.n31 a_n2650_13878.n141 70.6783
R7739 a_n2650_13878.n29 a_n2650_13878.n80 70.6783
R7740 a_n2650_13878.n28 a_n2650_13878.n79 70.6783
R7741 a_n2650_13878.n28 a_n2650_13878.n78 70.6783
R7742 a_n2650_13878.n27 a_n2650_13878.n77 70.6783
R7743 a_n2650_13878.n136 a_n2650_13878.n135 48.2005
R7744 a_n2650_13878.n66 a_n2650_13878.n133 20.9683
R7745 a_n2650_13878.n132 a_n2650_13878.n72 48.2005
R7746 a_n2650_13878.t14 a_n2650_13878.n70 533.335
R7747 a_n2650_13878.n118 a_n2650_13878.n117 48.2005
R7748 a_n2650_13878.n59 a_n2650_13878.n115 20.9683
R7749 a_n2650_13878.n114 a_n2650_13878.n75 48.2005
R7750 a_n2650_13878.t69 a_n2650_13878.n63 533.335
R7751 a_n2650_13878.n93 a_n2650_13878.n92 48.2005
R7752 a_n2650_13878.n95 a_n2650_13878.n44 20.9683
R7753 a_n2650_13878.n97 a_n2650_13878.n96 48.2005
R7754 a_n2650_13878.t44 a_n2650_13878.n48 533.335
R7755 a_n2650_13878.n86 a_n2650_13878.n85 48.2005
R7756 a_n2650_13878.n88 a_n2650_13878.n37 20.9683
R7757 a_n2650_13878.n90 a_n2650_13878.n89 48.2005
R7758 a_n2650_13878.t67 a_n2650_13878.n41 533.335
R7759 a_n2650_13878.n110 a_n2650_13878.n100 48.2005
R7760 a_n2650_13878.t89 a_n2650_13878.n56 533.335
R7761 a_n2650_13878.n108 a_n2650_13878.n101 48.2005
R7762 a_n2650_13878.t97 a_n2650_13878.n54 533.335
R7763 a_n2650_13878.n106 a_n2650_13878.n102 48.2005
R7764 a_n2650_13878.t83 a_n2650_13878.n52 533.335
R7765 a_n2650_13878.n104 a_n2650_13878.n103 48.2005
R7766 a_n2650_13878.t78 a_n2650_13878.n50 533.335
R7767 a_n2650_13878.n134 a_n2650_13878.n65 21.4216
R7768 a_n2650_13878.n116 a_n2650_13878.n58 21.4216
R7769 a_n2650_13878.n94 a_n2650_13878.n43 21.4216
R7770 a_n2650_13878.n87 a_n2650_13878.n36 21.4216
R7771 a_n2650_13878.n25 a_n2650_13878.n24 31.7747
R7772 a_n2650_13878.n69 a_n2650_13878.n73 34.4824
R7773 a_n2650_13878.n62 a_n2650_13878.n76 34.4824
R7774 a_n2650_13878.n98 a_n2650_13878.n47 34.4824
R7775 a_n2650_13878.n91 a_n2650_13878.n40 34.4824
R7776 a_n2650_13878.n133 a_n2650_13878.n67 35.3134
R7777 a_n2650_13878.n67 a_n2650_13878.n72 11.2134
R7778 a_n2650_13878.n115 a_n2650_13878.n60 35.3134
R7779 a_n2650_13878.n60 a_n2650_13878.n75 11.2134
R7780 a_n2650_13878.n95 a_n2650_13878.n45 35.3134
R7781 a_n2650_13878.n96 a_n2650_13878.n45 11.2134
R7782 a_n2650_13878.n88 a_n2650_13878.n38 35.3134
R7783 a_n2650_13878.n89 a_n2650_13878.n38 11.2134
R7784 a_n2650_13878.n111 a_n2650_13878.n55 35.3134
R7785 a_n2650_13878.n109 a_n2650_13878.n53 35.3134
R7786 a_n2650_13878.n107 a_n2650_13878.n51 35.3134
R7787 a_n2650_13878.n105 a_n2650_13878.n49 35.3134
R7788 a_n2650_13878.n34 a_n2650_13878.n26 23.891
R7789 a_n2650_13878.n64 a_n2650_13878.n71 36.139
R7790 a_n2650_13878.n57 a_n2650_13878.n74 36.139
R7791 a_n2650_13878.n82 a_n2650_13878.n42 36.139
R7792 a_n2650_13878.n84 a_n2650_13878.n35 36.139
R7793 a_n2650_13878.n23 a_n2650_13878.n13 13.3641
R7794 a_n2650_13878.n4 a_n2650_13878.n112 13.1596
R7795 a_n2650_13878.n137 a_n2650_13878.n2 11.8547
R7796 a_n2650_13878.n99 a_n2650_13878.n29 10.2167
R7797 a_n2650_13878.n15 a_n2650_13878.n13 9.99103
R7798 a_n2650_13878.n112 a_n2650_13878.n7 9.99103
R7799 a_n2650_13878.n99 a_n2650_13878.n17 8.01944
R7800 a_n2650_13878.n142 a_n2650_13878.n137 6.37334
R7801 a_n2650_13878.n112 a_n2650_13878.n99 5.3452
R7802 a_n2650_13878.n19 a_n2650_13878.n21 4.07247
R7803 a_n2650_13878.n34 a_n2650_13878.n6 4.06674
R7804 a_n2650_13878.n138 a_n2650_13878.t29 3.61217
R7805 a_n2650_13878.n138 a_n2650_13878.t13 3.61217
R7806 a_n2650_13878.n139 a_n2650_13878.t31 3.61217
R7807 a_n2650_13878.n139 a_n2650_13878.t23 3.61217
R7808 a_n2650_13878.n140 a_n2650_13878.t43 3.61217
R7809 a_n2650_13878.n140 a_n2650_13878.t19 3.61217
R7810 a_n2650_13878.n141 a_n2650_13878.t41 3.61217
R7811 a_n2650_13878.n141 a_n2650_13878.t39 3.61217
R7812 a_n2650_13878.n80 a_n2650_13878.t35 3.61217
R7813 a_n2650_13878.n80 a_n2650_13878.t9 3.61217
R7814 a_n2650_13878.n79 a_n2650_13878.t25 3.61217
R7815 a_n2650_13878.n79 a_n2650_13878.t37 3.61217
R7816 a_n2650_13878.n78 a_n2650_13878.t33 3.61217
R7817 a_n2650_13878.n78 a_n2650_13878.t17 3.61217
R7818 a_n2650_13878.n77 a_n2650_13878.t11 3.61217
R7819 a_n2650_13878.n77 a_n2650_13878.t27 3.61217
R7820 a_n2650_13878.n128 a_n2650_13878.t4 2.82907
R7821 a_n2650_13878.n128 a_n2650_13878.t52 2.82907
R7822 a_n2650_13878.n129 a_n2650_13878.t3 2.82907
R7823 a_n2650_13878.n129 a_n2650_13878.t53 2.82907
R7824 a_n2650_13878.n130 a_n2650_13878.t55 2.82907
R7825 a_n2650_13878.n130 a_n2650_13878.t58 2.82907
R7826 a_n2650_13878.n127 a_n2650_13878.t47 2.82907
R7827 a_n2650_13878.n127 a_n2650_13878.t60 2.82907
R7828 a_n2650_13878.n126 a_n2650_13878.t49 2.82907
R7829 a_n2650_13878.n126 a_n2650_13878.t2 2.82907
R7830 a_n2650_13878.n125 a_n2650_13878.t5 2.82907
R7831 a_n2650_13878.n125 a_n2650_13878.t50 2.82907
R7832 a_n2650_13878.n122 a_n2650_13878.t0 2.82907
R7833 a_n2650_13878.n122 a_n2650_13878.t48 2.82907
R7834 a_n2650_13878.n123 a_n2650_13878.t57 2.82907
R7835 a_n2650_13878.n123 a_n2650_13878.t46 2.82907
R7836 a_n2650_13878.n124 a_n2650_13878.t54 2.82907
R7837 a_n2650_13878.n124 a_n2650_13878.t62 2.82907
R7838 a_n2650_13878.n121 a_n2650_13878.t51 2.82907
R7839 a_n2650_13878.n121 a_n2650_13878.t56 2.82907
R7840 a_n2650_13878.n120 a_n2650_13878.t1 2.82907
R7841 a_n2650_13878.n120 a_n2650_13878.t59 2.82907
R7842 a_n2650_13878.n119 a_n2650_13878.t63 2.82907
R7843 a_n2650_13878.n119 a_n2650_13878.t61 2.82907
R7844 a_n2650_13878.n137 a_n2650_13878.n13 1.30542
R7845 a_n2650_13878.n10 a_n2650_13878.n11 1.04595
R7846 a_n2650_13878.n68 a_n2650_13878.n131 47.835
R7847 a_n2650_13878.n61 a_n2650_13878.n113 47.835
R7848 a_n2650_13878.n81 a_n2650_13878.n46 47.835
R7849 a_n2650_13878.n83 a_n2650_13878.n39 47.835
R7850 a_n2650_13878.n21 a_n2650_13878.n20 1.13686
R7851 a_n2650_13878.n17 a_n2650_13878.n16 1.13686
R7852 a_n2650_13878.n4 a_n2650_13878.n3 1.13686
R7853 a_n2650_13878.n34 a_n2650_13878.n1 1.10471
R7854 a_n2650_13878.n24 a_n2650_13878.n33 1.07378
R7855 a_n2650_13878.n22 a_n2650_13878.n23 0.758076
R7856 a_n2650_13878.n20 a_n2650_13878.n22 0.758076
R7857 a_n2650_13878.n18 a_n2650_13878.n19 0.758076
R7858 a_n2650_13878.n16 a_n2650_13878.n18 0.758076
R7859 a_n2650_13878.n15 a_n2650_13878.n14 0.758076
R7860 a_n2650_13878.n12 a_n2650_13878.n11 0.758076
R7861 a_n2650_13878.n10 a_n2650_13878.n9 0.758076
R7862 a_n2650_13878.n8 a_n2650_13878.n7 0.758076
R7863 a_n2650_13878.n6 a_n2650_13878.n5 0.758076
R7864 a_n2650_13878.n3 a_n2650_13878.n5 0.758076
R7865 a_n2650_13878.n2 a_n2650_13878.n0 0.758076
R7866 a_n2650_13878.n1 a_n2650_13878.n0 0.758076
R7867 a_n2650_13878.n26 a_n2650_13878.n32 0.716017
R7868 a_n2650_13878.n31 a_n2650_13878.n30 0.716017
R7869 a_n2650_13878.n142 a_n2650_13878.n31 0.716017
R7870 a_n2650_13878.n29 a_n2650_13878.n28 0.716017
R7871 a_n2650_13878.n28 a_n2650_13878.n27 0.716017
R7872 a_n2650_13878.n26 a_n2650_13878.n25 0.716017
R7873 a_n2650_13878.n12 a_n2650_13878.n14 0.67853
R7874 a_n2650_13878.n8 a_n2650_13878.n9 0.67853
R7875 a_n2472_13878.n25 a_n2472_13878.n24 98.9632
R7876 a_n2472_13878.n2 a_n2472_13878.n0 98.7517
R7877 a_n2472_13878.n20 a_n2472_13878.n19 98.6055
R7878 a_n2472_13878.n22 a_n2472_13878.n21 98.6055
R7879 a_n2472_13878.n24 a_n2472_13878.n23 98.6055
R7880 a_n2472_13878.n8 a_n2472_13878.n7 98.6055
R7881 a_n2472_13878.n6 a_n2472_13878.n5 98.6055
R7882 a_n2472_13878.n4 a_n2472_13878.n3 98.6055
R7883 a_n2472_13878.n2 a_n2472_13878.n1 98.6055
R7884 a_n2472_13878.n18 a_n2472_13878.n17 98.6054
R7885 a_n2472_13878.n10 a_n2472_13878.t21 74.6477
R7886 a_n2472_13878.n15 a_n2472_13878.t22 74.2899
R7887 a_n2472_13878.n12 a_n2472_13878.t23 74.2899
R7888 a_n2472_13878.n11 a_n2472_13878.t20 74.2899
R7889 a_n2472_13878.n14 a_n2472_13878.n13 70.6783
R7890 a_n2472_13878.n10 a_n2472_13878.n9 70.6783
R7891 a_n2472_13878.n16 a_n2472_13878.n8 15.0004
R7892 a_n2472_13878.n18 a_n2472_13878.n16 12.2917
R7893 a_n2472_13878.n16 a_n2472_13878.n15 7.67184
R7894 a_n2472_13878.n17 a_n2472_13878.t16 3.61217
R7895 a_n2472_13878.n17 a_n2472_13878.t5 3.61217
R7896 a_n2472_13878.n19 a_n2472_13878.t8 3.61217
R7897 a_n2472_13878.n19 a_n2472_13878.t9 3.61217
R7898 a_n2472_13878.n21 a_n2472_13878.t17 3.61217
R7899 a_n2472_13878.n21 a_n2472_13878.t18 3.61217
R7900 a_n2472_13878.n23 a_n2472_13878.t0 3.61217
R7901 a_n2472_13878.n23 a_n2472_13878.t10 3.61217
R7902 a_n2472_13878.n13 a_n2472_13878.t26 3.61217
R7903 a_n2472_13878.n13 a_n2472_13878.t27 3.61217
R7904 a_n2472_13878.n9 a_n2472_13878.t24 3.61217
R7905 a_n2472_13878.n9 a_n2472_13878.t25 3.61217
R7906 a_n2472_13878.n7 a_n2472_13878.t11 3.61217
R7907 a_n2472_13878.n7 a_n2472_13878.t1 3.61217
R7908 a_n2472_13878.n5 a_n2472_13878.t14 3.61217
R7909 a_n2472_13878.n5 a_n2472_13878.t3 3.61217
R7910 a_n2472_13878.n3 a_n2472_13878.t2 3.61217
R7911 a_n2472_13878.n3 a_n2472_13878.t4 3.61217
R7912 a_n2472_13878.n1 a_n2472_13878.t12 3.61217
R7913 a_n2472_13878.n1 a_n2472_13878.t6 3.61217
R7914 a_n2472_13878.n0 a_n2472_13878.t15 3.61217
R7915 a_n2472_13878.n0 a_n2472_13878.t7 3.61217
R7916 a_n2472_13878.n25 a_n2472_13878.t13 3.61217
R7917 a_n2472_13878.t19 a_n2472_13878.n25 3.61217
R7918 a_n2472_13878.n11 a_n2472_13878.n10 0.358259
R7919 a_n2472_13878.n14 a_n2472_13878.n12 0.358259
R7920 a_n2472_13878.n15 a_n2472_13878.n14 0.358259
R7921 a_n2472_13878.n24 a_n2472_13878.n22 0.358259
R7922 a_n2472_13878.n22 a_n2472_13878.n20 0.358259
R7923 a_n2472_13878.n20 a_n2472_13878.n18 0.358259
R7924 a_n2472_13878.n4 a_n2472_13878.n2 0.146627
R7925 a_n2472_13878.n6 a_n2472_13878.n4 0.146627
R7926 a_n2472_13878.n8 a_n2472_13878.n6 0.146627
R7927 a_n2472_13878.n12 a_n2472_13878.n11 0.101793
R7928 commonsourceibias.n35 commonsourceibias.t58 223.028
R7929 commonsourceibias.n128 commonsourceibias.t85 223.028
R7930 commonsourceibias.n217 commonsourceibias.t75 223.028
R7931 commonsourceibias.n364 commonsourceibias.t30 223.028
R7932 commonsourceibias.n305 commonsourceibias.t91 223.028
R7933 commonsourceibias.n499 commonsourceibias.t78 223.028
R7934 commonsourceibias.n99 commonsourceibias.t60 207.983
R7935 commonsourceibias.n192 commonsourceibias.t92 207.983
R7936 commonsourceibias.n281 commonsourceibias.t81 207.983
R7937 commonsourceibias.n430 commonsourceibias.t20 207.983
R7938 commonsourceibias.n476 commonsourceibias.t110 207.983
R7939 commonsourceibias.n565 commonsourceibias.t97 207.983
R7940 commonsourceibias.n97 commonsourceibias.t28 168.701
R7941 commonsourceibias.n91 commonsourceibias.t0 168.701
R7942 commonsourceibias.n17 commonsourceibias.t18 168.701
R7943 commonsourceibias.n83 commonsourceibias.t50 168.701
R7944 commonsourceibias.n77 commonsourceibias.t62 168.701
R7945 commonsourceibias.n22 commonsourceibias.t8 168.701
R7946 commonsourceibias.n69 commonsourceibias.t48 168.701
R7947 commonsourceibias.n63 commonsourceibias.t22 168.701
R7948 commonsourceibias.n25 commonsourceibias.t54 168.701
R7949 commonsourceibias.n27 commonsourceibias.t36 168.701
R7950 commonsourceibias.n29 commonsourceibias.t10 168.701
R7951 commonsourceibias.n46 commonsourceibias.t52 168.701
R7952 commonsourceibias.n40 commonsourceibias.t34 168.701
R7953 commonsourceibias.n34 commonsourceibias.t14 168.701
R7954 commonsourceibias.n190 commonsourceibias.t106 168.701
R7955 commonsourceibias.n184 commonsourceibias.t119 168.701
R7956 commonsourceibias.n5 commonsourceibias.t84 168.701
R7957 commonsourceibias.n176 commonsourceibias.t100 168.701
R7958 commonsourceibias.n170 commonsourceibias.t114 168.701
R7959 commonsourceibias.n10 commonsourceibias.t80 168.701
R7960 commonsourceibias.n162 commonsourceibias.t76 168.701
R7961 commonsourceibias.n156 commonsourceibias.t105 168.701
R7962 commonsourceibias.n118 commonsourceibias.t121 168.701
R7963 commonsourceibias.n120 commonsourceibias.t71 168.701
R7964 commonsourceibias.n122 commonsourceibias.t99 168.701
R7965 commonsourceibias.n139 commonsourceibias.t95 168.701
R7966 commonsourceibias.n133 commonsourceibias.t109 168.701
R7967 commonsourceibias.n127 commonsourceibias.t89 168.701
R7968 commonsourceibias.n216 commonsourceibias.t77 168.701
R7969 commonsourceibias.n222 commonsourceibias.t96 168.701
R7970 commonsourceibias.n228 commonsourceibias.t82 168.701
R7971 commonsourceibias.n211 commonsourceibias.t86 168.701
R7972 commonsourceibias.n209 commonsourceibias.t127 168.701
R7973 commonsourceibias.n207 commonsourceibias.t108 168.701
R7974 commonsourceibias.n245 commonsourceibias.t93 168.701
R7975 commonsourceibias.n251 commonsourceibias.t67 168.701
R7976 commonsourceibias.n204 commonsourceibias.t70 168.701
R7977 commonsourceibias.n259 commonsourceibias.t101 168.701
R7978 commonsourceibias.n265 commonsourceibias.t87 168.701
R7979 commonsourceibias.n199 commonsourceibias.t74 168.701
R7980 commonsourceibias.n273 commonsourceibias.t107 168.701
R7981 commonsourceibias.n279 commonsourceibias.t94 168.701
R7982 commonsourceibias.n363 commonsourceibias.t46 168.701
R7983 commonsourceibias.n369 commonsourceibias.t24 168.701
R7984 commonsourceibias.n375 commonsourceibias.t42 168.701
R7985 commonsourceibias.n358 commonsourceibias.t2 168.701
R7986 commonsourceibias.n356 commonsourceibias.t32 168.701
R7987 commonsourceibias.n354 commonsourceibias.t44 168.701
R7988 commonsourceibias.n392 commonsourceibias.t6 168.701
R7989 commonsourceibias.n398 commonsourceibias.t38 168.701
R7990 commonsourceibias.n400 commonsourceibias.t4 168.701
R7991 commonsourceibias.n407 commonsourceibias.t16 168.701
R7992 commonsourceibias.n413 commonsourceibias.t40 168.701
R7993 commonsourceibias.n415 commonsourceibias.t12 168.701
R7994 commonsourceibias.n422 commonsourceibias.t26 168.701
R7995 commonsourceibias.n428 commonsourceibias.t56 168.701
R7996 commonsourceibias.n474 commonsourceibias.t123 168.701
R7997 commonsourceibias.n468 commonsourceibias.t68 168.701
R7998 commonsourceibias.n461 commonsourceibias.t102 168.701
R7999 commonsourceibias.n459 commonsourceibias.t117 168.701
R8000 commonsourceibias.n453 commonsourceibias.t64 168.701
R8001 commonsourceibias.n446 commonsourceibias.t72 168.701
R8002 commonsourceibias.n444 commonsourceibias.t90 168.701
R8003 commonsourceibias.n304 commonsourceibias.t83 168.701
R8004 commonsourceibias.n310 commonsourceibias.t126 168.701
R8005 commonsourceibias.n316 commonsourceibias.t113 168.701
R8006 commonsourceibias.n299 commonsourceibias.t116 168.701
R8007 commonsourceibias.n297 commonsourceibias.t66 168.701
R8008 commonsourceibias.n295 commonsourceibias.t69 168.701
R8009 commonsourceibias.n333 commonsourceibias.t122 168.701
R8010 commonsourceibias.n498 commonsourceibias.t73 168.701
R8011 commonsourceibias.n504 commonsourceibias.t115 168.701
R8012 commonsourceibias.n510 commonsourceibias.t98 168.701
R8013 commonsourceibias.n493 commonsourceibias.t103 168.701
R8014 commonsourceibias.n491 commonsourceibias.t120 168.701
R8015 commonsourceibias.n489 commonsourceibias.t125 168.701
R8016 commonsourceibias.n527 commonsourceibias.t111 168.701
R8017 commonsourceibias.n533 commonsourceibias.t79 168.701
R8018 commonsourceibias.n535 commonsourceibias.t65 168.701
R8019 commonsourceibias.n542 commonsourceibias.t118 168.701
R8020 commonsourceibias.n548 commonsourceibias.t104 168.701
R8021 commonsourceibias.n550 commonsourceibias.t88 168.701
R8022 commonsourceibias.n557 commonsourceibias.t124 168.701
R8023 commonsourceibias.n563 commonsourceibias.t112 168.701
R8024 commonsourceibias.n36 commonsourceibias.n33 161.3
R8025 commonsourceibias.n38 commonsourceibias.n37 161.3
R8026 commonsourceibias.n39 commonsourceibias.n32 161.3
R8027 commonsourceibias.n42 commonsourceibias.n41 161.3
R8028 commonsourceibias.n43 commonsourceibias.n31 161.3
R8029 commonsourceibias.n45 commonsourceibias.n44 161.3
R8030 commonsourceibias.n47 commonsourceibias.n30 161.3
R8031 commonsourceibias.n49 commonsourceibias.n48 161.3
R8032 commonsourceibias.n51 commonsourceibias.n50 161.3
R8033 commonsourceibias.n52 commonsourceibias.n28 161.3
R8034 commonsourceibias.n54 commonsourceibias.n53 161.3
R8035 commonsourceibias.n56 commonsourceibias.n55 161.3
R8036 commonsourceibias.n57 commonsourceibias.n26 161.3
R8037 commonsourceibias.n59 commonsourceibias.n58 161.3
R8038 commonsourceibias.n61 commonsourceibias.n60 161.3
R8039 commonsourceibias.n62 commonsourceibias.n24 161.3
R8040 commonsourceibias.n65 commonsourceibias.n64 161.3
R8041 commonsourceibias.n66 commonsourceibias.n23 161.3
R8042 commonsourceibias.n68 commonsourceibias.n67 161.3
R8043 commonsourceibias.n70 commonsourceibias.n21 161.3
R8044 commonsourceibias.n72 commonsourceibias.n71 161.3
R8045 commonsourceibias.n73 commonsourceibias.n20 161.3
R8046 commonsourceibias.n75 commonsourceibias.n74 161.3
R8047 commonsourceibias.n76 commonsourceibias.n19 161.3
R8048 commonsourceibias.n79 commonsourceibias.n78 161.3
R8049 commonsourceibias.n80 commonsourceibias.n18 161.3
R8050 commonsourceibias.n82 commonsourceibias.n81 161.3
R8051 commonsourceibias.n84 commonsourceibias.n16 161.3
R8052 commonsourceibias.n86 commonsourceibias.n85 161.3
R8053 commonsourceibias.n87 commonsourceibias.n15 161.3
R8054 commonsourceibias.n89 commonsourceibias.n88 161.3
R8055 commonsourceibias.n90 commonsourceibias.n14 161.3
R8056 commonsourceibias.n93 commonsourceibias.n92 161.3
R8057 commonsourceibias.n94 commonsourceibias.n13 161.3
R8058 commonsourceibias.n96 commonsourceibias.n95 161.3
R8059 commonsourceibias.n98 commonsourceibias.n12 161.3
R8060 commonsourceibias.n129 commonsourceibias.n126 161.3
R8061 commonsourceibias.n131 commonsourceibias.n130 161.3
R8062 commonsourceibias.n132 commonsourceibias.n125 161.3
R8063 commonsourceibias.n135 commonsourceibias.n134 161.3
R8064 commonsourceibias.n136 commonsourceibias.n124 161.3
R8065 commonsourceibias.n138 commonsourceibias.n137 161.3
R8066 commonsourceibias.n140 commonsourceibias.n123 161.3
R8067 commonsourceibias.n142 commonsourceibias.n141 161.3
R8068 commonsourceibias.n144 commonsourceibias.n143 161.3
R8069 commonsourceibias.n145 commonsourceibias.n121 161.3
R8070 commonsourceibias.n147 commonsourceibias.n146 161.3
R8071 commonsourceibias.n149 commonsourceibias.n148 161.3
R8072 commonsourceibias.n150 commonsourceibias.n119 161.3
R8073 commonsourceibias.n152 commonsourceibias.n151 161.3
R8074 commonsourceibias.n154 commonsourceibias.n153 161.3
R8075 commonsourceibias.n155 commonsourceibias.n117 161.3
R8076 commonsourceibias.n158 commonsourceibias.n157 161.3
R8077 commonsourceibias.n159 commonsourceibias.n11 161.3
R8078 commonsourceibias.n161 commonsourceibias.n160 161.3
R8079 commonsourceibias.n163 commonsourceibias.n9 161.3
R8080 commonsourceibias.n165 commonsourceibias.n164 161.3
R8081 commonsourceibias.n166 commonsourceibias.n8 161.3
R8082 commonsourceibias.n168 commonsourceibias.n167 161.3
R8083 commonsourceibias.n169 commonsourceibias.n7 161.3
R8084 commonsourceibias.n172 commonsourceibias.n171 161.3
R8085 commonsourceibias.n173 commonsourceibias.n6 161.3
R8086 commonsourceibias.n175 commonsourceibias.n174 161.3
R8087 commonsourceibias.n177 commonsourceibias.n4 161.3
R8088 commonsourceibias.n179 commonsourceibias.n178 161.3
R8089 commonsourceibias.n180 commonsourceibias.n3 161.3
R8090 commonsourceibias.n182 commonsourceibias.n181 161.3
R8091 commonsourceibias.n183 commonsourceibias.n2 161.3
R8092 commonsourceibias.n186 commonsourceibias.n185 161.3
R8093 commonsourceibias.n187 commonsourceibias.n1 161.3
R8094 commonsourceibias.n189 commonsourceibias.n188 161.3
R8095 commonsourceibias.n191 commonsourceibias.n0 161.3
R8096 commonsourceibias.n280 commonsourceibias.n194 161.3
R8097 commonsourceibias.n278 commonsourceibias.n277 161.3
R8098 commonsourceibias.n276 commonsourceibias.n195 161.3
R8099 commonsourceibias.n275 commonsourceibias.n274 161.3
R8100 commonsourceibias.n272 commonsourceibias.n196 161.3
R8101 commonsourceibias.n271 commonsourceibias.n270 161.3
R8102 commonsourceibias.n269 commonsourceibias.n197 161.3
R8103 commonsourceibias.n268 commonsourceibias.n267 161.3
R8104 commonsourceibias.n266 commonsourceibias.n198 161.3
R8105 commonsourceibias.n264 commonsourceibias.n263 161.3
R8106 commonsourceibias.n262 commonsourceibias.n200 161.3
R8107 commonsourceibias.n261 commonsourceibias.n260 161.3
R8108 commonsourceibias.n258 commonsourceibias.n201 161.3
R8109 commonsourceibias.n257 commonsourceibias.n256 161.3
R8110 commonsourceibias.n255 commonsourceibias.n202 161.3
R8111 commonsourceibias.n254 commonsourceibias.n253 161.3
R8112 commonsourceibias.n252 commonsourceibias.n203 161.3
R8113 commonsourceibias.n250 commonsourceibias.n249 161.3
R8114 commonsourceibias.n248 commonsourceibias.n205 161.3
R8115 commonsourceibias.n247 commonsourceibias.n246 161.3
R8116 commonsourceibias.n244 commonsourceibias.n206 161.3
R8117 commonsourceibias.n243 commonsourceibias.n242 161.3
R8118 commonsourceibias.n241 commonsourceibias.n240 161.3
R8119 commonsourceibias.n239 commonsourceibias.n208 161.3
R8120 commonsourceibias.n238 commonsourceibias.n237 161.3
R8121 commonsourceibias.n236 commonsourceibias.n235 161.3
R8122 commonsourceibias.n234 commonsourceibias.n210 161.3
R8123 commonsourceibias.n233 commonsourceibias.n232 161.3
R8124 commonsourceibias.n231 commonsourceibias.n230 161.3
R8125 commonsourceibias.n229 commonsourceibias.n212 161.3
R8126 commonsourceibias.n227 commonsourceibias.n226 161.3
R8127 commonsourceibias.n225 commonsourceibias.n213 161.3
R8128 commonsourceibias.n224 commonsourceibias.n223 161.3
R8129 commonsourceibias.n221 commonsourceibias.n214 161.3
R8130 commonsourceibias.n220 commonsourceibias.n219 161.3
R8131 commonsourceibias.n218 commonsourceibias.n215 161.3
R8132 commonsourceibias.n429 commonsourceibias.n343 161.3
R8133 commonsourceibias.n427 commonsourceibias.n426 161.3
R8134 commonsourceibias.n425 commonsourceibias.n344 161.3
R8135 commonsourceibias.n424 commonsourceibias.n423 161.3
R8136 commonsourceibias.n421 commonsourceibias.n345 161.3
R8137 commonsourceibias.n420 commonsourceibias.n419 161.3
R8138 commonsourceibias.n418 commonsourceibias.n346 161.3
R8139 commonsourceibias.n417 commonsourceibias.n416 161.3
R8140 commonsourceibias.n414 commonsourceibias.n347 161.3
R8141 commonsourceibias.n412 commonsourceibias.n411 161.3
R8142 commonsourceibias.n410 commonsourceibias.n348 161.3
R8143 commonsourceibias.n409 commonsourceibias.n408 161.3
R8144 commonsourceibias.n406 commonsourceibias.n349 161.3
R8145 commonsourceibias.n405 commonsourceibias.n404 161.3
R8146 commonsourceibias.n403 commonsourceibias.n350 161.3
R8147 commonsourceibias.n402 commonsourceibias.n401 161.3
R8148 commonsourceibias.n399 commonsourceibias.n351 161.3
R8149 commonsourceibias.n397 commonsourceibias.n396 161.3
R8150 commonsourceibias.n395 commonsourceibias.n352 161.3
R8151 commonsourceibias.n394 commonsourceibias.n393 161.3
R8152 commonsourceibias.n391 commonsourceibias.n353 161.3
R8153 commonsourceibias.n390 commonsourceibias.n389 161.3
R8154 commonsourceibias.n388 commonsourceibias.n387 161.3
R8155 commonsourceibias.n386 commonsourceibias.n355 161.3
R8156 commonsourceibias.n385 commonsourceibias.n384 161.3
R8157 commonsourceibias.n383 commonsourceibias.n382 161.3
R8158 commonsourceibias.n381 commonsourceibias.n357 161.3
R8159 commonsourceibias.n380 commonsourceibias.n379 161.3
R8160 commonsourceibias.n378 commonsourceibias.n377 161.3
R8161 commonsourceibias.n376 commonsourceibias.n359 161.3
R8162 commonsourceibias.n374 commonsourceibias.n373 161.3
R8163 commonsourceibias.n372 commonsourceibias.n360 161.3
R8164 commonsourceibias.n371 commonsourceibias.n370 161.3
R8165 commonsourceibias.n368 commonsourceibias.n361 161.3
R8166 commonsourceibias.n367 commonsourceibias.n366 161.3
R8167 commonsourceibias.n365 commonsourceibias.n362 161.3
R8168 commonsourceibias.n335 commonsourceibias.n334 161.3
R8169 commonsourceibias.n332 commonsourceibias.n294 161.3
R8170 commonsourceibias.n331 commonsourceibias.n330 161.3
R8171 commonsourceibias.n329 commonsourceibias.n328 161.3
R8172 commonsourceibias.n327 commonsourceibias.n296 161.3
R8173 commonsourceibias.n326 commonsourceibias.n325 161.3
R8174 commonsourceibias.n324 commonsourceibias.n323 161.3
R8175 commonsourceibias.n322 commonsourceibias.n298 161.3
R8176 commonsourceibias.n321 commonsourceibias.n320 161.3
R8177 commonsourceibias.n319 commonsourceibias.n318 161.3
R8178 commonsourceibias.n317 commonsourceibias.n300 161.3
R8179 commonsourceibias.n315 commonsourceibias.n314 161.3
R8180 commonsourceibias.n313 commonsourceibias.n301 161.3
R8181 commonsourceibias.n312 commonsourceibias.n311 161.3
R8182 commonsourceibias.n309 commonsourceibias.n302 161.3
R8183 commonsourceibias.n308 commonsourceibias.n307 161.3
R8184 commonsourceibias.n306 commonsourceibias.n303 161.3
R8185 commonsourceibias.n441 commonsourceibias.n293 161.3
R8186 commonsourceibias.n475 commonsourceibias.n284 161.3
R8187 commonsourceibias.n473 commonsourceibias.n472 161.3
R8188 commonsourceibias.n471 commonsourceibias.n285 161.3
R8189 commonsourceibias.n470 commonsourceibias.n469 161.3
R8190 commonsourceibias.n467 commonsourceibias.n286 161.3
R8191 commonsourceibias.n466 commonsourceibias.n465 161.3
R8192 commonsourceibias.n464 commonsourceibias.n287 161.3
R8193 commonsourceibias.n463 commonsourceibias.n462 161.3
R8194 commonsourceibias.n460 commonsourceibias.n288 161.3
R8195 commonsourceibias.n458 commonsourceibias.n457 161.3
R8196 commonsourceibias.n456 commonsourceibias.n289 161.3
R8197 commonsourceibias.n455 commonsourceibias.n454 161.3
R8198 commonsourceibias.n452 commonsourceibias.n290 161.3
R8199 commonsourceibias.n451 commonsourceibias.n450 161.3
R8200 commonsourceibias.n449 commonsourceibias.n291 161.3
R8201 commonsourceibias.n448 commonsourceibias.n447 161.3
R8202 commonsourceibias.n445 commonsourceibias.n292 161.3
R8203 commonsourceibias.n443 commonsourceibias.n442 161.3
R8204 commonsourceibias.n564 commonsourceibias.n478 161.3
R8205 commonsourceibias.n562 commonsourceibias.n561 161.3
R8206 commonsourceibias.n560 commonsourceibias.n479 161.3
R8207 commonsourceibias.n559 commonsourceibias.n558 161.3
R8208 commonsourceibias.n556 commonsourceibias.n480 161.3
R8209 commonsourceibias.n555 commonsourceibias.n554 161.3
R8210 commonsourceibias.n553 commonsourceibias.n481 161.3
R8211 commonsourceibias.n552 commonsourceibias.n551 161.3
R8212 commonsourceibias.n549 commonsourceibias.n482 161.3
R8213 commonsourceibias.n547 commonsourceibias.n546 161.3
R8214 commonsourceibias.n545 commonsourceibias.n483 161.3
R8215 commonsourceibias.n544 commonsourceibias.n543 161.3
R8216 commonsourceibias.n541 commonsourceibias.n484 161.3
R8217 commonsourceibias.n540 commonsourceibias.n539 161.3
R8218 commonsourceibias.n538 commonsourceibias.n485 161.3
R8219 commonsourceibias.n537 commonsourceibias.n536 161.3
R8220 commonsourceibias.n534 commonsourceibias.n486 161.3
R8221 commonsourceibias.n532 commonsourceibias.n531 161.3
R8222 commonsourceibias.n530 commonsourceibias.n487 161.3
R8223 commonsourceibias.n529 commonsourceibias.n528 161.3
R8224 commonsourceibias.n526 commonsourceibias.n488 161.3
R8225 commonsourceibias.n525 commonsourceibias.n524 161.3
R8226 commonsourceibias.n523 commonsourceibias.n522 161.3
R8227 commonsourceibias.n521 commonsourceibias.n490 161.3
R8228 commonsourceibias.n520 commonsourceibias.n519 161.3
R8229 commonsourceibias.n518 commonsourceibias.n517 161.3
R8230 commonsourceibias.n516 commonsourceibias.n492 161.3
R8231 commonsourceibias.n515 commonsourceibias.n514 161.3
R8232 commonsourceibias.n513 commonsourceibias.n512 161.3
R8233 commonsourceibias.n511 commonsourceibias.n494 161.3
R8234 commonsourceibias.n509 commonsourceibias.n508 161.3
R8235 commonsourceibias.n507 commonsourceibias.n495 161.3
R8236 commonsourceibias.n506 commonsourceibias.n505 161.3
R8237 commonsourceibias.n503 commonsourceibias.n496 161.3
R8238 commonsourceibias.n502 commonsourceibias.n501 161.3
R8239 commonsourceibias.n500 commonsourceibias.n497 161.3
R8240 commonsourceibias.n111 commonsourceibias.n109 81.5057
R8241 commonsourceibias.n338 commonsourceibias.n336 81.5057
R8242 commonsourceibias.n111 commonsourceibias.n110 80.9324
R8243 commonsourceibias.n113 commonsourceibias.n112 80.9324
R8244 commonsourceibias.n115 commonsourceibias.n114 80.9324
R8245 commonsourceibias.n108 commonsourceibias.n107 80.9324
R8246 commonsourceibias.n106 commonsourceibias.n105 80.9324
R8247 commonsourceibias.n104 commonsourceibias.n103 80.9324
R8248 commonsourceibias.n102 commonsourceibias.n101 80.9324
R8249 commonsourceibias.n433 commonsourceibias.n432 80.9324
R8250 commonsourceibias.n435 commonsourceibias.n434 80.9324
R8251 commonsourceibias.n437 commonsourceibias.n436 80.9324
R8252 commonsourceibias.n439 commonsourceibias.n438 80.9324
R8253 commonsourceibias.n342 commonsourceibias.n341 80.9324
R8254 commonsourceibias.n340 commonsourceibias.n339 80.9324
R8255 commonsourceibias.n338 commonsourceibias.n337 80.9324
R8256 commonsourceibias.n100 commonsourceibias.n99 80.6037
R8257 commonsourceibias.n193 commonsourceibias.n192 80.6037
R8258 commonsourceibias.n282 commonsourceibias.n281 80.6037
R8259 commonsourceibias.n431 commonsourceibias.n430 80.6037
R8260 commonsourceibias.n477 commonsourceibias.n476 80.6037
R8261 commonsourceibias.n566 commonsourceibias.n565 80.6037
R8262 commonsourceibias.n85 commonsourceibias.n84 56.5617
R8263 commonsourceibias.n71 commonsourceibias.n70 56.5617
R8264 commonsourceibias.n62 commonsourceibias.n61 56.5617
R8265 commonsourceibias.n48 commonsourceibias.n47 56.5617
R8266 commonsourceibias.n178 commonsourceibias.n177 56.5617
R8267 commonsourceibias.n164 commonsourceibias.n163 56.5617
R8268 commonsourceibias.n155 commonsourceibias.n154 56.5617
R8269 commonsourceibias.n141 commonsourceibias.n140 56.5617
R8270 commonsourceibias.n230 commonsourceibias.n229 56.5617
R8271 commonsourceibias.n244 commonsourceibias.n243 56.5617
R8272 commonsourceibias.n253 commonsourceibias.n252 56.5617
R8273 commonsourceibias.n267 commonsourceibias.n266 56.5617
R8274 commonsourceibias.n377 commonsourceibias.n376 56.5617
R8275 commonsourceibias.n391 commonsourceibias.n390 56.5617
R8276 commonsourceibias.n401 commonsourceibias.n399 56.5617
R8277 commonsourceibias.n416 commonsourceibias.n414 56.5617
R8278 commonsourceibias.n462 commonsourceibias.n460 56.5617
R8279 commonsourceibias.n447 commonsourceibias.n445 56.5617
R8280 commonsourceibias.n318 commonsourceibias.n317 56.5617
R8281 commonsourceibias.n332 commonsourceibias.n331 56.5617
R8282 commonsourceibias.n512 commonsourceibias.n511 56.5617
R8283 commonsourceibias.n526 commonsourceibias.n525 56.5617
R8284 commonsourceibias.n536 commonsourceibias.n534 56.5617
R8285 commonsourceibias.n551 commonsourceibias.n549 56.5617
R8286 commonsourceibias.n76 commonsourceibias.n75 56.0773
R8287 commonsourceibias.n57 commonsourceibias.n56 56.0773
R8288 commonsourceibias.n169 commonsourceibias.n168 56.0773
R8289 commonsourceibias.n150 commonsourceibias.n149 56.0773
R8290 commonsourceibias.n239 commonsourceibias.n238 56.0773
R8291 commonsourceibias.n258 commonsourceibias.n257 56.0773
R8292 commonsourceibias.n386 commonsourceibias.n385 56.0773
R8293 commonsourceibias.n406 commonsourceibias.n405 56.0773
R8294 commonsourceibias.n452 commonsourceibias.n451 56.0773
R8295 commonsourceibias.n327 commonsourceibias.n326 56.0773
R8296 commonsourceibias.n521 commonsourceibias.n520 56.0773
R8297 commonsourceibias.n541 commonsourceibias.n540 56.0773
R8298 commonsourceibias.n99 commonsourceibias.n98 55.3321
R8299 commonsourceibias.n192 commonsourceibias.n191 55.3321
R8300 commonsourceibias.n281 commonsourceibias.n280 55.3321
R8301 commonsourceibias.n430 commonsourceibias.n429 55.3321
R8302 commonsourceibias.n476 commonsourceibias.n475 55.3321
R8303 commonsourceibias.n565 commonsourceibias.n564 55.3321
R8304 commonsourceibias.n90 commonsourceibias.n89 55.1086
R8305 commonsourceibias.n41 commonsourceibias.n31 55.1086
R8306 commonsourceibias.n183 commonsourceibias.n182 55.1086
R8307 commonsourceibias.n134 commonsourceibias.n124 55.1086
R8308 commonsourceibias.n223 commonsourceibias.n213 55.1086
R8309 commonsourceibias.n272 commonsourceibias.n271 55.1086
R8310 commonsourceibias.n370 commonsourceibias.n360 55.1086
R8311 commonsourceibias.n421 commonsourceibias.n420 55.1086
R8312 commonsourceibias.n467 commonsourceibias.n466 55.1086
R8313 commonsourceibias.n311 commonsourceibias.n301 55.1086
R8314 commonsourceibias.n505 commonsourceibias.n495 55.1086
R8315 commonsourceibias.n556 commonsourceibias.n555 55.1086
R8316 commonsourceibias.n35 commonsourceibias.n34 47.4592
R8317 commonsourceibias.n128 commonsourceibias.n127 47.4592
R8318 commonsourceibias.n217 commonsourceibias.n216 47.4592
R8319 commonsourceibias.n364 commonsourceibias.n363 47.4592
R8320 commonsourceibias.n305 commonsourceibias.n304 47.4592
R8321 commonsourceibias.n499 commonsourceibias.n498 47.4592
R8322 commonsourceibias.n218 commonsourceibias.n217 44.0436
R8323 commonsourceibias.n365 commonsourceibias.n364 44.0436
R8324 commonsourceibias.n306 commonsourceibias.n305 44.0436
R8325 commonsourceibias.n500 commonsourceibias.n499 44.0436
R8326 commonsourceibias.n36 commonsourceibias.n35 44.0436
R8327 commonsourceibias.n129 commonsourceibias.n128 44.0436
R8328 commonsourceibias.n92 commonsourceibias.n13 42.5146
R8329 commonsourceibias.n39 commonsourceibias.n38 42.5146
R8330 commonsourceibias.n185 commonsourceibias.n1 42.5146
R8331 commonsourceibias.n132 commonsourceibias.n131 42.5146
R8332 commonsourceibias.n221 commonsourceibias.n220 42.5146
R8333 commonsourceibias.n274 commonsourceibias.n195 42.5146
R8334 commonsourceibias.n368 commonsourceibias.n367 42.5146
R8335 commonsourceibias.n423 commonsourceibias.n344 42.5146
R8336 commonsourceibias.n469 commonsourceibias.n285 42.5146
R8337 commonsourceibias.n309 commonsourceibias.n308 42.5146
R8338 commonsourceibias.n503 commonsourceibias.n502 42.5146
R8339 commonsourceibias.n558 commonsourceibias.n479 42.5146
R8340 commonsourceibias.n78 commonsourceibias.n18 41.5458
R8341 commonsourceibias.n53 commonsourceibias.n52 41.5458
R8342 commonsourceibias.n171 commonsourceibias.n6 41.5458
R8343 commonsourceibias.n146 commonsourceibias.n145 41.5458
R8344 commonsourceibias.n235 commonsourceibias.n234 41.5458
R8345 commonsourceibias.n260 commonsourceibias.n200 41.5458
R8346 commonsourceibias.n382 commonsourceibias.n381 41.5458
R8347 commonsourceibias.n408 commonsourceibias.n348 41.5458
R8348 commonsourceibias.n454 commonsourceibias.n289 41.5458
R8349 commonsourceibias.n323 commonsourceibias.n322 41.5458
R8350 commonsourceibias.n517 commonsourceibias.n516 41.5458
R8351 commonsourceibias.n543 commonsourceibias.n483 41.5458
R8352 commonsourceibias.n68 commonsourceibias.n23 40.577
R8353 commonsourceibias.n64 commonsourceibias.n23 40.577
R8354 commonsourceibias.n161 commonsourceibias.n11 40.577
R8355 commonsourceibias.n157 commonsourceibias.n11 40.577
R8356 commonsourceibias.n246 commonsourceibias.n205 40.577
R8357 commonsourceibias.n250 commonsourceibias.n205 40.577
R8358 commonsourceibias.n393 commonsourceibias.n352 40.577
R8359 commonsourceibias.n397 commonsourceibias.n352 40.577
R8360 commonsourceibias.n443 commonsourceibias.n293 40.577
R8361 commonsourceibias.n334 commonsourceibias.n293 40.577
R8362 commonsourceibias.n528 commonsourceibias.n487 40.577
R8363 commonsourceibias.n532 commonsourceibias.n487 40.577
R8364 commonsourceibias.n82 commonsourceibias.n18 39.6083
R8365 commonsourceibias.n52 commonsourceibias.n51 39.6083
R8366 commonsourceibias.n175 commonsourceibias.n6 39.6083
R8367 commonsourceibias.n145 commonsourceibias.n144 39.6083
R8368 commonsourceibias.n234 commonsourceibias.n233 39.6083
R8369 commonsourceibias.n264 commonsourceibias.n200 39.6083
R8370 commonsourceibias.n381 commonsourceibias.n380 39.6083
R8371 commonsourceibias.n412 commonsourceibias.n348 39.6083
R8372 commonsourceibias.n458 commonsourceibias.n289 39.6083
R8373 commonsourceibias.n322 commonsourceibias.n321 39.6083
R8374 commonsourceibias.n516 commonsourceibias.n515 39.6083
R8375 commonsourceibias.n547 commonsourceibias.n483 39.6083
R8376 commonsourceibias.n96 commonsourceibias.n13 38.6395
R8377 commonsourceibias.n38 commonsourceibias.n33 38.6395
R8378 commonsourceibias.n189 commonsourceibias.n1 38.6395
R8379 commonsourceibias.n131 commonsourceibias.n126 38.6395
R8380 commonsourceibias.n220 commonsourceibias.n215 38.6395
R8381 commonsourceibias.n278 commonsourceibias.n195 38.6395
R8382 commonsourceibias.n367 commonsourceibias.n362 38.6395
R8383 commonsourceibias.n427 commonsourceibias.n344 38.6395
R8384 commonsourceibias.n473 commonsourceibias.n285 38.6395
R8385 commonsourceibias.n308 commonsourceibias.n303 38.6395
R8386 commonsourceibias.n502 commonsourceibias.n497 38.6395
R8387 commonsourceibias.n562 commonsourceibias.n479 38.6395
R8388 commonsourceibias.n89 commonsourceibias.n15 26.0455
R8389 commonsourceibias.n45 commonsourceibias.n31 26.0455
R8390 commonsourceibias.n182 commonsourceibias.n3 26.0455
R8391 commonsourceibias.n138 commonsourceibias.n124 26.0455
R8392 commonsourceibias.n227 commonsourceibias.n213 26.0455
R8393 commonsourceibias.n271 commonsourceibias.n197 26.0455
R8394 commonsourceibias.n374 commonsourceibias.n360 26.0455
R8395 commonsourceibias.n420 commonsourceibias.n346 26.0455
R8396 commonsourceibias.n466 commonsourceibias.n287 26.0455
R8397 commonsourceibias.n315 commonsourceibias.n301 26.0455
R8398 commonsourceibias.n509 commonsourceibias.n495 26.0455
R8399 commonsourceibias.n555 commonsourceibias.n481 26.0455
R8400 commonsourceibias.n75 commonsourceibias.n20 25.0767
R8401 commonsourceibias.n58 commonsourceibias.n57 25.0767
R8402 commonsourceibias.n168 commonsourceibias.n8 25.0767
R8403 commonsourceibias.n151 commonsourceibias.n150 25.0767
R8404 commonsourceibias.n240 commonsourceibias.n239 25.0767
R8405 commonsourceibias.n257 commonsourceibias.n202 25.0767
R8406 commonsourceibias.n387 commonsourceibias.n386 25.0767
R8407 commonsourceibias.n405 commonsourceibias.n350 25.0767
R8408 commonsourceibias.n451 commonsourceibias.n291 25.0767
R8409 commonsourceibias.n328 commonsourceibias.n327 25.0767
R8410 commonsourceibias.n522 commonsourceibias.n521 25.0767
R8411 commonsourceibias.n540 commonsourceibias.n485 25.0767
R8412 commonsourceibias.n71 commonsourceibias.n22 24.3464
R8413 commonsourceibias.n61 commonsourceibias.n25 24.3464
R8414 commonsourceibias.n164 commonsourceibias.n10 24.3464
R8415 commonsourceibias.n154 commonsourceibias.n118 24.3464
R8416 commonsourceibias.n243 commonsourceibias.n207 24.3464
R8417 commonsourceibias.n253 commonsourceibias.n204 24.3464
R8418 commonsourceibias.n390 commonsourceibias.n354 24.3464
R8419 commonsourceibias.n401 commonsourceibias.n400 24.3464
R8420 commonsourceibias.n447 commonsourceibias.n446 24.3464
R8421 commonsourceibias.n331 commonsourceibias.n295 24.3464
R8422 commonsourceibias.n525 commonsourceibias.n489 24.3464
R8423 commonsourceibias.n536 commonsourceibias.n535 24.3464
R8424 commonsourceibias.n85 commonsourceibias.n17 23.8546
R8425 commonsourceibias.n47 commonsourceibias.n46 23.8546
R8426 commonsourceibias.n178 commonsourceibias.n5 23.8546
R8427 commonsourceibias.n140 commonsourceibias.n139 23.8546
R8428 commonsourceibias.n229 commonsourceibias.n228 23.8546
R8429 commonsourceibias.n267 commonsourceibias.n199 23.8546
R8430 commonsourceibias.n376 commonsourceibias.n375 23.8546
R8431 commonsourceibias.n416 commonsourceibias.n415 23.8546
R8432 commonsourceibias.n462 commonsourceibias.n461 23.8546
R8433 commonsourceibias.n317 commonsourceibias.n316 23.8546
R8434 commonsourceibias.n511 commonsourceibias.n510 23.8546
R8435 commonsourceibias.n551 commonsourceibias.n550 23.8546
R8436 commonsourceibias.n98 commonsourceibias.n97 17.4607
R8437 commonsourceibias.n191 commonsourceibias.n190 17.4607
R8438 commonsourceibias.n280 commonsourceibias.n279 17.4607
R8439 commonsourceibias.n429 commonsourceibias.n428 17.4607
R8440 commonsourceibias.n475 commonsourceibias.n474 17.4607
R8441 commonsourceibias.n564 commonsourceibias.n563 17.4607
R8442 commonsourceibias.n84 commonsourceibias.n83 16.9689
R8443 commonsourceibias.n48 commonsourceibias.n29 16.9689
R8444 commonsourceibias.n177 commonsourceibias.n176 16.9689
R8445 commonsourceibias.n141 commonsourceibias.n122 16.9689
R8446 commonsourceibias.n230 commonsourceibias.n211 16.9689
R8447 commonsourceibias.n266 commonsourceibias.n265 16.9689
R8448 commonsourceibias.n377 commonsourceibias.n358 16.9689
R8449 commonsourceibias.n414 commonsourceibias.n413 16.9689
R8450 commonsourceibias.n460 commonsourceibias.n459 16.9689
R8451 commonsourceibias.n318 commonsourceibias.n299 16.9689
R8452 commonsourceibias.n512 commonsourceibias.n493 16.9689
R8453 commonsourceibias.n549 commonsourceibias.n548 16.9689
R8454 commonsourceibias.n70 commonsourceibias.n69 16.477
R8455 commonsourceibias.n63 commonsourceibias.n62 16.477
R8456 commonsourceibias.n163 commonsourceibias.n162 16.477
R8457 commonsourceibias.n156 commonsourceibias.n155 16.477
R8458 commonsourceibias.n245 commonsourceibias.n244 16.477
R8459 commonsourceibias.n252 commonsourceibias.n251 16.477
R8460 commonsourceibias.n392 commonsourceibias.n391 16.477
R8461 commonsourceibias.n399 commonsourceibias.n398 16.477
R8462 commonsourceibias.n445 commonsourceibias.n444 16.477
R8463 commonsourceibias.n333 commonsourceibias.n332 16.477
R8464 commonsourceibias.n527 commonsourceibias.n526 16.477
R8465 commonsourceibias.n534 commonsourceibias.n533 16.477
R8466 commonsourceibias.n77 commonsourceibias.n76 15.9852
R8467 commonsourceibias.n56 commonsourceibias.n27 15.9852
R8468 commonsourceibias.n170 commonsourceibias.n169 15.9852
R8469 commonsourceibias.n149 commonsourceibias.n120 15.9852
R8470 commonsourceibias.n238 commonsourceibias.n209 15.9852
R8471 commonsourceibias.n259 commonsourceibias.n258 15.9852
R8472 commonsourceibias.n385 commonsourceibias.n356 15.9852
R8473 commonsourceibias.n407 commonsourceibias.n406 15.9852
R8474 commonsourceibias.n453 commonsourceibias.n452 15.9852
R8475 commonsourceibias.n326 commonsourceibias.n297 15.9852
R8476 commonsourceibias.n520 commonsourceibias.n491 15.9852
R8477 commonsourceibias.n542 commonsourceibias.n541 15.9852
R8478 commonsourceibias.n91 commonsourceibias.n90 15.4934
R8479 commonsourceibias.n41 commonsourceibias.n40 15.4934
R8480 commonsourceibias.n184 commonsourceibias.n183 15.4934
R8481 commonsourceibias.n134 commonsourceibias.n133 15.4934
R8482 commonsourceibias.n223 commonsourceibias.n222 15.4934
R8483 commonsourceibias.n273 commonsourceibias.n272 15.4934
R8484 commonsourceibias.n370 commonsourceibias.n369 15.4934
R8485 commonsourceibias.n422 commonsourceibias.n421 15.4934
R8486 commonsourceibias.n468 commonsourceibias.n467 15.4934
R8487 commonsourceibias.n311 commonsourceibias.n310 15.4934
R8488 commonsourceibias.n505 commonsourceibias.n504 15.4934
R8489 commonsourceibias.n557 commonsourceibias.n556 15.4934
R8490 commonsourceibias.n102 commonsourceibias.n100 13.2663
R8491 commonsourceibias.n433 commonsourceibias.n431 13.2663
R8492 commonsourceibias.n568 commonsourceibias.n283 12.2777
R8493 commonsourceibias.n568 commonsourceibias.n567 10.3347
R8494 commonsourceibias.n159 commonsourceibias.n116 9.50363
R8495 commonsourceibias.n441 commonsourceibias.n440 9.50363
R8496 commonsourceibias.n92 commonsourceibias.n91 9.09948
R8497 commonsourceibias.n40 commonsourceibias.n39 9.09948
R8498 commonsourceibias.n185 commonsourceibias.n184 9.09948
R8499 commonsourceibias.n133 commonsourceibias.n132 9.09948
R8500 commonsourceibias.n222 commonsourceibias.n221 9.09948
R8501 commonsourceibias.n274 commonsourceibias.n273 9.09948
R8502 commonsourceibias.n369 commonsourceibias.n368 9.09948
R8503 commonsourceibias.n423 commonsourceibias.n422 9.09948
R8504 commonsourceibias.n469 commonsourceibias.n468 9.09948
R8505 commonsourceibias.n310 commonsourceibias.n309 9.09948
R8506 commonsourceibias.n504 commonsourceibias.n503 9.09948
R8507 commonsourceibias.n558 commonsourceibias.n557 9.09948
R8508 commonsourceibias.n283 commonsourceibias.n193 8.79261
R8509 commonsourceibias.n567 commonsourceibias.n477 8.79261
R8510 commonsourceibias.n78 commonsourceibias.n77 8.60764
R8511 commonsourceibias.n53 commonsourceibias.n27 8.60764
R8512 commonsourceibias.n171 commonsourceibias.n170 8.60764
R8513 commonsourceibias.n146 commonsourceibias.n120 8.60764
R8514 commonsourceibias.n235 commonsourceibias.n209 8.60764
R8515 commonsourceibias.n260 commonsourceibias.n259 8.60764
R8516 commonsourceibias.n382 commonsourceibias.n356 8.60764
R8517 commonsourceibias.n408 commonsourceibias.n407 8.60764
R8518 commonsourceibias.n454 commonsourceibias.n453 8.60764
R8519 commonsourceibias.n323 commonsourceibias.n297 8.60764
R8520 commonsourceibias.n517 commonsourceibias.n491 8.60764
R8521 commonsourceibias.n543 commonsourceibias.n542 8.60764
R8522 commonsourceibias.n69 commonsourceibias.n68 8.11581
R8523 commonsourceibias.n64 commonsourceibias.n63 8.11581
R8524 commonsourceibias.n162 commonsourceibias.n161 8.11581
R8525 commonsourceibias.n157 commonsourceibias.n156 8.11581
R8526 commonsourceibias.n246 commonsourceibias.n245 8.11581
R8527 commonsourceibias.n251 commonsourceibias.n250 8.11581
R8528 commonsourceibias.n393 commonsourceibias.n392 8.11581
R8529 commonsourceibias.n398 commonsourceibias.n397 8.11581
R8530 commonsourceibias.n444 commonsourceibias.n443 8.11581
R8531 commonsourceibias.n334 commonsourceibias.n333 8.11581
R8532 commonsourceibias.n528 commonsourceibias.n527 8.11581
R8533 commonsourceibias.n533 commonsourceibias.n532 8.11581
R8534 commonsourceibias.n83 commonsourceibias.n82 7.62397
R8535 commonsourceibias.n51 commonsourceibias.n29 7.62397
R8536 commonsourceibias.n176 commonsourceibias.n175 7.62397
R8537 commonsourceibias.n144 commonsourceibias.n122 7.62397
R8538 commonsourceibias.n233 commonsourceibias.n211 7.62397
R8539 commonsourceibias.n265 commonsourceibias.n264 7.62397
R8540 commonsourceibias.n380 commonsourceibias.n358 7.62397
R8541 commonsourceibias.n413 commonsourceibias.n412 7.62397
R8542 commonsourceibias.n459 commonsourceibias.n458 7.62397
R8543 commonsourceibias.n321 commonsourceibias.n299 7.62397
R8544 commonsourceibias.n515 commonsourceibias.n493 7.62397
R8545 commonsourceibias.n548 commonsourceibias.n547 7.62397
R8546 commonsourceibias.n97 commonsourceibias.n96 7.13213
R8547 commonsourceibias.n34 commonsourceibias.n33 7.13213
R8548 commonsourceibias.n190 commonsourceibias.n189 7.13213
R8549 commonsourceibias.n127 commonsourceibias.n126 7.13213
R8550 commonsourceibias.n216 commonsourceibias.n215 7.13213
R8551 commonsourceibias.n279 commonsourceibias.n278 7.13213
R8552 commonsourceibias.n363 commonsourceibias.n362 7.13213
R8553 commonsourceibias.n428 commonsourceibias.n427 7.13213
R8554 commonsourceibias.n474 commonsourceibias.n473 7.13213
R8555 commonsourceibias.n304 commonsourceibias.n303 7.13213
R8556 commonsourceibias.n498 commonsourceibias.n497 7.13213
R8557 commonsourceibias.n563 commonsourceibias.n562 7.13213
R8558 commonsourceibias.n283 commonsourceibias.n282 5.06534
R8559 commonsourceibias.n567 commonsourceibias.n566 5.06534
R8560 commonsourceibias commonsourceibias.n568 4.04308
R8561 commonsourceibias.n109 commonsourceibias.t15 2.82907
R8562 commonsourceibias.n109 commonsourceibias.t59 2.82907
R8563 commonsourceibias.n110 commonsourceibias.t53 2.82907
R8564 commonsourceibias.n110 commonsourceibias.t35 2.82907
R8565 commonsourceibias.n112 commonsourceibias.t37 2.82907
R8566 commonsourceibias.n112 commonsourceibias.t11 2.82907
R8567 commonsourceibias.n114 commonsourceibias.t23 2.82907
R8568 commonsourceibias.n114 commonsourceibias.t55 2.82907
R8569 commonsourceibias.n107 commonsourceibias.t9 2.82907
R8570 commonsourceibias.n107 commonsourceibias.t49 2.82907
R8571 commonsourceibias.n105 commonsourceibias.t51 2.82907
R8572 commonsourceibias.n105 commonsourceibias.t63 2.82907
R8573 commonsourceibias.n103 commonsourceibias.t1 2.82907
R8574 commonsourceibias.n103 commonsourceibias.t19 2.82907
R8575 commonsourceibias.n101 commonsourceibias.t61 2.82907
R8576 commonsourceibias.n101 commonsourceibias.t29 2.82907
R8577 commonsourceibias.n432 commonsourceibias.t57 2.82907
R8578 commonsourceibias.n432 commonsourceibias.t21 2.82907
R8579 commonsourceibias.n434 commonsourceibias.t13 2.82907
R8580 commonsourceibias.n434 commonsourceibias.t27 2.82907
R8581 commonsourceibias.n436 commonsourceibias.t17 2.82907
R8582 commonsourceibias.n436 commonsourceibias.t41 2.82907
R8583 commonsourceibias.n438 commonsourceibias.t39 2.82907
R8584 commonsourceibias.n438 commonsourceibias.t5 2.82907
R8585 commonsourceibias.n341 commonsourceibias.t45 2.82907
R8586 commonsourceibias.n341 commonsourceibias.t7 2.82907
R8587 commonsourceibias.n339 commonsourceibias.t3 2.82907
R8588 commonsourceibias.n339 commonsourceibias.t33 2.82907
R8589 commonsourceibias.n337 commonsourceibias.t25 2.82907
R8590 commonsourceibias.n337 commonsourceibias.t43 2.82907
R8591 commonsourceibias.n336 commonsourceibias.t31 2.82907
R8592 commonsourceibias.n336 commonsourceibias.t47 2.82907
R8593 commonsourceibias.n17 commonsourceibias.n15 0.738255
R8594 commonsourceibias.n46 commonsourceibias.n45 0.738255
R8595 commonsourceibias.n5 commonsourceibias.n3 0.738255
R8596 commonsourceibias.n139 commonsourceibias.n138 0.738255
R8597 commonsourceibias.n228 commonsourceibias.n227 0.738255
R8598 commonsourceibias.n199 commonsourceibias.n197 0.738255
R8599 commonsourceibias.n375 commonsourceibias.n374 0.738255
R8600 commonsourceibias.n415 commonsourceibias.n346 0.738255
R8601 commonsourceibias.n461 commonsourceibias.n287 0.738255
R8602 commonsourceibias.n316 commonsourceibias.n315 0.738255
R8603 commonsourceibias.n510 commonsourceibias.n509 0.738255
R8604 commonsourceibias.n550 commonsourceibias.n481 0.738255
R8605 commonsourceibias.n104 commonsourceibias.n102 0.573776
R8606 commonsourceibias.n106 commonsourceibias.n104 0.573776
R8607 commonsourceibias.n108 commonsourceibias.n106 0.573776
R8608 commonsourceibias.n115 commonsourceibias.n113 0.573776
R8609 commonsourceibias.n113 commonsourceibias.n111 0.573776
R8610 commonsourceibias.n340 commonsourceibias.n338 0.573776
R8611 commonsourceibias.n342 commonsourceibias.n340 0.573776
R8612 commonsourceibias.n439 commonsourceibias.n437 0.573776
R8613 commonsourceibias.n437 commonsourceibias.n435 0.573776
R8614 commonsourceibias.n435 commonsourceibias.n433 0.573776
R8615 commonsourceibias.n116 commonsourceibias.n108 0.287138
R8616 commonsourceibias.n116 commonsourceibias.n115 0.287138
R8617 commonsourceibias.n440 commonsourceibias.n342 0.287138
R8618 commonsourceibias.n440 commonsourceibias.n439 0.287138
R8619 commonsourceibias.n100 commonsourceibias.n12 0.285035
R8620 commonsourceibias.n193 commonsourceibias.n0 0.285035
R8621 commonsourceibias.n282 commonsourceibias.n194 0.285035
R8622 commonsourceibias.n431 commonsourceibias.n343 0.285035
R8623 commonsourceibias.n477 commonsourceibias.n284 0.285035
R8624 commonsourceibias.n566 commonsourceibias.n478 0.285035
R8625 commonsourceibias.n22 commonsourceibias.n20 0.246418
R8626 commonsourceibias.n58 commonsourceibias.n25 0.246418
R8627 commonsourceibias.n10 commonsourceibias.n8 0.246418
R8628 commonsourceibias.n151 commonsourceibias.n118 0.246418
R8629 commonsourceibias.n240 commonsourceibias.n207 0.246418
R8630 commonsourceibias.n204 commonsourceibias.n202 0.246418
R8631 commonsourceibias.n387 commonsourceibias.n354 0.246418
R8632 commonsourceibias.n400 commonsourceibias.n350 0.246418
R8633 commonsourceibias.n446 commonsourceibias.n291 0.246418
R8634 commonsourceibias.n328 commonsourceibias.n295 0.246418
R8635 commonsourceibias.n522 commonsourceibias.n489 0.246418
R8636 commonsourceibias.n535 commonsourceibias.n485 0.246418
R8637 commonsourceibias.n95 commonsourceibias.n12 0.189894
R8638 commonsourceibias.n95 commonsourceibias.n94 0.189894
R8639 commonsourceibias.n94 commonsourceibias.n93 0.189894
R8640 commonsourceibias.n93 commonsourceibias.n14 0.189894
R8641 commonsourceibias.n88 commonsourceibias.n14 0.189894
R8642 commonsourceibias.n88 commonsourceibias.n87 0.189894
R8643 commonsourceibias.n87 commonsourceibias.n86 0.189894
R8644 commonsourceibias.n86 commonsourceibias.n16 0.189894
R8645 commonsourceibias.n81 commonsourceibias.n16 0.189894
R8646 commonsourceibias.n81 commonsourceibias.n80 0.189894
R8647 commonsourceibias.n80 commonsourceibias.n79 0.189894
R8648 commonsourceibias.n79 commonsourceibias.n19 0.189894
R8649 commonsourceibias.n74 commonsourceibias.n19 0.189894
R8650 commonsourceibias.n74 commonsourceibias.n73 0.189894
R8651 commonsourceibias.n73 commonsourceibias.n72 0.189894
R8652 commonsourceibias.n72 commonsourceibias.n21 0.189894
R8653 commonsourceibias.n67 commonsourceibias.n21 0.189894
R8654 commonsourceibias.n67 commonsourceibias.n66 0.189894
R8655 commonsourceibias.n66 commonsourceibias.n65 0.189894
R8656 commonsourceibias.n65 commonsourceibias.n24 0.189894
R8657 commonsourceibias.n60 commonsourceibias.n24 0.189894
R8658 commonsourceibias.n60 commonsourceibias.n59 0.189894
R8659 commonsourceibias.n59 commonsourceibias.n26 0.189894
R8660 commonsourceibias.n55 commonsourceibias.n26 0.189894
R8661 commonsourceibias.n55 commonsourceibias.n54 0.189894
R8662 commonsourceibias.n54 commonsourceibias.n28 0.189894
R8663 commonsourceibias.n50 commonsourceibias.n28 0.189894
R8664 commonsourceibias.n50 commonsourceibias.n49 0.189894
R8665 commonsourceibias.n49 commonsourceibias.n30 0.189894
R8666 commonsourceibias.n44 commonsourceibias.n30 0.189894
R8667 commonsourceibias.n44 commonsourceibias.n43 0.189894
R8668 commonsourceibias.n43 commonsourceibias.n42 0.189894
R8669 commonsourceibias.n42 commonsourceibias.n32 0.189894
R8670 commonsourceibias.n37 commonsourceibias.n32 0.189894
R8671 commonsourceibias.n37 commonsourceibias.n36 0.189894
R8672 commonsourceibias.n158 commonsourceibias.n117 0.189894
R8673 commonsourceibias.n153 commonsourceibias.n117 0.189894
R8674 commonsourceibias.n153 commonsourceibias.n152 0.189894
R8675 commonsourceibias.n152 commonsourceibias.n119 0.189894
R8676 commonsourceibias.n148 commonsourceibias.n119 0.189894
R8677 commonsourceibias.n148 commonsourceibias.n147 0.189894
R8678 commonsourceibias.n147 commonsourceibias.n121 0.189894
R8679 commonsourceibias.n143 commonsourceibias.n121 0.189894
R8680 commonsourceibias.n143 commonsourceibias.n142 0.189894
R8681 commonsourceibias.n142 commonsourceibias.n123 0.189894
R8682 commonsourceibias.n137 commonsourceibias.n123 0.189894
R8683 commonsourceibias.n137 commonsourceibias.n136 0.189894
R8684 commonsourceibias.n136 commonsourceibias.n135 0.189894
R8685 commonsourceibias.n135 commonsourceibias.n125 0.189894
R8686 commonsourceibias.n130 commonsourceibias.n125 0.189894
R8687 commonsourceibias.n130 commonsourceibias.n129 0.189894
R8688 commonsourceibias.n188 commonsourceibias.n0 0.189894
R8689 commonsourceibias.n188 commonsourceibias.n187 0.189894
R8690 commonsourceibias.n187 commonsourceibias.n186 0.189894
R8691 commonsourceibias.n186 commonsourceibias.n2 0.189894
R8692 commonsourceibias.n181 commonsourceibias.n2 0.189894
R8693 commonsourceibias.n181 commonsourceibias.n180 0.189894
R8694 commonsourceibias.n180 commonsourceibias.n179 0.189894
R8695 commonsourceibias.n179 commonsourceibias.n4 0.189894
R8696 commonsourceibias.n174 commonsourceibias.n4 0.189894
R8697 commonsourceibias.n174 commonsourceibias.n173 0.189894
R8698 commonsourceibias.n173 commonsourceibias.n172 0.189894
R8699 commonsourceibias.n172 commonsourceibias.n7 0.189894
R8700 commonsourceibias.n167 commonsourceibias.n7 0.189894
R8701 commonsourceibias.n167 commonsourceibias.n166 0.189894
R8702 commonsourceibias.n166 commonsourceibias.n165 0.189894
R8703 commonsourceibias.n165 commonsourceibias.n9 0.189894
R8704 commonsourceibias.n160 commonsourceibias.n9 0.189894
R8705 commonsourceibias.n277 commonsourceibias.n194 0.189894
R8706 commonsourceibias.n277 commonsourceibias.n276 0.189894
R8707 commonsourceibias.n276 commonsourceibias.n275 0.189894
R8708 commonsourceibias.n275 commonsourceibias.n196 0.189894
R8709 commonsourceibias.n270 commonsourceibias.n196 0.189894
R8710 commonsourceibias.n270 commonsourceibias.n269 0.189894
R8711 commonsourceibias.n269 commonsourceibias.n268 0.189894
R8712 commonsourceibias.n268 commonsourceibias.n198 0.189894
R8713 commonsourceibias.n263 commonsourceibias.n198 0.189894
R8714 commonsourceibias.n263 commonsourceibias.n262 0.189894
R8715 commonsourceibias.n262 commonsourceibias.n261 0.189894
R8716 commonsourceibias.n261 commonsourceibias.n201 0.189894
R8717 commonsourceibias.n256 commonsourceibias.n201 0.189894
R8718 commonsourceibias.n256 commonsourceibias.n255 0.189894
R8719 commonsourceibias.n255 commonsourceibias.n254 0.189894
R8720 commonsourceibias.n254 commonsourceibias.n203 0.189894
R8721 commonsourceibias.n249 commonsourceibias.n203 0.189894
R8722 commonsourceibias.n249 commonsourceibias.n248 0.189894
R8723 commonsourceibias.n248 commonsourceibias.n247 0.189894
R8724 commonsourceibias.n247 commonsourceibias.n206 0.189894
R8725 commonsourceibias.n242 commonsourceibias.n206 0.189894
R8726 commonsourceibias.n242 commonsourceibias.n241 0.189894
R8727 commonsourceibias.n241 commonsourceibias.n208 0.189894
R8728 commonsourceibias.n237 commonsourceibias.n208 0.189894
R8729 commonsourceibias.n237 commonsourceibias.n236 0.189894
R8730 commonsourceibias.n236 commonsourceibias.n210 0.189894
R8731 commonsourceibias.n232 commonsourceibias.n210 0.189894
R8732 commonsourceibias.n232 commonsourceibias.n231 0.189894
R8733 commonsourceibias.n231 commonsourceibias.n212 0.189894
R8734 commonsourceibias.n226 commonsourceibias.n212 0.189894
R8735 commonsourceibias.n226 commonsourceibias.n225 0.189894
R8736 commonsourceibias.n225 commonsourceibias.n224 0.189894
R8737 commonsourceibias.n224 commonsourceibias.n214 0.189894
R8738 commonsourceibias.n219 commonsourceibias.n214 0.189894
R8739 commonsourceibias.n219 commonsourceibias.n218 0.189894
R8740 commonsourceibias.n366 commonsourceibias.n365 0.189894
R8741 commonsourceibias.n366 commonsourceibias.n361 0.189894
R8742 commonsourceibias.n371 commonsourceibias.n361 0.189894
R8743 commonsourceibias.n372 commonsourceibias.n371 0.189894
R8744 commonsourceibias.n373 commonsourceibias.n372 0.189894
R8745 commonsourceibias.n373 commonsourceibias.n359 0.189894
R8746 commonsourceibias.n378 commonsourceibias.n359 0.189894
R8747 commonsourceibias.n379 commonsourceibias.n378 0.189894
R8748 commonsourceibias.n379 commonsourceibias.n357 0.189894
R8749 commonsourceibias.n383 commonsourceibias.n357 0.189894
R8750 commonsourceibias.n384 commonsourceibias.n383 0.189894
R8751 commonsourceibias.n384 commonsourceibias.n355 0.189894
R8752 commonsourceibias.n388 commonsourceibias.n355 0.189894
R8753 commonsourceibias.n389 commonsourceibias.n388 0.189894
R8754 commonsourceibias.n389 commonsourceibias.n353 0.189894
R8755 commonsourceibias.n394 commonsourceibias.n353 0.189894
R8756 commonsourceibias.n395 commonsourceibias.n394 0.189894
R8757 commonsourceibias.n396 commonsourceibias.n395 0.189894
R8758 commonsourceibias.n396 commonsourceibias.n351 0.189894
R8759 commonsourceibias.n402 commonsourceibias.n351 0.189894
R8760 commonsourceibias.n403 commonsourceibias.n402 0.189894
R8761 commonsourceibias.n404 commonsourceibias.n403 0.189894
R8762 commonsourceibias.n404 commonsourceibias.n349 0.189894
R8763 commonsourceibias.n409 commonsourceibias.n349 0.189894
R8764 commonsourceibias.n410 commonsourceibias.n409 0.189894
R8765 commonsourceibias.n411 commonsourceibias.n410 0.189894
R8766 commonsourceibias.n411 commonsourceibias.n347 0.189894
R8767 commonsourceibias.n417 commonsourceibias.n347 0.189894
R8768 commonsourceibias.n418 commonsourceibias.n417 0.189894
R8769 commonsourceibias.n419 commonsourceibias.n418 0.189894
R8770 commonsourceibias.n419 commonsourceibias.n345 0.189894
R8771 commonsourceibias.n424 commonsourceibias.n345 0.189894
R8772 commonsourceibias.n425 commonsourceibias.n424 0.189894
R8773 commonsourceibias.n426 commonsourceibias.n425 0.189894
R8774 commonsourceibias.n426 commonsourceibias.n343 0.189894
R8775 commonsourceibias.n307 commonsourceibias.n306 0.189894
R8776 commonsourceibias.n307 commonsourceibias.n302 0.189894
R8777 commonsourceibias.n312 commonsourceibias.n302 0.189894
R8778 commonsourceibias.n313 commonsourceibias.n312 0.189894
R8779 commonsourceibias.n314 commonsourceibias.n313 0.189894
R8780 commonsourceibias.n314 commonsourceibias.n300 0.189894
R8781 commonsourceibias.n319 commonsourceibias.n300 0.189894
R8782 commonsourceibias.n320 commonsourceibias.n319 0.189894
R8783 commonsourceibias.n320 commonsourceibias.n298 0.189894
R8784 commonsourceibias.n324 commonsourceibias.n298 0.189894
R8785 commonsourceibias.n325 commonsourceibias.n324 0.189894
R8786 commonsourceibias.n325 commonsourceibias.n296 0.189894
R8787 commonsourceibias.n329 commonsourceibias.n296 0.189894
R8788 commonsourceibias.n330 commonsourceibias.n329 0.189894
R8789 commonsourceibias.n330 commonsourceibias.n294 0.189894
R8790 commonsourceibias.n335 commonsourceibias.n294 0.189894
R8791 commonsourceibias.n442 commonsourceibias.n292 0.189894
R8792 commonsourceibias.n448 commonsourceibias.n292 0.189894
R8793 commonsourceibias.n449 commonsourceibias.n448 0.189894
R8794 commonsourceibias.n450 commonsourceibias.n449 0.189894
R8795 commonsourceibias.n450 commonsourceibias.n290 0.189894
R8796 commonsourceibias.n455 commonsourceibias.n290 0.189894
R8797 commonsourceibias.n456 commonsourceibias.n455 0.189894
R8798 commonsourceibias.n457 commonsourceibias.n456 0.189894
R8799 commonsourceibias.n457 commonsourceibias.n288 0.189894
R8800 commonsourceibias.n463 commonsourceibias.n288 0.189894
R8801 commonsourceibias.n464 commonsourceibias.n463 0.189894
R8802 commonsourceibias.n465 commonsourceibias.n464 0.189894
R8803 commonsourceibias.n465 commonsourceibias.n286 0.189894
R8804 commonsourceibias.n470 commonsourceibias.n286 0.189894
R8805 commonsourceibias.n471 commonsourceibias.n470 0.189894
R8806 commonsourceibias.n472 commonsourceibias.n471 0.189894
R8807 commonsourceibias.n472 commonsourceibias.n284 0.189894
R8808 commonsourceibias.n501 commonsourceibias.n500 0.189894
R8809 commonsourceibias.n501 commonsourceibias.n496 0.189894
R8810 commonsourceibias.n506 commonsourceibias.n496 0.189894
R8811 commonsourceibias.n507 commonsourceibias.n506 0.189894
R8812 commonsourceibias.n508 commonsourceibias.n507 0.189894
R8813 commonsourceibias.n508 commonsourceibias.n494 0.189894
R8814 commonsourceibias.n513 commonsourceibias.n494 0.189894
R8815 commonsourceibias.n514 commonsourceibias.n513 0.189894
R8816 commonsourceibias.n514 commonsourceibias.n492 0.189894
R8817 commonsourceibias.n518 commonsourceibias.n492 0.189894
R8818 commonsourceibias.n519 commonsourceibias.n518 0.189894
R8819 commonsourceibias.n519 commonsourceibias.n490 0.189894
R8820 commonsourceibias.n523 commonsourceibias.n490 0.189894
R8821 commonsourceibias.n524 commonsourceibias.n523 0.189894
R8822 commonsourceibias.n524 commonsourceibias.n488 0.189894
R8823 commonsourceibias.n529 commonsourceibias.n488 0.189894
R8824 commonsourceibias.n530 commonsourceibias.n529 0.189894
R8825 commonsourceibias.n531 commonsourceibias.n530 0.189894
R8826 commonsourceibias.n531 commonsourceibias.n486 0.189894
R8827 commonsourceibias.n537 commonsourceibias.n486 0.189894
R8828 commonsourceibias.n538 commonsourceibias.n537 0.189894
R8829 commonsourceibias.n539 commonsourceibias.n538 0.189894
R8830 commonsourceibias.n539 commonsourceibias.n484 0.189894
R8831 commonsourceibias.n544 commonsourceibias.n484 0.189894
R8832 commonsourceibias.n545 commonsourceibias.n544 0.189894
R8833 commonsourceibias.n546 commonsourceibias.n545 0.189894
R8834 commonsourceibias.n546 commonsourceibias.n482 0.189894
R8835 commonsourceibias.n552 commonsourceibias.n482 0.189894
R8836 commonsourceibias.n553 commonsourceibias.n552 0.189894
R8837 commonsourceibias.n554 commonsourceibias.n553 0.189894
R8838 commonsourceibias.n554 commonsourceibias.n480 0.189894
R8839 commonsourceibias.n559 commonsourceibias.n480 0.189894
R8840 commonsourceibias.n560 commonsourceibias.n559 0.189894
R8841 commonsourceibias.n561 commonsourceibias.n560 0.189894
R8842 commonsourceibias.n561 commonsourceibias.n478 0.189894
R8843 commonsourceibias.n159 commonsourceibias.n158 0.170955
R8844 commonsourceibias.n160 commonsourceibias.n159 0.170955
R8845 commonsourceibias.n441 commonsourceibias.n335 0.170955
R8846 commonsourceibias.n442 commonsourceibias.n441 0.170955
R8847 gnd.n6886 gnd.n454 1305.8
R8848 gnd.n4833 gnd.n4832 939.716
R8849 gnd.n7298 gnd.n107 795.207
R8850 gnd.n7462 gnd.n103 795.207
R8851 gnd.n1498 gnd.n1445 795.207
R8852 gnd.n4348 gnd.n1500 795.207
R8853 gnd.n4593 gnd.n1274 795.207
R8854 gnd.n3672 gnd.n1272 795.207
R8855 gnd.n2456 gnd.n960 795.207
R8856 gnd.n2518 gnd.n2457 795.207
R8857 gnd.n7460 gnd.n109 775.989
R8858 gnd.n177 gnd.n105 775.989
R8859 gnd.n4351 gnd.n4350 775.989
R8860 gnd.n4423 gnd.n1449 775.989
R8861 gnd.n4595 gnd.n1269 775.989
R8862 gnd.n2310 gnd.n1271 775.989
R8863 gnd.n4754 gnd.n4753 775.989
R8864 gnd.n4830 gnd.n964 775.989
R8865 gnd.n6238 gnd.n929 766.379
R8866 gnd.n6154 gnd.n931 766.379
R8867 gnd.n5342 gnd.n5245 766.379
R8868 gnd.n5338 gnd.n5243 766.379
R8869 gnd.n6235 gnd.n4835 756.769
R8870 gnd.n6204 gnd.n932 756.769
R8871 gnd.n5521 gnd.n5152 756.769
R8872 gnd.n5519 gnd.n5155 756.769
R8873 gnd.n3718 gnd.n1279 711.122
R8874 gnd.n4435 gnd.n1405 711.122
R8875 gnd.n3722 gnd.n2160 711.122
R8876 gnd.n4136 gnd.n1408 711.122
R8877 gnd.n6428 gnd.n727 670.282
R8878 gnd.n6885 gnd.n455 670.282
R8879 gnd.n7099 gnd.n7097 670.282
R8880 gnd.n2396 gnd.n895 670.282
R8881 gnd.n730 gnd.n727 585
R8882 gnd.n6426 gnd.n727 585
R8883 gnd.n6424 gnd.n6423 585
R8884 gnd.n6425 gnd.n6424 585
R8885 gnd.n6422 gnd.n729 585
R8886 gnd.n729 gnd.n728 585
R8887 gnd.n6421 gnd.n6420 585
R8888 gnd.n6420 gnd.n6419 585
R8889 gnd.n735 gnd.n734 585
R8890 gnd.n6418 gnd.n735 585
R8891 gnd.n6416 gnd.n6415 585
R8892 gnd.n6417 gnd.n6416 585
R8893 gnd.n6414 gnd.n737 585
R8894 gnd.n737 gnd.n736 585
R8895 gnd.n6413 gnd.n6412 585
R8896 gnd.n6412 gnd.n6411 585
R8897 gnd.n743 gnd.n742 585
R8898 gnd.n6410 gnd.n743 585
R8899 gnd.n6408 gnd.n6407 585
R8900 gnd.n6409 gnd.n6408 585
R8901 gnd.n6406 gnd.n745 585
R8902 gnd.n745 gnd.n744 585
R8903 gnd.n6405 gnd.n6404 585
R8904 gnd.n6404 gnd.n6403 585
R8905 gnd.n751 gnd.n750 585
R8906 gnd.n6402 gnd.n751 585
R8907 gnd.n6400 gnd.n6399 585
R8908 gnd.n6401 gnd.n6400 585
R8909 gnd.n6398 gnd.n753 585
R8910 gnd.n753 gnd.n752 585
R8911 gnd.n6397 gnd.n6396 585
R8912 gnd.n6396 gnd.n6395 585
R8913 gnd.n759 gnd.n758 585
R8914 gnd.n6394 gnd.n759 585
R8915 gnd.n6392 gnd.n6391 585
R8916 gnd.n6393 gnd.n6392 585
R8917 gnd.n6390 gnd.n761 585
R8918 gnd.n761 gnd.n760 585
R8919 gnd.n6389 gnd.n6388 585
R8920 gnd.n6388 gnd.n6387 585
R8921 gnd.n767 gnd.n766 585
R8922 gnd.n6386 gnd.n767 585
R8923 gnd.n6384 gnd.n6383 585
R8924 gnd.n6385 gnd.n6384 585
R8925 gnd.n6382 gnd.n769 585
R8926 gnd.n769 gnd.n768 585
R8927 gnd.n6381 gnd.n6380 585
R8928 gnd.n6380 gnd.n6379 585
R8929 gnd.n775 gnd.n774 585
R8930 gnd.n6378 gnd.n775 585
R8931 gnd.n6376 gnd.n6375 585
R8932 gnd.n6377 gnd.n6376 585
R8933 gnd.n6374 gnd.n777 585
R8934 gnd.n777 gnd.n776 585
R8935 gnd.n6373 gnd.n6372 585
R8936 gnd.n6372 gnd.n6371 585
R8937 gnd.n783 gnd.n782 585
R8938 gnd.n6370 gnd.n783 585
R8939 gnd.n6368 gnd.n6367 585
R8940 gnd.n6369 gnd.n6368 585
R8941 gnd.n6366 gnd.n785 585
R8942 gnd.n785 gnd.n784 585
R8943 gnd.n6365 gnd.n6364 585
R8944 gnd.n6364 gnd.n6363 585
R8945 gnd.n791 gnd.n790 585
R8946 gnd.n6362 gnd.n791 585
R8947 gnd.n6360 gnd.n6359 585
R8948 gnd.n6361 gnd.n6360 585
R8949 gnd.n6358 gnd.n793 585
R8950 gnd.n793 gnd.n792 585
R8951 gnd.n6357 gnd.n6356 585
R8952 gnd.n6356 gnd.n6355 585
R8953 gnd.n799 gnd.n798 585
R8954 gnd.n6354 gnd.n799 585
R8955 gnd.n6352 gnd.n6351 585
R8956 gnd.n6353 gnd.n6352 585
R8957 gnd.n6350 gnd.n801 585
R8958 gnd.n801 gnd.n800 585
R8959 gnd.n6349 gnd.n6348 585
R8960 gnd.n6348 gnd.n6347 585
R8961 gnd.n807 gnd.n806 585
R8962 gnd.n6346 gnd.n807 585
R8963 gnd.n6344 gnd.n6343 585
R8964 gnd.n6345 gnd.n6344 585
R8965 gnd.n6342 gnd.n809 585
R8966 gnd.n809 gnd.n808 585
R8967 gnd.n6341 gnd.n6340 585
R8968 gnd.n6340 gnd.n6339 585
R8969 gnd.n815 gnd.n814 585
R8970 gnd.n6338 gnd.n815 585
R8971 gnd.n6336 gnd.n6335 585
R8972 gnd.n6337 gnd.n6336 585
R8973 gnd.n6334 gnd.n817 585
R8974 gnd.n817 gnd.n816 585
R8975 gnd.n6333 gnd.n6332 585
R8976 gnd.n6332 gnd.n6331 585
R8977 gnd.n823 gnd.n822 585
R8978 gnd.n6330 gnd.n823 585
R8979 gnd.n6328 gnd.n6327 585
R8980 gnd.n6329 gnd.n6328 585
R8981 gnd.n6326 gnd.n825 585
R8982 gnd.n825 gnd.n824 585
R8983 gnd.n6325 gnd.n6324 585
R8984 gnd.n6324 gnd.n6323 585
R8985 gnd.n831 gnd.n830 585
R8986 gnd.n6322 gnd.n831 585
R8987 gnd.n6320 gnd.n6319 585
R8988 gnd.n6321 gnd.n6320 585
R8989 gnd.n6318 gnd.n833 585
R8990 gnd.n833 gnd.n832 585
R8991 gnd.n6317 gnd.n6316 585
R8992 gnd.n6316 gnd.n6315 585
R8993 gnd.n839 gnd.n838 585
R8994 gnd.n6314 gnd.n839 585
R8995 gnd.n6312 gnd.n6311 585
R8996 gnd.n6313 gnd.n6312 585
R8997 gnd.n6310 gnd.n841 585
R8998 gnd.n841 gnd.n840 585
R8999 gnd.n6309 gnd.n6308 585
R9000 gnd.n6308 gnd.n6307 585
R9001 gnd.n847 gnd.n846 585
R9002 gnd.n6306 gnd.n847 585
R9003 gnd.n6304 gnd.n6303 585
R9004 gnd.n6305 gnd.n6304 585
R9005 gnd.n6302 gnd.n849 585
R9006 gnd.n849 gnd.n848 585
R9007 gnd.n6301 gnd.n6300 585
R9008 gnd.n6300 gnd.n6299 585
R9009 gnd.n855 gnd.n854 585
R9010 gnd.n6298 gnd.n855 585
R9011 gnd.n6296 gnd.n6295 585
R9012 gnd.n6297 gnd.n6296 585
R9013 gnd.n6294 gnd.n857 585
R9014 gnd.n857 gnd.n856 585
R9015 gnd.n6293 gnd.n6292 585
R9016 gnd.n6292 gnd.n6291 585
R9017 gnd.n863 gnd.n862 585
R9018 gnd.n6290 gnd.n863 585
R9019 gnd.n6288 gnd.n6287 585
R9020 gnd.n6289 gnd.n6288 585
R9021 gnd.n6286 gnd.n865 585
R9022 gnd.n865 gnd.n864 585
R9023 gnd.n6285 gnd.n6284 585
R9024 gnd.n6284 gnd.n6283 585
R9025 gnd.n871 gnd.n870 585
R9026 gnd.n6282 gnd.n871 585
R9027 gnd.n6280 gnd.n6279 585
R9028 gnd.n6281 gnd.n6280 585
R9029 gnd.n6278 gnd.n873 585
R9030 gnd.n873 gnd.n872 585
R9031 gnd.n6277 gnd.n6276 585
R9032 gnd.n6276 gnd.n6275 585
R9033 gnd.n879 gnd.n878 585
R9034 gnd.n6274 gnd.n879 585
R9035 gnd.n6272 gnd.n6271 585
R9036 gnd.n6273 gnd.n6272 585
R9037 gnd.n6270 gnd.n881 585
R9038 gnd.n881 gnd.n880 585
R9039 gnd.n6269 gnd.n6268 585
R9040 gnd.n6268 gnd.n6267 585
R9041 gnd.n887 gnd.n886 585
R9042 gnd.n6266 gnd.n887 585
R9043 gnd.n6264 gnd.n6263 585
R9044 gnd.n6265 gnd.n6264 585
R9045 gnd.n6262 gnd.n889 585
R9046 gnd.n889 gnd.n888 585
R9047 gnd.n6261 gnd.n6260 585
R9048 gnd.n6260 gnd.n6259 585
R9049 gnd.n6429 gnd.n6428 585
R9050 gnd.n6428 gnd.n6427 585
R9051 gnd.n725 gnd.n724 585
R9052 gnd.n724 gnd.n723 585
R9053 gnd.n6434 gnd.n6433 585
R9054 gnd.n6435 gnd.n6434 585
R9055 gnd.n722 gnd.n721 585
R9056 gnd.n6436 gnd.n722 585
R9057 gnd.n6439 gnd.n6438 585
R9058 gnd.n6438 gnd.n6437 585
R9059 gnd.n719 gnd.n718 585
R9060 gnd.n718 gnd.n717 585
R9061 gnd.n6444 gnd.n6443 585
R9062 gnd.n6445 gnd.n6444 585
R9063 gnd.n716 gnd.n715 585
R9064 gnd.n6446 gnd.n716 585
R9065 gnd.n6449 gnd.n6448 585
R9066 gnd.n6448 gnd.n6447 585
R9067 gnd.n713 gnd.n712 585
R9068 gnd.n712 gnd.n711 585
R9069 gnd.n6454 gnd.n6453 585
R9070 gnd.n6455 gnd.n6454 585
R9071 gnd.n710 gnd.n709 585
R9072 gnd.n6456 gnd.n710 585
R9073 gnd.n6459 gnd.n6458 585
R9074 gnd.n6458 gnd.n6457 585
R9075 gnd.n707 gnd.n706 585
R9076 gnd.n706 gnd.n705 585
R9077 gnd.n6464 gnd.n6463 585
R9078 gnd.n6465 gnd.n6464 585
R9079 gnd.n704 gnd.n703 585
R9080 gnd.n6466 gnd.n704 585
R9081 gnd.n6469 gnd.n6468 585
R9082 gnd.n6468 gnd.n6467 585
R9083 gnd.n701 gnd.n700 585
R9084 gnd.n700 gnd.n699 585
R9085 gnd.n6474 gnd.n6473 585
R9086 gnd.n6475 gnd.n6474 585
R9087 gnd.n698 gnd.n697 585
R9088 gnd.n6476 gnd.n698 585
R9089 gnd.n6479 gnd.n6478 585
R9090 gnd.n6478 gnd.n6477 585
R9091 gnd.n695 gnd.n694 585
R9092 gnd.n694 gnd.n693 585
R9093 gnd.n6484 gnd.n6483 585
R9094 gnd.n6485 gnd.n6484 585
R9095 gnd.n692 gnd.n691 585
R9096 gnd.n6486 gnd.n692 585
R9097 gnd.n6489 gnd.n6488 585
R9098 gnd.n6488 gnd.n6487 585
R9099 gnd.n689 gnd.n688 585
R9100 gnd.n688 gnd.n687 585
R9101 gnd.n6494 gnd.n6493 585
R9102 gnd.n6495 gnd.n6494 585
R9103 gnd.n686 gnd.n685 585
R9104 gnd.n6496 gnd.n686 585
R9105 gnd.n6499 gnd.n6498 585
R9106 gnd.n6498 gnd.n6497 585
R9107 gnd.n683 gnd.n682 585
R9108 gnd.n682 gnd.n681 585
R9109 gnd.n6504 gnd.n6503 585
R9110 gnd.n6505 gnd.n6504 585
R9111 gnd.n680 gnd.n679 585
R9112 gnd.n6506 gnd.n680 585
R9113 gnd.n6509 gnd.n6508 585
R9114 gnd.n6508 gnd.n6507 585
R9115 gnd.n677 gnd.n676 585
R9116 gnd.n676 gnd.n675 585
R9117 gnd.n6514 gnd.n6513 585
R9118 gnd.n6515 gnd.n6514 585
R9119 gnd.n674 gnd.n673 585
R9120 gnd.n6516 gnd.n674 585
R9121 gnd.n6519 gnd.n6518 585
R9122 gnd.n6518 gnd.n6517 585
R9123 gnd.n671 gnd.n670 585
R9124 gnd.n670 gnd.n669 585
R9125 gnd.n6524 gnd.n6523 585
R9126 gnd.n6525 gnd.n6524 585
R9127 gnd.n668 gnd.n667 585
R9128 gnd.n6526 gnd.n668 585
R9129 gnd.n6529 gnd.n6528 585
R9130 gnd.n6528 gnd.n6527 585
R9131 gnd.n665 gnd.n664 585
R9132 gnd.n664 gnd.n663 585
R9133 gnd.n6534 gnd.n6533 585
R9134 gnd.n6535 gnd.n6534 585
R9135 gnd.n662 gnd.n661 585
R9136 gnd.n6536 gnd.n662 585
R9137 gnd.n6539 gnd.n6538 585
R9138 gnd.n6538 gnd.n6537 585
R9139 gnd.n659 gnd.n658 585
R9140 gnd.n658 gnd.n657 585
R9141 gnd.n6544 gnd.n6543 585
R9142 gnd.n6545 gnd.n6544 585
R9143 gnd.n656 gnd.n655 585
R9144 gnd.n6546 gnd.n656 585
R9145 gnd.n6549 gnd.n6548 585
R9146 gnd.n6548 gnd.n6547 585
R9147 gnd.n653 gnd.n652 585
R9148 gnd.n652 gnd.n651 585
R9149 gnd.n6554 gnd.n6553 585
R9150 gnd.n6555 gnd.n6554 585
R9151 gnd.n650 gnd.n649 585
R9152 gnd.n6556 gnd.n650 585
R9153 gnd.n6559 gnd.n6558 585
R9154 gnd.n6558 gnd.n6557 585
R9155 gnd.n647 gnd.n646 585
R9156 gnd.n646 gnd.n645 585
R9157 gnd.n6564 gnd.n6563 585
R9158 gnd.n6565 gnd.n6564 585
R9159 gnd.n644 gnd.n643 585
R9160 gnd.n6566 gnd.n644 585
R9161 gnd.n6569 gnd.n6568 585
R9162 gnd.n6568 gnd.n6567 585
R9163 gnd.n641 gnd.n640 585
R9164 gnd.n640 gnd.n639 585
R9165 gnd.n6574 gnd.n6573 585
R9166 gnd.n6575 gnd.n6574 585
R9167 gnd.n638 gnd.n637 585
R9168 gnd.n6576 gnd.n638 585
R9169 gnd.n6579 gnd.n6578 585
R9170 gnd.n6578 gnd.n6577 585
R9171 gnd.n635 gnd.n634 585
R9172 gnd.n634 gnd.n633 585
R9173 gnd.n6584 gnd.n6583 585
R9174 gnd.n6585 gnd.n6584 585
R9175 gnd.n632 gnd.n631 585
R9176 gnd.n6586 gnd.n632 585
R9177 gnd.n6589 gnd.n6588 585
R9178 gnd.n6588 gnd.n6587 585
R9179 gnd.n629 gnd.n628 585
R9180 gnd.n628 gnd.n627 585
R9181 gnd.n6594 gnd.n6593 585
R9182 gnd.n6595 gnd.n6594 585
R9183 gnd.n626 gnd.n625 585
R9184 gnd.n6596 gnd.n626 585
R9185 gnd.n6599 gnd.n6598 585
R9186 gnd.n6598 gnd.n6597 585
R9187 gnd.n623 gnd.n622 585
R9188 gnd.n622 gnd.n621 585
R9189 gnd.n6604 gnd.n6603 585
R9190 gnd.n6605 gnd.n6604 585
R9191 gnd.n620 gnd.n619 585
R9192 gnd.n6606 gnd.n620 585
R9193 gnd.n6609 gnd.n6608 585
R9194 gnd.n6608 gnd.n6607 585
R9195 gnd.n617 gnd.n616 585
R9196 gnd.n616 gnd.n615 585
R9197 gnd.n6614 gnd.n6613 585
R9198 gnd.n6615 gnd.n6614 585
R9199 gnd.n614 gnd.n613 585
R9200 gnd.n6616 gnd.n614 585
R9201 gnd.n6619 gnd.n6618 585
R9202 gnd.n6618 gnd.n6617 585
R9203 gnd.n611 gnd.n610 585
R9204 gnd.n610 gnd.n609 585
R9205 gnd.n6624 gnd.n6623 585
R9206 gnd.n6625 gnd.n6624 585
R9207 gnd.n608 gnd.n607 585
R9208 gnd.n6626 gnd.n608 585
R9209 gnd.n6629 gnd.n6628 585
R9210 gnd.n6628 gnd.n6627 585
R9211 gnd.n605 gnd.n604 585
R9212 gnd.n604 gnd.n603 585
R9213 gnd.n6634 gnd.n6633 585
R9214 gnd.n6635 gnd.n6634 585
R9215 gnd.n602 gnd.n601 585
R9216 gnd.n6636 gnd.n602 585
R9217 gnd.n6639 gnd.n6638 585
R9218 gnd.n6638 gnd.n6637 585
R9219 gnd.n599 gnd.n598 585
R9220 gnd.n598 gnd.n597 585
R9221 gnd.n6644 gnd.n6643 585
R9222 gnd.n6645 gnd.n6644 585
R9223 gnd.n596 gnd.n595 585
R9224 gnd.n6646 gnd.n596 585
R9225 gnd.n6649 gnd.n6648 585
R9226 gnd.n6648 gnd.n6647 585
R9227 gnd.n593 gnd.n592 585
R9228 gnd.n592 gnd.n591 585
R9229 gnd.n6654 gnd.n6653 585
R9230 gnd.n6655 gnd.n6654 585
R9231 gnd.n590 gnd.n589 585
R9232 gnd.n6656 gnd.n590 585
R9233 gnd.n6659 gnd.n6658 585
R9234 gnd.n6658 gnd.n6657 585
R9235 gnd.n587 gnd.n586 585
R9236 gnd.n586 gnd.n585 585
R9237 gnd.n6664 gnd.n6663 585
R9238 gnd.n6665 gnd.n6664 585
R9239 gnd.n584 gnd.n583 585
R9240 gnd.n6666 gnd.n584 585
R9241 gnd.n6669 gnd.n6668 585
R9242 gnd.n6668 gnd.n6667 585
R9243 gnd.n581 gnd.n580 585
R9244 gnd.n580 gnd.n579 585
R9245 gnd.n6674 gnd.n6673 585
R9246 gnd.n6675 gnd.n6674 585
R9247 gnd.n578 gnd.n577 585
R9248 gnd.n6676 gnd.n578 585
R9249 gnd.n6679 gnd.n6678 585
R9250 gnd.n6678 gnd.n6677 585
R9251 gnd.n575 gnd.n574 585
R9252 gnd.n574 gnd.n573 585
R9253 gnd.n6684 gnd.n6683 585
R9254 gnd.n6685 gnd.n6684 585
R9255 gnd.n572 gnd.n571 585
R9256 gnd.n6686 gnd.n572 585
R9257 gnd.n6689 gnd.n6688 585
R9258 gnd.n6688 gnd.n6687 585
R9259 gnd.n569 gnd.n568 585
R9260 gnd.n568 gnd.n567 585
R9261 gnd.n6694 gnd.n6693 585
R9262 gnd.n6695 gnd.n6694 585
R9263 gnd.n566 gnd.n565 585
R9264 gnd.n6696 gnd.n566 585
R9265 gnd.n6699 gnd.n6698 585
R9266 gnd.n6698 gnd.n6697 585
R9267 gnd.n563 gnd.n562 585
R9268 gnd.n562 gnd.n561 585
R9269 gnd.n6704 gnd.n6703 585
R9270 gnd.n6705 gnd.n6704 585
R9271 gnd.n560 gnd.n559 585
R9272 gnd.n6706 gnd.n560 585
R9273 gnd.n6709 gnd.n6708 585
R9274 gnd.n6708 gnd.n6707 585
R9275 gnd.n557 gnd.n556 585
R9276 gnd.n556 gnd.n555 585
R9277 gnd.n6714 gnd.n6713 585
R9278 gnd.n6715 gnd.n6714 585
R9279 gnd.n554 gnd.n553 585
R9280 gnd.n6716 gnd.n554 585
R9281 gnd.n6719 gnd.n6718 585
R9282 gnd.n6718 gnd.n6717 585
R9283 gnd.n551 gnd.n550 585
R9284 gnd.n550 gnd.n549 585
R9285 gnd.n6724 gnd.n6723 585
R9286 gnd.n6725 gnd.n6724 585
R9287 gnd.n548 gnd.n547 585
R9288 gnd.n6726 gnd.n548 585
R9289 gnd.n6729 gnd.n6728 585
R9290 gnd.n6728 gnd.n6727 585
R9291 gnd.n545 gnd.n544 585
R9292 gnd.n544 gnd.n543 585
R9293 gnd.n6734 gnd.n6733 585
R9294 gnd.n6735 gnd.n6734 585
R9295 gnd.n542 gnd.n541 585
R9296 gnd.n6736 gnd.n542 585
R9297 gnd.n6739 gnd.n6738 585
R9298 gnd.n6738 gnd.n6737 585
R9299 gnd.n539 gnd.n538 585
R9300 gnd.n538 gnd.n537 585
R9301 gnd.n6744 gnd.n6743 585
R9302 gnd.n6745 gnd.n6744 585
R9303 gnd.n536 gnd.n535 585
R9304 gnd.n6746 gnd.n536 585
R9305 gnd.n6749 gnd.n6748 585
R9306 gnd.n6748 gnd.n6747 585
R9307 gnd.n533 gnd.n532 585
R9308 gnd.n532 gnd.n531 585
R9309 gnd.n6754 gnd.n6753 585
R9310 gnd.n6755 gnd.n6754 585
R9311 gnd.n530 gnd.n529 585
R9312 gnd.n6756 gnd.n530 585
R9313 gnd.n6759 gnd.n6758 585
R9314 gnd.n6758 gnd.n6757 585
R9315 gnd.n527 gnd.n526 585
R9316 gnd.n526 gnd.n525 585
R9317 gnd.n6764 gnd.n6763 585
R9318 gnd.n6765 gnd.n6764 585
R9319 gnd.n524 gnd.n523 585
R9320 gnd.n6766 gnd.n524 585
R9321 gnd.n6769 gnd.n6768 585
R9322 gnd.n6768 gnd.n6767 585
R9323 gnd.n521 gnd.n520 585
R9324 gnd.n520 gnd.n519 585
R9325 gnd.n6774 gnd.n6773 585
R9326 gnd.n6775 gnd.n6774 585
R9327 gnd.n518 gnd.n517 585
R9328 gnd.n6776 gnd.n518 585
R9329 gnd.n6779 gnd.n6778 585
R9330 gnd.n6778 gnd.n6777 585
R9331 gnd.n515 gnd.n514 585
R9332 gnd.n514 gnd.n513 585
R9333 gnd.n6784 gnd.n6783 585
R9334 gnd.n6785 gnd.n6784 585
R9335 gnd.n512 gnd.n511 585
R9336 gnd.n6786 gnd.n512 585
R9337 gnd.n6789 gnd.n6788 585
R9338 gnd.n6788 gnd.n6787 585
R9339 gnd.n509 gnd.n508 585
R9340 gnd.n508 gnd.n507 585
R9341 gnd.n6794 gnd.n6793 585
R9342 gnd.n6795 gnd.n6794 585
R9343 gnd.n506 gnd.n505 585
R9344 gnd.n6796 gnd.n506 585
R9345 gnd.n6799 gnd.n6798 585
R9346 gnd.n6798 gnd.n6797 585
R9347 gnd.n503 gnd.n502 585
R9348 gnd.n502 gnd.n501 585
R9349 gnd.n6804 gnd.n6803 585
R9350 gnd.n6805 gnd.n6804 585
R9351 gnd.n500 gnd.n499 585
R9352 gnd.n6806 gnd.n500 585
R9353 gnd.n6809 gnd.n6808 585
R9354 gnd.n6808 gnd.n6807 585
R9355 gnd.n497 gnd.n496 585
R9356 gnd.n496 gnd.n495 585
R9357 gnd.n6814 gnd.n6813 585
R9358 gnd.n6815 gnd.n6814 585
R9359 gnd.n494 gnd.n493 585
R9360 gnd.n6816 gnd.n494 585
R9361 gnd.n6819 gnd.n6818 585
R9362 gnd.n6818 gnd.n6817 585
R9363 gnd.n491 gnd.n490 585
R9364 gnd.n490 gnd.n489 585
R9365 gnd.n6824 gnd.n6823 585
R9366 gnd.n6825 gnd.n6824 585
R9367 gnd.n488 gnd.n487 585
R9368 gnd.n6826 gnd.n488 585
R9369 gnd.n6829 gnd.n6828 585
R9370 gnd.n6828 gnd.n6827 585
R9371 gnd.n485 gnd.n484 585
R9372 gnd.n484 gnd.n483 585
R9373 gnd.n6834 gnd.n6833 585
R9374 gnd.n6835 gnd.n6834 585
R9375 gnd.n482 gnd.n481 585
R9376 gnd.n6836 gnd.n482 585
R9377 gnd.n6839 gnd.n6838 585
R9378 gnd.n6838 gnd.n6837 585
R9379 gnd.n479 gnd.n478 585
R9380 gnd.n478 gnd.n477 585
R9381 gnd.n6844 gnd.n6843 585
R9382 gnd.n6845 gnd.n6844 585
R9383 gnd.n476 gnd.n475 585
R9384 gnd.n6846 gnd.n476 585
R9385 gnd.n6849 gnd.n6848 585
R9386 gnd.n6848 gnd.n6847 585
R9387 gnd.n473 gnd.n472 585
R9388 gnd.n472 gnd.n471 585
R9389 gnd.n6854 gnd.n6853 585
R9390 gnd.n6855 gnd.n6854 585
R9391 gnd.n470 gnd.n469 585
R9392 gnd.n6856 gnd.n470 585
R9393 gnd.n6859 gnd.n6858 585
R9394 gnd.n6858 gnd.n6857 585
R9395 gnd.n467 gnd.n466 585
R9396 gnd.n466 gnd.n465 585
R9397 gnd.n6864 gnd.n6863 585
R9398 gnd.n6865 gnd.n6864 585
R9399 gnd.n464 gnd.n463 585
R9400 gnd.n6866 gnd.n464 585
R9401 gnd.n6869 gnd.n6868 585
R9402 gnd.n6868 gnd.n6867 585
R9403 gnd.n461 gnd.n460 585
R9404 gnd.n460 gnd.n459 585
R9405 gnd.n6875 gnd.n6874 585
R9406 gnd.n6876 gnd.n6875 585
R9407 gnd.n458 gnd.n457 585
R9408 gnd.n6877 gnd.n458 585
R9409 gnd.n6880 gnd.n6879 585
R9410 gnd.n6879 gnd.n6878 585
R9411 gnd.n6881 gnd.n455 585
R9412 gnd.n455 gnd.n454 585
R9413 gnd.n330 gnd.n329 585
R9414 gnd.n7088 gnd.n329 585
R9415 gnd.n7091 gnd.n7090 585
R9416 gnd.n7090 gnd.n7089 585
R9417 gnd.n333 gnd.n332 585
R9418 gnd.n7087 gnd.n333 585
R9419 gnd.n7085 gnd.n7084 585
R9420 gnd.n7086 gnd.n7085 585
R9421 gnd.n336 gnd.n335 585
R9422 gnd.n335 gnd.n334 585
R9423 gnd.n7080 gnd.n7079 585
R9424 gnd.n7079 gnd.n7078 585
R9425 gnd.n339 gnd.n338 585
R9426 gnd.n7077 gnd.n339 585
R9427 gnd.n7075 gnd.n7074 585
R9428 gnd.n7076 gnd.n7075 585
R9429 gnd.n342 gnd.n341 585
R9430 gnd.n341 gnd.n340 585
R9431 gnd.n7070 gnd.n7069 585
R9432 gnd.n7069 gnd.n7068 585
R9433 gnd.n345 gnd.n344 585
R9434 gnd.n7067 gnd.n345 585
R9435 gnd.n7065 gnd.n7064 585
R9436 gnd.n7066 gnd.n7065 585
R9437 gnd.n348 gnd.n347 585
R9438 gnd.n347 gnd.n346 585
R9439 gnd.n7060 gnd.n7059 585
R9440 gnd.n7059 gnd.n7058 585
R9441 gnd.n351 gnd.n350 585
R9442 gnd.n7057 gnd.n351 585
R9443 gnd.n7055 gnd.n7054 585
R9444 gnd.n7056 gnd.n7055 585
R9445 gnd.n354 gnd.n353 585
R9446 gnd.n353 gnd.n352 585
R9447 gnd.n7050 gnd.n7049 585
R9448 gnd.n7049 gnd.n7048 585
R9449 gnd.n357 gnd.n356 585
R9450 gnd.n7047 gnd.n357 585
R9451 gnd.n7045 gnd.n7044 585
R9452 gnd.n7046 gnd.n7045 585
R9453 gnd.n360 gnd.n359 585
R9454 gnd.n359 gnd.n358 585
R9455 gnd.n7040 gnd.n7039 585
R9456 gnd.n7039 gnd.n7038 585
R9457 gnd.n363 gnd.n362 585
R9458 gnd.n7037 gnd.n363 585
R9459 gnd.n7035 gnd.n7034 585
R9460 gnd.n7036 gnd.n7035 585
R9461 gnd.n366 gnd.n365 585
R9462 gnd.n365 gnd.n364 585
R9463 gnd.n7030 gnd.n7029 585
R9464 gnd.n7029 gnd.n7028 585
R9465 gnd.n369 gnd.n368 585
R9466 gnd.n7027 gnd.n369 585
R9467 gnd.n7025 gnd.n7024 585
R9468 gnd.n7026 gnd.n7025 585
R9469 gnd.n372 gnd.n371 585
R9470 gnd.n371 gnd.n370 585
R9471 gnd.n7020 gnd.n7019 585
R9472 gnd.n7019 gnd.n7018 585
R9473 gnd.n375 gnd.n374 585
R9474 gnd.n7017 gnd.n375 585
R9475 gnd.n7015 gnd.n7014 585
R9476 gnd.n7016 gnd.n7015 585
R9477 gnd.n378 gnd.n377 585
R9478 gnd.n377 gnd.n376 585
R9479 gnd.n7010 gnd.n7009 585
R9480 gnd.n7009 gnd.n7008 585
R9481 gnd.n381 gnd.n380 585
R9482 gnd.n7007 gnd.n381 585
R9483 gnd.n7005 gnd.n7004 585
R9484 gnd.n7006 gnd.n7005 585
R9485 gnd.n384 gnd.n383 585
R9486 gnd.n383 gnd.n382 585
R9487 gnd.n7000 gnd.n6999 585
R9488 gnd.n6999 gnd.n6998 585
R9489 gnd.n387 gnd.n386 585
R9490 gnd.n6997 gnd.n387 585
R9491 gnd.n6995 gnd.n6994 585
R9492 gnd.n6996 gnd.n6995 585
R9493 gnd.n390 gnd.n389 585
R9494 gnd.n389 gnd.n388 585
R9495 gnd.n6990 gnd.n6989 585
R9496 gnd.n6989 gnd.n6988 585
R9497 gnd.n393 gnd.n392 585
R9498 gnd.n6987 gnd.n393 585
R9499 gnd.n6985 gnd.n6984 585
R9500 gnd.n6986 gnd.n6985 585
R9501 gnd.n396 gnd.n395 585
R9502 gnd.n395 gnd.n394 585
R9503 gnd.n6980 gnd.n6979 585
R9504 gnd.n6979 gnd.n6978 585
R9505 gnd.n399 gnd.n398 585
R9506 gnd.n6977 gnd.n399 585
R9507 gnd.n6975 gnd.n6974 585
R9508 gnd.n6976 gnd.n6975 585
R9509 gnd.n402 gnd.n401 585
R9510 gnd.n401 gnd.n400 585
R9511 gnd.n6970 gnd.n6969 585
R9512 gnd.n6969 gnd.n6968 585
R9513 gnd.n405 gnd.n404 585
R9514 gnd.n6967 gnd.n405 585
R9515 gnd.n6965 gnd.n6964 585
R9516 gnd.n6966 gnd.n6965 585
R9517 gnd.n408 gnd.n407 585
R9518 gnd.n407 gnd.n406 585
R9519 gnd.n6960 gnd.n6959 585
R9520 gnd.n6959 gnd.n6958 585
R9521 gnd.n411 gnd.n410 585
R9522 gnd.n6957 gnd.n411 585
R9523 gnd.n6955 gnd.n6954 585
R9524 gnd.n6956 gnd.n6955 585
R9525 gnd.n414 gnd.n413 585
R9526 gnd.n413 gnd.n412 585
R9527 gnd.n6950 gnd.n6949 585
R9528 gnd.n6949 gnd.n6948 585
R9529 gnd.n417 gnd.n416 585
R9530 gnd.n6947 gnd.n417 585
R9531 gnd.n6945 gnd.n6944 585
R9532 gnd.n6946 gnd.n6945 585
R9533 gnd.n420 gnd.n419 585
R9534 gnd.n419 gnd.n418 585
R9535 gnd.n6940 gnd.n6939 585
R9536 gnd.n6939 gnd.n6938 585
R9537 gnd.n423 gnd.n422 585
R9538 gnd.n6937 gnd.n423 585
R9539 gnd.n6935 gnd.n6934 585
R9540 gnd.n6936 gnd.n6935 585
R9541 gnd.n426 gnd.n425 585
R9542 gnd.n425 gnd.n424 585
R9543 gnd.n6930 gnd.n6929 585
R9544 gnd.n6929 gnd.n6928 585
R9545 gnd.n429 gnd.n428 585
R9546 gnd.n6927 gnd.n429 585
R9547 gnd.n6925 gnd.n6924 585
R9548 gnd.n6926 gnd.n6925 585
R9549 gnd.n432 gnd.n431 585
R9550 gnd.n431 gnd.n430 585
R9551 gnd.n6920 gnd.n6919 585
R9552 gnd.n6919 gnd.n6918 585
R9553 gnd.n435 gnd.n434 585
R9554 gnd.n6917 gnd.n435 585
R9555 gnd.n6915 gnd.n6914 585
R9556 gnd.n6916 gnd.n6915 585
R9557 gnd.n438 gnd.n437 585
R9558 gnd.n437 gnd.n436 585
R9559 gnd.n6910 gnd.n6909 585
R9560 gnd.n6909 gnd.n6908 585
R9561 gnd.n441 gnd.n440 585
R9562 gnd.n6907 gnd.n441 585
R9563 gnd.n6905 gnd.n6904 585
R9564 gnd.n6906 gnd.n6905 585
R9565 gnd.n444 gnd.n443 585
R9566 gnd.n443 gnd.n442 585
R9567 gnd.n6900 gnd.n6899 585
R9568 gnd.n6899 gnd.n6898 585
R9569 gnd.n447 gnd.n446 585
R9570 gnd.n6897 gnd.n447 585
R9571 gnd.n6895 gnd.n6894 585
R9572 gnd.n6896 gnd.n6895 585
R9573 gnd.n450 gnd.n449 585
R9574 gnd.n449 gnd.n448 585
R9575 gnd.n6890 gnd.n6889 585
R9576 gnd.n6889 gnd.n6888 585
R9577 gnd.n453 gnd.n452 585
R9578 gnd.n6887 gnd.n453 585
R9579 gnd.n6885 gnd.n6884 585
R9580 gnd.n6886 gnd.n6885 585
R9581 gnd.n4593 gnd.n4592 585
R9582 gnd.n4594 gnd.n4593 585
R9583 gnd.n1260 gnd.n1259 585
R9584 gnd.n2821 gnd.n1260 585
R9585 gnd.n4602 gnd.n4601 585
R9586 gnd.n4601 gnd.n4600 585
R9587 gnd.n4603 gnd.n1254 585
R9588 gnd.n2781 gnd.n1254 585
R9589 gnd.n4605 gnd.n4604 585
R9590 gnd.n4606 gnd.n4605 585
R9591 gnd.n1239 gnd.n1238 585
R9592 gnd.n2772 gnd.n1239 585
R9593 gnd.n4614 gnd.n4613 585
R9594 gnd.n4613 gnd.n4612 585
R9595 gnd.n4615 gnd.n1233 585
R9596 gnd.n2764 gnd.n1233 585
R9597 gnd.n4617 gnd.n4616 585
R9598 gnd.n4618 gnd.n4617 585
R9599 gnd.n1217 gnd.n1216 585
R9600 gnd.n2694 gnd.n1217 585
R9601 gnd.n4626 gnd.n4625 585
R9602 gnd.n4625 gnd.n4624 585
R9603 gnd.n4627 gnd.n1211 585
R9604 gnd.n2682 gnd.n1211 585
R9605 gnd.n4629 gnd.n4628 585
R9606 gnd.n4630 gnd.n4629 585
R9607 gnd.n1197 gnd.n1196 585
R9608 gnd.n2677 gnd.n1197 585
R9609 gnd.n4638 gnd.n4637 585
R9610 gnd.n4637 gnd.n4636 585
R9611 gnd.n4639 gnd.n1191 585
R9612 gnd.n2708 gnd.n1191 585
R9613 gnd.n4641 gnd.n4640 585
R9614 gnd.n4642 gnd.n4641 585
R9615 gnd.n1175 gnd.n1174 585
R9616 gnd.n2669 gnd.n1175 585
R9617 gnd.n4650 gnd.n4649 585
R9618 gnd.n4649 gnd.n4648 585
R9619 gnd.n4651 gnd.n1169 585
R9620 gnd.n2661 gnd.n1169 585
R9621 gnd.n4653 gnd.n4652 585
R9622 gnd.n4654 gnd.n4653 585
R9623 gnd.n1156 gnd.n1155 585
R9624 gnd.n2652 gnd.n1156 585
R9625 gnd.n4662 gnd.n4661 585
R9626 gnd.n4661 gnd.n4660 585
R9627 gnd.n4663 gnd.n1150 585
R9628 gnd.n2644 gnd.n1150 585
R9629 gnd.n4665 gnd.n4664 585
R9630 gnd.n4666 gnd.n4665 585
R9631 gnd.n1137 gnd.n1136 585
R9632 gnd.n2612 gnd.n1137 585
R9633 gnd.n4675 gnd.n4674 585
R9634 gnd.n4674 gnd.n4673 585
R9635 gnd.n4676 gnd.n1131 585
R9636 gnd.n2621 gnd.n1131 585
R9637 gnd.n4678 gnd.n4677 585
R9638 gnd.n4679 gnd.n4678 585
R9639 gnd.n1119 gnd.n1118 585
R9640 gnd.n2627 gnd.n1119 585
R9641 gnd.n4687 gnd.n4686 585
R9642 gnd.n4686 gnd.n4685 585
R9643 gnd.n4688 gnd.n1113 585
R9644 gnd.n2633 gnd.n1113 585
R9645 gnd.n4690 gnd.n4689 585
R9646 gnd.n4691 gnd.n4690 585
R9647 gnd.n1096 gnd.n1095 585
R9648 gnd.n2577 gnd.n1096 585
R9649 gnd.n4699 gnd.n4698 585
R9650 gnd.n4698 gnd.n4697 585
R9651 gnd.n4700 gnd.n1090 585
R9652 gnd.n1098 gnd.n1090 585
R9653 gnd.n4702 gnd.n4701 585
R9654 gnd.n4703 gnd.n4702 585
R9655 gnd.n1077 gnd.n1076 585
R9656 gnd.n1080 gnd.n1077 585
R9657 gnd.n4711 gnd.n4710 585
R9658 gnd.n4710 gnd.n4709 585
R9659 gnd.n4712 gnd.n1071 585
R9660 gnd.n1071 gnd.n1070 585
R9661 gnd.n4714 gnd.n4713 585
R9662 gnd.n4715 gnd.n4714 585
R9663 gnd.n1056 gnd.n1055 585
R9664 gnd.n1067 gnd.n1056 585
R9665 gnd.n4723 gnd.n4722 585
R9666 gnd.n4722 gnd.n4721 585
R9667 gnd.n4724 gnd.n1050 585
R9668 gnd.n1057 gnd.n1050 585
R9669 gnd.n4726 gnd.n4725 585
R9670 gnd.n4727 gnd.n4726 585
R9671 gnd.n1037 gnd.n1036 585
R9672 gnd.n1040 gnd.n1037 585
R9673 gnd.n4735 gnd.n4734 585
R9674 gnd.n4734 gnd.n4733 585
R9675 gnd.n4736 gnd.n1031 585
R9676 gnd.n1031 gnd.n1029 585
R9677 gnd.n4738 gnd.n4737 585
R9678 gnd.n4739 gnd.n4738 585
R9679 gnd.n1032 gnd.n1030 585
R9680 gnd.n1030 gnd.n1017 585
R9681 gnd.n2523 gnd.n1018 585
R9682 gnd.n4745 gnd.n1018 585
R9683 gnd.n2460 gnd.n2458 585
R9684 gnd.n2458 gnd.n1015 585
R9685 gnd.n2528 gnd.n2527 585
R9686 gnd.n2535 gnd.n2528 585
R9687 gnd.n2459 gnd.n2457 585
R9688 gnd.n2457 gnd.n961 585
R9689 gnd.n2519 gnd.n2518 585
R9690 gnd.n2517 gnd.n2516 585
R9691 gnd.n2515 gnd.n2514 585
R9692 gnd.n2513 gnd.n2512 585
R9693 gnd.n2511 gnd.n2510 585
R9694 gnd.n2509 gnd.n2508 585
R9695 gnd.n2507 gnd.n2506 585
R9696 gnd.n2505 gnd.n2504 585
R9697 gnd.n2503 gnd.n2502 585
R9698 gnd.n2501 gnd.n2500 585
R9699 gnd.n2499 gnd.n2498 585
R9700 gnd.n2497 gnd.n2496 585
R9701 gnd.n2495 gnd.n2494 585
R9702 gnd.n2493 gnd.n2492 585
R9703 gnd.n2491 gnd.n2490 585
R9704 gnd.n2489 gnd.n2488 585
R9705 gnd.n2487 gnd.n2486 585
R9706 gnd.n2479 gnd.n2476 585
R9707 gnd.n2482 gnd.n960 585
R9708 gnd.n4832 gnd.n960 585
R9709 gnd.n3673 gnd.n3672 585
R9710 gnd.n2233 gnd.n2225 585
R9711 gnd.n3680 gnd.n2222 585
R9712 gnd.n3681 gnd.n2221 585
R9713 gnd.n2247 gnd.n2215 585
R9714 gnd.n3688 gnd.n2214 585
R9715 gnd.n3689 gnd.n2213 585
R9716 gnd.n2245 gnd.n2205 585
R9717 gnd.n3696 gnd.n2204 585
R9718 gnd.n3697 gnd.n2203 585
R9719 gnd.n2242 gnd.n2197 585
R9720 gnd.n3704 gnd.n2196 585
R9721 gnd.n3705 gnd.n2195 585
R9722 gnd.n2240 gnd.n2188 585
R9723 gnd.n3712 gnd.n2187 585
R9724 gnd.n3713 gnd.n2186 585
R9725 gnd.n2237 gnd.n2185 585
R9726 gnd.n2236 gnd.n2235 585
R9727 gnd.n1276 gnd.n1274 585
R9728 gnd.n3670 gnd.n1274 585
R9729 gnd.n2318 gnd.n1272 585
R9730 gnd.n4594 gnd.n1272 585
R9731 gnd.n2820 gnd.n2819 585
R9732 gnd.n2821 gnd.n2820 585
R9733 gnd.n2317 gnd.n1263 585
R9734 gnd.n4600 gnd.n1263 585
R9735 gnd.n2783 gnd.n2782 585
R9736 gnd.n2782 gnd.n2781 585
R9737 gnd.n2320 gnd.n1252 585
R9738 gnd.n4606 gnd.n1252 585
R9739 gnd.n2771 gnd.n2770 585
R9740 gnd.n2772 gnd.n2771 585
R9741 gnd.n2324 gnd.n1241 585
R9742 gnd.n4612 gnd.n1241 585
R9743 gnd.n2766 gnd.n2765 585
R9744 gnd.n2765 gnd.n2764 585
R9745 gnd.n2326 gnd.n1231 585
R9746 gnd.n4618 gnd.n1231 585
R9747 gnd.n2696 gnd.n2695 585
R9748 gnd.n2695 gnd.n2694 585
R9749 gnd.n2346 gnd.n1220 585
R9750 gnd.n4624 gnd.n1220 585
R9751 gnd.n2700 gnd.n2345 585
R9752 gnd.n2682 gnd.n2345 585
R9753 gnd.n2701 gnd.n1210 585
R9754 gnd.n4630 gnd.n1210 585
R9755 gnd.n2702 gnd.n2344 585
R9756 gnd.n2677 gnd.n2344 585
R9757 gnd.n2341 gnd.n1199 585
R9758 gnd.n4636 gnd.n1199 585
R9759 gnd.n2707 gnd.n2706 585
R9760 gnd.n2708 gnd.n2707 585
R9761 gnd.n2340 gnd.n1189 585
R9762 gnd.n4642 gnd.n1189 585
R9763 gnd.n2668 gnd.n2667 585
R9764 gnd.n2669 gnd.n2668 585
R9765 gnd.n2353 gnd.n1178 585
R9766 gnd.n4648 gnd.n1178 585
R9767 gnd.n2663 gnd.n2662 585
R9768 gnd.n2662 gnd.n2661 585
R9769 gnd.n2355 gnd.n1168 585
R9770 gnd.n4654 gnd.n1168 585
R9771 gnd.n2651 gnd.n2650 585
R9772 gnd.n2652 gnd.n2651 585
R9773 gnd.n2360 gnd.n1158 585
R9774 gnd.n4660 gnd.n1158 585
R9775 gnd.n2646 gnd.n2645 585
R9776 gnd.n2645 gnd.n2644 585
R9777 gnd.n2362 gnd.n1148 585
R9778 gnd.n4666 gnd.n1148 585
R9779 gnd.n2614 gnd.n2613 585
R9780 gnd.n2613 gnd.n2612 585
R9781 gnd.n2618 gnd.n1140 585
R9782 gnd.n4673 gnd.n1140 585
R9783 gnd.n2620 gnd.n2619 585
R9784 gnd.n2621 gnd.n2620 585
R9785 gnd.n2404 gnd.n1130 585
R9786 gnd.n4679 gnd.n1130 585
R9787 gnd.n2629 gnd.n2628 585
R9788 gnd.n2628 gnd.n2627 585
R9789 gnd.n2630 gnd.n1121 585
R9790 gnd.n4685 gnd.n1121 585
R9791 gnd.n2632 gnd.n2631 585
R9792 gnd.n2633 gnd.n2632 585
R9793 gnd.n2400 gnd.n1111 585
R9794 gnd.n4691 gnd.n1111 585
R9795 gnd.n2576 gnd.n2575 585
R9796 gnd.n2577 gnd.n2576 585
R9797 gnd.n2445 gnd.n1100 585
R9798 gnd.n4697 gnd.n1100 585
R9799 gnd.n2570 gnd.n2569 585
R9800 gnd.n2569 gnd.n1098 585
R9801 gnd.n2568 gnd.n1089 585
R9802 gnd.n4703 gnd.n1089 585
R9803 gnd.n2567 gnd.n2566 585
R9804 gnd.n2566 gnd.n1080 585
R9805 gnd.n2447 gnd.n1079 585
R9806 gnd.n4709 gnd.n1079 585
R9807 gnd.n2562 gnd.n2561 585
R9808 gnd.n2561 gnd.n1070 585
R9809 gnd.n2560 gnd.n1069 585
R9810 gnd.n4715 gnd.n1069 585
R9811 gnd.n2559 gnd.n2558 585
R9812 gnd.n2558 gnd.n1067 585
R9813 gnd.n2449 gnd.n1059 585
R9814 gnd.n4721 gnd.n1059 585
R9815 gnd.n2554 gnd.n2553 585
R9816 gnd.n2553 gnd.n1057 585
R9817 gnd.n2552 gnd.n1049 585
R9818 gnd.n4727 gnd.n1049 585
R9819 gnd.n2551 gnd.n2550 585
R9820 gnd.n2550 gnd.n1040 585
R9821 gnd.n2451 gnd.n1039 585
R9822 gnd.n4733 gnd.n1039 585
R9823 gnd.n2546 gnd.n2545 585
R9824 gnd.n2545 gnd.n1029 585
R9825 gnd.n2544 gnd.n1028 585
R9826 gnd.n4739 gnd.n1028 585
R9827 gnd.n2543 gnd.n2542 585
R9828 gnd.n2542 gnd.n1017 585
R9829 gnd.n2453 gnd.n1016 585
R9830 gnd.n4745 gnd.n1016 585
R9831 gnd.n2538 gnd.n2537 585
R9832 gnd.n2537 gnd.n1015 585
R9833 gnd.n2536 gnd.n2455 585
R9834 gnd.n2536 gnd.n2535 585
R9835 gnd.n2480 gnd.n2456 585
R9836 gnd.n2456 gnd.n961 585
R9837 gnd.n7365 gnd.n107 585
R9838 gnd.n7461 gnd.n107 585
R9839 gnd.n7366 gnd.n7296 585
R9840 gnd.n7296 gnd.n104 585
R9841 gnd.n7367 gnd.n187 585
R9842 gnd.n7381 gnd.n187 585
R9843 gnd.n198 gnd.n196 585
R9844 gnd.n196 gnd.n185 585
R9845 gnd.n7372 gnd.n7371 585
R9846 gnd.n7373 gnd.n7372 585
R9847 gnd.n197 gnd.n195 585
R9848 gnd.n195 gnd.n193 585
R9849 gnd.n7292 gnd.n7291 585
R9850 gnd.n7291 gnd.n7290 585
R9851 gnd.n201 gnd.n200 585
R9852 gnd.n211 gnd.n201 585
R9853 gnd.n7281 gnd.n7280 585
R9854 gnd.n7282 gnd.n7281 585
R9855 gnd.n213 gnd.n212 585
R9856 gnd.n212 gnd.n208 585
R9857 gnd.n7276 gnd.n7275 585
R9858 gnd.n7275 gnd.n7274 585
R9859 gnd.n216 gnd.n215 585
R9860 gnd.n218 gnd.n216 585
R9861 gnd.n7265 gnd.n7264 585
R9862 gnd.n7266 gnd.n7265 585
R9863 gnd.n228 gnd.n227 585
R9864 gnd.n227 gnd.n225 585
R9865 gnd.n7260 gnd.n7259 585
R9866 gnd.n7259 gnd.n7258 585
R9867 gnd.n231 gnd.n230 585
R9868 gnd.n241 gnd.n231 585
R9869 gnd.n7249 gnd.n7248 585
R9870 gnd.n7250 gnd.n7249 585
R9871 gnd.n243 gnd.n242 585
R9872 gnd.n242 gnd.n238 585
R9873 gnd.n7244 gnd.n7243 585
R9874 gnd.n7243 gnd.n7242 585
R9875 gnd.n246 gnd.n245 585
R9876 gnd.n248 gnd.n246 585
R9877 gnd.n7233 gnd.n7232 585
R9878 gnd.n7234 gnd.n7233 585
R9879 gnd.n259 gnd.n258 585
R9880 gnd.n7187 gnd.n258 585
R9881 gnd.n7228 gnd.n7227 585
R9882 gnd.n7227 gnd.n7226 585
R9883 gnd.n262 gnd.n261 585
R9884 gnd.n7192 gnd.n262 585
R9885 gnd.n7205 gnd.n7204 585
R9886 gnd.n7204 gnd.n7203 585
R9887 gnd.n7206 gnd.n293 585
R9888 gnd.n7198 gnd.n293 585
R9889 gnd.n319 gnd.n290 585
R9890 gnd.n320 gnd.n319 585
R9891 gnd.n7211 gnd.n289 585
R9892 gnd.n7132 gnd.n289 585
R9893 gnd.n7212 gnd.n288 585
R9894 gnd.n7127 gnd.n288 585
R9895 gnd.n7213 gnd.n287 585
R9896 gnd.n314 gnd.n287 585
R9897 gnd.n284 gnd.n282 585
R9898 gnd.n7119 gnd.n282 585
R9899 gnd.n7218 gnd.n7217 585
R9900 gnd.n7219 gnd.n7218 585
R9901 gnd.n283 gnd.n281 585
R9902 gnd.n4276 gnd.n281 585
R9903 gnd.n4317 gnd.n4315 585
R9904 gnd.n4315 gnd.n4314 585
R9905 gnd.n4318 gnd.n1526 585
R9906 gnd.n1538 gnd.n1526 585
R9907 gnd.n4319 gnd.n1525 585
R9908 gnd.n4306 gnd.n1525 585
R9909 gnd.n4287 gnd.n1523 585
R9910 gnd.n4288 gnd.n4287 585
R9911 gnd.n4323 gnd.n1522 585
R9912 gnd.n1546 gnd.n1522 585
R9913 gnd.n4324 gnd.n1521 585
R9914 gnd.n4253 gnd.n1521 585
R9915 gnd.n4325 gnd.n1520 585
R9916 gnd.n1573 gnd.n1520 585
R9917 gnd.n4242 gnd.n1518 585
R9918 gnd.n4243 gnd.n4242 585
R9919 gnd.n4329 gnd.n1517 585
R9920 gnd.n4230 gnd.n1517 585
R9921 gnd.n4330 gnd.n1516 585
R9922 gnd.n1580 gnd.n1516 585
R9923 gnd.n4331 gnd.n1515 585
R9924 gnd.n4216 gnd.n1515 585
R9925 gnd.n1600 gnd.n1513 585
R9926 gnd.n1601 gnd.n1600 585
R9927 gnd.n4335 gnd.n1512 585
R9928 gnd.n4206 gnd.n1512 585
R9929 gnd.n4336 gnd.n1511 585
R9930 gnd.n4194 gnd.n1511 585
R9931 gnd.n4337 gnd.n1510 585
R9932 gnd.n1671 gnd.n1510 585
R9933 gnd.n1618 gnd.n1508 585
R9934 gnd.n4185 gnd.n1618 585
R9935 gnd.n4341 gnd.n1507 585
R9936 gnd.n1628 gnd.n1507 585
R9937 gnd.n4342 gnd.n1506 585
R9938 gnd.n4175 gnd.n1506 585
R9939 gnd.n4343 gnd.n1505 585
R9940 gnd.n4163 gnd.n1505 585
R9941 gnd.n1502 gnd.n1501 585
R9942 gnd.n1647 gnd.n1501 585
R9943 gnd.n4348 gnd.n4347 585
R9944 gnd.n4349 gnd.n4348 585
R9945 gnd.n1722 gnd.n1500 585
R9946 gnd.n1727 gnd.n1726 585
R9947 gnd.n1729 gnd.n1728 585
R9948 gnd.n1732 gnd.n1731 585
R9949 gnd.n1730 gnd.n1715 585
R9950 gnd.n1746 gnd.n1745 585
R9951 gnd.n1748 gnd.n1747 585
R9952 gnd.n1751 gnd.n1750 585
R9953 gnd.n1749 gnd.n1708 585
R9954 gnd.n1765 gnd.n1764 585
R9955 gnd.n1767 gnd.n1766 585
R9956 gnd.n1770 gnd.n1769 585
R9957 gnd.n1768 gnd.n1701 585
R9958 gnd.n1783 gnd.n1782 585
R9959 gnd.n1785 gnd.n1784 585
R9960 gnd.n1694 gnd.n1693 585
R9961 gnd.n1798 gnd.n1695 585
R9962 gnd.n1799 gnd.n1690 585
R9963 gnd.n1800 gnd.n1445 585
R9964 gnd.n4425 gnd.n1445 585
R9965 gnd.n7336 gnd.n103 585
R9966 gnd.n7337 gnd.n7334 585
R9967 gnd.n7338 gnd.n7330 585
R9968 gnd.n7328 gnd.n7326 585
R9969 gnd.n7342 gnd.n7325 585
R9970 gnd.n7343 gnd.n7323 585
R9971 gnd.n7344 gnd.n7322 585
R9972 gnd.n7320 gnd.n7318 585
R9973 gnd.n7348 gnd.n7317 585
R9974 gnd.n7349 gnd.n7315 585
R9975 gnd.n7350 gnd.n7314 585
R9976 gnd.n7312 gnd.n7310 585
R9977 gnd.n7354 gnd.n7309 585
R9978 gnd.n7355 gnd.n7307 585
R9979 gnd.n7356 gnd.n7306 585
R9980 gnd.n7304 gnd.n7302 585
R9981 gnd.n7360 gnd.n7301 585
R9982 gnd.n7361 gnd.n7299 585
R9983 gnd.n7362 gnd.n7298 585
R9984 gnd.n7298 gnd.n106 585
R9985 gnd.n7463 gnd.n7462 585
R9986 gnd.n7462 gnd.n7461 585
R9987 gnd.n7464 gnd.n101 585
R9988 gnd.n104 gnd.n101 585
R9989 gnd.n7465 gnd.n100 585
R9990 gnd.n7381 gnd.n100 585
R9991 gnd.n184 gnd.n98 585
R9992 gnd.n185 gnd.n184 585
R9993 gnd.n7469 gnd.n97 585
R9994 gnd.n7373 gnd.n97 585
R9995 gnd.n7470 gnd.n96 585
R9996 gnd.n193 gnd.n96 585
R9997 gnd.n7471 gnd.n95 585
R9998 gnd.n7290 gnd.n95 585
R9999 gnd.n210 gnd.n93 585
R10000 gnd.n211 gnd.n210 585
R10001 gnd.n7475 gnd.n92 585
R10002 gnd.n7282 gnd.n92 585
R10003 gnd.n7476 gnd.n91 585
R10004 gnd.n208 gnd.n91 585
R10005 gnd.n7477 gnd.n90 585
R10006 gnd.n7274 gnd.n90 585
R10007 gnd.n217 gnd.n88 585
R10008 gnd.n218 gnd.n217 585
R10009 gnd.n7481 gnd.n87 585
R10010 gnd.n7266 gnd.n87 585
R10011 gnd.n7482 gnd.n86 585
R10012 gnd.n225 gnd.n86 585
R10013 gnd.n7483 gnd.n85 585
R10014 gnd.n7258 gnd.n85 585
R10015 gnd.n240 gnd.n83 585
R10016 gnd.n241 gnd.n240 585
R10017 gnd.n7487 gnd.n82 585
R10018 gnd.n7250 gnd.n82 585
R10019 gnd.n7488 gnd.n81 585
R10020 gnd.n238 gnd.n81 585
R10021 gnd.n7489 gnd.n80 585
R10022 gnd.n7242 gnd.n80 585
R10023 gnd.n247 gnd.n78 585
R10024 gnd.n248 gnd.n247 585
R10025 gnd.n7493 gnd.n77 585
R10026 gnd.n7234 gnd.n77 585
R10027 gnd.n7494 gnd.n76 585
R10028 gnd.n7187 gnd.n76 585
R10029 gnd.n7495 gnd.n75 585
R10030 gnd.n7226 gnd.n75 585
R10031 gnd.n7191 gnd.n73 585
R10032 gnd.n7192 gnd.n7191 585
R10033 gnd.n7499 gnd.n72 585
R10034 gnd.n7203 gnd.n72 585
R10035 gnd.n7500 gnd.n71 585
R10036 gnd.n7198 gnd.n71 585
R10037 gnd.n7501 gnd.n70 585
R10038 gnd.n320 gnd.n70 585
R10039 gnd.n303 gnd.n69 585
R10040 gnd.n7132 gnd.n303 585
R10041 gnd.n7126 gnd.n7125 585
R10042 gnd.n7127 gnd.n7126 585
R10043 gnd.n309 gnd.n308 585
R10044 gnd.n314 gnd.n308 585
R10045 gnd.n7121 gnd.n7120 585
R10046 gnd.n7120 gnd.n7119 585
R10047 gnd.n311 gnd.n280 585
R10048 gnd.n7219 gnd.n280 585
R10049 gnd.n4279 gnd.n4277 585
R10050 gnd.n4277 gnd.n4276 585
R10051 gnd.n4280 gnd.n1528 585
R10052 gnd.n4314 gnd.n1528 585
R10053 gnd.n4281 gnd.n1553 585
R10054 gnd.n1553 gnd.n1538 585
R10055 gnd.n1550 gnd.n1537 585
R10056 gnd.n4306 gnd.n1537 585
R10057 gnd.n4286 gnd.n4285 585
R10058 gnd.n4288 gnd.n4286 585
R10059 gnd.n1549 gnd.n1548 585
R10060 gnd.n1548 gnd.n1546 585
R10061 gnd.n4223 gnd.n1562 585
R10062 gnd.n4253 gnd.n1562 585
R10063 gnd.n4224 gnd.n4222 585
R10064 gnd.n4222 gnd.n1573 585
R10065 gnd.n1584 gnd.n1572 585
R10066 gnd.n4243 gnd.n1572 585
R10067 gnd.n4229 gnd.n4228 585
R10068 gnd.n4230 gnd.n4229 585
R10069 gnd.n1583 gnd.n1582 585
R10070 gnd.n1582 gnd.n1580 585
R10071 gnd.n4218 gnd.n4217 585
R10072 gnd.n4217 gnd.n4216 585
R10073 gnd.n1587 gnd.n1586 585
R10074 gnd.n1601 gnd.n1587 585
R10075 gnd.n1611 gnd.n1599 585
R10076 gnd.n4206 gnd.n1599 585
R10077 gnd.n4193 gnd.n4192 585
R10078 gnd.n4194 gnd.n4193 585
R10079 gnd.n1610 gnd.n1609 585
R10080 gnd.n1671 gnd.n1609 585
R10081 gnd.n4187 gnd.n4186 585
R10082 gnd.n4186 gnd.n4185 585
R10083 gnd.n1614 gnd.n1613 585
R10084 gnd.n1628 gnd.n1614 585
R10085 gnd.n1682 gnd.n1627 585
R10086 gnd.n4175 gnd.n1627 585
R10087 gnd.n4162 gnd.n4161 585
R10088 gnd.n4163 gnd.n4162 585
R10089 gnd.n1681 gnd.n1680 585
R10090 gnd.n1680 gnd.n1647 585
R10091 gnd.n4156 gnd.n1498 585
R10092 gnd.n4349 gnd.n1498 585
R10093 gnd.n6239 gnd.n6238 585
R10094 gnd.n6238 gnd.n6237 585
R10095 gnd.n6240 gnd.n924 585
R10096 gnd.n6147 gnd.n924 585
R10097 gnd.n6242 gnd.n6241 585
R10098 gnd.n6243 gnd.n6242 585
R10099 gnd.n925 gnd.n923 585
R10100 gnd.n923 gnd.n919 585
R10101 gnd.n906 gnd.n905 585
R10102 gnd.n910 gnd.n906 585
R10103 gnd.n6253 gnd.n6252 585
R10104 gnd.n6252 gnd.n6251 585
R10105 gnd.n6254 gnd.n900 585
R10106 gnd.n6136 gnd.n900 585
R10107 gnd.n6256 gnd.n6255 585
R10108 gnd.n6257 gnd.n6256 585
R10109 gnd.n901 gnd.n899 585
R10110 gnd.n6130 gnd.n899 585
R10111 gnd.n6111 gnd.n4936 585
R10112 gnd.n4936 gnd.n4935 585
R10113 gnd.n6113 gnd.n6112 585
R10114 gnd.n6114 gnd.n6113 585
R10115 gnd.n4937 gnd.n4934 585
R10116 gnd.n4934 gnd.n4930 585
R10117 gnd.n5818 gnd.n5817 585
R10118 gnd.n5817 gnd.n5816 585
R10119 gnd.n4944 gnd.n4943 585
R10120 gnd.n4953 gnd.n4944 585
R10121 gnd.n5807 gnd.n5806 585
R10122 gnd.n5806 gnd.n5805 585
R10123 gnd.n4951 gnd.n4950 585
R10124 gnd.n5793 gnd.n4951 585
R10125 gnd.n5768 gnd.n4968 585
R10126 gnd.n5761 gnd.n4968 585
R10127 gnd.n5770 gnd.n5769 585
R10128 gnd.n5771 gnd.n5770 585
R10129 gnd.n4969 gnd.n4967 585
R10130 gnd.n4977 gnd.n4967 585
R10131 gnd.n5744 gnd.n4989 585
R10132 gnd.n4989 gnd.n4976 585
R10133 gnd.n5746 gnd.n5745 585
R10134 gnd.n5747 gnd.n5746 585
R10135 gnd.n4990 gnd.n4988 585
R10136 gnd.n4988 gnd.n4984 585
R10137 gnd.n5732 gnd.n5731 585
R10138 gnd.n5731 gnd.n5730 585
R10139 gnd.n4995 gnd.n4994 585
R10140 gnd.n4999 gnd.n4995 585
R10141 gnd.n5716 gnd.n5715 585
R10142 gnd.n5717 gnd.n5716 585
R10143 gnd.n5009 gnd.n5008 585
R10144 gnd.n5707 gnd.n5008 585
R10145 gnd.n5681 gnd.n5024 585
R10146 gnd.n5024 gnd.n5016 585
R10147 gnd.n5683 gnd.n5682 585
R10148 gnd.n5684 gnd.n5683 585
R10149 gnd.n5025 gnd.n5023 585
R10150 gnd.n5029 gnd.n5023 585
R10151 gnd.n5662 gnd.n5661 585
R10152 gnd.n5663 gnd.n5662 585
R10153 gnd.n5041 gnd.n5040 585
R10154 gnd.n5040 gnd.n5036 585
R10155 gnd.n5652 gnd.n5651 585
R10156 gnd.n5653 gnd.n5652 585
R10157 gnd.n5049 gnd.n5048 585
R10158 gnd.n5053 gnd.n5048 585
R10159 gnd.n5630 gnd.n5065 585
R10160 gnd.n5409 gnd.n5065 585
R10161 gnd.n5632 gnd.n5631 585
R10162 gnd.n5633 gnd.n5632 585
R10163 gnd.n5066 gnd.n5064 585
R10164 gnd.n5064 gnd.n5060 585
R10165 gnd.n5621 gnd.n5620 585
R10166 gnd.n5622 gnd.n5621 585
R10167 gnd.n5074 gnd.n5073 585
R10168 gnd.n5079 gnd.n5073 585
R10169 gnd.n5599 gnd.n5091 585
R10170 gnd.n5091 gnd.n5078 585
R10171 gnd.n5601 gnd.n5600 585
R10172 gnd.n5602 gnd.n5601 585
R10173 gnd.n5092 gnd.n5090 585
R10174 gnd.n5090 gnd.n5086 585
R10175 gnd.n5590 gnd.n5589 585
R10176 gnd.n5591 gnd.n5590 585
R10177 gnd.n5100 gnd.n5099 585
R10178 gnd.n5474 gnd.n5099 585
R10179 gnd.n5568 gnd.n5116 585
R10180 gnd.n5116 gnd.n5104 585
R10181 gnd.n5570 gnd.n5569 585
R10182 gnd.n5571 gnd.n5570 585
R10183 gnd.n5117 gnd.n5115 585
R10184 gnd.n5115 gnd.n5111 585
R10185 gnd.n5559 gnd.n5558 585
R10186 gnd.n5560 gnd.n5559 585
R10187 gnd.n5124 gnd.n5123 585
R10188 gnd.n5129 gnd.n5123 585
R10189 gnd.n5537 gnd.n5142 585
R10190 gnd.n5142 gnd.n5128 585
R10191 gnd.n5539 gnd.n5538 585
R10192 gnd.n5540 gnd.n5539 585
R10193 gnd.n5143 gnd.n5141 585
R10194 gnd.n5141 gnd.n5137 585
R10195 gnd.n5528 gnd.n5527 585
R10196 gnd.n5529 gnd.n5528 585
R10197 gnd.n5150 gnd.n5149 585
R10198 gnd.n5154 gnd.n5149 585
R10199 gnd.n5505 gnd.n5171 585
R10200 gnd.n5171 gnd.n5153 585
R10201 gnd.n5507 gnd.n5506 585
R10202 gnd.n5508 gnd.n5507 585
R10203 gnd.n5172 gnd.n5170 585
R10204 gnd.n5170 gnd.n5161 585
R10205 gnd.n5500 gnd.n5499 585
R10206 gnd.n5499 gnd.n5498 585
R10207 gnd.n5219 gnd.n5218 585
R10208 gnd.n5220 gnd.n5219 585
R10209 gnd.n5373 gnd.n5372 585
R10210 gnd.n5374 gnd.n5373 585
R10211 gnd.n5229 gnd.n5228 585
R10212 gnd.n5228 gnd.n5227 585
R10213 gnd.n5368 gnd.n5367 585
R10214 gnd.n5367 gnd.n5366 585
R10215 gnd.n5232 gnd.n5231 585
R10216 gnd.n5233 gnd.n5232 585
R10217 gnd.n5357 gnd.n5356 585
R10218 gnd.n5358 gnd.n5357 585
R10219 gnd.n5240 gnd.n5239 585
R10220 gnd.n5349 gnd.n5239 585
R10221 gnd.n5352 gnd.n5351 585
R10222 gnd.n5351 gnd.n5350 585
R10223 gnd.n5243 gnd.n5242 585
R10224 gnd.n5244 gnd.n5243 585
R10225 gnd.n5338 gnd.n5337 585
R10226 gnd.n5336 gnd.n5262 585
R10227 gnd.n5335 gnd.n5261 585
R10228 gnd.n5340 gnd.n5261 585
R10229 gnd.n5334 gnd.n5333 585
R10230 gnd.n5332 gnd.n5331 585
R10231 gnd.n5330 gnd.n5329 585
R10232 gnd.n5328 gnd.n5327 585
R10233 gnd.n5326 gnd.n5325 585
R10234 gnd.n5324 gnd.n5323 585
R10235 gnd.n5322 gnd.n5321 585
R10236 gnd.n5320 gnd.n5319 585
R10237 gnd.n5318 gnd.n5317 585
R10238 gnd.n5316 gnd.n5315 585
R10239 gnd.n5314 gnd.n5313 585
R10240 gnd.n5312 gnd.n5311 585
R10241 gnd.n5310 gnd.n5309 585
R10242 gnd.n5308 gnd.n5307 585
R10243 gnd.n5306 gnd.n5305 585
R10244 gnd.n5304 gnd.n5303 585
R10245 gnd.n5302 gnd.n5301 585
R10246 gnd.n5300 gnd.n5299 585
R10247 gnd.n5298 gnd.n5297 585
R10248 gnd.n5296 gnd.n5295 585
R10249 gnd.n5294 gnd.n5293 585
R10250 gnd.n5292 gnd.n5291 585
R10251 gnd.n5249 gnd.n5248 585
R10252 gnd.n5343 gnd.n5342 585
R10253 gnd.n6155 gnd.n6154 585
R10254 gnd.n6156 gnd.n4912 585
R10255 gnd.n6158 gnd.n6157 585
R10256 gnd.n6160 gnd.n4911 585
R10257 gnd.n6162 gnd.n6161 585
R10258 gnd.n6163 gnd.n4902 585
R10259 gnd.n6165 gnd.n6164 585
R10260 gnd.n6167 gnd.n4900 585
R10261 gnd.n6169 gnd.n6168 585
R10262 gnd.n6170 gnd.n4895 585
R10263 gnd.n6172 gnd.n6171 585
R10264 gnd.n6174 gnd.n4893 585
R10265 gnd.n6176 gnd.n6175 585
R10266 gnd.n6177 gnd.n4888 585
R10267 gnd.n6179 gnd.n6178 585
R10268 gnd.n6181 gnd.n4886 585
R10269 gnd.n6183 gnd.n6182 585
R10270 gnd.n6184 gnd.n4881 585
R10271 gnd.n6186 gnd.n6185 585
R10272 gnd.n6188 gnd.n4879 585
R10273 gnd.n6190 gnd.n6189 585
R10274 gnd.n6191 gnd.n4874 585
R10275 gnd.n6193 gnd.n6192 585
R10276 gnd.n6195 gnd.n4872 585
R10277 gnd.n6197 gnd.n6196 585
R10278 gnd.n6198 gnd.n4870 585
R10279 gnd.n6199 gnd.n929 585
R10280 gnd.n4833 gnd.n929 585
R10281 gnd.n6150 gnd.n931 585
R10282 gnd.n6237 gnd.n931 585
R10283 gnd.n6149 gnd.n6148 585
R10284 gnd.n6148 gnd.n6147 585
R10285 gnd.n6146 gnd.n921 585
R10286 gnd.n6243 gnd.n921 585
R10287 gnd.n6140 gnd.n4917 585
R10288 gnd.n6140 gnd.n919 585
R10289 gnd.n6142 gnd.n6141 585
R10290 gnd.n6141 gnd.n910 585
R10291 gnd.n6139 gnd.n908 585
R10292 gnd.n6251 gnd.n908 585
R10293 gnd.n6138 gnd.n6137 585
R10294 gnd.n6137 gnd.n6136 585
R10295 gnd.n4919 gnd.n897 585
R10296 gnd.n6257 gnd.n897 585
R10297 gnd.n6132 gnd.n6131 585
R10298 gnd.n6131 gnd.n6130 585
R10299 gnd.n4922 gnd.n4921 585
R10300 gnd.n4935 gnd.n4922 585
R10301 gnd.n5782 gnd.n4932 585
R10302 gnd.n6114 gnd.n4932 585
R10303 gnd.n5784 gnd.n5783 585
R10304 gnd.n5783 gnd.n4930 585
R10305 gnd.n5785 gnd.n4946 585
R10306 gnd.n5816 gnd.n4946 585
R10307 gnd.n5787 gnd.n5786 585
R10308 gnd.n5786 gnd.n4953 585
R10309 gnd.n5788 gnd.n4952 585
R10310 gnd.n5805 gnd.n4952 585
R10311 gnd.n5790 gnd.n5789 585
R10312 gnd.n5793 gnd.n5790 585
R10313 gnd.n4962 gnd.n4961 585
R10314 gnd.n5761 gnd.n4961 585
R10315 gnd.n5773 gnd.n5772 585
R10316 gnd.n5772 gnd.n5771 585
R10317 gnd.n4965 gnd.n4964 585
R10318 gnd.n4977 gnd.n4965 585
R10319 gnd.n5697 gnd.n5696 585
R10320 gnd.n5696 gnd.n4976 585
R10321 gnd.n5698 gnd.n4986 585
R10322 gnd.n5747 gnd.n4986 585
R10323 gnd.n5700 gnd.n5699 585
R10324 gnd.n5699 gnd.n4984 585
R10325 gnd.n5701 gnd.n4996 585
R10326 gnd.n5730 gnd.n4996 585
R10327 gnd.n5703 gnd.n5702 585
R10328 gnd.n5702 gnd.n4999 585
R10329 gnd.n5704 gnd.n5006 585
R10330 gnd.n5717 gnd.n5006 585
R10331 gnd.n5706 gnd.n5705 585
R10332 gnd.n5707 gnd.n5706 585
R10333 gnd.n5018 gnd.n5017 585
R10334 gnd.n5017 gnd.n5016 585
R10335 gnd.n5686 gnd.n5685 585
R10336 gnd.n5685 gnd.n5684 585
R10337 gnd.n5021 gnd.n5020 585
R10338 gnd.n5029 gnd.n5021 585
R10339 gnd.n5401 gnd.n5038 585
R10340 gnd.n5663 gnd.n5038 585
R10341 gnd.n5404 gnd.n5403 585
R10342 gnd.n5403 gnd.n5036 585
R10343 gnd.n5405 gnd.n5047 585
R10344 gnd.n5653 gnd.n5047 585
R10345 gnd.n5408 gnd.n5407 585
R10346 gnd.n5408 gnd.n5053 585
R10347 gnd.n5411 gnd.n5410 585
R10348 gnd.n5410 gnd.n5409 585
R10349 gnd.n5412 gnd.n5062 585
R10350 gnd.n5633 gnd.n5062 585
R10351 gnd.n5400 gnd.n5399 585
R10352 gnd.n5399 gnd.n5060 585
R10353 gnd.n5464 gnd.n5072 585
R10354 gnd.n5622 gnd.n5072 585
R10355 gnd.n5466 gnd.n5465 585
R10356 gnd.n5466 gnd.n5079 585
R10357 gnd.n5468 gnd.n5467 585
R10358 gnd.n5467 gnd.n5078 585
R10359 gnd.n5469 gnd.n5088 585
R10360 gnd.n5602 gnd.n5088 585
R10361 gnd.n5471 gnd.n5470 585
R10362 gnd.n5470 gnd.n5086 585
R10363 gnd.n5472 gnd.n5098 585
R10364 gnd.n5591 gnd.n5098 585
R10365 gnd.n5475 gnd.n5473 585
R10366 gnd.n5475 gnd.n5474 585
R10367 gnd.n5477 gnd.n5476 585
R10368 gnd.n5476 gnd.n5104 585
R10369 gnd.n5478 gnd.n5113 585
R10370 gnd.n5571 gnd.n5113 585
R10371 gnd.n5480 gnd.n5479 585
R10372 gnd.n5479 gnd.n5111 585
R10373 gnd.n5481 gnd.n5122 585
R10374 gnd.n5560 gnd.n5122 585
R10375 gnd.n5483 gnd.n5482 585
R10376 gnd.n5483 gnd.n5129 585
R10377 gnd.n5485 gnd.n5484 585
R10378 gnd.n5484 gnd.n5128 585
R10379 gnd.n5486 gnd.n5139 585
R10380 gnd.n5540 gnd.n5139 585
R10381 gnd.n5488 gnd.n5487 585
R10382 gnd.n5487 gnd.n5137 585
R10383 gnd.n5489 gnd.n5148 585
R10384 gnd.n5529 gnd.n5148 585
R10385 gnd.n5491 gnd.n5490 585
R10386 gnd.n5491 gnd.n5154 585
R10387 gnd.n5493 gnd.n5492 585
R10388 gnd.n5492 gnd.n5153 585
R10389 gnd.n5494 gnd.n5169 585
R10390 gnd.n5508 gnd.n5169 585
R10391 gnd.n5495 gnd.n5222 585
R10392 gnd.n5222 gnd.n5161 585
R10393 gnd.n5497 gnd.n5496 585
R10394 gnd.n5498 gnd.n5497 585
R10395 gnd.n5223 gnd.n5221 585
R10396 gnd.n5221 gnd.n5220 585
R10397 gnd.n5376 gnd.n5375 585
R10398 gnd.n5375 gnd.n5374 585
R10399 gnd.n5226 gnd.n5225 585
R10400 gnd.n5227 gnd.n5226 585
R10401 gnd.n5365 gnd.n5364 585
R10402 gnd.n5366 gnd.n5365 585
R10403 gnd.n5235 gnd.n5234 585
R10404 gnd.n5234 gnd.n5233 585
R10405 gnd.n5360 gnd.n5359 585
R10406 gnd.n5359 gnd.n5358 585
R10407 gnd.n5238 gnd.n5237 585
R10408 gnd.n5349 gnd.n5238 585
R10409 gnd.n5348 gnd.n5347 585
R10410 gnd.n5350 gnd.n5348 585
R10411 gnd.n5246 gnd.n5245 585
R10412 gnd.n5245 gnd.n5244 585
R10413 gnd.n6235 gnd.n6234 585
R10414 gnd.n6236 gnd.n6235 585
R10415 gnd.n4836 gnd.n4834 585
R10416 gnd.n4834 gnd.n930 585
R10417 gnd.n918 gnd.n917 585
R10418 gnd.n922 gnd.n918 585
R10419 gnd.n6246 gnd.n6245 585
R10420 gnd.n6245 gnd.n6244 585
R10421 gnd.n6247 gnd.n912 585
R10422 gnd.n6099 gnd.n912 585
R10423 gnd.n6249 gnd.n6248 585
R10424 gnd.n6250 gnd.n6249 585
R10425 gnd.n913 gnd.n911 585
R10426 gnd.n911 gnd.n907 585
R10427 gnd.n6125 gnd.n6124 585
R10428 gnd.n6124 gnd.n898 585
R10429 gnd.n6126 gnd.n4925 585
R10430 gnd.n4925 gnd.n896 585
R10431 gnd.n6128 gnd.n6127 585
R10432 gnd.n6129 gnd.n6128 585
R10433 gnd.n4926 gnd.n4924 585
R10434 gnd.n4933 gnd.n4924 585
R10435 gnd.n6117 gnd.n6116 585
R10436 gnd.n6116 gnd.n6115 585
R10437 gnd.n4929 gnd.n4928 585
R10438 gnd.n5815 gnd.n4929 585
R10439 gnd.n5801 gnd.n4955 585
R10440 gnd.n4955 gnd.n4945 585
R10441 gnd.n5803 gnd.n5802 585
R10442 gnd.n5804 gnd.n5803 585
R10443 gnd.n4956 gnd.n4954 585
R10444 gnd.n5792 gnd.n4954 585
R10445 gnd.n5796 gnd.n5795 585
R10446 gnd.n5795 gnd.n5794 585
R10447 gnd.n4959 gnd.n4958 585
R10448 gnd.n5762 gnd.n4959 585
R10449 gnd.n5755 gnd.n4979 585
R10450 gnd.n4979 gnd.n4966 585
R10451 gnd.n5757 gnd.n5756 585
R10452 gnd.n5758 gnd.n5757 585
R10453 gnd.n4980 gnd.n4978 585
R10454 gnd.n4987 gnd.n4978 585
R10455 gnd.n5750 gnd.n5749 585
R10456 gnd.n5749 gnd.n5748 585
R10457 gnd.n4983 gnd.n4982 585
R10458 gnd.n5729 gnd.n4983 585
R10459 gnd.n5725 gnd.n5724 585
R10460 gnd.n5726 gnd.n5725 585
R10461 gnd.n5001 gnd.n5000 585
R10462 gnd.n5007 gnd.n5000 585
R10463 gnd.n5720 gnd.n5719 585
R10464 gnd.n5719 gnd.n5718 585
R10465 gnd.n5004 gnd.n5003 585
R10466 gnd.n5708 gnd.n5004 585
R10467 gnd.n5671 gnd.n5031 585
R10468 gnd.n5031 gnd.n5022 585
R10469 gnd.n5673 gnd.n5672 585
R10470 gnd.n5674 gnd.n5673 585
R10471 gnd.n5032 gnd.n5030 585
R10472 gnd.n5039 gnd.n5030 585
R10473 gnd.n5666 gnd.n5665 585
R10474 gnd.n5665 gnd.n5664 585
R10475 gnd.n5035 gnd.n5034 585
R10476 gnd.n5654 gnd.n5035 585
R10477 gnd.n5641 gnd.n5055 585
R10478 gnd.n5055 gnd.n5046 585
R10479 gnd.n5643 gnd.n5642 585
R10480 gnd.n5644 gnd.n5643 585
R10481 gnd.n5056 gnd.n5054 585
R10482 gnd.n5063 gnd.n5054 585
R10483 gnd.n5636 gnd.n5635 585
R10484 gnd.n5635 gnd.n5634 585
R10485 gnd.n5059 gnd.n5058 585
R10486 gnd.n5623 gnd.n5059 585
R10487 gnd.n5610 gnd.n5081 585
R10488 gnd.n5081 gnd.n5071 585
R10489 gnd.n5612 gnd.n5611 585
R10490 gnd.n5613 gnd.n5612 585
R10491 gnd.n5082 gnd.n5080 585
R10492 gnd.n5089 gnd.n5080 585
R10493 gnd.n5605 gnd.n5604 585
R10494 gnd.n5604 gnd.n5603 585
R10495 gnd.n5085 gnd.n5084 585
R10496 gnd.n5592 gnd.n5085 585
R10497 gnd.n5579 gnd.n5106 585
R10498 gnd.n5106 gnd.n5097 585
R10499 gnd.n5581 gnd.n5580 585
R10500 gnd.n5582 gnd.n5581 585
R10501 gnd.n5107 gnd.n5105 585
R10502 gnd.n5114 gnd.n5105 585
R10503 gnd.n5574 gnd.n5573 585
R10504 gnd.n5573 gnd.n5572 585
R10505 gnd.n5110 gnd.n5109 585
R10506 gnd.n5561 gnd.n5110 585
R10507 gnd.n5548 gnd.n5132 585
R10508 gnd.n5132 gnd.n5131 585
R10509 gnd.n5550 gnd.n5549 585
R10510 gnd.n5551 gnd.n5550 585
R10511 gnd.n5133 gnd.n5130 585
R10512 gnd.n5140 gnd.n5130 585
R10513 gnd.n5543 gnd.n5542 585
R10514 gnd.n5542 gnd.n5541 585
R10515 gnd.n5136 gnd.n5135 585
R10516 gnd.n5530 gnd.n5136 585
R10517 gnd.n5517 gnd.n5157 585
R10518 gnd.n5157 gnd.n5156 585
R10519 gnd.n5519 gnd.n5518 585
R10520 gnd.n5520 gnd.n5519 585
R10521 gnd.n5513 gnd.n5155 585
R10522 gnd.n5512 gnd.n5511 585
R10523 gnd.n5160 gnd.n5159 585
R10524 gnd.n5509 gnd.n5160 585
R10525 gnd.n5182 gnd.n5181 585
R10526 gnd.n5185 gnd.n5184 585
R10527 gnd.n5183 gnd.n5178 585
R10528 gnd.n5190 gnd.n5189 585
R10529 gnd.n5192 gnd.n5191 585
R10530 gnd.n5195 gnd.n5194 585
R10531 gnd.n5193 gnd.n5176 585
R10532 gnd.n5200 gnd.n5199 585
R10533 gnd.n5202 gnd.n5201 585
R10534 gnd.n5205 gnd.n5204 585
R10535 gnd.n5203 gnd.n5174 585
R10536 gnd.n5210 gnd.n5209 585
R10537 gnd.n5214 gnd.n5211 585
R10538 gnd.n5215 gnd.n5152 585
R10539 gnd.n6204 gnd.n6203 585
R10540 gnd.n6206 gnd.n4865 585
R10541 gnd.n6208 gnd.n6207 585
R10542 gnd.n6209 gnd.n4858 585
R10543 gnd.n6211 gnd.n6210 585
R10544 gnd.n6213 gnd.n4856 585
R10545 gnd.n6215 gnd.n6214 585
R10546 gnd.n6216 gnd.n4851 585
R10547 gnd.n6218 gnd.n6217 585
R10548 gnd.n6220 gnd.n4849 585
R10549 gnd.n6222 gnd.n6221 585
R10550 gnd.n6223 gnd.n4844 585
R10551 gnd.n6225 gnd.n6224 585
R10552 gnd.n6227 gnd.n4842 585
R10553 gnd.n6229 gnd.n6228 585
R10554 gnd.n6230 gnd.n4840 585
R10555 gnd.n6231 gnd.n4835 585
R10556 gnd.n4835 gnd.n4833 585
R10557 gnd.n6093 gnd.n932 585
R10558 gnd.n6236 gnd.n932 585
R10559 gnd.n6095 gnd.n6094 585
R10560 gnd.n6095 gnd.n930 585
R10561 gnd.n6097 gnd.n6096 585
R10562 gnd.n6096 gnd.n922 585
R10563 gnd.n6098 gnd.n920 585
R10564 gnd.n6244 gnd.n920 585
R10565 gnd.n6101 gnd.n6100 585
R10566 gnd.n6100 gnd.n6099 585
R10567 gnd.n6102 gnd.n909 585
R10568 gnd.n6250 gnd.n909 585
R10569 gnd.n6104 gnd.n6103 585
R10570 gnd.n6104 gnd.n907 585
R10571 gnd.n6105 gnd.n5828 585
R10572 gnd.n6105 gnd.n898 585
R10573 gnd.n6107 gnd.n6106 585
R10574 gnd.n6106 gnd.n896 585
R10575 gnd.n6108 gnd.n4923 585
R10576 gnd.n6129 gnd.n4923 585
R10577 gnd.n5825 gnd.n5824 585
R10578 gnd.n5824 gnd.n4933 585
R10579 gnd.n5823 gnd.n4931 585
R10580 gnd.n6115 gnd.n4931 585
R10581 gnd.n5814 gnd.n4941 585
R10582 gnd.n5815 gnd.n5814 585
R10583 gnd.n5813 gnd.n5812 585
R10584 gnd.n5813 gnd.n4945 585
R10585 gnd.n5811 gnd.n4947 585
R10586 gnd.n5804 gnd.n4947 585
R10587 gnd.n5791 gnd.n4948 585
R10588 gnd.n5792 gnd.n5791 585
R10589 gnd.n5765 gnd.n4960 585
R10590 gnd.n5794 gnd.n4960 585
R10591 gnd.n5764 gnd.n5763 585
R10592 gnd.n5763 gnd.n5762 585
R10593 gnd.n5760 gnd.n4973 585
R10594 gnd.n5760 gnd.n4966 585
R10595 gnd.n5759 gnd.n4975 585
R10596 gnd.n5759 gnd.n5758 585
R10597 gnd.n5738 gnd.n4974 585
R10598 gnd.n4987 gnd.n4974 585
R10599 gnd.n5737 gnd.n4985 585
R10600 gnd.n5748 gnd.n4985 585
R10601 gnd.n5728 gnd.n4992 585
R10602 gnd.n5729 gnd.n5728 585
R10603 gnd.n5727 gnd.n4998 585
R10604 gnd.n5727 gnd.n5726 585
R10605 gnd.n5712 gnd.n4997 585
R10606 gnd.n5007 gnd.n4997 585
R10607 gnd.n5711 gnd.n5005 585
R10608 gnd.n5718 gnd.n5005 585
R10609 gnd.n5710 gnd.n5709 585
R10610 gnd.n5709 gnd.n5708 585
R10611 gnd.n5015 gnd.n5012 585
R10612 gnd.n5022 gnd.n5015 585
R10613 gnd.n5676 gnd.n5675 585
R10614 gnd.n5675 gnd.n5674 585
R10615 gnd.n5028 gnd.n5027 585
R10616 gnd.n5039 gnd.n5028 585
R10617 gnd.n5657 gnd.n5037 585
R10618 gnd.n5664 gnd.n5037 585
R10619 gnd.n5656 gnd.n5655 585
R10620 gnd.n5655 gnd.n5654 585
R10621 gnd.n5045 gnd.n5043 585
R10622 gnd.n5046 gnd.n5045 585
R10623 gnd.n5646 gnd.n5645 585
R10624 gnd.n5645 gnd.n5644 585
R10625 gnd.n5052 gnd.n5051 585
R10626 gnd.n5063 gnd.n5052 585
R10627 gnd.n5626 gnd.n5061 585
R10628 gnd.n5634 gnd.n5061 585
R10629 gnd.n5625 gnd.n5624 585
R10630 gnd.n5624 gnd.n5623 585
R10631 gnd.n5070 gnd.n5068 585
R10632 gnd.n5071 gnd.n5070 585
R10633 gnd.n5615 gnd.n5614 585
R10634 gnd.n5614 gnd.n5613 585
R10635 gnd.n5077 gnd.n5076 585
R10636 gnd.n5089 gnd.n5077 585
R10637 gnd.n5595 gnd.n5087 585
R10638 gnd.n5603 gnd.n5087 585
R10639 gnd.n5594 gnd.n5593 585
R10640 gnd.n5593 gnd.n5592 585
R10641 gnd.n5096 gnd.n5094 585
R10642 gnd.n5097 gnd.n5096 585
R10643 gnd.n5584 gnd.n5583 585
R10644 gnd.n5583 gnd.n5582 585
R10645 gnd.n5103 gnd.n5102 585
R10646 gnd.n5114 gnd.n5103 585
R10647 gnd.n5564 gnd.n5112 585
R10648 gnd.n5572 gnd.n5112 585
R10649 gnd.n5563 gnd.n5562 585
R10650 gnd.n5562 gnd.n5561 585
R10651 gnd.n5121 gnd.n5119 585
R10652 gnd.n5131 gnd.n5121 585
R10653 gnd.n5553 gnd.n5552 585
R10654 gnd.n5552 gnd.n5551 585
R10655 gnd.n5127 gnd.n5126 585
R10656 gnd.n5140 gnd.n5127 585
R10657 gnd.n5533 gnd.n5138 585
R10658 gnd.n5541 gnd.n5138 585
R10659 gnd.n5532 gnd.n5531 585
R10660 gnd.n5531 gnd.n5530 585
R10661 gnd.n5147 gnd.n5145 585
R10662 gnd.n5156 gnd.n5147 585
R10663 gnd.n5522 gnd.n5521 585
R10664 gnd.n5521 gnd.n5520 585
R10665 gnd.n4596 gnd.n4595 585
R10666 gnd.n4595 gnd.n4594 585
R10667 gnd.n4597 gnd.n1264 585
R10668 gnd.n2821 gnd.n1264 585
R10669 gnd.n4599 gnd.n4598 585
R10670 gnd.n4600 gnd.n4599 585
R10671 gnd.n1249 gnd.n1248 585
R10672 gnd.n2781 gnd.n1249 585
R10673 gnd.n4608 gnd.n4607 585
R10674 gnd.n4607 gnd.n4606 585
R10675 gnd.n4609 gnd.n1243 585
R10676 gnd.n2772 gnd.n1243 585
R10677 gnd.n4611 gnd.n4610 585
R10678 gnd.n4612 gnd.n4611 585
R10679 gnd.n1228 gnd.n1227 585
R10680 gnd.n2764 gnd.n1228 585
R10681 gnd.n4620 gnd.n4619 585
R10682 gnd.n4619 gnd.n4618 585
R10683 gnd.n4621 gnd.n1222 585
R10684 gnd.n2694 gnd.n1222 585
R10685 gnd.n4623 gnd.n4622 585
R10686 gnd.n4624 gnd.n4623 585
R10687 gnd.n1207 gnd.n1206 585
R10688 gnd.n2682 gnd.n1207 585
R10689 gnd.n4632 gnd.n4631 585
R10690 gnd.n4631 gnd.n4630 585
R10691 gnd.n4633 gnd.n1201 585
R10692 gnd.n2677 gnd.n1201 585
R10693 gnd.n4635 gnd.n4634 585
R10694 gnd.n4636 gnd.n4635 585
R10695 gnd.n1186 gnd.n1185 585
R10696 gnd.n2708 gnd.n1186 585
R10697 gnd.n4644 gnd.n4643 585
R10698 gnd.n4643 gnd.n4642 585
R10699 gnd.n4645 gnd.n1180 585
R10700 gnd.n2669 gnd.n1180 585
R10701 gnd.n4647 gnd.n4646 585
R10702 gnd.n4648 gnd.n4647 585
R10703 gnd.n1165 gnd.n1164 585
R10704 gnd.n2661 gnd.n1165 585
R10705 gnd.n4656 gnd.n4655 585
R10706 gnd.n4655 gnd.n4654 585
R10707 gnd.n4657 gnd.n1160 585
R10708 gnd.n2652 gnd.n1160 585
R10709 gnd.n4659 gnd.n4658 585
R10710 gnd.n4660 gnd.n4659 585
R10711 gnd.n1161 gnd.n1145 585
R10712 gnd.n2644 gnd.n1145 585
R10713 gnd.n4668 gnd.n4667 585
R10714 gnd.n4667 gnd.n4666 585
R10715 gnd.n4669 gnd.n1142 585
R10716 gnd.n2612 gnd.n1142 585
R10717 gnd.n4672 gnd.n4671 585
R10718 gnd.n4673 gnd.n4672 585
R10719 gnd.n1143 gnd.n1127 585
R10720 gnd.n2621 gnd.n1127 585
R10721 gnd.n4681 gnd.n4680 585
R10722 gnd.n4680 gnd.n4679 585
R10723 gnd.n4682 gnd.n1123 585
R10724 gnd.n2627 gnd.n1123 585
R10725 gnd.n4684 gnd.n4683 585
R10726 gnd.n4685 gnd.n4684 585
R10727 gnd.n1108 gnd.n1107 585
R10728 gnd.n2633 gnd.n1108 585
R10729 gnd.n4693 gnd.n4692 585
R10730 gnd.n4692 gnd.n4691 585
R10731 gnd.n4694 gnd.n1102 585
R10732 gnd.n2577 gnd.n1102 585
R10733 gnd.n4696 gnd.n4695 585
R10734 gnd.n4697 gnd.n4696 585
R10735 gnd.n1087 gnd.n1086 585
R10736 gnd.n1098 gnd.n1087 585
R10737 gnd.n4705 gnd.n4704 585
R10738 gnd.n4704 gnd.n4703 585
R10739 gnd.n4706 gnd.n1081 585
R10740 gnd.n1081 gnd.n1080 585
R10741 gnd.n4708 gnd.n4707 585
R10742 gnd.n4709 gnd.n4708 585
R10743 gnd.n1066 gnd.n1065 585
R10744 gnd.n1070 gnd.n1066 585
R10745 gnd.n4717 gnd.n4716 585
R10746 gnd.n4716 gnd.n4715 585
R10747 gnd.n4718 gnd.n1060 585
R10748 gnd.n1067 gnd.n1060 585
R10749 gnd.n4720 gnd.n4719 585
R10750 gnd.n4721 gnd.n4720 585
R10751 gnd.n1047 gnd.n1046 585
R10752 gnd.n1057 gnd.n1047 585
R10753 gnd.n4729 gnd.n4728 585
R10754 gnd.n4728 gnd.n4727 585
R10755 gnd.n4730 gnd.n1041 585
R10756 gnd.n1041 gnd.n1040 585
R10757 gnd.n4732 gnd.n4731 585
R10758 gnd.n4733 gnd.n4732 585
R10759 gnd.n1026 gnd.n1025 585
R10760 gnd.n1029 gnd.n1026 585
R10761 gnd.n4741 gnd.n4740 585
R10762 gnd.n4740 gnd.n4739 585
R10763 gnd.n4742 gnd.n1020 585
R10764 gnd.n1020 gnd.n1017 585
R10765 gnd.n4744 gnd.n4743 585
R10766 gnd.n4745 gnd.n4744 585
R10767 gnd.n1021 gnd.n1019 585
R10768 gnd.n1019 gnd.n1015 585
R10769 gnd.n2534 gnd.n2533 585
R10770 gnd.n2535 gnd.n2534 585
R10771 gnd.n2529 gnd.n964 585
R10772 gnd.n964 gnd.n961 585
R10773 gnd.n4830 gnd.n4829 585
R10774 gnd.n4828 gnd.n963 585
R10775 gnd.n4827 gnd.n962 585
R10776 gnd.n4832 gnd.n962 585
R10777 gnd.n4826 gnd.n4825 585
R10778 gnd.n4824 gnd.n4823 585
R10779 gnd.n4822 gnd.n4821 585
R10780 gnd.n4820 gnd.n4819 585
R10781 gnd.n4818 gnd.n4817 585
R10782 gnd.n4816 gnd.n4815 585
R10783 gnd.n4814 gnd.n4813 585
R10784 gnd.n4812 gnd.n4811 585
R10785 gnd.n4810 gnd.n4809 585
R10786 gnd.n4808 gnd.n4807 585
R10787 gnd.n4806 gnd.n4805 585
R10788 gnd.n4804 gnd.n4803 585
R10789 gnd.n4802 gnd.n4801 585
R10790 gnd.n4800 gnd.n4799 585
R10791 gnd.n4798 gnd.n4797 585
R10792 gnd.n4795 gnd.n4794 585
R10793 gnd.n4793 gnd.n4792 585
R10794 gnd.n4791 gnd.n4790 585
R10795 gnd.n4789 gnd.n4788 585
R10796 gnd.n4787 gnd.n4786 585
R10797 gnd.n4785 gnd.n4784 585
R10798 gnd.n4783 gnd.n4782 585
R10799 gnd.n4781 gnd.n4780 585
R10800 gnd.n4779 gnd.n4778 585
R10801 gnd.n4777 gnd.n4776 585
R10802 gnd.n4775 gnd.n4774 585
R10803 gnd.n4773 gnd.n4772 585
R10804 gnd.n4771 gnd.n4770 585
R10805 gnd.n4769 gnd.n4768 585
R10806 gnd.n4767 gnd.n4766 585
R10807 gnd.n4765 gnd.n4764 585
R10808 gnd.n4763 gnd.n4762 585
R10809 gnd.n4761 gnd.n4760 585
R10810 gnd.n4759 gnd.n1003 585
R10811 gnd.n1007 gnd.n1004 585
R10812 gnd.n4755 gnd.n4754 585
R10813 gnd.n2311 gnd.n2310 585
R10814 gnd.n2829 gnd.n2828 585
R10815 gnd.n2831 gnd.n2830 585
R10816 gnd.n2833 gnd.n2832 585
R10817 gnd.n2835 gnd.n2834 585
R10818 gnd.n2837 gnd.n2836 585
R10819 gnd.n2839 gnd.n2838 585
R10820 gnd.n2841 gnd.n2840 585
R10821 gnd.n2843 gnd.n2842 585
R10822 gnd.n2845 gnd.n2844 585
R10823 gnd.n2847 gnd.n2846 585
R10824 gnd.n2849 gnd.n2848 585
R10825 gnd.n2851 gnd.n2850 585
R10826 gnd.n2853 gnd.n2852 585
R10827 gnd.n2855 gnd.n2854 585
R10828 gnd.n2857 gnd.n2856 585
R10829 gnd.n2859 gnd.n2858 585
R10830 gnd.n2861 gnd.n2860 585
R10831 gnd.n2863 gnd.n2862 585
R10832 gnd.n2866 gnd.n2865 585
R10833 gnd.n2864 gnd.n2289 585
R10834 gnd.n3643 gnd.n3642 585
R10835 gnd.n3645 gnd.n3644 585
R10836 gnd.n3647 gnd.n3646 585
R10837 gnd.n3649 gnd.n3648 585
R10838 gnd.n3651 gnd.n3650 585
R10839 gnd.n3653 gnd.n3652 585
R10840 gnd.n3655 gnd.n3654 585
R10841 gnd.n3657 gnd.n3656 585
R10842 gnd.n3659 gnd.n3658 585
R10843 gnd.n3661 gnd.n3660 585
R10844 gnd.n3663 gnd.n3662 585
R10845 gnd.n3665 gnd.n3664 585
R10846 gnd.n3666 gnd.n2270 585
R10847 gnd.n3668 gnd.n3667 585
R10848 gnd.n2271 gnd.n2269 585
R10849 gnd.n2272 gnd.n1269 585
R10850 gnd.n3670 gnd.n1269 585
R10851 gnd.n2824 gnd.n1271 585
R10852 gnd.n4594 gnd.n1271 585
R10853 gnd.n2823 gnd.n2822 585
R10854 gnd.n2822 gnd.n2821 585
R10855 gnd.n2315 gnd.n1262 585
R10856 gnd.n4600 gnd.n1262 585
R10857 gnd.n2780 gnd.n2779 585
R10858 gnd.n2781 gnd.n2780 585
R10859 gnd.n2321 gnd.n1251 585
R10860 gnd.n4606 gnd.n1251 585
R10861 gnd.n2774 gnd.n2773 585
R10862 gnd.n2773 gnd.n2772 585
R10863 gnd.n2323 gnd.n1240 585
R10864 gnd.n4612 gnd.n1240 585
R10865 gnd.n2690 gnd.n2327 585
R10866 gnd.n2764 gnd.n2327 585
R10867 gnd.n2691 gnd.n1230 585
R10868 gnd.n4618 gnd.n1230 585
R10869 gnd.n2693 gnd.n2692 585
R10870 gnd.n2694 gnd.n2693 585
R10871 gnd.n2347 gnd.n1219 585
R10872 gnd.n4624 gnd.n1219 585
R10873 gnd.n2684 gnd.n2683 585
R10874 gnd.n2683 gnd.n2682 585
R10875 gnd.n2680 gnd.n1209 585
R10876 gnd.n4630 gnd.n1209 585
R10877 gnd.n2679 gnd.n2678 585
R10878 gnd.n2678 gnd.n2677 585
R10879 gnd.n2349 gnd.n1198 585
R10880 gnd.n4636 gnd.n1198 585
R10881 gnd.n2673 gnd.n2339 585
R10882 gnd.n2708 gnd.n2339 585
R10883 gnd.n2672 gnd.n1188 585
R10884 gnd.n4642 gnd.n1188 585
R10885 gnd.n2671 gnd.n2670 585
R10886 gnd.n2670 gnd.n2669 585
R10887 gnd.n2351 gnd.n1177 585
R10888 gnd.n4648 gnd.n1177 585
R10889 gnd.n2660 gnd.n2659 585
R10890 gnd.n2661 gnd.n2660 585
R10891 gnd.n2357 gnd.n1167 585
R10892 gnd.n4654 gnd.n1167 585
R10893 gnd.n2654 gnd.n2653 585
R10894 gnd.n2653 gnd.n2652 585
R10895 gnd.n2359 gnd.n1157 585
R10896 gnd.n4660 gnd.n1157 585
R10897 gnd.n2608 gnd.n2363 585
R10898 gnd.n2644 gnd.n2363 585
R10899 gnd.n2609 gnd.n1147 585
R10900 gnd.n4666 gnd.n1147 585
R10901 gnd.n2611 gnd.n2610 585
R10902 gnd.n2612 gnd.n2611 585
R10903 gnd.n2587 gnd.n1139 585
R10904 gnd.n4673 gnd.n1139 585
R10905 gnd.n2623 gnd.n2622 585
R10906 gnd.n2622 gnd.n2621 585
R10907 gnd.n2624 gnd.n1129 585
R10908 gnd.n4679 gnd.n1129 585
R10909 gnd.n2626 gnd.n2625 585
R10910 gnd.n2627 gnd.n2626 585
R10911 gnd.n2405 gnd.n1120 585
R10912 gnd.n4685 gnd.n1120 585
R10913 gnd.n2581 gnd.n2399 585
R10914 gnd.n2633 gnd.n2399 585
R10915 gnd.n2580 gnd.n1110 585
R10916 gnd.n4691 gnd.n1110 585
R10917 gnd.n2579 gnd.n2578 585
R10918 gnd.n2578 gnd.n2577 585
R10919 gnd.n2407 gnd.n1099 585
R10920 gnd.n4697 gnd.n1099 585
R10921 gnd.n2441 gnd.n2440 585
R10922 gnd.n2440 gnd.n1098 585
R10923 gnd.n2439 gnd.n1088 585
R10924 gnd.n4703 gnd.n1088 585
R10925 gnd.n2438 gnd.n2437 585
R10926 gnd.n2437 gnd.n1080 585
R10927 gnd.n2409 gnd.n1078 585
R10928 gnd.n4709 gnd.n1078 585
R10929 gnd.n2433 gnd.n2432 585
R10930 gnd.n2432 gnd.n1070 585
R10931 gnd.n2431 gnd.n1068 585
R10932 gnd.n4715 gnd.n1068 585
R10933 gnd.n2430 gnd.n2429 585
R10934 gnd.n2429 gnd.n1067 585
R10935 gnd.n2411 gnd.n1058 585
R10936 gnd.n4721 gnd.n1058 585
R10937 gnd.n2425 gnd.n2424 585
R10938 gnd.n2424 gnd.n1057 585
R10939 gnd.n2423 gnd.n1048 585
R10940 gnd.n4727 gnd.n1048 585
R10941 gnd.n2422 gnd.n2421 585
R10942 gnd.n2421 gnd.n1040 585
R10943 gnd.n2413 gnd.n1038 585
R10944 gnd.n4733 gnd.n1038 585
R10945 gnd.n2417 gnd.n2416 585
R10946 gnd.n2416 gnd.n1029 585
R10947 gnd.n2415 gnd.n1027 585
R10948 gnd.n4739 gnd.n1027 585
R10949 gnd.n1014 gnd.n1012 585
R10950 gnd.n1017 gnd.n1014 585
R10951 gnd.n4747 gnd.n4746 585
R10952 gnd.n4746 gnd.n4745 585
R10953 gnd.n1013 gnd.n1010 585
R10954 gnd.n1015 gnd.n1013 585
R10955 gnd.n4751 gnd.n1009 585
R10956 gnd.n2535 gnd.n1009 585
R10957 gnd.n4753 gnd.n4752 585
R10958 gnd.n4753 gnd.n961 585
R10959 gnd.n7460 gnd.n7459 585
R10960 gnd.n7461 gnd.n7460 585
R10961 gnd.n110 gnd.n108 585
R10962 gnd.n108 gnd.n104 585
R10963 gnd.n7380 gnd.n7379 585
R10964 gnd.n7381 gnd.n7380 585
R10965 gnd.n189 gnd.n188 585
R10966 gnd.n188 gnd.n185 585
R10967 gnd.n7375 gnd.n7374 585
R10968 gnd.n7374 gnd.n7373 585
R10969 gnd.n192 gnd.n191 585
R10970 gnd.n193 gnd.n192 585
R10971 gnd.n7289 gnd.n7288 585
R10972 gnd.n7290 gnd.n7289 585
R10973 gnd.n204 gnd.n203 585
R10974 gnd.n211 gnd.n203 585
R10975 gnd.n7284 gnd.n7283 585
R10976 gnd.n7283 gnd.n7282 585
R10977 gnd.n207 gnd.n206 585
R10978 gnd.n208 gnd.n207 585
R10979 gnd.n7273 gnd.n7272 585
R10980 gnd.n7274 gnd.n7273 585
R10981 gnd.n221 gnd.n220 585
R10982 gnd.n220 gnd.n218 585
R10983 gnd.n7268 gnd.n7267 585
R10984 gnd.n7267 gnd.n7266 585
R10985 gnd.n224 gnd.n223 585
R10986 gnd.n225 gnd.n224 585
R10987 gnd.n7257 gnd.n7256 585
R10988 gnd.n7258 gnd.n7257 585
R10989 gnd.n234 gnd.n233 585
R10990 gnd.n241 gnd.n233 585
R10991 gnd.n7252 gnd.n7251 585
R10992 gnd.n7251 gnd.n7250 585
R10993 gnd.n237 gnd.n236 585
R10994 gnd.n238 gnd.n237 585
R10995 gnd.n7241 gnd.n7240 585
R10996 gnd.n7242 gnd.n7241 585
R10997 gnd.n252 gnd.n251 585
R10998 gnd.n251 gnd.n248 585
R10999 gnd.n7236 gnd.n7235 585
R11000 gnd.n7235 gnd.n7234 585
R11001 gnd.n255 gnd.n254 585
R11002 gnd.n7187 gnd.n255 585
R11003 gnd.n7225 gnd.n7224 585
R11004 gnd.n7226 gnd.n7225 585
R11005 gnd.n267 gnd.n266 585
R11006 gnd.n7192 gnd.n266 585
R11007 gnd.n7202 gnd.n7201 585
R11008 gnd.n7203 gnd.n7202 585
R11009 gnd.n7200 gnd.n7199 585
R11010 gnd.n7199 gnd.n7198 585
R11011 gnd.n7129 gnd.n297 585
R11012 gnd.n320 gnd.n297 585
R11013 gnd.n7131 gnd.n7130 585
R11014 gnd.n7132 gnd.n7131 585
R11015 gnd.n7128 gnd.n306 585
R11016 gnd.n7128 gnd.n7127 585
R11017 gnd.n305 gnd.n273 585
R11018 gnd.n314 gnd.n305 585
R11019 gnd.n277 gnd.n274 585
R11020 gnd.n7119 gnd.n277 585
R11021 gnd.n7221 gnd.n7220 585
R11022 gnd.n7220 gnd.n7219 585
R11023 gnd.n276 gnd.n275 585
R11024 gnd.n4276 gnd.n276 585
R11025 gnd.n4313 gnd.n4312 585
R11026 gnd.n4314 gnd.n4313 585
R11027 gnd.n1531 gnd.n1530 585
R11028 gnd.n1538 gnd.n1530 585
R11029 gnd.n4308 gnd.n4307 585
R11030 gnd.n4307 gnd.n4306 585
R11031 gnd.n1534 gnd.n1533 585
R11032 gnd.n4288 gnd.n1534 585
R11033 gnd.n4250 gnd.n1565 585
R11034 gnd.n1565 gnd.n1546 585
R11035 gnd.n4252 gnd.n4251 585
R11036 gnd.n4253 gnd.n4252 585
R11037 gnd.n1566 gnd.n1564 585
R11038 gnd.n1573 gnd.n1564 585
R11039 gnd.n4245 gnd.n4244 585
R11040 gnd.n4244 gnd.n4243 585
R11041 gnd.n1569 gnd.n1568 585
R11042 gnd.n4230 gnd.n1569 585
R11043 gnd.n4213 gnd.n1592 585
R11044 gnd.n1592 gnd.n1580 585
R11045 gnd.n4215 gnd.n4214 585
R11046 gnd.n4216 gnd.n4215 585
R11047 gnd.n1593 gnd.n1591 585
R11048 gnd.n1601 gnd.n1591 585
R11049 gnd.n4208 gnd.n4207 585
R11050 gnd.n4207 gnd.n4206 585
R11051 gnd.n1596 gnd.n1595 585
R11052 gnd.n4194 gnd.n1596 585
R11053 gnd.n4182 gnd.n1620 585
R11054 gnd.n1671 gnd.n1620 585
R11055 gnd.n4184 gnd.n4183 585
R11056 gnd.n4185 gnd.n4184 585
R11057 gnd.n1621 gnd.n1619 585
R11058 gnd.n1628 gnd.n1619 585
R11059 gnd.n4177 gnd.n4176 585
R11060 gnd.n4176 gnd.n4175 585
R11061 gnd.n1624 gnd.n1623 585
R11062 gnd.n4163 gnd.n1624 585
R11063 gnd.n1646 gnd.n1645 585
R11064 gnd.n1647 gnd.n1646 585
R11065 gnd.n1642 gnd.n1449 585
R11066 gnd.n4349 gnd.n1449 585
R11067 gnd.n4423 gnd.n4422 585
R11068 gnd.n4421 gnd.n1448 585
R11069 gnd.n4420 gnd.n1447 585
R11070 gnd.n4425 gnd.n1447 585
R11071 gnd.n4419 gnd.n4418 585
R11072 gnd.n4417 gnd.n4416 585
R11073 gnd.n4415 gnd.n4414 585
R11074 gnd.n4413 gnd.n4412 585
R11075 gnd.n4411 gnd.n4410 585
R11076 gnd.n4409 gnd.n4408 585
R11077 gnd.n4407 gnd.n4406 585
R11078 gnd.n4405 gnd.n4404 585
R11079 gnd.n4403 gnd.n4402 585
R11080 gnd.n4401 gnd.n4400 585
R11081 gnd.n4399 gnd.n4398 585
R11082 gnd.n4397 gnd.n4396 585
R11083 gnd.n4395 gnd.n4394 585
R11084 gnd.n4392 gnd.n4391 585
R11085 gnd.n4390 gnd.n4389 585
R11086 gnd.n4388 gnd.n4387 585
R11087 gnd.n4386 gnd.n4385 585
R11088 gnd.n4384 gnd.n4383 585
R11089 gnd.n4382 gnd.n4381 585
R11090 gnd.n4380 gnd.n4379 585
R11091 gnd.n4378 gnd.n4377 585
R11092 gnd.n4376 gnd.n4375 585
R11093 gnd.n4374 gnd.n4373 585
R11094 gnd.n4372 gnd.n4371 585
R11095 gnd.n4370 gnd.n4369 585
R11096 gnd.n4368 gnd.n4367 585
R11097 gnd.n4366 gnd.n4365 585
R11098 gnd.n4364 gnd.n4363 585
R11099 gnd.n4362 gnd.n4361 585
R11100 gnd.n4360 gnd.n4359 585
R11101 gnd.n4358 gnd.n4357 585
R11102 gnd.n4356 gnd.n1489 585
R11103 gnd.n1493 gnd.n1490 585
R11104 gnd.n4352 gnd.n4351 585
R11105 gnd.n178 gnd.n177 585
R11106 gnd.n7389 gnd.n173 585
R11107 gnd.n7391 gnd.n7390 585
R11108 gnd.n7393 gnd.n171 585
R11109 gnd.n7395 gnd.n7394 585
R11110 gnd.n7396 gnd.n166 585
R11111 gnd.n7398 gnd.n7397 585
R11112 gnd.n7400 gnd.n164 585
R11113 gnd.n7402 gnd.n7401 585
R11114 gnd.n7403 gnd.n159 585
R11115 gnd.n7405 gnd.n7404 585
R11116 gnd.n7407 gnd.n157 585
R11117 gnd.n7409 gnd.n7408 585
R11118 gnd.n7410 gnd.n152 585
R11119 gnd.n7412 gnd.n7411 585
R11120 gnd.n7414 gnd.n150 585
R11121 gnd.n7416 gnd.n7415 585
R11122 gnd.n7417 gnd.n145 585
R11123 gnd.n7419 gnd.n7418 585
R11124 gnd.n7421 gnd.n143 585
R11125 gnd.n7423 gnd.n7422 585
R11126 gnd.n7427 gnd.n138 585
R11127 gnd.n7429 gnd.n7428 585
R11128 gnd.n7431 gnd.n136 585
R11129 gnd.n7433 gnd.n7432 585
R11130 gnd.n7434 gnd.n131 585
R11131 gnd.n7436 gnd.n7435 585
R11132 gnd.n7438 gnd.n129 585
R11133 gnd.n7440 gnd.n7439 585
R11134 gnd.n7441 gnd.n124 585
R11135 gnd.n7443 gnd.n7442 585
R11136 gnd.n7445 gnd.n122 585
R11137 gnd.n7447 gnd.n7446 585
R11138 gnd.n7448 gnd.n117 585
R11139 gnd.n7450 gnd.n7449 585
R11140 gnd.n7452 gnd.n115 585
R11141 gnd.n7454 gnd.n7453 585
R11142 gnd.n7455 gnd.n113 585
R11143 gnd.n7456 gnd.n109 585
R11144 gnd.n109 gnd.n106 585
R11145 gnd.n7385 gnd.n105 585
R11146 gnd.n7461 gnd.n105 585
R11147 gnd.n7384 gnd.n7383 585
R11148 gnd.n7383 gnd.n104 585
R11149 gnd.n7382 gnd.n182 585
R11150 gnd.n7382 gnd.n7381 585
R11151 gnd.n7161 gnd.n183 585
R11152 gnd.n185 gnd.n183 585
R11153 gnd.n7162 gnd.n194 585
R11154 gnd.n7373 gnd.n194 585
R11155 gnd.n7164 gnd.n7163 585
R11156 gnd.n7163 gnd.n193 585
R11157 gnd.n7165 gnd.n202 585
R11158 gnd.n7290 gnd.n202 585
R11159 gnd.n7167 gnd.n7166 585
R11160 gnd.n7166 gnd.n211 585
R11161 gnd.n7168 gnd.n209 585
R11162 gnd.n7282 gnd.n209 585
R11163 gnd.n7170 gnd.n7169 585
R11164 gnd.n7169 gnd.n208 585
R11165 gnd.n7171 gnd.n219 585
R11166 gnd.n7274 gnd.n219 585
R11167 gnd.n7173 gnd.n7172 585
R11168 gnd.n7172 gnd.n218 585
R11169 gnd.n7174 gnd.n226 585
R11170 gnd.n7266 gnd.n226 585
R11171 gnd.n7176 gnd.n7175 585
R11172 gnd.n7175 gnd.n225 585
R11173 gnd.n7177 gnd.n232 585
R11174 gnd.n7258 gnd.n232 585
R11175 gnd.n7179 gnd.n7178 585
R11176 gnd.n7178 gnd.n241 585
R11177 gnd.n7180 gnd.n239 585
R11178 gnd.n7250 gnd.n239 585
R11179 gnd.n7182 gnd.n7181 585
R11180 gnd.n7181 gnd.n238 585
R11181 gnd.n7183 gnd.n249 585
R11182 gnd.n7242 gnd.n249 585
R11183 gnd.n7185 gnd.n7184 585
R11184 gnd.n7184 gnd.n248 585
R11185 gnd.n7186 gnd.n257 585
R11186 gnd.n7234 gnd.n257 585
R11187 gnd.n7189 gnd.n7188 585
R11188 gnd.n7188 gnd.n7187 585
R11189 gnd.n7190 gnd.n264 585
R11190 gnd.n7226 gnd.n264 585
R11191 gnd.n7194 gnd.n7193 585
R11192 gnd.n7193 gnd.n7192 585
R11193 gnd.n7195 gnd.n295 585
R11194 gnd.n7203 gnd.n295 585
R11195 gnd.n7197 gnd.n7196 585
R11196 gnd.n7198 gnd.n7197 585
R11197 gnd.n7135 gnd.n298 585
R11198 gnd.n320 gnd.n298 585
R11199 gnd.n7134 gnd.n7133 585
R11200 gnd.n7133 gnd.n7132 585
R11201 gnd.n301 gnd.n299 585
R11202 gnd.n7127 gnd.n301 585
R11203 gnd.n4271 gnd.n4270 585
R11204 gnd.n4270 gnd.n314 585
R11205 gnd.n4272 gnd.n313 585
R11206 gnd.n7119 gnd.n313 585
R11207 gnd.n4273 gnd.n279 585
R11208 gnd.n7219 gnd.n279 585
R11209 gnd.n4275 gnd.n4274 585
R11210 gnd.n4276 gnd.n4275 585
R11211 gnd.n1554 gnd.n1527 585
R11212 gnd.n4314 gnd.n1527 585
R11213 gnd.n4262 gnd.n4261 585
R11214 gnd.n4261 gnd.n1538 585
R11215 gnd.n4260 gnd.n1536 585
R11216 gnd.n4306 gnd.n1536 585
R11217 gnd.n4259 gnd.n1547 585
R11218 gnd.n4288 gnd.n1547 585
R11219 gnd.n1560 gnd.n1556 585
R11220 gnd.n1560 gnd.n1546 585
R11221 gnd.n4255 gnd.n4254 585
R11222 gnd.n4254 gnd.n4253 585
R11223 gnd.n1559 gnd.n1558 585
R11224 gnd.n1573 gnd.n1559 585
R11225 gnd.n1662 gnd.n1571 585
R11226 gnd.n4243 gnd.n1571 585
R11227 gnd.n1663 gnd.n1581 585
R11228 gnd.n4230 gnd.n1581 585
R11229 gnd.n1665 gnd.n1664 585
R11230 gnd.n1664 gnd.n1580 585
R11231 gnd.n1666 gnd.n1589 585
R11232 gnd.n4216 gnd.n1589 585
R11233 gnd.n1668 gnd.n1667 585
R11234 gnd.n1667 gnd.n1601 585
R11235 gnd.n1669 gnd.n1598 585
R11236 gnd.n4206 gnd.n1598 585
R11237 gnd.n1670 gnd.n1608 585
R11238 gnd.n4194 gnd.n1608 585
R11239 gnd.n1673 gnd.n1672 585
R11240 gnd.n1672 gnd.n1671 585
R11241 gnd.n1674 gnd.n1616 585
R11242 gnd.n4185 gnd.n1616 585
R11243 gnd.n1676 gnd.n1675 585
R11244 gnd.n1675 gnd.n1628 585
R11245 gnd.n1677 gnd.n1626 585
R11246 gnd.n4175 gnd.n1626 585
R11247 gnd.n1679 gnd.n1678 585
R11248 gnd.n4163 gnd.n1679 585
R11249 gnd.n1648 gnd.n1495 585
R11250 gnd.n1647 gnd.n1495 585
R11251 gnd.n4350 gnd.n1496 585
R11252 gnd.n4350 gnd.n4349 585
R11253 gnd.n3378 gnd.n3175 585
R11254 gnd.n3256 gnd.n3175 585
R11255 gnd.n3380 gnd.n3379 585
R11256 gnd.n3380 gnd.n1897 585
R11257 gnd.n3381 gnd.n3174 585
R11258 gnd.n3381 gnd.n1896 585
R11259 gnd.n3383 gnd.n3382 585
R11260 gnd.n3382 gnd.t131 585
R11261 gnd.n3384 gnd.n3169 585
R11262 gnd.n3169 gnd.n1903 585
R11263 gnd.n3386 gnd.n3385 585
R11264 gnd.n3387 gnd.n3386 585
R11265 gnd.n3173 gnd.n3168 585
R11266 gnd.n3168 gnd.n1912 585
R11267 gnd.n3172 gnd.n3171 585
R11268 gnd.n3171 gnd.n1911 585
R11269 gnd.n3170 gnd.n3160 585
R11270 gnd.n3394 gnd.n3160 585
R11271 gnd.n3397 gnd.n3159 585
R11272 gnd.n3397 gnd.n3396 585
R11273 gnd.n3399 gnd.n3398 585
R11274 gnd.n3398 gnd.n1918 585
R11275 gnd.n3400 gnd.n3157 585
R11276 gnd.n3157 gnd.n3156 585
R11277 gnd.n3402 gnd.n3401 585
R11278 gnd.n3403 gnd.n3402 585
R11279 gnd.n3158 gnd.n3155 585
R11280 gnd.n3155 gnd.n1925 585
R11281 gnd.n3147 gnd.n3146 585
R11282 gnd.n3409 gnd.n3147 585
R11283 gnd.n3413 gnd.n3412 585
R11284 gnd.n3412 gnd.n3411 585
R11285 gnd.n3414 gnd.n3143 585
R11286 gnd.n3143 gnd.n1931 585
R11287 gnd.n3416 gnd.n3415 585
R11288 gnd.n3417 gnd.n3416 585
R11289 gnd.n3145 gnd.n3142 585
R11290 gnd.n3142 gnd.n1939 585
R11291 gnd.n3144 gnd.n3134 585
R11292 gnd.n3134 gnd.n1938 585
R11293 gnd.n3425 gnd.n3133 585
R11294 gnd.n3425 gnd.n3424 585
R11295 gnd.n3427 gnd.n3426 585
R11296 gnd.n3426 gnd.n1947 585
R11297 gnd.n3428 gnd.n3132 585
R11298 gnd.n3132 gnd.n1945 585
R11299 gnd.n3430 gnd.n3429 585
R11300 gnd.n3431 gnd.n3430 585
R11301 gnd.n3126 gnd.n3125 585
R11302 gnd.n3126 gnd.n1953 585
R11303 gnd.n3439 gnd.n3438 585
R11304 gnd.n3438 gnd.n3437 585
R11305 gnd.n3440 gnd.n3123 585
R11306 gnd.n3127 gnd.n3123 585
R11307 gnd.n3442 gnd.n3441 585
R11308 gnd.n3443 gnd.n3442 585
R11309 gnd.n3124 gnd.n3115 585
R11310 gnd.n3115 gnd.n1959 585
R11311 gnd.n3451 gnd.n3114 585
R11312 gnd.n3451 gnd.n3450 585
R11313 gnd.n3453 gnd.n3452 585
R11314 gnd.n3452 gnd.n1967 585
R11315 gnd.n3454 gnd.n3111 585
R11316 gnd.n3111 gnd.n1966 585
R11317 gnd.n3456 gnd.n3455 585
R11318 gnd.n3457 gnd.n3456 585
R11319 gnd.n3113 gnd.n3110 585
R11320 gnd.n3110 gnd.n1975 585
R11321 gnd.n3112 gnd.n3102 585
R11322 gnd.n3102 gnd.n1973 585
R11323 gnd.n3466 gnd.n3101 585
R11324 gnd.n3466 gnd.n3465 585
R11325 gnd.n3468 gnd.n3467 585
R11326 gnd.n3467 gnd.n1981 585
R11327 gnd.n3469 gnd.n3098 585
R11328 gnd.n3098 gnd.n3097 585
R11329 gnd.n3471 gnd.n3470 585
R11330 gnd.n3472 gnd.n3471 585
R11331 gnd.n3100 gnd.n3096 585
R11332 gnd.n3096 gnd.n1989 585
R11333 gnd.n3099 gnd.n3089 585
R11334 gnd.n3089 gnd.n1987 585
R11335 gnd.n3481 gnd.n3088 585
R11336 gnd.n3481 gnd.n3480 585
R11337 gnd.n3483 gnd.n3482 585
R11338 gnd.n3482 gnd.n1995 585
R11339 gnd.n3484 gnd.n3085 585
R11340 gnd.n3085 gnd.n3084 585
R11341 gnd.n3486 gnd.n3485 585
R11342 gnd.n3487 gnd.n3486 585
R11343 gnd.n3087 gnd.n3083 585
R11344 gnd.n3083 gnd.n2002 585
R11345 gnd.n3086 gnd.n3061 585
R11346 gnd.n3493 gnd.n3061 585
R11347 gnd.n3496 gnd.n3062 585
R11348 gnd.n3496 gnd.n3495 585
R11349 gnd.n3497 gnd.n3060 585
R11350 gnd.n3497 gnd.n2009 585
R11351 gnd.n3499 gnd.n3498 585
R11352 gnd.n3498 gnd.n2008 585
R11353 gnd.n3500 gnd.n3059 585
R11354 gnd.n3074 gnd.n3059 585
R11355 gnd.n3502 gnd.n3501 585
R11356 gnd.n3502 gnd.n2017 585
R11357 gnd.n3503 gnd.n3058 585
R11358 gnd.n3503 gnd.n2015 585
R11359 gnd.n3505 gnd.n3504 585
R11360 gnd.n3504 gnd.n2025 585
R11361 gnd.n3506 gnd.n3056 585
R11362 gnd.n3056 gnd.n2023 585
R11363 gnd.n3508 gnd.n3507 585
R11364 gnd.n3509 gnd.n3508 585
R11365 gnd.n3057 gnd.n3055 585
R11366 gnd.n3055 gnd.n2032 585
R11367 gnd.n3041 gnd.n3040 585
R11368 gnd.n3515 gnd.n3041 585
R11369 gnd.n3518 gnd.n3517 585
R11370 gnd.n3517 gnd.n3516 585
R11371 gnd.n3519 gnd.n3039 585
R11372 gnd.n3039 gnd.n2038 585
R11373 gnd.n3521 gnd.n3520 585
R11374 gnd.n3522 gnd.n3521 585
R11375 gnd.n3035 gnd.n3034 585
R11376 gnd.n3523 gnd.n3035 585
R11377 gnd.n3527 gnd.n3526 585
R11378 gnd.n3526 gnd.n3525 585
R11379 gnd.n3528 gnd.n3031 585
R11380 gnd.n3031 gnd.n2044 585
R11381 gnd.n3530 gnd.n3529 585
R11382 gnd.n3531 gnd.n3530 585
R11383 gnd.n3033 gnd.n3030 585
R11384 gnd.n3030 gnd.n2052 585
R11385 gnd.n3032 gnd.n3021 585
R11386 gnd.n3021 gnd.n2051 585
R11387 gnd.n3539 gnd.n3020 585
R11388 gnd.n3539 gnd.n3538 585
R11389 gnd.n3541 gnd.n3540 585
R11390 gnd.n3540 gnd.n2060 585
R11391 gnd.n3542 gnd.n3017 585
R11392 gnd.n3017 gnd.n2058 585
R11393 gnd.n3544 gnd.n3543 585
R11394 gnd.n3545 gnd.n3544 585
R11395 gnd.n3019 gnd.n3016 585
R11396 gnd.n3016 gnd.n2067 585
R11397 gnd.n3018 gnd.n3008 585
R11398 gnd.n3008 gnd.n2066 585
R11399 gnd.n3553 gnd.n3007 585
R11400 gnd.n3553 gnd.n3552 585
R11401 gnd.n3555 gnd.n3554 585
R11402 gnd.n3554 gnd.n2075 585
R11403 gnd.n3556 gnd.n3006 585
R11404 gnd.n3006 gnd.n2073 585
R11405 gnd.n3558 gnd.n3557 585
R11406 gnd.n3559 gnd.n3558 585
R11407 gnd.n2998 gnd.n2997 585
R11408 gnd.n3004 gnd.n2998 585
R11409 gnd.n3567 gnd.n3566 585
R11410 gnd.n3566 gnd.n3565 585
R11411 gnd.n3568 gnd.n2894 585
R11412 gnd.n2894 gnd.n2892 585
R11413 gnd.n3570 gnd.n3569 585
R11414 gnd.n3571 gnd.n3570 585
R11415 gnd.n2995 gnd.n2893 585
R11416 gnd.n2994 gnd.n2993 585
R11417 gnd.n2991 gnd.n2915 585
R11418 gnd.n2991 gnd.n2086 585
R11419 gnd.n2990 gnd.n2989 585
R11420 gnd.n2988 gnd.n2987 585
R11421 gnd.n2986 gnd.n2917 585
R11422 gnd.n2984 gnd.n2983 585
R11423 gnd.n2982 gnd.n2918 585
R11424 gnd.n2981 gnd.n2980 585
R11425 gnd.n2978 gnd.n2919 585
R11426 gnd.n2976 gnd.n2975 585
R11427 gnd.n2974 gnd.n2920 585
R11428 gnd.n2973 gnd.n2972 585
R11429 gnd.n2970 gnd.n2921 585
R11430 gnd.n2968 gnd.n2967 585
R11431 gnd.n2966 gnd.n2922 585
R11432 gnd.n2965 gnd.n2964 585
R11433 gnd.n2962 gnd.n2923 585
R11434 gnd.n2960 gnd.n2959 585
R11435 gnd.n2958 gnd.n2924 585
R11436 gnd.n2957 gnd.n2956 585
R11437 gnd.n2954 gnd.n2925 585
R11438 gnd.n2952 gnd.n2951 585
R11439 gnd.n2950 gnd.n2926 585
R11440 gnd.n2949 gnd.n2948 585
R11441 gnd.n2946 gnd.n2927 585
R11442 gnd.n2944 gnd.n2943 585
R11443 gnd.n2942 gnd.n2928 585
R11444 gnd.n2941 gnd.n2940 585
R11445 gnd.n2938 gnd.n2937 585
R11446 gnd.n2936 gnd.n2935 585
R11447 gnd.n2934 gnd.n2871 585
R11448 gnd.n3640 gnd.n3639 585
R11449 gnd.n3637 gnd.n2870 585
R11450 gnd.n3635 gnd.n3634 585
R11451 gnd.n3633 gnd.n2873 585
R11452 gnd.n3631 gnd.n3630 585
R11453 gnd.n3628 gnd.n2876 585
R11454 gnd.n3626 gnd.n3625 585
R11455 gnd.n3624 gnd.n2877 585
R11456 gnd.n3623 gnd.n3622 585
R11457 gnd.n3620 gnd.n2878 585
R11458 gnd.n3618 gnd.n3617 585
R11459 gnd.n3616 gnd.n2879 585
R11460 gnd.n3615 gnd.n3614 585
R11461 gnd.n3612 gnd.n2880 585
R11462 gnd.n3610 gnd.n3609 585
R11463 gnd.n3608 gnd.n2881 585
R11464 gnd.n3607 gnd.n3606 585
R11465 gnd.n3604 gnd.n2882 585
R11466 gnd.n3602 gnd.n3601 585
R11467 gnd.n3600 gnd.n2883 585
R11468 gnd.n3599 gnd.n3598 585
R11469 gnd.n3596 gnd.n2884 585
R11470 gnd.n3594 gnd.n3593 585
R11471 gnd.n3592 gnd.n2885 585
R11472 gnd.n3591 gnd.n3590 585
R11473 gnd.n3588 gnd.n2886 585
R11474 gnd.n3586 gnd.n3585 585
R11475 gnd.n3584 gnd.n2887 585
R11476 gnd.n3583 gnd.n3582 585
R11477 gnd.n3580 gnd.n2888 585
R11478 gnd.n3578 gnd.n3577 585
R11479 gnd.n3576 gnd.n2889 585
R11480 gnd.n3575 gnd.n3574 585
R11481 gnd.n3259 gnd.n3258 585
R11482 gnd.n3260 gnd.n3245 585
R11483 gnd.n3262 gnd.n3261 585
R11484 gnd.n3264 gnd.n3243 585
R11485 gnd.n3266 gnd.n3265 585
R11486 gnd.n3267 gnd.n3242 585
R11487 gnd.n3269 gnd.n3268 585
R11488 gnd.n3271 gnd.n3240 585
R11489 gnd.n3273 gnd.n3272 585
R11490 gnd.n3274 gnd.n3239 585
R11491 gnd.n3276 gnd.n3275 585
R11492 gnd.n3278 gnd.n3237 585
R11493 gnd.n3280 gnd.n3279 585
R11494 gnd.n3281 gnd.n3236 585
R11495 gnd.n3283 gnd.n3282 585
R11496 gnd.n3285 gnd.n3234 585
R11497 gnd.n3287 gnd.n3286 585
R11498 gnd.n3288 gnd.n3233 585
R11499 gnd.n3290 gnd.n3289 585
R11500 gnd.n3292 gnd.n3231 585
R11501 gnd.n3294 gnd.n3293 585
R11502 gnd.n3295 gnd.n3230 585
R11503 gnd.n3297 gnd.n3296 585
R11504 gnd.n3299 gnd.n3228 585
R11505 gnd.n3301 gnd.n3300 585
R11506 gnd.n3302 gnd.n3227 585
R11507 gnd.n3304 gnd.n3303 585
R11508 gnd.n3306 gnd.n3225 585
R11509 gnd.n3308 gnd.n3307 585
R11510 gnd.n3310 gnd.n3222 585
R11511 gnd.n3312 gnd.n3311 585
R11512 gnd.n3314 gnd.n3221 585
R11513 gnd.n3315 gnd.n3196 585
R11514 gnd.n3318 gnd.n1466 585
R11515 gnd.n3320 gnd.n3319 585
R11516 gnd.n3322 gnd.n3219 585
R11517 gnd.n3324 gnd.n3323 585
R11518 gnd.n3326 gnd.n3216 585
R11519 gnd.n3328 gnd.n3327 585
R11520 gnd.n3330 gnd.n3214 585
R11521 gnd.n3332 gnd.n3331 585
R11522 gnd.n3333 gnd.n3213 585
R11523 gnd.n3335 gnd.n3334 585
R11524 gnd.n3337 gnd.n3211 585
R11525 gnd.n3339 gnd.n3338 585
R11526 gnd.n3340 gnd.n3210 585
R11527 gnd.n3342 gnd.n3341 585
R11528 gnd.n3344 gnd.n3208 585
R11529 gnd.n3346 gnd.n3345 585
R11530 gnd.n3347 gnd.n3207 585
R11531 gnd.n3349 gnd.n3348 585
R11532 gnd.n3351 gnd.n3205 585
R11533 gnd.n3353 gnd.n3352 585
R11534 gnd.n3354 gnd.n3204 585
R11535 gnd.n3356 gnd.n3355 585
R11536 gnd.n3358 gnd.n3202 585
R11537 gnd.n3360 gnd.n3359 585
R11538 gnd.n3361 gnd.n3201 585
R11539 gnd.n3363 gnd.n3362 585
R11540 gnd.n3365 gnd.n3199 585
R11541 gnd.n3367 gnd.n3366 585
R11542 gnd.n3368 gnd.n3198 585
R11543 gnd.n3370 gnd.n3369 585
R11544 gnd.n3372 gnd.n3197 585
R11545 gnd.n3373 gnd.n3195 585
R11546 gnd.n3376 gnd.n3375 585
R11547 gnd.n3257 gnd.n3246 585
R11548 gnd.n3257 gnd.n3256 585
R11549 gnd.n3254 gnd.n3253 585
R11550 gnd.n3254 gnd.n1897 585
R11551 gnd.n3252 gnd.n3248 585
R11552 gnd.n3248 gnd.n1896 585
R11553 gnd.n3251 gnd.n3250 585
R11554 gnd.n3250 gnd.t131 585
R11555 gnd.n3249 gnd.n3167 585
R11556 gnd.n3167 gnd.n1903 585
R11557 gnd.n3388 gnd.n3166 585
R11558 gnd.n3388 gnd.n3387 585
R11559 gnd.n3390 gnd.n3389 585
R11560 gnd.n3389 gnd.n1912 585
R11561 gnd.n3391 gnd.n3162 585
R11562 gnd.n3162 gnd.n1911 585
R11563 gnd.n3393 gnd.n3392 585
R11564 gnd.n3394 gnd.n3393 585
R11565 gnd.n3165 gnd.n3161 585
R11566 gnd.n3396 gnd.n3161 585
R11567 gnd.n3164 gnd.n3163 585
R11568 gnd.n3163 gnd.n1918 585
R11569 gnd.n3153 gnd.n3152 585
R11570 gnd.n3156 gnd.n3153 585
R11571 gnd.n3405 gnd.n3404 585
R11572 gnd.n3404 gnd.n3403 585
R11573 gnd.n3406 gnd.n3149 585
R11574 gnd.n3149 gnd.n1925 585
R11575 gnd.n3408 gnd.n3407 585
R11576 gnd.n3409 gnd.n3408 585
R11577 gnd.n3151 gnd.n3148 585
R11578 gnd.n3411 gnd.n3148 585
R11579 gnd.n3150 gnd.n3140 585
R11580 gnd.n3140 gnd.n1931 585
R11581 gnd.n3418 gnd.n3139 585
R11582 gnd.n3418 gnd.n3417 585
R11583 gnd.n3420 gnd.n3419 585
R11584 gnd.n3419 gnd.n1939 585
R11585 gnd.n3421 gnd.n3137 585
R11586 gnd.n3137 gnd.n1938 585
R11587 gnd.n3423 gnd.n3422 585
R11588 gnd.n3424 gnd.n3423 585
R11589 gnd.n3138 gnd.n3136 585
R11590 gnd.n3136 gnd.n1947 585
R11591 gnd.n3130 gnd.n3129 585
R11592 gnd.n3130 gnd.n1945 585
R11593 gnd.n3433 gnd.n3432 585
R11594 gnd.n3432 gnd.n3431 585
R11595 gnd.n3434 gnd.n3128 585
R11596 gnd.n3128 gnd.n1953 585
R11597 gnd.n3436 gnd.n3435 585
R11598 gnd.n3437 gnd.n3436 585
R11599 gnd.n3121 gnd.n3120 585
R11600 gnd.n3127 gnd.n3121 585
R11601 gnd.n3445 gnd.n3444 585
R11602 gnd.n3444 gnd.n3443 585
R11603 gnd.n3446 gnd.n3117 585
R11604 gnd.n3117 gnd.n1959 585
R11605 gnd.n3448 gnd.n3447 585
R11606 gnd.n3450 gnd.n3448 585
R11607 gnd.n3119 gnd.n3116 585
R11608 gnd.n3116 gnd.n1967 585
R11609 gnd.n3118 gnd.n3108 585
R11610 gnd.n3108 gnd.n1966 585
R11611 gnd.n3458 gnd.n3107 585
R11612 gnd.n3458 gnd.n3457 585
R11613 gnd.n3460 gnd.n3459 585
R11614 gnd.n3459 gnd.n1975 585
R11615 gnd.n3461 gnd.n3104 585
R11616 gnd.n3104 gnd.n1973 585
R11617 gnd.n3463 gnd.n3462 585
R11618 gnd.n3465 gnd.n3463 585
R11619 gnd.n3106 gnd.n3103 585
R11620 gnd.n3103 gnd.n1981 585
R11621 gnd.n3105 gnd.n3094 585
R11622 gnd.n3097 gnd.n3094 585
R11623 gnd.n3473 gnd.n3093 585
R11624 gnd.n3473 gnd.n3472 585
R11625 gnd.n3475 gnd.n3474 585
R11626 gnd.n3474 gnd.n1989 585
R11627 gnd.n3476 gnd.n3091 585
R11628 gnd.n3091 gnd.n1987 585
R11629 gnd.n3478 gnd.n3477 585
R11630 gnd.n3480 gnd.n3478 585
R11631 gnd.n3092 gnd.n3090 585
R11632 gnd.n3090 gnd.n1995 585
R11633 gnd.n3081 gnd.n3080 585
R11634 gnd.n3084 gnd.n3081 585
R11635 gnd.n3489 gnd.n3488 585
R11636 gnd.n3488 gnd.n3487 585
R11637 gnd.n3490 gnd.n3064 585
R11638 gnd.n3064 gnd.n2002 585
R11639 gnd.n3492 gnd.n3491 585
R11640 gnd.n3493 gnd.n3492 585
R11641 gnd.n3079 gnd.n3063 585
R11642 gnd.n3495 gnd.n3063 585
R11643 gnd.n3078 gnd.n3077 585
R11644 gnd.n3077 gnd.n2009 585
R11645 gnd.n3076 gnd.n3065 585
R11646 gnd.n3076 gnd.n2008 585
R11647 gnd.n3075 gnd.n3072 585
R11648 gnd.n3075 gnd.n3074 585
R11649 gnd.n3071 gnd.n3066 585
R11650 gnd.n3066 gnd.n2017 585
R11651 gnd.n3070 gnd.n3069 585
R11652 gnd.n3069 gnd.n2015 585
R11653 gnd.n3068 gnd.n3067 585
R11654 gnd.n3068 gnd.n2025 585
R11655 gnd.n3053 gnd.n3052 585
R11656 gnd.n3053 gnd.n2023 585
R11657 gnd.n3511 gnd.n3510 585
R11658 gnd.n3510 gnd.n3509 585
R11659 gnd.n3512 gnd.n3044 585
R11660 gnd.n3044 gnd.n2032 585
R11661 gnd.n3514 gnd.n3513 585
R11662 gnd.n3515 gnd.n3514 585
R11663 gnd.n3051 gnd.n3043 585
R11664 gnd.n3516 gnd.n3043 585
R11665 gnd.n3050 gnd.n3049 585
R11666 gnd.n3049 gnd.n2038 585
R11667 gnd.n3048 gnd.n3038 585
R11668 gnd.n3522 gnd.n3038 585
R11669 gnd.n3047 gnd.n3037 585
R11670 gnd.n3523 gnd.n3037 585
R11671 gnd.n3046 gnd.n3036 585
R11672 gnd.n3525 gnd.n3036 585
R11673 gnd.n3045 gnd.n3028 585
R11674 gnd.n3028 gnd.n2044 585
R11675 gnd.n3532 gnd.n3027 585
R11676 gnd.n3532 gnd.n3531 585
R11677 gnd.n3534 gnd.n3533 585
R11678 gnd.n3533 gnd.n2052 585
R11679 gnd.n3535 gnd.n3024 585
R11680 gnd.n3024 gnd.n2051 585
R11681 gnd.n3537 gnd.n3536 585
R11682 gnd.n3538 gnd.n3537 585
R11683 gnd.n3026 gnd.n3023 585
R11684 gnd.n3023 gnd.n2060 585
R11685 gnd.n3025 gnd.n3014 585
R11686 gnd.n3014 gnd.n2058 585
R11687 gnd.n3546 gnd.n3013 585
R11688 gnd.n3546 gnd.n3545 585
R11689 gnd.n3548 gnd.n3547 585
R11690 gnd.n3547 gnd.n2067 585
R11691 gnd.n3549 gnd.n3011 585
R11692 gnd.n3011 gnd.n2066 585
R11693 gnd.n3551 gnd.n3550 585
R11694 gnd.n3552 gnd.n3551 585
R11695 gnd.n3012 gnd.n3010 585
R11696 gnd.n3010 gnd.n2075 585
R11697 gnd.n3003 gnd.n3002 585
R11698 gnd.n3003 gnd.n2073 585
R11699 gnd.n3561 gnd.n3560 585
R11700 gnd.n3560 gnd.n3559 585
R11701 gnd.n3562 gnd.n3000 585
R11702 gnd.n3004 gnd.n3000 585
R11703 gnd.n3564 gnd.n3563 585
R11704 gnd.n3565 gnd.n3564 585
R11705 gnd.n3001 gnd.n2891 585
R11706 gnd.n2892 gnd.n2891 585
R11707 gnd.n3572 gnd.n2890 585
R11708 gnd.n3572 gnd.n3571 585
R11709 gnd.n895 gnd.n894 585
R11710 gnd.n1097 gnd.n895 585
R11711 gnd.n7097 gnd.n7096 585
R11712 gnd.n7097 gnd.n250 585
R11713 gnd.n7099 gnd.n328 585
R11714 gnd.n7099 gnd.n7098 585
R11715 gnd.n7101 gnd.n7100 585
R11716 gnd.n7100 gnd.n256 585
R11717 gnd.n7102 gnd.n324 585
R11718 gnd.n324 gnd.n265 585
R11719 gnd.n7104 gnd.n7103 585
R11720 gnd.n7104 gnd.n263 585
R11721 gnd.n7105 gnd.n323 585
R11722 gnd.n7105 gnd.n296 585
R11723 gnd.n7107 gnd.n7106 585
R11724 gnd.n7106 gnd.n294 585
R11725 gnd.n7109 gnd.n322 585
R11726 gnd.n322 gnd.n321 585
R11727 gnd.n7111 gnd.n7110 585
R11728 gnd.n7111 gnd.n304 585
R11729 gnd.n7113 gnd.n7112 585
R11730 gnd.n7112 gnd.n302 585
R11731 gnd.n7114 gnd.n316 585
R11732 gnd.n316 gnd.n307 585
R11733 gnd.n7117 gnd.n7116 585
R11734 gnd.n7118 gnd.n7117 585
R11735 gnd.n317 gnd.n315 585
R11736 gnd.n315 gnd.n312 585
R11737 gnd.n4299 gnd.n4298 585
R11738 gnd.n4299 gnd.n278 585
R11739 gnd.n4301 gnd.n4300 585
R11740 gnd.n4300 gnd.n1529 585
R11741 gnd.n4302 gnd.n1541 585
R11742 gnd.n1541 gnd.n1540 585
R11743 gnd.n4304 gnd.n4303 585
R11744 gnd.n4305 gnd.n4304 585
R11745 gnd.n1542 gnd.n1539 585
R11746 gnd.n1539 gnd.n1535 585
R11747 gnd.n4291 gnd.n4290 585
R11748 gnd.n4290 gnd.n4289 585
R11749 gnd.n1545 gnd.n1544 585
R11750 gnd.n1563 gnd.n1545 585
R11751 gnd.n4238 gnd.n1575 585
R11752 gnd.n1575 gnd.n1561 585
R11753 gnd.n4240 gnd.n4239 585
R11754 gnd.n4241 gnd.n4240 585
R11755 gnd.n1576 gnd.n1574 585
R11756 gnd.n1574 gnd.n1570 585
R11757 gnd.n4233 gnd.n4232 585
R11758 gnd.n4232 gnd.n4231 585
R11759 gnd.n1579 gnd.n1578 585
R11760 gnd.n1590 gnd.n1579 585
R11761 gnd.n4202 gnd.n1603 585
R11762 gnd.n1603 gnd.n1588 585
R11763 gnd.n4204 gnd.n4203 585
R11764 gnd.n4205 gnd.n4204 585
R11765 gnd.n1604 gnd.n1602 585
R11766 gnd.n1602 gnd.n1597 585
R11767 gnd.n4197 gnd.n4196 585
R11768 gnd.n4196 gnd.n4195 585
R11769 gnd.n1607 gnd.n1606 585
R11770 gnd.n1617 gnd.n1607 585
R11771 gnd.n4171 gnd.n1630 585
R11772 gnd.n1630 gnd.n1615 585
R11773 gnd.n4173 gnd.n4172 585
R11774 gnd.n4174 gnd.n4173 585
R11775 gnd.n1631 gnd.n1629 585
R11776 gnd.n1629 gnd.n1625 585
R11777 gnd.n4166 gnd.n4165 585
R11778 gnd.n4165 gnd.n4164 585
R11779 gnd.n1641 gnd.n1633 585
R11780 gnd.n1641 gnd.n1499 585
R11781 gnd.n1640 gnd.n1639 585
R11782 gnd.n1640 gnd.n1497 585
R11783 gnd.n1635 gnd.n1634 585
R11784 gnd.n1634 gnd.n1446 585
R11785 gnd.n1416 gnd.n1415 585
R11786 gnd.n4426 gnd.n1416 585
R11787 gnd.n4429 gnd.n4428 585
R11788 gnd.n4428 gnd.n4427 585
R11789 gnd.n4430 gnd.n1410 585
R11790 gnd.n1417 gnd.n1410 585
R11791 gnd.n4432 gnd.n4431 585
R11792 gnd.n4433 gnd.n4432 585
R11793 gnd.n1411 gnd.n1407 585
R11794 gnd.n4434 gnd.n1407 585
R11795 gnd.n4123 gnd.n1826 585
R11796 gnd.n1826 gnd.n1406 585
R11797 gnd.n4125 gnd.n4124 585
R11798 gnd.n4126 gnd.n4125 585
R11799 gnd.n1827 gnd.n1825 585
R11800 gnd.n1825 gnd.n1823 585
R11801 gnd.n4117 gnd.n4116 585
R11802 gnd.n4116 gnd.n4115 585
R11803 gnd.n1830 gnd.n1829 585
R11804 gnd.n1831 gnd.n1830 585
R11805 gnd.n4104 gnd.n4103 585
R11806 gnd.n4105 gnd.n4104 585
R11807 gnd.n1840 gnd.n1839 585
R11808 gnd.n1845 gnd.n1839 585
R11809 gnd.n4099 gnd.n4098 585
R11810 gnd.n4098 gnd.n4097 585
R11811 gnd.n1843 gnd.n1842 585
R11812 gnd.n1844 gnd.n1843 585
R11813 gnd.n4088 gnd.n4087 585
R11814 gnd.n4089 gnd.n4088 585
R11815 gnd.n1854 gnd.n1853 585
R11816 gnd.n1853 gnd.n1851 585
R11817 gnd.n4083 gnd.n4082 585
R11818 gnd.n4082 gnd.n4081 585
R11819 gnd.n1857 gnd.n1856 585
R11820 gnd.n1858 gnd.n1857 585
R11821 gnd.n4072 gnd.n4071 585
R11822 gnd.n4073 gnd.n4072 585
R11823 gnd.n1867 gnd.n1866 585
R11824 gnd.n1866 gnd.n1864 585
R11825 gnd.n4067 gnd.n4066 585
R11826 gnd.n4066 gnd.n4065 585
R11827 gnd.n1870 gnd.n1869 585
R11828 gnd.n1871 gnd.n1870 585
R11829 gnd.n4056 gnd.n4055 585
R11830 gnd.n4057 gnd.n4056 585
R11831 gnd.n1880 gnd.n1879 585
R11832 gnd.n1879 gnd.n1877 585
R11833 gnd.n4051 gnd.n4050 585
R11834 gnd.n4050 gnd.n4049 585
R11835 gnd.n1883 gnd.n1882 585
R11836 gnd.n1890 gnd.n1883 585
R11837 gnd.n4040 gnd.n4039 585
R11838 gnd.n4041 gnd.n4040 585
R11839 gnd.n1892 gnd.n1891 585
R11840 gnd.n3255 gnd.n1891 585
R11841 gnd.n4035 gnd.n4034 585
R11842 gnd.n4034 gnd.n4033 585
R11843 gnd.n1895 gnd.n1894 585
R11844 gnd.n1905 gnd.n1895 585
R11845 gnd.n4024 gnd.n4023 585
R11846 gnd.n4025 gnd.n4024 585
R11847 gnd.n1907 gnd.n1906 585
R11848 gnd.t156 gnd.n1906 585
R11849 gnd.n4019 gnd.n4018 585
R11850 gnd.n4018 gnd.n4017 585
R11851 gnd.n1910 gnd.n1909 585
R11852 gnd.n3395 gnd.n1910 585
R11853 gnd.n4008 gnd.n4007 585
R11854 gnd.n4009 gnd.n4008 585
R11855 gnd.n1921 gnd.n1920 585
R11856 gnd.n3154 gnd.n1920 585
R11857 gnd.n4003 gnd.n4002 585
R11858 gnd.n4002 gnd.n4001 585
R11859 gnd.n1924 gnd.n1923 585
R11860 gnd.n3410 gnd.n1924 585
R11861 gnd.n3992 gnd.n3991 585
R11862 gnd.n3993 gnd.n3992 585
R11863 gnd.n1934 gnd.n1933 585
R11864 gnd.n3141 gnd.n1933 585
R11865 gnd.n3987 gnd.n3986 585
R11866 gnd.n3986 gnd.n3985 585
R11867 gnd.n1937 gnd.n1936 585
R11868 gnd.n3135 gnd.n1937 585
R11869 gnd.n3976 gnd.n3975 585
R11870 gnd.n3977 gnd.n3976 585
R11871 gnd.n1949 gnd.n1948 585
R11872 gnd.n3131 gnd.n1948 585
R11873 gnd.n3971 gnd.n3970 585
R11874 gnd.n3970 gnd.n3969 585
R11875 gnd.n1952 gnd.n1951 585
R11876 gnd.n3122 gnd.n1952 585
R11877 gnd.n3960 gnd.n3959 585
R11878 gnd.n3961 gnd.n3960 585
R11879 gnd.n1962 gnd.n1961 585
R11880 gnd.n3449 gnd.n1961 585
R11881 gnd.n3955 gnd.n3954 585
R11882 gnd.n3954 gnd.n3953 585
R11883 gnd.n1965 gnd.n1964 585
R11884 gnd.n3109 gnd.n1965 585
R11885 gnd.n3944 gnd.n3943 585
R11886 gnd.n3945 gnd.n3944 585
R11887 gnd.n1977 gnd.n1976 585
R11888 gnd.n3464 gnd.n1976 585
R11889 gnd.n3939 gnd.n3938 585
R11890 gnd.n3938 gnd.n3937 585
R11891 gnd.n1980 gnd.n1979 585
R11892 gnd.n3095 gnd.n1980 585
R11893 gnd.n3928 gnd.n3927 585
R11894 gnd.n3929 gnd.n3928 585
R11895 gnd.n1991 gnd.n1990 585
R11896 gnd.n3479 gnd.n1990 585
R11897 gnd.n3923 gnd.n3922 585
R11898 gnd.n3922 gnd.n3921 585
R11899 gnd.n1994 gnd.n1993 585
R11900 gnd.n3082 gnd.n1994 585
R11901 gnd.n3912 gnd.n3911 585
R11902 gnd.n3913 gnd.n3912 585
R11903 gnd.n2004 gnd.n2003 585
R11904 gnd.n3494 gnd.n2003 585
R11905 gnd.n3907 gnd.n3906 585
R11906 gnd.n3906 gnd.n3905 585
R11907 gnd.n2007 gnd.n2006 585
R11908 gnd.n3073 gnd.n2007 585
R11909 gnd.n3896 gnd.n3895 585
R11910 gnd.n3897 gnd.n3896 585
R11911 gnd.n2019 gnd.n2018 585
R11912 gnd.n2024 gnd.n2018 585
R11913 gnd.n3891 gnd.n3890 585
R11914 gnd.n3890 gnd.n3889 585
R11915 gnd.n2022 gnd.n2021 585
R11916 gnd.n3054 gnd.n2022 585
R11917 gnd.n3880 gnd.n3879 585
R11918 gnd.n3881 gnd.n3880 585
R11919 gnd.n2034 gnd.n2033 585
R11920 gnd.n3042 gnd.n2033 585
R11921 gnd.n3875 gnd.n3874 585
R11922 gnd.n3874 gnd.n3873 585
R11923 gnd.n2037 gnd.n2036 585
R11924 gnd.n3524 gnd.n2037 585
R11925 gnd.n3864 gnd.n3863 585
R11926 gnd.n3865 gnd.n3864 585
R11927 gnd.n2047 gnd.n2046 585
R11928 gnd.n3029 gnd.n2046 585
R11929 gnd.n3859 gnd.n3858 585
R11930 gnd.n3858 gnd.n3857 585
R11931 gnd.n2050 gnd.n2049 585
R11932 gnd.n3022 gnd.n2050 585
R11933 gnd.n3848 gnd.n3847 585
R11934 gnd.n3849 gnd.n3848 585
R11935 gnd.n2062 gnd.n2061 585
R11936 gnd.n3015 gnd.n2061 585
R11937 gnd.n3843 gnd.n3842 585
R11938 gnd.n3842 gnd.n3841 585
R11939 gnd.n2065 gnd.n2064 585
R11940 gnd.n3009 gnd.n2065 585
R11941 gnd.n3832 gnd.n3831 585
R11942 gnd.n3833 gnd.n3832 585
R11943 gnd.n2077 gnd.n2076 585
R11944 gnd.n3005 gnd.n2076 585
R11945 gnd.n3827 gnd.n3826 585
R11946 gnd.n3826 gnd.n3825 585
R11947 gnd.n2080 gnd.n2079 585
R11948 gnd.n2999 gnd.n2080 585
R11949 gnd.n3816 gnd.n3815 585
R11950 gnd.n3817 gnd.n3816 585
R11951 gnd.n2089 gnd.n2088 585
R11952 gnd.n2093 gnd.n2088 585
R11953 gnd.n3811 gnd.n3810 585
R11954 gnd.n3810 gnd.n3809 585
R11955 gnd.n2092 gnd.n2091 585
R11956 gnd.n2101 gnd.n2092 585
R11957 gnd.n3800 gnd.n3799 585
R11958 gnd.n3801 gnd.n3800 585
R11959 gnd.n2103 gnd.n2102 585
R11960 gnd.n2102 gnd.n2099 585
R11961 gnd.n3795 gnd.n3794 585
R11962 gnd.n3794 gnd.n3793 585
R11963 gnd.n2106 gnd.n2105 585
R11964 gnd.n2107 gnd.n2106 585
R11965 gnd.n3784 gnd.n3783 585
R11966 gnd.n3785 gnd.n3784 585
R11967 gnd.n2116 gnd.n2115 585
R11968 gnd.n2115 gnd.n2113 585
R11969 gnd.n3779 gnd.n3778 585
R11970 gnd.n3778 gnd.n3777 585
R11971 gnd.n2119 gnd.n2118 585
R11972 gnd.n2120 gnd.n2119 585
R11973 gnd.n3768 gnd.n3767 585
R11974 gnd.n3769 gnd.n3768 585
R11975 gnd.n2129 gnd.n2128 585
R11976 gnd.n2128 gnd.n2126 585
R11977 gnd.n3763 gnd.n3762 585
R11978 gnd.n3762 gnd.n3761 585
R11979 gnd.n2132 gnd.n2131 585
R11980 gnd.n2133 gnd.n2132 585
R11981 gnd.n3752 gnd.n3751 585
R11982 gnd.n3753 gnd.n3752 585
R11983 gnd.n2141 gnd.n2140 585
R11984 gnd.n2146 gnd.n2140 585
R11985 gnd.n3747 gnd.n3746 585
R11986 gnd.n3746 gnd.n3745 585
R11987 gnd.n2144 gnd.n2143 585
R11988 gnd.n2145 gnd.n2144 585
R11989 gnd.n3736 gnd.n3735 585
R11990 gnd.n3737 gnd.n3736 585
R11991 gnd.n2155 gnd.n2154 585
R11992 gnd.n2154 gnd.n2152 585
R11993 gnd.n3731 gnd.n3730 585
R11994 gnd.n3730 gnd.n3729 585
R11995 gnd.n2158 gnd.n2157 585
R11996 gnd.n2159 gnd.n2158 585
R11997 gnd.n2743 gnd.n2742 585
R11998 gnd.n2743 gnd.n2178 585
R11999 gnd.n2744 gnd.n2739 585
R12000 gnd.n2744 gnd.n2165 585
R12001 gnd.n2747 gnd.n2746 585
R12002 gnd.n2746 gnd.n2745 585
R12003 gnd.n2748 gnd.n2734 585
R12004 gnd.n2734 gnd.n2250 585
R12005 gnd.n2750 gnd.n2749 585
R12006 gnd.n2750 gnd.n2234 585
R12007 gnd.n2751 gnd.n2733 585
R12008 gnd.n2751 gnd.n1273 585
R12009 gnd.n2753 gnd.n2752 585
R12010 gnd.n2752 gnd.n1270 585
R12011 gnd.n2754 gnd.n2728 585
R12012 gnd.n2728 gnd.n2316 585
R12013 gnd.n2756 gnd.n2755 585
R12014 gnd.n2756 gnd.n1261 585
R12015 gnd.n2757 gnd.n2727 585
R12016 gnd.n2757 gnd.n1253 585
R12017 gnd.n2759 gnd.n2758 585
R12018 gnd.n2758 gnd.n1250 585
R12019 gnd.n2760 gnd.n2329 585
R12020 gnd.n2329 gnd.n1242 585
R12021 gnd.n2762 gnd.n2761 585
R12022 gnd.n2763 gnd.n2762 585
R12023 gnd.n2330 gnd.n2328 585
R12024 gnd.n2328 gnd.n1232 585
R12025 gnd.n2721 gnd.n2720 585
R12026 gnd.n2720 gnd.n1229 585
R12027 gnd.n2719 gnd.n2332 585
R12028 gnd.n2719 gnd.n1221 585
R12029 gnd.n2718 gnd.n2717 585
R12030 gnd.n2718 gnd.n1218 585
R12031 gnd.n2334 gnd.n2333 585
R12032 gnd.n2681 gnd.n2333 585
R12033 gnd.n2713 gnd.n2712 585
R12034 gnd.n2712 gnd.n1208 585
R12035 gnd.n2711 gnd.n2336 585
R12036 gnd.n2711 gnd.n1200 585
R12037 gnd.n2710 gnd.n2338 585
R12038 gnd.n2710 gnd.n2709 585
R12039 gnd.n2376 gnd.n2337 585
R12040 gnd.n2337 gnd.n1190 585
R12041 gnd.n2378 gnd.n2377 585
R12042 gnd.n2377 gnd.n1187 585
R12043 gnd.n2379 gnd.n2370 585
R12044 gnd.n2370 gnd.n1179 585
R12045 gnd.n2381 gnd.n2380 585
R12046 gnd.n2381 gnd.n1176 585
R12047 gnd.n2382 gnd.n2369 585
R12048 gnd.n2382 gnd.n2356 585
R12049 gnd.n2384 gnd.n2383 585
R12050 gnd.n2383 gnd.n1166 585
R12051 gnd.n2367 gnd.n2365 585
R12052 gnd.n2365 gnd.n1159 585
R12053 gnd.n2642 gnd.n2641 585
R12054 gnd.n2643 gnd.n2642 585
R12055 gnd.n2366 gnd.n2364 585
R12056 gnd.n2364 gnd.n1149 585
R12057 gnd.n2592 gnd.n2591 585
R12058 gnd.n2591 gnd.n1146 585
R12059 gnd.n2594 gnd.n2593 585
R12060 gnd.n2594 gnd.n1141 585
R12061 gnd.n2596 gnd.n2595 585
R12062 gnd.n2595 gnd.n1138 585
R12063 gnd.n2598 gnd.n2597 585
R12064 gnd.n2599 gnd.n2598 585
R12065 gnd.n2590 gnd.n2589 585
R12066 gnd.n2590 gnd.n1128 585
R12067 gnd.n2588 gnd.n2398 585
R12068 gnd.n2398 gnd.n1122 585
R12069 gnd.n2635 gnd.n2392 585
R12070 gnd.n2635 gnd.n2634 585
R12071 gnd.n2637 gnd.n2636 585
R12072 gnd.n2636 gnd.n1112 585
R12073 gnd.n2397 gnd.n2391 585
R12074 gnd.n2397 gnd.n1109 585
R12075 gnd.n2396 gnd.n2395 585
R12076 gnd.n2396 gnd.n1101 585
R12077 gnd.n4436 gnd.n4435 585
R12078 gnd.n4435 gnd.n4434 585
R12079 gnd.n4437 gnd.n1404 585
R12080 gnd.n1406 gnd.n1404 585
R12081 gnd.n1824 gnd.n1402 585
R12082 gnd.n4126 gnd.n1824 585
R12083 gnd.n4441 gnd.n1401 585
R12084 gnd.n1823 gnd.n1401 585
R12085 gnd.n4442 gnd.n1400 585
R12086 gnd.n4115 gnd.n1400 585
R12087 gnd.n4443 gnd.n1399 585
R12088 gnd.n1831 gnd.n1399 585
R12089 gnd.n1838 gnd.n1397 585
R12090 gnd.n4105 gnd.n1838 585
R12091 gnd.n4447 gnd.n1396 585
R12092 gnd.n1845 gnd.n1396 585
R12093 gnd.n4448 gnd.n1395 585
R12094 gnd.n4097 gnd.n1395 585
R12095 gnd.n4449 gnd.n1394 585
R12096 gnd.n1844 gnd.n1394 585
R12097 gnd.n1852 gnd.n1392 585
R12098 gnd.n4089 gnd.n1852 585
R12099 gnd.n4453 gnd.n1391 585
R12100 gnd.n1851 gnd.n1391 585
R12101 gnd.n4454 gnd.n1390 585
R12102 gnd.n4081 gnd.n1390 585
R12103 gnd.n4455 gnd.n1389 585
R12104 gnd.n1858 gnd.n1389 585
R12105 gnd.n1865 gnd.n1387 585
R12106 gnd.n4073 gnd.n1865 585
R12107 gnd.n4459 gnd.n1386 585
R12108 gnd.n1864 gnd.n1386 585
R12109 gnd.n4460 gnd.n1385 585
R12110 gnd.n4065 gnd.n1385 585
R12111 gnd.n4461 gnd.n1384 585
R12112 gnd.n1871 gnd.n1384 585
R12113 gnd.n1878 gnd.n1382 585
R12114 gnd.n4057 gnd.n1878 585
R12115 gnd.n4465 gnd.n1381 585
R12116 gnd.n1877 gnd.n1381 585
R12117 gnd.n4466 gnd.n1380 585
R12118 gnd.n4049 gnd.n1380 585
R12119 gnd.n4467 gnd.n1379 585
R12120 gnd.n1890 gnd.n1379 585
R12121 gnd.n1889 gnd.n1377 585
R12122 gnd.n4041 gnd.n1889 585
R12123 gnd.n4471 gnd.n1376 585
R12124 gnd.n3255 gnd.n1376 585
R12125 gnd.n4472 gnd.n1375 585
R12126 gnd.n4033 gnd.n1375 585
R12127 gnd.n4473 gnd.n1374 585
R12128 gnd.n1905 gnd.n1374 585
R12129 gnd.n1904 gnd.n1372 585
R12130 gnd.n4025 gnd.n1904 585
R12131 gnd.n4477 gnd.n1371 585
R12132 gnd.t156 gnd.n1371 585
R12133 gnd.n4478 gnd.n1370 585
R12134 gnd.n4017 gnd.n1370 585
R12135 gnd.n4479 gnd.n1369 585
R12136 gnd.n3395 gnd.n1369 585
R12137 gnd.n1919 gnd.n1367 585
R12138 gnd.n4009 gnd.n1919 585
R12139 gnd.n4483 gnd.n1366 585
R12140 gnd.n3154 gnd.n1366 585
R12141 gnd.n4484 gnd.n1365 585
R12142 gnd.n4001 gnd.n1365 585
R12143 gnd.n4485 gnd.n1364 585
R12144 gnd.n3410 gnd.n1364 585
R12145 gnd.n1932 gnd.n1362 585
R12146 gnd.n3993 gnd.n1932 585
R12147 gnd.n4489 gnd.n1361 585
R12148 gnd.n3141 gnd.n1361 585
R12149 gnd.n4490 gnd.n1360 585
R12150 gnd.n3985 gnd.n1360 585
R12151 gnd.n4491 gnd.n1359 585
R12152 gnd.n3135 gnd.n1359 585
R12153 gnd.n1946 gnd.n1357 585
R12154 gnd.n3977 gnd.n1946 585
R12155 gnd.n4495 gnd.n1356 585
R12156 gnd.n3131 gnd.n1356 585
R12157 gnd.n4496 gnd.n1355 585
R12158 gnd.n3969 gnd.n1355 585
R12159 gnd.n4497 gnd.n1354 585
R12160 gnd.n3122 gnd.n1354 585
R12161 gnd.n1960 gnd.n1352 585
R12162 gnd.n3961 gnd.n1960 585
R12163 gnd.n4501 gnd.n1351 585
R12164 gnd.n3449 gnd.n1351 585
R12165 gnd.n4502 gnd.n1350 585
R12166 gnd.n3953 gnd.n1350 585
R12167 gnd.n4503 gnd.n1349 585
R12168 gnd.n3109 gnd.n1349 585
R12169 gnd.n1974 gnd.n1347 585
R12170 gnd.n3945 gnd.n1974 585
R12171 gnd.n4507 gnd.n1346 585
R12172 gnd.n3464 gnd.n1346 585
R12173 gnd.n4508 gnd.n1345 585
R12174 gnd.n3937 gnd.n1345 585
R12175 gnd.n4509 gnd.n1344 585
R12176 gnd.n3095 gnd.n1344 585
R12177 gnd.n1988 gnd.n1342 585
R12178 gnd.n3929 gnd.n1988 585
R12179 gnd.n4513 gnd.n1341 585
R12180 gnd.n3479 gnd.n1341 585
R12181 gnd.n4514 gnd.n1340 585
R12182 gnd.n3921 gnd.n1340 585
R12183 gnd.n4515 gnd.n1339 585
R12184 gnd.n3082 gnd.n1339 585
R12185 gnd.n2001 gnd.n1337 585
R12186 gnd.n3913 gnd.n2001 585
R12187 gnd.n4519 gnd.n1336 585
R12188 gnd.n3494 gnd.n1336 585
R12189 gnd.n4520 gnd.n1335 585
R12190 gnd.n3905 gnd.n1335 585
R12191 gnd.n4521 gnd.n1334 585
R12192 gnd.n3073 gnd.n1334 585
R12193 gnd.n2016 gnd.n1332 585
R12194 gnd.n3897 gnd.n2016 585
R12195 gnd.n4525 gnd.n1331 585
R12196 gnd.n2024 gnd.n1331 585
R12197 gnd.n4526 gnd.n1330 585
R12198 gnd.n3889 gnd.n1330 585
R12199 gnd.n4527 gnd.n1329 585
R12200 gnd.n3054 gnd.n1329 585
R12201 gnd.n2031 gnd.n1327 585
R12202 gnd.n3881 gnd.n2031 585
R12203 gnd.n4531 gnd.n1326 585
R12204 gnd.n3042 gnd.n1326 585
R12205 gnd.n4532 gnd.n1325 585
R12206 gnd.n3873 gnd.n1325 585
R12207 gnd.n4533 gnd.n1324 585
R12208 gnd.n3524 gnd.n1324 585
R12209 gnd.n2045 gnd.n1322 585
R12210 gnd.n3865 gnd.n2045 585
R12211 gnd.n4537 gnd.n1321 585
R12212 gnd.n3029 gnd.n1321 585
R12213 gnd.n4538 gnd.n1320 585
R12214 gnd.n3857 gnd.n1320 585
R12215 gnd.n4539 gnd.n1319 585
R12216 gnd.n3022 gnd.n1319 585
R12217 gnd.n2059 gnd.n1317 585
R12218 gnd.n3849 gnd.n2059 585
R12219 gnd.n4543 gnd.n1316 585
R12220 gnd.n3015 gnd.n1316 585
R12221 gnd.n4544 gnd.n1315 585
R12222 gnd.n3841 gnd.n1315 585
R12223 gnd.n4545 gnd.n1314 585
R12224 gnd.n3009 gnd.n1314 585
R12225 gnd.n2074 gnd.n1312 585
R12226 gnd.n3833 gnd.n2074 585
R12227 gnd.n4549 gnd.n1311 585
R12228 gnd.n3005 gnd.n1311 585
R12229 gnd.n4550 gnd.n1310 585
R12230 gnd.n3825 gnd.n1310 585
R12231 gnd.n4551 gnd.n1309 585
R12232 gnd.n2999 gnd.n1309 585
R12233 gnd.n2087 gnd.n1307 585
R12234 gnd.n3817 gnd.n2087 585
R12235 gnd.n4555 gnd.n1306 585
R12236 gnd.n2093 gnd.n1306 585
R12237 gnd.n4556 gnd.n1305 585
R12238 gnd.n3809 gnd.n1305 585
R12239 gnd.n4557 gnd.n1304 585
R12240 gnd.n2101 gnd.n1304 585
R12241 gnd.n2100 gnd.n1302 585
R12242 gnd.n3801 gnd.n2100 585
R12243 gnd.n4561 gnd.n1301 585
R12244 gnd.n2099 gnd.n1301 585
R12245 gnd.n4562 gnd.n1300 585
R12246 gnd.n3793 gnd.n1300 585
R12247 gnd.n4563 gnd.n1299 585
R12248 gnd.n2107 gnd.n1299 585
R12249 gnd.n2114 gnd.n1297 585
R12250 gnd.n3785 gnd.n2114 585
R12251 gnd.n4567 gnd.n1296 585
R12252 gnd.n2113 gnd.n1296 585
R12253 gnd.n4568 gnd.n1295 585
R12254 gnd.n3777 gnd.n1295 585
R12255 gnd.n4569 gnd.n1294 585
R12256 gnd.n2120 gnd.n1294 585
R12257 gnd.n2127 gnd.n1292 585
R12258 gnd.n3769 gnd.n2127 585
R12259 gnd.n4573 gnd.n1291 585
R12260 gnd.n2126 gnd.n1291 585
R12261 gnd.n4574 gnd.n1290 585
R12262 gnd.n3761 gnd.n1290 585
R12263 gnd.n4575 gnd.n1289 585
R12264 gnd.n2133 gnd.n1289 585
R12265 gnd.n2139 gnd.n1287 585
R12266 gnd.n3753 gnd.n2139 585
R12267 gnd.n4579 gnd.n1286 585
R12268 gnd.n2146 gnd.n1286 585
R12269 gnd.n4580 gnd.n1285 585
R12270 gnd.n3745 gnd.n1285 585
R12271 gnd.n4581 gnd.n1284 585
R12272 gnd.n2145 gnd.n1284 585
R12273 gnd.n2153 gnd.n1282 585
R12274 gnd.n3737 gnd.n2153 585
R12275 gnd.n4585 gnd.n1281 585
R12276 gnd.n2152 gnd.n1281 585
R12277 gnd.n4586 gnd.n1280 585
R12278 gnd.n3729 gnd.n1280 585
R12279 gnd.n4587 gnd.n1279 585
R12280 gnd.n2159 gnd.n1279 585
R12281 gnd.n3718 gnd.n3717 585
R12282 gnd.n3716 gnd.n2180 585
R12283 gnd.n2182 gnd.n2179 585
R12284 gnd.n3720 gnd.n2179 585
R12285 gnd.n3709 gnd.n2190 585
R12286 gnd.n3708 gnd.n2191 585
R12287 gnd.n2193 gnd.n2192 585
R12288 gnd.n3701 gnd.n2199 585
R12289 gnd.n3700 gnd.n2200 585
R12290 gnd.n2207 gnd.n2201 585
R12291 gnd.n3693 gnd.n2208 585
R12292 gnd.n3692 gnd.n2209 585
R12293 gnd.n2211 gnd.n2210 585
R12294 gnd.n3685 gnd.n2217 585
R12295 gnd.n3684 gnd.n2218 585
R12296 gnd.n2227 gnd.n2219 585
R12297 gnd.n3677 gnd.n2228 585
R12298 gnd.n3676 gnd.n2229 585
R12299 gnd.n2231 gnd.n2230 585
R12300 gnd.n2814 gnd.n2787 585
R12301 gnd.n2813 gnd.n2788 585
R12302 gnd.n2812 gnd.n2789 585
R12303 gnd.n2791 gnd.n2790 585
R12304 gnd.n2808 gnd.n2793 585
R12305 gnd.n2807 gnd.n2794 585
R12306 gnd.n2806 gnd.n2795 585
R12307 gnd.n2803 gnd.n2800 585
R12308 gnd.n2802 gnd.n2801 585
R12309 gnd.n2164 gnd.n2163 585
R12310 gnd.n3723 gnd.n3722 585
R12311 gnd.n4130 gnd.n1408 585
R12312 gnd.n4434 gnd.n1408 585
R12313 gnd.n4129 gnd.n4128 585
R12314 gnd.n4128 gnd.n1406 585
R12315 gnd.n4127 gnd.n1821 585
R12316 gnd.n4127 gnd.n4126 585
R12317 gnd.n1834 gnd.n1822 585
R12318 gnd.n1823 gnd.n1822 585
R12319 gnd.n4114 gnd.n4113 585
R12320 gnd.n4115 gnd.n4114 585
R12321 gnd.n1833 gnd.n1832 585
R12322 gnd.n1832 gnd.n1831 585
R12323 gnd.n4107 gnd.n4106 585
R12324 gnd.n4106 gnd.n4105 585
R12325 gnd.n1837 gnd.n1836 585
R12326 gnd.n1845 gnd.n1837 585
R12327 gnd.n4096 gnd.n4095 585
R12328 gnd.n4097 gnd.n4096 585
R12329 gnd.n1847 gnd.n1846 585
R12330 gnd.n1846 gnd.n1844 585
R12331 gnd.n4091 gnd.n4090 585
R12332 gnd.n4090 gnd.n4089 585
R12333 gnd.n1850 gnd.n1849 585
R12334 gnd.n1851 gnd.n1850 585
R12335 gnd.n4080 gnd.n4079 585
R12336 gnd.n4081 gnd.n4080 585
R12337 gnd.n1860 gnd.n1859 585
R12338 gnd.n1859 gnd.n1858 585
R12339 gnd.n4075 gnd.n4074 585
R12340 gnd.n4074 gnd.n4073 585
R12341 gnd.n1863 gnd.n1862 585
R12342 gnd.n1864 gnd.n1863 585
R12343 gnd.n4064 gnd.n4063 585
R12344 gnd.n4065 gnd.n4064 585
R12345 gnd.n1873 gnd.n1872 585
R12346 gnd.n1872 gnd.n1871 585
R12347 gnd.n4059 gnd.n4058 585
R12348 gnd.n4058 gnd.n4057 585
R12349 gnd.n1876 gnd.n1875 585
R12350 gnd.n1877 gnd.n1876 585
R12351 gnd.n4048 gnd.n4047 585
R12352 gnd.n4049 gnd.n4048 585
R12353 gnd.n1885 gnd.n1884 585
R12354 gnd.n1890 gnd.n1884 585
R12355 gnd.n4043 gnd.n4042 585
R12356 gnd.n4042 gnd.n4041 585
R12357 gnd.n1888 gnd.n1887 585
R12358 gnd.n3255 gnd.n1888 585
R12359 gnd.n4032 gnd.n4031 585
R12360 gnd.n4033 gnd.n4032 585
R12361 gnd.n1899 gnd.n1898 585
R12362 gnd.n1905 gnd.n1898 585
R12363 gnd.n4027 gnd.n4026 585
R12364 gnd.n4026 gnd.n4025 585
R12365 gnd.n1902 gnd.n1901 585
R12366 gnd.t156 gnd.n1902 585
R12367 gnd.n4016 gnd.n4015 585
R12368 gnd.n4017 gnd.n4016 585
R12369 gnd.n1914 gnd.n1913 585
R12370 gnd.n3395 gnd.n1913 585
R12371 gnd.n4011 gnd.n4010 585
R12372 gnd.n4010 gnd.n4009 585
R12373 gnd.n1917 gnd.n1916 585
R12374 gnd.n3154 gnd.n1917 585
R12375 gnd.n4000 gnd.n3999 585
R12376 gnd.n4001 gnd.n4000 585
R12377 gnd.n1927 gnd.n1926 585
R12378 gnd.n3410 gnd.n1926 585
R12379 gnd.n3995 gnd.n3994 585
R12380 gnd.n3994 gnd.n3993 585
R12381 gnd.n1930 gnd.n1929 585
R12382 gnd.n3141 gnd.n1930 585
R12383 gnd.n3984 gnd.n3983 585
R12384 gnd.n3985 gnd.n3984 585
R12385 gnd.n1941 gnd.n1940 585
R12386 gnd.n3135 gnd.n1940 585
R12387 gnd.n3979 gnd.n3978 585
R12388 gnd.n3978 gnd.n3977 585
R12389 gnd.n1944 gnd.n1943 585
R12390 gnd.n3131 gnd.n1944 585
R12391 gnd.n3968 gnd.n3967 585
R12392 gnd.n3969 gnd.n3968 585
R12393 gnd.n1955 gnd.n1954 585
R12394 gnd.n3122 gnd.n1954 585
R12395 gnd.n3963 gnd.n3962 585
R12396 gnd.n3962 gnd.n3961 585
R12397 gnd.n1958 gnd.n1957 585
R12398 gnd.n3449 gnd.n1958 585
R12399 gnd.n3952 gnd.n3951 585
R12400 gnd.n3953 gnd.n3952 585
R12401 gnd.n1969 gnd.n1968 585
R12402 gnd.n3109 gnd.n1968 585
R12403 gnd.n3947 gnd.n3946 585
R12404 gnd.n3946 gnd.n3945 585
R12405 gnd.n1972 gnd.n1971 585
R12406 gnd.n3464 gnd.n1972 585
R12407 gnd.n3936 gnd.n3935 585
R12408 gnd.n3937 gnd.n3936 585
R12409 gnd.n1983 gnd.n1982 585
R12410 gnd.n3095 gnd.n1982 585
R12411 gnd.n3931 gnd.n3930 585
R12412 gnd.n3930 gnd.n3929 585
R12413 gnd.n1986 gnd.n1985 585
R12414 gnd.n3479 gnd.n1986 585
R12415 gnd.n3920 gnd.n3919 585
R12416 gnd.n3921 gnd.n3920 585
R12417 gnd.n1997 gnd.n1996 585
R12418 gnd.n3082 gnd.n1996 585
R12419 gnd.n3915 gnd.n3914 585
R12420 gnd.n3914 gnd.n3913 585
R12421 gnd.n2000 gnd.n1999 585
R12422 gnd.n3494 gnd.n2000 585
R12423 gnd.n3904 gnd.n3903 585
R12424 gnd.n3905 gnd.n3904 585
R12425 gnd.n2011 gnd.n2010 585
R12426 gnd.n3073 gnd.n2010 585
R12427 gnd.n3899 gnd.n3898 585
R12428 gnd.n3898 gnd.n3897 585
R12429 gnd.n2014 gnd.n2013 585
R12430 gnd.n2024 gnd.n2014 585
R12431 gnd.n3888 gnd.n3887 585
R12432 gnd.n3889 gnd.n3888 585
R12433 gnd.n2027 gnd.n2026 585
R12434 gnd.n3054 gnd.n2026 585
R12435 gnd.n3883 gnd.n3882 585
R12436 gnd.n3882 gnd.n3881 585
R12437 gnd.n2030 gnd.n2029 585
R12438 gnd.n3042 gnd.n2030 585
R12439 gnd.n3872 gnd.n3871 585
R12440 gnd.n3873 gnd.n3872 585
R12441 gnd.n2040 gnd.n2039 585
R12442 gnd.n3524 gnd.n2039 585
R12443 gnd.n3867 gnd.n3866 585
R12444 gnd.n3866 gnd.n3865 585
R12445 gnd.n2043 gnd.n2042 585
R12446 gnd.n3029 gnd.n2043 585
R12447 gnd.n3856 gnd.n3855 585
R12448 gnd.n3857 gnd.n3856 585
R12449 gnd.n2054 gnd.n2053 585
R12450 gnd.n3022 gnd.n2053 585
R12451 gnd.n3851 gnd.n3850 585
R12452 gnd.n3850 gnd.n3849 585
R12453 gnd.n2057 gnd.n2056 585
R12454 gnd.n3015 gnd.n2057 585
R12455 gnd.n3840 gnd.n3839 585
R12456 gnd.n3841 gnd.n3840 585
R12457 gnd.n2069 gnd.n2068 585
R12458 gnd.n3009 gnd.n2068 585
R12459 gnd.n3835 gnd.n3834 585
R12460 gnd.n3834 gnd.n3833 585
R12461 gnd.n2072 gnd.n2071 585
R12462 gnd.n3005 gnd.n2072 585
R12463 gnd.n3824 gnd.n3823 585
R12464 gnd.n3825 gnd.n3824 585
R12465 gnd.n2082 gnd.n2081 585
R12466 gnd.n2999 gnd.n2081 585
R12467 gnd.n3819 gnd.n3818 585
R12468 gnd.n3818 gnd.n3817 585
R12469 gnd.n2085 gnd.n2084 585
R12470 gnd.n2093 gnd.n2085 585
R12471 gnd.n3808 gnd.n3807 585
R12472 gnd.n3809 gnd.n3808 585
R12473 gnd.n2095 gnd.n2094 585
R12474 gnd.n2101 gnd.n2094 585
R12475 gnd.n3803 gnd.n3802 585
R12476 gnd.n3802 gnd.n3801 585
R12477 gnd.n2098 gnd.n2097 585
R12478 gnd.n2099 gnd.n2098 585
R12479 gnd.n3792 gnd.n3791 585
R12480 gnd.n3793 gnd.n3792 585
R12481 gnd.n2109 gnd.n2108 585
R12482 gnd.n2108 gnd.n2107 585
R12483 gnd.n3787 gnd.n3786 585
R12484 gnd.n3786 gnd.n3785 585
R12485 gnd.n2112 gnd.n2111 585
R12486 gnd.n2113 gnd.n2112 585
R12487 gnd.n3776 gnd.n3775 585
R12488 gnd.n3777 gnd.n3776 585
R12489 gnd.n2122 gnd.n2121 585
R12490 gnd.n2121 gnd.n2120 585
R12491 gnd.n3771 gnd.n3770 585
R12492 gnd.n3770 gnd.n3769 585
R12493 gnd.n2125 gnd.n2124 585
R12494 gnd.n2126 gnd.n2125 585
R12495 gnd.n3760 gnd.n3759 585
R12496 gnd.n3761 gnd.n3760 585
R12497 gnd.n2135 gnd.n2134 585
R12498 gnd.n2134 gnd.n2133 585
R12499 gnd.n3755 gnd.n3754 585
R12500 gnd.n3754 gnd.n3753 585
R12501 gnd.n2138 gnd.n2137 585
R12502 gnd.n2146 gnd.n2138 585
R12503 gnd.n3744 gnd.n3743 585
R12504 gnd.n3745 gnd.n3744 585
R12505 gnd.n2148 gnd.n2147 585
R12506 gnd.n2147 gnd.n2145 585
R12507 gnd.n3739 gnd.n3738 585
R12508 gnd.n3738 gnd.n3737 585
R12509 gnd.n2151 gnd.n2150 585
R12510 gnd.n2152 gnd.n2151 585
R12511 gnd.n3728 gnd.n3727 585
R12512 gnd.n3729 gnd.n3728 585
R12513 gnd.n2161 gnd.n2160 585
R12514 gnd.n2160 gnd.n2159 585
R12515 gnd.n4137 gnd.n4136 585
R12516 gnd.n4136 gnd.n1409 585
R12517 gnd.n4138 gnd.n4135 585
R12518 gnd.n4133 gnd.n1819 585
R12519 gnd.n4142 gnd.n1818 585
R12520 gnd.n4146 gnd.n1816 585
R12521 gnd.n4147 gnd.n1815 585
R12522 gnd.n1813 gnd.n1811 585
R12523 gnd.n4151 gnd.n1810 585
R12524 gnd.n4152 gnd.n1808 585
R12525 gnd.n4153 gnd.n1807 585
R12526 gnd.n1805 gnd.n1685 585
R12527 gnd.n1804 gnd.n1803 585
R12528 gnd.n1793 gnd.n1687 585
R12529 gnd.n1795 gnd.n1794 585
R12530 gnd.n1791 gnd.n1697 585
R12531 gnd.n1790 gnd.n1789 585
R12532 gnd.n1777 gnd.n1699 585
R12533 gnd.n1779 gnd.n1778 585
R12534 gnd.n1775 gnd.n1703 585
R12535 gnd.n1774 gnd.n1773 585
R12536 gnd.n1758 gnd.n1705 585
R12537 gnd.n1760 gnd.n1759 585
R12538 gnd.n1756 gnd.n1710 585
R12539 gnd.n1755 gnd.n1754 585
R12540 gnd.n1739 gnd.n1712 585
R12541 gnd.n1741 gnd.n1740 585
R12542 gnd.n1737 gnd.n1717 585
R12543 gnd.n1736 gnd.n1735 585
R12544 gnd.n1719 gnd.n1405 585
R12545 gnd.n2874 gnd.t166 543.808
R12546 gnd.n3223 gnd.t163 543.808
R12547 gnd.n2929 gnd.t119 543.808
R12548 gnd.n3217 gnd.t112 543.808
R12549 gnd.n3375 gnd.n3175 458.866
R12550 gnd.n3258 gnd.n3257 458.866
R12551 gnd.n3574 gnd.n3572 458.866
R12552 gnd.n3570 gnd.n2893 458.866
R12553 gnd.n6427 gnd.n6426 404.397
R12554 gnd.n2796 gnd.t126 371.625
R12555 gnd.n7331 gnd.t142 371.625
R12556 gnd.n1691 gnd.t136 371.625
R12557 gnd.n2223 gnd.t158 371.625
R12558 gnd.n1469 gnd.t109 371.625
R12559 gnd.n1491 gnd.t98 371.625
R12560 gnd.n179 gnd.t172 371.625
R12561 gnd.n7424 gnd.t94 371.625
R12562 gnd.n983 gnd.t72 371.625
R12563 gnd.n1005 gnd.t152 371.625
R12564 gnd.n2312 gnd.t169 371.625
R12565 gnd.n2290 gnd.t86 371.625
R12566 gnd.n2477 gnd.t102 371.625
R12567 gnd.n4143 gnd.t82 371.625
R12568 gnd.n5212 gnd.t148 323.425
R12569 gnd.n4863 gnd.t90 323.425
R12570 gnd.n6079 gnd.n6053 289.615
R12571 gnd.n6047 gnd.n6021 289.615
R12572 gnd.n6015 gnd.n5989 289.615
R12573 gnd.n5984 gnd.n5958 289.615
R12574 gnd.n5952 gnd.n5926 289.615
R12575 gnd.n5920 gnd.n5894 289.615
R12576 gnd.n5888 gnd.n5862 289.615
R12577 gnd.n5857 gnd.n5831 289.615
R12578 gnd.n5286 gnd.t105 279.217
R12579 gnd.n4907 gnd.t68 279.217
R12580 gnd.n2901 gnd.t81 260.649
R12581 gnd.n3187 gnd.t118 260.649
R12582 gnd.n2992 gnd.n2086 256.663
R12583 gnd.n2916 gnd.n2086 256.663
R12584 gnd.n2985 gnd.n2086 256.663
R12585 gnd.n2979 gnd.n2086 256.663
R12586 gnd.n2977 gnd.n2086 256.663
R12587 gnd.n2971 gnd.n2086 256.663
R12588 gnd.n2969 gnd.n2086 256.663
R12589 gnd.n2963 gnd.n2086 256.663
R12590 gnd.n2961 gnd.n2086 256.663
R12591 gnd.n2955 gnd.n2086 256.663
R12592 gnd.n2953 gnd.n2086 256.663
R12593 gnd.n2947 gnd.n2086 256.663
R12594 gnd.n2945 gnd.n2086 256.663
R12595 gnd.n2939 gnd.n2086 256.663
R12596 gnd.n2932 gnd.n2086 256.663
R12597 gnd.n2933 gnd.n2086 256.663
R12598 gnd.n3640 gnd.n2872 256.663
R12599 gnd.n3638 gnd.n2086 256.663
R12600 gnd.n3636 gnd.n2086 256.663
R12601 gnd.n3629 gnd.n2086 256.663
R12602 gnd.n3627 gnd.n2086 256.663
R12603 gnd.n3621 gnd.n2086 256.663
R12604 gnd.n3619 gnd.n2086 256.663
R12605 gnd.n3613 gnd.n2086 256.663
R12606 gnd.n3611 gnd.n2086 256.663
R12607 gnd.n3605 gnd.n2086 256.663
R12608 gnd.n3603 gnd.n2086 256.663
R12609 gnd.n3597 gnd.n2086 256.663
R12610 gnd.n3595 gnd.n2086 256.663
R12611 gnd.n3589 gnd.n2086 256.663
R12612 gnd.n3587 gnd.n2086 256.663
R12613 gnd.n3581 gnd.n2086 256.663
R12614 gnd.n3579 gnd.n2086 256.663
R12615 gnd.n3573 gnd.n2086 256.663
R12616 gnd.n3247 gnd.n3196 256.663
R12617 gnd.n3263 gnd.n3196 256.663
R12618 gnd.n3244 gnd.n3196 256.663
R12619 gnd.n3270 gnd.n3196 256.663
R12620 gnd.n3241 gnd.n3196 256.663
R12621 gnd.n3277 gnd.n3196 256.663
R12622 gnd.n3238 gnd.n3196 256.663
R12623 gnd.n3284 gnd.n3196 256.663
R12624 gnd.n3235 gnd.n3196 256.663
R12625 gnd.n3291 gnd.n3196 256.663
R12626 gnd.n3232 gnd.n3196 256.663
R12627 gnd.n3298 gnd.n3196 256.663
R12628 gnd.n3229 gnd.n3196 256.663
R12629 gnd.n3305 gnd.n3196 256.663
R12630 gnd.n3226 gnd.n3196 256.663
R12631 gnd.n3313 gnd.n3196 256.663
R12632 gnd.n3316 gnd.n1466 256.663
R12633 gnd.n3317 gnd.n3196 256.663
R12634 gnd.n3321 gnd.n3196 256.663
R12635 gnd.n3220 gnd.n3196 256.663
R12636 gnd.n3329 gnd.n3196 256.663
R12637 gnd.n3215 gnd.n3196 256.663
R12638 gnd.n3336 gnd.n3196 256.663
R12639 gnd.n3212 gnd.n3196 256.663
R12640 gnd.n3343 gnd.n3196 256.663
R12641 gnd.n3209 gnd.n3196 256.663
R12642 gnd.n3350 gnd.n3196 256.663
R12643 gnd.n3206 gnd.n3196 256.663
R12644 gnd.n3357 gnd.n3196 256.663
R12645 gnd.n3203 gnd.n3196 256.663
R12646 gnd.n3364 gnd.n3196 256.663
R12647 gnd.n3200 gnd.n3196 256.663
R12648 gnd.n3371 gnd.n3196 256.663
R12649 gnd.n3374 gnd.n3196 256.663
R12650 gnd.n4832 gnd.n951 242.672
R12651 gnd.n4832 gnd.n952 242.672
R12652 gnd.n4832 gnd.n953 242.672
R12653 gnd.n4832 gnd.n954 242.672
R12654 gnd.n4832 gnd.n955 242.672
R12655 gnd.n4832 gnd.n956 242.672
R12656 gnd.n4832 gnd.n957 242.672
R12657 gnd.n4832 gnd.n958 242.672
R12658 gnd.n4832 gnd.n959 242.672
R12659 gnd.n3671 gnd.n3670 242.672
R12660 gnd.n3670 gnd.n2249 242.672
R12661 gnd.n3670 gnd.n2248 242.672
R12662 gnd.n3670 gnd.n2246 242.672
R12663 gnd.n3670 gnd.n2244 242.672
R12664 gnd.n3670 gnd.n2243 242.672
R12665 gnd.n3670 gnd.n2241 242.672
R12666 gnd.n3670 gnd.n2239 242.672
R12667 gnd.n3670 gnd.n2238 242.672
R12668 gnd.n4425 gnd.n1436 242.672
R12669 gnd.n4425 gnd.n1437 242.672
R12670 gnd.n4425 gnd.n1438 242.672
R12671 gnd.n4425 gnd.n1439 242.672
R12672 gnd.n4425 gnd.n1440 242.672
R12673 gnd.n4425 gnd.n1441 242.672
R12674 gnd.n4425 gnd.n1442 242.672
R12675 gnd.n4425 gnd.n1443 242.672
R12676 gnd.n4425 gnd.n1444 242.672
R12677 gnd.n7333 gnd.n106 242.672
R12678 gnd.n7329 gnd.n106 242.672
R12679 gnd.n7324 gnd.n106 242.672
R12680 gnd.n7321 gnd.n106 242.672
R12681 gnd.n7316 gnd.n106 242.672
R12682 gnd.n7313 gnd.n106 242.672
R12683 gnd.n7308 gnd.n106 242.672
R12684 gnd.n7305 gnd.n106 242.672
R12685 gnd.n7300 gnd.n106 242.672
R12686 gnd.n5340 gnd.n5339 242.672
R12687 gnd.n5340 gnd.n5250 242.672
R12688 gnd.n5340 gnd.n5251 242.672
R12689 gnd.n5340 gnd.n5252 242.672
R12690 gnd.n5340 gnd.n5253 242.672
R12691 gnd.n5340 gnd.n5254 242.672
R12692 gnd.n5340 gnd.n5255 242.672
R12693 gnd.n5340 gnd.n5256 242.672
R12694 gnd.n5340 gnd.n5257 242.672
R12695 gnd.n5340 gnd.n5258 242.672
R12696 gnd.n5340 gnd.n5259 242.672
R12697 gnd.n5340 gnd.n5260 242.672
R12698 gnd.n5341 gnd.n5340 242.672
R12699 gnd.n6153 gnd.n4833 242.672
R12700 gnd.n6159 gnd.n4833 242.672
R12701 gnd.n4910 gnd.n4833 242.672
R12702 gnd.n6166 gnd.n4833 242.672
R12703 gnd.n4901 gnd.n4833 242.672
R12704 gnd.n6173 gnd.n4833 242.672
R12705 gnd.n4894 gnd.n4833 242.672
R12706 gnd.n6180 gnd.n4833 242.672
R12707 gnd.n4887 gnd.n4833 242.672
R12708 gnd.n6187 gnd.n4833 242.672
R12709 gnd.n4880 gnd.n4833 242.672
R12710 gnd.n6194 gnd.n4833 242.672
R12711 gnd.n4873 gnd.n4833 242.672
R12712 gnd.n5510 gnd.n5509 242.672
R12713 gnd.n5509 gnd.n5162 242.672
R12714 gnd.n5509 gnd.n5163 242.672
R12715 gnd.n5509 gnd.n5164 242.672
R12716 gnd.n5509 gnd.n5165 242.672
R12717 gnd.n5509 gnd.n5166 242.672
R12718 gnd.n5509 gnd.n5167 242.672
R12719 gnd.n5509 gnd.n5168 242.672
R12720 gnd.n6205 gnd.n4833 242.672
R12721 gnd.n4866 gnd.n4833 242.672
R12722 gnd.n6212 gnd.n4833 242.672
R12723 gnd.n4857 gnd.n4833 242.672
R12724 gnd.n6219 gnd.n4833 242.672
R12725 gnd.n4850 gnd.n4833 242.672
R12726 gnd.n6226 gnd.n4833 242.672
R12727 gnd.n4843 gnd.n4833 242.672
R12728 gnd.n4832 gnd.n4831 242.672
R12729 gnd.n4832 gnd.n933 242.672
R12730 gnd.n4832 gnd.n934 242.672
R12731 gnd.n4832 gnd.n935 242.672
R12732 gnd.n4832 gnd.n936 242.672
R12733 gnd.n4832 gnd.n937 242.672
R12734 gnd.n4832 gnd.n938 242.672
R12735 gnd.n4832 gnd.n939 242.672
R12736 gnd.n4832 gnd.n940 242.672
R12737 gnd.n4832 gnd.n941 242.672
R12738 gnd.n4832 gnd.n942 242.672
R12739 gnd.n4832 gnd.n943 242.672
R12740 gnd.n4832 gnd.n944 242.672
R12741 gnd.n4832 gnd.n945 242.672
R12742 gnd.n4832 gnd.n946 242.672
R12743 gnd.n4832 gnd.n947 242.672
R12744 gnd.n4832 gnd.n948 242.672
R12745 gnd.n4832 gnd.n949 242.672
R12746 gnd.n4832 gnd.n950 242.672
R12747 gnd.n3670 gnd.n2251 242.672
R12748 gnd.n3670 gnd.n2252 242.672
R12749 gnd.n3670 gnd.n2253 242.672
R12750 gnd.n3670 gnd.n2254 242.672
R12751 gnd.n3670 gnd.n2255 242.672
R12752 gnd.n3670 gnd.n2256 242.672
R12753 gnd.n3670 gnd.n2257 242.672
R12754 gnd.n3670 gnd.n2258 242.672
R12755 gnd.n3670 gnd.n2259 242.672
R12756 gnd.n3670 gnd.n2260 242.672
R12757 gnd.n3670 gnd.n2261 242.672
R12758 gnd.n3641 gnd.n2292 242.672
R12759 gnd.n3670 gnd.n2262 242.672
R12760 gnd.n3670 gnd.n2263 242.672
R12761 gnd.n3670 gnd.n2264 242.672
R12762 gnd.n3670 gnd.n2265 242.672
R12763 gnd.n3670 gnd.n2266 242.672
R12764 gnd.n3670 gnd.n2267 242.672
R12765 gnd.n3670 gnd.n2268 242.672
R12766 gnd.n3670 gnd.n3669 242.672
R12767 gnd.n4425 gnd.n4424 242.672
R12768 gnd.n4425 gnd.n1418 242.672
R12769 gnd.n4425 gnd.n1419 242.672
R12770 gnd.n4425 gnd.n1420 242.672
R12771 gnd.n4425 gnd.n1421 242.672
R12772 gnd.n4425 gnd.n1422 242.672
R12773 gnd.n4425 gnd.n1423 242.672
R12774 gnd.n4425 gnd.n1424 242.672
R12775 gnd.n4393 gnd.n1467 242.672
R12776 gnd.n4425 gnd.n1425 242.672
R12777 gnd.n4425 gnd.n1426 242.672
R12778 gnd.n4425 gnd.n1427 242.672
R12779 gnd.n4425 gnd.n1428 242.672
R12780 gnd.n4425 gnd.n1429 242.672
R12781 gnd.n4425 gnd.n1430 242.672
R12782 gnd.n4425 gnd.n1431 242.672
R12783 gnd.n4425 gnd.n1432 242.672
R12784 gnd.n4425 gnd.n1433 242.672
R12785 gnd.n4425 gnd.n1434 242.672
R12786 gnd.n4425 gnd.n1435 242.672
R12787 gnd.n176 gnd.n106 242.672
R12788 gnd.n7392 gnd.n106 242.672
R12789 gnd.n172 gnd.n106 242.672
R12790 gnd.n7399 gnd.n106 242.672
R12791 gnd.n165 gnd.n106 242.672
R12792 gnd.n7406 gnd.n106 242.672
R12793 gnd.n158 gnd.n106 242.672
R12794 gnd.n7413 gnd.n106 242.672
R12795 gnd.n151 gnd.n106 242.672
R12796 gnd.n7420 gnd.n106 242.672
R12797 gnd.n144 gnd.n106 242.672
R12798 gnd.n7430 gnd.n106 242.672
R12799 gnd.n137 gnd.n106 242.672
R12800 gnd.n7437 gnd.n106 242.672
R12801 gnd.n130 gnd.n106 242.672
R12802 gnd.n7444 gnd.n106 242.672
R12803 gnd.n123 gnd.n106 242.672
R12804 gnd.n7451 gnd.n106 242.672
R12805 gnd.n116 gnd.n106 242.672
R12806 gnd.n3720 gnd.n3719 242.672
R12807 gnd.n3720 gnd.n2166 242.672
R12808 gnd.n3720 gnd.n2167 242.672
R12809 gnd.n3720 gnd.n2168 242.672
R12810 gnd.n3720 gnd.n2169 242.672
R12811 gnd.n3720 gnd.n2170 242.672
R12812 gnd.n3720 gnd.n2171 242.672
R12813 gnd.n3720 gnd.n2172 242.672
R12814 gnd.n3720 gnd.n2173 242.672
R12815 gnd.n3720 gnd.n2174 242.672
R12816 gnd.n3720 gnd.n2175 242.672
R12817 gnd.n3720 gnd.n2176 242.672
R12818 gnd.n3720 gnd.n2177 242.672
R12819 gnd.n3721 gnd.n3720 242.672
R12820 gnd.n4134 gnd.n1409 242.672
R12821 gnd.n1817 gnd.n1409 242.672
R12822 gnd.n1814 gnd.n1409 242.672
R12823 gnd.n1809 gnd.n1409 242.672
R12824 gnd.n1806 gnd.n1409 242.672
R12825 gnd.n1686 gnd.n1409 242.672
R12826 gnd.n1792 gnd.n1409 242.672
R12827 gnd.n1698 gnd.n1409 242.672
R12828 gnd.n1776 gnd.n1409 242.672
R12829 gnd.n1704 gnd.n1409 242.672
R12830 gnd.n1757 gnd.n1409 242.672
R12831 gnd.n1711 gnd.n1409 242.672
R12832 gnd.n1738 gnd.n1409 242.672
R12833 gnd.n1718 gnd.n1409 242.672
R12834 gnd.n113 gnd.n109 240.244
R12835 gnd.n7453 gnd.n7452 240.244
R12836 gnd.n7450 gnd.n117 240.244
R12837 gnd.n7446 gnd.n7445 240.244
R12838 gnd.n7443 gnd.n124 240.244
R12839 gnd.n7439 gnd.n7438 240.244
R12840 gnd.n7436 gnd.n131 240.244
R12841 gnd.n7432 gnd.n7431 240.244
R12842 gnd.n7429 gnd.n138 240.244
R12843 gnd.n7422 gnd.n7421 240.244
R12844 gnd.n7419 gnd.n145 240.244
R12845 gnd.n7415 gnd.n7414 240.244
R12846 gnd.n7412 gnd.n152 240.244
R12847 gnd.n7408 gnd.n7407 240.244
R12848 gnd.n7405 gnd.n159 240.244
R12849 gnd.n7401 gnd.n7400 240.244
R12850 gnd.n7398 gnd.n166 240.244
R12851 gnd.n7394 gnd.n7393 240.244
R12852 gnd.n7391 gnd.n173 240.244
R12853 gnd.n4350 gnd.n1495 240.244
R12854 gnd.n1679 gnd.n1495 240.244
R12855 gnd.n1679 gnd.n1626 240.244
R12856 gnd.n1675 gnd.n1626 240.244
R12857 gnd.n1675 gnd.n1616 240.244
R12858 gnd.n1672 gnd.n1616 240.244
R12859 gnd.n1672 gnd.n1608 240.244
R12860 gnd.n1608 gnd.n1598 240.244
R12861 gnd.n1667 gnd.n1598 240.244
R12862 gnd.n1667 gnd.n1589 240.244
R12863 gnd.n1664 gnd.n1589 240.244
R12864 gnd.n1664 gnd.n1581 240.244
R12865 gnd.n1581 gnd.n1571 240.244
R12866 gnd.n1571 gnd.n1559 240.244
R12867 gnd.n4254 gnd.n1559 240.244
R12868 gnd.n4254 gnd.n1560 240.244
R12869 gnd.n1560 gnd.n1547 240.244
R12870 gnd.n1547 gnd.n1536 240.244
R12871 gnd.n4261 gnd.n1536 240.244
R12872 gnd.n4261 gnd.n1527 240.244
R12873 gnd.n4275 gnd.n1527 240.244
R12874 gnd.n4275 gnd.n279 240.244
R12875 gnd.n313 gnd.n279 240.244
R12876 gnd.n4270 gnd.n313 240.244
R12877 gnd.n4270 gnd.n301 240.244
R12878 gnd.n7133 gnd.n301 240.244
R12879 gnd.n7133 gnd.n298 240.244
R12880 gnd.n7197 gnd.n298 240.244
R12881 gnd.n7197 gnd.n295 240.244
R12882 gnd.n7193 gnd.n295 240.244
R12883 gnd.n7193 gnd.n264 240.244
R12884 gnd.n7188 gnd.n264 240.244
R12885 gnd.n7188 gnd.n257 240.244
R12886 gnd.n7184 gnd.n257 240.244
R12887 gnd.n7184 gnd.n249 240.244
R12888 gnd.n7181 gnd.n249 240.244
R12889 gnd.n7181 gnd.n239 240.244
R12890 gnd.n7178 gnd.n239 240.244
R12891 gnd.n7178 gnd.n232 240.244
R12892 gnd.n7175 gnd.n232 240.244
R12893 gnd.n7175 gnd.n226 240.244
R12894 gnd.n7172 gnd.n226 240.244
R12895 gnd.n7172 gnd.n219 240.244
R12896 gnd.n7169 gnd.n219 240.244
R12897 gnd.n7169 gnd.n209 240.244
R12898 gnd.n7166 gnd.n209 240.244
R12899 gnd.n7166 gnd.n202 240.244
R12900 gnd.n7163 gnd.n202 240.244
R12901 gnd.n7163 gnd.n194 240.244
R12902 gnd.n194 gnd.n183 240.244
R12903 gnd.n7382 gnd.n183 240.244
R12904 gnd.n7383 gnd.n7382 240.244
R12905 gnd.n7383 gnd.n105 240.244
R12906 gnd.n1448 gnd.n1447 240.244
R12907 gnd.n4418 gnd.n1447 240.244
R12908 gnd.n4416 gnd.n4415 240.244
R12909 gnd.n4412 gnd.n4411 240.244
R12910 gnd.n4408 gnd.n4407 240.244
R12911 gnd.n4404 gnd.n4403 240.244
R12912 gnd.n4400 gnd.n4399 240.244
R12913 gnd.n4396 gnd.n4395 240.244
R12914 gnd.n4391 gnd.n4390 240.244
R12915 gnd.n4387 gnd.n4386 240.244
R12916 gnd.n4383 gnd.n4382 240.244
R12917 gnd.n4379 gnd.n4378 240.244
R12918 gnd.n4375 gnd.n4374 240.244
R12919 gnd.n4371 gnd.n4370 240.244
R12920 gnd.n4367 gnd.n4366 240.244
R12921 gnd.n4363 gnd.n4362 240.244
R12922 gnd.n4359 gnd.n4358 240.244
R12923 gnd.n1490 gnd.n1489 240.244
R12924 gnd.n1646 gnd.n1449 240.244
R12925 gnd.n1646 gnd.n1624 240.244
R12926 gnd.n4176 gnd.n1624 240.244
R12927 gnd.n4176 gnd.n1619 240.244
R12928 gnd.n4184 gnd.n1619 240.244
R12929 gnd.n4184 gnd.n1620 240.244
R12930 gnd.n1620 gnd.n1596 240.244
R12931 gnd.n4207 gnd.n1596 240.244
R12932 gnd.n4207 gnd.n1591 240.244
R12933 gnd.n4215 gnd.n1591 240.244
R12934 gnd.n4215 gnd.n1592 240.244
R12935 gnd.n1592 gnd.n1569 240.244
R12936 gnd.n4244 gnd.n1569 240.244
R12937 gnd.n4244 gnd.n1564 240.244
R12938 gnd.n4252 gnd.n1564 240.244
R12939 gnd.n4252 gnd.n1565 240.244
R12940 gnd.n1565 gnd.n1534 240.244
R12941 gnd.n4307 gnd.n1534 240.244
R12942 gnd.n4307 gnd.n1530 240.244
R12943 gnd.n4313 gnd.n1530 240.244
R12944 gnd.n4313 gnd.n276 240.244
R12945 gnd.n7220 gnd.n276 240.244
R12946 gnd.n7220 gnd.n277 240.244
R12947 gnd.n305 gnd.n277 240.244
R12948 gnd.n7128 gnd.n305 240.244
R12949 gnd.n7131 gnd.n7128 240.244
R12950 gnd.n7131 gnd.n297 240.244
R12951 gnd.n7199 gnd.n297 240.244
R12952 gnd.n7202 gnd.n7199 240.244
R12953 gnd.n7202 gnd.n266 240.244
R12954 gnd.n7225 gnd.n266 240.244
R12955 gnd.n7225 gnd.n255 240.244
R12956 gnd.n7235 gnd.n255 240.244
R12957 gnd.n7235 gnd.n251 240.244
R12958 gnd.n7241 gnd.n251 240.244
R12959 gnd.n7241 gnd.n237 240.244
R12960 gnd.n7251 gnd.n237 240.244
R12961 gnd.n7251 gnd.n233 240.244
R12962 gnd.n7257 gnd.n233 240.244
R12963 gnd.n7257 gnd.n224 240.244
R12964 gnd.n7267 gnd.n224 240.244
R12965 gnd.n7267 gnd.n220 240.244
R12966 gnd.n7273 gnd.n220 240.244
R12967 gnd.n7273 gnd.n207 240.244
R12968 gnd.n7283 gnd.n207 240.244
R12969 gnd.n7283 gnd.n203 240.244
R12970 gnd.n7289 gnd.n203 240.244
R12971 gnd.n7289 gnd.n192 240.244
R12972 gnd.n7374 gnd.n192 240.244
R12973 gnd.n7374 gnd.n188 240.244
R12974 gnd.n7380 gnd.n188 240.244
R12975 gnd.n7380 gnd.n108 240.244
R12976 gnd.n7460 gnd.n108 240.244
R12977 gnd.n2269 gnd.n1269 240.244
R12978 gnd.n3668 gnd.n2270 240.244
R12979 gnd.n3664 gnd.n3663 240.244
R12980 gnd.n3660 gnd.n3659 240.244
R12981 gnd.n3656 gnd.n3655 240.244
R12982 gnd.n3652 gnd.n3651 240.244
R12983 gnd.n3648 gnd.n3647 240.244
R12984 gnd.n3644 gnd.n3643 240.244
R12985 gnd.n2865 gnd.n2864 240.244
R12986 gnd.n2862 gnd.n2861 240.244
R12987 gnd.n2858 gnd.n2857 240.244
R12988 gnd.n2854 gnd.n2853 240.244
R12989 gnd.n2850 gnd.n2849 240.244
R12990 gnd.n2846 gnd.n2845 240.244
R12991 gnd.n2842 gnd.n2841 240.244
R12992 gnd.n2838 gnd.n2837 240.244
R12993 gnd.n2834 gnd.n2833 240.244
R12994 gnd.n2830 gnd.n2829 240.244
R12995 gnd.n4753 gnd.n1009 240.244
R12996 gnd.n1013 gnd.n1009 240.244
R12997 gnd.n4746 gnd.n1013 240.244
R12998 gnd.n4746 gnd.n1014 240.244
R12999 gnd.n1027 gnd.n1014 240.244
R13000 gnd.n2416 gnd.n1027 240.244
R13001 gnd.n2416 gnd.n1038 240.244
R13002 gnd.n2421 gnd.n1038 240.244
R13003 gnd.n2421 gnd.n1048 240.244
R13004 gnd.n2424 gnd.n1048 240.244
R13005 gnd.n2424 gnd.n1058 240.244
R13006 gnd.n2429 gnd.n1058 240.244
R13007 gnd.n2429 gnd.n1068 240.244
R13008 gnd.n2432 gnd.n1068 240.244
R13009 gnd.n2432 gnd.n1078 240.244
R13010 gnd.n2437 gnd.n1078 240.244
R13011 gnd.n2437 gnd.n1088 240.244
R13012 gnd.n2440 gnd.n1088 240.244
R13013 gnd.n2440 gnd.n1099 240.244
R13014 gnd.n2578 gnd.n1099 240.244
R13015 gnd.n2578 gnd.n1110 240.244
R13016 gnd.n2399 gnd.n1110 240.244
R13017 gnd.n2399 gnd.n1120 240.244
R13018 gnd.n2626 gnd.n1120 240.244
R13019 gnd.n2626 gnd.n1129 240.244
R13020 gnd.n2622 gnd.n1129 240.244
R13021 gnd.n2622 gnd.n1139 240.244
R13022 gnd.n2611 gnd.n1139 240.244
R13023 gnd.n2611 gnd.n1147 240.244
R13024 gnd.n2363 gnd.n1147 240.244
R13025 gnd.n2363 gnd.n1157 240.244
R13026 gnd.n2653 gnd.n1157 240.244
R13027 gnd.n2653 gnd.n1167 240.244
R13028 gnd.n2660 gnd.n1167 240.244
R13029 gnd.n2660 gnd.n1177 240.244
R13030 gnd.n2670 gnd.n1177 240.244
R13031 gnd.n2670 gnd.n1188 240.244
R13032 gnd.n2339 gnd.n1188 240.244
R13033 gnd.n2339 gnd.n1198 240.244
R13034 gnd.n2678 gnd.n1198 240.244
R13035 gnd.n2678 gnd.n1209 240.244
R13036 gnd.n2683 gnd.n1209 240.244
R13037 gnd.n2683 gnd.n1219 240.244
R13038 gnd.n2693 gnd.n1219 240.244
R13039 gnd.n2693 gnd.n1230 240.244
R13040 gnd.n2327 gnd.n1230 240.244
R13041 gnd.n2327 gnd.n1240 240.244
R13042 gnd.n2773 gnd.n1240 240.244
R13043 gnd.n2773 gnd.n1251 240.244
R13044 gnd.n2780 gnd.n1251 240.244
R13045 gnd.n2780 gnd.n1262 240.244
R13046 gnd.n2822 gnd.n1262 240.244
R13047 gnd.n2822 gnd.n1271 240.244
R13048 gnd.n963 gnd.n962 240.244
R13049 gnd.n4825 gnd.n962 240.244
R13050 gnd.n4823 gnd.n4822 240.244
R13051 gnd.n4819 gnd.n4818 240.244
R13052 gnd.n4815 gnd.n4814 240.244
R13053 gnd.n4811 gnd.n4810 240.244
R13054 gnd.n4807 gnd.n4806 240.244
R13055 gnd.n4803 gnd.n4802 240.244
R13056 gnd.n4799 gnd.n4798 240.244
R13057 gnd.n4794 gnd.n4793 240.244
R13058 gnd.n4790 gnd.n4789 240.244
R13059 gnd.n4786 gnd.n4785 240.244
R13060 gnd.n4782 gnd.n4781 240.244
R13061 gnd.n4778 gnd.n4777 240.244
R13062 gnd.n4774 gnd.n4773 240.244
R13063 gnd.n4770 gnd.n4769 240.244
R13064 gnd.n4766 gnd.n4765 240.244
R13065 gnd.n4762 gnd.n4761 240.244
R13066 gnd.n1004 gnd.n1003 240.244
R13067 gnd.n2534 gnd.n964 240.244
R13068 gnd.n2534 gnd.n1019 240.244
R13069 gnd.n4744 gnd.n1019 240.244
R13070 gnd.n4744 gnd.n1020 240.244
R13071 gnd.n4740 gnd.n1020 240.244
R13072 gnd.n4740 gnd.n1026 240.244
R13073 gnd.n4732 gnd.n1026 240.244
R13074 gnd.n4732 gnd.n1041 240.244
R13075 gnd.n4728 gnd.n1041 240.244
R13076 gnd.n4728 gnd.n1047 240.244
R13077 gnd.n4720 gnd.n1047 240.244
R13078 gnd.n4720 gnd.n1060 240.244
R13079 gnd.n4716 gnd.n1060 240.244
R13080 gnd.n4716 gnd.n1066 240.244
R13081 gnd.n4708 gnd.n1066 240.244
R13082 gnd.n4708 gnd.n1081 240.244
R13083 gnd.n4704 gnd.n1081 240.244
R13084 gnd.n4704 gnd.n1087 240.244
R13085 gnd.n4696 gnd.n1087 240.244
R13086 gnd.n4696 gnd.n1102 240.244
R13087 gnd.n4692 gnd.n1102 240.244
R13088 gnd.n4692 gnd.n1108 240.244
R13089 gnd.n4684 gnd.n1108 240.244
R13090 gnd.n4684 gnd.n1123 240.244
R13091 gnd.n4680 gnd.n1123 240.244
R13092 gnd.n4680 gnd.n1127 240.244
R13093 gnd.n4672 gnd.n1127 240.244
R13094 gnd.n4672 gnd.n1142 240.244
R13095 gnd.n4667 gnd.n1142 240.244
R13096 gnd.n4667 gnd.n1145 240.244
R13097 gnd.n4659 gnd.n1145 240.244
R13098 gnd.n4659 gnd.n1160 240.244
R13099 gnd.n4655 gnd.n1160 240.244
R13100 gnd.n4655 gnd.n1165 240.244
R13101 gnd.n4647 gnd.n1165 240.244
R13102 gnd.n4647 gnd.n1180 240.244
R13103 gnd.n4643 gnd.n1180 240.244
R13104 gnd.n4643 gnd.n1186 240.244
R13105 gnd.n4635 gnd.n1186 240.244
R13106 gnd.n4635 gnd.n1201 240.244
R13107 gnd.n4631 gnd.n1201 240.244
R13108 gnd.n4631 gnd.n1207 240.244
R13109 gnd.n4623 gnd.n1207 240.244
R13110 gnd.n4623 gnd.n1222 240.244
R13111 gnd.n4619 gnd.n1222 240.244
R13112 gnd.n4619 gnd.n1228 240.244
R13113 gnd.n4611 gnd.n1228 240.244
R13114 gnd.n4611 gnd.n1243 240.244
R13115 gnd.n4607 gnd.n1243 240.244
R13116 gnd.n4607 gnd.n1249 240.244
R13117 gnd.n4599 gnd.n1249 240.244
R13118 gnd.n4599 gnd.n1264 240.244
R13119 gnd.n4595 gnd.n1264 240.244
R13120 gnd.n4840 gnd.n4835 240.244
R13121 gnd.n6228 gnd.n6227 240.244
R13122 gnd.n6225 gnd.n4844 240.244
R13123 gnd.n6221 gnd.n6220 240.244
R13124 gnd.n6218 gnd.n4851 240.244
R13125 gnd.n6214 gnd.n6213 240.244
R13126 gnd.n6211 gnd.n4858 240.244
R13127 gnd.n6207 gnd.n6206 240.244
R13128 gnd.n5521 gnd.n5147 240.244
R13129 gnd.n5531 gnd.n5147 240.244
R13130 gnd.n5531 gnd.n5138 240.244
R13131 gnd.n5138 gnd.n5127 240.244
R13132 gnd.n5552 gnd.n5127 240.244
R13133 gnd.n5552 gnd.n5121 240.244
R13134 gnd.n5562 gnd.n5121 240.244
R13135 gnd.n5562 gnd.n5112 240.244
R13136 gnd.n5112 gnd.n5103 240.244
R13137 gnd.n5583 gnd.n5103 240.244
R13138 gnd.n5583 gnd.n5096 240.244
R13139 gnd.n5593 gnd.n5096 240.244
R13140 gnd.n5593 gnd.n5087 240.244
R13141 gnd.n5087 gnd.n5077 240.244
R13142 gnd.n5614 gnd.n5077 240.244
R13143 gnd.n5614 gnd.n5070 240.244
R13144 gnd.n5624 gnd.n5070 240.244
R13145 gnd.n5624 gnd.n5061 240.244
R13146 gnd.n5061 gnd.n5052 240.244
R13147 gnd.n5645 gnd.n5052 240.244
R13148 gnd.n5645 gnd.n5045 240.244
R13149 gnd.n5655 gnd.n5045 240.244
R13150 gnd.n5655 gnd.n5037 240.244
R13151 gnd.n5037 gnd.n5028 240.244
R13152 gnd.n5675 gnd.n5028 240.244
R13153 gnd.n5675 gnd.n5015 240.244
R13154 gnd.n5709 gnd.n5015 240.244
R13155 gnd.n5709 gnd.n5005 240.244
R13156 gnd.n5005 gnd.n4997 240.244
R13157 gnd.n5727 gnd.n4997 240.244
R13158 gnd.n5728 gnd.n5727 240.244
R13159 gnd.n5728 gnd.n4985 240.244
R13160 gnd.n4985 gnd.n4974 240.244
R13161 gnd.n5759 gnd.n4974 240.244
R13162 gnd.n5760 gnd.n5759 240.244
R13163 gnd.n5763 gnd.n5760 240.244
R13164 gnd.n5763 gnd.n4960 240.244
R13165 gnd.n5791 gnd.n4960 240.244
R13166 gnd.n5791 gnd.n4947 240.244
R13167 gnd.n5813 gnd.n4947 240.244
R13168 gnd.n5814 gnd.n5813 240.244
R13169 gnd.n5814 gnd.n4931 240.244
R13170 gnd.n5824 gnd.n4931 240.244
R13171 gnd.n5824 gnd.n4923 240.244
R13172 gnd.n6106 gnd.n4923 240.244
R13173 gnd.n6106 gnd.n6105 240.244
R13174 gnd.n6105 gnd.n6104 240.244
R13175 gnd.n6104 gnd.n909 240.244
R13176 gnd.n6100 gnd.n909 240.244
R13177 gnd.n6100 gnd.n920 240.244
R13178 gnd.n6096 gnd.n920 240.244
R13179 gnd.n6096 gnd.n6095 240.244
R13180 gnd.n6095 gnd.n932 240.244
R13181 gnd.n5511 gnd.n5160 240.244
R13182 gnd.n5181 gnd.n5160 240.244
R13183 gnd.n5184 gnd.n5183 240.244
R13184 gnd.n5191 gnd.n5190 240.244
R13185 gnd.n5194 gnd.n5193 240.244
R13186 gnd.n5201 gnd.n5200 240.244
R13187 gnd.n5204 gnd.n5203 240.244
R13188 gnd.n5211 gnd.n5210 240.244
R13189 gnd.n5519 gnd.n5157 240.244
R13190 gnd.n5157 gnd.n5136 240.244
R13191 gnd.n5542 gnd.n5136 240.244
R13192 gnd.n5542 gnd.n5130 240.244
R13193 gnd.n5550 gnd.n5130 240.244
R13194 gnd.n5550 gnd.n5132 240.244
R13195 gnd.n5132 gnd.n5110 240.244
R13196 gnd.n5573 gnd.n5110 240.244
R13197 gnd.n5573 gnd.n5105 240.244
R13198 gnd.n5581 gnd.n5105 240.244
R13199 gnd.n5581 gnd.n5106 240.244
R13200 gnd.n5106 gnd.n5085 240.244
R13201 gnd.n5604 gnd.n5085 240.244
R13202 gnd.n5604 gnd.n5080 240.244
R13203 gnd.n5612 gnd.n5080 240.244
R13204 gnd.n5612 gnd.n5081 240.244
R13205 gnd.n5081 gnd.n5059 240.244
R13206 gnd.n5635 gnd.n5059 240.244
R13207 gnd.n5635 gnd.n5054 240.244
R13208 gnd.n5643 gnd.n5054 240.244
R13209 gnd.n5643 gnd.n5055 240.244
R13210 gnd.n5055 gnd.n5035 240.244
R13211 gnd.n5665 gnd.n5035 240.244
R13212 gnd.n5665 gnd.n5030 240.244
R13213 gnd.n5673 gnd.n5030 240.244
R13214 gnd.n5673 gnd.n5031 240.244
R13215 gnd.n5031 gnd.n5004 240.244
R13216 gnd.n5719 gnd.n5004 240.244
R13217 gnd.n5719 gnd.n5000 240.244
R13218 gnd.n5725 gnd.n5000 240.244
R13219 gnd.n5725 gnd.n4983 240.244
R13220 gnd.n5749 gnd.n4983 240.244
R13221 gnd.n5749 gnd.n4978 240.244
R13222 gnd.n5757 gnd.n4978 240.244
R13223 gnd.n5757 gnd.n4979 240.244
R13224 gnd.n4979 gnd.n4959 240.244
R13225 gnd.n5795 gnd.n4959 240.244
R13226 gnd.n5795 gnd.n4954 240.244
R13227 gnd.n5803 gnd.n4954 240.244
R13228 gnd.n5803 gnd.n4955 240.244
R13229 gnd.n4955 gnd.n4929 240.244
R13230 gnd.n6116 gnd.n4929 240.244
R13231 gnd.n6116 gnd.n4924 240.244
R13232 gnd.n6128 gnd.n4924 240.244
R13233 gnd.n6128 gnd.n4925 240.244
R13234 gnd.n6124 gnd.n4925 240.244
R13235 gnd.n6124 gnd.n911 240.244
R13236 gnd.n6249 gnd.n911 240.244
R13237 gnd.n6249 gnd.n912 240.244
R13238 gnd.n6245 gnd.n912 240.244
R13239 gnd.n6245 gnd.n918 240.244
R13240 gnd.n4834 gnd.n918 240.244
R13241 gnd.n6235 gnd.n4834 240.244
R13242 gnd.n4870 gnd.n929 240.244
R13243 gnd.n6196 gnd.n6195 240.244
R13244 gnd.n6193 gnd.n4874 240.244
R13245 gnd.n6189 gnd.n6188 240.244
R13246 gnd.n6186 gnd.n4881 240.244
R13247 gnd.n6182 gnd.n6181 240.244
R13248 gnd.n6179 gnd.n4888 240.244
R13249 gnd.n6175 gnd.n6174 240.244
R13250 gnd.n6172 gnd.n4895 240.244
R13251 gnd.n6168 gnd.n6167 240.244
R13252 gnd.n6165 gnd.n4902 240.244
R13253 gnd.n6161 gnd.n6160 240.244
R13254 gnd.n6158 gnd.n4912 240.244
R13255 gnd.n5348 gnd.n5245 240.244
R13256 gnd.n5348 gnd.n5238 240.244
R13257 gnd.n5359 gnd.n5238 240.244
R13258 gnd.n5359 gnd.n5234 240.244
R13259 gnd.n5365 gnd.n5234 240.244
R13260 gnd.n5365 gnd.n5226 240.244
R13261 gnd.n5375 gnd.n5226 240.244
R13262 gnd.n5375 gnd.n5221 240.244
R13263 gnd.n5497 gnd.n5221 240.244
R13264 gnd.n5497 gnd.n5222 240.244
R13265 gnd.n5222 gnd.n5169 240.244
R13266 gnd.n5492 gnd.n5169 240.244
R13267 gnd.n5492 gnd.n5491 240.244
R13268 gnd.n5491 gnd.n5148 240.244
R13269 gnd.n5487 gnd.n5148 240.244
R13270 gnd.n5487 gnd.n5139 240.244
R13271 gnd.n5484 gnd.n5139 240.244
R13272 gnd.n5484 gnd.n5483 240.244
R13273 gnd.n5483 gnd.n5122 240.244
R13274 gnd.n5479 gnd.n5122 240.244
R13275 gnd.n5479 gnd.n5113 240.244
R13276 gnd.n5476 gnd.n5113 240.244
R13277 gnd.n5476 gnd.n5475 240.244
R13278 gnd.n5475 gnd.n5098 240.244
R13279 gnd.n5470 gnd.n5098 240.244
R13280 gnd.n5470 gnd.n5088 240.244
R13281 gnd.n5467 gnd.n5088 240.244
R13282 gnd.n5467 gnd.n5466 240.244
R13283 gnd.n5466 gnd.n5072 240.244
R13284 gnd.n5399 gnd.n5072 240.244
R13285 gnd.n5399 gnd.n5062 240.244
R13286 gnd.n5410 gnd.n5062 240.244
R13287 gnd.n5410 gnd.n5408 240.244
R13288 gnd.n5408 gnd.n5047 240.244
R13289 gnd.n5403 gnd.n5047 240.244
R13290 gnd.n5403 gnd.n5038 240.244
R13291 gnd.n5038 gnd.n5021 240.244
R13292 gnd.n5685 gnd.n5021 240.244
R13293 gnd.n5685 gnd.n5017 240.244
R13294 gnd.n5706 gnd.n5017 240.244
R13295 gnd.n5706 gnd.n5006 240.244
R13296 gnd.n5702 gnd.n5006 240.244
R13297 gnd.n5702 gnd.n4996 240.244
R13298 gnd.n5699 gnd.n4996 240.244
R13299 gnd.n5699 gnd.n4986 240.244
R13300 gnd.n5696 gnd.n4986 240.244
R13301 gnd.n5696 gnd.n4965 240.244
R13302 gnd.n5772 gnd.n4965 240.244
R13303 gnd.n5772 gnd.n4961 240.244
R13304 gnd.n5790 gnd.n4961 240.244
R13305 gnd.n5790 gnd.n4952 240.244
R13306 gnd.n5786 gnd.n4952 240.244
R13307 gnd.n5786 gnd.n4946 240.244
R13308 gnd.n5783 gnd.n4946 240.244
R13309 gnd.n5783 gnd.n4932 240.244
R13310 gnd.n4932 gnd.n4922 240.244
R13311 gnd.n6131 gnd.n4922 240.244
R13312 gnd.n6131 gnd.n897 240.244
R13313 gnd.n6137 gnd.n897 240.244
R13314 gnd.n6137 gnd.n908 240.244
R13315 gnd.n6141 gnd.n908 240.244
R13316 gnd.n6141 gnd.n6140 240.244
R13317 gnd.n6140 gnd.n921 240.244
R13318 gnd.n6148 gnd.n921 240.244
R13319 gnd.n6148 gnd.n931 240.244
R13320 gnd.n5262 gnd.n5261 240.244
R13321 gnd.n5333 gnd.n5261 240.244
R13322 gnd.n5331 gnd.n5330 240.244
R13323 gnd.n5327 gnd.n5326 240.244
R13324 gnd.n5323 gnd.n5322 240.244
R13325 gnd.n5319 gnd.n5318 240.244
R13326 gnd.n5315 gnd.n5314 240.244
R13327 gnd.n5311 gnd.n5310 240.244
R13328 gnd.n5307 gnd.n5306 240.244
R13329 gnd.n5303 gnd.n5302 240.244
R13330 gnd.n5299 gnd.n5298 240.244
R13331 gnd.n5295 gnd.n5294 240.244
R13332 gnd.n5291 gnd.n5249 240.244
R13333 gnd.n5351 gnd.n5243 240.244
R13334 gnd.n5351 gnd.n5239 240.244
R13335 gnd.n5357 gnd.n5239 240.244
R13336 gnd.n5357 gnd.n5232 240.244
R13337 gnd.n5367 gnd.n5232 240.244
R13338 gnd.n5367 gnd.n5228 240.244
R13339 gnd.n5373 gnd.n5228 240.244
R13340 gnd.n5373 gnd.n5219 240.244
R13341 gnd.n5499 gnd.n5219 240.244
R13342 gnd.n5499 gnd.n5170 240.244
R13343 gnd.n5507 gnd.n5170 240.244
R13344 gnd.n5507 gnd.n5171 240.244
R13345 gnd.n5171 gnd.n5149 240.244
R13346 gnd.n5528 gnd.n5149 240.244
R13347 gnd.n5528 gnd.n5141 240.244
R13348 gnd.n5539 gnd.n5141 240.244
R13349 gnd.n5539 gnd.n5142 240.244
R13350 gnd.n5142 gnd.n5123 240.244
R13351 gnd.n5559 gnd.n5123 240.244
R13352 gnd.n5559 gnd.n5115 240.244
R13353 gnd.n5570 gnd.n5115 240.244
R13354 gnd.n5570 gnd.n5116 240.244
R13355 gnd.n5116 gnd.n5099 240.244
R13356 gnd.n5590 gnd.n5099 240.244
R13357 gnd.n5590 gnd.n5090 240.244
R13358 gnd.n5601 gnd.n5090 240.244
R13359 gnd.n5601 gnd.n5091 240.244
R13360 gnd.n5091 gnd.n5073 240.244
R13361 gnd.n5621 gnd.n5073 240.244
R13362 gnd.n5621 gnd.n5064 240.244
R13363 gnd.n5632 gnd.n5064 240.244
R13364 gnd.n5632 gnd.n5065 240.244
R13365 gnd.n5065 gnd.n5048 240.244
R13366 gnd.n5652 gnd.n5048 240.244
R13367 gnd.n5652 gnd.n5040 240.244
R13368 gnd.n5662 gnd.n5040 240.244
R13369 gnd.n5662 gnd.n5023 240.244
R13370 gnd.n5683 gnd.n5023 240.244
R13371 gnd.n5683 gnd.n5024 240.244
R13372 gnd.n5024 gnd.n5008 240.244
R13373 gnd.n5716 gnd.n5008 240.244
R13374 gnd.n5716 gnd.n4995 240.244
R13375 gnd.n5731 gnd.n4995 240.244
R13376 gnd.n5731 gnd.n4988 240.244
R13377 gnd.n5746 gnd.n4988 240.244
R13378 gnd.n5746 gnd.n4989 240.244
R13379 gnd.n4989 gnd.n4967 240.244
R13380 gnd.n5770 gnd.n4967 240.244
R13381 gnd.n5770 gnd.n4968 240.244
R13382 gnd.n4968 gnd.n4951 240.244
R13383 gnd.n5806 gnd.n4951 240.244
R13384 gnd.n5806 gnd.n4944 240.244
R13385 gnd.n5817 gnd.n4944 240.244
R13386 gnd.n5817 gnd.n4934 240.244
R13387 gnd.n6113 gnd.n4934 240.244
R13388 gnd.n6113 gnd.n4936 240.244
R13389 gnd.n4936 gnd.n899 240.244
R13390 gnd.n6256 gnd.n899 240.244
R13391 gnd.n6256 gnd.n900 240.244
R13392 gnd.n6252 gnd.n900 240.244
R13393 gnd.n6252 gnd.n906 240.244
R13394 gnd.n923 gnd.n906 240.244
R13395 gnd.n6242 gnd.n923 240.244
R13396 gnd.n6242 gnd.n924 240.244
R13397 gnd.n6238 gnd.n924 240.244
R13398 gnd.n7299 gnd.n7298 240.244
R13399 gnd.n7304 gnd.n7301 240.244
R13400 gnd.n7307 gnd.n7306 240.244
R13401 gnd.n7312 gnd.n7309 240.244
R13402 gnd.n7315 gnd.n7314 240.244
R13403 gnd.n7320 gnd.n7317 240.244
R13404 gnd.n7323 gnd.n7322 240.244
R13405 gnd.n7328 gnd.n7325 240.244
R13406 gnd.n7334 gnd.n7330 240.244
R13407 gnd.n1680 gnd.n1498 240.244
R13408 gnd.n4162 gnd.n1680 240.244
R13409 gnd.n4162 gnd.n1627 240.244
R13410 gnd.n1627 gnd.n1614 240.244
R13411 gnd.n4186 gnd.n1614 240.244
R13412 gnd.n4186 gnd.n1609 240.244
R13413 gnd.n4193 gnd.n1609 240.244
R13414 gnd.n4193 gnd.n1599 240.244
R13415 gnd.n1599 gnd.n1587 240.244
R13416 gnd.n4217 gnd.n1587 240.244
R13417 gnd.n4217 gnd.n1582 240.244
R13418 gnd.n4229 gnd.n1582 240.244
R13419 gnd.n4229 gnd.n1572 240.244
R13420 gnd.n4222 gnd.n1572 240.244
R13421 gnd.n4222 gnd.n1562 240.244
R13422 gnd.n1562 gnd.n1548 240.244
R13423 gnd.n4286 gnd.n1548 240.244
R13424 gnd.n4286 gnd.n1537 240.244
R13425 gnd.n1553 gnd.n1537 240.244
R13426 gnd.n1553 gnd.n1528 240.244
R13427 gnd.n4277 gnd.n1528 240.244
R13428 gnd.n4277 gnd.n280 240.244
R13429 gnd.n7120 gnd.n280 240.244
R13430 gnd.n7120 gnd.n308 240.244
R13431 gnd.n7126 gnd.n308 240.244
R13432 gnd.n7126 gnd.n303 240.244
R13433 gnd.n303 gnd.n70 240.244
R13434 gnd.n71 gnd.n70 240.244
R13435 gnd.n72 gnd.n71 240.244
R13436 gnd.n7191 gnd.n72 240.244
R13437 gnd.n7191 gnd.n75 240.244
R13438 gnd.n76 gnd.n75 240.244
R13439 gnd.n77 gnd.n76 240.244
R13440 gnd.n247 gnd.n77 240.244
R13441 gnd.n247 gnd.n80 240.244
R13442 gnd.n81 gnd.n80 240.244
R13443 gnd.n82 gnd.n81 240.244
R13444 gnd.n240 gnd.n82 240.244
R13445 gnd.n240 gnd.n85 240.244
R13446 gnd.n86 gnd.n85 240.244
R13447 gnd.n87 gnd.n86 240.244
R13448 gnd.n217 gnd.n87 240.244
R13449 gnd.n217 gnd.n90 240.244
R13450 gnd.n91 gnd.n90 240.244
R13451 gnd.n92 gnd.n91 240.244
R13452 gnd.n210 gnd.n92 240.244
R13453 gnd.n210 gnd.n95 240.244
R13454 gnd.n96 gnd.n95 240.244
R13455 gnd.n97 gnd.n96 240.244
R13456 gnd.n184 gnd.n97 240.244
R13457 gnd.n184 gnd.n100 240.244
R13458 gnd.n101 gnd.n100 240.244
R13459 gnd.n7462 gnd.n101 240.244
R13460 gnd.n1728 gnd.n1727 240.244
R13461 gnd.n1731 gnd.n1730 240.244
R13462 gnd.n1747 gnd.n1746 240.244
R13463 gnd.n1750 gnd.n1749 240.244
R13464 gnd.n1766 gnd.n1765 240.244
R13465 gnd.n1769 gnd.n1768 240.244
R13466 gnd.n1784 gnd.n1783 240.244
R13467 gnd.n1695 gnd.n1694 240.244
R13468 gnd.n1690 gnd.n1445 240.244
R13469 gnd.n4348 gnd.n1501 240.244
R13470 gnd.n1505 gnd.n1501 240.244
R13471 gnd.n1506 gnd.n1505 240.244
R13472 gnd.n1507 gnd.n1506 240.244
R13473 gnd.n1618 gnd.n1507 240.244
R13474 gnd.n1618 gnd.n1510 240.244
R13475 gnd.n1511 gnd.n1510 240.244
R13476 gnd.n1512 gnd.n1511 240.244
R13477 gnd.n1600 gnd.n1512 240.244
R13478 gnd.n1600 gnd.n1515 240.244
R13479 gnd.n1516 gnd.n1515 240.244
R13480 gnd.n1517 gnd.n1516 240.244
R13481 gnd.n4242 gnd.n1517 240.244
R13482 gnd.n4242 gnd.n1520 240.244
R13483 gnd.n1521 gnd.n1520 240.244
R13484 gnd.n1522 gnd.n1521 240.244
R13485 gnd.n4287 gnd.n1522 240.244
R13486 gnd.n4287 gnd.n1525 240.244
R13487 gnd.n1526 gnd.n1525 240.244
R13488 gnd.n4315 gnd.n1526 240.244
R13489 gnd.n4315 gnd.n281 240.244
R13490 gnd.n7218 gnd.n281 240.244
R13491 gnd.n7218 gnd.n282 240.244
R13492 gnd.n287 gnd.n282 240.244
R13493 gnd.n288 gnd.n287 240.244
R13494 gnd.n289 gnd.n288 240.244
R13495 gnd.n319 gnd.n289 240.244
R13496 gnd.n319 gnd.n293 240.244
R13497 gnd.n7204 gnd.n293 240.244
R13498 gnd.n7204 gnd.n262 240.244
R13499 gnd.n7227 gnd.n262 240.244
R13500 gnd.n7227 gnd.n258 240.244
R13501 gnd.n7233 gnd.n258 240.244
R13502 gnd.n7233 gnd.n246 240.244
R13503 gnd.n7243 gnd.n246 240.244
R13504 gnd.n7243 gnd.n242 240.244
R13505 gnd.n7249 gnd.n242 240.244
R13506 gnd.n7249 gnd.n231 240.244
R13507 gnd.n7259 gnd.n231 240.244
R13508 gnd.n7259 gnd.n227 240.244
R13509 gnd.n7265 gnd.n227 240.244
R13510 gnd.n7265 gnd.n216 240.244
R13511 gnd.n7275 gnd.n216 240.244
R13512 gnd.n7275 gnd.n212 240.244
R13513 gnd.n7281 gnd.n212 240.244
R13514 gnd.n7281 gnd.n201 240.244
R13515 gnd.n7291 gnd.n201 240.244
R13516 gnd.n7291 gnd.n195 240.244
R13517 gnd.n7372 gnd.n195 240.244
R13518 gnd.n7372 gnd.n196 240.244
R13519 gnd.n196 gnd.n187 240.244
R13520 gnd.n7296 gnd.n187 240.244
R13521 gnd.n7296 gnd.n107 240.244
R13522 gnd.n2236 gnd.n1274 240.244
R13523 gnd.n2237 gnd.n2186 240.244
R13524 gnd.n2240 gnd.n2187 240.244
R13525 gnd.n2196 gnd.n2195 240.244
R13526 gnd.n2242 gnd.n2203 240.244
R13527 gnd.n2245 gnd.n2204 240.244
R13528 gnd.n2214 gnd.n2213 240.244
R13529 gnd.n2247 gnd.n2221 240.244
R13530 gnd.n2233 gnd.n2222 240.244
R13531 gnd.n2536 gnd.n2456 240.244
R13532 gnd.n2537 gnd.n2536 240.244
R13533 gnd.n2537 gnd.n1016 240.244
R13534 gnd.n2542 gnd.n1016 240.244
R13535 gnd.n2542 gnd.n1028 240.244
R13536 gnd.n2545 gnd.n1028 240.244
R13537 gnd.n2545 gnd.n1039 240.244
R13538 gnd.n2550 gnd.n1039 240.244
R13539 gnd.n2550 gnd.n1049 240.244
R13540 gnd.n2553 gnd.n1049 240.244
R13541 gnd.n2553 gnd.n1059 240.244
R13542 gnd.n2558 gnd.n1059 240.244
R13543 gnd.n2558 gnd.n1069 240.244
R13544 gnd.n2561 gnd.n1069 240.244
R13545 gnd.n2561 gnd.n1079 240.244
R13546 gnd.n2566 gnd.n1079 240.244
R13547 gnd.n2566 gnd.n1089 240.244
R13548 gnd.n2569 gnd.n1089 240.244
R13549 gnd.n2569 gnd.n1100 240.244
R13550 gnd.n2576 gnd.n1100 240.244
R13551 gnd.n2576 gnd.n1111 240.244
R13552 gnd.n2632 gnd.n1111 240.244
R13553 gnd.n2632 gnd.n1121 240.244
R13554 gnd.n2628 gnd.n1121 240.244
R13555 gnd.n2628 gnd.n1130 240.244
R13556 gnd.n2620 gnd.n1130 240.244
R13557 gnd.n2620 gnd.n1140 240.244
R13558 gnd.n2613 gnd.n1140 240.244
R13559 gnd.n2613 gnd.n1148 240.244
R13560 gnd.n2645 gnd.n1148 240.244
R13561 gnd.n2645 gnd.n1158 240.244
R13562 gnd.n2651 gnd.n1158 240.244
R13563 gnd.n2651 gnd.n1168 240.244
R13564 gnd.n2662 gnd.n1168 240.244
R13565 gnd.n2662 gnd.n1178 240.244
R13566 gnd.n2668 gnd.n1178 240.244
R13567 gnd.n2668 gnd.n1189 240.244
R13568 gnd.n2707 gnd.n1189 240.244
R13569 gnd.n2707 gnd.n1199 240.244
R13570 gnd.n2344 gnd.n1199 240.244
R13571 gnd.n2344 gnd.n1210 240.244
R13572 gnd.n2345 gnd.n1210 240.244
R13573 gnd.n2345 gnd.n1220 240.244
R13574 gnd.n2695 gnd.n1220 240.244
R13575 gnd.n2695 gnd.n1231 240.244
R13576 gnd.n2765 gnd.n1231 240.244
R13577 gnd.n2765 gnd.n1241 240.244
R13578 gnd.n2771 gnd.n1241 240.244
R13579 gnd.n2771 gnd.n1252 240.244
R13580 gnd.n2782 gnd.n1252 240.244
R13581 gnd.n2782 gnd.n1263 240.244
R13582 gnd.n2820 gnd.n1263 240.244
R13583 gnd.n2820 gnd.n1272 240.244
R13584 gnd.n2516 gnd.n2515 240.244
R13585 gnd.n2512 gnd.n2511 240.244
R13586 gnd.n2508 gnd.n2507 240.244
R13587 gnd.n2504 gnd.n2503 240.244
R13588 gnd.n2500 gnd.n2499 240.244
R13589 gnd.n2496 gnd.n2495 240.244
R13590 gnd.n2492 gnd.n2491 240.244
R13591 gnd.n2488 gnd.n2487 240.244
R13592 gnd.n2476 gnd.n960 240.244
R13593 gnd.n2528 gnd.n2457 240.244
R13594 gnd.n2528 gnd.n2458 240.244
R13595 gnd.n2458 gnd.n1018 240.244
R13596 gnd.n1030 gnd.n1018 240.244
R13597 gnd.n4738 gnd.n1030 240.244
R13598 gnd.n4738 gnd.n1031 240.244
R13599 gnd.n4734 gnd.n1031 240.244
R13600 gnd.n4734 gnd.n1037 240.244
R13601 gnd.n4726 gnd.n1037 240.244
R13602 gnd.n4726 gnd.n1050 240.244
R13603 gnd.n4722 gnd.n1050 240.244
R13604 gnd.n4722 gnd.n1056 240.244
R13605 gnd.n4714 gnd.n1056 240.244
R13606 gnd.n4714 gnd.n1071 240.244
R13607 gnd.n4710 gnd.n1071 240.244
R13608 gnd.n4710 gnd.n1077 240.244
R13609 gnd.n4702 gnd.n1077 240.244
R13610 gnd.n4702 gnd.n1090 240.244
R13611 gnd.n4698 gnd.n1090 240.244
R13612 gnd.n4698 gnd.n1096 240.244
R13613 gnd.n4690 gnd.n1096 240.244
R13614 gnd.n4690 gnd.n1113 240.244
R13615 gnd.n4686 gnd.n1113 240.244
R13616 gnd.n4686 gnd.n1119 240.244
R13617 gnd.n4678 gnd.n1119 240.244
R13618 gnd.n4678 gnd.n1131 240.244
R13619 gnd.n4674 gnd.n1131 240.244
R13620 gnd.n4674 gnd.n1137 240.244
R13621 gnd.n4665 gnd.n1137 240.244
R13622 gnd.n4665 gnd.n1150 240.244
R13623 gnd.n4661 gnd.n1150 240.244
R13624 gnd.n4661 gnd.n1156 240.244
R13625 gnd.n4653 gnd.n1156 240.244
R13626 gnd.n4653 gnd.n1169 240.244
R13627 gnd.n4649 gnd.n1169 240.244
R13628 gnd.n4649 gnd.n1175 240.244
R13629 gnd.n4641 gnd.n1175 240.244
R13630 gnd.n4641 gnd.n1191 240.244
R13631 gnd.n4637 gnd.n1191 240.244
R13632 gnd.n4637 gnd.n1197 240.244
R13633 gnd.n4629 gnd.n1197 240.244
R13634 gnd.n4629 gnd.n1211 240.244
R13635 gnd.n4625 gnd.n1211 240.244
R13636 gnd.n4625 gnd.n1217 240.244
R13637 gnd.n4617 gnd.n1217 240.244
R13638 gnd.n4617 gnd.n1233 240.244
R13639 gnd.n4613 gnd.n1233 240.244
R13640 gnd.n4613 gnd.n1239 240.244
R13641 gnd.n4605 gnd.n1239 240.244
R13642 gnd.n4605 gnd.n1254 240.244
R13643 gnd.n4601 gnd.n1254 240.244
R13644 gnd.n4601 gnd.n1260 240.244
R13645 gnd.n4593 gnd.n1260 240.244
R13646 gnd.n6428 gnd.n724 240.244
R13647 gnd.n6434 gnd.n724 240.244
R13648 gnd.n6434 gnd.n722 240.244
R13649 gnd.n6438 gnd.n722 240.244
R13650 gnd.n6438 gnd.n718 240.244
R13651 gnd.n6444 gnd.n718 240.244
R13652 gnd.n6444 gnd.n716 240.244
R13653 gnd.n6448 gnd.n716 240.244
R13654 gnd.n6448 gnd.n712 240.244
R13655 gnd.n6454 gnd.n712 240.244
R13656 gnd.n6454 gnd.n710 240.244
R13657 gnd.n6458 gnd.n710 240.244
R13658 gnd.n6458 gnd.n706 240.244
R13659 gnd.n6464 gnd.n706 240.244
R13660 gnd.n6464 gnd.n704 240.244
R13661 gnd.n6468 gnd.n704 240.244
R13662 gnd.n6468 gnd.n700 240.244
R13663 gnd.n6474 gnd.n700 240.244
R13664 gnd.n6474 gnd.n698 240.244
R13665 gnd.n6478 gnd.n698 240.244
R13666 gnd.n6478 gnd.n694 240.244
R13667 gnd.n6484 gnd.n694 240.244
R13668 gnd.n6484 gnd.n692 240.244
R13669 gnd.n6488 gnd.n692 240.244
R13670 gnd.n6488 gnd.n688 240.244
R13671 gnd.n6494 gnd.n688 240.244
R13672 gnd.n6494 gnd.n686 240.244
R13673 gnd.n6498 gnd.n686 240.244
R13674 gnd.n6498 gnd.n682 240.244
R13675 gnd.n6504 gnd.n682 240.244
R13676 gnd.n6504 gnd.n680 240.244
R13677 gnd.n6508 gnd.n680 240.244
R13678 gnd.n6508 gnd.n676 240.244
R13679 gnd.n6514 gnd.n676 240.244
R13680 gnd.n6514 gnd.n674 240.244
R13681 gnd.n6518 gnd.n674 240.244
R13682 gnd.n6518 gnd.n670 240.244
R13683 gnd.n6524 gnd.n670 240.244
R13684 gnd.n6524 gnd.n668 240.244
R13685 gnd.n6528 gnd.n668 240.244
R13686 gnd.n6528 gnd.n664 240.244
R13687 gnd.n6534 gnd.n664 240.244
R13688 gnd.n6534 gnd.n662 240.244
R13689 gnd.n6538 gnd.n662 240.244
R13690 gnd.n6538 gnd.n658 240.244
R13691 gnd.n6544 gnd.n658 240.244
R13692 gnd.n6544 gnd.n656 240.244
R13693 gnd.n6548 gnd.n656 240.244
R13694 gnd.n6548 gnd.n652 240.244
R13695 gnd.n6554 gnd.n652 240.244
R13696 gnd.n6554 gnd.n650 240.244
R13697 gnd.n6558 gnd.n650 240.244
R13698 gnd.n6558 gnd.n646 240.244
R13699 gnd.n6564 gnd.n646 240.244
R13700 gnd.n6564 gnd.n644 240.244
R13701 gnd.n6568 gnd.n644 240.244
R13702 gnd.n6568 gnd.n640 240.244
R13703 gnd.n6574 gnd.n640 240.244
R13704 gnd.n6574 gnd.n638 240.244
R13705 gnd.n6578 gnd.n638 240.244
R13706 gnd.n6578 gnd.n634 240.244
R13707 gnd.n6584 gnd.n634 240.244
R13708 gnd.n6584 gnd.n632 240.244
R13709 gnd.n6588 gnd.n632 240.244
R13710 gnd.n6588 gnd.n628 240.244
R13711 gnd.n6594 gnd.n628 240.244
R13712 gnd.n6594 gnd.n626 240.244
R13713 gnd.n6598 gnd.n626 240.244
R13714 gnd.n6598 gnd.n622 240.244
R13715 gnd.n6604 gnd.n622 240.244
R13716 gnd.n6604 gnd.n620 240.244
R13717 gnd.n6608 gnd.n620 240.244
R13718 gnd.n6608 gnd.n616 240.244
R13719 gnd.n6614 gnd.n616 240.244
R13720 gnd.n6614 gnd.n614 240.244
R13721 gnd.n6618 gnd.n614 240.244
R13722 gnd.n6618 gnd.n610 240.244
R13723 gnd.n6624 gnd.n610 240.244
R13724 gnd.n6624 gnd.n608 240.244
R13725 gnd.n6628 gnd.n608 240.244
R13726 gnd.n6628 gnd.n604 240.244
R13727 gnd.n6634 gnd.n604 240.244
R13728 gnd.n6634 gnd.n602 240.244
R13729 gnd.n6638 gnd.n602 240.244
R13730 gnd.n6638 gnd.n598 240.244
R13731 gnd.n6644 gnd.n598 240.244
R13732 gnd.n6644 gnd.n596 240.244
R13733 gnd.n6648 gnd.n596 240.244
R13734 gnd.n6648 gnd.n592 240.244
R13735 gnd.n6654 gnd.n592 240.244
R13736 gnd.n6654 gnd.n590 240.244
R13737 gnd.n6658 gnd.n590 240.244
R13738 gnd.n6658 gnd.n586 240.244
R13739 gnd.n6664 gnd.n586 240.244
R13740 gnd.n6664 gnd.n584 240.244
R13741 gnd.n6668 gnd.n584 240.244
R13742 gnd.n6668 gnd.n580 240.244
R13743 gnd.n6674 gnd.n580 240.244
R13744 gnd.n6674 gnd.n578 240.244
R13745 gnd.n6678 gnd.n578 240.244
R13746 gnd.n6678 gnd.n574 240.244
R13747 gnd.n6684 gnd.n574 240.244
R13748 gnd.n6684 gnd.n572 240.244
R13749 gnd.n6688 gnd.n572 240.244
R13750 gnd.n6688 gnd.n568 240.244
R13751 gnd.n6694 gnd.n568 240.244
R13752 gnd.n6694 gnd.n566 240.244
R13753 gnd.n6698 gnd.n566 240.244
R13754 gnd.n6698 gnd.n562 240.244
R13755 gnd.n6704 gnd.n562 240.244
R13756 gnd.n6704 gnd.n560 240.244
R13757 gnd.n6708 gnd.n560 240.244
R13758 gnd.n6708 gnd.n556 240.244
R13759 gnd.n6714 gnd.n556 240.244
R13760 gnd.n6714 gnd.n554 240.244
R13761 gnd.n6718 gnd.n554 240.244
R13762 gnd.n6718 gnd.n550 240.244
R13763 gnd.n6724 gnd.n550 240.244
R13764 gnd.n6724 gnd.n548 240.244
R13765 gnd.n6728 gnd.n548 240.244
R13766 gnd.n6728 gnd.n544 240.244
R13767 gnd.n6734 gnd.n544 240.244
R13768 gnd.n6734 gnd.n542 240.244
R13769 gnd.n6738 gnd.n542 240.244
R13770 gnd.n6738 gnd.n538 240.244
R13771 gnd.n6744 gnd.n538 240.244
R13772 gnd.n6744 gnd.n536 240.244
R13773 gnd.n6748 gnd.n536 240.244
R13774 gnd.n6748 gnd.n532 240.244
R13775 gnd.n6754 gnd.n532 240.244
R13776 gnd.n6754 gnd.n530 240.244
R13777 gnd.n6758 gnd.n530 240.244
R13778 gnd.n6758 gnd.n526 240.244
R13779 gnd.n6764 gnd.n526 240.244
R13780 gnd.n6764 gnd.n524 240.244
R13781 gnd.n6768 gnd.n524 240.244
R13782 gnd.n6768 gnd.n520 240.244
R13783 gnd.n6774 gnd.n520 240.244
R13784 gnd.n6774 gnd.n518 240.244
R13785 gnd.n6778 gnd.n518 240.244
R13786 gnd.n6778 gnd.n514 240.244
R13787 gnd.n6784 gnd.n514 240.244
R13788 gnd.n6784 gnd.n512 240.244
R13789 gnd.n6788 gnd.n512 240.244
R13790 gnd.n6788 gnd.n508 240.244
R13791 gnd.n6794 gnd.n508 240.244
R13792 gnd.n6794 gnd.n506 240.244
R13793 gnd.n6798 gnd.n506 240.244
R13794 gnd.n6798 gnd.n502 240.244
R13795 gnd.n6804 gnd.n502 240.244
R13796 gnd.n6804 gnd.n500 240.244
R13797 gnd.n6808 gnd.n500 240.244
R13798 gnd.n6808 gnd.n496 240.244
R13799 gnd.n6814 gnd.n496 240.244
R13800 gnd.n6814 gnd.n494 240.244
R13801 gnd.n6818 gnd.n494 240.244
R13802 gnd.n6818 gnd.n490 240.244
R13803 gnd.n6824 gnd.n490 240.244
R13804 gnd.n6824 gnd.n488 240.244
R13805 gnd.n6828 gnd.n488 240.244
R13806 gnd.n6828 gnd.n484 240.244
R13807 gnd.n6834 gnd.n484 240.244
R13808 gnd.n6834 gnd.n482 240.244
R13809 gnd.n6838 gnd.n482 240.244
R13810 gnd.n6838 gnd.n478 240.244
R13811 gnd.n6844 gnd.n478 240.244
R13812 gnd.n6844 gnd.n476 240.244
R13813 gnd.n6848 gnd.n476 240.244
R13814 gnd.n6848 gnd.n472 240.244
R13815 gnd.n6854 gnd.n472 240.244
R13816 gnd.n6854 gnd.n470 240.244
R13817 gnd.n6858 gnd.n470 240.244
R13818 gnd.n6858 gnd.n466 240.244
R13819 gnd.n6864 gnd.n466 240.244
R13820 gnd.n6864 gnd.n464 240.244
R13821 gnd.n6868 gnd.n464 240.244
R13822 gnd.n6868 gnd.n460 240.244
R13823 gnd.n6875 gnd.n460 240.244
R13824 gnd.n6875 gnd.n458 240.244
R13825 gnd.n6879 gnd.n458 240.244
R13826 gnd.n6879 gnd.n455 240.244
R13827 gnd.n6885 gnd.n453 240.244
R13828 gnd.n6889 gnd.n453 240.244
R13829 gnd.n6889 gnd.n449 240.244
R13830 gnd.n6895 gnd.n449 240.244
R13831 gnd.n6895 gnd.n447 240.244
R13832 gnd.n6899 gnd.n447 240.244
R13833 gnd.n6899 gnd.n443 240.244
R13834 gnd.n6905 gnd.n443 240.244
R13835 gnd.n6905 gnd.n441 240.244
R13836 gnd.n6909 gnd.n441 240.244
R13837 gnd.n6909 gnd.n437 240.244
R13838 gnd.n6915 gnd.n437 240.244
R13839 gnd.n6915 gnd.n435 240.244
R13840 gnd.n6919 gnd.n435 240.244
R13841 gnd.n6919 gnd.n431 240.244
R13842 gnd.n6925 gnd.n431 240.244
R13843 gnd.n6925 gnd.n429 240.244
R13844 gnd.n6929 gnd.n429 240.244
R13845 gnd.n6929 gnd.n425 240.244
R13846 gnd.n6935 gnd.n425 240.244
R13847 gnd.n6935 gnd.n423 240.244
R13848 gnd.n6939 gnd.n423 240.244
R13849 gnd.n6939 gnd.n419 240.244
R13850 gnd.n6945 gnd.n419 240.244
R13851 gnd.n6945 gnd.n417 240.244
R13852 gnd.n6949 gnd.n417 240.244
R13853 gnd.n6949 gnd.n413 240.244
R13854 gnd.n6955 gnd.n413 240.244
R13855 gnd.n6955 gnd.n411 240.244
R13856 gnd.n6959 gnd.n411 240.244
R13857 gnd.n6959 gnd.n407 240.244
R13858 gnd.n6965 gnd.n407 240.244
R13859 gnd.n6965 gnd.n405 240.244
R13860 gnd.n6969 gnd.n405 240.244
R13861 gnd.n6969 gnd.n401 240.244
R13862 gnd.n6975 gnd.n401 240.244
R13863 gnd.n6975 gnd.n399 240.244
R13864 gnd.n6979 gnd.n399 240.244
R13865 gnd.n6979 gnd.n395 240.244
R13866 gnd.n6985 gnd.n395 240.244
R13867 gnd.n6985 gnd.n393 240.244
R13868 gnd.n6989 gnd.n393 240.244
R13869 gnd.n6989 gnd.n389 240.244
R13870 gnd.n6995 gnd.n389 240.244
R13871 gnd.n6995 gnd.n387 240.244
R13872 gnd.n6999 gnd.n387 240.244
R13873 gnd.n6999 gnd.n383 240.244
R13874 gnd.n7005 gnd.n383 240.244
R13875 gnd.n7005 gnd.n381 240.244
R13876 gnd.n7009 gnd.n381 240.244
R13877 gnd.n7009 gnd.n377 240.244
R13878 gnd.n7015 gnd.n377 240.244
R13879 gnd.n7015 gnd.n375 240.244
R13880 gnd.n7019 gnd.n375 240.244
R13881 gnd.n7019 gnd.n371 240.244
R13882 gnd.n7025 gnd.n371 240.244
R13883 gnd.n7025 gnd.n369 240.244
R13884 gnd.n7029 gnd.n369 240.244
R13885 gnd.n7029 gnd.n365 240.244
R13886 gnd.n7035 gnd.n365 240.244
R13887 gnd.n7035 gnd.n363 240.244
R13888 gnd.n7039 gnd.n363 240.244
R13889 gnd.n7039 gnd.n359 240.244
R13890 gnd.n7045 gnd.n359 240.244
R13891 gnd.n7045 gnd.n357 240.244
R13892 gnd.n7049 gnd.n357 240.244
R13893 gnd.n7049 gnd.n353 240.244
R13894 gnd.n7055 gnd.n353 240.244
R13895 gnd.n7055 gnd.n351 240.244
R13896 gnd.n7059 gnd.n351 240.244
R13897 gnd.n7059 gnd.n347 240.244
R13898 gnd.n7065 gnd.n347 240.244
R13899 gnd.n7065 gnd.n345 240.244
R13900 gnd.n7069 gnd.n345 240.244
R13901 gnd.n7069 gnd.n341 240.244
R13902 gnd.n7075 gnd.n341 240.244
R13903 gnd.n7075 gnd.n339 240.244
R13904 gnd.n7079 gnd.n339 240.244
R13905 gnd.n7079 gnd.n335 240.244
R13906 gnd.n7085 gnd.n335 240.244
R13907 gnd.n7085 gnd.n333 240.244
R13908 gnd.n7090 gnd.n333 240.244
R13909 gnd.n7090 gnd.n329 240.244
R13910 gnd.n7097 gnd.n329 240.244
R13911 gnd.n2397 gnd.n2396 240.244
R13912 gnd.n2636 gnd.n2397 240.244
R13913 gnd.n2636 gnd.n2635 240.244
R13914 gnd.n2635 gnd.n2398 240.244
R13915 gnd.n2590 gnd.n2398 240.244
R13916 gnd.n2598 gnd.n2590 240.244
R13917 gnd.n2598 gnd.n2595 240.244
R13918 gnd.n2595 gnd.n2594 240.244
R13919 gnd.n2594 gnd.n2591 240.244
R13920 gnd.n2591 gnd.n2364 240.244
R13921 gnd.n2642 gnd.n2364 240.244
R13922 gnd.n2642 gnd.n2365 240.244
R13923 gnd.n2383 gnd.n2365 240.244
R13924 gnd.n2383 gnd.n2382 240.244
R13925 gnd.n2382 gnd.n2381 240.244
R13926 gnd.n2381 gnd.n2370 240.244
R13927 gnd.n2377 gnd.n2370 240.244
R13928 gnd.n2377 gnd.n2337 240.244
R13929 gnd.n2710 gnd.n2337 240.244
R13930 gnd.n2711 gnd.n2710 240.244
R13931 gnd.n2712 gnd.n2711 240.244
R13932 gnd.n2712 gnd.n2333 240.244
R13933 gnd.n2718 gnd.n2333 240.244
R13934 gnd.n2719 gnd.n2718 240.244
R13935 gnd.n2720 gnd.n2719 240.244
R13936 gnd.n2720 gnd.n2328 240.244
R13937 gnd.n2762 gnd.n2328 240.244
R13938 gnd.n2762 gnd.n2329 240.244
R13939 gnd.n2758 gnd.n2329 240.244
R13940 gnd.n2758 gnd.n2757 240.244
R13941 gnd.n2757 gnd.n2756 240.244
R13942 gnd.n2756 gnd.n2728 240.244
R13943 gnd.n2752 gnd.n2728 240.244
R13944 gnd.n2752 gnd.n2751 240.244
R13945 gnd.n2751 gnd.n2750 240.244
R13946 gnd.n2750 gnd.n2734 240.244
R13947 gnd.n2746 gnd.n2734 240.244
R13948 gnd.n2746 gnd.n2744 240.244
R13949 gnd.n2744 gnd.n2743 240.244
R13950 gnd.n2743 gnd.n2158 240.244
R13951 gnd.n3730 gnd.n2158 240.244
R13952 gnd.n3730 gnd.n2154 240.244
R13953 gnd.n3736 gnd.n2154 240.244
R13954 gnd.n3736 gnd.n2144 240.244
R13955 gnd.n3746 gnd.n2144 240.244
R13956 gnd.n3746 gnd.n2140 240.244
R13957 gnd.n3752 gnd.n2140 240.244
R13958 gnd.n3752 gnd.n2132 240.244
R13959 gnd.n3762 gnd.n2132 240.244
R13960 gnd.n3762 gnd.n2128 240.244
R13961 gnd.n3768 gnd.n2128 240.244
R13962 gnd.n3768 gnd.n2119 240.244
R13963 gnd.n3778 gnd.n2119 240.244
R13964 gnd.n3778 gnd.n2115 240.244
R13965 gnd.n3784 gnd.n2115 240.244
R13966 gnd.n3784 gnd.n2106 240.244
R13967 gnd.n3794 gnd.n2106 240.244
R13968 gnd.n3794 gnd.n2102 240.244
R13969 gnd.n3800 gnd.n2102 240.244
R13970 gnd.n3800 gnd.n2092 240.244
R13971 gnd.n3810 gnd.n2092 240.244
R13972 gnd.n3810 gnd.n2088 240.244
R13973 gnd.n3816 gnd.n2088 240.244
R13974 gnd.n3816 gnd.n2080 240.244
R13975 gnd.n3826 gnd.n2080 240.244
R13976 gnd.n3826 gnd.n2076 240.244
R13977 gnd.n3832 gnd.n2076 240.244
R13978 gnd.n3832 gnd.n2065 240.244
R13979 gnd.n3842 gnd.n2065 240.244
R13980 gnd.n3842 gnd.n2061 240.244
R13981 gnd.n3848 gnd.n2061 240.244
R13982 gnd.n3848 gnd.n2050 240.244
R13983 gnd.n3858 gnd.n2050 240.244
R13984 gnd.n3858 gnd.n2046 240.244
R13985 gnd.n3864 gnd.n2046 240.244
R13986 gnd.n3864 gnd.n2037 240.244
R13987 gnd.n3874 gnd.n2037 240.244
R13988 gnd.n3874 gnd.n2033 240.244
R13989 gnd.n3880 gnd.n2033 240.244
R13990 gnd.n3880 gnd.n2022 240.244
R13991 gnd.n3890 gnd.n2022 240.244
R13992 gnd.n3890 gnd.n2018 240.244
R13993 gnd.n3896 gnd.n2018 240.244
R13994 gnd.n3896 gnd.n2007 240.244
R13995 gnd.n3906 gnd.n2007 240.244
R13996 gnd.n3906 gnd.n2003 240.244
R13997 gnd.n3912 gnd.n2003 240.244
R13998 gnd.n3912 gnd.n1994 240.244
R13999 gnd.n3922 gnd.n1994 240.244
R14000 gnd.n3922 gnd.n1990 240.244
R14001 gnd.n3928 gnd.n1990 240.244
R14002 gnd.n3928 gnd.n1980 240.244
R14003 gnd.n3938 gnd.n1980 240.244
R14004 gnd.n3938 gnd.n1976 240.244
R14005 gnd.n3944 gnd.n1976 240.244
R14006 gnd.n3944 gnd.n1965 240.244
R14007 gnd.n3954 gnd.n1965 240.244
R14008 gnd.n3954 gnd.n1961 240.244
R14009 gnd.n3960 gnd.n1961 240.244
R14010 gnd.n3960 gnd.n1952 240.244
R14011 gnd.n3970 gnd.n1952 240.244
R14012 gnd.n3970 gnd.n1948 240.244
R14013 gnd.n3976 gnd.n1948 240.244
R14014 gnd.n3976 gnd.n1937 240.244
R14015 gnd.n3986 gnd.n1937 240.244
R14016 gnd.n3986 gnd.n1933 240.244
R14017 gnd.n3992 gnd.n1933 240.244
R14018 gnd.n3992 gnd.n1924 240.244
R14019 gnd.n4002 gnd.n1924 240.244
R14020 gnd.n4002 gnd.n1920 240.244
R14021 gnd.n4008 gnd.n1920 240.244
R14022 gnd.n4008 gnd.n1910 240.244
R14023 gnd.n4018 gnd.n1910 240.244
R14024 gnd.n4018 gnd.n1906 240.244
R14025 gnd.n4024 gnd.n1906 240.244
R14026 gnd.n4024 gnd.n1895 240.244
R14027 gnd.n4034 gnd.n1895 240.244
R14028 gnd.n4034 gnd.n1891 240.244
R14029 gnd.n4040 gnd.n1891 240.244
R14030 gnd.n4040 gnd.n1883 240.244
R14031 gnd.n4050 gnd.n1883 240.244
R14032 gnd.n4050 gnd.n1879 240.244
R14033 gnd.n4056 gnd.n1879 240.244
R14034 gnd.n4056 gnd.n1870 240.244
R14035 gnd.n4066 gnd.n1870 240.244
R14036 gnd.n4066 gnd.n1866 240.244
R14037 gnd.n4072 gnd.n1866 240.244
R14038 gnd.n4072 gnd.n1857 240.244
R14039 gnd.n4082 gnd.n1857 240.244
R14040 gnd.n4082 gnd.n1853 240.244
R14041 gnd.n4088 gnd.n1853 240.244
R14042 gnd.n4088 gnd.n1843 240.244
R14043 gnd.n4098 gnd.n1843 240.244
R14044 gnd.n4098 gnd.n1839 240.244
R14045 gnd.n4104 gnd.n1839 240.244
R14046 gnd.n4104 gnd.n1830 240.244
R14047 gnd.n4116 gnd.n1830 240.244
R14048 gnd.n4116 gnd.n1825 240.244
R14049 gnd.n4125 gnd.n1825 240.244
R14050 gnd.n4125 gnd.n1826 240.244
R14051 gnd.n1826 gnd.n1407 240.244
R14052 gnd.n4432 gnd.n1407 240.244
R14053 gnd.n4432 gnd.n1410 240.244
R14054 gnd.n4428 gnd.n1410 240.244
R14055 gnd.n4428 gnd.n1416 240.244
R14056 gnd.n1634 gnd.n1416 240.244
R14057 gnd.n1640 gnd.n1634 240.244
R14058 gnd.n1641 gnd.n1640 240.244
R14059 gnd.n4165 gnd.n1641 240.244
R14060 gnd.n4165 gnd.n1629 240.244
R14061 gnd.n4173 gnd.n1629 240.244
R14062 gnd.n4173 gnd.n1630 240.244
R14063 gnd.n1630 gnd.n1607 240.244
R14064 gnd.n4196 gnd.n1607 240.244
R14065 gnd.n4196 gnd.n1602 240.244
R14066 gnd.n4204 gnd.n1602 240.244
R14067 gnd.n4204 gnd.n1603 240.244
R14068 gnd.n1603 gnd.n1579 240.244
R14069 gnd.n4232 gnd.n1579 240.244
R14070 gnd.n4232 gnd.n1574 240.244
R14071 gnd.n4240 gnd.n1574 240.244
R14072 gnd.n4240 gnd.n1575 240.244
R14073 gnd.n1575 gnd.n1545 240.244
R14074 gnd.n4290 gnd.n1545 240.244
R14075 gnd.n4290 gnd.n1539 240.244
R14076 gnd.n4304 gnd.n1539 240.244
R14077 gnd.n4304 gnd.n1541 240.244
R14078 gnd.n4300 gnd.n1541 240.244
R14079 gnd.n4300 gnd.n4299 240.244
R14080 gnd.n4299 gnd.n315 240.244
R14081 gnd.n7117 gnd.n315 240.244
R14082 gnd.n7117 gnd.n316 240.244
R14083 gnd.n7112 gnd.n316 240.244
R14084 gnd.n7112 gnd.n7111 240.244
R14085 gnd.n7111 gnd.n322 240.244
R14086 gnd.n7106 gnd.n322 240.244
R14087 gnd.n7106 gnd.n7105 240.244
R14088 gnd.n7105 gnd.n7104 240.244
R14089 gnd.n7104 gnd.n324 240.244
R14090 gnd.n7100 gnd.n324 240.244
R14091 gnd.n7100 gnd.n7099 240.244
R14092 gnd.n6424 gnd.n727 240.244
R14093 gnd.n6424 gnd.n729 240.244
R14094 gnd.n6420 gnd.n729 240.244
R14095 gnd.n6420 gnd.n735 240.244
R14096 gnd.n6416 gnd.n735 240.244
R14097 gnd.n6416 gnd.n737 240.244
R14098 gnd.n6412 gnd.n737 240.244
R14099 gnd.n6412 gnd.n743 240.244
R14100 gnd.n6408 gnd.n743 240.244
R14101 gnd.n6408 gnd.n745 240.244
R14102 gnd.n6404 gnd.n745 240.244
R14103 gnd.n6404 gnd.n751 240.244
R14104 gnd.n6400 gnd.n751 240.244
R14105 gnd.n6400 gnd.n753 240.244
R14106 gnd.n6396 gnd.n753 240.244
R14107 gnd.n6396 gnd.n759 240.244
R14108 gnd.n6392 gnd.n759 240.244
R14109 gnd.n6392 gnd.n761 240.244
R14110 gnd.n6388 gnd.n761 240.244
R14111 gnd.n6388 gnd.n767 240.244
R14112 gnd.n6384 gnd.n767 240.244
R14113 gnd.n6384 gnd.n769 240.244
R14114 gnd.n6380 gnd.n769 240.244
R14115 gnd.n6380 gnd.n775 240.244
R14116 gnd.n6376 gnd.n775 240.244
R14117 gnd.n6376 gnd.n777 240.244
R14118 gnd.n6372 gnd.n777 240.244
R14119 gnd.n6372 gnd.n783 240.244
R14120 gnd.n6368 gnd.n783 240.244
R14121 gnd.n6368 gnd.n785 240.244
R14122 gnd.n6364 gnd.n785 240.244
R14123 gnd.n6364 gnd.n791 240.244
R14124 gnd.n6360 gnd.n791 240.244
R14125 gnd.n6360 gnd.n793 240.244
R14126 gnd.n6356 gnd.n793 240.244
R14127 gnd.n6356 gnd.n799 240.244
R14128 gnd.n6352 gnd.n799 240.244
R14129 gnd.n6352 gnd.n801 240.244
R14130 gnd.n6348 gnd.n801 240.244
R14131 gnd.n6348 gnd.n807 240.244
R14132 gnd.n6344 gnd.n807 240.244
R14133 gnd.n6344 gnd.n809 240.244
R14134 gnd.n6340 gnd.n809 240.244
R14135 gnd.n6340 gnd.n815 240.244
R14136 gnd.n6336 gnd.n815 240.244
R14137 gnd.n6336 gnd.n817 240.244
R14138 gnd.n6332 gnd.n817 240.244
R14139 gnd.n6332 gnd.n823 240.244
R14140 gnd.n6328 gnd.n823 240.244
R14141 gnd.n6328 gnd.n825 240.244
R14142 gnd.n6324 gnd.n825 240.244
R14143 gnd.n6324 gnd.n831 240.244
R14144 gnd.n6320 gnd.n831 240.244
R14145 gnd.n6320 gnd.n833 240.244
R14146 gnd.n6316 gnd.n833 240.244
R14147 gnd.n6316 gnd.n839 240.244
R14148 gnd.n6312 gnd.n839 240.244
R14149 gnd.n6312 gnd.n841 240.244
R14150 gnd.n6308 gnd.n841 240.244
R14151 gnd.n6308 gnd.n847 240.244
R14152 gnd.n6304 gnd.n847 240.244
R14153 gnd.n6304 gnd.n849 240.244
R14154 gnd.n6300 gnd.n849 240.244
R14155 gnd.n6300 gnd.n855 240.244
R14156 gnd.n6296 gnd.n855 240.244
R14157 gnd.n6296 gnd.n857 240.244
R14158 gnd.n6292 gnd.n857 240.244
R14159 gnd.n6292 gnd.n863 240.244
R14160 gnd.n6288 gnd.n863 240.244
R14161 gnd.n6288 gnd.n865 240.244
R14162 gnd.n6284 gnd.n865 240.244
R14163 gnd.n6284 gnd.n871 240.244
R14164 gnd.n6280 gnd.n871 240.244
R14165 gnd.n6280 gnd.n873 240.244
R14166 gnd.n6276 gnd.n873 240.244
R14167 gnd.n6276 gnd.n879 240.244
R14168 gnd.n6272 gnd.n879 240.244
R14169 gnd.n6272 gnd.n881 240.244
R14170 gnd.n6268 gnd.n881 240.244
R14171 gnd.n6268 gnd.n887 240.244
R14172 gnd.n6264 gnd.n887 240.244
R14173 gnd.n6264 gnd.n889 240.244
R14174 gnd.n6260 gnd.n889 240.244
R14175 gnd.n6260 gnd.n895 240.244
R14176 gnd.n1280 gnd.n1279 240.244
R14177 gnd.n1281 gnd.n1280 240.244
R14178 gnd.n2153 gnd.n1281 240.244
R14179 gnd.n2153 gnd.n1284 240.244
R14180 gnd.n1285 gnd.n1284 240.244
R14181 gnd.n1286 gnd.n1285 240.244
R14182 gnd.n2139 gnd.n1286 240.244
R14183 gnd.n2139 gnd.n1289 240.244
R14184 gnd.n1290 gnd.n1289 240.244
R14185 gnd.n1291 gnd.n1290 240.244
R14186 gnd.n2127 gnd.n1291 240.244
R14187 gnd.n2127 gnd.n1294 240.244
R14188 gnd.n1295 gnd.n1294 240.244
R14189 gnd.n1296 gnd.n1295 240.244
R14190 gnd.n2114 gnd.n1296 240.244
R14191 gnd.n2114 gnd.n1299 240.244
R14192 gnd.n1300 gnd.n1299 240.244
R14193 gnd.n1301 gnd.n1300 240.244
R14194 gnd.n2100 gnd.n1301 240.244
R14195 gnd.n2100 gnd.n1304 240.244
R14196 gnd.n1305 gnd.n1304 240.244
R14197 gnd.n1306 gnd.n1305 240.244
R14198 gnd.n2087 gnd.n1306 240.244
R14199 gnd.n2087 gnd.n1309 240.244
R14200 gnd.n1310 gnd.n1309 240.244
R14201 gnd.n1311 gnd.n1310 240.244
R14202 gnd.n2074 gnd.n1311 240.244
R14203 gnd.n2074 gnd.n1314 240.244
R14204 gnd.n1315 gnd.n1314 240.244
R14205 gnd.n1316 gnd.n1315 240.244
R14206 gnd.n2059 gnd.n1316 240.244
R14207 gnd.n2059 gnd.n1319 240.244
R14208 gnd.n1320 gnd.n1319 240.244
R14209 gnd.n1321 gnd.n1320 240.244
R14210 gnd.n2045 gnd.n1321 240.244
R14211 gnd.n2045 gnd.n1324 240.244
R14212 gnd.n1325 gnd.n1324 240.244
R14213 gnd.n1326 gnd.n1325 240.244
R14214 gnd.n2031 gnd.n1326 240.244
R14215 gnd.n2031 gnd.n1329 240.244
R14216 gnd.n1330 gnd.n1329 240.244
R14217 gnd.n1331 gnd.n1330 240.244
R14218 gnd.n2016 gnd.n1331 240.244
R14219 gnd.n2016 gnd.n1334 240.244
R14220 gnd.n1335 gnd.n1334 240.244
R14221 gnd.n1336 gnd.n1335 240.244
R14222 gnd.n2001 gnd.n1336 240.244
R14223 gnd.n2001 gnd.n1339 240.244
R14224 gnd.n1340 gnd.n1339 240.244
R14225 gnd.n1341 gnd.n1340 240.244
R14226 gnd.n1988 gnd.n1341 240.244
R14227 gnd.n1988 gnd.n1344 240.244
R14228 gnd.n1345 gnd.n1344 240.244
R14229 gnd.n1346 gnd.n1345 240.244
R14230 gnd.n1974 gnd.n1346 240.244
R14231 gnd.n1974 gnd.n1349 240.244
R14232 gnd.n1350 gnd.n1349 240.244
R14233 gnd.n1351 gnd.n1350 240.244
R14234 gnd.n1960 gnd.n1351 240.244
R14235 gnd.n1960 gnd.n1354 240.244
R14236 gnd.n1355 gnd.n1354 240.244
R14237 gnd.n1356 gnd.n1355 240.244
R14238 gnd.n1946 gnd.n1356 240.244
R14239 gnd.n1946 gnd.n1359 240.244
R14240 gnd.n1360 gnd.n1359 240.244
R14241 gnd.n1361 gnd.n1360 240.244
R14242 gnd.n1932 gnd.n1361 240.244
R14243 gnd.n1932 gnd.n1364 240.244
R14244 gnd.n1365 gnd.n1364 240.244
R14245 gnd.n1366 gnd.n1365 240.244
R14246 gnd.n1919 gnd.n1366 240.244
R14247 gnd.n1919 gnd.n1369 240.244
R14248 gnd.n1370 gnd.n1369 240.244
R14249 gnd.n1371 gnd.n1370 240.244
R14250 gnd.n1904 gnd.n1371 240.244
R14251 gnd.n1904 gnd.n1374 240.244
R14252 gnd.n1375 gnd.n1374 240.244
R14253 gnd.n1376 gnd.n1375 240.244
R14254 gnd.n1889 gnd.n1376 240.244
R14255 gnd.n1889 gnd.n1379 240.244
R14256 gnd.n1380 gnd.n1379 240.244
R14257 gnd.n1381 gnd.n1380 240.244
R14258 gnd.n1878 gnd.n1381 240.244
R14259 gnd.n1878 gnd.n1384 240.244
R14260 gnd.n1385 gnd.n1384 240.244
R14261 gnd.n1386 gnd.n1385 240.244
R14262 gnd.n1865 gnd.n1386 240.244
R14263 gnd.n1865 gnd.n1389 240.244
R14264 gnd.n1390 gnd.n1389 240.244
R14265 gnd.n1391 gnd.n1390 240.244
R14266 gnd.n1852 gnd.n1391 240.244
R14267 gnd.n1852 gnd.n1394 240.244
R14268 gnd.n1395 gnd.n1394 240.244
R14269 gnd.n1396 gnd.n1395 240.244
R14270 gnd.n1838 gnd.n1396 240.244
R14271 gnd.n1838 gnd.n1399 240.244
R14272 gnd.n1400 gnd.n1399 240.244
R14273 gnd.n1401 gnd.n1400 240.244
R14274 gnd.n1824 gnd.n1401 240.244
R14275 gnd.n1824 gnd.n1404 240.244
R14276 gnd.n4435 gnd.n1404 240.244
R14277 gnd.n2180 gnd.n2179 240.244
R14278 gnd.n2190 gnd.n2179 240.244
R14279 gnd.n2192 gnd.n2191 240.244
R14280 gnd.n2200 gnd.n2199 240.244
R14281 gnd.n2208 gnd.n2207 240.244
R14282 gnd.n2210 gnd.n2209 240.244
R14283 gnd.n2218 gnd.n2217 240.244
R14284 gnd.n2228 gnd.n2227 240.244
R14285 gnd.n2230 gnd.n2229 240.244
R14286 gnd.n2788 gnd.n2787 240.244
R14287 gnd.n2790 gnd.n2789 240.244
R14288 gnd.n2794 gnd.n2793 240.244
R14289 gnd.n2800 gnd.n2795 240.244
R14290 gnd.n2801 gnd.n2164 240.244
R14291 gnd.n3728 gnd.n2160 240.244
R14292 gnd.n3728 gnd.n2151 240.244
R14293 gnd.n3738 gnd.n2151 240.244
R14294 gnd.n3738 gnd.n2147 240.244
R14295 gnd.n3744 gnd.n2147 240.244
R14296 gnd.n3744 gnd.n2138 240.244
R14297 gnd.n3754 gnd.n2138 240.244
R14298 gnd.n3754 gnd.n2134 240.244
R14299 gnd.n3760 gnd.n2134 240.244
R14300 gnd.n3760 gnd.n2125 240.244
R14301 gnd.n3770 gnd.n2125 240.244
R14302 gnd.n3770 gnd.n2121 240.244
R14303 gnd.n3776 gnd.n2121 240.244
R14304 gnd.n3776 gnd.n2112 240.244
R14305 gnd.n3786 gnd.n2112 240.244
R14306 gnd.n3786 gnd.n2108 240.244
R14307 gnd.n3792 gnd.n2108 240.244
R14308 gnd.n3792 gnd.n2098 240.244
R14309 gnd.n3802 gnd.n2098 240.244
R14310 gnd.n3802 gnd.n2094 240.244
R14311 gnd.n3808 gnd.n2094 240.244
R14312 gnd.n3808 gnd.n2085 240.244
R14313 gnd.n3818 gnd.n2085 240.244
R14314 gnd.n3818 gnd.n2081 240.244
R14315 gnd.n3824 gnd.n2081 240.244
R14316 gnd.n3824 gnd.n2072 240.244
R14317 gnd.n3834 gnd.n2072 240.244
R14318 gnd.n3834 gnd.n2068 240.244
R14319 gnd.n3840 gnd.n2068 240.244
R14320 gnd.n3840 gnd.n2057 240.244
R14321 gnd.n3850 gnd.n2057 240.244
R14322 gnd.n3850 gnd.n2053 240.244
R14323 gnd.n3856 gnd.n2053 240.244
R14324 gnd.n3856 gnd.n2043 240.244
R14325 gnd.n3866 gnd.n2043 240.244
R14326 gnd.n3866 gnd.n2039 240.244
R14327 gnd.n3872 gnd.n2039 240.244
R14328 gnd.n3872 gnd.n2030 240.244
R14329 gnd.n3882 gnd.n2030 240.244
R14330 gnd.n3882 gnd.n2026 240.244
R14331 gnd.n3888 gnd.n2026 240.244
R14332 gnd.n3888 gnd.n2014 240.244
R14333 gnd.n3898 gnd.n2014 240.244
R14334 gnd.n3898 gnd.n2010 240.244
R14335 gnd.n3904 gnd.n2010 240.244
R14336 gnd.n3904 gnd.n2000 240.244
R14337 gnd.n3914 gnd.n2000 240.244
R14338 gnd.n3914 gnd.n1996 240.244
R14339 gnd.n3920 gnd.n1996 240.244
R14340 gnd.n3920 gnd.n1986 240.244
R14341 gnd.n3930 gnd.n1986 240.244
R14342 gnd.n3930 gnd.n1982 240.244
R14343 gnd.n3936 gnd.n1982 240.244
R14344 gnd.n3936 gnd.n1972 240.244
R14345 gnd.n3946 gnd.n1972 240.244
R14346 gnd.n3946 gnd.n1968 240.244
R14347 gnd.n3952 gnd.n1968 240.244
R14348 gnd.n3952 gnd.n1958 240.244
R14349 gnd.n3962 gnd.n1958 240.244
R14350 gnd.n3962 gnd.n1954 240.244
R14351 gnd.n3968 gnd.n1954 240.244
R14352 gnd.n3968 gnd.n1944 240.244
R14353 gnd.n3978 gnd.n1944 240.244
R14354 gnd.n3978 gnd.n1940 240.244
R14355 gnd.n3984 gnd.n1940 240.244
R14356 gnd.n3984 gnd.n1930 240.244
R14357 gnd.n3994 gnd.n1930 240.244
R14358 gnd.n3994 gnd.n1926 240.244
R14359 gnd.n4000 gnd.n1926 240.244
R14360 gnd.n4000 gnd.n1917 240.244
R14361 gnd.n4010 gnd.n1917 240.244
R14362 gnd.n4010 gnd.n1913 240.244
R14363 gnd.n4016 gnd.n1913 240.244
R14364 gnd.n4016 gnd.n1902 240.244
R14365 gnd.n4026 gnd.n1902 240.244
R14366 gnd.n4026 gnd.n1898 240.244
R14367 gnd.n4032 gnd.n1898 240.244
R14368 gnd.n4032 gnd.n1888 240.244
R14369 gnd.n4042 gnd.n1888 240.244
R14370 gnd.n4042 gnd.n1884 240.244
R14371 gnd.n4048 gnd.n1884 240.244
R14372 gnd.n4048 gnd.n1876 240.244
R14373 gnd.n4058 gnd.n1876 240.244
R14374 gnd.n4058 gnd.n1872 240.244
R14375 gnd.n4064 gnd.n1872 240.244
R14376 gnd.n4064 gnd.n1863 240.244
R14377 gnd.n4074 gnd.n1863 240.244
R14378 gnd.n4074 gnd.n1859 240.244
R14379 gnd.n4080 gnd.n1859 240.244
R14380 gnd.n4080 gnd.n1850 240.244
R14381 gnd.n4090 gnd.n1850 240.244
R14382 gnd.n4090 gnd.n1846 240.244
R14383 gnd.n4096 gnd.n1846 240.244
R14384 gnd.n4096 gnd.n1837 240.244
R14385 gnd.n4106 gnd.n1837 240.244
R14386 gnd.n4106 gnd.n1832 240.244
R14387 gnd.n4114 gnd.n1832 240.244
R14388 gnd.n4114 gnd.n1822 240.244
R14389 gnd.n4127 gnd.n1822 240.244
R14390 gnd.n4128 gnd.n4127 240.244
R14391 gnd.n4128 gnd.n1408 240.244
R14392 gnd.n1737 gnd.n1736 240.244
R14393 gnd.n1740 gnd.n1739 240.244
R14394 gnd.n1756 gnd.n1755 240.244
R14395 gnd.n1759 gnd.n1758 240.244
R14396 gnd.n1775 gnd.n1774 240.244
R14397 gnd.n1778 gnd.n1777 240.244
R14398 gnd.n1791 gnd.n1790 240.244
R14399 gnd.n1794 gnd.n1793 240.244
R14400 gnd.n1805 gnd.n1804 240.244
R14401 gnd.n1808 gnd.n1807 240.244
R14402 gnd.n1813 gnd.n1810 240.244
R14403 gnd.n1816 gnd.n1815 240.244
R14404 gnd.n4133 gnd.n1818 240.244
R14405 gnd.n4136 gnd.n4135 240.244
R14406 gnd.n2901 gnd.n2900 240.132
R14407 gnd.n3187 gnd.n3186 240.132
R14408 gnd.n6427 gnd.n723 225.874
R14409 gnd.n6435 gnd.n723 225.874
R14410 gnd.n6436 gnd.n6435 225.874
R14411 gnd.n6437 gnd.n6436 225.874
R14412 gnd.n6437 gnd.n717 225.874
R14413 gnd.n6445 gnd.n717 225.874
R14414 gnd.n6446 gnd.n6445 225.874
R14415 gnd.n6447 gnd.n6446 225.874
R14416 gnd.n6447 gnd.n711 225.874
R14417 gnd.n6455 gnd.n711 225.874
R14418 gnd.n6456 gnd.n6455 225.874
R14419 gnd.n6457 gnd.n6456 225.874
R14420 gnd.n6457 gnd.n705 225.874
R14421 gnd.n6465 gnd.n705 225.874
R14422 gnd.n6466 gnd.n6465 225.874
R14423 gnd.n6467 gnd.n6466 225.874
R14424 gnd.n6467 gnd.n699 225.874
R14425 gnd.n6475 gnd.n699 225.874
R14426 gnd.n6476 gnd.n6475 225.874
R14427 gnd.n6477 gnd.n6476 225.874
R14428 gnd.n6477 gnd.n693 225.874
R14429 gnd.n6485 gnd.n693 225.874
R14430 gnd.n6486 gnd.n6485 225.874
R14431 gnd.n6487 gnd.n6486 225.874
R14432 gnd.n6487 gnd.n687 225.874
R14433 gnd.n6495 gnd.n687 225.874
R14434 gnd.n6496 gnd.n6495 225.874
R14435 gnd.n6497 gnd.n6496 225.874
R14436 gnd.n6497 gnd.n681 225.874
R14437 gnd.n6505 gnd.n681 225.874
R14438 gnd.n6506 gnd.n6505 225.874
R14439 gnd.n6507 gnd.n6506 225.874
R14440 gnd.n6507 gnd.n675 225.874
R14441 gnd.n6515 gnd.n675 225.874
R14442 gnd.n6516 gnd.n6515 225.874
R14443 gnd.n6517 gnd.n6516 225.874
R14444 gnd.n6517 gnd.n669 225.874
R14445 gnd.n6525 gnd.n669 225.874
R14446 gnd.n6526 gnd.n6525 225.874
R14447 gnd.n6527 gnd.n6526 225.874
R14448 gnd.n6527 gnd.n663 225.874
R14449 gnd.n6535 gnd.n663 225.874
R14450 gnd.n6536 gnd.n6535 225.874
R14451 gnd.n6537 gnd.n6536 225.874
R14452 gnd.n6537 gnd.n657 225.874
R14453 gnd.n6545 gnd.n657 225.874
R14454 gnd.n6546 gnd.n6545 225.874
R14455 gnd.n6547 gnd.n6546 225.874
R14456 gnd.n6547 gnd.n651 225.874
R14457 gnd.n6555 gnd.n651 225.874
R14458 gnd.n6556 gnd.n6555 225.874
R14459 gnd.n6557 gnd.n6556 225.874
R14460 gnd.n6557 gnd.n645 225.874
R14461 gnd.n6565 gnd.n645 225.874
R14462 gnd.n6566 gnd.n6565 225.874
R14463 gnd.n6567 gnd.n6566 225.874
R14464 gnd.n6567 gnd.n639 225.874
R14465 gnd.n6575 gnd.n639 225.874
R14466 gnd.n6576 gnd.n6575 225.874
R14467 gnd.n6577 gnd.n6576 225.874
R14468 gnd.n6577 gnd.n633 225.874
R14469 gnd.n6585 gnd.n633 225.874
R14470 gnd.n6586 gnd.n6585 225.874
R14471 gnd.n6587 gnd.n6586 225.874
R14472 gnd.n6587 gnd.n627 225.874
R14473 gnd.n6595 gnd.n627 225.874
R14474 gnd.n6596 gnd.n6595 225.874
R14475 gnd.n6597 gnd.n6596 225.874
R14476 gnd.n6597 gnd.n621 225.874
R14477 gnd.n6605 gnd.n621 225.874
R14478 gnd.n6606 gnd.n6605 225.874
R14479 gnd.n6607 gnd.n6606 225.874
R14480 gnd.n6607 gnd.n615 225.874
R14481 gnd.n6615 gnd.n615 225.874
R14482 gnd.n6616 gnd.n6615 225.874
R14483 gnd.n6617 gnd.n6616 225.874
R14484 gnd.n6617 gnd.n609 225.874
R14485 gnd.n6625 gnd.n609 225.874
R14486 gnd.n6626 gnd.n6625 225.874
R14487 gnd.n6627 gnd.n6626 225.874
R14488 gnd.n6627 gnd.n603 225.874
R14489 gnd.n6635 gnd.n603 225.874
R14490 gnd.n6636 gnd.n6635 225.874
R14491 gnd.n6637 gnd.n6636 225.874
R14492 gnd.n6637 gnd.n597 225.874
R14493 gnd.n6645 gnd.n597 225.874
R14494 gnd.n6646 gnd.n6645 225.874
R14495 gnd.n6647 gnd.n6646 225.874
R14496 gnd.n6647 gnd.n591 225.874
R14497 gnd.n6655 gnd.n591 225.874
R14498 gnd.n6656 gnd.n6655 225.874
R14499 gnd.n6657 gnd.n6656 225.874
R14500 gnd.n6657 gnd.n585 225.874
R14501 gnd.n6665 gnd.n585 225.874
R14502 gnd.n6666 gnd.n6665 225.874
R14503 gnd.n6667 gnd.n6666 225.874
R14504 gnd.n6667 gnd.n579 225.874
R14505 gnd.n6675 gnd.n579 225.874
R14506 gnd.n6676 gnd.n6675 225.874
R14507 gnd.n6677 gnd.n6676 225.874
R14508 gnd.n6677 gnd.n573 225.874
R14509 gnd.n6685 gnd.n573 225.874
R14510 gnd.n6686 gnd.n6685 225.874
R14511 gnd.n6687 gnd.n6686 225.874
R14512 gnd.n6687 gnd.n567 225.874
R14513 gnd.n6695 gnd.n567 225.874
R14514 gnd.n6696 gnd.n6695 225.874
R14515 gnd.n6697 gnd.n6696 225.874
R14516 gnd.n6697 gnd.n561 225.874
R14517 gnd.n6705 gnd.n561 225.874
R14518 gnd.n6706 gnd.n6705 225.874
R14519 gnd.n6707 gnd.n6706 225.874
R14520 gnd.n6707 gnd.n555 225.874
R14521 gnd.n6715 gnd.n555 225.874
R14522 gnd.n6716 gnd.n6715 225.874
R14523 gnd.n6717 gnd.n6716 225.874
R14524 gnd.n6717 gnd.n549 225.874
R14525 gnd.n6725 gnd.n549 225.874
R14526 gnd.n6726 gnd.n6725 225.874
R14527 gnd.n6727 gnd.n6726 225.874
R14528 gnd.n6727 gnd.n543 225.874
R14529 gnd.n6735 gnd.n543 225.874
R14530 gnd.n6736 gnd.n6735 225.874
R14531 gnd.n6737 gnd.n6736 225.874
R14532 gnd.n6737 gnd.n537 225.874
R14533 gnd.n6745 gnd.n537 225.874
R14534 gnd.n6746 gnd.n6745 225.874
R14535 gnd.n6747 gnd.n6746 225.874
R14536 gnd.n6747 gnd.n531 225.874
R14537 gnd.n6755 gnd.n531 225.874
R14538 gnd.n6756 gnd.n6755 225.874
R14539 gnd.n6757 gnd.n6756 225.874
R14540 gnd.n6757 gnd.n525 225.874
R14541 gnd.n6765 gnd.n525 225.874
R14542 gnd.n6766 gnd.n6765 225.874
R14543 gnd.n6767 gnd.n6766 225.874
R14544 gnd.n6767 gnd.n519 225.874
R14545 gnd.n6775 gnd.n519 225.874
R14546 gnd.n6776 gnd.n6775 225.874
R14547 gnd.n6777 gnd.n6776 225.874
R14548 gnd.n6777 gnd.n513 225.874
R14549 gnd.n6785 gnd.n513 225.874
R14550 gnd.n6786 gnd.n6785 225.874
R14551 gnd.n6787 gnd.n6786 225.874
R14552 gnd.n6787 gnd.n507 225.874
R14553 gnd.n6795 gnd.n507 225.874
R14554 gnd.n6796 gnd.n6795 225.874
R14555 gnd.n6797 gnd.n6796 225.874
R14556 gnd.n6797 gnd.n501 225.874
R14557 gnd.n6805 gnd.n501 225.874
R14558 gnd.n6806 gnd.n6805 225.874
R14559 gnd.n6807 gnd.n6806 225.874
R14560 gnd.n6807 gnd.n495 225.874
R14561 gnd.n6815 gnd.n495 225.874
R14562 gnd.n6816 gnd.n6815 225.874
R14563 gnd.n6817 gnd.n6816 225.874
R14564 gnd.n6817 gnd.n489 225.874
R14565 gnd.n6825 gnd.n489 225.874
R14566 gnd.n6826 gnd.n6825 225.874
R14567 gnd.n6827 gnd.n6826 225.874
R14568 gnd.n6827 gnd.n483 225.874
R14569 gnd.n6835 gnd.n483 225.874
R14570 gnd.n6836 gnd.n6835 225.874
R14571 gnd.n6837 gnd.n6836 225.874
R14572 gnd.n6837 gnd.n477 225.874
R14573 gnd.n6845 gnd.n477 225.874
R14574 gnd.n6846 gnd.n6845 225.874
R14575 gnd.n6847 gnd.n6846 225.874
R14576 gnd.n6847 gnd.n471 225.874
R14577 gnd.n6855 gnd.n471 225.874
R14578 gnd.n6856 gnd.n6855 225.874
R14579 gnd.n6857 gnd.n6856 225.874
R14580 gnd.n6857 gnd.n465 225.874
R14581 gnd.n6865 gnd.n465 225.874
R14582 gnd.n6866 gnd.n6865 225.874
R14583 gnd.n6867 gnd.n6866 225.874
R14584 gnd.n6867 gnd.n459 225.874
R14585 gnd.n6876 gnd.n459 225.874
R14586 gnd.n6877 gnd.n6876 225.874
R14587 gnd.n6878 gnd.n6877 225.874
R14588 gnd.n6878 gnd.n454 225.874
R14589 gnd.n5286 gnd.t108 224.174
R14590 gnd.n4907 gnd.t70 224.174
R14591 gnd.n1467 gnd.n1424 199.319
R14592 gnd.n1467 gnd.n1425 199.319
R14593 gnd.n2292 gnd.n2262 199.319
R14594 gnd.n2292 gnd.n2261 199.319
R14595 gnd.n2902 gnd.n2899 186.49
R14596 gnd.n3188 gnd.n3185 186.49
R14597 gnd.n6080 gnd.n6079 185
R14598 gnd.n6078 gnd.n6077 185
R14599 gnd.n6057 gnd.n6056 185
R14600 gnd.n6072 gnd.n6071 185
R14601 gnd.n6070 gnd.n6069 185
R14602 gnd.n6061 gnd.n6060 185
R14603 gnd.n6064 gnd.n6063 185
R14604 gnd.n6048 gnd.n6047 185
R14605 gnd.n6046 gnd.n6045 185
R14606 gnd.n6025 gnd.n6024 185
R14607 gnd.n6040 gnd.n6039 185
R14608 gnd.n6038 gnd.n6037 185
R14609 gnd.n6029 gnd.n6028 185
R14610 gnd.n6032 gnd.n6031 185
R14611 gnd.n6016 gnd.n6015 185
R14612 gnd.n6014 gnd.n6013 185
R14613 gnd.n5993 gnd.n5992 185
R14614 gnd.n6008 gnd.n6007 185
R14615 gnd.n6006 gnd.n6005 185
R14616 gnd.n5997 gnd.n5996 185
R14617 gnd.n6000 gnd.n5999 185
R14618 gnd.n5985 gnd.n5984 185
R14619 gnd.n5983 gnd.n5982 185
R14620 gnd.n5962 gnd.n5961 185
R14621 gnd.n5977 gnd.n5976 185
R14622 gnd.n5975 gnd.n5974 185
R14623 gnd.n5966 gnd.n5965 185
R14624 gnd.n5969 gnd.n5968 185
R14625 gnd.n5953 gnd.n5952 185
R14626 gnd.n5951 gnd.n5950 185
R14627 gnd.n5930 gnd.n5929 185
R14628 gnd.n5945 gnd.n5944 185
R14629 gnd.n5943 gnd.n5942 185
R14630 gnd.n5934 gnd.n5933 185
R14631 gnd.n5937 gnd.n5936 185
R14632 gnd.n5921 gnd.n5920 185
R14633 gnd.n5919 gnd.n5918 185
R14634 gnd.n5898 gnd.n5897 185
R14635 gnd.n5913 gnd.n5912 185
R14636 gnd.n5911 gnd.n5910 185
R14637 gnd.n5902 gnd.n5901 185
R14638 gnd.n5905 gnd.n5904 185
R14639 gnd.n5889 gnd.n5888 185
R14640 gnd.n5887 gnd.n5886 185
R14641 gnd.n5866 gnd.n5865 185
R14642 gnd.n5881 gnd.n5880 185
R14643 gnd.n5879 gnd.n5878 185
R14644 gnd.n5870 gnd.n5869 185
R14645 gnd.n5873 gnd.n5872 185
R14646 gnd.n5858 gnd.n5857 185
R14647 gnd.n5856 gnd.n5855 185
R14648 gnd.n5835 gnd.n5834 185
R14649 gnd.n5850 gnd.n5849 185
R14650 gnd.n5848 gnd.n5847 185
R14651 gnd.n5839 gnd.n5838 185
R14652 gnd.n5842 gnd.n5841 185
R14653 gnd.n5287 gnd.t107 178.987
R14654 gnd.n4908 gnd.t71 178.987
R14655 gnd.n4393 gnd.n1466 171.457
R14656 gnd.n3641 gnd.n3640 171.457
R14657 gnd.n1 gnd.t15 170.774
R14658 gnd.n9 gnd.t34 170.103
R14659 gnd.n8 gnd.t29 170.103
R14660 gnd.n7 gnd.t44 170.103
R14661 gnd.n6 gnd.t3 170.103
R14662 gnd.n5 gnd.t48 170.103
R14663 gnd.n4 gnd.t25 170.103
R14664 gnd.n3 gnd.t53 170.103
R14665 gnd.n2 gnd.t50 170.103
R14666 gnd.n1 gnd.t13 170.103
R14667 gnd.n3373 gnd.n3372 163.367
R14668 gnd.n3370 gnd.n3198 163.367
R14669 gnd.n3366 gnd.n3365 163.367
R14670 gnd.n3363 gnd.n3201 163.367
R14671 gnd.n3359 gnd.n3358 163.367
R14672 gnd.n3356 gnd.n3204 163.367
R14673 gnd.n3352 gnd.n3351 163.367
R14674 gnd.n3349 gnd.n3207 163.367
R14675 gnd.n3345 gnd.n3344 163.367
R14676 gnd.n3342 gnd.n3210 163.367
R14677 gnd.n3338 gnd.n3337 163.367
R14678 gnd.n3335 gnd.n3213 163.367
R14679 gnd.n3331 gnd.n3330 163.367
R14680 gnd.n3328 gnd.n3216 163.367
R14681 gnd.n3323 gnd.n3322 163.367
R14682 gnd.n3320 gnd.n3318 163.367
R14683 gnd.n3315 gnd.n3314 163.367
R14684 gnd.n3312 gnd.n3222 163.367
R14685 gnd.n3307 gnd.n3306 163.367
R14686 gnd.n3304 gnd.n3227 163.367
R14687 gnd.n3300 gnd.n3299 163.367
R14688 gnd.n3297 gnd.n3230 163.367
R14689 gnd.n3293 gnd.n3292 163.367
R14690 gnd.n3290 gnd.n3233 163.367
R14691 gnd.n3286 gnd.n3285 163.367
R14692 gnd.n3283 gnd.n3236 163.367
R14693 gnd.n3279 gnd.n3278 163.367
R14694 gnd.n3276 gnd.n3239 163.367
R14695 gnd.n3272 gnd.n3271 163.367
R14696 gnd.n3269 gnd.n3242 163.367
R14697 gnd.n3265 gnd.n3264 163.367
R14698 gnd.n3262 gnd.n3245 163.367
R14699 gnd.n3572 gnd.n2891 163.367
R14700 gnd.n3564 gnd.n2891 163.367
R14701 gnd.n3564 gnd.n3000 163.367
R14702 gnd.n3560 gnd.n3000 163.367
R14703 gnd.n3560 gnd.n3003 163.367
R14704 gnd.n3010 gnd.n3003 163.367
R14705 gnd.n3551 gnd.n3010 163.367
R14706 gnd.n3551 gnd.n3011 163.367
R14707 gnd.n3547 gnd.n3011 163.367
R14708 gnd.n3547 gnd.n3546 163.367
R14709 gnd.n3546 gnd.n3014 163.367
R14710 gnd.n3023 gnd.n3014 163.367
R14711 gnd.n3537 gnd.n3023 163.367
R14712 gnd.n3537 gnd.n3024 163.367
R14713 gnd.n3533 gnd.n3024 163.367
R14714 gnd.n3533 gnd.n3532 163.367
R14715 gnd.n3532 gnd.n3028 163.367
R14716 gnd.n3036 gnd.n3028 163.367
R14717 gnd.n3037 gnd.n3036 163.367
R14718 gnd.n3038 gnd.n3037 163.367
R14719 gnd.n3049 gnd.n3038 163.367
R14720 gnd.n3049 gnd.n3043 163.367
R14721 gnd.n3514 gnd.n3043 163.367
R14722 gnd.n3514 gnd.n3044 163.367
R14723 gnd.n3510 gnd.n3044 163.367
R14724 gnd.n3510 gnd.n3053 163.367
R14725 gnd.n3068 gnd.n3053 163.367
R14726 gnd.n3069 gnd.n3068 163.367
R14727 gnd.n3069 gnd.n3066 163.367
R14728 gnd.n3075 gnd.n3066 163.367
R14729 gnd.n3076 gnd.n3075 163.367
R14730 gnd.n3077 gnd.n3076 163.367
R14731 gnd.n3077 gnd.n3063 163.367
R14732 gnd.n3492 gnd.n3063 163.367
R14733 gnd.n3492 gnd.n3064 163.367
R14734 gnd.n3488 gnd.n3064 163.367
R14735 gnd.n3488 gnd.n3081 163.367
R14736 gnd.n3090 gnd.n3081 163.367
R14737 gnd.n3478 gnd.n3090 163.367
R14738 gnd.n3478 gnd.n3091 163.367
R14739 gnd.n3474 gnd.n3091 163.367
R14740 gnd.n3474 gnd.n3473 163.367
R14741 gnd.n3473 gnd.n3094 163.367
R14742 gnd.n3103 gnd.n3094 163.367
R14743 gnd.n3463 gnd.n3103 163.367
R14744 gnd.n3463 gnd.n3104 163.367
R14745 gnd.n3459 gnd.n3104 163.367
R14746 gnd.n3459 gnd.n3458 163.367
R14747 gnd.n3458 gnd.n3108 163.367
R14748 gnd.n3116 gnd.n3108 163.367
R14749 gnd.n3448 gnd.n3116 163.367
R14750 gnd.n3448 gnd.n3117 163.367
R14751 gnd.n3444 gnd.n3117 163.367
R14752 gnd.n3444 gnd.n3121 163.367
R14753 gnd.n3436 gnd.n3121 163.367
R14754 gnd.n3436 gnd.n3128 163.367
R14755 gnd.n3432 gnd.n3128 163.367
R14756 gnd.n3432 gnd.n3130 163.367
R14757 gnd.n3136 gnd.n3130 163.367
R14758 gnd.n3423 gnd.n3136 163.367
R14759 gnd.n3423 gnd.n3137 163.367
R14760 gnd.n3419 gnd.n3137 163.367
R14761 gnd.n3419 gnd.n3418 163.367
R14762 gnd.n3418 gnd.n3140 163.367
R14763 gnd.n3148 gnd.n3140 163.367
R14764 gnd.n3408 gnd.n3148 163.367
R14765 gnd.n3408 gnd.n3149 163.367
R14766 gnd.n3404 gnd.n3149 163.367
R14767 gnd.n3404 gnd.n3153 163.367
R14768 gnd.n3163 gnd.n3153 163.367
R14769 gnd.n3163 gnd.n3161 163.367
R14770 gnd.n3393 gnd.n3161 163.367
R14771 gnd.n3393 gnd.n3162 163.367
R14772 gnd.n3389 gnd.n3162 163.367
R14773 gnd.n3389 gnd.n3388 163.367
R14774 gnd.n3388 gnd.n3167 163.367
R14775 gnd.n3250 gnd.n3167 163.367
R14776 gnd.n3250 gnd.n3248 163.367
R14777 gnd.n3254 gnd.n3248 163.367
R14778 gnd.n3257 gnd.n3254 163.367
R14779 gnd.n2993 gnd.n2991 163.367
R14780 gnd.n2991 gnd.n2990 163.367
R14781 gnd.n2987 gnd.n2986 163.367
R14782 gnd.n2984 gnd.n2918 163.367
R14783 gnd.n2980 gnd.n2978 163.367
R14784 gnd.n2976 gnd.n2920 163.367
R14785 gnd.n2972 gnd.n2970 163.367
R14786 gnd.n2968 gnd.n2922 163.367
R14787 gnd.n2964 gnd.n2962 163.367
R14788 gnd.n2960 gnd.n2924 163.367
R14789 gnd.n2956 gnd.n2954 163.367
R14790 gnd.n2952 gnd.n2926 163.367
R14791 gnd.n2948 gnd.n2946 163.367
R14792 gnd.n2944 gnd.n2928 163.367
R14793 gnd.n2940 gnd.n2938 163.367
R14794 gnd.n2935 gnd.n2934 163.367
R14795 gnd.n3639 gnd.n3637 163.367
R14796 gnd.n3635 gnd.n2873 163.367
R14797 gnd.n3630 gnd.n3628 163.367
R14798 gnd.n3626 gnd.n2877 163.367
R14799 gnd.n3622 gnd.n3620 163.367
R14800 gnd.n3618 gnd.n2879 163.367
R14801 gnd.n3614 gnd.n3612 163.367
R14802 gnd.n3610 gnd.n2881 163.367
R14803 gnd.n3606 gnd.n3604 163.367
R14804 gnd.n3602 gnd.n2883 163.367
R14805 gnd.n3598 gnd.n3596 163.367
R14806 gnd.n3594 gnd.n2885 163.367
R14807 gnd.n3590 gnd.n3588 163.367
R14808 gnd.n3586 gnd.n2887 163.367
R14809 gnd.n3582 gnd.n3580 163.367
R14810 gnd.n3578 gnd.n2889 163.367
R14811 gnd.n3570 gnd.n2894 163.367
R14812 gnd.n3566 gnd.n2894 163.367
R14813 gnd.n3566 gnd.n2998 163.367
R14814 gnd.n3558 gnd.n2998 163.367
R14815 gnd.n3558 gnd.n3006 163.367
R14816 gnd.n3554 gnd.n3006 163.367
R14817 gnd.n3554 gnd.n3553 163.367
R14818 gnd.n3553 gnd.n3008 163.367
R14819 gnd.n3016 gnd.n3008 163.367
R14820 gnd.n3544 gnd.n3016 163.367
R14821 gnd.n3544 gnd.n3017 163.367
R14822 gnd.n3540 gnd.n3017 163.367
R14823 gnd.n3540 gnd.n3539 163.367
R14824 gnd.n3539 gnd.n3021 163.367
R14825 gnd.n3030 gnd.n3021 163.367
R14826 gnd.n3530 gnd.n3030 163.367
R14827 gnd.n3530 gnd.n3031 163.367
R14828 gnd.n3526 gnd.n3031 163.367
R14829 gnd.n3526 gnd.n3035 163.367
R14830 gnd.n3521 gnd.n3035 163.367
R14831 gnd.n3521 gnd.n3039 163.367
R14832 gnd.n3517 gnd.n3039 163.367
R14833 gnd.n3517 gnd.n3041 163.367
R14834 gnd.n3055 gnd.n3041 163.367
R14835 gnd.n3508 gnd.n3055 163.367
R14836 gnd.n3508 gnd.n3056 163.367
R14837 gnd.n3504 gnd.n3056 163.367
R14838 gnd.n3504 gnd.n3503 163.367
R14839 gnd.n3503 gnd.n3502 163.367
R14840 gnd.n3502 gnd.n3059 163.367
R14841 gnd.n3498 gnd.n3059 163.367
R14842 gnd.n3498 gnd.n3497 163.367
R14843 gnd.n3497 gnd.n3496 163.367
R14844 gnd.n3496 gnd.n3061 163.367
R14845 gnd.n3083 gnd.n3061 163.367
R14846 gnd.n3486 gnd.n3083 163.367
R14847 gnd.n3486 gnd.n3085 163.367
R14848 gnd.n3482 gnd.n3085 163.367
R14849 gnd.n3482 gnd.n3481 163.367
R14850 gnd.n3481 gnd.n3089 163.367
R14851 gnd.n3096 gnd.n3089 163.367
R14852 gnd.n3471 gnd.n3096 163.367
R14853 gnd.n3471 gnd.n3098 163.367
R14854 gnd.n3467 gnd.n3098 163.367
R14855 gnd.n3467 gnd.n3466 163.367
R14856 gnd.n3466 gnd.n3102 163.367
R14857 gnd.n3110 gnd.n3102 163.367
R14858 gnd.n3456 gnd.n3110 163.367
R14859 gnd.n3456 gnd.n3111 163.367
R14860 gnd.n3452 gnd.n3111 163.367
R14861 gnd.n3452 gnd.n3451 163.367
R14862 gnd.n3451 gnd.n3115 163.367
R14863 gnd.n3442 gnd.n3115 163.367
R14864 gnd.n3442 gnd.n3123 163.367
R14865 gnd.n3438 gnd.n3123 163.367
R14866 gnd.n3438 gnd.n3126 163.367
R14867 gnd.n3430 gnd.n3126 163.367
R14868 gnd.n3430 gnd.n3132 163.367
R14869 gnd.n3426 gnd.n3132 163.367
R14870 gnd.n3426 gnd.n3425 163.367
R14871 gnd.n3425 gnd.n3134 163.367
R14872 gnd.n3142 gnd.n3134 163.367
R14873 gnd.n3416 gnd.n3142 163.367
R14874 gnd.n3416 gnd.n3143 163.367
R14875 gnd.n3412 gnd.n3143 163.367
R14876 gnd.n3412 gnd.n3147 163.367
R14877 gnd.n3155 gnd.n3147 163.367
R14878 gnd.n3402 gnd.n3155 163.367
R14879 gnd.n3402 gnd.n3157 163.367
R14880 gnd.n3398 gnd.n3157 163.367
R14881 gnd.n3398 gnd.n3397 163.367
R14882 gnd.n3397 gnd.n3160 163.367
R14883 gnd.n3171 gnd.n3160 163.367
R14884 gnd.n3171 gnd.n3168 163.367
R14885 gnd.n3386 gnd.n3168 163.367
R14886 gnd.n3386 gnd.n3169 163.367
R14887 gnd.n3382 gnd.n3169 163.367
R14888 gnd.n3382 gnd.n3381 163.367
R14889 gnd.n3381 gnd.n3380 163.367
R14890 gnd.n3380 gnd.n3175 163.367
R14891 gnd.n3194 gnd.n3193 156.462
R14892 gnd.n6020 gnd.n5988 153.042
R14893 gnd.n6084 gnd.n6083 152.079
R14894 gnd.n6052 gnd.n6051 152.079
R14895 gnd.n6020 gnd.n6019 152.079
R14896 gnd.n2907 gnd.n2906 152
R14897 gnd.n2908 gnd.n2897 152
R14898 gnd.n2910 gnd.n2909 152
R14899 gnd.n2912 gnd.n2895 152
R14900 gnd.n2914 gnd.n2913 152
R14901 gnd.n3192 gnd.n3176 152
R14902 gnd.n3184 gnd.n3177 152
R14903 gnd.n3183 gnd.n3182 152
R14904 gnd.n3181 gnd.n3178 152
R14905 gnd.n3179 gnd.t116 150.546
R14906 gnd.t58 gnd.n6062 147.661
R14907 gnd.t330 gnd.n6030 147.661
R14908 gnd.t22 gnd.n5998 147.661
R14909 gnd.t27 gnd.n5967 147.661
R14910 gnd.t37 gnd.n5935 147.661
R14911 gnd.t42 gnd.n5903 147.661
R14912 gnd.t64 gnd.n5871 147.661
R14913 gnd.t326 gnd.n5840 147.661
R14914 gnd.n3317 gnd.n3316 143.351
R14915 gnd.n2933 gnd.n2872 143.351
R14916 gnd.n3638 gnd.n2872 143.351
R14917 gnd.n2904 gnd.t145 130.484
R14918 gnd.n6887 gnd.n6886 127.278
R14919 gnd.n6888 gnd.n6887 127.278
R14920 gnd.n6888 gnd.n448 127.278
R14921 gnd.n6896 gnd.n448 127.278
R14922 gnd.n6897 gnd.n6896 127.278
R14923 gnd.n6898 gnd.n6897 127.278
R14924 gnd.n6898 gnd.n442 127.278
R14925 gnd.n6906 gnd.n442 127.278
R14926 gnd.n6907 gnd.n6906 127.278
R14927 gnd.n6908 gnd.n6907 127.278
R14928 gnd.n6908 gnd.n436 127.278
R14929 gnd.n6916 gnd.n436 127.278
R14930 gnd.n6917 gnd.n6916 127.278
R14931 gnd.n6918 gnd.n6917 127.278
R14932 gnd.n6918 gnd.n430 127.278
R14933 gnd.n6926 gnd.n430 127.278
R14934 gnd.n6927 gnd.n6926 127.278
R14935 gnd.n6928 gnd.n6927 127.278
R14936 gnd.n6928 gnd.n424 127.278
R14937 gnd.n6936 gnd.n424 127.278
R14938 gnd.n6937 gnd.n6936 127.278
R14939 gnd.n6938 gnd.n6937 127.278
R14940 gnd.n6938 gnd.n418 127.278
R14941 gnd.n6946 gnd.n418 127.278
R14942 gnd.n6947 gnd.n6946 127.278
R14943 gnd.n6948 gnd.n6947 127.278
R14944 gnd.n6948 gnd.n412 127.278
R14945 gnd.n6956 gnd.n412 127.278
R14946 gnd.n6957 gnd.n6956 127.278
R14947 gnd.n6958 gnd.n6957 127.278
R14948 gnd.n6958 gnd.n406 127.278
R14949 gnd.n6966 gnd.n406 127.278
R14950 gnd.n6967 gnd.n6966 127.278
R14951 gnd.n6968 gnd.n6967 127.278
R14952 gnd.n6968 gnd.n400 127.278
R14953 gnd.n6976 gnd.n400 127.278
R14954 gnd.n6977 gnd.n6976 127.278
R14955 gnd.n6978 gnd.n6977 127.278
R14956 gnd.n6978 gnd.n394 127.278
R14957 gnd.n6986 gnd.n394 127.278
R14958 gnd.n6987 gnd.n6986 127.278
R14959 gnd.n6988 gnd.n6987 127.278
R14960 gnd.n6988 gnd.n388 127.278
R14961 gnd.n6996 gnd.n388 127.278
R14962 gnd.n6997 gnd.n6996 127.278
R14963 gnd.n6998 gnd.n6997 127.278
R14964 gnd.n6998 gnd.n382 127.278
R14965 gnd.n7006 gnd.n382 127.278
R14966 gnd.n7007 gnd.n7006 127.278
R14967 gnd.n7008 gnd.n7007 127.278
R14968 gnd.n7008 gnd.n376 127.278
R14969 gnd.n7016 gnd.n376 127.278
R14970 gnd.n7017 gnd.n7016 127.278
R14971 gnd.n7018 gnd.n7017 127.278
R14972 gnd.n7018 gnd.n370 127.278
R14973 gnd.n7026 gnd.n370 127.278
R14974 gnd.n7027 gnd.n7026 127.278
R14975 gnd.n7028 gnd.n7027 127.278
R14976 gnd.n7028 gnd.n364 127.278
R14977 gnd.n7036 gnd.n364 127.278
R14978 gnd.n7037 gnd.n7036 127.278
R14979 gnd.n7038 gnd.n7037 127.278
R14980 gnd.n7038 gnd.n358 127.278
R14981 gnd.n7046 gnd.n358 127.278
R14982 gnd.n7047 gnd.n7046 127.278
R14983 gnd.n7048 gnd.n7047 127.278
R14984 gnd.n7048 gnd.n352 127.278
R14985 gnd.n7056 gnd.n352 127.278
R14986 gnd.n7057 gnd.n7056 127.278
R14987 gnd.n7058 gnd.n7057 127.278
R14988 gnd.n7058 gnd.n346 127.278
R14989 gnd.n7066 gnd.n346 127.278
R14990 gnd.n7067 gnd.n7066 127.278
R14991 gnd.n7068 gnd.n7067 127.278
R14992 gnd.n7068 gnd.n340 127.278
R14993 gnd.n7076 gnd.n340 127.278
R14994 gnd.n7077 gnd.n7076 127.278
R14995 gnd.n7078 gnd.n7077 127.278
R14996 gnd.n7078 gnd.n334 127.278
R14997 gnd.n7086 gnd.n334 127.278
R14998 gnd.n7087 gnd.n7086 127.278
R14999 gnd.n7089 gnd.n7087 127.278
R15000 gnd.n7089 gnd.n7088 127.278
R15001 gnd.n2913 gnd.t79 126.766
R15002 gnd.n2911 gnd.t139 126.766
R15003 gnd.n2897 gnd.t161 126.766
R15004 gnd.n2905 gnd.t123 126.766
R15005 gnd.n3180 gnd.t155 126.766
R15006 gnd.n3182 gnd.t130 126.766
R15007 gnd.n3191 gnd.t76 126.766
R15008 gnd.n3193 gnd.t133 126.766
R15009 gnd.n6079 gnd.n6078 104.615
R15010 gnd.n6078 gnd.n6056 104.615
R15011 gnd.n6071 gnd.n6056 104.615
R15012 gnd.n6071 gnd.n6070 104.615
R15013 gnd.n6070 gnd.n6060 104.615
R15014 gnd.n6063 gnd.n6060 104.615
R15015 gnd.n6047 gnd.n6046 104.615
R15016 gnd.n6046 gnd.n6024 104.615
R15017 gnd.n6039 gnd.n6024 104.615
R15018 gnd.n6039 gnd.n6038 104.615
R15019 gnd.n6038 gnd.n6028 104.615
R15020 gnd.n6031 gnd.n6028 104.615
R15021 gnd.n6015 gnd.n6014 104.615
R15022 gnd.n6014 gnd.n5992 104.615
R15023 gnd.n6007 gnd.n5992 104.615
R15024 gnd.n6007 gnd.n6006 104.615
R15025 gnd.n6006 gnd.n5996 104.615
R15026 gnd.n5999 gnd.n5996 104.615
R15027 gnd.n5984 gnd.n5983 104.615
R15028 gnd.n5983 gnd.n5961 104.615
R15029 gnd.n5976 gnd.n5961 104.615
R15030 gnd.n5976 gnd.n5975 104.615
R15031 gnd.n5975 gnd.n5965 104.615
R15032 gnd.n5968 gnd.n5965 104.615
R15033 gnd.n5952 gnd.n5951 104.615
R15034 gnd.n5951 gnd.n5929 104.615
R15035 gnd.n5944 gnd.n5929 104.615
R15036 gnd.n5944 gnd.n5943 104.615
R15037 gnd.n5943 gnd.n5933 104.615
R15038 gnd.n5936 gnd.n5933 104.615
R15039 gnd.n5920 gnd.n5919 104.615
R15040 gnd.n5919 gnd.n5897 104.615
R15041 gnd.n5912 gnd.n5897 104.615
R15042 gnd.n5912 gnd.n5911 104.615
R15043 gnd.n5911 gnd.n5901 104.615
R15044 gnd.n5904 gnd.n5901 104.615
R15045 gnd.n5888 gnd.n5887 104.615
R15046 gnd.n5887 gnd.n5865 104.615
R15047 gnd.n5880 gnd.n5865 104.615
R15048 gnd.n5880 gnd.n5879 104.615
R15049 gnd.n5879 gnd.n5869 104.615
R15050 gnd.n5872 gnd.n5869 104.615
R15051 gnd.n5857 gnd.n5856 104.615
R15052 gnd.n5856 gnd.n5834 104.615
R15053 gnd.n5849 gnd.n5834 104.615
R15054 gnd.n5849 gnd.n5848 104.615
R15055 gnd.n5848 gnd.n5838 104.615
R15056 gnd.n5841 gnd.n5838 104.615
R15057 gnd.n5212 gnd.t151 100.632
R15058 gnd.n4863 gnd.t92 100.632
R15059 gnd.n7453 gnd.n116 99.6594
R15060 gnd.n7451 gnd.n7450 99.6594
R15061 gnd.n7446 gnd.n123 99.6594
R15062 gnd.n7444 gnd.n7443 99.6594
R15063 gnd.n7439 gnd.n130 99.6594
R15064 gnd.n7437 gnd.n7436 99.6594
R15065 gnd.n7432 gnd.n137 99.6594
R15066 gnd.n7430 gnd.n7429 99.6594
R15067 gnd.n7422 gnd.n144 99.6594
R15068 gnd.n7420 gnd.n7419 99.6594
R15069 gnd.n7415 gnd.n151 99.6594
R15070 gnd.n7413 gnd.n7412 99.6594
R15071 gnd.n7408 gnd.n158 99.6594
R15072 gnd.n7406 gnd.n7405 99.6594
R15073 gnd.n7401 gnd.n165 99.6594
R15074 gnd.n7399 gnd.n7398 99.6594
R15075 gnd.n7394 gnd.n172 99.6594
R15076 gnd.n7392 gnd.n7391 99.6594
R15077 gnd.n177 gnd.n176 99.6594
R15078 gnd.n4424 gnd.n4423 99.6594
R15079 gnd.n4418 gnd.n1418 99.6594
R15080 gnd.n4415 gnd.n1419 99.6594
R15081 gnd.n4411 gnd.n1420 99.6594
R15082 gnd.n4407 gnd.n1421 99.6594
R15083 gnd.n4403 gnd.n1422 99.6594
R15084 gnd.n4399 gnd.n1423 99.6594
R15085 gnd.n4395 gnd.n1424 99.6594
R15086 gnd.n4390 gnd.n1426 99.6594
R15087 gnd.n4386 gnd.n1427 99.6594
R15088 gnd.n4382 gnd.n1428 99.6594
R15089 gnd.n4378 gnd.n1429 99.6594
R15090 gnd.n4374 gnd.n1430 99.6594
R15091 gnd.n4370 gnd.n1431 99.6594
R15092 gnd.n4366 gnd.n1432 99.6594
R15093 gnd.n4362 gnd.n1433 99.6594
R15094 gnd.n4358 gnd.n1434 99.6594
R15095 gnd.n1490 gnd.n1435 99.6594
R15096 gnd.n3669 gnd.n3668 99.6594
R15097 gnd.n3664 gnd.n2268 99.6594
R15098 gnd.n3660 gnd.n2267 99.6594
R15099 gnd.n3656 gnd.n2266 99.6594
R15100 gnd.n3652 gnd.n2265 99.6594
R15101 gnd.n3648 gnd.n2264 99.6594
R15102 gnd.n3644 gnd.n2263 99.6594
R15103 gnd.n2864 gnd.n2261 99.6594
R15104 gnd.n2862 gnd.n2260 99.6594
R15105 gnd.n2858 gnd.n2259 99.6594
R15106 gnd.n2854 gnd.n2258 99.6594
R15107 gnd.n2850 gnd.n2257 99.6594
R15108 gnd.n2846 gnd.n2256 99.6594
R15109 gnd.n2842 gnd.n2255 99.6594
R15110 gnd.n2838 gnd.n2254 99.6594
R15111 gnd.n2834 gnd.n2253 99.6594
R15112 gnd.n2830 gnd.n2252 99.6594
R15113 gnd.n2310 gnd.n2251 99.6594
R15114 gnd.n4831 gnd.n4830 99.6594
R15115 gnd.n4825 gnd.n933 99.6594
R15116 gnd.n4822 gnd.n934 99.6594
R15117 gnd.n4818 gnd.n935 99.6594
R15118 gnd.n4814 gnd.n936 99.6594
R15119 gnd.n4810 gnd.n937 99.6594
R15120 gnd.n4806 gnd.n938 99.6594
R15121 gnd.n4802 gnd.n939 99.6594
R15122 gnd.n4798 gnd.n940 99.6594
R15123 gnd.n4793 gnd.n941 99.6594
R15124 gnd.n4789 gnd.n942 99.6594
R15125 gnd.n4785 gnd.n943 99.6594
R15126 gnd.n4781 gnd.n944 99.6594
R15127 gnd.n4777 gnd.n945 99.6594
R15128 gnd.n4773 gnd.n946 99.6594
R15129 gnd.n4769 gnd.n947 99.6594
R15130 gnd.n4765 gnd.n948 99.6594
R15131 gnd.n4761 gnd.n949 99.6594
R15132 gnd.n1004 gnd.n950 99.6594
R15133 gnd.n6228 gnd.n4843 99.6594
R15134 gnd.n6226 gnd.n6225 99.6594
R15135 gnd.n6221 gnd.n4850 99.6594
R15136 gnd.n6219 gnd.n6218 99.6594
R15137 gnd.n6214 gnd.n4857 99.6594
R15138 gnd.n6212 gnd.n6211 99.6594
R15139 gnd.n6207 gnd.n4866 99.6594
R15140 gnd.n6205 gnd.n6204 99.6594
R15141 gnd.n5510 gnd.n5155 99.6594
R15142 gnd.n5181 gnd.n5162 99.6594
R15143 gnd.n5183 gnd.n5163 99.6594
R15144 gnd.n5191 gnd.n5164 99.6594
R15145 gnd.n5193 gnd.n5165 99.6594
R15146 gnd.n5201 gnd.n5166 99.6594
R15147 gnd.n5203 gnd.n5167 99.6594
R15148 gnd.n5211 gnd.n5168 99.6594
R15149 gnd.n6196 gnd.n4873 99.6594
R15150 gnd.n6194 gnd.n6193 99.6594
R15151 gnd.n6189 gnd.n4880 99.6594
R15152 gnd.n6187 gnd.n6186 99.6594
R15153 gnd.n6182 gnd.n4887 99.6594
R15154 gnd.n6180 gnd.n6179 99.6594
R15155 gnd.n6175 gnd.n4894 99.6594
R15156 gnd.n6173 gnd.n6172 99.6594
R15157 gnd.n6168 gnd.n4901 99.6594
R15158 gnd.n6166 gnd.n6165 99.6594
R15159 gnd.n6161 gnd.n4910 99.6594
R15160 gnd.n6159 gnd.n6158 99.6594
R15161 gnd.n6154 gnd.n6153 99.6594
R15162 gnd.n5339 gnd.n5338 99.6594
R15163 gnd.n5333 gnd.n5250 99.6594
R15164 gnd.n5330 gnd.n5251 99.6594
R15165 gnd.n5326 gnd.n5252 99.6594
R15166 gnd.n5322 gnd.n5253 99.6594
R15167 gnd.n5318 gnd.n5254 99.6594
R15168 gnd.n5314 gnd.n5255 99.6594
R15169 gnd.n5310 gnd.n5256 99.6594
R15170 gnd.n5306 gnd.n5257 99.6594
R15171 gnd.n5302 gnd.n5258 99.6594
R15172 gnd.n5298 gnd.n5259 99.6594
R15173 gnd.n5294 gnd.n5260 99.6594
R15174 gnd.n5341 gnd.n5249 99.6594
R15175 gnd.n7301 gnd.n7300 99.6594
R15176 gnd.n7306 gnd.n7305 99.6594
R15177 gnd.n7309 gnd.n7308 99.6594
R15178 gnd.n7314 gnd.n7313 99.6594
R15179 gnd.n7317 gnd.n7316 99.6594
R15180 gnd.n7322 gnd.n7321 99.6594
R15181 gnd.n7325 gnd.n7324 99.6594
R15182 gnd.n7330 gnd.n7329 99.6594
R15183 gnd.n7333 gnd.n103 99.6594
R15184 gnd.n1500 gnd.n1436 99.6594
R15185 gnd.n1728 gnd.n1437 99.6594
R15186 gnd.n1730 gnd.n1438 99.6594
R15187 gnd.n1747 gnd.n1439 99.6594
R15188 gnd.n1749 gnd.n1440 99.6594
R15189 gnd.n1766 gnd.n1441 99.6594
R15190 gnd.n1768 gnd.n1442 99.6594
R15191 gnd.n1784 gnd.n1443 99.6594
R15192 gnd.n1695 gnd.n1444 99.6594
R15193 gnd.n2238 gnd.n2237 99.6594
R15194 gnd.n2239 gnd.n2187 99.6594
R15195 gnd.n2241 gnd.n2195 99.6594
R15196 gnd.n2243 gnd.n2242 99.6594
R15197 gnd.n2244 gnd.n2204 99.6594
R15198 gnd.n2246 gnd.n2213 99.6594
R15199 gnd.n2248 gnd.n2247 99.6594
R15200 gnd.n2249 gnd.n2222 99.6594
R15201 gnd.n3672 gnd.n3671 99.6594
R15202 gnd.n2518 gnd.n951 99.6594
R15203 gnd.n2515 gnd.n952 99.6594
R15204 gnd.n2511 gnd.n953 99.6594
R15205 gnd.n2507 gnd.n954 99.6594
R15206 gnd.n2503 gnd.n955 99.6594
R15207 gnd.n2499 gnd.n956 99.6594
R15208 gnd.n2495 gnd.n957 99.6594
R15209 gnd.n2491 gnd.n958 99.6594
R15210 gnd.n2487 gnd.n959 99.6594
R15211 gnd.n2516 gnd.n951 99.6594
R15212 gnd.n2512 gnd.n952 99.6594
R15213 gnd.n2508 gnd.n953 99.6594
R15214 gnd.n2504 gnd.n954 99.6594
R15215 gnd.n2500 gnd.n955 99.6594
R15216 gnd.n2496 gnd.n956 99.6594
R15217 gnd.n2492 gnd.n957 99.6594
R15218 gnd.n2488 gnd.n958 99.6594
R15219 gnd.n2476 gnd.n959 99.6594
R15220 gnd.n3671 gnd.n2233 99.6594
R15221 gnd.n2249 gnd.n2221 99.6594
R15222 gnd.n2248 gnd.n2214 99.6594
R15223 gnd.n2246 gnd.n2245 99.6594
R15224 gnd.n2244 gnd.n2203 99.6594
R15225 gnd.n2243 gnd.n2196 99.6594
R15226 gnd.n2241 gnd.n2240 99.6594
R15227 gnd.n2239 gnd.n2186 99.6594
R15228 gnd.n2238 gnd.n2236 99.6594
R15229 gnd.n1727 gnd.n1436 99.6594
R15230 gnd.n1731 gnd.n1437 99.6594
R15231 gnd.n1746 gnd.n1438 99.6594
R15232 gnd.n1750 gnd.n1439 99.6594
R15233 gnd.n1765 gnd.n1440 99.6594
R15234 gnd.n1769 gnd.n1441 99.6594
R15235 gnd.n1783 gnd.n1442 99.6594
R15236 gnd.n1694 gnd.n1443 99.6594
R15237 gnd.n1690 gnd.n1444 99.6594
R15238 gnd.n7334 gnd.n7333 99.6594
R15239 gnd.n7329 gnd.n7328 99.6594
R15240 gnd.n7324 gnd.n7323 99.6594
R15241 gnd.n7321 gnd.n7320 99.6594
R15242 gnd.n7316 gnd.n7315 99.6594
R15243 gnd.n7313 gnd.n7312 99.6594
R15244 gnd.n7308 gnd.n7307 99.6594
R15245 gnd.n7305 gnd.n7304 99.6594
R15246 gnd.n7300 gnd.n7299 99.6594
R15247 gnd.n5339 gnd.n5262 99.6594
R15248 gnd.n5331 gnd.n5250 99.6594
R15249 gnd.n5327 gnd.n5251 99.6594
R15250 gnd.n5323 gnd.n5252 99.6594
R15251 gnd.n5319 gnd.n5253 99.6594
R15252 gnd.n5315 gnd.n5254 99.6594
R15253 gnd.n5311 gnd.n5255 99.6594
R15254 gnd.n5307 gnd.n5256 99.6594
R15255 gnd.n5303 gnd.n5257 99.6594
R15256 gnd.n5299 gnd.n5258 99.6594
R15257 gnd.n5295 gnd.n5259 99.6594
R15258 gnd.n5291 gnd.n5260 99.6594
R15259 gnd.n5342 gnd.n5341 99.6594
R15260 gnd.n6153 gnd.n4912 99.6594
R15261 gnd.n6160 gnd.n6159 99.6594
R15262 gnd.n4910 gnd.n4902 99.6594
R15263 gnd.n6167 gnd.n6166 99.6594
R15264 gnd.n4901 gnd.n4895 99.6594
R15265 gnd.n6174 gnd.n6173 99.6594
R15266 gnd.n4894 gnd.n4888 99.6594
R15267 gnd.n6181 gnd.n6180 99.6594
R15268 gnd.n4887 gnd.n4881 99.6594
R15269 gnd.n6188 gnd.n6187 99.6594
R15270 gnd.n4880 gnd.n4874 99.6594
R15271 gnd.n6195 gnd.n6194 99.6594
R15272 gnd.n4873 gnd.n4870 99.6594
R15273 gnd.n5511 gnd.n5510 99.6594
R15274 gnd.n5184 gnd.n5162 99.6594
R15275 gnd.n5190 gnd.n5163 99.6594
R15276 gnd.n5194 gnd.n5164 99.6594
R15277 gnd.n5200 gnd.n5165 99.6594
R15278 gnd.n5204 gnd.n5166 99.6594
R15279 gnd.n5210 gnd.n5167 99.6594
R15280 gnd.n5168 gnd.n5152 99.6594
R15281 gnd.n6206 gnd.n6205 99.6594
R15282 gnd.n4866 gnd.n4858 99.6594
R15283 gnd.n6213 gnd.n6212 99.6594
R15284 gnd.n4857 gnd.n4851 99.6594
R15285 gnd.n6220 gnd.n6219 99.6594
R15286 gnd.n4850 gnd.n4844 99.6594
R15287 gnd.n6227 gnd.n6226 99.6594
R15288 gnd.n4843 gnd.n4840 99.6594
R15289 gnd.n4831 gnd.n963 99.6594
R15290 gnd.n4823 gnd.n933 99.6594
R15291 gnd.n4819 gnd.n934 99.6594
R15292 gnd.n4815 gnd.n935 99.6594
R15293 gnd.n4811 gnd.n936 99.6594
R15294 gnd.n4807 gnd.n937 99.6594
R15295 gnd.n4803 gnd.n938 99.6594
R15296 gnd.n4799 gnd.n939 99.6594
R15297 gnd.n4794 gnd.n940 99.6594
R15298 gnd.n4790 gnd.n941 99.6594
R15299 gnd.n4786 gnd.n942 99.6594
R15300 gnd.n4782 gnd.n943 99.6594
R15301 gnd.n4778 gnd.n944 99.6594
R15302 gnd.n4774 gnd.n945 99.6594
R15303 gnd.n4770 gnd.n946 99.6594
R15304 gnd.n4766 gnd.n947 99.6594
R15305 gnd.n4762 gnd.n948 99.6594
R15306 gnd.n1003 gnd.n949 99.6594
R15307 gnd.n4754 gnd.n950 99.6594
R15308 gnd.n2829 gnd.n2251 99.6594
R15309 gnd.n2833 gnd.n2252 99.6594
R15310 gnd.n2837 gnd.n2253 99.6594
R15311 gnd.n2841 gnd.n2254 99.6594
R15312 gnd.n2845 gnd.n2255 99.6594
R15313 gnd.n2849 gnd.n2256 99.6594
R15314 gnd.n2853 gnd.n2257 99.6594
R15315 gnd.n2857 gnd.n2258 99.6594
R15316 gnd.n2861 gnd.n2259 99.6594
R15317 gnd.n2865 gnd.n2260 99.6594
R15318 gnd.n3643 gnd.n2262 99.6594
R15319 gnd.n3647 gnd.n2263 99.6594
R15320 gnd.n3651 gnd.n2264 99.6594
R15321 gnd.n3655 gnd.n2265 99.6594
R15322 gnd.n3659 gnd.n2266 99.6594
R15323 gnd.n3663 gnd.n2267 99.6594
R15324 gnd.n2270 gnd.n2268 99.6594
R15325 gnd.n3669 gnd.n2269 99.6594
R15326 gnd.n4424 gnd.n1448 99.6594
R15327 gnd.n4416 gnd.n1418 99.6594
R15328 gnd.n4412 gnd.n1419 99.6594
R15329 gnd.n4408 gnd.n1420 99.6594
R15330 gnd.n4404 gnd.n1421 99.6594
R15331 gnd.n4400 gnd.n1422 99.6594
R15332 gnd.n4396 gnd.n1423 99.6594
R15333 gnd.n4391 gnd.n1425 99.6594
R15334 gnd.n4387 gnd.n1426 99.6594
R15335 gnd.n4383 gnd.n1427 99.6594
R15336 gnd.n4379 gnd.n1428 99.6594
R15337 gnd.n4375 gnd.n1429 99.6594
R15338 gnd.n4371 gnd.n1430 99.6594
R15339 gnd.n4367 gnd.n1431 99.6594
R15340 gnd.n4363 gnd.n1432 99.6594
R15341 gnd.n4359 gnd.n1433 99.6594
R15342 gnd.n1489 gnd.n1434 99.6594
R15343 gnd.n4351 gnd.n1435 99.6594
R15344 gnd.n176 gnd.n173 99.6594
R15345 gnd.n7393 gnd.n7392 99.6594
R15346 gnd.n172 gnd.n166 99.6594
R15347 gnd.n7400 gnd.n7399 99.6594
R15348 gnd.n165 gnd.n159 99.6594
R15349 gnd.n7407 gnd.n7406 99.6594
R15350 gnd.n158 gnd.n152 99.6594
R15351 gnd.n7414 gnd.n7413 99.6594
R15352 gnd.n151 gnd.n145 99.6594
R15353 gnd.n7421 gnd.n7420 99.6594
R15354 gnd.n144 gnd.n138 99.6594
R15355 gnd.n7431 gnd.n7430 99.6594
R15356 gnd.n137 gnd.n131 99.6594
R15357 gnd.n7438 gnd.n7437 99.6594
R15358 gnd.n130 gnd.n124 99.6594
R15359 gnd.n7445 gnd.n7444 99.6594
R15360 gnd.n123 gnd.n117 99.6594
R15361 gnd.n7452 gnd.n7451 99.6594
R15362 gnd.n116 gnd.n113 99.6594
R15363 gnd.n3719 gnd.n3718 99.6594
R15364 gnd.n2190 gnd.n2166 99.6594
R15365 gnd.n2192 gnd.n2167 99.6594
R15366 gnd.n2200 gnd.n2168 99.6594
R15367 gnd.n2208 gnd.n2169 99.6594
R15368 gnd.n2210 gnd.n2170 99.6594
R15369 gnd.n2218 gnd.n2171 99.6594
R15370 gnd.n2228 gnd.n2172 99.6594
R15371 gnd.n2230 gnd.n2173 99.6594
R15372 gnd.n2788 gnd.n2174 99.6594
R15373 gnd.n2790 gnd.n2175 99.6594
R15374 gnd.n2794 gnd.n2176 99.6594
R15375 gnd.n2800 gnd.n2177 99.6594
R15376 gnd.n3721 gnd.n2164 99.6594
R15377 gnd.n3719 gnd.n2180 99.6594
R15378 gnd.n2191 gnd.n2166 99.6594
R15379 gnd.n2199 gnd.n2167 99.6594
R15380 gnd.n2207 gnd.n2168 99.6594
R15381 gnd.n2209 gnd.n2169 99.6594
R15382 gnd.n2217 gnd.n2170 99.6594
R15383 gnd.n2227 gnd.n2171 99.6594
R15384 gnd.n2229 gnd.n2172 99.6594
R15385 gnd.n2787 gnd.n2173 99.6594
R15386 gnd.n2789 gnd.n2174 99.6594
R15387 gnd.n2793 gnd.n2175 99.6594
R15388 gnd.n2795 gnd.n2176 99.6594
R15389 gnd.n2801 gnd.n2177 99.6594
R15390 gnd.n3722 gnd.n3721 99.6594
R15391 gnd.n1736 gnd.n1718 99.6594
R15392 gnd.n1740 gnd.n1738 99.6594
R15393 gnd.n1755 gnd.n1711 99.6594
R15394 gnd.n1759 gnd.n1757 99.6594
R15395 gnd.n1774 gnd.n1704 99.6594
R15396 gnd.n1778 gnd.n1776 99.6594
R15397 gnd.n1790 gnd.n1698 99.6594
R15398 gnd.n1794 gnd.n1792 99.6594
R15399 gnd.n1804 gnd.n1686 99.6594
R15400 gnd.n1807 gnd.n1806 99.6594
R15401 gnd.n1810 gnd.n1809 99.6594
R15402 gnd.n1815 gnd.n1814 99.6594
R15403 gnd.n1818 gnd.n1817 99.6594
R15404 gnd.n4135 gnd.n4134 99.6594
R15405 gnd.n4134 gnd.n4133 99.6594
R15406 gnd.n1817 gnd.n1816 99.6594
R15407 gnd.n1814 gnd.n1813 99.6594
R15408 gnd.n1809 gnd.n1808 99.6594
R15409 gnd.n1806 gnd.n1805 99.6594
R15410 gnd.n1793 gnd.n1686 99.6594
R15411 gnd.n1792 gnd.n1791 99.6594
R15412 gnd.n1777 gnd.n1698 99.6594
R15413 gnd.n1776 gnd.n1775 99.6594
R15414 gnd.n1758 gnd.n1704 99.6594
R15415 gnd.n1757 gnd.n1756 99.6594
R15416 gnd.n1739 gnd.n1711 99.6594
R15417 gnd.n1738 gnd.n1737 99.6594
R15418 gnd.n1718 gnd.n1405 99.6594
R15419 gnd.n2796 gnd.t129 98.63
R15420 gnd.n7331 gnd.t143 98.63
R15421 gnd.n1691 gnd.t138 98.63
R15422 gnd.n2223 gnd.t159 98.63
R15423 gnd.n1469 gnd.t111 98.63
R15424 gnd.n1491 gnd.t101 98.63
R15425 gnd.n179 gnd.t173 98.63
R15426 gnd.n7424 gnd.t96 98.63
R15427 gnd.n983 gnd.t75 98.63
R15428 gnd.n1005 gnd.t154 98.63
R15429 gnd.n2312 gnd.t170 98.63
R15430 gnd.n2290 gnd.t88 98.63
R15431 gnd.n2477 gnd.t104 98.63
R15432 gnd.n4143 gnd.t84 98.63
R15433 gnd.n2874 gnd.t168 88.9408
R15434 gnd.n3223 gnd.t164 88.9408
R15435 gnd.n2929 gnd.t122 88.933
R15436 gnd.n3217 gnd.t114 88.933
R15437 gnd.n2904 gnd.n2903 81.8399
R15438 gnd.n7088 gnd.n186 76.3673
R15439 gnd.n5213 gnd.t150 74.8376
R15440 gnd.n4864 gnd.t93 74.8376
R15441 gnd.n2875 gnd.t167 72.8438
R15442 gnd.n3224 gnd.t165 72.8438
R15443 gnd.n2905 gnd.n2898 72.8411
R15444 gnd.n2911 gnd.n2896 72.8411
R15445 gnd.n3191 gnd.n3190 72.8411
R15446 gnd.n2797 gnd.t128 72.836
R15447 gnd.n2930 gnd.t121 72.836
R15448 gnd.n3218 gnd.t115 72.836
R15449 gnd.n7332 gnd.t144 72.836
R15450 gnd.n1692 gnd.t137 72.836
R15451 gnd.n2224 gnd.t160 72.836
R15452 gnd.n1470 gnd.t110 72.836
R15453 gnd.n1492 gnd.t100 72.836
R15454 gnd.n180 gnd.t174 72.836
R15455 gnd.n7425 gnd.t97 72.836
R15456 gnd.n984 gnd.t74 72.836
R15457 gnd.n1006 gnd.t153 72.836
R15458 gnd.n2313 gnd.t171 72.836
R15459 gnd.n2291 gnd.t89 72.836
R15460 gnd.n2478 gnd.t103 72.836
R15461 gnd.n4144 gnd.t85 72.836
R15462 gnd.n3374 gnd.n3373 71.676
R15463 gnd.n3371 gnd.n3370 71.676
R15464 gnd.n3366 gnd.n3200 71.676
R15465 gnd.n3364 gnd.n3363 71.676
R15466 gnd.n3359 gnd.n3203 71.676
R15467 gnd.n3357 gnd.n3356 71.676
R15468 gnd.n3352 gnd.n3206 71.676
R15469 gnd.n3350 gnd.n3349 71.676
R15470 gnd.n3345 gnd.n3209 71.676
R15471 gnd.n3343 gnd.n3342 71.676
R15472 gnd.n3338 gnd.n3212 71.676
R15473 gnd.n3336 gnd.n3335 71.676
R15474 gnd.n3331 gnd.n3215 71.676
R15475 gnd.n3329 gnd.n3328 71.676
R15476 gnd.n3323 gnd.n3220 71.676
R15477 gnd.n3321 gnd.n3320 71.676
R15478 gnd.n3316 gnd.n3315 71.676
R15479 gnd.n3313 gnd.n3312 71.676
R15480 gnd.n3307 gnd.n3226 71.676
R15481 gnd.n3305 gnd.n3304 71.676
R15482 gnd.n3300 gnd.n3229 71.676
R15483 gnd.n3298 gnd.n3297 71.676
R15484 gnd.n3293 gnd.n3232 71.676
R15485 gnd.n3291 gnd.n3290 71.676
R15486 gnd.n3286 gnd.n3235 71.676
R15487 gnd.n3284 gnd.n3283 71.676
R15488 gnd.n3279 gnd.n3238 71.676
R15489 gnd.n3277 gnd.n3276 71.676
R15490 gnd.n3272 gnd.n3241 71.676
R15491 gnd.n3270 gnd.n3269 71.676
R15492 gnd.n3265 gnd.n3244 71.676
R15493 gnd.n3263 gnd.n3262 71.676
R15494 gnd.n3258 gnd.n3247 71.676
R15495 gnd.n2992 gnd.n2893 71.676
R15496 gnd.n2990 gnd.n2916 71.676
R15497 gnd.n2986 gnd.n2985 71.676
R15498 gnd.n2979 gnd.n2918 71.676
R15499 gnd.n2978 gnd.n2977 71.676
R15500 gnd.n2971 gnd.n2920 71.676
R15501 gnd.n2970 gnd.n2969 71.676
R15502 gnd.n2963 gnd.n2922 71.676
R15503 gnd.n2962 gnd.n2961 71.676
R15504 gnd.n2955 gnd.n2924 71.676
R15505 gnd.n2954 gnd.n2953 71.676
R15506 gnd.n2947 gnd.n2926 71.676
R15507 gnd.n2946 gnd.n2945 71.676
R15508 gnd.n2939 gnd.n2928 71.676
R15509 gnd.n2938 gnd.n2932 71.676
R15510 gnd.n2934 gnd.n2933 71.676
R15511 gnd.n3637 gnd.n3636 71.676
R15512 gnd.n3629 gnd.n2873 71.676
R15513 gnd.n3628 gnd.n3627 71.676
R15514 gnd.n3621 gnd.n2877 71.676
R15515 gnd.n3620 gnd.n3619 71.676
R15516 gnd.n3613 gnd.n2879 71.676
R15517 gnd.n3612 gnd.n3611 71.676
R15518 gnd.n3605 gnd.n2881 71.676
R15519 gnd.n3604 gnd.n3603 71.676
R15520 gnd.n3597 gnd.n2883 71.676
R15521 gnd.n3596 gnd.n3595 71.676
R15522 gnd.n3589 gnd.n2885 71.676
R15523 gnd.n3588 gnd.n3587 71.676
R15524 gnd.n3581 gnd.n2887 71.676
R15525 gnd.n3580 gnd.n3579 71.676
R15526 gnd.n3573 gnd.n2889 71.676
R15527 gnd.n2993 gnd.n2992 71.676
R15528 gnd.n2987 gnd.n2916 71.676
R15529 gnd.n2985 gnd.n2984 71.676
R15530 gnd.n2980 gnd.n2979 71.676
R15531 gnd.n2977 gnd.n2976 71.676
R15532 gnd.n2972 gnd.n2971 71.676
R15533 gnd.n2969 gnd.n2968 71.676
R15534 gnd.n2964 gnd.n2963 71.676
R15535 gnd.n2961 gnd.n2960 71.676
R15536 gnd.n2956 gnd.n2955 71.676
R15537 gnd.n2953 gnd.n2952 71.676
R15538 gnd.n2948 gnd.n2947 71.676
R15539 gnd.n2945 gnd.n2944 71.676
R15540 gnd.n2940 gnd.n2939 71.676
R15541 gnd.n2935 gnd.n2932 71.676
R15542 gnd.n3639 gnd.n3638 71.676
R15543 gnd.n3636 gnd.n3635 71.676
R15544 gnd.n3630 gnd.n3629 71.676
R15545 gnd.n3627 gnd.n3626 71.676
R15546 gnd.n3622 gnd.n3621 71.676
R15547 gnd.n3619 gnd.n3618 71.676
R15548 gnd.n3614 gnd.n3613 71.676
R15549 gnd.n3611 gnd.n3610 71.676
R15550 gnd.n3606 gnd.n3605 71.676
R15551 gnd.n3603 gnd.n3602 71.676
R15552 gnd.n3598 gnd.n3597 71.676
R15553 gnd.n3595 gnd.n3594 71.676
R15554 gnd.n3590 gnd.n3589 71.676
R15555 gnd.n3587 gnd.n3586 71.676
R15556 gnd.n3582 gnd.n3581 71.676
R15557 gnd.n3579 gnd.n3578 71.676
R15558 gnd.n3574 gnd.n3573 71.676
R15559 gnd.n3247 gnd.n3245 71.676
R15560 gnd.n3264 gnd.n3263 71.676
R15561 gnd.n3244 gnd.n3242 71.676
R15562 gnd.n3271 gnd.n3270 71.676
R15563 gnd.n3241 gnd.n3239 71.676
R15564 gnd.n3278 gnd.n3277 71.676
R15565 gnd.n3238 gnd.n3236 71.676
R15566 gnd.n3285 gnd.n3284 71.676
R15567 gnd.n3235 gnd.n3233 71.676
R15568 gnd.n3292 gnd.n3291 71.676
R15569 gnd.n3232 gnd.n3230 71.676
R15570 gnd.n3299 gnd.n3298 71.676
R15571 gnd.n3229 gnd.n3227 71.676
R15572 gnd.n3306 gnd.n3305 71.676
R15573 gnd.n3226 gnd.n3222 71.676
R15574 gnd.n3314 gnd.n3313 71.676
R15575 gnd.n3318 gnd.n3317 71.676
R15576 gnd.n3322 gnd.n3321 71.676
R15577 gnd.n3220 gnd.n3216 71.676
R15578 gnd.n3330 gnd.n3329 71.676
R15579 gnd.n3215 gnd.n3213 71.676
R15580 gnd.n3337 gnd.n3336 71.676
R15581 gnd.n3212 gnd.n3210 71.676
R15582 gnd.n3344 gnd.n3343 71.676
R15583 gnd.n3209 gnd.n3207 71.676
R15584 gnd.n3351 gnd.n3350 71.676
R15585 gnd.n3206 gnd.n3204 71.676
R15586 gnd.n3358 gnd.n3357 71.676
R15587 gnd.n3203 gnd.n3201 71.676
R15588 gnd.n3365 gnd.n3364 71.676
R15589 gnd.n3200 gnd.n3198 71.676
R15590 gnd.n3372 gnd.n3371 71.676
R15591 gnd.n3375 gnd.n3374 71.676
R15592 gnd.n10 gnd.t323 69.1507
R15593 gnd.n18 gnd.t17 68.4792
R15594 gnd.n17 gnd.t46 68.4792
R15595 gnd.n16 gnd.t60 68.4792
R15596 gnd.n15 gnd.t304 68.4792
R15597 gnd.n14 gnd.t31 68.4792
R15598 gnd.n13 gnd.t11 68.4792
R15599 gnd.n12 gnd.t39 68.4792
R15600 gnd.n11 gnd.t328 68.4792
R15601 gnd.n10 gnd.t62 68.4792
R15602 gnd.n5340 gnd.n5244 64.369
R15603 gnd.n3632 gnd.n2875 59.5399
R15604 gnd.n3309 gnd.n3224 59.5399
R15605 gnd.n2931 gnd.n2930 59.5399
R15606 gnd.n3325 gnd.n3218 59.5399
R15607 gnd.n2996 gnd.n2914 59.1804
R15608 gnd.n6236 gnd.n4833 57.3586
R15609 gnd.n4832 gnd.n961 57.3586
R15610 gnd.n7461 gnd.n106 57.3586
R15611 gnd.n5446 gnd.t204 56.607
R15612 gnd.n52 gnd.t299 56.607
R15613 gnd.n5415 gnd.t238 56.407
R15614 gnd.n5430 gnd.t217 56.407
R15615 gnd.n21 gnd.t272 56.407
R15616 gnd.n36 gnd.t250 56.407
R15617 gnd.n5459 gnd.t292 55.8337
R15618 gnd.n5428 gnd.t275 55.8337
R15619 gnd.n5443 gnd.t252 55.8337
R15620 gnd.n65 gnd.t231 55.8337
R15621 gnd.n34 gnd.t280 55.8337
R15622 gnd.n49 gnd.t265 55.8337
R15623 gnd.n2902 gnd.n2901 54.358
R15624 gnd.n3188 gnd.n3187 54.358
R15625 gnd.n5446 gnd.n5445 53.0052
R15626 gnd.n5448 gnd.n5447 53.0052
R15627 gnd.n5450 gnd.n5449 53.0052
R15628 gnd.n5452 gnd.n5451 53.0052
R15629 gnd.n5454 gnd.n5453 53.0052
R15630 gnd.n5456 gnd.n5455 53.0052
R15631 gnd.n5458 gnd.n5457 53.0052
R15632 gnd.n5415 gnd.n5414 53.0052
R15633 gnd.n5417 gnd.n5416 53.0052
R15634 gnd.n5419 gnd.n5418 53.0052
R15635 gnd.n5421 gnd.n5420 53.0052
R15636 gnd.n5423 gnd.n5422 53.0052
R15637 gnd.n5425 gnd.n5424 53.0052
R15638 gnd.n5427 gnd.n5426 53.0052
R15639 gnd.n5430 gnd.n5429 53.0052
R15640 gnd.n5432 gnd.n5431 53.0052
R15641 gnd.n5434 gnd.n5433 53.0052
R15642 gnd.n5436 gnd.n5435 53.0052
R15643 gnd.n5438 gnd.n5437 53.0052
R15644 gnd.n5440 gnd.n5439 53.0052
R15645 gnd.n5442 gnd.n5441 53.0052
R15646 gnd.n64 gnd.n63 53.0052
R15647 gnd.n62 gnd.n61 53.0052
R15648 gnd.n60 gnd.n59 53.0052
R15649 gnd.n58 gnd.n57 53.0052
R15650 gnd.n56 gnd.n55 53.0052
R15651 gnd.n54 gnd.n53 53.0052
R15652 gnd.n52 gnd.n51 53.0052
R15653 gnd.n33 gnd.n32 53.0052
R15654 gnd.n31 gnd.n30 53.0052
R15655 gnd.n29 gnd.n28 53.0052
R15656 gnd.n27 gnd.n26 53.0052
R15657 gnd.n25 gnd.n24 53.0052
R15658 gnd.n23 gnd.n22 53.0052
R15659 gnd.n21 gnd.n20 53.0052
R15660 gnd.n48 gnd.n47 53.0052
R15661 gnd.n46 gnd.n45 53.0052
R15662 gnd.n44 gnd.n43 53.0052
R15663 gnd.n42 gnd.n41 53.0052
R15664 gnd.n40 gnd.n39 53.0052
R15665 gnd.n38 gnd.n37 53.0052
R15666 gnd.n36 gnd.n35 53.0052
R15667 gnd.n3179 gnd.n3178 52.4801
R15668 gnd.n6063 gnd.t58 52.3082
R15669 gnd.n6031 gnd.t330 52.3082
R15670 gnd.n5999 gnd.t22 52.3082
R15671 gnd.n5968 gnd.t27 52.3082
R15672 gnd.n5936 gnd.t37 52.3082
R15673 gnd.n5904 gnd.t42 52.3082
R15674 gnd.n5872 gnd.t64 52.3082
R15675 gnd.n5841 gnd.t326 52.3082
R15676 gnd.n5893 gnd.n5861 51.4173
R15677 gnd.n5957 gnd.n5956 50.455
R15678 gnd.n5925 gnd.n5924 50.455
R15679 gnd.n5893 gnd.n5892 50.455
R15680 gnd.n5287 gnd.n5286 45.1884
R15681 gnd.n4908 gnd.n4907 45.1884
R15682 gnd.n3377 gnd.n3194 44.3322
R15683 gnd.n2905 gnd.n2904 44.3189
R15684 gnd.n2798 gnd.n2797 42.4732
R15685 gnd.n4145 gnd.n4144 42.4732
R15686 gnd.n5288 gnd.n5287 42.2793
R15687 gnd.n4909 gnd.n4908 42.2793
R15688 gnd.n5214 gnd.n5213 42.2793
R15689 gnd.n4865 gnd.n4864 42.2793
R15690 gnd.n7337 gnd.n7332 42.2793
R15691 gnd.n1799 gnd.n1692 42.2793
R15692 gnd.n2225 gnd.n2224 42.2793
R15693 gnd.n1493 gnd.n1492 42.2793
R15694 gnd.n7389 gnd.n180 42.2793
R15695 gnd.n7426 gnd.n7425 42.2793
R15696 gnd.n4796 gnd.n984 42.2793
R15697 gnd.n1007 gnd.n1006 42.2793
R15698 gnd.n2828 gnd.n2313 42.2793
R15699 gnd.n2479 gnd.n2478 42.2793
R15700 gnd.n2903 gnd.n2902 41.6274
R15701 gnd.n3189 gnd.n3188 41.6274
R15702 gnd.n2912 gnd.n2911 40.8975
R15703 gnd.n3192 gnd.n3191 40.8975
R15704 gnd.n4393 gnd.n1470 36.9518
R15705 gnd.n3641 gnd.n2291 36.9518
R15706 gnd.n6426 gnd.n6425 36.594
R15707 gnd.n6425 gnd.n728 36.594
R15708 gnd.n6419 gnd.n728 36.594
R15709 gnd.n6419 gnd.n6418 36.594
R15710 gnd.n6418 gnd.n6417 36.594
R15711 gnd.n6417 gnd.n736 36.594
R15712 gnd.n6411 gnd.n736 36.594
R15713 gnd.n6411 gnd.n6410 36.594
R15714 gnd.n6410 gnd.n6409 36.594
R15715 gnd.n6409 gnd.n744 36.594
R15716 gnd.n6403 gnd.n744 36.594
R15717 gnd.n6403 gnd.n6402 36.594
R15718 gnd.n6402 gnd.n6401 36.594
R15719 gnd.n6401 gnd.n752 36.594
R15720 gnd.n6395 gnd.n752 36.594
R15721 gnd.n6395 gnd.n6394 36.594
R15722 gnd.n6394 gnd.n6393 36.594
R15723 gnd.n6393 gnd.n760 36.594
R15724 gnd.n6387 gnd.n760 36.594
R15725 gnd.n6387 gnd.n6386 36.594
R15726 gnd.n6386 gnd.n6385 36.594
R15727 gnd.n6385 gnd.n768 36.594
R15728 gnd.n6379 gnd.n768 36.594
R15729 gnd.n6379 gnd.n6378 36.594
R15730 gnd.n6378 gnd.n6377 36.594
R15731 gnd.n6377 gnd.n776 36.594
R15732 gnd.n6371 gnd.n776 36.594
R15733 gnd.n6371 gnd.n6370 36.594
R15734 gnd.n6370 gnd.n6369 36.594
R15735 gnd.n6369 gnd.n784 36.594
R15736 gnd.n6363 gnd.n784 36.594
R15737 gnd.n6363 gnd.n6362 36.594
R15738 gnd.n6362 gnd.n6361 36.594
R15739 gnd.n6361 gnd.n792 36.594
R15740 gnd.n6355 gnd.n792 36.594
R15741 gnd.n6355 gnd.n6354 36.594
R15742 gnd.n6354 gnd.n6353 36.594
R15743 gnd.n6353 gnd.n800 36.594
R15744 gnd.n6347 gnd.n800 36.594
R15745 gnd.n6347 gnd.n6346 36.594
R15746 gnd.n6346 gnd.n6345 36.594
R15747 gnd.n6345 gnd.n808 36.594
R15748 gnd.n6339 gnd.n808 36.594
R15749 gnd.n6339 gnd.n6338 36.594
R15750 gnd.n6338 gnd.n6337 36.594
R15751 gnd.n6337 gnd.n816 36.594
R15752 gnd.n6331 gnd.n816 36.594
R15753 gnd.n6331 gnd.n6330 36.594
R15754 gnd.n6330 gnd.n6329 36.594
R15755 gnd.n6329 gnd.n824 36.594
R15756 gnd.n6323 gnd.n824 36.594
R15757 gnd.n6323 gnd.n6322 36.594
R15758 gnd.n6322 gnd.n6321 36.594
R15759 gnd.n6321 gnd.n832 36.594
R15760 gnd.n6315 gnd.n832 36.594
R15761 gnd.n6315 gnd.n6314 36.594
R15762 gnd.n6314 gnd.n6313 36.594
R15763 gnd.n6313 gnd.n840 36.594
R15764 gnd.n6307 gnd.n840 36.594
R15765 gnd.n6307 gnd.n6306 36.594
R15766 gnd.n6306 gnd.n6305 36.594
R15767 gnd.n6305 gnd.n848 36.594
R15768 gnd.n6299 gnd.n848 36.594
R15769 gnd.n6299 gnd.n6298 36.594
R15770 gnd.n6298 gnd.n6297 36.594
R15771 gnd.n6297 gnd.n856 36.594
R15772 gnd.n6291 gnd.n856 36.594
R15773 gnd.n6291 gnd.n6290 36.594
R15774 gnd.n6290 gnd.n6289 36.594
R15775 gnd.n6289 gnd.n864 36.594
R15776 gnd.n6283 gnd.n864 36.594
R15777 gnd.n6283 gnd.n6282 36.594
R15778 gnd.n6282 gnd.n6281 36.594
R15779 gnd.n6281 gnd.n872 36.594
R15780 gnd.n6275 gnd.n872 36.594
R15781 gnd.n6275 gnd.n6274 36.594
R15782 gnd.n6274 gnd.n6273 36.594
R15783 gnd.n6273 gnd.n880 36.594
R15784 gnd.n6267 gnd.n880 36.594
R15785 gnd.n6267 gnd.n6266 36.594
R15786 gnd.n6266 gnd.n6265 36.594
R15787 gnd.n6265 gnd.n888 36.594
R15788 gnd.n6259 gnd.n888 36.594
R15789 gnd.n2911 gnd.n2910 35.055
R15790 gnd.n2906 gnd.n2905 35.055
R15791 gnd.n3181 gnd.n3180 35.055
R15792 gnd.n3191 gnd.n3177 35.055
R15793 gnd.n5350 gnd.n5244 31.8661
R15794 gnd.n5350 gnd.n5349 31.8661
R15795 gnd.n5358 gnd.n5233 31.8661
R15796 gnd.n5366 gnd.n5233 31.8661
R15797 gnd.n5366 gnd.n5227 31.8661
R15798 gnd.n5374 gnd.n5227 31.8661
R15799 gnd.n5374 gnd.n5220 31.8661
R15800 gnd.n5498 gnd.n5220 31.8661
R15801 gnd.n5508 gnd.n5153 31.8661
R15802 gnd.n2535 gnd.n961 31.8661
R15803 gnd.n4745 gnd.n1015 31.8661
R15804 gnd.n4745 gnd.n1017 31.8661
R15805 gnd.n4739 gnd.n1017 31.8661
R15806 gnd.n4739 gnd.n1029 31.8661
R15807 gnd.n4733 gnd.n1040 31.8661
R15808 gnd.n4727 gnd.n1040 31.8661
R15809 gnd.n4721 gnd.n1057 31.8661
R15810 gnd.n4715 gnd.n1067 31.8661
R15811 gnd.n4715 gnd.n1070 31.8661
R15812 gnd.n4709 gnd.n1080 31.8661
R15813 gnd.n4703 gnd.n1080 31.8661
R15814 gnd.n4697 gnd.n1098 31.8661
R15815 gnd.n2234 gnd.n1273 31.8661
R15816 gnd.n2745 gnd.n2250 31.8661
R15817 gnd.n2745 gnd.n2165 31.8661
R15818 gnd.n2178 gnd.n2159 31.8661
R15819 gnd.n3729 gnd.n2159 31.8661
R15820 gnd.n3737 gnd.n2152 31.8661
R15821 gnd.n3737 gnd.n2145 31.8661
R15822 gnd.n3745 gnd.n2145 31.8661
R15823 gnd.n3745 gnd.n2146 31.8661
R15824 gnd.n3753 gnd.n2133 31.8661
R15825 gnd.n3761 gnd.n2133 31.8661
R15826 gnd.n3761 gnd.n2126 31.8661
R15827 gnd.n3769 gnd.n2126 31.8661
R15828 gnd.n3777 gnd.n2120 31.8661
R15829 gnd.n3777 gnd.n2113 31.8661
R15830 gnd.n3785 gnd.n2113 31.8661
R15831 gnd.n3793 gnd.n2107 31.8661
R15832 gnd.n3793 gnd.n2099 31.8661
R15833 gnd.n3801 gnd.n2099 31.8661
R15834 gnd.n3801 gnd.n2101 31.8661
R15835 gnd.n3809 gnd.n2093 31.8661
R15836 gnd.n4041 gnd.n1890 31.8661
R15837 gnd.n4049 gnd.n1877 31.8661
R15838 gnd.n4057 gnd.n1877 31.8661
R15839 gnd.n4057 gnd.n1871 31.8661
R15840 gnd.n4065 gnd.n1871 31.8661
R15841 gnd.n4073 gnd.n1864 31.8661
R15842 gnd.n4073 gnd.n1858 31.8661
R15843 gnd.n4081 gnd.n1858 31.8661
R15844 gnd.n4089 gnd.n1851 31.8661
R15845 gnd.n4089 gnd.n1844 31.8661
R15846 gnd.n4097 gnd.n1844 31.8661
R15847 gnd.n4097 gnd.n1845 31.8661
R15848 gnd.n4105 gnd.n1831 31.8661
R15849 gnd.n4115 gnd.n1831 31.8661
R15850 gnd.n4115 gnd.n1823 31.8661
R15851 gnd.n4126 gnd.n1823 31.8661
R15852 gnd.n4434 gnd.n1406 31.8661
R15853 gnd.n4434 gnd.n4433 31.8661
R15854 gnd.n4427 gnd.n1417 31.8661
R15855 gnd.n4427 gnd.n4426 31.8661
R15856 gnd.n1497 gnd.n1446 31.8661
R15857 gnd.n7242 gnd.n248 31.8661
R15858 gnd.n7250 gnd.n238 31.8661
R15859 gnd.n7250 gnd.n241 31.8661
R15860 gnd.n7258 gnd.n225 31.8661
R15861 gnd.n7266 gnd.n225 31.8661
R15862 gnd.n7274 gnd.n218 31.8661
R15863 gnd.n7282 gnd.n208 31.8661
R15864 gnd.n7282 gnd.n211 31.8661
R15865 gnd.n7290 gnd.n193 31.8661
R15866 gnd.n7373 gnd.n193 31.8661
R15867 gnd.n7373 gnd.n185 31.8661
R15868 gnd.n7381 gnd.n185 31.8661
R15869 gnd.n7461 gnd.n104 31.8661
R15870 gnd.n3259 gnd.n3246 29.8151
R15871 gnd.n3575 gnd.n2890 29.8151
R15872 gnd.n4721 gnd.t179 27.7236
R15873 gnd.t218 gnd.n218 27.7236
R15874 gnd.n3785 gnd.t12 27.0862
R15875 gnd.t45 gnd.n1864 27.0862
R15876 gnd.n3817 gnd.n2086 26.4489
R15877 gnd.n3255 gnd.n3196 26.4489
R15878 gnd.n2797 gnd.n2796 25.7944
R15879 gnd.n5213 gnd.n5212 25.7944
R15880 gnd.n4864 gnd.n4863 25.7944
R15881 gnd.n7332 gnd.n7331 25.7944
R15882 gnd.n1692 gnd.n1691 25.7944
R15883 gnd.n2224 gnd.n2223 25.7944
R15884 gnd.n1470 gnd.n1469 25.7944
R15885 gnd.n1492 gnd.n1491 25.7944
R15886 gnd.n180 gnd.n179 25.7944
R15887 gnd.n7425 gnd.n7424 25.7944
R15888 gnd.n984 gnd.n983 25.7944
R15889 gnd.n1006 gnd.n1005 25.7944
R15890 gnd.n2313 gnd.n2312 25.7944
R15891 gnd.n2291 gnd.n2290 25.7944
R15892 gnd.n2478 gnd.n2477 25.7944
R15893 gnd.n4144 gnd.n4143 25.7944
R15894 gnd.n1057 gnd.t269 25.1743
R15895 gnd.n7274 gnd.t214 25.1743
R15896 gnd.n5520 gnd.n5154 24.8557
R15897 gnd.n5530 gnd.n5137 24.8557
R15898 gnd.n5140 gnd.n5128 24.8557
R15899 gnd.n5551 gnd.n5129 24.8557
R15900 gnd.n5561 gnd.n5111 24.8557
R15901 gnd.n5572 gnd.n5571 24.8557
R15902 gnd.n5591 gnd.n5097 24.8557
R15903 gnd.n5592 gnd.n5086 24.8557
R15904 gnd.n5603 gnd.n5602 24.8557
R15905 gnd.n5613 gnd.n5079 24.8557
R15906 gnd.n5622 gnd.n5071 24.8557
R15907 gnd.n5634 gnd.n5633 24.8557
R15908 gnd.n5409 gnd.n5063 24.8557
R15909 gnd.n5644 gnd.n5053 24.8557
R15910 gnd.n5653 gnd.n5046 24.8557
R15911 gnd.n5039 gnd.n5029 24.8557
R15912 gnd.n5022 gnd.n5016 24.8557
R15913 gnd.n5708 gnd.n5707 24.8557
R15914 gnd.n5718 gnd.n5717 24.8557
R15915 gnd.n5007 gnd.n4999 24.8557
R15916 gnd.n5729 gnd.n4984 24.8557
R15917 gnd.n5748 gnd.n5747 24.8557
R15918 gnd.n5758 gnd.n4977 24.8557
R15919 gnd.n5771 gnd.n4966 24.8557
R15920 gnd.n5762 gnd.n5761 24.8557
R15921 gnd.n5794 gnd.n5793 24.8557
R15922 gnd.n5804 gnd.n4953 24.8557
R15923 gnd.n5816 gnd.n4945 24.8557
R15924 gnd.n6115 gnd.n6114 24.8557
R15925 gnd.n6130 gnd.n6129 24.8557
R15926 gnd.n6251 gnd.n907 24.8557
R15927 gnd.n6250 gnd.n910 24.8557
R15928 gnd.n6099 gnd.n919 24.8557
R15929 gnd.n6237 gnd.n930 24.8557
R15930 gnd.n3729 gnd.t127 24.537
R15931 gnd.t322 gnd.n2120 24.537
R15932 gnd.n4081 gnd.t33 24.537
R15933 gnd.t83 gnd.n1406 24.537
R15934 gnd.n3720 gnd.n2178 23.8997
R15935 gnd.n4433 gnd.n1409 23.8997
R15936 gnd.n5541 gnd.t325 23.2624
R15937 gnd.n5156 gnd.t149 22.6251
R15938 gnd.n2535 gnd.t73 22.6251
R15939 gnd.t95 gnd.n104 22.6251
R15940 gnd.n6259 gnd.n6258 21.9566
R15941 gnd.n3571 gnd.n2892 21.6691
R15942 gnd.n3538 gnd.n2051 21.6691
R15943 gnd.n3523 gnd.n3522 21.6691
R15944 gnd.n3509 gnd.n2023 21.6691
R15945 gnd.n3487 gnd.n2002 21.6691
R15946 gnd.n3480 gnd.n1995 21.6691
R15947 gnd.n3472 gnd.n1989 21.6691
R15948 gnd.n3465 gnd.n1981 21.6691
R15949 gnd.n3437 gnd.n3127 21.6691
R15950 gnd.n3424 gnd.n1938 21.6691
R15951 gnd.n3409 gnd.n1925 21.6691
R15952 gnd.t26 gnd.n5161 21.3504
R15953 gnd.n3565 gnd.n2999 21.0318
R15954 gnd.n3005 gnd.n3004 21.0318
R15955 gnd.n3889 gnd.n2025 21.0318
R15956 gnd.n3897 gnd.n2015 21.0318
R15957 gnd.n3449 gnd.n1959 21.0318
R15958 gnd.n3443 gnd.n3122 21.0318
R15959 gnd.n4025 gnd.t131 21.0318
R15960 gnd.n4033 gnd.n1896 21.0318
R15961 gnd.t308 gnd.n4930 20.7131
R15962 gnd.n1097 gnd.t198 20.3945
R15963 gnd.n250 gnd.t235 20.3945
R15964 gnd.t310 gnd.n4976 20.0758
R15965 gnd.n2899 gnd.t125 19.8005
R15966 gnd.n2899 gnd.t147 19.8005
R15967 gnd.n2900 gnd.t141 19.8005
R15968 gnd.n2900 gnd.t162 19.8005
R15969 gnd.n3185 gnd.t78 19.8005
R15970 gnd.n3185 gnd.t135 19.8005
R15971 gnd.n3186 gnd.t157 19.8005
R15972 gnd.n3186 gnd.t132 19.8005
R15973 gnd.n3670 gnd.n2250 19.7572
R15974 gnd.n3009 gnd.n2075 19.7572
R15975 gnd.n3881 gnd.n2032 19.7572
R15976 gnd.n3905 gnd.n2008 19.7572
R15977 gnd.n3109 gnd.n1966 19.7572
R15978 gnd.n3131 gnd.n1953 19.7572
R15979 gnd.n4017 gnd.n1912 19.7572
R15980 gnd.n4426 gnd.n4425 19.7572
R15981 gnd.n2896 gnd.n2895 19.5087
R15982 gnd.n2909 gnd.n2896 19.5087
R15983 gnd.n2907 gnd.n2898 19.5087
R15984 gnd.n3190 gnd.n3184 19.5087
R15985 gnd.n5684 gnd.t314 19.4385
R15986 gnd.n2146 gnd.t14 19.4385
R15987 gnd.n4105 gnd.t16 19.4385
R15988 gnd.n3727 gnd.n2161 19.3944
R15989 gnd.n3727 gnd.n2150 19.3944
R15990 gnd.n3739 gnd.n2150 19.3944
R15991 gnd.n3739 gnd.n2148 19.3944
R15992 gnd.n3743 gnd.n2148 19.3944
R15993 gnd.n3743 gnd.n2137 19.3944
R15994 gnd.n3755 gnd.n2137 19.3944
R15995 gnd.n3755 gnd.n2135 19.3944
R15996 gnd.n3759 gnd.n2135 19.3944
R15997 gnd.n3759 gnd.n2124 19.3944
R15998 gnd.n3771 gnd.n2124 19.3944
R15999 gnd.n3771 gnd.n2122 19.3944
R16000 gnd.n3775 gnd.n2122 19.3944
R16001 gnd.n3775 gnd.n2111 19.3944
R16002 gnd.n3787 gnd.n2111 19.3944
R16003 gnd.n3787 gnd.n2109 19.3944
R16004 gnd.n3791 gnd.n2109 19.3944
R16005 gnd.n3791 gnd.n2097 19.3944
R16006 gnd.n3803 gnd.n2097 19.3944
R16007 gnd.n3803 gnd.n2095 19.3944
R16008 gnd.n3807 gnd.n2095 19.3944
R16009 gnd.n3807 gnd.n2084 19.3944
R16010 gnd.n3819 gnd.n2084 19.3944
R16011 gnd.n3819 gnd.n2082 19.3944
R16012 gnd.n3823 gnd.n2082 19.3944
R16013 gnd.n3823 gnd.n2071 19.3944
R16014 gnd.n3835 gnd.n2071 19.3944
R16015 gnd.n3835 gnd.n2069 19.3944
R16016 gnd.n3839 gnd.n2069 19.3944
R16017 gnd.n3839 gnd.n2056 19.3944
R16018 gnd.n3851 gnd.n2056 19.3944
R16019 gnd.n3851 gnd.n2054 19.3944
R16020 gnd.n3855 gnd.n2054 19.3944
R16021 gnd.n3855 gnd.n2042 19.3944
R16022 gnd.n3867 gnd.n2042 19.3944
R16023 gnd.n3867 gnd.n2040 19.3944
R16024 gnd.n3871 gnd.n2040 19.3944
R16025 gnd.n3871 gnd.n2029 19.3944
R16026 gnd.n3883 gnd.n2029 19.3944
R16027 gnd.n3883 gnd.n2027 19.3944
R16028 gnd.n3887 gnd.n2027 19.3944
R16029 gnd.n3887 gnd.n2013 19.3944
R16030 gnd.n3899 gnd.n2013 19.3944
R16031 gnd.n3899 gnd.n2011 19.3944
R16032 gnd.n3903 gnd.n2011 19.3944
R16033 gnd.n3903 gnd.n1999 19.3944
R16034 gnd.n3915 gnd.n1999 19.3944
R16035 gnd.n3915 gnd.n1997 19.3944
R16036 gnd.n3919 gnd.n1997 19.3944
R16037 gnd.n3919 gnd.n1985 19.3944
R16038 gnd.n3931 gnd.n1985 19.3944
R16039 gnd.n3931 gnd.n1983 19.3944
R16040 gnd.n3935 gnd.n1983 19.3944
R16041 gnd.n3935 gnd.n1971 19.3944
R16042 gnd.n3947 gnd.n1971 19.3944
R16043 gnd.n3947 gnd.n1969 19.3944
R16044 gnd.n3951 gnd.n1969 19.3944
R16045 gnd.n3951 gnd.n1957 19.3944
R16046 gnd.n3963 gnd.n1957 19.3944
R16047 gnd.n3963 gnd.n1955 19.3944
R16048 gnd.n3967 gnd.n1955 19.3944
R16049 gnd.n3967 gnd.n1943 19.3944
R16050 gnd.n3979 gnd.n1943 19.3944
R16051 gnd.n3979 gnd.n1941 19.3944
R16052 gnd.n3983 gnd.n1941 19.3944
R16053 gnd.n3983 gnd.n1929 19.3944
R16054 gnd.n3995 gnd.n1929 19.3944
R16055 gnd.n3995 gnd.n1927 19.3944
R16056 gnd.n3999 gnd.n1927 19.3944
R16057 gnd.n3999 gnd.n1916 19.3944
R16058 gnd.n4011 gnd.n1916 19.3944
R16059 gnd.n4011 gnd.n1914 19.3944
R16060 gnd.n4015 gnd.n1914 19.3944
R16061 gnd.n4015 gnd.n1901 19.3944
R16062 gnd.n4027 gnd.n1901 19.3944
R16063 gnd.n4027 gnd.n1899 19.3944
R16064 gnd.n4031 gnd.n1899 19.3944
R16065 gnd.n4031 gnd.n1887 19.3944
R16066 gnd.n4043 gnd.n1887 19.3944
R16067 gnd.n4043 gnd.n1885 19.3944
R16068 gnd.n4047 gnd.n1885 19.3944
R16069 gnd.n4047 gnd.n1875 19.3944
R16070 gnd.n4059 gnd.n1875 19.3944
R16071 gnd.n4059 gnd.n1873 19.3944
R16072 gnd.n4063 gnd.n1873 19.3944
R16073 gnd.n4063 gnd.n1862 19.3944
R16074 gnd.n4075 gnd.n1862 19.3944
R16075 gnd.n4075 gnd.n1860 19.3944
R16076 gnd.n4079 gnd.n1860 19.3944
R16077 gnd.n4079 gnd.n1849 19.3944
R16078 gnd.n4091 gnd.n1849 19.3944
R16079 gnd.n4091 gnd.n1847 19.3944
R16080 gnd.n4095 gnd.n1847 19.3944
R16081 gnd.n4095 gnd.n1836 19.3944
R16082 gnd.n4107 gnd.n1836 19.3944
R16083 gnd.n4107 gnd.n1833 19.3944
R16084 gnd.n4113 gnd.n1833 19.3944
R16085 gnd.n4113 gnd.n1834 19.3944
R16086 gnd.n1834 gnd.n1821 19.3944
R16087 gnd.n4129 gnd.n1821 19.3944
R16088 gnd.n4130 gnd.n4129 19.3944
R16089 gnd.n2803 gnd.n2802 19.3944
R16090 gnd.n2802 gnd.n2163 19.3944
R16091 gnd.n3723 gnd.n2163 19.3944
R16092 gnd.n3717 gnd.n3716 19.3944
R16093 gnd.n3716 gnd.n2182 19.3944
R16094 gnd.n3709 gnd.n2182 19.3944
R16095 gnd.n3709 gnd.n3708 19.3944
R16096 gnd.n3708 gnd.n2193 19.3944
R16097 gnd.n3701 gnd.n2193 19.3944
R16098 gnd.n3701 gnd.n3700 19.3944
R16099 gnd.n3700 gnd.n2201 19.3944
R16100 gnd.n3693 gnd.n2201 19.3944
R16101 gnd.n3693 gnd.n3692 19.3944
R16102 gnd.n3692 gnd.n2211 19.3944
R16103 gnd.n3685 gnd.n2211 19.3944
R16104 gnd.n3685 gnd.n3684 19.3944
R16105 gnd.n3684 gnd.n2219 19.3944
R16106 gnd.n3677 gnd.n2219 19.3944
R16107 gnd.n3677 gnd.n3676 19.3944
R16108 gnd.n3676 gnd.n2231 19.3944
R16109 gnd.n2814 gnd.n2231 19.3944
R16110 gnd.n2814 gnd.n2813 19.3944
R16111 gnd.n2813 gnd.n2812 19.3944
R16112 gnd.n2812 gnd.n2791 19.3944
R16113 gnd.n2808 gnd.n2791 19.3944
R16114 gnd.n2808 gnd.n2807 19.3944
R16115 gnd.n2807 gnd.n2806 19.3944
R16116 gnd.n5337 gnd.n5336 19.3944
R16117 gnd.n5336 gnd.n5335 19.3944
R16118 gnd.n5335 gnd.n5334 19.3944
R16119 gnd.n5334 gnd.n5332 19.3944
R16120 gnd.n5332 gnd.n5329 19.3944
R16121 gnd.n5329 gnd.n5328 19.3944
R16122 gnd.n5328 gnd.n5325 19.3944
R16123 gnd.n5325 gnd.n5324 19.3944
R16124 gnd.n5324 gnd.n5321 19.3944
R16125 gnd.n5321 gnd.n5320 19.3944
R16126 gnd.n5320 gnd.n5317 19.3944
R16127 gnd.n5317 gnd.n5316 19.3944
R16128 gnd.n5316 gnd.n5313 19.3944
R16129 gnd.n5313 gnd.n5312 19.3944
R16130 gnd.n5312 gnd.n5309 19.3944
R16131 gnd.n5309 gnd.n5308 19.3944
R16132 gnd.n5308 gnd.n5305 19.3944
R16133 gnd.n5305 gnd.n5304 19.3944
R16134 gnd.n5304 gnd.n5301 19.3944
R16135 gnd.n5301 gnd.n5300 19.3944
R16136 gnd.n5300 gnd.n5297 19.3944
R16137 gnd.n5297 gnd.n5296 19.3944
R16138 gnd.n5293 gnd.n5292 19.3944
R16139 gnd.n5292 gnd.n5248 19.3944
R16140 gnd.n5343 gnd.n5248 19.3944
R16141 gnd.n6157 gnd.n4911 19.3944
R16142 gnd.n6157 gnd.n6156 19.3944
R16143 gnd.n6156 gnd.n6155 19.3944
R16144 gnd.n6199 gnd.n6198 19.3944
R16145 gnd.n6198 gnd.n6197 19.3944
R16146 gnd.n6197 gnd.n4872 19.3944
R16147 gnd.n6192 gnd.n4872 19.3944
R16148 gnd.n6192 gnd.n6191 19.3944
R16149 gnd.n6191 gnd.n6190 19.3944
R16150 gnd.n6190 gnd.n4879 19.3944
R16151 gnd.n6185 gnd.n4879 19.3944
R16152 gnd.n6185 gnd.n6184 19.3944
R16153 gnd.n6184 gnd.n6183 19.3944
R16154 gnd.n6183 gnd.n4886 19.3944
R16155 gnd.n6178 gnd.n4886 19.3944
R16156 gnd.n6178 gnd.n6177 19.3944
R16157 gnd.n6177 gnd.n6176 19.3944
R16158 gnd.n6176 gnd.n4893 19.3944
R16159 gnd.n6171 gnd.n4893 19.3944
R16160 gnd.n6171 gnd.n6170 19.3944
R16161 gnd.n6170 gnd.n6169 19.3944
R16162 gnd.n6169 gnd.n4900 19.3944
R16163 gnd.n6164 gnd.n4900 19.3944
R16164 gnd.n6164 gnd.n6163 19.3944
R16165 gnd.n6163 gnd.n6162 19.3944
R16166 gnd.n5522 gnd.n5145 19.3944
R16167 gnd.n5532 gnd.n5145 19.3944
R16168 gnd.n5533 gnd.n5532 19.3944
R16169 gnd.n5533 gnd.n5126 19.3944
R16170 gnd.n5553 gnd.n5126 19.3944
R16171 gnd.n5553 gnd.n5119 19.3944
R16172 gnd.n5563 gnd.n5119 19.3944
R16173 gnd.n5564 gnd.n5563 19.3944
R16174 gnd.n5564 gnd.n5102 19.3944
R16175 gnd.n5584 gnd.n5102 19.3944
R16176 gnd.n5584 gnd.n5094 19.3944
R16177 gnd.n5594 gnd.n5094 19.3944
R16178 gnd.n5595 gnd.n5594 19.3944
R16179 gnd.n5595 gnd.n5076 19.3944
R16180 gnd.n5615 gnd.n5076 19.3944
R16181 gnd.n5615 gnd.n5068 19.3944
R16182 gnd.n5625 gnd.n5068 19.3944
R16183 gnd.n5626 gnd.n5625 19.3944
R16184 gnd.n5626 gnd.n5051 19.3944
R16185 gnd.n5646 gnd.n5051 19.3944
R16186 gnd.n5646 gnd.n5043 19.3944
R16187 gnd.n5656 gnd.n5043 19.3944
R16188 gnd.n5657 gnd.n5656 19.3944
R16189 gnd.n5657 gnd.n5027 19.3944
R16190 gnd.n5676 gnd.n5027 19.3944
R16191 gnd.n5676 gnd.n5012 19.3944
R16192 gnd.n5710 gnd.n5012 19.3944
R16193 gnd.n5711 gnd.n5710 19.3944
R16194 gnd.n5712 gnd.n5711 19.3944
R16195 gnd.n5712 gnd.n4998 19.3944
R16196 gnd.n4998 gnd.n4992 19.3944
R16197 gnd.n5737 gnd.n4992 19.3944
R16198 gnd.n5738 gnd.n5737 19.3944
R16199 gnd.n5738 gnd.n4975 19.3944
R16200 gnd.n4975 gnd.n4973 19.3944
R16201 gnd.n5764 gnd.n4973 19.3944
R16202 gnd.n5765 gnd.n5764 19.3944
R16203 gnd.n5765 gnd.n4948 19.3944
R16204 gnd.n5811 gnd.n4948 19.3944
R16205 gnd.n5812 gnd.n5811 19.3944
R16206 gnd.n5812 gnd.n4941 19.3944
R16207 gnd.n5823 gnd.n4941 19.3944
R16208 gnd.n5825 gnd.n5823 19.3944
R16209 gnd.n6108 gnd.n5825 19.3944
R16210 gnd.n6108 gnd.n6107 19.3944
R16211 gnd.n6107 gnd.n5828 19.3944
R16212 gnd.n6103 gnd.n5828 19.3944
R16213 gnd.n6103 gnd.n6102 19.3944
R16214 gnd.n6102 gnd.n6101 19.3944
R16215 gnd.n6101 gnd.n6098 19.3944
R16216 gnd.n6098 gnd.n6097 19.3944
R16217 gnd.n6097 gnd.n6094 19.3944
R16218 gnd.n6094 gnd.n6093 19.3944
R16219 gnd.n5513 gnd.n5512 19.3944
R16220 gnd.n5512 gnd.n5159 19.3944
R16221 gnd.n5182 gnd.n5159 19.3944
R16222 gnd.n5185 gnd.n5182 19.3944
R16223 gnd.n5185 gnd.n5178 19.3944
R16224 gnd.n5189 gnd.n5178 19.3944
R16225 gnd.n5192 gnd.n5189 19.3944
R16226 gnd.n5195 gnd.n5192 19.3944
R16227 gnd.n5195 gnd.n5176 19.3944
R16228 gnd.n5199 gnd.n5176 19.3944
R16229 gnd.n5202 gnd.n5199 19.3944
R16230 gnd.n5205 gnd.n5202 19.3944
R16231 gnd.n5205 gnd.n5174 19.3944
R16232 gnd.n5209 gnd.n5174 19.3944
R16233 gnd.n5518 gnd.n5517 19.3944
R16234 gnd.n5517 gnd.n5135 19.3944
R16235 gnd.n5543 gnd.n5135 19.3944
R16236 gnd.n5543 gnd.n5133 19.3944
R16237 gnd.n5549 gnd.n5133 19.3944
R16238 gnd.n5549 gnd.n5548 19.3944
R16239 gnd.n5548 gnd.n5109 19.3944
R16240 gnd.n5574 gnd.n5109 19.3944
R16241 gnd.n5574 gnd.n5107 19.3944
R16242 gnd.n5580 gnd.n5107 19.3944
R16243 gnd.n5580 gnd.n5579 19.3944
R16244 gnd.n5579 gnd.n5084 19.3944
R16245 gnd.n5605 gnd.n5084 19.3944
R16246 gnd.n5605 gnd.n5082 19.3944
R16247 gnd.n5611 gnd.n5082 19.3944
R16248 gnd.n5611 gnd.n5610 19.3944
R16249 gnd.n5610 gnd.n5058 19.3944
R16250 gnd.n5636 gnd.n5058 19.3944
R16251 gnd.n5636 gnd.n5056 19.3944
R16252 gnd.n5642 gnd.n5056 19.3944
R16253 gnd.n5642 gnd.n5641 19.3944
R16254 gnd.n5641 gnd.n5034 19.3944
R16255 gnd.n5666 gnd.n5034 19.3944
R16256 gnd.n5666 gnd.n5032 19.3944
R16257 gnd.n5672 gnd.n5032 19.3944
R16258 gnd.n5672 gnd.n5671 19.3944
R16259 gnd.n5671 gnd.n5003 19.3944
R16260 gnd.n5720 gnd.n5003 19.3944
R16261 gnd.n5720 gnd.n5001 19.3944
R16262 gnd.n5724 gnd.n5001 19.3944
R16263 gnd.n5724 gnd.n4982 19.3944
R16264 gnd.n5750 gnd.n4982 19.3944
R16265 gnd.n5750 gnd.n4980 19.3944
R16266 gnd.n5756 gnd.n4980 19.3944
R16267 gnd.n5756 gnd.n5755 19.3944
R16268 gnd.n5755 gnd.n4958 19.3944
R16269 gnd.n5796 gnd.n4958 19.3944
R16270 gnd.n5796 gnd.n4956 19.3944
R16271 gnd.n5802 gnd.n4956 19.3944
R16272 gnd.n5802 gnd.n5801 19.3944
R16273 gnd.n5801 gnd.n4928 19.3944
R16274 gnd.n6117 gnd.n4928 19.3944
R16275 gnd.n6117 gnd.n4926 19.3944
R16276 gnd.n6127 gnd.n4926 19.3944
R16277 gnd.n6127 gnd.n6126 19.3944
R16278 gnd.n6126 gnd.n6125 19.3944
R16279 gnd.n6125 gnd.n913 19.3944
R16280 gnd.n6248 gnd.n913 19.3944
R16281 gnd.n6248 gnd.n6247 19.3944
R16282 gnd.n6247 gnd.n6246 19.3944
R16283 gnd.n6246 gnd.n917 19.3944
R16284 gnd.n4836 gnd.n917 19.3944
R16285 gnd.n6234 gnd.n4836 19.3944
R16286 gnd.n6231 gnd.n6230 19.3944
R16287 gnd.n6230 gnd.n6229 19.3944
R16288 gnd.n6229 gnd.n4842 19.3944
R16289 gnd.n6224 gnd.n4842 19.3944
R16290 gnd.n6224 gnd.n6223 19.3944
R16291 gnd.n6223 gnd.n6222 19.3944
R16292 gnd.n6222 gnd.n4849 19.3944
R16293 gnd.n6217 gnd.n4849 19.3944
R16294 gnd.n6217 gnd.n6216 19.3944
R16295 gnd.n6216 gnd.n6215 19.3944
R16296 gnd.n6215 gnd.n4856 19.3944
R16297 gnd.n6210 gnd.n4856 19.3944
R16298 gnd.n6210 gnd.n6209 19.3944
R16299 gnd.n6209 gnd.n6208 19.3944
R16300 gnd.n5347 gnd.n5246 19.3944
R16301 gnd.n5347 gnd.n5237 19.3944
R16302 gnd.n5360 gnd.n5237 19.3944
R16303 gnd.n5360 gnd.n5235 19.3944
R16304 gnd.n5364 gnd.n5235 19.3944
R16305 gnd.n5364 gnd.n5225 19.3944
R16306 gnd.n5376 gnd.n5225 19.3944
R16307 gnd.n5376 gnd.n5223 19.3944
R16308 gnd.n5496 gnd.n5223 19.3944
R16309 gnd.n5496 gnd.n5495 19.3944
R16310 gnd.n5495 gnd.n5494 19.3944
R16311 gnd.n5494 gnd.n5493 19.3944
R16312 gnd.n5493 gnd.n5490 19.3944
R16313 gnd.n5490 gnd.n5489 19.3944
R16314 gnd.n5489 gnd.n5488 19.3944
R16315 gnd.n5488 gnd.n5486 19.3944
R16316 gnd.n5486 gnd.n5485 19.3944
R16317 gnd.n5485 gnd.n5482 19.3944
R16318 gnd.n5482 gnd.n5481 19.3944
R16319 gnd.n5481 gnd.n5480 19.3944
R16320 gnd.n5480 gnd.n5478 19.3944
R16321 gnd.n5478 gnd.n5477 19.3944
R16322 gnd.n5477 gnd.n5473 19.3944
R16323 gnd.n5473 gnd.n5472 19.3944
R16324 gnd.n5472 gnd.n5471 19.3944
R16325 gnd.n5471 gnd.n5469 19.3944
R16326 gnd.n5469 gnd.n5468 19.3944
R16327 gnd.n5468 gnd.n5465 19.3944
R16328 gnd.n5465 gnd.n5464 19.3944
R16329 gnd.n5412 gnd.n5400 19.3944
R16330 gnd.n5411 gnd.n5407 19.3944
R16331 gnd.n5405 gnd.n5404 19.3944
R16332 gnd.n5401 gnd.n5020 19.3944
R16333 gnd.n5686 gnd.n5020 19.3944
R16334 gnd.n5686 gnd.n5018 19.3944
R16335 gnd.n5705 gnd.n5018 19.3944
R16336 gnd.n5705 gnd.n5704 19.3944
R16337 gnd.n5704 gnd.n5703 19.3944
R16338 gnd.n5703 gnd.n5701 19.3944
R16339 gnd.n5701 gnd.n5700 19.3944
R16340 gnd.n5700 gnd.n5698 19.3944
R16341 gnd.n5698 gnd.n5697 19.3944
R16342 gnd.n5697 gnd.n4964 19.3944
R16343 gnd.n5773 gnd.n4964 19.3944
R16344 gnd.n5773 gnd.n4962 19.3944
R16345 gnd.n5789 gnd.n4962 19.3944
R16346 gnd.n5789 gnd.n5788 19.3944
R16347 gnd.n5788 gnd.n5787 19.3944
R16348 gnd.n5787 gnd.n5785 19.3944
R16349 gnd.n5785 gnd.n5784 19.3944
R16350 gnd.n5784 gnd.n5782 19.3944
R16351 gnd.n5782 gnd.n4921 19.3944
R16352 gnd.n6132 gnd.n4921 19.3944
R16353 gnd.n6132 gnd.n4919 19.3944
R16354 gnd.n6138 gnd.n4919 19.3944
R16355 gnd.n6139 gnd.n6138 19.3944
R16356 gnd.n6142 gnd.n6139 19.3944
R16357 gnd.n6142 gnd.n4917 19.3944
R16358 gnd.n6146 gnd.n4917 19.3944
R16359 gnd.n6149 gnd.n6146 19.3944
R16360 gnd.n6150 gnd.n6149 19.3944
R16361 gnd.n5352 gnd.n5242 19.3944
R16362 gnd.n5352 gnd.n5240 19.3944
R16363 gnd.n5356 gnd.n5240 19.3944
R16364 gnd.n5356 gnd.n5231 19.3944
R16365 gnd.n5368 gnd.n5231 19.3944
R16366 gnd.n5368 gnd.n5229 19.3944
R16367 gnd.n5372 gnd.n5229 19.3944
R16368 gnd.n5372 gnd.n5218 19.3944
R16369 gnd.n5500 gnd.n5218 19.3944
R16370 gnd.n5500 gnd.n5172 19.3944
R16371 gnd.n5506 gnd.n5172 19.3944
R16372 gnd.n5506 gnd.n5505 19.3944
R16373 gnd.n5505 gnd.n5150 19.3944
R16374 gnd.n5527 gnd.n5150 19.3944
R16375 gnd.n5527 gnd.n5143 19.3944
R16376 gnd.n5538 gnd.n5143 19.3944
R16377 gnd.n5538 gnd.n5537 19.3944
R16378 gnd.n5537 gnd.n5124 19.3944
R16379 gnd.n5558 gnd.n5124 19.3944
R16380 gnd.n5558 gnd.n5117 19.3944
R16381 gnd.n5569 gnd.n5117 19.3944
R16382 gnd.n5569 gnd.n5568 19.3944
R16383 gnd.n5568 gnd.n5100 19.3944
R16384 gnd.n5589 gnd.n5100 19.3944
R16385 gnd.n5589 gnd.n5092 19.3944
R16386 gnd.n5600 gnd.n5092 19.3944
R16387 gnd.n5600 gnd.n5599 19.3944
R16388 gnd.n5599 gnd.n5074 19.3944
R16389 gnd.n5620 gnd.n5074 19.3944
R16390 gnd.n5620 gnd.n5066 19.3944
R16391 gnd.n5631 gnd.n5066 19.3944
R16392 gnd.n5631 gnd.n5630 19.3944
R16393 gnd.n5630 gnd.n5049 19.3944
R16394 gnd.n5651 gnd.n5049 19.3944
R16395 gnd.n5651 gnd.n5041 19.3944
R16396 gnd.n5661 gnd.n5041 19.3944
R16397 gnd.n5661 gnd.n5025 19.3944
R16398 gnd.n5682 gnd.n5025 19.3944
R16399 gnd.n5682 gnd.n5681 19.3944
R16400 gnd.n5681 gnd.n5009 19.3944
R16401 gnd.n5715 gnd.n5009 19.3944
R16402 gnd.n5715 gnd.n4994 19.3944
R16403 gnd.n5732 gnd.n4994 19.3944
R16404 gnd.n5732 gnd.n4990 19.3944
R16405 gnd.n5745 gnd.n4990 19.3944
R16406 gnd.n5745 gnd.n5744 19.3944
R16407 gnd.n5744 gnd.n4969 19.3944
R16408 gnd.n5769 gnd.n4969 19.3944
R16409 gnd.n5769 gnd.n5768 19.3944
R16410 gnd.n5768 gnd.n4950 19.3944
R16411 gnd.n5807 gnd.n4950 19.3944
R16412 gnd.n5807 gnd.n4943 19.3944
R16413 gnd.n5818 gnd.n4943 19.3944
R16414 gnd.n5818 gnd.n4937 19.3944
R16415 gnd.n6112 gnd.n4937 19.3944
R16416 gnd.n6112 gnd.n6111 19.3944
R16417 gnd.n6111 gnd.n901 19.3944
R16418 gnd.n6255 gnd.n901 19.3944
R16419 gnd.n6255 gnd.n6254 19.3944
R16420 gnd.n6254 gnd.n6253 19.3944
R16421 gnd.n6253 gnd.n905 19.3944
R16422 gnd.n925 gnd.n905 19.3944
R16423 gnd.n6241 gnd.n925 19.3944
R16424 gnd.n6241 gnd.n6240 19.3944
R16425 gnd.n6240 gnd.n6239 19.3944
R16426 gnd.n4156 gnd.n1681 19.3944
R16427 gnd.n4161 gnd.n1681 19.3944
R16428 gnd.n4161 gnd.n1682 19.3944
R16429 gnd.n1682 gnd.n1613 19.3944
R16430 gnd.n4187 gnd.n1613 19.3944
R16431 gnd.n4187 gnd.n1610 19.3944
R16432 gnd.n4192 gnd.n1610 19.3944
R16433 gnd.n4192 gnd.n1611 19.3944
R16434 gnd.n1611 gnd.n1586 19.3944
R16435 gnd.n4218 gnd.n1586 19.3944
R16436 gnd.n4218 gnd.n1583 19.3944
R16437 gnd.n4228 gnd.n1583 19.3944
R16438 gnd.n4228 gnd.n1584 19.3944
R16439 gnd.n4224 gnd.n1584 19.3944
R16440 gnd.n4224 gnd.n4223 19.3944
R16441 gnd.n4223 gnd.n1549 19.3944
R16442 gnd.n4285 gnd.n1549 19.3944
R16443 gnd.n4285 gnd.n1550 19.3944
R16444 gnd.n4281 gnd.n1550 19.3944
R16445 gnd.n4281 gnd.n4280 19.3944
R16446 gnd.n4280 gnd.n4279 19.3944
R16447 gnd.n4279 gnd.n311 19.3944
R16448 gnd.n7121 gnd.n311 19.3944
R16449 gnd.n7121 gnd.n309 19.3944
R16450 gnd.n7125 gnd.n309 19.3944
R16451 gnd.n7125 gnd.n69 19.3944
R16452 gnd.n7501 gnd.n69 19.3944
R16453 gnd.n7501 gnd.n7500 19.3944
R16454 gnd.n7500 gnd.n7499 19.3944
R16455 gnd.n7499 gnd.n73 19.3944
R16456 gnd.n7495 gnd.n73 19.3944
R16457 gnd.n7495 gnd.n7494 19.3944
R16458 gnd.n7494 gnd.n7493 19.3944
R16459 gnd.n7493 gnd.n78 19.3944
R16460 gnd.n7489 gnd.n78 19.3944
R16461 gnd.n7489 gnd.n7488 19.3944
R16462 gnd.n7488 gnd.n7487 19.3944
R16463 gnd.n7487 gnd.n83 19.3944
R16464 gnd.n7483 gnd.n83 19.3944
R16465 gnd.n7483 gnd.n7482 19.3944
R16466 gnd.n7482 gnd.n7481 19.3944
R16467 gnd.n7481 gnd.n88 19.3944
R16468 gnd.n7477 gnd.n88 19.3944
R16469 gnd.n7477 gnd.n7476 19.3944
R16470 gnd.n7476 gnd.n7475 19.3944
R16471 gnd.n7475 gnd.n93 19.3944
R16472 gnd.n7471 gnd.n93 19.3944
R16473 gnd.n7471 gnd.n7470 19.3944
R16474 gnd.n7470 gnd.n7469 19.3944
R16475 gnd.n7469 gnd.n98 19.3944
R16476 gnd.n7465 gnd.n98 19.3944
R16477 gnd.n7465 gnd.n7464 19.3944
R16478 gnd.n7464 gnd.n7463 19.3944
R16479 gnd.n7362 gnd.n7361 19.3944
R16480 gnd.n7361 gnd.n7360 19.3944
R16481 gnd.n7360 gnd.n7302 19.3944
R16482 gnd.n7356 gnd.n7302 19.3944
R16483 gnd.n7356 gnd.n7355 19.3944
R16484 gnd.n7355 gnd.n7354 19.3944
R16485 gnd.n7354 gnd.n7310 19.3944
R16486 gnd.n7350 gnd.n7310 19.3944
R16487 gnd.n7350 gnd.n7349 19.3944
R16488 gnd.n7349 gnd.n7348 19.3944
R16489 gnd.n7348 gnd.n7318 19.3944
R16490 gnd.n7344 gnd.n7318 19.3944
R16491 gnd.n7344 gnd.n7343 19.3944
R16492 gnd.n7343 gnd.n7342 19.3944
R16493 gnd.n7342 gnd.n7326 19.3944
R16494 gnd.n7338 gnd.n7326 19.3944
R16495 gnd.n1726 gnd.n1722 19.3944
R16496 gnd.n1729 gnd.n1726 19.3944
R16497 gnd.n1732 gnd.n1729 19.3944
R16498 gnd.n1732 gnd.n1715 19.3944
R16499 gnd.n1745 gnd.n1715 19.3944
R16500 gnd.n1748 gnd.n1745 19.3944
R16501 gnd.n1751 gnd.n1748 19.3944
R16502 gnd.n1751 gnd.n1708 19.3944
R16503 gnd.n1764 gnd.n1708 19.3944
R16504 gnd.n1767 gnd.n1764 19.3944
R16505 gnd.n1770 gnd.n1767 19.3944
R16506 gnd.n1770 gnd.n1701 19.3944
R16507 gnd.n1782 gnd.n1701 19.3944
R16508 gnd.n1785 gnd.n1782 19.3944
R16509 gnd.n1785 gnd.n1693 19.3944
R16510 gnd.n1798 gnd.n1693 19.3944
R16511 gnd.n4347 gnd.n1502 19.3944
R16512 gnd.n4343 gnd.n1502 19.3944
R16513 gnd.n4343 gnd.n4342 19.3944
R16514 gnd.n4342 gnd.n4341 19.3944
R16515 gnd.n4341 gnd.n1508 19.3944
R16516 gnd.n4337 gnd.n1508 19.3944
R16517 gnd.n4337 gnd.n4336 19.3944
R16518 gnd.n4336 gnd.n4335 19.3944
R16519 gnd.n4335 gnd.n1513 19.3944
R16520 gnd.n4331 gnd.n1513 19.3944
R16521 gnd.n4331 gnd.n4330 19.3944
R16522 gnd.n4330 gnd.n4329 19.3944
R16523 gnd.n4329 gnd.n1518 19.3944
R16524 gnd.n4325 gnd.n1518 19.3944
R16525 gnd.n4325 gnd.n4324 19.3944
R16526 gnd.n4324 gnd.n4323 19.3944
R16527 gnd.n4323 gnd.n1523 19.3944
R16528 gnd.n4319 gnd.n1523 19.3944
R16529 gnd.n4319 gnd.n4318 19.3944
R16530 gnd.n4318 gnd.n4317 19.3944
R16531 gnd.n4317 gnd.n283 19.3944
R16532 gnd.n7217 gnd.n283 19.3944
R16533 gnd.n7217 gnd.n284 19.3944
R16534 gnd.n7213 gnd.n284 19.3944
R16535 gnd.n7213 gnd.n7212 19.3944
R16536 gnd.n7212 gnd.n7211 19.3944
R16537 gnd.n7211 gnd.n290 19.3944
R16538 gnd.n7206 gnd.n290 19.3944
R16539 gnd.n7206 gnd.n7205 19.3944
R16540 gnd.n7205 gnd.n261 19.3944
R16541 gnd.n7228 gnd.n261 19.3944
R16542 gnd.n7228 gnd.n259 19.3944
R16543 gnd.n7232 gnd.n259 19.3944
R16544 gnd.n7232 gnd.n245 19.3944
R16545 gnd.n7244 gnd.n245 19.3944
R16546 gnd.n7244 gnd.n243 19.3944
R16547 gnd.n7248 gnd.n243 19.3944
R16548 gnd.n7248 gnd.n230 19.3944
R16549 gnd.n7260 gnd.n230 19.3944
R16550 gnd.n7260 gnd.n228 19.3944
R16551 gnd.n7264 gnd.n228 19.3944
R16552 gnd.n7264 gnd.n215 19.3944
R16553 gnd.n7276 gnd.n215 19.3944
R16554 gnd.n7276 gnd.n213 19.3944
R16555 gnd.n7280 gnd.n213 19.3944
R16556 gnd.n7280 gnd.n200 19.3944
R16557 gnd.n7292 gnd.n200 19.3944
R16558 gnd.n7292 gnd.n197 19.3944
R16559 gnd.n7371 gnd.n197 19.3944
R16560 gnd.n7371 gnd.n198 19.3944
R16561 gnd.n7367 gnd.n198 19.3944
R16562 gnd.n7367 gnd.n7366 19.3944
R16563 gnd.n7366 gnd.n7365 19.3944
R16564 gnd.n2235 gnd.n1276 19.3944
R16565 gnd.n2235 gnd.n2185 19.3944
R16566 gnd.n3713 gnd.n2185 19.3944
R16567 gnd.n3713 gnd.n3712 19.3944
R16568 gnd.n3712 gnd.n2188 19.3944
R16569 gnd.n3705 gnd.n2188 19.3944
R16570 gnd.n3705 gnd.n3704 19.3944
R16571 gnd.n3704 gnd.n2197 19.3944
R16572 gnd.n3697 gnd.n2197 19.3944
R16573 gnd.n3697 gnd.n3696 19.3944
R16574 gnd.n3696 gnd.n2205 19.3944
R16575 gnd.n3689 gnd.n2205 19.3944
R16576 gnd.n3689 gnd.n3688 19.3944
R16577 gnd.n3688 gnd.n2215 19.3944
R16578 gnd.n3681 gnd.n2215 19.3944
R16579 gnd.n3681 gnd.n3680 19.3944
R16580 gnd.n6884 gnd.n452 19.3944
R16581 gnd.n6890 gnd.n452 19.3944
R16582 gnd.n6890 gnd.n450 19.3944
R16583 gnd.n6894 gnd.n450 19.3944
R16584 gnd.n6894 gnd.n446 19.3944
R16585 gnd.n6900 gnd.n446 19.3944
R16586 gnd.n6900 gnd.n444 19.3944
R16587 gnd.n6904 gnd.n444 19.3944
R16588 gnd.n6904 gnd.n440 19.3944
R16589 gnd.n6910 gnd.n440 19.3944
R16590 gnd.n6910 gnd.n438 19.3944
R16591 gnd.n6914 gnd.n438 19.3944
R16592 gnd.n6914 gnd.n434 19.3944
R16593 gnd.n6920 gnd.n434 19.3944
R16594 gnd.n6920 gnd.n432 19.3944
R16595 gnd.n6924 gnd.n432 19.3944
R16596 gnd.n6924 gnd.n428 19.3944
R16597 gnd.n6930 gnd.n428 19.3944
R16598 gnd.n6930 gnd.n426 19.3944
R16599 gnd.n6934 gnd.n426 19.3944
R16600 gnd.n6934 gnd.n422 19.3944
R16601 gnd.n6940 gnd.n422 19.3944
R16602 gnd.n6940 gnd.n420 19.3944
R16603 gnd.n6944 gnd.n420 19.3944
R16604 gnd.n6944 gnd.n416 19.3944
R16605 gnd.n6950 gnd.n416 19.3944
R16606 gnd.n6950 gnd.n414 19.3944
R16607 gnd.n6954 gnd.n414 19.3944
R16608 gnd.n6954 gnd.n410 19.3944
R16609 gnd.n6960 gnd.n410 19.3944
R16610 gnd.n6960 gnd.n408 19.3944
R16611 gnd.n6964 gnd.n408 19.3944
R16612 gnd.n6964 gnd.n404 19.3944
R16613 gnd.n6970 gnd.n404 19.3944
R16614 gnd.n6970 gnd.n402 19.3944
R16615 gnd.n6974 gnd.n402 19.3944
R16616 gnd.n6974 gnd.n398 19.3944
R16617 gnd.n6980 gnd.n398 19.3944
R16618 gnd.n6980 gnd.n396 19.3944
R16619 gnd.n6984 gnd.n396 19.3944
R16620 gnd.n6984 gnd.n392 19.3944
R16621 gnd.n6990 gnd.n392 19.3944
R16622 gnd.n6990 gnd.n390 19.3944
R16623 gnd.n6994 gnd.n390 19.3944
R16624 gnd.n6994 gnd.n386 19.3944
R16625 gnd.n7000 gnd.n386 19.3944
R16626 gnd.n7000 gnd.n384 19.3944
R16627 gnd.n7004 gnd.n384 19.3944
R16628 gnd.n7004 gnd.n380 19.3944
R16629 gnd.n7010 gnd.n380 19.3944
R16630 gnd.n7010 gnd.n378 19.3944
R16631 gnd.n7014 gnd.n378 19.3944
R16632 gnd.n7014 gnd.n374 19.3944
R16633 gnd.n7020 gnd.n374 19.3944
R16634 gnd.n7020 gnd.n372 19.3944
R16635 gnd.n7024 gnd.n372 19.3944
R16636 gnd.n7024 gnd.n368 19.3944
R16637 gnd.n7030 gnd.n368 19.3944
R16638 gnd.n7030 gnd.n366 19.3944
R16639 gnd.n7034 gnd.n366 19.3944
R16640 gnd.n7034 gnd.n362 19.3944
R16641 gnd.n7040 gnd.n362 19.3944
R16642 gnd.n7040 gnd.n360 19.3944
R16643 gnd.n7044 gnd.n360 19.3944
R16644 gnd.n7044 gnd.n356 19.3944
R16645 gnd.n7050 gnd.n356 19.3944
R16646 gnd.n7050 gnd.n354 19.3944
R16647 gnd.n7054 gnd.n354 19.3944
R16648 gnd.n7054 gnd.n350 19.3944
R16649 gnd.n7060 gnd.n350 19.3944
R16650 gnd.n7060 gnd.n348 19.3944
R16651 gnd.n7064 gnd.n348 19.3944
R16652 gnd.n7064 gnd.n344 19.3944
R16653 gnd.n7070 gnd.n344 19.3944
R16654 gnd.n7070 gnd.n342 19.3944
R16655 gnd.n7074 gnd.n342 19.3944
R16656 gnd.n7074 gnd.n338 19.3944
R16657 gnd.n7080 gnd.n338 19.3944
R16658 gnd.n7080 gnd.n336 19.3944
R16659 gnd.n7084 gnd.n336 19.3944
R16660 gnd.n7084 gnd.n332 19.3944
R16661 gnd.n7091 gnd.n332 19.3944
R16662 gnd.n7091 gnd.n330 19.3944
R16663 gnd.n7096 gnd.n330 19.3944
R16664 gnd.n6429 gnd.n725 19.3944
R16665 gnd.n6433 gnd.n725 19.3944
R16666 gnd.n6433 gnd.n721 19.3944
R16667 gnd.n6439 gnd.n721 19.3944
R16668 gnd.n6439 gnd.n719 19.3944
R16669 gnd.n6443 gnd.n719 19.3944
R16670 gnd.n6443 gnd.n715 19.3944
R16671 gnd.n6449 gnd.n715 19.3944
R16672 gnd.n6449 gnd.n713 19.3944
R16673 gnd.n6453 gnd.n713 19.3944
R16674 gnd.n6453 gnd.n709 19.3944
R16675 gnd.n6459 gnd.n709 19.3944
R16676 gnd.n6459 gnd.n707 19.3944
R16677 gnd.n6463 gnd.n707 19.3944
R16678 gnd.n6463 gnd.n703 19.3944
R16679 gnd.n6469 gnd.n703 19.3944
R16680 gnd.n6469 gnd.n701 19.3944
R16681 gnd.n6473 gnd.n701 19.3944
R16682 gnd.n6473 gnd.n697 19.3944
R16683 gnd.n6479 gnd.n697 19.3944
R16684 gnd.n6479 gnd.n695 19.3944
R16685 gnd.n6483 gnd.n695 19.3944
R16686 gnd.n6483 gnd.n691 19.3944
R16687 gnd.n6489 gnd.n691 19.3944
R16688 gnd.n6489 gnd.n689 19.3944
R16689 gnd.n6493 gnd.n689 19.3944
R16690 gnd.n6493 gnd.n685 19.3944
R16691 gnd.n6499 gnd.n685 19.3944
R16692 gnd.n6499 gnd.n683 19.3944
R16693 gnd.n6503 gnd.n683 19.3944
R16694 gnd.n6503 gnd.n679 19.3944
R16695 gnd.n6509 gnd.n679 19.3944
R16696 gnd.n6509 gnd.n677 19.3944
R16697 gnd.n6513 gnd.n677 19.3944
R16698 gnd.n6513 gnd.n673 19.3944
R16699 gnd.n6519 gnd.n673 19.3944
R16700 gnd.n6519 gnd.n671 19.3944
R16701 gnd.n6523 gnd.n671 19.3944
R16702 gnd.n6523 gnd.n667 19.3944
R16703 gnd.n6529 gnd.n667 19.3944
R16704 gnd.n6529 gnd.n665 19.3944
R16705 gnd.n6533 gnd.n665 19.3944
R16706 gnd.n6533 gnd.n661 19.3944
R16707 gnd.n6539 gnd.n661 19.3944
R16708 gnd.n6539 gnd.n659 19.3944
R16709 gnd.n6543 gnd.n659 19.3944
R16710 gnd.n6543 gnd.n655 19.3944
R16711 gnd.n6549 gnd.n655 19.3944
R16712 gnd.n6549 gnd.n653 19.3944
R16713 gnd.n6553 gnd.n653 19.3944
R16714 gnd.n6553 gnd.n649 19.3944
R16715 gnd.n6559 gnd.n649 19.3944
R16716 gnd.n6559 gnd.n647 19.3944
R16717 gnd.n6563 gnd.n647 19.3944
R16718 gnd.n6563 gnd.n643 19.3944
R16719 gnd.n6569 gnd.n643 19.3944
R16720 gnd.n6569 gnd.n641 19.3944
R16721 gnd.n6573 gnd.n641 19.3944
R16722 gnd.n6573 gnd.n637 19.3944
R16723 gnd.n6579 gnd.n637 19.3944
R16724 gnd.n6579 gnd.n635 19.3944
R16725 gnd.n6583 gnd.n635 19.3944
R16726 gnd.n6583 gnd.n631 19.3944
R16727 gnd.n6589 gnd.n631 19.3944
R16728 gnd.n6589 gnd.n629 19.3944
R16729 gnd.n6593 gnd.n629 19.3944
R16730 gnd.n6593 gnd.n625 19.3944
R16731 gnd.n6599 gnd.n625 19.3944
R16732 gnd.n6599 gnd.n623 19.3944
R16733 gnd.n6603 gnd.n623 19.3944
R16734 gnd.n6603 gnd.n619 19.3944
R16735 gnd.n6609 gnd.n619 19.3944
R16736 gnd.n6609 gnd.n617 19.3944
R16737 gnd.n6613 gnd.n617 19.3944
R16738 gnd.n6613 gnd.n613 19.3944
R16739 gnd.n6619 gnd.n613 19.3944
R16740 gnd.n6619 gnd.n611 19.3944
R16741 gnd.n6623 gnd.n611 19.3944
R16742 gnd.n6623 gnd.n607 19.3944
R16743 gnd.n6629 gnd.n607 19.3944
R16744 gnd.n6629 gnd.n605 19.3944
R16745 gnd.n6633 gnd.n605 19.3944
R16746 gnd.n6633 gnd.n601 19.3944
R16747 gnd.n6639 gnd.n601 19.3944
R16748 gnd.n6639 gnd.n599 19.3944
R16749 gnd.n6643 gnd.n599 19.3944
R16750 gnd.n6643 gnd.n595 19.3944
R16751 gnd.n6649 gnd.n595 19.3944
R16752 gnd.n6649 gnd.n593 19.3944
R16753 gnd.n6653 gnd.n593 19.3944
R16754 gnd.n6653 gnd.n589 19.3944
R16755 gnd.n6659 gnd.n589 19.3944
R16756 gnd.n6659 gnd.n587 19.3944
R16757 gnd.n6663 gnd.n587 19.3944
R16758 gnd.n6663 gnd.n583 19.3944
R16759 gnd.n6669 gnd.n583 19.3944
R16760 gnd.n6669 gnd.n581 19.3944
R16761 gnd.n6673 gnd.n581 19.3944
R16762 gnd.n6673 gnd.n577 19.3944
R16763 gnd.n6679 gnd.n577 19.3944
R16764 gnd.n6679 gnd.n575 19.3944
R16765 gnd.n6683 gnd.n575 19.3944
R16766 gnd.n6683 gnd.n571 19.3944
R16767 gnd.n6689 gnd.n571 19.3944
R16768 gnd.n6689 gnd.n569 19.3944
R16769 gnd.n6693 gnd.n569 19.3944
R16770 gnd.n6693 gnd.n565 19.3944
R16771 gnd.n6699 gnd.n565 19.3944
R16772 gnd.n6699 gnd.n563 19.3944
R16773 gnd.n6703 gnd.n563 19.3944
R16774 gnd.n6703 gnd.n559 19.3944
R16775 gnd.n6709 gnd.n559 19.3944
R16776 gnd.n6709 gnd.n557 19.3944
R16777 gnd.n6713 gnd.n557 19.3944
R16778 gnd.n6713 gnd.n553 19.3944
R16779 gnd.n6719 gnd.n553 19.3944
R16780 gnd.n6719 gnd.n551 19.3944
R16781 gnd.n6723 gnd.n551 19.3944
R16782 gnd.n6723 gnd.n547 19.3944
R16783 gnd.n6729 gnd.n547 19.3944
R16784 gnd.n6729 gnd.n545 19.3944
R16785 gnd.n6733 gnd.n545 19.3944
R16786 gnd.n6733 gnd.n541 19.3944
R16787 gnd.n6739 gnd.n541 19.3944
R16788 gnd.n6739 gnd.n539 19.3944
R16789 gnd.n6743 gnd.n539 19.3944
R16790 gnd.n6743 gnd.n535 19.3944
R16791 gnd.n6749 gnd.n535 19.3944
R16792 gnd.n6749 gnd.n533 19.3944
R16793 gnd.n6753 gnd.n533 19.3944
R16794 gnd.n6753 gnd.n529 19.3944
R16795 gnd.n6759 gnd.n529 19.3944
R16796 gnd.n6759 gnd.n527 19.3944
R16797 gnd.n6763 gnd.n527 19.3944
R16798 gnd.n6763 gnd.n523 19.3944
R16799 gnd.n6769 gnd.n523 19.3944
R16800 gnd.n6769 gnd.n521 19.3944
R16801 gnd.n6773 gnd.n521 19.3944
R16802 gnd.n6773 gnd.n517 19.3944
R16803 gnd.n6779 gnd.n517 19.3944
R16804 gnd.n6779 gnd.n515 19.3944
R16805 gnd.n6783 gnd.n515 19.3944
R16806 gnd.n6783 gnd.n511 19.3944
R16807 gnd.n6789 gnd.n511 19.3944
R16808 gnd.n6789 gnd.n509 19.3944
R16809 gnd.n6793 gnd.n509 19.3944
R16810 gnd.n6793 gnd.n505 19.3944
R16811 gnd.n6799 gnd.n505 19.3944
R16812 gnd.n6799 gnd.n503 19.3944
R16813 gnd.n6803 gnd.n503 19.3944
R16814 gnd.n6803 gnd.n499 19.3944
R16815 gnd.n6809 gnd.n499 19.3944
R16816 gnd.n6809 gnd.n497 19.3944
R16817 gnd.n6813 gnd.n497 19.3944
R16818 gnd.n6813 gnd.n493 19.3944
R16819 gnd.n6819 gnd.n493 19.3944
R16820 gnd.n6819 gnd.n491 19.3944
R16821 gnd.n6823 gnd.n491 19.3944
R16822 gnd.n6823 gnd.n487 19.3944
R16823 gnd.n6829 gnd.n487 19.3944
R16824 gnd.n6829 gnd.n485 19.3944
R16825 gnd.n6833 gnd.n485 19.3944
R16826 gnd.n6833 gnd.n481 19.3944
R16827 gnd.n6839 gnd.n481 19.3944
R16828 gnd.n6839 gnd.n479 19.3944
R16829 gnd.n6843 gnd.n479 19.3944
R16830 gnd.n6843 gnd.n475 19.3944
R16831 gnd.n6849 gnd.n475 19.3944
R16832 gnd.n6849 gnd.n473 19.3944
R16833 gnd.n6853 gnd.n473 19.3944
R16834 gnd.n6853 gnd.n469 19.3944
R16835 gnd.n6859 gnd.n469 19.3944
R16836 gnd.n6859 gnd.n467 19.3944
R16837 gnd.n6863 gnd.n467 19.3944
R16838 gnd.n6863 gnd.n463 19.3944
R16839 gnd.n6869 gnd.n463 19.3944
R16840 gnd.n6869 gnd.n461 19.3944
R16841 gnd.n6874 gnd.n461 19.3944
R16842 gnd.n6874 gnd.n457 19.3944
R16843 gnd.n6880 gnd.n457 19.3944
R16844 gnd.n6881 gnd.n6880 19.3944
R16845 gnd.n4422 gnd.n4421 19.3944
R16846 gnd.n4421 gnd.n4420 19.3944
R16847 gnd.n4420 gnd.n4419 19.3944
R16848 gnd.n4419 gnd.n4417 19.3944
R16849 gnd.n4417 gnd.n4414 19.3944
R16850 gnd.n4414 gnd.n4413 19.3944
R16851 gnd.n4413 gnd.n4410 19.3944
R16852 gnd.n4410 gnd.n4409 19.3944
R16853 gnd.n4409 gnd.n4406 19.3944
R16854 gnd.n4406 gnd.n4405 19.3944
R16855 gnd.n4405 gnd.n4402 19.3944
R16856 gnd.n4402 gnd.n4401 19.3944
R16857 gnd.n4401 gnd.n4398 19.3944
R16858 gnd.n4398 gnd.n4397 19.3944
R16859 gnd.n4397 gnd.n4394 19.3944
R16860 gnd.n4392 gnd.n4389 19.3944
R16861 gnd.n4389 gnd.n4388 19.3944
R16862 gnd.n4388 gnd.n4385 19.3944
R16863 gnd.n4385 gnd.n4384 19.3944
R16864 gnd.n4384 gnd.n4381 19.3944
R16865 gnd.n4381 gnd.n4380 19.3944
R16866 gnd.n4380 gnd.n4377 19.3944
R16867 gnd.n4377 gnd.n4376 19.3944
R16868 gnd.n4376 gnd.n4373 19.3944
R16869 gnd.n4373 gnd.n4372 19.3944
R16870 gnd.n4372 gnd.n4369 19.3944
R16871 gnd.n4369 gnd.n4368 19.3944
R16872 gnd.n4368 gnd.n4365 19.3944
R16873 gnd.n4365 gnd.n4364 19.3944
R16874 gnd.n4364 gnd.n4361 19.3944
R16875 gnd.n4361 gnd.n4360 19.3944
R16876 gnd.n4360 gnd.n4357 19.3944
R16877 gnd.n4357 gnd.n4356 19.3944
R16878 gnd.n1648 gnd.n1496 19.3944
R16879 gnd.n1678 gnd.n1648 19.3944
R16880 gnd.n1678 gnd.n1677 19.3944
R16881 gnd.n1677 gnd.n1676 19.3944
R16882 gnd.n1676 gnd.n1674 19.3944
R16883 gnd.n1674 gnd.n1673 19.3944
R16884 gnd.n1673 gnd.n1670 19.3944
R16885 gnd.n1670 gnd.n1669 19.3944
R16886 gnd.n1669 gnd.n1668 19.3944
R16887 gnd.n1668 gnd.n1666 19.3944
R16888 gnd.n1666 gnd.n1665 19.3944
R16889 gnd.n1665 gnd.n1663 19.3944
R16890 gnd.n1663 gnd.n1662 19.3944
R16891 gnd.n1662 gnd.n1558 19.3944
R16892 gnd.n4255 gnd.n1558 19.3944
R16893 gnd.n4255 gnd.n1556 19.3944
R16894 gnd.n4259 gnd.n1556 19.3944
R16895 gnd.n4260 gnd.n4259 19.3944
R16896 gnd.n4262 gnd.n4260 19.3944
R16897 gnd.n4262 gnd.n1554 19.3944
R16898 gnd.n4274 gnd.n1554 19.3944
R16899 gnd.n4274 gnd.n4273 19.3944
R16900 gnd.n4273 gnd.n4272 19.3944
R16901 gnd.n4272 gnd.n4271 19.3944
R16902 gnd.n4271 gnd.n299 19.3944
R16903 gnd.n7134 gnd.n299 19.3944
R16904 gnd.n7135 gnd.n7134 19.3944
R16905 gnd.n7196 gnd.n7135 19.3944
R16906 gnd.n7196 gnd.n7195 19.3944
R16907 gnd.n7195 gnd.n7194 19.3944
R16908 gnd.n7194 gnd.n7190 19.3944
R16909 gnd.n7190 gnd.n7189 19.3944
R16910 gnd.n7189 gnd.n7186 19.3944
R16911 gnd.n7186 gnd.n7185 19.3944
R16912 gnd.n7185 gnd.n7183 19.3944
R16913 gnd.n7183 gnd.n7182 19.3944
R16914 gnd.n7182 gnd.n7180 19.3944
R16915 gnd.n7180 gnd.n7179 19.3944
R16916 gnd.n7179 gnd.n7177 19.3944
R16917 gnd.n7177 gnd.n7176 19.3944
R16918 gnd.n7176 gnd.n7174 19.3944
R16919 gnd.n7174 gnd.n7173 19.3944
R16920 gnd.n7173 gnd.n7171 19.3944
R16921 gnd.n7171 gnd.n7170 19.3944
R16922 gnd.n7170 gnd.n7168 19.3944
R16923 gnd.n7168 gnd.n7167 19.3944
R16924 gnd.n7167 gnd.n7165 19.3944
R16925 gnd.n7165 gnd.n7164 19.3944
R16926 gnd.n7164 gnd.n7162 19.3944
R16927 gnd.n7162 gnd.n7161 19.3944
R16928 gnd.n7161 gnd.n182 19.3944
R16929 gnd.n7384 gnd.n182 19.3944
R16930 gnd.n7385 gnd.n7384 19.3944
R16931 gnd.n7423 gnd.n143 19.3944
R16932 gnd.n7418 gnd.n143 19.3944
R16933 gnd.n7418 gnd.n7417 19.3944
R16934 gnd.n7417 gnd.n7416 19.3944
R16935 gnd.n7416 gnd.n150 19.3944
R16936 gnd.n7411 gnd.n150 19.3944
R16937 gnd.n7411 gnd.n7410 19.3944
R16938 gnd.n7410 gnd.n7409 19.3944
R16939 gnd.n7409 gnd.n157 19.3944
R16940 gnd.n7404 gnd.n157 19.3944
R16941 gnd.n7404 gnd.n7403 19.3944
R16942 gnd.n7403 gnd.n7402 19.3944
R16943 gnd.n7402 gnd.n164 19.3944
R16944 gnd.n7397 gnd.n164 19.3944
R16945 gnd.n7397 gnd.n7396 19.3944
R16946 gnd.n7396 gnd.n7395 19.3944
R16947 gnd.n7395 gnd.n171 19.3944
R16948 gnd.n7390 gnd.n171 19.3944
R16949 gnd.n7456 gnd.n7455 19.3944
R16950 gnd.n7455 gnd.n7454 19.3944
R16951 gnd.n7454 gnd.n115 19.3944
R16952 gnd.n7449 gnd.n115 19.3944
R16953 gnd.n7449 gnd.n7448 19.3944
R16954 gnd.n7448 gnd.n7447 19.3944
R16955 gnd.n7447 gnd.n122 19.3944
R16956 gnd.n7442 gnd.n122 19.3944
R16957 gnd.n7442 gnd.n7441 19.3944
R16958 gnd.n7441 gnd.n7440 19.3944
R16959 gnd.n7440 gnd.n129 19.3944
R16960 gnd.n7435 gnd.n129 19.3944
R16961 gnd.n7435 gnd.n7434 19.3944
R16962 gnd.n7434 gnd.n7433 19.3944
R16963 gnd.n7433 gnd.n136 19.3944
R16964 gnd.n7428 gnd.n136 19.3944
R16965 gnd.n7428 gnd.n7427 19.3944
R16966 gnd.n1645 gnd.n1642 19.3944
R16967 gnd.n1645 gnd.n1623 19.3944
R16968 gnd.n4177 gnd.n1623 19.3944
R16969 gnd.n4177 gnd.n1621 19.3944
R16970 gnd.n4183 gnd.n1621 19.3944
R16971 gnd.n4183 gnd.n4182 19.3944
R16972 gnd.n4182 gnd.n1595 19.3944
R16973 gnd.n4208 gnd.n1595 19.3944
R16974 gnd.n4208 gnd.n1593 19.3944
R16975 gnd.n4214 gnd.n1593 19.3944
R16976 gnd.n4214 gnd.n4213 19.3944
R16977 gnd.n4213 gnd.n1568 19.3944
R16978 gnd.n4245 gnd.n1568 19.3944
R16979 gnd.n4245 gnd.n1566 19.3944
R16980 gnd.n4251 gnd.n1566 19.3944
R16981 gnd.n4251 gnd.n4250 19.3944
R16982 gnd.n4250 gnd.n1533 19.3944
R16983 gnd.n4308 gnd.n1533 19.3944
R16984 gnd.n4308 gnd.n1531 19.3944
R16985 gnd.n4312 gnd.n1531 19.3944
R16986 gnd.n4312 gnd.n275 19.3944
R16987 gnd.n7221 gnd.n275 19.3944
R16988 gnd.n274 gnd.n273 19.3944
R16989 gnd.n306 gnd.n273 19.3944
R16990 gnd.n7130 gnd.n7129 19.3944
R16991 gnd.n7201 gnd.n7200 19.3944
R16992 gnd.n7224 gnd.n267 19.3944
R16993 gnd.n7224 gnd.n254 19.3944
R16994 gnd.n7236 gnd.n254 19.3944
R16995 gnd.n7236 gnd.n252 19.3944
R16996 gnd.n7240 gnd.n252 19.3944
R16997 gnd.n7240 gnd.n236 19.3944
R16998 gnd.n7252 gnd.n236 19.3944
R16999 gnd.n7252 gnd.n234 19.3944
R17000 gnd.n7256 gnd.n234 19.3944
R17001 gnd.n7256 gnd.n223 19.3944
R17002 gnd.n7268 gnd.n223 19.3944
R17003 gnd.n7268 gnd.n221 19.3944
R17004 gnd.n7272 gnd.n221 19.3944
R17005 gnd.n7272 gnd.n206 19.3944
R17006 gnd.n7284 gnd.n206 19.3944
R17007 gnd.n7284 gnd.n204 19.3944
R17008 gnd.n7288 gnd.n204 19.3944
R17009 gnd.n7288 gnd.n191 19.3944
R17010 gnd.n7375 gnd.n191 19.3944
R17011 gnd.n7375 gnd.n189 19.3944
R17012 gnd.n7379 gnd.n189 19.3944
R17013 gnd.n7379 gnd.n110 19.3944
R17014 gnd.n7459 gnd.n110 19.3944
R17015 gnd.n2395 gnd.n2391 19.3944
R17016 gnd.n2637 gnd.n2391 19.3944
R17017 gnd.n2637 gnd.n2392 19.3944
R17018 gnd.n2589 gnd.n2588 19.3944
R17019 gnd.n2597 gnd.n2596 19.3944
R17020 gnd.n2593 gnd.n2592 19.3944
R17021 gnd.n2641 gnd.n2366 19.3944
R17022 gnd.n2384 gnd.n2367 19.3944
R17023 gnd.n2384 gnd.n2369 19.3944
R17024 gnd.n2380 gnd.n2369 19.3944
R17025 gnd.n2380 gnd.n2379 19.3944
R17026 gnd.n2379 gnd.n2378 19.3944
R17027 gnd.n2378 gnd.n2376 19.3944
R17028 gnd.n2376 gnd.n2338 19.3944
R17029 gnd.n2338 gnd.n2336 19.3944
R17030 gnd.n2713 gnd.n2336 19.3944
R17031 gnd.n2713 gnd.n2334 19.3944
R17032 gnd.n2717 gnd.n2334 19.3944
R17033 gnd.n2717 gnd.n2332 19.3944
R17034 gnd.n2721 gnd.n2332 19.3944
R17035 gnd.n2721 gnd.n2330 19.3944
R17036 gnd.n2761 gnd.n2330 19.3944
R17037 gnd.n2761 gnd.n2760 19.3944
R17038 gnd.n2760 gnd.n2759 19.3944
R17039 gnd.n2759 gnd.n2727 19.3944
R17040 gnd.n2755 gnd.n2727 19.3944
R17041 gnd.n2755 gnd.n2754 19.3944
R17042 gnd.n2754 gnd.n2753 19.3944
R17043 gnd.n2753 gnd.n2733 19.3944
R17044 gnd.n2749 gnd.n2733 19.3944
R17045 gnd.n2749 gnd.n2748 19.3944
R17046 gnd.n2748 gnd.n2747 19.3944
R17047 gnd.n2747 gnd.n2739 19.3944
R17048 gnd.n2742 gnd.n2739 19.3944
R17049 gnd.n2742 gnd.n2157 19.3944
R17050 gnd.n3731 gnd.n2157 19.3944
R17051 gnd.n3731 gnd.n2155 19.3944
R17052 gnd.n3735 gnd.n2155 19.3944
R17053 gnd.n3735 gnd.n2143 19.3944
R17054 gnd.n3747 gnd.n2143 19.3944
R17055 gnd.n3747 gnd.n2141 19.3944
R17056 gnd.n3751 gnd.n2141 19.3944
R17057 gnd.n3751 gnd.n2131 19.3944
R17058 gnd.n3763 gnd.n2131 19.3944
R17059 gnd.n3763 gnd.n2129 19.3944
R17060 gnd.n3767 gnd.n2129 19.3944
R17061 gnd.n3767 gnd.n2118 19.3944
R17062 gnd.n3779 gnd.n2118 19.3944
R17063 gnd.n3779 gnd.n2116 19.3944
R17064 gnd.n3783 gnd.n2116 19.3944
R17065 gnd.n3783 gnd.n2105 19.3944
R17066 gnd.n3795 gnd.n2105 19.3944
R17067 gnd.n3795 gnd.n2103 19.3944
R17068 gnd.n3799 gnd.n2103 19.3944
R17069 gnd.n3799 gnd.n2091 19.3944
R17070 gnd.n3811 gnd.n2091 19.3944
R17071 gnd.n3811 gnd.n2089 19.3944
R17072 gnd.n3815 gnd.n2089 19.3944
R17073 gnd.n3815 gnd.n2079 19.3944
R17074 gnd.n3827 gnd.n2079 19.3944
R17075 gnd.n3827 gnd.n2077 19.3944
R17076 gnd.n3831 gnd.n2077 19.3944
R17077 gnd.n3831 gnd.n2064 19.3944
R17078 gnd.n3843 gnd.n2064 19.3944
R17079 gnd.n3843 gnd.n2062 19.3944
R17080 gnd.n3847 gnd.n2062 19.3944
R17081 gnd.n3847 gnd.n2049 19.3944
R17082 gnd.n3859 gnd.n2049 19.3944
R17083 gnd.n3859 gnd.n2047 19.3944
R17084 gnd.n3863 gnd.n2047 19.3944
R17085 gnd.n3863 gnd.n2036 19.3944
R17086 gnd.n3875 gnd.n2036 19.3944
R17087 gnd.n3875 gnd.n2034 19.3944
R17088 gnd.n3879 gnd.n2034 19.3944
R17089 gnd.n3879 gnd.n2021 19.3944
R17090 gnd.n3891 gnd.n2021 19.3944
R17091 gnd.n3891 gnd.n2019 19.3944
R17092 gnd.n3895 gnd.n2019 19.3944
R17093 gnd.n3895 gnd.n2006 19.3944
R17094 gnd.n3907 gnd.n2006 19.3944
R17095 gnd.n3907 gnd.n2004 19.3944
R17096 gnd.n3911 gnd.n2004 19.3944
R17097 gnd.n3911 gnd.n1993 19.3944
R17098 gnd.n3923 gnd.n1993 19.3944
R17099 gnd.n3923 gnd.n1991 19.3944
R17100 gnd.n3927 gnd.n1991 19.3944
R17101 gnd.n3927 gnd.n1979 19.3944
R17102 gnd.n3939 gnd.n1979 19.3944
R17103 gnd.n3939 gnd.n1977 19.3944
R17104 gnd.n3943 gnd.n1977 19.3944
R17105 gnd.n3943 gnd.n1964 19.3944
R17106 gnd.n3955 gnd.n1964 19.3944
R17107 gnd.n3955 gnd.n1962 19.3944
R17108 gnd.n3959 gnd.n1962 19.3944
R17109 gnd.n3959 gnd.n1951 19.3944
R17110 gnd.n3971 gnd.n1951 19.3944
R17111 gnd.n3971 gnd.n1949 19.3944
R17112 gnd.n3975 gnd.n1949 19.3944
R17113 gnd.n3975 gnd.n1936 19.3944
R17114 gnd.n3987 gnd.n1936 19.3944
R17115 gnd.n3987 gnd.n1934 19.3944
R17116 gnd.n3991 gnd.n1934 19.3944
R17117 gnd.n3991 gnd.n1923 19.3944
R17118 gnd.n4003 gnd.n1923 19.3944
R17119 gnd.n4003 gnd.n1921 19.3944
R17120 gnd.n4007 gnd.n1921 19.3944
R17121 gnd.n4007 gnd.n1909 19.3944
R17122 gnd.n4019 gnd.n1909 19.3944
R17123 gnd.n4019 gnd.n1907 19.3944
R17124 gnd.n4023 gnd.n1907 19.3944
R17125 gnd.n4023 gnd.n1894 19.3944
R17126 gnd.n4035 gnd.n1894 19.3944
R17127 gnd.n4035 gnd.n1892 19.3944
R17128 gnd.n4039 gnd.n1892 19.3944
R17129 gnd.n4039 gnd.n1882 19.3944
R17130 gnd.n4051 gnd.n1882 19.3944
R17131 gnd.n4051 gnd.n1880 19.3944
R17132 gnd.n4055 gnd.n1880 19.3944
R17133 gnd.n4055 gnd.n1869 19.3944
R17134 gnd.n4067 gnd.n1869 19.3944
R17135 gnd.n4067 gnd.n1867 19.3944
R17136 gnd.n4071 gnd.n1867 19.3944
R17137 gnd.n4071 gnd.n1856 19.3944
R17138 gnd.n4083 gnd.n1856 19.3944
R17139 gnd.n4083 gnd.n1854 19.3944
R17140 gnd.n4087 gnd.n1854 19.3944
R17141 gnd.n4087 gnd.n1842 19.3944
R17142 gnd.n4099 gnd.n1842 19.3944
R17143 gnd.n4099 gnd.n1840 19.3944
R17144 gnd.n4103 gnd.n1840 19.3944
R17145 gnd.n4103 gnd.n1829 19.3944
R17146 gnd.n4117 gnd.n1829 19.3944
R17147 gnd.n4117 gnd.n1827 19.3944
R17148 gnd.n4124 gnd.n1827 19.3944
R17149 gnd.n4124 gnd.n4123 19.3944
R17150 gnd.n4123 gnd.n1411 19.3944
R17151 gnd.n4431 gnd.n1411 19.3944
R17152 gnd.n4431 gnd.n4430 19.3944
R17153 gnd.n4430 gnd.n4429 19.3944
R17154 gnd.n4429 gnd.n1415 19.3944
R17155 gnd.n1635 gnd.n1415 19.3944
R17156 gnd.n1639 gnd.n1635 19.3944
R17157 gnd.n1639 gnd.n1633 19.3944
R17158 gnd.n4166 gnd.n1633 19.3944
R17159 gnd.n4166 gnd.n1631 19.3944
R17160 gnd.n4172 gnd.n1631 19.3944
R17161 gnd.n4172 gnd.n4171 19.3944
R17162 gnd.n4171 gnd.n1606 19.3944
R17163 gnd.n4197 gnd.n1606 19.3944
R17164 gnd.n4197 gnd.n1604 19.3944
R17165 gnd.n4203 gnd.n1604 19.3944
R17166 gnd.n4203 gnd.n4202 19.3944
R17167 gnd.n4202 gnd.n1578 19.3944
R17168 gnd.n4233 gnd.n1578 19.3944
R17169 gnd.n4233 gnd.n1576 19.3944
R17170 gnd.n4239 gnd.n1576 19.3944
R17171 gnd.n4239 gnd.n4238 19.3944
R17172 gnd.n4238 gnd.n1544 19.3944
R17173 gnd.n4291 gnd.n1544 19.3944
R17174 gnd.n4291 gnd.n1542 19.3944
R17175 gnd.n4303 gnd.n1542 19.3944
R17176 gnd.n4303 gnd.n4302 19.3944
R17177 gnd.n4302 gnd.n4301 19.3944
R17178 gnd.n4301 gnd.n4298 19.3944
R17179 gnd.n7116 gnd.n317 19.3944
R17180 gnd.n7114 gnd.n7113 19.3944
R17181 gnd.n7110 gnd.n7109 19.3944
R17182 gnd.n7107 gnd.n323 19.3944
R17183 gnd.n7103 gnd.n7102 19.3944
R17184 gnd.n7102 gnd.n7101 19.3944
R17185 gnd.n7101 gnd.n328 19.3944
R17186 gnd.n4829 gnd.n4828 19.3944
R17187 gnd.n4828 gnd.n4827 19.3944
R17188 gnd.n4827 gnd.n4826 19.3944
R17189 gnd.n4826 gnd.n4824 19.3944
R17190 gnd.n4824 gnd.n4821 19.3944
R17191 gnd.n4821 gnd.n4820 19.3944
R17192 gnd.n4820 gnd.n4817 19.3944
R17193 gnd.n4817 gnd.n4816 19.3944
R17194 gnd.n4816 gnd.n4813 19.3944
R17195 gnd.n4813 gnd.n4812 19.3944
R17196 gnd.n4812 gnd.n4809 19.3944
R17197 gnd.n4809 gnd.n4808 19.3944
R17198 gnd.n4808 gnd.n4805 19.3944
R17199 gnd.n4805 gnd.n4804 19.3944
R17200 gnd.n4804 gnd.n4801 19.3944
R17201 gnd.n4801 gnd.n4800 19.3944
R17202 gnd.n4800 gnd.n4797 19.3944
R17203 gnd.n4795 gnd.n4792 19.3944
R17204 gnd.n4792 gnd.n4791 19.3944
R17205 gnd.n4791 gnd.n4788 19.3944
R17206 gnd.n4788 gnd.n4787 19.3944
R17207 gnd.n4787 gnd.n4784 19.3944
R17208 gnd.n4784 gnd.n4783 19.3944
R17209 gnd.n4783 gnd.n4780 19.3944
R17210 gnd.n4780 gnd.n4779 19.3944
R17211 gnd.n4779 gnd.n4776 19.3944
R17212 gnd.n4776 gnd.n4775 19.3944
R17213 gnd.n4775 gnd.n4772 19.3944
R17214 gnd.n4772 gnd.n4771 19.3944
R17215 gnd.n4771 gnd.n4768 19.3944
R17216 gnd.n4768 gnd.n4767 19.3944
R17217 gnd.n4767 gnd.n4764 19.3944
R17218 gnd.n4764 gnd.n4763 19.3944
R17219 gnd.n4763 gnd.n4760 19.3944
R17220 gnd.n4760 gnd.n4759 19.3944
R17221 gnd.n4752 gnd.n4751 19.3944
R17222 gnd.n4751 gnd.n1010 19.3944
R17223 gnd.n4747 gnd.n1010 19.3944
R17224 gnd.n4747 gnd.n1012 19.3944
R17225 gnd.n2415 gnd.n1012 19.3944
R17226 gnd.n2417 gnd.n2415 19.3944
R17227 gnd.n2417 gnd.n2413 19.3944
R17228 gnd.n2422 gnd.n2413 19.3944
R17229 gnd.n2423 gnd.n2422 19.3944
R17230 gnd.n2425 gnd.n2423 19.3944
R17231 gnd.n2425 gnd.n2411 19.3944
R17232 gnd.n2430 gnd.n2411 19.3944
R17233 gnd.n2431 gnd.n2430 19.3944
R17234 gnd.n2433 gnd.n2431 19.3944
R17235 gnd.n2433 gnd.n2409 19.3944
R17236 gnd.n2438 gnd.n2409 19.3944
R17237 gnd.n2439 gnd.n2438 19.3944
R17238 gnd.n2441 gnd.n2439 19.3944
R17239 gnd.n2441 gnd.n2407 19.3944
R17240 gnd.n2579 gnd.n2407 19.3944
R17241 gnd.n2580 gnd.n2579 19.3944
R17242 gnd.n2581 gnd.n2580 19.3944
R17243 gnd.n2581 gnd.n2405 19.3944
R17244 gnd.n2625 gnd.n2405 19.3944
R17245 gnd.n2625 gnd.n2624 19.3944
R17246 gnd.n2624 gnd.n2623 19.3944
R17247 gnd.n2623 gnd.n2587 19.3944
R17248 gnd.n2610 gnd.n2587 19.3944
R17249 gnd.n2610 gnd.n2609 19.3944
R17250 gnd.n2609 gnd.n2608 19.3944
R17251 gnd.n2608 gnd.n2359 19.3944
R17252 gnd.n2654 gnd.n2359 19.3944
R17253 gnd.n2654 gnd.n2357 19.3944
R17254 gnd.n2659 gnd.n2357 19.3944
R17255 gnd.n2659 gnd.n2351 19.3944
R17256 gnd.n2671 gnd.n2351 19.3944
R17257 gnd.n2672 gnd.n2671 19.3944
R17258 gnd.n2673 gnd.n2672 19.3944
R17259 gnd.n2673 gnd.n2349 19.3944
R17260 gnd.n2679 gnd.n2349 19.3944
R17261 gnd.n2680 gnd.n2679 19.3944
R17262 gnd.n2684 gnd.n2680 19.3944
R17263 gnd.n2684 gnd.n2347 19.3944
R17264 gnd.n2692 gnd.n2347 19.3944
R17265 gnd.n2692 gnd.n2691 19.3944
R17266 gnd.n2691 gnd.n2690 19.3944
R17267 gnd.n2690 gnd.n2323 19.3944
R17268 gnd.n2774 gnd.n2323 19.3944
R17269 gnd.n2774 gnd.n2321 19.3944
R17270 gnd.n2779 gnd.n2321 19.3944
R17271 gnd.n2779 gnd.n2315 19.3944
R17272 gnd.n2823 gnd.n2315 19.3944
R17273 gnd.n2824 gnd.n2823 19.3944
R17274 gnd.n2866 gnd.n2289 19.3944
R17275 gnd.n2866 gnd.n2863 19.3944
R17276 gnd.n2863 gnd.n2860 19.3944
R17277 gnd.n2860 gnd.n2859 19.3944
R17278 gnd.n2859 gnd.n2856 19.3944
R17279 gnd.n2856 gnd.n2855 19.3944
R17280 gnd.n2855 gnd.n2852 19.3944
R17281 gnd.n2852 gnd.n2851 19.3944
R17282 gnd.n2851 gnd.n2848 19.3944
R17283 gnd.n2848 gnd.n2847 19.3944
R17284 gnd.n2847 gnd.n2844 19.3944
R17285 gnd.n2844 gnd.n2843 19.3944
R17286 gnd.n2843 gnd.n2840 19.3944
R17287 gnd.n2840 gnd.n2839 19.3944
R17288 gnd.n2839 gnd.n2836 19.3944
R17289 gnd.n2836 gnd.n2835 19.3944
R17290 gnd.n2835 gnd.n2832 19.3944
R17291 gnd.n2832 gnd.n2831 19.3944
R17292 gnd.n2272 gnd.n2271 19.3944
R17293 gnd.n3667 gnd.n2271 19.3944
R17294 gnd.n3667 gnd.n3666 19.3944
R17295 gnd.n3666 gnd.n3665 19.3944
R17296 gnd.n3665 gnd.n3662 19.3944
R17297 gnd.n3662 gnd.n3661 19.3944
R17298 gnd.n3661 gnd.n3658 19.3944
R17299 gnd.n3658 gnd.n3657 19.3944
R17300 gnd.n3657 gnd.n3654 19.3944
R17301 gnd.n3654 gnd.n3653 19.3944
R17302 gnd.n3653 gnd.n3650 19.3944
R17303 gnd.n3650 gnd.n3649 19.3944
R17304 gnd.n3649 gnd.n3646 19.3944
R17305 gnd.n3646 gnd.n3645 19.3944
R17306 gnd.n3645 gnd.n3642 19.3944
R17307 gnd.n2527 gnd.n2459 19.3944
R17308 gnd.n2527 gnd.n2460 19.3944
R17309 gnd.n2523 gnd.n2460 19.3944
R17310 gnd.n2523 gnd.n1032 19.3944
R17311 gnd.n4737 gnd.n1032 19.3944
R17312 gnd.n4737 gnd.n4736 19.3944
R17313 gnd.n4736 gnd.n4735 19.3944
R17314 gnd.n4735 gnd.n1036 19.3944
R17315 gnd.n4725 gnd.n1036 19.3944
R17316 gnd.n4725 gnd.n4724 19.3944
R17317 gnd.n4724 gnd.n4723 19.3944
R17318 gnd.n4723 gnd.n1055 19.3944
R17319 gnd.n4713 gnd.n1055 19.3944
R17320 gnd.n4713 gnd.n4712 19.3944
R17321 gnd.n4712 gnd.n4711 19.3944
R17322 gnd.n4711 gnd.n1076 19.3944
R17323 gnd.n4701 gnd.n1076 19.3944
R17324 gnd.n4701 gnd.n4700 19.3944
R17325 gnd.n4700 gnd.n4699 19.3944
R17326 gnd.n4699 gnd.n1095 19.3944
R17327 gnd.n4689 gnd.n1095 19.3944
R17328 gnd.n4689 gnd.n4688 19.3944
R17329 gnd.n4688 gnd.n4687 19.3944
R17330 gnd.n4687 gnd.n1118 19.3944
R17331 gnd.n4677 gnd.n1118 19.3944
R17332 gnd.n4677 gnd.n4676 19.3944
R17333 gnd.n4676 gnd.n4675 19.3944
R17334 gnd.n4675 gnd.n1136 19.3944
R17335 gnd.n4664 gnd.n1136 19.3944
R17336 gnd.n4664 gnd.n4663 19.3944
R17337 gnd.n4663 gnd.n4662 19.3944
R17338 gnd.n4662 gnd.n1155 19.3944
R17339 gnd.n4652 gnd.n1155 19.3944
R17340 gnd.n4652 gnd.n4651 19.3944
R17341 gnd.n4651 gnd.n4650 19.3944
R17342 gnd.n4650 gnd.n1174 19.3944
R17343 gnd.n4640 gnd.n1174 19.3944
R17344 gnd.n4640 gnd.n4639 19.3944
R17345 gnd.n4639 gnd.n4638 19.3944
R17346 gnd.n4638 gnd.n1196 19.3944
R17347 gnd.n4628 gnd.n1196 19.3944
R17348 gnd.n4628 gnd.n4627 19.3944
R17349 gnd.n4627 gnd.n4626 19.3944
R17350 gnd.n4626 gnd.n1216 19.3944
R17351 gnd.n4616 gnd.n1216 19.3944
R17352 gnd.n4616 gnd.n4615 19.3944
R17353 gnd.n4615 gnd.n4614 19.3944
R17354 gnd.n4614 gnd.n1238 19.3944
R17355 gnd.n4604 gnd.n1238 19.3944
R17356 gnd.n4604 gnd.n4603 19.3944
R17357 gnd.n4603 gnd.n4602 19.3944
R17358 gnd.n4602 gnd.n1259 19.3944
R17359 gnd.n4592 gnd.n1259 19.3944
R17360 gnd.n2519 gnd.n2517 19.3944
R17361 gnd.n2517 gnd.n2514 19.3944
R17362 gnd.n2514 gnd.n2513 19.3944
R17363 gnd.n2513 gnd.n2510 19.3944
R17364 gnd.n2510 gnd.n2509 19.3944
R17365 gnd.n2509 gnd.n2506 19.3944
R17366 gnd.n2506 gnd.n2505 19.3944
R17367 gnd.n2505 gnd.n2502 19.3944
R17368 gnd.n2502 gnd.n2501 19.3944
R17369 gnd.n2501 gnd.n2498 19.3944
R17370 gnd.n2498 gnd.n2497 19.3944
R17371 gnd.n2497 gnd.n2494 19.3944
R17372 gnd.n2494 gnd.n2493 19.3944
R17373 gnd.n2493 gnd.n2490 19.3944
R17374 gnd.n2490 gnd.n2489 19.3944
R17375 gnd.n2489 gnd.n2486 19.3944
R17376 gnd.n2480 gnd.n2455 19.3944
R17377 gnd.n2538 gnd.n2455 19.3944
R17378 gnd.n2538 gnd.n2453 19.3944
R17379 gnd.n2543 gnd.n2453 19.3944
R17380 gnd.n2544 gnd.n2543 19.3944
R17381 gnd.n2546 gnd.n2544 19.3944
R17382 gnd.n2546 gnd.n2451 19.3944
R17383 gnd.n2551 gnd.n2451 19.3944
R17384 gnd.n2552 gnd.n2551 19.3944
R17385 gnd.n2554 gnd.n2552 19.3944
R17386 gnd.n2554 gnd.n2449 19.3944
R17387 gnd.n2559 gnd.n2449 19.3944
R17388 gnd.n2560 gnd.n2559 19.3944
R17389 gnd.n2562 gnd.n2560 19.3944
R17390 gnd.n2562 gnd.n2447 19.3944
R17391 gnd.n2567 gnd.n2447 19.3944
R17392 gnd.n2568 gnd.n2567 19.3944
R17393 gnd.n2570 gnd.n2568 19.3944
R17394 gnd.n2570 gnd.n2445 19.3944
R17395 gnd.n2575 gnd.n2445 19.3944
R17396 gnd.n2575 gnd.n2400 19.3944
R17397 gnd.n2631 gnd.n2400 19.3944
R17398 gnd.n2631 gnd.n2630 19.3944
R17399 gnd.n2630 gnd.n2629 19.3944
R17400 gnd.n2629 gnd.n2404 19.3944
R17401 gnd.n2619 gnd.n2404 19.3944
R17402 gnd.n2619 gnd.n2618 19.3944
R17403 gnd.n2618 gnd.n2614 19.3944
R17404 gnd.n2614 gnd.n2362 19.3944
R17405 gnd.n2646 gnd.n2362 19.3944
R17406 gnd.n2646 gnd.n2360 19.3944
R17407 gnd.n2650 gnd.n2360 19.3944
R17408 gnd.n2650 gnd.n2355 19.3944
R17409 gnd.n2663 gnd.n2355 19.3944
R17410 gnd.n2663 gnd.n2353 19.3944
R17411 gnd.n2667 gnd.n2353 19.3944
R17412 gnd.n2667 gnd.n2340 19.3944
R17413 gnd.n2706 gnd.n2340 19.3944
R17414 gnd.n2706 gnd.n2341 19.3944
R17415 gnd.n2702 gnd.n2341 19.3944
R17416 gnd.n2702 gnd.n2701 19.3944
R17417 gnd.n2701 gnd.n2700 19.3944
R17418 gnd.n2700 gnd.n2346 19.3944
R17419 gnd.n2696 gnd.n2346 19.3944
R17420 gnd.n2696 gnd.n2326 19.3944
R17421 gnd.n2766 gnd.n2326 19.3944
R17422 gnd.n2766 gnd.n2324 19.3944
R17423 gnd.n2770 gnd.n2324 19.3944
R17424 gnd.n2770 gnd.n2320 19.3944
R17425 gnd.n2783 gnd.n2320 19.3944
R17426 gnd.n2783 gnd.n2317 19.3944
R17427 gnd.n2819 gnd.n2317 19.3944
R17428 gnd.n2819 gnd.n2318 19.3944
R17429 gnd.n2533 gnd.n2529 19.3944
R17430 gnd.n2533 gnd.n1021 19.3944
R17431 gnd.n4743 gnd.n1021 19.3944
R17432 gnd.n4743 gnd.n4742 19.3944
R17433 gnd.n4742 gnd.n4741 19.3944
R17434 gnd.n4741 gnd.n1025 19.3944
R17435 gnd.n4731 gnd.n1025 19.3944
R17436 gnd.n4731 gnd.n4730 19.3944
R17437 gnd.n4730 gnd.n4729 19.3944
R17438 gnd.n4729 gnd.n1046 19.3944
R17439 gnd.n4719 gnd.n1046 19.3944
R17440 gnd.n4719 gnd.n4718 19.3944
R17441 gnd.n4718 gnd.n4717 19.3944
R17442 gnd.n4717 gnd.n1065 19.3944
R17443 gnd.n4707 gnd.n1065 19.3944
R17444 gnd.n4707 gnd.n4706 19.3944
R17445 gnd.n4706 gnd.n4705 19.3944
R17446 gnd.n4705 gnd.n1086 19.3944
R17447 gnd.n4695 gnd.n1086 19.3944
R17448 gnd.n4695 gnd.n4694 19.3944
R17449 gnd.n4694 gnd.n4693 19.3944
R17450 gnd.n4693 gnd.n1107 19.3944
R17451 gnd.n4683 gnd.n4682 19.3944
R17452 gnd.n4682 gnd.n4681 19.3944
R17453 gnd.n4671 gnd.n1143 19.3944
R17454 gnd.n4669 gnd.n4668 19.3944
R17455 gnd.n4658 gnd.n1161 19.3944
R17456 gnd.n4658 gnd.n4657 19.3944
R17457 gnd.n4657 gnd.n4656 19.3944
R17458 gnd.n4656 gnd.n1164 19.3944
R17459 gnd.n4646 gnd.n1164 19.3944
R17460 gnd.n4646 gnd.n4645 19.3944
R17461 gnd.n4645 gnd.n4644 19.3944
R17462 gnd.n4644 gnd.n1185 19.3944
R17463 gnd.n4634 gnd.n1185 19.3944
R17464 gnd.n4634 gnd.n4633 19.3944
R17465 gnd.n4633 gnd.n4632 19.3944
R17466 gnd.n4632 gnd.n1206 19.3944
R17467 gnd.n4622 gnd.n1206 19.3944
R17468 gnd.n4622 gnd.n4621 19.3944
R17469 gnd.n4621 gnd.n4620 19.3944
R17470 gnd.n4620 gnd.n1227 19.3944
R17471 gnd.n4610 gnd.n1227 19.3944
R17472 gnd.n4610 gnd.n4609 19.3944
R17473 gnd.n4609 gnd.n4608 19.3944
R17474 gnd.n4608 gnd.n1248 19.3944
R17475 gnd.n4598 gnd.n1248 19.3944
R17476 gnd.n4598 gnd.n4597 19.3944
R17477 gnd.n4597 gnd.n4596 19.3944
R17478 gnd.n6423 gnd.n730 19.3944
R17479 gnd.n6423 gnd.n6422 19.3944
R17480 gnd.n6422 gnd.n6421 19.3944
R17481 gnd.n6421 gnd.n734 19.3944
R17482 gnd.n6415 gnd.n734 19.3944
R17483 gnd.n6415 gnd.n6414 19.3944
R17484 gnd.n6414 gnd.n6413 19.3944
R17485 gnd.n6413 gnd.n742 19.3944
R17486 gnd.n6407 gnd.n742 19.3944
R17487 gnd.n6407 gnd.n6406 19.3944
R17488 gnd.n6406 gnd.n6405 19.3944
R17489 gnd.n6405 gnd.n750 19.3944
R17490 gnd.n6399 gnd.n750 19.3944
R17491 gnd.n6399 gnd.n6398 19.3944
R17492 gnd.n6398 gnd.n6397 19.3944
R17493 gnd.n6397 gnd.n758 19.3944
R17494 gnd.n6391 gnd.n758 19.3944
R17495 gnd.n6391 gnd.n6390 19.3944
R17496 gnd.n6390 gnd.n6389 19.3944
R17497 gnd.n6389 gnd.n766 19.3944
R17498 gnd.n6383 gnd.n766 19.3944
R17499 gnd.n6383 gnd.n6382 19.3944
R17500 gnd.n6382 gnd.n6381 19.3944
R17501 gnd.n6381 gnd.n774 19.3944
R17502 gnd.n6375 gnd.n774 19.3944
R17503 gnd.n6375 gnd.n6374 19.3944
R17504 gnd.n6374 gnd.n6373 19.3944
R17505 gnd.n6373 gnd.n782 19.3944
R17506 gnd.n6367 gnd.n782 19.3944
R17507 gnd.n6367 gnd.n6366 19.3944
R17508 gnd.n6366 gnd.n6365 19.3944
R17509 gnd.n6365 gnd.n790 19.3944
R17510 gnd.n6359 gnd.n790 19.3944
R17511 gnd.n6359 gnd.n6358 19.3944
R17512 gnd.n6358 gnd.n6357 19.3944
R17513 gnd.n6357 gnd.n798 19.3944
R17514 gnd.n6351 gnd.n798 19.3944
R17515 gnd.n6351 gnd.n6350 19.3944
R17516 gnd.n6350 gnd.n6349 19.3944
R17517 gnd.n6349 gnd.n806 19.3944
R17518 gnd.n6343 gnd.n806 19.3944
R17519 gnd.n6343 gnd.n6342 19.3944
R17520 gnd.n6342 gnd.n6341 19.3944
R17521 gnd.n6341 gnd.n814 19.3944
R17522 gnd.n6335 gnd.n814 19.3944
R17523 gnd.n6335 gnd.n6334 19.3944
R17524 gnd.n6334 gnd.n6333 19.3944
R17525 gnd.n6333 gnd.n822 19.3944
R17526 gnd.n6327 gnd.n822 19.3944
R17527 gnd.n6327 gnd.n6326 19.3944
R17528 gnd.n6326 gnd.n6325 19.3944
R17529 gnd.n6325 gnd.n830 19.3944
R17530 gnd.n6319 gnd.n830 19.3944
R17531 gnd.n6319 gnd.n6318 19.3944
R17532 gnd.n6318 gnd.n6317 19.3944
R17533 gnd.n6317 gnd.n838 19.3944
R17534 gnd.n6311 gnd.n838 19.3944
R17535 gnd.n6311 gnd.n6310 19.3944
R17536 gnd.n6310 gnd.n6309 19.3944
R17537 gnd.n6309 gnd.n846 19.3944
R17538 gnd.n6303 gnd.n846 19.3944
R17539 gnd.n6303 gnd.n6302 19.3944
R17540 gnd.n6302 gnd.n6301 19.3944
R17541 gnd.n6301 gnd.n854 19.3944
R17542 gnd.n6295 gnd.n854 19.3944
R17543 gnd.n6295 gnd.n6294 19.3944
R17544 gnd.n6294 gnd.n6293 19.3944
R17545 gnd.n6293 gnd.n862 19.3944
R17546 gnd.n6287 gnd.n862 19.3944
R17547 gnd.n6287 gnd.n6286 19.3944
R17548 gnd.n6286 gnd.n6285 19.3944
R17549 gnd.n6285 gnd.n870 19.3944
R17550 gnd.n6279 gnd.n870 19.3944
R17551 gnd.n6279 gnd.n6278 19.3944
R17552 gnd.n6278 gnd.n6277 19.3944
R17553 gnd.n6277 gnd.n878 19.3944
R17554 gnd.n6271 gnd.n878 19.3944
R17555 gnd.n6271 gnd.n6270 19.3944
R17556 gnd.n6270 gnd.n6269 19.3944
R17557 gnd.n6269 gnd.n886 19.3944
R17558 gnd.n6263 gnd.n886 19.3944
R17559 gnd.n6263 gnd.n6262 19.3944
R17560 gnd.n6262 gnd.n6261 19.3944
R17561 gnd.n6261 gnd.n894 19.3944
R17562 gnd.n4587 gnd.n4586 19.3944
R17563 gnd.n4586 gnd.n4585 19.3944
R17564 gnd.n4585 gnd.n1282 19.3944
R17565 gnd.n4581 gnd.n1282 19.3944
R17566 gnd.n4581 gnd.n4580 19.3944
R17567 gnd.n4580 gnd.n4579 19.3944
R17568 gnd.n4579 gnd.n1287 19.3944
R17569 gnd.n4575 gnd.n1287 19.3944
R17570 gnd.n4575 gnd.n4574 19.3944
R17571 gnd.n4574 gnd.n4573 19.3944
R17572 gnd.n4573 gnd.n1292 19.3944
R17573 gnd.n4569 gnd.n1292 19.3944
R17574 gnd.n4569 gnd.n4568 19.3944
R17575 gnd.n4568 gnd.n4567 19.3944
R17576 gnd.n4567 gnd.n1297 19.3944
R17577 gnd.n4563 gnd.n1297 19.3944
R17578 gnd.n4563 gnd.n4562 19.3944
R17579 gnd.n4562 gnd.n4561 19.3944
R17580 gnd.n4561 gnd.n1302 19.3944
R17581 gnd.n4557 gnd.n1302 19.3944
R17582 gnd.n4557 gnd.n4556 19.3944
R17583 gnd.n4556 gnd.n4555 19.3944
R17584 gnd.n4555 gnd.n1307 19.3944
R17585 gnd.n4551 gnd.n1307 19.3944
R17586 gnd.n4551 gnd.n4550 19.3944
R17587 gnd.n4550 gnd.n4549 19.3944
R17588 gnd.n4549 gnd.n1312 19.3944
R17589 gnd.n4545 gnd.n1312 19.3944
R17590 gnd.n4545 gnd.n4544 19.3944
R17591 gnd.n4544 gnd.n4543 19.3944
R17592 gnd.n4543 gnd.n1317 19.3944
R17593 gnd.n4539 gnd.n1317 19.3944
R17594 gnd.n4539 gnd.n4538 19.3944
R17595 gnd.n4538 gnd.n4537 19.3944
R17596 gnd.n4537 gnd.n1322 19.3944
R17597 gnd.n4533 gnd.n1322 19.3944
R17598 gnd.n4533 gnd.n4532 19.3944
R17599 gnd.n4532 gnd.n4531 19.3944
R17600 gnd.n4531 gnd.n1327 19.3944
R17601 gnd.n4527 gnd.n1327 19.3944
R17602 gnd.n4527 gnd.n4526 19.3944
R17603 gnd.n4526 gnd.n4525 19.3944
R17604 gnd.n4525 gnd.n1332 19.3944
R17605 gnd.n4521 gnd.n1332 19.3944
R17606 gnd.n4521 gnd.n4520 19.3944
R17607 gnd.n4520 gnd.n4519 19.3944
R17608 gnd.n4519 gnd.n1337 19.3944
R17609 gnd.n4515 gnd.n1337 19.3944
R17610 gnd.n4515 gnd.n4514 19.3944
R17611 gnd.n4514 gnd.n4513 19.3944
R17612 gnd.n4513 gnd.n1342 19.3944
R17613 gnd.n4509 gnd.n1342 19.3944
R17614 gnd.n4509 gnd.n4508 19.3944
R17615 gnd.n4508 gnd.n4507 19.3944
R17616 gnd.n4507 gnd.n1347 19.3944
R17617 gnd.n4503 gnd.n1347 19.3944
R17618 gnd.n4503 gnd.n4502 19.3944
R17619 gnd.n4502 gnd.n4501 19.3944
R17620 gnd.n4501 gnd.n1352 19.3944
R17621 gnd.n4497 gnd.n1352 19.3944
R17622 gnd.n4497 gnd.n4496 19.3944
R17623 gnd.n4496 gnd.n4495 19.3944
R17624 gnd.n4495 gnd.n1357 19.3944
R17625 gnd.n4491 gnd.n1357 19.3944
R17626 gnd.n4491 gnd.n4490 19.3944
R17627 gnd.n4490 gnd.n4489 19.3944
R17628 gnd.n4489 gnd.n1362 19.3944
R17629 gnd.n4485 gnd.n1362 19.3944
R17630 gnd.n4485 gnd.n4484 19.3944
R17631 gnd.n4484 gnd.n4483 19.3944
R17632 gnd.n4483 gnd.n1367 19.3944
R17633 gnd.n4479 gnd.n1367 19.3944
R17634 gnd.n4479 gnd.n4478 19.3944
R17635 gnd.n4478 gnd.n4477 19.3944
R17636 gnd.n4477 gnd.n1372 19.3944
R17637 gnd.n4473 gnd.n1372 19.3944
R17638 gnd.n4473 gnd.n4472 19.3944
R17639 gnd.n4472 gnd.n4471 19.3944
R17640 gnd.n4471 gnd.n1377 19.3944
R17641 gnd.n4467 gnd.n1377 19.3944
R17642 gnd.n4467 gnd.n4466 19.3944
R17643 gnd.n4466 gnd.n4465 19.3944
R17644 gnd.n4465 gnd.n1382 19.3944
R17645 gnd.n4461 gnd.n1382 19.3944
R17646 gnd.n4461 gnd.n4460 19.3944
R17647 gnd.n4460 gnd.n4459 19.3944
R17648 gnd.n4459 gnd.n1387 19.3944
R17649 gnd.n4455 gnd.n1387 19.3944
R17650 gnd.n4455 gnd.n4454 19.3944
R17651 gnd.n4454 gnd.n4453 19.3944
R17652 gnd.n4453 gnd.n1392 19.3944
R17653 gnd.n4449 gnd.n1392 19.3944
R17654 gnd.n4449 gnd.n4448 19.3944
R17655 gnd.n4448 gnd.n4447 19.3944
R17656 gnd.n4447 gnd.n1397 19.3944
R17657 gnd.n4443 gnd.n1397 19.3944
R17658 gnd.n4443 gnd.n4442 19.3944
R17659 gnd.n4442 gnd.n4441 19.3944
R17660 gnd.n4441 gnd.n1402 19.3944
R17661 gnd.n4437 gnd.n1402 19.3944
R17662 gnd.n4437 gnd.n4436 19.3944
R17663 gnd.n4142 gnd.n1819 19.3944
R17664 gnd.n4138 gnd.n1819 19.3944
R17665 gnd.n4138 gnd.n4137 19.3944
R17666 gnd.n1735 gnd.n1719 19.3944
R17667 gnd.n1735 gnd.n1717 19.3944
R17668 gnd.n1741 gnd.n1717 19.3944
R17669 gnd.n1741 gnd.n1712 19.3944
R17670 gnd.n1754 gnd.n1712 19.3944
R17671 gnd.n1754 gnd.n1710 19.3944
R17672 gnd.n1760 gnd.n1710 19.3944
R17673 gnd.n1760 gnd.n1705 19.3944
R17674 gnd.n1773 gnd.n1705 19.3944
R17675 gnd.n1773 gnd.n1703 19.3944
R17676 gnd.n1779 gnd.n1703 19.3944
R17677 gnd.n1779 gnd.n1699 19.3944
R17678 gnd.n1789 gnd.n1699 19.3944
R17679 gnd.n1789 gnd.n1697 19.3944
R17680 gnd.n1795 gnd.n1697 19.3944
R17681 gnd.n1795 gnd.n1687 19.3944
R17682 gnd.n1803 gnd.n1687 19.3944
R17683 gnd.n1803 gnd.n1685 19.3944
R17684 gnd.n4153 gnd.n1685 19.3944
R17685 gnd.n4153 gnd.n4152 19.3944
R17686 gnd.n4152 gnd.n4151 19.3944
R17687 gnd.n4151 gnd.n1811 19.3944
R17688 gnd.n4147 gnd.n1811 19.3944
R17689 gnd.n4147 gnd.n4146 19.3944
R17690 gnd.t124 gnd.n2066 19.1199
R17691 gnd.t117 gnd.n1911 19.1199
R17692 gnd.t316 gnd.n5060 18.8012
R17693 gnd.n5664 gnd.t329 18.8012
R17694 gnd.n5509 gnd.n5508 18.4825
R17695 gnd.n4691 gnd.n1109 18.4825
R17696 gnd.n2633 gnd.n1112 18.4825
R17697 gnd.n2627 gnd.n1122 18.4825
R17698 gnd.n4679 gnd.n1128 18.4825
R17699 gnd.n2621 gnd.n2599 18.4825
R17700 gnd.n4673 gnd.n1138 18.4825
R17701 gnd.n4666 gnd.n1146 18.4825
R17702 gnd.n2644 gnd.n1149 18.4825
R17703 gnd.n2652 gnd.n1159 18.4825
R17704 gnd.n4654 gnd.n1166 18.4825
R17705 gnd.n2661 gnd.n2356 18.4825
R17706 gnd.n4648 gnd.n1176 18.4825
R17707 gnd.n4642 gnd.n1187 18.4825
R17708 gnd.n2708 gnd.n1190 18.4825
R17709 gnd.n2677 gnd.n1200 18.4825
R17710 gnd.n4630 gnd.n1208 18.4825
R17711 gnd.n2682 gnd.n2681 18.4825
R17712 gnd.n4624 gnd.n1218 18.4825
R17713 gnd.n4618 gnd.n1229 18.4825
R17714 gnd.n2764 gnd.n1232 18.4825
R17715 gnd.n2772 gnd.n1242 18.4825
R17716 gnd.n4606 gnd.n1250 18.4825
R17717 gnd.n2781 gnd.n1253 18.4825
R17718 gnd.n4600 gnd.n1261 18.4825
R17719 gnd.n2821 gnd.n2316 18.4825
R17720 gnd.n4594 gnd.n1270 18.4825
R17721 gnd.n3873 gnd.n2038 18.4825
R17722 gnd.n3135 gnd.n1947 18.4825
R17723 gnd.n4349 gnd.n1499 18.4825
R17724 gnd.n4164 gnd.n1647 18.4825
R17725 gnd.n4163 gnd.n1625 18.4825
R17726 gnd.n4175 gnd.n4174 18.4825
R17727 gnd.n1628 gnd.n1615 18.4825
R17728 gnd.n4185 gnd.n1617 18.4825
R17729 gnd.n4194 gnd.n1597 18.4825
R17730 gnd.n4206 gnd.n4205 18.4825
R17731 gnd.n4216 gnd.n1590 18.4825
R17732 gnd.n4231 gnd.n1580 18.4825
R17733 gnd.n4230 gnd.n1570 18.4825
R17734 gnd.n4243 gnd.n4241 18.4825
R17735 gnd.n4253 gnd.n1563 18.4825
R17736 gnd.n4289 gnd.n1546 18.4825
R17737 gnd.n4306 gnd.n4305 18.4825
R17738 gnd.n1540 gnd.n1538 18.4825
R17739 gnd.n4314 gnd.n1529 18.4825
R17740 gnd.n4276 gnd.n278 18.4825
R17741 gnd.n7119 gnd.n7118 18.4825
R17742 gnd.n314 gnd.n307 18.4825
R17743 gnd.n7132 gnd.n304 18.4825
R17744 gnd.n321 gnd.n320 18.4825
R17745 gnd.n7198 gnd.n294 18.4825
R17746 gnd.n7203 gnd.n296 18.4825
R17747 gnd.n7226 gnd.n265 18.4825
R17748 gnd.n7187 gnd.n256 18.4825
R17749 gnd.n4394 gnd.n4393 18.4247
R17750 gnd.n3642 gnd.n3641 18.4247
R17751 gnd.n7338 gnd.n7337 18.2308
R17752 gnd.n1799 gnd.n1798 18.2308
R17753 gnd.n3680 gnd.n2225 18.2308
R17754 gnd.n2486 gnd.n2479 18.2308
R17755 gnd.t317 gnd.n5104 18.1639
R17756 gnd.n6258 gnd.n6257 18.1639
R17757 gnd.n3569 gnd.n2996 17.6395
R17758 gnd.n3378 gnd.n3377 17.6395
R17759 gnd.n5131 gnd.t319 17.5266
R17760 gnd.t251 gnd.n1029 17.5266
R17761 gnd.n4612 gnd.t203 17.5266
R17762 gnd.t24 gnd.n2017 17.5266
R17763 gnd.n3450 gnd.t30 17.5266
R17764 gnd.n1671 gnd.t249 17.5266
R17765 gnd.n7290 gnd.t230 17.5266
R17766 gnd.n5089 gnd.t313 16.8893
R17767 gnd.t210 gnd.n1070 16.8893
R17768 gnd.n4636 gnd.t228 16.8893
R17769 gnd.n3809 gnd.t61 16.8893
R17770 gnd.t52 gnd.n2044 16.8893
R17771 gnd.n3417 gnd.t303 16.8893
R17772 gnd.n1890 gnd.t28 16.8893
R17773 gnd.n1573 gnd.t201 16.8893
R17774 gnd.n7258 gnd.t244 16.8893
R17775 gnd.t54 gnd.n2060 16.5706
R17776 gnd.n3403 gnd.t6 16.5706
R17777 gnd.n5358 gnd.t106 16.2519
R17778 gnd.n5654 gnd.t307 16.2519
R17779 gnd.n4660 gnd.t267 16.2519
R17780 gnd.n7219 gnd.t239 16.2519
R17781 gnd.n2875 gnd.n2874 16.0975
R17782 gnd.n3224 gnd.n3223 16.0975
R17783 gnd.n2930 gnd.n2929 16.0975
R17784 gnd.n3218 gnd.n3217 16.0975
R17785 gnd.n3857 gnd.n2052 15.9333
R17786 gnd.n3493 gnd.t5 15.9333
R17787 gnd.n3479 gnd.n1987 15.9333
R17788 gnd.n3929 gnd.n1987 15.9333
R17789 gnd.t66 gnd.n1973 15.9333
R17790 gnd.n3411 gnd.n3410 15.9333
R17791 gnd.n6064 gnd.n6062 15.6674
R17792 gnd.n6032 gnd.n6030 15.6674
R17793 gnd.n6000 gnd.n5998 15.6674
R17794 gnd.n5969 gnd.n5967 15.6674
R17795 gnd.n5937 gnd.n5935 15.6674
R17796 gnd.n5905 gnd.n5903 15.6674
R17797 gnd.n5873 gnd.n5871 15.6674
R17798 gnd.n5842 gnd.n5840 15.6674
R17799 gnd.n5349 gnd.t106 15.6146
R17800 gnd.t69 gnd.n6243 15.6146
R17801 gnd.n6147 gnd.t91 15.6146
R17802 gnd.n4685 gnd.t181 15.6146
R17803 gnd.n7192 gnd.t188 15.6146
R17804 gnd.n3495 gnd.t67 15.296
R17805 gnd.t7 gnd.n1975 15.296
R17806 gnd.n3180 gnd.n3179 15.0827
R17807 gnd.n2903 gnd.n2898 15.0481
R17808 gnd.n3190 gnd.n3189 15.0481
R17809 gnd.n5792 gnd.t320 14.9773
R17810 gnd.n4709 gnd.t210 14.9773
R17811 gnd.n2101 gnd.t61 14.9773
R17812 gnd.n4049 gnd.t28 14.9773
R17813 gnd.n241 gnd.t244 14.9773
R17814 gnd.n3559 gnd.t120 14.6587
R17815 gnd.t4 gnd.n2058 14.6587
R17816 gnd.n3849 gnd.n2060 14.6587
R17817 gnd.n3525 gnd.n3524 14.6587
R17818 gnd.n3985 gnd.n1939 14.6587
R17819 gnd.n3403 gnd.n3154 14.6587
R17820 gnd.n3156 gnd.t20 14.6587
R17821 gnd.t113 gnd.n1903 14.6587
R17822 gnd.t36 gnd.n4933 14.34
R17823 gnd.t318 gnd.n898 14.34
R17824 gnd.n4733 gnd.t251 14.34
R17825 gnd.n211 gnd.t230 14.34
R17826 gnd.n5474 gnd.t21 13.7027
R17827 gnd.t190 gnd.n1101 13.7027
R17828 gnd.n7098 gnd.t177 13.7027
R17829 gnd.n5215 gnd.n5214 13.5763
R17830 gnd.n6203 gnd.n4865 13.5763
R17831 gnd.n4356 gnd.n1493 13.5763
R17832 gnd.n7390 gnd.n7389 13.5763
R17833 gnd.n4759 gnd.n1007 13.5763
R17834 gnd.n2831 gnd.n2828 13.5763
R17835 gnd.n5509 gnd.n5161 13.384
R17836 gnd.n4697 gnd.n1101 13.384
R17837 gnd.n2577 gnd.n1109 13.384
R17838 gnd.n4691 gnd.n1112 13.384
R17839 gnd.n2634 gnd.n2633 13.384
R17840 gnd.n4685 gnd.n1122 13.384
R17841 gnd.n2627 gnd.n1128 13.384
R17842 gnd.n2621 gnd.n1138 13.384
R17843 gnd.n4673 gnd.n1141 13.384
R17844 gnd.n2612 gnd.n1146 13.384
R17845 gnd.n4666 gnd.n1149 13.384
R17846 gnd.n2644 gnd.n2643 13.384
R17847 gnd.n4660 gnd.n1159 13.384
R17848 gnd.n2652 gnd.n1166 13.384
R17849 gnd.n2661 gnd.n1176 13.384
R17850 gnd.n4648 gnd.n1179 13.384
R17851 gnd.n2669 gnd.n1187 13.384
R17852 gnd.n4642 gnd.n1190 13.384
R17853 gnd.n2709 gnd.n2708 13.384
R17854 gnd.n4636 gnd.n1200 13.384
R17855 gnd.n2677 gnd.n1208 13.384
R17856 gnd.n2682 gnd.n1218 13.384
R17857 gnd.n4624 gnd.n1221 13.384
R17858 gnd.n2694 gnd.n1229 13.384
R17859 gnd.n4618 gnd.n1232 13.384
R17860 gnd.n2764 gnd.n2763 13.384
R17861 gnd.n4612 gnd.n1242 13.384
R17862 gnd.n2772 gnd.n1250 13.384
R17863 gnd.n4606 gnd.n1253 13.384
R17864 gnd.n2781 gnd.n1261 13.384
R17865 gnd.n2821 gnd.n1270 13.384
R17866 gnd.n4594 gnd.n1273 13.384
R17867 gnd.n3841 gnd.n2067 13.384
R17868 gnd.n3042 gnd.n2038 13.384
R17869 gnd.n3494 gnd.n3493 13.384
R17870 gnd.n3921 gnd.t40 13.384
R17871 gnd.t0 gnd.n3095 13.384
R17872 gnd.n3945 gnd.n1973 13.384
R17873 gnd.n3977 gnd.n1947 13.384
R17874 gnd.n3396 gnd.n3395 13.384
R17875 gnd.n4349 gnd.n1497 13.384
R17876 gnd.n1647 gnd.n1499 13.384
R17877 gnd.n4175 gnd.n1625 13.384
R17878 gnd.n4174 gnd.n1628 13.384
R17879 gnd.n4185 gnd.n1615 13.384
R17880 gnd.n1671 gnd.n1617 13.384
R17881 gnd.n4195 gnd.n4194 13.384
R17882 gnd.n4206 gnd.n1597 13.384
R17883 gnd.n4205 gnd.n1601 13.384
R17884 gnd.n4216 gnd.n1588 13.384
R17885 gnd.n1590 gnd.n1580 13.384
R17886 gnd.n4243 gnd.n1570 13.384
R17887 gnd.n4241 gnd.n1573 13.384
R17888 gnd.n4253 gnd.n1561 13.384
R17889 gnd.n1563 gnd.n1546 13.384
R17890 gnd.n4289 gnd.n4288 13.384
R17891 gnd.n4306 gnd.n1535 13.384
R17892 gnd.n4305 gnd.n1538 13.384
R17893 gnd.n4276 gnd.n1529 13.384
R17894 gnd.n7219 gnd.n278 13.384
R17895 gnd.n7119 gnd.n312 13.384
R17896 gnd.n7118 gnd.n314 13.384
R17897 gnd.n7127 gnd.n307 13.384
R17898 gnd.n7132 gnd.n302 13.384
R17899 gnd.n320 gnd.n304 13.384
R17900 gnd.n7203 gnd.n294 13.384
R17901 gnd.n7192 gnd.n296 13.384
R17902 gnd.n7226 gnd.n263 13.384
R17903 gnd.n7187 gnd.n265 13.384
R17904 gnd.n7234 gnd.n256 13.384
R17905 gnd.n7098 gnd.n248 13.384
R17906 gnd.n2914 gnd.n2895 13.1884
R17907 gnd.n2909 gnd.n2908 13.1884
R17908 gnd.n2908 gnd.n2907 13.1884
R17909 gnd.n3183 gnd.n3178 13.1884
R17910 gnd.n3184 gnd.n3183 13.1884
R17911 gnd.n2910 gnd.n2897 13.146
R17912 gnd.n2906 gnd.n2897 13.146
R17913 gnd.n3182 gnd.n3181 13.146
R17914 gnd.n3182 gnd.n3177 13.146
R17915 gnd.t253 gnd.n1141 13.0654
R17916 gnd.t257 gnd.n302 13.0654
R17917 gnd.n6065 gnd.n6061 12.8005
R17918 gnd.n6033 gnd.n6029 12.8005
R17919 gnd.n6001 gnd.n5997 12.8005
R17920 gnd.n5970 gnd.n5966 12.8005
R17921 gnd.n5938 gnd.n5934 12.8005
R17922 gnd.n5906 gnd.n5902 12.8005
R17923 gnd.n5874 gnd.n5870 12.8005
R17924 gnd.n5843 gnd.n5839 12.8005
R17925 gnd.t196 gnd.n1179 12.4281
R17926 gnd.n3753 gnd.t14 12.4281
R17927 gnd.n1845 gnd.t16 12.4281
R17928 gnd.t233 gnd.n1535 12.4281
R17929 gnd.n5214 gnd.n5209 12.4126
R17930 gnd.n6208 gnd.n4865 12.4126
R17931 gnd.n4352 gnd.n1493 12.4126
R17932 gnd.n7389 gnd.n178 12.4126
R17933 gnd.n4755 gnd.n1007 12.4126
R17934 gnd.n2828 gnd.n2311 12.4126
R17935 gnd.n2996 gnd.n2995 12.1761
R17936 gnd.n3377 gnd.n3376 12.1761
R17937 gnd.n3670 gnd.n2234 12.1094
R17938 gnd.n3833 gnd.n2075 12.1094
R17939 gnd.n3054 gnd.n2032 12.1094
R17940 gnd.n3073 gnd.n2008 12.1094
R17941 gnd.n3953 gnd.n1966 12.1094
R17942 gnd.n3969 gnd.n1953 12.1094
R17943 gnd.t156 gnd.n1912 12.1094
R17944 gnd.n3256 gnd.t77 12.1094
R17945 gnd.n4425 gnd.n1446 12.1094
R17946 gnd.n6069 gnd.n6068 12.0247
R17947 gnd.n6037 gnd.n6036 12.0247
R17948 gnd.n6005 gnd.n6004 12.0247
R17949 gnd.n5974 gnd.n5973 12.0247
R17950 gnd.n5942 gnd.n5941 12.0247
R17951 gnd.n5910 gnd.n5909 12.0247
R17952 gnd.n5878 gnd.n5877 12.0247
R17953 gnd.n5847 gnd.n5846 12.0247
R17954 gnd.t184 gnd.n1221 11.7908
R17955 gnd.t222 gnd.n1588 11.7908
R17956 gnd.n3029 gnd.t23 11.4721
R17957 gnd.n3516 gnd.t51 11.4721
R17958 gnd.t305 gnd.n1945 11.4721
R17959 gnd.n3993 gnd.t18 11.4721
R17960 gnd.n6072 gnd.n6059 11.249
R17961 gnd.n6040 gnd.n6027 11.249
R17962 gnd.n6008 gnd.n5995 11.249
R17963 gnd.n5977 gnd.n5964 11.249
R17964 gnd.n5945 gnd.n5932 11.249
R17965 gnd.n5913 gnd.n5900 11.249
R17966 gnd.n5881 gnd.n5868 11.249
R17967 gnd.n5850 gnd.n5837 11.249
R17968 gnd.n5582 gnd.t21 11.1535
R17969 gnd.n2024 gnd.n2015 10.8348
R17970 gnd.n3961 gnd.n1959 10.8348
R17971 gnd.n1905 gnd.n1896 10.8348
R17972 gnd.n3311 gnd.n3221 10.6151
R17973 gnd.n3311 gnd.n3310 10.6151
R17974 gnd.n3308 gnd.n3225 10.6151
R17975 gnd.n3303 gnd.n3225 10.6151
R17976 gnd.n3303 gnd.n3302 10.6151
R17977 gnd.n3302 gnd.n3301 10.6151
R17978 gnd.n3301 gnd.n3228 10.6151
R17979 gnd.n3296 gnd.n3228 10.6151
R17980 gnd.n3296 gnd.n3295 10.6151
R17981 gnd.n3295 gnd.n3294 10.6151
R17982 gnd.n3294 gnd.n3231 10.6151
R17983 gnd.n3289 gnd.n3231 10.6151
R17984 gnd.n3289 gnd.n3288 10.6151
R17985 gnd.n3288 gnd.n3287 10.6151
R17986 gnd.n3287 gnd.n3234 10.6151
R17987 gnd.n3282 gnd.n3234 10.6151
R17988 gnd.n3282 gnd.n3281 10.6151
R17989 gnd.n3281 gnd.n3280 10.6151
R17990 gnd.n3280 gnd.n3237 10.6151
R17991 gnd.n3275 gnd.n3237 10.6151
R17992 gnd.n3275 gnd.n3274 10.6151
R17993 gnd.n3274 gnd.n3273 10.6151
R17994 gnd.n3273 gnd.n3240 10.6151
R17995 gnd.n3268 gnd.n3240 10.6151
R17996 gnd.n3268 gnd.n3267 10.6151
R17997 gnd.n3267 gnd.n3266 10.6151
R17998 gnd.n3266 gnd.n3243 10.6151
R17999 gnd.n3261 gnd.n3243 10.6151
R18000 gnd.n3261 gnd.n3260 10.6151
R18001 gnd.n3260 gnd.n3259 10.6151
R18002 gnd.n3001 gnd.n2890 10.6151
R18003 gnd.n3563 gnd.n3001 10.6151
R18004 gnd.n3563 gnd.n3562 10.6151
R18005 gnd.n3562 gnd.n3561 10.6151
R18006 gnd.n3561 gnd.n3002 10.6151
R18007 gnd.n3012 gnd.n3002 10.6151
R18008 gnd.n3550 gnd.n3012 10.6151
R18009 gnd.n3550 gnd.n3549 10.6151
R18010 gnd.n3549 gnd.n3548 10.6151
R18011 gnd.n3548 gnd.n3013 10.6151
R18012 gnd.n3025 gnd.n3013 10.6151
R18013 gnd.n3026 gnd.n3025 10.6151
R18014 gnd.n3536 gnd.n3026 10.6151
R18015 gnd.n3536 gnd.n3535 10.6151
R18016 gnd.n3535 gnd.n3534 10.6151
R18017 gnd.n3534 gnd.n3027 10.6151
R18018 gnd.n3045 gnd.n3027 10.6151
R18019 gnd.n3046 gnd.n3045 10.6151
R18020 gnd.n3047 gnd.n3046 10.6151
R18021 gnd.n3048 gnd.n3047 10.6151
R18022 gnd.n3050 gnd.n3048 10.6151
R18023 gnd.n3051 gnd.n3050 10.6151
R18024 gnd.n3513 gnd.n3051 10.6151
R18025 gnd.n3513 gnd.n3512 10.6151
R18026 gnd.n3512 gnd.n3511 10.6151
R18027 gnd.n3511 gnd.n3052 10.6151
R18028 gnd.n3067 gnd.n3052 10.6151
R18029 gnd.n3070 gnd.n3067 10.6151
R18030 gnd.n3071 gnd.n3070 10.6151
R18031 gnd.n3072 gnd.n3071 10.6151
R18032 gnd.n3072 gnd.n3065 10.6151
R18033 gnd.n3078 gnd.n3065 10.6151
R18034 gnd.n3079 gnd.n3078 10.6151
R18035 gnd.n3491 gnd.n3079 10.6151
R18036 gnd.n3491 gnd.n3490 10.6151
R18037 gnd.n3490 gnd.n3489 10.6151
R18038 gnd.n3489 gnd.n3080 10.6151
R18039 gnd.n3092 gnd.n3080 10.6151
R18040 gnd.n3477 gnd.n3092 10.6151
R18041 gnd.n3477 gnd.n3476 10.6151
R18042 gnd.n3476 gnd.n3475 10.6151
R18043 gnd.n3475 gnd.n3093 10.6151
R18044 gnd.n3105 gnd.n3093 10.6151
R18045 gnd.n3106 gnd.n3105 10.6151
R18046 gnd.n3462 gnd.n3106 10.6151
R18047 gnd.n3462 gnd.n3461 10.6151
R18048 gnd.n3461 gnd.n3460 10.6151
R18049 gnd.n3460 gnd.n3107 10.6151
R18050 gnd.n3118 gnd.n3107 10.6151
R18051 gnd.n3119 gnd.n3118 10.6151
R18052 gnd.n3447 gnd.n3119 10.6151
R18053 gnd.n3447 gnd.n3446 10.6151
R18054 gnd.n3446 gnd.n3445 10.6151
R18055 gnd.n3445 gnd.n3120 10.6151
R18056 gnd.n3435 gnd.n3120 10.6151
R18057 gnd.n3435 gnd.n3434 10.6151
R18058 gnd.n3434 gnd.n3433 10.6151
R18059 gnd.n3433 gnd.n3129 10.6151
R18060 gnd.n3138 gnd.n3129 10.6151
R18061 gnd.n3422 gnd.n3138 10.6151
R18062 gnd.n3422 gnd.n3421 10.6151
R18063 gnd.n3421 gnd.n3420 10.6151
R18064 gnd.n3420 gnd.n3139 10.6151
R18065 gnd.n3150 gnd.n3139 10.6151
R18066 gnd.n3151 gnd.n3150 10.6151
R18067 gnd.n3407 gnd.n3151 10.6151
R18068 gnd.n3407 gnd.n3406 10.6151
R18069 gnd.n3406 gnd.n3405 10.6151
R18070 gnd.n3405 gnd.n3152 10.6151
R18071 gnd.n3164 gnd.n3152 10.6151
R18072 gnd.n3165 gnd.n3164 10.6151
R18073 gnd.n3392 gnd.n3165 10.6151
R18074 gnd.n3392 gnd.n3391 10.6151
R18075 gnd.n3391 gnd.n3390 10.6151
R18076 gnd.n3390 gnd.n3166 10.6151
R18077 gnd.n3249 gnd.n3166 10.6151
R18078 gnd.n3251 gnd.n3249 10.6151
R18079 gnd.n3252 gnd.n3251 10.6151
R18080 gnd.n3253 gnd.n3252 10.6151
R18081 gnd.n3253 gnd.n3246 10.6151
R18082 gnd.n3634 gnd.n2870 10.6151
R18083 gnd.n3634 gnd.n3633 10.6151
R18084 gnd.n3631 gnd.n2876 10.6151
R18085 gnd.n3625 gnd.n2876 10.6151
R18086 gnd.n3625 gnd.n3624 10.6151
R18087 gnd.n3624 gnd.n3623 10.6151
R18088 gnd.n3623 gnd.n2878 10.6151
R18089 gnd.n3617 gnd.n2878 10.6151
R18090 gnd.n3617 gnd.n3616 10.6151
R18091 gnd.n3616 gnd.n3615 10.6151
R18092 gnd.n3615 gnd.n2880 10.6151
R18093 gnd.n3609 gnd.n2880 10.6151
R18094 gnd.n3609 gnd.n3608 10.6151
R18095 gnd.n3608 gnd.n3607 10.6151
R18096 gnd.n3607 gnd.n2882 10.6151
R18097 gnd.n3601 gnd.n2882 10.6151
R18098 gnd.n3601 gnd.n3600 10.6151
R18099 gnd.n3600 gnd.n3599 10.6151
R18100 gnd.n3599 gnd.n2884 10.6151
R18101 gnd.n3593 gnd.n2884 10.6151
R18102 gnd.n3593 gnd.n3592 10.6151
R18103 gnd.n3592 gnd.n3591 10.6151
R18104 gnd.n3591 gnd.n2886 10.6151
R18105 gnd.n3585 gnd.n2886 10.6151
R18106 gnd.n3585 gnd.n3584 10.6151
R18107 gnd.n3584 gnd.n3583 10.6151
R18108 gnd.n3583 gnd.n2888 10.6151
R18109 gnd.n3577 gnd.n2888 10.6151
R18110 gnd.n3577 gnd.n3576 10.6151
R18111 gnd.n3576 gnd.n3575 10.6151
R18112 gnd.n2995 gnd.n2994 10.6151
R18113 gnd.n2994 gnd.n2915 10.6151
R18114 gnd.n2989 gnd.n2915 10.6151
R18115 gnd.n2989 gnd.n2988 10.6151
R18116 gnd.n2988 gnd.n2917 10.6151
R18117 gnd.n2983 gnd.n2917 10.6151
R18118 gnd.n2983 gnd.n2982 10.6151
R18119 gnd.n2982 gnd.n2981 10.6151
R18120 gnd.n2981 gnd.n2919 10.6151
R18121 gnd.n2975 gnd.n2919 10.6151
R18122 gnd.n2975 gnd.n2974 10.6151
R18123 gnd.n2974 gnd.n2973 10.6151
R18124 gnd.n2973 gnd.n2921 10.6151
R18125 gnd.n2967 gnd.n2921 10.6151
R18126 gnd.n2967 gnd.n2966 10.6151
R18127 gnd.n2966 gnd.n2965 10.6151
R18128 gnd.n2965 gnd.n2923 10.6151
R18129 gnd.n2959 gnd.n2923 10.6151
R18130 gnd.n2959 gnd.n2958 10.6151
R18131 gnd.n2958 gnd.n2957 10.6151
R18132 gnd.n2957 gnd.n2925 10.6151
R18133 gnd.n2951 gnd.n2925 10.6151
R18134 gnd.n2951 gnd.n2950 10.6151
R18135 gnd.n2950 gnd.n2949 10.6151
R18136 gnd.n2949 gnd.n2927 10.6151
R18137 gnd.n2943 gnd.n2927 10.6151
R18138 gnd.n2943 gnd.n2942 10.6151
R18139 gnd.n2942 gnd.n2941 10.6151
R18140 gnd.n2937 gnd.n2936 10.6151
R18141 gnd.n2936 gnd.n2871 10.6151
R18142 gnd.n3376 gnd.n3195 10.6151
R18143 gnd.n3197 gnd.n3195 10.6151
R18144 gnd.n3369 gnd.n3197 10.6151
R18145 gnd.n3369 gnd.n3368 10.6151
R18146 gnd.n3368 gnd.n3367 10.6151
R18147 gnd.n3367 gnd.n3199 10.6151
R18148 gnd.n3362 gnd.n3199 10.6151
R18149 gnd.n3362 gnd.n3361 10.6151
R18150 gnd.n3361 gnd.n3360 10.6151
R18151 gnd.n3360 gnd.n3202 10.6151
R18152 gnd.n3355 gnd.n3202 10.6151
R18153 gnd.n3355 gnd.n3354 10.6151
R18154 gnd.n3354 gnd.n3353 10.6151
R18155 gnd.n3353 gnd.n3205 10.6151
R18156 gnd.n3348 gnd.n3205 10.6151
R18157 gnd.n3348 gnd.n3347 10.6151
R18158 gnd.n3347 gnd.n3346 10.6151
R18159 gnd.n3346 gnd.n3208 10.6151
R18160 gnd.n3341 gnd.n3208 10.6151
R18161 gnd.n3341 gnd.n3340 10.6151
R18162 gnd.n3340 gnd.n3339 10.6151
R18163 gnd.n3339 gnd.n3211 10.6151
R18164 gnd.n3334 gnd.n3211 10.6151
R18165 gnd.n3334 gnd.n3333 10.6151
R18166 gnd.n3333 gnd.n3332 10.6151
R18167 gnd.n3332 gnd.n3214 10.6151
R18168 gnd.n3327 gnd.n3214 10.6151
R18169 gnd.n3327 gnd.n3326 10.6151
R18170 gnd.n3324 gnd.n3219 10.6151
R18171 gnd.n3319 gnd.n3219 10.6151
R18172 gnd.n3569 gnd.n3568 10.6151
R18173 gnd.n3568 gnd.n3567 10.6151
R18174 gnd.n3567 gnd.n2997 10.6151
R18175 gnd.n3557 gnd.n2997 10.6151
R18176 gnd.n3557 gnd.n3556 10.6151
R18177 gnd.n3556 gnd.n3555 10.6151
R18178 gnd.n3555 gnd.n3007 10.6151
R18179 gnd.n3018 gnd.n3007 10.6151
R18180 gnd.n3019 gnd.n3018 10.6151
R18181 gnd.n3543 gnd.n3019 10.6151
R18182 gnd.n3543 gnd.n3542 10.6151
R18183 gnd.n3542 gnd.n3541 10.6151
R18184 gnd.n3541 gnd.n3020 10.6151
R18185 gnd.n3032 gnd.n3020 10.6151
R18186 gnd.n3033 gnd.n3032 10.6151
R18187 gnd.n3529 gnd.n3033 10.6151
R18188 gnd.n3529 gnd.n3528 10.6151
R18189 gnd.n3528 gnd.n3527 10.6151
R18190 gnd.n3527 gnd.n3034 10.6151
R18191 gnd.n3520 gnd.n3034 10.6151
R18192 gnd.n3520 gnd.n3519 10.6151
R18193 gnd.n3519 gnd.n3518 10.6151
R18194 gnd.n3518 gnd.n3040 10.6151
R18195 gnd.n3057 gnd.n3040 10.6151
R18196 gnd.n3507 gnd.n3057 10.6151
R18197 gnd.n3507 gnd.n3506 10.6151
R18198 gnd.n3506 gnd.n3505 10.6151
R18199 gnd.n3505 gnd.n3058 10.6151
R18200 gnd.n3501 gnd.n3058 10.6151
R18201 gnd.n3501 gnd.n3500 10.6151
R18202 gnd.n3500 gnd.n3499 10.6151
R18203 gnd.n3499 gnd.n3060 10.6151
R18204 gnd.n3062 gnd.n3060 10.6151
R18205 gnd.n3086 gnd.n3062 10.6151
R18206 gnd.n3087 gnd.n3086 10.6151
R18207 gnd.n3485 gnd.n3087 10.6151
R18208 gnd.n3485 gnd.n3484 10.6151
R18209 gnd.n3484 gnd.n3483 10.6151
R18210 gnd.n3483 gnd.n3088 10.6151
R18211 gnd.n3099 gnd.n3088 10.6151
R18212 gnd.n3100 gnd.n3099 10.6151
R18213 gnd.n3470 gnd.n3100 10.6151
R18214 gnd.n3470 gnd.n3469 10.6151
R18215 gnd.n3469 gnd.n3468 10.6151
R18216 gnd.n3468 gnd.n3101 10.6151
R18217 gnd.n3112 gnd.n3101 10.6151
R18218 gnd.n3113 gnd.n3112 10.6151
R18219 gnd.n3455 gnd.n3113 10.6151
R18220 gnd.n3455 gnd.n3454 10.6151
R18221 gnd.n3454 gnd.n3453 10.6151
R18222 gnd.n3453 gnd.n3114 10.6151
R18223 gnd.n3124 gnd.n3114 10.6151
R18224 gnd.n3441 gnd.n3124 10.6151
R18225 gnd.n3441 gnd.n3440 10.6151
R18226 gnd.n3440 gnd.n3439 10.6151
R18227 gnd.n3439 gnd.n3125 10.6151
R18228 gnd.n3429 gnd.n3125 10.6151
R18229 gnd.n3429 gnd.n3428 10.6151
R18230 gnd.n3428 gnd.n3427 10.6151
R18231 gnd.n3427 gnd.n3133 10.6151
R18232 gnd.n3144 gnd.n3133 10.6151
R18233 gnd.n3145 gnd.n3144 10.6151
R18234 gnd.n3415 gnd.n3145 10.6151
R18235 gnd.n3415 gnd.n3414 10.6151
R18236 gnd.n3414 gnd.n3413 10.6151
R18237 gnd.n3413 gnd.n3146 10.6151
R18238 gnd.n3158 gnd.n3146 10.6151
R18239 gnd.n3401 gnd.n3158 10.6151
R18240 gnd.n3401 gnd.n3400 10.6151
R18241 gnd.n3400 gnd.n3399 10.6151
R18242 gnd.n3399 gnd.n3159 10.6151
R18243 gnd.n3170 gnd.n3159 10.6151
R18244 gnd.n3172 gnd.n3170 10.6151
R18245 gnd.n3173 gnd.n3172 10.6151
R18246 gnd.n3385 gnd.n3173 10.6151
R18247 gnd.n3385 gnd.n3384 10.6151
R18248 gnd.n3384 gnd.n3383 10.6151
R18249 gnd.n3383 gnd.n3174 10.6151
R18250 gnd.n3379 gnd.n3174 10.6151
R18251 gnd.n3379 gnd.n3378 10.6151
R18252 gnd.n5498 gnd.t26 10.5161
R18253 gnd.n4935 gnd.t36 10.5161
R18254 gnd.n6136 gnd.t318 10.5161
R18255 gnd.n6073 gnd.n6057 10.4732
R18256 gnd.n6041 gnd.n6025 10.4732
R18257 gnd.n6009 gnd.n5993 10.4732
R18258 gnd.n5978 gnd.n5962 10.4732
R18259 gnd.n5946 gnd.n5930 10.4732
R18260 gnd.n5914 gnd.n5898 10.4732
R18261 gnd.n5882 gnd.n5866 10.4732
R18262 gnd.n5851 gnd.n5835 10.4732
R18263 gnd.t51 gnd.n3515 10.1975
R18264 gnd.n3431 gnd.t305 10.1975
R18265 gnd.n5805 gnd.t320 9.87883
R18266 gnd.n7504 gnd.n66 9.73455
R18267 gnd.n6077 gnd.n6076 9.69747
R18268 gnd.n6045 gnd.n6044 9.69747
R18269 gnd.n6013 gnd.n6012 9.69747
R18270 gnd.n5982 gnd.n5981 9.69747
R18271 gnd.n5950 gnd.n5949 9.69747
R18272 gnd.n5918 gnd.n5917 9.69747
R18273 gnd.n5886 gnd.n5885 9.69747
R18274 gnd.n5855 gnd.n5854 9.69747
R18275 gnd.n3833 gnd.n2073 9.56018
R18276 gnd.n3865 gnd.t8 9.56018
R18277 gnd.n3074 gnd.n3073 9.56018
R18278 gnd.n3953 gnd.n1967 9.56018
R18279 gnd.n3141 gnd.t324 9.56018
R18280 gnd.n3387 gnd.t156 9.56018
R18281 gnd.t77 gnd.n1897 9.56018
R18282 gnd.n3256 gnd.n3255 9.56018
R18283 gnd.n4590 gnd.n1276 9.45751
R18284 gnd.n1722 gnd.n1503 9.45599
R18285 gnd.n6083 gnd.n6082 9.45567
R18286 gnd.n6051 gnd.n6050 9.45567
R18287 gnd.n6019 gnd.n6018 9.45567
R18288 gnd.n5988 gnd.n5987 9.45567
R18289 gnd.n5956 gnd.n5955 9.45567
R18290 gnd.n5924 gnd.n5923 9.45567
R18291 gnd.n5892 gnd.n5891 9.45567
R18292 gnd.n5861 gnd.n5860 9.45567
R18293 gnd.n5461 gnd.n5460 9.39724
R18294 gnd.n6082 gnd.n6081 9.3005
R18295 gnd.n6055 gnd.n6054 9.3005
R18296 gnd.n6076 gnd.n6075 9.3005
R18297 gnd.n6074 gnd.n6073 9.3005
R18298 gnd.n6059 gnd.n6058 9.3005
R18299 gnd.n6068 gnd.n6067 9.3005
R18300 gnd.n6066 gnd.n6065 9.3005
R18301 gnd.n6050 gnd.n6049 9.3005
R18302 gnd.n6023 gnd.n6022 9.3005
R18303 gnd.n6044 gnd.n6043 9.3005
R18304 gnd.n6042 gnd.n6041 9.3005
R18305 gnd.n6027 gnd.n6026 9.3005
R18306 gnd.n6036 gnd.n6035 9.3005
R18307 gnd.n6034 gnd.n6033 9.3005
R18308 gnd.n6018 gnd.n6017 9.3005
R18309 gnd.n5991 gnd.n5990 9.3005
R18310 gnd.n6012 gnd.n6011 9.3005
R18311 gnd.n6010 gnd.n6009 9.3005
R18312 gnd.n5995 gnd.n5994 9.3005
R18313 gnd.n6004 gnd.n6003 9.3005
R18314 gnd.n6002 gnd.n6001 9.3005
R18315 gnd.n5987 gnd.n5986 9.3005
R18316 gnd.n5960 gnd.n5959 9.3005
R18317 gnd.n5981 gnd.n5980 9.3005
R18318 gnd.n5979 gnd.n5978 9.3005
R18319 gnd.n5964 gnd.n5963 9.3005
R18320 gnd.n5973 gnd.n5972 9.3005
R18321 gnd.n5971 gnd.n5970 9.3005
R18322 gnd.n5955 gnd.n5954 9.3005
R18323 gnd.n5928 gnd.n5927 9.3005
R18324 gnd.n5949 gnd.n5948 9.3005
R18325 gnd.n5947 gnd.n5946 9.3005
R18326 gnd.n5932 gnd.n5931 9.3005
R18327 gnd.n5941 gnd.n5940 9.3005
R18328 gnd.n5939 gnd.n5938 9.3005
R18329 gnd.n5923 gnd.n5922 9.3005
R18330 gnd.n5896 gnd.n5895 9.3005
R18331 gnd.n5917 gnd.n5916 9.3005
R18332 gnd.n5915 gnd.n5914 9.3005
R18333 gnd.n5900 gnd.n5899 9.3005
R18334 gnd.n5909 gnd.n5908 9.3005
R18335 gnd.n5907 gnd.n5906 9.3005
R18336 gnd.n5891 gnd.n5890 9.3005
R18337 gnd.n5864 gnd.n5863 9.3005
R18338 gnd.n5885 gnd.n5884 9.3005
R18339 gnd.n5883 gnd.n5882 9.3005
R18340 gnd.n5868 gnd.n5867 9.3005
R18341 gnd.n5877 gnd.n5876 9.3005
R18342 gnd.n5875 gnd.n5874 9.3005
R18343 gnd.n5860 gnd.n5859 9.3005
R18344 gnd.n5833 gnd.n5832 9.3005
R18345 gnd.n5854 gnd.n5853 9.3005
R18346 gnd.n5852 gnd.n5851 9.3005
R18347 gnd.n5837 gnd.n5836 9.3005
R18348 gnd.n5846 gnd.n5845 9.3005
R18349 gnd.n5844 gnd.n5843 9.3005
R18350 gnd.n6230 gnd.n4839 9.3005
R18351 gnd.n6229 gnd.n4841 9.3005
R18352 gnd.n4845 gnd.n4842 9.3005
R18353 gnd.n6224 gnd.n4846 9.3005
R18354 gnd.n6223 gnd.n4847 9.3005
R18355 gnd.n6222 gnd.n4848 9.3005
R18356 gnd.n4852 gnd.n4849 9.3005
R18357 gnd.n6217 gnd.n4853 9.3005
R18358 gnd.n6216 gnd.n4854 9.3005
R18359 gnd.n6215 gnd.n4855 9.3005
R18360 gnd.n4859 gnd.n4856 9.3005
R18361 gnd.n6210 gnd.n4860 9.3005
R18362 gnd.n6209 gnd.n4861 9.3005
R18363 gnd.n6208 gnd.n4862 9.3005
R18364 gnd.n4867 gnd.n4865 9.3005
R18365 gnd.n6203 gnd.n6202 9.3005
R18366 gnd.n6232 gnd.n6231 9.3005
R18367 gnd.n5517 gnd.n5516 9.3005
R18368 gnd.n5135 gnd.n5134 9.3005
R18369 gnd.n5544 gnd.n5543 9.3005
R18370 gnd.n5545 gnd.n5133 9.3005
R18371 gnd.n5549 gnd.n5546 9.3005
R18372 gnd.n5548 gnd.n5547 9.3005
R18373 gnd.n5109 gnd.n5108 9.3005
R18374 gnd.n5575 gnd.n5574 9.3005
R18375 gnd.n5576 gnd.n5107 9.3005
R18376 gnd.n5580 gnd.n5577 9.3005
R18377 gnd.n5579 gnd.n5578 9.3005
R18378 gnd.n5084 gnd.n5083 9.3005
R18379 gnd.n5606 gnd.n5605 9.3005
R18380 gnd.n5607 gnd.n5082 9.3005
R18381 gnd.n5611 gnd.n5608 9.3005
R18382 gnd.n5610 gnd.n5609 9.3005
R18383 gnd.n5058 gnd.n5057 9.3005
R18384 gnd.n5637 gnd.n5636 9.3005
R18385 gnd.n5638 gnd.n5056 9.3005
R18386 gnd.n5642 gnd.n5639 9.3005
R18387 gnd.n5641 gnd.n5640 9.3005
R18388 gnd.n5034 gnd.n5033 9.3005
R18389 gnd.n5667 gnd.n5666 9.3005
R18390 gnd.n5668 gnd.n5032 9.3005
R18391 gnd.n5672 gnd.n5669 9.3005
R18392 gnd.n5671 gnd.n5670 9.3005
R18393 gnd.n5003 gnd.n5002 9.3005
R18394 gnd.n5721 gnd.n5720 9.3005
R18395 gnd.n5722 gnd.n5001 9.3005
R18396 gnd.n5724 gnd.n5723 9.3005
R18397 gnd.n4982 gnd.n4981 9.3005
R18398 gnd.n5751 gnd.n5750 9.3005
R18399 gnd.n5752 gnd.n4980 9.3005
R18400 gnd.n5756 gnd.n5753 9.3005
R18401 gnd.n5755 gnd.n5754 9.3005
R18402 gnd.n4958 gnd.n4957 9.3005
R18403 gnd.n5797 gnd.n5796 9.3005
R18404 gnd.n5798 gnd.n4956 9.3005
R18405 gnd.n5802 gnd.n5799 9.3005
R18406 gnd.n5801 gnd.n5800 9.3005
R18407 gnd.n4928 gnd.n4927 9.3005
R18408 gnd.n6118 gnd.n6117 9.3005
R18409 gnd.n6119 gnd.n4926 9.3005
R18410 gnd.n6127 gnd.n6120 9.3005
R18411 gnd.n6126 gnd.n6121 9.3005
R18412 gnd.n6125 gnd.n6123 9.3005
R18413 gnd.n6122 gnd.n913 9.3005
R18414 gnd.n6248 gnd.n914 9.3005
R18415 gnd.n6247 gnd.n915 9.3005
R18416 gnd.n6246 gnd.n916 9.3005
R18417 gnd.n4837 gnd.n917 9.3005
R18418 gnd.n4838 gnd.n4836 9.3005
R18419 gnd.n6234 gnd.n6233 9.3005
R18420 gnd.n5518 gnd.n5515 9.3005
R18421 gnd.n5214 gnd.n5173 9.3005
R18422 gnd.n5209 gnd.n5208 9.3005
R18423 gnd.n5207 gnd.n5174 9.3005
R18424 gnd.n5206 gnd.n5205 9.3005
R18425 gnd.n5202 gnd.n5175 9.3005
R18426 gnd.n5199 gnd.n5198 9.3005
R18427 gnd.n5197 gnd.n5176 9.3005
R18428 gnd.n5196 gnd.n5195 9.3005
R18429 gnd.n5192 gnd.n5177 9.3005
R18430 gnd.n5189 gnd.n5188 9.3005
R18431 gnd.n5187 gnd.n5178 9.3005
R18432 gnd.n5186 gnd.n5185 9.3005
R18433 gnd.n5182 gnd.n5180 9.3005
R18434 gnd.n5179 gnd.n5159 9.3005
R18435 gnd.n5512 gnd.n5158 9.3005
R18436 gnd.n5514 gnd.n5513 9.3005
R18437 gnd.n5216 gnd.n5215 9.3005
R18438 gnd.n5525 gnd.n5145 9.3005
R18439 gnd.n5532 gnd.n5146 9.3005
R18440 gnd.n5534 gnd.n5533 9.3005
R18441 gnd.n5535 gnd.n5126 9.3005
R18442 gnd.n5554 gnd.n5553 9.3005
R18443 gnd.n5556 gnd.n5119 9.3005
R18444 gnd.n5563 gnd.n5120 9.3005
R18445 gnd.n5565 gnd.n5564 9.3005
R18446 gnd.n5566 gnd.n5102 9.3005
R18447 gnd.n5585 gnd.n5584 9.3005
R18448 gnd.n5587 gnd.n5094 9.3005
R18449 gnd.n5594 gnd.n5095 9.3005
R18450 gnd.n5596 gnd.n5595 9.3005
R18451 gnd.n5597 gnd.n5076 9.3005
R18452 gnd.n5616 gnd.n5615 9.3005
R18453 gnd.n5618 gnd.n5068 9.3005
R18454 gnd.n5625 gnd.n5069 9.3005
R18455 gnd.n5627 gnd.n5626 9.3005
R18456 gnd.n5628 gnd.n5051 9.3005
R18457 gnd.n5647 gnd.n5646 9.3005
R18458 gnd.n5649 gnd.n5043 9.3005
R18459 gnd.n5656 gnd.n5044 9.3005
R18460 gnd.n5658 gnd.n5657 9.3005
R18461 gnd.n5659 gnd.n5027 9.3005
R18462 gnd.n5677 gnd.n5676 9.3005
R18463 gnd.n5679 gnd.n5012 9.3005
R18464 gnd.n5710 gnd.n5014 9.3005
R18465 gnd.n5711 gnd.n5010 9.3005
R18466 gnd.n5713 gnd.n5712 9.3005
R18467 gnd.n4998 gnd.n4993 9.3005
R18468 gnd.n5734 gnd.n4992 9.3005
R18469 gnd.n5737 gnd.n5736 9.3005
R18470 gnd.n5739 gnd.n5738 9.3005
R18471 gnd.n5742 gnd.n4975 9.3005
R18472 gnd.n5740 gnd.n4973 9.3005
R18473 gnd.n5764 gnd.n4971 9.3005
R18474 gnd.n5766 gnd.n5765 9.3005
R18475 gnd.n4949 gnd.n4948 9.3005
R18476 gnd.n5811 gnd.n5810 9.3005
R18477 gnd.n5812 gnd.n4942 9.3005
R18478 gnd.n5820 gnd.n4941 9.3005
R18479 gnd.n5823 gnd.n5822 9.3005
R18480 gnd.n5825 gnd.n4939 9.3005
R18481 gnd.n6109 gnd.n6108 9.3005
R18482 gnd.n6107 gnd.n5826 9.3005
R18483 gnd.n5828 gnd.n5827 9.3005
R18484 gnd.n6103 gnd.n5829 9.3005
R18485 gnd.n6102 gnd.n5830 9.3005
R18486 gnd.n6101 gnd.n6088 9.3005
R18487 gnd.n6098 gnd.n6090 9.3005
R18488 gnd.n6097 gnd.n6091 9.3005
R18489 gnd.n6094 gnd.n6092 9.3005
R18490 gnd.n6093 gnd.n4868 9.3005
R18491 gnd.n5523 gnd.n5522 9.3005
R18492 gnd.n6198 gnd.n4869 9.3005
R18493 gnd.n6197 gnd.n4871 9.3005
R18494 gnd.n4875 gnd.n4872 9.3005
R18495 gnd.n6192 gnd.n4876 9.3005
R18496 gnd.n6191 gnd.n4877 9.3005
R18497 gnd.n6190 gnd.n4878 9.3005
R18498 gnd.n4882 gnd.n4879 9.3005
R18499 gnd.n6185 gnd.n4883 9.3005
R18500 gnd.n6184 gnd.n4884 9.3005
R18501 gnd.n6183 gnd.n4885 9.3005
R18502 gnd.n4889 gnd.n4886 9.3005
R18503 gnd.n6178 gnd.n4890 9.3005
R18504 gnd.n6177 gnd.n4891 9.3005
R18505 gnd.n6176 gnd.n4892 9.3005
R18506 gnd.n4896 gnd.n4893 9.3005
R18507 gnd.n6171 gnd.n4897 9.3005
R18508 gnd.n6170 gnd.n4898 9.3005
R18509 gnd.n6169 gnd.n4899 9.3005
R18510 gnd.n4903 gnd.n4900 9.3005
R18511 gnd.n6164 gnd.n4904 9.3005
R18512 gnd.n6163 gnd.n4905 9.3005
R18513 gnd.n6162 gnd.n4906 9.3005
R18514 gnd.n4913 gnd.n4911 9.3005
R18515 gnd.n6157 gnd.n4914 9.3005
R18516 gnd.n6156 gnd.n4915 9.3005
R18517 gnd.n6155 gnd.n6152 9.3005
R18518 gnd.n6200 gnd.n6199 9.3005
R18519 gnd.n5020 gnd.n5019 9.3005
R18520 gnd.n5687 gnd.n5686 9.3005
R18521 gnd.n5688 gnd.n5018 9.3005
R18522 gnd.n5705 gnd.n5689 9.3005
R18523 gnd.n5704 gnd.n5690 9.3005
R18524 gnd.n5703 gnd.n5691 9.3005
R18525 gnd.n5701 gnd.n5692 9.3005
R18526 gnd.n5700 gnd.n5693 9.3005
R18527 gnd.n5698 gnd.n5694 9.3005
R18528 gnd.n5697 gnd.n5695 9.3005
R18529 gnd.n4964 gnd.n4963 9.3005
R18530 gnd.n5774 gnd.n5773 9.3005
R18531 gnd.n5775 gnd.n4962 9.3005
R18532 gnd.n5789 gnd.n5776 9.3005
R18533 gnd.n5788 gnd.n5777 9.3005
R18534 gnd.n5787 gnd.n5778 9.3005
R18535 gnd.n5785 gnd.n5779 9.3005
R18536 gnd.n5784 gnd.n5780 9.3005
R18537 gnd.n5782 gnd.n5781 9.3005
R18538 gnd.n4921 gnd.n4920 9.3005
R18539 gnd.n6133 gnd.n6132 9.3005
R18540 gnd.n6134 gnd.n4919 9.3005
R18541 gnd.n6138 gnd.n6135 9.3005
R18542 gnd.n6139 gnd.n4918 9.3005
R18543 gnd.n6143 gnd.n6142 9.3005
R18544 gnd.n6144 gnd.n4917 9.3005
R18545 gnd.n6146 gnd.n6145 9.3005
R18546 gnd.n6149 gnd.n4916 9.3005
R18547 gnd.n6151 gnd.n6150 9.3005
R18548 gnd.n5347 gnd.n5346 9.3005
R18549 gnd.n5237 gnd.n5236 9.3005
R18550 gnd.n5361 gnd.n5360 9.3005
R18551 gnd.n5362 gnd.n5235 9.3005
R18552 gnd.n5364 gnd.n5363 9.3005
R18553 gnd.n5225 gnd.n5224 9.3005
R18554 gnd.n5377 gnd.n5376 9.3005
R18555 gnd.n5378 gnd.n5223 9.3005
R18556 gnd.n5496 gnd.n5379 9.3005
R18557 gnd.n5495 gnd.n5380 9.3005
R18558 gnd.n5494 gnd.n5381 9.3005
R18559 gnd.n5493 gnd.n5382 9.3005
R18560 gnd.n5490 gnd.n5383 9.3005
R18561 gnd.n5489 gnd.n5384 9.3005
R18562 gnd.n5488 gnd.n5385 9.3005
R18563 gnd.n5486 gnd.n5386 9.3005
R18564 gnd.n5485 gnd.n5387 9.3005
R18565 gnd.n5482 gnd.n5388 9.3005
R18566 gnd.n5481 gnd.n5389 9.3005
R18567 gnd.n5480 gnd.n5390 9.3005
R18568 gnd.n5478 gnd.n5391 9.3005
R18569 gnd.n5477 gnd.n5392 9.3005
R18570 gnd.n5473 gnd.n5393 9.3005
R18571 gnd.n5472 gnd.n5394 9.3005
R18572 gnd.n5471 gnd.n5395 9.3005
R18573 gnd.n5469 gnd.n5396 9.3005
R18574 gnd.n5468 gnd.n5397 9.3005
R18575 gnd.n5465 gnd.n5398 9.3005
R18576 gnd.n5345 gnd.n5246 9.3005
R18577 gnd.n5248 gnd.n5247 9.3005
R18578 gnd.n5292 gnd.n5290 9.3005
R18579 gnd.n5293 gnd.n5289 9.3005
R18580 gnd.n5296 gnd.n5285 9.3005
R18581 gnd.n5297 gnd.n5284 9.3005
R18582 gnd.n5300 gnd.n5283 9.3005
R18583 gnd.n5301 gnd.n5282 9.3005
R18584 gnd.n5304 gnd.n5281 9.3005
R18585 gnd.n5305 gnd.n5280 9.3005
R18586 gnd.n5308 gnd.n5279 9.3005
R18587 gnd.n5309 gnd.n5278 9.3005
R18588 gnd.n5312 gnd.n5277 9.3005
R18589 gnd.n5313 gnd.n5276 9.3005
R18590 gnd.n5316 gnd.n5275 9.3005
R18591 gnd.n5317 gnd.n5274 9.3005
R18592 gnd.n5320 gnd.n5273 9.3005
R18593 gnd.n5321 gnd.n5272 9.3005
R18594 gnd.n5324 gnd.n5271 9.3005
R18595 gnd.n5325 gnd.n5270 9.3005
R18596 gnd.n5328 gnd.n5269 9.3005
R18597 gnd.n5329 gnd.n5268 9.3005
R18598 gnd.n5332 gnd.n5267 9.3005
R18599 gnd.n5334 gnd.n5266 9.3005
R18600 gnd.n5335 gnd.n5265 9.3005
R18601 gnd.n5336 gnd.n5264 9.3005
R18602 gnd.n5337 gnd.n5263 9.3005
R18603 gnd.n5344 gnd.n5343 9.3005
R18604 gnd.n5353 gnd.n5352 9.3005
R18605 gnd.n5354 gnd.n5240 9.3005
R18606 gnd.n5356 gnd.n5355 9.3005
R18607 gnd.n5231 gnd.n5230 9.3005
R18608 gnd.n5369 gnd.n5368 9.3005
R18609 gnd.n5370 gnd.n5229 9.3005
R18610 gnd.n5372 gnd.n5371 9.3005
R18611 gnd.n5218 gnd.n5217 9.3005
R18612 gnd.n5501 gnd.n5500 9.3005
R18613 gnd.n5502 gnd.n5172 9.3005
R18614 gnd.n5506 gnd.n5504 9.3005
R18615 gnd.n5505 gnd.n5151 9.3005
R18616 gnd.n5524 gnd.n5150 9.3005
R18617 gnd.n5527 gnd.n5526 9.3005
R18618 gnd.n5144 gnd.n5143 9.3005
R18619 gnd.n5538 gnd.n5536 9.3005
R18620 gnd.n5537 gnd.n5125 9.3005
R18621 gnd.n5555 gnd.n5124 9.3005
R18622 gnd.n5558 gnd.n5557 9.3005
R18623 gnd.n5118 gnd.n5117 9.3005
R18624 gnd.n5569 gnd.n5567 9.3005
R18625 gnd.n5568 gnd.n5101 9.3005
R18626 gnd.n5586 gnd.n5100 9.3005
R18627 gnd.n5589 gnd.n5588 9.3005
R18628 gnd.n5093 gnd.n5092 9.3005
R18629 gnd.n5600 gnd.n5598 9.3005
R18630 gnd.n5599 gnd.n5075 9.3005
R18631 gnd.n5617 gnd.n5074 9.3005
R18632 gnd.n5620 gnd.n5619 9.3005
R18633 gnd.n5067 gnd.n5066 9.3005
R18634 gnd.n5631 gnd.n5629 9.3005
R18635 gnd.n5630 gnd.n5050 9.3005
R18636 gnd.n5648 gnd.n5049 9.3005
R18637 gnd.n5651 gnd.n5650 9.3005
R18638 gnd.n5042 gnd.n5041 9.3005
R18639 gnd.n5661 gnd.n5660 9.3005
R18640 gnd.n5026 gnd.n5025 9.3005
R18641 gnd.n5682 gnd.n5678 9.3005
R18642 gnd.n5681 gnd.n5680 9.3005
R18643 gnd.n5013 gnd.n5009 9.3005
R18644 gnd.n5715 gnd.n5714 9.3005
R18645 gnd.n5011 gnd.n4994 9.3005
R18646 gnd.n5733 gnd.n5732 9.3005
R18647 gnd.n5735 gnd.n4990 9.3005
R18648 gnd.n5745 gnd.n4991 9.3005
R18649 gnd.n5744 gnd.n5743 9.3005
R18650 gnd.n5741 gnd.n4969 9.3005
R18651 gnd.n5769 gnd.n4970 9.3005
R18652 gnd.n5768 gnd.n5767 9.3005
R18653 gnd.n4972 gnd.n4950 9.3005
R18654 gnd.n5808 gnd.n5807 9.3005
R18655 gnd.n5809 gnd.n4943 9.3005
R18656 gnd.n5819 gnd.n5818 9.3005
R18657 gnd.n5821 gnd.n4937 9.3005
R18658 gnd.n6112 gnd.n4938 9.3005
R18659 gnd.n6111 gnd.n6110 9.3005
R18660 gnd.n4940 gnd.n901 9.3005
R18661 gnd.n6255 gnd.n902 9.3005
R18662 gnd.n6254 gnd.n903 9.3005
R18663 gnd.n6253 gnd.n904 9.3005
R18664 gnd.n6087 gnd.n905 9.3005
R18665 gnd.n6089 gnd.n925 9.3005
R18666 gnd.n6241 gnd.n926 9.3005
R18667 gnd.n6240 gnd.n927 9.3005
R18668 gnd.n6239 gnd.n928 9.3005
R18669 gnd.n5242 gnd.n5241 9.3005
R18670 gnd.n6430 gnd.n6429 9.3005
R18671 gnd.n6431 gnd.n725 9.3005
R18672 gnd.n6433 gnd.n6432 9.3005
R18673 gnd.n721 gnd.n720 9.3005
R18674 gnd.n6440 gnd.n6439 9.3005
R18675 gnd.n6441 gnd.n719 9.3005
R18676 gnd.n6443 gnd.n6442 9.3005
R18677 gnd.n715 gnd.n714 9.3005
R18678 gnd.n6450 gnd.n6449 9.3005
R18679 gnd.n6451 gnd.n713 9.3005
R18680 gnd.n6453 gnd.n6452 9.3005
R18681 gnd.n709 gnd.n708 9.3005
R18682 gnd.n6460 gnd.n6459 9.3005
R18683 gnd.n6461 gnd.n707 9.3005
R18684 gnd.n6463 gnd.n6462 9.3005
R18685 gnd.n703 gnd.n702 9.3005
R18686 gnd.n6470 gnd.n6469 9.3005
R18687 gnd.n6471 gnd.n701 9.3005
R18688 gnd.n6473 gnd.n6472 9.3005
R18689 gnd.n697 gnd.n696 9.3005
R18690 gnd.n6480 gnd.n6479 9.3005
R18691 gnd.n6481 gnd.n695 9.3005
R18692 gnd.n6483 gnd.n6482 9.3005
R18693 gnd.n691 gnd.n690 9.3005
R18694 gnd.n6490 gnd.n6489 9.3005
R18695 gnd.n6491 gnd.n689 9.3005
R18696 gnd.n6493 gnd.n6492 9.3005
R18697 gnd.n685 gnd.n684 9.3005
R18698 gnd.n6500 gnd.n6499 9.3005
R18699 gnd.n6501 gnd.n683 9.3005
R18700 gnd.n6503 gnd.n6502 9.3005
R18701 gnd.n679 gnd.n678 9.3005
R18702 gnd.n6510 gnd.n6509 9.3005
R18703 gnd.n6511 gnd.n677 9.3005
R18704 gnd.n6513 gnd.n6512 9.3005
R18705 gnd.n673 gnd.n672 9.3005
R18706 gnd.n6520 gnd.n6519 9.3005
R18707 gnd.n6521 gnd.n671 9.3005
R18708 gnd.n6523 gnd.n6522 9.3005
R18709 gnd.n667 gnd.n666 9.3005
R18710 gnd.n6530 gnd.n6529 9.3005
R18711 gnd.n6531 gnd.n665 9.3005
R18712 gnd.n6533 gnd.n6532 9.3005
R18713 gnd.n661 gnd.n660 9.3005
R18714 gnd.n6540 gnd.n6539 9.3005
R18715 gnd.n6541 gnd.n659 9.3005
R18716 gnd.n6543 gnd.n6542 9.3005
R18717 gnd.n655 gnd.n654 9.3005
R18718 gnd.n6550 gnd.n6549 9.3005
R18719 gnd.n6551 gnd.n653 9.3005
R18720 gnd.n6553 gnd.n6552 9.3005
R18721 gnd.n649 gnd.n648 9.3005
R18722 gnd.n6560 gnd.n6559 9.3005
R18723 gnd.n6561 gnd.n647 9.3005
R18724 gnd.n6563 gnd.n6562 9.3005
R18725 gnd.n643 gnd.n642 9.3005
R18726 gnd.n6570 gnd.n6569 9.3005
R18727 gnd.n6571 gnd.n641 9.3005
R18728 gnd.n6573 gnd.n6572 9.3005
R18729 gnd.n637 gnd.n636 9.3005
R18730 gnd.n6580 gnd.n6579 9.3005
R18731 gnd.n6581 gnd.n635 9.3005
R18732 gnd.n6583 gnd.n6582 9.3005
R18733 gnd.n631 gnd.n630 9.3005
R18734 gnd.n6590 gnd.n6589 9.3005
R18735 gnd.n6591 gnd.n629 9.3005
R18736 gnd.n6593 gnd.n6592 9.3005
R18737 gnd.n625 gnd.n624 9.3005
R18738 gnd.n6600 gnd.n6599 9.3005
R18739 gnd.n6601 gnd.n623 9.3005
R18740 gnd.n6603 gnd.n6602 9.3005
R18741 gnd.n619 gnd.n618 9.3005
R18742 gnd.n6610 gnd.n6609 9.3005
R18743 gnd.n6611 gnd.n617 9.3005
R18744 gnd.n6613 gnd.n6612 9.3005
R18745 gnd.n613 gnd.n612 9.3005
R18746 gnd.n6620 gnd.n6619 9.3005
R18747 gnd.n6621 gnd.n611 9.3005
R18748 gnd.n6623 gnd.n6622 9.3005
R18749 gnd.n607 gnd.n606 9.3005
R18750 gnd.n6630 gnd.n6629 9.3005
R18751 gnd.n6631 gnd.n605 9.3005
R18752 gnd.n6633 gnd.n6632 9.3005
R18753 gnd.n601 gnd.n600 9.3005
R18754 gnd.n6640 gnd.n6639 9.3005
R18755 gnd.n6641 gnd.n599 9.3005
R18756 gnd.n6643 gnd.n6642 9.3005
R18757 gnd.n595 gnd.n594 9.3005
R18758 gnd.n6650 gnd.n6649 9.3005
R18759 gnd.n6651 gnd.n593 9.3005
R18760 gnd.n6653 gnd.n6652 9.3005
R18761 gnd.n589 gnd.n588 9.3005
R18762 gnd.n6660 gnd.n6659 9.3005
R18763 gnd.n6661 gnd.n587 9.3005
R18764 gnd.n6663 gnd.n6662 9.3005
R18765 gnd.n583 gnd.n582 9.3005
R18766 gnd.n6670 gnd.n6669 9.3005
R18767 gnd.n6671 gnd.n581 9.3005
R18768 gnd.n6673 gnd.n6672 9.3005
R18769 gnd.n577 gnd.n576 9.3005
R18770 gnd.n6680 gnd.n6679 9.3005
R18771 gnd.n6681 gnd.n575 9.3005
R18772 gnd.n6683 gnd.n6682 9.3005
R18773 gnd.n571 gnd.n570 9.3005
R18774 gnd.n6690 gnd.n6689 9.3005
R18775 gnd.n6691 gnd.n569 9.3005
R18776 gnd.n6693 gnd.n6692 9.3005
R18777 gnd.n565 gnd.n564 9.3005
R18778 gnd.n6700 gnd.n6699 9.3005
R18779 gnd.n6701 gnd.n563 9.3005
R18780 gnd.n6703 gnd.n6702 9.3005
R18781 gnd.n559 gnd.n558 9.3005
R18782 gnd.n6710 gnd.n6709 9.3005
R18783 gnd.n6711 gnd.n557 9.3005
R18784 gnd.n6713 gnd.n6712 9.3005
R18785 gnd.n553 gnd.n552 9.3005
R18786 gnd.n6720 gnd.n6719 9.3005
R18787 gnd.n6721 gnd.n551 9.3005
R18788 gnd.n6723 gnd.n6722 9.3005
R18789 gnd.n547 gnd.n546 9.3005
R18790 gnd.n6730 gnd.n6729 9.3005
R18791 gnd.n6731 gnd.n545 9.3005
R18792 gnd.n6733 gnd.n6732 9.3005
R18793 gnd.n541 gnd.n540 9.3005
R18794 gnd.n6740 gnd.n6739 9.3005
R18795 gnd.n6741 gnd.n539 9.3005
R18796 gnd.n6743 gnd.n6742 9.3005
R18797 gnd.n535 gnd.n534 9.3005
R18798 gnd.n6750 gnd.n6749 9.3005
R18799 gnd.n6751 gnd.n533 9.3005
R18800 gnd.n6753 gnd.n6752 9.3005
R18801 gnd.n529 gnd.n528 9.3005
R18802 gnd.n6760 gnd.n6759 9.3005
R18803 gnd.n6761 gnd.n527 9.3005
R18804 gnd.n6763 gnd.n6762 9.3005
R18805 gnd.n523 gnd.n522 9.3005
R18806 gnd.n6770 gnd.n6769 9.3005
R18807 gnd.n6771 gnd.n521 9.3005
R18808 gnd.n6773 gnd.n6772 9.3005
R18809 gnd.n517 gnd.n516 9.3005
R18810 gnd.n6780 gnd.n6779 9.3005
R18811 gnd.n6781 gnd.n515 9.3005
R18812 gnd.n6783 gnd.n6782 9.3005
R18813 gnd.n511 gnd.n510 9.3005
R18814 gnd.n6790 gnd.n6789 9.3005
R18815 gnd.n6791 gnd.n509 9.3005
R18816 gnd.n6793 gnd.n6792 9.3005
R18817 gnd.n505 gnd.n504 9.3005
R18818 gnd.n6800 gnd.n6799 9.3005
R18819 gnd.n6801 gnd.n503 9.3005
R18820 gnd.n6803 gnd.n6802 9.3005
R18821 gnd.n499 gnd.n498 9.3005
R18822 gnd.n6810 gnd.n6809 9.3005
R18823 gnd.n6811 gnd.n497 9.3005
R18824 gnd.n6813 gnd.n6812 9.3005
R18825 gnd.n493 gnd.n492 9.3005
R18826 gnd.n6820 gnd.n6819 9.3005
R18827 gnd.n6821 gnd.n491 9.3005
R18828 gnd.n6823 gnd.n6822 9.3005
R18829 gnd.n487 gnd.n486 9.3005
R18830 gnd.n6830 gnd.n6829 9.3005
R18831 gnd.n6831 gnd.n485 9.3005
R18832 gnd.n6833 gnd.n6832 9.3005
R18833 gnd.n481 gnd.n480 9.3005
R18834 gnd.n6840 gnd.n6839 9.3005
R18835 gnd.n6841 gnd.n479 9.3005
R18836 gnd.n6843 gnd.n6842 9.3005
R18837 gnd.n475 gnd.n474 9.3005
R18838 gnd.n6850 gnd.n6849 9.3005
R18839 gnd.n6851 gnd.n473 9.3005
R18840 gnd.n6853 gnd.n6852 9.3005
R18841 gnd.n469 gnd.n468 9.3005
R18842 gnd.n6860 gnd.n6859 9.3005
R18843 gnd.n6861 gnd.n467 9.3005
R18844 gnd.n6863 gnd.n6862 9.3005
R18845 gnd.n463 gnd.n462 9.3005
R18846 gnd.n6870 gnd.n6869 9.3005
R18847 gnd.n6871 gnd.n461 9.3005
R18848 gnd.n6874 gnd.n6873 9.3005
R18849 gnd.n6872 gnd.n457 9.3005
R18850 gnd.n6880 gnd.n456 9.3005
R18851 gnd.n6882 gnd.n6881 9.3005
R18852 gnd.n452 gnd.n451 9.3005
R18853 gnd.n6891 gnd.n6890 9.3005
R18854 gnd.n6892 gnd.n450 9.3005
R18855 gnd.n6894 gnd.n6893 9.3005
R18856 gnd.n446 gnd.n445 9.3005
R18857 gnd.n6901 gnd.n6900 9.3005
R18858 gnd.n6902 gnd.n444 9.3005
R18859 gnd.n6904 gnd.n6903 9.3005
R18860 gnd.n440 gnd.n439 9.3005
R18861 gnd.n6911 gnd.n6910 9.3005
R18862 gnd.n6912 gnd.n438 9.3005
R18863 gnd.n6914 gnd.n6913 9.3005
R18864 gnd.n434 gnd.n433 9.3005
R18865 gnd.n6921 gnd.n6920 9.3005
R18866 gnd.n6922 gnd.n432 9.3005
R18867 gnd.n6924 gnd.n6923 9.3005
R18868 gnd.n428 gnd.n427 9.3005
R18869 gnd.n6931 gnd.n6930 9.3005
R18870 gnd.n6932 gnd.n426 9.3005
R18871 gnd.n6934 gnd.n6933 9.3005
R18872 gnd.n422 gnd.n421 9.3005
R18873 gnd.n6941 gnd.n6940 9.3005
R18874 gnd.n6942 gnd.n420 9.3005
R18875 gnd.n6944 gnd.n6943 9.3005
R18876 gnd.n416 gnd.n415 9.3005
R18877 gnd.n6951 gnd.n6950 9.3005
R18878 gnd.n6952 gnd.n414 9.3005
R18879 gnd.n6954 gnd.n6953 9.3005
R18880 gnd.n410 gnd.n409 9.3005
R18881 gnd.n6961 gnd.n6960 9.3005
R18882 gnd.n6962 gnd.n408 9.3005
R18883 gnd.n6964 gnd.n6963 9.3005
R18884 gnd.n404 gnd.n403 9.3005
R18885 gnd.n6971 gnd.n6970 9.3005
R18886 gnd.n6972 gnd.n402 9.3005
R18887 gnd.n6974 gnd.n6973 9.3005
R18888 gnd.n398 gnd.n397 9.3005
R18889 gnd.n6981 gnd.n6980 9.3005
R18890 gnd.n6982 gnd.n396 9.3005
R18891 gnd.n6984 gnd.n6983 9.3005
R18892 gnd.n392 gnd.n391 9.3005
R18893 gnd.n6991 gnd.n6990 9.3005
R18894 gnd.n6992 gnd.n390 9.3005
R18895 gnd.n6994 gnd.n6993 9.3005
R18896 gnd.n386 gnd.n385 9.3005
R18897 gnd.n7001 gnd.n7000 9.3005
R18898 gnd.n7002 gnd.n384 9.3005
R18899 gnd.n7004 gnd.n7003 9.3005
R18900 gnd.n380 gnd.n379 9.3005
R18901 gnd.n7011 gnd.n7010 9.3005
R18902 gnd.n7012 gnd.n378 9.3005
R18903 gnd.n7014 gnd.n7013 9.3005
R18904 gnd.n374 gnd.n373 9.3005
R18905 gnd.n7021 gnd.n7020 9.3005
R18906 gnd.n7022 gnd.n372 9.3005
R18907 gnd.n7024 gnd.n7023 9.3005
R18908 gnd.n368 gnd.n367 9.3005
R18909 gnd.n7031 gnd.n7030 9.3005
R18910 gnd.n7032 gnd.n366 9.3005
R18911 gnd.n7034 gnd.n7033 9.3005
R18912 gnd.n362 gnd.n361 9.3005
R18913 gnd.n7041 gnd.n7040 9.3005
R18914 gnd.n7042 gnd.n360 9.3005
R18915 gnd.n7044 gnd.n7043 9.3005
R18916 gnd.n356 gnd.n355 9.3005
R18917 gnd.n7051 gnd.n7050 9.3005
R18918 gnd.n7052 gnd.n354 9.3005
R18919 gnd.n7054 gnd.n7053 9.3005
R18920 gnd.n350 gnd.n349 9.3005
R18921 gnd.n7061 gnd.n7060 9.3005
R18922 gnd.n7062 gnd.n348 9.3005
R18923 gnd.n7064 gnd.n7063 9.3005
R18924 gnd.n344 gnd.n343 9.3005
R18925 gnd.n7071 gnd.n7070 9.3005
R18926 gnd.n7072 gnd.n342 9.3005
R18927 gnd.n7074 gnd.n7073 9.3005
R18928 gnd.n338 gnd.n337 9.3005
R18929 gnd.n7081 gnd.n7080 9.3005
R18930 gnd.n7082 gnd.n336 9.3005
R18931 gnd.n7084 gnd.n7083 9.3005
R18932 gnd.n332 gnd.n331 9.3005
R18933 gnd.n7092 gnd.n7091 9.3005
R18934 gnd.n7093 gnd.n330 9.3005
R18935 gnd.n7096 gnd.n7095 9.3005
R18936 gnd.n6884 gnd.n6883 9.3005
R18937 gnd.n7455 gnd.n112 9.3005
R18938 gnd.n7454 gnd.n114 9.3005
R18939 gnd.n118 gnd.n115 9.3005
R18940 gnd.n7449 gnd.n119 9.3005
R18941 gnd.n7448 gnd.n120 9.3005
R18942 gnd.n7447 gnd.n121 9.3005
R18943 gnd.n125 gnd.n122 9.3005
R18944 gnd.n7442 gnd.n126 9.3005
R18945 gnd.n7441 gnd.n127 9.3005
R18946 gnd.n7440 gnd.n128 9.3005
R18947 gnd.n132 gnd.n129 9.3005
R18948 gnd.n7435 gnd.n133 9.3005
R18949 gnd.n7434 gnd.n134 9.3005
R18950 gnd.n7433 gnd.n135 9.3005
R18951 gnd.n139 gnd.n136 9.3005
R18952 gnd.n7428 gnd.n140 9.3005
R18953 gnd.n7427 gnd.n141 9.3005
R18954 gnd.n7423 gnd.n142 9.3005
R18955 gnd.n146 gnd.n143 9.3005
R18956 gnd.n7418 gnd.n147 9.3005
R18957 gnd.n7417 gnd.n148 9.3005
R18958 gnd.n7416 gnd.n149 9.3005
R18959 gnd.n153 gnd.n150 9.3005
R18960 gnd.n7411 gnd.n154 9.3005
R18961 gnd.n7410 gnd.n155 9.3005
R18962 gnd.n7409 gnd.n156 9.3005
R18963 gnd.n160 gnd.n157 9.3005
R18964 gnd.n7404 gnd.n161 9.3005
R18965 gnd.n7403 gnd.n162 9.3005
R18966 gnd.n7402 gnd.n163 9.3005
R18967 gnd.n167 gnd.n164 9.3005
R18968 gnd.n7397 gnd.n168 9.3005
R18969 gnd.n7396 gnd.n169 9.3005
R18970 gnd.n7395 gnd.n170 9.3005
R18971 gnd.n174 gnd.n171 9.3005
R18972 gnd.n7390 gnd.n175 9.3005
R18973 gnd.n7389 gnd.n7388 9.3005
R18974 gnd.n7387 gnd.n178 9.3005
R18975 gnd.n7457 gnd.n7456 9.3005
R18976 gnd.n1649 gnd.n1648 9.3005
R18977 gnd.n1678 gnd.n1650 9.3005
R18978 gnd.n1677 gnd.n1651 9.3005
R18979 gnd.n1676 gnd.n1652 9.3005
R18980 gnd.n1674 gnd.n1653 9.3005
R18981 gnd.n1673 gnd.n1654 9.3005
R18982 gnd.n1670 gnd.n1655 9.3005
R18983 gnd.n1669 gnd.n1656 9.3005
R18984 gnd.n1668 gnd.n1657 9.3005
R18985 gnd.n1666 gnd.n1658 9.3005
R18986 gnd.n1665 gnd.n1659 9.3005
R18987 gnd.n1663 gnd.n1660 9.3005
R18988 gnd.n1662 gnd.n1661 9.3005
R18989 gnd.n1558 gnd.n1557 9.3005
R18990 gnd.n4256 gnd.n4255 9.3005
R18991 gnd.n4257 gnd.n1556 9.3005
R18992 gnd.n4259 gnd.n4258 9.3005
R18993 gnd.n4260 gnd.n1555 9.3005
R18994 gnd.n4263 gnd.n4262 9.3005
R18995 gnd.n4264 gnd.n1554 9.3005
R18996 gnd.n4274 gnd.n4265 9.3005
R18997 gnd.n4273 gnd.n4266 9.3005
R18998 gnd.n4272 gnd.n4267 9.3005
R18999 gnd.n4271 gnd.n4269 9.3005
R19000 gnd.n4268 gnd.n299 9.3005
R19001 gnd.n7134 gnd.n300 9.3005
R19002 gnd.n7136 gnd.n7135 9.3005
R19003 gnd.n7196 gnd.n7137 9.3005
R19004 gnd.n7195 gnd.n7138 9.3005
R19005 gnd.n7194 gnd.n7139 9.3005
R19006 gnd.n7190 gnd.n7140 9.3005
R19007 gnd.n7189 gnd.n7141 9.3005
R19008 gnd.n7186 gnd.n7142 9.3005
R19009 gnd.n7185 gnd.n7143 9.3005
R19010 gnd.n7183 gnd.n7144 9.3005
R19011 gnd.n7182 gnd.n7145 9.3005
R19012 gnd.n7180 gnd.n7146 9.3005
R19013 gnd.n7179 gnd.n7147 9.3005
R19014 gnd.n7177 gnd.n7148 9.3005
R19015 gnd.n7176 gnd.n7149 9.3005
R19016 gnd.n7174 gnd.n7150 9.3005
R19017 gnd.n7173 gnd.n7151 9.3005
R19018 gnd.n7171 gnd.n7152 9.3005
R19019 gnd.n7170 gnd.n7153 9.3005
R19020 gnd.n7168 gnd.n7154 9.3005
R19021 gnd.n7167 gnd.n7155 9.3005
R19022 gnd.n7165 gnd.n7156 9.3005
R19023 gnd.n7164 gnd.n7157 9.3005
R19024 gnd.n7162 gnd.n7158 9.3005
R19025 gnd.n7161 gnd.n7160 9.3005
R19026 gnd.n7159 gnd.n182 9.3005
R19027 gnd.n7384 gnd.n181 9.3005
R19028 gnd.n7386 gnd.n7385 9.3005
R19029 gnd.n1496 gnd.n1494 9.3005
R19030 gnd.n4356 gnd.n4355 9.3005
R19031 gnd.n4357 gnd.n1488 9.3005
R19032 gnd.n4360 gnd.n1487 9.3005
R19033 gnd.n4361 gnd.n1486 9.3005
R19034 gnd.n4364 gnd.n1485 9.3005
R19035 gnd.n4365 gnd.n1484 9.3005
R19036 gnd.n4368 gnd.n1483 9.3005
R19037 gnd.n4369 gnd.n1482 9.3005
R19038 gnd.n4372 gnd.n1481 9.3005
R19039 gnd.n4373 gnd.n1480 9.3005
R19040 gnd.n4376 gnd.n1479 9.3005
R19041 gnd.n4377 gnd.n1478 9.3005
R19042 gnd.n4380 gnd.n1477 9.3005
R19043 gnd.n4381 gnd.n1476 9.3005
R19044 gnd.n4384 gnd.n1475 9.3005
R19045 gnd.n4385 gnd.n1474 9.3005
R19046 gnd.n4388 gnd.n1473 9.3005
R19047 gnd.n4389 gnd.n1472 9.3005
R19048 gnd.n4392 gnd.n1471 9.3005
R19049 gnd.n4394 gnd.n1465 9.3005
R19050 gnd.n4397 gnd.n1464 9.3005
R19051 gnd.n4398 gnd.n1463 9.3005
R19052 gnd.n4401 gnd.n1462 9.3005
R19053 gnd.n4402 gnd.n1461 9.3005
R19054 gnd.n4405 gnd.n1460 9.3005
R19055 gnd.n4406 gnd.n1459 9.3005
R19056 gnd.n4409 gnd.n1458 9.3005
R19057 gnd.n4410 gnd.n1457 9.3005
R19058 gnd.n4413 gnd.n1456 9.3005
R19059 gnd.n4414 gnd.n1455 9.3005
R19060 gnd.n4417 gnd.n1454 9.3005
R19061 gnd.n4419 gnd.n1453 9.3005
R19062 gnd.n4420 gnd.n1452 9.3005
R19063 gnd.n4421 gnd.n1451 9.3005
R19064 gnd.n4422 gnd.n1450 9.3005
R19065 gnd.n4354 gnd.n1493 9.3005
R19066 gnd.n4353 gnd.n4352 9.3005
R19067 gnd.n1645 gnd.n1644 9.3005
R19068 gnd.n1623 gnd.n1622 9.3005
R19069 gnd.n4178 gnd.n4177 9.3005
R19070 gnd.n4179 gnd.n1621 9.3005
R19071 gnd.n4183 gnd.n4180 9.3005
R19072 gnd.n4182 gnd.n4181 9.3005
R19073 gnd.n1595 gnd.n1594 9.3005
R19074 gnd.n4209 gnd.n4208 9.3005
R19075 gnd.n4210 gnd.n1593 9.3005
R19076 gnd.n4214 gnd.n4211 9.3005
R19077 gnd.n4213 gnd.n4212 9.3005
R19078 gnd.n1568 gnd.n1567 9.3005
R19079 gnd.n4246 gnd.n4245 9.3005
R19080 gnd.n4247 gnd.n1566 9.3005
R19081 gnd.n4251 gnd.n4248 9.3005
R19082 gnd.n4250 gnd.n4249 9.3005
R19083 gnd.n1533 gnd.n1532 9.3005
R19084 gnd.n4309 gnd.n4308 9.3005
R19085 gnd.n4310 gnd.n1531 9.3005
R19086 gnd.n4312 gnd.n4311 9.3005
R19087 gnd.n275 gnd.n268 9.3005
R19088 gnd.n254 gnd.n253 9.3005
R19089 gnd.n7237 gnd.n7236 9.3005
R19090 gnd.n7238 gnd.n252 9.3005
R19091 gnd.n7240 gnd.n7239 9.3005
R19092 gnd.n236 gnd.n235 9.3005
R19093 gnd.n7253 gnd.n7252 9.3005
R19094 gnd.n7254 gnd.n234 9.3005
R19095 gnd.n7256 gnd.n7255 9.3005
R19096 gnd.n223 gnd.n222 9.3005
R19097 gnd.n7269 gnd.n7268 9.3005
R19098 gnd.n7270 gnd.n221 9.3005
R19099 gnd.n7272 gnd.n7271 9.3005
R19100 gnd.n206 gnd.n205 9.3005
R19101 gnd.n7285 gnd.n7284 9.3005
R19102 gnd.n7286 gnd.n204 9.3005
R19103 gnd.n7288 gnd.n7287 9.3005
R19104 gnd.n191 gnd.n190 9.3005
R19105 gnd.n7376 gnd.n7375 9.3005
R19106 gnd.n7377 gnd.n189 9.3005
R19107 gnd.n7379 gnd.n7378 9.3005
R19108 gnd.n111 gnd.n110 9.3005
R19109 gnd.n7459 gnd.n7458 9.3005
R19110 gnd.n1643 gnd.n1642 9.3005
R19111 gnd.n7223 gnd.n273 9.3005
R19112 gnd.n7224 gnd.n7223 9.3005
R19113 gnd.n2385 gnd.n2384 9.3005
R19114 gnd.n2369 gnd.n2368 9.3005
R19115 gnd.n2380 gnd.n2371 9.3005
R19116 gnd.n2379 gnd.n2372 9.3005
R19117 gnd.n2378 gnd.n2373 9.3005
R19118 gnd.n2376 gnd.n2375 9.3005
R19119 gnd.n2374 gnd.n2338 9.3005
R19120 gnd.n2336 gnd.n2335 9.3005
R19121 gnd.n2714 gnd.n2713 9.3005
R19122 gnd.n2715 gnd.n2334 9.3005
R19123 gnd.n2717 gnd.n2716 9.3005
R19124 gnd.n2332 gnd.n2331 9.3005
R19125 gnd.n2722 gnd.n2721 9.3005
R19126 gnd.n2723 gnd.n2330 9.3005
R19127 gnd.n2761 gnd.n2724 9.3005
R19128 gnd.n2760 gnd.n2725 9.3005
R19129 gnd.n2759 gnd.n2726 9.3005
R19130 gnd.n2729 gnd.n2727 9.3005
R19131 gnd.n2755 gnd.n2730 9.3005
R19132 gnd.n2754 gnd.n2731 9.3005
R19133 gnd.n2753 gnd.n2732 9.3005
R19134 gnd.n2735 gnd.n2733 9.3005
R19135 gnd.n2749 gnd.n2736 9.3005
R19136 gnd.n2748 gnd.n2737 9.3005
R19137 gnd.n2747 gnd.n2738 9.3005
R19138 gnd.n2740 gnd.n2739 9.3005
R19139 gnd.n2742 gnd.n2741 9.3005
R19140 gnd.n2157 gnd.n2156 9.3005
R19141 gnd.n3732 gnd.n3731 9.3005
R19142 gnd.n3733 gnd.n2155 9.3005
R19143 gnd.n3735 gnd.n3734 9.3005
R19144 gnd.n2143 gnd.n2142 9.3005
R19145 gnd.n3748 gnd.n3747 9.3005
R19146 gnd.n3749 gnd.n2141 9.3005
R19147 gnd.n3751 gnd.n3750 9.3005
R19148 gnd.n2131 gnd.n2130 9.3005
R19149 gnd.n3764 gnd.n3763 9.3005
R19150 gnd.n3765 gnd.n2129 9.3005
R19151 gnd.n3767 gnd.n3766 9.3005
R19152 gnd.n2118 gnd.n2117 9.3005
R19153 gnd.n3780 gnd.n3779 9.3005
R19154 gnd.n3781 gnd.n2116 9.3005
R19155 gnd.n3783 gnd.n3782 9.3005
R19156 gnd.n2105 gnd.n2104 9.3005
R19157 gnd.n3796 gnd.n3795 9.3005
R19158 gnd.n3797 gnd.n2103 9.3005
R19159 gnd.n3799 gnd.n3798 9.3005
R19160 gnd.n2091 gnd.n2090 9.3005
R19161 gnd.n3812 gnd.n3811 9.3005
R19162 gnd.n3813 gnd.n2089 9.3005
R19163 gnd.n3815 gnd.n3814 9.3005
R19164 gnd.n2079 gnd.n2078 9.3005
R19165 gnd.n3828 gnd.n3827 9.3005
R19166 gnd.n3829 gnd.n2077 9.3005
R19167 gnd.n3831 gnd.n3830 9.3005
R19168 gnd.n2064 gnd.n2063 9.3005
R19169 gnd.n3844 gnd.n3843 9.3005
R19170 gnd.n3845 gnd.n2062 9.3005
R19171 gnd.n3847 gnd.n3846 9.3005
R19172 gnd.n2049 gnd.n2048 9.3005
R19173 gnd.n3860 gnd.n3859 9.3005
R19174 gnd.n3861 gnd.n2047 9.3005
R19175 gnd.n3863 gnd.n3862 9.3005
R19176 gnd.n2036 gnd.n2035 9.3005
R19177 gnd.n3876 gnd.n3875 9.3005
R19178 gnd.n3877 gnd.n2034 9.3005
R19179 gnd.n3879 gnd.n3878 9.3005
R19180 gnd.n2021 gnd.n2020 9.3005
R19181 gnd.n3892 gnd.n3891 9.3005
R19182 gnd.n3893 gnd.n2019 9.3005
R19183 gnd.n3895 gnd.n3894 9.3005
R19184 gnd.n2006 gnd.n2005 9.3005
R19185 gnd.n3908 gnd.n3907 9.3005
R19186 gnd.n3909 gnd.n2004 9.3005
R19187 gnd.n3911 gnd.n3910 9.3005
R19188 gnd.n1993 gnd.n1992 9.3005
R19189 gnd.n3924 gnd.n3923 9.3005
R19190 gnd.n3925 gnd.n1991 9.3005
R19191 gnd.n3927 gnd.n3926 9.3005
R19192 gnd.n1979 gnd.n1978 9.3005
R19193 gnd.n3940 gnd.n3939 9.3005
R19194 gnd.n3941 gnd.n1977 9.3005
R19195 gnd.n3943 gnd.n3942 9.3005
R19196 gnd.n1964 gnd.n1963 9.3005
R19197 gnd.n3956 gnd.n3955 9.3005
R19198 gnd.n3957 gnd.n1962 9.3005
R19199 gnd.n3959 gnd.n3958 9.3005
R19200 gnd.n1951 gnd.n1950 9.3005
R19201 gnd.n3972 gnd.n3971 9.3005
R19202 gnd.n3973 gnd.n1949 9.3005
R19203 gnd.n3975 gnd.n3974 9.3005
R19204 gnd.n1936 gnd.n1935 9.3005
R19205 gnd.n3988 gnd.n3987 9.3005
R19206 gnd.n3989 gnd.n1934 9.3005
R19207 gnd.n3991 gnd.n3990 9.3005
R19208 gnd.n1923 gnd.n1922 9.3005
R19209 gnd.n4004 gnd.n4003 9.3005
R19210 gnd.n4005 gnd.n1921 9.3005
R19211 gnd.n4007 gnd.n4006 9.3005
R19212 gnd.n1909 gnd.n1908 9.3005
R19213 gnd.n4020 gnd.n4019 9.3005
R19214 gnd.n4021 gnd.n1907 9.3005
R19215 gnd.n4023 gnd.n4022 9.3005
R19216 gnd.n1894 gnd.n1893 9.3005
R19217 gnd.n4036 gnd.n4035 9.3005
R19218 gnd.n4037 gnd.n1892 9.3005
R19219 gnd.n4039 gnd.n4038 9.3005
R19220 gnd.n1882 gnd.n1881 9.3005
R19221 gnd.n4052 gnd.n4051 9.3005
R19222 gnd.n4053 gnd.n1880 9.3005
R19223 gnd.n4055 gnd.n4054 9.3005
R19224 gnd.n1869 gnd.n1868 9.3005
R19225 gnd.n4068 gnd.n4067 9.3005
R19226 gnd.n4069 gnd.n1867 9.3005
R19227 gnd.n4071 gnd.n4070 9.3005
R19228 gnd.n1856 gnd.n1855 9.3005
R19229 gnd.n4084 gnd.n4083 9.3005
R19230 gnd.n4085 gnd.n1854 9.3005
R19231 gnd.n4087 gnd.n4086 9.3005
R19232 gnd.n1842 gnd.n1841 9.3005
R19233 gnd.n4100 gnd.n4099 9.3005
R19234 gnd.n4101 gnd.n1840 9.3005
R19235 gnd.n4103 gnd.n4102 9.3005
R19236 gnd.n1829 gnd.n1828 9.3005
R19237 gnd.n4118 gnd.n4117 9.3005
R19238 gnd.n4119 gnd.n1827 9.3005
R19239 gnd.n4124 gnd.n4120 9.3005
R19240 gnd.n4123 gnd.n4122 9.3005
R19241 gnd.n4121 gnd.n1411 9.3005
R19242 gnd.n4431 gnd.n1412 9.3005
R19243 gnd.n4430 gnd.n1413 9.3005
R19244 gnd.n4429 gnd.n1414 9.3005
R19245 gnd.n1636 gnd.n1415 9.3005
R19246 gnd.n1637 gnd.n1635 9.3005
R19247 gnd.n1639 gnd.n1638 9.3005
R19248 gnd.n1633 gnd.n1632 9.3005
R19249 gnd.n4167 gnd.n4166 9.3005
R19250 gnd.n4168 gnd.n1631 9.3005
R19251 gnd.n4172 gnd.n4169 9.3005
R19252 gnd.n4171 gnd.n4170 9.3005
R19253 gnd.n1606 gnd.n1605 9.3005
R19254 gnd.n4198 gnd.n4197 9.3005
R19255 gnd.n4199 gnd.n1604 9.3005
R19256 gnd.n4203 gnd.n4200 9.3005
R19257 gnd.n4202 gnd.n4201 9.3005
R19258 gnd.n1578 gnd.n1577 9.3005
R19259 gnd.n4234 gnd.n4233 9.3005
R19260 gnd.n4235 gnd.n1576 9.3005
R19261 gnd.n4239 gnd.n4236 9.3005
R19262 gnd.n4238 gnd.n4237 9.3005
R19263 gnd.n1544 gnd.n1543 9.3005
R19264 gnd.n4292 gnd.n4291 9.3005
R19265 gnd.n4293 gnd.n1542 9.3005
R19266 gnd.n4303 gnd.n4294 9.3005
R19267 gnd.n4302 gnd.n4295 9.3005
R19268 gnd.n4301 gnd.n4296 9.3005
R19269 gnd.n7102 gnd.n326 9.3005
R19270 gnd.n7101 gnd.n327 9.3005
R19271 gnd.n7094 gnd.n328 9.3005
R19272 gnd.n3642 gnd.n2288 9.3005
R19273 gnd.n3645 gnd.n2287 9.3005
R19274 gnd.n3646 gnd.n2286 9.3005
R19275 gnd.n3649 gnd.n2285 9.3005
R19276 gnd.n3650 gnd.n2284 9.3005
R19277 gnd.n3653 gnd.n2283 9.3005
R19278 gnd.n3654 gnd.n2282 9.3005
R19279 gnd.n3657 gnd.n2281 9.3005
R19280 gnd.n3658 gnd.n2280 9.3005
R19281 gnd.n3661 gnd.n2279 9.3005
R19282 gnd.n3662 gnd.n2278 9.3005
R19283 gnd.n3665 gnd.n2277 9.3005
R19284 gnd.n3666 gnd.n2276 9.3005
R19285 gnd.n3667 gnd.n2275 9.3005
R19286 gnd.n2274 gnd.n2271 9.3005
R19287 gnd.n2273 gnd.n2272 9.3005
R19288 gnd.n2867 gnd.n2866 9.3005
R19289 gnd.n2863 gnd.n2293 9.3005
R19290 gnd.n2860 gnd.n2294 9.3005
R19291 gnd.n2859 gnd.n2295 9.3005
R19292 gnd.n2856 gnd.n2296 9.3005
R19293 gnd.n2855 gnd.n2297 9.3005
R19294 gnd.n2852 gnd.n2298 9.3005
R19295 gnd.n2851 gnd.n2299 9.3005
R19296 gnd.n2848 gnd.n2300 9.3005
R19297 gnd.n2847 gnd.n2301 9.3005
R19298 gnd.n2844 gnd.n2302 9.3005
R19299 gnd.n2843 gnd.n2303 9.3005
R19300 gnd.n2840 gnd.n2304 9.3005
R19301 gnd.n2839 gnd.n2305 9.3005
R19302 gnd.n2836 gnd.n2306 9.3005
R19303 gnd.n2835 gnd.n2307 9.3005
R19304 gnd.n2832 gnd.n2308 9.3005
R19305 gnd.n2831 gnd.n2309 9.3005
R19306 gnd.n2828 gnd.n2827 9.3005
R19307 gnd.n2826 gnd.n2311 9.3005
R19308 gnd.n2868 gnd.n2289 9.3005
R19309 gnd.n2455 gnd.n2454 9.3005
R19310 gnd.n2539 gnd.n2538 9.3005
R19311 gnd.n2540 gnd.n2453 9.3005
R19312 gnd.n2543 gnd.n2541 9.3005
R19313 gnd.n2544 gnd.n2452 9.3005
R19314 gnd.n2547 gnd.n2546 9.3005
R19315 gnd.n2548 gnd.n2451 9.3005
R19316 gnd.n2551 gnd.n2549 9.3005
R19317 gnd.n2552 gnd.n2450 9.3005
R19318 gnd.n2555 gnd.n2554 9.3005
R19319 gnd.n2556 gnd.n2449 9.3005
R19320 gnd.n2559 gnd.n2557 9.3005
R19321 gnd.n2560 gnd.n2448 9.3005
R19322 gnd.n2563 gnd.n2562 9.3005
R19323 gnd.n2564 gnd.n2447 9.3005
R19324 gnd.n2567 gnd.n2565 9.3005
R19325 gnd.n2568 gnd.n2446 9.3005
R19326 gnd.n2571 gnd.n2570 9.3005
R19327 gnd.n2572 gnd.n2445 9.3005
R19328 gnd.n2575 gnd.n2574 9.3005
R19329 gnd.n2573 gnd.n2400 9.3005
R19330 gnd.n2631 gnd.n2401 9.3005
R19331 gnd.n2630 gnd.n2402 9.3005
R19332 gnd.n2629 gnd.n2403 9.3005
R19333 gnd.n2600 gnd.n2404 9.3005
R19334 gnd.n2619 gnd.n2601 9.3005
R19335 gnd.n2481 gnd.n2480 9.3005
R19336 gnd.n2486 gnd.n2485 9.3005
R19337 gnd.n2489 gnd.n2475 9.3005
R19338 gnd.n2490 gnd.n2474 9.3005
R19339 gnd.n2493 gnd.n2473 9.3005
R19340 gnd.n2494 gnd.n2472 9.3005
R19341 gnd.n2497 gnd.n2471 9.3005
R19342 gnd.n2498 gnd.n2470 9.3005
R19343 gnd.n2501 gnd.n2469 9.3005
R19344 gnd.n2502 gnd.n2468 9.3005
R19345 gnd.n2505 gnd.n2467 9.3005
R19346 gnd.n2506 gnd.n2466 9.3005
R19347 gnd.n2509 gnd.n2465 9.3005
R19348 gnd.n2510 gnd.n2464 9.3005
R19349 gnd.n2513 gnd.n2463 9.3005
R19350 gnd.n2514 gnd.n2462 9.3005
R19351 gnd.n2517 gnd.n2461 9.3005
R19352 gnd.n2520 gnd.n2519 9.3005
R19353 gnd.n2484 gnd.n2479 9.3005
R19354 gnd.n2483 gnd.n2482 9.3005
R19355 gnd.n2527 gnd.n2526 9.3005
R19356 gnd.n2525 gnd.n2460 9.3005
R19357 gnd.n2524 gnd.n2523 9.3005
R19358 gnd.n2522 gnd.n1032 9.3005
R19359 gnd.n4737 gnd.n1033 9.3005
R19360 gnd.n4736 gnd.n1034 9.3005
R19361 gnd.n4735 gnd.n1035 9.3005
R19362 gnd.n1051 gnd.n1036 9.3005
R19363 gnd.n4725 gnd.n1052 9.3005
R19364 gnd.n4724 gnd.n1053 9.3005
R19365 gnd.n4723 gnd.n1054 9.3005
R19366 gnd.n1072 gnd.n1055 9.3005
R19367 gnd.n4713 gnd.n1073 9.3005
R19368 gnd.n4712 gnd.n1074 9.3005
R19369 gnd.n4711 gnd.n1075 9.3005
R19370 gnd.n1091 gnd.n1076 9.3005
R19371 gnd.n4701 gnd.n1092 9.3005
R19372 gnd.n4700 gnd.n1093 9.3005
R19373 gnd.n4699 gnd.n1094 9.3005
R19374 gnd.n1114 gnd.n1095 9.3005
R19375 gnd.n4689 gnd.n1115 9.3005
R19376 gnd.n4688 gnd.n1116 9.3005
R19377 gnd.n4687 gnd.n1117 9.3005
R19378 gnd.n1132 gnd.n1118 9.3005
R19379 gnd.n4677 gnd.n1133 9.3005
R19380 gnd.n4676 gnd.n1134 9.3005
R19381 gnd.n4675 gnd.n1135 9.3005
R19382 gnd.n1151 gnd.n1136 9.3005
R19383 gnd.n4664 gnd.n1152 9.3005
R19384 gnd.n4663 gnd.n1153 9.3005
R19385 gnd.n4662 gnd.n1154 9.3005
R19386 gnd.n1170 gnd.n1155 9.3005
R19387 gnd.n4652 gnd.n1171 9.3005
R19388 gnd.n4651 gnd.n1172 9.3005
R19389 gnd.n4650 gnd.n1173 9.3005
R19390 gnd.n1192 gnd.n1174 9.3005
R19391 gnd.n4640 gnd.n1193 9.3005
R19392 gnd.n4639 gnd.n1194 9.3005
R19393 gnd.n4638 gnd.n1195 9.3005
R19394 gnd.n1212 gnd.n1196 9.3005
R19395 gnd.n4628 gnd.n1213 9.3005
R19396 gnd.n4627 gnd.n1214 9.3005
R19397 gnd.n4626 gnd.n1215 9.3005
R19398 gnd.n1234 gnd.n1216 9.3005
R19399 gnd.n4616 gnd.n1235 9.3005
R19400 gnd.n4615 gnd.n1236 9.3005
R19401 gnd.n4614 gnd.n1237 9.3005
R19402 gnd.n1255 gnd.n1238 9.3005
R19403 gnd.n4604 gnd.n1256 9.3005
R19404 gnd.n4603 gnd.n1257 9.3005
R19405 gnd.n4602 gnd.n1258 9.3005
R19406 gnd.n1275 gnd.n1259 9.3005
R19407 gnd.n4592 gnd.n4591 9.3005
R19408 gnd.n2521 gnd.n2459 9.3005
R19409 gnd.n4751 gnd.n4750 9.3005
R19410 gnd.n4749 gnd.n1010 9.3005
R19411 gnd.n4748 gnd.n4747 9.3005
R19412 gnd.n1012 gnd.n1011 9.3005
R19413 gnd.n2415 gnd.n2414 9.3005
R19414 gnd.n2418 gnd.n2417 9.3005
R19415 gnd.n2419 gnd.n2413 9.3005
R19416 gnd.n2422 gnd.n2420 9.3005
R19417 gnd.n2423 gnd.n2412 9.3005
R19418 gnd.n2426 gnd.n2425 9.3005
R19419 gnd.n2427 gnd.n2411 9.3005
R19420 gnd.n2430 gnd.n2428 9.3005
R19421 gnd.n2431 gnd.n2410 9.3005
R19422 gnd.n2434 gnd.n2433 9.3005
R19423 gnd.n2435 gnd.n2409 9.3005
R19424 gnd.n2438 gnd.n2436 9.3005
R19425 gnd.n2439 gnd.n2408 9.3005
R19426 gnd.n2442 gnd.n2441 9.3005
R19427 gnd.n2443 gnd.n2407 9.3005
R19428 gnd.n2579 gnd.n2444 9.3005
R19429 gnd.n2580 gnd.n2406 9.3005
R19430 gnd.n2582 gnd.n2581 9.3005
R19431 gnd.n2583 gnd.n2405 9.3005
R19432 gnd.n2625 gnd.n2584 9.3005
R19433 gnd.n2624 gnd.n2585 9.3005
R19434 gnd.n2623 gnd.n2586 9.3005
R19435 gnd.n2604 gnd.n2587 9.3005
R19436 gnd.n2610 gnd.n2605 9.3005
R19437 gnd.n2609 gnd.n2606 9.3005
R19438 gnd.n2608 gnd.n2607 9.3005
R19439 gnd.n2359 gnd.n2358 9.3005
R19440 gnd.n2655 gnd.n2654 9.3005
R19441 gnd.n2656 gnd.n2357 9.3005
R19442 gnd.n2659 gnd.n2658 9.3005
R19443 gnd.n2657 gnd.n2351 9.3005
R19444 gnd.n2671 gnd.n2352 9.3005
R19445 gnd.n2672 gnd.n2350 9.3005
R19446 gnd.n2674 gnd.n2673 9.3005
R19447 gnd.n2675 gnd.n2349 9.3005
R19448 gnd.n2679 gnd.n2676 9.3005
R19449 gnd.n2680 gnd.n2348 9.3005
R19450 gnd.n2685 gnd.n2684 9.3005
R19451 gnd.n2686 gnd.n2347 9.3005
R19452 gnd.n2692 gnd.n2687 9.3005
R19453 gnd.n2691 gnd.n2688 9.3005
R19454 gnd.n2690 gnd.n2689 9.3005
R19455 gnd.n2323 gnd.n2322 9.3005
R19456 gnd.n2775 gnd.n2774 9.3005
R19457 gnd.n2776 gnd.n2321 9.3005
R19458 gnd.n2779 gnd.n2778 9.3005
R19459 gnd.n2777 gnd.n2315 9.3005
R19460 gnd.n2823 gnd.n2314 9.3005
R19461 gnd.n2825 gnd.n2824 9.3005
R19462 gnd.n4752 gnd.n1008 9.3005
R19463 gnd.n4759 gnd.n4758 9.3005
R19464 gnd.n4760 gnd.n1002 9.3005
R19465 gnd.n4763 gnd.n1001 9.3005
R19466 gnd.n4764 gnd.n1000 9.3005
R19467 gnd.n4767 gnd.n999 9.3005
R19468 gnd.n4768 gnd.n998 9.3005
R19469 gnd.n4771 gnd.n997 9.3005
R19470 gnd.n4772 gnd.n996 9.3005
R19471 gnd.n4775 gnd.n995 9.3005
R19472 gnd.n4776 gnd.n994 9.3005
R19473 gnd.n4779 gnd.n993 9.3005
R19474 gnd.n4780 gnd.n992 9.3005
R19475 gnd.n4783 gnd.n991 9.3005
R19476 gnd.n4784 gnd.n990 9.3005
R19477 gnd.n4787 gnd.n989 9.3005
R19478 gnd.n4788 gnd.n988 9.3005
R19479 gnd.n4791 gnd.n987 9.3005
R19480 gnd.n4792 gnd.n986 9.3005
R19481 gnd.n4795 gnd.n985 9.3005
R19482 gnd.n4797 gnd.n982 9.3005
R19483 gnd.n4800 gnd.n981 9.3005
R19484 gnd.n4801 gnd.n980 9.3005
R19485 gnd.n4804 gnd.n979 9.3005
R19486 gnd.n4805 gnd.n978 9.3005
R19487 gnd.n4808 gnd.n977 9.3005
R19488 gnd.n4809 gnd.n976 9.3005
R19489 gnd.n4812 gnd.n975 9.3005
R19490 gnd.n4813 gnd.n974 9.3005
R19491 gnd.n4816 gnd.n973 9.3005
R19492 gnd.n4817 gnd.n972 9.3005
R19493 gnd.n4820 gnd.n971 9.3005
R19494 gnd.n4821 gnd.n970 9.3005
R19495 gnd.n4824 gnd.n969 9.3005
R19496 gnd.n4826 gnd.n968 9.3005
R19497 gnd.n4827 gnd.n967 9.3005
R19498 gnd.n4828 gnd.n966 9.3005
R19499 gnd.n4829 gnd.n965 9.3005
R19500 gnd.n4757 gnd.n1007 9.3005
R19501 gnd.n4756 gnd.n4755 9.3005
R19502 gnd.n2533 gnd.n2532 9.3005
R19503 gnd.n2531 gnd.n1021 9.3005
R19504 gnd.n4743 gnd.n1022 9.3005
R19505 gnd.n4742 gnd.n1023 9.3005
R19506 gnd.n4741 gnd.n1024 9.3005
R19507 gnd.n1042 gnd.n1025 9.3005
R19508 gnd.n4731 gnd.n1043 9.3005
R19509 gnd.n4730 gnd.n1044 9.3005
R19510 gnd.n4729 gnd.n1045 9.3005
R19511 gnd.n1061 gnd.n1046 9.3005
R19512 gnd.n4719 gnd.n1062 9.3005
R19513 gnd.n4718 gnd.n1063 9.3005
R19514 gnd.n4717 gnd.n1064 9.3005
R19515 gnd.n1082 gnd.n1065 9.3005
R19516 gnd.n4707 gnd.n1083 9.3005
R19517 gnd.n4706 gnd.n1084 9.3005
R19518 gnd.n4705 gnd.n1085 9.3005
R19519 gnd.n1103 gnd.n1086 9.3005
R19520 gnd.n4695 gnd.n1104 9.3005
R19521 gnd.n4694 gnd.n1105 9.3005
R19522 gnd.n4693 gnd.n1106 9.3005
R19523 gnd.n4657 gnd.n1162 9.3005
R19524 gnd.n4656 gnd.n1163 9.3005
R19525 gnd.n1181 gnd.n1164 9.3005
R19526 gnd.n4646 gnd.n1182 9.3005
R19527 gnd.n4645 gnd.n1183 9.3005
R19528 gnd.n4644 gnd.n1184 9.3005
R19529 gnd.n1202 gnd.n1185 9.3005
R19530 gnd.n4634 gnd.n1203 9.3005
R19531 gnd.n4633 gnd.n1204 9.3005
R19532 gnd.n4632 gnd.n1205 9.3005
R19533 gnd.n1223 gnd.n1206 9.3005
R19534 gnd.n4622 gnd.n1224 9.3005
R19535 gnd.n4621 gnd.n1225 9.3005
R19536 gnd.n4620 gnd.n1226 9.3005
R19537 gnd.n1244 gnd.n1227 9.3005
R19538 gnd.n4610 gnd.n1245 9.3005
R19539 gnd.n4609 gnd.n1246 9.3005
R19540 gnd.n4608 gnd.n1247 9.3005
R19541 gnd.n1265 gnd.n1248 9.3005
R19542 gnd.n4598 gnd.n1266 9.3005
R19543 gnd.n4597 gnd.n1267 9.3005
R19544 gnd.n4596 gnd.n1268 9.3005
R19545 gnd.n2530 gnd.n2529 9.3005
R19546 gnd.n4682 gnd.n1125 9.3005
R19547 gnd.n4658 gnd.n1125 9.3005
R19548 gnd.n2391 gnd.n2390 9.3005
R19549 gnd.n2638 gnd.n2637 9.3005
R19550 gnd.n2395 gnd.n2394 9.3005
R19551 gnd.n6261 gnd.n893 9.3005
R19552 gnd.n6262 gnd.n892 9.3005
R19553 gnd.n6263 gnd.n891 9.3005
R19554 gnd.n890 gnd.n886 9.3005
R19555 gnd.n6269 gnd.n885 9.3005
R19556 gnd.n6270 gnd.n884 9.3005
R19557 gnd.n6271 gnd.n883 9.3005
R19558 gnd.n882 gnd.n878 9.3005
R19559 gnd.n6277 gnd.n877 9.3005
R19560 gnd.n6278 gnd.n876 9.3005
R19561 gnd.n6279 gnd.n875 9.3005
R19562 gnd.n874 gnd.n870 9.3005
R19563 gnd.n6285 gnd.n869 9.3005
R19564 gnd.n6286 gnd.n868 9.3005
R19565 gnd.n6287 gnd.n867 9.3005
R19566 gnd.n866 gnd.n862 9.3005
R19567 gnd.n6293 gnd.n861 9.3005
R19568 gnd.n6294 gnd.n860 9.3005
R19569 gnd.n6295 gnd.n859 9.3005
R19570 gnd.n858 gnd.n854 9.3005
R19571 gnd.n6301 gnd.n853 9.3005
R19572 gnd.n6302 gnd.n852 9.3005
R19573 gnd.n6303 gnd.n851 9.3005
R19574 gnd.n850 gnd.n846 9.3005
R19575 gnd.n6309 gnd.n845 9.3005
R19576 gnd.n6310 gnd.n844 9.3005
R19577 gnd.n6311 gnd.n843 9.3005
R19578 gnd.n842 gnd.n838 9.3005
R19579 gnd.n6317 gnd.n837 9.3005
R19580 gnd.n6318 gnd.n836 9.3005
R19581 gnd.n6319 gnd.n835 9.3005
R19582 gnd.n834 gnd.n830 9.3005
R19583 gnd.n6325 gnd.n829 9.3005
R19584 gnd.n6326 gnd.n828 9.3005
R19585 gnd.n6327 gnd.n827 9.3005
R19586 gnd.n826 gnd.n822 9.3005
R19587 gnd.n6333 gnd.n821 9.3005
R19588 gnd.n6334 gnd.n820 9.3005
R19589 gnd.n6335 gnd.n819 9.3005
R19590 gnd.n818 gnd.n814 9.3005
R19591 gnd.n6341 gnd.n813 9.3005
R19592 gnd.n6342 gnd.n812 9.3005
R19593 gnd.n6343 gnd.n811 9.3005
R19594 gnd.n810 gnd.n806 9.3005
R19595 gnd.n6349 gnd.n805 9.3005
R19596 gnd.n6350 gnd.n804 9.3005
R19597 gnd.n6351 gnd.n803 9.3005
R19598 gnd.n802 gnd.n798 9.3005
R19599 gnd.n6357 gnd.n797 9.3005
R19600 gnd.n6358 gnd.n796 9.3005
R19601 gnd.n6359 gnd.n795 9.3005
R19602 gnd.n794 gnd.n790 9.3005
R19603 gnd.n6365 gnd.n789 9.3005
R19604 gnd.n6366 gnd.n788 9.3005
R19605 gnd.n6367 gnd.n787 9.3005
R19606 gnd.n786 gnd.n782 9.3005
R19607 gnd.n6373 gnd.n781 9.3005
R19608 gnd.n6374 gnd.n780 9.3005
R19609 gnd.n6375 gnd.n779 9.3005
R19610 gnd.n778 gnd.n774 9.3005
R19611 gnd.n6381 gnd.n773 9.3005
R19612 gnd.n6382 gnd.n772 9.3005
R19613 gnd.n6383 gnd.n771 9.3005
R19614 gnd.n770 gnd.n766 9.3005
R19615 gnd.n6389 gnd.n765 9.3005
R19616 gnd.n6390 gnd.n764 9.3005
R19617 gnd.n6391 gnd.n763 9.3005
R19618 gnd.n762 gnd.n758 9.3005
R19619 gnd.n6397 gnd.n757 9.3005
R19620 gnd.n6398 gnd.n756 9.3005
R19621 gnd.n6399 gnd.n755 9.3005
R19622 gnd.n754 gnd.n750 9.3005
R19623 gnd.n6405 gnd.n749 9.3005
R19624 gnd.n6406 gnd.n748 9.3005
R19625 gnd.n6407 gnd.n747 9.3005
R19626 gnd.n746 gnd.n742 9.3005
R19627 gnd.n6413 gnd.n741 9.3005
R19628 gnd.n6414 gnd.n740 9.3005
R19629 gnd.n6415 gnd.n739 9.3005
R19630 gnd.n738 gnd.n734 9.3005
R19631 gnd.n6421 gnd.n733 9.3005
R19632 gnd.n6422 gnd.n732 9.3005
R19633 gnd.n6423 gnd.n731 9.3005
R19634 gnd.n730 gnd.n726 9.3005
R19635 gnd.n2393 gnd.n894 9.3005
R19636 gnd.n1735 gnd.n1734 9.3005
R19637 gnd.n1721 gnd.n1717 9.3005
R19638 gnd.n1742 gnd.n1741 9.3005
R19639 gnd.n1743 gnd.n1712 9.3005
R19640 gnd.n1754 gnd.n1753 9.3005
R19641 gnd.n1714 gnd.n1710 9.3005
R19642 gnd.n1761 gnd.n1760 9.3005
R19643 gnd.n1762 gnd.n1705 9.3005
R19644 gnd.n1773 gnd.n1772 9.3005
R19645 gnd.n1707 gnd.n1703 9.3005
R19646 gnd.n1780 gnd.n1779 9.3005
R19647 gnd.n1700 gnd.n1699 9.3005
R19648 gnd.n1789 gnd.n1788 9.3005
R19649 gnd.n1697 gnd.n1696 9.3005
R19650 gnd.n1796 gnd.n1795 9.3005
R19651 gnd.n1688 gnd.n1687 9.3005
R19652 gnd.n1803 gnd.n1802 9.3005
R19653 gnd.n1685 gnd.n1683 9.3005
R19654 gnd.n1724 gnd.n1719 9.3005
R19655 gnd.n1798 gnd.n1797 9.3005
R19656 gnd.n1787 gnd.n1693 9.3005
R19657 gnd.n1786 gnd.n1785 9.3005
R19658 gnd.n1782 gnd.n1781 9.3005
R19659 gnd.n1702 gnd.n1701 9.3005
R19660 gnd.n1771 gnd.n1770 9.3005
R19661 gnd.n1767 gnd.n1706 9.3005
R19662 gnd.n1764 gnd.n1763 9.3005
R19663 gnd.n1709 gnd.n1708 9.3005
R19664 gnd.n1752 gnd.n1751 9.3005
R19665 gnd.n1748 gnd.n1713 9.3005
R19666 gnd.n1745 gnd.n1744 9.3005
R19667 gnd.n1716 gnd.n1715 9.3005
R19668 gnd.n1733 gnd.n1732 9.3005
R19669 gnd.n1729 gnd.n1720 9.3005
R19670 gnd.n1726 gnd.n1725 9.3005
R19671 gnd.n1799 gnd.n1689 9.3005
R19672 gnd.n1801 gnd.n1800 9.3005
R19673 gnd.n4154 gnd.n4153 9.3005
R19674 gnd.n4152 gnd.n1684 9.3005
R19675 gnd.n4151 gnd.n4150 9.3005
R19676 gnd.n4149 gnd.n1811 9.3005
R19677 gnd.n4148 gnd.n4147 9.3005
R19678 gnd.n4146 gnd.n1812 9.3005
R19679 gnd.n4142 gnd.n4141 9.3005
R19680 gnd.n4140 gnd.n1819 9.3005
R19681 gnd.n4139 gnd.n4138 9.3005
R19682 gnd.n4137 gnd.n4132 9.3005
R19683 gnd.n3727 gnd.n3726 9.3005
R19684 gnd.n2150 gnd.n2149 9.3005
R19685 gnd.n3740 gnd.n3739 9.3005
R19686 gnd.n3741 gnd.n2148 9.3005
R19687 gnd.n3743 gnd.n3742 9.3005
R19688 gnd.n2137 gnd.n2136 9.3005
R19689 gnd.n3756 gnd.n3755 9.3005
R19690 gnd.n3757 gnd.n2135 9.3005
R19691 gnd.n3759 gnd.n3758 9.3005
R19692 gnd.n2124 gnd.n2123 9.3005
R19693 gnd.n3772 gnd.n3771 9.3005
R19694 gnd.n3773 gnd.n2122 9.3005
R19695 gnd.n3775 gnd.n3774 9.3005
R19696 gnd.n2111 gnd.n2110 9.3005
R19697 gnd.n3788 gnd.n3787 9.3005
R19698 gnd.n3789 gnd.n2109 9.3005
R19699 gnd.n3791 gnd.n3790 9.3005
R19700 gnd.n2097 gnd.n2096 9.3005
R19701 gnd.n3804 gnd.n3803 9.3005
R19702 gnd.n3805 gnd.n2095 9.3005
R19703 gnd.n3807 gnd.n3806 9.3005
R19704 gnd.n2084 gnd.n2083 9.3005
R19705 gnd.n3820 gnd.n3819 9.3005
R19706 gnd.n3821 gnd.n2082 9.3005
R19707 gnd.n3823 gnd.n3822 9.3005
R19708 gnd.n2071 gnd.n2070 9.3005
R19709 gnd.n3836 gnd.n3835 9.3005
R19710 gnd.n3837 gnd.n2069 9.3005
R19711 gnd.n3839 gnd.n3838 9.3005
R19712 gnd.n2056 gnd.n2055 9.3005
R19713 gnd.n3852 gnd.n3851 9.3005
R19714 gnd.n3853 gnd.n2054 9.3005
R19715 gnd.n3855 gnd.n3854 9.3005
R19716 gnd.n2042 gnd.n2041 9.3005
R19717 gnd.n3868 gnd.n3867 9.3005
R19718 gnd.n3869 gnd.n2040 9.3005
R19719 gnd.n3871 gnd.n3870 9.3005
R19720 gnd.n2029 gnd.n2028 9.3005
R19721 gnd.n3884 gnd.n3883 9.3005
R19722 gnd.n3885 gnd.n2027 9.3005
R19723 gnd.n3887 gnd.n3886 9.3005
R19724 gnd.n2013 gnd.n2012 9.3005
R19725 gnd.n3900 gnd.n3899 9.3005
R19726 gnd.n3901 gnd.n2011 9.3005
R19727 gnd.n3903 gnd.n3902 9.3005
R19728 gnd.n1999 gnd.n1998 9.3005
R19729 gnd.n3916 gnd.n3915 9.3005
R19730 gnd.n3917 gnd.n1997 9.3005
R19731 gnd.n3919 gnd.n3918 9.3005
R19732 gnd.n1985 gnd.n1984 9.3005
R19733 gnd.n3932 gnd.n3931 9.3005
R19734 gnd.n3933 gnd.n1983 9.3005
R19735 gnd.n3935 gnd.n3934 9.3005
R19736 gnd.n1971 gnd.n1970 9.3005
R19737 gnd.n3948 gnd.n3947 9.3005
R19738 gnd.n3949 gnd.n1969 9.3005
R19739 gnd.n3951 gnd.n3950 9.3005
R19740 gnd.n1957 gnd.n1956 9.3005
R19741 gnd.n3964 gnd.n3963 9.3005
R19742 gnd.n3965 gnd.n1955 9.3005
R19743 gnd.n3967 gnd.n3966 9.3005
R19744 gnd.n1943 gnd.n1942 9.3005
R19745 gnd.n3980 gnd.n3979 9.3005
R19746 gnd.n3981 gnd.n1941 9.3005
R19747 gnd.n3983 gnd.n3982 9.3005
R19748 gnd.n1929 gnd.n1928 9.3005
R19749 gnd.n3996 gnd.n3995 9.3005
R19750 gnd.n3997 gnd.n1927 9.3005
R19751 gnd.n3999 gnd.n3998 9.3005
R19752 gnd.n1916 gnd.n1915 9.3005
R19753 gnd.n4012 gnd.n4011 9.3005
R19754 gnd.n4013 gnd.n1914 9.3005
R19755 gnd.n4015 gnd.n4014 9.3005
R19756 gnd.n1901 gnd.n1900 9.3005
R19757 gnd.n4028 gnd.n4027 9.3005
R19758 gnd.n4029 gnd.n1899 9.3005
R19759 gnd.n4031 gnd.n4030 9.3005
R19760 gnd.n1887 gnd.n1886 9.3005
R19761 gnd.n4044 gnd.n4043 9.3005
R19762 gnd.n4045 gnd.n1885 9.3005
R19763 gnd.n4047 gnd.n4046 9.3005
R19764 gnd.n1875 gnd.n1874 9.3005
R19765 gnd.n4060 gnd.n4059 9.3005
R19766 gnd.n4061 gnd.n1873 9.3005
R19767 gnd.n4063 gnd.n4062 9.3005
R19768 gnd.n1862 gnd.n1861 9.3005
R19769 gnd.n4076 gnd.n4075 9.3005
R19770 gnd.n4077 gnd.n1860 9.3005
R19771 gnd.n4079 gnd.n4078 9.3005
R19772 gnd.n1849 gnd.n1848 9.3005
R19773 gnd.n4092 gnd.n4091 9.3005
R19774 gnd.n4093 gnd.n1847 9.3005
R19775 gnd.n4095 gnd.n4094 9.3005
R19776 gnd.n1836 gnd.n1835 9.3005
R19777 gnd.n4108 gnd.n4107 9.3005
R19778 gnd.n4109 gnd.n1833 9.3005
R19779 gnd.n4113 gnd.n4112 9.3005
R19780 gnd.n4111 gnd.n1834 9.3005
R19781 gnd.n4110 gnd.n1821 9.3005
R19782 gnd.n4129 gnd.n1820 9.3005
R19783 gnd.n4131 gnd.n4130 9.3005
R19784 gnd.n3725 gnd.n2161 9.3005
R19785 gnd.n2163 gnd.n2162 9.3005
R19786 gnd.n2802 gnd.n2799 9.3005
R19787 gnd.n2804 gnd.n2803 9.3005
R19788 gnd.n2806 gnd.n2805 9.3005
R19789 gnd.n2807 gnd.n2792 9.3005
R19790 gnd.n2809 gnd.n2808 9.3005
R19791 gnd.n2810 gnd.n2791 9.3005
R19792 gnd.n2812 gnd.n2811 9.3005
R19793 gnd.n2813 gnd.n2786 9.3005
R19794 gnd.n3724 gnd.n3723 9.3005
R19795 gnd.n2618 gnd.n2617 9.3005
R19796 gnd.n2616 gnd.n2614 9.3005
R19797 gnd.n2362 gnd.n2361 9.3005
R19798 gnd.n2647 gnd.n2646 9.3005
R19799 gnd.n2648 gnd.n2360 9.3005
R19800 gnd.n2650 gnd.n2649 9.3005
R19801 gnd.n2355 gnd.n2354 9.3005
R19802 gnd.n2664 gnd.n2663 9.3005
R19803 gnd.n2665 gnd.n2353 9.3005
R19804 gnd.n2667 gnd.n2666 9.3005
R19805 gnd.n2342 gnd.n2340 9.3005
R19806 gnd.n2706 gnd.n2705 9.3005
R19807 gnd.n2704 gnd.n2341 9.3005
R19808 gnd.n2703 gnd.n2702 9.3005
R19809 gnd.n2701 gnd.n2343 9.3005
R19810 gnd.n2700 gnd.n2699 9.3005
R19811 gnd.n2698 gnd.n2346 9.3005
R19812 gnd.n2697 gnd.n2696 9.3005
R19813 gnd.n2326 gnd.n2325 9.3005
R19814 gnd.n2767 gnd.n2766 9.3005
R19815 gnd.n2768 gnd.n2324 9.3005
R19816 gnd.n2770 gnd.n2769 9.3005
R19817 gnd.n2320 gnd.n2319 9.3005
R19818 gnd.n2784 gnd.n2783 9.3005
R19819 gnd.n2785 gnd.n2317 9.3005
R19820 gnd.n2819 gnd.n2818 9.3005
R19821 gnd.n2817 gnd.n2318 9.3005
R19822 gnd.n2815 gnd.n2814 9.3005
R19823 gnd.n2232 gnd.n2231 9.3005
R19824 gnd.n3676 gnd.n3675 9.3005
R19825 gnd.n3678 gnd.n3677 9.3005
R19826 gnd.n2220 gnd.n2219 9.3005
R19827 gnd.n3684 gnd.n3683 9.3005
R19828 gnd.n3686 gnd.n3685 9.3005
R19829 gnd.n2212 gnd.n2211 9.3005
R19830 gnd.n3692 gnd.n3691 9.3005
R19831 gnd.n3694 gnd.n3693 9.3005
R19832 gnd.n2202 gnd.n2201 9.3005
R19833 gnd.n3700 gnd.n3699 9.3005
R19834 gnd.n3702 gnd.n3701 9.3005
R19835 gnd.n2194 gnd.n2193 9.3005
R19836 gnd.n3708 gnd.n3707 9.3005
R19837 gnd.n3710 gnd.n3709 9.3005
R19838 gnd.n2184 gnd.n2182 9.3005
R19839 gnd.n3716 gnd.n3715 9.3005
R19840 gnd.n3717 gnd.n2181 9.3005
R19841 gnd.n2235 gnd.n1277 9.3005
R19842 gnd.n2185 gnd.n2183 9.3005
R19843 gnd.n3714 gnd.n3713 9.3005
R19844 gnd.n3712 gnd.n3711 9.3005
R19845 gnd.n2189 gnd.n2188 9.3005
R19846 gnd.n3706 gnd.n3705 9.3005
R19847 gnd.n3704 gnd.n3703 9.3005
R19848 gnd.n2198 gnd.n2197 9.3005
R19849 gnd.n3698 gnd.n3697 9.3005
R19850 gnd.n3696 gnd.n3695 9.3005
R19851 gnd.n2206 gnd.n2205 9.3005
R19852 gnd.n3690 gnd.n3689 9.3005
R19853 gnd.n3688 gnd.n3687 9.3005
R19854 gnd.n2216 gnd.n2215 9.3005
R19855 gnd.n3682 gnd.n3681 9.3005
R19856 gnd.n3680 gnd.n3679 9.3005
R19857 gnd.n2226 gnd.n2225 9.3005
R19858 gnd.n3674 gnd.n3673 9.3005
R19859 gnd.n4586 gnd.n1278 9.3005
R19860 gnd.n4585 gnd.n4584 9.3005
R19861 gnd.n4583 gnd.n1282 9.3005
R19862 gnd.n4582 gnd.n4581 9.3005
R19863 gnd.n4580 gnd.n1283 9.3005
R19864 gnd.n4579 gnd.n4578 9.3005
R19865 gnd.n4577 gnd.n1287 9.3005
R19866 gnd.n4576 gnd.n4575 9.3005
R19867 gnd.n4574 gnd.n1288 9.3005
R19868 gnd.n4573 gnd.n4572 9.3005
R19869 gnd.n4571 gnd.n1292 9.3005
R19870 gnd.n4570 gnd.n4569 9.3005
R19871 gnd.n4568 gnd.n1293 9.3005
R19872 gnd.n4567 gnd.n4566 9.3005
R19873 gnd.n4565 gnd.n1297 9.3005
R19874 gnd.n4564 gnd.n4563 9.3005
R19875 gnd.n4562 gnd.n1298 9.3005
R19876 gnd.n4561 gnd.n4560 9.3005
R19877 gnd.n4559 gnd.n1302 9.3005
R19878 gnd.n4558 gnd.n4557 9.3005
R19879 gnd.n4556 gnd.n1303 9.3005
R19880 gnd.n4555 gnd.n4554 9.3005
R19881 gnd.n4553 gnd.n1307 9.3005
R19882 gnd.n4552 gnd.n4551 9.3005
R19883 gnd.n4550 gnd.n1308 9.3005
R19884 gnd.n4549 gnd.n4548 9.3005
R19885 gnd.n4547 gnd.n1312 9.3005
R19886 gnd.n4546 gnd.n4545 9.3005
R19887 gnd.n4544 gnd.n1313 9.3005
R19888 gnd.n4543 gnd.n4542 9.3005
R19889 gnd.n4541 gnd.n1317 9.3005
R19890 gnd.n4540 gnd.n4539 9.3005
R19891 gnd.n4538 gnd.n1318 9.3005
R19892 gnd.n4537 gnd.n4536 9.3005
R19893 gnd.n4535 gnd.n1322 9.3005
R19894 gnd.n4534 gnd.n4533 9.3005
R19895 gnd.n4532 gnd.n1323 9.3005
R19896 gnd.n4531 gnd.n4530 9.3005
R19897 gnd.n4529 gnd.n1327 9.3005
R19898 gnd.n4528 gnd.n4527 9.3005
R19899 gnd.n4526 gnd.n1328 9.3005
R19900 gnd.n4525 gnd.n4524 9.3005
R19901 gnd.n4523 gnd.n1332 9.3005
R19902 gnd.n4522 gnd.n4521 9.3005
R19903 gnd.n4520 gnd.n1333 9.3005
R19904 gnd.n4519 gnd.n4518 9.3005
R19905 gnd.n4517 gnd.n1337 9.3005
R19906 gnd.n4516 gnd.n4515 9.3005
R19907 gnd.n4514 gnd.n1338 9.3005
R19908 gnd.n4513 gnd.n4512 9.3005
R19909 gnd.n4511 gnd.n1342 9.3005
R19910 gnd.n4510 gnd.n4509 9.3005
R19911 gnd.n4508 gnd.n1343 9.3005
R19912 gnd.n4507 gnd.n4506 9.3005
R19913 gnd.n4505 gnd.n1347 9.3005
R19914 gnd.n4504 gnd.n4503 9.3005
R19915 gnd.n4502 gnd.n1348 9.3005
R19916 gnd.n4501 gnd.n4500 9.3005
R19917 gnd.n4499 gnd.n1352 9.3005
R19918 gnd.n4498 gnd.n4497 9.3005
R19919 gnd.n4496 gnd.n1353 9.3005
R19920 gnd.n4495 gnd.n4494 9.3005
R19921 gnd.n4493 gnd.n1357 9.3005
R19922 gnd.n4492 gnd.n4491 9.3005
R19923 gnd.n4490 gnd.n1358 9.3005
R19924 gnd.n4489 gnd.n4488 9.3005
R19925 gnd.n4487 gnd.n1362 9.3005
R19926 gnd.n4486 gnd.n4485 9.3005
R19927 gnd.n4484 gnd.n1363 9.3005
R19928 gnd.n4483 gnd.n4482 9.3005
R19929 gnd.n4481 gnd.n1367 9.3005
R19930 gnd.n4480 gnd.n4479 9.3005
R19931 gnd.n4478 gnd.n1368 9.3005
R19932 gnd.n4477 gnd.n4476 9.3005
R19933 gnd.n4475 gnd.n1372 9.3005
R19934 gnd.n4474 gnd.n4473 9.3005
R19935 gnd.n4472 gnd.n1373 9.3005
R19936 gnd.n4471 gnd.n4470 9.3005
R19937 gnd.n4469 gnd.n1377 9.3005
R19938 gnd.n4468 gnd.n4467 9.3005
R19939 gnd.n4466 gnd.n1378 9.3005
R19940 gnd.n4465 gnd.n4464 9.3005
R19941 gnd.n4463 gnd.n1382 9.3005
R19942 gnd.n4462 gnd.n4461 9.3005
R19943 gnd.n4460 gnd.n1383 9.3005
R19944 gnd.n4459 gnd.n4458 9.3005
R19945 gnd.n4457 gnd.n1387 9.3005
R19946 gnd.n4456 gnd.n4455 9.3005
R19947 gnd.n4454 gnd.n1388 9.3005
R19948 gnd.n4453 gnd.n4452 9.3005
R19949 gnd.n4451 gnd.n1392 9.3005
R19950 gnd.n4450 gnd.n4449 9.3005
R19951 gnd.n4448 gnd.n1393 9.3005
R19952 gnd.n4447 gnd.n4446 9.3005
R19953 gnd.n4445 gnd.n1397 9.3005
R19954 gnd.n4444 gnd.n4443 9.3005
R19955 gnd.n4442 gnd.n1398 9.3005
R19956 gnd.n4441 gnd.n4440 9.3005
R19957 gnd.n4439 gnd.n1402 9.3005
R19958 gnd.n4438 gnd.n4437 9.3005
R19959 gnd.n4436 gnd.n1403 9.3005
R19960 gnd.n4588 gnd.n4587 9.3005
R19961 gnd.n4345 gnd.n1502 9.3005
R19962 gnd.n4344 gnd.n4343 9.3005
R19963 gnd.n4342 gnd.n1504 9.3005
R19964 gnd.n4341 gnd.n4340 9.3005
R19965 gnd.n4339 gnd.n1508 9.3005
R19966 gnd.n4338 gnd.n4337 9.3005
R19967 gnd.n4336 gnd.n1509 9.3005
R19968 gnd.n4335 gnd.n4334 9.3005
R19969 gnd.n4333 gnd.n1513 9.3005
R19970 gnd.n4332 gnd.n4331 9.3005
R19971 gnd.n4330 gnd.n1514 9.3005
R19972 gnd.n4329 gnd.n4328 9.3005
R19973 gnd.n4327 gnd.n1518 9.3005
R19974 gnd.n4326 gnd.n4325 9.3005
R19975 gnd.n4324 gnd.n1519 9.3005
R19976 gnd.n4323 gnd.n4322 9.3005
R19977 gnd.n4321 gnd.n1523 9.3005
R19978 gnd.n4320 gnd.n4319 9.3005
R19979 gnd.n4318 gnd.n1524 9.3005
R19980 gnd.n4317 gnd.n4316 9.3005
R19981 gnd.n285 gnd.n283 9.3005
R19982 gnd.n7217 gnd.n7216 9.3005
R19983 gnd.n7215 gnd.n284 9.3005
R19984 gnd.n7214 gnd.n7213 9.3005
R19985 gnd.n7212 gnd.n286 9.3005
R19986 gnd.n7211 gnd.n7210 9.3005
R19987 gnd.n7208 gnd.n290 9.3005
R19988 gnd.n7207 gnd.n7206 9.3005
R19989 gnd.n7205 gnd.n292 9.3005
R19990 gnd.n261 gnd.n260 9.3005
R19991 gnd.n7229 gnd.n7228 9.3005
R19992 gnd.n7230 gnd.n259 9.3005
R19993 gnd.n7232 gnd.n7231 9.3005
R19994 gnd.n245 gnd.n244 9.3005
R19995 gnd.n7245 gnd.n7244 9.3005
R19996 gnd.n7246 gnd.n243 9.3005
R19997 gnd.n7248 gnd.n7247 9.3005
R19998 gnd.n230 gnd.n229 9.3005
R19999 gnd.n7261 gnd.n7260 9.3005
R20000 gnd.n7262 gnd.n228 9.3005
R20001 gnd.n7264 gnd.n7263 9.3005
R20002 gnd.n215 gnd.n214 9.3005
R20003 gnd.n7277 gnd.n7276 9.3005
R20004 gnd.n7278 gnd.n213 9.3005
R20005 gnd.n7280 gnd.n7279 9.3005
R20006 gnd.n200 gnd.n199 9.3005
R20007 gnd.n7293 gnd.n7292 9.3005
R20008 gnd.n7294 gnd.n197 9.3005
R20009 gnd.n7371 gnd.n7370 9.3005
R20010 gnd.n7369 gnd.n198 9.3005
R20011 gnd.n7368 gnd.n7367 9.3005
R20012 gnd.n7366 gnd.n7295 9.3005
R20013 gnd.n7365 gnd.n7364 9.3005
R20014 gnd.n4347 gnd.n4346 9.3005
R20015 gnd.n7361 gnd.n7297 9.3005
R20016 gnd.n7360 gnd.n7359 9.3005
R20017 gnd.n7358 gnd.n7302 9.3005
R20018 gnd.n7357 gnd.n7356 9.3005
R20019 gnd.n7355 gnd.n7303 9.3005
R20020 gnd.n7354 gnd.n7353 9.3005
R20021 gnd.n7352 gnd.n7310 9.3005
R20022 gnd.n7351 gnd.n7350 9.3005
R20023 gnd.n7349 gnd.n7311 9.3005
R20024 gnd.n7348 gnd.n7347 9.3005
R20025 gnd.n7346 gnd.n7318 9.3005
R20026 gnd.n7345 gnd.n7344 9.3005
R20027 gnd.n7343 gnd.n7319 9.3005
R20028 gnd.n7342 gnd.n7341 9.3005
R20029 gnd.n7340 gnd.n7326 9.3005
R20030 gnd.n7339 gnd.n7338 9.3005
R20031 gnd.n7337 gnd.n7327 9.3005
R20032 gnd.n7336 gnd.n7335 9.3005
R20033 gnd.n7363 gnd.n7362 9.3005
R20034 gnd.n4158 gnd.n1681 9.3005
R20035 gnd.n4161 gnd.n4160 9.3005
R20036 gnd.n4159 gnd.n1682 9.3005
R20037 gnd.n1613 gnd.n1612 9.3005
R20038 gnd.n4188 gnd.n4187 9.3005
R20039 gnd.n4189 gnd.n1610 9.3005
R20040 gnd.n4192 gnd.n4191 9.3005
R20041 gnd.n4190 gnd.n1611 9.3005
R20042 gnd.n1586 gnd.n1585 9.3005
R20043 gnd.n4219 gnd.n4218 9.3005
R20044 gnd.n4220 gnd.n1583 9.3005
R20045 gnd.n4228 gnd.n4227 9.3005
R20046 gnd.n4226 gnd.n1584 9.3005
R20047 gnd.n4225 gnd.n4224 9.3005
R20048 gnd.n4223 gnd.n4221 9.3005
R20049 gnd.n1551 gnd.n1549 9.3005
R20050 gnd.n4285 gnd.n4284 9.3005
R20051 gnd.n4283 gnd.n1550 9.3005
R20052 gnd.n4282 gnd.n4281 9.3005
R20053 gnd.n4280 gnd.n1552 9.3005
R20054 gnd.n4279 gnd.n4278 9.3005
R20055 gnd.n311 gnd.n310 9.3005
R20056 gnd.n7122 gnd.n7121 9.3005
R20057 gnd.n7123 gnd.n309 9.3005
R20058 gnd.n7125 gnd.n7124 9.3005
R20059 gnd.n69 gnd.n67 9.3005
R20060 gnd.n7502 gnd.n7501 9.3005
R20061 gnd.n7500 gnd.n68 9.3005
R20062 gnd.n7499 gnd.n7498 9.3005
R20063 gnd.n7497 gnd.n73 9.3005
R20064 gnd.n7496 gnd.n7495 9.3005
R20065 gnd.n7494 gnd.n74 9.3005
R20066 gnd.n7493 gnd.n7492 9.3005
R20067 gnd.n7491 gnd.n78 9.3005
R20068 gnd.n7490 gnd.n7489 9.3005
R20069 gnd.n7488 gnd.n79 9.3005
R20070 gnd.n7487 gnd.n7486 9.3005
R20071 gnd.n7485 gnd.n83 9.3005
R20072 gnd.n7484 gnd.n7483 9.3005
R20073 gnd.n7482 gnd.n84 9.3005
R20074 gnd.n7481 gnd.n7480 9.3005
R20075 gnd.n7479 gnd.n88 9.3005
R20076 gnd.n7478 gnd.n7477 9.3005
R20077 gnd.n7476 gnd.n89 9.3005
R20078 gnd.n7475 gnd.n7474 9.3005
R20079 gnd.n7473 gnd.n93 9.3005
R20080 gnd.n7472 gnd.n7471 9.3005
R20081 gnd.n7470 gnd.n94 9.3005
R20082 gnd.n7469 gnd.n7468 9.3005
R20083 gnd.n7467 gnd.n98 9.3005
R20084 gnd.n7466 gnd.n7465 9.3005
R20085 gnd.n7464 gnd.n99 9.3005
R20086 gnd.n7463 gnd.n102 9.3005
R20087 gnd.n4157 gnd.n4156 9.3005
R20088 gnd.n5730 gnd.t321 9.24152
R20089 gnd.n6244 gnd.t69 9.24152
R20090 gnd.t91 gnd.n922 9.24152
R20091 gnd.t73 gnd.n1015 9.24152
R20092 gnd.n2681 gnd.t175 9.24152
R20093 gnd.n4600 gnd.t87 9.24152
R20094 gnd.t327 gnd.n2067 9.24152
R20095 gnd.n4009 gnd.t43 9.24152
R20096 gnd.n3396 gnd.t43 9.24152
R20097 gnd.t99 gnd.n4163 9.24152
R20098 gnd.n4231 gnd.t192 9.24152
R20099 gnd.t41 gnd.t321 8.92286
R20100 gnd.t1 gnd.n3054 8.92286
R20101 gnd.n2025 gnd.t55 8.92286
R20102 gnd.n3443 gnd.t35 8.92286
R20103 gnd.n3969 gnd.t56 8.92286
R20104 gnd.n6080 gnd.n6055 8.92171
R20105 gnd.n6048 gnd.n6023 8.92171
R20106 gnd.n6016 gnd.n5991 8.92171
R20107 gnd.n5985 gnd.n5960 8.92171
R20108 gnd.n5953 gnd.n5928 8.92171
R20109 gnd.n5921 gnd.n5896 8.92171
R20110 gnd.n5889 gnd.n5864 8.92171
R20111 gnd.n5858 gnd.n5833 8.92171
R20112 gnd.n3194 gnd.n3176 8.72777
R20113 gnd.t307 gnd.n5036 8.60421
R20114 gnd.n2356 gnd.t194 8.60421
R20115 gnd.n3084 gnd.t10 8.60421
R20116 gnd.n3097 gnd.t47 8.60421
R20117 gnd.n1540 gnd.t208 8.60421
R20118 gnd.n5444 gnd.n5428 8.43467
R20119 gnd.n50 gnd.n34 8.43467
R20120 gnd.n2615 gnd.n0 8.41456
R20121 gnd.n7504 gnd.n7503 8.41456
R20122 gnd.n3841 gnd.n2066 8.28555
R20123 gnd.n3516 gnd.n3042 8.28555
R20124 gnd.n3495 gnd.n3494 8.28555
R20125 gnd.n3945 gnd.n1975 8.28555
R20126 gnd.n3977 gnd.n1945 8.28555
R20127 gnd.n3395 gnd.n3394 8.28555
R20128 gnd.n6081 gnd.n6053 8.14595
R20129 gnd.n6049 gnd.n6021 8.14595
R20130 gnd.n6017 gnd.n5989 8.14595
R20131 gnd.n5986 gnd.n5958 8.14595
R20132 gnd.n5954 gnd.n5926 8.14595
R20133 gnd.n5922 gnd.n5894 8.14595
R20134 gnd.n5890 gnd.n5862 8.14595
R20135 gnd.n5859 gnd.n5831 8.14595
R20136 gnd.n6086 gnd.n6085 7.97301
R20137 gnd.t313 gnd.n5078 7.9669
R20138 gnd.n2599 gnd.t186 7.9669
R20139 gnd.n3720 gnd.n2165 7.9669
R20140 gnd.n3004 gnd.t49 7.9669
R20141 gnd.t131 gnd.t59 7.9669
R20142 gnd.n1417 gnd.n1409 7.9669
R20143 gnd.n321 gnd.t206 7.9669
R20144 gnd.n7337 gnd.n7336 7.75808
R20145 gnd.n1800 gnd.n1799 7.75808
R20146 gnd.n3673 gnd.n2225 7.75808
R20147 gnd.n2482 gnd.n2479 7.75808
R20148 gnd.n3525 gnd.t8 7.64824
R20149 gnd.t324 gnd.n1939 7.64824
R20150 gnd.n186 gnd.t95 7.64824
R20151 gnd.n5560 gnd.t319 7.32958
R20152 gnd.t127 gnd.n2152 7.32958
R20153 gnd.n3769 gnd.t322 7.32958
R20154 gnd.t33 gnd.n1851 7.32958
R20155 gnd.n4126 gnd.t83 7.32958
R20156 gnd.n2913 gnd.n2912 7.30353
R20157 gnd.n3193 gnd.n3192 7.30353
R20158 gnd.n5520 gnd.n5153 7.01093
R20159 gnd.n5156 gnd.n5154 7.01093
R20160 gnd.n5530 gnd.n5529 7.01093
R20161 gnd.n5541 gnd.n5137 7.01093
R20162 gnd.n5540 gnd.n5140 7.01093
R20163 gnd.n5551 gnd.n5128 7.01093
R20164 gnd.n5131 gnd.n5129 7.01093
R20165 gnd.n5561 gnd.n5560 7.01093
R20166 gnd.n5572 gnd.n5111 7.01093
R20167 gnd.n5571 gnd.n5114 7.01093
R20168 gnd.n5582 gnd.n5104 7.01093
R20169 gnd.n5474 gnd.n5097 7.01093
R20170 gnd.n5603 gnd.n5086 7.01093
R20171 gnd.n5602 gnd.n5089 7.01093
R20172 gnd.n5613 gnd.n5078 7.01093
R20173 gnd.n5079 gnd.n5071 7.01093
R20174 gnd.n5634 gnd.n5060 7.01093
R20175 gnd.n5633 gnd.n5063 7.01093
R20176 gnd.n5053 gnd.n5046 7.01093
R20177 gnd.n5654 gnd.n5653 7.01093
R20178 gnd.n5664 gnd.n5036 7.01093
R20179 gnd.n5663 gnd.n5039 7.01093
R20180 gnd.n5674 gnd.n5029 7.01093
R20181 gnd.n5684 gnd.n5022 7.01093
R20182 gnd.n5708 gnd.n5016 7.01093
R20183 gnd.n5717 gnd.n5007 7.01093
R20184 gnd.n5726 gnd.n4999 7.01093
R20185 gnd.n5730 gnd.n5729 7.01093
R20186 gnd.n5748 gnd.n4984 7.01093
R20187 gnd.n5747 gnd.n4987 7.01093
R20188 gnd.n5758 gnd.n4976 7.01093
R20189 gnd.n4977 gnd.n4966 7.01093
R20190 gnd.n5793 gnd.n5792 7.01093
R20191 gnd.n5805 gnd.n5804 7.01093
R20192 gnd.n4953 gnd.n4945 7.01093
R20193 gnd.n5816 gnd.n5815 7.01093
R20194 gnd.n6115 gnd.n4930 7.01093
R20195 gnd.n6114 gnd.n4933 7.01093
R20196 gnd.n6130 gnd.n896 7.01093
R20197 gnd.n6257 gnd.n898 7.01093
R20198 gnd.n6136 gnd.n907 7.01093
R20199 gnd.n6251 gnd.n6250 7.01093
R20200 gnd.n6099 gnd.n910 7.01093
R20201 gnd.n6244 gnd.n919 7.01093
R20202 gnd.n6243 gnd.n922 7.01093
R20203 gnd.n6147 gnd.n930 7.01093
R20204 gnd.n6237 gnd.n6236 7.01093
R20205 gnd.t120 gnd.n2073 7.01093
R20206 gnd.n3545 gnd.t4 7.01093
R20207 gnd.n3849 gnd.n2058 7.01093
R20208 gnd.n3524 gnd.n3523 7.01093
R20209 gnd.n3487 gnd.n3082 7.01093
R20210 gnd.n3937 gnd.n1981 7.01093
R20211 gnd.n3985 gnd.n1938 7.01093
R20212 gnd.n3156 gnd.n3154 7.01093
R20213 gnd.t20 gnd.n1918 7.01093
R20214 gnd.n3387 gnd.t113 7.01093
R20215 gnd.n5114 gnd.t317 6.69227
R20216 gnd.n5726 gnd.t41 6.69227
R20217 gnd.n6129 gnd.t312 6.69227
R20218 gnd.n6258 gnd.n896 6.69227
R20219 gnd.n4727 gnd.t269 6.69227
R20220 gnd.n2694 gnd.t184 6.69227
R20221 gnd.n1601 gnd.t222 6.69227
R20222 gnd.t214 gnd.n208 6.69227
R20223 gnd.n3310 gnd.n3309 6.5566
R20224 gnd.n3633 gnd.n3632 6.5566
R20225 gnd.n2937 gnd.n2931 6.5566
R20226 gnd.n3325 gnd.n3324 6.5566
R20227 gnd.n3015 gnd.t146 6.37362
R20228 gnd.t67 gnd.n2009 6.37362
R20229 gnd.n3457 gnd.t7 6.37362
R20230 gnd.n2803 gnd.n2798 6.20656
R20231 gnd.n7426 gnd.n7423 6.20656
R20232 gnd.n4796 gnd.n4795 6.20656
R20233 gnd.n4145 gnd.n4142 6.20656
R20234 gnd.t63 gnd.n5622 6.05496
R20235 gnd.n5623 gnd.t316 6.05496
R20236 gnd.t329 gnd.n5663 6.05496
R20237 gnd.n5762 gnd.t315 6.05496
R20238 gnd.n4703 gnd.t198 6.05496
R20239 gnd.n2669 gnd.t196 6.05496
R20240 gnd.t10 gnd.n3082 6.05496
R20241 gnd.n3937 gnd.t47 6.05496
R20242 gnd.n4288 gnd.t233 6.05496
R20243 gnd.t235 gnd.n238 6.05496
R20244 gnd.n6083 gnd.n6053 5.81868
R20245 gnd.n6051 gnd.n6021 5.81868
R20246 gnd.n6019 gnd.n5989 5.81868
R20247 gnd.n5988 gnd.n5958 5.81868
R20248 gnd.n5956 gnd.n5926 5.81868
R20249 gnd.n5924 gnd.n5894 5.81868
R20250 gnd.n5892 gnd.n5862 5.81868
R20251 gnd.n5861 gnd.n5831 5.81868
R20252 gnd.n3825 gnd.t140 5.73631
R20253 gnd.n3857 gnd.n2051 5.73631
R20254 gnd.n3531 gnd.n3029 5.73631
R20255 gnd.n3480 gnd.n3479 5.73631
R20256 gnd.n3929 gnd.n1989 5.73631
R20257 gnd.n3993 gnd.n1931 5.73631
R20258 gnd.n3410 gnd.n3409 5.73631
R20259 gnd.n3221 gnd.n1466 5.62001
R20260 gnd.n3640 gnd.n2870 5.62001
R20261 gnd.n3640 gnd.n2871 5.62001
R20262 gnd.n3319 gnd.n1466 5.62001
R20263 gnd.n5293 gnd.n5288 5.4308
R20264 gnd.n4911 gnd.n4909 5.4308
R20265 gnd.n5674 gnd.t314 5.41765
R20266 gnd.n5718 gnd.t306 5.41765
R20267 gnd.n5794 gnd.t57 5.41765
R20268 gnd.n1098 gnd.n1097 5.41765
R20269 gnd.n4679 gnd.t186 5.41765
R20270 gnd.n2612 gnd.t253 5.41765
R20271 gnd.n2093 gnd.n2086 5.41765
R20272 gnd.n7127 gnd.t257 5.41765
R20273 gnd.n7198 gnd.t206 5.41765
R20274 gnd.n7242 gnd.n250 5.41765
R20275 gnd.n3817 gnd.t80 5.09899
R20276 gnd.n3565 gnd.t140 5.09899
R20277 gnd.n6081 gnd.n6080 5.04292
R20278 gnd.n6049 gnd.n6048 5.04292
R20279 gnd.n6017 gnd.n6016 5.04292
R20280 gnd.n5986 gnd.n5985 5.04292
R20281 gnd.n5954 gnd.n5953 5.04292
R20282 gnd.n5922 gnd.n5921 5.04292
R20283 gnd.n5890 gnd.n5889 5.04292
R20284 gnd.n5859 gnd.n5858 5.04292
R20285 gnd.n5460 gnd.n5459 4.82753
R20286 gnd.n66 gnd.n65 4.82753
R20287 gnd.n5644 gnd.t309 4.78034
R20288 gnd.n4987 gnd.t310 4.78034
R20289 gnd.n2577 gnd.t190 4.78034
R20290 gnd.n4654 gnd.t194 4.78034
R20291 gnd.t12 gnd.n2107 4.78034
R20292 gnd.n3531 gnd.t52 4.78034
R20293 gnd.t303 gnd.n1931 4.78034
R20294 gnd.n3196 gnd.t134 4.78034
R20295 gnd.n4065 gnd.t45 4.78034
R20296 gnd.n4314 gnd.t208 4.78034
R20297 gnd.n7234 gnd.t177 4.78034
R20298 gnd.n5464 gnd.n5463 4.74817
R20299 gnd.n5413 gnd.n5411 4.74817
R20300 gnd.n5406 gnd.n5405 4.74817
R20301 gnd.n5402 gnd.n5401 4.74817
R20302 gnd.n5463 gnd.n5400 4.74817
R20303 gnd.n5413 gnd.n5412 4.74817
R20304 gnd.n5407 gnd.n5406 4.74817
R20305 gnd.n5404 gnd.n5402 4.74817
R20306 gnd.n7222 gnd.n7221 4.74817
R20307 gnd.n7130 gnd.n272 4.74817
R20308 gnd.n7200 gnd.n271 4.74817
R20309 gnd.n270 gnd.n267 4.74817
R20310 gnd.n7222 gnd.n274 4.74817
R20311 gnd.n306 gnd.n272 4.74817
R20312 gnd.n7129 gnd.n271 4.74817
R20313 gnd.n7201 gnd.n270 4.74817
R20314 gnd.n2392 gnd.n2389 4.74817
R20315 gnd.n2597 gnd.n2388 4.74817
R20316 gnd.n2593 gnd.n2387 4.74817
R20317 gnd.n2386 gnd.n2366 4.74817
R20318 gnd.n2640 gnd.n2367 4.74817
R20319 gnd.n4297 gnd.n317 4.74817
R20320 gnd.n7115 gnd.n7114 4.74817
R20321 gnd.n7110 gnd.n318 4.74817
R20322 gnd.n7108 gnd.n7107 4.74817
R20323 gnd.n7103 gnd.n325 4.74817
R20324 gnd.n4298 gnd.n4297 4.74817
R20325 gnd.n7116 gnd.n7115 4.74817
R20326 gnd.n7113 gnd.n318 4.74817
R20327 gnd.n7109 gnd.n7108 4.74817
R20328 gnd.n325 gnd.n323 4.74817
R20329 gnd.n1124 gnd.n1107 4.74817
R20330 gnd.n1143 gnd.n1126 4.74817
R20331 gnd.n4670 gnd.n4669 4.74817
R20332 gnd.n1161 gnd.n1144 4.74817
R20333 gnd.n4683 gnd.n1124 4.74817
R20334 gnd.n4681 gnd.n1126 4.74817
R20335 gnd.n4671 gnd.n4670 4.74817
R20336 gnd.n4668 gnd.n1144 4.74817
R20337 gnd.n2588 gnd.n2389 4.74817
R20338 gnd.n2589 gnd.n2388 4.74817
R20339 gnd.n2596 gnd.n2387 4.74817
R20340 gnd.n2592 gnd.n2386 4.74817
R20341 gnd.n2641 gnd.n2640 4.74817
R20342 gnd.n5444 gnd.n5443 4.7074
R20343 gnd.n50 gnd.n49 4.7074
R20344 gnd.n5460 gnd.n5444 4.65959
R20345 gnd.n66 gnd.n50 4.65959
R20346 gnd.n4393 gnd.n1468 4.6132
R20347 gnd.n3641 gnd.n2869 4.6132
R20348 gnd.n3571 gnd.t80 4.46168
R20349 gnd.n3538 gnd.n3022 4.46168
R20350 gnd.t23 gnd.n2052 4.46168
R20351 gnd.n3865 gnd.n2044 4.46168
R20352 gnd.n3921 gnd.n1995 4.46168
R20353 gnd.n3472 gnd.n3095 4.46168
R20354 gnd.n3417 gnd.n3141 4.46168
R20355 gnd.n3411 gnd.t18 4.46168
R20356 gnd.n4001 gnd.n1925 4.46168
R20357 gnd.n3189 gnd.n3176 4.46111
R20358 gnd.n6066 gnd.n6062 4.38594
R20359 gnd.n6034 gnd.n6030 4.38594
R20360 gnd.n6002 gnd.n5998 4.38594
R20361 gnd.n5971 gnd.n5967 4.38594
R20362 gnd.n5939 gnd.n5935 4.38594
R20363 gnd.n5907 gnd.n5903 4.38594
R20364 gnd.n5875 gnd.n5871 4.38594
R20365 gnd.n5844 gnd.n5840 4.38594
R20366 gnd.n6077 gnd.n6055 4.26717
R20367 gnd.n6045 gnd.n6023 4.26717
R20368 gnd.n6013 gnd.n5991 4.26717
R20369 gnd.n5982 gnd.n5960 4.26717
R20370 gnd.n5950 gnd.n5928 4.26717
R20371 gnd.n5918 gnd.n5896 4.26717
R20372 gnd.n5886 gnd.n5864 4.26717
R20373 gnd.n5855 gnd.n5833 4.26717
R20374 gnd.n5592 gnd.t311 4.14303
R20375 gnd.n5815 gnd.t308 4.14303
R20376 gnd.n1067 gnd.t179 4.14303
R20377 gnd.n4630 gnd.t175 4.14303
R20378 gnd.n2316 gnd.t87 4.14303
R20379 gnd.n4164 gnd.t99 4.14303
R20380 gnd.t192 gnd.n4230 4.14303
R20381 gnd.n7266 gnd.t218 4.14303
R20382 gnd.n6085 gnd.n6084 4.08274
R20383 gnd.n3309 gnd.n3308 4.05904
R20384 gnd.n3632 gnd.n3631 4.05904
R20385 gnd.n2941 gnd.n2931 4.05904
R20386 gnd.n3326 gnd.n3325 4.05904
R20387 gnd.n19 gnd.n9 3.99943
R20388 gnd.n3084 gnd.t40 3.82437
R20389 gnd.n3097 gnd.t0 3.82437
R20390 gnd.n6085 gnd.n5957 3.70378
R20391 gnd.n5462 gnd.n5461 3.65935
R20392 gnd.n19 gnd.n18 3.60163
R20393 gnd.n6076 gnd.n6057 3.49141
R20394 gnd.n6044 gnd.n6025 3.49141
R20395 gnd.n6012 gnd.n5993 3.49141
R20396 gnd.n5981 gnd.n5962 3.49141
R20397 gnd.n5949 gnd.n5930 3.49141
R20398 gnd.n5917 gnd.n5898 3.49141
R20399 gnd.n5885 gnd.n5866 3.49141
R20400 gnd.n5854 gnd.n5835 3.49141
R20401 gnd.n3545 gnd.n3015 3.18706
R20402 gnd.n3074 gnd.t9 3.18706
R20403 gnd.n3913 gnd.n2002 3.18706
R20404 gnd.n3465 gnd.n3464 3.18706
R20405 gnd.t32 gnd.n1967 3.18706
R20406 gnd.n4009 gnd.n1918 3.18706
R20407 gnd.t311 gnd.n5591 2.8684
R20408 gnd.n2634 gnd.t181 2.8684
R20409 gnd.n3825 gnd.t49 2.8684
R20410 gnd.t146 gnd.t327 2.8684
R20411 gnd.t59 gnd.n1905 2.8684
R20412 gnd.t188 gnd.n263 2.8684
R20413 gnd.n5445 gnd.t176 2.82907
R20414 gnd.n5445 gnd.t262 2.82907
R20415 gnd.n5447 gnd.t286 2.82907
R20416 gnd.n5447 gnd.t243 2.82907
R20417 gnd.n5449 gnd.t268 2.82907
R20418 gnd.n5449 gnd.t216 2.82907
R20419 gnd.n5451 gnd.t248 2.82907
R20420 gnd.n5451 gnd.t285 2.82907
R20421 gnd.n5453 gnd.t295 2.82907
R20422 gnd.n5453 gnd.t288 2.82907
R20423 gnd.n5455 gnd.t287 2.82907
R20424 gnd.n5455 gnd.t278 2.82907
R20425 gnd.n5457 gnd.t290 2.82907
R20426 gnd.n5457 gnd.t200 2.82907
R20427 gnd.n5414 gnd.t183 2.82907
R20428 gnd.n5414 gnd.t212 2.82907
R20429 gnd.n5416 gnd.t226 2.82907
R20430 gnd.n5416 gnd.t256 2.82907
R20431 gnd.n5418 gnd.t300 2.82907
R20432 gnd.n5418 gnd.t195 2.82907
R20433 gnd.n5420 gnd.t213 2.82907
R20434 gnd.n5420 gnd.t274 2.82907
R20435 gnd.n5422 gnd.t191 2.82907
R20436 gnd.n5422 gnd.t182 2.82907
R20437 gnd.n5424 gnd.t237 2.82907
R20438 gnd.n5424 gnd.t227 2.82907
R20439 gnd.n5426 gnd.t282 2.82907
R20440 gnd.n5426 gnd.t205 2.82907
R20441 gnd.n5429 gnd.t294 2.82907
R20442 gnd.n5429 gnd.t185 2.82907
R20443 gnd.n5431 gnd.t197 2.82907
R20444 gnd.n5431 gnd.t229 2.82907
R20445 gnd.n5433 gnd.t284 2.82907
R20446 gnd.n5433 gnd.t302 2.82907
R20447 gnd.n5435 gnd.t187 2.82907
R20448 gnd.n5435 gnd.t254 2.82907
R20449 gnd.n5437 gnd.t298 2.82907
R20450 gnd.n5437 gnd.t293 2.82907
R20451 gnd.n5439 gnd.t211 2.82907
R20452 gnd.n5439 gnd.t199 2.82907
R20453 gnd.n5441 gnd.t270 2.82907
R20454 gnd.n5441 gnd.t180 2.82907
R20455 gnd.n63 gnd.t296 2.82907
R20456 gnd.n63 gnd.t215 2.82907
R20457 gnd.n61 gnd.t242 2.82907
R20458 gnd.n61 gnd.t260 2.82907
R20459 gnd.n59 gnd.t261 2.82907
R20460 gnd.n59 gnd.t283 2.82907
R20461 gnd.n57 gnd.t258 2.82907
R20462 gnd.n57 gnd.t207 2.82907
R20463 gnd.n55 gnd.t301 2.82907
R20464 gnd.n55 gnd.t240 2.82907
R20465 gnd.n53 gnd.t202 2.82907
R20466 gnd.n53 gnd.t259 2.82907
R20467 gnd.n51 gnd.t223 2.82907
R20468 gnd.n51 gnd.t277 2.82907
R20469 gnd.n32 gnd.t241 2.82907
R20470 gnd.n32 gnd.t276 2.82907
R20471 gnd.n30 gnd.t264 2.82907
R20472 gnd.n30 gnd.t271 2.82907
R20473 gnd.n28 gnd.t220 2.82907
R20474 gnd.n28 gnd.t178 2.82907
R20475 gnd.n26 gnd.t297 2.82907
R20476 gnd.n26 gnd.t247 2.82907
R20477 gnd.n24 gnd.t232 2.82907
R20478 gnd.n24 gnd.t291 2.82907
R20479 gnd.n22 gnd.t281 2.82907
R20480 gnd.n22 gnd.t263 2.82907
R20481 gnd.n20 gnd.t246 2.82907
R20482 gnd.n20 gnd.t221 2.82907
R20483 gnd.n47 gnd.t219 2.82907
R20484 gnd.n47 gnd.t255 2.82907
R20485 gnd.n45 gnd.t236 2.82907
R20486 gnd.n45 gnd.t245 2.82907
R20487 gnd.n43 gnd.t189 2.82907
R20488 gnd.n43 gnd.t289 2.82907
R20489 gnd.n41 gnd.t279 2.82907
R20490 gnd.n41 gnd.t225 2.82907
R20491 gnd.n39 gnd.t209 2.82907
R20492 gnd.n39 gnd.t273 2.82907
R20493 gnd.n37 gnd.t266 2.82907
R20494 gnd.n37 gnd.t234 2.82907
R20495 gnd.n35 gnd.t224 2.82907
R20496 gnd.n35 gnd.t193 2.82907
R20497 gnd.n6073 gnd.n6072 2.71565
R20498 gnd.n6041 gnd.n6040 2.71565
R20499 gnd.n6009 gnd.n6008 2.71565
R20500 gnd.n5978 gnd.n5977 2.71565
R20501 gnd.n5946 gnd.n5945 2.71565
R20502 gnd.n5914 gnd.n5913 2.71565
R20503 gnd.n5882 gnd.n5881 2.71565
R20504 gnd.n5851 gnd.n5850 2.71565
R20505 gnd.n3552 gnd.t124 2.54975
R20506 gnd.n3913 gnd.t5 2.54975
R20507 gnd.n3464 gnd.t66 2.54975
R20508 gnd.n3394 gnd.t117 2.54975
R20509 gnd.n5463 gnd.n5462 2.27742
R20510 gnd.n5462 gnd.n5413 2.27742
R20511 gnd.n5462 gnd.n5406 2.27742
R20512 gnd.n5462 gnd.n5402 2.27742
R20513 gnd.n7223 gnd.n7222 2.27742
R20514 gnd.n7223 gnd.n272 2.27742
R20515 gnd.n7223 gnd.n271 2.27742
R20516 gnd.n7223 gnd.n270 2.27742
R20517 gnd.n4297 gnd.n269 2.27742
R20518 gnd.n7115 gnd.n269 2.27742
R20519 gnd.n318 gnd.n269 2.27742
R20520 gnd.n7108 gnd.n269 2.27742
R20521 gnd.n325 gnd.n269 2.27742
R20522 gnd.n1125 gnd.n1124 2.27742
R20523 gnd.n1126 gnd.n1125 2.27742
R20524 gnd.n4670 gnd.n1125 2.27742
R20525 gnd.n1144 gnd.n1125 2.27742
R20526 gnd.n2639 gnd.n2389 2.27742
R20527 gnd.n2639 gnd.n2388 2.27742
R20528 gnd.n2639 gnd.n2387 2.27742
R20529 gnd.n2639 gnd.n2386 2.27742
R20530 gnd.n2640 gnd.n2639 2.27742
R20531 gnd.n5529 gnd.t149 2.23109
R20532 gnd.n5409 gnd.t309 2.23109
R20533 gnd.n2643 gnd.t267 2.23109
R20534 gnd.n312 gnd.t239 2.23109
R20535 gnd.n6069 gnd.n6059 1.93989
R20536 gnd.n6037 gnd.n6027 1.93989
R20537 gnd.n6005 gnd.n5995 1.93989
R20538 gnd.n5974 gnd.n5964 1.93989
R20539 gnd.n5942 gnd.n5932 1.93989
R20540 gnd.n5910 gnd.n5900 1.93989
R20541 gnd.n5878 gnd.n5868 1.93989
R20542 gnd.n5847 gnd.n5837 1.93989
R20543 gnd.n3552 gnd.n3009 1.91244
R20544 gnd.n3522 gnd.t19 1.91244
R20545 gnd.t55 gnd.n2024 1.91244
R20546 gnd.n3905 gnd.n2009 1.91244
R20547 gnd.n3457 gnd.n3109 1.91244
R20548 gnd.n3961 gnd.t35 1.91244
R20549 gnd.n3424 gnd.t65 1.91244
R20550 gnd.n4017 gnd.n1911 1.91244
R20551 gnd.t325 gnd.n5540 1.59378
R20552 gnd.n5707 gnd.t306 1.59378
R20553 gnd.n5761 gnd.t57 1.59378
R20554 gnd.n2709 gnd.t228 1.59378
R20555 gnd.n3881 gnd.t38 1.59378
R20556 gnd.t2 gnd.n3131 1.59378
R20557 gnd.t201 gnd.n1561 1.59378
R20558 gnd.n7381 gnd.n186 1.59378
R20559 gnd.n3873 gnd.t19 1.27512
R20560 gnd.t65 gnd.n3135 1.27512
R20561 gnd.n5296 gnd.n5288 1.16414
R20562 gnd.n6162 gnd.n4909 1.16414
R20563 gnd.n6068 gnd.n6061 1.16414
R20564 gnd.n6036 gnd.n6029 1.16414
R20565 gnd.n6004 gnd.n5997 1.16414
R20566 gnd.n5973 gnd.n5966 1.16414
R20567 gnd.n5941 gnd.n5934 1.16414
R20568 gnd.n5909 gnd.n5902 1.16414
R20569 gnd.n5877 gnd.n5870 1.16414
R20570 gnd.n5846 gnd.n5839 1.16414
R20571 gnd.n4393 gnd.n4392 0.970197
R20572 gnd.n3641 gnd.n2289 0.970197
R20573 gnd.n6052 gnd.n6020 0.962709
R20574 gnd.n6084 gnd.n6052 0.962709
R20575 gnd.n5925 gnd.n5893 0.962709
R20576 gnd.n5957 gnd.n5925 0.962709
R20577 gnd.n5623 gnd.t63 0.956468
R20578 gnd.n5771 gnd.t315 0.956468
R20579 gnd.n2763 gnd.t203 0.956468
R20580 gnd.t9 gnd.t24 0.956468
R20581 gnd.t30 gnd.t32 0.956468
R20582 gnd.n4195 gnd.t249 0.956468
R20583 gnd.n5454 gnd.n5452 0.773756
R20584 gnd.n60 gnd.n58 0.773756
R20585 gnd.n5459 gnd.n5458 0.773756
R20586 gnd.n5458 gnd.n5456 0.773756
R20587 gnd.n5456 gnd.n5454 0.773756
R20588 gnd.n5452 gnd.n5450 0.773756
R20589 gnd.n5450 gnd.n5448 0.773756
R20590 gnd.n5448 gnd.n5446 0.773756
R20591 gnd.n54 gnd.n52 0.773756
R20592 gnd.n56 gnd.n54 0.773756
R20593 gnd.n58 gnd.n56 0.773756
R20594 gnd.n62 gnd.n60 0.773756
R20595 gnd.n64 gnd.n62 0.773756
R20596 gnd.n65 gnd.n64 0.773756
R20597 gnd.n2 gnd.n1 0.672012
R20598 gnd.n3 gnd.n2 0.672012
R20599 gnd.n4 gnd.n3 0.672012
R20600 gnd.n5 gnd.n4 0.672012
R20601 gnd.n6 gnd.n5 0.672012
R20602 gnd.n7 gnd.n6 0.672012
R20603 gnd.n8 gnd.n7 0.672012
R20604 gnd.n9 gnd.n8 0.672012
R20605 gnd.n11 gnd.n10 0.672012
R20606 gnd.n12 gnd.n11 0.672012
R20607 gnd.n13 gnd.n12 0.672012
R20608 gnd.n14 gnd.n13 0.672012
R20609 gnd.n15 gnd.n14 0.672012
R20610 gnd.n16 gnd.n15 0.672012
R20611 gnd.n17 gnd.n16 0.672012
R20612 gnd.n18 gnd.n17 0.672012
R20613 gnd gnd.n0 0.665707
R20614 gnd.n2999 gnd.n2892 0.637812
R20615 gnd.n3559 gnd.n3005 0.637812
R20616 gnd.n3022 gnd.t54 0.637812
R20617 gnd.n3509 gnd.t1 0.637812
R20618 gnd.n3889 gnd.n2023 0.637812
R20619 gnd.n3897 gnd.n2017 0.637812
R20620 gnd.n3450 gnd.n3449 0.637812
R20621 gnd.n3127 gnd.n3122 0.637812
R20622 gnd.n3437 gnd.t56 0.637812
R20623 gnd.n4001 gnd.t6 0.637812
R20624 gnd.n4025 gnd.n1903 0.637812
R20625 gnd.n4033 gnd.n1897 0.637812
R20626 gnd.n4041 gnd.t134 0.637812
R20627 gnd.n5428 gnd.n5427 0.573776
R20628 gnd.n5427 gnd.n5425 0.573776
R20629 gnd.n5425 gnd.n5423 0.573776
R20630 gnd.n5423 gnd.n5421 0.573776
R20631 gnd.n5421 gnd.n5419 0.573776
R20632 gnd.n5419 gnd.n5417 0.573776
R20633 gnd.n5417 gnd.n5415 0.573776
R20634 gnd.n5443 gnd.n5442 0.573776
R20635 gnd.n5442 gnd.n5440 0.573776
R20636 gnd.n5440 gnd.n5438 0.573776
R20637 gnd.n5438 gnd.n5436 0.573776
R20638 gnd.n5436 gnd.n5434 0.573776
R20639 gnd.n5434 gnd.n5432 0.573776
R20640 gnd.n5432 gnd.n5430 0.573776
R20641 gnd.n23 gnd.n21 0.573776
R20642 gnd.n25 gnd.n23 0.573776
R20643 gnd.n27 gnd.n25 0.573776
R20644 gnd.n29 gnd.n27 0.573776
R20645 gnd.n31 gnd.n29 0.573776
R20646 gnd.n33 gnd.n31 0.573776
R20647 gnd.n34 gnd.n33 0.573776
R20648 gnd.n38 gnd.n36 0.573776
R20649 gnd.n40 gnd.n38 0.573776
R20650 gnd.n42 gnd.n40 0.573776
R20651 gnd.n44 gnd.n42 0.573776
R20652 gnd.n46 gnd.n44 0.573776
R20653 gnd.n48 gnd.n46 0.573776
R20654 gnd.n49 gnd.n48 0.573776
R20655 gnd.n7505 gnd.n7504 0.553847
R20656 gnd.n7223 gnd.n269 0.548625
R20657 gnd.n2639 gnd.n1125 0.548625
R20658 gnd.n2483 gnd.n2481 0.505073
R20659 gnd.n2521 gnd.n2520 0.505073
R20660 gnd.n7364 gnd.n7363 0.505073
R20661 gnd.n7335 gnd.n102 0.505073
R20662 gnd.n7458 gnd.n7457 0.492878
R20663 gnd.n7387 gnd.n7386 0.492878
R20664 gnd.n4353 gnd.n1494 0.492878
R20665 gnd.n1643 gnd.n1450 0.492878
R20666 gnd.n2273 gnd.n1268 0.492878
R20667 gnd.n2826 gnd.n2825 0.492878
R20668 gnd.n4756 gnd.n1008 0.492878
R20669 gnd.n2530 gnd.n965 0.492878
R20670 gnd.n6152 gnd.n6151 0.486781
R20671 gnd.n1723 gnd.n1403 0.486781
R20672 gnd.n5345 gnd.n5344 0.48678
R20673 gnd.n4589 gnd.n4588 0.485256
R20674 gnd.n6233 gnd.n6232 0.480683
R20675 gnd.n5515 gnd.n5514 0.480683
R20676 gnd.n4132 gnd.n4131 0.451719
R20677 gnd.n3725 gnd.n3724 0.451719
R20678 gnd.n6430 gnd.n726 0.425805
R20679 gnd.n6883 gnd.n6882 0.425805
R20680 gnd.n7095 gnd.n7094 0.425805
R20681 gnd.n2394 gnd.n2393 0.425805
R20682 gnd.n4591 gnd.n4590 0.406268
R20683 gnd.n4346 gnd.n1503 0.404992
R20684 gnd.n2806 gnd.n2798 0.388379
R20685 gnd.n6065 gnd.n6064 0.388379
R20686 gnd.n6033 gnd.n6032 0.388379
R20687 gnd.n6001 gnd.n6000 0.388379
R20688 gnd.n5970 gnd.n5969 0.388379
R20689 gnd.n5938 gnd.n5937 0.388379
R20690 gnd.n5906 gnd.n5905 0.388379
R20691 gnd.n5874 gnd.n5873 0.388379
R20692 gnd.n5843 gnd.n5842 0.388379
R20693 gnd.n7427 gnd.n7426 0.388379
R20694 gnd.n4797 gnd.n4796 0.388379
R20695 gnd.n4146 gnd.n4145 0.388379
R20696 gnd.n7505 gnd.n19 0.374463
R20697 gnd gnd.n7505 0.367492
R20698 gnd.n4935 gnd.t312 0.319156
R20699 gnd.n3515 gnd.t38 0.319156
R20700 gnd.n3431 gnd.t2 0.319156
R20701 gnd.n5263 gnd.n5241 0.311721
R20702 gnd.n2817 gnd.n2816 0.27489
R20703 gnd.n4157 gnd.n4155 0.27489
R20704 gnd.n6202 gnd.n6201 0.268793
R20705 gnd.n6201 gnd.n6200 0.241354
R20706 gnd.n1468 gnd.n1465 0.229039
R20707 gnd.n1471 gnd.n1468 0.229039
R20708 gnd.n2869 gnd.n2288 0.229039
R20709 gnd.n2869 gnd.n2868 0.229039
R20710 gnd.n5503 gnd.n5216 0.206293
R20711 gnd.n5461 gnd.n0 0.169152
R20712 gnd.n6082 gnd.n6054 0.155672
R20713 gnd.n6075 gnd.n6054 0.155672
R20714 gnd.n6075 gnd.n6074 0.155672
R20715 gnd.n6074 gnd.n6058 0.155672
R20716 gnd.n6067 gnd.n6058 0.155672
R20717 gnd.n6067 gnd.n6066 0.155672
R20718 gnd.n6050 gnd.n6022 0.155672
R20719 gnd.n6043 gnd.n6022 0.155672
R20720 gnd.n6043 gnd.n6042 0.155672
R20721 gnd.n6042 gnd.n6026 0.155672
R20722 gnd.n6035 gnd.n6026 0.155672
R20723 gnd.n6035 gnd.n6034 0.155672
R20724 gnd.n6018 gnd.n5990 0.155672
R20725 gnd.n6011 gnd.n5990 0.155672
R20726 gnd.n6011 gnd.n6010 0.155672
R20727 gnd.n6010 gnd.n5994 0.155672
R20728 gnd.n6003 gnd.n5994 0.155672
R20729 gnd.n6003 gnd.n6002 0.155672
R20730 gnd.n5987 gnd.n5959 0.155672
R20731 gnd.n5980 gnd.n5959 0.155672
R20732 gnd.n5980 gnd.n5979 0.155672
R20733 gnd.n5979 gnd.n5963 0.155672
R20734 gnd.n5972 gnd.n5963 0.155672
R20735 gnd.n5972 gnd.n5971 0.155672
R20736 gnd.n5955 gnd.n5927 0.155672
R20737 gnd.n5948 gnd.n5927 0.155672
R20738 gnd.n5948 gnd.n5947 0.155672
R20739 gnd.n5947 gnd.n5931 0.155672
R20740 gnd.n5940 gnd.n5931 0.155672
R20741 gnd.n5940 gnd.n5939 0.155672
R20742 gnd.n5923 gnd.n5895 0.155672
R20743 gnd.n5916 gnd.n5895 0.155672
R20744 gnd.n5916 gnd.n5915 0.155672
R20745 gnd.n5915 gnd.n5899 0.155672
R20746 gnd.n5908 gnd.n5899 0.155672
R20747 gnd.n5908 gnd.n5907 0.155672
R20748 gnd.n5891 gnd.n5863 0.155672
R20749 gnd.n5884 gnd.n5863 0.155672
R20750 gnd.n5884 gnd.n5883 0.155672
R20751 gnd.n5883 gnd.n5867 0.155672
R20752 gnd.n5876 gnd.n5867 0.155672
R20753 gnd.n5876 gnd.n5875 0.155672
R20754 gnd.n5860 gnd.n5832 0.155672
R20755 gnd.n5853 gnd.n5832 0.155672
R20756 gnd.n5853 gnd.n5852 0.155672
R20757 gnd.n5852 gnd.n5836 0.155672
R20758 gnd.n5845 gnd.n5836 0.155672
R20759 gnd.n5845 gnd.n5844 0.155672
R20760 gnd.n6232 gnd.n4839 0.152939
R20761 gnd.n4841 gnd.n4839 0.152939
R20762 gnd.n4845 gnd.n4841 0.152939
R20763 gnd.n4846 gnd.n4845 0.152939
R20764 gnd.n4847 gnd.n4846 0.152939
R20765 gnd.n4848 gnd.n4847 0.152939
R20766 gnd.n4852 gnd.n4848 0.152939
R20767 gnd.n4853 gnd.n4852 0.152939
R20768 gnd.n4854 gnd.n4853 0.152939
R20769 gnd.n4855 gnd.n4854 0.152939
R20770 gnd.n4859 gnd.n4855 0.152939
R20771 gnd.n4860 gnd.n4859 0.152939
R20772 gnd.n4861 gnd.n4860 0.152939
R20773 gnd.n4862 gnd.n4861 0.152939
R20774 gnd.n4867 gnd.n4862 0.152939
R20775 gnd.n6202 gnd.n4867 0.152939
R20776 gnd.n5516 gnd.n5515 0.152939
R20777 gnd.n5516 gnd.n5134 0.152939
R20778 gnd.n5544 gnd.n5134 0.152939
R20779 gnd.n5545 gnd.n5544 0.152939
R20780 gnd.n5546 gnd.n5545 0.152939
R20781 gnd.n5547 gnd.n5546 0.152939
R20782 gnd.n5547 gnd.n5108 0.152939
R20783 gnd.n5575 gnd.n5108 0.152939
R20784 gnd.n5576 gnd.n5575 0.152939
R20785 gnd.n5577 gnd.n5576 0.152939
R20786 gnd.n5578 gnd.n5577 0.152939
R20787 gnd.n5578 gnd.n5083 0.152939
R20788 gnd.n5606 gnd.n5083 0.152939
R20789 gnd.n5607 gnd.n5606 0.152939
R20790 gnd.n5608 gnd.n5607 0.152939
R20791 gnd.n5609 gnd.n5608 0.152939
R20792 gnd.n5609 gnd.n5057 0.152939
R20793 gnd.n5637 gnd.n5057 0.152939
R20794 gnd.n5638 gnd.n5637 0.152939
R20795 gnd.n5639 gnd.n5638 0.152939
R20796 gnd.n5640 gnd.n5639 0.152939
R20797 gnd.n5640 gnd.n5033 0.152939
R20798 gnd.n5667 gnd.n5033 0.152939
R20799 gnd.n5668 gnd.n5667 0.152939
R20800 gnd.n5669 gnd.n5668 0.152939
R20801 gnd.n5670 gnd.n5669 0.152939
R20802 gnd.n5670 gnd.n5002 0.152939
R20803 gnd.n5721 gnd.n5002 0.152939
R20804 gnd.n5722 gnd.n5721 0.152939
R20805 gnd.n5723 gnd.n5722 0.152939
R20806 gnd.n5723 gnd.n4981 0.152939
R20807 gnd.n5751 gnd.n4981 0.152939
R20808 gnd.n5752 gnd.n5751 0.152939
R20809 gnd.n5753 gnd.n5752 0.152939
R20810 gnd.n5754 gnd.n5753 0.152939
R20811 gnd.n5754 gnd.n4957 0.152939
R20812 gnd.n5797 gnd.n4957 0.152939
R20813 gnd.n5798 gnd.n5797 0.152939
R20814 gnd.n5799 gnd.n5798 0.152939
R20815 gnd.n5800 gnd.n5799 0.152939
R20816 gnd.n5800 gnd.n4927 0.152939
R20817 gnd.n6118 gnd.n4927 0.152939
R20818 gnd.n6119 gnd.n6118 0.152939
R20819 gnd.n6120 gnd.n6119 0.152939
R20820 gnd.n6121 gnd.n6120 0.152939
R20821 gnd.n6123 gnd.n6121 0.152939
R20822 gnd.n6123 gnd.n6122 0.152939
R20823 gnd.n6122 gnd.n914 0.152939
R20824 gnd.n915 gnd.n914 0.152939
R20825 gnd.n916 gnd.n915 0.152939
R20826 gnd.n4837 gnd.n916 0.152939
R20827 gnd.n4838 gnd.n4837 0.152939
R20828 gnd.n6233 gnd.n4838 0.152939
R20829 gnd.n5514 gnd.n5158 0.152939
R20830 gnd.n5179 gnd.n5158 0.152939
R20831 gnd.n5180 gnd.n5179 0.152939
R20832 gnd.n5186 gnd.n5180 0.152939
R20833 gnd.n5187 gnd.n5186 0.152939
R20834 gnd.n5188 gnd.n5187 0.152939
R20835 gnd.n5188 gnd.n5177 0.152939
R20836 gnd.n5196 gnd.n5177 0.152939
R20837 gnd.n5197 gnd.n5196 0.152939
R20838 gnd.n5198 gnd.n5197 0.152939
R20839 gnd.n5198 gnd.n5175 0.152939
R20840 gnd.n5206 gnd.n5175 0.152939
R20841 gnd.n5207 gnd.n5206 0.152939
R20842 gnd.n5208 gnd.n5207 0.152939
R20843 gnd.n5208 gnd.n5173 0.152939
R20844 gnd.n5216 gnd.n5173 0.152939
R20845 gnd.n6200 gnd.n4869 0.152939
R20846 gnd.n4871 gnd.n4869 0.152939
R20847 gnd.n4875 gnd.n4871 0.152939
R20848 gnd.n4876 gnd.n4875 0.152939
R20849 gnd.n4877 gnd.n4876 0.152939
R20850 gnd.n4878 gnd.n4877 0.152939
R20851 gnd.n4882 gnd.n4878 0.152939
R20852 gnd.n4883 gnd.n4882 0.152939
R20853 gnd.n4884 gnd.n4883 0.152939
R20854 gnd.n4885 gnd.n4884 0.152939
R20855 gnd.n4889 gnd.n4885 0.152939
R20856 gnd.n4890 gnd.n4889 0.152939
R20857 gnd.n4891 gnd.n4890 0.152939
R20858 gnd.n4892 gnd.n4891 0.152939
R20859 gnd.n4896 gnd.n4892 0.152939
R20860 gnd.n4897 gnd.n4896 0.152939
R20861 gnd.n4898 gnd.n4897 0.152939
R20862 gnd.n4899 gnd.n4898 0.152939
R20863 gnd.n4903 gnd.n4899 0.152939
R20864 gnd.n4904 gnd.n4903 0.152939
R20865 gnd.n4905 gnd.n4904 0.152939
R20866 gnd.n4906 gnd.n4905 0.152939
R20867 gnd.n4913 gnd.n4906 0.152939
R20868 gnd.n4914 gnd.n4913 0.152939
R20869 gnd.n4915 gnd.n4914 0.152939
R20870 gnd.n6152 gnd.n4915 0.152939
R20871 gnd.n5687 gnd.n5019 0.152939
R20872 gnd.n5688 gnd.n5687 0.152939
R20873 gnd.n5689 gnd.n5688 0.152939
R20874 gnd.n5690 gnd.n5689 0.152939
R20875 gnd.n5691 gnd.n5690 0.152939
R20876 gnd.n5692 gnd.n5691 0.152939
R20877 gnd.n5693 gnd.n5692 0.152939
R20878 gnd.n5694 gnd.n5693 0.152939
R20879 gnd.n5695 gnd.n5694 0.152939
R20880 gnd.n5695 gnd.n4963 0.152939
R20881 gnd.n5774 gnd.n4963 0.152939
R20882 gnd.n5775 gnd.n5774 0.152939
R20883 gnd.n5776 gnd.n5775 0.152939
R20884 gnd.n5777 gnd.n5776 0.152939
R20885 gnd.n5778 gnd.n5777 0.152939
R20886 gnd.n5779 gnd.n5778 0.152939
R20887 gnd.n5780 gnd.n5779 0.152939
R20888 gnd.n5781 gnd.n5780 0.152939
R20889 gnd.n5781 gnd.n4920 0.152939
R20890 gnd.n6133 gnd.n4920 0.152939
R20891 gnd.n6134 gnd.n6133 0.152939
R20892 gnd.n6135 gnd.n6134 0.152939
R20893 gnd.n6135 gnd.n4918 0.152939
R20894 gnd.n6143 gnd.n4918 0.152939
R20895 gnd.n6144 gnd.n6143 0.152939
R20896 gnd.n6145 gnd.n6144 0.152939
R20897 gnd.n6145 gnd.n4916 0.152939
R20898 gnd.n6151 gnd.n4916 0.152939
R20899 gnd.n5346 gnd.n5345 0.152939
R20900 gnd.n5346 gnd.n5236 0.152939
R20901 gnd.n5361 gnd.n5236 0.152939
R20902 gnd.n5362 gnd.n5361 0.152939
R20903 gnd.n5363 gnd.n5362 0.152939
R20904 gnd.n5363 gnd.n5224 0.152939
R20905 gnd.n5377 gnd.n5224 0.152939
R20906 gnd.n5378 gnd.n5377 0.152939
R20907 gnd.n5379 gnd.n5378 0.152939
R20908 gnd.n5380 gnd.n5379 0.152939
R20909 gnd.n5381 gnd.n5380 0.152939
R20910 gnd.n5382 gnd.n5381 0.152939
R20911 gnd.n5383 gnd.n5382 0.152939
R20912 gnd.n5384 gnd.n5383 0.152939
R20913 gnd.n5385 gnd.n5384 0.152939
R20914 gnd.n5386 gnd.n5385 0.152939
R20915 gnd.n5387 gnd.n5386 0.152939
R20916 gnd.n5388 gnd.n5387 0.152939
R20917 gnd.n5389 gnd.n5388 0.152939
R20918 gnd.n5390 gnd.n5389 0.152939
R20919 gnd.n5391 gnd.n5390 0.152939
R20920 gnd.n5392 gnd.n5391 0.152939
R20921 gnd.n5393 gnd.n5392 0.152939
R20922 gnd.n5394 gnd.n5393 0.152939
R20923 gnd.n5395 gnd.n5394 0.152939
R20924 gnd.n5396 gnd.n5395 0.152939
R20925 gnd.n5397 gnd.n5396 0.152939
R20926 gnd.n5398 gnd.n5397 0.152939
R20927 gnd.n5264 gnd.n5263 0.152939
R20928 gnd.n5265 gnd.n5264 0.152939
R20929 gnd.n5266 gnd.n5265 0.152939
R20930 gnd.n5267 gnd.n5266 0.152939
R20931 gnd.n5268 gnd.n5267 0.152939
R20932 gnd.n5269 gnd.n5268 0.152939
R20933 gnd.n5270 gnd.n5269 0.152939
R20934 gnd.n5271 gnd.n5270 0.152939
R20935 gnd.n5272 gnd.n5271 0.152939
R20936 gnd.n5273 gnd.n5272 0.152939
R20937 gnd.n5274 gnd.n5273 0.152939
R20938 gnd.n5275 gnd.n5274 0.152939
R20939 gnd.n5276 gnd.n5275 0.152939
R20940 gnd.n5277 gnd.n5276 0.152939
R20941 gnd.n5278 gnd.n5277 0.152939
R20942 gnd.n5279 gnd.n5278 0.152939
R20943 gnd.n5280 gnd.n5279 0.152939
R20944 gnd.n5281 gnd.n5280 0.152939
R20945 gnd.n5282 gnd.n5281 0.152939
R20946 gnd.n5283 gnd.n5282 0.152939
R20947 gnd.n5284 gnd.n5283 0.152939
R20948 gnd.n5285 gnd.n5284 0.152939
R20949 gnd.n5289 gnd.n5285 0.152939
R20950 gnd.n5290 gnd.n5289 0.152939
R20951 gnd.n5290 gnd.n5247 0.152939
R20952 gnd.n5344 gnd.n5247 0.152939
R20953 gnd.n6431 gnd.n6430 0.152939
R20954 gnd.n6432 gnd.n6431 0.152939
R20955 gnd.n6432 gnd.n720 0.152939
R20956 gnd.n6440 gnd.n720 0.152939
R20957 gnd.n6441 gnd.n6440 0.152939
R20958 gnd.n6442 gnd.n6441 0.152939
R20959 gnd.n6442 gnd.n714 0.152939
R20960 gnd.n6450 gnd.n714 0.152939
R20961 gnd.n6451 gnd.n6450 0.152939
R20962 gnd.n6452 gnd.n6451 0.152939
R20963 gnd.n6452 gnd.n708 0.152939
R20964 gnd.n6460 gnd.n708 0.152939
R20965 gnd.n6461 gnd.n6460 0.152939
R20966 gnd.n6462 gnd.n6461 0.152939
R20967 gnd.n6462 gnd.n702 0.152939
R20968 gnd.n6470 gnd.n702 0.152939
R20969 gnd.n6471 gnd.n6470 0.152939
R20970 gnd.n6472 gnd.n6471 0.152939
R20971 gnd.n6472 gnd.n696 0.152939
R20972 gnd.n6480 gnd.n696 0.152939
R20973 gnd.n6481 gnd.n6480 0.152939
R20974 gnd.n6482 gnd.n6481 0.152939
R20975 gnd.n6482 gnd.n690 0.152939
R20976 gnd.n6490 gnd.n690 0.152939
R20977 gnd.n6491 gnd.n6490 0.152939
R20978 gnd.n6492 gnd.n6491 0.152939
R20979 gnd.n6492 gnd.n684 0.152939
R20980 gnd.n6500 gnd.n684 0.152939
R20981 gnd.n6501 gnd.n6500 0.152939
R20982 gnd.n6502 gnd.n6501 0.152939
R20983 gnd.n6502 gnd.n678 0.152939
R20984 gnd.n6510 gnd.n678 0.152939
R20985 gnd.n6511 gnd.n6510 0.152939
R20986 gnd.n6512 gnd.n6511 0.152939
R20987 gnd.n6512 gnd.n672 0.152939
R20988 gnd.n6520 gnd.n672 0.152939
R20989 gnd.n6521 gnd.n6520 0.152939
R20990 gnd.n6522 gnd.n6521 0.152939
R20991 gnd.n6522 gnd.n666 0.152939
R20992 gnd.n6530 gnd.n666 0.152939
R20993 gnd.n6531 gnd.n6530 0.152939
R20994 gnd.n6532 gnd.n6531 0.152939
R20995 gnd.n6532 gnd.n660 0.152939
R20996 gnd.n6540 gnd.n660 0.152939
R20997 gnd.n6541 gnd.n6540 0.152939
R20998 gnd.n6542 gnd.n6541 0.152939
R20999 gnd.n6542 gnd.n654 0.152939
R21000 gnd.n6550 gnd.n654 0.152939
R21001 gnd.n6551 gnd.n6550 0.152939
R21002 gnd.n6552 gnd.n6551 0.152939
R21003 gnd.n6552 gnd.n648 0.152939
R21004 gnd.n6560 gnd.n648 0.152939
R21005 gnd.n6561 gnd.n6560 0.152939
R21006 gnd.n6562 gnd.n6561 0.152939
R21007 gnd.n6562 gnd.n642 0.152939
R21008 gnd.n6570 gnd.n642 0.152939
R21009 gnd.n6571 gnd.n6570 0.152939
R21010 gnd.n6572 gnd.n6571 0.152939
R21011 gnd.n6572 gnd.n636 0.152939
R21012 gnd.n6580 gnd.n636 0.152939
R21013 gnd.n6581 gnd.n6580 0.152939
R21014 gnd.n6582 gnd.n6581 0.152939
R21015 gnd.n6582 gnd.n630 0.152939
R21016 gnd.n6590 gnd.n630 0.152939
R21017 gnd.n6591 gnd.n6590 0.152939
R21018 gnd.n6592 gnd.n6591 0.152939
R21019 gnd.n6592 gnd.n624 0.152939
R21020 gnd.n6600 gnd.n624 0.152939
R21021 gnd.n6601 gnd.n6600 0.152939
R21022 gnd.n6602 gnd.n6601 0.152939
R21023 gnd.n6602 gnd.n618 0.152939
R21024 gnd.n6610 gnd.n618 0.152939
R21025 gnd.n6611 gnd.n6610 0.152939
R21026 gnd.n6612 gnd.n6611 0.152939
R21027 gnd.n6612 gnd.n612 0.152939
R21028 gnd.n6620 gnd.n612 0.152939
R21029 gnd.n6621 gnd.n6620 0.152939
R21030 gnd.n6622 gnd.n6621 0.152939
R21031 gnd.n6622 gnd.n606 0.152939
R21032 gnd.n6630 gnd.n606 0.152939
R21033 gnd.n6631 gnd.n6630 0.152939
R21034 gnd.n6632 gnd.n6631 0.152939
R21035 gnd.n6632 gnd.n600 0.152939
R21036 gnd.n6640 gnd.n600 0.152939
R21037 gnd.n6641 gnd.n6640 0.152939
R21038 gnd.n6642 gnd.n6641 0.152939
R21039 gnd.n6642 gnd.n594 0.152939
R21040 gnd.n6650 gnd.n594 0.152939
R21041 gnd.n6651 gnd.n6650 0.152939
R21042 gnd.n6652 gnd.n6651 0.152939
R21043 gnd.n6652 gnd.n588 0.152939
R21044 gnd.n6660 gnd.n588 0.152939
R21045 gnd.n6661 gnd.n6660 0.152939
R21046 gnd.n6662 gnd.n6661 0.152939
R21047 gnd.n6662 gnd.n582 0.152939
R21048 gnd.n6670 gnd.n582 0.152939
R21049 gnd.n6671 gnd.n6670 0.152939
R21050 gnd.n6672 gnd.n6671 0.152939
R21051 gnd.n6672 gnd.n576 0.152939
R21052 gnd.n6680 gnd.n576 0.152939
R21053 gnd.n6681 gnd.n6680 0.152939
R21054 gnd.n6682 gnd.n6681 0.152939
R21055 gnd.n6682 gnd.n570 0.152939
R21056 gnd.n6690 gnd.n570 0.152939
R21057 gnd.n6691 gnd.n6690 0.152939
R21058 gnd.n6692 gnd.n6691 0.152939
R21059 gnd.n6692 gnd.n564 0.152939
R21060 gnd.n6700 gnd.n564 0.152939
R21061 gnd.n6701 gnd.n6700 0.152939
R21062 gnd.n6702 gnd.n6701 0.152939
R21063 gnd.n6702 gnd.n558 0.152939
R21064 gnd.n6710 gnd.n558 0.152939
R21065 gnd.n6711 gnd.n6710 0.152939
R21066 gnd.n6712 gnd.n6711 0.152939
R21067 gnd.n6712 gnd.n552 0.152939
R21068 gnd.n6720 gnd.n552 0.152939
R21069 gnd.n6721 gnd.n6720 0.152939
R21070 gnd.n6722 gnd.n6721 0.152939
R21071 gnd.n6722 gnd.n546 0.152939
R21072 gnd.n6730 gnd.n546 0.152939
R21073 gnd.n6731 gnd.n6730 0.152939
R21074 gnd.n6732 gnd.n6731 0.152939
R21075 gnd.n6732 gnd.n540 0.152939
R21076 gnd.n6740 gnd.n540 0.152939
R21077 gnd.n6741 gnd.n6740 0.152939
R21078 gnd.n6742 gnd.n6741 0.152939
R21079 gnd.n6742 gnd.n534 0.152939
R21080 gnd.n6750 gnd.n534 0.152939
R21081 gnd.n6751 gnd.n6750 0.152939
R21082 gnd.n6752 gnd.n6751 0.152939
R21083 gnd.n6752 gnd.n528 0.152939
R21084 gnd.n6760 gnd.n528 0.152939
R21085 gnd.n6761 gnd.n6760 0.152939
R21086 gnd.n6762 gnd.n6761 0.152939
R21087 gnd.n6762 gnd.n522 0.152939
R21088 gnd.n6770 gnd.n522 0.152939
R21089 gnd.n6771 gnd.n6770 0.152939
R21090 gnd.n6772 gnd.n6771 0.152939
R21091 gnd.n6772 gnd.n516 0.152939
R21092 gnd.n6780 gnd.n516 0.152939
R21093 gnd.n6781 gnd.n6780 0.152939
R21094 gnd.n6782 gnd.n6781 0.152939
R21095 gnd.n6782 gnd.n510 0.152939
R21096 gnd.n6790 gnd.n510 0.152939
R21097 gnd.n6791 gnd.n6790 0.152939
R21098 gnd.n6792 gnd.n6791 0.152939
R21099 gnd.n6792 gnd.n504 0.152939
R21100 gnd.n6800 gnd.n504 0.152939
R21101 gnd.n6801 gnd.n6800 0.152939
R21102 gnd.n6802 gnd.n6801 0.152939
R21103 gnd.n6802 gnd.n498 0.152939
R21104 gnd.n6810 gnd.n498 0.152939
R21105 gnd.n6811 gnd.n6810 0.152939
R21106 gnd.n6812 gnd.n6811 0.152939
R21107 gnd.n6812 gnd.n492 0.152939
R21108 gnd.n6820 gnd.n492 0.152939
R21109 gnd.n6821 gnd.n6820 0.152939
R21110 gnd.n6822 gnd.n6821 0.152939
R21111 gnd.n6822 gnd.n486 0.152939
R21112 gnd.n6830 gnd.n486 0.152939
R21113 gnd.n6831 gnd.n6830 0.152939
R21114 gnd.n6832 gnd.n6831 0.152939
R21115 gnd.n6832 gnd.n480 0.152939
R21116 gnd.n6840 gnd.n480 0.152939
R21117 gnd.n6841 gnd.n6840 0.152939
R21118 gnd.n6842 gnd.n6841 0.152939
R21119 gnd.n6842 gnd.n474 0.152939
R21120 gnd.n6850 gnd.n474 0.152939
R21121 gnd.n6851 gnd.n6850 0.152939
R21122 gnd.n6852 gnd.n6851 0.152939
R21123 gnd.n6852 gnd.n468 0.152939
R21124 gnd.n6860 gnd.n468 0.152939
R21125 gnd.n6861 gnd.n6860 0.152939
R21126 gnd.n6862 gnd.n6861 0.152939
R21127 gnd.n6862 gnd.n462 0.152939
R21128 gnd.n6870 gnd.n462 0.152939
R21129 gnd.n6871 gnd.n6870 0.152939
R21130 gnd.n6873 gnd.n6871 0.152939
R21131 gnd.n6873 gnd.n6872 0.152939
R21132 gnd.n6872 gnd.n456 0.152939
R21133 gnd.n6882 gnd.n456 0.152939
R21134 gnd.n6883 gnd.n451 0.152939
R21135 gnd.n6891 gnd.n451 0.152939
R21136 gnd.n6892 gnd.n6891 0.152939
R21137 gnd.n6893 gnd.n6892 0.152939
R21138 gnd.n6893 gnd.n445 0.152939
R21139 gnd.n6901 gnd.n445 0.152939
R21140 gnd.n6902 gnd.n6901 0.152939
R21141 gnd.n6903 gnd.n6902 0.152939
R21142 gnd.n6903 gnd.n439 0.152939
R21143 gnd.n6911 gnd.n439 0.152939
R21144 gnd.n6912 gnd.n6911 0.152939
R21145 gnd.n6913 gnd.n6912 0.152939
R21146 gnd.n6913 gnd.n433 0.152939
R21147 gnd.n6921 gnd.n433 0.152939
R21148 gnd.n6922 gnd.n6921 0.152939
R21149 gnd.n6923 gnd.n6922 0.152939
R21150 gnd.n6923 gnd.n427 0.152939
R21151 gnd.n6931 gnd.n427 0.152939
R21152 gnd.n6932 gnd.n6931 0.152939
R21153 gnd.n6933 gnd.n6932 0.152939
R21154 gnd.n6933 gnd.n421 0.152939
R21155 gnd.n6941 gnd.n421 0.152939
R21156 gnd.n6942 gnd.n6941 0.152939
R21157 gnd.n6943 gnd.n6942 0.152939
R21158 gnd.n6943 gnd.n415 0.152939
R21159 gnd.n6951 gnd.n415 0.152939
R21160 gnd.n6952 gnd.n6951 0.152939
R21161 gnd.n6953 gnd.n6952 0.152939
R21162 gnd.n6953 gnd.n409 0.152939
R21163 gnd.n6961 gnd.n409 0.152939
R21164 gnd.n6962 gnd.n6961 0.152939
R21165 gnd.n6963 gnd.n6962 0.152939
R21166 gnd.n6963 gnd.n403 0.152939
R21167 gnd.n6971 gnd.n403 0.152939
R21168 gnd.n6972 gnd.n6971 0.152939
R21169 gnd.n6973 gnd.n6972 0.152939
R21170 gnd.n6973 gnd.n397 0.152939
R21171 gnd.n6981 gnd.n397 0.152939
R21172 gnd.n6982 gnd.n6981 0.152939
R21173 gnd.n6983 gnd.n6982 0.152939
R21174 gnd.n6983 gnd.n391 0.152939
R21175 gnd.n6991 gnd.n391 0.152939
R21176 gnd.n6992 gnd.n6991 0.152939
R21177 gnd.n6993 gnd.n6992 0.152939
R21178 gnd.n6993 gnd.n385 0.152939
R21179 gnd.n7001 gnd.n385 0.152939
R21180 gnd.n7002 gnd.n7001 0.152939
R21181 gnd.n7003 gnd.n7002 0.152939
R21182 gnd.n7003 gnd.n379 0.152939
R21183 gnd.n7011 gnd.n379 0.152939
R21184 gnd.n7012 gnd.n7011 0.152939
R21185 gnd.n7013 gnd.n7012 0.152939
R21186 gnd.n7013 gnd.n373 0.152939
R21187 gnd.n7021 gnd.n373 0.152939
R21188 gnd.n7022 gnd.n7021 0.152939
R21189 gnd.n7023 gnd.n7022 0.152939
R21190 gnd.n7023 gnd.n367 0.152939
R21191 gnd.n7031 gnd.n367 0.152939
R21192 gnd.n7032 gnd.n7031 0.152939
R21193 gnd.n7033 gnd.n7032 0.152939
R21194 gnd.n7033 gnd.n361 0.152939
R21195 gnd.n7041 gnd.n361 0.152939
R21196 gnd.n7042 gnd.n7041 0.152939
R21197 gnd.n7043 gnd.n7042 0.152939
R21198 gnd.n7043 gnd.n355 0.152939
R21199 gnd.n7051 gnd.n355 0.152939
R21200 gnd.n7052 gnd.n7051 0.152939
R21201 gnd.n7053 gnd.n7052 0.152939
R21202 gnd.n7053 gnd.n349 0.152939
R21203 gnd.n7061 gnd.n349 0.152939
R21204 gnd.n7062 gnd.n7061 0.152939
R21205 gnd.n7063 gnd.n7062 0.152939
R21206 gnd.n7063 gnd.n343 0.152939
R21207 gnd.n7071 gnd.n343 0.152939
R21208 gnd.n7072 gnd.n7071 0.152939
R21209 gnd.n7073 gnd.n7072 0.152939
R21210 gnd.n7073 gnd.n337 0.152939
R21211 gnd.n7081 gnd.n337 0.152939
R21212 gnd.n7082 gnd.n7081 0.152939
R21213 gnd.n7083 gnd.n7082 0.152939
R21214 gnd.n7083 gnd.n331 0.152939
R21215 gnd.n7092 gnd.n331 0.152939
R21216 gnd.n7093 gnd.n7092 0.152939
R21217 gnd.n7095 gnd.n7093 0.152939
R21218 gnd.n327 gnd.n326 0.152939
R21219 gnd.n7094 gnd.n327 0.152939
R21220 gnd.n7237 gnd.n253 0.152939
R21221 gnd.n7238 gnd.n7237 0.152939
R21222 gnd.n7239 gnd.n7238 0.152939
R21223 gnd.n7239 gnd.n235 0.152939
R21224 gnd.n7253 gnd.n235 0.152939
R21225 gnd.n7254 gnd.n7253 0.152939
R21226 gnd.n7255 gnd.n7254 0.152939
R21227 gnd.n7255 gnd.n222 0.152939
R21228 gnd.n7269 gnd.n222 0.152939
R21229 gnd.n7270 gnd.n7269 0.152939
R21230 gnd.n7271 gnd.n7270 0.152939
R21231 gnd.n7271 gnd.n205 0.152939
R21232 gnd.n7285 gnd.n205 0.152939
R21233 gnd.n7286 gnd.n7285 0.152939
R21234 gnd.n7287 gnd.n7286 0.152939
R21235 gnd.n7287 gnd.n190 0.152939
R21236 gnd.n7376 gnd.n190 0.152939
R21237 gnd.n7377 gnd.n7376 0.152939
R21238 gnd.n7378 gnd.n7377 0.152939
R21239 gnd.n7378 gnd.n111 0.152939
R21240 gnd.n7458 gnd.n111 0.152939
R21241 gnd.n7457 gnd.n112 0.152939
R21242 gnd.n114 gnd.n112 0.152939
R21243 gnd.n118 gnd.n114 0.152939
R21244 gnd.n119 gnd.n118 0.152939
R21245 gnd.n120 gnd.n119 0.152939
R21246 gnd.n121 gnd.n120 0.152939
R21247 gnd.n125 gnd.n121 0.152939
R21248 gnd.n126 gnd.n125 0.152939
R21249 gnd.n127 gnd.n126 0.152939
R21250 gnd.n128 gnd.n127 0.152939
R21251 gnd.n132 gnd.n128 0.152939
R21252 gnd.n133 gnd.n132 0.152939
R21253 gnd.n134 gnd.n133 0.152939
R21254 gnd.n135 gnd.n134 0.152939
R21255 gnd.n139 gnd.n135 0.152939
R21256 gnd.n140 gnd.n139 0.152939
R21257 gnd.n141 gnd.n140 0.152939
R21258 gnd.n142 gnd.n141 0.152939
R21259 gnd.n146 gnd.n142 0.152939
R21260 gnd.n147 gnd.n146 0.152939
R21261 gnd.n148 gnd.n147 0.152939
R21262 gnd.n149 gnd.n148 0.152939
R21263 gnd.n153 gnd.n149 0.152939
R21264 gnd.n154 gnd.n153 0.152939
R21265 gnd.n155 gnd.n154 0.152939
R21266 gnd.n156 gnd.n155 0.152939
R21267 gnd.n160 gnd.n156 0.152939
R21268 gnd.n161 gnd.n160 0.152939
R21269 gnd.n162 gnd.n161 0.152939
R21270 gnd.n163 gnd.n162 0.152939
R21271 gnd.n167 gnd.n163 0.152939
R21272 gnd.n168 gnd.n167 0.152939
R21273 gnd.n169 gnd.n168 0.152939
R21274 gnd.n170 gnd.n169 0.152939
R21275 gnd.n174 gnd.n170 0.152939
R21276 gnd.n175 gnd.n174 0.152939
R21277 gnd.n7388 gnd.n175 0.152939
R21278 gnd.n7388 gnd.n7387 0.152939
R21279 gnd.n1649 gnd.n1494 0.152939
R21280 gnd.n1650 gnd.n1649 0.152939
R21281 gnd.n1651 gnd.n1650 0.152939
R21282 gnd.n1652 gnd.n1651 0.152939
R21283 gnd.n1653 gnd.n1652 0.152939
R21284 gnd.n1654 gnd.n1653 0.152939
R21285 gnd.n1655 gnd.n1654 0.152939
R21286 gnd.n1656 gnd.n1655 0.152939
R21287 gnd.n1657 gnd.n1656 0.152939
R21288 gnd.n1658 gnd.n1657 0.152939
R21289 gnd.n1659 gnd.n1658 0.152939
R21290 gnd.n1660 gnd.n1659 0.152939
R21291 gnd.n1661 gnd.n1660 0.152939
R21292 gnd.n1661 gnd.n1557 0.152939
R21293 gnd.n4256 gnd.n1557 0.152939
R21294 gnd.n4257 gnd.n4256 0.152939
R21295 gnd.n4258 gnd.n4257 0.152939
R21296 gnd.n4258 gnd.n1555 0.152939
R21297 gnd.n4263 gnd.n1555 0.152939
R21298 gnd.n4264 gnd.n4263 0.152939
R21299 gnd.n4265 gnd.n4264 0.152939
R21300 gnd.n4266 gnd.n4265 0.152939
R21301 gnd.n4267 gnd.n4266 0.152939
R21302 gnd.n4269 gnd.n4267 0.152939
R21303 gnd.n4269 gnd.n4268 0.152939
R21304 gnd.n4268 gnd.n300 0.152939
R21305 gnd.n7137 gnd.n7136 0.152939
R21306 gnd.n7138 gnd.n7137 0.152939
R21307 gnd.n7139 gnd.n7138 0.152939
R21308 gnd.n7140 gnd.n7139 0.152939
R21309 gnd.n7141 gnd.n7140 0.152939
R21310 gnd.n7142 gnd.n7141 0.152939
R21311 gnd.n7143 gnd.n7142 0.152939
R21312 gnd.n7144 gnd.n7143 0.152939
R21313 gnd.n7145 gnd.n7144 0.152939
R21314 gnd.n7146 gnd.n7145 0.152939
R21315 gnd.n7147 gnd.n7146 0.152939
R21316 gnd.n7148 gnd.n7147 0.152939
R21317 gnd.n7149 gnd.n7148 0.152939
R21318 gnd.n7150 gnd.n7149 0.152939
R21319 gnd.n7151 gnd.n7150 0.152939
R21320 gnd.n7152 gnd.n7151 0.152939
R21321 gnd.n7153 gnd.n7152 0.152939
R21322 gnd.n7154 gnd.n7153 0.152939
R21323 gnd.n7155 gnd.n7154 0.152939
R21324 gnd.n7156 gnd.n7155 0.152939
R21325 gnd.n7157 gnd.n7156 0.152939
R21326 gnd.n7158 gnd.n7157 0.152939
R21327 gnd.n7160 gnd.n7158 0.152939
R21328 gnd.n7160 gnd.n7159 0.152939
R21329 gnd.n7159 gnd.n181 0.152939
R21330 gnd.n7386 gnd.n181 0.152939
R21331 gnd.n1451 gnd.n1450 0.152939
R21332 gnd.n1452 gnd.n1451 0.152939
R21333 gnd.n1453 gnd.n1452 0.152939
R21334 gnd.n1454 gnd.n1453 0.152939
R21335 gnd.n1455 gnd.n1454 0.152939
R21336 gnd.n1456 gnd.n1455 0.152939
R21337 gnd.n1457 gnd.n1456 0.152939
R21338 gnd.n1458 gnd.n1457 0.152939
R21339 gnd.n1459 gnd.n1458 0.152939
R21340 gnd.n1460 gnd.n1459 0.152939
R21341 gnd.n1461 gnd.n1460 0.152939
R21342 gnd.n1462 gnd.n1461 0.152939
R21343 gnd.n1463 gnd.n1462 0.152939
R21344 gnd.n1464 gnd.n1463 0.152939
R21345 gnd.n1465 gnd.n1464 0.152939
R21346 gnd.n1472 gnd.n1471 0.152939
R21347 gnd.n1473 gnd.n1472 0.152939
R21348 gnd.n1474 gnd.n1473 0.152939
R21349 gnd.n1475 gnd.n1474 0.152939
R21350 gnd.n1476 gnd.n1475 0.152939
R21351 gnd.n1477 gnd.n1476 0.152939
R21352 gnd.n1478 gnd.n1477 0.152939
R21353 gnd.n1479 gnd.n1478 0.152939
R21354 gnd.n1480 gnd.n1479 0.152939
R21355 gnd.n1481 gnd.n1480 0.152939
R21356 gnd.n1482 gnd.n1481 0.152939
R21357 gnd.n1483 gnd.n1482 0.152939
R21358 gnd.n1484 gnd.n1483 0.152939
R21359 gnd.n1485 gnd.n1484 0.152939
R21360 gnd.n1486 gnd.n1485 0.152939
R21361 gnd.n1487 gnd.n1486 0.152939
R21362 gnd.n1488 gnd.n1487 0.152939
R21363 gnd.n4355 gnd.n1488 0.152939
R21364 gnd.n4355 gnd.n4354 0.152939
R21365 gnd.n4354 gnd.n4353 0.152939
R21366 gnd.n1644 gnd.n1643 0.152939
R21367 gnd.n1644 gnd.n1622 0.152939
R21368 gnd.n4178 gnd.n1622 0.152939
R21369 gnd.n4179 gnd.n4178 0.152939
R21370 gnd.n4180 gnd.n4179 0.152939
R21371 gnd.n4181 gnd.n4180 0.152939
R21372 gnd.n4181 gnd.n1594 0.152939
R21373 gnd.n4209 gnd.n1594 0.152939
R21374 gnd.n4210 gnd.n4209 0.152939
R21375 gnd.n4211 gnd.n4210 0.152939
R21376 gnd.n4212 gnd.n4211 0.152939
R21377 gnd.n4212 gnd.n1567 0.152939
R21378 gnd.n4246 gnd.n1567 0.152939
R21379 gnd.n4247 gnd.n4246 0.152939
R21380 gnd.n4248 gnd.n4247 0.152939
R21381 gnd.n4249 gnd.n4248 0.152939
R21382 gnd.n4249 gnd.n1532 0.152939
R21383 gnd.n4309 gnd.n1532 0.152939
R21384 gnd.n4310 gnd.n4309 0.152939
R21385 gnd.n4311 gnd.n4310 0.152939
R21386 gnd.n4311 gnd.n268 0.152939
R21387 gnd.n2385 gnd.n2368 0.152939
R21388 gnd.n2371 gnd.n2368 0.152939
R21389 gnd.n2372 gnd.n2371 0.152939
R21390 gnd.n2373 gnd.n2372 0.152939
R21391 gnd.n2375 gnd.n2373 0.152939
R21392 gnd.n2375 gnd.n2374 0.152939
R21393 gnd.n2374 gnd.n2335 0.152939
R21394 gnd.n2714 gnd.n2335 0.152939
R21395 gnd.n2715 gnd.n2714 0.152939
R21396 gnd.n2716 gnd.n2715 0.152939
R21397 gnd.n2716 gnd.n2331 0.152939
R21398 gnd.n2722 gnd.n2331 0.152939
R21399 gnd.n2723 gnd.n2722 0.152939
R21400 gnd.n2724 gnd.n2723 0.152939
R21401 gnd.n2725 gnd.n2724 0.152939
R21402 gnd.n2726 gnd.n2725 0.152939
R21403 gnd.n2729 gnd.n2726 0.152939
R21404 gnd.n2730 gnd.n2729 0.152939
R21405 gnd.n2731 gnd.n2730 0.152939
R21406 gnd.n2732 gnd.n2731 0.152939
R21407 gnd.n2735 gnd.n2732 0.152939
R21408 gnd.n2736 gnd.n2735 0.152939
R21409 gnd.n2737 gnd.n2736 0.152939
R21410 gnd.n2738 gnd.n2737 0.152939
R21411 gnd.n2740 gnd.n2738 0.152939
R21412 gnd.n2741 gnd.n2740 0.152939
R21413 gnd.n2741 gnd.n2156 0.152939
R21414 gnd.n3732 gnd.n2156 0.152939
R21415 gnd.n3733 gnd.n3732 0.152939
R21416 gnd.n3734 gnd.n3733 0.152939
R21417 gnd.n3734 gnd.n2142 0.152939
R21418 gnd.n3748 gnd.n2142 0.152939
R21419 gnd.n3749 gnd.n3748 0.152939
R21420 gnd.n3750 gnd.n3749 0.152939
R21421 gnd.n3750 gnd.n2130 0.152939
R21422 gnd.n3764 gnd.n2130 0.152939
R21423 gnd.n3765 gnd.n3764 0.152939
R21424 gnd.n3766 gnd.n3765 0.152939
R21425 gnd.n3766 gnd.n2117 0.152939
R21426 gnd.n3780 gnd.n2117 0.152939
R21427 gnd.n3781 gnd.n3780 0.152939
R21428 gnd.n3782 gnd.n3781 0.152939
R21429 gnd.n3782 gnd.n2104 0.152939
R21430 gnd.n3796 gnd.n2104 0.152939
R21431 gnd.n3797 gnd.n3796 0.152939
R21432 gnd.n3798 gnd.n3797 0.152939
R21433 gnd.n3798 gnd.n2090 0.152939
R21434 gnd.n3812 gnd.n2090 0.152939
R21435 gnd.n3813 gnd.n3812 0.152939
R21436 gnd.n3814 gnd.n3813 0.152939
R21437 gnd.n3814 gnd.n2078 0.152939
R21438 gnd.n3828 gnd.n2078 0.152939
R21439 gnd.n3829 gnd.n3828 0.152939
R21440 gnd.n3830 gnd.n3829 0.152939
R21441 gnd.n3830 gnd.n2063 0.152939
R21442 gnd.n3844 gnd.n2063 0.152939
R21443 gnd.n3845 gnd.n3844 0.152939
R21444 gnd.n3846 gnd.n3845 0.152939
R21445 gnd.n3846 gnd.n2048 0.152939
R21446 gnd.n3860 gnd.n2048 0.152939
R21447 gnd.n3861 gnd.n3860 0.152939
R21448 gnd.n3862 gnd.n3861 0.152939
R21449 gnd.n3862 gnd.n2035 0.152939
R21450 gnd.n3876 gnd.n2035 0.152939
R21451 gnd.n3877 gnd.n3876 0.152939
R21452 gnd.n3878 gnd.n3877 0.152939
R21453 gnd.n3878 gnd.n2020 0.152939
R21454 gnd.n3892 gnd.n2020 0.152939
R21455 gnd.n3893 gnd.n3892 0.152939
R21456 gnd.n3894 gnd.n3893 0.152939
R21457 gnd.n3894 gnd.n2005 0.152939
R21458 gnd.n3908 gnd.n2005 0.152939
R21459 gnd.n3909 gnd.n3908 0.152939
R21460 gnd.n3910 gnd.n3909 0.152939
R21461 gnd.n3910 gnd.n1992 0.152939
R21462 gnd.n3924 gnd.n1992 0.152939
R21463 gnd.n3925 gnd.n3924 0.152939
R21464 gnd.n3926 gnd.n3925 0.152939
R21465 gnd.n3926 gnd.n1978 0.152939
R21466 gnd.n3940 gnd.n1978 0.152939
R21467 gnd.n3941 gnd.n3940 0.152939
R21468 gnd.n3942 gnd.n3941 0.152939
R21469 gnd.n3942 gnd.n1963 0.152939
R21470 gnd.n3956 gnd.n1963 0.152939
R21471 gnd.n3957 gnd.n3956 0.152939
R21472 gnd.n3958 gnd.n3957 0.152939
R21473 gnd.n3958 gnd.n1950 0.152939
R21474 gnd.n3972 gnd.n1950 0.152939
R21475 gnd.n3973 gnd.n3972 0.152939
R21476 gnd.n3974 gnd.n3973 0.152939
R21477 gnd.n3974 gnd.n1935 0.152939
R21478 gnd.n3988 gnd.n1935 0.152939
R21479 gnd.n3989 gnd.n3988 0.152939
R21480 gnd.n3990 gnd.n3989 0.152939
R21481 gnd.n3990 gnd.n1922 0.152939
R21482 gnd.n4004 gnd.n1922 0.152939
R21483 gnd.n4005 gnd.n4004 0.152939
R21484 gnd.n4006 gnd.n4005 0.152939
R21485 gnd.n4006 gnd.n1908 0.152939
R21486 gnd.n4020 gnd.n1908 0.152939
R21487 gnd.n4021 gnd.n4020 0.152939
R21488 gnd.n4022 gnd.n4021 0.152939
R21489 gnd.n4022 gnd.n1893 0.152939
R21490 gnd.n4036 gnd.n1893 0.152939
R21491 gnd.n4037 gnd.n4036 0.152939
R21492 gnd.n4038 gnd.n4037 0.152939
R21493 gnd.n4038 gnd.n1881 0.152939
R21494 gnd.n4052 gnd.n1881 0.152939
R21495 gnd.n4053 gnd.n4052 0.152939
R21496 gnd.n4054 gnd.n4053 0.152939
R21497 gnd.n4054 gnd.n1868 0.152939
R21498 gnd.n4068 gnd.n1868 0.152939
R21499 gnd.n4069 gnd.n4068 0.152939
R21500 gnd.n4070 gnd.n4069 0.152939
R21501 gnd.n4070 gnd.n1855 0.152939
R21502 gnd.n4084 gnd.n1855 0.152939
R21503 gnd.n4085 gnd.n4084 0.152939
R21504 gnd.n4086 gnd.n4085 0.152939
R21505 gnd.n4086 gnd.n1841 0.152939
R21506 gnd.n4100 gnd.n1841 0.152939
R21507 gnd.n4101 gnd.n4100 0.152939
R21508 gnd.n4102 gnd.n4101 0.152939
R21509 gnd.n4102 gnd.n1828 0.152939
R21510 gnd.n4118 gnd.n1828 0.152939
R21511 gnd.n4119 gnd.n4118 0.152939
R21512 gnd.n4120 gnd.n4119 0.152939
R21513 gnd.n4122 gnd.n4120 0.152939
R21514 gnd.n4122 gnd.n4121 0.152939
R21515 gnd.n4121 gnd.n1412 0.152939
R21516 gnd.n1413 gnd.n1412 0.152939
R21517 gnd.n1414 gnd.n1413 0.152939
R21518 gnd.n1636 gnd.n1414 0.152939
R21519 gnd.n1637 gnd.n1636 0.152939
R21520 gnd.n1638 gnd.n1637 0.152939
R21521 gnd.n1638 gnd.n1632 0.152939
R21522 gnd.n4167 gnd.n1632 0.152939
R21523 gnd.n4168 gnd.n4167 0.152939
R21524 gnd.n4169 gnd.n4168 0.152939
R21525 gnd.n4170 gnd.n4169 0.152939
R21526 gnd.n4170 gnd.n1605 0.152939
R21527 gnd.n4198 gnd.n1605 0.152939
R21528 gnd.n4199 gnd.n4198 0.152939
R21529 gnd.n4200 gnd.n4199 0.152939
R21530 gnd.n4201 gnd.n4200 0.152939
R21531 gnd.n4201 gnd.n1577 0.152939
R21532 gnd.n4234 gnd.n1577 0.152939
R21533 gnd.n4235 gnd.n4234 0.152939
R21534 gnd.n4236 gnd.n4235 0.152939
R21535 gnd.n4237 gnd.n4236 0.152939
R21536 gnd.n4237 gnd.n1543 0.152939
R21537 gnd.n4292 gnd.n1543 0.152939
R21538 gnd.n4293 gnd.n4292 0.152939
R21539 gnd.n4294 gnd.n4293 0.152939
R21540 gnd.n4295 gnd.n4294 0.152939
R21541 gnd.n4296 gnd.n4295 0.152939
R21542 gnd.n1163 gnd.n1162 0.152939
R21543 gnd.n1181 gnd.n1163 0.152939
R21544 gnd.n1182 gnd.n1181 0.152939
R21545 gnd.n1183 gnd.n1182 0.152939
R21546 gnd.n1184 gnd.n1183 0.152939
R21547 gnd.n1202 gnd.n1184 0.152939
R21548 gnd.n1203 gnd.n1202 0.152939
R21549 gnd.n1204 gnd.n1203 0.152939
R21550 gnd.n1205 gnd.n1204 0.152939
R21551 gnd.n1223 gnd.n1205 0.152939
R21552 gnd.n1224 gnd.n1223 0.152939
R21553 gnd.n1225 gnd.n1224 0.152939
R21554 gnd.n1226 gnd.n1225 0.152939
R21555 gnd.n1244 gnd.n1226 0.152939
R21556 gnd.n1245 gnd.n1244 0.152939
R21557 gnd.n1246 gnd.n1245 0.152939
R21558 gnd.n1247 gnd.n1246 0.152939
R21559 gnd.n1265 gnd.n1247 0.152939
R21560 gnd.n1266 gnd.n1265 0.152939
R21561 gnd.n1267 gnd.n1266 0.152939
R21562 gnd.n1268 gnd.n1267 0.152939
R21563 gnd.n2274 gnd.n2273 0.152939
R21564 gnd.n2275 gnd.n2274 0.152939
R21565 gnd.n2276 gnd.n2275 0.152939
R21566 gnd.n2277 gnd.n2276 0.152939
R21567 gnd.n2278 gnd.n2277 0.152939
R21568 gnd.n2279 gnd.n2278 0.152939
R21569 gnd.n2280 gnd.n2279 0.152939
R21570 gnd.n2281 gnd.n2280 0.152939
R21571 gnd.n2282 gnd.n2281 0.152939
R21572 gnd.n2283 gnd.n2282 0.152939
R21573 gnd.n2284 gnd.n2283 0.152939
R21574 gnd.n2285 gnd.n2284 0.152939
R21575 gnd.n2286 gnd.n2285 0.152939
R21576 gnd.n2287 gnd.n2286 0.152939
R21577 gnd.n2288 gnd.n2287 0.152939
R21578 gnd.n2868 gnd.n2867 0.152939
R21579 gnd.n2867 gnd.n2293 0.152939
R21580 gnd.n2294 gnd.n2293 0.152939
R21581 gnd.n2295 gnd.n2294 0.152939
R21582 gnd.n2296 gnd.n2295 0.152939
R21583 gnd.n2297 gnd.n2296 0.152939
R21584 gnd.n2298 gnd.n2297 0.152939
R21585 gnd.n2299 gnd.n2298 0.152939
R21586 gnd.n2300 gnd.n2299 0.152939
R21587 gnd.n2301 gnd.n2300 0.152939
R21588 gnd.n2302 gnd.n2301 0.152939
R21589 gnd.n2303 gnd.n2302 0.152939
R21590 gnd.n2304 gnd.n2303 0.152939
R21591 gnd.n2305 gnd.n2304 0.152939
R21592 gnd.n2306 gnd.n2305 0.152939
R21593 gnd.n2307 gnd.n2306 0.152939
R21594 gnd.n2308 gnd.n2307 0.152939
R21595 gnd.n2309 gnd.n2308 0.152939
R21596 gnd.n2827 gnd.n2309 0.152939
R21597 gnd.n2827 gnd.n2826 0.152939
R21598 gnd.n2481 gnd.n2454 0.152939
R21599 gnd.n2539 gnd.n2454 0.152939
R21600 gnd.n2540 gnd.n2539 0.152939
R21601 gnd.n2541 gnd.n2540 0.152939
R21602 gnd.n2541 gnd.n2452 0.152939
R21603 gnd.n2547 gnd.n2452 0.152939
R21604 gnd.n2548 gnd.n2547 0.152939
R21605 gnd.n2549 gnd.n2548 0.152939
R21606 gnd.n2549 gnd.n2450 0.152939
R21607 gnd.n2555 gnd.n2450 0.152939
R21608 gnd.n2556 gnd.n2555 0.152939
R21609 gnd.n2557 gnd.n2556 0.152939
R21610 gnd.n2557 gnd.n2448 0.152939
R21611 gnd.n2563 gnd.n2448 0.152939
R21612 gnd.n2564 gnd.n2563 0.152939
R21613 gnd.n2565 gnd.n2564 0.152939
R21614 gnd.n2565 gnd.n2446 0.152939
R21615 gnd.n2571 gnd.n2446 0.152939
R21616 gnd.n2572 gnd.n2571 0.152939
R21617 gnd.n2574 gnd.n2572 0.152939
R21618 gnd.n2574 gnd.n2573 0.152939
R21619 gnd.n2573 gnd.n2401 0.152939
R21620 gnd.n2402 gnd.n2401 0.152939
R21621 gnd.n2403 gnd.n2402 0.152939
R21622 gnd.n2600 gnd.n2403 0.152939
R21623 gnd.n2601 gnd.n2600 0.152939
R21624 gnd.n2520 gnd.n2461 0.152939
R21625 gnd.n2462 gnd.n2461 0.152939
R21626 gnd.n2463 gnd.n2462 0.152939
R21627 gnd.n2464 gnd.n2463 0.152939
R21628 gnd.n2465 gnd.n2464 0.152939
R21629 gnd.n2466 gnd.n2465 0.152939
R21630 gnd.n2467 gnd.n2466 0.152939
R21631 gnd.n2468 gnd.n2467 0.152939
R21632 gnd.n2469 gnd.n2468 0.152939
R21633 gnd.n2470 gnd.n2469 0.152939
R21634 gnd.n2471 gnd.n2470 0.152939
R21635 gnd.n2472 gnd.n2471 0.152939
R21636 gnd.n2473 gnd.n2472 0.152939
R21637 gnd.n2474 gnd.n2473 0.152939
R21638 gnd.n2475 gnd.n2474 0.152939
R21639 gnd.n2485 gnd.n2475 0.152939
R21640 gnd.n2485 gnd.n2484 0.152939
R21641 gnd.n2484 gnd.n2483 0.152939
R21642 gnd.n2526 gnd.n2521 0.152939
R21643 gnd.n2526 gnd.n2525 0.152939
R21644 gnd.n2525 gnd.n2524 0.152939
R21645 gnd.n2524 gnd.n2522 0.152939
R21646 gnd.n2522 gnd.n1033 0.152939
R21647 gnd.n1034 gnd.n1033 0.152939
R21648 gnd.n1035 gnd.n1034 0.152939
R21649 gnd.n1051 gnd.n1035 0.152939
R21650 gnd.n1052 gnd.n1051 0.152939
R21651 gnd.n1053 gnd.n1052 0.152939
R21652 gnd.n1054 gnd.n1053 0.152939
R21653 gnd.n1072 gnd.n1054 0.152939
R21654 gnd.n1073 gnd.n1072 0.152939
R21655 gnd.n1074 gnd.n1073 0.152939
R21656 gnd.n1075 gnd.n1074 0.152939
R21657 gnd.n1091 gnd.n1075 0.152939
R21658 gnd.n1092 gnd.n1091 0.152939
R21659 gnd.n1093 gnd.n1092 0.152939
R21660 gnd.n1094 gnd.n1093 0.152939
R21661 gnd.n1114 gnd.n1094 0.152939
R21662 gnd.n1115 gnd.n1114 0.152939
R21663 gnd.n1116 gnd.n1115 0.152939
R21664 gnd.n1117 gnd.n1116 0.152939
R21665 gnd.n1132 gnd.n1117 0.152939
R21666 gnd.n1133 gnd.n1132 0.152939
R21667 gnd.n1134 gnd.n1133 0.152939
R21668 gnd.n1151 gnd.n1135 0.152939
R21669 gnd.n1152 gnd.n1151 0.152939
R21670 gnd.n1153 gnd.n1152 0.152939
R21671 gnd.n1154 gnd.n1153 0.152939
R21672 gnd.n1170 gnd.n1154 0.152939
R21673 gnd.n1171 gnd.n1170 0.152939
R21674 gnd.n1172 gnd.n1171 0.152939
R21675 gnd.n1173 gnd.n1172 0.152939
R21676 gnd.n1192 gnd.n1173 0.152939
R21677 gnd.n1193 gnd.n1192 0.152939
R21678 gnd.n1194 gnd.n1193 0.152939
R21679 gnd.n1195 gnd.n1194 0.152939
R21680 gnd.n1212 gnd.n1195 0.152939
R21681 gnd.n1213 gnd.n1212 0.152939
R21682 gnd.n1214 gnd.n1213 0.152939
R21683 gnd.n1215 gnd.n1214 0.152939
R21684 gnd.n1234 gnd.n1215 0.152939
R21685 gnd.n1235 gnd.n1234 0.152939
R21686 gnd.n1236 gnd.n1235 0.152939
R21687 gnd.n1237 gnd.n1236 0.152939
R21688 gnd.n1255 gnd.n1237 0.152939
R21689 gnd.n1256 gnd.n1255 0.152939
R21690 gnd.n1257 gnd.n1256 0.152939
R21691 gnd.n1258 gnd.n1257 0.152939
R21692 gnd.n1275 gnd.n1258 0.152939
R21693 gnd.n4591 gnd.n1275 0.152939
R21694 gnd.n4750 gnd.n1008 0.152939
R21695 gnd.n4750 gnd.n4749 0.152939
R21696 gnd.n4749 gnd.n4748 0.152939
R21697 gnd.n4748 gnd.n1011 0.152939
R21698 gnd.n2414 gnd.n1011 0.152939
R21699 gnd.n2418 gnd.n2414 0.152939
R21700 gnd.n2419 gnd.n2418 0.152939
R21701 gnd.n2420 gnd.n2419 0.152939
R21702 gnd.n2420 gnd.n2412 0.152939
R21703 gnd.n2426 gnd.n2412 0.152939
R21704 gnd.n2427 gnd.n2426 0.152939
R21705 gnd.n2428 gnd.n2427 0.152939
R21706 gnd.n2428 gnd.n2410 0.152939
R21707 gnd.n2434 gnd.n2410 0.152939
R21708 gnd.n2435 gnd.n2434 0.152939
R21709 gnd.n2436 gnd.n2435 0.152939
R21710 gnd.n2436 gnd.n2408 0.152939
R21711 gnd.n2442 gnd.n2408 0.152939
R21712 gnd.n2443 gnd.n2442 0.152939
R21713 gnd.n2444 gnd.n2443 0.152939
R21714 gnd.n2444 gnd.n2406 0.152939
R21715 gnd.n2582 gnd.n2406 0.152939
R21716 gnd.n2583 gnd.n2582 0.152939
R21717 gnd.n2584 gnd.n2583 0.152939
R21718 gnd.n2585 gnd.n2584 0.152939
R21719 gnd.n2586 gnd.n2585 0.152939
R21720 gnd.n2605 gnd.n2604 0.152939
R21721 gnd.n2606 gnd.n2605 0.152939
R21722 gnd.n2607 gnd.n2606 0.152939
R21723 gnd.n2607 gnd.n2358 0.152939
R21724 gnd.n2655 gnd.n2358 0.152939
R21725 gnd.n2656 gnd.n2655 0.152939
R21726 gnd.n2658 gnd.n2656 0.152939
R21727 gnd.n2658 gnd.n2657 0.152939
R21728 gnd.n2657 gnd.n2352 0.152939
R21729 gnd.n2352 gnd.n2350 0.152939
R21730 gnd.n2674 gnd.n2350 0.152939
R21731 gnd.n2675 gnd.n2674 0.152939
R21732 gnd.n2676 gnd.n2675 0.152939
R21733 gnd.n2676 gnd.n2348 0.152939
R21734 gnd.n2685 gnd.n2348 0.152939
R21735 gnd.n2686 gnd.n2685 0.152939
R21736 gnd.n2687 gnd.n2686 0.152939
R21737 gnd.n2688 gnd.n2687 0.152939
R21738 gnd.n2689 gnd.n2688 0.152939
R21739 gnd.n2689 gnd.n2322 0.152939
R21740 gnd.n2775 gnd.n2322 0.152939
R21741 gnd.n2776 gnd.n2775 0.152939
R21742 gnd.n2778 gnd.n2776 0.152939
R21743 gnd.n2778 gnd.n2777 0.152939
R21744 gnd.n2777 gnd.n2314 0.152939
R21745 gnd.n2825 gnd.n2314 0.152939
R21746 gnd.n966 gnd.n965 0.152939
R21747 gnd.n967 gnd.n966 0.152939
R21748 gnd.n968 gnd.n967 0.152939
R21749 gnd.n969 gnd.n968 0.152939
R21750 gnd.n970 gnd.n969 0.152939
R21751 gnd.n971 gnd.n970 0.152939
R21752 gnd.n972 gnd.n971 0.152939
R21753 gnd.n973 gnd.n972 0.152939
R21754 gnd.n974 gnd.n973 0.152939
R21755 gnd.n975 gnd.n974 0.152939
R21756 gnd.n976 gnd.n975 0.152939
R21757 gnd.n977 gnd.n976 0.152939
R21758 gnd.n978 gnd.n977 0.152939
R21759 gnd.n979 gnd.n978 0.152939
R21760 gnd.n980 gnd.n979 0.152939
R21761 gnd.n981 gnd.n980 0.152939
R21762 gnd.n982 gnd.n981 0.152939
R21763 gnd.n985 gnd.n982 0.152939
R21764 gnd.n986 gnd.n985 0.152939
R21765 gnd.n987 gnd.n986 0.152939
R21766 gnd.n988 gnd.n987 0.152939
R21767 gnd.n989 gnd.n988 0.152939
R21768 gnd.n990 gnd.n989 0.152939
R21769 gnd.n991 gnd.n990 0.152939
R21770 gnd.n992 gnd.n991 0.152939
R21771 gnd.n993 gnd.n992 0.152939
R21772 gnd.n994 gnd.n993 0.152939
R21773 gnd.n995 gnd.n994 0.152939
R21774 gnd.n996 gnd.n995 0.152939
R21775 gnd.n997 gnd.n996 0.152939
R21776 gnd.n998 gnd.n997 0.152939
R21777 gnd.n999 gnd.n998 0.152939
R21778 gnd.n1000 gnd.n999 0.152939
R21779 gnd.n1001 gnd.n1000 0.152939
R21780 gnd.n1002 gnd.n1001 0.152939
R21781 gnd.n4758 gnd.n1002 0.152939
R21782 gnd.n4758 gnd.n4757 0.152939
R21783 gnd.n4757 gnd.n4756 0.152939
R21784 gnd.n2532 gnd.n2530 0.152939
R21785 gnd.n2532 gnd.n2531 0.152939
R21786 gnd.n2531 gnd.n1022 0.152939
R21787 gnd.n1023 gnd.n1022 0.152939
R21788 gnd.n1024 gnd.n1023 0.152939
R21789 gnd.n1042 gnd.n1024 0.152939
R21790 gnd.n1043 gnd.n1042 0.152939
R21791 gnd.n1044 gnd.n1043 0.152939
R21792 gnd.n1045 gnd.n1044 0.152939
R21793 gnd.n1061 gnd.n1045 0.152939
R21794 gnd.n1062 gnd.n1061 0.152939
R21795 gnd.n1063 gnd.n1062 0.152939
R21796 gnd.n1064 gnd.n1063 0.152939
R21797 gnd.n1082 gnd.n1064 0.152939
R21798 gnd.n1083 gnd.n1082 0.152939
R21799 gnd.n1084 gnd.n1083 0.152939
R21800 gnd.n1085 gnd.n1084 0.152939
R21801 gnd.n1103 gnd.n1085 0.152939
R21802 gnd.n1104 gnd.n1103 0.152939
R21803 gnd.n1105 gnd.n1104 0.152939
R21804 gnd.n1106 gnd.n1105 0.152939
R21805 gnd.n2394 gnd.n2390 0.152939
R21806 gnd.n2638 gnd.n2390 0.152939
R21807 gnd.n731 gnd.n726 0.152939
R21808 gnd.n732 gnd.n731 0.152939
R21809 gnd.n733 gnd.n732 0.152939
R21810 gnd.n738 gnd.n733 0.152939
R21811 gnd.n739 gnd.n738 0.152939
R21812 gnd.n740 gnd.n739 0.152939
R21813 gnd.n741 gnd.n740 0.152939
R21814 gnd.n746 gnd.n741 0.152939
R21815 gnd.n747 gnd.n746 0.152939
R21816 gnd.n748 gnd.n747 0.152939
R21817 gnd.n749 gnd.n748 0.152939
R21818 gnd.n754 gnd.n749 0.152939
R21819 gnd.n755 gnd.n754 0.152939
R21820 gnd.n756 gnd.n755 0.152939
R21821 gnd.n757 gnd.n756 0.152939
R21822 gnd.n762 gnd.n757 0.152939
R21823 gnd.n763 gnd.n762 0.152939
R21824 gnd.n764 gnd.n763 0.152939
R21825 gnd.n765 gnd.n764 0.152939
R21826 gnd.n770 gnd.n765 0.152939
R21827 gnd.n771 gnd.n770 0.152939
R21828 gnd.n772 gnd.n771 0.152939
R21829 gnd.n773 gnd.n772 0.152939
R21830 gnd.n778 gnd.n773 0.152939
R21831 gnd.n779 gnd.n778 0.152939
R21832 gnd.n780 gnd.n779 0.152939
R21833 gnd.n781 gnd.n780 0.152939
R21834 gnd.n786 gnd.n781 0.152939
R21835 gnd.n787 gnd.n786 0.152939
R21836 gnd.n788 gnd.n787 0.152939
R21837 gnd.n789 gnd.n788 0.152939
R21838 gnd.n794 gnd.n789 0.152939
R21839 gnd.n795 gnd.n794 0.152939
R21840 gnd.n796 gnd.n795 0.152939
R21841 gnd.n797 gnd.n796 0.152939
R21842 gnd.n802 gnd.n797 0.152939
R21843 gnd.n803 gnd.n802 0.152939
R21844 gnd.n804 gnd.n803 0.152939
R21845 gnd.n805 gnd.n804 0.152939
R21846 gnd.n810 gnd.n805 0.152939
R21847 gnd.n811 gnd.n810 0.152939
R21848 gnd.n812 gnd.n811 0.152939
R21849 gnd.n813 gnd.n812 0.152939
R21850 gnd.n818 gnd.n813 0.152939
R21851 gnd.n819 gnd.n818 0.152939
R21852 gnd.n820 gnd.n819 0.152939
R21853 gnd.n821 gnd.n820 0.152939
R21854 gnd.n826 gnd.n821 0.152939
R21855 gnd.n827 gnd.n826 0.152939
R21856 gnd.n828 gnd.n827 0.152939
R21857 gnd.n829 gnd.n828 0.152939
R21858 gnd.n834 gnd.n829 0.152939
R21859 gnd.n835 gnd.n834 0.152939
R21860 gnd.n836 gnd.n835 0.152939
R21861 gnd.n837 gnd.n836 0.152939
R21862 gnd.n842 gnd.n837 0.152939
R21863 gnd.n843 gnd.n842 0.152939
R21864 gnd.n844 gnd.n843 0.152939
R21865 gnd.n845 gnd.n844 0.152939
R21866 gnd.n850 gnd.n845 0.152939
R21867 gnd.n851 gnd.n850 0.152939
R21868 gnd.n852 gnd.n851 0.152939
R21869 gnd.n853 gnd.n852 0.152939
R21870 gnd.n858 gnd.n853 0.152939
R21871 gnd.n859 gnd.n858 0.152939
R21872 gnd.n860 gnd.n859 0.152939
R21873 gnd.n861 gnd.n860 0.152939
R21874 gnd.n866 gnd.n861 0.152939
R21875 gnd.n867 gnd.n866 0.152939
R21876 gnd.n868 gnd.n867 0.152939
R21877 gnd.n869 gnd.n868 0.152939
R21878 gnd.n874 gnd.n869 0.152939
R21879 gnd.n875 gnd.n874 0.152939
R21880 gnd.n876 gnd.n875 0.152939
R21881 gnd.n877 gnd.n876 0.152939
R21882 gnd.n882 gnd.n877 0.152939
R21883 gnd.n883 gnd.n882 0.152939
R21884 gnd.n884 gnd.n883 0.152939
R21885 gnd.n885 gnd.n884 0.152939
R21886 gnd.n890 gnd.n885 0.152939
R21887 gnd.n891 gnd.n890 0.152939
R21888 gnd.n892 gnd.n891 0.152939
R21889 gnd.n893 gnd.n892 0.152939
R21890 gnd.n2393 gnd.n893 0.152939
R21891 gnd.n4154 gnd.n1684 0.152939
R21892 gnd.n4150 gnd.n1684 0.152939
R21893 gnd.n4150 gnd.n4149 0.152939
R21894 gnd.n4149 gnd.n4148 0.152939
R21895 gnd.n4148 gnd.n1812 0.152939
R21896 gnd.n4141 gnd.n1812 0.152939
R21897 gnd.n4141 gnd.n4140 0.152939
R21898 gnd.n4140 gnd.n4139 0.152939
R21899 gnd.n4139 gnd.n4132 0.152939
R21900 gnd.n3726 gnd.n3725 0.152939
R21901 gnd.n3726 gnd.n2149 0.152939
R21902 gnd.n3740 gnd.n2149 0.152939
R21903 gnd.n3741 gnd.n3740 0.152939
R21904 gnd.n3742 gnd.n3741 0.152939
R21905 gnd.n3742 gnd.n2136 0.152939
R21906 gnd.n3756 gnd.n2136 0.152939
R21907 gnd.n3757 gnd.n3756 0.152939
R21908 gnd.n3758 gnd.n3757 0.152939
R21909 gnd.n3758 gnd.n2123 0.152939
R21910 gnd.n3772 gnd.n2123 0.152939
R21911 gnd.n3773 gnd.n3772 0.152939
R21912 gnd.n3774 gnd.n3773 0.152939
R21913 gnd.n3774 gnd.n2110 0.152939
R21914 gnd.n3788 gnd.n2110 0.152939
R21915 gnd.n3789 gnd.n3788 0.152939
R21916 gnd.n3790 gnd.n3789 0.152939
R21917 gnd.n3790 gnd.n2096 0.152939
R21918 gnd.n3804 gnd.n2096 0.152939
R21919 gnd.n3805 gnd.n3804 0.152939
R21920 gnd.n3806 gnd.n3805 0.152939
R21921 gnd.n3806 gnd.n2083 0.152939
R21922 gnd.n3820 gnd.n2083 0.152939
R21923 gnd.n3821 gnd.n3820 0.152939
R21924 gnd.n3822 gnd.n3821 0.152939
R21925 gnd.n3822 gnd.n2070 0.152939
R21926 gnd.n3836 gnd.n2070 0.152939
R21927 gnd.n3837 gnd.n3836 0.152939
R21928 gnd.n3838 gnd.n3837 0.152939
R21929 gnd.n3838 gnd.n2055 0.152939
R21930 gnd.n3852 gnd.n2055 0.152939
R21931 gnd.n3853 gnd.n3852 0.152939
R21932 gnd.n3854 gnd.n3853 0.152939
R21933 gnd.n3854 gnd.n2041 0.152939
R21934 gnd.n3868 gnd.n2041 0.152939
R21935 gnd.n3869 gnd.n3868 0.152939
R21936 gnd.n3870 gnd.n3869 0.152939
R21937 gnd.n3870 gnd.n2028 0.152939
R21938 gnd.n3884 gnd.n2028 0.152939
R21939 gnd.n3885 gnd.n3884 0.152939
R21940 gnd.n3886 gnd.n3885 0.152939
R21941 gnd.n3886 gnd.n2012 0.152939
R21942 gnd.n3900 gnd.n2012 0.152939
R21943 gnd.n3901 gnd.n3900 0.152939
R21944 gnd.n3902 gnd.n3901 0.152939
R21945 gnd.n3902 gnd.n1998 0.152939
R21946 gnd.n3916 gnd.n1998 0.152939
R21947 gnd.n3917 gnd.n3916 0.152939
R21948 gnd.n3918 gnd.n3917 0.152939
R21949 gnd.n3918 gnd.n1984 0.152939
R21950 gnd.n3932 gnd.n1984 0.152939
R21951 gnd.n3933 gnd.n3932 0.152939
R21952 gnd.n3934 gnd.n3933 0.152939
R21953 gnd.n3934 gnd.n1970 0.152939
R21954 gnd.n3948 gnd.n1970 0.152939
R21955 gnd.n3949 gnd.n3948 0.152939
R21956 gnd.n3950 gnd.n3949 0.152939
R21957 gnd.n3950 gnd.n1956 0.152939
R21958 gnd.n3964 gnd.n1956 0.152939
R21959 gnd.n3965 gnd.n3964 0.152939
R21960 gnd.n3966 gnd.n3965 0.152939
R21961 gnd.n3966 gnd.n1942 0.152939
R21962 gnd.n3980 gnd.n1942 0.152939
R21963 gnd.n3981 gnd.n3980 0.152939
R21964 gnd.n3982 gnd.n3981 0.152939
R21965 gnd.n3982 gnd.n1928 0.152939
R21966 gnd.n3996 gnd.n1928 0.152939
R21967 gnd.n3997 gnd.n3996 0.152939
R21968 gnd.n3998 gnd.n3997 0.152939
R21969 gnd.n3998 gnd.n1915 0.152939
R21970 gnd.n4012 gnd.n1915 0.152939
R21971 gnd.n4013 gnd.n4012 0.152939
R21972 gnd.n4014 gnd.n4013 0.152939
R21973 gnd.n4014 gnd.n1900 0.152939
R21974 gnd.n4028 gnd.n1900 0.152939
R21975 gnd.n4029 gnd.n4028 0.152939
R21976 gnd.n4030 gnd.n4029 0.152939
R21977 gnd.n4030 gnd.n1886 0.152939
R21978 gnd.n4044 gnd.n1886 0.152939
R21979 gnd.n4045 gnd.n4044 0.152939
R21980 gnd.n4046 gnd.n4045 0.152939
R21981 gnd.n4046 gnd.n1874 0.152939
R21982 gnd.n4060 gnd.n1874 0.152939
R21983 gnd.n4061 gnd.n4060 0.152939
R21984 gnd.n4062 gnd.n4061 0.152939
R21985 gnd.n4062 gnd.n1861 0.152939
R21986 gnd.n4076 gnd.n1861 0.152939
R21987 gnd.n4077 gnd.n4076 0.152939
R21988 gnd.n4078 gnd.n4077 0.152939
R21989 gnd.n4078 gnd.n1848 0.152939
R21990 gnd.n4092 gnd.n1848 0.152939
R21991 gnd.n4093 gnd.n4092 0.152939
R21992 gnd.n4094 gnd.n4093 0.152939
R21993 gnd.n4094 gnd.n1835 0.152939
R21994 gnd.n4108 gnd.n1835 0.152939
R21995 gnd.n4109 gnd.n4108 0.152939
R21996 gnd.n4112 gnd.n4109 0.152939
R21997 gnd.n4112 gnd.n4111 0.152939
R21998 gnd.n4111 gnd.n4110 0.152939
R21999 gnd.n4110 gnd.n1820 0.152939
R22000 gnd.n4131 gnd.n1820 0.152939
R22001 gnd.n2811 gnd.n2786 0.152939
R22002 gnd.n2811 gnd.n2810 0.152939
R22003 gnd.n2810 gnd.n2809 0.152939
R22004 gnd.n2809 gnd.n2792 0.152939
R22005 gnd.n2805 gnd.n2792 0.152939
R22006 gnd.n2805 gnd.n2804 0.152939
R22007 gnd.n2804 gnd.n2799 0.152939
R22008 gnd.n2799 gnd.n2162 0.152939
R22009 gnd.n3724 gnd.n2162 0.152939
R22010 gnd.n2617 gnd.n2616 0.152939
R22011 gnd.n2616 gnd.n2361 0.152939
R22012 gnd.n2647 gnd.n2361 0.152939
R22013 gnd.n2648 gnd.n2647 0.152939
R22014 gnd.n2649 gnd.n2648 0.152939
R22015 gnd.n2649 gnd.n2354 0.152939
R22016 gnd.n2664 gnd.n2354 0.152939
R22017 gnd.n2665 gnd.n2664 0.152939
R22018 gnd.n2666 gnd.n2665 0.152939
R22019 gnd.n2666 gnd.n2342 0.152939
R22020 gnd.n2705 gnd.n2342 0.152939
R22021 gnd.n2705 gnd.n2704 0.152939
R22022 gnd.n2704 gnd.n2703 0.152939
R22023 gnd.n2703 gnd.n2343 0.152939
R22024 gnd.n2699 gnd.n2343 0.152939
R22025 gnd.n2699 gnd.n2698 0.152939
R22026 gnd.n2698 gnd.n2697 0.152939
R22027 gnd.n2697 gnd.n2325 0.152939
R22028 gnd.n2767 gnd.n2325 0.152939
R22029 gnd.n2768 gnd.n2767 0.152939
R22030 gnd.n2769 gnd.n2768 0.152939
R22031 gnd.n2769 gnd.n2319 0.152939
R22032 gnd.n2784 gnd.n2319 0.152939
R22033 gnd.n2785 gnd.n2784 0.152939
R22034 gnd.n2818 gnd.n2785 0.152939
R22035 gnd.n2818 gnd.n2817 0.152939
R22036 gnd.n4588 gnd.n1278 0.152939
R22037 gnd.n4584 gnd.n1278 0.152939
R22038 gnd.n4584 gnd.n4583 0.152939
R22039 gnd.n4583 gnd.n4582 0.152939
R22040 gnd.n4582 gnd.n1283 0.152939
R22041 gnd.n4578 gnd.n1283 0.152939
R22042 gnd.n4578 gnd.n4577 0.152939
R22043 gnd.n4577 gnd.n4576 0.152939
R22044 gnd.n4576 gnd.n1288 0.152939
R22045 gnd.n4572 gnd.n1288 0.152939
R22046 gnd.n4572 gnd.n4571 0.152939
R22047 gnd.n4571 gnd.n4570 0.152939
R22048 gnd.n4570 gnd.n1293 0.152939
R22049 gnd.n4566 gnd.n1293 0.152939
R22050 gnd.n4566 gnd.n4565 0.152939
R22051 gnd.n4565 gnd.n4564 0.152939
R22052 gnd.n4564 gnd.n1298 0.152939
R22053 gnd.n4560 gnd.n1298 0.152939
R22054 gnd.n4560 gnd.n4559 0.152939
R22055 gnd.n4559 gnd.n4558 0.152939
R22056 gnd.n4558 gnd.n1303 0.152939
R22057 gnd.n4554 gnd.n1303 0.152939
R22058 gnd.n4554 gnd.n4553 0.152939
R22059 gnd.n4553 gnd.n4552 0.152939
R22060 gnd.n4552 gnd.n1308 0.152939
R22061 gnd.n4548 gnd.n1308 0.152939
R22062 gnd.n4548 gnd.n4547 0.152939
R22063 gnd.n4547 gnd.n4546 0.152939
R22064 gnd.n4546 gnd.n1313 0.152939
R22065 gnd.n4542 gnd.n1313 0.152939
R22066 gnd.n4542 gnd.n4541 0.152939
R22067 gnd.n4541 gnd.n4540 0.152939
R22068 gnd.n4540 gnd.n1318 0.152939
R22069 gnd.n4536 gnd.n1318 0.152939
R22070 gnd.n4536 gnd.n4535 0.152939
R22071 gnd.n4535 gnd.n4534 0.152939
R22072 gnd.n4534 gnd.n1323 0.152939
R22073 gnd.n4530 gnd.n1323 0.152939
R22074 gnd.n4530 gnd.n4529 0.152939
R22075 gnd.n4529 gnd.n4528 0.152939
R22076 gnd.n4528 gnd.n1328 0.152939
R22077 gnd.n4524 gnd.n1328 0.152939
R22078 gnd.n4524 gnd.n4523 0.152939
R22079 gnd.n4523 gnd.n4522 0.152939
R22080 gnd.n4522 gnd.n1333 0.152939
R22081 gnd.n4518 gnd.n1333 0.152939
R22082 gnd.n4518 gnd.n4517 0.152939
R22083 gnd.n4517 gnd.n4516 0.152939
R22084 gnd.n4516 gnd.n1338 0.152939
R22085 gnd.n4512 gnd.n1338 0.152939
R22086 gnd.n4512 gnd.n4511 0.152939
R22087 gnd.n4511 gnd.n4510 0.152939
R22088 gnd.n4510 gnd.n1343 0.152939
R22089 gnd.n4506 gnd.n1343 0.152939
R22090 gnd.n4506 gnd.n4505 0.152939
R22091 gnd.n4505 gnd.n4504 0.152939
R22092 gnd.n4504 gnd.n1348 0.152939
R22093 gnd.n4500 gnd.n1348 0.152939
R22094 gnd.n4500 gnd.n4499 0.152939
R22095 gnd.n4499 gnd.n4498 0.152939
R22096 gnd.n4498 gnd.n1353 0.152939
R22097 gnd.n4494 gnd.n1353 0.152939
R22098 gnd.n4494 gnd.n4493 0.152939
R22099 gnd.n4493 gnd.n4492 0.152939
R22100 gnd.n4492 gnd.n1358 0.152939
R22101 gnd.n4488 gnd.n1358 0.152939
R22102 gnd.n4488 gnd.n4487 0.152939
R22103 gnd.n4487 gnd.n4486 0.152939
R22104 gnd.n4486 gnd.n1363 0.152939
R22105 gnd.n4482 gnd.n1363 0.152939
R22106 gnd.n4482 gnd.n4481 0.152939
R22107 gnd.n4481 gnd.n4480 0.152939
R22108 gnd.n4480 gnd.n1368 0.152939
R22109 gnd.n4476 gnd.n1368 0.152939
R22110 gnd.n4476 gnd.n4475 0.152939
R22111 gnd.n4475 gnd.n4474 0.152939
R22112 gnd.n4474 gnd.n1373 0.152939
R22113 gnd.n4470 gnd.n1373 0.152939
R22114 gnd.n4470 gnd.n4469 0.152939
R22115 gnd.n4469 gnd.n4468 0.152939
R22116 gnd.n4468 gnd.n1378 0.152939
R22117 gnd.n4464 gnd.n1378 0.152939
R22118 gnd.n4464 gnd.n4463 0.152939
R22119 gnd.n4463 gnd.n4462 0.152939
R22120 gnd.n4462 gnd.n1383 0.152939
R22121 gnd.n4458 gnd.n1383 0.152939
R22122 gnd.n4458 gnd.n4457 0.152939
R22123 gnd.n4457 gnd.n4456 0.152939
R22124 gnd.n4456 gnd.n1388 0.152939
R22125 gnd.n4452 gnd.n1388 0.152939
R22126 gnd.n4452 gnd.n4451 0.152939
R22127 gnd.n4451 gnd.n4450 0.152939
R22128 gnd.n4450 gnd.n1393 0.152939
R22129 gnd.n4446 gnd.n1393 0.152939
R22130 gnd.n4446 gnd.n4445 0.152939
R22131 gnd.n4445 gnd.n4444 0.152939
R22132 gnd.n4444 gnd.n1398 0.152939
R22133 gnd.n4440 gnd.n1398 0.152939
R22134 gnd.n4440 gnd.n4439 0.152939
R22135 gnd.n4439 gnd.n4438 0.152939
R22136 gnd.n4438 gnd.n1403 0.152939
R22137 gnd.n4346 gnd.n4345 0.152939
R22138 gnd.n4345 gnd.n4344 0.152939
R22139 gnd.n4344 gnd.n1504 0.152939
R22140 gnd.n4340 gnd.n1504 0.152939
R22141 gnd.n4340 gnd.n4339 0.152939
R22142 gnd.n4339 gnd.n4338 0.152939
R22143 gnd.n4338 gnd.n1509 0.152939
R22144 gnd.n4334 gnd.n1509 0.152939
R22145 gnd.n4334 gnd.n4333 0.152939
R22146 gnd.n4333 gnd.n4332 0.152939
R22147 gnd.n4332 gnd.n1514 0.152939
R22148 gnd.n4328 gnd.n1514 0.152939
R22149 gnd.n4328 gnd.n4327 0.152939
R22150 gnd.n4327 gnd.n4326 0.152939
R22151 gnd.n4326 gnd.n1519 0.152939
R22152 gnd.n4322 gnd.n1519 0.152939
R22153 gnd.n4322 gnd.n4321 0.152939
R22154 gnd.n4321 gnd.n4320 0.152939
R22155 gnd.n4320 gnd.n1524 0.152939
R22156 gnd.n4316 gnd.n1524 0.152939
R22157 gnd.n4316 gnd.n285 0.152939
R22158 gnd.n7216 gnd.n285 0.152939
R22159 gnd.n7216 gnd.n7215 0.152939
R22160 gnd.n7215 gnd.n7214 0.152939
R22161 gnd.n7214 gnd.n286 0.152939
R22162 gnd.n7210 gnd.n286 0.152939
R22163 gnd.n7208 gnd.n7207 0.152939
R22164 gnd.n7207 gnd.n292 0.152939
R22165 gnd.n292 gnd.n260 0.152939
R22166 gnd.n7229 gnd.n260 0.152939
R22167 gnd.n7230 gnd.n7229 0.152939
R22168 gnd.n7231 gnd.n7230 0.152939
R22169 gnd.n7231 gnd.n244 0.152939
R22170 gnd.n7245 gnd.n244 0.152939
R22171 gnd.n7246 gnd.n7245 0.152939
R22172 gnd.n7247 gnd.n7246 0.152939
R22173 gnd.n7247 gnd.n229 0.152939
R22174 gnd.n7261 gnd.n229 0.152939
R22175 gnd.n7262 gnd.n7261 0.152939
R22176 gnd.n7263 gnd.n7262 0.152939
R22177 gnd.n7263 gnd.n214 0.152939
R22178 gnd.n7277 gnd.n214 0.152939
R22179 gnd.n7278 gnd.n7277 0.152939
R22180 gnd.n7279 gnd.n7278 0.152939
R22181 gnd.n7279 gnd.n199 0.152939
R22182 gnd.n7293 gnd.n199 0.152939
R22183 gnd.n7294 gnd.n7293 0.152939
R22184 gnd.n7370 gnd.n7294 0.152939
R22185 gnd.n7370 gnd.n7369 0.152939
R22186 gnd.n7369 gnd.n7368 0.152939
R22187 gnd.n7368 gnd.n7295 0.152939
R22188 gnd.n7364 gnd.n7295 0.152939
R22189 gnd.n7363 gnd.n7297 0.152939
R22190 gnd.n7359 gnd.n7297 0.152939
R22191 gnd.n7359 gnd.n7358 0.152939
R22192 gnd.n7358 gnd.n7357 0.152939
R22193 gnd.n7357 gnd.n7303 0.152939
R22194 gnd.n7353 gnd.n7303 0.152939
R22195 gnd.n7353 gnd.n7352 0.152939
R22196 gnd.n7352 gnd.n7351 0.152939
R22197 gnd.n7351 gnd.n7311 0.152939
R22198 gnd.n7347 gnd.n7311 0.152939
R22199 gnd.n7347 gnd.n7346 0.152939
R22200 gnd.n7346 gnd.n7345 0.152939
R22201 gnd.n7345 gnd.n7319 0.152939
R22202 gnd.n7341 gnd.n7319 0.152939
R22203 gnd.n7341 gnd.n7340 0.152939
R22204 gnd.n7340 gnd.n7339 0.152939
R22205 gnd.n7339 gnd.n7327 0.152939
R22206 gnd.n7335 gnd.n7327 0.152939
R22207 gnd.n4158 gnd.n4157 0.152939
R22208 gnd.n4160 gnd.n4158 0.152939
R22209 gnd.n4160 gnd.n4159 0.152939
R22210 gnd.n4159 gnd.n1612 0.152939
R22211 gnd.n4188 gnd.n1612 0.152939
R22212 gnd.n4189 gnd.n4188 0.152939
R22213 gnd.n4191 gnd.n4189 0.152939
R22214 gnd.n4191 gnd.n4190 0.152939
R22215 gnd.n4190 gnd.n1585 0.152939
R22216 gnd.n4219 gnd.n1585 0.152939
R22217 gnd.n4220 gnd.n4219 0.152939
R22218 gnd.n4227 gnd.n4220 0.152939
R22219 gnd.n4227 gnd.n4226 0.152939
R22220 gnd.n4226 gnd.n4225 0.152939
R22221 gnd.n4225 gnd.n4221 0.152939
R22222 gnd.n4221 gnd.n1551 0.152939
R22223 gnd.n4284 gnd.n1551 0.152939
R22224 gnd.n4284 gnd.n4283 0.152939
R22225 gnd.n4283 gnd.n4282 0.152939
R22226 gnd.n4282 gnd.n1552 0.152939
R22227 gnd.n4278 gnd.n1552 0.152939
R22228 gnd.n4278 gnd.n310 0.152939
R22229 gnd.n7122 gnd.n310 0.152939
R22230 gnd.n7123 gnd.n7122 0.152939
R22231 gnd.n7124 gnd.n7123 0.152939
R22232 gnd.n7124 gnd.n67 0.152939
R22233 gnd.n7502 gnd.n68 0.152939
R22234 gnd.n7498 gnd.n68 0.152939
R22235 gnd.n7498 gnd.n7497 0.152939
R22236 gnd.n7497 gnd.n7496 0.152939
R22237 gnd.n7496 gnd.n74 0.152939
R22238 gnd.n7492 gnd.n74 0.152939
R22239 gnd.n7492 gnd.n7491 0.152939
R22240 gnd.n7491 gnd.n7490 0.152939
R22241 gnd.n7490 gnd.n79 0.152939
R22242 gnd.n7486 gnd.n79 0.152939
R22243 gnd.n7486 gnd.n7485 0.152939
R22244 gnd.n7485 gnd.n7484 0.152939
R22245 gnd.n7484 gnd.n84 0.152939
R22246 gnd.n7480 gnd.n84 0.152939
R22247 gnd.n7480 gnd.n7479 0.152939
R22248 gnd.n7479 gnd.n7478 0.152939
R22249 gnd.n7478 gnd.n89 0.152939
R22250 gnd.n7474 gnd.n89 0.152939
R22251 gnd.n7474 gnd.n7473 0.152939
R22252 gnd.n7473 gnd.n7472 0.152939
R22253 gnd.n7472 gnd.n94 0.152939
R22254 gnd.n7468 gnd.n94 0.152939
R22255 gnd.n7468 gnd.n7467 0.152939
R22256 gnd.n7467 gnd.n7466 0.152939
R22257 gnd.n7466 gnd.n99 0.152939
R22258 gnd.n102 gnd.n99 0.152939
R22259 gnd.n4155 gnd.n4154 0.151415
R22260 gnd.n2816 gnd.n2786 0.151415
R22261 gnd.n2639 gnd.n2385 0.140744
R22262 gnd.n4296 gnd.n269 0.140744
R22263 gnd.n5462 gnd.n5019 0.0767195
R22264 gnd.n5462 gnd.n5398 0.0767195
R22265 gnd.n7223 gnd.n253 0.0767195
R22266 gnd.n300 gnd.n291 0.0767195
R22267 gnd.n7136 gnd.n291 0.0767195
R22268 gnd.n7223 gnd.n268 0.0767195
R22269 gnd.n1162 gnd.n1125 0.0767195
R22270 gnd.n2602 gnd.n1134 0.0767195
R22271 gnd.n2602 gnd.n1135 0.0767195
R22272 gnd.n2603 gnd.n2586 0.0767195
R22273 gnd.n2604 gnd.n2603 0.0767195
R22274 gnd.n1125 gnd.n1106 0.0767195
R22275 gnd.n7210 gnd.n7209 0.0767195
R22276 gnd.n7209 gnd.n7208 0.0767195
R22277 gnd.n7503 gnd.n67 0.0767195
R22278 gnd.n7503 gnd.n7502 0.0767195
R22279 gnd.n2615 gnd.n2601 0.0695946
R22280 gnd.n2617 gnd.n2615 0.0695946
R22281 gnd.n4590 gnd.n4589 0.063
R22282 gnd.n1723 gnd.n1503 0.063
R22283 gnd.n6201 gnd.n4868 0.0477147
R22284 gnd.n5353 gnd.n5241 0.0442063
R22285 gnd.n5354 gnd.n5353 0.0442063
R22286 gnd.n5355 gnd.n5354 0.0442063
R22287 gnd.n5355 gnd.n5230 0.0442063
R22288 gnd.n5369 gnd.n5230 0.0442063
R22289 gnd.n5370 gnd.n5369 0.0442063
R22290 gnd.n5371 gnd.n5370 0.0442063
R22291 gnd.n5371 gnd.n5217 0.0442063
R22292 gnd.n5501 gnd.n5217 0.0442063
R22293 gnd.n5502 gnd.n5501 0.0442063
R22294 gnd.n5504 gnd.n5151 0.0344674
R22295 gnd.n1802 gnd.n1683 0.0343753
R22296 gnd.n2815 gnd.n2232 0.0343753
R22297 gnd.n5524 gnd.n5523 0.0269946
R22298 gnd.n5526 gnd.n5525 0.0269946
R22299 gnd.n5146 gnd.n5144 0.0269946
R22300 gnd.n5536 gnd.n5534 0.0269946
R22301 gnd.n5535 gnd.n5125 0.0269946
R22302 gnd.n5555 gnd.n5554 0.0269946
R22303 gnd.n5557 gnd.n5556 0.0269946
R22304 gnd.n5120 gnd.n5118 0.0269946
R22305 gnd.n5567 gnd.n5565 0.0269946
R22306 gnd.n5566 gnd.n5101 0.0269946
R22307 gnd.n5586 gnd.n5585 0.0269946
R22308 gnd.n5588 gnd.n5587 0.0269946
R22309 gnd.n5095 gnd.n5093 0.0269946
R22310 gnd.n5598 gnd.n5596 0.0269946
R22311 gnd.n5597 gnd.n5075 0.0269946
R22312 gnd.n5617 gnd.n5616 0.0269946
R22313 gnd.n5619 gnd.n5618 0.0269946
R22314 gnd.n5069 gnd.n5067 0.0269946
R22315 gnd.n5629 gnd.n5627 0.0269946
R22316 gnd.n5628 gnd.n5050 0.0269946
R22317 gnd.n5648 gnd.n5647 0.0269946
R22318 gnd.n5650 gnd.n5649 0.0269946
R22319 gnd.n5044 gnd.n5042 0.0269946
R22320 gnd.n5660 gnd.n5658 0.0269946
R22321 gnd.n5659 gnd.n5026 0.0269946
R22322 gnd.n5678 gnd.n5677 0.0269946
R22323 gnd.n5680 gnd.n5679 0.0269946
R22324 gnd.n5014 gnd.n5013 0.0269946
R22325 gnd.n5714 gnd.n5010 0.0269946
R22326 gnd.n5713 gnd.n5011 0.0269946
R22327 gnd.n5733 gnd.n4993 0.0269946
R22328 gnd.n5735 gnd.n5734 0.0269946
R22329 gnd.n5736 gnd.n4991 0.0269946
R22330 gnd.n5743 gnd.n5739 0.0269946
R22331 gnd.n5742 gnd.n5741 0.0269946
R22332 gnd.n5740 gnd.n4970 0.0269946
R22333 gnd.n5767 gnd.n4971 0.0269946
R22334 gnd.n5766 gnd.n4972 0.0269946
R22335 gnd.n5808 gnd.n4949 0.0269946
R22336 gnd.n5810 gnd.n5809 0.0269946
R22337 gnd.n5819 gnd.n4942 0.0269946
R22338 gnd.n5821 gnd.n5820 0.0269946
R22339 gnd.n5822 gnd.n4938 0.0269946
R22340 gnd.n6110 gnd.n4939 0.0269946
R22341 gnd.n6109 gnd.n4940 0.0269946
R22342 gnd.n5826 gnd.n902 0.0269946
R22343 gnd.n5827 gnd.n903 0.0269946
R22344 gnd.n5829 gnd.n904 0.0269946
R22345 gnd.n6089 gnd.n6088 0.0269946
R22346 gnd.n6090 gnd.n926 0.0269946
R22347 gnd.n6091 gnd.n927 0.0269946
R22348 gnd.n6092 gnd.n928 0.0269946
R22349 gnd.n1725 gnd.n1723 0.0245515
R22350 gnd.n4589 gnd.n1277 0.0245515
R22351 gnd.n5504 gnd.n5503 0.0202011
R22352 gnd.n1725 gnd.n1724 0.0174377
R22353 gnd.n1724 gnd.n1720 0.0174377
R22354 gnd.n1734 gnd.n1720 0.0174377
R22355 gnd.n1734 gnd.n1733 0.0174377
R22356 gnd.n1733 gnd.n1721 0.0174377
R22357 gnd.n1721 gnd.n1716 0.0174377
R22358 gnd.n1742 gnd.n1716 0.0174377
R22359 gnd.n1744 gnd.n1742 0.0174377
R22360 gnd.n1744 gnd.n1743 0.0174377
R22361 gnd.n1743 gnd.n1713 0.0174377
R22362 gnd.n1753 gnd.n1713 0.0174377
R22363 gnd.n1753 gnd.n1752 0.0174377
R22364 gnd.n1752 gnd.n1714 0.0174377
R22365 gnd.n1714 gnd.n1709 0.0174377
R22366 gnd.n1761 gnd.n1709 0.0174377
R22367 gnd.n1763 gnd.n1761 0.0174377
R22368 gnd.n1763 gnd.n1762 0.0174377
R22369 gnd.n1762 gnd.n1706 0.0174377
R22370 gnd.n1772 gnd.n1706 0.0174377
R22371 gnd.n1772 gnd.n1771 0.0174377
R22372 gnd.n1771 gnd.n1707 0.0174377
R22373 gnd.n1707 gnd.n1702 0.0174377
R22374 gnd.n1780 gnd.n1702 0.0174377
R22375 gnd.n1781 gnd.n1780 0.0174377
R22376 gnd.n1781 gnd.n1700 0.0174377
R22377 gnd.n1786 gnd.n1700 0.0174377
R22378 gnd.n1788 gnd.n1786 0.0174377
R22379 gnd.n1788 gnd.n1787 0.0174377
R22380 gnd.n1787 gnd.n1696 0.0174377
R22381 gnd.n1797 gnd.n1696 0.0174377
R22382 gnd.n1797 gnd.n1796 0.0174377
R22383 gnd.n1796 gnd.n1689 0.0174377
R22384 gnd.n1689 gnd.n1688 0.0174377
R22385 gnd.n1801 gnd.n1688 0.0174377
R22386 gnd.n1802 gnd.n1801 0.0174377
R22387 gnd.n2181 gnd.n1277 0.0174377
R22388 gnd.n2183 gnd.n2181 0.0174377
R22389 gnd.n3715 gnd.n2183 0.0174377
R22390 gnd.n3715 gnd.n3714 0.0174377
R22391 gnd.n3714 gnd.n2184 0.0174377
R22392 gnd.n3711 gnd.n2184 0.0174377
R22393 gnd.n3711 gnd.n3710 0.0174377
R22394 gnd.n3710 gnd.n2189 0.0174377
R22395 gnd.n3707 gnd.n2189 0.0174377
R22396 gnd.n3707 gnd.n3706 0.0174377
R22397 gnd.n3706 gnd.n2194 0.0174377
R22398 gnd.n3703 gnd.n2194 0.0174377
R22399 gnd.n3703 gnd.n3702 0.0174377
R22400 gnd.n3702 gnd.n2198 0.0174377
R22401 gnd.n3699 gnd.n2198 0.0174377
R22402 gnd.n3699 gnd.n3698 0.0174377
R22403 gnd.n3698 gnd.n2202 0.0174377
R22404 gnd.n3695 gnd.n2202 0.0174377
R22405 gnd.n3695 gnd.n3694 0.0174377
R22406 gnd.n3694 gnd.n2206 0.0174377
R22407 gnd.n3691 gnd.n2206 0.0174377
R22408 gnd.n3691 gnd.n3690 0.0174377
R22409 gnd.n3690 gnd.n2212 0.0174377
R22410 gnd.n3687 gnd.n2212 0.0174377
R22411 gnd.n3687 gnd.n3686 0.0174377
R22412 gnd.n3686 gnd.n2216 0.0174377
R22413 gnd.n3683 gnd.n2216 0.0174377
R22414 gnd.n3683 gnd.n3682 0.0174377
R22415 gnd.n3682 gnd.n2220 0.0174377
R22416 gnd.n3679 gnd.n2220 0.0174377
R22417 gnd.n3679 gnd.n3678 0.0174377
R22418 gnd.n3678 gnd.n2226 0.0174377
R22419 gnd.n3675 gnd.n2226 0.0174377
R22420 gnd.n3675 gnd.n3674 0.0174377
R22421 gnd.n3674 gnd.n2232 0.0174377
R22422 gnd.n5503 gnd.n5502 0.0148637
R22423 gnd.n6086 gnd.n5830 0.0144266
R22424 gnd.n6087 gnd.n6086 0.0130679
R22425 gnd.n326 gnd.n269 0.0126951
R22426 gnd.n2639 gnd.n2638 0.0126951
R22427 gnd.n5523 gnd.n5151 0.00797283
R22428 gnd.n5525 gnd.n5524 0.00797283
R22429 gnd.n5526 gnd.n5146 0.00797283
R22430 gnd.n5534 gnd.n5144 0.00797283
R22431 gnd.n5536 gnd.n5535 0.00797283
R22432 gnd.n5554 gnd.n5125 0.00797283
R22433 gnd.n5556 gnd.n5555 0.00797283
R22434 gnd.n5557 gnd.n5120 0.00797283
R22435 gnd.n5565 gnd.n5118 0.00797283
R22436 gnd.n5567 gnd.n5566 0.00797283
R22437 gnd.n5585 gnd.n5101 0.00797283
R22438 gnd.n5587 gnd.n5586 0.00797283
R22439 gnd.n5588 gnd.n5095 0.00797283
R22440 gnd.n5596 gnd.n5093 0.00797283
R22441 gnd.n5598 gnd.n5597 0.00797283
R22442 gnd.n5616 gnd.n5075 0.00797283
R22443 gnd.n5618 gnd.n5617 0.00797283
R22444 gnd.n5619 gnd.n5069 0.00797283
R22445 gnd.n5627 gnd.n5067 0.00797283
R22446 gnd.n5629 gnd.n5628 0.00797283
R22447 gnd.n5647 gnd.n5050 0.00797283
R22448 gnd.n5649 gnd.n5648 0.00797283
R22449 gnd.n5650 gnd.n5044 0.00797283
R22450 gnd.n5658 gnd.n5042 0.00797283
R22451 gnd.n5660 gnd.n5659 0.00797283
R22452 gnd.n5677 gnd.n5026 0.00797283
R22453 gnd.n5679 gnd.n5678 0.00797283
R22454 gnd.n5680 gnd.n5014 0.00797283
R22455 gnd.n5013 gnd.n5010 0.00797283
R22456 gnd.n5714 gnd.n5713 0.00797283
R22457 gnd.n5011 gnd.n4993 0.00797283
R22458 gnd.n5734 gnd.n5733 0.00797283
R22459 gnd.n5736 gnd.n5735 0.00797283
R22460 gnd.n5739 gnd.n4991 0.00797283
R22461 gnd.n5743 gnd.n5742 0.00797283
R22462 gnd.n5741 gnd.n5740 0.00797283
R22463 gnd.n4971 gnd.n4970 0.00797283
R22464 gnd.n5767 gnd.n5766 0.00797283
R22465 gnd.n4972 gnd.n4949 0.00797283
R22466 gnd.n5810 gnd.n5808 0.00797283
R22467 gnd.n5809 gnd.n4942 0.00797283
R22468 gnd.n5820 gnd.n5819 0.00797283
R22469 gnd.n5822 gnd.n5821 0.00797283
R22470 gnd.n4939 gnd.n4938 0.00797283
R22471 gnd.n6110 gnd.n6109 0.00797283
R22472 gnd.n5826 gnd.n4940 0.00797283
R22473 gnd.n5827 gnd.n902 0.00797283
R22474 gnd.n5829 gnd.n903 0.00797283
R22475 gnd.n5830 gnd.n904 0.00797283
R22476 gnd.n6088 gnd.n6087 0.00797283
R22477 gnd.n6090 gnd.n6089 0.00797283
R22478 gnd.n6091 gnd.n926 0.00797283
R22479 gnd.n6092 gnd.n927 0.00797283
R22480 gnd.n4868 gnd.n928 0.00797283
R22481 gnd.n7209 gnd.n291 0.00507153
R22482 gnd.n2603 gnd.n2602 0.00507153
R22483 gnd.n4155 gnd.n1683 0.000838753
R22484 gnd.n2816 gnd.n2815 0.000838753
R22485 diffpairibias.n0 diffpairibias.t27 436.822
R22486 diffpairibias.n27 diffpairibias.t24 435.479
R22487 diffpairibias.n26 diffpairibias.t21 435.479
R22488 diffpairibias.n25 diffpairibias.t22 435.479
R22489 diffpairibias.n24 diffpairibias.t26 435.479
R22490 diffpairibias.n23 diffpairibias.t20 435.479
R22491 diffpairibias.n0 diffpairibias.t23 435.479
R22492 diffpairibias.n1 diffpairibias.t28 435.479
R22493 diffpairibias.n2 diffpairibias.t25 435.479
R22494 diffpairibias.n3 diffpairibias.t29 435.479
R22495 diffpairibias.n13 diffpairibias.t14 377.536
R22496 diffpairibias.n13 diffpairibias.t0 376.193
R22497 diffpairibias.n14 diffpairibias.t10 376.193
R22498 diffpairibias.n15 diffpairibias.t12 376.193
R22499 diffpairibias.n16 diffpairibias.t6 376.193
R22500 diffpairibias.n17 diffpairibias.t2 376.193
R22501 diffpairibias.n18 diffpairibias.t16 376.193
R22502 diffpairibias.n19 diffpairibias.t4 376.193
R22503 diffpairibias.n20 diffpairibias.t18 376.193
R22504 diffpairibias.n21 diffpairibias.t8 376.193
R22505 diffpairibias.n4 diffpairibias.t15 113.368
R22506 diffpairibias.n4 diffpairibias.t1 112.698
R22507 diffpairibias.n5 diffpairibias.t11 112.698
R22508 diffpairibias.n6 diffpairibias.t13 112.698
R22509 diffpairibias.n7 diffpairibias.t7 112.698
R22510 diffpairibias.n8 diffpairibias.t3 112.698
R22511 diffpairibias.n9 diffpairibias.t17 112.698
R22512 diffpairibias.n10 diffpairibias.t5 112.698
R22513 diffpairibias.n11 diffpairibias.t19 112.698
R22514 diffpairibias.n12 diffpairibias.t9 112.698
R22515 diffpairibias.n22 diffpairibias.n21 4.77242
R22516 diffpairibias.n22 diffpairibias.n12 4.30807
R22517 diffpairibias.n23 diffpairibias.n22 4.13945
R22518 diffpairibias.n21 diffpairibias.n20 1.34352
R22519 diffpairibias.n20 diffpairibias.n19 1.34352
R22520 diffpairibias.n19 diffpairibias.n18 1.34352
R22521 diffpairibias.n18 diffpairibias.n17 1.34352
R22522 diffpairibias.n17 diffpairibias.n16 1.34352
R22523 diffpairibias.n16 diffpairibias.n15 1.34352
R22524 diffpairibias.n15 diffpairibias.n14 1.34352
R22525 diffpairibias.n14 diffpairibias.n13 1.34352
R22526 diffpairibias.n3 diffpairibias.n2 1.34352
R22527 diffpairibias.n2 diffpairibias.n1 1.34352
R22528 diffpairibias.n1 diffpairibias.n0 1.34352
R22529 diffpairibias.n24 diffpairibias.n23 1.34352
R22530 diffpairibias.n25 diffpairibias.n24 1.34352
R22531 diffpairibias.n26 diffpairibias.n25 1.34352
R22532 diffpairibias.n27 diffpairibias.n26 1.34352
R22533 diffpairibias.n28 diffpairibias.n27 0.862419
R22534 diffpairibias diffpairibias.n28 0.684875
R22535 diffpairibias.n12 diffpairibias.n11 0.672012
R22536 diffpairibias.n11 diffpairibias.n10 0.672012
R22537 diffpairibias.n10 diffpairibias.n9 0.672012
R22538 diffpairibias.n9 diffpairibias.n8 0.672012
R22539 diffpairibias.n8 diffpairibias.n7 0.672012
R22540 diffpairibias.n7 diffpairibias.n6 0.672012
R22541 diffpairibias.n6 diffpairibias.n5 0.672012
R22542 diffpairibias.n5 diffpairibias.n4 0.672012
R22543 diffpairibias.n28 diffpairibias.n3 0.190907
R22544 a_n3827_n3924.n51 a_n3827_n3924.t13 214.994
R22545 a_n3827_n3924.t20 a_n3827_n3924.n58 214.994
R22546 a_n3827_n3924.n51 a_n3827_n3924.t17 214.321
R22547 a_n3827_n3924.n53 a_n3827_n3924.t12 214.321
R22548 a_n3827_n3924.n54 a_n3827_n3924.t15 214.321
R22549 a_n3827_n3924.n55 a_n3827_n3924.t11 214.321
R22550 a_n3827_n3924.n56 a_n3827_n3924.t16 214.321
R22551 a_n3827_n3924.n57 a_n3827_n3924.t19 214.321
R22552 a_n3827_n3924.n0 a_n3827_n3924.t18 214.321
R22553 a_n3827_n3924.n58 a_n3827_n3924.t14 214.321
R22554 a_n3827_n3924.n14 a_n3827_n3924.t0 55.8337
R22555 a_n3827_n3924.n13 a_n3827_n3924.t39 55.8337
R22556 a_n3827_n3924.n2 a_n3827_n3924.t9 55.8337
R22557 a_n3827_n3924.n25 a_n3827_n3924.t36 55.8335
R22558 a_n3827_n3924.n49 a_n3827_n3924.t24 55.8335
R22559 a_n3827_n3924.n38 a_n3827_n3924.t51 55.8335
R22560 a_n3827_n3924.n37 a_n3827_n3924.t28 55.8335
R22561 a_n3827_n3924.n26 a_n3827_n3924.t2 55.8335
R22562 a_n3827_n3924.n24 a_n3827_n3924.n23 53.0052
R22563 a_n3827_n3924.n22 a_n3827_n3924.n21 53.0052
R22564 a_n3827_n3924.n20 a_n3827_n3924.n19 53.0052
R22565 a_n3827_n3924.n18 a_n3827_n3924.n17 53.0052
R22566 a_n3827_n3924.n16 a_n3827_n3924.n15 53.0052
R22567 a_n3827_n3924.n12 a_n3827_n3924.n11 53.0052
R22568 a_n3827_n3924.n10 a_n3827_n3924.n9 53.0052
R22569 a_n3827_n3924.n8 a_n3827_n3924.n7 53.0052
R22570 a_n3827_n3924.n6 a_n3827_n3924.n5 53.0052
R22571 a_n3827_n3924.n4 a_n3827_n3924.n3 53.0052
R22572 a_n3827_n3924.n48 a_n3827_n3924.n47 53.0051
R22573 a_n3827_n3924.n46 a_n3827_n3924.n45 53.0051
R22574 a_n3827_n3924.n44 a_n3827_n3924.n43 53.0051
R22575 a_n3827_n3924.n42 a_n3827_n3924.n41 53.0051
R22576 a_n3827_n3924.n40 a_n3827_n3924.n39 53.0051
R22577 a_n3827_n3924.n36 a_n3827_n3924.n35 53.0051
R22578 a_n3827_n3924.n34 a_n3827_n3924.n33 53.0051
R22579 a_n3827_n3924.n32 a_n3827_n3924.n31 53.0051
R22580 a_n3827_n3924.n30 a_n3827_n3924.n29 53.0051
R22581 a_n3827_n3924.n28 a_n3827_n3924.n27 53.0051
R22582 a_n3827_n3924.n2 a_n3827_n3924.n1 12.1555
R22583 a_n3827_n3924.n50 a_n3827_n3924.n25 12.1555
R22584 a_n3827_n3924.n26 a_n3827_n3924.n1 5.07593
R22585 a_n3827_n3924.n50 a_n3827_n3924.n49 5.07593
R22586 a_n3827_n3924.n47 a_n3827_n3924.t21 2.82907
R22587 a_n3827_n3924.n47 a_n3827_n3924.t4 2.82907
R22588 a_n3827_n3924.n45 a_n3827_n3924.t50 2.82907
R22589 a_n3827_n3924.n45 a_n3827_n3924.t45 2.82907
R22590 a_n3827_n3924.n43 a_n3827_n3924.t43 2.82907
R22591 a_n3827_n3924.n43 a_n3827_n3924.t41 2.82907
R22592 a_n3827_n3924.n41 a_n3827_n3924.t47 2.82907
R22593 a_n3827_n3924.n41 a_n3827_n3924.t32 2.82907
R22594 a_n3827_n3924.n39 a_n3827_n3924.t49 2.82907
R22595 a_n3827_n3924.n39 a_n3827_n3924.t5 2.82907
R22596 a_n3827_n3924.n35 a_n3827_n3924.t54 2.82907
R22597 a_n3827_n3924.n35 a_n3827_n3924.t3 2.82907
R22598 a_n3827_n3924.n33 a_n3827_n3924.t33 2.82907
R22599 a_n3827_n3924.n33 a_n3827_n3924.t30 2.82907
R22600 a_n3827_n3924.n31 a_n3827_n3924.t29 2.82907
R22601 a_n3827_n3924.n31 a_n3827_n3924.t1 2.82907
R22602 a_n3827_n3924.n29 a_n3827_n3924.t10 2.82907
R22603 a_n3827_n3924.n29 a_n3827_n3924.t57 2.82907
R22604 a_n3827_n3924.n27 a_n3827_n3924.t44 2.82907
R22605 a_n3827_n3924.n27 a_n3827_n3924.t52 2.82907
R22606 a_n3827_n3924.n23 a_n3827_n3924.t23 2.82907
R22607 a_n3827_n3924.n23 a_n3827_n3924.t55 2.82907
R22608 a_n3827_n3924.n21 a_n3827_n3924.t37 2.82907
R22609 a_n3827_n3924.n21 a_n3827_n3924.t53 2.82907
R22610 a_n3827_n3924.n19 a_n3827_n3924.t35 2.82907
R22611 a_n3827_n3924.n19 a_n3827_n3924.t56 2.82907
R22612 a_n3827_n3924.n17 a_n3827_n3924.t26 2.82907
R22613 a_n3827_n3924.n17 a_n3827_n3924.t27 2.82907
R22614 a_n3827_n3924.n15 a_n3827_n3924.t38 2.82907
R22615 a_n3827_n3924.n15 a_n3827_n3924.t34 2.82907
R22616 a_n3827_n3924.n11 a_n3827_n3924.t40 2.82907
R22617 a_n3827_n3924.n11 a_n3827_n3924.t8 2.82907
R22618 a_n3827_n3924.n9 a_n3827_n3924.t46 2.82907
R22619 a_n3827_n3924.n9 a_n3827_n3924.t7 2.82907
R22620 a_n3827_n3924.n7 a_n3827_n3924.t48 2.82907
R22621 a_n3827_n3924.n7 a_n3827_n3924.t42 2.82907
R22622 a_n3827_n3924.n5 a_n3827_n3924.t6 2.82907
R22623 a_n3827_n3924.n5 a_n3827_n3924.t22 2.82907
R22624 a_n3827_n3924.n3 a_n3827_n3924.t31 2.82907
R22625 a_n3827_n3924.n3 a_n3827_n3924.t25 2.82907
R22626 a_n3827_n3924.n0 a_n3827_n3924.n1 1.95694
R22627 a_n3827_n3924.n52 a_n3827_n3924.n50 1.95694
R22628 a_n3827_n3924.n58 a_n3827_n3924.n0 0.672012
R22629 a_n3827_n3924.n57 a_n3827_n3924.n56 0.672012
R22630 a_n3827_n3924.n56 a_n3827_n3924.n55 0.672012
R22631 a_n3827_n3924.n55 a_n3827_n3924.n54 0.672012
R22632 a_n3827_n3924.n54 a_n3827_n3924.n53 0.672012
R22633 a_n3827_n3924.n0 a_n3827_n3924.n57 0.672012
R22634 a_n3827_n3924.n53 a_n3827_n3924.n52 0.501227
R22635 a_n3827_n3924.n4 a_n3827_n3924.n2 0.358259
R22636 a_n3827_n3924.n6 a_n3827_n3924.n4 0.358259
R22637 a_n3827_n3924.n8 a_n3827_n3924.n6 0.358259
R22638 a_n3827_n3924.n10 a_n3827_n3924.n8 0.358259
R22639 a_n3827_n3924.n12 a_n3827_n3924.n10 0.358259
R22640 a_n3827_n3924.n13 a_n3827_n3924.n12 0.358259
R22641 a_n3827_n3924.n16 a_n3827_n3924.n14 0.358259
R22642 a_n3827_n3924.n18 a_n3827_n3924.n16 0.358259
R22643 a_n3827_n3924.n20 a_n3827_n3924.n18 0.358259
R22644 a_n3827_n3924.n22 a_n3827_n3924.n20 0.358259
R22645 a_n3827_n3924.n24 a_n3827_n3924.n22 0.358259
R22646 a_n3827_n3924.n25 a_n3827_n3924.n24 0.358259
R22647 a_n3827_n3924.n28 a_n3827_n3924.n26 0.358259
R22648 a_n3827_n3924.n30 a_n3827_n3924.n28 0.358259
R22649 a_n3827_n3924.n32 a_n3827_n3924.n30 0.358259
R22650 a_n3827_n3924.n34 a_n3827_n3924.n32 0.358259
R22651 a_n3827_n3924.n36 a_n3827_n3924.n34 0.358259
R22652 a_n3827_n3924.n37 a_n3827_n3924.n36 0.358259
R22653 a_n3827_n3924.n40 a_n3827_n3924.n38 0.358259
R22654 a_n3827_n3924.n42 a_n3827_n3924.n40 0.358259
R22655 a_n3827_n3924.n44 a_n3827_n3924.n42 0.358259
R22656 a_n3827_n3924.n46 a_n3827_n3924.n44 0.358259
R22657 a_n3827_n3924.n48 a_n3827_n3924.n46 0.358259
R22658 a_n3827_n3924.n49 a_n3827_n3924.n48 0.358259
R22659 a_n3827_n3924.n14 a_n3827_n3924.n13 0.235414
R22660 a_n3827_n3924.n38 a_n3827_n3924.n37 0.235414
R22661 a_n3827_n3924.n52 a_n3827_n3924.n51 0.171285
R22662 output.n41 output.n15 289.615
R22663 output.n72 output.n46 289.615
R22664 output.n104 output.n78 289.615
R22665 output.n136 output.n110 289.615
R22666 output.n77 output.n45 197.26
R22667 output.n77 output.n76 196.298
R22668 output.n109 output.n108 196.298
R22669 output.n141 output.n140 196.298
R22670 output.n42 output.n41 185
R22671 output.n40 output.n39 185
R22672 output.n19 output.n18 185
R22673 output.n34 output.n33 185
R22674 output.n32 output.n31 185
R22675 output.n23 output.n22 185
R22676 output.n26 output.n25 185
R22677 output.n73 output.n72 185
R22678 output.n71 output.n70 185
R22679 output.n50 output.n49 185
R22680 output.n65 output.n64 185
R22681 output.n63 output.n62 185
R22682 output.n54 output.n53 185
R22683 output.n57 output.n56 185
R22684 output.n105 output.n104 185
R22685 output.n103 output.n102 185
R22686 output.n82 output.n81 185
R22687 output.n97 output.n96 185
R22688 output.n95 output.n94 185
R22689 output.n86 output.n85 185
R22690 output.n89 output.n88 185
R22691 output.n137 output.n136 185
R22692 output.n135 output.n134 185
R22693 output.n114 output.n113 185
R22694 output.n129 output.n128 185
R22695 output.n127 output.n126 185
R22696 output.n118 output.n117 185
R22697 output.n121 output.n120 185
R22698 output.t2 output.n24 147.661
R22699 output.t19 output.n55 147.661
R22700 output.t0 output.n87 147.661
R22701 output.t1 output.n119 147.661
R22702 output.n41 output.n40 104.615
R22703 output.n40 output.n18 104.615
R22704 output.n33 output.n18 104.615
R22705 output.n33 output.n32 104.615
R22706 output.n32 output.n22 104.615
R22707 output.n25 output.n22 104.615
R22708 output.n72 output.n71 104.615
R22709 output.n71 output.n49 104.615
R22710 output.n64 output.n49 104.615
R22711 output.n64 output.n63 104.615
R22712 output.n63 output.n53 104.615
R22713 output.n56 output.n53 104.615
R22714 output.n104 output.n103 104.615
R22715 output.n103 output.n81 104.615
R22716 output.n96 output.n81 104.615
R22717 output.n96 output.n95 104.615
R22718 output.n95 output.n85 104.615
R22719 output.n88 output.n85 104.615
R22720 output.n136 output.n135 104.615
R22721 output.n135 output.n113 104.615
R22722 output.n128 output.n113 104.615
R22723 output.n128 output.n127 104.615
R22724 output.n127 output.n117 104.615
R22725 output.n120 output.n117 104.615
R22726 output.n1 output.t15 77.056
R22727 output.n14 output.t16 76.6694
R22728 output.n1 output.n0 72.7095
R22729 output.n3 output.n2 72.7095
R22730 output.n5 output.n4 72.7095
R22731 output.n7 output.n6 72.7095
R22732 output.n9 output.n8 72.7095
R22733 output.n11 output.n10 72.7095
R22734 output.n13 output.n12 72.7095
R22735 output.n25 output.t2 52.3082
R22736 output.n56 output.t19 52.3082
R22737 output.n88 output.t0 52.3082
R22738 output.n120 output.t1 52.3082
R22739 output.n26 output.n24 15.6674
R22740 output.n57 output.n55 15.6674
R22741 output.n89 output.n87 15.6674
R22742 output.n121 output.n119 15.6674
R22743 output.n27 output.n23 12.8005
R22744 output.n58 output.n54 12.8005
R22745 output.n90 output.n86 12.8005
R22746 output.n122 output.n118 12.8005
R22747 output.n31 output.n30 12.0247
R22748 output.n62 output.n61 12.0247
R22749 output.n94 output.n93 12.0247
R22750 output.n126 output.n125 12.0247
R22751 output.n34 output.n21 11.249
R22752 output.n65 output.n52 11.249
R22753 output.n97 output.n84 11.249
R22754 output.n129 output.n116 11.249
R22755 output.n35 output.n19 10.4732
R22756 output.n66 output.n50 10.4732
R22757 output.n98 output.n82 10.4732
R22758 output.n130 output.n114 10.4732
R22759 output.n39 output.n38 9.69747
R22760 output.n70 output.n69 9.69747
R22761 output.n102 output.n101 9.69747
R22762 output.n134 output.n133 9.69747
R22763 output.n45 output.n44 9.45567
R22764 output.n76 output.n75 9.45567
R22765 output.n108 output.n107 9.45567
R22766 output.n140 output.n139 9.45567
R22767 output.n44 output.n43 9.3005
R22768 output.n17 output.n16 9.3005
R22769 output.n38 output.n37 9.3005
R22770 output.n36 output.n35 9.3005
R22771 output.n21 output.n20 9.3005
R22772 output.n30 output.n29 9.3005
R22773 output.n28 output.n27 9.3005
R22774 output.n75 output.n74 9.3005
R22775 output.n48 output.n47 9.3005
R22776 output.n69 output.n68 9.3005
R22777 output.n67 output.n66 9.3005
R22778 output.n52 output.n51 9.3005
R22779 output.n61 output.n60 9.3005
R22780 output.n59 output.n58 9.3005
R22781 output.n107 output.n106 9.3005
R22782 output.n80 output.n79 9.3005
R22783 output.n101 output.n100 9.3005
R22784 output.n99 output.n98 9.3005
R22785 output.n84 output.n83 9.3005
R22786 output.n93 output.n92 9.3005
R22787 output.n91 output.n90 9.3005
R22788 output.n139 output.n138 9.3005
R22789 output.n112 output.n111 9.3005
R22790 output.n133 output.n132 9.3005
R22791 output.n131 output.n130 9.3005
R22792 output.n116 output.n115 9.3005
R22793 output.n125 output.n124 9.3005
R22794 output.n123 output.n122 9.3005
R22795 output.n42 output.n17 8.92171
R22796 output.n73 output.n48 8.92171
R22797 output.n105 output.n80 8.92171
R22798 output.n137 output.n112 8.92171
R22799 output output.n141 8.15037
R22800 output.n43 output.n15 8.14595
R22801 output.n74 output.n46 8.14595
R22802 output.n106 output.n78 8.14595
R22803 output.n138 output.n110 8.14595
R22804 output.n45 output.n15 5.81868
R22805 output.n76 output.n46 5.81868
R22806 output.n108 output.n78 5.81868
R22807 output.n140 output.n110 5.81868
R22808 output.n43 output.n42 5.04292
R22809 output.n74 output.n73 5.04292
R22810 output.n106 output.n105 5.04292
R22811 output.n138 output.n137 5.04292
R22812 output.n28 output.n24 4.38594
R22813 output.n59 output.n55 4.38594
R22814 output.n91 output.n87 4.38594
R22815 output.n123 output.n119 4.38594
R22816 output.n39 output.n17 4.26717
R22817 output.n70 output.n48 4.26717
R22818 output.n102 output.n80 4.26717
R22819 output.n134 output.n112 4.26717
R22820 output.n0 output.t5 3.9605
R22821 output.n0 output.t9 3.9605
R22822 output.n2 output.t12 3.9605
R22823 output.n2 output.t17 3.9605
R22824 output.n4 output.t18 3.9605
R22825 output.n4 output.t7 3.9605
R22826 output.n6 output.t11 3.9605
R22827 output.n6 output.t3 3.9605
R22828 output.n8 output.t6 3.9605
R22829 output.n8 output.t4 3.9605
R22830 output.n10 output.t10 3.9605
R22831 output.n10 output.t13 3.9605
R22832 output.n12 output.t14 3.9605
R22833 output.n12 output.t8 3.9605
R22834 output.n38 output.n19 3.49141
R22835 output.n69 output.n50 3.49141
R22836 output.n101 output.n82 3.49141
R22837 output.n133 output.n114 3.49141
R22838 output.n35 output.n34 2.71565
R22839 output.n66 output.n65 2.71565
R22840 output.n98 output.n97 2.71565
R22841 output.n130 output.n129 2.71565
R22842 output.n31 output.n21 1.93989
R22843 output.n62 output.n52 1.93989
R22844 output.n94 output.n84 1.93989
R22845 output.n126 output.n116 1.93989
R22846 output.n30 output.n23 1.16414
R22847 output.n61 output.n54 1.16414
R22848 output.n93 output.n86 1.16414
R22849 output.n125 output.n118 1.16414
R22850 output.n141 output.n109 0.962709
R22851 output.n109 output.n77 0.962709
R22852 output.n27 output.n26 0.388379
R22853 output.n58 output.n57 0.388379
R22854 output.n90 output.n89 0.388379
R22855 output.n122 output.n121 0.388379
R22856 output.n14 output.n13 0.387128
R22857 output.n13 output.n11 0.387128
R22858 output.n11 output.n9 0.387128
R22859 output.n9 output.n7 0.387128
R22860 output.n7 output.n5 0.387128
R22861 output.n5 output.n3 0.387128
R22862 output.n3 output.n1 0.387128
R22863 output.n44 output.n16 0.155672
R22864 output.n37 output.n16 0.155672
R22865 output.n37 output.n36 0.155672
R22866 output.n36 output.n20 0.155672
R22867 output.n29 output.n20 0.155672
R22868 output.n29 output.n28 0.155672
R22869 output.n75 output.n47 0.155672
R22870 output.n68 output.n47 0.155672
R22871 output.n68 output.n67 0.155672
R22872 output.n67 output.n51 0.155672
R22873 output.n60 output.n51 0.155672
R22874 output.n60 output.n59 0.155672
R22875 output.n107 output.n79 0.155672
R22876 output.n100 output.n79 0.155672
R22877 output.n100 output.n99 0.155672
R22878 output.n99 output.n83 0.155672
R22879 output.n92 output.n83 0.155672
R22880 output.n92 output.n91 0.155672
R22881 output.n139 output.n111 0.155672
R22882 output.n132 output.n111 0.155672
R22883 output.n132 output.n131 0.155672
R22884 output.n131 output.n115 0.155672
R22885 output.n124 output.n115 0.155672
R22886 output.n124 output.n123 0.155672
R22887 output output.n14 0.126227
R22888 a_n2650_8322.n10 a_n2650_8322.t3 74.6477
R22889 a_n2650_8322.n1 a_n2650_8322.t23 74.6477
R22890 a_n2650_8322.n24 a_n2650_8322.t25 74.6474
R22891 a_n2650_8322.n18 a_n2650_8322.t22 74.2899
R22892 a_n2650_8322.n11 a_n2650_8322.t1 74.2899
R22893 a_n2650_8322.n12 a_n2650_8322.t4 74.2899
R22894 a_n2650_8322.n15 a_n2650_8322.t5 74.2899
R22895 a_n2650_8322.n8 a_n2650_8322.t8 74.2899
R22896 a_n2650_8322.n24 a_n2650_8322.n23 70.6783
R22897 a_n2650_8322.n22 a_n2650_8322.n21 70.6783
R22898 a_n2650_8322.n20 a_n2650_8322.n19 70.6783
R22899 a_n2650_8322.n10 a_n2650_8322.n9 70.6783
R22900 a_n2650_8322.n14 a_n2650_8322.n13 70.6783
R22901 a_n2650_8322.n1 a_n2650_8322.n0 70.6783
R22902 a_n2650_8322.n3 a_n2650_8322.n2 70.6783
R22903 a_n2650_8322.n5 a_n2650_8322.n4 70.6783
R22904 a_n2650_8322.n7 a_n2650_8322.n6 70.6783
R22905 a_n2650_8322.n26 a_n2650_8322.n25 70.6782
R22906 a_n2650_8322.n16 a_n2650_8322.n8 24.1867
R22907 a_n2650_8322.n17 a_n2650_8322.t28 9.90091
R22908 a_n2650_8322.n16 a_n2650_8322.n15 7.67184
R22909 a_n2650_8322.n18 a_n2650_8322.n17 6.55222
R22910 a_n2650_8322.n17 a_n2650_8322.n16 5.3452
R22911 a_n2650_8322.n23 a_n2650_8322.t20 3.61217
R22912 a_n2650_8322.n23 a_n2650_8322.t16 3.61217
R22913 a_n2650_8322.n21 a_n2650_8322.t24 3.61217
R22914 a_n2650_8322.n21 a_n2650_8322.t14 3.61217
R22915 a_n2650_8322.n19 a_n2650_8322.t12 3.61217
R22916 a_n2650_8322.n19 a_n2650_8322.t11 3.61217
R22917 a_n2650_8322.n9 a_n2650_8322.t7 3.61217
R22918 a_n2650_8322.n9 a_n2650_8322.t6 3.61217
R22919 a_n2650_8322.n13 a_n2650_8322.t2 3.61217
R22920 a_n2650_8322.n13 a_n2650_8322.t0 3.61217
R22921 a_n2650_8322.n0 a_n2650_8322.t26 3.61217
R22922 a_n2650_8322.n0 a_n2650_8322.t18 3.61217
R22923 a_n2650_8322.n2 a_n2650_8322.t10 3.61217
R22924 a_n2650_8322.n2 a_n2650_8322.t9 3.61217
R22925 a_n2650_8322.n4 a_n2650_8322.t21 3.61217
R22926 a_n2650_8322.n4 a_n2650_8322.t15 3.61217
R22927 a_n2650_8322.n6 a_n2650_8322.t19 3.61217
R22928 a_n2650_8322.n6 a_n2650_8322.t17 3.61217
R22929 a_n2650_8322.n26 a_n2650_8322.t13 3.61217
R22930 a_n2650_8322.t27 a_n2650_8322.n26 3.61217
R22931 a_n2650_8322.n15 a_n2650_8322.n14 0.358259
R22932 a_n2650_8322.n14 a_n2650_8322.n12 0.358259
R22933 a_n2650_8322.n11 a_n2650_8322.n10 0.358259
R22934 a_n2650_8322.n8 a_n2650_8322.n7 0.358259
R22935 a_n2650_8322.n7 a_n2650_8322.n5 0.358259
R22936 a_n2650_8322.n5 a_n2650_8322.n3 0.358259
R22937 a_n2650_8322.n3 a_n2650_8322.n1 0.358259
R22938 a_n2650_8322.n20 a_n2650_8322.n18 0.358259
R22939 a_n2650_8322.n22 a_n2650_8322.n20 0.358259
R22940 a_n2650_8322.n25 a_n2650_8322.n22 0.358259
R22941 a_n2650_8322.n25 a_n2650_8322.n24 0.358259
R22942 a_n2650_8322.n12 a_n2650_8322.n11 0.101793
R22943 a_n2650_8322.t30 a_n2650_8322.t33 0.0788333
R22944 a_n2650_8322.t29 a_n2650_8322.t31 0.0788333
R22945 a_n2650_8322.t28 a_n2650_8322.t32 0.0788333
R22946 a_n2650_8322.t29 a_n2650_8322.t30 0.0318333
R22947 a_n2650_8322.t28 a_n2650_8322.t31 0.0318333
R22948 a_n2650_8322.t33 a_n2650_8322.t31 0.0318333
R22949 a_n2650_8322.t32 a_n2650_8322.t29 0.0318333
R22950 plus.n43 plus.t25 442.325
R22951 plus.n11 plus.t12 442.325
R22952 plus.n42 plus.t5 415.966
R22953 plus.n41 plus.t20 415.966
R22954 plus.n47 plus.t26 415.966
R22955 plus.n39 plus.t11 415.966
R22956 plus.n52 plus.t6 415.966
R22957 plus.n54 plus.t10 415.966
R22958 plus.n37 plus.t19 415.966
R22959 plus.n59 plus.t8 415.966
R22960 plus.n35 plus.t16 415.966
R22961 plus.n64 plus.t28 415.966
R22962 plus.n66 plus.t21 415.966
R22963 plus.n32 plus.t23 415.966
R22964 plus.n30 plus.t13 415.966
R22965 plus.n29 plus.t27 415.966
R22966 plus.n3 plus.t22 415.966
R22967 plus.n23 plus.t7 415.966
R22968 plus.n22 plus.t18 415.966
R22969 plus.n6 plus.t14 415.966
R22970 plus.n17 plus.t24 415.966
R22971 plus.n15 plus.t17 415.966
R22972 plus.n9 plus.t9 415.966
R22973 plus.n10 plus.t15 415.966
R22974 plus.n70 plus.t3 243.97
R22975 plus.n70 plus.n69 223.454
R22976 plus.n72 plus.n71 223.454
R22977 plus.n67 plus.n66 161.3
R22978 plus.n65 plus.n34 161.3
R22979 plus.n64 plus.n63 161.3
R22980 plus.n62 plus.n35 161.3
R22981 plus.n61 plus.n60 161.3
R22982 plus.n59 plus.n36 161.3
R22983 plus.n58 plus.n57 161.3
R22984 plus.n56 plus.n37 161.3
R22985 plus.n55 plus.n54 161.3
R22986 plus.n53 plus.n38 161.3
R22987 plus.n52 plus.n51 161.3
R22988 plus.n50 plus.n39 161.3
R22989 plus.n49 plus.n48 161.3
R22990 plus.n47 plus.n40 161.3
R22991 plus.n46 plus.n45 161.3
R22992 plus.n44 plus.n41 161.3
R22993 plus.n12 plus.n9 161.3
R22994 plus.n14 plus.n13 161.3
R22995 plus.n15 plus.n8 161.3
R22996 plus.n16 plus.n7 161.3
R22997 plus.n18 plus.n17 161.3
R22998 plus.n19 plus.n6 161.3
R22999 plus.n21 plus.n20 161.3
R23000 plus.n22 plus.n5 161.3
R23001 plus.n23 plus.n4 161.3
R23002 plus.n25 plus.n24 161.3
R23003 plus.n26 plus.n3 161.3
R23004 plus.n28 plus.n27 161.3
R23005 plus.n29 plus.n2 161.3
R23006 plus.n30 plus.n1 161.3
R23007 plus.n31 plus.n0 161.3
R23008 plus.n33 plus.n32 161.3
R23009 plus.n42 plus.n41 48.2005
R23010 plus.n52 plus.n39 48.2005
R23011 plus.n54 plus.n37 48.2005
R23012 plus.n64 plus.n35 48.2005
R23013 plus.n30 plus.n29 48.2005
R23014 plus.n23 plus.n22 48.2005
R23015 plus.n17 plus.n6 48.2005
R23016 plus.n10 plus.n9 48.2005
R23017 plus.n48 plus.n47 47.4702
R23018 plus.n59 plus.n58 47.4702
R23019 plus.n24 plus.n3 47.4702
R23020 plus.n16 plus.n15 47.4702
R23021 plus.n66 plus.n65 46.0096
R23022 plus.n32 plus.n31 46.0096
R23023 plus.n44 plus.n43 45.0871
R23024 plus.n12 plus.n11 45.0871
R23025 plus.n68 plus.n67 31.0554
R23026 plus.n47 plus.n46 25.5611
R23027 plus.n60 plus.n59 25.5611
R23028 plus.n28 plus.n3 25.5611
R23029 plus.n15 plus.n14 25.5611
R23030 plus.n53 plus.n52 24.1005
R23031 plus.n54 plus.n53 24.1005
R23032 plus.n22 plus.n21 24.1005
R23033 plus.n21 plus.n6 24.1005
R23034 plus.n46 plus.n41 22.6399
R23035 plus.n60 plus.n35 22.6399
R23036 plus.n29 plus.n28 22.6399
R23037 plus.n14 plus.n9 22.6399
R23038 plus.n69 plus.t4 19.8005
R23039 plus.n69 plus.t1 19.8005
R23040 plus.n71 plus.t0 19.8005
R23041 plus.n71 plus.t2 19.8005
R23042 plus plus.n73 14.7003
R23043 plus.n43 plus.n42 14.1472
R23044 plus.n11 plus.n10 14.1472
R23045 plus.n68 plus.n33 11.7259
R23046 plus.n73 plus.n72 5.40567
R23047 plus.n65 plus.n64 2.19141
R23048 plus.n31 plus.n30 2.19141
R23049 plus.n73 plus.n68 1.188
R23050 plus.n48 plus.n39 0.730803
R23051 plus.n58 plus.n37 0.730803
R23052 plus.n24 plus.n23 0.730803
R23053 plus.n17 plus.n16 0.730803
R23054 plus.n72 plus.n70 0.716017
R23055 plus.n45 plus.n44 0.189894
R23056 plus.n45 plus.n40 0.189894
R23057 plus.n49 plus.n40 0.189894
R23058 plus.n50 plus.n49 0.189894
R23059 plus.n51 plus.n50 0.189894
R23060 plus.n51 plus.n38 0.189894
R23061 plus.n55 plus.n38 0.189894
R23062 plus.n56 plus.n55 0.189894
R23063 plus.n57 plus.n56 0.189894
R23064 plus.n57 plus.n36 0.189894
R23065 plus.n61 plus.n36 0.189894
R23066 plus.n62 plus.n61 0.189894
R23067 plus.n63 plus.n62 0.189894
R23068 plus.n63 plus.n34 0.189894
R23069 plus.n67 plus.n34 0.189894
R23070 plus.n33 plus.n0 0.189894
R23071 plus.n1 plus.n0 0.189894
R23072 plus.n2 plus.n1 0.189894
R23073 plus.n27 plus.n2 0.189894
R23074 plus.n27 plus.n26 0.189894
R23075 plus.n26 plus.n25 0.189894
R23076 plus.n25 plus.n4 0.189894
R23077 plus.n5 plus.n4 0.189894
R23078 plus.n20 plus.n5 0.189894
R23079 plus.n20 plus.n19 0.189894
R23080 plus.n19 plus.n18 0.189894
R23081 plus.n18 plus.n7 0.189894
R23082 plus.n8 plus.n7 0.189894
R23083 plus.n13 plus.n8 0.189894
R23084 plus.n13 plus.n12 0.189894
R23085 minus.n45 minus.t26 442.325
R23086 minus.n9 minus.t12 442.325
R23087 minus.n66 minus.t16 415.966
R23088 minus.n64 minus.t28 415.966
R23089 minus.n63 minus.t21 415.966
R23090 minus.n37 minus.t14 415.966
R23091 minus.n57 minus.t23 415.966
R23092 minus.n56 minus.t11 415.966
R23093 minus.n40 minus.t5 415.966
R23094 minus.n51 minus.t17 415.966
R23095 minus.n49 minus.t10 415.966
R23096 minus.n43 minus.t25 415.966
R23097 minus.n44 minus.t7 415.966
R23098 minus.n8 minus.t18 415.966
R23099 minus.n7 minus.t8 415.966
R23100 minus.n13 minus.t13 415.966
R23101 minus.n5 minus.t24 415.966
R23102 minus.n18 minus.t19 415.966
R23103 minus.n20 minus.t22 415.966
R23104 minus.n3 minus.t6 415.966
R23105 minus.n25 minus.t20 415.966
R23106 minus.n1 minus.t27 415.966
R23107 minus.n30 minus.t15 415.966
R23108 minus.n32 minus.t9 415.966
R23109 minus.n72 minus.t3 243.255
R23110 minus.n71 minus.n69 224.169
R23111 minus.n71 minus.n70 223.454
R23112 minus.n46 minus.n43 161.3
R23113 minus.n48 minus.n47 161.3
R23114 minus.n49 minus.n42 161.3
R23115 minus.n50 minus.n41 161.3
R23116 minus.n52 minus.n51 161.3
R23117 minus.n53 minus.n40 161.3
R23118 minus.n55 minus.n54 161.3
R23119 minus.n56 minus.n39 161.3
R23120 minus.n57 minus.n38 161.3
R23121 minus.n59 minus.n58 161.3
R23122 minus.n60 minus.n37 161.3
R23123 minus.n62 minus.n61 161.3
R23124 minus.n63 minus.n36 161.3
R23125 minus.n64 minus.n35 161.3
R23126 minus.n65 minus.n34 161.3
R23127 minus.n67 minus.n66 161.3
R23128 minus.n33 minus.n32 161.3
R23129 minus.n31 minus.n0 161.3
R23130 minus.n30 minus.n29 161.3
R23131 minus.n28 minus.n1 161.3
R23132 minus.n27 minus.n26 161.3
R23133 minus.n25 minus.n2 161.3
R23134 minus.n24 minus.n23 161.3
R23135 minus.n22 minus.n3 161.3
R23136 minus.n21 minus.n20 161.3
R23137 minus.n19 minus.n4 161.3
R23138 minus.n18 minus.n17 161.3
R23139 minus.n16 minus.n5 161.3
R23140 minus.n15 minus.n14 161.3
R23141 minus.n13 minus.n6 161.3
R23142 minus.n12 minus.n11 161.3
R23143 minus.n10 minus.n7 161.3
R23144 minus.n64 minus.n63 48.2005
R23145 minus.n57 minus.n56 48.2005
R23146 minus.n51 minus.n40 48.2005
R23147 minus.n44 minus.n43 48.2005
R23148 minus.n8 minus.n7 48.2005
R23149 minus.n18 minus.n5 48.2005
R23150 minus.n20 minus.n3 48.2005
R23151 minus.n30 minus.n1 48.2005
R23152 minus.n58 minus.n37 47.4702
R23153 minus.n50 minus.n49 47.4702
R23154 minus.n14 minus.n13 47.4702
R23155 minus.n25 minus.n24 47.4702
R23156 minus.n66 minus.n65 46.0096
R23157 minus.n32 minus.n31 46.0096
R23158 minus.n10 minus.n9 45.0871
R23159 minus.n46 minus.n45 45.0871
R23160 minus.n68 minus.n67 31.2713
R23161 minus.n62 minus.n37 25.5611
R23162 minus.n49 minus.n48 25.5611
R23163 minus.n13 minus.n12 25.5611
R23164 minus.n26 minus.n25 25.5611
R23165 minus.n56 minus.n55 24.1005
R23166 minus.n55 minus.n40 24.1005
R23167 minus.n19 minus.n18 24.1005
R23168 minus.n20 minus.n19 24.1005
R23169 minus.n63 minus.n62 22.6399
R23170 minus.n48 minus.n43 22.6399
R23171 minus.n12 minus.n7 22.6399
R23172 minus.n26 minus.n1 22.6399
R23173 minus.n70 minus.t2 19.8005
R23174 minus.n70 minus.t0 19.8005
R23175 minus.n69 minus.t1 19.8005
R23176 minus.n69 minus.t4 19.8005
R23177 minus.n45 minus.n44 14.1472
R23178 minus.n9 minus.n8 14.1472
R23179 minus.n68 minus.n33 11.9418
R23180 minus minus.n73 11.8631
R23181 minus.n73 minus.n72 4.80222
R23182 minus.n65 minus.n64 2.19141
R23183 minus.n31 minus.n30 2.19141
R23184 minus.n73 minus.n68 0.972091
R23185 minus.n58 minus.n57 0.730803
R23186 minus.n51 minus.n50 0.730803
R23187 minus.n14 minus.n5 0.730803
R23188 minus.n24 minus.n3 0.730803
R23189 minus.n72 minus.n71 0.716017
R23190 minus.n67 minus.n34 0.189894
R23191 minus.n35 minus.n34 0.189894
R23192 minus.n36 minus.n35 0.189894
R23193 minus.n61 minus.n36 0.189894
R23194 minus.n61 minus.n60 0.189894
R23195 minus.n60 minus.n59 0.189894
R23196 minus.n59 minus.n38 0.189894
R23197 minus.n39 minus.n38 0.189894
R23198 minus.n54 minus.n39 0.189894
R23199 minus.n54 minus.n53 0.189894
R23200 minus.n53 minus.n52 0.189894
R23201 minus.n52 minus.n41 0.189894
R23202 minus.n42 minus.n41 0.189894
R23203 minus.n47 minus.n42 0.189894
R23204 minus.n47 minus.n46 0.189894
R23205 minus.n11 minus.n10 0.189894
R23206 minus.n11 minus.n6 0.189894
R23207 minus.n15 minus.n6 0.189894
R23208 minus.n16 minus.n15 0.189894
R23209 minus.n17 minus.n16 0.189894
R23210 minus.n17 minus.n4 0.189894
R23211 minus.n21 minus.n4 0.189894
R23212 minus.n22 minus.n21 0.189894
R23213 minus.n23 minus.n22 0.189894
R23214 minus.n23 minus.n2 0.189894
R23215 minus.n27 minus.n2 0.189894
R23216 minus.n28 minus.n27 0.189894
R23217 minus.n29 minus.n28 0.189894
R23218 minus.n29 minus.n0 0.189894
R23219 minus.n33 minus.n0 0.189894
R23220 outputibias.n27 outputibias.n1 289.615
R23221 outputibias.n58 outputibias.n32 289.615
R23222 outputibias.n90 outputibias.n64 289.615
R23223 outputibias.n122 outputibias.n96 289.615
R23224 outputibias.n28 outputibias.n27 185
R23225 outputibias.n26 outputibias.n25 185
R23226 outputibias.n5 outputibias.n4 185
R23227 outputibias.n20 outputibias.n19 185
R23228 outputibias.n18 outputibias.n17 185
R23229 outputibias.n9 outputibias.n8 185
R23230 outputibias.n12 outputibias.n11 185
R23231 outputibias.n59 outputibias.n58 185
R23232 outputibias.n57 outputibias.n56 185
R23233 outputibias.n36 outputibias.n35 185
R23234 outputibias.n51 outputibias.n50 185
R23235 outputibias.n49 outputibias.n48 185
R23236 outputibias.n40 outputibias.n39 185
R23237 outputibias.n43 outputibias.n42 185
R23238 outputibias.n91 outputibias.n90 185
R23239 outputibias.n89 outputibias.n88 185
R23240 outputibias.n68 outputibias.n67 185
R23241 outputibias.n83 outputibias.n82 185
R23242 outputibias.n81 outputibias.n80 185
R23243 outputibias.n72 outputibias.n71 185
R23244 outputibias.n75 outputibias.n74 185
R23245 outputibias.n123 outputibias.n122 185
R23246 outputibias.n121 outputibias.n120 185
R23247 outputibias.n100 outputibias.n99 185
R23248 outputibias.n115 outputibias.n114 185
R23249 outputibias.n113 outputibias.n112 185
R23250 outputibias.n104 outputibias.n103 185
R23251 outputibias.n107 outputibias.n106 185
R23252 outputibias.n0 outputibias.t8 178.945
R23253 outputibias.n133 outputibias.t11 177.018
R23254 outputibias.n132 outputibias.t9 177.018
R23255 outputibias.n0 outputibias.t10 177.018
R23256 outputibias.t5 outputibias.n10 147.661
R23257 outputibias.t7 outputibias.n41 147.661
R23258 outputibias.t1 outputibias.n73 147.661
R23259 outputibias.t3 outputibias.n105 147.661
R23260 outputibias.n128 outputibias.t4 132.363
R23261 outputibias.n128 outputibias.t6 130.436
R23262 outputibias.n129 outputibias.t0 130.436
R23263 outputibias.n130 outputibias.t2 130.436
R23264 outputibias.n27 outputibias.n26 104.615
R23265 outputibias.n26 outputibias.n4 104.615
R23266 outputibias.n19 outputibias.n4 104.615
R23267 outputibias.n19 outputibias.n18 104.615
R23268 outputibias.n18 outputibias.n8 104.615
R23269 outputibias.n11 outputibias.n8 104.615
R23270 outputibias.n58 outputibias.n57 104.615
R23271 outputibias.n57 outputibias.n35 104.615
R23272 outputibias.n50 outputibias.n35 104.615
R23273 outputibias.n50 outputibias.n49 104.615
R23274 outputibias.n49 outputibias.n39 104.615
R23275 outputibias.n42 outputibias.n39 104.615
R23276 outputibias.n90 outputibias.n89 104.615
R23277 outputibias.n89 outputibias.n67 104.615
R23278 outputibias.n82 outputibias.n67 104.615
R23279 outputibias.n82 outputibias.n81 104.615
R23280 outputibias.n81 outputibias.n71 104.615
R23281 outputibias.n74 outputibias.n71 104.615
R23282 outputibias.n122 outputibias.n121 104.615
R23283 outputibias.n121 outputibias.n99 104.615
R23284 outputibias.n114 outputibias.n99 104.615
R23285 outputibias.n114 outputibias.n113 104.615
R23286 outputibias.n113 outputibias.n103 104.615
R23287 outputibias.n106 outputibias.n103 104.615
R23288 outputibias.n63 outputibias.n31 95.6354
R23289 outputibias.n63 outputibias.n62 94.6732
R23290 outputibias.n95 outputibias.n94 94.6732
R23291 outputibias.n127 outputibias.n126 94.6732
R23292 outputibias.n11 outputibias.t5 52.3082
R23293 outputibias.n42 outputibias.t7 52.3082
R23294 outputibias.n74 outputibias.t1 52.3082
R23295 outputibias.n106 outputibias.t3 52.3082
R23296 outputibias.n12 outputibias.n10 15.6674
R23297 outputibias.n43 outputibias.n41 15.6674
R23298 outputibias.n75 outputibias.n73 15.6674
R23299 outputibias.n107 outputibias.n105 15.6674
R23300 outputibias.n13 outputibias.n9 12.8005
R23301 outputibias.n44 outputibias.n40 12.8005
R23302 outputibias.n76 outputibias.n72 12.8005
R23303 outputibias.n108 outputibias.n104 12.8005
R23304 outputibias.n17 outputibias.n16 12.0247
R23305 outputibias.n48 outputibias.n47 12.0247
R23306 outputibias.n80 outputibias.n79 12.0247
R23307 outputibias.n112 outputibias.n111 12.0247
R23308 outputibias.n20 outputibias.n7 11.249
R23309 outputibias.n51 outputibias.n38 11.249
R23310 outputibias.n83 outputibias.n70 11.249
R23311 outputibias.n115 outputibias.n102 11.249
R23312 outputibias.n21 outputibias.n5 10.4732
R23313 outputibias.n52 outputibias.n36 10.4732
R23314 outputibias.n84 outputibias.n68 10.4732
R23315 outputibias.n116 outputibias.n100 10.4732
R23316 outputibias.n25 outputibias.n24 9.69747
R23317 outputibias.n56 outputibias.n55 9.69747
R23318 outputibias.n88 outputibias.n87 9.69747
R23319 outputibias.n120 outputibias.n119 9.69747
R23320 outputibias.n31 outputibias.n30 9.45567
R23321 outputibias.n62 outputibias.n61 9.45567
R23322 outputibias.n94 outputibias.n93 9.45567
R23323 outputibias.n126 outputibias.n125 9.45567
R23324 outputibias.n30 outputibias.n29 9.3005
R23325 outputibias.n3 outputibias.n2 9.3005
R23326 outputibias.n24 outputibias.n23 9.3005
R23327 outputibias.n22 outputibias.n21 9.3005
R23328 outputibias.n7 outputibias.n6 9.3005
R23329 outputibias.n16 outputibias.n15 9.3005
R23330 outputibias.n14 outputibias.n13 9.3005
R23331 outputibias.n61 outputibias.n60 9.3005
R23332 outputibias.n34 outputibias.n33 9.3005
R23333 outputibias.n55 outputibias.n54 9.3005
R23334 outputibias.n53 outputibias.n52 9.3005
R23335 outputibias.n38 outputibias.n37 9.3005
R23336 outputibias.n47 outputibias.n46 9.3005
R23337 outputibias.n45 outputibias.n44 9.3005
R23338 outputibias.n93 outputibias.n92 9.3005
R23339 outputibias.n66 outputibias.n65 9.3005
R23340 outputibias.n87 outputibias.n86 9.3005
R23341 outputibias.n85 outputibias.n84 9.3005
R23342 outputibias.n70 outputibias.n69 9.3005
R23343 outputibias.n79 outputibias.n78 9.3005
R23344 outputibias.n77 outputibias.n76 9.3005
R23345 outputibias.n125 outputibias.n124 9.3005
R23346 outputibias.n98 outputibias.n97 9.3005
R23347 outputibias.n119 outputibias.n118 9.3005
R23348 outputibias.n117 outputibias.n116 9.3005
R23349 outputibias.n102 outputibias.n101 9.3005
R23350 outputibias.n111 outputibias.n110 9.3005
R23351 outputibias.n109 outputibias.n108 9.3005
R23352 outputibias.n28 outputibias.n3 8.92171
R23353 outputibias.n59 outputibias.n34 8.92171
R23354 outputibias.n91 outputibias.n66 8.92171
R23355 outputibias.n123 outputibias.n98 8.92171
R23356 outputibias.n29 outputibias.n1 8.14595
R23357 outputibias.n60 outputibias.n32 8.14595
R23358 outputibias.n92 outputibias.n64 8.14595
R23359 outputibias.n124 outputibias.n96 8.14595
R23360 outputibias.n31 outputibias.n1 5.81868
R23361 outputibias.n62 outputibias.n32 5.81868
R23362 outputibias.n94 outputibias.n64 5.81868
R23363 outputibias.n126 outputibias.n96 5.81868
R23364 outputibias.n131 outputibias.n130 5.20947
R23365 outputibias.n29 outputibias.n28 5.04292
R23366 outputibias.n60 outputibias.n59 5.04292
R23367 outputibias.n92 outputibias.n91 5.04292
R23368 outputibias.n124 outputibias.n123 5.04292
R23369 outputibias.n131 outputibias.n127 4.42209
R23370 outputibias.n14 outputibias.n10 4.38594
R23371 outputibias.n45 outputibias.n41 4.38594
R23372 outputibias.n77 outputibias.n73 4.38594
R23373 outputibias.n109 outputibias.n105 4.38594
R23374 outputibias.n132 outputibias.n131 4.28454
R23375 outputibias.n25 outputibias.n3 4.26717
R23376 outputibias.n56 outputibias.n34 4.26717
R23377 outputibias.n88 outputibias.n66 4.26717
R23378 outputibias.n120 outputibias.n98 4.26717
R23379 outputibias.n24 outputibias.n5 3.49141
R23380 outputibias.n55 outputibias.n36 3.49141
R23381 outputibias.n87 outputibias.n68 3.49141
R23382 outputibias.n119 outputibias.n100 3.49141
R23383 outputibias.n21 outputibias.n20 2.71565
R23384 outputibias.n52 outputibias.n51 2.71565
R23385 outputibias.n84 outputibias.n83 2.71565
R23386 outputibias.n116 outputibias.n115 2.71565
R23387 outputibias.n17 outputibias.n7 1.93989
R23388 outputibias.n48 outputibias.n38 1.93989
R23389 outputibias.n80 outputibias.n70 1.93989
R23390 outputibias.n112 outputibias.n102 1.93989
R23391 outputibias.n130 outputibias.n129 1.9266
R23392 outputibias.n129 outputibias.n128 1.9266
R23393 outputibias.n133 outputibias.n132 1.92658
R23394 outputibias.n134 outputibias.n133 1.29913
R23395 outputibias.n16 outputibias.n9 1.16414
R23396 outputibias.n47 outputibias.n40 1.16414
R23397 outputibias.n79 outputibias.n72 1.16414
R23398 outputibias.n111 outputibias.n104 1.16414
R23399 outputibias.n127 outputibias.n95 0.962709
R23400 outputibias.n95 outputibias.n63 0.962709
R23401 outputibias.n13 outputibias.n12 0.388379
R23402 outputibias.n44 outputibias.n43 0.388379
R23403 outputibias.n76 outputibias.n75 0.388379
R23404 outputibias.n108 outputibias.n107 0.388379
R23405 outputibias.n134 outputibias.n0 0.337251
R23406 outputibias outputibias.n134 0.302375
R23407 outputibias.n30 outputibias.n2 0.155672
R23408 outputibias.n23 outputibias.n2 0.155672
R23409 outputibias.n23 outputibias.n22 0.155672
R23410 outputibias.n22 outputibias.n6 0.155672
R23411 outputibias.n15 outputibias.n6 0.155672
R23412 outputibias.n15 outputibias.n14 0.155672
R23413 outputibias.n61 outputibias.n33 0.155672
R23414 outputibias.n54 outputibias.n33 0.155672
R23415 outputibias.n54 outputibias.n53 0.155672
R23416 outputibias.n53 outputibias.n37 0.155672
R23417 outputibias.n46 outputibias.n37 0.155672
R23418 outputibias.n46 outputibias.n45 0.155672
R23419 outputibias.n93 outputibias.n65 0.155672
R23420 outputibias.n86 outputibias.n65 0.155672
R23421 outputibias.n86 outputibias.n85 0.155672
R23422 outputibias.n85 outputibias.n69 0.155672
R23423 outputibias.n78 outputibias.n69 0.155672
R23424 outputibias.n78 outputibias.n77 0.155672
R23425 outputibias.n125 outputibias.n97 0.155672
R23426 outputibias.n118 outputibias.n97 0.155672
R23427 outputibias.n118 outputibias.n117 0.155672
R23428 outputibias.n117 outputibias.n101 0.155672
R23429 outputibias.n110 outputibias.n101 0.155672
R23430 outputibias.n110 outputibias.n109 0.155672
C0 output outputibias 2.34152f
C1 vdd output 7.23429f
C2 CSoutput output 6.13571f
C3 CSoutput outputibias 0.032386f
C4 vdd CSoutput 0.116919p
C5 minus diffpairibias 2.98e-19
C6 commonsourceibias output 0.006808f
C7 vdd plus 0.08876f
C8 CSoutput minus 3.02748f
C9 plus diffpairibias 2.75e-19
C10 commonsourceibias outputibias 0.003832f
C11 vdd commonsourceibias 0.004218f
C12 CSoutput plus 0.872047f
C13 commonsourceibias diffpairibias 0.052527f
C14 CSoutput commonsourceibias 37.4715f
C15 minus plus 9.47051f
C16 minus commonsourceibias 0.331305f
C17 plus commonsourceibias 0.276969f
C18 diffpairibias gnd 59.991135f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.150748p
C22 plus gnd 34.01f
C23 minus gnd 28.691391f
C24 CSoutput gnd 0.102317p
C25 vdd gnd 0.477765p
C26 outputibias.t10 gnd 0.11477f
C27 outputibias.t8 gnd 0.115567f
C28 outputibias.n0 gnd 0.130108f
C29 outputibias.n1 gnd 0.001372f
C30 outputibias.n2 gnd 9.76e-19
C31 outputibias.n3 gnd 5.24e-19
C32 outputibias.n4 gnd 0.001239f
C33 outputibias.n5 gnd 5.55e-19
C34 outputibias.n6 gnd 9.76e-19
C35 outputibias.n7 gnd 5.24e-19
C36 outputibias.n8 gnd 0.001239f
C37 outputibias.n9 gnd 5.55e-19
C38 outputibias.n10 gnd 0.004176f
C39 outputibias.t5 gnd 0.00202f
C40 outputibias.n11 gnd 9.3e-19
C41 outputibias.n12 gnd 7.32e-19
C42 outputibias.n13 gnd 5.24e-19
C43 outputibias.n14 gnd 0.02322f
C44 outputibias.n15 gnd 9.76e-19
C45 outputibias.n16 gnd 5.24e-19
C46 outputibias.n17 gnd 5.55e-19
C47 outputibias.n18 gnd 0.001239f
C48 outputibias.n19 gnd 0.001239f
C49 outputibias.n20 gnd 5.55e-19
C50 outputibias.n21 gnd 5.24e-19
C51 outputibias.n22 gnd 9.76e-19
C52 outputibias.n23 gnd 9.76e-19
C53 outputibias.n24 gnd 5.24e-19
C54 outputibias.n25 gnd 5.55e-19
C55 outputibias.n26 gnd 0.001239f
C56 outputibias.n27 gnd 0.002683f
C57 outputibias.n28 gnd 5.55e-19
C58 outputibias.n29 gnd 5.24e-19
C59 outputibias.n30 gnd 0.002256f
C60 outputibias.n31 gnd 0.005781f
C61 outputibias.n32 gnd 0.001372f
C62 outputibias.n33 gnd 9.76e-19
C63 outputibias.n34 gnd 5.24e-19
C64 outputibias.n35 gnd 0.001239f
C65 outputibias.n36 gnd 5.55e-19
C66 outputibias.n37 gnd 9.76e-19
C67 outputibias.n38 gnd 5.24e-19
C68 outputibias.n39 gnd 0.001239f
C69 outputibias.n40 gnd 5.55e-19
C70 outputibias.n41 gnd 0.004176f
C71 outputibias.t7 gnd 0.00202f
C72 outputibias.n42 gnd 9.3e-19
C73 outputibias.n43 gnd 7.32e-19
C74 outputibias.n44 gnd 5.24e-19
C75 outputibias.n45 gnd 0.02322f
C76 outputibias.n46 gnd 9.76e-19
C77 outputibias.n47 gnd 5.24e-19
C78 outputibias.n48 gnd 5.55e-19
C79 outputibias.n49 gnd 0.001239f
C80 outputibias.n50 gnd 0.001239f
C81 outputibias.n51 gnd 5.55e-19
C82 outputibias.n52 gnd 5.24e-19
C83 outputibias.n53 gnd 9.76e-19
C84 outputibias.n54 gnd 9.76e-19
C85 outputibias.n55 gnd 5.24e-19
C86 outputibias.n56 gnd 5.55e-19
C87 outputibias.n57 gnd 0.001239f
C88 outputibias.n58 gnd 0.002683f
C89 outputibias.n59 gnd 5.55e-19
C90 outputibias.n60 gnd 5.24e-19
C91 outputibias.n61 gnd 0.002256f
C92 outputibias.n62 gnd 0.005197f
C93 outputibias.n63 gnd 0.121892f
C94 outputibias.n64 gnd 0.001372f
C95 outputibias.n65 gnd 9.76e-19
C96 outputibias.n66 gnd 5.24e-19
C97 outputibias.n67 gnd 0.001239f
C98 outputibias.n68 gnd 5.55e-19
C99 outputibias.n69 gnd 9.76e-19
C100 outputibias.n70 gnd 5.24e-19
C101 outputibias.n71 gnd 0.001239f
C102 outputibias.n72 gnd 5.55e-19
C103 outputibias.n73 gnd 0.004176f
C104 outputibias.t1 gnd 0.00202f
C105 outputibias.n74 gnd 9.3e-19
C106 outputibias.n75 gnd 7.32e-19
C107 outputibias.n76 gnd 5.24e-19
C108 outputibias.n77 gnd 0.02322f
C109 outputibias.n78 gnd 9.76e-19
C110 outputibias.n79 gnd 5.24e-19
C111 outputibias.n80 gnd 5.55e-19
C112 outputibias.n81 gnd 0.001239f
C113 outputibias.n82 gnd 0.001239f
C114 outputibias.n83 gnd 5.55e-19
C115 outputibias.n84 gnd 5.24e-19
C116 outputibias.n85 gnd 9.76e-19
C117 outputibias.n86 gnd 9.76e-19
C118 outputibias.n87 gnd 5.24e-19
C119 outputibias.n88 gnd 5.55e-19
C120 outputibias.n89 gnd 0.001239f
C121 outputibias.n90 gnd 0.002683f
C122 outputibias.n91 gnd 5.55e-19
C123 outputibias.n92 gnd 5.24e-19
C124 outputibias.n93 gnd 0.002256f
C125 outputibias.n94 gnd 0.005197f
C126 outputibias.n95 gnd 0.064513f
C127 outputibias.n96 gnd 0.001372f
C128 outputibias.n97 gnd 9.76e-19
C129 outputibias.n98 gnd 5.24e-19
C130 outputibias.n99 gnd 0.001239f
C131 outputibias.n100 gnd 5.55e-19
C132 outputibias.n101 gnd 9.76e-19
C133 outputibias.n102 gnd 5.24e-19
C134 outputibias.n103 gnd 0.001239f
C135 outputibias.n104 gnd 5.55e-19
C136 outputibias.n105 gnd 0.004176f
C137 outputibias.t3 gnd 0.00202f
C138 outputibias.n106 gnd 9.3e-19
C139 outputibias.n107 gnd 7.32e-19
C140 outputibias.n108 gnd 5.24e-19
C141 outputibias.n109 gnd 0.02322f
C142 outputibias.n110 gnd 9.76e-19
C143 outputibias.n111 gnd 5.24e-19
C144 outputibias.n112 gnd 5.55e-19
C145 outputibias.n113 gnd 0.001239f
C146 outputibias.n114 gnd 0.001239f
C147 outputibias.n115 gnd 5.55e-19
C148 outputibias.n116 gnd 5.24e-19
C149 outputibias.n117 gnd 9.76e-19
C150 outputibias.n118 gnd 9.76e-19
C151 outputibias.n119 gnd 5.24e-19
C152 outputibias.n120 gnd 5.55e-19
C153 outputibias.n121 gnd 0.001239f
C154 outputibias.n122 gnd 0.002683f
C155 outputibias.n123 gnd 5.55e-19
C156 outputibias.n124 gnd 5.24e-19
C157 outputibias.n125 gnd 0.002256f
C158 outputibias.n126 gnd 0.005197f
C159 outputibias.n127 gnd 0.084814f
C160 outputibias.t2 gnd 0.108319f
C161 outputibias.t0 gnd 0.108319f
C162 outputibias.t6 gnd 0.108319f
C163 outputibias.t4 gnd 0.109238f
C164 outputibias.n128 gnd 0.134674f
C165 outputibias.n129 gnd 0.07244f
C166 outputibias.n130 gnd 0.079818f
C167 outputibias.n131 gnd 0.164901f
C168 outputibias.t9 gnd 0.11477f
C169 outputibias.n132 gnd 0.067481f
C170 outputibias.t11 gnd 0.11477f
C171 outputibias.n133 gnd 0.065115f
C172 outputibias.n134 gnd 0.029159f
C173 minus.n0 gnd 0.032264f
C174 minus.t27 gnd 0.325958f
C175 minus.n1 gnd 0.150402f
C176 minus.n2 gnd 0.032264f
C177 minus.t6 gnd 0.325958f
C178 minus.n3 gnd 0.147418f
C179 minus.n4 gnd 0.032264f
C180 minus.t24 gnd 0.325958f
C181 minus.n5 gnd 0.147418f
C182 minus.n6 gnd 0.032264f
C183 minus.t8 gnd 0.325958f
C184 minus.n7 gnd 0.150402f
C185 minus.t12 gnd 0.334734f
C186 minus.t18 gnd 0.325958f
C187 minus.n8 gnd 0.15422f
C188 minus.n9 gnd 0.1396f
C189 minus.n10 gnd 0.131004f
C190 minus.n11 gnd 0.032264f
C191 minus.n12 gnd 0.007321f
C192 minus.t13 gnd 0.325958f
C193 minus.n13 gnd 0.1507f
C194 minus.n14 gnd 0.007321f
C195 minus.n15 gnd 0.032264f
C196 minus.n16 gnd 0.032264f
C197 minus.n17 gnd 0.032264f
C198 minus.t19 gnd 0.325958f
C199 minus.n18 gnd 0.150601f
C200 minus.n19 gnd 0.007321f
C201 minus.t22 gnd 0.325958f
C202 minus.n20 gnd 0.150601f
C203 minus.n21 gnd 0.032264f
C204 minus.n22 gnd 0.032264f
C205 minus.n23 gnd 0.032264f
C206 minus.n24 gnd 0.007321f
C207 minus.t20 gnd 0.325958f
C208 minus.n25 gnd 0.1507f
C209 minus.n26 gnd 0.007321f
C210 minus.n27 gnd 0.032264f
C211 minus.n28 gnd 0.032264f
C212 minus.n29 gnd 0.032264f
C213 minus.t15 gnd 0.325958f
C214 minus.n30 gnd 0.147617f
C215 minus.n31 gnd 0.007321f
C216 minus.t9 gnd 0.325958f
C217 minus.n32 gnd 0.14702f
C218 minus.n33 gnd 0.362089f
C219 minus.n34 gnd 0.032264f
C220 minus.t16 gnd 0.325958f
C221 minus.t28 gnd 0.325958f
C222 minus.n35 gnd 0.032264f
C223 minus.t21 gnd 0.325958f
C224 minus.n36 gnd 0.032264f
C225 minus.t14 gnd 0.325958f
C226 minus.n37 gnd 0.1507f
C227 minus.n38 gnd 0.032264f
C228 minus.t23 gnd 0.325958f
C229 minus.t11 gnd 0.325958f
C230 minus.n39 gnd 0.032264f
C231 minus.t5 gnd 0.325958f
C232 minus.n40 gnd 0.150601f
C233 minus.n41 gnd 0.032264f
C234 minus.t17 gnd 0.325958f
C235 minus.t10 gnd 0.325958f
C236 minus.n42 gnd 0.032264f
C237 minus.t25 gnd 0.325958f
C238 minus.n43 gnd 0.150402f
C239 minus.t26 gnd 0.334734f
C240 minus.t7 gnd 0.325958f
C241 minus.n44 gnd 0.15422f
C242 minus.n45 gnd 0.1396f
C243 minus.n46 gnd 0.131004f
C244 minus.n47 gnd 0.032264f
C245 minus.n48 gnd 0.007321f
C246 minus.n49 gnd 0.1507f
C247 minus.n50 gnd 0.007321f
C248 minus.n51 gnd 0.147418f
C249 minus.n52 gnd 0.032264f
C250 minus.n53 gnd 0.032264f
C251 minus.n54 gnd 0.032264f
C252 minus.n55 gnd 0.007321f
C253 minus.n56 gnd 0.150601f
C254 minus.n57 gnd 0.147418f
C255 minus.n58 gnd 0.007321f
C256 minus.n59 gnd 0.032264f
C257 minus.n60 gnd 0.032264f
C258 minus.n61 gnd 0.032264f
C259 minus.n62 gnd 0.007321f
C260 minus.n63 gnd 0.150402f
C261 minus.n64 gnd 0.147617f
C262 minus.n65 gnd 0.007321f
C263 minus.n66 gnd 0.14702f
C264 minus.n67 gnd 0.979055f
C265 minus.n68 gnd 1.48514f
C266 minus.t1 gnd 0.009946f
C267 minus.t4 gnd 0.009946f
C268 minus.n69 gnd 0.032705f
C269 minus.t2 gnd 0.009946f
C270 minus.t0 gnd 0.009946f
C271 minus.n70 gnd 0.032256f
C272 minus.n71 gnd 0.275295f
C273 minus.t3 gnd 0.055358f
C274 minus.n72 gnd 0.150226f
C275 minus.n73 gnd 2.26062f
C276 plus.n0 gnd 0.023469f
C277 plus.t23 gnd 0.237103f
C278 plus.n1 gnd 0.023469f
C279 plus.t13 gnd 0.237103f
C280 plus.n2 gnd 0.023469f
C281 plus.t27 gnd 0.237103f
C282 plus.t22 gnd 0.237103f
C283 plus.n3 gnd 0.10962f
C284 plus.n4 gnd 0.023469f
C285 plus.t7 gnd 0.237103f
C286 plus.n5 gnd 0.023469f
C287 plus.t18 gnd 0.237103f
C288 plus.t14 gnd 0.237103f
C289 plus.n6 gnd 0.109548f
C290 plus.n7 gnd 0.023469f
C291 plus.t24 gnd 0.237103f
C292 plus.n8 gnd 0.023469f
C293 plus.t17 gnd 0.237103f
C294 plus.t9 gnd 0.237103f
C295 plus.n9 gnd 0.109403f
C296 plus.t12 gnd 0.243487f
C297 plus.t15 gnd 0.237103f
C298 plus.n10 gnd 0.11218f
C299 plus.n11 gnd 0.101546f
C300 plus.n12 gnd 0.095293f
C301 plus.n13 gnd 0.023469f
C302 plus.n14 gnd 0.005326f
C303 plus.n15 gnd 0.10962f
C304 plus.n16 gnd 0.005326f
C305 plus.n17 gnd 0.107233f
C306 plus.n18 gnd 0.023469f
C307 plus.n19 gnd 0.023469f
C308 plus.n20 gnd 0.023469f
C309 plus.n21 gnd 0.005326f
C310 plus.n22 gnd 0.109548f
C311 plus.n23 gnd 0.107233f
C312 plus.n24 gnd 0.005326f
C313 plus.n25 gnd 0.023469f
C314 plus.n26 gnd 0.023469f
C315 plus.n27 gnd 0.023469f
C316 plus.n28 gnd 0.005326f
C317 plus.n29 gnd 0.109403f
C318 plus.n30 gnd 0.107377f
C319 plus.n31 gnd 0.005326f
C320 plus.n32 gnd 0.106943f
C321 plus.n33 gnd 0.257321f
C322 plus.n34 gnd 0.023469f
C323 plus.t16 gnd 0.237103f
C324 plus.n35 gnd 0.109403f
C325 plus.t28 gnd 0.237103f
C326 plus.n36 gnd 0.023469f
C327 plus.t19 gnd 0.237103f
C328 plus.n37 gnd 0.107233f
C329 plus.n38 gnd 0.023469f
C330 plus.t11 gnd 0.237103f
C331 plus.n39 gnd 0.107233f
C332 plus.t6 gnd 0.237103f
C333 plus.n40 gnd 0.023469f
C334 plus.t20 gnd 0.237103f
C335 plus.n41 gnd 0.109403f
C336 plus.t25 gnd 0.243487f
C337 plus.t5 gnd 0.237103f
C338 plus.n42 gnd 0.11218f
C339 plus.n43 gnd 0.101546f
C340 plus.n44 gnd 0.095293f
C341 plus.n45 gnd 0.023469f
C342 plus.n46 gnd 0.005326f
C343 plus.t26 gnd 0.237103f
C344 plus.n47 gnd 0.10962f
C345 plus.n48 gnd 0.005326f
C346 plus.n49 gnd 0.023469f
C347 plus.n50 gnd 0.023469f
C348 plus.n51 gnd 0.023469f
C349 plus.n52 gnd 0.109548f
C350 plus.n53 gnd 0.005326f
C351 plus.t10 gnd 0.237103f
C352 plus.n54 gnd 0.109548f
C353 plus.n55 gnd 0.023469f
C354 plus.n56 gnd 0.023469f
C355 plus.n57 gnd 0.023469f
C356 plus.n58 gnd 0.005326f
C357 plus.t8 gnd 0.237103f
C358 plus.n59 gnd 0.10962f
C359 plus.n60 gnd 0.005326f
C360 plus.n61 gnd 0.023469f
C361 plus.n62 gnd 0.023469f
C362 plus.n63 gnd 0.023469f
C363 plus.n64 gnd 0.107377f
C364 plus.n65 gnd 0.005326f
C365 plus.t21 gnd 0.237103f
C366 plus.n66 gnd 0.106943f
C367 plus.n67 gnd 0.702732f
C368 plus.n68 gnd 1.07105f
C369 plus.t3 gnd 0.040514f
C370 plus.t4 gnd 0.007235f
C371 plus.t1 gnd 0.007235f
C372 plus.n69 gnd 0.023463f
C373 plus.n70 gnd 0.182149f
C374 plus.t0 gnd 0.007235f
C375 plus.t2 gnd 0.007235f
C376 plus.n71 gnd 0.023463f
C377 plus.n72 gnd 0.136725f
C378 plus.n73 gnd 2.83731f
C379 a_n2650_8322.t13 gnd 0.097992f
C380 a_n2650_8322.t31 gnd 20.329401f
C381 a_n2650_8322.t33 gnd 20.186901f
C382 a_n2650_8322.t30 gnd 20.186901f
C383 a_n2650_8322.t29 gnd 20.329401f
C384 a_n2650_8322.t32 gnd 20.186901f
C385 a_n2650_8322.t28 gnd 29.294302f
C386 a_n2650_8322.t23 gnd 0.917551f
C387 a_n2650_8322.t26 gnd 0.097992f
C388 a_n2650_8322.t18 gnd 0.097992f
C389 a_n2650_8322.n0 gnd 0.690258f
C390 a_n2650_8322.n1 gnd 0.771262f
C391 a_n2650_8322.t10 gnd 0.097992f
C392 a_n2650_8322.t9 gnd 0.097992f
C393 a_n2650_8322.n2 gnd 0.690258f
C394 a_n2650_8322.n3 gnd 0.391868f
C395 a_n2650_8322.t21 gnd 0.097992f
C396 a_n2650_8322.t15 gnd 0.097992f
C397 a_n2650_8322.n4 gnd 0.690258f
C398 a_n2650_8322.n5 gnd 0.391868f
C399 a_n2650_8322.t19 gnd 0.097992f
C400 a_n2650_8322.t17 gnd 0.097992f
C401 a_n2650_8322.n6 gnd 0.690258f
C402 a_n2650_8322.n7 gnd 0.391868f
C403 a_n2650_8322.t8 gnd 0.915724f
C404 a_n2650_8322.n8 gnd 1.70884f
C405 a_n2650_8322.t3 gnd 0.917551f
C406 a_n2650_8322.t7 gnd 0.097992f
C407 a_n2650_8322.t6 gnd 0.097992f
C408 a_n2650_8322.n9 gnd 0.690258f
C409 a_n2650_8322.n10 gnd 0.771262f
C410 a_n2650_8322.t1 gnd 0.915724f
C411 a_n2650_8322.n11 gnd 0.38811f
C412 a_n2650_8322.t4 gnd 0.915724f
C413 a_n2650_8322.n12 gnd 0.38811f
C414 a_n2650_8322.t2 gnd 0.097992f
C415 a_n2650_8322.t0 gnd 0.097992f
C416 a_n2650_8322.n13 gnd 0.690258f
C417 a_n2650_8322.n14 gnd 0.391868f
C418 a_n2650_8322.t5 gnd 0.915724f
C419 a_n2650_8322.n15 gnd 1.27333f
C420 a_n2650_8322.n16 gnd 2.0805f
C421 a_n2650_8322.n17 gnd 3.60069f
C422 a_n2650_8322.t22 gnd 0.915724f
C423 a_n2650_8322.n18 gnd 0.996043f
C424 a_n2650_8322.t12 gnd 0.097992f
C425 a_n2650_8322.t11 gnd 0.097992f
C426 a_n2650_8322.n19 gnd 0.690258f
C427 a_n2650_8322.n20 gnd 0.391868f
C428 a_n2650_8322.t24 gnd 0.097992f
C429 a_n2650_8322.t14 gnd 0.097992f
C430 a_n2650_8322.n21 gnd 0.690258f
C431 a_n2650_8322.n22 gnd 0.391868f
C432 a_n2650_8322.t25 gnd 0.917548f
C433 a_n2650_8322.t20 gnd 0.097992f
C434 a_n2650_8322.t16 gnd 0.097992f
C435 a_n2650_8322.n23 gnd 0.690258f
C436 a_n2650_8322.n24 gnd 0.771264f
C437 a_n2650_8322.n25 gnd 0.391867f
C438 a_n2650_8322.n26 gnd 0.69026f
C439 a_n2650_8322.t27 gnd 0.097992f
C440 output.t15 gnd 0.464308f
C441 output.t5 gnd 0.044422f
C442 output.t9 gnd 0.044422f
C443 output.n0 gnd 0.364624f
C444 output.n1 gnd 0.614102f
C445 output.t12 gnd 0.044422f
C446 output.t17 gnd 0.044422f
C447 output.n2 gnd 0.364624f
C448 output.n3 gnd 0.350265f
C449 output.t18 gnd 0.044422f
C450 output.t7 gnd 0.044422f
C451 output.n4 gnd 0.364624f
C452 output.n5 gnd 0.350265f
C453 output.t11 gnd 0.044422f
C454 output.t3 gnd 0.044422f
C455 output.n6 gnd 0.364624f
C456 output.n7 gnd 0.350265f
C457 output.t6 gnd 0.044422f
C458 output.t4 gnd 0.044422f
C459 output.n8 gnd 0.364624f
C460 output.n9 gnd 0.350265f
C461 output.t10 gnd 0.044422f
C462 output.t13 gnd 0.044422f
C463 output.n10 gnd 0.364624f
C464 output.n11 gnd 0.350265f
C465 output.t14 gnd 0.044422f
C466 output.t8 gnd 0.044422f
C467 output.n12 gnd 0.364624f
C468 output.n13 gnd 0.350265f
C469 output.t16 gnd 0.462979f
C470 output.n14 gnd 0.28994f
C471 output.n15 gnd 0.015803f
C472 output.n16 gnd 0.011243f
C473 output.n17 gnd 0.006041f
C474 output.n18 gnd 0.01428f
C475 output.n19 gnd 0.006397f
C476 output.n20 gnd 0.011243f
C477 output.n21 gnd 0.006041f
C478 output.n22 gnd 0.01428f
C479 output.n23 gnd 0.006397f
C480 output.n24 gnd 0.048111f
C481 output.t2 gnd 0.023274f
C482 output.n25 gnd 0.01071f
C483 output.n26 gnd 0.008435f
C484 output.n27 gnd 0.006041f
C485 output.n28 gnd 0.267512f
C486 output.n29 gnd 0.011243f
C487 output.n30 gnd 0.006041f
C488 output.n31 gnd 0.006397f
C489 output.n32 gnd 0.01428f
C490 output.n33 gnd 0.01428f
C491 output.n34 gnd 0.006397f
C492 output.n35 gnd 0.006041f
C493 output.n36 gnd 0.011243f
C494 output.n37 gnd 0.011243f
C495 output.n38 gnd 0.006041f
C496 output.n39 gnd 0.006397f
C497 output.n40 gnd 0.01428f
C498 output.n41 gnd 0.030913f
C499 output.n42 gnd 0.006397f
C500 output.n43 gnd 0.006041f
C501 output.n44 gnd 0.025987f
C502 output.n45 gnd 0.097665f
C503 output.n46 gnd 0.015803f
C504 output.n47 gnd 0.011243f
C505 output.n48 gnd 0.006041f
C506 output.n49 gnd 0.01428f
C507 output.n50 gnd 0.006397f
C508 output.n51 gnd 0.011243f
C509 output.n52 gnd 0.006041f
C510 output.n53 gnd 0.01428f
C511 output.n54 gnd 0.006397f
C512 output.n55 gnd 0.048111f
C513 output.t19 gnd 0.023274f
C514 output.n56 gnd 0.01071f
C515 output.n57 gnd 0.008435f
C516 output.n58 gnd 0.006041f
C517 output.n59 gnd 0.267512f
C518 output.n60 gnd 0.011243f
C519 output.n61 gnd 0.006041f
C520 output.n62 gnd 0.006397f
C521 output.n63 gnd 0.01428f
C522 output.n64 gnd 0.01428f
C523 output.n65 gnd 0.006397f
C524 output.n66 gnd 0.006041f
C525 output.n67 gnd 0.011243f
C526 output.n68 gnd 0.011243f
C527 output.n69 gnd 0.006041f
C528 output.n70 gnd 0.006397f
C529 output.n71 gnd 0.01428f
C530 output.n72 gnd 0.030913f
C531 output.n73 gnd 0.006397f
C532 output.n74 gnd 0.006041f
C533 output.n75 gnd 0.025987f
C534 output.n76 gnd 0.09306f
C535 output.n77 gnd 1.65264f
C536 output.n78 gnd 0.015803f
C537 output.n79 gnd 0.011243f
C538 output.n80 gnd 0.006041f
C539 output.n81 gnd 0.01428f
C540 output.n82 gnd 0.006397f
C541 output.n83 gnd 0.011243f
C542 output.n84 gnd 0.006041f
C543 output.n85 gnd 0.01428f
C544 output.n86 gnd 0.006397f
C545 output.n87 gnd 0.048111f
C546 output.t0 gnd 0.023274f
C547 output.n88 gnd 0.01071f
C548 output.n89 gnd 0.008435f
C549 output.n90 gnd 0.006041f
C550 output.n91 gnd 0.267512f
C551 output.n92 gnd 0.011243f
C552 output.n93 gnd 0.006041f
C553 output.n94 gnd 0.006397f
C554 output.n95 gnd 0.01428f
C555 output.n96 gnd 0.01428f
C556 output.n97 gnd 0.006397f
C557 output.n98 gnd 0.006041f
C558 output.n99 gnd 0.011243f
C559 output.n100 gnd 0.011243f
C560 output.n101 gnd 0.006041f
C561 output.n102 gnd 0.006397f
C562 output.n103 gnd 0.01428f
C563 output.n104 gnd 0.030913f
C564 output.n105 gnd 0.006397f
C565 output.n106 gnd 0.006041f
C566 output.n107 gnd 0.025987f
C567 output.n108 gnd 0.09306f
C568 output.n109 gnd 0.713089f
C569 output.n110 gnd 0.015803f
C570 output.n111 gnd 0.011243f
C571 output.n112 gnd 0.006041f
C572 output.n113 gnd 0.01428f
C573 output.n114 gnd 0.006397f
C574 output.n115 gnd 0.011243f
C575 output.n116 gnd 0.006041f
C576 output.n117 gnd 0.01428f
C577 output.n118 gnd 0.006397f
C578 output.n119 gnd 0.048111f
C579 output.t1 gnd 0.023274f
C580 output.n120 gnd 0.01071f
C581 output.n121 gnd 0.008435f
C582 output.n122 gnd 0.006041f
C583 output.n123 gnd 0.267512f
C584 output.n124 gnd 0.011243f
C585 output.n125 gnd 0.006041f
C586 output.n126 gnd 0.006397f
C587 output.n127 gnd 0.01428f
C588 output.n128 gnd 0.01428f
C589 output.n129 gnd 0.006397f
C590 output.n130 gnd 0.006041f
C591 output.n131 gnd 0.011243f
C592 output.n132 gnd 0.011243f
C593 output.n133 gnd 0.006041f
C594 output.n134 gnd 0.006397f
C595 output.n135 gnd 0.01428f
C596 output.n136 gnd 0.030913f
C597 output.n137 gnd 0.006397f
C598 output.n138 gnd 0.006041f
C599 output.n139 gnd 0.025987f
C600 output.n140 gnd 0.09306f
C601 output.n141 gnd 1.67353f
C602 a_n3827_n3924.n0 gnd 1.10033f
C603 a_n3827_n3924.n1 gnd 0.958536f
C604 a_n3827_n3924.t9 gnd 1.06719f
C605 a_n3827_n3924.n2 gnd 0.920943f
C606 a_n3827_n3924.t31 gnd 0.102682f
C607 a_n3827_n3924.t25 gnd 0.102682f
C608 a_n3827_n3924.n3 gnd 0.838616f
C609 a_n3827_n3924.n4 gnd 0.340114f
C610 a_n3827_n3924.t6 gnd 0.102682f
C611 a_n3827_n3924.t22 gnd 0.102682f
C612 a_n3827_n3924.n5 gnd 0.838616f
C613 a_n3827_n3924.n6 gnd 0.340114f
C614 a_n3827_n3924.t48 gnd 0.102682f
C615 a_n3827_n3924.t42 gnd 0.102682f
C616 a_n3827_n3924.n7 gnd 0.838616f
C617 a_n3827_n3924.n8 gnd 0.340114f
C618 a_n3827_n3924.t46 gnd 0.102682f
C619 a_n3827_n3924.t7 gnd 0.102682f
C620 a_n3827_n3924.n9 gnd 0.838616f
C621 a_n3827_n3924.n10 gnd 0.340114f
C622 a_n3827_n3924.t40 gnd 0.102682f
C623 a_n3827_n3924.t8 gnd 0.102682f
C624 a_n3827_n3924.n11 gnd 0.838616f
C625 a_n3827_n3924.n12 gnd 0.340114f
C626 a_n3827_n3924.t39 gnd 1.06719f
C627 a_n3827_n3924.n13 gnd 0.362194f
C628 a_n3827_n3924.t0 gnd 1.06719f
C629 a_n3827_n3924.n14 gnd 0.362194f
C630 a_n3827_n3924.t38 gnd 0.102682f
C631 a_n3827_n3924.t34 gnd 0.102682f
C632 a_n3827_n3924.n15 gnd 0.838616f
C633 a_n3827_n3924.n16 gnd 0.340114f
C634 a_n3827_n3924.t26 gnd 0.102682f
C635 a_n3827_n3924.t27 gnd 0.102682f
C636 a_n3827_n3924.n17 gnd 0.838616f
C637 a_n3827_n3924.n18 gnd 0.340114f
C638 a_n3827_n3924.t35 gnd 0.102682f
C639 a_n3827_n3924.t56 gnd 0.102682f
C640 a_n3827_n3924.n19 gnd 0.838616f
C641 a_n3827_n3924.n20 gnd 0.340114f
C642 a_n3827_n3924.t37 gnd 0.102682f
C643 a_n3827_n3924.t53 gnd 0.102682f
C644 a_n3827_n3924.n21 gnd 0.838616f
C645 a_n3827_n3924.n22 gnd 0.340114f
C646 a_n3827_n3924.t23 gnd 0.102682f
C647 a_n3827_n3924.t55 gnd 0.102682f
C648 a_n3827_n3924.n23 gnd 0.838616f
C649 a_n3827_n3924.n24 gnd 0.340114f
C650 a_n3827_n3924.t36 gnd 1.06718f
C651 a_n3827_n3924.n25 gnd 0.920947f
C652 a_n3827_n3924.t2 gnd 1.06718f
C653 a_n3827_n3924.n26 gnd 0.58539f
C654 a_n3827_n3924.t44 gnd 0.102682f
C655 a_n3827_n3924.t52 gnd 0.102682f
C656 a_n3827_n3924.n27 gnd 0.838615f
C657 a_n3827_n3924.n28 gnd 0.340116f
C658 a_n3827_n3924.t10 gnd 0.102682f
C659 a_n3827_n3924.t57 gnd 0.102682f
C660 a_n3827_n3924.n29 gnd 0.838615f
C661 a_n3827_n3924.n30 gnd 0.340116f
C662 a_n3827_n3924.t29 gnd 0.102682f
C663 a_n3827_n3924.t1 gnd 0.102682f
C664 a_n3827_n3924.n31 gnd 0.838615f
C665 a_n3827_n3924.n32 gnd 0.340116f
C666 a_n3827_n3924.t33 gnd 0.102682f
C667 a_n3827_n3924.t30 gnd 0.102682f
C668 a_n3827_n3924.n33 gnd 0.838615f
C669 a_n3827_n3924.n34 gnd 0.340116f
C670 a_n3827_n3924.t54 gnd 0.102682f
C671 a_n3827_n3924.t3 gnd 0.102682f
C672 a_n3827_n3924.n35 gnd 0.838615f
C673 a_n3827_n3924.n36 gnd 0.340116f
C674 a_n3827_n3924.t28 gnd 1.06718f
C675 a_n3827_n3924.n37 gnd 0.362198f
C676 a_n3827_n3924.t51 gnd 1.06718f
C677 a_n3827_n3924.n38 gnd 0.362198f
C678 a_n3827_n3924.t49 gnd 0.102682f
C679 a_n3827_n3924.t5 gnd 0.102682f
C680 a_n3827_n3924.n39 gnd 0.838615f
C681 a_n3827_n3924.n40 gnd 0.340116f
C682 a_n3827_n3924.t47 gnd 0.102682f
C683 a_n3827_n3924.t32 gnd 0.102682f
C684 a_n3827_n3924.n41 gnd 0.838615f
C685 a_n3827_n3924.n42 gnd 0.340116f
C686 a_n3827_n3924.t43 gnd 0.102682f
C687 a_n3827_n3924.t41 gnd 0.102682f
C688 a_n3827_n3924.n43 gnd 0.838615f
C689 a_n3827_n3924.n44 gnd 0.340116f
C690 a_n3827_n3924.t50 gnd 0.102682f
C691 a_n3827_n3924.t45 gnd 0.102682f
C692 a_n3827_n3924.n45 gnd 0.838615f
C693 a_n3827_n3924.n46 gnd 0.340116f
C694 a_n3827_n3924.t21 gnd 0.102682f
C695 a_n3827_n3924.t4 gnd 0.102682f
C696 a_n3827_n3924.n47 gnd 0.838615f
C697 a_n3827_n3924.n48 gnd 0.340116f
C698 a_n3827_n3924.t24 gnd 1.06718f
C699 a_n3827_n3924.n49 gnd 0.58539f
C700 a_n3827_n3924.n50 gnd 0.958536f
C701 a_n3827_n3924.t13 gnd 1.32959f
C702 a_n3827_n3924.t17 gnd 1.32595f
C703 a_n3827_n3924.n51 gnd 1.82937f
C704 a_n3827_n3924.n52 gnd 0.504753f
C705 a_n3827_n3924.t12 gnd 1.32595f
C706 a_n3827_n3924.n53 gnd 0.844057f
C707 a_n3827_n3924.t15 gnd 1.32595f
C708 a_n3827_n3924.n54 gnd 0.933892f
C709 a_n3827_n3924.t11 gnd 1.32595f
C710 a_n3827_n3924.n55 gnd 0.933892f
C711 a_n3827_n3924.t16 gnd 1.32595f
C712 a_n3827_n3924.n56 gnd 0.933892f
C713 a_n3827_n3924.t19 gnd 1.32595f
C714 a_n3827_n3924.n57 gnd 0.918983f
C715 a_n3827_n3924.t18 gnd 1.32595f
C716 a_n3827_n3924.t14 gnd 1.32595f
C717 a_n3827_n3924.n58 gnd 1.5379f
C718 a_n3827_n3924.t20 gnd 1.32785f
C719 diffpairibias.t27 gnd 0.090128f
C720 diffpairibias.t23 gnd 0.08996f
C721 diffpairibias.n0 gnd 0.105991f
C722 diffpairibias.t28 gnd 0.08996f
C723 diffpairibias.n1 gnd 0.051736f
C724 diffpairibias.t25 gnd 0.08996f
C725 diffpairibias.n2 gnd 0.051736f
C726 diffpairibias.t29 gnd 0.08996f
C727 diffpairibias.n3 gnd 0.041084f
C728 diffpairibias.t15 gnd 0.086371f
C729 diffpairibias.t1 gnd 0.085993f
C730 diffpairibias.n4 gnd 0.13579f
C731 diffpairibias.t11 gnd 0.085993f
C732 diffpairibias.n5 gnd 0.072463f
C733 diffpairibias.t13 gnd 0.085993f
C734 diffpairibias.n6 gnd 0.072463f
C735 diffpairibias.t7 gnd 0.085993f
C736 diffpairibias.n7 gnd 0.072463f
C737 diffpairibias.t3 gnd 0.085993f
C738 diffpairibias.n8 gnd 0.072463f
C739 diffpairibias.t17 gnd 0.085993f
C740 diffpairibias.n9 gnd 0.072463f
C741 diffpairibias.t5 gnd 0.085993f
C742 diffpairibias.n10 gnd 0.072463f
C743 diffpairibias.t19 gnd 0.085993f
C744 diffpairibias.n11 gnd 0.072463f
C745 diffpairibias.t9 gnd 0.085993f
C746 diffpairibias.n12 gnd 0.102883f
C747 diffpairibias.t14 gnd 0.086899f
C748 diffpairibias.t0 gnd 0.086748f
C749 diffpairibias.n13 gnd 0.094648f
C750 diffpairibias.t10 gnd 0.086748f
C751 diffpairibias.n14 gnd 0.052262f
C752 diffpairibias.t12 gnd 0.086748f
C753 diffpairibias.n15 gnd 0.052262f
C754 diffpairibias.t6 gnd 0.086748f
C755 diffpairibias.n16 gnd 0.052262f
C756 diffpairibias.t2 gnd 0.086748f
C757 diffpairibias.n17 gnd 0.052262f
C758 diffpairibias.t16 gnd 0.086748f
C759 diffpairibias.n18 gnd 0.052262f
C760 diffpairibias.t4 gnd 0.086748f
C761 diffpairibias.n19 gnd 0.052262f
C762 diffpairibias.t18 gnd 0.086748f
C763 diffpairibias.n20 gnd 0.052262f
C764 diffpairibias.t8 gnd 0.086748f
C765 diffpairibias.n21 gnd 0.061849f
C766 diffpairibias.n22 gnd 0.233513f
C767 diffpairibias.t20 gnd 0.08996f
C768 diffpairibias.n23 gnd 0.051747f
C769 diffpairibias.t26 gnd 0.08996f
C770 diffpairibias.n24 gnd 0.051736f
C771 diffpairibias.t22 gnd 0.08996f
C772 diffpairibias.n25 gnd 0.051736f
C773 diffpairibias.t21 gnd 0.08996f
C774 diffpairibias.n26 gnd 0.051736f
C775 diffpairibias.t24 gnd 0.08996f
C776 diffpairibias.n27 gnd 0.04729f
C777 diffpairibias.n28 gnd 0.047711f
C778 commonsourceibias.n0 gnd 0.010571f
C779 commonsourceibias.t92 gnd 0.160069f
C780 commonsourceibias.t106 gnd 0.148006f
C781 commonsourceibias.n1 gnd 0.006439f
C782 commonsourceibias.n2 gnd 0.007922f
C783 commonsourceibias.t119 gnd 0.148006f
C784 commonsourceibias.n3 gnd 0.008036f
C785 commonsourceibias.n4 gnd 0.007922f
C786 commonsourceibias.t84 gnd 0.148006f
C787 commonsourceibias.n5 gnd 0.059054f
C788 commonsourceibias.t100 gnd 0.148006f
C789 commonsourceibias.n6 gnd 0.006408f
C790 commonsourceibias.n7 gnd 0.007922f
C791 commonsourceibias.t114 gnd 0.148006f
C792 commonsourceibias.n8 gnd 0.007648f
C793 commonsourceibias.n9 gnd 0.007922f
C794 commonsourceibias.t80 gnd 0.148006f
C795 commonsourceibias.n10 gnd 0.059054f
C796 commonsourceibias.t76 gnd 0.148006f
C797 commonsourceibias.n11 gnd 0.006398f
C798 commonsourceibias.n12 gnd 0.010571f
C799 commonsourceibias.t60 gnd 0.160069f
C800 commonsourceibias.t28 gnd 0.148006f
C801 commonsourceibias.n13 gnd 0.006439f
C802 commonsourceibias.n14 gnd 0.007922f
C803 commonsourceibias.t0 gnd 0.148006f
C804 commonsourceibias.n15 gnd 0.008036f
C805 commonsourceibias.n16 gnd 0.007922f
C806 commonsourceibias.t18 gnd 0.148006f
C807 commonsourceibias.n17 gnd 0.059054f
C808 commonsourceibias.t50 gnd 0.148006f
C809 commonsourceibias.n18 gnd 0.006408f
C810 commonsourceibias.n19 gnd 0.007922f
C811 commonsourceibias.t62 gnd 0.148006f
C812 commonsourceibias.n20 gnd 0.007648f
C813 commonsourceibias.n21 gnd 0.007922f
C814 commonsourceibias.t8 gnd 0.148006f
C815 commonsourceibias.n22 gnd 0.059054f
C816 commonsourceibias.t48 gnd 0.148006f
C817 commonsourceibias.n23 gnd 0.006398f
C818 commonsourceibias.n24 gnd 0.007922f
C819 commonsourceibias.t22 gnd 0.148006f
C820 commonsourceibias.t54 gnd 0.148006f
C821 commonsourceibias.n25 gnd 0.059054f
C822 commonsourceibias.n26 gnd 0.007922f
C823 commonsourceibias.t36 gnd 0.148006f
C824 commonsourceibias.n27 gnd 0.059054f
C825 commonsourceibias.n28 gnd 0.007922f
C826 commonsourceibias.t10 gnd 0.148006f
C827 commonsourceibias.n29 gnd 0.059054f
C828 commonsourceibias.n30 gnd 0.007922f
C829 commonsourceibias.t52 gnd 0.148006f
C830 commonsourceibias.n31 gnd 0.009005f
C831 commonsourceibias.n32 gnd 0.007922f
C832 commonsourceibias.t34 gnd 0.148006f
C833 commonsourceibias.n33 gnd 0.010649f
C834 commonsourceibias.t58 gnd 0.164876f
C835 commonsourceibias.t14 gnd 0.148006f
C836 commonsourceibias.n34 gnd 0.065802f
C837 commonsourceibias.n35 gnd 0.070497f
C838 commonsourceibias.n36 gnd 0.03372f
C839 commonsourceibias.n37 gnd 0.007922f
C840 commonsourceibias.n38 gnd 0.006439f
C841 commonsourceibias.n39 gnd 0.010916f
C842 commonsourceibias.n40 gnd 0.059054f
C843 commonsourceibias.n41 gnd 0.010963f
C844 commonsourceibias.n42 gnd 0.007922f
C845 commonsourceibias.n43 gnd 0.007922f
C846 commonsourceibias.n44 gnd 0.007922f
C847 commonsourceibias.n45 gnd 0.008036f
C848 commonsourceibias.n46 gnd 0.059054f
C849 commonsourceibias.n47 gnd 0.009764f
C850 commonsourceibias.n48 gnd 0.010802f
C851 commonsourceibias.n49 gnd 0.007922f
C852 commonsourceibias.n50 gnd 0.007922f
C853 commonsourceibias.n51 gnd 0.010731f
C854 commonsourceibias.n52 gnd 0.006408f
C855 commonsourceibias.n53 gnd 0.010864f
C856 commonsourceibias.n54 gnd 0.007922f
C857 commonsourceibias.n55 gnd 0.007922f
C858 commonsourceibias.n56 gnd 0.010931f
C859 commonsourceibias.n57 gnd 0.009425f
C860 commonsourceibias.n58 gnd 0.007648f
C861 commonsourceibias.n59 gnd 0.007922f
C862 commonsourceibias.n60 gnd 0.007922f
C863 commonsourceibias.n61 gnd 0.00969f
C864 commonsourceibias.n62 gnd 0.010876f
C865 commonsourceibias.n63 gnd 0.059054f
C866 commonsourceibias.n64 gnd 0.010803f
C867 commonsourceibias.n65 gnd 0.007922f
C868 commonsourceibias.n66 gnd 0.007922f
C869 commonsourceibias.n67 gnd 0.007922f
C870 commonsourceibias.n68 gnd 0.010803f
C871 commonsourceibias.n69 gnd 0.059054f
C872 commonsourceibias.n70 gnd 0.010876f
C873 commonsourceibias.n71 gnd 0.00969f
C874 commonsourceibias.n72 gnd 0.007922f
C875 commonsourceibias.n73 gnd 0.007922f
C876 commonsourceibias.n74 gnd 0.007922f
C877 commonsourceibias.n75 gnd 0.009425f
C878 commonsourceibias.n76 gnd 0.010931f
C879 commonsourceibias.n77 gnd 0.059054f
C880 commonsourceibias.n78 gnd 0.010864f
C881 commonsourceibias.n79 gnd 0.007922f
C882 commonsourceibias.n80 gnd 0.007922f
C883 commonsourceibias.n81 gnd 0.007922f
C884 commonsourceibias.n82 gnd 0.010731f
C885 commonsourceibias.n83 gnd 0.059054f
C886 commonsourceibias.n84 gnd 0.010802f
C887 commonsourceibias.n85 gnd 0.009764f
C888 commonsourceibias.n86 gnd 0.007922f
C889 commonsourceibias.n87 gnd 0.007922f
C890 commonsourceibias.n88 gnd 0.007922f
C891 commonsourceibias.n89 gnd 0.009005f
C892 commonsourceibias.n90 gnd 0.010963f
C893 commonsourceibias.n91 gnd 0.059054f
C894 commonsourceibias.n92 gnd 0.010916f
C895 commonsourceibias.n93 gnd 0.007922f
C896 commonsourceibias.n94 gnd 0.007922f
C897 commonsourceibias.n95 gnd 0.007922f
C898 commonsourceibias.n96 gnd 0.010649f
C899 commonsourceibias.n97 gnd 0.059054f
C900 commonsourceibias.n98 gnd 0.010674f
C901 commonsourceibias.n99 gnd 0.071211f
C902 commonsourceibias.n100 gnd 0.079625f
C903 commonsourceibias.t61 gnd 0.017095f
C904 commonsourceibias.t29 gnd 0.017095f
C905 commonsourceibias.n101 gnd 0.151055f
C906 commonsourceibias.n102 gnd 0.130846f
C907 commonsourceibias.t1 gnd 0.017095f
C908 commonsourceibias.t19 gnd 0.017095f
C909 commonsourceibias.n103 gnd 0.151055f
C910 commonsourceibias.n104 gnd 0.069385f
C911 commonsourceibias.t51 gnd 0.017095f
C912 commonsourceibias.t63 gnd 0.017095f
C913 commonsourceibias.n105 gnd 0.151055f
C914 commonsourceibias.n106 gnd 0.069385f
C915 commonsourceibias.t9 gnd 0.017095f
C916 commonsourceibias.t49 gnd 0.017095f
C917 commonsourceibias.n107 gnd 0.151055f
C918 commonsourceibias.n108 gnd 0.057968f
C919 commonsourceibias.t15 gnd 0.017095f
C920 commonsourceibias.t59 gnd 0.017095f
C921 commonsourceibias.n109 gnd 0.15156f
C922 commonsourceibias.t53 gnd 0.017095f
C923 commonsourceibias.t35 gnd 0.017095f
C924 commonsourceibias.n110 gnd 0.151055f
C925 commonsourceibias.n111 gnd 0.140755f
C926 commonsourceibias.t37 gnd 0.017095f
C927 commonsourceibias.t11 gnd 0.017095f
C928 commonsourceibias.n112 gnd 0.151055f
C929 commonsourceibias.n113 gnd 0.069385f
C930 commonsourceibias.t23 gnd 0.017095f
C931 commonsourceibias.t55 gnd 0.017095f
C932 commonsourceibias.n114 gnd 0.151055f
C933 commonsourceibias.n115 gnd 0.057968f
C934 commonsourceibias.n116 gnd 0.070193f
C935 commonsourceibias.n117 gnd 0.007922f
C936 commonsourceibias.t105 gnd 0.148006f
C937 commonsourceibias.t121 gnd 0.148006f
C938 commonsourceibias.n118 gnd 0.059054f
C939 commonsourceibias.n119 gnd 0.007922f
C940 commonsourceibias.t71 gnd 0.148006f
C941 commonsourceibias.n120 gnd 0.059054f
C942 commonsourceibias.n121 gnd 0.007922f
C943 commonsourceibias.t99 gnd 0.148006f
C944 commonsourceibias.n122 gnd 0.059054f
C945 commonsourceibias.n123 gnd 0.007922f
C946 commonsourceibias.t95 gnd 0.148006f
C947 commonsourceibias.n124 gnd 0.009005f
C948 commonsourceibias.n125 gnd 0.007922f
C949 commonsourceibias.t109 gnd 0.148006f
C950 commonsourceibias.n126 gnd 0.010649f
C951 commonsourceibias.t85 gnd 0.164876f
C952 commonsourceibias.t89 gnd 0.148006f
C953 commonsourceibias.n127 gnd 0.065802f
C954 commonsourceibias.n128 gnd 0.070497f
C955 commonsourceibias.n129 gnd 0.03372f
C956 commonsourceibias.n130 gnd 0.007922f
C957 commonsourceibias.n131 gnd 0.006439f
C958 commonsourceibias.n132 gnd 0.010916f
C959 commonsourceibias.n133 gnd 0.059054f
C960 commonsourceibias.n134 gnd 0.010963f
C961 commonsourceibias.n135 gnd 0.007922f
C962 commonsourceibias.n136 gnd 0.007922f
C963 commonsourceibias.n137 gnd 0.007922f
C964 commonsourceibias.n138 gnd 0.008036f
C965 commonsourceibias.n139 gnd 0.059054f
C966 commonsourceibias.n140 gnd 0.009764f
C967 commonsourceibias.n141 gnd 0.010802f
C968 commonsourceibias.n142 gnd 0.007922f
C969 commonsourceibias.n143 gnd 0.007922f
C970 commonsourceibias.n144 gnd 0.010731f
C971 commonsourceibias.n145 gnd 0.006408f
C972 commonsourceibias.n146 gnd 0.010864f
C973 commonsourceibias.n147 gnd 0.007922f
C974 commonsourceibias.n148 gnd 0.007922f
C975 commonsourceibias.n149 gnd 0.010931f
C976 commonsourceibias.n150 gnd 0.009425f
C977 commonsourceibias.n151 gnd 0.007648f
C978 commonsourceibias.n152 gnd 0.007922f
C979 commonsourceibias.n153 gnd 0.007922f
C980 commonsourceibias.n154 gnd 0.00969f
C981 commonsourceibias.n155 gnd 0.010876f
C982 commonsourceibias.n156 gnd 0.059054f
C983 commonsourceibias.n157 gnd 0.010803f
C984 commonsourceibias.n158 gnd 0.007884f
C985 commonsourceibias.n159 gnd 0.057266f
C986 commonsourceibias.n160 gnd 0.007884f
C987 commonsourceibias.n161 gnd 0.010803f
C988 commonsourceibias.n162 gnd 0.059054f
C989 commonsourceibias.n163 gnd 0.010876f
C990 commonsourceibias.n164 gnd 0.00969f
C991 commonsourceibias.n165 gnd 0.007922f
C992 commonsourceibias.n166 gnd 0.007922f
C993 commonsourceibias.n167 gnd 0.007922f
C994 commonsourceibias.n168 gnd 0.009425f
C995 commonsourceibias.n169 gnd 0.010931f
C996 commonsourceibias.n170 gnd 0.059054f
C997 commonsourceibias.n171 gnd 0.010864f
C998 commonsourceibias.n172 gnd 0.007922f
C999 commonsourceibias.n173 gnd 0.007922f
C1000 commonsourceibias.n174 gnd 0.007922f
C1001 commonsourceibias.n175 gnd 0.010731f
C1002 commonsourceibias.n176 gnd 0.059054f
C1003 commonsourceibias.n177 gnd 0.010802f
C1004 commonsourceibias.n178 gnd 0.009764f
C1005 commonsourceibias.n179 gnd 0.007922f
C1006 commonsourceibias.n180 gnd 0.007922f
C1007 commonsourceibias.n181 gnd 0.007922f
C1008 commonsourceibias.n182 gnd 0.009005f
C1009 commonsourceibias.n183 gnd 0.010963f
C1010 commonsourceibias.n184 gnd 0.059054f
C1011 commonsourceibias.n185 gnd 0.010916f
C1012 commonsourceibias.n186 gnd 0.007922f
C1013 commonsourceibias.n187 gnd 0.007922f
C1014 commonsourceibias.n188 gnd 0.007922f
C1015 commonsourceibias.n189 gnd 0.010649f
C1016 commonsourceibias.n190 gnd 0.059054f
C1017 commonsourceibias.n191 gnd 0.010674f
C1018 commonsourceibias.n192 gnd 0.071211f
C1019 commonsourceibias.n193 gnd 0.047027f
C1020 commonsourceibias.n194 gnd 0.010571f
C1021 commonsourceibias.t94 gnd 0.148006f
C1022 commonsourceibias.n195 gnd 0.006439f
C1023 commonsourceibias.n196 gnd 0.007922f
C1024 commonsourceibias.t107 gnd 0.148006f
C1025 commonsourceibias.n197 gnd 0.008036f
C1026 commonsourceibias.n198 gnd 0.007922f
C1027 commonsourceibias.t74 gnd 0.148006f
C1028 commonsourceibias.n199 gnd 0.059054f
C1029 commonsourceibias.t87 gnd 0.148006f
C1030 commonsourceibias.n200 gnd 0.006408f
C1031 commonsourceibias.n201 gnd 0.007922f
C1032 commonsourceibias.t101 gnd 0.148006f
C1033 commonsourceibias.n202 gnd 0.007648f
C1034 commonsourceibias.n203 gnd 0.007922f
C1035 commonsourceibias.t70 gnd 0.148006f
C1036 commonsourceibias.n204 gnd 0.059054f
C1037 commonsourceibias.t67 gnd 0.148006f
C1038 commonsourceibias.n205 gnd 0.006398f
C1039 commonsourceibias.n206 gnd 0.007922f
C1040 commonsourceibias.t93 gnd 0.148006f
C1041 commonsourceibias.t108 gnd 0.148006f
C1042 commonsourceibias.n207 gnd 0.059054f
C1043 commonsourceibias.n208 gnd 0.007922f
C1044 commonsourceibias.t127 gnd 0.148006f
C1045 commonsourceibias.n209 gnd 0.059054f
C1046 commonsourceibias.n210 gnd 0.007922f
C1047 commonsourceibias.t86 gnd 0.148006f
C1048 commonsourceibias.n211 gnd 0.059054f
C1049 commonsourceibias.n212 gnd 0.007922f
C1050 commonsourceibias.t82 gnd 0.148006f
C1051 commonsourceibias.n213 gnd 0.009005f
C1052 commonsourceibias.n214 gnd 0.007922f
C1053 commonsourceibias.t96 gnd 0.148006f
C1054 commonsourceibias.n215 gnd 0.010649f
C1055 commonsourceibias.t75 gnd 0.164876f
C1056 commonsourceibias.t77 gnd 0.148006f
C1057 commonsourceibias.n216 gnd 0.065802f
C1058 commonsourceibias.n217 gnd 0.070497f
C1059 commonsourceibias.n218 gnd 0.03372f
C1060 commonsourceibias.n219 gnd 0.007922f
C1061 commonsourceibias.n220 gnd 0.006439f
C1062 commonsourceibias.n221 gnd 0.010916f
C1063 commonsourceibias.n222 gnd 0.059054f
C1064 commonsourceibias.n223 gnd 0.010963f
C1065 commonsourceibias.n224 gnd 0.007922f
C1066 commonsourceibias.n225 gnd 0.007922f
C1067 commonsourceibias.n226 gnd 0.007922f
C1068 commonsourceibias.n227 gnd 0.008036f
C1069 commonsourceibias.n228 gnd 0.059054f
C1070 commonsourceibias.n229 gnd 0.009764f
C1071 commonsourceibias.n230 gnd 0.010802f
C1072 commonsourceibias.n231 gnd 0.007922f
C1073 commonsourceibias.n232 gnd 0.007922f
C1074 commonsourceibias.n233 gnd 0.010731f
C1075 commonsourceibias.n234 gnd 0.006408f
C1076 commonsourceibias.n235 gnd 0.010864f
C1077 commonsourceibias.n236 gnd 0.007922f
C1078 commonsourceibias.n237 gnd 0.007922f
C1079 commonsourceibias.n238 gnd 0.010931f
C1080 commonsourceibias.n239 gnd 0.009425f
C1081 commonsourceibias.n240 gnd 0.007648f
C1082 commonsourceibias.n241 gnd 0.007922f
C1083 commonsourceibias.n242 gnd 0.007922f
C1084 commonsourceibias.n243 gnd 0.00969f
C1085 commonsourceibias.n244 gnd 0.010876f
C1086 commonsourceibias.n245 gnd 0.059054f
C1087 commonsourceibias.n246 gnd 0.010803f
C1088 commonsourceibias.n247 gnd 0.007922f
C1089 commonsourceibias.n248 gnd 0.007922f
C1090 commonsourceibias.n249 gnd 0.007922f
C1091 commonsourceibias.n250 gnd 0.010803f
C1092 commonsourceibias.n251 gnd 0.059054f
C1093 commonsourceibias.n252 gnd 0.010876f
C1094 commonsourceibias.n253 gnd 0.00969f
C1095 commonsourceibias.n254 gnd 0.007922f
C1096 commonsourceibias.n255 gnd 0.007922f
C1097 commonsourceibias.n256 gnd 0.007922f
C1098 commonsourceibias.n257 gnd 0.009425f
C1099 commonsourceibias.n258 gnd 0.010931f
C1100 commonsourceibias.n259 gnd 0.059054f
C1101 commonsourceibias.n260 gnd 0.010864f
C1102 commonsourceibias.n261 gnd 0.007922f
C1103 commonsourceibias.n262 gnd 0.007922f
C1104 commonsourceibias.n263 gnd 0.007922f
C1105 commonsourceibias.n264 gnd 0.010731f
C1106 commonsourceibias.n265 gnd 0.059054f
C1107 commonsourceibias.n266 gnd 0.010802f
C1108 commonsourceibias.n267 gnd 0.009764f
C1109 commonsourceibias.n268 gnd 0.007922f
C1110 commonsourceibias.n269 gnd 0.007922f
C1111 commonsourceibias.n270 gnd 0.007922f
C1112 commonsourceibias.n271 gnd 0.009005f
C1113 commonsourceibias.n272 gnd 0.010963f
C1114 commonsourceibias.n273 gnd 0.059054f
C1115 commonsourceibias.n274 gnd 0.010916f
C1116 commonsourceibias.n275 gnd 0.007922f
C1117 commonsourceibias.n276 gnd 0.007922f
C1118 commonsourceibias.n277 gnd 0.007922f
C1119 commonsourceibias.n278 gnd 0.010649f
C1120 commonsourceibias.n279 gnd 0.059054f
C1121 commonsourceibias.n280 gnd 0.010674f
C1122 commonsourceibias.t81 gnd 0.160069f
C1123 commonsourceibias.n281 gnd 0.071211f
C1124 commonsourceibias.n282 gnd 0.025411f
C1125 commonsourceibias.n283 gnd 0.458519f
C1126 commonsourceibias.n284 gnd 0.010571f
C1127 commonsourceibias.t110 gnd 0.160069f
C1128 commonsourceibias.t123 gnd 0.148006f
C1129 commonsourceibias.n285 gnd 0.006439f
C1130 commonsourceibias.n286 gnd 0.007922f
C1131 commonsourceibias.t68 gnd 0.148006f
C1132 commonsourceibias.n287 gnd 0.008036f
C1133 commonsourceibias.n288 gnd 0.007922f
C1134 commonsourceibias.t117 gnd 0.148006f
C1135 commonsourceibias.n289 gnd 0.006408f
C1136 commonsourceibias.n290 gnd 0.007922f
C1137 commonsourceibias.t64 gnd 0.148006f
C1138 commonsourceibias.n291 gnd 0.007648f
C1139 commonsourceibias.n292 gnd 0.007922f
C1140 commonsourceibias.t90 gnd 0.148006f
C1141 commonsourceibias.n293 gnd 0.006398f
C1142 commonsourceibias.n294 gnd 0.007922f
C1143 commonsourceibias.t122 gnd 0.148006f
C1144 commonsourceibias.t69 gnd 0.148006f
C1145 commonsourceibias.n295 gnd 0.059054f
C1146 commonsourceibias.n296 gnd 0.007922f
C1147 commonsourceibias.t66 gnd 0.148006f
C1148 commonsourceibias.n297 gnd 0.059054f
C1149 commonsourceibias.n298 gnd 0.007922f
C1150 commonsourceibias.t116 gnd 0.148006f
C1151 commonsourceibias.n299 gnd 0.059054f
C1152 commonsourceibias.n300 gnd 0.007922f
C1153 commonsourceibias.t113 gnd 0.148006f
C1154 commonsourceibias.n301 gnd 0.009005f
C1155 commonsourceibias.n302 gnd 0.007922f
C1156 commonsourceibias.t126 gnd 0.148006f
C1157 commonsourceibias.n303 gnd 0.010649f
C1158 commonsourceibias.t91 gnd 0.164876f
C1159 commonsourceibias.t83 gnd 0.148006f
C1160 commonsourceibias.n304 gnd 0.065802f
C1161 commonsourceibias.n305 gnd 0.070497f
C1162 commonsourceibias.n306 gnd 0.03372f
C1163 commonsourceibias.n307 gnd 0.007922f
C1164 commonsourceibias.n308 gnd 0.006439f
C1165 commonsourceibias.n309 gnd 0.010916f
C1166 commonsourceibias.n310 gnd 0.059054f
C1167 commonsourceibias.n311 gnd 0.010963f
C1168 commonsourceibias.n312 gnd 0.007922f
C1169 commonsourceibias.n313 gnd 0.007922f
C1170 commonsourceibias.n314 gnd 0.007922f
C1171 commonsourceibias.n315 gnd 0.008036f
C1172 commonsourceibias.n316 gnd 0.059054f
C1173 commonsourceibias.n317 gnd 0.009764f
C1174 commonsourceibias.n318 gnd 0.010802f
C1175 commonsourceibias.n319 gnd 0.007922f
C1176 commonsourceibias.n320 gnd 0.007922f
C1177 commonsourceibias.n321 gnd 0.010731f
C1178 commonsourceibias.n322 gnd 0.006408f
C1179 commonsourceibias.n323 gnd 0.010864f
C1180 commonsourceibias.n324 gnd 0.007922f
C1181 commonsourceibias.n325 gnd 0.007922f
C1182 commonsourceibias.n326 gnd 0.010931f
C1183 commonsourceibias.n327 gnd 0.009425f
C1184 commonsourceibias.n328 gnd 0.007648f
C1185 commonsourceibias.n329 gnd 0.007922f
C1186 commonsourceibias.n330 gnd 0.007922f
C1187 commonsourceibias.n331 gnd 0.00969f
C1188 commonsourceibias.n332 gnd 0.010876f
C1189 commonsourceibias.n333 gnd 0.059054f
C1190 commonsourceibias.n334 gnd 0.010803f
C1191 commonsourceibias.n335 gnd 0.007884f
C1192 commonsourceibias.t31 gnd 0.017095f
C1193 commonsourceibias.t47 gnd 0.017095f
C1194 commonsourceibias.n336 gnd 0.15156f
C1195 commonsourceibias.t25 gnd 0.017095f
C1196 commonsourceibias.t43 gnd 0.017095f
C1197 commonsourceibias.n337 gnd 0.151055f
C1198 commonsourceibias.n338 gnd 0.140755f
C1199 commonsourceibias.t3 gnd 0.017095f
C1200 commonsourceibias.t33 gnd 0.017095f
C1201 commonsourceibias.n339 gnd 0.151055f
C1202 commonsourceibias.n340 gnd 0.069385f
C1203 commonsourceibias.t45 gnd 0.017095f
C1204 commonsourceibias.t7 gnd 0.017095f
C1205 commonsourceibias.n341 gnd 0.151055f
C1206 commonsourceibias.n342 gnd 0.057968f
C1207 commonsourceibias.n343 gnd 0.010571f
C1208 commonsourceibias.t56 gnd 0.148006f
C1209 commonsourceibias.n344 gnd 0.006439f
C1210 commonsourceibias.n345 gnd 0.007922f
C1211 commonsourceibias.t26 gnd 0.148006f
C1212 commonsourceibias.n346 gnd 0.008036f
C1213 commonsourceibias.n347 gnd 0.007922f
C1214 commonsourceibias.t40 gnd 0.148006f
C1215 commonsourceibias.n348 gnd 0.006408f
C1216 commonsourceibias.n349 gnd 0.007922f
C1217 commonsourceibias.t16 gnd 0.148006f
C1218 commonsourceibias.n350 gnd 0.007648f
C1219 commonsourceibias.n351 gnd 0.007922f
C1220 commonsourceibias.t38 gnd 0.148006f
C1221 commonsourceibias.n352 gnd 0.006398f
C1222 commonsourceibias.n353 gnd 0.007922f
C1223 commonsourceibias.t6 gnd 0.148006f
C1224 commonsourceibias.t44 gnd 0.148006f
C1225 commonsourceibias.n354 gnd 0.059054f
C1226 commonsourceibias.n355 gnd 0.007922f
C1227 commonsourceibias.t32 gnd 0.148006f
C1228 commonsourceibias.n356 gnd 0.059054f
C1229 commonsourceibias.n357 gnd 0.007922f
C1230 commonsourceibias.t2 gnd 0.148006f
C1231 commonsourceibias.n358 gnd 0.059054f
C1232 commonsourceibias.n359 gnd 0.007922f
C1233 commonsourceibias.t42 gnd 0.148006f
C1234 commonsourceibias.n360 gnd 0.009005f
C1235 commonsourceibias.n361 gnd 0.007922f
C1236 commonsourceibias.t24 gnd 0.148006f
C1237 commonsourceibias.n362 gnd 0.010649f
C1238 commonsourceibias.t30 gnd 0.164876f
C1239 commonsourceibias.t46 gnd 0.148006f
C1240 commonsourceibias.n363 gnd 0.065802f
C1241 commonsourceibias.n364 gnd 0.070497f
C1242 commonsourceibias.n365 gnd 0.03372f
C1243 commonsourceibias.n366 gnd 0.007922f
C1244 commonsourceibias.n367 gnd 0.006439f
C1245 commonsourceibias.n368 gnd 0.010916f
C1246 commonsourceibias.n369 gnd 0.059054f
C1247 commonsourceibias.n370 gnd 0.010963f
C1248 commonsourceibias.n371 gnd 0.007922f
C1249 commonsourceibias.n372 gnd 0.007922f
C1250 commonsourceibias.n373 gnd 0.007922f
C1251 commonsourceibias.n374 gnd 0.008036f
C1252 commonsourceibias.n375 gnd 0.059054f
C1253 commonsourceibias.n376 gnd 0.009764f
C1254 commonsourceibias.n377 gnd 0.010802f
C1255 commonsourceibias.n378 gnd 0.007922f
C1256 commonsourceibias.n379 gnd 0.007922f
C1257 commonsourceibias.n380 gnd 0.010731f
C1258 commonsourceibias.n381 gnd 0.006408f
C1259 commonsourceibias.n382 gnd 0.010864f
C1260 commonsourceibias.n383 gnd 0.007922f
C1261 commonsourceibias.n384 gnd 0.007922f
C1262 commonsourceibias.n385 gnd 0.010931f
C1263 commonsourceibias.n386 gnd 0.009425f
C1264 commonsourceibias.n387 gnd 0.007648f
C1265 commonsourceibias.n388 gnd 0.007922f
C1266 commonsourceibias.n389 gnd 0.007922f
C1267 commonsourceibias.n390 gnd 0.00969f
C1268 commonsourceibias.n391 gnd 0.010876f
C1269 commonsourceibias.n392 gnd 0.059054f
C1270 commonsourceibias.n393 gnd 0.010803f
C1271 commonsourceibias.n394 gnd 0.007922f
C1272 commonsourceibias.n395 gnd 0.007922f
C1273 commonsourceibias.n396 gnd 0.007922f
C1274 commonsourceibias.n397 gnd 0.010803f
C1275 commonsourceibias.n398 gnd 0.059054f
C1276 commonsourceibias.n399 gnd 0.010876f
C1277 commonsourceibias.t4 gnd 0.148006f
C1278 commonsourceibias.n400 gnd 0.059054f
C1279 commonsourceibias.n401 gnd 0.00969f
C1280 commonsourceibias.n402 gnd 0.007922f
C1281 commonsourceibias.n403 gnd 0.007922f
C1282 commonsourceibias.n404 gnd 0.007922f
C1283 commonsourceibias.n405 gnd 0.009425f
C1284 commonsourceibias.n406 gnd 0.010931f
C1285 commonsourceibias.n407 gnd 0.059054f
C1286 commonsourceibias.n408 gnd 0.010864f
C1287 commonsourceibias.n409 gnd 0.007922f
C1288 commonsourceibias.n410 gnd 0.007922f
C1289 commonsourceibias.n411 gnd 0.007922f
C1290 commonsourceibias.n412 gnd 0.010731f
C1291 commonsourceibias.n413 gnd 0.059054f
C1292 commonsourceibias.n414 gnd 0.010802f
C1293 commonsourceibias.t12 gnd 0.148006f
C1294 commonsourceibias.n415 gnd 0.059054f
C1295 commonsourceibias.n416 gnd 0.009764f
C1296 commonsourceibias.n417 gnd 0.007922f
C1297 commonsourceibias.n418 gnd 0.007922f
C1298 commonsourceibias.n419 gnd 0.007922f
C1299 commonsourceibias.n420 gnd 0.009005f
C1300 commonsourceibias.n421 gnd 0.010963f
C1301 commonsourceibias.n422 gnd 0.059054f
C1302 commonsourceibias.n423 gnd 0.010916f
C1303 commonsourceibias.n424 gnd 0.007922f
C1304 commonsourceibias.n425 gnd 0.007922f
C1305 commonsourceibias.n426 gnd 0.007922f
C1306 commonsourceibias.n427 gnd 0.010649f
C1307 commonsourceibias.n428 gnd 0.059054f
C1308 commonsourceibias.n429 gnd 0.010674f
C1309 commonsourceibias.t20 gnd 0.160069f
C1310 commonsourceibias.n430 gnd 0.071211f
C1311 commonsourceibias.n431 gnd 0.079625f
C1312 commonsourceibias.t57 gnd 0.017095f
C1313 commonsourceibias.t21 gnd 0.017095f
C1314 commonsourceibias.n432 gnd 0.151055f
C1315 commonsourceibias.n433 gnd 0.130846f
C1316 commonsourceibias.t13 gnd 0.017095f
C1317 commonsourceibias.t27 gnd 0.017095f
C1318 commonsourceibias.n434 gnd 0.151055f
C1319 commonsourceibias.n435 gnd 0.069385f
C1320 commonsourceibias.t17 gnd 0.017095f
C1321 commonsourceibias.t41 gnd 0.017095f
C1322 commonsourceibias.n436 gnd 0.151055f
C1323 commonsourceibias.n437 gnd 0.069385f
C1324 commonsourceibias.t39 gnd 0.017095f
C1325 commonsourceibias.t5 gnd 0.017095f
C1326 commonsourceibias.n438 gnd 0.151055f
C1327 commonsourceibias.n439 gnd 0.057968f
C1328 commonsourceibias.n440 gnd 0.070193f
C1329 commonsourceibias.n441 gnd 0.057266f
C1330 commonsourceibias.n442 gnd 0.007884f
C1331 commonsourceibias.n443 gnd 0.010803f
C1332 commonsourceibias.n444 gnd 0.059054f
C1333 commonsourceibias.n445 gnd 0.010876f
C1334 commonsourceibias.t72 gnd 0.148006f
C1335 commonsourceibias.n446 gnd 0.059054f
C1336 commonsourceibias.n447 gnd 0.00969f
C1337 commonsourceibias.n448 gnd 0.007922f
C1338 commonsourceibias.n449 gnd 0.007922f
C1339 commonsourceibias.n450 gnd 0.007922f
C1340 commonsourceibias.n451 gnd 0.009425f
C1341 commonsourceibias.n452 gnd 0.010931f
C1342 commonsourceibias.n453 gnd 0.059054f
C1343 commonsourceibias.n454 gnd 0.010864f
C1344 commonsourceibias.n455 gnd 0.007922f
C1345 commonsourceibias.n456 gnd 0.007922f
C1346 commonsourceibias.n457 gnd 0.007922f
C1347 commonsourceibias.n458 gnd 0.010731f
C1348 commonsourceibias.n459 gnd 0.059054f
C1349 commonsourceibias.n460 gnd 0.010802f
C1350 commonsourceibias.t102 gnd 0.148006f
C1351 commonsourceibias.n461 gnd 0.059054f
C1352 commonsourceibias.n462 gnd 0.009764f
C1353 commonsourceibias.n463 gnd 0.007922f
C1354 commonsourceibias.n464 gnd 0.007922f
C1355 commonsourceibias.n465 gnd 0.007922f
C1356 commonsourceibias.n466 gnd 0.009005f
C1357 commonsourceibias.n467 gnd 0.010963f
C1358 commonsourceibias.n468 gnd 0.059054f
C1359 commonsourceibias.n469 gnd 0.010916f
C1360 commonsourceibias.n470 gnd 0.007922f
C1361 commonsourceibias.n471 gnd 0.007922f
C1362 commonsourceibias.n472 gnd 0.007922f
C1363 commonsourceibias.n473 gnd 0.010649f
C1364 commonsourceibias.n474 gnd 0.059054f
C1365 commonsourceibias.n475 gnd 0.010674f
C1366 commonsourceibias.n476 gnd 0.071211f
C1367 commonsourceibias.n477 gnd 0.047027f
C1368 commonsourceibias.n478 gnd 0.010571f
C1369 commonsourceibias.t112 gnd 0.148006f
C1370 commonsourceibias.n479 gnd 0.006439f
C1371 commonsourceibias.n480 gnd 0.007922f
C1372 commonsourceibias.t124 gnd 0.148006f
C1373 commonsourceibias.n481 gnd 0.008036f
C1374 commonsourceibias.n482 gnd 0.007922f
C1375 commonsourceibias.t104 gnd 0.148006f
C1376 commonsourceibias.n483 gnd 0.006408f
C1377 commonsourceibias.n484 gnd 0.007922f
C1378 commonsourceibias.t118 gnd 0.148006f
C1379 commonsourceibias.n485 gnd 0.007648f
C1380 commonsourceibias.n486 gnd 0.007922f
C1381 commonsourceibias.t79 gnd 0.148006f
C1382 commonsourceibias.n487 gnd 0.006398f
C1383 commonsourceibias.n488 gnd 0.007922f
C1384 commonsourceibias.t111 gnd 0.148006f
C1385 commonsourceibias.t125 gnd 0.148006f
C1386 commonsourceibias.n489 gnd 0.059054f
C1387 commonsourceibias.n490 gnd 0.007922f
C1388 commonsourceibias.t120 gnd 0.148006f
C1389 commonsourceibias.n491 gnd 0.059054f
C1390 commonsourceibias.n492 gnd 0.007922f
C1391 commonsourceibias.t103 gnd 0.148006f
C1392 commonsourceibias.n493 gnd 0.059054f
C1393 commonsourceibias.n494 gnd 0.007922f
C1394 commonsourceibias.t98 gnd 0.148006f
C1395 commonsourceibias.n495 gnd 0.009005f
C1396 commonsourceibias.n496 gnd 0.007922f
C1397 commonsourceibias.t115 gnd 0.148006f
C1398 commonsourceibias.n497 gnd 0.010649f
C1399 commonsourceibias.t78 gnd 0.164876f
C1400 commonsourceibias.t73 gnd 0.148006f
C1401 commonsourceibias.n498 gnd 0.065802f
C1402 commonsourceibias.n499 gnd 0.070497f
C1403 commonsourceibias.n500 gnd 0.03372f
C1404 commonsourceibias.n501 gnd 0.007922f
C1405 commonsourceibias.n502 gnd 0.006439f
C1406 commonsourceibias.n503 gnd 0.010916f
C1407 commonsourceibias.n504 gnd 0.059054f
C1408 commonsourceibias.n505 gnd 0.010963f
C1409 commonsourceibias.n506 gnd 0.007922f
C1410 commonsourceibias.n507 gnd 0.007922f
C1411 commonsourceibias.n508 gnd 0.007922f
C1412 commonsourceibias.n509 gnd 0.008036f
C1413 commonsourceibias.n510 gnd 0.059054f
C1414 commonsourceibias.n511 gnd 0.009764f
C1415 commonsourceibias.n512 gnd 0.010802f
C1416 commonsourceibias.n513 gnd 0.007922f
C1417 commonsourceibias.n514 gnd 0.007922f
C1418 commonsourceibias.n515 gnd 0.010731f
C1419 commonsourceibias.n516 gnd 0.006408f
C1420 commonsourceibias.n517 gnd 0.010864f
C1421 commonsourceibias.n518 gnd 0.007922f
C1422 commonsourceibias.n519 gnd 0.007922f
C1423 commonsourceibias.n520 gnd 0.010931f
C1424 commonsourceibias.n521 gnd 0.009425f
C1425 commonsourceibias.n522 gnd 0.007648f
C1426 commonsourceibias.n523 gnd 0.007922f
C1427 commonsourceibias.n524 gnd 0.007922f
C1428 commonsourceibias.n525 gnd 0.00969f
C1429 commonsourceibias.n526 gnd 0.010876f
C1430 commonsourceibias.n527 gnd 0.059054f
C1431 commonsourceibias.n528 gnd 0.010803f
C1432 commonsourceibias.n529 gnd 0.007922f
C1433 commonsourceibias.n530 gnd 0.007922f
C1434 commonsourceibias.n531 gnd 0.007922f
C1435 commonsourceibias.n532 gnd 0.010803f
C1436 commonsourceibias.n533 gnd 0.059054f
C1437 commonsourceibias.n534 gnd 0.010876f
C1438 commonsourceibias.t65 gnd 0.148006f
C1439 commonsourceibias.n535 gnd 0.059054f
C1440 commonsourceibias.n536 gnd 0.00969f
C1441 commonsourceibias.n537 gnd 0.007922f
C1442 commonsourceibias.n538 gnd 0.007922f
C1443 commonsourceibias.n539 gnd 0.007922f
C1444 commonsourceibias.n540 gnd 0.009425f
C1445 commonsourceibias.n541 gnd 0.010931f
C1446 commonsourceibias.n542 gnd 0.059054f
C1447 commonsourceibias.n543 gnd 0.010864f
C1448 commonsourceibias.n544 gnd 0.007922f
C1449 commonsourceibias.n545 gnd 0.007922f
C1450 commonsourceibias.n546 gnd 0.007922f
C1451 commonsourceibias.n547 gnd 0.010731f
C1452 commonsourceibias.n548 gnd 0.059054f
C1453 commonsourceibias.n549 gnd 0.010802f
C1454 commonsourceibias.t88 gnd 0.148006f
C1455 commonsourceibias.n550 gnd 0.059054f
C1456 commonsourceibias.n551 gnd 0.009764f
C1457 commonsourceibias.n552 gnd 0.007922f
C1458 commonsourceibias.n553 gnd 0.007922f
C1459 commonsourceibias.n554 gnd 0.007922f
C1460 commonsourceibias.n555 gnd 0.009005f
C1461 commonsourceibias.n556 gnd 0.010963f
C1462 commonsourceibias.n557 gnd 0.059054f
C1463 commonsourceibias.n558 gnd 0.010916f
C1464 commonsourceibias.n559 gnd 0.007922f
C1465 commonsourceibias.n560 gnd 0.007922f
C1466 commonsourceibias.n561 gnd 0.007922f
C1467 commonsourceibias.n562 gnd 0.010649f
C1468 commonsourceibias.n563 gnd 0.059054f
C1469 commonsourceibias.n564 gnd 0.010674f
C1470 commonsourceibias.t97 gnd 0.160069f
C1471 commonsourceibias.n565 gnd 0.071211f
C1472 commonsourceibias.n566 gnd 0.025411f
C1473 commonsourceibias.n567 gnd 0.219034f
C1474 commonsourceibias.n568 gnd 4.63083f
C1475 a_n2472_13878.t13 gnd 0.187752f
C1476 a_n2472_13878.t15 gnd 0.187752f
C1477 a_n2472_13878.t7 gnd 0.187752f
C1478 a_n2472_13878.n0 gnd 1.47995f
C1479 a_n2472_13878.t12 gnd 0.187752f
C1480 a_n2472_13878.t6 gnd 0.187752f
C1481 a_n2472_13878.n1 gnd 1.47838f
C1482 a_n2472_13878.n2 gnd 2.06575f
C1483 a_n2472_13878.t2 gnd 0.187752f
C1484 a_n2472_13878.t4 gnd 0.187752f
C1485 a_n2472_13878.n3 gnd 1.47838f
C1486 a_n2472_13878.n4 gnd 1.00763f
C1487 a_n2472_13878.t14 gnd 0.187752f
C1488 a_n2472_13878.t3 gnd 0.187752f
C1489 a_n2472_13878.n5 gnd 1.47838f
C1490 a_n2472_13878.n6 gnd 1.00763f
C1491 a_n2472_13878.t11 gnd 0.187752f
C1492 a_n2472_13878.t1 gnd 0.187752f
C1493 a_n2472_13878.n7 gnd 1.47838f
C1494 a_n2472_13878.n8 gnd 4.40971f
C1495 a_n2472_13878.t21 gnd 1.75801f
C1496 a_n2472_13878.t24 gnd 0.187752f
C1497 a_n2472_13878.t25 gnd 0.187752f
C1498 a_n2472_13878.n9 gnd 1.32252f
C1499 a_n2472_13878.n10 gnd 1.47772f
C1500 a_n2472_13878.t20 gnd 1.75451f
C1501 a_n2472_13878.n11 gnd 0.743612f
C1502 a_n2472_13878.t23 gnd 1.75451f
C1503 a_n2472_13878.n12 gnd 0.743612f
C1504 a_n2472_13878.t26 gnd 0.187752f
C1505 a_n2472_13878.t27 gnd 0.187752f
C1506 a_n2472_13878.n13 gnd 1.32252f
C1507 a_n2472_13878.n14 gnd 0.750813f
C1508 a_n2472_13878.t22 gnd 1.75451f
C1509 a_n2472_13878.n15 gnd 2.43968f
C1510 a_n2472_13878.n16 gnd 3.23176f
C1511 a_n2472_13878.t16 gnd 0.187752f
C1512 a_n2472_13878.t5 gnd 0.187752f
C1513 a_n2472_13878.n17 gnd 1.47838f
C1514 a_n2472_13878.n18 gnd 2.22265f
C1515 a_n2472_13878.t8 gnd 0.187752f
C1516 a_n2472_13878.t9 gnd 0.187752f
C1517 a_n2472_13878.n19 gnd 1.47838f
C1518 a_n2472_13878.n20 gnd 0.655033f
C1519 a_n2472_13878.t17 gnd 0.187752f
C1520 a_n2472_13878.t18 gnd 0.187752f
C1521 a_n2472_13878.n21 gnd 1.47838f
C1522 a_n2472_13878.n22 gnd 0.655033f
C1523 a_n2472_13878.t0 gnd 0.187752f
C1524 a_n2472_13878.t10 gnd 0.187752f
C1525 a_n2472_13878.n23 gnd 1.47838f
C1526 a_n2472_13878.n24 gnd 1.32888f
C1527 a_n2472_13878.n25 gnd 1.48083f
C1528 a_n2472_13878.t19 gnd 0.187752f
C1529 a_n2650_13878.n0 gnd 0.21772f
C1530 a_n2650_13878.n1 gnd 0.21772f
C1531 a_n2650_13878.n2 gnd 0.809668f
C1532 a_n2650_13878.n3 gnd 0.21772f
C1533 a_n2650_13878.n4 gnd 0.942749f
C1534 a_n2650_13878.n5 gnd 0.21772f
C1535 a_n2650_13878.n6 gnd 0.506761f
C1536 a_n2650_13878.n7 gnd 0.809584f
C1537 a_n2650_13878.n8 gnd 0.20658f
C1538 a_n2650_13878.n9 gnd 0.15215f
C1539 a_n2650_13878.n10 gnd 0.239132f
C1540 a_n2650_13878.n11 gnd 0.184702f
C1541 a_n2650_13878.n12 gnd 0.20658f
C1542 a_n2650_13878.n13 gnd 1.25084f
C1543 a_n2650_13878.n14 gnd 0.15215f
C1544 a_n2650_13878.n15 gnd 0.864014f
C1545 a_n2650_13878.n16 gnd 0.21772f
C1546 a_n2650_13878.n17 gnd 0.702566f
C1547 a_n2650_13878.n18 gnd 0.21772f
C1548 a_n2650_13878.n19 gnd 0.507263f
C1549 a_n2650_13878.n20 gnd 0.21772f
C1550 a_n2650_13878.n21 gnd 0.561693f
C1551 a_n2650_13878.n22 gnd 0.21772f
C1552 a_n2650_13878.n23 gnd 0.901301f
C1553 a_n2650_13878.n24 gnd 3.52187f
C1554 a_n2650_13878.n25 gnd 2.68251f
C1555 a_n2650_13878.n26 gnd 3.77855f
C1556 a_n2650_13878.n27 gnd 1.18856f
C1557 a_n2650_13878.n28 gnd 1.20779f
C1558 a_n2650_13878.n29 gnd 2.25634f
C1559 a_n2650_13878.n30 gnd 1.79246f
C1560 a_n2650_13878.n31 gnd 1.20779f
C1561 a_n2650_13878.n32 gnd 0.732992f
C1562 a_n2650_13878.n33 gnd 0.732995f
C1563 a_n2650_13878.n34 gnd 3.25198f
C1564 a_n2650_13878.n35 gnd 0.008736f
C1565 a_n2650_13878.n36 gnd 4.21e-19
C1566 a_n2650_13878.n38 gnd 0.008429f
C1567 a_n2650_13878.n39 gnd 0.012257f
C1568 a_n2650_13878.n40 gnd 0.008109f
C1569 a_n2650_13878.n41 gnd 0.287607f
C1570 a_n2650_13878.n42 gnd 0.008736f
C1571 a_n2650_13878.n43 gnd 4.21e-19
C1572 a_n2650_13878.n45 gnd 0.008429f
C1573 a_n2650_13878.n46 gnd 0.012257f
C1574 a_n2650_13878.n47 gnd 0.008109f
C1575 a_n2650_13878.n48 gnd 0.287607f
C1576 a_n2650_13878.n49 gnd 0.008429f
C1577 a_n2650_13878.n50 gnd 0.287607f
C1578 a_n2650_13878.n51 gnd 0.008429f
C1579 a_n2650_13878.n52 gnd 0.287607f
C1580 a_n2650_13878.n53 gnd 0.008429f
C1581 a_n2650_13878.n54 gnd 0.287607f
C1582 a_n2650_13878.n55 gnd 0.008429f
C1583 a_n2650_13878.n56 gnd 0.287607f
C1584 a_n2650_13878.n57 gnd 0.008736f
C1585 a_n2650_13878.n58 gnd 4.21e-19
C1586 a_n2650_13878.n60 gnd 0.008429f
C1587 a_n2650_13878.n61 gnd 0.012257f
C1588 a_n2650_13878.n62 gnd 0.008109f
C1589 a_n2650_13878.n63 gnd 0.287607f
C1590 a_n2650_13878.n64 gnd 0.008736f
C1591 a_n2650_13878.n65 gnd 4.21e-19
C1592 a_n2650_13878.n67 gnd 0.008429f
C1593 a_n2650_13878.n68 gnd 0.012257f
C1594 a_n2650_13878.n69 gnd 0.008109f
C1595 a_n2650_13878.n70 gnd 0.287607f
C1596 a_n2650_13878.t6 gnd 0.702438f
C1597 a_n2650_13878.t40 gnd 0.702438f
C1598 a_n2650_13878.t38 gnd 0.702438f
C1599 a_n2650_13878.n71 gnd 0.308697f
C1600 a_n2650_13878.t42 gnd 0.702438f
C1601 a_n2650_13878.t18 gnd 0.702438f
C1602 a_n2650_13878.t30 gnd 0.702438f
C1603 a_n2650_13878.n72 gnd 0.304914f
C1604 a_n2650_13878.t22 gnd 0.702438f
C1605 a_n2650_13878.t28 gnd 0.702438f
C1606 a_n2650_13878.t12 gnd 0.702438f
C1607 a_n2650_13878.n73 gnd 0.308821f
C1608 a_n2650_13878.t98 gnd 0.702438f
C1609 a_n2650_13878.t77 gnd 0.702438f
C1610 a_n2650_13878.t82 gnd 0.702438f
C1611 a_n2650_13878.n74 gnd 0.308697f
C1612 a_n2650_13878.t71 gnd 0.702438f
C1613 a_n2650_13878.t87 gnd 0.702438f
C1614 a_n2650_13878.t95 gnd 0.702438f
C1615 a_n2650_13878.n75 gnd 0.304914f
C1616 a_n2650_13878.t96 gnd 0.702438f
C1617 a_n2650_13878.t66 gnd 0.702438f
C1618 a_n2650_13878.t79 gnd 0.702438f
C1619 a_n2650_13878.n76 gnd 0.308821f
C1620 a_n2650_13878.t21 gnd 1.41401f
C1621 a_n2650_13878.t11 gnd 0.151013f
C1622 a_n2650_13878.t27 gnd 0.151013f
C1623 a_n2650_13878.n77 gnd 1.06373f
C1624 a_n2650_13878.t33 gnd 0.151013f
C1625 a_n2650_13878.t17 gnd 0.151013f
C1626 a_n2650_13878.n78 gnd 1.06373f
C1627 a_n2650_13878.t25 gnd 0.151013f
C1628 a_n2650_13878.t37 gnd 0.151013f
C1629 a_n2650_13878.n79 gnd 1.06373f
C1630 a_n2650_13878.t35 gnd 0.151013f
C1631 a_n2650_13878.t9 gnd 0.151013f
C1632 a_n2650_13878.n80 gnd 1.06373f
C1633 a_n2650_13878.t45 gnd 1.41119f
C1634 a_n2650_13878.t34 gnd 0.702438f
C1635 a_n2650_13878.n81 gnd 0.305176f
C1636 a_n2650_13878.t24 gnd 0.702438f
C1637 a_n2650_13878.t26 gnd 0.702438f
C1638 a_n2650_13878.n82 gnd 0.308697f
C1639 a_n2650_13878.t20 gnd 0.702438f
C1640 a_n2650_13878.t76 gnd 0.702438f
C1641 a_n2650_13878.n83 gnd 0.305176f
C1642 a_n2650_13878.t91 gnd 0.702438f
C1643 a_n2650_13878.t94 gnd 0.702438f
C1644 a_n2650_13878.n84 gnd 0.308697f
C1645 a_n2650_13878.t70 gnd 0.702438f
C1646 a_n2650_13878.n85 gnd 0.299377f
C1647 a_n2650_13878.t93 gnd 0.702438f
C1648 a_n2650_13878.n86 gnd 0.304579f
C1649 a_n2650_13878.t68 gnd 0.702438f
C1650 a_n2650_13878.n87 gnd 0.311475f
C1651 a_n2650_13878.t90 gnd 0.702438f
C1652 a_n2650_13878.n88 gnd 0.308836f
C1653 a_n2650_13878.n89 gnd 0.304914f
C1654 a_n2650_13878.t65 gnd 0.702438f
C1655 a_n2650_13878.n90 gnd 0.299545f
C1656 a_n2650_13878.t86 gnd 0.702438f
C1657 a_n2650_13878.n91 gnd 0.308821f
C1658 a_n2650_13878.t67 gnd 0.714208f
C1659 a_n2650_13878.n92 gnd 0.299377f
C1660 a_n2650_13878.t10 gnd 0.702438f
C1661 a_n2650_13878.n93 gnd 0.304579f
C1662 a_n2650_13878.t32 gnd 0.702438f
C1663 a_n2650_13878.n94 gnd 0.311475f
C1664 a_n2650_13878.t16 gnd 0.702438f
C1665 a_n2650_13878.n95 gnd 0.308836f
C1666 a_n2650_13878.n96 gnd 0.304914f
C1667 a_n2650_13878.t36 gnd 0.702438f
C1668 a_n2650_13878.n97 gnd 0.299545f
C1669 a_n2650_13878.t8 gnd 0.702438f
C1670 a_n2650_13878.n98 gnd 0.308821f
C1671 a_n2650_13878.t44 gnd 0.714208f
C1672 a_n2650_13878.n99 gnd 1.28381f
C1673 a_n2650_13878.t74 gnd 0.702438f
C1674 a_n2650_13878.n100 gnd 0.304914f
C1675 a_n2650_13878.t81 gnd 0.702438f
C1676 a_n2650_13878.n101 gnd 0.304914f
C1677 a_n2650_13878.t72 gnd 0.702438f
C1678 a_n2650_13878.n102 gnd 0.304914f
C1679 a_n2650_13878.t85 gnd 0.702438f
C1680 a_n2650_13878.n103 gnd 0.304914f
C1681 a_n2650_13878.t75 gnd 0.702438f
C1682 a_n2650_13878.n104 gnd 0.299377f
C1683 a_n2650_13878.t99 gnd 0.702438f
C1684 a_n2650_13878.n105 gnd 0.308836f
C1685 a_n2650_13878.t78 gnd 0.714208f
C1686 a_n2650_13878.t88 gnd 0.702438f
C1687 a_n2650_13878.n106 gnd 0.299377f
C1688 a_n2650_13878.t73 gnd 0.702438f
C1689 a_n2650_13878.n107 gnd 0.308836f
C1690 a_n2650_13878.t83 gnd 0.714208f
C1691 a_n2650_13878.t92 gnd 0.702438f
C1692 a_n2650_13878.n108 gnd 0.299377f
C1693 a_n2650_13878.t80 gnd 0.702438f
C1694 a_n2650_13878.n109 gnd 0.308836f
C1695 a_n2650_13878.t97 gnd 0.714208f
C1696 a_n2650_13878.t84 gnd 0.702438f
C1697 a_n2650_13878.n110 gnd 0.299377f
C1698 a_n2650_13878.t64 gnd 0.702438f
C1699 a_n2650_13878.n111 gnd 0.308836f
C1700 a_n2650_13878.t89 gnd 0.714208f
C1701 a_n2650_13878.n112 gnd 1.58548f
C1702 a_n2650_13878.t69 gnd 0.714208f
C1703 a_n2650_13878.n113 gnd 0.305176f
C1704 a_n2650_13878.n114 gnd 0.299545f
C1705 a_n2650_13878.n115 gnd 0.308836f
C1706 a_n2650_13878.n116 gnd 0.311475f
C1707 a_n2650_13878.n117 gnd 0.304579f
C1708 a_n2650_13878.n118 gnd 0.299377f
C1709 a_n2650_13878.t14 gnd 0.714208f
C1710 a_n2650_13878.t63 gnd 0.117454f
C1711 a_n2650_13878.t61 gnd 0.117454f
C1712 a_n2650_13878.n119 gnd 1.03952f
C1713 a_n2650_13878.t1 gnd 0.117454f
C1714 a_n2650_13878.t59 gnd 0.117454f
C1715 a_n2650_13878.n120 gnd 1.03787f
C1716 a_n2650_13878.t51 gnd 0.117454f
C1717 a_n2650_13878.t56 gnd 0.117454f
C1718 a_n2650_13878.n121 gnd 1.03787f
C1719 a_n2650_13878.t0 gnd 0.117454f
C1720 a_n2650_13878.t48 gnd 0.117454f
C1721 a_n2650_13878.n122 gnd 1.03952f
C1722 a_n2650_13878.t57 gnd 0.117454f
C1723 a_n2650_13878.t46 gnd 0.117454f
C1724 a_n2650_13878.n123 gnd 1.03787f
C1725 a_n2650_13878.t54 gnd 0.117454f
C1726 a_n2650_13878.t62 gnd 0.117454f
C1727 a_n2650_13878.n124 gnd 1.03787f
C1728 a_n2650_13878.t5 gnd 0.117454f
C1729 a_n2650_13878.t50 gnd 0.117454f
C1730 a_n2650_13878.n125 gnd 1.03787f
C1731 a_n2650_13878.t49 gnd 0.117454f
C1732 a_n2650_13878.t2 gnd 0.117454f
C1733 a_n2650_13878.n126 gnd 1.03787f
C1734 a_n2650_13878.t47 gnd 0.117454f
C1735 a_n2650_13878.t60 gnd 0.117454f
C1736 a_n2650_13878.n127 gnd 1.03787f
C1737 a_n2650_13878.t4 gnd 0.117454f
C1738 a_n2650_13878.t52 gnd 0.117454f
C1739 a_n2650_13878.n128 gnd 1.03952f
C1740 a_n2650_13878.t3 gnd 0.117454f
C1741 a_n2650_13878.t53 gnd 0.117454f
C1742 a_n2650_13878.n129 gnd 1.03787f
C1743 a_n2650_13878.t55 gnd 0.117454f
C1744 a_n2650_13878.t58 gnd 0.117454f
C1745 a_n2650_13878.n130 gnd 1.03787f
C1746 a_n2650_13878.n131 gnd 0.305176f
C1747 a_n2650_13878.n132 gnd 0.299545f
C1748 a_n2650_13878.n133 gnd 0.308836f
C1749 a_n2650_13878.n134 gnd 0.311475f
C1750 a_n2650_13878.n135 gnd 0.304579f
C1751 a_n2650_13878.n136 gnd 0.299377f
C1752 a_n2650_13878.n137 gnd 0.949281f
C1753 a_n2650_13878.t15 gnd 1.41401f
C1754 a_n2650_13878.t29 gnd 0.151013f
C1755 a_n2650_13878.t13 gnd 0.151013f
C1756 a_n2650_13878.n138 gnd 1.06373f
C1757 a_n2650_13878.t31 gnd 0.151013f
C1758 a_n2650_13878.t23 gnd 0.151013f
C1759 a_n2650_13878.n139 gnd 1.06373f
C1760 a_n2650_13878.t43 gnd 0.151013f
C1761 a_n2650_13878.t19 gnd 0.151013f
C1762 a_n2650_13878.n140 gnd 1.06373f
C1763 a_n2650_13878.t41 gnd 0.151013f
C1764 a_n2650_13878.t39 gnd 0.151013f
C1765 a_n2650_13878.n141 gnd 1.06373f
C1766 a_n2650_13878.n142 gnd 1.45813f
C1767 a_n2650_13878.t7 gnd 1.41119f
C1768 CSoutput.n0 gnd 0.044585f
C1769 CSoutput.t173 gnd 0.294918f
C1770 CSoutput.n1 gnd 0.13317f
C1771 CSoutput.n2 gnd 0.044585f
C1772 CSoutput.t179 gnd 0.294918f
C1773 CSoutput.n3 gnd 0.035337f
C1774 CSoutput.n4 gnd 0.044585f
C1775 CSoutput.t168 gnd 0.294918f
C1776 CSoutput.n5 gnd 0.030471f
C1777 CSoutput.n6 gnd 0.044585f
C1778 CSoutput.t176 gnd 0.294918f
C1779 CSoutput.t160 gnd 0.294918f
C1780 CSoutput.n7 gnd 0.131719f
C1781 CSoutput.n8 gnd 0.044585f
C1782 CSoutput.t181 gnd 0.294918f
C1783 CSoutput.n9 gnd 0.029053f
C1784 CSoutput.n10 gnd 0.044585f
C1785 CSoutput.t169 gnd 0.294918f
C1786 CSoutput.t180 gnd 0.294918f
C1787 CSoutput.n11 gnd 0.131719f
C1788 CSoutput.n12 gnd 0.044585f
C1789 CSoutput.t177 gnd 0.294918f
C1790 CSoutput.n13 gnd 0.030471f
C1791 CSoutput.n14 gnd 0.044585f
C1792 CSoutput.t167 gnd 0.294918f
C1793 CSoutput.t170 gnd 0.294918f
C1794 CSoutput.n15 gnd 0.131719f
C1795 CSoutput.n16 gnd 0.044585f
C1796 CSoutput.t174 gnd 0.294918f
C1797 CSoutput.n17 gnd 0.032545f
C1798 CSoutput.t164 gnd 0.352435f
C1799 CSoutput.t166 gnd 0.294918f
C1800 CSoutput.n18 gnd 0.168154f
C1801 CSoutput.n19 gnd 0.163167f
C1802 CSoutput.n20 gnd 0.189294f
C1803 CSoutput.n21 gnd 0.044585f
C1804 CSoutput.n22 gnd 0.037211f
C1805 CSoutput.n23 gnd 0.131719f
C1806 CSoutput.n24 gnd 0.03587f
C1807 CSoutput.n25 gnd 0.035337f
C1808 CSoutput.n26 gnd 0.044585f
C1809 CSoutput.n27 gnd 0.044585f
C1810 CSoutput.n28 gnd 0.036925f
C1811 CSoutput.n29 gnd 0.03135f
C1812 CSoutput.n30 gnd 0.134651f
C1813 CSoutput.n31 gnd 0.031782f
C1814 CSoutput.n32 gnd 0.044585f
C1815 CSoutput.n33 gnd 0.044585f
C1816 CSoutput.n34 gnd 0.044585f
C1817 CSoutput.n35 gnd 0.036532f
C1818 CSoutput.n36 gnd 0.131719f
C1819 CSoutput.n37 gnd 0.034937f
C1820 CSoutput.n38 gnd 0.03627f
C1821 CSoutput.n39 gnd 0.044585f
C1822 CSoutput.n40 gnd 0.044585f
C1823 CSoutput.n41 gnd 0.037203f
C1824 CSoutput.n42 gnd 0.034004f
C1825 CSoutput.n43 gnd 0.131719f
C1826 CSoutput.n44 gnd 0.034866f
C1827 CSoutput.n45 gnd 0.044585f
C1828 CSoutput.n46 gnd 0.044585f
C1829 CSoutput.n47 gnd 0.044585f
C1830 CSoutput.n48 gnd 0.034866f
C1831 CSoutput.n49 gnd 0.131719f
C1832 CSoutput.n50 gnd 0.034004f
C1833 CSoutput.n51 gnd 0.037203f
C1834 CSoutput.n52 gnd 0.044585f
C1835 CSoutput.n53 gnd 0.044585f
C1836 CSoutput.n54 gnd 0.03627f
C1837 CSoutput.n55 gnd 0.034937f
C1838 CSoutput.n56 gnd 0.131719f
C1839 CSoutput.n57 gnd 0.036532f
C1840 CSoutput.n58 gnd 0.044585f
C1841 CSoutput.n59 gnd 0.044585f
C1842 CSoutput.n60 gnd 0.044585f
C1843 CSoutput.n61 gnd 0.031782f
C1844 CSoutput.n62 gnd 0.134651f
C1845 CSoutput.n63 gnd 0.03135f
C1846 CSoutput.t162 gnd 0.294918f
C1847 CSoutput.n64 gnd 0.131719f
C1848 CSoutput.n65 gnd 0.036925f
C1849 CSoutput.n66 gnd 0.044585f
C1850 CSoutput.n67 gnd 0.044585f
C1851 CSoutput.n68 gnd 0.044585f
C1852 CSoutput.n69 gnd 0.03587f
C1853 CSoutput.n70 gnd 0.131719f
C1854 CSoutput.n71 gnd 0.037211f
C1855 CSoutput.n72 gnd 0.032545f
C1856 CSoutput.n73 gnd 0.044585f
C1857 CSoutput.n74 gnd 0.044585f
C1858 CSoutput.n75 gnd 0.033751f
C1859 CSoutput.n76 gnd 0.020045f
C1860 CSoutput.t165 gnd 0.331362f
C1861 CSoutput.n77 gnd 0.164607f
C1862 CSoutput.n78 gnd 0.704339f
C1863 CSoutput.t54 gnd 0.055613f
C1864 CSoutput.t103 gnd 0.055613f
C1865 CSoutput.n79 gnd 0.430575f
C1866 CSoutput.t60 gnd 0.055613f
C1867 CSoutput.t83 gnd 0.055613f
C1868 CSoutput.n80 gnd 0.429808f
C1869 CSoutput.n81 gnd 0.436254f
C1870 CSoutput.t142 gnd 0.055613f
C1871 CSoutput.t97 gnd 0.055613f
C1872 CSoutput.n82 gnd 0.429808f
C1873 CSoutput.n83 gnd 0.214968f
C1874 CSoutput.t62 gnd 0.055613f
C1875 CSoutput.t129 gnd 0.055613f
C1876 CSoutput.n84 gnd 0.429808f
C1877 CSoutput.n85 gnd 0.214968f
C1878 CSoutput.t69 gnd 0.055613f
C1879 CSoutput.t112 gnd 0.055613f
C1880 CSoutput.n86 gnd 0.429808f
C1881 CSoutput.n87 gnd 0.214968f
C1882 CSoutput.t87 gnd 0.055613f
C1883 CSoutput.t104 gnd 0.055613f
C1884 CSoutput.n88 gnd 0.429808f
C1885 CSoutput.n89 gnd 0.214968f
C1886 CSoutput.t100 gnd 0.055613f
C1887 CSoutput.t134 gnd 0.055613f
C1888 CSoutput.n90 gnd 0.429808f
C1889 CSoutput.n91 gnd 0.214968f
C1890 CSoutput.t76 gnd 0.055613f
C1891 CSoutput.t117 gnd 0.055613f
C1892 CSoutput.n92 gnd 0.429808f
C1893 CSoutput.n93 gnd 0.394201f
C1894 CSoutput.t72 gnd 0.055613f
C1895 CSoutput.t135 gnd 0.055613f
C1896 CSoutput.n94 gnd 0.430575f
C1897 CSoutput.t110 gnd 0.055613f
C1898 CSoutput.t109 gnd 0.055613f
C1899 CSoutput.n95 gnd 0.429808f
C1900 CSoutput.n96 gnd 0.436254f
C1901 CSoutput.t101 gnd 0.055613f
C1902 CSoutput.t70 gnd 0.055613f
C1903 CSoutput.n97 gnd 0.429808f
C1904 CSoutput.n98 gnd 0.214968f
C1905 CSoutput.t53 gnd 0.055613f
C1906 CSoutput.t102 gnd 0.055613f
C1907 CSoutput.n99 gnd 0.429808f
C1908 CSoutput.n100 gnd 0.214968f
C1909 CSoutput.t98 gnd 0.055613f
C1910 CSoutput.t68 gnd 0.055613f
C1911 CSoutput.n101 gnd 0.429808f
C1912 CSoutput.n102 gnd 0.214968f
C1913 CSoutput.t51 gnd 0.055613f
C1914 CSoutput.t49 gnd 0.055613f
C1915 CSoutput.n103 gnd 0.429808f
C1916 CSoutput.n104 gnd 0.214968f
C1917 CSoutput.t113 gnd 0.055613f
C1918 CSoutput.t84 gnd 0.055613f
C1919 CSoutput.n105 gnd 0.429808f
C1920 CSoutput.n106 gnd 0.214968f
C1921 CSoutput.t78 gnd 0.055613f
C1922 CSoutput.t48 gnd 0.055613f
C1923 CSoutput.n107 gnd 0.429808f
C1924 CSoutput.n108 gnd 0.320571f
C1925 CSoutput.n109 gnd 0.404238f
C1926 CSoutput.t88 gnd 0.055613f
C1927 CSoutput.t143 gnd 0.055613f
C1928 CSoutput.n110 gnd 0.430575f
C1929 CSoutput.t120 gnd 0.055613f
C1930 CSoutput.t119 gnd 0.055613f
C1931 CSoutput.n111 gnd 0.429808f
C1932 CSoutput.n112 gnd 0.436254f
C1933 CSoutput.t107 gnd 0.055613f
C1934 CSoutput.t85 gnd 0.055613f
C1935 CSoutput.n113 gnd 0.429808f
C1936 CSoutput.n114 gnd 0.214968f
C1937 CSoutput.t65 gnd 0.055613f
C1938 CSoutput.t108 gnd 0.055613f
C1939 CSoutput.n115 gnd 0.429808f
C1940 CSoutput.n116 gnd 0.214968f
C1941 CSoutput.t106 gnd 0.055613f
C1942 CSoutput.t82 gnd 0.055613f
C1943 CSoutput.n117 gnd 0.429808f
C1944 CSoutput.n118 gnd 0.214968f
C1945 CSoutput.t64 gnd 0.055613f
C1946 CSoutput.t63 gnd 0.055613f
C1947 CSoutput.n119 gnd 0.429808f
C1948 CSoutput.n120 gnd 0.214968f
C1949 CSoutput.t121 gnd 0.055613f
C1950 CSoutput.t94 gnd 0.055613f
C1951 CSoutput.n121 gnd 0.429808f
C1952 CSoutput.n122 gnd 0.214968f
C1953 CSoutput.t91 gnd 0.055613f
C1954 CSoutput.t59 gnd 0.055613f
C1955 CSoutput.n123 gnd 0.429808f
C1956 CSoutput.n124 gnd 0.320571f
C1957 CSoutput.n125 gnd 0.451834f
C1958 CSoutput.n126 gnd 8.919849f
C1959 CSoutput.n128 gnd 0.788695f
C1960 CSoutput.n129 gnd 0.591522f
C1961 CSoutput.n130 gnd 0.788695f
C1962 CSoutput.n131 gnd 0.788695f
C1963 CSoutput.n132 gnd 2.12341f
C1964 CSoutput.n133 gnd 0.788695f
C1965 CSoutput.n134 gnd 0.788695f
C1966 CSoutput.t161 gnd 0.985869f
C1967 CSoutput.n135 gnd 0.788695f
C1968 CSoutput.n136 gnd 0.788695f
C1969 CSoutput.n140 gnd 0.788695f
C1970 CSoutput.n144 gnd 0.788695f
C1971 CSoutput.n145 gnd 0.788695f
C1972 CSoutput.n147 gnd 0.788695f
C1973 CSoutput.n152 gnd 0.788695f
C1974 CSoutput.n154 gnd 0.788695f
C1975 CSoutput.n155 gnd 0.788695f
C1976 CSoutput.n157 gnd 0.788695f
C1977 CSoutput.n158 gnd 0.788695f
C1978 CSoutput.n160 gnd 0.788695f
C1979 CSoutput.t172 gnd 13.179f
C1980 CSoutput.n162 gnd 0.788695f
C1981 CSoutput.n163 gnd 0.591522f
C1982 CSoutput.n164 gnd 0.788695f
C1983 CSoutput.n165 gnd 0.788695f
C1984 CSoutput.n166 gnd 2.12341f
C1985 CSoutput.n167 gnd 0.788695f
C1986 CSoutput.n168 gnd 0.788695f
C1987 CSoutput.t175 gnd 0.985869f
C1988 CSoutput.n169 gnd 0.788695f
C1989 CSoutput.n170 gnd 0.788695f
C1990 CSoutput.n174 gnd 0.788695f
C1991 CSoutput.n178 gnd 0.788695f
C1992 CSoutput.n179 gnd 0.788695f
C1993 CSoutput.n181 gnd 0.788695f
C1994 CSoutput.n186 gnd 0.788695f
C1995 CSoutput.n188 gnd 0.788695f
C1996 CSoutput.n189 gnd 0.788695f
C1997 CSoutput.n191 gnd 0.788695f
C1998 CSoutput.n192 gnd 0.788695f
C1999 CSoutput.n194 gnd 0.788695f
C2000 CSoutput.n195 gnd 0.591522f
C2001 CSoutput.n197 gnd 0.788695f
C2002 CSoutput.n198 gnd 0.591522f
C2003 CSoutput.n199 gnd 0.788695f
C2004 CSoutput.n200 gnd 0.788695f
C2005 CSoutput.n201 gnd 2.12341f
C2006 CSoutput.n202 gnd 0.788695f
C2007 CSoutput.n203 gnd 0.788695f
C2008 CSoutput.t171 gnd 0.985869f
C2009 CSoutput.n204 gnd 0.788695f
C2010 CSoutput.n205 gnd 2.12341f
C2011 CSoutput.n207 gnd 0.788695f
C2012 CSoutput.n208 gnd 0.788695f
C2013 CSoutput.n210 gnd 0.788695f
C2014 CSoutput.n211 gnd 0.788695f
C2015 CSoutput.t178 gnd 12.9642f
C2016 CSoutput.t163 gnd 13.179f
C2017 CSoutput.n217 gnd 2.47425f
C2018 CSoutput.n218 gnd 10.0792f
C2019 CSoutput.n219 gnd 10.501f
C2020 CSoutput.n224 gnd 2.68028f
C2021 CSoutput.n230 gnd 0.788695f
C2022 CSoutput.n232 gnd 0.788695f
C2023 CSoutput.n234 gnd 0.788695f
C2024 CSoutput.n236 gnd 0.788695f
C2025 CSoutput.n238 gnd 0.788695f
C2026 CSoutput.n244 gnd 0.788695f
C2027 CSoutput.n251 gnd 1.44695f
C2028 CSoutput.n252 gnd 1.44695f
C2029 CSoutput.n253 gnd 0.788695f
C2030 CSoutput.n254 gnd 0.788695f
C2031 CSoutput.n256 gnd 0.591522f
C2032 CSoutput.n257 gnd 0.506585f
C2033 CSoutput.n259 gnd 0.591522f
C2034 CSoutput.n260 gnd 0.506585f
C2035 CSoutput.n261 gnd 0.591522f
C2036 CSoutput.n263 gnd 0.788695f
C2037 CSoutput.n265 gnd 2.12341f
C2038 CSoutput.n266 gnd 2.47425f
C2039 CSoutput.n267 gnd 9.27028f
C2040 CSoutput.n269 gnd 0.591522f
C2041 CSoutput.n270 gnd 1.52202f
C2042 CSoutput.n271 gnd 0.591522f
C2043 CSoutput.n273 gnd 0.788695f
C2044 CSoutput.n275 gnd 2.12341f
C2045 CSoutput.n276 gnd 4.62513f
C2046 CSoutput.t122 gnd 0.055613f
C2047 CSoutput.t52 gnd 0.055613f
C2048 CSoutput.n277 gnd 0.430575f
C2049 CSoutput.t81 gnd 0.055613f
C2050 CSoutput.t58 gnd 0.055613f
C2051 CSoutput.n278 gnd 0.429808f
C2052 CSoutput.n279 gnd 0.436254f
C2053 CSoutput.t96 gnd 0.055613f
C2054 CSoutput.t75 gnd 0.055613f
C2055 CSoutput.n280 gnd 0.429808f
C2056 CSoutput.n281 gnd 0.214968f
C2057 CSoutput.t128 gnd 0.055613f
C2058 CSoutput.t61 gnd 0.055613f
C2059 CSoutput.n282 gnd 0.429808f
C2060 CSoutput.n283 gnd 0.214968f
C2061 CSoutput.t111 gnd 0.055613f
C2062 CSoutput.t66 gnd 0.055613f
C2063 CSoutput.n284 gnd 0.429808f
C2064 CSoutput.n285 gnd 0.214968f
C2065 CSoutput.t124 gnd 0.055613f
C2066 CSoutput.t86 gnd 0.055613f
C2067 CSoutput.n286 gnd 0.429808f
C2068 CSoutput.n287 gnd 0.214968f
C2069 CSoutput.t133 gnd 0.055613f
C2070 CSoutput.t99 gnd 0.055613f
C2071 CSoutput.n288 gnd 0.429808f
C2072 CSoutput.n289 gnd 0.214968f
C2073 CSoutput.t116 gnd 0.055613f
C2074 CSoutput.t77 gnd 0.055613f
C2075 CSoutput.n290 gnd 0.429808f
C2076 CSoutput.n291 gnd 0.394201f
C2077 CSoutput.t80 gnd 0.055613f
C2078 CSoutput.t132 gnd 0.055613f
C2079 CSoutput.n292 gnd 0.430575f
C2080 CSoutput.t73 gnd 0.055613f
C2081 CSoutput.t74 gnd 0.055613f
C2082 CSoutput.n293 gnd 0.429808f
C2083 CSoutput.n294 gnd 0.436254f
C2084 CSoutput.t130 gnd 0.055613f
C2085 CSoutput.t131 gnd 0.055613f
C2086 CSoutput.n295 gnd 0.429808f
C2087 CSoutput.n296 gnd 0.214968f
C2088 CSoutput.t57 gnd 0.055613f
C2089 CSoutput.t118 gnd 0.055613f
C2090 CSoutput.n297 gnd 0.429808f
C2091 CSoutput.n298 gnd 0.214968f
C2092 CSoutput.t127 gnd 0.055613f
C2093 CSoutput.t55 gnd 0.055613f
C2094 CSoutput.n299 gnd 0.429808f
C2095 CSoutput.n300 gnd 0.214968f
C2096 CSoutput.t95 gnd 0.055613f
C2097 CSoutput.t115 gnd 0.055613f
C2098 CSoutput.n301 gnd 0.429808f
C2099 CSoutput.n302 gnd 0.214968f
C2100 CSoutput.t137 gnd 0.055613f
C2101 CSoutput.t79 gnd 0.055613f
C2102 CSoutput.n303 gnd 0.429808f
C2103 CSoutput.n304 gnd 0.214968f
C2104 CSoutput.t114 gnd 0.055613f
C2105 CSoutput.t141 gnd 0.055613f
C2106 CSoutput.n305 gnd 0.429808f
C2107 CSoutput.n306 gnd 0.320571f
C2108 CSoutput.n307 gnd 0.404238f
C2109 CSoutput.t93 gnd 0.055613f
C2110 CSoutput.t140 gnd 0.055613f
C2111 CSoutput.n308 gnd 0.430575f
C2112 CSoutput.t89 gnd 0.055613f
C2113 CSoutput.t90 gnd 0.055613f
C2114 CSoutput.n309 gnd 0.429808f
C2115 CSoutput.n310 gnd 0.436254f
C2116 CSoutput.t138 gnd 0.055613f
C2117 CSoutput.t139 gnd 0.055613f
C2118 CSoutput.n311 gnd 0.429808f
C2119 CSoutput.n312 gnd 0.214968f
C2120 CSoutput.t71 gnd 0.055613f
C2121 CSoutput.t126 gnd 0.055613f
C2122 CSoutput.n313 gnd 0.429808f
C2123 CSoutput.n314 gnd 0.214968f
C2124 CSoutput.t136 gnd 0.055613f
C2125 CSoutput.t67 gnd 0.055613f
C2126 CSoutput.n315 gnd 0.429808f
C2127 CSoutput.n316 gnd 0.214968f
C2128 CSoutput.t105 gnd 0.055613f
C2129 CSoutput.t125 gnd 0.055613f
C2130 CSoutput.n317 gnd 0.429808f
C2131 CSoutput.n318 gnd 0.214968f
C2132 CSoutput.t50 gnd 0.055613f
C2133 CSoutput.t92 gnd 0.055613f
C2134 CSoutput.n319 gnd 0.429808f
C2135 CSoutput.n320 gnd 0.214968f
C2136 CSoutput.t123 gnd 0.055613f
C2137 CSoutput.t56 gnd 0.055613f
C2138 CSoutput.n321 gnd 0.429806f
C2139 CSoutput.n322 gnd 0.320572f
C2140 CSoutput.n323 gnd 0.451834f
C2141 CSoutput.n324 gnd 12.496f
C2142 CSoutput.t7 gnd 0.048662f
C2143 CSoutput.t25 gnd 0.048662f
C2144 CSoutput.n325 gnd 0.431429f
C2145 CSoutput.t27 gnd 0.048662f
C2146 CSoutput.t147 gnd 0.048662f
C2147 CSoutput.n326 gnd 0.42999f
C2148 CSoutput.n327 gnd 0.40067f
C2149 CSoutput.t8 gnd 0.048662f
C2150 CSoutput.t150 gnd 0.048662f
C2151 CSoutput.n328 gnd 0.42999f
C2152 CSoutput.n329 gnd 0.197512f
C2153 CSoutput.t15 gnd 0.048662f
C2154 CSoutput.t43 gnd 0.048662f
C2155 CSoutput.n330 gnd 0.42999f
C2156 CSoutput.n331 gnd 0.197512f
C2157 CSoutput.t46 gnd 0.048662f
C2158 CSoutput.t152 gnd 0.048662f
C2159 CSoutput.n332 gnd 0.42999f
C2160 CSoutput.n333 gnd 0.197512f
C2161 CSoutput.t153 gnd 0.048662f
C2162 CSoutput.t16 gnd 0.048662f
C2163 CSoutput.n334 gnd 0.42999f
C2164 CSoutput.n335 gnd 0.197512f
C2165 CSoutput.t44 gnd 0.048662f
C2166 CSoutput.t10 gnd 0.048662f
C2167 CSoutput.n336 gnd 0.42999f
C2168 CSoutput.n337 gnd 0.197512f
C2169 CSoutput.t0 gnd 0.048662f
C2170 CSoutput.t20 gnd 0.048662f
C2171 CSoutput.n338 gnd 0.42999f
C2172 CSoutput.n339 gnd 0.364251f
C2173 CSoutput.t144 gnd 0.048662f
C2174 CSoutput.t36 gnd 0.048662f
C2175 CSoutput.n340 gnd 0.431429f
C2176 CSoutput.t32 gnd 0.048662f
C2177 CSoutput.t13 gnd 0.048662f
C2178 CSoutput.n341 gnd 0.42999f
C2179 CSoutput.n342 gnd 0.40067f
C2180 CSoutput.t33 gnd 0.048662f
C2181 CSoutput.t37 gnd 0.048662f
C2182 CSoutput.n343 gnd 0.42999f
C2183 CSoutput.n344 gnd 0.197512f
C2184 CSoutput.t159 gnd 0.048662f
C2185 CSoutput.t18 gnd 0.048662f
C2186 CSoutput.n345 gnd 0.42999f
C2187 CSoutput.n346 gnd 0.197512f
C2188 CSoutput.t35 gnd 0.048662f
C2189 CSoutput.t17 gnd 0.048662f
C2190 CSoutput.n347 gnd 0.42999f
C2191 CSoutput.n348 gnd 0.197512f
C2192 CSoutput.t28 gnd 0.048662f
C2193 CSoutput.t21 gnd 0.048662f
C2194 CSoutput.n349 gnd 0.42999f
C2195 CSoutput.n350 gnd 0.197512f
C2196 CSoutput.t145 gnd 0.048662f
C2197 CSoutput.t45 gnd 0.048662f
C2198 CSoutput.n351 gnd 0.42999f
C2199 CSoutput.n352 gnd 0.197512f
C2200 CSoutput.t29 gnd 0.048662f
C2201 CSoutput.t42 gnd 0.048662f
C2202 CSoutput.n353 gnd 0.42999f
C2203 CSoutput.n354 gnd 0.299865f
C2204 CSoutput.n355 gnd 0.557172f
C2205 CSoutput.n356 gnd 12.9547f
C2206 CSoutput.t3 gnd 0.048662f
C2207 CSoutput.t148 gnd 0.048662f
C2208 CSoutput.n357 gnd 0.431429f
C2209 CSoutput.t2 gnd 0.048662f
C2210 CSoutput.t19 gnd 0.048662f
C2211 CSoutput.n358 gnd 0.42999f
C2212 CSoutput.n359 gnd 0.40067f
C2213 CSoutput.t149 gnd 0.048662f
C2214 CSoutput.t151 gnd 0.048662f
C2215 CSoutput.n360 gnd 0.42999f
C2216 CSoutput.n361 gnd 0.197512f
C2217 CSoutput.t1 gnd 0.048662f
C2218 CSoutput.t154 gnd 0.048662f
C2219 CSoutput.n362 gnd 0.42999f
C2220 CSoutput.n363 gnd 0.197512f
C2221 CSoutput.t158 gnd 0.048662f
C2222 CSoutput.t40 gnd 0.048662f
C2223 CSoutput.n364 gnd 0.42999f
C2224 CSoutput.n365 gnd 0.197512f
C2225 CSoutput.t156 gnd 0.048662f
C2226 CSoutput.t5 gnd 0.048662f
C2227 CSoutput.n366 gnd 0.42999f
C2228 CSoutput.n367 gnd 0.197512f
C2229 CSoutput.t47 gnd 0.048662f
C2230 CSoutput.t155 gnd 0.048662f
C2231 CSoutput.n368 gnd 0.42999f
C2232 CSoutput.n369 gnd 0.197512f
C2233 CSoutput.t6 gnd 0.048662f
C2234 CSoutput.t146 gnd 0.048662f
C2235 CSoutput.n370 gnd 0.42999f
C2236 CSoutput.n371 gnd 0.364251f
C2237 CSoutput.t22 gnd 0.048662f
C2238 CSoutput.t24 gnd 0.048662f
C2239 CSoutput.n372 gnd 0.431429f
C2240 CSoutput.t34 gnd 0.048662f
C2241 CSoutput.t11 gnd 0.048662f
C2242 CSoutput.n373 gnd 0.42999f
C2243 CSoutput.n374 gnd 0.40067f
C2244 CSoutput.t39 gnd 0.048662f
C2245 CSoutput.t38 gnd 0.048662f
C2246 CSoutput.n375 gnd 0.42999f
C2247 CSoutput.n376 gnd 0.197512f
C2248 CSoutput.t14 gnd 0.048662f
C2249 CSoutput.t4 gnd 0.048662f
C2250 CSoutput.n377 gnd 0.42999f
C2251 CSoutput.n378 gnd 0.197512f
C2252 CSoutput.t41 gnd 0.048662f
C2253 CSoutput.t23 gnd 0.048662f
C2254 CSoutput.n379 gnd 0.42999f
C2255 CSoutput.n380 gnd 0.197512f
C2256 CSoutput.t9 gnd 0.048662f
C2257 CSoutput.t157 gnd 0.048662f
C2258 CSoutput.n381 gnd 0.42999f
C2259 CSoutput.n382 gnd 0.197512f
C2260 CSoutput.t26 gnd 0.048662f
C2261 CSoutput.t31 gnd 0.048662f
C2262 CSoutput.n383 gnd 0.42999f
C2263 CSoutput.n384 gnd 0.197512f
C2264 CSoutput.t30 gnd 0.048662f
C2265 CSoutput.t12 gnd 0.048662f
C2266 CSoutput.n385 gnd 0.42999f
C2267 CSoutput.n386 gnd 0.299865f
C2268 CSoutput.n387 gnd 0.557172f
C2269 CSoutput.n388 gnd 7.74668f
C2270 CSoutput.n389 gnd 14.352401f
C2271 vdd.t267 gnd 0.035806f
C2272 vdd.t271 gnd 0.035806f
C2273 vdd.n0 gnd 0.282409f
C2274 vdd.t263 gnd 0.035806f
C2275 vdd.t6 gnd 0.035806f
C2276 vdd.n1 gnd 0.281942f
C2277 vdd.n2 gnd 0.260005f
C2278 vdd.t15 gnd 0.035806f
C2279 vdd.t259 gnd 0.035806f
C2280 vdd.n3 gnd 0.281942f
C2281 vdd.n4 gnd 0.131494f
C2282 vdd.t261 gnd 0.035806f
C2283 vdd.t112 gnd 0.035806f
C2284 vdd.n5 gnd 0.281942f
C2285 vdd.n6 gnd 0.123383f
C2286 vdd.t22 gnd 0.035806f
C2287 vdd.t17 gnd 0.035806f
C2288 vdd.n7 gnd 0.282409f
C2289 vdd.t269 gnd 0.035806f
C2290 vdd.t265 gnd 0.035806f
C2291 vdd.n8 gnd 0.281942f
C2292 vdd.n9 gnd 0.260005f
C2293 vdd.t115 gnd 0.035806f
C2294 vdd.t2 gnd 0.035806f
C2295 vdd.n10 gnd 0.281942f
C2296 vdd.n11 gnd 0.131494f
C2297 vdd.t120 gnd 0.035806f
C2298 vdd.t117 gnd 0.035806f
C2299 vdd.n12 gnd 0.281942f
C2300 vdd.n13 gnd 0.123383f
C2301 vdd.n14 gnd 0.087229f
C2302 vdd.t127 gnd 0.019892f
C2303 vdd.t121 gnd 0.019892f
C2304 vdd.n15 gnd 0.1831f
C2305 vdd.t128 gnd 0.019892f
C2306 vdd.t125 gnd 0.019892f
C2307 vdd.n16 gnd 0.182564f
C2308 vdd.n17 gnd 0.317719f
C2309 vdd.t33 gnd 0.019892f
C2310 vdd.t10 gnd 0.019892f
C2311 vdd.n18 gnd 0.182564f
C2312 vdd.n19 gnd 0.131444f
C2313 vdd.t129 gnd 0.019892f
C2314 vdd.t122 gnd 0.019892f
C2315 vdd.n20 gnd 0.1831f
C2316 vdd.t32 gnd 0.019892f
C2317 vdd.t12 gnd 0.019892f
C2318 vdd.n21 gnd 0.182564f
C2319 vdd.n22 gnd 0.317719f
C2320 vdd.t123 gnd 0.019892f
C2321 vdd.t124 gnd 0.019892f
C2322 vdd.n23 gnd 0.182564f
C2323 vdd.n24 gnd 0.131444f
C2324 vdd.t24 gnd 0.019892f
C2325 vdd.t11 gnd 0.019892f
C2326 vdd.n25 gnd 0.182564f
C2327 vdd.t25 gnd 0.019892f
C2328 vdd.t126 gnd 0.019892f
C2329 vdd.n26 gnd 0.182564f
C2330 vdd.n27 gnd 21.2232f
C2331 vdd.n28 gnd 8.1529f
C2332 vdd.n29 gnd 0.005425f
C2333 vdd.n30 gnd 0.005035f
C2334 vdd.n31 gnd 0.002785f
C2335 vdd.n32 gnd 0.006394f
C2336 vdd.n33 gnd 0.002705f
C2337 vdd.n34 gnd 0.002864f
C2338 vdd.n35 gnd 0.005035f
C2339 vdd.n36 gnd 0.002705f
C2340 vdd.n37 gnd 0.006394f
C2341 vdd.n38 gnd 0.002864f
C2342 vdd.n39 gnd 0.005035f
C2343 vdd.n40 gnd 0.002705f
C2344 vdd.n41 gnd 0.004796f
C2345 vdd.n42 gnd 0.00481f
C2346 vdd.t239 gnd 0.013738f
C2347 vdd.n43 gnd 0.030567f
C2348 vdd.n44 gnd 0.159077f
C2349 vdd.n45 gnd 0.002705f
C2350 vdd.n46 gnd 0.002864f
C2351 vdd.n47 gnd 0.006394f
C2352 vdd.n48 gnd 0.006394f
C2353 vdd.n49 gnd 0.002864f
C2354 vdd.n50 gnd 0.002705f
C2355 vdd.n51 gnd 0.005035f
C2356 vdd.n52 gnd 0.005035f
C2357 vdd.n53 gnd 0.002705f
C2358 vdd.n54 gnd 0.002864f
C2359 vdd.n55 gnd 0.006394f
C2360 vdd.n56 gnd 0.006394f
C2361 vdd.n57 gnd 0.002864f
C2362 vdd.n58 gnd 0.002705f
C2363 vdd.n59 gnd 0.005035f
C2364 vdd.n60 gnd 0.005035f
C2365 vdd.n61 gnd 0.002705f
C2366 vdd.n62 gnd 0.002864f
C2367 vdd.n63 gnd 0.006394f
C2368 vdd.n64 gnd 0.006394f
C2369 vdd.n65 gnd 0.015118f
C2370 vdd.n66 gnd 0.002785f
C2371 vdd.n67 gnd 0.002705f
C2372 vdd.n68 gnd 0.013013f
C2373 vdd.n69 gnd 0.009085f
C2374 vdd.t139 gnd 0.031828f
C2375 vdd.t184 gnd 0.031828f
C2376 vdd.n70 gnd 0.218742f
C2377 vdd.n71 gnd 0.172007f
C2378 vdd.t152 gnd 0.031828f
C2379 vdd.t204 gnd 0.031828f
C2380 vdd.n72 gnd 0.218742f
C2381 vdd.n73 gnd 0.138808f
C2382 vdd.t175 gnd 0.031828f
C2383 vdd.t243 gnd 0.031828f
C2384 vdd.n74 gnd 0.218742f
C2385 vdd.n75 gnd 0.138808f
C2386 vdd.t156 gnd 0.031828f
C2387 vdd.t224 gnd 0.031828f
C2388 vdd.n76 gnd 0.218742f
C2389 vdd.n77 gnd 0.138808f
C2390 vdd.t163 gnd 0.031828f
C2391 vdd.t235 gnd 0.031828f
C2392 vdd.n78 gnd 0.218742f
C2393 vdd.n79 gnd 0.138808f
C2394 vdd.t192 gnd 0.031828f
C2395 vdd.t247 gnd 0.031828f
C2396 vdd.n80 gnd 0.218742f
C2397 vdd.n81 gnd 0.138808f
C2398 vdd.t207 gnd 0.031828f
C2399 vdd.t230 gnd 0.031828f
C2400 vdd.n82 gnd 0.218742f
C2401 vdd.n83 gnd 0.138808f
C2402 vdd.n84 gnd 0.005425f
C2403 vdd.n85 gnd 0.005035f
C2404 vdd.n86 gnd 0.002785f
C2405 vdd.n87 gnd 0.006394f
C2406 vdd.n88 gnd 0.002705f
C2407 vdd.n89 gnd 0.002864f
C2408 vdd.n90 gnd 0.005035f
C2409 vdd.n91 gnd 0.002705f
C2410 vdd.n92 gnd 0.006394f
C2411 vdd.n93 gnd 0.002864f
C2412 vdd.n94 gnd 0.005035f
C2413 vdd.n95 gnd 0.002705f
C2414 vdd.n96 gnd 0.004796f
C2415 vdd.n97 gnd 0.00481f
C2416 vdd.t178 gnd 0.013738f
C2417 vdd.n98 gnd 0.030567f
C2418 vdd.n99 gnd 0.159077f
C2419 vdd.n100 gnd 0.002705f
C2420 vdd.n101 gnd 0.002864f
C2421 vdd.n102 gnd 0.006394f
C2422 vdd.n103 gnd 0.006394f
C2423 vdd.n104 gnd 0.002864f
C2424 vdd.n105 gnd 0.002705f
C2425 vdd.n106 gnd 0.005035f
C2426 vdd.n107 gnd 0.005035f
C2427 vdd.n108 gnd 0.002705f
C2428 vdd.n109 gnd 0.002864f
C2429 vdd.n110 gnd 0.006394f
C2430 vdd.n111 gnd 0.006394f
C2431 vdd.n112 gnd 0.002864f
C2432 vdd.n113 gnd 0.002705f
C2433 vdd.n114 gnd 0.005035f
C2434 vdd.n115 gnd 0.005035f
C2435 vdd.n116 gnd 0.002705f
C2436 vdd.n117 gnd 0.002864f
C2437 vdd.n118 gnd 0.006394f
C2438 vdd.n119 gnd 0.006394f
C2439 vdd.n120 gnd 0.015118f
C2440 vdd.n121 gnd 0.002785f
C2441 vdd.n122 gnd 0.002705f
C2442 vdd.n123 gnd 0.013013f
C2443 vdd.n124 gnd 0.0088f
C2444 vdd.n125 gnd 0.103274f
C2445 vdd.n126 gnd 0.005425f
C2446 vdd.n127 gnd 0.005035f
C2447 vdd.n128 gnd 0.002785f
C2448 vdd.n129 gnd 0.006394f
C2449 vdd.n130 gnd 0.002705f
C2450 vdd.n131 gnd 0.002864f
C2451 vdd.n132 gnd 0.005035f
C2452 vdd.n133 gnd 0.002705f
C2453 vdd.n134 gnd 0.006394f
C2454 vdd.n135 gnd 0.002864f
C2455 vdd.n136 gnd 0.005035f
C2456 vdd.n137 gnd 0.002705f
C2457 vdd.n138 gnd 0.004796f
C2458 vdd.n139 gnd 0.00481f
C2459 vdd.t183 gnd 0.013738f
C2460 vdd.n140 gnd 0.030567f
C2461 vdd.n141 gnd 0.159077f
C2462 vdd.n142 gnd 0.002705f
C2463 vdd.n143 gnd 0.002864f
C2464 vdd.n144 gnd 0.006394f
C2465 vdd.n145 gnd 0.006394f
C2466 vdd.n146 gnd 0.002864f
C2467 vdd.n147 gnd 0.002705f
C2468 vdd.n148 gnd 0.005035f
C2469 vdd.n149 gnd 0.005035f
C2470 vdd.n150 gnd 0.002705f
C2471 vdd.n151 gnd 0.002864f
C2472 vdd.n152 gnd 0.006394f
C2473 vdd.n153 gnd 0.006394f
C2474 vdd.n154 gnd 0.002864f
C2475 vdd.n155 gnd 0.002705f
C2476 vdd.n156 gnd 0.005035f
C2477 vdd.n157 gnd 0.005035f
C2478 vdd.n158 gnd 0.002705f
C2479 vdd.n159 gnd 0.002864f
C2480 vdd.n160 gnd 0.006394f
C2481 vdd.n161 gnd 0.006394f
C2482 vdd.n162 gnd 0.015118f
C2483 vdd.n163 gnd 0.002785f
C2484 vdd.n164 gnd 0.002705f
C2485 vdd.n165 gnd 0.013013f
C2486 vdd.n166 gnd 0.009085f
C2487 vdd.t246 gnd 0.031828f
C2488 vdd.t172 gnd 0.031828f
C2489 vdd.n167 gnd 0.218742f
C2490 vdd.n168 gnd 0.172007f
C2491 vdd.t173 gnd 0.031828f
C2492 vdd.t234 gnd 0.031828f
C2493 vdd.n169 gnd 0.218742f
C2494 vdd.n170 gnd 0.138808f
C2495 vdd.t245 gnd 0.031828f
C2496 vdd.t150 gnd 0.031828f
C2497 vdd.n171 gnd 0.218742f
C2498 vdd.n172 gnd 0.138808f
C2499 vdd.t232 gnd 0.031828f
C2500 vdd.t242 gnd 0.031828f
C2501 vdd.n173 gnd 0.218742f
C2502 vdd.n174 gnd 0.138808f
C2503 vdd.t146 gnd 0.031828f
C2504 vdd.t202 gnd 0.031828f
C2505 vdd.n175 gnd 0.218742f
C2506 vdd.n176 gnd 0.138808f
C2507 vdd.t229 gnd 0.031828f
C2508 vdd.t251 gnd 0.031828f
C2509 vdd.n177 gnd 0.218742f
C2510 vdd.n178 gnd 0.138808f
C2511 vdd.t181 gnd 0.031828f
C2512 vdd.t228 gnd 0.031828f
C2513 vdd.n179 gnd 0.218742f
C2514 vdd.n180 gnd 0.138808f
C2515 vdd.n181 gnd 0.005425f
C2516 vdd.n182 gnd 0.005035f
C2517 vdd.n183 gnd 0.002785f
C2518 vdd.n184 gnd 0.006394f
C2519 vdd.n185 gnd 0.002705f
C2520 vdd.n186 gnd 0.002864f
C2521 vdd.n187 gnd 0.005035f
C2522 vdd.n188 gnd 0.002705f
C2523 vdd.n189 gnd 0.006394f
C2524 vdd.n190 gnd 0.002864f
C2525 vdd.n191 gnd 0.005035f
C2526 vdd.n192 gnd 0.002705f
C2527 vdd.n193 gnd 0.004796f
C2528 vdd.n194 gnd 0.00481f
C2529 vdd.t255 gnd 0.013738f
C2530 vdd.n195 gnd 0.030567f
C2531 vdd.n196 gnd 0.159077f
C2532 vdd.n197 gnd 0.002705f
C2533 vdd.n198 gnd 0.002864f
C2534 vdd.n199 gnd 0.006394f
C2535 vdd.n200 gnd 0.006394f
C2536 vdd.n201 gnd 0.002864f
C2537 vdd.n202 gnd 0.002705f
C2538 vdd.n203 gnd 0.005035f
C2539 vdd.n204 gnd 0.005035f
C2540 vdd.n205 gnd 0.002705f
C2541 vdd.n206 gnd 0.002864f
C2542 vdd.n207 gnd 0.006394f
C2543 vdd.n208 gnd 0.006394f
C2544 vdd.n209 gnd 0.002864f
C2545 vdd.n210 gnd 0.002705f
C2546 vdd.n211 gnd 0.005035f
C2547 vdd.n212 gnd 0.005035f
C2548 vdd.n213 gnd 0.002705f
C2549 vdd.n214 gnd 0.002864f
C2550 vdd.n215 gnd 0.006394f
C2551 vdd.n216 gnd 0.006394f
C2552 vdd.n217 gnd 0.015118f
C2553 vdd.n218 gnd 0.002785f
C2554 vdd.n219 gnd 0.002705f
C2555 vdd.n220 gnd 0.013013f
C2556 vdd.n221 gnd 0.0088f
C2557 vdd.n222 gnd 0.061438f
C2558 vdd.n223 gnd 0.221376f
C2559 vdd.n224 gnd 0.005425f
C2560 vdd.n225 gnd 0.005035f
C2561 vdd.n226 gnd 0.002785f
C2562 vdd.n227 gnd 0.006394f
C2563 vdd.n228 gnd 0.002705f
C2564 vdd.n229 gnd 0.002864f
C2565 vdd.n230 gnd 0.005035f
C2566 vdd.n231 gnd 0.002705f
C2567 vdd.n232 gnd 0.006394f
C2568 vdd.n233 gnd 0.002864f
C2569 vdd.n234 gnd 0.005035f
C2570 vdd.n235 gnd 0.002705f
C2571 vdd.n236 gnd 0.004796f
C2572 vdd.n237 gnd 0.00481f
C2573 vdd.t199 gnd 0.013738f
C2574 vdd.n238 gnd 0.030567f
C2575 vdd.n239 gnd 0.159077f
C2576 vdd.n240 gnd 0.002705f
C2577 vdd.n241 gnd 0.002864f
C2578 vdd.n242 gnd 0.006394f
C2579 vdd.n243 gnd 0.006394f
C2580 vdd.n244 gnd 0.002864f
C2581 vdd.n245 gnd 0.002705f
C2582 vdd.n246 gnd 0.005035f
C2583 vdd.n247 gnd 0.005035f
C2584 vdd.n248 gnd 0.002705f
C2585 vdd.n249 gnd 0.002864f
C2586 vdd.n250 gnd 0.006394f
C2587 vdd.n251 gnd 0.006394f
C2588 vdd.n252 gnd 0.002864f
C2589 vdd.n253 gnd 0.002705f
C2590 vdd.n254 gnd 0.005035f
C2591 vdd.n255 gnd 0.005035f
C2592 vdd.n256 gnd 0.002705f
C2593 vdd.n257 gnd 0.002864f
C2594 vdd.n258 gnd 0.006394f
C2595 vdd.n259 gnd 0.006394f
C2596 vdd.n260 gnd 0.015118f
C2597 vdd.n261 gnd 0.002785f
C2598 vdd.n262 gnd 0.002705f
C2599 vdd.n263 gnd 0.013013f
C2600 vdd.n264 gnd 0.009085f
C2601 vdd.t254 gnd 0.031828f
C2602 vdd.t195 gnd 0.031828f
C2603 vdd.n265 gnd 0.218742f
C2604 vdd.n266 gnd 0.172007f
C2605 vdd.t196 gnd 0.031828f
C2606 vdd.t252 gnd 0.031828f
C2607 vdd.n267 gnd 0.218742f
C2608 vdd.n268 gnd 0.138808f
C2609 vdd.t253 gnd 0.031828f
C2610 vdd.t169 gnd 0.031828f
C2611 vdd.n269 gnd 0.218742f
C2612 vdd.n270 gnd 0.138808f
C2613 vdd.t233 gnd 0.031828f
C2614 vdd.t250 gnd 0.031828f
C2615 vdd.n271 gnd 0.218742f
C2616 vdd.n272 gnd 0.138808f
C2617 vdd.t164 gnd 0.031828f
C2618 vdd.t217 gnd 0.031828f
C2619 vdd.n273 gnd 0.218742f
C2620 vdd.n274 gnd 0.138808f
C2621 vdd.t241 gnd 0.031828f
C2622 vdd.t135 gnd 0.031828f
C2623 vdd.n275 gnd 0.218742f
C2624 vdd.n276 gnd 0.138808f
C2625 vdd.t198 gnd 0.031828f
C2626 vdd.t240 gnd 0.031828f
C2627 vdd.n277 gnd 0.218742f
C2628 vdd.n278 gnd 0.138808f
C2629 vdd.n279 gnd 0.005425f
C2630 vdd.n280 gnd 0.005035f
C2631 vdd.n281 gnd 0.002785f
C2632 vdd.n282 gnd 0.006394f
C2633 vdd.n283 gnd 0.002705f
C2634 vdd.n284 gnd 0.002864f
C2635 vdd.n285 gnd 0.005035f
C2636 vdd.n286 gnd 0.002705f
C2637 vdd.n287 gnd 0.006394f
C2638 vdd.n288 gnd 0.002864f
C2639 vdd.n289 gnd 0.005035f
C2640 vdd.n290 gnd 0.002705f
C2641 vdd.n291 gnd 0.004796f
C2642 vdd.n292 gnd 0.00481f
C2643 vdd.t148 gnd 0.013738f
C2644 vdd.n293 gnd 0.030567f
C2645 vdd.n294 gnd 0.159077f
C2646 vdd.n295 gnd 0.002705f
C2647 vdd.n296 gnd 0.002864f
C2648 vdd.n297 gnd 0.006394f
C2649 vdd.n298 gnd 0.006394f
C2650 vdd.n299 gnd 0.002864f
C2651 vdd.n300 gnd 0.002705f
C2652 vdd.n301 gnd 0.005035f
C2653 vdd.n302 gnd 0.005035f
C2654 vdd.n303 gnd 0.002705f
C2655 vdd.n304 gnd 0.002864f
C2656 vdd.n305 gnd 0.006394f
C2657 vdd.n306 gnd 0.006394f
C2658 vdd.n307 gnd 0.002864f
C2659 vdd.n308 gnd 0.002705f
C2660 vdd.n309 gnd 0.005035f
C2661 vdd.n310 gnd 0.005035f
C2662 vdd.n311 gnd 0.002705f
C2663 vdd.n312 gnd 0.002864f
C2664 vdd.n313 gnd 0.006394f
C2665 vdd.n314 gnd 0.006394f
C2666 vdd.n315 gnd 0.015118f
C2667 vdd.n316 gnd 0.002785f
C2668 vdd.n317 gnd 0.002705f
C2669 vdd.n318 gnd 0.013013f
C2670 vdd.n319 gnd 0.0088f
C2671 vdd.n320 gnd 0.061438f
C2672 vdd.n321 gnd 0.247912f
C2673 vdd.n322 gnd 0.007598f
C2674 vdd.n323 gnd 0.009886f
C2675 vdd.n324 gnd 0.007957f
C2676 vdd.n325 gnd 0.007957f
C2677 vdd.n326 gnd 0.009886f
C2678 vdd.n327 gnd 0.009886f
C2679 vdd.n328 gnd 0.722355f
C2680 vdd.n329 gnd 0.009886f
C2681 vdd.n330 gnd 0.009886f
C2682 vdd.n331 gnd 0.009886f
C2683 vdd.n332 gnd 0.782973f
C2684 vdd.n333 gnd 0.009886f
C2685 vdd.n334 gnd 0.009886f
C2686 vdd.n335 gnd 0.009886f
C2687 vdd.n336 gnd 0.009886f
C2688 vdd.n337 gnd 0.007957f
C2689 vdd.n338 gnd 0.009886f
C2690 vdd.t201 gnd 0.505144f
C2691 vdd.n339 gnd 0.009886f
C2692 vdd.n340 gnd 0.009886f
C2693 vdd.n341 gnd 0.009886f
C2694 vdd.t134 gnd 0.505144f
C2695 vdd.n342 gnd 0.009886f
C2696 vdd.n343 gnd 0.009886f
C2697 vdd.n344 gnd 0.009886f
C2698 vdd.n345 gnd 0.009886f
C2699 vdd.n346 gnd 0.009886f
C2700 vdd.n347 gnd 0.007957f
C2701 vdd.n348 gnd 0.009886f
C2702 vdd.n349 gnd 0.570812f
C2703 vdd.n350 gnd 0.009886f
C2704 vdd.n351 gnd 0.009886f
C2705 vdd.n352 gnd 0.009886f
C2706 vdd.t227 gnd 0.505144f
C2707 vdd.n353 gnd 0.009886f
C2708 vdd.n354 gnd 0.009886f
C2709 vdd.n355 gnd 0.009886f
C2710 vdd.n356 gnd 0.009886f
C2711 vdd.n357 gnd 0.009886f
C2712 vdd.n358 gnd 0.007957f
C2713 vdd.n359 gnd 0.009886f
C2714 vdd.t147 gnd 0.505144f
C2715 vdd.n360 gnd 0.009886f
C2716 vdd.n361 gnd 0.009886f
C2717 vdd.n362 gnd 0.009886f
C2718 vdd.n363 gnd 0.853693f
C2719 vdd.n364 gnd 0.009886f
C2720 vdd.n365 gnd 0.009886f
C2721 vdd.n366 gnd 0.009886f
C2722 vdd.n367 gnd 0.009886f
C2723 vdd.n368 gnd 0.009886f
C2724 vdd.n369 gnd 0.006604f
C2725 vdd.n370 gnd 0.022512f
C2726 vdd.t51 gnd 0.505144f
C2727 vdd.n371 gnd 0.009886f
C2728 vdd.n372 gnd 0.022512f
C2729 vdd.n404 gnd 0.009886f
C2730 vdd.t67 gnd 0.121622f
C2731 vdd.t66 gnd 0.12998f
C2732 vdd.t65 gnd 0.158837f
C2733 vdd.n405 gnd 0.203606f
C2734 vdd.n406 gnd 0.171862f
C2735 vdd.n407 gnd 0.013049f
C2736 vdd.n408 gnd 0.009886f
C2737 vdd.n409 gnd 0.007957f
C2738 vdd.n410 gnd 0.009886f
C2739 vdd.n411 gnd 0.007957f
C2740 vdd.n412 gnd 0.009886f
C2741 vdd.n413 gnd 0.007957f
C2742 vdd.n414 gnd 0.009886f
C2743 vdd.n415 gnd 0.007957f
C2744 vdd.n416 gnd 0.009886f
C2745 vdd.n417 gnd 0.007957f
C2746 vdd.n418 gnd 0.009886f
C2747 vdd.t53 gnd 0.121622f
C2748 vdd.t52 gnd 0.12998f
C2749 vdd.t50 gnd 0.158837f
C2750 vdd.n419 gnd 0.203606f
C2751 vdd.n420 gnd 0.171862f
C2752 vdd.n421 gnd 0.007957f
C2753 vdd.n422 gnd 0.009886f
C2754 vdd.n423 gnd 0.007957f
C2755 vdd.n424 gnd 0.009886f
C2756 vdd.n425 gnd 0.007957f
C2757 vdd.n426 gnd 0.009886f
C2758 vdd.n427 gnd 0.007957f
C2759 vdd.n428 gnd 0.009886f
C2760 vdd.n429 gnd 0.007957f
C2761 vdd.n430 gnd 0.009886f
C2762 vdd.t74 gnd 0.121622f
C2763 vdd.t73 gnd 0.12998f
C2764 vdd.t72 gnd 0.158837f
C2765 vdd.n431 gnd 0.203606f
C2766 vdd.n432 gnd 0.171862f
C2767 vdd.n433 gnd 0.017028f
C2768 vdd.n434 gnd 0.009886f
C2769 vdd.n435 gnd 0.007957f
C2770 vdd.n436 gnd 0.009886f
C2771 vdd.n437 gnd 0.007957f
C2772 vdd.n438 gnd 0.009886f
C2773 vdd.n439 gnd 0.007957f
C2774 vdd.n440 gnd 0.009886f
C2775 vdd.n441 gnd 0.007957f
C2776 vdd.n442 gnd 0.009886f
C2777 vdd.n443 gnd 0.022512f
C2778 vdd.n444 gnd 0.022666f
C2779 vdd.n445 gnd 0.022666f
C2780 vdd.n446 gnd 0.006604f
C2781 vdd.n447 gnd 0.007957f
C2782 vdd.n448 gnd 0.009886f
C2783 vdd.n449 gnd 0.009886f
C2784 vdd.n450 gnd 0.007957f
C2785 vdd.n451 gnd 0.009886f
C2786 vdd.n452 gnd 0.009886f
C2787 vdd.n453 gnd 0.009886f
C2788 vdd.n454 gnd 0.009886f
C2789 vdd.n455 gnd 0.009886f
C2790 vdd.n456 gnd 0.007957f
C2791 vdd.n457 gnd 0.007957f
C2792 vdd.n458 gnd 0.009886f
C2793 vdd.n459 gnd 0.009886f
C2794 vdd.n460 gnd 0.007957f
C2795 vdd.n461 gnd 0.009886f
C2796 vdd.n462 gnd 0.009886f
C2797 vdd.n463 gnd 0.009886f
C2798 vdd.n464 gnd 0.009886f
C2799 vdd.n465 gnd 0.009886f
C2800 vdd.n466 gnd 0.007957f
C2801 vdd.n467 gnd 0.007957f
C2802 vdd.n468 gnd 0.009886f
C2803 vdd.n469 gnd 0.009886f
C2804 vdd.n470 gnd 0.007957f
C2805 vdd.n471 gnd 0.009886f
C2806 vdd.n472 gnd 0.009886f
C2807 vdd.n473 gnd 0.009886f
C2808 vdd.n474 gnd 0.009886f
C2809 vdd.n475 gnd 0.009886f
C2810 vdd.n476 gnd 0.007957f
C2811 vdd.n477 gnd 0.007957f
C2812 vdd.n478 gnd 0.009886f
C2813 vdd.n479 gnd 0.009886f
C2814 vdd.n480 gnd 0.007957f
C2815 vdd.n481 gnd 0.009886f
C2816 vdd.n482 gnd 0.009886f
C2817 vdd.n483 gnd 0.009886f
C2818 vdd.n484 gnd 0.009886f
C2819 vdd.n485 gnd 0.009886f
C2820 vdd.n486 gnd 0.007957f
C2821 vdd.n487 gnd 0.007957f
C2822 vdd.n488 gnd 0.009886f
C2823 vdd.n489 gnd 0.009886f
C2824 vdd.n490 gnd 0.006644f
C2825 vdd.n491 gnd 0.009886f
C2826 vdd.n492 gnd 0.009886f
C2827 vdd.n493 gnd 0.009886f
C2828 vdd.n494 gnd 0.009886f
C2829 vdd.n495 gnd 0.009886f
C2830 vdd.n496 gnd 0.006644f
C2831 vdd.n497 gnd 0.007957f
C2832 vdd.n498 gnd 0.009886f
C2833 vdd.n499 gnd 0.009886f
C2834 vdd.n500 gnd 0.007957f
C2835 vdd.n501 gnd 0.009886f
C2836 vdd.n502 gnd 0.009886f
C2837 vdd.n503 gnd 0.009886f
C2838 vdd.n504 gnd 0.009886f
C2839 vdd.n505 gnd 0.009886f
C2840 vdd.n506 gnd 0.007957f
C2841 vdd.n507 gnd 0.007957f
C2842 vdd.n508 gnd 0.009886f
C2843 vdd.n509 gnd 0.009886f
C2844 vdd.n510 gnd 0.007957f
C2845 vdd.n511 gnd 0.009886f
C2846 vdd.n512 gnd 0.009886f
C2847 vdd.n513 gnd 0.009886f
C2848 vdd.n514 gnd 0.009886f
C2849 vdd.n515 gnd 0.009886f
C2850 vdd.n516 gnd 0.007957f
C2851 vdd.n517 gnd 0.007957f
C2852 vdd.n518 gnd 0.009886f
C2853 vdd.n519 gnd 0.009886f
C2854 vdd.n520 gnd 0.007957f
C2855 vdd.n521 gnd 0.009886f
C2856 vdd.n522 gnd 0.009886f
C2857 vdd.n523 gnd 0.009886f
C2858 vdd.n524 gnd 0.009886f
C2859 vdd.n525 gnd 0.009886f
C2860 vdd.n526 gnd 0.007957f
C2861 vdd.n527 gnd 0.007957f
C2862 vdd.n528 gnd 0.009886f
C2863 vdd.n529 gnd 0.009886f
C2864 vdd.n530 gnd 0.007957f
C2865 vdd.n531 gnd 0.009886f
C2866 vdd.n532 gnd 0.009886f
C2867 vdd.n533 gnd 0.009886f
C2868 vdd.n534 gnd 0.009886f
C2869 vdd.n535 gnd 0.009886f
C2870 vdd.n536 gnd 0.007957f
C2871 vdd.n537 gnd 0.007957f
C2872 vdd.n538 gnd 0.009886f
C2873 vdd.n539 gnd 0.009886f
C2874 vdd.n540 gnd 0.007957f
C2875 vdd.n541 gnd 0.009886f
C2876 vdd.n542 gnd 0.009886f
C2877 vdd.n543 gnd 0.009886f
C2878 vdd.n544 gnd 0.009886f
C2879 vdd.n545 gnd 0.009886f
C2880 vdd.n546 gnd 0.005411f
C2881 vdd.n547 gnd 0.017028f
C2882 vdd.n548 gnd 0.009886f
C2883 vdd.n549 gnd 0.009886f
C2884 vdd.n550 gnd 0.007877f
C2885 vdd.n551 gnd 0.009886f
C2886 vdd.n552 gnd 0.009886f
C2887 vdd.n553 gnd 0.009886f
C2888 vdd.n554 gnd 0.009886f
C2889 vdd.n555 gnd 0.009886f
C2890 vdd.n556 gnd 0.007957f
C2891 vdd.n557 gnd 0.007957f
C2892 vdd.n558 gnd 0.009886f
C2893 vdd.n559 gnd 0.009886f
C2894 vdd.n560 gnd 0.007957f
C2895 vdd.n561 gnd 0.009886f
C2896 vdd.n562 gnd 0.009886f
C2897 vdd.n563 gnd 0.009886f
C2898 vdd.n564 gnd 0.009886f
C2899 vdd.n565 gnd 0.009886f
C2900 vdd.n566 gnd 0.007957f
C2901 vdd.n567 gnd 0.007957f
C2902 vdd.n568 gnd 0.009886f
C2903 vdd.n569 gnd 0.009886f
C2904 vdd.n570 gnd 0.007957f
C2905 vdd.n571 gnd 0.009886f
C2906 vdd.n572 gnd 0.009886f
C2907 vdd.n573 gnd 0.009886f
C2908 vdd.n574 gnd 0.009886f
C2909 vdd.n575 gnd 0.009886f
C2910 vdd.n576 gnd 0.007957f
C2911 vdd.n577 gnd 0.007957f
C2912 vdd.n578 gnd 0.009886f
C2913 vdd.n579 gnd 0.009886f
C2914 vdd.n580 gnd 0.007957f
C2915 vdd.n581 gnd 0.009886f
C2916 vdd.n582 gnd 0.009886f
C2917 vdd.n583 gnd 0.009886f
C2918 vdd.n584 gnd 0.009886f
C2919 vdd.n585 gnd 0.009886f
C2920 vdd.n586 gnd 0.007957f
C2921 vdd.n587 gnd 0.007957f
C2922 vdd.n588 gnd 0.009886f
C2923 vdd.n589 gnd 0.009886f
C2924 vdd.n590 gnd 0.007957f
C2925 vdd.n591 gnd 0.009886f
C2926 vdd.n592 gnd 0.009886f
C2927 vdd.n593 gnd 0.009886f
C2928 vdd.n594 gnd 0.009886f
C2929 vdd.n595 gnd 0.009886f
C2930 vdd.n596 gnd 0.007957f
C2931 vdd.n597 gnd 0.009886f
C2932 vdd.n598 gnd 0.007957f
C2933 vdd.n599 gnd 0.004177f
C2934 vdd.n600 gnd 0.009886f
C2935 vdd.n601 gnd 0.009886f
C2936 vdd.n602 gnd 0.007957f
C2937 vdd.n603 gnd 0.009886f
C2938 vdd.n604 gnd 0.007957f
C2939 vdd.n605 gnd 0.009886f
C2940 vdd.n606 gnd 0.007957f
C2941 vdd.n607 gnd 0.009886f
C2942 vdd.n608 gnd 0.007957f
C2943 vdd.n609 gnd 0.009886f
C2944 vdd.n610 gnd 0.007957f
C2945 vdd.n611 gnd 0.009886f
C2946 vdd.n612 gnd 0.009886f
C2947 vdd.n613 gnd 0.550607f
C2948 vdd.t155 gnd 0.505144f
C2949 vdd.n614 gnd 0.009886f
C2950 vdd.n615 gnd 0.007957f
C2951 vdd.n616 gnd 0.009886f
C2952 vdd.n617 gnd 0.007957f
C2953 vdd.n618 gnd 0.009886f
C2954 vdd.t174 gnd 0.505144f
C2955 vdd.n619 gnd 0.009886f
C2956 vdd.n620 gnd 0.007957f
C2957 vdd.n621 gnd 0.009886f
C2958 vdd.n622 gnd 0.007957f
C2959 vdd.n623 gnd 0.009886f
C2960 vdd.t203 gnd 0.505144f
C2961 vdd.n624 gnd 0.631429f
C2962 vdd.n625 gnd 0.009886f
C2963 vdd.n626 gnd 0.007957f
C2964 vdd.n627 gnd 0.009886f
C2965 vdd.n628 gnd 0.007957f
C2966 vdd.n629 gnd 0.009886f
C2967 vdd.t151 gnd 0.505144f
C2968 vdd.n630 gnd 0.009886f
C2969 vdd.n631 gnd 0.007957f
C2970 vdd.n632 gnd 0.009886f
C2971 vdd.n633 gnd 0.007957f
C2972 vdd.n634 gnd 0.009886f
C2973 vdd.n635 gnd 0.70215f
C2974 vdd.n636 gnd 0.838538f
C2975 vdd.t171 gnd 0.505144f
C2976 vdd.n637 gnd 0.009886f
C2977 vdd.n638 gnd 0.007957f
C2978 vdd.n639 gnd 0.009886f
C2979 vdd.n640 gnd 0.007957f
C2980 vdd.n641 gnd 0.009886f
C2981 vdd.n642 gnd 0.530401f
C2982 vdd.n643 gnd 0.009886f
C2983 vdd.n644 gnd 0.007957f
C2984 vdd.n645 gnd 0.009886f
C2985 vdd.n646 gnd 0.007957f
C2986 vdd.n647 gnd 0.009886f
C2987 vdd.n648 gnd 1.01029f
C2988 vdd.t182 gnd 0.505144f
C2989 vdd.n649 gnd 0.009886f
C2990 vdd.n650 gnd 0.007957f
C2991 vdd.n651 gnd 0.009886f
C2992 vdd.n652 gnd 0.007957f
C2993 vdd.n653 gnd 0.009886f
C2994 vdd.t36 gnd 0.505144f
C2995 vdd.n654 gnd 0.009886f
C2996 vdd.n655 gnd 0.007957f
C2997 vdd.n656 gnd 0.022666f
C2998 vdd.n657 gnd 0.022666f
C2999 vdd.n658 gnd 10.496901f
C3000 vdd.n659 gnd 0.560709f
C3001 vdd.n660 gnd 0.022666f
C3002 vdd.n661 gnd 0.008502f
C3003 vdd.n662 gnd 0.007957f
C3004 vdd.n667 gnd 0.006327f
C3005 vdd.n668 gnd 0.007957f
C3006 vdd.n669 gnd 0.009886f
C3007 vdd.n670 gnd 0.009886f
C3008 vdd.n671 gnd 0.009886f
C3009 vdd.n672 gnd 0.009886f
C3010 vdd.n673 gnd 0.009886f
C3011 vdd.n674 gnd 0.007957f
C3012 vdd.n675 gnd 0.009886f
C3013 vdd.n676 gnd 0.009886f
C3014 vdd.n677 gnd 0.009886f
C3015 vdd.n678 gnd 0.009886f
C3016 vdd.n679 gnd 0.009886f
C3017 vdd.n680 gnd 0.007957f
C3018 vdd.n681 gnd 0.009886f
C3019 vdd.n682 gnd 0.009886f
C3020 vdd.n683 gnd 0.009886f
C3021 vdd.n684 gnd 0.009886f
C3022 vdd.n685 gnd 0.009886f
C3023 vdd.t48 gnd 0.121622f
C3024 vdd.t49 gnd 0.12998f
C3025 vdd.t47 gnd 0.158837f
C3026 vdd.n686 gnd 0.203606f
C3027 vdd.n687 gnd 0.171066f
C3028 vdd.n688 gnd 0.016232f
C3029 vdd.n689 gnd 0.009886f
C3030 vdd.n690 gnd 0.009886f
C3031 vdd.n691 gnd 0.009886f
C3032 vdd.n692 gnd 0.009886f
C3033 vdd.n693 gnd 0.009886f
C3034 vdd.n694 gnd 0.007957f
C3035 vdd.n695 gnd 0.009886f
C3036 vdd.n696 gnd 0.009886f
C3037 vdd.n697 gnd 0.009886f
C3038 vdd.n698 gnd 0.009886f
C3039 vdd.n699 gnd 0.009886f
C3040 vdd.n700 gnd 0.007957f
C3041 vdd.n701 gnd 0.009886f
C3042 vdd.n702 gnd 0.009886f
C3043 vdd.n703 gnd 0.009886f
C3044 vdd.n704 gnd 0.009886f
C3045 vdd.n705 gnd 0.009886f
C3046 vdd.n706 gnd 0.007957f
C3047 vdd.n707 gnd 0.009886f
C3048 vdd.n708 gnd 0.009886f
C3049 vdd.n709 gnd 0.009886f
C3050 vdd.n710 gnd 0.009886f
C3051 vdd.n711 gnd 0.009886f
C3052 vdd.n712 gnd 0.007957f
C3053 vdd.n713 gnd 0.009886f
C3054 vdd.n714 gnd 0.009886f
C3055 vdd.n715 gnd 0.009886f
C3056 vdd.n716 gnd 0.009886f
C3057 vdd.n717 gnd 0.009886f
C3058 vdd.n718 gnd 0.007957f
C3059 vdd.n719 gnd 0.009886f
C3060 vdd.n720 gnd 0.009886f
C3061 vdd.n721 gnd 0.009886f
C3062 vdd.n722 gnd 0.007877f
C3063 vdd.t37 gnd 0.121622f
C3064 vdd.t38 gnd 0.12998f
C3065 vdd.t35 gnd 0.158837f
C3066 vdd.n723 gnd 0.203606f
C3067 vdd.n724 gnd 0.171066f
C3068 vdd.n725 gnd 0.009886f
C3069 vdd.n726 gnd 0.007957f
C3070 vdd.n728 gnd 0.009886f
C3071 vdd.n730 gnd 0.009886f
C3072 vdd.n731 gnd 0.009886f
C3073 vdd.n732 gnd 0.007957f
C3074 vdd.n733 gnd 0.009886f
C3075 vdd.n734 gnd 0.009886f
C3076 vdd.n735 gnd 0.009886f
C3077 vdd.n736 gnd 0.009886f
C3078 vdd.n737 gnd 0.009886f
C3079 vdd.n738 gnd 0.007957f
C3080 vdd.n739 gnd 0.009886f
C3081 vdd.n740 gnd 0.009886f
C3082 vdd.n741 gnd 0.009886f
C3083 vdd.n742 gnd 0.009886f
C3084 vdd.n743 gnd 0.009886f
C3085 vdd.n744 gnd 0.007957f
C3086 vdd.n745 gnd 0.009886f
C3087 vdd.n746 gnd 0.009886f
C3088 vdd.n747 gnd 0.009886f
C3089 vdd.n748 gnd 0.006327f
C3090 vdd.n753 gnd 0.006722f
C3091 vdd.n754 gnd 0.006722f
C3092 vdd.n755 gnd 0.006722f
C3093 vdd.n756 gnd 10.274599f
C3094 vdd.n757 gnd 0.006722f
C3095 vdd.n758 gnd 0.006722f
C3096 vdd.n759 gnd 0.006722f
C3097 vdd.n761 gnd 0.006722f
C3098 vdd.n762 gnd 0.006722f
C3099 vdd.n764 gnd 0.006722f
C3100 vdd.n765 gnd 0.004893f
C3101 vdd.n767 gnd 0.006722f
C3102 vdd.t42 gnd 0.27165f
C3103 vdd.t41 gnd 0.278068f
C3104 vdd.t39 gnd 0.177344f
C3105 vdd.n768 gnd 0.095845f
C3106 vdd.n769 gnd 0.054366f
C3107 vdd.n770 gnd 0.009607f
C3108 vdd.n771 gnd 0.015411f
C3109 vdd.n773 gnd 0.006722f
C3110 vdd.n774 gnd 0.686995f
C3111 vdd.n775 gnd 0.014559f
C3112 vdd.n776 gnd 0.014559f
C3113 vdd.n777 gnd 0.006722f
C3114 vdd.n778 gnd 0.015494f
C3115 vdd.n779 gnd 0.006722f
C3116 vdd.n780 gnd 0.006722f
C3117 vdd.n781 gnd 0.006722f
C3118 vdd.n782 gnd 0.006722f
C3119 vdd.n783 gnd 0.006722f
C3120 vdd.n785 gnd 0.006722f
C3121 vdd.n786 gnd 0.006722f
C3122 vdd.n788 gnd 0.006722f
C3123 vdd.n789 gnd 0.006722f
C3124 vdd.n791 gnd 0.006722f
C3125 vdd.n792 gnd 0.006722f
C3126 vdd.n794 gnd 0.006722f
C3127 vdd.n795 gnd 0.006722f
C3128 vdd.n797 gnd 0.006722f
C3129 vdd.n798 gnd 0.006722f
C3130 vdd.n800 gnd 0.006722f
C3131 vdd.n801 gnd 0.004893f
C3132 vdd.n803 gnd 0.006722f
C3133 vdd.t77 gnd 0.27165f
C3134 vdd.t76 gnd 0.278068f
C3135 vdd.t75 gnd 0.177344f
C3136 vdd.n804 gnd 0.095845f
C3137 vdd.n805 gnd 0.054366f
C3138 vdd.n806 gnd 0.009607f
C3139 vdd.n807 gnd 0.006722f
C3140 vdd.n808 gnd 0.006722f
C3141 vdd.t40 gnd 0.343498f
C3142 vdd.n809 gnd 0.006722f
C3143 vdd.n810 gnd 0.006722f
C3144 vdd.n811 gnd 0.006722f
C3145 vdd.n812 gnd 0.006722f
C3146 vdd.n813 gnd 0.006722f
C3147 vdd.n814 gnd 0.686995f
C3148 vdd.n815 gnd 0.006722f
C3149 vdd.n816 gnd 0.006722f
C3150 vdd.n817 gnd 0.560709f
C3151 vdd.n818 gnd 0.006722f
C3152 vdd.n819 gnd 0.006722f
C3153 vdd.n820 gnd 0.006722f
C3154 vdd.n821 gnd 0.006722f
C3155 vdd.n822 gnd 0.686995f
C3156 vdd.n823 gnd 0.006722f
C3157 vdd.n824 gnd 0.006722f
C3158 vdd.n825 gnd 0.006722f
C3159 vdd.n826 gnd 0.006722f
C3160 vdd.n827 gnd 0.006722f
C3161 vdd.t28 gnd 0.343498f
C3162 vdd.n828 gnd 0.006722f
C3163 vdd.n829 gnd 0.006722f
C3164 vdd.n830 gnd 0.006722f
C3165 vdd.n831 gnd 0.006722f
C3166 vdd.n832 gnd 0.006722f
C3167 vdd.t7 gnd 0.343498f
C3168 vdd.n833 gnd 0.006722f
C3169 vdd.n834 gnd 0.006722f
C3170 vdd.n835 gnd 0.681944f
C3171 vdd.n836 gnd 0.006722f
C3172 vdd.n837 gnd 0.006722f
C3173 vdd.n838 gnd 0.006722f
C3174 vdd.t3 gnd 0.343498f
C3175 vdd.n839 gnd 0.006722f
C3176 vdd.n840 gnd 0.006722f
C3177 vdd.n841 gnd 0.530401f
C3178 vdd.n842 gnd 0.006722f
C3179 vdd.n843 gnd 0.006722f
C3180 vdd.n844 gnd 0.006722f
C3181 vdd.n845 gnd 0.459681f
C3182 vdd.n846 gnd 0.006722f
C3183 vdd.n847 gnd 0.006722f
C3184 vdd.n848 gnd 0.378858f
C3185 vdd.n849 gnd 0.006722f
C3186 vdd.n850 gnd 0.006722f
C3187 vdd.n851 gnd 0.006722f
C3188 vdd.n852 gnd 0.565761f
C3189 vdd.n853 gnd 0.006722f
C3190 vdd.n854 gnd 0.006722f
C3191 vdd.t0 gnd 0.343498f
C3192 vdd.n855 gnd 0.006722f
C3193 vdd.t56 gnd 0.278068f
C3194 vdd.t54 gnd 0.177344f
C3195 vdd.t57 gnd 0.278068f
C3196 vdd.n856 gnd 0.156286f
C3197 vdd.n857 gnd 0.006722f
C3198 vdd.n858 gnd 0.006722f
C3199 vdd.n859 gnd 0.686995f
C3200 vdd.n860 gnd 0.006722f
C3201 vdd.n861 gnd 0.006722f
C3202 vdd.t55 gnd 0.267726f
C3203 vdd.t13 gnd 0.121234f
C3204 vdd.n862 gnd 0.006722f
C3205 vdd.n863 gnd 0.006722f
C3206 vdd.n864 gnd 0.006722f
C3207 vdd.t113 gnd 0.343498f
C3208 vdd.n865 gnd 0.006722f
C3209 vdd.n866 gnd 0.006722f
C3210 vdd.n867 gnd 0.006722f
C3211 vdd.n868 gnd 0.006722f
C3212 vdd.n869 gnd 0.006722f
C3213 vdd.t118 gnd 0.343498f
C3214 vdd.n870 gnd 0.006722f
C3215 vdd.n871 gnd 0.006722f
C3216 vdd.n872 gnd 0.611224f
C3217 vdd.n873 gnd 0.006722f
C3218 vdd.n874 gnd 0.006722f
C3219 vdd.n875 gnd 0.006722f
C3220 vdd.n876 gnd 0.378858f
C3221 vdd.n877 gnd 0.006722f
C3222 vdd.n878 gnd 0.006722f
C3223 vdd.t16 gnd 0.343498f
C3224 vdd.n879 gnd 0.006722f
C3225 vdd.n880 gnd 0.006722f
C3226 vdd.n881 gnd 0.006722f
C3227 vdd.n882 gnd 0.530401f
C3228 vdd.n883 gnd 0.006722f
C3229 vdd.n884 gnd 0.006722f
C3230 vdd.t29 gnd 0.252572f
C3231 vdd.t21 gnd 0.308138f
C3232 vdd.n885 gnd 0.006722f
C3233 vdd.n886 gnd 0.006722f
C3234 vdd.n887 gnd 0.006722f
C3235 vdd.t264 gnd 0.343498f
C3236 vdd.n888 gnd 0.006722f
C3237 vdd.n889 gnd 0.006722f
C3238 vdd.t9 gnd 0.343498f
C3239 vdd.n890 gnd 0.006722f
C3240 vdd.n891 gnd 0.006722f
C3241 vdd.n892 gnd 0.006722f
C3242 vdd.t268 gnd 0.343498f
C3243 vdd.n893 gnd 0.006722f
C3244 vdd.n894 gnd 0.006722f
C3245 vdd.t18 gnd 0.343498f
C3246 vdd.n895 gnd 0.006722f
C3247 vdd.n896 gnd 0.006722f
C3248 vdd.n897 gnd 0.006722f
C3249 vdd.n898 gnd 0.686995f
C3250 vdd.n899 gnd 0.006722f
C3251 vdd.n900 gnd 0.006722f
C3252 vdd.n901 gnd 0.474835f
C3253 vdd.n902 gnd 0.006722f
C3254 vdd.n903 gnd 0.006722f
C3255 vdd.n904 gnd 0.006722f
C3256 vdd.t1 gnd 0.343498f
C3257 vdd.n905 gnd 0.006722f
C3258 vdd.n906 gnd 0.006722f
C3259 vdd.n907 gnd 0.006722f
C3260 vdd.n908 gnd 0.006722f
C3261 vdd.n909 gnd 0.006722f
C3262 vdd.t114 gnd 0.343498f
C3263 vdd.n910 gnd 0.006722f
C3264 vdd.n911 gnd 0.006722f
C3265 vdd.t86 gnd 0.343498f
C3266 vdd.n912 gnd 0.006722f
C3267 vdd.n913 gnd 0.015494f
C3268 vdd.n914 gnd 0.015494f
C3269 vdd.t116 gnd 0.606172f
C3270 vdd.n915 gnd 0.014559f
C3271 vdd.n916 gnd 0.014559f
C3272 vdd.n917 gnd 0.383909f
C3273 vdd.n918 gnd 0.015494f
C3274 vdd.n919 gnd 0.006722f
C3275 vdd.n920 gnd 0.006722f
C3276 vdd.t260 gnd 0.606172f
C3277 vdd.n938 gnd 0.015494f
C3278 vdd.n956 gnd 0.014559f
C3279 vdd.n957 gnd 0.006722f
C3280 vdd.n958 gnd 0.014559f
C3281 vdd.t107 gnd 0.27165f
C3282 vdd.t106 gnd 0.278068f
C3283 vdd.t105 gnd 0.177344f
C3284 vdd.n959 gnd 0.095845f
C3285 vdd.n960 gnd 0.054366f
C3286 vdd.n961 gnd 0.015411f
C3287 vdd.n962 gnd 0.006722f
C3288 vdd.n963 gnd 0.383909f
C3289 vdd.n964 gnd 0.014559f
C3290 vdd.n965 gnd 0.006722f
C3291 vdd.n966 gnd 0.015494f
C3292 vdd.n967 gnd 0.006722f
C3293 vdd.t84 gnd 0.27165f
C3294 vdd.t83 gnd 0.278068f
C3295 vdd.t81 gnd 0.177344f
C3296 vdd.n968 gnd 0.095845f
C3297 vdd.n969 gnd 0.054366f
C3298 vdd.n970 gnd 0.009607f
C3299 vdd.n971 gnd 0.006722f
C3300 vdd.n972 gnd 0.006722f
C3301 vdd.t82 gnd 0.343498f
C3302 vdd.n973 gnd 0.006722f
C3303 vdd.t258 gnd 0.343498f
C3304 vdd.n974 gnd 0.006722f
C3305 vdd.n975 gnd 0.006722f
C3306 vdd.n976 gnd 0.006722f
C3307 vdd.n977 gnd 0.006722f
C3308 vdd.n978 gnd 0.006722f
C3309 vdd.n979 gnd 0.686995f
C3310 vdd.n980 gnd 0.006722f
C3311 vdd.n981 gnd 0.006722f
C3312 vdd.t14 gnd 0.343498f
C3313 vdd.n982 gnd 0.006722f
C3314 vdd.n983 gnd 0.006722f
C3315 vdd.n984 gnd 0.006722f
C3316 vdd.n985 gnd 0.006722f
C3317 vdd.n986 gnd 0.474835f
C3318 vdd.n987 gnd 0.006722f
C3319 vdd.n988 gnd 0.006722f
C3320 vdd.n989 gnd 0.006722f
C3321 vdd.n990 gnd 0.006722f
C3322 vdd.n991 gnd 0.006722f
C3323 vdd.t4 gnd 0.343498f
C3324 vdd.n992 gnd 0.006722f
C3325 vdd.n993 gnd 0.006722f
C3326 vdd.t5 gnd 0.343498f
C3327 vdd.n994 gnd 0.006722f
C3328 vdd.n995 gnd 0.006722f
C3329 vdd.n996 gnd 0.006722f
C3330 vdd.t26 gnd 0.343498f
C3331 vdd.n997 gnd 0.006722f
C3332 vdd.n998 gnd 0.006722f
C3333 vdd.t262 gnd 0.343498f
C3334 vdd.n999 gnd 0.006722f
C3335 vdd.n1000 gnd 0.006722f
C3336 vdd.n1001 gnd 0.006722f
C3337 vdd.t270 gnd 0.308138f
C3338 vdd.n1002 gnd 0.006722f
C3339 vdd.n1003 gnd 0.006722f
C3340 vdd.n1004 gnd 0.530401f
C3341 vdd.n1005 gnd 0.006722f
C3342 vdd.n1006 gnd 0.006722f
C3343 vdd.n1007 gnd 0.006722f
C3344 vdd.t266 gnd 0.343498f
C3345 vdd.n1008 gnd 0.006722f
C3346 vdd.n1009 gnd 0.006722f
C3347 vdd.t8 gnd 0.252572f
C3348 vdd.n1010 gnd 0.378858f
C3349 vdd.n1011 gnd 0.006722f
C3350 vdd.n1012 gnd 0.006722f
C3351 vdd.n1013 gnd 0.006722f
C3352 vdd.n1014 gnd 0.611224f
C3353 vdd.n1015 gnd 0.006722f
C3354 vdd.n1016 gnd 0.006722f
C3355 vdd.t23 gnd 0.343498f
C3356 vdd.n1017 gnd 0.006722f
C3357 vdd.n1018 gnd 0.006722f
C3358 vdd.n1019 gnd 0.006722f
C3359 vdd.n1020 gnd 0.686995f
C3360 vdd.n1021 gnd 0.006722f
C3361 vdd.n1022 gnd 0.006722f
C3362 vdd.t30 gnd 0.343498f
C3363 vdd.n1023 gnd 0.006722f
C3364 vdd.n1024 gnd 0.006722f
C3365 vdd.n1025 gnd 0.006722f
C3366 vdd.t31 gnd 0.121234f
C3367 vdd.n1026 gnd 0.006722f
C3368 vdd.n1027 gnd 0.006722f
C3369 vdd.n1028 gnd 0.006722f
C3370 vdd.t97 gnd 0.278068f
C3371 vdd.t95 gnd 0.177344f
C3372 vdd.t98 gnd 0.278068f
C3373 vdd.n1029 gnd 0.156286f
C3374 vdd.n1030 gnd 0.006722f
C3375 vdd.n1031 gnd 0.006722f
C3376 vdd.t27 gnd 0.343498f
C3377 vdd.n1032 gnd 0.006722f
C3378 vdd.n1033 gnd 0.006722f
C3379 vdd.t96 gnd 0.267726f
C3380 vdd.n1034 gnd 0.565761f
C3381 vdd.n1035 gnd 0.006722f
C3382 vdd.n1036 gnd 0.006722f
C3383 vdd.n1037 gnd 0.006722f
C3384 vdd.n1038 gnd 0.378858f
C3385 vdd.n1039 gnd 0.006722f
C3386 vdd.n1040 gnd 0.006722f
C3387 vdd.n1041 gnd 0.459681f
C3388 vdd.n1042 gnd 0.006722f
C3389 vdd.n1043 gnd 0.006722f
C3390 vdd.n1044 gnd 0.006722f
C3391 vdd.n1045 gnd 0.530401f
C3392 vdd.n1046 gnd 0.006722f
C3393 vdd.n1047 gnd 0.006722f
C3394 vdd.t19 gnd 0.343498f
C3395 vdd.n1048 gnd 0.006722f
C3396 vdd.n1049 gnd 0.006722f
C3397 vdd.n1050 gnd 0.006722f
C3398 vdd.n1051 gnd 0.681944f
C3399 vdd.n1052 gnd 0.006722f
C3400 vdd.n1053 gnd 0.006722f
C3401 vdd.t34 gnd 0.343498f
C3402 vdd.n1054 gnd 0.006722f
C3403 vdd.n1055 gnd 0.006722f
C3404 vdd.n1056 gnd 0.006722f
C3405 vdd.n1057 gnd 0.686995f
C3406 vdd.n1058 gnd 0.006722f
C3407 vdd.n1059 gnd 0.006722f
C3408 vdd.t20 gnd 0.343498f
C3409 vdd.n1060 gnd 0.006722f
C3410 vdd.n1061 gnd 0.006722f
C3411 vdd.n1062 gnd 0.006722f
C3412 vdd.n1063 gnd 0.686995f
C3413 vdd.n1064 gnd 0.006722f
C3414 vdd.n1065 gnd 0.006722f
C3415 vdd.n1066 gnd 0.006722f
C3416 vdd.n1067 gnd 0.006722f
C3417 vdd.n1068 gnd 0.006722f
C3418 vdd.n1069 gnd 0.560709f
C3419 vdd.n1070 gnd 0.006722f
C3420 vdd.n1071 gnd 0.006722f
C3421 vdd.n1072 gnd 0.006722f
C3422 vdd.n1073 gnd 0.006722f
C3423 vdd.n1074 gnd 0.006722f
C3424 vdd.n1075 gnd 0.686995f
C3425 vdd.n1076 gnd 0.006722f
C3426 vdd.n1077 gnd 0.006722f
C3427 vdd.t44 gnd 0.343498f
C3428 vdd.n1078 gnd 0.006722f
C3429 vdd.n1079 gnd 0.015494f
C3430 vdd.n1080 gnd 0.015494f
C3431 vdd.n1081 gnd 10.274599f
C3432 vdd.n1082 gnd 0.014559f
C3433 vdd.n1083 gnd 0.014559f
C3434 vdd.n1084 gnd 0.015494f
C3435 vdd.n1085 gnd 0.006722f
C3436 vdd.n1087 gnd 0.006722f
C3437 vdd.n1088 gnd 0.006722f
C3438 vdd.n1089 gnd 0.006722f
C3439 vdd.n1090 gnd 0.006722f
C3440 vdd.n1091 gnd 0.006722f
C3441 vdd.n1092 gnd 0.006722f
C3442 vdd.n1093 gnd 0.03537f
C3443 vdd.n1094 gnd 0.006722f
C3444 vdd.n1095 gnd 0.006722f
C3445 vdd.n1096 gnd 0.006722f
C3446 vdd.n1097 gnd 0.006722f
C3447 vdd.n1098 gnd 0.006722f
C3448 vdd.n1099 gnd 0.006722f
C3449 vdd.n1100 gnd 0.006722f
C3450 vdd.t109 gnd 0.27165f
C3451 vdd.t110 gnd 0.278068f
C3452 vdd.t108 gnd 0.177344f
C3453 vdd.n1101 gnd 0.095845f
C3454 vdd.n1102 gnd 0.054366f
C3455 vdd.n1103 gnd 0.006722f
C3456 vdd.n1104 gnd 0.006722f
C3457 vdd.n1105 gnd 0.006722f
C3458 vdd.n1106 gnd 0.006722f
C3459 vdd.t45 gnd 0.27165f
C3460 vdd.t46 gnd 0.278068f
C3461 vdd.t43 gnd 0.177344f
C3462 vdd.n1107 gnd 0.095845f
C3463 vdd.n1108 gnd 0.054366f
C3464 vdd.n1109 gnd 0.006722f
C3465 vdd.n1110 gnd 0.006722f
C3466 vdd.n1111 gnd 0.006722f
C3467 vdd.n1112 gnd 0.006722f
C3468 vdd.n1113 gnd 0.006722f
C3469 vdd.n1114 gnd 0.006722f
C3470 vdd.n1115 gnd 0.006327f
C3471 vdd.n1118 gnd 0.022666f
C3472 vdd.n1119 gnd 0.007957f
C3473 vdd.n1120 gnd 0.009886f
C3474 vdd.n1122 gnd 0.009886f
C3475 vdd.n1123 gnd 0.006604f
C3476 vdd.n1124 gnd 0.560709f
C3477 vdd.n1125 gnd 10.496901f
C3478 vdd.n1126 gnd 0.009886f
C3479 vdd.n1127 gnd 0.022666f
C3480 vdd.n1128 gnd 0.007957f
C3481 vdd.n1129 gnd 0.009886f
C3482 vdd.n1130 gnd 0.007957f
C3483 vdd.n1131 gnd 0.009886f
C3484 vdd.n1132 gnd 1.01029f
C3485 vdd.n1133 gnd 0.009886f
C3486 vdd.n1134 gnd 0.007957f
C3487 vdd.n1135 gnd 0.007957f
C3488 vdd.n1136 gnd 0.009886f
C3489 vdd.n1137 gnd 0.007957f
C3490 vdd.n1138 gnd 0.009886f
C3491 vdd.t214 gnd 0.505144f
C3492 vdd.n1139 gnd 0.009886f
C3493 vdd.n1140 gnd 0.007957f
C3494 vdd.n1141 gnd 0.009886f
C3495 vdd.n1142 gnd 0.007957f
C3496 vdd.n1143 gnd 0.009886f
C3497 vdd.t142 gnd 0.505144f
C3498 vdd.n1144 gnd 0.009886f
C3499 vdd.n1145 gnd 0.007957f
C3500 vdd.n1146 gnd 0.009886f
C3501 vdd.n1147 gnd 0.007957f
C3502 vdd.n1148 gnd 0.009886f
C3503 vdd.t186 gnd 0.505144f
C3504 vdd.n1149 gnd 0.70215f
C3505 vdd.n1150 gnd 0.009886f
C3506 vdd.n1151 gnd 0.007957f
C3507 vdd.n1152 gnd 0.009886f
C3508 vdd.n1153 gnd 0.007957f
C3509 vdd.n1154 gnd 0.009886f
C3510 vdd.n1155 gnd 0.803178f
C3511 vdd.n1156 gnd 0.009886f
C3512 vdd.n1157 gnd 0.007957f
C3513 vdd.n1158 gnd 0.009886f
C3514 vdd.n1159 gnd 0.007957f
C3515 vdd.n1160 gnd 0.009886f
C3516 vdd.n1161 gnd 0.631429f
C3517 vdd.t167 gnd 0.505144f
C3518 vdd.n1162 gnd 0.009886f
C3519 vdd.n1163 gnd 0.007957f
C3520 vdd.n1164 gnd 0.009886f
C3521 vdd.n1165 gnd 0.007957f
C3522 vdd.n1166 gnd 0.009886f
C3523 vdd.t212 gnd 0.505144f
C3524 vdd.n1167 gnd 0.009886f
C3525 vdd.n1168 gnd 0.007957f
C3526 vdd.n1169 gnd 0.009886f
C3527 vdd.n1170 gnd 0.007957f
C3528 vdd.n1171 gnd 0.009886f
C3529 vdd.t140 gnd 0.505144f
C3530 vdd.n1172 gnd 0.550607f
C3531 vdd.n1173 gnd 0.009886f
C3532 vdd.n1174 gnd 0.007957f
C3533 vdd.n1175 gnd 0.009886f
C3534 vdd.n1176 gnd 0.007957f
C3535 vdd.n1177 gnd 0.009886f
C3536 vdd.t160 gnd 0.505144f
C3537 vdd.n1178 gnd 0.009886f
C3538 vdd.n1179 gnd 0.007957f
C3539 vdd.n1180 gnd 0.009886f
C3540 vdd.n1181 gnd 0.007957f
C3541 vdd.n1182 gnd 0.009886f
C3542 vdd.n1183 gnd 0.782973f
C3543 vdd.n1184 gnd 0.838538f
C3544 vdd.t165 gnd 0.505144f
C3545 vdd.n1185 gnd 0.009886f
C3546 vdd.n1186 gnd 0.007957f
C3547 vdd.n1187 gnd 0.009886f
C3548 vdd.n1188 gnd 0.007957f
C3549 vdd.n1189 gnd 0.009886f
C3550 vdd.n1190 gnd 0.611224f
C3551 vdd.n1191 gnd 0.009886f
C3552 vdd.n1192 gnd 0.007957f
C3553 vdd.n1193 gnd 0.009886f
C3554 vdd.n1194 gnd 0.007957f
C3555 vdd.n1195 gnd 0.009886f
C3556 vdd.t188 gnd 0.505144f
C3557 vdd.t136 gnd 0.505144f
C3558 vdd.n1196 gnd 0.009886f
C3559 vdd.n1197 gnd 0.007957f
C3560 vdd.n1198 gnd 0.009886f
C3561 vdd.n1199 gnd 0.007957f
C3562 vdd.n1200 gnd 0.009886f
C3563 vdd.t208 gnd 0.505144f
C3564 vdd.n1201 gnd 0.009886f
C3565 vdd.n1202 gnd 0.007957f
C3566 vdd.n1203 gnd 0.009886f
C3567 vdd.n1204 gnd 0.007957f
C3568 vdd.n1205 gnd 0.009886f
C3569 vdd.t130 gnd 0.505144f
C3570 vdd.n1206 gnd 0.742561f
C3571 vdd.n1207 gnd 0.009886f
C3572 vdd.n1208 gnd 0.007957f
C3573 vdd.n1209 gnd 0.009886f
C3574 vdd.n1210 gnd 0.007957f
C3575 vdd.n1211 gnd 0.009886f
C3576 vdd.n1212 gnd 1.01029f
C3577 vdd.n1213 gnd 0.009886f
C3578 vdd.n1214 gnd 0.007957f
C3579 vdd.n1215 gnd 0.009886f
C3580 vdd.n1216 gnd 0.007957f
C3581 vdd.n1217 gnd 0.009886f
C3582 vdd.n1218 gnd 0.853693f
C3583 vdd.n1219 gnd 0.009886f
C3584 vdd.n1220 gnd 0.007957f
C3585 vdd.n1221 gnd 0.022512f
C3586 vdd.n1222 gnd 0.006604f
C3587 vdd.n1223 gnd 0.022512f
C3588 vdd.n1224 gnd 1.33358f
C3589 vdd.n1225 gnd 0.022512f
C3590 vdd.n1226 gnd 0.006604f
C3591 vdd.n1227 gnd 0.009886f
C3592 vdd.t70 gnd 0.121622f
C3593 vdd.t71 gnd 0.12998f
C3594 vdd.t68 gnd 0.158837f
C3595 vdd.n1228 gnd 0.203606f
C3596 vdd.n1229 gnd 0.171862f
C3597 vdd.n1230 gnd 0.013049f
C3598 vdd.n1231 gnd 0.009886f
C3599 vdd.n1262 gnd 0.009886f
C3600 vdd.n1263 gnd 0.009886f
C3601 vdd.n1264 gnd 0.022666f
C3602 vdd.n1265 gnd 0.007957f
C3603 vdd.n1266 gnd 0.009886f
C3604 vdd.n1267 gnd 0.009886f
C3605 vdd.n1268 gnd 0.009886f
C3606 vdd.n1269 gnd 0.009886f
C3607 vdd.n1270 gnd 0.007957f
C3608 vdd.n1271 gnd 0.009886f
C3609 vdd.n1272 gnd 0.009886f
C3610 vdd.n1273 gnd 0.009886f
C3611 vdd.n1274 gnd 0.009886f
C3612 vdd.n1275 gnd 0.009886f
C3613 vdd.n1276 gnd 0.007957f
C3614 vdd.n1277 gnd 0.009886f
C3615 vdd.n1278 gnd 0.009886f
C3616 vdd.n1279 gnd 0.009886f
C3617 vdd.n1280 gnd 0.009886f
C3618 vdd.n1281 gnd 0.009886f
C3619 vdd.n1282 gnd 0.007957f
C3620 vdd.n1283 gnd 0.009886f
C3621 vdd.n1284 gnd 0.009886f
C3622 vdd.n1285 gnd 0.009886f
C3623 vdd.n1286 gnd 0.009886f
C3624 vdd.n1287 gnd 0.009886f
C3625 vdd.n1288 gnd 0.006644f
C3626 vdd.n1289 gnd 0.009886f
C3627 vdd.n1290 gnd 0.009886f
C3628 vdd.n1291 gnd 0.009886f
C3629 vdd.n1292 gnd 0.007957f
C3630 vdd.n1293 gnd 0.009886f
C3631 vdd.n1294 gnd 0.009886f
C3632 vdd.n1295 gnd 0.009886f
C3633 vdd.n1296 gnd 0.009886f
C3634 vdd.n1297 gnd 0.009886f
C3635 vdd.n1298 gnd 0.007957f
C3636 vdd.n1299 gnd 0.009886f
C3637 vdd.n1300 gnd 0.009886f
C3638 vdd.n1301 gnd 0.009886f
C3639 vdd.n1302 gnd 0.009886f
C3640 vdd.n1303 gnd 0.009886f
C3641 vdd.n1304 gnd 0.007957f
C3642 vdd.n1305 gnd 0.009886f
C3643 vdd.n1306 gnd 0.009886f
C3644 vdd.n1307 gnd 0.009886f
C3645 vdd.n1308 gnd 0.009886f
C3646 vdd.n1309 gnd 0.009886f
C3647 vdd.n1310 gnd 0.007957f
C3648 vdd.n1311 gnd 0.009886f
C3649 vdd.n1312 gnd 0.009886f
C3650 vdd.n1313 gnd 0.009886f
C3651 vdd.n1314 gnd 0.009886f
C3652 vdd.n1315 gnd 0.009886f
C3653 vdd.n1316 gnd 0.007957f
C3654 vdd.n1317 gnd 0.009886f
C3655 vdd.n1318 gnd 0.009886f
C3656 vdd.n1319 gnd 0.009886f
C3657 vdd.n1320 gnd 0.009886f
C3658 vdd.n1321 gnd 0.007877f
C3659 vdd.n1322 gnd 0.009886f
C3660 vdd.n1323 gnd 0.009886f
C3661 vdd.n1324 gnd 0.009886f
C3662 vdd.n1325 gnd 0.009886f
C3663 vdd.n1326 gnd 0.009886f
C3664 vdd.n1327 gnd 0.007957f
C3665 vdd.n1328 gnd 0.009886f
C3666 vdd.n1329 gnd 0.009886f
C3667 vdd.n1330 gnd 0.009886f
C3668 vdd.n1331 gnd 0.009886f
C3669 vdd.n1332 gnd 0.009886f
C3670 vdd.n1333 gnd 0.007957f
C3671 vdd.n1334 gnd 0.009886f
C3672 vdd.n1335 gnd 0.009886f
C3673 vdd.n1336 gnd 0.009886f
C3674 vdd.n1337 gnd 0.009886f
C3675 vdd.n1338 gnd 0.009886f
C3676 vdd.n1339 gnd 0.007957f
C3677 vdd.n1340 gnd 0.009886f
C3678 vdd.n1341 gnd 0.009886f
C3679 vdd.n1342 gnd 0.009886f
C3680 vdd.n1343 gnd 0.009886f
C3681 vdd.n1344 gnd 0.009886f
C3682 vdd.n1345 gnd 0.007957f
C3683 vdd.n1346 gnd 0.009886f
C3684 vdd.n1347 gnd 0.009886f
C3685 vdd.n1348 gnd 0.009886f
C3686 vdd.n1349 gnd 0.009886f
C3687 vdd.n1350 gnd 0.009886f
C3688 vdd.n1351 gnd 0.004177f
C3689 vdd.n1352 gnd 0.009886f
C3690 vdd.n1353 gnd 0.007957f
C3691 vdd.n1354 gnd 0.007957f
C3692 vdd.n1355 gnd 0.007957f
C3693 vdd.n1356 gnd 0.009886f
C3694 vdd.n1357 gnd 0.009886f
C3695 vdd.n1358 gnd 0.009886f
C3696 vdd.n1359 gnd 0.007957f
C3697 vdd.n1360 gnd 0.007957f
C3698 vdd.n1361 gnd 0.007957f
C3699 vdd.n1362 gnd 0.009886f
C3700 vdd.n1363 gnd 0.009886f
C3701 vdd.n1364 gnd 0.009886f
C3702 vdd.n1365 gnd 0.007957f
C3703 vdd.n1366 gnd 0.007957f
C3704 vdd.n1367 gnd 0.007957f
C3705 vdd.n1368 gnd 0.009886f
C3706 vdd.n1369 gnd 0.009886f
C3707 vdd.n1370 gnd 0.009886f
C3708 vdd.n1371 gnd 0.007957f
C3709 vdd.n1372 gnd 0.007957f
C3710 vdd.n1373 gnd 0.007957f
C3711 vdd.n1374 gnd 0.009886f
C3712 vdd.n1375 gnd 0.009886f
C3713 vdd.n1376 gnd 0.009886f
C3714 vdd.n1377 gnd 0.007957f
C3715 vdd.n1378 gnd 0.007957f
C3716 vdd.n1379 gnd 0.007957f
C3717 vdd.n1380 gnd 0.009886f
C3718 vdd.n1381 gnd 0.009886f
C3719 vdd.n1382 gnd 0.009886f
C3720 vdd.n1383 gnd 0.009886f
C3721 vdd.t93 gnd 0.121622f
C3722 vdd.t94 gnd 0.12998f
C3723 vdd.t92 gnd 0.158837f
C3724 vdd.n1384 gnd 0.203606f
C3725 vdd.n1385 gnd 0.171862f
C3726 vdd.n1386 gnd 0.017028f
C3727 vdd.n1387 gnd 0.005411f
C3728 vdd.n1388 gnd 0.007957f
C3729 vdd.n1389 gnd 0.009886f
C3730 vdd.n1390 gnd 0.009886f
C3731 vdd.n1391 gnd 0.009886f
C3732 vdd.n1392 gnd 0.007957f
C3733 vdd.n1393 gnd 0.007957f
C3734 vdd.n1394 gnd 0.007957f
C3735 vdd.n1395 gnd 0.009886f
C3736 vdd.n1396 gnd 0.009886f
C3737 vdd.n1397 gnd 0.009886f
C3738 vdd.n1398 gnd 0.007957f
C3739 vdd.n1399 gnd 0.007957f
C3740 vdd.n1400 gnd 0.007957f
C3741 vdd.n1401 gnd 0.009886f
C3742 vdd.n1402 gnd 0.009886f
C3743 vdd.n1403 gnd 0.009886f
C3744 vdd.n1404 gnd 0.007957f
C3745 vdd.n1405 gnd 0.007957f
C3746 vdd.n1406 gnd 0.007957f
C3747 vdd.n1407 gnd 0.009886f
C3748 vdd.n1408 gnd 0.009886f
C3749 vdd.n1409 gnd 0.009886f
C3750 vdd.n1410 gnd 0.007957f
C3751 vdd.n1411 gnd 0.007957f
C3752 vdd.n1412 gnd 0.007957f
C3753 vdd.n1413 gnd 0.009886f
C3754 vdd.n1414 gnd 0.009886f
C3755 vdd.n1415 gnd 0.009886f
C3756 vdd.n1416 gnd 0.007957f
C3757 vdd.n1417 gnd 0.006644f
C3758 vdd.n1418 gnd 0.009886f
C3759 vdd.n1419 gnd 0.009886f
C3760 vdd.t103 gnd 0.121622f
C3761 vdd.t104 gnd 0.12998f
C3762 vdd.t102 gnd 0.158837f
C3763 vdd.n1420 gnd 0.203606f
C3764 vdd.n1421 gnd 0.171862f
C3765 vdd.n1422 gnd 0.017028f
C3766 vdd.n1423 gnd 0.009886f
C3767 vdd.n1424 gnd 0.009886f
C3768 vdd.n1425 gnd 0.009886f
C3769 vdd.n1426 gnd 0.007957f
C3770 vdd.n1427 gnd 0.007957f
C3771 vdd.n1428 gnd 0.007957f
C3772 vdd.n1429 gnd 0.009886f
C3773 vdd.n1430 gnd 0.009886f
C3774 vdd.n1431 gnd 0.009886f
C3775 vdd.n1432 gnd 0.007957f
C3776 vdd.n1433 gnd 0.007957f
C3777 vdd.n1434 gnd 0.007957f
C3778 vdd.n1435 gnd 0.009886f
C3779 vdd.n1436 gnd 0.009886f
C3780 vdd.n1437 gnd 0.009886f
C3781 vdd.n1438 gnd 0.007957f
C3782 vdd.n1439 gnd 0.007957f
C3783 vdd.n1440 gnd 0.007957f
C3784 vdd.n1441 gnd 0.009886f
C3785 vdd.n1442 gnd 0.009886f
C3786 vdd.n1443 gnd 0.009886f
C3787 vdd.n1444 gnd 0.007957f
C3788 vdd.n1445 gnd 0.007957f
C3789 vdd.n1446 gnd 0.007957f
C3790 vdd.n1447 gnd 0.009886f
C3791 vdd.n1448 gnd 0.009886f
C3792 vdd.n1449 gnd 0.009886f
C3793 vdd.n1450 gnd 0.007957f
C3794 vdd.n1451 gnd 0.006604f
C3795 vdd.n1452 gnd 0.022666f
C3796 vdd.n1454 gnd 2.23273f
C3797 vdd.n1455 gnd 0.022666f
C3798 vdd.n1456 gnd 0.00378f
C3799 vdd.n1457 gnd 0.022666f
C3800 vdd.n1458 gnd 0.022512f
C3801 vdd.n1459 gnd 0.009886f
C3802 vdd.n1460 gnd 0.007957f
C3803 vdd.n1461 gnd 0.009886f
C3804 vdd.t69 gnd 0.505144f
C3805 vdd.n1462 gnd 0.661738f
C3806 vdd.n1463 gnd 0.009886f
C3807 vdd.n1464 gnd 0.007957f
C3808 vdd.n1465 gnd 0.009886f
C3809 vdd.n1466 gnd 0.009886f
C3810 vdd.n1467 gnd 0.009886f
C3811 vdd.n1468 gnd 0.007957f
C3812 vdd.n1469 gnd 0.009886f
C3813 vdd.n1470 gnd 1.01029f
C3814 vdd.n1471 gnd 0.009886f
C3815 vdd.n1472 gnd 0.007957f
C3816 vdd.n1473 gnd 0.009886f
C3817 vdd.n1474 gnd 0.009886f
C3818 vdd.n1475 gnd 0.009886f
C3819 vdd.n1476 gnd 0.007957f
C3820 vdd.n1477 gnd 0.009886f
C3821 vdd.n1478 gnd 0.838538f
C3822 vdd.t176 gnd 0.505144f
C3823 vdd.n1479 gnd 0.580915f
C3824 vdd.n1480 gnd 0.009886f
C3825 vdd.n1481 gnd 0.007957f
C3826 vdd.n1482 gnd 0.009886f
C3827 vdd.n1483 gnd 0.009886f
C3828 vdd.n1484 gnd 0.009886f
C3829 vdd.n1485 gnd 0.007957f
C3830 vdd.n1486 gnd 0.009886f
C3831 vdd.n1487 gnd 0.601121f
C3832 vdd.n1488 gnd 0.009886f
C3833 vdd.n1489 gnd 0.007957f
C3834 vdd.n1490 gnd 0.009886f
C3835 vdd.n1491 gnd 0.009886f
C3836 vdd.n1492 gnd 0.009886f
C3837 vdd.n1493 gnd 0.007957f
C3838 vdd.n1494 gnd 0.009886f
C3839 vdd.n1495 gnd 0.570812f
C3840 vdd.n1496 gnd 0.77287f
C3841 vdd.n1497 gnd 0.009886f
C3842 vdd.n1498 gnd 0.007957f
C3843 vdd.n1499 gnd 0.009886f
C3844 vdd.n1500 gnd 0.009886f
C3845 vdd.n1501 gnd 0.009886f
C3846 vdd.n1502 gnd 0.007957f
C3847 vdd.n1503 gnd 0.009886f
C3848 vdd.n1504 gnd 0.838538f
C3849 vdd.n1505 gnd 0.009886f
C3850 vdd.n1506 gnd 0.007957f
C3851 vdd.n1507 gnd 0.009886f
C3852 vdd.n1508 gnd 0.009886f
C3853 vdd.n1509 gnd 0.009886f
C3854 vdd.n1510 gnd 0.007957f
C3855 vdd.n1511 gnd 0.009886f
C3856 vdd.t132 gnd 0.505144f
C3857 vdd.n1512 gnd 0.732458f
C3858 vdd.n1513 gnd 0.009886f
C3859 vdd.n1514 gnd 0.007957f
C3860 vdd.n1515 gnd 0.009886f
C3861 vdd.n1516 gnd 0.009886f
C3862 vdd.n1517 gnd 0.009886f
C3863 vdd.n1518 gnd 0.007957f
C3864 vdd.n1519 gnd 0.009886f
C3865 vdd.n1520 gnd 0.560709f
C3866 vdd.n1521 gnd 0.009886f
C3867 vdd.n1522 gnd 0.007957f
C3868 vdd.n1523 gnd 0.009886f
C3869 vdd.n1524 gnd 0.009886f
C3870 vdd.n1525 gnd 0.009886f
C3871 vdd.n1526 gnd 0.007957f
C3872 vdd.n1527 gnd 0.009886f
C3873 vdd.n1528 gnd 0.722355f
C3874 vdd.n1529 gnd 0.621327f
C3875 vdd.n1530 gnd 0.009886f
C3876 vdd.n1531 gnd 0.007957f
C3877 vdd.n1532 gnd 0.007598f
C3878 vdd.n1533 gnd 0.005425f
C3879 vdd.n1534 gnd 0.005035f
C3880 vdd.n1535 gnd 0.002785f
C3881 vdd.n1536 gnd 0.006394f
C3882 vdd.n1537 gnd 0.002705f
C3883 vdd.n1538 gnd 0.002864f
C3884 vdd.n1539 gnd 0.005035f
C3885 vdd.n1540 gnd 0.002705f
C3886 vdd.n1541 gnd 0.006394f
C3887 vdd.n1542 gnd 0.002864f
C3888 vdd.n1543 gnd 0.005035f
C3889 vdd.n1544 gnd 0.002705f
C3890 vdd.n1545 gnd 0.004796f
C3891 vdd.n1546 gnd 0.00481f
C3892 vdd.t215 gnd 0.013738f
C3893 vdd.n1547 gnd 0.030567f
C3894 vdd.n1548 gnd 0.159077f
C3895 vdd.n1549 gnd 0.002705f
C3896 vdd.n1550 gnd 0.002864f
C3897 vdd.n1551 gnd 0.006394f
C3898 vdd.n1552 gnd 0.006394f
C3899 vdd.n1553 gnd 0.002864f
C3900 vdd.n1554 gnd 0.002705f
C3901 vdd.n1555 gnd 0.005035f
C3902 vdd.n1556 gnd 0.005035f
C3903 vdd.n1557 gnd 0.002705f
C3904 vdd.n1558 gnd 0.002864f
C3905 vdd.n1559 gnd 0.006394f
C3906 vdd.n1560 gnd 0.006394f
C3907 vdd.n1561 gnd 0.002864f
C3908 vdd.n1562 gnd 0.002705f
C3909 vdd.n1563 gnd 0.005035f
C3910 vdd.n1564 gnd 0.005035f
C3911 vdd.n1565 gnd 0.002705f
C3912 vdd.n1566 gnd 0.002864f
C3913 vdd.n1567 gnd 0.006394f
C3914 vdd.n1568 gnd 0.006394f
C3915 vdd.n1569 gnd 0.015118f
C3916 vdd.n1570 gnd 0.002785f
C3917 vdd.n1571 gnd 0.002705f
C3918 vdd.n1572 gnd 0.013013f
C3919 vdd.n1573 gnd 0.009085f
C3920 vdd.t187 gnd 0.031828f
C3921 vdd.t143 gnd 0.031828f
C3922 vdd.n1574 gnd 0.218742f
C3923 vdd.n1575 gnd 0.172007f
C3924 vdd.t205 gnd 0.031828f
C3925 vdd.t154 gnd 0.031828f
C3926 vdd.n1576 gnd 0.218742f
C3927 vdd.n1577 gnd 0.138808f
C3928 vdd.t244 gnd 0.031828f
C3929 vdd.t256 gnd 0.031828f
C3930 vdd.n1578 gnd 0.218742f
C3931 vdd.n1579 gnd 0.138808f
C3932 vdd.t225 gnd 0.031828f
C3933 vdd.t157 gnd 0.031828f
C3934 vdd.n1580 gnd 0.218742f
C3935 vdd.n1581 gnd 0.138808f
C3936 vdd.t216 gnd 0.031828f
C3937 vdd.t166 gnd 0.031828f
C3938 vdd.n1582 gnd 0.218742f
C3939 vdd.n1583 gnd 0.138808f
C3940 vdd.t248 gnd 0.031828f
C3941 vdd.t193 gnd 0.031828f
C3942 vdd.n1584 gnd 0.218742f
C3943 vdd.n1585 gnd 0.138808f
C3944 vdd.t231 gnd 0.031828f
C3945 vdd.t209 gnd 0.031828f
C3946 vdd.n1586 gnd 0.218742f
C3947 vdd.n1587 gnd 0.138808f
C3948 vdd.n1588 gnd 0.005425f
C3949 vdd.n1589 gnd 0.005035f
C3950 vdd.n1590 gnd 0.002785f
C3951 vdd.n1591 gnd 0.006394f
C3952 vdd.n1592 gnd 0.002705f
C3953 vdd.n1593 gnd 0.002864f
C3954 vdd.n1594 gnd 0.005035f
C3955 vdd.n1595 gnd 0.002705f
C3956 vdd.n1596 gnd 0.006394f
C3957 vdd.n1597 gnd 0.002864f
C3958 vdd.n1598 gnd 0.005035f
C3959 vdd.n1599 gnd 0.002705f
C3960 vdd.n1600 gnd 0.004796f
C3961 vdd.n1601 gnd 0.00481f
C3962 vdd.t177 gnd 0.013738f
C3963 vdd.n1602 gnd 0.030567f
C3964 vdd.n1603 gnd 0.159077f
C3965 vdd.n1604 gnd 0.002705f
C3966 vdd.n1605 gnd 0.002864f
C3967 vdd.n1606 gnd 0.006394f
C3968 vdd.n1607 gnd 0.006394f
C3969 vdd.n1608 gnd 0.002864f
C3970 vdd.n1609 gnd 0.002705f
C3971 vdd.n1610 gnd 0.005035f
C3972 vdd.n1611 gnd 0.005035f
C3973 vdd.n1612 gnd 0.002705f
C3974 vdd.n1613 gnd 0.002864f
C3975 vdd.n1614 gnd 0.006394f
C3976 vdd.n1615 gnd 0.006394f
C3977 vdd.n1616 gnd 0.002864f
C3978 vdd.n1617 gnd 0.002705f
C3979 vdd.n1618 gnd 0.005035f
C3980 vdd.n1619 gnd 0.005035f
C3981 vdd.n1620 gnd 0.002705f
C3982 vdd.n1621 gnd 0.002864f
C3983 vdd.n1622 gnd 0.006394f
C3984 vdd.n1623 gnd 0.006394f
C3985 vdd.n1624 gnd 0.015118f
C3986 vdd.n1625 gnd 0.002785f
C3987 vdd.n1626 gnd 0.002705f
C3988 vdd.n1627 gnd 0.013013f
C3989 vdd.n1628 gnd 0.0088f
C3990 vdd.n1629 gnd 0.103274f
C3991 vdd.n1630 gnd 0.005425f
C3992 vdd.n1631 gnd 0.005035f
C3993 vdd.n1632 gnd 0.002785f
C3994 vdd.n1633 gnd 0.006394f
C3995 vdd.n1634 gnd 0.002705f
C3996 vdd.n1635 gnd 0.002864f
C3997 vdd.n1636 gnd 0.005035f
C3998 vdd.n1637 gnd 0.002705f
C3999 vdd.n1638 gnd 0.006394f
C4000 vdd.n1639 gnd 0.002864f
C4001 vdd.n1640 gnd 0.005035f
C4002 vdd.n1641 gnd 0.002705f
C4003 vdd.n1642 gnd 0.004796f
C4004 vdd.n1643 gnd 0.00481f
C4005 vdd.t249 gnd 0.013738f
C4006 vdd.n1644 gnd 0.030567f
C4007 vdd.n1645 gnd 0.159077f
C4008 vdd.n1646 gnd 0.002705f
C4009 vdd.n1647 gnd 0.002864f
C4010 vdd.n1648 gnd 0.006394f
C4011 vdd.n1649 gnd 0.006394f
C4012 vdd.n1650 gnd 0.002864f
C4013 vdd.n1651 gnd 0.002705f
C4014 vdd.n1652 gnd 0.005035f
C4015 vdd.n1653 gnd 0.005035f
C4016 vdd.n1654 gnd 0.002705f
C4017 vdd.n1655 gnd 0.002864f
C4018 vdd.n1656 gnd 0.006394f
C4019 vdd.n1657 gnd 0.006394f
C4020 vdd.n1658 gnd 0.002864f
C4021 vdd.n1659 gnd 0.002705f
C4022 vdd.n1660 gnd 0.005035f
C4023 vdd.n1661 gnd 0.005035f
C4024 vdd.n1662 gnd 0.002705f
C4025 vdd.n1663 gnd 0.002864f
C4026 vdd.n1664 gnd 0.006394f
C4027 vdd.n1665 gnd 0.006394f
C4028 vdd.n1666 gnd 0.015118f
C4029 vdd.n1667 gnd 0.002785f
C4030 vdd.n1668 gnd 0.002705f
C4031 vdd.n1669 gnd 0.013013f
C4032 vdd.n1670 gnd 0.009085f
C4033 vdd.t221 gnd 0.031828f
C4034 vdd.t170 gnd 0.031828f
C4035 vdd.n1671 gnd 0.218742f
C4036 vdd.n1672 gnd 0.172007f
C4037 vdd.t168 gnd 0.031828f
C4038 vdd.t222 gnd 0.031828f
C4039 vdd.n1673 gnd 0.218742f
C4040 vdd.n1674 gnd 0.138808f
C4041 vdd.t213 gnd 0.031828f
C4042 vdd.t211 gnd 0.031828f
C4043 vdd.n1675 gnd 0.218742f
C4044 vdd.n1676 gnd 0.138808f
C4045 vdd.t161 gnd 0.031828f
C4046 vdd.t141 gnd 0.031828f
C4047 vdd.n1677 gnd 0.218742f
C4048 vdd.n1678 gnd 0.138808f
C4049 vdd.t133 gnd 0.031828f
C4050 vdd.t206 gnd 0.031828f
C4051 vdd.n1679 gnd 0.218742f
C4052 vdd.n1680 gnd 0.138808f
C4053 vdd.t189 gnd 0.031828f
C4054 vdd.t137 gnd 0.031828f
C4055 vdd.n1681 gnd 0.218742f
C4056 vdd.n1682 gnd 0.138808f
C4057 vdd.t131 gnd 0.031828f
C4058 vdd.t226 gnd 0.031828f
C4059 vdd.n1683 gnd 0.218742f
C4060 vdd.n1684 gnd 0.138808f
C4061 vdd.n1685 gnd 0.005425f
C4062 vdd.n1686 gnd 0.005035f
C4063 vdd.n1687 gnd 0.002785f
C4064 vdd.n1688 gnd 0.006394f
C4065 vdd.n1689 gnd 0.002705f
C4066 vdd.n1690 gnd 0.002864f
C4067 vdd.n1691 gnd 0.005035f
C4068 vdd.n1692 gnd 0.002705f
C4069 vdd.n1693 gnd 0.006394f
C4070 vdd.n1694 gnd 0.002864f
C4071 vdd.n1695 gnd 0.005035f
C4072 vdd.n1696 gnd 0.002705f
C4073 vdd.n1697 gnd 0.004796f
C4074 vdd.n1698 gnd 0.00481f
C4075 vdd.t179 gnd 0.013738f
C4076 vdd.n1699 gnd 0.030567f
C4077 vdd.n1700 gnd 0.159077f
C4078 vdd.n1701 gnd 0.002705f
C4079 vdd.n1702 gnd 0.002864f
C4080 vdd.n1703 gnd 0.006394f
C4081 vdd.n1704 gnd 0.006394f
C4082 vdd.n1705 gnd 0.002864f
C4083 vdd.n1706 gnd 0.002705f
C4084 vdd.n1707 gnd 0.005035f
C4085 vdd.n1708 gnd 0.005035f
C4086 vdd.n1709 gnd 0.002705f
C4087 vdd.n1710 gnd 0.002864f
C4088 vdd.n1711 gnd 0.006394f
C4089 vdd.n1712 gnd 0.006394f
C4090 vdd.n1713 gnd 0.002864f
C4091 vdd.n1714 gnd 0.002705f
C4092 vdd.n1715 gnd 0.005035f
C4093 vdd.n1716 gnd 0.005035f
C4094 vdd.n1717 gnd 0.002705f
C4095 vdd.n1718 gnd 0.002864f
C4096 vdd.n1719 gnd 0.006394f
C4097 vdd.n1720 gnd 0.006394f
C4098 vdd.n1721 gnd 0.015118f
C4099 vdd.n1722 gnd 0.002785f
C4100 vdd.n1723 gnd 0.002705f
C4101 vdd.n1724 gnd 0.013013f
C4102 vdd.n1725 gnd 0.0088f
C4103 vdd.n1726 gnd 0.061438f
C4104 vdd.n1727 gnd 0.221376f
C4105 vdd.n1728 gnd 0.005425f
C4106 vdd.n1729 gnd 0.005035f
C4107 vdd.n1730 gnd 0.002785f
C4108 vdd.n1731 gnd 0.006394f
C4109 vdd.n1732 gnd 0.002705f
C4110 vdd.n1733 gnd 0.002864f
C4111 vdd.n1734 gnd 0.005035f
C4112 vdd.n1735 gnd 0.002705f
C4113 vdd.n1736 gnd 0.006394f
C4114 vdd.n1737 gnd 0.002864f
C4115 vdd.n1738 gnd 0.005035f
C4116 vdd.n1739 gnd 0.002705f
C4117 vdd.n1740 gnd 0.004796f
C4118 vdd.n1741 gnd 0.00481f
C4119 vdd.t257 gnd 0.013738f
C4120 vdd.n1742 gnd 0.030567f
C4121 vdd.n1743 gnd 0.159077f
C4122 vdd.n1744 gnd 0.002705f
C4123 vdd.n1745 gnd 0.002864f
C4124 vdd.n1746 gnd 0.006394f
C4125 vdd.n1747 gnd 0.006394f
C4126 vdd.n1748 gnd 0.002864f
C4127 vdd.n1749 gnd 0.002705f
C4128 vdd.n1750 gnd 0.005035f
C4129 vdd.n1751 gnd 0.005035f
C4130 vdd.n1752 gnd 0.002705f
C4131 vdd.n1753 gnd 0.002864f
C4132 vdd.n1754 gnd 0.006394f
C4133 vdd.n1755 gnd 0.006394f
C4134 vdd.n1756 gnd 0.002864f
C4135 vdd.n1757 gnd 0.002705f
C4136 vdd.n1758 gnd 0.005035f
C4137 vdd.n1759 gnd 0.005035f
C4138 vdd.n1760 gnd 0.002705f
C4139 vdd.n1761 gnd 0.002864f
C4140 vdd.n1762 gnd 0.006394f
C4141 vdd.n1763 gnd 0.006394f
C4142 vdd.n1764 gnd 0.015118f
C4143 vdd.n1765 gnd 0.002785f
C4144 vdd.n1766 gnd 0.002705f
C4145 vdd.n1767 gnd 0.013013f
C4146 vdd.n1768 gnd 0.009085f
C4147 vdd.t236 gnd 0.031828f
C4148 vdd.t194 gnd 0.031828f
C4149 vdd.n1769 gnd 0.218742f
C4150 vdd.n1770 gnd 0.172007f
C4151 vdd.t190 gnd 0.031828f
C4152 vdd.t237 gnd 0.031828f
C4153 vdd.n1771 gnd 0.218742f
C4154 vdd.n1772 gnd 0.138808f
C4155 vdd.t220 gnd 0.031828f
C4156 vdd.t219 gnd 0.031828f
C4157 vdd.n1773 gnd 0.218742f
C4158 vdd.n1774 gnd 0.138808f
C4159 vdd.t185 gnd 0.031828f
C4160 vdd.t162 gnd 0.031828f
C4161 vdd.n1775 gnd 0.218742f
C4162 vdd.n1776 gnd 0.138808f
C4163 vdd.t158 gnd 0.031828f
C4164 vdd.t218 gnd 0.031828f
C4165 vdd.n1777 gnd 0.218742f
C4166 vdd.n1778 gnd 0.138808f
C4167 vdd.t200 gnd 0.031828f
C4168 vdd.t159 gnd 0.031828f
C4169 vdd.n1779 gnd 0.218742f
C4170 vdd.n1780 gnd 0.138808f
C4171 vdd.t144 gnd 0.031828f
C4172 vdd.t238 gnd 0.031828f
C4173 vdd.n1781 gnd 0.218742f
C4174 vdd.n1782 gnd 0.138808f
C4175 vdd.n1783 gnd 0.005425f
C4176 vdd.n1784 gnd 0.005035f
C4177 vdd.n1785 gnd 0.002785f
C4178 vdd.n1786 gnd 0.006394f
C4179 vdd.n1787 gnd 0.002705f
C4180 vdd.n1788 gnd 0.002864f
C4181 vdd.n1789 gnd 0.005035f
C4182 vdd.n1790 gnd 0.002705f
C4183 vdd.n1791 gnd 0.006394f
C4184 vdd.n1792 gnd 0.002864f
C4185 vdd.n1793 gnd 0.005035f
C4186 vdd.n1794 gnd 0.002705f
C4187 vdd.n1795 gnd 0.004796f
C4188 vdd.n1796 gnd 0.00481f
C4189 vdd.t197 gnd 0.013738f
C4190 vdd.n1797 gnd 0.030567f
C4191 vdd.n1798 gnd 0.159077f
C4192 vdd.n1799 gnd 0.002705f
C4193 vdd.n1800 gnd 0.002864f
C4194 vdd.n1801 gnd 0.006394f
C4195 vdd.n1802 gnd 0.006394f
C4196 vdd.n1803 gnd 0.002864f
C4197 vdd.n1804 gnd 0.002705f
C4198 vdd.n1805 gnd 0.005035f
C4199 vdd.n1806 gnd 0.005035f
C4200 vdd.n1807 gnd 0.002705f
C4201 vdd.n1808 gnd 0.002864f
C4202 vdd.n1809 gnd 0.006394f
C4203 vdd.n1810 gnd 0.006394f
C4204 vdd.n1811 gnd 0.002864f
C4205 vdd.n1812 gnd 0.002705f
C4206 vdd.n1813 gnd 0.005035f
C4207 vdd.n1814 gnd 0.005035f
C4208 vdd.n1815 gnd 0.002705f
C4209 vdd.n1816 gnd 0.002864f
C4210 vdd.n1817 gnd 0.006394f
C4211 vdd.n1818 gnd 0.006394f
C4212 vdd.n1819 gnd 0.015118f
C4213 vdd.n1820 gnd 0.002785f
C4214 vdd.n1821 gnd 0.002705f
C4215 vdd.n1822 gnd 0.013013f
C4216 vdd.n1823 gnd 0.0088f
C4217 vdd.n1824 gnd 0.061438f
C4218 vdd.n1825 gnd 0.247912f
C4219 vdd.n1826 gnd 2.60377f
C4220 vdd.n1827 gnd 0.583105f
C4221 vdd.n1828 gnd 0.007598f
C4222 vdd.n1829 gnd 0.009886f
C4223 vdd.n1830 gnd 0.007957f
C4224 vdd.n1831 gnd 0.009886f
C4225 vdd.n1832 gnd 0.793075f
C4226 vdd.n1833 gnd 0.009886f
C4227 vdd.n1834 gnd 0.007957f
C4228 vdd.n1835 gnd 0.009886f
C4229 vdd.n1836 gnd 0.009886f
C4230 vdd.n1837 gnd 0.009886f
C4231 vdd.n1838 gnd 0.007957f
C4232 vdd.n1839 gnd 0.009886f
C4233 vdd.t210 gnd 0.505144f
C4234 vdd.n1840 gnd 0.838538f
C4235 vdd.n1841 gnd 0.009886f
C4236 vdd.n1842 gnd 0.007957f
C4237 vdd.n1843 gnd 0.009886f
C4238 vdd.n1844 gnd 0.009886f
C4239 vdd.n1845 gnd 0.009886f
C4240 vdd.n1846 gnd 0.007957f
C4241 vdd.n1847 gnd 0.009886f
C4242 vdd.n1848 gnd 0.712252f
C4243 vdd.n1849 gnd 0.009886f
C4244 vdd.n1850 gnd 0.007957f
C4245 vdd.n1851 gnd 0.009886f
C4246 vdd.n1852 gnd 0.009886f
C4247 vdd.n1853 gnd 0.009886f
C4248 vdd.n1854 gnd 0.007957f
C4249 vdd.n1855 gnd 0.009886f
C4250 vdd.n1856 gnd 0.838538f
C4251 vdd.t153 gnd 0.505144f
C4252 vdd.n1857 gnd 0.540504f
C4253 vdd.n1858 gnd 0.009886f
C4254 vdd.n1859 gnd 0.007957f
C4255 vdd.n1860 gnd 0.009886f
C4256 vdd.n1861 gnd 0.009886f
C4257 vdd.n1862 gnd 0.009886f
C4258 vdd.n1863 gnd 0.007957f
C4259 vdd.n1864 gnd 0.009886f
C4260 vdd.n1865 gnd 0.641532f
C4261 vdd.n1866 gnd 0.009886f
C4262 vdd.n1867 gnd 0.007957f
C4263 vdd.n1868 gnd 0.009886f
C4264 vdd.n1869 gnd 0.009886f
C4265 vdd.n1870 gnd 0.009886f
C4266 vdd.n1871 gnd 0.007957f
C4267 vdd.n1872 gnd 0.009886f
C4268 vdd.n1873 gnd 0.530401f
C4269 vdd.n1874 gnd 0.813281f
C4270 vdd.n1875 gnd 0.009886f
C4271 vdd.n1876 gnd 0.007957f
C4272 vdd.n1877 gnd 0.009886f
C4273 vdd.n1878 gnd 0.009886f
C4274 vdd.n1879 gnd 0.009886f
C4275 vdd.n1880 gnd 0.007957f
C4276 vdd.n1881 gnd 0.009886f
C4277 vdd.n1882 gnd 0.98503f
C4278 vdd.n1883 gnd 0.009886f
C4279 vdd.n1884 gnd 0.007957f
C4280 vdd.n1885 gnd 0.009886f
C4281 vdd.n1886 gnd 0.009886f
C4282 vdd.n1887 gnd 0.022512f
C4283 vdd.n1888 gnd 0.009886f
C4284 vdd.n1889 gnd 0.009886f
C4285 vdd.n1890 gnd 0.007957f
C4286 vdd.n1891 gnd 0.009886f
C4287 vdd.t62 gnd 0.505144f
C4288 vdd.n1892 gnd 0.954721f
C4289 vdd.n1893 gnd 0.009886f
C4290 vdd.n1894 gnd 0.007957f
C4291 vdd.n1895 gnd 0.009886f
C4292 vdd.n1896 gnd 0.009886f
C4293 vdd.n1897 gnd 0.008502f
C4294 vdd.n1898 gnd 0.007957f
C4295 vdd.n1900 gnd 0.009886f
C4296 vdd.n1902 gnd 0.007957f
C4297 vdd.n1903 gnd 0.009886f
C4298 vdd.n1904 gnd 0.007957f
C4299 vdd.n1906 gnd 0.009886f
C4300 vdd.n1907 gnd 0.007957f
C4301 vdd.n1908 gnd 0.009886f
C4302 vdd.n1909 gnd 0.009886f
C4303 vdd.n1910 gnd 0.009886f
C4304 vdd.n1911 gnd 0.009886f
C4305 vdd.n1912 gnd 0.009886f
C4306 vdd.n1913 gnd 0.007957f
C4307 vdd.n1915 gnd 0.009886f
C4308 vdd.n1916 gnd 0.009886f
C4309 vdd.n1917 gnd 0.009886f
C4310 vdd.n1918 gnd 0.009886f
C4311 vdd.n1919 gnd 0.009886f
C4312 vdd.n1920 gnd 0.007957f
C4313 vdd.n1922 gnd 0.009886f
C4314 vdd.n1923 gnd 0.009886f
C4315 vdd.n1924 gnd 0.009886f
C4316 vdd.n1925 gnd 0.009886f
C4317 vdd.n1926 gnd 0.006644f
C4318 vdd.t91 gnd 0.121622f
C4319 vdd.t90 gnd 0.12998f
C4320 vdd.t89 gnd 0.158837f
C4321 vdd.n1927 gnd 0.203606f
C4322 vdd.n1928 gnd 0.171066f
C4323 vdd.n1930 gnd 0.009886f
C4324 vdd.n1931 gnd 0.009886f
C4325 vdd.n1932 gnd 0.007957f
C4326 vdd.n1933 gnd 0.009886f
C4327 vdd.n1935 gnd 0.009886f
C4328 vdd.n1936 gnd 0.009886f
C4329 vdd.n1937 gnd 0.009886f
C4330 vdd.n1938 gnd 0.009886f
C4331 vdd.n1939 gnd 0.007957f
C4332 vdd.n1941 gnd 0.009886f
C4333 vdd.n1942 gnd 0.009886f
C4334 vdd.n1943 gnd 0.009886f
C4335 vdd.n1944 gnd 0.009886f
C4336 vdd.n1945 gnd 0.009886f
C4337 vdd.n1946 gnd 0.007957f
C4338 vdd.n1948 gnd 0.009886f
C4339 vdd.n1949 gnd 0.009886f
C4340 vdd.n1950 gnd 0.009886f
C4341 vdd.n1951 gnd 0.009886f
C4342 vdd.n1952 gnd 0.009886f
C4343 vdd.n1953 gnd 0.007957f
C4344 vdd.n1955 gnd 0.009886f
C4345 vdd.n1956 gnd 0.009886f
C4346 vdd.n1957 gnd 0.009886f
C4347 vdd.n1958 gnd 0.009886f
C4348 vdd.n1959 gnd 0.009886f
C4349 vdd.n1960 gnd 0.007957f
C4350 vdd.n1962 gnd 0.009886f
C4351 vdd.n1963 gnd 0.009886f
C4352 vdd.n1964 gnd 0.009886f
C4353 vdd.n1965 gnd 0.009886f
C4354 vdd.n1966 gnd 0.007877f
C4355 vdd.t80 gnd 0.121622f
C4356 vdd.t79 gnd 0.12998f
C4357 vdd.t78 gnd 0.158837f
C4358 vdd.n1967 gnd 0.203606f
C4359 vdd.n1968 gnd 0.171066f
C4360 vdd.n1970 gnd 0.009886f
C4361 vdd.n1971 gnd 0.009886f
C4362 vdd.n1972 gnd 0.007957f
C4363 vdd.n1973 gnd 0.009886f
C4364 vdd.n1975 gnd 0.009886f
C4365 vdd.n1976 gnd 0.009886f
C4366 vdd.n1977 gnd 0.009886f
C4367 vdd.n1978 gnd 0.009886f
C4368 vdd.n1979 gnd 0.007957f
C4369 vdd.n1981 gnd 0.009886f
C4370 vdd.n1982 gnd 0.009886f
C4371 vdd.n1983 gnd 0.009886f
C4372 vdd.n1984 gnd 0.009886f
C4373 vdd.n1985 gnd 0.009886f
C4374 vdd.n1986 gnd 0.007957f
C4375 vdd.n1988 gnd 0.009886f
C4376 vdd.n1989 gnd 0.009886f
C4377 vdd.n1990 gnd 0.009886f
C4378 vdd.n1991 gnd 0.009886f
C4379 vdd.n1992 gnd 0.009886f
C4380 vdd.n1993 gnd 0.009886f
C4381 vdd.n1994 gnd 0.007957f
C4382 vdd.n1996 gnd 0.009886f
C4383 vdd.n1998 gnd 0.009886f
C4384 vdd.n1999 gnd 0.007957f
C4385 vdd.n2000 gnd 0.007957f
C4386 vdd.n2001 gnd 0.009886f
C4387 vdd.n2003 gnd 0.009886f
C4388 vdd.n2004 gnd 0.007957f
C4389 vdd.n2005 gnd 0.007957f
C4390 vdd.n2006 gnd 0.009886f
C4391 vdd.n2008 gnd 0.009886f
C4392 vdd.n2009 gnd 0.009886f
C4393 vdd.n2010 gnd 0.007957f
C4394 vdd.n2011 gnd 0.007957f
C4395 vdd.n2012 gnd 0.007957f
C4396 vdd.n2013 gnd 0.009886f
C4397 vdd.n2015 gnd 0.009886f
C4398 vdd.n2016 gnd 0.009886f
C4399 vdd.n2017 gnd 0.007957f
C4400 vdd.n2018 gnd 0.007957f
C4401 vdd.n2019 gnd 0.007957f
C4402 vdd.n2020 gnd 0.009886f
C4403 vdd.n2022 gnd 0.009886f
C4404 vdd.n2023 gnd 0.009886f
C4405 vdd.n2024 gnd 0.007957f
C4406 vdd.n2025 gnd 0.007957f
C4407 vdd.n2026 gnd 0.007957f
C4408 vdd.n2027 gnd 0.009886f
C4409 vdd.n2029 gnd 0.009886f
C4410 vdd.n2030 gnd 0.009886f
C4411 vdd.n2031 gnd 0.007957f
C4412 vdd.n2032 gnd 0.009886f
C4413 vdd.n2033 gnd 0.009886f
C4414 vdd.n2034 gnd 0.009886f
C4415 vdd.n2035 gnd 0.016232f
C4416 vdd.n2036 gnd 0.005411f
C4417 vdd.n2037 gnd 0.007957f
C4418 vdd.n2038 gnd 0.009886f
C4419 vdd.n2040 gnd 0.009886f
C4420 vdd.n2041 gnd 0.009886f
C4421 vdd.n2042 gnd 0.007957f
C4422 vdd.n2043 gnd 0.007957f
C4423 vdd.n2044 gnd 0.007957f
C4424 vdd.n2045 gnd 0.009886f
C4425 vdd.n2047 gnd 0.009886f
C4426 vdd.n2048 gnd 0.009886f
C4427 vdd.n2049 gnd 0.007957f
C4428 vdd.n2050 gnd 0.007957f
C4429 vdd.n2051 gnd 0.007957f
C4430 vdd.n2052 gnd 0.009886f
C4431 vdd.n2054 gnd 0.009886f
C4432 vdd.n2055 gnd 0.009886f
C4433 vdd.n2056 gnd 0.007957f
C4434 vdd.n2057 gnd 0.007957f
C4435 vdd.n2058 gnd 0.007957f
C4436 vdd.n2059 gnd 0.009886f
C4437 vdd.n2061 gnd 0.009886f
C4438 vdd.n2062 gnd 0.009886f
C4439 vdd.n2063 gnd 0.007957f
C4440 vdd.n2064 gnd 0.007957f
C4441 vdd.n2065 gnd 0.007957f
C4442 vdd.n2066 gnd 0.009886f
C4443 vdd.n2068 gnd 0.009886f
C4444 vdd.n2069 gnd 0.009886f
C4445 vdd.n2070 gnd 0.007957f
C4446 vdd.n2071 gnd 0.009886f
C4447 vdd.n2072 gnd 0.009886f
C4448 vdd.n2073 gnd 0.009886f
C4449 vdd.n2074 gnd 0.016232f
C4450 vdd.n2075 gnd 0.006644f
C4451 vdd.n2076 gnd 0.007957f
C4452 vdd.n2077 gnd 0.009886f
C4453 vdd.n2079 gnd 0.009886f
C4454 vdd.n2080 gnd 0.009886f
C4455 vdd.n2081 gnd 0.007957f
C4456 vdd.n2082 gnd 0.007957f
C4457 vdd.n2083 gnd 0.007957f
C4458 vdd.n2084 gnd 0.009886f
C4459 vdd.n2086 gnd 0.009886f
C4460 vdd.n2087 gnd 0.009886f
C4461 vdd.n2088 gnd 0.007957f
C4462 vdd.n2089 gnd 0.007957f
C4463 vdd.n2090 gnd 0.007957f
C4464 vdd.n2091 gnd 0.009886f
C4465 vdd.n2093 gnd 0.009886f
C4466 vdd.n2094 gnd 0.009886f
C4467 vdd.n2096 gnd 0.009886f
C4468 vdd.n2097 gnd 0.007957f
C4469 vdd.n2098 gnd 0.006327f
C4470 vdd.n2099 gnd 0.899297f
C4471 vdd.n2101 gnd 0.007957f
C4472 vdd.n2102 gnd 0.007957f
C4473 vdd.n2103 gnd 0.009886f
C4474 vdd.n2105 gnd 0.009886f
C4475 vdd.n2106 gnd 0.009886f
C4476 vdd.n2107 gnd 0.007957f
C4477 vdd.n2108 gnd 0.006604f
C4478 vdd.n2109 gnd 0.022666f
C4479 vdd.n2110 gnd 0.022512f
C4480 vdd.n2111 gnd 0.006604f
C4481 vdd.n2112 gnd 0.022512f
C4482 vdd.n2113 gnd 1.33358f
C4483 vdd.n2114 gnd 0.022512f
C4484 vdd.n2115 gnd 0.022666f
C4485 vdd.n2116 gnd 0.00378f
C4486 vdd.t64 gnd 0.121622f
C4487 vdd.t63 gnd 0.12998f
C4488 vdd.t61 gnd 0.158837f
C4489 vdd.n2117 gnd 0.203606f
C4490 vdd.n2118 gnd 0.171066f
C4491 vdd.n2119 gnd 0.012254f
C4492 vdd.n2120 gnd 0.004177f
C4493 vdd.n2121 gnd 0.008502f
C4494 vdd.n2122 gnd 0.899297f
C4495 vdd.n2123 gnd 0.03537f
C4496 vdd.n2124 gnd 0.006722f
C4497 vdd.n2125 gnd 0.006722f
C4498 vdd.n2126 gnd 0.006722f
C4499 vdd.n2127 gnd 0.006722f
C4500 vdd.n2128 gnd 0.006722f
C4501 vdd.n2129 gnd 0.006722f
C4502 vdd.n2130 gnd 0.006722f
C4503 vdd.n2131 gnd 0.006722f
C4504 vdd.n2133 gnd 0.006722f
C4505 vdd.n2135 gnd 0.006722f
C4506 vdd.n2136 gnd 0.006722f
C4507 vdd.n2137 gnd 0.006722f
C4508 vdd.n2138 gnd 0.006722f
C4509 vdd.n2139 gnd 0.006722f
C4510 vdd.n2141 gnd 0.006722f
C4511 vdd.n2143 gnd 0.006722f
C4512 vdd.n2144 gnd 0.006722f
C4513 vdd.n2145 gnd 0.006722f
C4514 vdd.n2146 gnd 0.006722f
C4515 vdd.n2147 gnd 0.006722f
C4516 vdd.n2149 gnd 0.006722f
C4517 vdd.n2151 gnd 0.006722f
C4518 vdd.n2152 gnd 0.006722f
C4519 vdd.n2153 gnd 0.006722f
C4520 vdd.n2154 gnd 0.006722f
C4521 vdd.n2155 gnd 0.006722f
C4522 vdd.n2157 gnd 0.006722f
C4523 vdd.n2159 gnd 0.006722f
C4524 vdd.n2160 gnd 0.006722f
C4525 vdd.n2161 gnd 0.006722f
C4526 vdd.n2162 gnd 0.006722f
C4527 vdd.n2163 gnd 0.006722f
C4528 vdd.n2165 gnd 0.006722f
C4529 vdd.n2167 gnd 0.006722f
C4530 vdd.n2168 gnd 0.006722f
C4531 vdd.n2169 gnd 0.006722f
C4532 vdd.n2170 gnd 0.006722f
C4533 vdd.n2171 gnd 0.006722f
C4534 vdd.n2173 gnd 0.006722f
C4535 vdd.n2175 gnd 0.006722f
C4536 vdd.n2176 gnd 0.006722f
C4537 vdd.n2177 gnd 0.006722f
C4538 vdd.n2178 gnd 0.006722f
C4539 vdd.n2179 gnd 0.006722f
C4540 vdd.n2181 gnd 0.006722f
C4541 vdd.n2183 gnd 0.006722f
C4542 vdd.n2184 gnd 0.006722f
C4543 vdd.n2185 gnd 0.006722f
C4544 vdd.n2186 gnd 0.006722f
C4545 vdd.n2187 gnd 0.006722f
C4546 vdd.n2189 gnd 0.006722f
C4547 vdd.n2191 gnd 0.006722f
C4548 vdd.n2192 gnd 0.006722f
C4549 vdd.n2193 gnd 0.004893f
C4550 vdd.n2194 gnd 0.009607f
C4551 vdd.n2195 gnd 0.00519f
C4552 vdd.n2196 gnd 0.006722f
C4553 vdd.n2198 gnd 0.006722f
C4554 vdd.n2199 gnd 0.015494f
C4555 vdd.n2200 gnd 0.015494f
C4556 vdd.n2201 gnd 0.014559f
C4557 vdd.n2202 gnd 0.006722f
C4558 vdd.n2203 gnd 0.006722f
C4559 vdd.n2204 gnd 0.006722f
C4560 vdd.n2205 gnd 0.006722f
C4561 vdd.n2206 gnd 0.006722f
C4562 vdd.n2207 gnd 0.006722f
C4563 vdd.n2208 gnd 0.006722f
C4564 vdd.n2209 gnd 0.006722f
C4565 vdd.n2210 gnd 0.006722f
C4566 vdd.n2211 gnd 0.006722f
C4567 vdd.n2212 gnd 0.006722f
C4568 vdd.n2213 gnd 0.006722f
C4569 vdd.n2214 gnd 0.006722f
C4570 vdd.n2215 gnd 0.006722f
C4571 vdd.n2216 gnd 0.006722f
C4572 vdd.n2217 gnd 0.006722f
C4573 vdd.n2218 gnd 0.006722f
C4574 vdd.n2219 gnd 0.006722f
C4575 vdd.n2220 gnd 0.006722f
C4576 vdd.n2221 gnd 0.006722f
C4577 vdd.n2222 gnd 0.006722f
C4578 vdd.n2223 gnd 0.006722f
C4579 vdd.n2224 gnd 0.006722f
C4580 vdd.n2225 gnd 0.006722f
C4581 vdd.n2226 gnd 0.006722f
C4582 vdd.n2227 gnd 0.006722f
C4583 vdd.n2228 gnd 0.006722f
C4584 vdd.n2229 gnd 0.006722f
C4585 vdd.n2230 gnd 0.006722f
C4586 vdd.n2231 gnd 0.006722f
C4587 vdd.n2232 gnd 0.006722f
C4588 vdd.n2233 gnd 0.006722f
C4589 vdd.n2234 gnd 0.006722f
C4590 vdd.n2235 gnd 0.006722f
C4591 vdd.n2236 gnd 0.006722f
C4592 vdd.n2237 gnd 0.006722f
C4593 vdd.n2238 gnd 0.006722f
C4594 vdd.n2239 gnd 0.006722f
C4595 vdd.n2240 gnd 0.006722f
C4596 vdd.n2241 gnd 0.006722f
C4597 vdd.n2242 gnd 0.006722f
C4598 vdd.n2243 gnd 0.006722f
C4599 vdd.n2244 gnd 0.006722f
C4600 vdd.n2245 gnd 0.006722f
C4601 vdd.n2246 gnd 0.006722f
C4602 vdd.n2247 gnd 0.006722f
C4603 vdd.n2248 gnd 0.006722f
C4604 vdd.n2249 gnd 0.006722f
C4605 vdd.n2250 gnd 0.006722f
C4606 vdd.n2251 gnd 0.409166f
C4607 vdd.n2252 gnd 0.006722f
C4608 vdd.n2253 gnd 0.006722f
C4609 vdd.n2254 gnd 0.006722f
C4610 vdd.n2255 gnd 0.006722f
C4611 vdd.n2256 gnd 0.006722f
C4612 vdd.n2257 gnd 0.006722f
C4613 vdd.n2258 gnd 0.006722f
C4614 vdd.n2259 gnd 0.006722f
C4615 vdd.n2260 gnd 0.006722f
C4616 vdd.n2261 gnd 0.006722f
C4617 vdd.n2262 gnd 0.006722f
C4618 vdd.n2263 gnd 0.621327f
C4619 vdd.n2264 gnd 0.006722f
C4620 vdd.n2265 gnd 0.006722f
C4621 vdd.n2266 gnd 0.006722f
C4622 vdd.n2267 gnd 0.006722f
C4623 vdd.n2268 gnd 0.006722f
C4624 vdd.n2269 gnd 0.006722f
C4625 vdd.n2270 gnd 0.006722f
C4626 vdd.n2271 gnd 0.006722f
C4627 vdd.n2272 gnd 0.006722f
C4628 vdd.n2273 gnd 0.006722f
C4629 vdd.n2274 gnd 0.006722f
C4630 vdd.n2275 gnd 0.217212f
C4631 vdd.n2276 gnd 0.006722f
C4632 vdd.n2277 gnd 0.006722f
C4633 vdd.n2278 gnd 0.006722f
C4634 vdd.n2279 gnd 0.006722f
C4635 vdd.n2280 gnd 0.006722f
C4636 vdd.n2281 gnd 0.006722f
C4637 vdd.n2282 gnd 0.006722f
C4638 vdd.n2283 gnd 0.006722f
C4639 vdd.n2284 gnd 0.006722f
C4640 vdd.n2285 gnd 0.006722f
C4641 vdd.n2286 gnd 0.006722f
C4642 vdd.n2287 gnd 0.006722f
C4643 vdd.n2288 gnd 0.006722f
C4644 vdd.n2289 gnd 0.006722f
C4645 vdd.n2290 gnd 0.006722f
C4646 vdd.n2291 gnd 0.006722f
C4647 vdd.n2292 gnd 0.006722f
C4648 vdd.n2293 gnd 0.006722f
C4649 vdd.n2294 gnd 0.006722f
C4650 vdd.n2295 gnd 0.006722f
C4651 vdd.n2296 gnd 0.006722f
C4652 vdd.n2297 gnd 0.006722f
C4653 vdd.n2298 gnd 0.006722f
C4654 vdd.n2299 gnd 0.006722f
C4655 vdd.n2300 gnd 0.006722f
C4656 vdd.n2301 gnd 0.006722f
C4657 vdd.n2302 gnd 0.006722f
C4658 vdd.n2303 gnd 0.006722f
C4659 vdd.n2304 gnd 0.006722f
C4660 vdd.n2305 gnd 0.006722f
C4661 vdd.n2306 gnd 0.006722f
C4662 vdd.n2307 gnd 0.006722f
C4663 vdd.n2308 gnd 0.006722f
C4664 vdd.n2309 gnd 0.006722f
C4665 vdd.n2310 gnd 0.006722f
C4666 vdd.n2311 gnd 0.014559f
C4667 vdd.n2312 gnd 0.015494f
C4668 vdd.n2313 gnd 0.015494f
C4669 vdd.n2315 gnd 0.006722f
C4670 vdd.n2317 gnd 0.006722f
C4671 vdd.n2318 gnd 0.00519f
C4672 vdd.n2319 gnd 0.009607f
C4673 vdd.n2320 gnd 0.004893f
C4674 vdd.n2321 gnd 0.006722f
C4675 vdd.n2322 gnd 0.006722f
C4676 vdd.n2324 gnd 0.006722f
C4677 vdd.n2326 gnd 0.006722f
C4678 vdd.n2327 gnd 0.006722f
C4679 vdd.n2328 gnd 0.006722f
C4680 vdd.n2329 gnd 0.006722f
C4681 vdd.n2330 gnd 0.006722f
C4682 vdd.n2332 gnd 0.006722f
C4683 vdd.n2334 gnd 0.006722f
C4684 vdd.n2335 gnd 0.006722f
C4685 vdd.n2336 gnd 0.006722f
C4686 vdd.n2337 gnd 0.006722f
C4687 vdd.n2338 gnd 0.006722f
C4688 vdd.n2340 gnd 0.006722f
C4689 vdd.n2342 gnd 0.006722f
C4690 vdd.n2343 gnd 0.006722f
C4691 vdd.n2344 gnd 0.006722f
C4692 vdd.n2345 gnd 0.006722f
C4693 vdd.n2346 gnd 0.006722f
C4694 vdd.n2348 gnd 0.006722f
C4695 vdd.n2350 gnd 0.006722f
C4696 vdd.n2351 gnd 0.006722f
C4697 vdd.n2352 gnd 0.006722f
C4698 vdd.n2353 gnd 0.006722f
C4699 vdd.n2354 gnd 0.006722f
C4700 vdd.n2356 gnd 0.006722f
C4701 vdd.n2358 gnd 0.006722f
C4702 vdd.n2359 gnd 0.006722f
C4703 vdd.n2360 gnd 0.006722f
C4704 vdd.n2361 gnd 0.006722f
C4705 vdd.n2362 gnd 0.006722f
C4706 vdd.n2364 gnd 0.006722f
C4707 vdd.n2366 gnd 0.006722f
C4708 vdd.n2367 gnd 0.006722f
C4709 vdd.n2368 gnd 0.006722f
C4710 vdd.n2369 gnd 0.006722f
C4711 vdd.n2370 gnd 0.006722f
C4712 vdd.n2372 gnd 0.006722f
C4713 vdd.n2373 gnd 0.006722f
C4714 vdd.n2374 gnd 0.006722f
C4715 vdd.n2375 gnd 0.006722f
C4716 vdd.n2376 gnd 0.006722f
C4717 vdd.n2377 gnd 0.006722f
C4718 vdd.n2379 gnd 0.006722f
C4719 vdd.n2380 gnd 0.006722f
C4720 vdd.n2381 gnd 0.015494f
C4721 vdd.n2382 gnd 0.014559f
C4722 vdd.n2383 gnd 0.014559f
C4723 vdd.n2384 gnd 0.94967f
C4724 vdd.n2385 gnd 0.014559f
C4725 vdd.n2386 gnd 0.014559f
C4726 vdd.n2387 gnd 0.006722f
C4727 vdd.n2388 gnd 0.006722f
C4728 vdd.n2389 gnd 0.006722f
C4729 vdd.n2390 gnd 0.469784f
C4730 vdd.n2391 gnd 0.006722f
C4731 vdd.n2392 gnd 0.006722f
C4732 vdd.n2393 gnd 0.006722f
C4733 vdd.n2394 gnd 0.006722f
C4734 vdd.n2395 gnd 0.006722f
C4735 vdd.n2396 gnd 0.686995f
C4736 vdd.n2397 gnd 0.006722f
C4737 vdd.n2398 gnd 0.006722f
C4738 vdd.n2399 gnd 0.006722f
C4739 vdd.n2400 gnd 0.006722f
C4740 vdd.n2401 gnd 0.006722f
C4741 vdd.n2402 gnd 0.686995f
C4742 vdd.n2403 gnd 0.006722f
C4743 vdd.n2404 gnd 0.006722f
C4744 vdd.n2405 gnd 0.006722f
C4745 vdd.n2406 gnd 0.006722f
C4746 vdd.n2407 gnd 0.006722f
C4747 vdd.n2408 gnd 0.348549f
C4748 vdd.n2409 gnd 0.006722f
C4749 vdd.n2410 gnd 0.006722f
C4750 vdd.n2411 gnd 0.006722f
C4751 vdd.n2412 gnd 0.006722f
C4752 vdd.n2413 gnd 0.006722f
C4753 vdd.n2414 gnd 0.500092f
C4754 vdd.n2415 gnd 0.006722f
C4755 vdd.n2416 gnd 0.006722f
C4756 vdd.n2417 gnd 0.006722f
C4757 vdd.n2418 gnd 0.006722f
C4758 vdd.n2419 gnd 0.006722f
C4759 vdd.n2420 gnd 0.651635f
C4760 vdd.n2421 gnd 0.006722f
C4761 vdd.n2422 gnd 0.006722f
C4762 vdd.n2423 gnd 0.006722f
C4763 vdd.n2424 gnd 0.006722f
C4764 vdd.n2425 gnd 0.006722f
C4765 vdd.n2426 gnd 0.686995f
C4766 vdd.n2427 gnd 0.006722f
C4767 vdd.n2428 gnd 0.006722f
C4768 vdd.n2429 gnd 0.006722f
C4769 vdd.n2430 gnd 0.006722f
C4770 vdd.n2431 gnd 0.006722f
C4771 vdd.n2432 gnd 0.570812f
C4772 vdd.n2433 gnd 0.006722f
C4773 vdd.n2434 gnd 0.006722f
C4774 vdd.n2435 gnd 0.005536f
C4775 vdd.n2436 gnd 0.019474f
C4776 vdd.n2437 gnd 0.004548f
C4777 vdd.n2438 gnd 0.006722f
C4778 vdd.n2439 gnd 0.419269f
C4779 vdd.n2440 gnd 0.006722f
C4780 vdd.n2441 gnd 0.006722f
C4781 vdd.n2442 gnd 0.006722f
C4782 vdd.n2443 gnd 0.006722f
C4783 vdd.n2444 gnd 0.006722f
C4784 vdd.n2445 gnd 0.419269f
C4785 vdd.n2446 gnd 0.006722f
C4786 vdd.n2447 gnd 0.006722f
C4787 vdd.n2448 gnd 0.006722f
C4788 vdd.n2449 gnd 0.006722f
C4789 vdd.n2450 gnd 0.006722f
C4790 vdd.n2451 gnd 0.570812f
C4791 vdd.n2452 gnd 0.006722f
C4792 vdd.n2453 gnd 0.006722f
C4793 vdd.n2454 gnd 0.006722f
C4794 vdd.n2455 gnd 0.006722f
C4795 vdd.n2456 gnd 0.006722f
C4796 vdd.n2457 gnd 0.585967f
C4797 vdd.n2458 gnd 0.006722f
C4798 vdd.n2459 gnd 0.006722f
C4799 vdd.n2460 gnd 0.006722f
C4800 vdd.n2461 gnd 0.006722f
C4801 vdd.n2462 gnd 0.006722f
C4802 vdd.n2463 gnd 0.434423f
C4803 vdd.n2464 gnd 0.006722f
C4804 vdd.n2465 gnd 0.006722f
C4805 vdd.n2466 gnd 0.006722f
C4806 vdd.n2467 gnd 0.006722f
C4807 vdd.n2468 gnd 0.006722f
C4808 vdd.n2469 gnd 0.217212f
C4809 vdd.n2470 gnd 0.006722f
C4810 vdd.n2471 gnd 0.006722f
C4811 vdd.n2472 gnd 0.006722f
C4812 vdd.n2473 gnd 0.006722f
C4813 vdd.n2474 gnd 0.006722f
C4814 vdd.n2475 gnd 0.217212f
C4815 vdd.n2476 gnd 0.006722f
C4816 vdd.n2477 gnd 0.006722f
C4817 vdd.n2478 gnd 0.006722f
C4818 vdd.n2479 gnd 0.006722f
C4819 vdd.n2480 gnd 0.006722f
C4820 vdd.n2481 gnd 0.686995f
C4821 vdd.n2482 gnd 0.006722f
C4822 vdd.n2483 gnd 0.006722f
C4823 vdd.n2484 gnd 0.006722f
C4824 vdd.n2485 gnd 0.006722f
C4825 vdd.n2486 gnd 0.006722f
C4826 vdd.n2487 gnd 0.006722f
C4827 vdd.n2488 gnd 0.006722f
C4828 vdd.n2489 gnd 0.495041f
C4829 vdd.n2490 gnd 0.006722f
C4830 vdd.n2491 gnd 0.006722f
C4831 vdd.n2492 gnd 0.006722f
C4832 vdd.n2493 gnd 0.006722f
C4833 vdd.n2494 gnd 0.006722f
C4834 vdd.n2495 gnd 0.006722f
C4835 vdd.n2496 gnd 0.429372f
C4836 vdd.n2497 gnd 0.006722f
C4837 vdd.n2498 gnd 0.006722f
C4838 vdd.n2499 gnd 0.006722f
C4839 vdd.n2500 gnd 0.015411f
C4840 vdd.n2501 gnd 0.014642f
C4841 vdd.n2502 gnd 0.006722f
C4842 vdd.n2503 gnd 0.006722f
C4843 vdd.n2504 gnd 0.00519f
C4844 vdd.n2505 gnd 0.006722f
C4845 vdd.n2506 gnd 0.006722f
C4846 vdd.n2507 gnd 0.004893f
C4847 vdd.n2508 gnd 0.006722f
C4848 vdd.n2509 gnd 0.006722f
C4849 vdd.n2510 gnd 0.006722f
C4850 vdd.n2511 gnd 0.006722f
C4851 vdd.n2512 gnd 0.006722f
C4852 vdd.n2513 gnd 0.006722f
C4853 vdd.n2514 gnd 0.006722f
C4854 vdd.n2515 gnd 0.006722f
C4855 vdd.n2516 gnd 0.006722f
C4856 vdd.n2517 gnd 0.006722f
C4857 vdd.n2518 gnd 0.006722f
C4858 vdd.n2519 gnd 0.006722f
C4859 vdd.n2520 gnd 0.006722f
C4860 vdd.n2521 gnd 0.006722f
C4861 vdd.n2522 gnd 0.006722f
C4862 vdd.n2523 gnd 0.006722f
C4863 vdd.n2524 gnd 0.006722f
C4864 vdd.n2525 gnd 0.006722f
C4865 vdd.n2526 gnd 0.006722f
C4866 vdd.n2527 gnd 0.006722f
C4867 vdd.n2528 gnd 0.006722f
C4868 vdd.n2529 gnd 0.006722f
C4869 vdd.n2530 gnd 0.006722f
C4870 vdd.n2531 gnd 0.006722f
C4871 vdd.n2532 gnd 0.006722f
C4872 vdd.n2533 gnd 0.006722f
C4873 vdd.n2534 gnd 0.006722f
C4874 vdd.n2535 gnd 0.006722f
C4875 vdd.n2536 gnd 0.006722f
C4876 vdd.n2537 gnd 0.006722f
C4877 vdd.n2538 gnd 0.006722f
C4878 vdd.n2539 gnd 0.006722f
C4879 vdd.n2540 gnd 0.006722f
C4880 vdd.n2541 gnd 0.006722f
C4881 vdd.n2542 gnd 0.006722f
C4882 vdd.n2543 gnd 0.006722f
C4883 vdd.n2544 gnd 0.006722f
C4884 vdd.n2545 gnd 0.006722f
C4885 vdd.n2546 gnd 0.006722f
C4886 vdd.n2547 gnd 0.006722f
C4887 vdd.n2548 gnd 0.006722f
C4888 vdd.n2549 gnd 0.006722f
C4889 vdd.n2550 gnd 0.006722f
C4890 vdd.n2551 gnd 0.006722f
C4891 vdd.n2552 gnd 0.006722f
C4892 vdd.n2553 gnd 0.006722f
C4893 vdd.n2554 gnd 0.006722f
C4894 vdd.n2555 gnd 0.006722f
C4895 vdd.n2556 gnd 0.006722f
C4896 vdd.n2557 gnd 0.006722f
C4897 vdd.n2558 gnd 0.006722f
C4898 vdd.n2559 gnd 0.006722f
C4899 vdd.n2560 gnd 0.006722f
C4900 vdd.n2561 gnd 0.006722f
C4901 vdd.n2562 gnd 0.006722f
C4902 vdd.n2563 gnd 0.006722f
C4903 vdd.n2564 gnd 0.006722f
C4904 vdd.n2565 gnd 0.006722f
C4905 vdd.n2566 gnd 0.006722f
C4906 vdd.n2567 gnd 0.006722f
C4907 vdd.n2568 gnd 0.015494f
C4908 vdd.n2569 gnd 0.014559f
C4909 vdd.n2570 gnd 0.014559f
C4910 vdd.n2571 gnd 0.798127f
C4911 vdd.n2572 gnd 0.014559f
C4912 vdd.n2573 gnd 0.015494f
C4913 vdd.n2574 gnd 0.014642f
C4914 vdd.n2575 gnd 0.006722f
C4915 vdd.n2576 gnd 0.006722f
C4916 vdd.n2577 gnd 0.006722f
C4917 vdd.n2578 gnd 0.00519f
C4918 vdd.n2579 gnd 0.009607f
C4919 vdd.n2580 gnd 0.004893f
C4920 vdd.n2581 gnd 0.006722f
C4921 vdd.n2582 gnd 0.006722f
C4922 vdd.n2583 gnd 0.006722f
C4923 vdd.n2584 gnd 0.006722f
C4924 vdd.n2585 gnd 0.006722f
C4925 vdd.n2586 gnd 0.006722f
C4926 vdd.n2587 gnd 0.006722f
C4927 vdd.n2588 gnd 0.006722f
C4928 vdd.n2589 gnd 0.006722f
C4929 vdd.n2590 gnd 0.006722f
C4930 vdd.n2591 gnd 0.006722f
C4931 vdd.n2592 gnd 0.006722f
C4932 vdd.n2593 gnd 0.006722f
C4933 vdd.n2594 gnd 0.006722f
C4934 vdd.n2595 gnd 0.006722f
C4935 vdd.n2596 gnd 0.006722f
C4936 vdd.n2597 gnd 0.006722f
C4937 vdd.n2598 gnd 0.006722f
C4938 vdd.n2599 gnd 0.006722f
C4939 vdd.n2600 gnd 0.006722f
C4940 vdd.n2601 gnd 0.006722f
C4941 vdd.n2602 gnd 0.006722f
C4942 vdd.n2603 gnd 0.006722f
C4943 vdd.n2604 gnd 0.006722f
C4944 vdd.n2605 gnd 0.006722f
C4945 vdd.n2606 gnd 0.006722f
C4946 vdd.n2607 gnd 0.006722f
C4947 vdd.n2608 gnd 0.006722f
C4948 vdd.n2609 gnd 0.006722f
C4949 vdd.n2610 gnd 0.006722f
C4950 vdd.n2611 gnd 0.006722f
C4951 vdd.n2612 gnd 0.006722f
C4952 vdd.n2613 gnd 0.006722f
C4953 vdd.n2614 gnd 0.006722f
C4954 vdd.n2615 gnd 0.006722f
C4955 vdd.n2616 gnd 0.006722f
C4956 vdd.n2617 gnd 0.006722f
C4957 vdd.n2618 gnd 0.006722f
C4958 vdd.n2619 gnd 0.006722f
C4959 vdd.n2620 gnd 0.006722f
C4960 vdd.n2621 gnd 0.006722f
C4961 vdd.n2622 gnd 0.006722f
C4962 vdd.n2623 gnd 0.006722f
C4963 vdd.n2624 gnd 0.006722f
C4964 vdd.n2625 gnd 0.006722f
C4965 vdd.n2626 gnd 0.006722f
C4966 vdd.n2627 gnd 0.006722f
C4967 vdd.n2628 gnd 0.006722f
C4968 vdd.n2629 gnd 0.006722f
C4969 vdd.n2630 gnd 0.006722f
C4970 vdd.n2631 gnd 0.006722f
C4971 vdd.n2632 gnd 0.006722f
C4972 vdd.n2633 gnd 0.006722f
C4973 vdd.n2634 gnd 0.006722f
C4974 vdd.n2635 gnd 0.006722f
C4975 vdd.n2636 gnd 0.006722f
C4976 vdd.n2637 gnd 0.006722f
C4977 vdd.n2638 gnd 0.006722f
C4978 vdd.n2639 gnd 0.006722f
C4979 vdd.n2640 gnd 0.006722f
C4980 vdd.n2641 gnd 0.015494f
C4981 vdd.n2642 gnd 0.015494f
C4982 vdd.n2643 gnd 0.838538f
C4983 vdd.t111 gnd 2.98035f
C4984 vdd.t119 gnd 2.98035f
C4985 vdd.n2677 gnd 0.006722f
C4986 vdd.t100 gnd 0.27165f
C4987 vdd.t101 gnd 0.278068f
C4988 vdd.t99 gnd 0.177344f
C4989 vdd.n2678 gnd 0.095845f
C4990 vdd.n2679 gnd 0.054366f
C4991 vdd.n2680 gnd 0.009607f
C4992 vdd.n2681 gnd 0.006722f
C4993 vdd.n2682 gnd 0.006722f
C4994 vdd.n2683 gnd 0.006722f
C4995 vdd.n2684 gnd 0.006722f
C4996 vdd.n2685 gnd 0.006722f
C4997 vdd.n2686 gnd 0.006722f
C4998 vdd.n2687 gnd 0.006722f
C4999 vdd.n2688 gnd 0.006722f
C5000 vdd.n2689 gnd 0.006722f
C5001 vdd.n2690 gnd 0.006722f
C5002 vdd.n2691 gnd 0.006722f
C5003 vdd.n2692 gnd 0.006722f
C5004 vdd.n2693 gnd 0.006722f
C5005 vdd.n2694 gnd 0.006722f
C5006 vdd.n2695 gnd 0.006722f
C5007 vdd.n2696 gnd 0.006722f
C5008 vdd.n2697 gnd 0.006722f
C5009 vdd.n2698 gnd 0.006722f
C5010 vdd.n2699 gnd 0.006722f
C5011 vdd.n2700 gnd 0.006722f
C5012 vdd.n2701 gnd 0.006722f
C5013 vdd.n2702 gnd 0.006722f
C5014 vdd.n2703 gnd 0.006722f
C5015 vdd.n2704 gnd 0.006722f
C5016 vdd.n2705 gnd 0.006722f
C5017 vdd.n2706 gnd 0.006722f
C5018 vdd.n2707 gnd 0.006722f
C5019 vdd.n2708 gnd 0.006722f
C5020 vdd.n2709 gnd 0.006722f
C5021 vdd.n2710 gnd 0.006722f
C5022 vdd.n2711 gnd 0.006722f
C5023 vdd.n2712 gnd 0.006722f
C5024 vdd.n2713 gnd 0.006722f
C5025 vdd.n2714 gnd 0.006722f
C5026 vdd.n2715 gnd 0.006722f
C5027 vdd.n2716 gnd 0.006722f
C5028 vdd.n2717 gnd 0.006722f
C5029 vdd.n2718 gnd 0.006722f
C5030 vdd.n2719 gnd 0.006722f
C5031 vdd.n2720 gnd 0.006722f
C5032 vdd.n2721 gnd 0.006722f
C5033 vdd.n2722 gnd 0.006722f
C5034 vdd.n2723 gnd 0.006722f
C5035 vdd.n2724 gnd 0.006722f
C5036 vdd.n2725 gnd 0.006722f
C5037 vdd.n2726 gnd 0.006722f
C5038 vdd.n2727 gnd 0.006722f
C5039 vdd.n2728 gnd 0.006722f
C5040 vdd.n2729 gnd 0.006722f
C5041 vdd.n2730 gnd 0.006722f
C5042 vdd.n2731 gnd 0.006722f
C5043 vdd.n2732 gnd 0.006722f
C5044 vdd.n2733 gnd 0.006722f
C5045 vdd.n2734 gnd 0.006722f
C5046 vdd.n2735 gnd 0.006722f
C5047 vdd.n2736 gnd 0.006722f
C5048 vdd.n2737 gnd 0.006722f
C5049 vdd.n2738 gnd 0.006722f
C5050 vdd.n2739 gnd 0.006722f
C5051 vdd.n2740 gnd 0.006722f
C5052 vdd.n2741 gnd 0.004893f
C5053 vdd.n2742 gnd 0.006722f
C5054 vdd.n2743 gnd 0.006722f
C5055 vdd.n2744 gnd 0.00519f
C5056 vdd.n2745 gnd 0.006722f
C5057 vdd.n2746 gnd 0.006722f
C5058 vdd.t87 gnd 0.27165f
C5059 vdd.t88 gnd 0.278068f
C5060 vdd.t85 gnd 0.177344f
C5061 vdd.n2747 gnd 0.095845f
C5062 vdd.n2748 gnd 0.054366f
C5063 vdd.n2749 gnd 0.006722f
C5064 vdd.n2750 gnd 0.006722f
C5065 vdd.n2751 gnd 0.006722f
C5066 vdd.n2752 gnd 0.006722f
C5067 vdd.n2753 gnd 0.006722f
C5068 vdd.n2754 gnd 0.006722f
C5069 vdd.n2755 gnd 0.006722f
C5070 vdd.n2756 gnd 0.006722f
C5071 vdd.n2757 gnd 0.006722f
C5072 vdd.n2758 gnd 0.006722f
C5073 vdd.n2759 gnd 0.006722f
C5074 vdd.n2760 gnd 0.006722f
C5075 vdd.n2761 gnd 0.006722f
C5076 vdd.n2762 gnd 0.006722f
C5077 vdd.n2763 gnd 0.006722f
C5078 vdd.n2764 gnd 0.006722f
C5079 vdd.n2765 gnd 0.006722f
C5080 vdd.n2766 gnd 0.006722f
C5081 vdd.n2767 gnd 0.006722f
C5082 vdd.n2768 gnd 0.006722f
C5083 vdd.n2769 gnd 0.006722f
C5084 vdd.n2770 gnd 0.006722f
C5085 vdd.n2771 gnd 0.006722f
C5086 vdd.n2772 gnd 0.006722f
C5087 vdd.n2773 gnd 0.006722f
C5088 vdd.n2774 gnd 0.006722f
C5089 vdd.n2775 gnd 0.006722f
C5090 vdd.n2776 gnd 0.006722f
C5091 vdd.n2777 gnd 0.006722f
C5092 vdd.n2778 gnd 0.006722f
C5093 vdd.n2779 gnd 0.006722f
C5094 vdd.n2780 gnd 0.006722f
C5095 vdd.n2781 gnd 0.006722f
C5096 vdd.n2782 gnd 0.006722f
C5097 vdd.n2783 gnd 0.006722f
C5098 vdd.n2784 gnd 0.006722f
C5099 vdd.n2785 gnd 0.006722f
C5100 vdd.n2786 gnd 0.006722f
C5101 vdd.n2787 gnd 0.006722f
C5102 vdd.n2788 gnd 0.006722f
C5103 vdd.n2789 gnd 0.006722f
C5104 vdd.n2790 gnd 0.006722f
C5105 vdd.n2791 gnd 0.006722f
C5106 vdd.n2792 gnd 0.006722f
C5107 vdd.n2793 gnd 0.006722f
C5108 vdd.n2794 gnd 0.006722f
C5109 vdd.n2795 gnd 0.006722f
C5110 vdd.n2796 gnd 0.006722f
C5111 vdd.n2797 gnd 0.006722f
C5112 vdd.n2798 gnd 0.006722f
C5113 vdd.n2799 gnd 0.006722f
C5114 vdd.n2800 gnd 0.006722f
C5115 vdd.n2801 gnd 0.006722f
C5116 vdd.n2802 gnd 0.006722f
C5117 vdd.n2803 gnd 0.006722f
C5118 vdd.n2804 gnd 0.006722f
C5119 vdd.n2805 gnd 0.006722f
C5120 vdd.n2806 gnd 0.004893f
C5121 vdd.n2807 gnd 0.009607f
C5122 vdd.n2808 gnd 0.00519f
C5123 vdd.n2809 gnd 0.006722f
C5124 vdd.n2810 gnd 0.006722f
C5125 vdd.n2811 gnd 0.006722f
C5126 vdd.n2812 gnd 0.015494f
C5127 vdd.n2813 gnd 0.015494f
C5128 vdd.n2814 gnd 0.014559f
C5129 vdd.n2815 gnd 0.006722f
C5130 vdd.n2816 gnd 0.006722f
C5131 vdd.n2817 gnd 0.006722f
C5132 vdd.n2818 gnd 0.006722f
C5133 vdd.n2819 gnd 0.006722f
C5134 vdd.n2820 gnd 0.006722f
C5135 vdd.n2821 gnd 0.006722f
C5136 vdd.n2822 gnd 0.006722f
C5137 vdd.n2823 gnd 0.006722f
C5138 vdd.n2824 gnd 0.006722f
C5139 vdd.n2825 gnd 0.006722f
C5140 vdd.n2826 gnd 0.006722f
C5141 vdd.n2827 gnd 0.006722f
C5142 vdd.n2828 gnd 0.006722f
C5143 vdd.n2829 gnd 0.006722f
C5144 vdd.n2830 gnd 0.006722f
C5145 vdd.n2831 gnd 0.006722f
C5146 vdd.n2832 gnd 0.006722f
C5147 vdd.n2833 gnd 0.006722f
C5148 vdd.n2834 gnd 0.006722f
C5149 vdd.n2835 gnd 0.006722f
C5150 vdd.n2836 gnd 0.006722f
C5151 vdd.n2837 gnd 0.006722f
C5152 vdd.n2838 gnd 0.006722f
C5153 vdd.n2839 gnd 0.006722f
C5154 vdd.n2840 gnd 0.006722f
C5155 vdd.n2841 gnd 0.006722f
C5156 vdd.n2842 gnd 0.006722f
C5157 vdd.n2843 gnd 0.006722f
C5158 vdd.n2844 gnd 0.006722f
C5159 vdd.n2845 gnd 0.006722f
C5160 vdd.n2846 gnd 0.006722f
C5161 vdd.n2847 gnd 0.006722f
C5162 vdd.n2848 gnd 0.006722f
C5163 vdd.n2849 gnd 0.006722f
C5164 vdd.n2850 gnd 0.006722f
C5165 vdd.n2851 gnd 0.006722f
C5166 vdd.n2852 gnd 0.006722f
C5167 vdd.n2853 gnd 0.006722f
C5168 vdd.n2854 gnd 0.006722f
C5169 vdd.n2855 gnd 0.006722f
C5170 vdd.n2856 gnd 0.006722f
C5171 vdd.n2857 gnd 0.006722f
C5172 vdd.n2858 gnd 0.006722f
C5173 vdd.n2859 gnd 0.006722f
C5174 vdd.n2860 gnd 0.006722f
C5175 vdd.n2861 gnd 0.006722f
C5176 vdd.n2862 gnd 0.006722f
C5177 vdd.n2863 gnd 0.006722f
C5178 vdd.n2864 gnd 0.006722f
C5179 vdd.n2865 gnd 0.006722f
C5180 vdd.n2866 gnd 0.006722f
C5181 vdd.n2867 gnd 0.006722f
C5182 vdd.n2868 gnd 0.006722f
C5183 vdd.n2869 gnd 0.006722f
C5184 vdd.n2870 gnd 0.006722f
C5185 vdd.n2871 gnd 0.006722f
C5186 vdd.n2872 gnd 0.006722f
C5187 vdd.n2873 gnd 0.006722f
C5188 vdd.n2874 gnd 0.006722f
C5189 vdd.n2875 gnd 0.006722f
C5190 vdd.n2876 gnd 0.006722f
C5191 vdd.n2877 gnd 0.006722f
C5192 vdd.n2878 gnd 0.006722f
C5193 vdd.n2879 gnd 0.006722f
C5194 vdd.n2880 gnd 0.006722f
C5195 vdd.n2881 gnd 0.006722f
C5196 vdd.n2882 gnd 0.006722f
C5197 vdd.n2883 gnd 0.006722f
C5198 vdd.n2884 gnd 0.006722f
C5199 vdd.n2885 gnd 0.006722f
C5200 vdd.n2886 gnd 0.006722f
C5201 vdd.n2887 gnd 0.006722f
C5202 vdd.n2888 gnd 0.006722f
C5203 vdd.n2889 gnd 0.006722f
C5204 vdd.n2890 gnd 0.006722f
C5205 vdd.n2891 gnd 0.006722f
C5206 vdd.n2892 gnd 0.006722f
C5207 vdd.n2893 gnd 0.006722f
C5208 vdd.n2894 gnd 0.217212f
C5209 vdd.n2895 gnd 0.006722f
C5210 vdd.n2896 gnd 0.006722f
C5211 vdd.n2897 gnd 0.006722f
C5212 vdd.n2898 gnd 0.006722f
C5213 vdd.n2899 gnd 0.006722f
C5214 vdd.n2900 gnd 0.006722f
C5215 vdd.n2901 gnd 0.006722f
C5216 vdd.n2902 gnd 0.006722f
C5217 vdd.n2903 gnd 0.006722f
C5218 vdd.n2904 gnd 0.006722f
C5219 vdd.n2905 gnd 0.006722f
C5220 vdd.n2906 gnd 0.621327f
C5221 vdd.n2907 gnd 0.006722f
C5222 vdd.n2908 gnd 0.006722f
C5223 vdd.n2909 gnd 0.006722f
C5224 vdd.n2910 gnd 0.006722f
C5225 vdd.n2911 gnd 0.006722f
C5226 vdd.n2912 gnd 0.006722f
C5227 vdd.n2913 gnd 0.006722f
C5228 vdd.n2914 gnd 0.006722f
C5229 vdd.n2915 gnd 0.006722f
C5230 vdd.n2916 gnd 0.006722f
C5231 vdd.n2917 gnd 0.006722f
C5232 vdd.n2918 gnd 0.409166f
C5233 vdd.n2919 gnd 0.006722f
C5234 vdd.n2920 gnd 0.006722f
C5235 vdd.n2921 gnd 0.006722f
C5236 vdd.n2922 gnd 0.006722f
C5237 vdd.n2923 gnd 0.006722f
C5238 vdd.n2924 gnd 0.014559f
C5239 vdd.n2925 gnd 0.015494f
C5240 vdd.n2926 gnd 0.015494f
C5241 vdd.n2927 gnd 0.838538f
C5242 vdd.n2929 gnd 0.006722f
C5243 vdd.n2930 gnd 0.006722f
C5244 vdd.n2931 gnd 0.015494f
C5245 vdd.n2932 gnd 0.014559f
C5246 vdd.n2933 gnd 0.014559f
C5247 vdd.n2934 gnd 0.798127f
C5248 vdd.n2935 gnd 0.014559f
C5249 vdd.n2936 gnd 0.014559f
C5250 vdd.n2937 gnd 0.006722f
C5251 vdd.n2938 gnd 0.006722f
C5252 vdd.n2939 gnd 0.006722f
C5253 vdd.n2940 gnd 0.429372f
C5254 vdd.n2941 gnd 0.006722f
C5255 vdd.n2942 gnd 0.006722f
C5256 vdd.n2943 gnd 0.006722f
C5257 vdd.n2944 gnd 0.006722f
C5258 vdd.n2945 gnd 0.006722f
C5259 vdd.n2946 gnd 0.495041f
C5260 vdd.n2947 gnd 0.006722f
C5261 vdd.n2948 gnd 0.006722f
C5262 vdd.n2949 gnd 0.006722f
C5263 vdd.n2950 gnd 0.006722f
C5264 vdd.n2951 gnd 0.006722f
C5265 vdd.n2952 gnd 0.686995f
C5266 vdd.n2953 gnd 0.006722f
C5267 vdd.n2954 gnd 0.006722f
C5268 vdd.n2955 gnd 0.006722f
C5269 vdd.n2956 gnd 0.006722f
C5270 vdd.n2957 gnd 0.006722f
C5271 vdd.n2958 gnd 0.217212f
C5272 vdd.n2959 gnd 0.006722f
C5273 vdd.n2960 gnd 0.006722f
C5274 vdd.n2961 gnd 0.006722f
C5275 vdd.n2962 gnd 0.006722f
C5276 vdd.n2963 gnd 0.006722f
C5277 vdd.n2964 gnd 0.217212f
C5278 vdd.n2965 gnd 0.006722f
C5279 vdd.n2966 gnd 0.006722f
C5280 vdd.n2967 gnd 0.006722f
C5281 vdd.n2968 gnd 0.006722f
C5282 vdd.n2969 gnd 0.006722f
C5283 vdd.n2970 gnd 0.434423f
C5284 vdd.n2971 gnd 0.006722f
C5285 vdd.n2972 gnd 0.006722f
C5286 vdd.n2973 gnd 0.006722f
C5287 vdd.n2974 gnd 0.006722f
C5288 vdd.n2975 gnd 0.006722f
C5289 vdd.n2976 gnd 0.585967f
C5290 vdd.n2977 gnd 0.006722f
C5291 vdd.n2978 gnd 0.006722f
C5292 vdd.n2979 gnd 0.006722f
C5293 vdd.n2980 gnd 0.006722f
C5294 vdd.n2981 gnd 0.006722f
C5295 vdd.n2982 gnd 0.570812f
C5296 vdd.n2983 gnd 0.006722f
C5297 vdd.n2984 gnd 0.006722f
C5298 vdd.n2985 gnd 0.006722f
C5299 vdd.n2986 gnd 0.006722f
C5300 vdd.n2987 gnd 0.006722f
C5301 vdd.n2988 gnd 0.419269f
C5302 vdd.n2989 gnd 0.006722f
C5303 vdd.n2990 gnd 0.006722f
C5304 vdd.n2991 gnd 0.006722f
C5305 vdd.n2992 gnd 0.006722f
C5306 vdd.n2993 gnd 0.006722f
C5307 vdd.n2994 gnd 0.419269f
C5308 vdd.n2995 gnd 0.006722f
C5309 vdd.n2996 gnd 0.004548f
C5310 vdd.n2997 gnd 0.019474f
C5311 vdd.n2998 gnd 0.005536f
C5312 vdd.n2999 gnd 0.006722f
C5313 vdd.n3000 gnd 0.006722f
C5314 vdd.n3001 gnd 0.570812f
C5315 vdd.n3002 gnd 0.006722f
C5316 vdd.n3003 gnd 0.006722f
C5317 vdd.n3004 gnd 0.006722f
C5318 vdd.n3005 gnd 0.006722f
C5319 vdd.n3006 gnd 0.006722f
C5320 vdd.n3007 gnd 0.686995f
C5321 vdd.n3008 gnd 0.006722f
C5322 vdd.n3009 gnd 0.006722f
C5323 vdd.n3010 gnd 0.006722f
C5324 vdd.n3011 gnd 0.006722f
C5325 vdd.n3012 gnd 0.006722f
C5326 vdd.n3013 gnd 0.651635f
C5327 vdd.n3014 gnd 0.006722f
C5328 vdd.n3015 gnd 0.006722f
C5329 vdd.n3016 gnd 0.006722f
C5330 vdd.n3017 gnd 0.006722f
C5331 vdd.n3018 gnd 0.006722f
C5332 vdd.n3019 gnd 0.500092f
C5333 vdd.n3020 gnd 0.006722f
C5334 vdd.n3021 gnd 0.006722f
C5335 vdd.n3022 gnd 0.006722f
C5336 vdd.n3023 gnd 0.006722f
C5337 vdd.n3024 gnd 0.006722f
C5338 vdd.n3025 gnd 0.348549f
C5339 vdd.n3026 gnd 0.006722f
C5340 vdd.n3027 gnd 0.006722f
C5341 vdd.n3028 gnd 0.006722f
C5342 vdd.n3029 gnd 0.006722f
C5343 vdd.n3030 gnd 0.006722f
C5344 vdd.n3031 gnd 0.686995f
C5345 vdd.n3032 gnd 0.006722f
C5346 vdd.n3033 gnd 0.006722f
C5347 vdd.n3034 gnd 0.006722f
C5348 vdd.n3035 gnd 0.006722f
C5349 vdd.n3036 gnd 0.006722f
C5350 vdd.n3037 gnd 0.006722f
C5351 vdd.n3039 gnd 0.006722f
C5352 vdd.n3040 gnd 0.006722f
C5353 vdd.n3042 gnd 0.006722f
C5354 vdd.n3043 gnd 0.006722f
C5355 vdd.n3046 gnd 0.006722f
C5356 vdd.n3047 gnd 0.006722f
C5357 vdd.n3048 gnd 0.006722f
C5358 vdd.n3049 gnd 0.006722f
C5359 vdd.n3051 gnd 0.006722f
C5360 vdd.n3052 gnd 0.006722f
C5361 vdd.n3053 gnd 0.006722f
C5362 vdd.n3054 gnd 0.006722f
C5363 vdd.n3055 gnd 0.006722f
C5364 vdd.n3056 gnd 0.006722f
C5365 vdd.n3058 gnd 0.006722f
C5366 vdd.n3059 gnd 0.006722f
C5367 vdd.n3060 gnd 0.006722f
C5368 vdd.n3061 gnd 0.006722f
C5369 vdd.n3062 gnd 0.006722f
C5370 vdd.n3063 gnd 0.006722f
C5371 vdd.n3065 gnd 0.006722f
C5372 vdd.n3066 gnd 0.006722f
C5373 vdd.n3067 gnd 0.006722f
C5374 vdd.n3068 gnd 0.006722f
C5375 vdd.n3069 gnd 0.006722f
C5376 vdd.n3070 gnd 0.006722f
C5377 vdd.n3072 gnd 0.006722f
C5378 vdd.n3073 gnd 0.015494f
C5379 vdd.n3074 gnd 0.015494f
C5380 vdd.n3075 gnd 0.014559f
C5381 vdd.n3076 gnd 0.006722f
C5382 vdd.n3077 gnd 0.006722f
C5383 vdd.n3078 gnd 0.006722f
C5384 vdd.n3079 gnd 0.006722f
C5385 vdd.n3080 gnd 0.006722f
C5386 vdd.n3081 gnd 0.006722f
C5387 vdd.n3082 gnd 0.686995f
C5388 vdd.n3083 gnd 0.006722f
C5389 vdd.n3084 gnd 0.006722f
C5390 vdd.n3085 gnd 0.006722f
C5391 vdd.n3086 gnd 0.006722f
C5392 vdd.n3087 gnd 0.006722f
C5393 vdd.n3088 gnd 0.469784f
C5394 vdd.n3089 gnd 0.006722f
C5395 vdd.n3090 gnd 0.006722f
C5396 vdd.n3091 gnd 0.006722f
C5397 vdd.n3092 gnd 0.015411f
C5398 vdd.n3094 gnd 0.015494f
C5399 vdd.n3095 gnd 0.014642f
C5400 vdd.n3096 gnd 0.006722f
C5401 vdd.n3097 gnd 0.00519f
C5402 vdd.n3098 gnd 0.006722f
C5403 vdd.n3100 gnd 0.006722f
C5404 vdd.n3101 gnd 0.006722f
C5405 vdd.n3102 gnd 0.006722f
C5406 vdd.n3103 gnd 0.006722f
C5407 vdd.n3104 gnd 0.006722f
C5408 vdd.n3105 gnd 0.006722f
C5409 vdd.n3107 gnd 0.006722f
C5410 vdd.n3108 gnd 0.006722f
C5411 vdd.n3109 gnd 0.006722f
C5412 vdd.n3110 gnd 0.006722f
C5413 vdd.n3111 gnd 0.006722f
C5414 vdd.n3112 gnd 0.006722f
C5415 vdd.n3114 gnd 0.006722f
C5416 vdd.n3115 gnd 0.006722f
C5417 vdd.n3116 gnd 0.006722f
C5418 vdd.n3117 gnd 0.006722f
C5419 vdd.n3118 gnd 0.006722f
C5420 vdd.n3119 gnd 0.006722f
C5421 vdd.n3121 gnd 0.006722f
C5422 vdd.n3122 gnd 0.006722f
C5423 vdd.n3123 gnd 0.006722f
C5424 vdd.n3124 gnd 0.903113f
C5425 vdd.n3125 gnd 0.031555f
C5426 vdd.n3126 gnd 0.006722f
C5427 vdd.n3127 gnd 0.006722f
C5428 vdd.n3129 gnd 0.006722f
C5429 vdd.n3130 gnd 0.006722f
C5430 vdd.n3131 gnd 0.006722f
C5431 vdd.n3132 gnd 0.006722f
C5432 vdd.n3133 gnd 0.006722f
C5433 vdd.n3134 gnd 0.006722f
C5434 vdd.n3136 gnd 0.006722f
C5435 vdd.n3137 gnd 0.006722f
C5436 vdd.n3138 gnd 0.006722f
C5437 vdd.n3139 gnd 0.006722f
C5438 vdd.n3140 gnd 0.006722f
C5439 vdd.n3141 gnd 0.006722f
C5440 vdd.n3143 gnd 0.006722f
C5441 vdd.n3144 gnd 0.006722f
C5442 vdd.n3145 gnd 0.006722f
C5443 vdd.n3146 gnd 0.006722f
C5444 vdd.n3147 gnd 0.006722f
C5445 vdd.n3148 gnd 0.006722f
C5446 vdd.n3150 gnd 0.006722f
C5447 vdd.n3151 gnd 0.006722f
C5448 vdd.n3153 gnd 0.006722f
C5449 vdd.n3154 gnd 0.006722f
C5450 vdd.n3155 gnd 0.015494f
C5451 vdd.n3156 gnd 0.014559f
C5452 vdd.n3157 gnd 0.014559f
C5453 vdd.n3158 gnd 0.94967f
C5454 vdd.n3159 gnd 0.014559f
C5455 vdd.n3160 gnd 0.015494f
C5456 vdd.n3161 gnd 0.014642f
C5457 vdd.n3162 gnd 0.006722f
C5458 vdd.n3163 gnd 0.00519f
C5459 vdd.n3164 gnd 0.006722f
C5460 vdd.n3166 gnd 0.006722f
C5461 vdd.n3167 gnd 0.006722f
C5462 vdd.n3168 gnd 0.006722f
C5463 vdd.n3169 gnd 0.006722f
C5464 vdd.n3170 gnd 0.006722f
C5465 vdd.n3171 gnd 0.006722f
C5466 vdd.n3173 gnd 0.006722f
C5467 vdd.n3174 gnd 0.006722f
C5468 vdd.n3175 gnd 0.006722f
C5469 vdd.n3176 gnd 0.006722f
C5470 vdd.n3177 gnd 0.006722f
C5471 vdd.n3178 gnd 0.006722f
C5472 vdd.n3180 gnd 0.006722f
C5473 vdd.n3181 gnd 0.006722f
C5474 vdd.n3182 gnd 0.006722f
C5475 vdd.n3183 gnd 0.006722f
C5476 vdd.n3184 gnd 0.006722f
C5477 vdd.n3185 gnd 0.006722f
C5478 vdd.n3187 gnd 0.006722f
C5479 vdd.n3188 gnd 0.006722f
C5480 vdd.n3190 gnd 0.006722f
C5481 vdd.n3191 gnd 0.031555f
C5482 vdd.n3192 gnd 0.903113f
C5483 vdd.n3193 gnd 0.008502f
C5484 vdd.n3194 gnd 0.00378f
C5485 vdd.t59 gnd 0.121622f
C5486 vdd.t60 gnd 0.12998f
C5487 vdd.t58 gnd 0.158837f
C5488 vdd.n3195 gnd 0.203606f
C5489 vdd.n3196 gnd 0.171066f
C5490 vdd.n3197 gnd 0.012254f
C5491 vdd.n3198 gnd 0.009886f
C5492 vdd.n3199 gnd 0.004177f
C5493 vdd.n3200 gnd 0.007957f
C5494 vdd.n3201 gnd 0.009886f
C5495 vdd.n3202 gnd 0.009886f
C5496 vdd.n3203 gnd 0.007957f
C5497 vdd.n3204 gnd 0.007957f
C5498 vdd.n3205 gnd 0.009886f
C5499 vdd.n3207 gnd 0.009886f
C5500 vdd.n3208 gnd 0.007957f
C5501 vdd.n3209 gnd 0.007957f
C5502 vdd.n3210 gnd 0.007957f
C5503 vdd.n3211 gnd 0.009886f
C5504 vdd.n3213 gnd 0.009886f
C5505 vdd.n3215 gnd 0.009886f
C5506 vdd.n3216 gnd 0.007957f
C5507 vdd.n3217 gnd 0.007957f
C5508 vdd.n3218 gnd 0.007957f
C5509 vdd.n3219 gnd 0.009886f
C5510 vdd.n3221 gnd 0.009886f
C5511 vdd.n3223 gnd 0.009886f
C5512 vdd.n3224 gnd 0.007957f
C5513 vdd.n3225 gnd 0.007957f
C5514 vdd.n3226 gnd 0.007957f
C5515 vdd.n3227 gnd 0.009886f
C5516 vdd.n3229 gnd 0.009886f
C5517 vdd.n3230 gnd 0.009886f
C5518 vdd.n3231 gnd 0.007957f
C5519 vdd.n3232 gnd 0.007957f
C5520 vdd.n3233 gnd 0.009886f
C5521 vdd.n3234 gnd 0.009886f
C5522 vdd.n3236 gnd 0.009886f
C5523 vdd.n3237 gnd 0.007957f
C5524 vdd.n3238 gnd 0.009886f
C5525 vdd.n3239 gnd 0.009886f
C5526 vdd.n3240 gnd 0.009886f
C5527 vdd.n3241 gnd 0.016232f
C5528 vdd.n3242 gnd 0.005411f
C5529 vdd.n3243 gnd 0.009886f
C5530 vdd.n3245 gnd 0.009886f
C5531 vdd.n3247 gnd 0.009886f
C5532 vdd.n3248 gnd 0.007957f
C5533 vdd.n3249 gnd 0.007957f
C5534 vdd.n3250 gnd 0.007957f
C5535 vdd.n3251 gnd 0.009886f
C5536 vdd.n3253 gnd 0.009886f
C5537 vdd.n3255 gnd 0.009886f
C5538 vdd.n3256 gnd 0.007957f
C5539 vdd.n3257 gnd 0.007957f
C5540 vdd.n3258 gnd 0.007957f
C5541 vdd.n3259 gnd 0.009886f
C5542 vdd.n3261 gnd 0.009886f
C5543 vdd.n3263 gnd 0.009886f
C5544 vdd.n3264 gnd 0.007957f
C5545 vdd.n3265 gnd 0.007957f
C5546 vdd.n3266 gnd 0.007957f
C5547 vdd.n3267 gnd 0.009886f
C5548 vdd.n3269 gnd 0.009886f
C5549 vdd.n3271 gnd 0.009886f
C5550 vdd.n3272 gnd 0.007957f
C5551 vdd.n3273 gnd 0.007957f
C5552 vdd.n3274 gnd 0.007957f
C5553 vdd.n3275 gnd 0.009886f
C5554 vdd.n3277 gnd 0.009886f
C5555 vdd.n3279 gnd 0.009886f
C5556 vdd.n3280 gnd 0.007957f
C5557 vdd.n3281 gnd 0.007957f
C5558 vdd.n3282 gnd 0.006644f
C5559 vdd.n3283 gnd 0.009886f
C5560 vdd.n3285 gnd 0.009886f
C5561 vdd.n3287 gnd 0.009886f
C5562 vdd.n3288 gnd 0.006644f
C5563 vdd.n3289 gnd 0.007957f
C5564 vdd.n3290 gnd 0.007957f
C5565 vdd.n3291 gnd 0.009886f
C5566 vdd.n3293 gnd 0.009886f
C5567 vdd.n3295 gnd 0.009886f
C5568 vdd.n3296 gnd 0.007957f
C5569 vdd.n3297 gnd 0.007957f
C5570 vdd.n3298 gnd 0.007957f
C5571 vdd.n3299 gnd 0.009886f
C5572 vdd.n3301 gnd 0.009886f
C5573 vdd.n3303 gnd 0.009886f
C5574 vdd.n3304 gnd 0.007957f
C5575 vdd.n3305 gnd 0.007957f
C5576 vdd.n3306 gnd 0.007957f
C5577 vdd.n3307 gnd 0.009886f
C5578 vdd.n3309 gnd 0.009886f
C5579 vdd.n3310 gnd 0.009886f
C5580 vdd.n3311 gnd 0.007957f
C5581 vdd.n3312 gnd 0.007957f
C5582 vdd.n3313 gnd 0.009886f
C5583 vdd.n3314 gnd 0.009886f
C5584 vdd.n3315 gnd 0.007957f
C5585 vdd.n3316 gnd 0.007957f
C5586 vdd.n3317 gnd 0.009886f
C5587 vdd.n3318 gnd 0.009886f
C5588 vdd.n3320 gnd 0.009886f
C5589 vdd.n3321 gnd 0.007957f
C5590 vdd.n3322 gnd 0.006604f
C5591 vdd.n3323 gnd 0.022666f
C5592 vdd.n3324 gnd 0.022512f
C5593 vdd.n3325 gnd 0.006604f
C5594 vdd.n3326 gnd 0.022512f
C5595 vdd.n3327 gnd 1.33358f
C5596 vdd.n3328 gnd 0.022512f
C5597 vdd.n3329 gnd 0.006604f
C5598 vdd.n3330 gnd 0.022512f
C5599 vdd.n3331 gnd 0.009886f
C5600 vdd.n3332 gnd 0.009886f
C5601 vdd.n3333 gnd 0.007957f
C5602 vdd.n3334 gnd 0.009886f
C5603 vdd.n3335 gnd 0.954721f
C5604 vdd.n3336 gnd 0.009886f
C5605 vdd.n3337 gnd 0.007957f
C5606 vdd.n3338 gnd 0.009886f
C5607 vdd.n3339 gnd 0.009886f
C5608 vdd.n3340 gnd 0.009886f
C5609 vdd.n3341 gnd 0.007957f
C5610 vdd.n3342 gnd 0.009886f
C5611 vdd.n3343 gnd 0.98503f
C5612 vdd.n3344 gnd 0.009886f
C5613 vdd.n3345 gnd 0.007957f
C5614 vdd.n3346 gnd 0.009886f
C5615 vdd.n3347 gnd 0.009886f
C5616 vdd.n3348 gnd 0.009886f
C5617 vdd.n3349 gnd 0.007957f
C5618 vdd.n3350 gnd 0.009886f
C5619 vdd.t138 gnd 0.505144f
C5620 vdd.n3351 gnd 0.813281f
C5621 vdd.n3352 gnd 0.009886f
C5622 vdd.n3353 gnd 0.007957f
C5623 vdd.n3354 gnd 0.009886f
C5624 vdd.n3355 gnd 0.009886f
C5625 vdd.n3356 gnd 0.009886f
C5626 vdd.n3357 gnd 0.007957f
C5627 vdd.n3358 gnd 0.009886f
C5628 vdd.n3359 gnd 0.641532f
C5629 vdd.n3360 gnd 0.009886f
C5630 vdd.n3361 gnd 0.007957f
C5631 vdd.n3362 gnd 0.009886f
C5632 vdd.n3363 gnd 0.009886f
C5633 vdd.n3364 gnd 0.009886f
C5634 vdd.n3365 gnd 0.007957f
C5635 vdd.n3366 gnd 0.009886f
C5636 vdd.n3367 gnd 0.803178f
C5637 vdd.n3368 gnd 0.540504f
C5638 vdd.n3369 gnd 0.009886f
C5639 vdd.n3370 gnd 0.007957f
C5640 vdd.n3371 gnd 0.009886f
C5641 vdd.n3372 gnd 0.009886f
C5642 vdd.n3373 gnd 0.009886f
C5643 vdd.n3374 gnd 0.007957f
C5644 vdd.n3375 gnd 0.009886f
C5645 vdd.n3376 gnd 0.712252f
C5646 vdd.n3377 gnd 0.009886f
C5647 vdd.n3378 gnd 0.007957f
C5648 vdd.n3379 gnd 0.009886f
C5649 vdd.n3380 gnd 0.009886f
C5650 vdd.n3381 gnd 0.009886f
C5651 vdd.n3382 gnd 0.009886f
C5652 vdd.n3383 gnd 0.009886f
C5653 vdd.n3384 gnd 0.007957f
C5654 vdd.n3385 gnd 0.007957f
C5655 vdd.n3386 gnd 0.009886f
C5656 vdd.t149 gnd 0.505144f
C5657 vdd.n3387 gnd 0.838538f
C5658 vdd.n3388 gnd 0.009886f
C5659 vdd.n3389 gnd 0.007957f
C5660 vdd.n3390 gnd 0.009886f
C5661 vdd.n3391 gnd 0.009886f
C5662 vdd.n3392 gnd 0.009886f
C5663 vdd.n3393 gnd 0.007957f
C5664 vdd.n3394 gnd 0.009886f
C5665 vdd.n3395 gnd 0.793075f
C5666 vdd.n3396 gnd 0.009886f
C5667 vdd.n3397 gnd 0.009886f
C5668 vdd.n3398 gnd 0.007957f
C5669 vdd.n3399 gnd 0.007957f
C5670 vdd.n3400 gnd 0.007957f
C5671 vdd.n3401 gnd 0.009886f
C5672 vdd.n3402 gnd 0.009886f
C5673 vdd.n3403 gnd 0.009886f
C5674 vdd.n3404 gnd 0.009886f
C5675 vdd.n3405 gnd 0.007957f
C5676 vdd.n3406 gnd 0.007957f
C5677 vdd.n3407 gnd 0.007957f
C5678 vdd.n3408 gnd 0.009886f
C5679 vdd.n3409 gnd 0.009886f
C5680 vdd.n3410 gnd 0.009886f
C5681 vdd.n3411 gnd 0.009886f
C5682 vdd.n3412 gnd 0.007957f
C5683 vdd.n3413 gnd 0.007957f
C5684 vdd.n3414 gnd 0.007957f
C5685 vdd.n3415 gnd 0.009886f
C5686 vdd.n3416 gnd 0.009886f
C5687 vdd.n3417 gnd 0.009886f
C5688 vdd.n3418 gnd 0.838538f
C5689 vdd.n3419 gnd 0.009886f
C5690 vdd.n3420 gnd 0.007957f
C5691 vdd.n3421 gnd 0.007957f
C5692 vdd.n3422 gnd 0.007957f
C5693 vdd.n3423 gnd 0.009886f
C5694 vdd.n3424 gnd 0.009886f
C5695 vdd.n3425 gnd 0.009886f
C5696 vdd.n3426 gnd 0.009886f
C5697 vdd.n3427 gnd 0.007957f
C5698 vdd.n3428 gnd 0.007957f
C5699 vdd.n3429 gnd 0.006604f
C5700 vdd.n3430 gnd 0.022512f
C5701 vdd.n3431 gnd 0.022666f
C5702 vdd.n3432 gnd 0.00378f
C5703 vdd.n3433 gnd 0.022666f
C5704 vdd.n3435 gnd 2.23273f
C5705 vdd.n3436 gnd 1.33358f
C5706 vdd.n3437 gnd 0.661738f
C5707 vdd.n3438 gnd 0.009886f
C5708 vdd.n3439 gnd 0.007957f
C5709 vdd.n3440 gnd 0.007957f
C5710 vdd.n3441 gnd 0.007957f
C5711 vdd.n3442 gnd 0.009886f
C5712 vdd.n3443 gnd 1.01029f
C5713 vdd.n3444 gnd 1.01029f
C5714 vdd.n3445 gnd 0.580915f
C5715 vdd.n3446 gnd 0.009886f
C5716 vdd.n3447 gnd 0.007957f
C5717 vdd.n3448 gnd 0.007957f
C5718 vdd.n3449 gnd 0.007957f
C5719 vdd.n3450 gnd 0.009886f
C5720 vdd.n3451 gnd 0.601121f
C5721 vdd.n3452 gnd 0.742561f
C5722 vdd.t180 gnd 0.505144f
C5723 vdd.n3453 gnd 0.77287f
C5724 vdd.n3454 gnd 0.009886f
C5725 vdd.n3455 gnd 0.007957f
C5726 vdd.n3456 gnd 0.007957f
C5727 vdd.n3457 gnd 0.007957f
C5728 vdd.n3458 gnd 0.009886f
C5729 vdd.n3459 gnd 0.838538f
C5730 vdd.t191 gnd 0.505144f
C5731 vdd.n3460 gnd 0.611224f
C5732 vdd.n3461 gnd 0.732458f
C5733 vdd.n3462 gnd 0.009886f
C5734 vdd.n3463 gnd 0.007957f
C5735 vdd.n3464 gnd 0.007957f
C5736 vdd.n3465 gnd 0.007957f
C5737 vdd.n3466 gnd 0.009886f
C5738 vdd.n3467 gnd 0.560709f
C5739 vdd.t145 gnd 0.505144f
C5740 vdd.n3468 gnd 0.838538f
C5741 vdd.t223 gnd 0.505144f
C5742 vdd.n3469 gnd 0.621327f
C5743 vdd.n3470 gnd 0.009886f
C5744 vdd.n3471 gnd 0.007957f
C5745 vdd.n3472 gnd 0.007598f
C5746 vdd.n3473 gnd 0.583105f
C5747 vdd.n3474 gnd 2.59295f
C5748 a_n8300_8799.n0 gnd 0.211582f
C5749 a_n8300_8799.n1 gnd 0.295727f
C5750 a_n8300_8799.n2 gnd 0.211582f
C5751 a_n8300_8799.n3 gnd 0.211582f
C5752 a_n8300_8799.n4 gnd 0.211582f
C5753 a_n8300_8799.n5 gnd 0.27875f
C5754 a_n8300_8799.n6 gnd 0.211582f
C5755 a_n8300_8799.n7 gnd 0.295727f
C5756 a_n8300_8799.n8 gnd 0.211582f
C5757 a_n8300_8799.n9 gnd 0.211582f
C5758 a_n8300_8799.n10 gnd 0.211582f
C5759 a_n8300_8799.n11 gnd 0.27875f
C5760 a_n8300_8799.n12 gnd 0.211582f
C5761 a_n8300_8799.n13 gnd 0.463461f
C5762 a_n8300_8799.n14 gnd 0.211582f
C5763 a_n8300_8799.n15 gnd 0.211582f
C5764 a_n8300_8799.n16 gnd 0.211582f
C5765 a_n8300_8799.n17 gnd 0.27875f
C5766 a_n8300_8799.n18 gnd 0.331646f
C5767 a_n8300_8799.n19 gnd 0.211582f
C5768 a_n8300_8799.n20 gnd 0.211582f
C5769 a_n8300_8799.n21 gnd 0.211582f
C5770 a_n8300_8799.n22 gnd 0.211582f
C5771 a_n8300_8799.n23 gnd 0.242831f
C5772 a_n8300_8799.n24 gnd 0.331646f
C5773 a_n8300_8799.n25 gnd 0.211582f
C5774 a_n8300_8799.n26 gnd 0.211582f
C5775 a_n8300_8799.n27 gnd 0.211582f
C5776 a_n8300_8799.n28 gnd 0.211582f
C5777 a_n8300_8799.n29 gnd 0.242831f
C5778 a_n8300_8799.n30 gnd 0.331646f
C5779 a_n8300_8799.n31 gnd 0.211582f
C5780 a_n8300_8799.n32 gnd 0.211582f
C5781 a_n8300_8799.n33 gnd 0.211582f
C5782 a_n8300_8799.n34 gnd 0.211582f
C5783 a_n8300_8799.n35 gnd 0.410566f
C5784 a_n8300_8799.n36 gnd 3.47236f
C5785 a_n8300_8799.n37 gnd 1.77052f
C5786 a_n8300_8799.n38 gnd 3.01244f
C5787 a_n8300_8799.n39 gnd 1.55073f
C5788 a_n8300_8799.n40 gnd 4.00706f
C5789 a_n8300_8799.n41 gnd 1.55073f
C5790 a_n8300_8799.n42 gnd 2.82921f
C5791 a_n8300_8799.n43 gnd 0.712333f
C5792 a_n8300_8799.n44 gnd 0.008776f
C5793 a_n8300_8799.n45 gnd 0.001178f
C5794 a_n8300_8799.n47 gnd 0.007881f
C5795 a_n8300_8799.n48 gnd 0.011912f
C5796 a_n8300_8799.n49 gnd 0.008192f
C5797 a_n8300_8799.n51 gnd 4.09e-19
C5798 a_n8300_8799.n52 gnd 0.00849f
C5799 a_n8300_8799.n53 gnd 0.011726f
C5800 a_n8300_8799.n54 gnd 0.007556f
C5801 a_n8300_8799.n55 gnd 0.008776f
C5802 a_n8300_8799.n56 gnd 0.001178f
C5803 a_n8300_8799.n58 gnd 0.007881f
C5804 a_n8300_8799.n59 gnd 0.011912f
C5805 a_n8300_8799.n60 gnd 0.008192f
C5806 a_n8300_8799.n62 gnd 4.09e-19
C5807 a_n8300_8799.n63 gnd 0.00849f
C5808 a_n8300_8799.n64 gnd 0.011726f
C5809 a_n8300_8799.n65 gnd 0.007556f
C5810 a_n8300_8799.n66 gnd 0.008776f
C5811 a_n8300_8799.n67 gnd 0.001178f
C5812 a_n8300_8799.n69 gnd 0.007881f
C5813 a_n8300_8799.n70 gnd 0.011912f
C5814 a_n8300_8799.n71 gnd 0.008192f
C5815 a_n8300_8799.n73 gnd 4.09e-19
C5816 a_n8300_8799.n74 gnd 0.00849f
C5817 a_n8300_8799.n75 gnd 0.011726f
C5818 a_n8300_8799.n76 gnd 0.007556f
C5819 a_n8300_8799.n77 gnd 0.001178f
C5820 a_n8300_8799.n79 gnd 0.007881f
C5821 a_n8300_8799.n80 gnd 0.011912f
C5822 a_n8300_8799.n81 gnd 0.008192f
C5823 a_n8300_8799.n83 gnd 4.09e-19
C5824 a_n8300_8799.n84 gnd 0.00849f
C5825 a_n8300_8799.n85 gnd 0.011726f
C5826 a_n8300_8799.n86 gnd 0.007556f
C5827 a_n8300_8799.n87 gnd 0.254725f
C5828 a_n8300_8799.n88 gnd 0.001178f
C5829 a_n8300_8799.n90 gnd 0.007881f
C5830 a_n8300_8799.n91 gnd 0.011912f
C5831 a_n8300_8799.n92 gnd 0.008192f
C5832 a_n8300_8799.n94 gnd 4.09e-19
C5833 a_n8300_8799.n95 gnd 0.00849f
C5834 a_n8300_8799.n96 gnd 0.011726f
C5835 a_n8300_8799.n97 gnd 0.007556f
C5836 a_n8300_8799.n98 gnd 0.254725f
C5837 a_n8300_8799.n99 gnd 0.001178f
C5838 a_n8300_8799.n101 gnd 0.007881f
C5839 a_n8300_8799.n102 gnd 0.011912f
C5840 a_n8300_8799.n103 gnd 0.008192f
C5841 a_n8300_8799.n105 gnd 4.09e-19
C5842 a_n8300_8799.n106 gnd 0.00849f
C5843 a_n8300_8799.n107 gnd 0.011726f
C5844 a_n8300_8799.n108 gnd 0.007556f
C5845 a_n8300_8799.n109 gnd 0.254725f
C5846 a_n8300_8799.t1 gnd 0.146756f
C5847 a_n8300_8799.t37 gnd 0.146756f
C5848 a_n8300_8799.t6 gnd 0.146756f
C5849 a_n8300_8799.n110 gnd 1.15749f
C5850 a_n8300_8799.t20 gnd 0.146756f
C5851 a_n8300_8799.t29 gnd 0.146756f
C5852 a_n8300_8799.n111 gnd 1.15558f
C5853 a_n8300_8799.t27 gnd 0.146756f
C5854 a_n8300_8799.t12 gnd 0.146756f
C5855 a_n8300_8799.n112 gnd 1.15558f
C5856 a_n8300_8799.t26 gnd 0.146756f
C5857 a_n8300_8799.t2 gnd 0.146756f
C5858 a_n8300_8799.n113 gnd 1.15748f
C5859 a_n8300_8799.t13 gnd 0.146756f
C5860 a_n8300_8799.t5 gnd 0.146756f
C5861 a_n8300_8799.n114 gnd 1.15558f
C5862 a_n8300_8799.t34 gnd 0.146756f
C5863 a_n8300_8799.t35 gnd 0.146756f
C5864 a_n8300_8799.n115 gnd 1.15558f
C5865 a_n8300_8799.t11 gnd 0.146756f
C5866 a_n8300_8799.t15 gnd 0.146756f
C5867 a_n8300_8799.n116 gnd 1.15558f
C5868 a_n8300_8799.t28 gnd 0.146756f
C5869 a_n8300_8799.t30 gnd 0.146756f
C5870 a_n8300_8799.n117 gnd 1.15558f
C5871 a_n8300_8799.t3 gnd 0.114143f
C5872 a_n8300_8799.t33 gnd 0.114143f
C5873 a_n8300_8799.n118 gnd 1.01022f
C5874 a_n8300_8799.t24 gnd 0.114143f
C5875 a_n8300_8799.t17 gnd 0.114143f
C5876 a_n8300_8799.n119 gnd 1.00861f
C5877 a_n8300_8799.t18 gnd 0.114143f
C5878 a_n8300_8799.t25 gnd 0.114143f
C5879 a_n8300_8799.n120 gnd 1.00861f
C5880 a_n8300_8799.t8 gnd 0.114143f
C5881 a_n8300_8799.t36 gnd 0.114143f
C5882 a_n8300_8799.n121 gnd 1.01022f
C5883 a_n8300_8799.t38 gnd 0.114143f
C5884 a_n8300_8799.t10 gnd 0.114143f
C5885 a_n8300_8799.n122 gnd 1.00861f
C5886 a_n8300_8799.t43 gnd 0.114143f
C5887 a_n8300_8799.t21 gnd 0.114143f
C5888 a_n8300_8799.n123 gnd 1.00861f
C5889 a_n8300_8799.t9 gnd 0.114143f
C5890 a_n8300_8799.t19 gnd 0.114143f
C5891 a_n8300_8799.n124 gnd 1.01022f
C5892 a_n8300_8799.t22 gnd 0.114143f
C5893 a_n8300_8799.t40 gnd 0.114143f
C5894 a_n8300_8799.n125 gnd 1.00861f
C5895 a_n8300_8799.t7 gnd 0.114143f
C5896 a_n8300_8799.t23 gnd 0.114143f
C5897 a_n8300_8799.n126 gnd 1.00861f
C5898 a_n8300_8799.t41 gnd 0.114143f
C5899 a_n8300_8799.t31 gnd 0.114143f
C5900 a_n8300_8799.n127 gnd 1.00861f
C5901 a_n8300_8799.t39 gnd 0.114143f
C5902 a_n8300_8799.t14 gnd 0.114143f
C5903 a_n8300_8799.n128 gnd 1.00861f
C5904 a_n8300_8799.t42 gnd 0.114143f
C5905 a_n8300_8799.t32 gnd 0.114143f
C5906 a_n8300_8799.n129 gnd 1.00861f
C5907 a_n8300_8799.t68 gnd 0.608518f
C5908 a_n8300_8799.n130 gnd 0.272053f
C5909 a_n8300_8799.t102 gnd 0.608518f
C5910 a_n8300_8799.t122 gnd 0.608518f
C5911 a_n8300_8799.n131 gnd 0.275424f
C5912 a_n8300_8799.t79 gnd 0.608518f
C5913 a_n8300_8799.t81 gnd 0.608518f
C5914 a_n8300_8799.t93 gnd 0.608518f
C5915 a_n8300_8799.n132 gnd 0.277546f
C5916 a_n8300_8799.t123 gnd 0.608518f
C5917 a_n8300_8799.t128 gnd 0.608518f
C5918 a_n8300_8799.n133 gnd 0.270961f
C5919 a_n8300_8799.t96 gnd 0.620035f
C5920 a_n8300_8799.n134 gnd 0.255117f
C5921 a_n8300_8799.n135 gnd 0.012003f
C5922 a_n8300_8799.t66 gnd 0.608518f
C5923 a_n8300_8799.n136 gnd 0.271776f
C5924 a_n8300_8799.n137 gnd 0.275409f
C5925 a_n8300_8799.t124 gnd 0.608518f
C5926 a_n8300_8799.n138 gnd 0.271867f
C5927 a_n8300_8799.n139 gnd 0.266395f
C5928 a_n8300_8799.t105 gnd 0.608518f
C5929 a_n8300_8799.n140 gnd 0.271613f
C5930 a_n8300_8799.n141 gnd 0.277989f
C5931 a_n8300_8799.t80 gnd 0.608518f
C5932 a_n8300_8799.n142 gnd 0.275289f
C5933 a_n8300_8799.n143 gnd 0.271287f
C5934 a_n8300_8799.t67 gnd 0.608518f
C5935 a_n8300_8799.n144 gnd 0.266721f
C5936 a_n8300_8799.t99 gnd 0.608518f
C5937 a_n8300_8799.n145 gnd 0.275408f
C5938 a_n8300_8799.t44 gnd 0.620025f
C5939 a_n8300_8799.t78 gnd 0.608518f
C5940 a_n8300_8799.n146 gnd 0.272053f
C5941 a_n8300_8799.t117 gnd 0.608518f
C5942 a_n8300_8799.t134 gnd 0.608518f
C5943 a_n8300_8799.n147 gnd 0.275424f
C5944 a_n8300_8799.t85 gnd 0.608518f
C5945 a_n8300_8799.t89 gnd 0.608518f
C5946 a_n8300_8799.t103 gnd 0.608518f
C5947 a_n8300_8799.n148 gnd 0.277546f
C5948 a_n8300_8799.t136 gnd 0.608518f
C5949 a_n8300_8799.t139 gnd 0.608518f
C5950 a_n8300_8799.n149 gnd 0.270961f
C5951 a_n8300_8799.t109 gnd 0.620035f
C5952 a_n8300_8799.n150 gnd 0.255117f
C5953 a_n8300_8799.n151 gnd 0.012003f
C5954 a_n8300_8799.t74 gnd 0.608518f
C5955 a_n8300_8799.n152 gnd 0.271776f
C5956 a_n8300_8799.n153 gnd 0.275409f
C5957 a_n8300_8799.t138 gnd 0.608518f
C5958 a_n8300_8799.n154 gnd 0.271867f
C5959 a_n8300_8799.n155 gnd 0.266395f
C5960 a_n8300_8799.t119 gnd 0.608518f
C5961 a_n8300_8799.n156 gnd 0.271613f
C5962 a_n8300_8799.n157 gnd 0.277989f
C5963 a_n8300_8799.t86 gnd 0.608518f
C5964 a_n8300_8799.n158 gnd 0.275289f
C5965 a_n8300_8799.n159 gnd 0.271287f
C5966 a_n8300_8799.t77 gnd 0.608518f
C5967 a_n8300_8799.n160 gnd 0.266721f
C5968 a_n8300_8799.t115 gnd 0.608518f
C5969 a_n8300_8799.n161 gnd 0.275408f
C5970 a_n8300_8799.t52 gnd 0.620025f
C5971 a_n8300_8799.n162 gnd 0.916496f
C5972 a_n8300_8799.t104 gnd 0.608518f
C5973 a_n8300_8799.n163 gnd 0.272053f
C5974 a_n8300_8799.t90 gnd 0.608518f
C5975 a_n8300_8799.t125 gnd 0.608518f
C5976 a_n8300_8799.n164 gnd 0.275424f
C5977 a_n8300_8799.t58 gnd 0.608518f
C5978 a_n8300_8799.t118 gnd 0.608518f
C5979 a_n8300_8799.t53 gnd 0.608518f
C5980 a_n8300_8799.n165 gnd 0.277546f
C5981 a_n8300_8799.t100 gnd 0.608518f
C5982 a_n8300_8799.t70 gnd 0.608518f
C5983 a_n8300_8799.n166 gnd 0.270961f
C5984 a_n8300_8799.t111 gnd 0.620035f
C5985 a_n8300_8799.n167 gnd 0.255117f
C5986 a_n8300_8799.n168 gnd 0.012003f
C5987 a_n8300_8799.t87 gnd 0.608518f
C5988 a_n8300_8799.n169 gnd 0.271776f
C5989 a_n8300_8799.n170 gnd 0.275409f
C5990 a_n8300_8799.t83 gnd 0.608518f
C5991 a_n8300_8799.n171 gnd 0.271867f
C5992 a_n8300_8799.n172 gnd 0.266395f
C5993 a_n8300_8799.t75 gnd 0.608518f
C5994 a_n8300_8799.n173 gnd 0.271613f
C5995 a_n8300_8799.n174 gnd 0.277989f
C5996 a_n8300_8799.t45 gnd 0.608518f
C5997 a_n8300_8799.n175 gnd 0.275289f
C5998 a_n8300_8799.n176 gnd 0.271287f
C5999 a_n8300_8799.t127 gnd 0.608518f
C6000 a_n8300_8799.n177 gnd 0.266721f
C6001 a_n8300_8799.t133 gnd 0.608518f
C6002 a_n8300_8799.n178 gnd 0.275408f
C6003 a_n8300_8799.t84 gnd 0.620025f
C6004 a_n8300_8799.n179 gnd 1.73585f
C6005 a_n8300_8799.t94 gnd 0.608518f
C6006 a_n8300_8799.t47 gnd 0.608518f
C6007 a_n8300_8799.t98 gnd 0.608518f
C6008 a_n8300_8799.n180 gnd 0.275003f
C6009 a_n8300_8799.t97 gnd 0.608518f
C6010 a_n8300_8799.t49 gnd 0.608518f
C6011 a_n8300_8799.t48 gnd 0.608518f
C6012 a_n8300_8799.n181 gnd 0.271867f
C6013 a_n8300_8799.t116 gnd 0.608518f
C6014 a_n8300_8799.t61 gnd 0.608518f
C6015 a_n8300_8799.t51 gnd 0.608518f
C6016 a_n8300_8799.n182 gnd 0.275424f
C6017 a_n8300_8799.t120 gnd 0.608518f
C6018 a_n8300_8799.t82 gnd 0.608518f
C6019 a_n8300_8799.t62 gnd 0.608518f
C6020 a_n8300_8799.n183 gnd 0.271287f
C6021 a_n8300_8799.t137 gnd 0.608518f
C6022 a_n8300_8799.t95 gnd 0.608518f
C6023 a_n8300_8799.t64 gnd 0.608518f
C6024 a_n8300_8799.n184 gnd 0.275408f
C6025 a_n8300_8799.t131 gnd 0.620035f
C6026 a_n8300_8799.n185 gnd 0.255117f
C6027 a_n8300_8799.n186 gnd 0.272053f
C6028 a_n8300_8799.n187 gnd 0.266721f
C6029 a_n8300_8799.n188 gnd 0.275289f
C6030 a_n8300_8799.n189 gnd 0.277989f
C6031 a_n8300_8799.n190 gnd 0.271613f
C6032 a_n8300_8799.n191 gnd 0.266395f
C6033 a_n8300_8799.n192 gnd 0.275409f
C6034 a_n8300_8799.n193 gnd 0.277546f
C6035 a_n8300_8799.n194 gnd 0.270961f
C6036 a_n8300_8799.n195 gnd 0.266232f
C6037 a_n8300_8799.t107 gnd 0.608518f
C6038 a_n8300_8799.t55 gnd 0.608518f
C6039 a_n8300_8799.t114 gnd 0.608518f
C6040 a_n8300_8799.n196 gnd 0.275003f
C6041 a_n8300_8799.t113 gnd 0.608518f
C6042 a_n8300_8799.t57 gnd 0.608518f
C6043 a_n8300_8799.t56 gnd 0.608518f
C6044 a_n8300_8799.n197 gnd 0.271867f
C6045 a_n8300_8799.t130 gnd 0.608518f
C6046 a_n8300_8799.t69 gnd 0.608518f
C6047 a_n8300_8799.t60 gnd 0.608518f
C6048 a_n8300_8799.n198 gnd 0.275424f
C6049 a_n8300_8799.t132 gnd 0.608518f
C6050 a_n8300_8799.t92 gnd 0.608518f
C6051 a_n8300_8799.t72 gnd 0.608518f
C6052 a_n8300_8799.n199 gnd 0.271287f
C6053 a_n8300_8799.t50 gnd 0.608518f
C6054 a_n8300_8799.t108 gnd 0.608518f
C6055 a_n8300_8799.t73 gnd 0.608518f
C6056 a_n8300_8799.n200 gnd 0.275408f
C6057 a_n8300_8799.t46 gnd 0.620035f
C6058 a_n8300_8799.n201 gnd 0.255117f
C6059 a_n8300_8799.n202 gnd 0.272053f
C6060 a_n8300_8799.n203 gnd 0.266721f
C6061 a_n8300_8799.n204 gnd 0.275289f
C6062 a_n8300_8799.n205 gnd 0.277989f
C6063 a_n8300_8799.n206 gnd 0.271613f
C6064 a_n8300_8799.n207 gnd 0.266395f
C6065 a_n8300_8799.n208 gnd 0.275409f
C6066 a_n8300_8799.n209 gnd 0.277546f
C6067 a_n8300_8799.n210 gnd 0.270961f
C6068 a_n8300_8799.n211 gnd 0.266232f
C6069 a_n8300_8799.n212 gnd 0.916496f
C6070 a_n8300_8799.t65 gnd 0.608518f
C6071 a_n8300_8799.t135 gnd 0.608518f
C6072 a_n8300_8799.t106 gnd 0.608518f
C6073 a_n8300_8799.n213 gnd 0.275003f
C6074 a_n8300_8799.t129 gnd 0.608518f
C6075 a_n8300_8799.t91 gnd 0.608518f
C6076 a_n8300_8799.t112 gnd 0.608518f
C6077 a_n8300_8799.n214 gnd 0.271867f
C6078 a_n8300_8799.t59 gnd 0.608518f
C6079 a_n8300_8799.t126 gnd 0.608518f
C6080 a_n8300_8799.t76 gnd 0.608518f
C6081 a_n8300_8799.n215 gnd 0.275424f
C6082 a_n8300_8799.t121 gnd 0.608518f
C6083 a_n8300_8799.t63 gnd 0.608518f
C6084 a_n8300_8799.t101 gnd 0.608518f
C6085 a_n8300_8799.n216 gnd 0.271287f
C6086 a_n8300_8799.t54 gnd 0.608518f
C6087 a_n8300_8799.t88 gnd 0.608518f
C6088 a_n8300_8799.t71 gnd 0.608518f
C6089 a_n8300_8799.n217 gnd 0.275408f
C6090 a_n8300_8799.t110 gnd 0.620035f
C6091 a_n8300_8799.n218 gnd 0.255117f
C6092 a_n8300_8799.n219 gnd 0.272053f
C6093 a_n8300_8799.n220 gnd 0.266721f
C6094 a_n8300_8799.n221 gnd 0.275289f
C6095 a_n8300_8799.n222 gnd 0.277989f
C6096 a_n8300_8799.n223 gnd 0.271613f
C6097 a_n8300_8799.n224 gnd 0.266395f
C6098 a_n8300_8799.n225 gnd 0.275409f
C6099 a_n8300_8799.n226 gnd 0.277546f
C6100 a_n8300_8799.n227 gnd 0.270961f
C6101 a_n8300_8799.n228 gnd 0.266232f
C6102 a_n8300_8799.n229 gnd 1.33515f
C6103 a_n8300_8799.n230 gnd 15.9687f
C6104 a_n8300_8799.n231 gnd 4.45347f
C6105 a_n8300_8799.n232 gnd 7.1166f
C6106 a_n8300_8799.t4 gnd 0.146756f
C6107 a_n8300_8799.t16 gnd 0.146756f
C6108 a_n8300_8799.n233 gnd 1.15558f
C6109 a_n8300_8799.n234 gnd 1.15558f
C6110 a_n8300_8799.t0 gnd 0.146756f
.ends

