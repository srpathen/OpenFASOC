* NGSPICE file created from opamp461.ext - technology: sky130A

.subckt opamp461 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 a_n8300_8799.t43 plus.t5 a_n3827_n3924.t28 gnd.t167 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X1 CSoutput.t97 a_n8300_8799.t44 vdd.t138 vdd.t95 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X2 a_n2472_13878.t27 a_n2650_13878.t11 a_n2650_13878.t12 vdd.t258 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 a_n2472_13878.t7 a_n2650_13878.t64 vdd.t140 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 gnd.t291 gnd.t289 gnd.t290 gnd.t241 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X5 vdd.t136 a_n8300_8799.t45 CSoutput.t96 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X6 outputibias.t7 outputibias.t6 gnd.t151 gnd.t150 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X7 gnd.t288 gnd.t286 minus.t4 gnd.t287 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X8 CSoutput.t95 a_n8300_8799.t46 vdd.t137 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X9 a_n3827_n3924.t15 diffpairibias.t20 gnd.t154 gnd.t153 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X10 gnd.t156 commonsourceibias.t80 CSoutput.t139 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X11 gnd.t285 gnd.t283 gnd.t284 gnd.t261 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X12 CSoutput.t94 a_n8300_8799.t47 vdd.t135 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X13 commonsourceibias.t79 commonsourceibias.t78 gnd.t155 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X14 a_n3827_n3924.t27 plus.t6 a_n8300_8799.t42 gnd.t338 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X15 commonsourceibias.t77 commonsourceibias.t76 gnd.t35 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X16 gnd.t282 gnd.t280 gnd.t281 gnd.t261 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X17 a_n3827_n3924.t5 minus.t5 a_n2650_13878.t2 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X18 a_n2650_8322.t25 a_n2650_13878.t65 a_n8300_8799.t1 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X19 vdd.t227 CSoutput.t176 output.t15 gnd.t48 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X20 gnd.t279 gnd.t277 gnd.t278 gnd.t196 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X21 CSoutput.t140 commonsourceibias.t81 gnd.t158 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X22 CSoutput.t93 a_n8300_8799.t48 vdd.t134 vdd.t57 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X23 gnd.t93 commonsourceibias.t74 commonsourceibias.t75 gnd.t86 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X24 CSoutput.t104 commonsourceibias.t82 gnd.t52 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X25 vdd.t133 a_n8300_8799.t49 CSoutput.t92 vdd.t84 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X26 gnd.t276 gnd.t274 gnd.t275 gnd.t196 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X27 a_n2650_13878.t0 minus.t6 a_n3827_n3924.t0 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X28 commonsourceibias.t73 commonsourceibias.t72 gnd.t94 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X29 vdd.t228 CSoutput.t177 output.t14 gnd.t49 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X30 a_n8300_8799.t17 a_n2650_13878.t66 a_n2650_8322.t24 vdd.t268 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X31 CSoutput.t105 commonsourceibias.t83 gnd.t54 gnd.t53 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 vdd.t132 a_n8300_8799.t50 CSoutput.t91 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X33 a_n2650_13878.t1 minus.t7 a_n3827_n3924.t4 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X34 vdd.t131 a_n8300_8799.t51 CSoutput.t90 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X35 a_n8300_8799.t18 a_n2650_13878.t67 a_n2650_8322.t23 vdd.t269 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X36 gnd.t273 gnd.t270 gnd.t272 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X37 commonsourceibias.t71 commonsourceibias.t70 gnd.t141 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X38 a_n3827_n3924.t10 minus.t8 a_n2650_13878.t47 gnd.t114 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X39 CSoutput.t89 a_n8300_8799.t52 vdd.t130 vdd.t95 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X40 a_n3827_n3924.t2 diffpairibias.t21 gnd.t4 gnd.t3 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X41 CSoutput.t164 commonsourceibias.t84 gnd.t323 gnd.t146 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X42 CSoutput.t88 a_n8300_8799.t53 vdd.t129 vdd.t69 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X43 gnd.t324 commonsourceibias.t85 CSoutput.t165 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X44 vdd.t128 a_n8300_8799.t54 CSoutput.t87 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X45 gnd.t269 gnd.t267 gnd.t268 gnd.t188 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X46 gnd.t308 commonsourceibias.t68 commonsourceibias.t69 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X47 CSoutput.t86 a_n8300_8799.t55 vdd.t127 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X48 commonsourceibias.t67 commonsourceibias.t66 gnd.t309 gnd.t132 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X49 a_n3827_n3924.t26 plus.t7 a_n8300_8799.t41 gnd.t166 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X50 vdd.t219 vdd.t217 vdd.t218 vdd.t153 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X51 gnd.t139 commonsourceibias.t86 CSoutput.t137 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 a_n2472_13878.t26 a_n2650_13878.t5 a_n2650_13878.t6 vdd.t262 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X53 a_n8300_8799.t40 plus.t8 a_n3827_n3924.t43 gnd.t337 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X54 gnd.t140 commonsourceibias.t87 CSoutput.t138 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X55 a_n2650_13878.t42 a_n2650_13878.t41 a_n2472_13878.t25 vdd.t263 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X56 gnd.t306 commonsourceibias.t88 CSoutput.t158 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X57 a_n8300_8799.t39 plus.t9 a_n3827_n3924.t42 gnd.t336 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X58 CSoutput.t85 a_n8300_8799.t56 vdd.t126 vdd.t57 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X59 vdd.t216 vdd.t214 vdd.t215 vdd.t191 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X60 output.t13 CSoutput.t178 vdd.t229 gnd.t50 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X61 vdd.t114 a_n8300_8799.t57 CSoutput.t84 vdd.t84 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X62 gnd.t163 commonsourceibias.t64 commonsourceibias.t65 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X63 diffpairibias.t19 diffpairibias.t18 gnd.t67 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X64 a_n3827_n3924.t41 plus.t10 a_n8300_8799.t38 gnd.t335 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X65 commonsourceibias.t63 commonsourceibias.t62 gnd.t161 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X66 a_n2650_13878.t63 minus.t9 a_n3827_n3924.t56 gnd.t331 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X67 a_n2650_13878.t40 a_n2650_13878.t39 a_n2472_13878.t24 vdd.t237 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X68 a_n8300_8799.t19 a_n2650_13878.t68 a_n2650_8322.t22 vdd.t259 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X69 CSoutput.t83 a_n8300_8799.t58 vdd.t125 vdd.t93 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X70 commonsourceibias.t61 commonsourceibias.t60 gnd.t95 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X71 gnd.t266 gnd.t264 plus.t4 gnd.t265 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X72 a_n2650_13878.t30 a_n2650_13878.t29 a_n2472_13878.t23 vdd.t253 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X73 vdd.t124 a_n8300_8799.t59 CSoutput.t82 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X74 vdd.t123 a_n8300_8799.t60 CSoutput.t81 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X75 a_n8300_8799.t8 a_n2650_13878.t69 a_n2650_8322.t21 vdd.t252 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X76 gnd.t263 gnd.t260 gnd.t262 gnd.t261 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X77 diffpairibias.t17 diffpairibias.t16 gnd.t319 gnd.t318 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X78 gnd.t142 commonsourceibias.t58 commonsourceibias.t59 gnd.t128 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X79 CSoutput.t80 a_n8300_8799.t61 vdd.t121 vdd.t38 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X80 CSoutput.t159 commonsourceibias.t89 gnd.t307 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X81 a_n2650_8322.t20 a_n2650_13878.t70 a_n8300_8799.t9 vdd.t253 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X82 CSoutput.t135 commonsourceibias.t90 gnd.t137 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X83 vdd.t213 vdd.t211 vdd.t212 vdd.t178 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X84 CSoutput.t79 a_n8300_8799.t62 vdd.t122 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X85 gnd.t144 commonsourceibias.t56 commonsourceibias.t57 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X86 vdd.t3 CSoutput.t179 output.t12 gnd.t14 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X87 CSoutput.t136 commonsourceibias.t91 gnd.t138 gnd.t132 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 CSoutput.t119 commonsourceibias.t92 gnd.t91 gnd.t90 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 gnd.t259 gnd.t257 gnd.t258 gnd.t203 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X90 gnd.t256 gnd.t254 plus.t3 gnd.t255 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X91 a_n3827_n3924.t40 plus.t11 a_n8300_8799.t37 gnd.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X92 CSoutput.t120 commonsourceibias.t93 gnd.t92 gnd.t55 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X93 CSoutput.t156 commonsourceibias.t94 gnd.t304 gnd.t53 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 a_n3827_n3924.t3 diffpairibias.t22 gnd.t6 gnd.t5 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X95 vdd.t120 a_n8300_8799.t63 CSoutput.t78 vdd.t82 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X96 vdd.t119 a_n8300_8799.t64 CSoutput.t77 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X97 a_n2650_13878.t10 a_n2650_13878.t9 a_n2472_13878.t22 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X98 vdd.t118 a_n8300_8799.t65 CSoutput.t76 vdd.t63 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X99 vdd.t117 a_n8300_8799.t66 CSoutput.t75 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X100 output.t11 CSoutput.t180 vdd.t4 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X101 a_n8300_8799.t10 a_n2650_13878.t71 a_n2650_8322.t19 vdd.t254 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X102 a_n2650_13878.t36 a_n2650_13878.t35 a_n2472_13878.t21 vdd.t223 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X103 gnd.t170 commonsourceibias.t54 commonsourceibias.t55 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X104 gnd.t361 commonsourceibias.t52 commonsourceibias.t53 gnd.t123 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X105 gnd.t356 commonsourceibias.t50 commonsourceibias.t51 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X106 output.t19 outputibias.t8 gnd.t22 gnd.t21 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X107 CSoutput.t181 a_n2650_8322.t5 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X108 vdd.t116 a_n8300_8799.t67 CSoutput.t74 vdd.t36 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X109 CSoutput.t73 a_n8300_8799.t68 vdd.t115 vdd.t67 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X110 gnd.t253 gnd.t250 gnd.t252 gnd.t251 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X111 diffpairibias.t15 diffpairibias.t14 gnd.t165 gnd.t164 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X112 a_n2650_13878.t60 minus.t10 a_n3827_n3924.t52 gnd.t330 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X113 output.t18 outputibias.t9 gnd.t175 gnd.t174 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X114 vdd.t210 vdd.t208 vdd.t209 vdd.t195 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X115 CSoutput.t72 a_n8300_8799.t69 vdd.t113 vdd.t38 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X116 gnd.t305 commonsourceibias.t95 CSoutput.t157 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X117 vdd.t207 vdd.t204 vdd.t206 vdd.t205 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X118 gnd.t302 commonsourceibias.t96 CSoutput.t154 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X119 gnd.t303 commonsourceibias.t97 CSoutput.t155 gnd.t128 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X120 gnd.t134 commonsourceibias.t98 CSoutput.t133 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X121 a_n3827_n3924.t49 minus.t11 a_n2650_13878.t57 gnd.t329 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X122 CSoutput.t71 a_n8300_8799.t70 vdd.t112 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X123 gnd.t136 commonsourceibias.t99 CSoutput.t134 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X124 output.t10 CSoutput.t182 vdd.t5 gnd.t16 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X125 vdd.t111 a_n8300_8799.t71 CSoutput.t70 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X126 vdd.t142 CSoutput.t183 output.t9 gnd.t33 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X127 vdd.t241 a_n2650_13878.t72 a_n2650_8322.t33 vdd.t240 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X128 a_n2650_13878.t26 a_n2650_13878.t25 a_n2472_13878.t20 vdd.t260 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X129 gnd.t87 commonsourceibias.t100 CSoutput.t117 gnd.t86 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X130 vdd.t203 vdd.t201 vdd.t202 vdd.t178 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X131 vdd.t200 vdd.t198 vdd.t199 vdd.t171 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X132 gnd.t249 gnd.t247 gnd.t248 gnd.t207 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X133 a_n2650_8322.t32 a_n2650_13878.t73 vdd.t243 vdd.t242 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X134 a_n3827_n3924.t20 diffpairibias.t23 gnd.t296 gnd.t295 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X135 CSoutput.t69 a_n8300_8799.t72 vdd.t110 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X136 CSoutput.t118 commonsourceibias.t101 gnd.t89 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X137 a_n3827_n3924.t13 minus.t12 a_n2650_13878.t49 gnd.t118 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X138 a_n3827_n3924.t7 minus.t13 a_n2650_13878.t44 gnd.t68 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X139 gnd.t74 commonsourceibias.t48 commonsourceibias.t49 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X140 vdd.t245 a_n2650_13878.t74 a_n2472_13878.t6 vdd.t244 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X141 a_n2650_13878.t45 minus.t14 a_n3827_n3924.t8 gnd.t110 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X142 a_n3827_n3924.t44 plus.t12 a_n8300_8799.t36 gnd.t334 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X143 a_n3827_n3924.t35 plus.t13 a_n8300_8799.t35 gnd.t294 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X144 gnd.t85 commonsourceibias.t102 CSoutput.t116 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X145 vdd.t197 vdd.t194 vdd.t196 vdd.t195 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X146 a_n2650_13878.t50 minus.t15 a_n3827_n3924.t14 gnd.t152 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X147 vdd.t109 a_n8300_8799.t73 CSoutput.t68 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X148 vdd.t107 a_n8300_8799.t74 CSoutput.t67 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X149 gnd.t315 commonsourceibias.t46 commonsourceibias.t47 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X150 gnd.t246 gnd.t244 plus.t2 gnd.t245 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X151 a_n8300_8799.t34 plus.t14 a_n3827_n3924.t39 gnd.t333 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X152 a_n8300_8799.t33 plus.t15 a_n3827_n3924.t36 gnd.t332 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X153 vdd.t193 vdd.t190 vdd.t192 vdd.t191 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X154 a_n2650_8322.t31 a_n2650_13878.t75 vdd.t256 vdd.t255 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X155 a_n8300_8799.t11 a_n2650_13878.t76 a_n2650_8322.t18 vdd.t257 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X156 CSoutput.t66 a_n8300_8799.t75 vdd.t106 vdd.t46 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X157 diffpairibias.t13 diffpairibias.t12 gnd.t342 gnd.t341 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X158 CSoutput.t184 a_n2650_8322.t4 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X159 vdd.t105 a_n8300_8799.t76 CSoutput.t65 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X160 CSoutput.t101 commonsourceibias.t103 gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X161 a_n2650_13878.t46 minus.t16 a_n3827_n3924.t9 gnd.t113 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X162 a_n2650_13878.t34 a_n2650_13878.t33 a_n2472_13878.t19 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X163 vdd.t103 a_n8300_8799.t77 CSoutput.t64 vdd.t36 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X164 a_n8300_8799.t12 a_n2650_13878.t77 a_n2650_8322.t17 vdd.t258 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X165 CSoutput.t63 a_n8300_8799.t78 vdd.t102 vdd.t67 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X166 CSoutput.t132 commonsourceibias.t104 gnd.t133 gnd.t132 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X167 a_n2472_13878.t18 a_n2650_13878.t23 a_n2650_13878.t24 vdd.t254 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X168 commonsourceibias.t45 commonsourceibias.t44 gnd.t182 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X169 CSoutput.t153 commonsourceibias.t105 gnd.t301 gnd.t90 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X170 gnd.t131 commonsourceibias.t106 CSoutput.t131 gnd.t130 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X171 a_n3827_n3924.t6 minus.t17 a_n2650_13878.t43 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X172 CSoutput.t115 commonsourceibias.t107 gnd.t83 gnd.t55 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X173 vdd.t143 CSoutput.t185 output.t8 gnd.t34 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X174 CSoutput.t152 commonsourceibias.t108 gnd.t300 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X175 gnd.t61 commonsourceibias.t109 CSoutput.t107 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X176 CSoutput.t62 a_n8300_8799.t79 vdd.t101 vdd.t93 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X177 gnd.t183 commonsourceibias.t42 commonsourceibias.t43 gnd.t125 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X178 gnd.t243 gnd.t240 gnd.t242 gnd.t241 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X179 vdd.t236 a_n2650_13878.t78 a_n2650_8322.t30 vdd.t235 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X180 a_n2472_13878.t17 a_n2650_13878.t15 a_n2650_13878.t16 vdd.t268 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X181 gnd.t82 commonsourceibias.t110 CSoutput.t114 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X182 vdd.t100 a_n8300_8799.t80 CSoutput.t61 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X183 vdd.t189 vdd.t187 vdd.t188 vdd.t171 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X184 a_n2650_13878.t22 a_n2650_13878.t21 a_n2472_13878.t16 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X185 commonsourceibias.t41 commonsourceibias.t40 gnd.t76 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X186 gnd.t326 commonsourceibias.t38 commonsourceibias.t39 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X187 minus.t3 gnd.t237 gnd.t239 gnd.t238 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X188 a_n3827_n3924.t34 plus.t16 a_n8300_8799.t32 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X189 vdd.t99 a_n8300_8799.t81 CSoutput.t60 vdd.t48 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X190 gnd.t58 commonsourceibias.t36 commonsourceibias.t37 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X191 a_n3827_n3924.t53 diffpairibias.t24 gnd.t360 gnd.t359 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X192 commonsourceibias.t35 commonsourceibias.t34 gnd.t106 gnd.t53 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X193 a_n3827_n3924.t1 diffpairibias.t25 gnd.t2 gnd.t1 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X194 gnd.t299 commonsourceibias.t111 CSoutput.t151 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X195 vdd.t98 a_n8300_8799.t82 CSoutput.t59 vdd.t82 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X196 a_n8300_8799.t31 plus.t17 a_n3827_n3924.t38 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X197 gnd.t298 commonsourceibias.t112 CSoutput.t150 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X198 gnd.t129 commonsourceibias.t113 CSoutput.t130 gnd.t128 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X199 gnd.t80 commonsourceibias.t114 CSoutput.t113 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X200 gnd.t127 commonsourceibias.t115 CSoutput.t129 gnd.t86 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X201 a_n2472_13878.t15 a_n2650_13878.t7 a_n2650_13878.t8 vdd.t261 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X202 vdd.t186 vdd.t184 vdd.t185 vdd.t149 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X203 CSoutput.t186 a_n2650_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X204 CSoutput.t112 commonsourceibias.t116 gnd.t78 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X205 a_n2650_8322.t16 a_n2650_13878.t79 a_n8300_8799.t5 vdd.t237 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X206 CSoutput.t58 a_n8300_8799.t83 vdd.t97 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X207 commonsourceibias.t33 commonsourceibias.t32 gnd.t172 gnd.t171 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X208 CSoutput.t149 commonsourceibias.t117 gnd.t297 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X209 CSoutput.t57 a_n8300_8799.t84 vdd.t96 vdd.t95 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X210 CSoutput.t187 a_n2650_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X211 gnd.t60 commonsourceibias.t118 CSoutput.t106 gnd.t59 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X212 CSoutput.t111 commonsourceibias.t119 gnd.t72 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X213 gnd.t236 gnd.t234 gnd.t235 gnd.t188 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X214 diffpairibias.t11 diffpairibias.t10 gnd.t112 gnd.t111 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X215 a_n2472_13878.t5 a_n2650_13878.t80 vdd.t239 vdd.t238 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X216 gnd.t314 commonsourceibias.t120 CSoutput.t162 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X217 vdd.t231 a_n2650_13878.t81 a_n2472_13878.t4 vdd.t230 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X218 output.t17 outputibias.t10 gnd.t293 gnd.t292 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X219 gnd.t37 commonsourceibias.t30 commonsourceibias.t31 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X220 CSoutput.t56 a_n8300_8799.t85 vdd.t94 vdd.t93 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X221 gnd.t357 commonsourceibias.t28 commonsourceibias.t29 gnd.t130 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X222 vdd.t92 a_n8300_8799.t86 CSoutput.t55 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X223 commonsourceibias.t27 commonsourceibias.t26 gnd.t64 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X224 vdd.t90 a_n8300_8799.t87 CSoutput.t54 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X225 CSoutput.t110 commonsourceibias.t121 gnd.t71 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X226 CSoutput.t53 a_n8300_8799.t88 vdd.t88 vdd.t61 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X227 plus.t1 gnd.t231 gnd.t233 gnd.t232 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X228 a_n2472_13878.t14 a_n2650_13878.t27 a_n2650_13878.t28 vdd.t259 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X229 diffpairibias.t9 diffpairibias.t8 gnd.t340 gnd.t339 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X230 a_n3827_n3924.t17 minus.t18 a_n2650_13878.t51 gnd.t166 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X231 vdd.t87 a_n8300_8799.t89 CSoutput.t52 vdd.t48 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X232 gnd.t18 commonsourceibias.t24 commonsourceibias.t25 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X233 CSoutput.t148 commonsourceibias.t122 gnd.t181 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X234 a_n2650_13878.t62 minus.t19 a_n3827_n3924.t55 gnd.t337 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X235 a_n2650_8322.t15 a_n2650_13878.t82 a_n8300_8799.t4 vdd.t232 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X236 CSoutput.t51 a_n8300_8799.t90 vdd.t86 vdd.t50 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X237 diffpairibias.t7 diffpairibias.t6 gnd.t101 gnd.t100 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X238 vdd.t85 a_n8300_8799.t91 CSoutput.t50 vdd.t84 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X239 a_n2472_13878.t13 a_n2650_13878.t31 a_n2650_13878.t32 vdd.t252 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X240 a_n2650_13878.t56 minus.t20 a_n3827_n3924.t48 gnd.t336 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X241 a_n2650_13878.t52 minus.t21 a_n3827_n3924.t18 gnd.t167 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X242 gnd.t313 commonsourceibias.t123 CSoutput.t161 gnd.t130 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X243 vdd.t183 vdd.t181 vdd.t182 vdd.t160 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X244 vdd.t234 a_n2650_13878.t83 a_n2650_8322.t29 vdd.t233 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X245 vdd.t83 a_n8300_8799.t92 CSoutput.t49 vdd.t82 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X246 a_n3827_n3924.t51 minus.t22 a_n2650_13878.t59 gnd.t335 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X247 vdd.t270 CSoutput.t188 output.t7 gnd.t321 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X248 CSoutput.t109 commonsourceibias.t124 gnd.t70 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X249 a_n8300_8799.t30 plus.t18 a_n3827_n3924.t45 gnd.t331 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X250 CSoutput.t147 commonsourceibias.t125 gnd.t180 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X251 gnd.t230 gnd.t227 gnd.t229 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X252 gnd.t312 commonsourceibias.t126 CSoutput.t160 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X253 a_n3827_n3924.t54 minus.t23 a_n2650_13878.t61 gnd.t338 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X254 CSoutput.t48 a_n8300_8799.t93 vdd.t81 vdd.t69 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X255 gnd.t226 gnd.t223 gnd.t225 gnd.t224 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X256 gnd.t351 commonsourceibias.t127 CSoutput.t173 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X257 a_n2472_13878.t3 a_n2650_13878.t84 vdd.t7 vdd.t6 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X258 vdd.t180 vdd.t177 vdd.t179 vdd.t178 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X259 CSoutput.t103 commonsourceibias.t128 gnd.t44 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X260 vdd.t176 vdd.t174 vdd.t175 vdd.t160 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X261 commonsourceibias.t23 commonsourceibias.t22 gnd.t56 gnd.t55 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X262 CSoutput.t1 commonsourceibias.t129 gnd.t10 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X263 vdd.t80 a_n8300_8799.t94 CSoutput.t47 vdd.t63 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X264 CSoutput.t46 a_n8300_8799.t95 vdd.t79 vdd.t61 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X265 gnd.t222 gnd.t220 minus.t2 gnd.t221 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X266 gnd.t219 gnd.t217 gnd.t218 gnd.t207 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X267 vdd.t78 a_n8300_8799.t96 CSoutput.t45 vdd.t13 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X268 a_n3827_n3924.t21 diffpairibias.t26 gnd.t317 gnd.t316 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X269 a_n2650_8322.t14 a_n2650_13878.t85 a_n8300_8799.t0 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X270 vdd.t10 a_n2650_13878.t86 a_n2650_8322.t28 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X271 gnd.t62 commonsourceibias.t130 CSoutput.t108 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X272 CSoutput.t44 a_n8300_8799.t97 vdd.t77 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 vdd.t173 vdd.t170 vdd.t172 vdd.t171 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X274 vdd.t169 vdd.t167 vdd.t168 vdd.t145 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X275 vdd.t76 a_n8300_8799.t98 CSoutput.t43 vdd.t54 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X276 vdd.t75 a_n8300_8799.t99 CSoutput.t42 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X277 a_n8300_8799.t29 plus.t19 a_n3827_n3924.t31 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X278 gnd.t355 commonsourceibias.t131 CSoutput.t175 gnd.t123 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X279 CSoutput.t100 commonsourceibias.t132 gnd.t30 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X280 vdd.t166 vdd.t163 vdd.t165 vdd.t164 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X281 CSoutput.t142 commonsourceibias.t133 gnd.t169 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X282 a_n3827_n3924.t23 plus.t20 a_n8300_8799.t28 gnd.t114 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X283 vdd.t74 a_n8300_8799.t100 CSoutput.t41 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X284 CSoutput.t40 a_n8300_8799.t101 vdd.t73 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X285 gnd.t105 commonsourceibias.t134 CSoutput.t122 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X286 gnd.t325 commonsourceibias.t135 CSoutput.t166 gnd.t59 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X287 a_n2472_13878.t12 a_n2650_13878.t3 a_n2650_13878.t4 vdd.t249 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X288 CSoutput.t39 a_n8300_8799.t102 vdd.t71 vdd.t50 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X289 vdd.t271 CSoutput.t189 output.t6 gnd.t322 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X290 CSoutput.t146 commonsourceibias.t136 gnd.t179 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X291 a_n2650_8322.t13 a_n2650_13878.t87 a_n8300_8799.t16 vdd.t263 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X292 vdd.t162 vdd.t159 vdd.t161 vdd.t160 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X293 vdd.t158 vdd.t156 vdd.t157 vdd.t145 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X294 diffpairibias.t5 diffpairibias.t4 gnd.t344 gnd.t343 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X295 commonsourceibias.t21 commonsourceibias.t20 gnd.t39 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X296 gnd.t216 gnd.t213 gnd.t215 gnd.t214 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X297 gnd.t20 commonsourceibias.t137 CSoutput.t98 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X298 CSoutput.t145 commonsourceibias.t138 gnd.t178 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X299 gnd.t97 commonsourceibias.t18 commonsourceibias.t19 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X300 CSoutput.t38 a_n8300_8799.t103 vdd.t70 vdd.t69 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X301 CSoutput.t37 a_n8300_8799.t104 vdd.t68 vdd.t67 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X302 CSoutput.t36 a_n8300_8799.t105 vdd.t66 vdd.t46 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X303 a_n3827_n3924.t57 diffpairibias.t27 gnd.t363 gnd.t362 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X304 vdd.t65 a_n8300_8799.t106 CSoutput.t35 vdd.t54 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X305 CSoutput.t102 commonsourceibias.t139 gnd.t43 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X306 CSoutput.t190 a_n2650_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X307 vdd.t64 a_n8300_8799.t107 CSoutput.t34 vdd.t63 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X308 a_n2650_8322.t27 a_n2650_13878.t88 vdd.t265 vdd.t264 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X309 CSoutput.t33 a_n8300_8799.t108 vdd.t62 vdd.t61 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X310 CSoutput.t0 commonsourceibias.t140 gnd.t8 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X311 vdd.t60 a_n8300_8799.t109 CSoutput.t32 vdd.t13 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X312 CSoutput.t31 a_n8300_8799.t110 vdd.t59 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X313 vdd.t267 a_n2650_13878.t89 a_n2472_13878.t2 vdd.t266 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X314 gnd.t99 commonsourceibias.t16 commonsourceibias.t17 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X315 output.t16 outputibias.t11 gnd.t24 gnd.t23 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X316 plus.t0 gnd.t210 gnd.t212 gnd.t211 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X317 vdd.t14 a_n8300_8799.t111 CSoutput.t30 vdd.t13 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X318 CSoutput.t29 a_n8300_8799.t112 vdd.t58 vdd.t57 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X319 CSoutput.t163 commonsourceibias.t141 gnd.t320 gnd.t171 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X320 CSoutput.t28 a_n8300_8799.t113 vdd.t56 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X321 gnd.t126 commonsourceibias.t142 CSoutput.t128 gnd.t125 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X322 a_n3827_n3924.t24 plus.t21 a_n8300_8799.t27 gnd.t68 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X323 vdd.t55 a_n8300_8799.t114 CSoutput.t27 vdd.t54 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X324 vdd.t53 a_n8300_8799.t115 CSoutput.t26 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X325 CSoutput.t174 commonsourceibias.t143 gnd.t354 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X326 commonsourceibias.t15 commonsourceibias.t14 gnd.t145 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X327 a_n3827_n3924.t50 minus.t24 a_n2650_13878.t58 gnd.t334 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X328 a_n2650_8322.t12 a_n2650_13878.t90 a_n8300_8799.t6 vdd.t248 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X329 commonsourceibias.t13 commonsourceibias.t12 gnd.t310 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X330 a_n8300_8799.t7 a_n2650_13878.t91 a_n2650_8322.t11 vdd.t249 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X331 CSoutput.t99 commonsourceibias.t144 gnd.t28 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X332 gnd.t107 commonsourceibias.t10 commonsourceibias.t11 gnd.t59 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X333 output.t5 CSoutput.t191 vdd.t224 gnd.t45 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X334 a_n8300_8799.t26 plus.t22 a_n3827_n3924.t22 gnd.t152 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X335 a_n2472_13878.t1 a_n2650_13878.t92 vdd.t251 vdd.t250 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X336 gnd.t168 commonsourceibias.t145 CSoutput.t141 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X337 CSoutput.t121 commonsourceibias.t146 gnd.t104 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X338 vdd.t155 vdd.t152 vdd.t154 vdd.t153 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X339 vdd.t52 a_n8300_8799.t116 CSoutput.t25 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X340 vdd.t151 vdd.t148 vdd.t150 vdd.t149 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X341 a_n2650_13878.t55 minus.t25 a_n3827_n3924.t47 gnd.t333 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X342 CSoutput.t24 a_n8300_8799.t117 vdd.t51 vdd.t50 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X343 gnd.t209 gnd.t206 gnd.t208 gnd.t207 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X344 vdd.t147 vdd.t144 vdd.t146 vdd.t145 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X345 a_n8300_8799.t13 a_n2650_13878.t93 a_n2650_8322.t10 vdd.t261 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X346 commonsourceibias.t9 commonsourceibias.t8 gnd.t173 gnd.t90 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X347 a_n2650_8322.t9 a_n2650_13878.t94 a_n8300_8799.t14 vdd.t260 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X348 a_n8300_8799.t25 plus.t23 a_n3827_n3924.t25 gnd.t113 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X349 gnd.t205 gnd.t202 gnd.t204 gnd.t203 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X350 gnd.t201 gnd.t199 minus.t1 gnd.t200 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X351 a_n3827_n3924.t12 minus.t26 a_n2650_13878.t48 gnd.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X352 vdd.t49 a_n8300_8799.t118 CSoutput.t23 vdd.t48 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X353 CSoutput.t22 a_n8300_8799.t119 vdd.t47 vdd.t46 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X354 CSoutput.t21 a_n8300_8799.t120 vdd.t45 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X355 gnd.t41 commonsourceibias.t6 commonsourceibias.t7 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X356 CSoutput.t20 a_n8300_8799.t121 vdd.t44 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X357 a_n2472_13878.t11 a_n2650_13878.t37 a_n2650_13878.t38 vdd.t257 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X358 commonsourceibias.t5 commonsourceibias.t4 gnd.t358 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X359 a_n3827_n3924.t37 plus.t24 a_n8300_8799.t24 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X360 vdd.t43 a_n8300_8799.t122 CSoutput.t19 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X361 gnd.t124 commonsourceibias.t147 CSoutput.t127 gnd.t123 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X362 CSoutput.t144 commonsourceibias.t148 gnd.t177 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X363 CSoutput.t192 a_n2650_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X364 output.t4 CSoutput.t193 vdd.t225 gnd.t46 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X365 gnd.t176 commonsourceibias.t149 CSoutput.t143 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X366 a_n3827_n3924.t11 diffpairibias.t28 gnd.t116 gnd.t115 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X367 vdd.t42 a_n8300_8799.t123 CSoutput.t18 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X368 gnd.t122 commonsourceibias.t150 CSoutput.t126 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X369 CSoutput.t17 a_n8300_8799.t124 vdd.t41 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X370 a_n2650_13878.t14 a_n2650_13878.t13 a_n2472_13878.t10 vdd.t248 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X371 gnd.t198 gnd.t195 gnd.t197 gnd.t196 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X372 a_n8300_8799.t15 a_n2650_13878.t95 a_n2650_8322.t8 vdd.t262 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X373 vdd.t40 a_n8300_8799.t125 CSoutput.t16 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X374 output.t3 CSoutput.t194 vdd.t226 gnd.t47 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X375 gnd.t121 commonsourceibias.t151 CSoutput.t125 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X376 CSoutput.t15 a_n8300_8799.t126 vdd.t39 vdd.t38 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X377 a_n8300_8799.t23 plus.t25 a_n3827_n3924.t33 gnd.t330 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X378 vdd.t0 CSoutput.t195 output.t2 gnd.t11 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X379 gnd.t194 gnd.t191 gnd.t193 gnd.t192 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X380 CSoutput.t124 commonsourceibias.t152 gnd.t120 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X381 CSoutput.t123 commonsourceibias.t153 gnd.t119 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X382 commonsourceibias.t3 commonsourceibias.t2 gnd.t311 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X383 outputibias.t5 outputibias.t4 gnd.t353 gnd.t352 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X384 diffpairibias.t3 diffpairibias.t2 gnd.t103 gnd.t102 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X385 vdd.t37 a_n8300_8799.t127 CSoutput.t14 vdd.t36 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X386 CSoutput.t13 a_n8300_8799.t128 vdd.t35 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X387 CSoutput.t12 a_n8300_8799.t129 vdd.t34 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X388 a_n2650_8322.t7 a_n2650_13878.t96 a_n8300_8799.t2 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X389 a_n3827_n3924.t32 plus.t26 a_n8300_8799.t22 gnd.t329 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X390 vdd.t32 a_n8300_8799.t130 CSoutput.t11 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X391 outputibias.t3 outputibias.t2 gnd.t109 gnd.t108 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X392 CSoutput.t10 a_n8300_8799.t131 vdd.t30 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X393 diffpairibias.t1 diffpairibias.t0 gnd.t328 gnd.t327 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X394 a_n3827_n3924.t29 plus.t27 a_n8300_8799.t21 gnd.t118 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X395 CSoutput.t172 commonsourceibias.t154 gnd.t350 gnd.t171 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X396 outputibias.t1 outputibias.t0 gnd.t149 gnd.t148 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X397 vdd.t222 a_n2650_13878.t97 a_n2472_13878.t0 vdd.t221 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X398 gnd.t349 commonsourceibias.t155 CSoutput.t171 gnd.t125 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X399 a_n8300_8799.t20 plus.t28 a_n3827_n3924.t30 gnd.t110 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X400 CSoutput.t9 a_n8300_8799.t132 vdd.t28 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X401 a_n3827_n3924.t19 minus.t27 a_n2650_13878.t53 gnd.t294 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X402 vdd.t26 a_n8300_8799.t133 CSoutput.t8 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X403 vdd.t24 a_n8300_8799.t134 CSoutput.t7 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X404 CSoutput.t170 commonsourceibias.t156 gnd.t348 gnd.t146 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X405 CSoutput.t6 a_n8300_8799.t135 vdd.t22 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X406 output.t1 CSoutput.t196 vdd.t1 gnd.t12 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X407 gnd.t345 commonsourceibias.t157 CSoutput.t167 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X408 gnd.t190 gnd.t187 gnd.t189 gnd.t188 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X409 a_n2650_13878.t54 minus.t28 a_n3827_n3924.t46 gnd.t332 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X410 gnd.t347 commonsourceibias.t158 CSoutput.t169 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X411 a_n2650_8322.t6 a_n2650_13878.t98 a_n8300_8799.t3 vdd.t223 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X412 vdd.t20 a_n8300_8799.t136 CSoutput.t5 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X413 vdd.t18 a_n8300_8799.t137 CSoutput.t4 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X414 CSoutput.t3 a_n8300_8799.t138 vdd.t16 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X415 output.t0 CSoutput.t197 vdd.t2 gnd.t13 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X416 gnd.t346 commonsourceibias.t159 CSoutput.t168 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X417 a_n2650_8322.t26 a_n2650_13878.t99 vdd.t247 vdd.t246 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X418 a_n2472_13878.t9 a_n2650_13878.t17 a_n2650_13878.t18 vdd.t269 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X419 minus.t0 gnd.t184 gnd.t186 gnd.t185 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X420 commonsourceibias.t1 commonsourceibias.t0 gnd.t147 gnd.t146 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X421 a_n3827_n3924.t16 diffpairibias.t29 gnd.t160 gnd.t159 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X422 CSoutput.t2 a_n8300_8799.t139 vdd.t12 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X423 a_n2650_13878.t20 a_n2650_13878.t19 a_n2472_13878.t8 vdd.t232 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 plus.n53 plus.t20 323.478
R1 plus.n11 plus.t15 323.478
R2 plus.n52 plus.t19 297.12
R3 plus.n56 plus.t26 297.12
R4 plus.n58 plus.t25 297.12
R5 plus.n62 plus.t27 297.12
R6 plus.n64 plus.t9 297.12
R7 plus.n68 plus.t7 297.12
R8 plus.n70 plus.t14 297.12
R9 plus.n74 plus.t12 297.12
R10 plus.n76 plus.t28 297.12
R11 plus.n80 plus.t10 297.12
R12 plus.n82 plus.t8 297.12
R13 plus.n40 plus.t21 297.12
R14 plus.n38 plus.t22 297.12
R15 plus.n2 plus.t16 297.12
R16 plus.n32 plus.t17 297.12
R17 plus.n4 plus.t11 297.12
R18 plus.n26 plus.t5 297.12
R19 plus.n6 plus.t6 297.12
R20 plus.n20 plus.t23 297.12
R21 plus.n8 plus.t24 297.12
R22 plus.n14 plus.t18 297.12
R23 plus.n10 plus.t13 297.12
R24 plus.n86 plus.t2 243.97
R25 plus.n86 plus.n85 223.454
R26 plus.n88 plus.n87 223.454
R27 plus.n83 plus.n82 161.3
R28 plus.n81 plus.n42 161.3
R29 plus.n80 plus.n79 161.3
R30 plus.n78 plus.n43 161.3
R31 plus.n77 plus.n76 161.3
R32 plus.n75 plus.n44 161.3
R33 plus.n74 plus.n73 161.3
R34 plus.n72 plus.n45 161.3
R35 plus.n71 plus.n70 161.3
R36 plus.n69 plus.n46 161.3
R37 plus.n68 plus.n67 161.3
R38 plus.n66 plus.n47 161.3
R39 plus.n65 plus.n64 161.3
R40 plus.n63 plus.n48 161.3
R41 plus.n62 plus.n61 161.3
R42 plus.n60 plus.n49 161.3
R43 plus.n59 plus.n58 161.3
R44 plus.n57 plus.n50 161.3
R45 plus.n56 plus.n55 161.3
R46 plus.n54 plus.n51 161.3
R47 plus.n13 plus.n12 161.3
R48 plus.n14 plus.n9 161.3
R49 plus.n16 plus.n15 161.3
R50 plus.n17 plus.n8 161.3
R51 plus.n19 plus.n18 161.3
R52 plus.n20 plus.n7 161.3
R53 plus.n22 plus.n21 161.3
R54 plus.n23 plus.n6 161.3
R55 plus.n25 plus.n24 161.3
R56 plus.n26 plus.n5 161.3
R57 plus.n28 plus.n27 161.3
R58 plus.n29 plus.n4 161.3
R59 plus.n31 plus.n30 161.3
R60 plus.n32 plus.n3 161.3
R61 plus.n34 plus.n33 161.3
R62 plus.n35 plus.n2 161.3
R63 plus.n37 plus.n36 161.3
R64 plus.n38 plus.n1 161.3
R65 plus.n39 plus.n0 161.3
R66 plus.n41 plus.n40 161.3
R67 plus.n82 plus.n81 46.0096
R68 plus.n40 plus.n39 46.0096
R69 plus.n54 plus.n53 45.0871
R70 plus.n12 plus.n11 45.0871
R71 plus.n52 plus.n51 41.6278
R72 plus.n80 plus.n43 41.6278
R73 plus.n38 plus.n37 41.6278
R74 plus.n13 plus.n10 41.6278
R75 plus.n57 plus.n56 37.246
R76 plus.n76 plus.n75 37.246
R77 plus.n33 plus.n2 37.246
R78 plus.n15 plus.n14 37.246
R79 plus.n84 plus.n83 33.1766
R80 plus.n58 plus.n49 32.8641
R81 plus.n74 plus.n45 32.8641
R82 plus.n32 plus.n31 32.8641
R83 plus.n19 plus.n8 32.8641
R84 plus.n63 plus.n62 28.4823
R85 plus.n70 plus.n69 28.4823
R86 plus.n27 plus.n4 28.4823
R87 plus.n21 plus.n20 28.4823
R88 plus.n64 plus.n47 24.1005
R89 plus.n68 plus.n47 24.1005
R90 plus.n26 plus.n25 24.1005
R91 plus.n25 plus.n6 24.1005
R92 plus.n85 plus.t3 19.8005
R93 plus.n85 plus.t1 19.8005
R94 plus.n87 plus.t4 19.8005
R95 plus.n87 plus.t0 19.8005
R96 plus.n64 plus.n63 19.7187
R97 plus.n69 plus.n68 19.7187
R98 plus.n27 plus.n26 19.7187
R99 plus.n21 plus.n6 19.7187
R100 plus.n62 plus.n49 15.3369
R101 plus.n70 plus.n45 15.3369
R102 plus.n31 plus.n4 15.3369
R103 plus.n20 plus.n19 15.3369
R104 plus plus.n89 15.1953
R105 plus.n53 plus.n52 14.1472
R106 plus.n11 plus.n10 14.1472
R107 plus.n84 plus.n41 11.8774
R108 plus.n58 plus.n57 10.955
R109 plus.n75 plus.n74 10.955
R110 plus.n33 plus.n32 10.955
R111 plus.n15 plus.n8 10.955
R112 plus.n56 plus.n51 6.57323
R113 plus.n76 plus.n43 6.57323
R114 plus.n37 plus.n2 6.57323
R115 plus.n14 plus.n13 6.57323
R116 plus.n89 plus.n88 5.40567
R117 plus.n81 plus.n80 2.19141
R118 plus.n39 plus.n38 2.19141
R119 plus.n89 plus.n84 1.188
R120 plus.n88 plus.n86 0.716017
R121 plus.n55 plus.n54 0.189894
R122 plus.n55 plus.n50 0.189894
R123 plus.n59 plus.n50 0.189894
R124 plus.n60 plus.n59 0.189894
R125 plus.n61 plus.n60 0.189894
R126 plus.n61 plus.n48 0.189894
R127 plus.n65 plus.n48 0.189894
R128 plus.n66 plus.n65 0.189894
R129 plus.n67 plus.n66 0.189894
R130 plus.n67 plus.n46 0.189894
R131 plus.n71 plus.n46 0.189894
R132 plus.n72 plus.n71 0.189894
R133 plus.n73 plus.n72 0.189894
R134 plus.n73 plus.n44 0.189894
R135 plus.n77 plus.n44 0.189894
R136 plus.n78 plus.n77 0.189894
R137 plus.n79 plus.n78 0.189894
R138 plus.n79 plus.n42 0.189894
R139 plus.n83 plus.n42 0.189894
R140 plus.n41 plus.n0 0.189894
R141 plus.n1 plus.n0 0.189894
R142 plus.n36 plus.n1 0.189894
R143 plus.n36 plus.n35 0.189894
R144 plus.n35 plus.n34 0.189894
R145 plus.n34 plus.n3 0.189894
R146 plus.n30 plus.n3 0.189894
R147 plus.n30 plus.n29 0.189894
R148 plus.n29 plus.n28 0.189894
R149 plus.n28 plus.n5 0.189894
R150 plus.n24 plus.n5 0.189894
R151 plus.n24 plus.n23 0.189894
R152 plus.n23 plus.n22 0.189894
R153 plus.n22 plus.n7 0.189894
R154 plus.n18 plus.n7 0.189894
R155 plus.n18 plus.n17 0.189894
R156 plus.n17 plus.n16 0.189894
R157 plus.n16 plus.n9 0.189894
R158 plus.n12 plus.n9 0.189894
R159 a_n3827_n3924.n8 a_n3827_n3924.t15 214.994
R160 a_n3827_n3924.n5 a_n3827_n3924.t57 214.786
R161 a_n3827_n3924.n5 a_n3827_n3924.t20 214.321
R162 a_n3827_n3924.n5 a_n3827_n3924.t11 214.321
R163 a_n3827_n3924.n5 a_n3827_n3924.t1 214.321
R164 a_n3827_n3924.n6 a_n3827_n3924.t16 214.321
R165 a_n3827_n3924.n6 a_n3827_n3924.t53 214.321
R166 a_n3827_n3924.n7 a_n3827_n3924.t2 214.321
R167 a_n3827_n3924.n8 a_n3827_n3924.t3 214.321
R168 a_n3827_n3924.n8 a_n3827_n3924.t21 214.321
R169 a_n3827_n3924.n1 a_n3827_n3924.t23 55.8337
R170 a_n3827_n3924.n1 a_n3827_n3924.t46 55.8337
R171 a_n3827_n3924.n10 a_n3827_n3924.t7 55.8337
R172 a_n3827_n3924.n0 a_n3827_n3924.t43 55.8335
R173 a_n3827_n3924.n9 a_n3827_n3924.t55 55.8335
R174 a_n3827_n3924.n4 a_n3827_n3924.t10 55.8335
R175 a_n3827_n3924.n4 a_n3827_n3924.t36 55.8335
R176 a_n3827_n3924.n3 a_n3827_n3924.t24 55.8335
R177 a_n3827_n3924.n0 a_n3827_n3924.n25 53.0052
R178 a_n3827_n3924.n0 a_n3827_n3924.n26 53.0052
R179 a_n3827_n3924.n0 a_n3827_n3924.n27 53.0052
R180 a_n3827_n3924.n1 a_n3827_n3924.n28 53.0052
R181 a_n3827_n3924.n1 a_n3827_n3924.n29 53.0052
R182 a_n3827_n3924.n1 a_n3827_n3924.n30 53.0052
R183 a_n3827_n3924.n1 a_n3827_n3924.n31 53.0052
R184 a_n3827_n3924.n11 a_n3827_n3924.n32 53.0052
R185 a_n3827_n3924.n10 a_n3827_n3924.n12 53.0052
R186 a_n3827_n3924.n9 a_n3827_n3924.n23 53.0051
R187 a_n3827_n3924.n2 a_n3827_n3924.n22 53.0051
R188 a_n3827_n3924.n2 a_n3827_n3924.n21 53.0051
R189 a_n3827_n3924.n2 a_n3827_n3924.n20 53.0051
R190 a_n3827_n3924.n2 a_n3827_n3924.n19 53.0051
R191 a_n3827_n3924.n4 a_n3827_n3924.n18 53.0051
R192 a_n3827_n3924.n4 a_n3827_n3924.n17 53.0051
R193 a_n3827_n3924.n4 a_n3827_n3924.n16 53.0051
R194 a_n3827_n3924.n3 a_n3827_n3924.n15 53.0051
R195 a_n3827_n3924.n3 a_n3827_n3924.n14 53.0051
R196 a_n3827_n3924.n33 a_n3827_n3924.n11 53.0051
R197 a_n3827_n3924.n13 a_n3827_n3924.n10 12.1986
R198 a_n3827_n3924.n0 a_n3827_n3924.n24 12.1986
R199 a_n3827_n3924.n3 a_n3827_n3924.n13 5.11903
R200 a_n3827_n3924.n24 a_n3827_n3924.n9 5.11903
R201 a_n3827_n3924.n25 a_n3827_n3924.t30 2.82907
R202 a_n3827_n3924.n25 a_n3827_n3924.t41 2.82907
R203 a_n3827_n3924.n26 a_n3827_n3924.t39 2.82907
R204 a_n3827_n3924.n26 a_n3827_n3924.t44 2.82907
R205 a_n3827_n3924.n27 a_n3827_n3924.t42 2.82907
R206 a_n3827_n3924.n27 a_n3827_n3924.t26 2.82907
R207 a_n3827_n3924.n28 a_n3827_n3924.t33 2.82907
R208 a_n3827_n3924.n28 a_n3827_n3924.t29 2.82907
R209 a_n3827_n3924.n29 a_n3827_n3924.t31 2.82907
R210 a_n3827_n3924.n29 a_n3827_n3924.t32 2.82907
R211 a_n3827_n3924.n30 a_n3827_n3924.t56 2.82907
R212 a_n3827_n3924.n30 a_n3827_n3924.t19 2.82907
R213 a_n3827_n3924.n31 a_n3827_n3924.t9 2.82907
R214 a_n3827_n3924.n31 a_n3827_n3924.t6 2.82907
R215 a_n3827_n3924.n32 a_n3827_n3924.t18 2.82907
R216 a_n3827_n3924.n32 a_n3827_n3924.t54 2.82907
R217 a_n3827_n3924.n12 a_n3827_n3924.t14 2.82907
R218 a_n3827_n3924.n12 a_n3827_n3924.t5 2.82907
R219 a_n3827_n3924.n23 a_n3827_n3924.t8 2.82907
R220 a_n3827_n3924.n23 a_n3827_n3924.t51 2.82907
R221 a_n3827_n3924.n22 a_n3827_n3924.t47 2.82907
R222 a_n3827_n3924.n22 a_n3827_n3924.t50 2.82907
R223 a_n3827_n3924.n21 a_n3827_n3924.t48 2.82907
R224 a_n3827_n3924.n21 a_n3827_n3924.t17 2.82907
R225 a_n3827_n3924.n20 a_n3827_n3924.t52 2.82907
R226 a_n3827_n3924.n20 a_n3827_n3924.t13 2.82907
R227 a_n3827_n3924.n19 a_n3827_n3924.t4 2.82907
R228 a_n3827_n3924.n19 a_n3827_n3924.t49 2.82907
R229 a_n3827_n3924.n18 a_n3827_n3924.t45 2.82907
R230 a_n3827_n3924.n18 a_n3827_n3924.t35 2.82907
R231 a_n3827_n3924.n17 a_n3827_n3924.t25 2.82907
R232 a_n3827_n3924.n17 a_n3827_n3924.t37 2.82907
R233 a_n3827_n3924.n16 a_n3827_n3924.t28 2.82907
R234 a_n3827_n3924.n16 a_n3827_n3924.t27 2.82907
R235 a_n3827_n3924.n15 a_n3827_n3924.t38 2.82907
R236 a_n3827_n3924.n15 a_n3827_n3924.t40 2.82907
R237 a_n3827_n3924.n14 a_n3827_n3924.t22 2.82907
R238 a_n3827_n3924.n14 a_n3827_n3924.t34 2.82907
R239 a_n3827_n3924.t0 a_n3827_n3924.n33 2.82907
R240 a_n3827_n3924.n33 a_n3827_n3924.t12 2.82907
R241 a_n3827_n3924.n1 a_n3827_n3924.n0 2.66429
R242 a_n3827_n3924.n6 a_n3827_n3924.n5 2.22216
R243 a_n3827_n3924.n2 a_n3827_n3924.n4 2.01128
R244 a_n3827_n3924.n24 a_n3827_n3924.n5 1.95694
R245 a_n3827_n3924.n13 a_n3827_n3924.n8 1.95694
R246 a_n3827_n3924.n4 a_n3827_n3924.n3 1.77636
R247 a_n3827_n3924.n9 a_n3827_n3924.n2 1.77636
R248 a_n3827_n3924.n11 a_n3827_n3924.n1 1.56731
R249 a_n3827_n3924.n7 a_n3827_n3924.n6 1.34352
R250 a_n3827_n3924.n8 a_n3827_n3924.n7 1.34352
R251 a_n3827_n3924.n11 a_n3827_n3924.n10 1.3324
R252 a_n8300_8799.n182 a_n8300_8799.t131 485.149
R253 a_n8300_8799.n230 a_n8300_8799.t46 485.149
R254 a_n8300_8799.n279 a_n8300_8799.t110 485.149
R255 a_n8300_8799.n34 a_n8300_8799.t96 485.149
R256 a_n8300_8799.n82 a_n8300_8799.t109 485.149
R257 a_n8300_8799.n131 a_n8300_8799.t111 485.149
R258 a_n8300_8799.n214 a_n8300_8799.t94 464.166
R259 a_n8300_8799.n213 a_n8300_8799.t47 464.166
R260 a_n8300_8799.n169 a_n8300_8799.t98 464.166
R261 a_n8300_8799.n207 a_n8300_8799.t97 464.166
R262 a_n8300_8799.n206 a_n8300_8799.t49 464.166
R263 a_n8300_8799.n172 a_n8300_8799.t48 464.166
R264 a_n8300_8799.n200 a_n8300_8799.t116 464.166
R265 a_n8300_8799.n199 a_n8300_8799.t61 464.166
R266 a_n8300_8799.n175 a_n8300_8799.t51 464.166
R267 a_n8300_8799.n194 a_n8300_8799.t120 464.166
R268 a_n8300_8799.n192 a_n8300_8799.t82 464.166
R269 a_n8300_8799.n178 a_n8300_8799.t62 464.166
R270 a_n8300_8799.n187 a_n8300_8799.t137 464.166
R271 a_n8300_8799.n185 a_n8300_8799.t95 464.166
R272 a_n8300_8799.n181 a_n8300_8799.t64 464.166
R273 a_n8300_8799.n262 a_n8300_8799.t107 464.166
R274 a_n8300_8799.n261 a_n8300_8799.t55 464.166
R275 a_n8300_8799.n217 a_n8300_8799.t114 464.166
R276 a_n8300_8799.n255 a_n8300_8799.t113 464.166
R277 a_n8300_8799.n254 a_n8300_8799.t57 464.166
R278 a_n8300_8799.n220 a_n8300_8799.t56 464.166
R279 a_n8300_8799.n248 a_n8300_8799.t130 464.166
R280 a_n8300_8799.n247 a_n8300_8799.t69 464.166
R281 a_n8300_8799.n223 a_n8300_8799.t60 464.166
R282 a_n8300_8799.n242 a_n8300_8799.t132 464.166
R283 a_n8300_8799.n240 a_n8300_8799.t92 464.166
R284 a_n8300_8799.n226 a_n8300_8799.t72 464.166
R285 a_n8300_8799.n235 a_n8300_8799.t50 464.166
R286 a_n8300_8799.n233 a_n8300_8799.t108 464.166
R287 a_n8300_8799.n229 a_n8300_8799.t73 464.166
R288 a_n8300_8799.n311 a_n8300_8799.t65 464.166
R289 a_n8300_8799.n310 a_n8300_8799.t135 464.166
R290 a_n8300_8799.n266 a_n8300_8799.t106 464.166
R291 a_n8300_8799.n304 a_n8300_8799.t129 464.166
R292 a_n8300_8799.n303 a_n8300_8799.t91 464.166
R293 a_n8300_8799.n269 a_n8300_8799.t112 464.166
R294 a_n8300_8799.n297 a_n8300_8799.t59 464.166
R295 a_n8300_8799.n296 a_n8300_8799.t126 464.166
R296 a_n8300_8799.n272 a_n8300_8799.t76 464.166
R297 a_n8300_8799.n291 a_n8300_8799.t121 464.166
R298 a_n8300_8799.n289 a_n8300_8799.t63 464.166
R299 a_n8300_8799.n275 a_n8300_8799.t101 464.166
R300 a_n8300_8799.n284 a_n8300_8799.t54 464.166
R301 a_n8300_8799.n282 a_n8300_8799.t88 464.166
R302 a_n8300_8799.n278 a_n8300_8799.t71 464.166
R303 a_n8300_8799.n33 a_n8300_8799.t128 464.166
R304 a_n8300_8799.n37 a_n8300_8799.t66 464.166
R305 a_n8300_8799.n31 a_n8300_8799.t93 464.166
R306 a_n8300_8799.n42 a_n8300_8799.t123 464.166
R307 a_n8300_8799.n44 a_n8300_8799.t124 464.166
R308 a_n8300_8799.n48 a_n8300_8799.t81 464.166
R309 a_n8300_8799.n49 a_n8300_8799.t105 464.166
R310 a_n8300_8799.n27 a_n8300_8799.t122 464.166
R311 a_n8300_8799.n54 a_n8300_8799.t79 464.166
R312 a_n8300_8799.n56 a_n8300_8799.t80 464.166
R313 a_n8300_8799.n60 a_n8300_8799.t102 464.166
R314 a_n8300_8799.n61 a_n8300_8799.t67 464.166
R315 a_n8300_8799.n23 a_n8300_8799.t68 464.166
R316 a_n8300_8799.n67 a_n8300_8799.t99 464.166
R317 a_n8300_8799.n68 a_n8300_8799.t44 464.166
R318 a_n8300_8799.n81 a_n8300_8799.t139 464.166
R319 a_n8300_8799.n85 a_n8300_8799.t74 464.166
R320 a_n8300_8799.n79 a_n8300_8799.t103 464.166
R321 a_n8300_8799.n90 a_n8300_8799.t136 464.166
R322 a_n8300_8799.n92 a_n8300_8799.t138 464.166
R323 a_n8300_8799.n96 a_n8300_8799.t89 464.166
R324 a_n8300_8799.n97 a_n8300_8799.t119 464.166
R325 a_n8300_8799.n75 a_n8300_8799.t134 464.166
R326 a_n8300_8799.n102 a_n8300_8799.t85 464.166
R327 a_n8300_8799.n104 a_n8300_8799.t86 464.166
R328 a_n8300_8799.n108 a_n8300_8799.t117 464.166
R329 a_n8300_8799.n109 a_n8300_8799.t77 464.166
R330 a_n8300_8799.n71 a_n8300_8799.t78 464.166
R331 a_n8300_8799.n115 a_n8300_8799.t115 464.166
R332 a_n8300_8799.n116 a_n8300_8799.t52 464.166
R333 a_n8300_8799.n130 a_n8300_8799.t70 464.166
R334 a_n8300_8799.n134 a_n8300_8799.t87 464.166
R335 a_n8300_8799.n128 a_n8300_8799.t53 464.166
R336 a_n8300_8799.n139 a_n8300_8799.t100 464.166
R337 a_n8300_8799.n141 a_n8300_8799.t83 464.166
R338 a_n8300_8799.n145 a_n8300_8799.t118 464.166
R339 a_n8300_8799.n146 a_n8300_8799.t75 464.166
R340 a_n8300_8799.n124 a_n8300_8799.t125 464.166
R341 a_n8300_8799.n151 a_n8300_8799.t58 464.166
R342 a_n8300_8799.n153 a_n8300_8799.t45 464.166
R343 a_n8300_8799.n157 a_n8300_8799.t90 464.166
R344 a_n8300_8799.n158 a_n8300_8799.t127 464.166
R345 a_n8300_8799.n120 a_n8300_8799.t104 464.166
R346 a_n8300_8799.n164 a_n8300_8799.t133 464.166
R347 a_n8300_8799.n165 a_n8300_8799.t84 464.166
R348 a_n8300_8799.n184 a_n8300_8799.n183 161.3
R349 a_n8300_8799.n185 a_n8300_8799.n180 161.3
R350 a_n8300_8799.n186 a_n8300_8799.n179 161.3
R351 a_n8300_8799.n188 a_n8300_8799.n187 161.3
R352 a_n8300_8799.n189 a_n8300_8799.n178 161.3
R353 a_n8300_8799.n191 a_n8300_8799.n190 161.3
R354 a_n8300_8799.n192 a_n8300_8799.n177 161.3
R355 a_n8300_8799.n193 a_n8300_8799.n176 161.3
R356 a_n8300_8799.n195 a_n8300_8799.n194 161.3
R357 a_n8300_8799.n196 a_n8300_8799.n175 161.3
R358 a_n8300_8799.n198 a_n8300_8799.n197 161.3
R359 a_n8300_8799.n199 a_n8300_8799.n174 161.3
R360 a_n8300_8799.n200 a_n8300_8799.n173 161.3
R361 a_n8300_8799.n202 a_n8300_8799.n201 161.3
R362 a_n8300_8799.n203 a_n8300_8799.n172 161.3
R363 a_n8300_8799.n205 a_n8300_8799.n204 161.3
R364 a_n8300_8799.n206 a_n8300_8799.n171 161.3
R365 a_n8300_8799.n207 a_n8300_8799.n170 161.3
R366 a_n8300_8799.n209 a_n8300_8799.n208 161.3
R367 a_n8300_8799.n210 a_n8300_8799.n169 161.3
R368 a_n8300_8799.n212 a_n8300_8799.n211 161.3
R369 a_n8300_8799.n213 a_n8300_8799.n168 161.3
R370 a_n8300_8799.n215 a_n8300_8799.n214 161.3
R371 a_n8300_8799.n232 a_n8300_8799.n231 161.3
R372 a_n8300_8799.n233 a_n8300_8799.n228 161.3
R373 a_n8300_8799.n234 a_n8300_8799.n227 161.3
R374 a_n8300_8799.n236 a_n8300_8799.n235 161.3
R375 a_n8300_8799.n237 a_n8300_8799.n226 161.3
R376 a_n8300_8799.n239 a_n8300_8799.n238 161.3
R377 a_n8300_8799.n240 a_n8300_8799.n225 161.3
R378 a_n8300_8799.n241 a_n8300_8799.n224 161.3
R379 a_n8300_8799.n243 a_n8300_8799.n242 161.3
R380 a_n8300_8799.n244 a_n8300_8799.n223 161.3
R381 a_n8300_8799.n246 a_n8300_8799.n245 161.3
R382 a_n8300_8799.n247 a_n8300_8799.n222 161.3
R383 a_n8300_8799.n248 a_n8300_8799.n221 161.3
R384 a_n8300_8799.n250 a_n8300_8799.n249 161.3
R385 a_n8300_8799.n251 a_n8300_8799.n220 161.3
R386 a_n8300_8799.n253 a_n8300_8799.n252 161.3
R387 a_n8300_8799.n254 a_n8300_8799.n219 161.3
R388 a_n8300_8799.n255 a_n8300_8799.n218 161.3
R389 a_n8300_8799.n257 a_n8300_8799.n256 161.3
R390 a_n8300_8799.n258 a_n8300_8799.n217 161.3
R391 a_n8300_8799.n260 a_n8300_8799.n259 161.3
R392 a_n8300_8799.n261 a_n8300_8799.n216 161.3
R393 a_n8300_8799.n263 a_n8300_8799.n262 161.3
R394 a_n8300_8799.n281 a_n8300_8799.n280 161.3
R395 a_n8300_8799.n282 a_n8300_8799.n277 161.3
R396 a_n8300_8799.n283 a_n8300_8799.n276 161.3
R397 a_n8300_8799.n285 a_n8300_8799.n284 161.3
R398 a_n8300_8799.n286 a_n8300_8799.n275 161.3
R399 a_n8300_8799.n288 a_n8300_8799.n287 161.3
R400 a_n8300_8799.n289 a_n8300_8799.n274 161.3
R401 a_n8300_8799.n290 a_n8300_8799.n273 161.3
R402 a_n8300_8799.n292 a_n8300_8799.n291 161.3
R403 a_n8300_8799.n293 a_n8300_8799.n272 161.3
R404 a_n8300_8799.n295 a_n8300_8799.n294 161.3
R405 a_n8300_8799.n296 a_n8300_8799.n271 161.3
R406 a_n8300_8799.n297 a_n8300_8799.n270 161.3
R407 a_n8300_8799.n299 a_n8300_8799.n298 161.3
R408 a_n8300_8799.n300 a_n8300_8799.n269 161.3
R409 a_n8300_8799.n302 a_n8300_8799.n301 161.3
R410 a_n8300_8799.n303 a_n8300_8799.n268 161.3
R411 a_n8300_8799.n304 a_n8300_8799.n267 161.3
R412 a_n8300_8799.n306 a_n8300_8799.n305 161.3
R413 a_n8300_8799.n307 a_n8300_8799.n266 161.3
R414 a_n8300_8799.n309 a_n8300_8799.n308 161.3
R415 a_n8300_8799.n310 a_n8300_8799.n265 161.3
R416 a_n8300_8799.n312 a_n8300_8799.n311 161.3
R417 a_n8300_8799.n69 a_n8300_8799.n68 161.3
R418 a_n8300_8799.n67 a_n8300_8799.n22 161.3
R419 a_n8300_8799.n66 a_n8300_8799.n65 161.3
R420 a_n8300_8799.n64 a_n8300_8799.n23 161.3
R421 a_n8300_8799.n63 a_n8300_8799.n62 161.3
R422 a_n8300_8799.n61 a_n8300_8799.n24 161.3
R423 a_n8300_8799.n60 a_n8300_8799.n59 161.3
R424 a_n8300_8799.n58 a_n8300_8799.n25 161.3
R425 a_n8300_8799.n57 a_n8300_8799.n56 161.3
R426 a_n8300_8799.n55 a_n8300_8799.n26 161.3
R427 a_n8300_8799.n54 a_n8300_8799.n53 161.3
R428 a_n8300_8799.n52 a_n8300_8799.n27 161.3
R429 a_n8300_8799.n51 a_n8300_8799.n50 161.3
R430 a_n8300_8799.n49 a_n8300_8799.n28 161.3
R431 a_n8300_8799.n48 a_n8300_8799.n47 161.3
R432 a_n8300_8799.n46 a_n8300_8799.n29 161.3
R433 a_n8300_8799.n45 a_n8300_8799.n44 161.3
R434 a_n8300_8799.n43 a_n8300_8799.n30 161.3
R435 a_n8300_8799.n42 a_n8300_8799.n41 161.3
R436 a_n8300_8799.n40 a_n8300_8799.n31 161.3
R437 a_n8300_8799.n39 a_n8300_8799.n38 161.3
R438 a_n8300_8799.n37 a_n8300_8799.n32 161.3
R439 a_n8300_8799.n36 a_n8300_8799.n35 161.3
R440 a_n8300_8799.n117 a_n8300_8799.n116 161.3
R441 a_n8300_8799.n115 a_n8300_8799.n70 161.3
R442 a_n8300_8799.n114 a_n8300_8799.n113 161.3
R443 a_n8300_8799.n112 a_n8300_8799.n71 161.3
R444 a_n8300_8799.n111 a_n8300_8799.n110 161.3
R445 a_n8300_8799.n109 a_n8300_8799.n72 161.3
R446 a_n8300_8799.n108 a_n8300_8799.n107 161.3
R447 a_n8300_8799.n106 a_n8300_8799.n73 161.3
R448 a_n8300_8799.n105 a_n8300_8799.n104 161.3
R449 a_n8300_8799.n103 a_n8300_8799.n74 161.3
R450 a_n8300_8799.n102 a_n8300_8799.n101 161.3
R451 a_n8300_8799.n100 a_n8300_8799.n75 161.3
R452 a_n8300_8799.n99 a_n8300_8799.n98 161.3
R453 a_n8300_8799.n97 a_n8300_8799.n76 161.3
R454 a_n8300_8799.n96 a_n8300_8799.n95 161.3
R455 a_n8300_8799.n94 a_n8300_8799.n77 161.3
R456 a_n8300_8799.n93 a_n8300_8799.n92 161.3
R457 a_n8300_8799.n91 a_n8300_8799.n78 161.3
R458 a_n8300_8799.n90 a_n8300_8799.n89 161.3
R459 a_n8300_8799.n88 a_n8300_8799.n79 161.3
R460 a_n8300_8799.n87 a_n8300_8799.n86 161.3
R461 a_n8300_8799.n85 a_n8300_8799.n80 161.3
R462 a_n8300_8799.n84 a_n8300_8799.n83 161.3
R463 a_n8300_8799.n166 a_n8300_8799.n165 161.3
R464 a_n8300_8799.n164 a_n8300_8799.n119 161.3
R465 a_n8300_8799.n163 a_n8300_8799.n162 161.3
R466 a_n8300_8799.n161 a_n8300_8799.n120 161.3
R467 a_n8300_8799.n160 a_n8300_8799.n159 161.3
R468 a_n8300_8799.n158 a_n8300_8799.n121 161.3
R469 a_n8300_8799.n157 a_n8300_8799.n156 161.3
R470 a_n8300_8799.n155 a_n8300_8799.n122 161.3
R471 a_n8300_8799.n154 a_n8300_8799.n153 161.3
R472 a_n8300_8799.n152 a_n8300_8799.n123 161.3
R473 a_n8300_8799.n151 a_n8300_8799.n150 161.3
R474 a_n8300_8799.n149 a_n8300_8799.n124 161.3
R475 a_n8300_8799.n148 a_n8300_8799.n147 161.3
R476 a_n8300_8799.n146 a_n8300_8799.n125 161.3
R477 a_n8300_8799.n145 a_n8300_8799.n144 161.3
R478 a_n8300_8799.n143 a_n8300_8799.n126 161.3
R479 a_n8300_8799.n142 a_n8300_8799.n141 161.3
R480 a_n8300_8799.n140 a_n8300_8799.n127 161.3
R481 a_n8300_8799.n139 a_n8300_8799.n138 161.3
R482 a_n8300_8799.n137 a_n8300_8799.n128 161.3
R483 a_n8300_8799.n136 a_n8300_8799.n135 161.3
R484 a_n8300_8799.n134 a_n8300_8799.n129 161.3
R485 a_n8300_8799.n133 a_n8300_8799.n132 161.3
R486 a_n8300_8799.n14 a_n8300_8799.n12 98.9633
R487 a_n8300_8799.n5 a_n8300_8799.n3 98.9631
R488 a_n8300_8799.n20 a_n8300_8799.n19 98.6055
R489 a_n8300_8799.n18 a_n8300_8799.n17 98.6055
R490 a_n8300_8799.n16 a_n8300_8799.n15 98.6055
R491 a_n8300_8799.n14 a_n8300_8799.n13 98.6055
R492 a_n8300_8799.n5 a_n8300_8799.n4 98.6055
R493 a_n8300_8799.n7 a_n8300_8799.n6 98.6055
R494 a_n8300_8799.n9 a_n8300_8799.n8 98.6055
R495 a_n8300_8799.n11 a_n8300_8799.n10 98.6055
R496 a_n8300_8799.n318 a_n8300_8799.n316 81.3764
R497 a_n8300_8799.n330 a_n8300_8799.n328 81.3764
R498 a_n8300_8799.n2 a_n8300_8799.n0 81.3764
R499 a_n8300_8799.n335 a_n8300_8799.n334 80.9326
R500 a_n8300_8799.n327 a_n8300_8799.n326 80.9324
R501 a_n8300_8799.n325 a_n8300_8799.n324 80.9324
R502 a_n8300_8799.n323 a_n8300_8799.n322 80.9324
R503 a_n8300_8799.n320 a_n8300_8799.n319 80.9324
R504 a_n8300_8799.n318 a_n8300_8799.n317 80.9324
R505 a_n8300_8799.n330 a_n8300_8799.n329 80.9324
R506 a_n8300_8799.n332 a_n8300_8799.n331 80.9324
R507 a_n8300_8799.n2 a_n8300_8799.n1 80.9324
R508 a_n8300_8799.n183 a_n8300_8799.n182 70.4033
R509 a_n8300_8799.n231 a_n8300_8799.n230 70.4033
R510 a_n8300_8799.n280 a_n8300_8799.n279 70.4033
R511 a_n8300_8799.n35 a_n8300_8799.n34 70.4033
R512 a_n8300_8799.n83 a_n8300_8799.n82 70.4033
R513 a_n8300_8799.n132 a_n8300_8799.n131 70.4033
R514 a_n8300_8799.n214 a_n8300_8799.n213 48.2005
R515 a_n8300_8799.n207 a_n8300_8799.n206 48.2005
R516 a_n8300_8799.n200 a_n8300_8799.n199 48.2005
R517 a_n8300_8799.n194 a_n8300_8799.n175 48.2005
R518 a_n8300_8799.n187 a_n8300_8799.n178 48.2005
R519 a_n8300_8799.n262 a_n8300_8799.n261 48.2005
R520 a_n8300_8799.n255 a_n8300_8799.n254 48.2005
R521 a_n8300_8799.n248 a_n8300_8799.n247 48.2005
R522 a_n8300_8799.n242 a_n8300_8799.n223 48.2005
R523 a_n8300_8799.n235 a_n8300_8799.n226 48.2005
R524 a_n8300_8799.n311 a_n8300_8799.n310 48.2005
R525 a_n8300_8799.n304 a_n8300_8799.n303 48.2005
R526 a_n8300_8799.n297 a_n8300_8799.n296 48.2005
R527 a_n8300_8799.n291 a_n8300_8799.n272 48.2005
R528 a_n8300_8799.n284 a_n8300_8799.n275 48.2005
R529 a_n8300_8799.n42 a_n8300_8799.n31 48.2005
R530 a_n8300_8799.n49 a_n8300_8799.n48 48.2005
R531 a_n8300_8799.n54 a_n8300_8799.n27 48.2005
R532 a_n8300_8799.n61 a_n8300_8799.n60 48.2005
R533 a_n8300_8799.n68 a_n8300_8799.n67 48.2005
R534 a_n8300_8799.n90 a_n8300_8799.n79 48.2005
R535 a_n8300_8799.n97 a_n8300_8799.n96 48.2005
R536 a_n8300_8799.n102 a_n8300_8799.n75 48.2005
R537 a_n8300_8799.n109 a_n8300_8799.n108 48.2005
R538 a_n8300_8799.n116 a_n8300_8799.n115 48.2005
R539 a_n8300_8799.n139 a_n8300_8799.n128 48.2005
R540 a_n8300_8799.n146 a_n8300_8799.n145 48.2005
R541 a_n8300_8799.n151 a_n8300_8799.n124 48.2005
R542 a_n8300_8799.n158 a_n8300_8799.n157 48.2005
R543 a_n8300_8799.n165 a_n8300_8799.n164 48.2005
R544 a_n8300_8799.n201 a_n8300_8799.n172 47.4702
R545 a_n8300_8799.n193 a_n8300_8799.n192 47.4702
R546 a_n8300_8799.n249 a_n8300_8799.n220 47.4702
R547 a_n8300_8799.n241 a_n8300_8799.n240 47.4702
R548 a_n8300_8799.n298 a_n8300_8799.n269 47.4702
R549 a_n8300_8799.n290 a_n8300_8799.n289 47.4702
R550 a_n8300_8799.n44 a_n8300_8799.n29 47.4702
R551 a_n8300_8799.n56 a_n8300_8799.n55 47.4702
R552 a_n8300_8799.n92 a_n8300_8799.n77 47.4702
R553 a_n8300_8799.n104 a_n8300_8799.n103 47.4702
R554 a_n8300_8799.n141 a_n8300_8799.n126 47.4702
R555 a_n8300_8799.n153 a_n8300_8799.n152 47.4702
R556 a_n8300_8799.n208 a_n8300_8799.n169 46.0096
R557 a_n8300_8799.n186 a_n8300_8799.n185 46.0096
R558 a_n8300_8799.n256 a_n8300_8799.n217 46.0096
R559 a_n8300_8799.n234 a_n8300_8799.n233 46.0096
R560 a_n8300_8799.n305 a_n8300_8799.n266 46.0096
R561 a_n8300_8799.n283 a_n8300_8799.n282 46.0096
R562 a_n8300_8799.n38 a_n8300_8799.n37 46.0096
R563 a_n8300_8799.n62 a_n8300_8799.n23 46.0096
R564 a_n8300_8799.n86 a_n8300_8799.n85 46.0096
R565 a_n8300_8799.n110 a_n8300_8799.n71 46.0096
R566 a_n8300_8799.n135 a_n8300_8799.n134 46.0096
R567 a_n8300_8799.n159 a_n8300_8799.n120 46.0096
R568 a_n8300_8799.n333 a_n8300_8799.n327 33.4185
R569 a_n8300_8799.n21 a_n8300_8799.n11 33.0821
R570 a_n8300_8799.n212 a_n8300_8799.n169 27.0217
R571 a_n8300_8799.n185 a_n8300_8799.n184 27.0217
R572 a_n8300_8799.n260 a_n8300_8799.n217 27.0217
R573 a_n8300_8799.n233 a_n8300_8799.n232 27.0217
R574 a_n8300_8799.n309 a_n8300_8799.n266 27.0217
R575 a_n8300_8799.n282 a_n8300_8799.n281 27.0217
R576 a_n8300_8799.n37 a_n8300_8799.n36 27.0217
R577 a_n8300_8799.n66 a_n8300_8799.n23 27.0217
R578 a_n8300_8799.n85 a_n8300_8799.n84 27.0217
R579 a_n8300_8799.n114 a_n8300_8799.n71 27.0217
R580 a_n8300_8799.n134 a_n8300_8799.n133 27.0217
R581 a_n8300_8799.n163 a_n8300_8799.n120 27.0217
R582 a_n8300_8799.n205 a_n8300_8799.n172 25.5611
R583 a_n8300_8799.n192 a_n8300_8799.n191 25.5611
R584 a_n8300_8799.n253 a_n8300_8799.n220 25.5611
R585 a_n8300_8799.n240 a_n8300_8799.n239 25.5611
R586 a_n8300_8799.n302 a_n8300_8799.n269 25.5611
R587 a_n8300_8799.n289 a_n8300_8799.n288 25.5611
R588 a_n8300_8799.n44 a_n8300_8799.n43 25.5611
R589 a_n8300_8799.n56 a_n8300_8799.n25 25.5611
R590 a_n8300_8799.n92 a_n8300_8799.n91 25.5611
R591 a_n8300_8799.n104 a_n8300_8799.n73 25.5611
R592 a_n8300_8799.n141 a_n8300_8799.n140 25.5611
R593 a_n8300_8799.n153 a_n8300_8799.n122 25.5611
R594 a_n8300_8799.n199 a_n8300_8799.n198 24.1005
R595 a_n8300_8799.n198 a_n8300_8799.n175 24.1005
R596 a_n8300_8799.n247 a_n8300_8799.n246 24.1005
R597 a_n8300_8799.n246 a_n8300_8799.n223 24.1005
R598 a_n8300_8799.n296 a_n8300_8799.n295 24.1005
R599 a_n8300_8799.n295 a_n8300_8799.n272 24.1005
R600 a_n8300_8799.n50 a_n8300_8799.n49 24.1005
R601 a_n8300_8799.n50 a_n8300_8799.n27 24.1005
R602 a_n8300_8799.n98 a_n8300_8799.n97 24.1005
R603 a_n8300_8799.n98 a_n8300_8799.n75 24.1005
R604 a_n8300_8799.n147 a_n8300_8799.n146 24.1005
R605 a_n8300_8799.n147 a_n8300_8799.n124 24.1005
R606 a_n8300_8799.n206 a_n8300_8799.n205 22.6399
R607 a_n8300_8799.n191 a_n8300_8799.n178 22.6399
R608 a_n8300_8799.n254 a_n8300_8799.n253 22.6399
R609 a_n8300_8799.n239 a_n8300_8799.n226 22.6399
R610 a_n8300_8799.n303 a_n8300_8799.n302 22.6399
R611 a_n8300_8799.n288 a_n8300_8799.n275 22.6399
R612 a_n8300_8799.n43 a_n8300_8799.n42 22.6399
R613 a_n8300_8799.n60 a_n8300_8799.n25 22.6399
R614 a_n8300_8799.n91 a_n8300_8799.n90 22.6399
R615 a_n8300_8799.n108 a_n8300_8799.n73 22.6399
R616 a_n8300_8799.n140 a_n8300_8799.n139 22.6399
R617 a_n8300_8799.n157 a_n8300_8799.n122 22.6399
R618 a_n8300_8799.n213 a_n8300_8799.n212 21.1793
R619 a_n8300_8799.n184 a_n8300_8799.n181 21.1793
R620 a_n8300_8799.n261 a_n8300_8799.n260 21.1793
R621 a_n8300_8799.n232 a_n8300_8799.n229 21.1793
R622 a_n8300_8799.n310 a_n8300_8799.n309 21.1793
R623 a_n8300_8799.n281 a_n8300_8799.n278 21.1793
R624 a_n8300_8799.n36 a_n8300_8799.n33 21.1793
R625 a_n8300_8799.n67 a_n8300_8799.n66 21.1793
R626 a_n8300_8799.n84 a_n8300_8799.n81 21.1793
R627 a_n8300_8799.n115 a_n8300_8799.n114 21.1793
R628 a_n8300_8799.n133 a_n8300_8799.n130 21.1793
R629 a_n8300_8799.n164 a_n8300_8799.n163 21.1793
R630 a_n8300_8799.n182 a_n8300_8799.n181 20.9576
R631 a_n8300_8799.n230 a_n8300_8799.n229 20.9576
R632 a_n8300_8799.n279 a_n8300_8799.n278 20.9576
R633 a_n8300_8799.n34 a_n8300_8799.n33 20.9576
R634 a_n8300_8799.n82 a_n8300_8799.n81 20.9576
R635 a_n8300_8799.n131 a_n8300_8799.n130 20.9576
R636 a_n8300_8799.n21 a_n8300_8799.n20 19.6606
R637 a_n8300_8799.n321 a_n8300_8799.n315 12.3339
R638 a_n8300_8799.n315 a_n8300_8799.n21 11.4887
R639 a_n8300_8799.n264 a_n8300_8799.n215 9.07815
R640 a_n8300_8799.n118 a_n8300_8799.n69 9.07815
R641 a_n8300_8799.n314 a_n8300_8799.n167 7.11017
R642 a_n8300_8799.n314 a_n8300_8799.n313 6.68874
R643 a_n8300_8799.n264 a_n8300_8799.n263 4.9702
R644 a_n8300_8799.n313 a_n8300_8799.n312 4.9702
R645 a_n8300_8799.n118 a_n8300_8799.n117 4.9702
R646 a_n8300_8799.n167 a_n8300_8799.n166 4.9702
R647 a_n8300_8799.n313 a_n8300_8799.n264 4.10845
R648 a_n8300_8799.n167 a_n8300_8799.n118 4.10845
R649 a_n8300_8799.n19 a_n8300_8799.t5 3.61217
R650 a_n8300_8799.n19 a_n8300_8799.t8 3.61217
R651 a_n8300_8799.n17 a_n8300_8799.t2 3.61217
R652 a_n8300_8799.n17 a_n8300_8799.t17 3.61217
R653 a_n8300_8799.n15 a_n8300_8799.t16 3.61217
R654 a_n8300_8799.n15 a_n8300_8799.t15 3.61217
R655 a_n8300_8799.n13 a_n8300_8799.t4 3.61217
R656 a_n8300_8799.n13 a_n8300_8799.t10 3.61217
R657 a_n8300_8799.n12 a_n8300_8799.t3 3.61217
R658 a_n8300_8799.n12 a_n8300_8799.t12 3.61217
R659 a_n8300_8799.n3 a_n8300_8799.t0 3.61217
R660 a_n8300_8799.n3 a_n8300_8799.t18 3.61217
R661 a_n8300_8799.n4 a_n8300_8799.t1 3.61217
R662 a_n8300_8799.n4 a_n8300_8799.t11 3.61217
R663 a_n8300_8799.n6 a_n8300_8799.t6 3.61217
R664 a_n8300_8799.n6 a_n8300_8799.t7 3.61217
R665 a_n8300_8799.n8 a_n8300_8799.t14 3.61217
R666 a_n8300_8799.n8 a_n8300_8799.t19 3.61217
R667 a_n8300_8799.n10 a_n8300_8799.t9 3.61217
R668 a_n8300_8799.n10 a_n8300_8799.t13 3.61217
R669 a_n8300_8799.n315 a_n8300_8799.n314 3.4105
R670 a_n8300_8799.n328 a_n8300_8799.t35 2.82907
R671 a_n8300_8799.n328 a_n8300_8799.t33 2.82907
R672 a_n8300_8799.n329 a_n8300_8799.t24 2.82907
R673 a_n8300_8799.n329 a_n8300_8799.t30 2.82907
R674 a_n8300_8799.n331 a_n8300_8799.t42 2.82907
R675 a_n8300_8799.n331 a_n8300_8799.t25 2.82907
R676 a_n8300_8799.n1 a_n8300_8799.t32 2.82907
R677 a_n8300_8799.n1 a_n8300_8799.t31 2.82907
R678 a_n8300_8799.n0 a_n8300_8799.t27 2.82907
R679 a_n8300_8799.n0 a_n8300_8799.t26 2.82907
R680 a_n8300_8799.n326 a_n8300_8799.t38 2.82907
R681 a_n8300_8799.n326 a_n8300_8799.t40 2.82907
R682 a_n8300_8799.n324 a_n8300_8799.t36 2.82907
R683 a_n8300_8799.n324 a_n8300_8799.t20 2.82907
R684 a_n8300_8799.n322 a_n8300_8799.t41 2.82907
R685 a_n8300_8799.n322 a_n8300_8799.t34 2.82907
R686 a_n8300_8799.n319 a_n8300_8799.t21 2.82907
R687 a_n8300_8799.n319 a_n8300_8799.t39 2.82907
R688 a_n8300_8799.n317 a_n8300_8799.t22 2.82907
R689 a_n8300_8799.n317 a_n8300_8799.t23 2.82907
R690 a_n8300_8799.n316 a_n8300_8799.t28 2.82907
R691 a_n8300_8799.n316 a_n8300_8799.t29 2.82907
R692 a_n8300_8799.n335 a_n8300_8799.t37 2.82907
R693 a_n8300_8799.t43 a_n8300_8799.n335 2.82907
R694 a_n8300_8799.n208 a_n8300_8799.n207 2.19141
R695 a_n8300_8799.n187 a_n8300_8799.n186 2.19141
R696 a_n8300_8799.n256 a_n8300_8799.n255 2.19141
R697 a_n8300_8799.n235 a_n8300_8799.n234 2.19141
R698 a_n8300_8799.n305 a_n8300_8799.n304 2.19141
R699 a_n8300_8799.n284 a_n8300_8799.n283 2.19141
R700 a_n8300_8799.n38 a_n8300_8799.n31 2.19141
R701 a_n8300_8799.n62 a_n8300_8799.n61 2.19141
R702 a_n8300_8799.n86 a_n8300_8799.n79 2.19141
R703 a_n8300_8799.n110 a_n8300_8799.n109 2.19141
R704 a_n8300_8799.n135 a_n8300_8799.n128 2.19141
R705 a_n8300_8799.n159 a_n8300_8799.n158 2.19141
R706 a_n8300_8799.n201 a_n8300_8799.n200 0.730803
R707 a_n8300_8799.n194 a_n8300_8799.n193 0.730803
R708 a_n8300_8799.n249 a_n8300_8799.n248 0.730803
R709 a_n8300_8799.n242 a_n8300_8799.n241 0.730803
R710 a_n8300_8799.n298 a_n8300_8799.n297 0.730803
R711 a_n8300_8799.n291 a_n8300_8799.n290 0.730803
R712 a_n8300_8799.n48 a_n8300_8799.n29 0.730803
R713 a_n8300_8799.n55 a_n8300_8799.n54 0.730803
R714 a_n8300_8799.n96 a_n8300_8799.n77 0.730803
R715 a_n8300_8799.n103 a_n8300_8799.n102 0.730803
R716 a_n8300_8799.n145 a_n8300_8799.n126 0.730803
R717 a_n8300_8799.n152 a_n8300_8799.n151 0.730803
R718 a_n8300_8799.n320 a_n8300_8799.n318 0.444466
R719 a_n8300_8799.n325 a_n8300_8799.n323 0.444466
R720 a_n8300_8799.n327 a_n8300_8799.n325 0.444466
R721 a_n8300_8799.n334 a_n8300_8799.n2 0.444466
R722 a_n8300_8799.n332 a_n8300_8799.n330 0.444466
R723 a_n8300_8799.n16 a_n8300_8799.n14 0.358259
R724 a_n8300_8799.n18 a_n8300_8799.n16 0.358259
R725 a_n8300_8799.n20 a_n8300_8799.n18 0.358259
R726 a_n8300_8799.n11 a_n8300_8799.n9 0.358259
R727 a_n8300_8799.n9 a_n8300_8799.n7 0.358259
R728 a_n8300_8799.n7 a_n8300_8799.n5 0.358259
R729 a_n8300_8799.n321 a_n8300_8799.n320 0.222483
R730 a_n8300_8799.n323 a_n8300_8799.n321 0.222483
R731 a_n8300_8799.n334 a_n8300_8799.n333 0.222483
R732 a_n8300_8799.n333 a_n8300_8799.n332 0.222483
R733 a_n8300_8799.n215 a_n8300_8799.n168 0.189894
R734 a_n8300_8799.n211 a_n8300_8799.n168 0.189894
R735 a_n8300_8799.n211 a_n8300_8799.n210 0.189894
R736 a_n8300_8799.n210 a_n8300_8799.n209 0.189894
R737 a_n8300_8799.n209 a_n8300_8799.n170 0.189894
R738 a_n8300_8799.n171 a_n8300_8799.n170 0.189894
R739 a_n8300_8799.n204 a_n8300_8799.n171 0.189894
R740 a_n8300_8799.n204 a_n8300_8799.n203 0.189894
R741 a_n8300_8799.n203 a_n8300_8799.n202 0.189894
R742 a_n8300_8799.n202 a_n8300_8799.n173 0.189894
R743 a_n8300_8799.n174 a_n8300_8799.n173 0.189894
R744 a_n8300_8799.n197 a_n8300_8799.n174 0.189894
R745 a_n8300_8799.n197 a_n8300_8799.n196 0.189894
R746 a_n8300_8799.n196 a_n8300_8799.n195 0.189894
R747 a_n8300_8799.n195 a_n8300_8799.n176 0.189894
R748 a_n8300_8799.n177 a_n8300_8799.n176 0.189894
R749 a_n8300_8799.n190 a_n8300_8799.n177 0.189894
R750 a_n8300_8799.n190 a_n8300_8799.n189 0.189894
R751 a_n8300_8799.n189 a_n8300_8799.n188 0.189894
R752 a_n8300_8799.n188 a_n8300_8799.n179 0.189894
R753 a_n8300_8799.n180 a_n8300_8799.n179 0.189894
R754 a_n8300_8799.n183 a_n8300_8799.n180 0.189894
R755 a_n8300_8799.n263 a_n8300_8799.n216 0.189894
R756 a_n8300_8799.n259 a_n8300_8799.n216 0.189894
R757 a_n8300_8799.n259 a_n8300_8799.n258 0.189894
R758 a_n8300_8799.n258 a_n8300_8799.n257 0.189894
R759 a_n8300_8799.n257 a_n8300_8799.n218 0.189894
R760 a_n8300_8799.n219 a_n8300_8799.n218 0.189894
R761 a_n8300_8799.n252 a_n8300_8799.n219 0.189894
R762 a_n8300_8799.n252 a_n8300_8799.n251 0.189894
R763 a_n8300_8799.n251 a_n8300_8799.n250 0.189894
R764 a_n8300_8799.n250 a_n8300_8799.n221 0.189894
R765 a_n8300_8799.n222 a_n8300_8799.n221 0.189894
R766 a_n8300_8799.n245 a_n8300_8799.n222 0.189894
R767 a_n8300_8799.n245 a_n8300_8799.n244 0.189894
R768 a_n8300_8799.n244 a_n8300_8799.n243 0.189894
R769 a_n8300_8799.n243 a_n8300_8799.n224 0.189894
R770 a_n8300_8799.n225 a_n8300_8799.n224 0.189894
R771 a_n8300_8799.n238 a_n8300_8799.n225 0.189894
R772 a_n8300_8799.n238 a_n8300_8799.n237 0.189894
R773 a_n8300_8799.n237 a_n8300_8799.n236 0.189894
R774 a_n8300_8799.n236 a_n8300_8799.n227 0.189894
R775 a_n8300_8799.n228 a_n8300_8799.n227 0.189894
R776 a_n8300_8799.n231 a_n8300_8799.n228 0.189894
R777 a_n8300_8799.n312 a_n8300_8799.n265 0.189894
R778 a_n8300_8799.n308 a_n8300_8799.n265 0.189894
R779 a_n8300_8799.n308 a_n8300_8799.n307 0.189894
R780 a_n8300_8799.n307 a_n8300_8799.n306 0.189894
R781 a_n8300_8799.n306 a_n8300_8799.n267 0.189894
R782 a_n8300_8799.n268 a_n8300_8799.n267 0.189894
R783 a_n8300_8799.n301 a_n8300_8799.n268 0.189894
R784 a_n8300_8799.n301 a_n8300_8799.n300 0.189894
R785 a_n8300_8799.n300 a_n8300_8799.n299 0.189894
R786 a_n8300_8799.n299 a_n8300_8799.n270 0.189894
R787 a_n8300_8799.n271 a_n8300_8799.n270 0.189894
R788 a_n8300_8799.n294 a_n8300_8799.n271 0.189894
R789 a_n8300_8799.n294 a_n8300_8799.n293 0.189894
R790 a_n8300_8799.n293 a_n8300_8799.n292 0.189894
R791 a_n8300_8799.n292 a_n8300_8799.n273 0.189894
R792 a_n8300_8799.n274 a_n8300_8799.n273 0.189894
R793 a_n8300_8799.n287 a_n8300_8799.n274 0.189894
R794 a_n8300_8799.n287 a_n8300_8799.n286 0.189894
R795 a_n8300_8799.n286 a_n8300_8799.n285 0.189894
R796 a_n8300_8799.n285 a_n8300_8799.n276 0.189894
R797 a_n8300_8799.n277 a_n8300_8799.n276 0.189894
R798 a_n8300_8799.n280 a_n8300_8799.n277 0.189894
R799 a_n8300_8799.n35 a_n8300_8799.n32 0.189894
R800 a_n8300_8799.n39 a_n8300_8799.n32 0.189894
R801 a_n8300_8799.n40 a_n8300_8799.n39 0.189894
R802 a_n8300_8799.n41 a_n8300_8799.n40 0.189894
R803 a_n8300_8799.n41 a_n8300_8799.n30 0.189894
R804 a_n8300_8799.n45 a_n8300_8799.n30 0.189894
R805 a_n8300_8799.n46 a_n8300_8799.n45 0.189894
R806 a_n8300_8799.n47 a_n8300_8799.n46 0.189894
R807 a_n8300_8799.n47 a_n8300_8799.n28 0.189894
R808 a_n8300_8799.n51 a_n8300_8799.n28 0.189894
R809 a_n8300_8799.n52 a_n8300_8799.n51 0.189894
R810 a_n8300_8799.n53 a_n8300_8799.n52 0.189894
R811 a_n8300_8799.n53 a_n8300_8799.n26 0.189894
R812 a_n8300_8799.n57 a_n8300_8799.n26 0.189894
R813 a_n8300_8799.n58 a_n8300_8799.n57 0.189894
R814 a_n8300_8799.n59 a_n8300_8799.n58 0.189894
R815 a_n8300_8799.n59 a_n8300_8799.n24 0.189894
R816 a_n8300_8799.n63 a_n8300_8799.n24 0.189894
R817 a_n8300_8799.n64 a_n8300_8799.n63 0.189894
R818 a_n8300_8799.n65 a_n8300_8799.n64 0.189894
R819 a_n8300_8799.n65 a_n8300_8799.n22 0.189894
R820 a_n8300_8799.n69 a_n8300_8799.n22 0.189894
R821 a_n8300_8799.n83 a_n8300_8799.n80 0.189894
R822 a_n8300_8799.n87 a_n8300_8799.n80 0.189894
R823 a_n8300_8799.n88 a_n8300_8799.n87 0.189894
R824 a_n8300_8799.n89 a_n8300_8799.n88 0.189894
R825 a_n8300_8799.n89 a_n8300_8799.n78 0.189894
R826 a_n8300_8799.n93 a_n8300_8799.n78 0.189894
R827 a_n8300_8799.n94 a_n8300_8799.n93 0.189894
R828 a_n8300_8799.n95 a_n8300_8799.n94 0.189894
R829 a_n8300_8799.n95 a_n8300_8799.n76 0.189894
R830 a_n8300_8799.n99 a_n8300_8799.n76 0.189894
R831 a_n8300_8799.n100 a_n8300_8799.n99 0.189894
R832 a_n8300_8799.n101 a_n8300_8799.n100 0.189894
R833 a_n8300_8799.n101 a_n8300_8799.n74 0.189894
R834 a_n8300_8799.n105 a_n8300_8799.n74 0.189894
R835 a_n8300_8799.n106 a_n8300_8799.n105 0.189894
R836 a_n8300_8799.n107 a_n8300_8799.n106 0.189894
R837 a_n8300_8799.n107 a_n8300_8799.n72 0.189894
R838 a_n8300_8799.n111 a_n8300_8799.n72 0.189894
R839 a_n8300_8799.n112 a_n8300_8799.n111 0.189894
R840 a_n8300_8799.n113 a_n8300_8799.n112 0.189894
R841 a_n8300_8799.n113 a_n8300_8799.n70 0.189894
R842 a_n8300_8799.n117 a_n8300_8799.n70 0.189894
R843 a_n8300_8799.n132 a_n8300_8799.n129 0.189894
R844 a_n8300_8799.n136 a_n8300_8799.n129 0.189894
R845 a_n8300_8799.n137 a_n8300_8799.n136 0.189894
R846 a_n8300_8799.n138 a_n8300_8799.n137 0.189894
R847 a_n8300_8799.n138 a_n8300_8799.n127 0.189894
R848 a_n8300_8799.n142 a_n8300_8799.n127 0.189894
R849 a_n8300_8799.n143 a_n8300_8799.n142 0.189894
R850 a_n8300_8799.n144 a_n8300_8799.n143 0.189894
R851 a_n8300_8799.n144 a_n8300_8799.n125 0.189894
R852 a_n8300_8799.n148 a_n8300_8799.n125 0.189894
R853 a_n8300_8799.n149 a_n8300_8799.n148 0.189894
R854 a_n8300_8799.n150 a_n8300_8799.n149 0.189894
R855 a_n8300_8799.n150 a_n8300_8799.n123 0.189894
R856 a_n8300_8799.n154 a_n8300_8799.n123 0.189894
R857 a_n8300_8799.n155 a_n8300_8799.n154 0.189894
R858 a_n8300_8799.n156 a_n8300_8799.n155 0.189894
R859 a_n8300_8799.n156 a_n8300_8799.n121 0.189894
R860 a_n8300_8799.n160 a_n8300_8799.n121 0.189894
R861 a_n8300_8799.n161 a_n8300_8799.n160 0.189894
R862 a_n8300_8799.n162 a_n8300_8799.n161 0.189894
R863 a_n8300_8799.n162 a_n8300_8799.n119 0.189894
R864 a_n8300_8799.n166 a_n8300_8799.n119 0.189894
R865 gnd.n2473 gnd.n2140 1008.05
R866 gnd.n4444 gnd.n4443 939.716
R867 gnd.n4351 gnd.n1565 766.379
R868 gnd.n4354 gnd.n4353 766.379
R869 gnd.n3593 gnd.n3496 766.379
R870 gnd.n3589 gnd.n3494 766.379
R871 gnd.n4442 gnd.n1587 756.769
R872 gnd.n4345 gnd.n4344 756.769
R873 gnd.n3686 gnd.n3403 756.769
R874 gnd.n3684 gnd.n3406 756.769
R875 gnd.n7681 gnd.n129 751.963
R876 gnd.n7839 gnd.n7838 751.963
R877 gnd.n7175 gnd.n531 751.963
R878 gnd.n7254 gnd.n499 751.963
R879 gnd.n5351 gnd.n1178 751.963
R880 gnd.n5743 gnd.n5742 751.963
R881 gnd.n4511 gnd.n4446 751.963
R882 gnd.n4759 gnd.n1563 751.963
R883 gnd.n7836 gnd.n131 732.745
R884 gnd.n199 gnd.n127 732.745
R885 gnd.n7178 gnd.n7177 732.745
R886 gnd.n7250 gnd.n494 732.745
R887 gnd.n5740 gnd.n1180 732.745
R888 gnd.n5671 gnd.n1176 732.745
R889 gnd.n4678 gnd.n4445 732.745
R890 gnd.n4757 gnd.n4567 732.745
R891 gnd.n5789 gnd.n1098 711.122
R892 gnd.n6733 gnd.n6732 711.122
R893 gnd.n5799 gnd.n1100 711.122
R894 gnd.n7075 gnd.n655 711.122
R895 gnd.n2842 gnd.n1782 670.282
R896 gnd.n2474 gnd.n2141 670.282
R897 gnd.n7563 gnd.n336 670.282
R898 gnd.n3053 gnd.n1658 670.282
R899 gnd.n1782 gnd.n1781 585
R900 gnd.n2844 gnd.n1782 585
R901 gnd.n2847 gnd.n2846 585
R902 gnd.n2846 gnd.n2845 585
R903 gnd.n1779 gnd.n1778 585
R904 gnd.n1778 gnd.n1777 585
R905 gnd.n2852 gnd.n2851 585
R906 gnd.n2853 gnd.n2852 585
R907 gnd.n1776 gnd.n1775 585
R908 gnd.n2854 gnd.n1776 585
R909 gnd.n2857 gnd.n2856 585
R910 gnd.n2856 gnd.n2855 585
R911 gnd.n1773 gnd.n1772 585
R912 gnd.n1772 gnd.n1771 585
R913 gnd.n2862 gnd.n2861 585
R914 gnd.n2863 gnd.n2862 585
R915 gnd.n1770 gnd.n1769 585
R916 gnd.n2864 gnd.n1770 585
R917 gnd.n2867 gnd.n2866 585
R918 gnd.n2866 gnd.n2865 585
R919 gnd.n1767 gnd.n1766 585
R920 gnd.n1766 gnd.n1765 585
R921 gnd.n2872 gnd.n2871 585
R922 gnd.n2873 gnd.n2872 585
R923 gnd.n1764 gnd.n1763 585
R924 gnd.n2874 gnd.n1764 585
R925 gnd.n2877 gnd.n2876 585
R926 gnd.n2876 gnd.n2875 585
R927 gnd.n1761 gnd.n1760 585
R928 gnd.n1760 gnd.n1759 585
R929 gnd.n2882 gnd.n2881 585
R930 gnd.n2883 gnd.n2882 585
R931 gnd.n1758 gnd.n1757 585
R932 gnd.n2884 gnd.n1758 585
R933 gnd.n2887 gnd.n2886 585
R934 gnd.n2886 gnd.n2885 585
R935 gnd.n1755 gnd.n1754 585
R936 gnd.n1754 gnd.n1753 585
R937 gnd.n2892 gnd.n2891 585
R938 gnd.n2893 gnd.n2892 585
R939 gnd.n1752 gnd.n1751 585
R940 gnd.n2894 gnd.n1752 585
R941 gnd.n2897 gnd.n2896 585
R942 gnd.n2896 gnd.n2895 585
R943 gnd.n1749 gnd.n1748 585
R944 gnd.n1748 gnd.n1747 585
R945 gnd.n2902 gnd.n2901 585
R946 gnd.n2903 gnd.n2902 585
R947 gnd.n1746 gnd.n1745 585
R948 gnd.n2904 gnd.n1746 585
R949 gnd.n2907 gnd.n2906 585
R950 gnd.n2906 gnd.n2905 585
R951 gnd.n1743 gnd.n1742 585
R952 gnd.n1742 gnd.n1741 585
R953 gnd.n2912 gnd.n2911 585
R954 gnd.n2913 gnd.n2912 585
R955 gnd.n1740 gnd.n1739 585
R956 gnd.n2914 gnd.n1740 585
R957 gnd.n2917 gnd.n2916 585
R958 gnd.n2916 gnd.n2915 585
R959 gnd.n1737 gnd.n1736 585
R960 gnd.n1736 gnd.n1735 585
R961 gnd.n2922 gnd.n2921 585
R962 gnd.n2923 gnd.n2922 585
R963 gnd.n1734 gnd.n1733 585
R964 gnd.n2924 gnd.n1734 585
R965 gnd.n2927 gnd.n2926 585
R966 gnd.n2926 gnd.n2925 585
R967 gnd.n1731 gnd.n1730 585
R968 gnd.n1730 gnd.n1729 585
R969 gnd.n2932 gnd.n2931 585
R970 gnd.n2933 gnd.n2932 585
R971 gnd.n1728 gnd.n1727 585
R972 gnd.n2934 gnd.n1728 585
R973 gnd.n2937 gnd.n2936 585
R974 gnd.n2936 gnd.n2935 585
R975 gnd.n1725 gnd.n1724 585
R976 gnd.n1724 gnd.n1723 585
R977 gnd.n2942 gnd.n2941 585
R978 gnd.n2943 gnd.n2942 585
R979 gnd.n1722 gnd.n1721 585
R980 gnd.n2944 gnd.n1722 585
R981 gnd.n2947 gnd.n2946 585
R982 gnd.n2946 gnd.n2945 585
R983 gnd.n1719 gnd.n1718 585
R984 gnd.n1718 gnd.n1717 585
R985 gnd.n2952 gnd.n2951 585
R986 gnd.n2953 gnd.n2952 585
R987 gnd.n1716 gnd.n1715 585
R988 gnd.n2954 gnd.n1716 585
R989 gnd.n2957 gnd.n2956 585
R990 gnd.n2956 gnd.n2955 585
R991 gnd.n1713 gnd.n1712 585
R992 gnd.n1712 gnd.n1711 585
R993 gnd.n2962 gnd.n2961 585
R994 gnd.n2963 gnd.n2962 585
R995 gnd.n1710 gnd.n1709 585
R996 gnd.n2964 gnd.n1710 585
R997 gnd.n2967 gnd.n2966 585
R998 gnd.n2966 gnd.n2965 585
R999 gnd.n1707 gnd.n1706 585
R1000 gnd.n1706 gnd.n1705 585
R1001 gnd.n2972 gnd.n2971 585
R1002 gnd.n2973 gnd.n2972 585
R1003 gnd.n1704 gnd.n1703 585
R1004 gnd.n2974 gnd.n1704 585
R1005 gnd.n2977 gnd.n2976 585
R1006 gnd.n2976 gnd.n2975 585
R1007 gnd.n1701 gnd.n1700 585
R1008 gnd.n1700 gnd.n1699 585
R1009 gnd.n2982 gnd.n2981 585
R1010 gnd.n2983 gnd.n2982 585
R1011 gnd.n1698 gnd.n1697 585
R1012 gnd.n2984 gnd.n1698 585
R1013 gnd.n2987 gnd.n2986 585
R1014 gnd.n2986 gnd.n2985 585
R1015 gnd.n1695 gnd.n1694 585
R1016 gnd.n1694 gnd.n1693 585
R1017 gnd.n2992 gnd.n2991 585
R1018 gnd.n2993 gnd.n2992 585
R1019 gnd.n1692 gnd.n1691 585
R1020 gnd.n2994 gnd.n1692 585
R1021 gnd.n2997 gnd.n2996 585
R1022 gnd.n2996 gnd.n2995 585
R1023 gnd.n1689 gnd.n1688 585
R1024 gnd.n1688 gnd.n1687 585
R1025 gnd.n3002 gnd.n3001 585
R1026 gnd.n3003 gnd.n3002 585
R1027 gnd.n1686 gnd.n1685 585
R1028 gnd.n3004 gnd.n1686 585
R1029 gnd.n3007 gnd.n3006 585
R1030 gnd.n3006 gnd.n3005 585
R1031 gnd.n1683 gnd.n1682 585
R1032 gnd.n1682 gnd.n1681 585
R1033 gnd.n3012 gnd.n3011 585
R1034 gnd.n3013 gnd.n3012 585
R1035 gnd.n1680 gnd.n1679 585
R1036 gnd.n3014 gnd.n1680 585
R1037 gnd.n3017 gnd.n3016 585
R1038 gnd.n3016 gnd.n3015 585
R1039 gnd.n1677 gnd.n1676 585
R1040 gnd.n1676 gnd.n1675 585
R1041 gnd.n3022 gnd.n3021 585
R1042 gnd.n3023 gnd.n3022 585
R1043 gnd.n1674 gnd.n1673 585
R1044 gnd.n3024 gnd.n1674 585
R1045 gnd.n3027 gnd.n3026 585
R1046 gnd.n3026 gnd.n3025 585
R1047 gnd.n1671 gnd.n1670 585
R1048 gnd.n1670 gnd.n1669 585
R1049 gnd.n3032 gnd.n3031 585
R1050 gnd.n3033 gnd.n3032 585
R1051 gnd.n1668 gnd.n1667 585
R1052 gnd.n3034 gnd.n1668 585
R1053 gnd.n3037 gnd.n3036 585
R1054 gnd.n3036 gnd.n3035 585
R1055 gnd.n1665 gnd.n1664 585
R1056 gnd.n1664 gnd.n1663 585
R1057 gnd.n3042 gnd.n3041 585
R1058 gnd.n3043 gnd.n3042 585
R1059 gnd.n1662 gnd.n1661 585
R1060 gnd.n3044 gnd.n1662 585
R1061 gnd.n3047 gnd.n3046 585
R1062 gnd.n3046 gnd.n3045 585
R1063 gnd.n1659 gnd.n1657 585
R1064 gnd.n1657 gnd.n1656 585
R1065 gnd.n3059 gnd.n3058 585
R1066 gnd.n3060 gnd.n3059 585
R1067 gnd.n2842 gnd.n2841 585
R1068 gnd.n2843 gnd.n2842 585
R1069 gnd.n1785 gnd.n1784 585
R1070 gnd.n1784 gnd.n1783 585
R1071 gnd.n2837 gnd.n2836 585
R1072 gnd.n2836 gnd.n2835 585
R1073 gnd.n1788 gnd.n1787 585
R1074 gnd.n2834 gnd.n1788 585
R1075 gnd.n2832 gnd.n2831 585
R1076 gnd.n2833 gnd.n2832 585
R1077 gnd.n2830 gnd.n1790 585
R1078 gnd.n1790 gnd.n1789 585
R1079 gnd.n2829 gnd.n2828 585
R1080 gnd.n2828 gnd.n2827 585
R1081 gnd.n1795 gnd.n1794 585
R1082 gnd.n2826 gnd.n1795 585
R1083 gnd.n2824 gnd.n2823 585
R1084 gnd.n2825 gnd.n2824 585
R1085 gnd.n2822 gnd.n1797 585
R1086 gnd.n1797 gnd.n1796 585
R1087 gnd.n2821 gnd.n2820 585
R1088 gnd.n2820 gnd.n2819 585
R1089 gnd.n1803 gnd.n1802 585
R1090 gnd.n2818 gnd.n1803 585
R1091 gnd.n2816 gnd.n2815 585
R1092 gnd.n2817 gnd.n2816 585
R1093 gnd.n2814 gnd.n1805 585
R1094 gnd.n1805 gnd.n1804 585
R1095 gnd.n2813 gnd.n2812 585
R1096 gnd.n2812 gnd.n2811 585
R1097 gnd.n1811 gnd.n1810 585
R1098 gnd.n2810 gnd.n1811 585
R1099 gnd.n2808 gnd.n2807 585
R1100 gnd.n2809 gnd.n2808 585
R1101 gnd.n2806 gnd.n1813 585
R1102 gnd.n1813 gnd.n1812 585
R1103 gnd.n2805 gnd.n2804 585
R1104 gnd.n2804 gnd.n2803 585
R1105 gnd.n1819 gnd.n1818 585
R1106 gnd.n2802 gnd.n1819 585
R1107 gnd.n2800 gnd.n2799 585
R1108 gnd.n2801 gnd.n2800 585
R1109 gnd.n2798 gnd.n1821 585
R1110 gnd.n1821 gnd.n1820 585
R1111 gnd.n2797 gnd.n2796 585
R1112 gnd.n2796 gnd.n2795 585
R1113 gnd.n1827 gnd.n1826 585
R1114 gnd.n2794 gnd.n1827 585
R1115 gnd.n2792 gnd.n2791 585
R1116 gnd.n2793 gnd.n2792 585
R1117 gnd.n2790 gnd.n1829 585
R1118 gnd.n1829 gnd.n1828 585
R1119 gnd.n2789 gnd.n2788 585
R1120 gnd.n2788 gnd.n2787 585
R1121 gnd.n1835 gnd.n1834 585
R1122 gnd.n2786 gnd.n1835 585
R1123 gnd.n2784 gnd.n2783 585
R1124 gnd.n2785 gnd.n2784 585
R1125 gnd.n2782 gnd.n1837 585
R1126 gnd.n1837 gnd.n1836 585
R1127 gnd.n2781 gnd.n2780 585
R1128 gnd.n2780 gnd.n2779 585
R1129 gnd.n1843 gnd.n1842 585
R1130 gnd.n2778 gnd.n1843 585
R1131 gnd.n2776 gnd.n2775 585
R1132 gnd.n2777 gnd.n2776 585
R1133 gnd.n2774 gnd.n1845 585
R1134 gnd.n1845 gnd.n1844 585
R1135 gnd.n2773 gnd.n2772 585
R1136 gnd.n2772 gnd.n2771 585
R1137 gnd.n1851 gnd.n1850 585
R1138 gnd.n2770 gnd.n1851 585
R1139 gnd.n2768 gnd.n2767 585
R1140 gnd.n2769 gnd.n2768 585
R1141 gnd.n2766 gnd.n1853 585
R1142 gnd.n1853 gnd.n1852 585
R1143 gnd.n2765 gnd.n2764 585
R1144 gnd.n2764 gnd.n2763 585
R1145 gnd.n1859 gnd.n1858 585
R1146 gnd.n2762 gnd.n1859 585
R1147 gnd.n2760 gnd.n2759 585
R1148 gnd.n2761 gnd.n2760 585
R1149 gnd.n2758 gnd.n1861 585
R1150 gnd.n1861 gnd.n1860 585
R1151 gnd.n2757 gnd.n2756 585
R1152 gnd.n2756 gnd.n2755 585
R1153 gnd.n1867 gnd.n1866 585
R1154 gnd.n2754 gnd.n1867 585
R1155 gnd.n2752 gnd.n2751 585
R1156 gnd.n2753 gnd.n2752 585
R1157 gnd.n2750 gnd.n1869 585
R1158 gnd.n1869 gnd.n1868 585
R1159 gnd.n2749 gnd.n2748 585
R1160 gnd.n2748 gnd.n2747 585
R1161 gnd.n1875 gnd.n1874 585
R1162 gnd.n2746 gnd.n1875 585
R1163 gnd.n2744 gnd.n2743 585
R1164 gnd.n2745 gnd.n2744 585
R1165 gnd.n2742 gnd.n1877 585
R1166 gnd.n1877 gnd.n1876 585
R1167 gnd.n2741 gnd.n2740 585
R1168 gnd.n2740 gnd.n2739 585
R1169 gnd.n1883 gnd.n1882 585
R1170 gnd.n2738 gnd.n1883 585
R1171 gnd.n2736 gnd.n2735 585
R1172 gnd.n2737 gnd.n2736 585
R1173 gnd.n2734 gnd.n1885 585
R1174 gnd.n1885 gnd.n1884 585
R1175 gnd.n2733 gnd.n2732 585
R1176 gnd.n2732 gnd.n2731 585
R1177 gnd.n1891 gnd.n1890 585
R1178 gnd.n2730 gnd.n1891 585
R1179 gnd.n2728 gnd.n2727 585
R1180 gnd.n2729 gnd.n2728 585
R1181 gnd.n2726 gnd.n1893 585
R1182 gnd.n1893 gnd.n1892 585
R1183 gnd.n2725 gnd.n2724 585
R1184 gnd.n2724 gnd.n2723 585
R1185 gnd.n1899 gnd.n1898 585
R1186 gnd.n2722 gnd.n1899 585
R1187 gnd.n2720 gnd.n2719 585
R1188 gnd.n2721 gnd.n2720 585
R1189 gnd.n2718 gnd.n1901 585
R1190 gnd.n1901 gnd.n1900 585
R1191 gnd.n2717 gnd.n2716 585
R1192 gnd.n2716 gnd.n2715 585
R1193 gnd.n1907 gnd.n1906 585
R1194 gnd.n2714 gnd.n1907 585
R1195 gnd.n2712 gnd.n2711 585
R1196 gnd.n2713 gnd.n2712 585
R1197 gnd.n2710 gnd.n1909 585
R1198 gnd.n1909 gnd.n1908 585
R1199 gnd.n2709 gnd.n2708 585
R1200 gnd.n2708 gnd.n2707 585
R1201 gnd.n1915 gnd.n1914 585
R1202 gnd.n2706 gnd.n1915 585
R1203 gnd.n2704 gnd.n2703 585
R1204 gnd.n2705 gnd.n2704 585
R1205 gnd.n2702 gnd.n1917 585
R1206 gnd.n1917 gnd.n1916 585
R1207 gnd.n2701 gnd.n2700 585
R1208 gnd.n2700 gnd.n2699 585
R1209 gnd.n1923 gnd.n1922 585
R1210 gnd.n2698 gnd.n1923 585
R1211 gnd.n2696 gnd.n2695 585
R1212 gnd.n2697 gnd.n2696 585
R1213 gnd.n2694 gnd.n1925 585
R1214 gnd.n1925 gnd.n1924 585
R1215 gnd.n2693 gnd.n2692 585
R1216 gnd.n2692 gnd.n2691 585
R1217 gnd.n1931 gnd.n1930 585
R1218 gnd.n2690 gnd.n1931 585
R1219 gnd.n2688 gnd.n2687 585
R1220 gnd.n2689 gnd.n2688 585
R1221 gnd.n2686 gnd.n1933 585
R1222 gnd.n1933 gnd.n1932 585
R1223 gnd.n2685 gnd.n2684 585
R1224 gnd.n2684 gnd.n2683 585
R1225 gnd.n1939 gnd.n1938 585
R1226 gnd.n2682 gnd.n1939 585
R1227 gnd.n2680 gnd.n2679 585
R1228 gnd.n2681 gnd.n2680 585
R1229 gnd.n2678 gnd.n1941 585
R1230 gnd.n1941 gnd.n1940 585
R1231 gnd.n2677 gnd.n2676 585
R1232 gnd.n2676 gnd.n2675 585
R1233 gnd.n1947 gnd.n1946 585
R1234 gnd.n2674 gnd.n1947 585
R1235 gnd.n2672 gnd.n2671 585
R1236 gnd.n2673 gnd.n2672 585
R1237 gnd.n2670 gnd.n1949 585
R1238 gnd.n1949 gnd.n1948 585
R1239 gnd.n2669 gnd.n2668 585
R1240 gnd.n2668 gnd.n2667 585
R1241 gnd.n1955 gnd.n1954 585
R1242 gnd.n2666 gnd.n1955 585
R1243 gnd.n2664 gnd.n2663 585
R1244 gnd.n2665 gnd.n2664 585
R1245 gnd.n2662 gnd.n1957 585
R1246 gnd.n1957 gnd.n1956 585
R1247 gnd.n2661 gnd.n2660 585
R1248 gnd.n2660 gnd.n2659 585
R1249 gnd.n1963 gnd.n1962 585
R1250 gnd.n2658 gnd.n1963 585
R1251 gnd.n2656 gnd.n2655 585
R1252 gnd.n2657 gnd.n2656 585
R1253 gnd.n2654 gnd.n1965 585
R1254 gnd.n1965 gnd.n1964 585
R1255 gnd.n2653 gnd.n2652 585
R1256 gnd.n2652 gnd.n2651 585
R1257 gnd.n1971 gnd.n1970 585
R1258 gnd.n2650 gnd.n1971 585
R1259 gnd.n2648 gnd.n2647 585
R1260 gnd.n2649 gnd.n2648 585
R1261 gnd.n2646 gnd.n1973 585
R1262 gnd.n1973 gnd.n1972 585
R1263 gnd.n2645 gnd.n2644 585
R1264 gnd.n2644 gnd.n2643 585
R1265 gnd.n1979 gnd.n1978 585
R1266 gnd.n2642 gnd.n1979 585
R1267 gnd.n2640 gnd.n2639 585
R1268 gnd.n2641 gnd.n2640 585
R1269 gnd.n2638 gnd.n1981 585
R1270 gnd.n1981 gnd.n1980 585
R1271 gnd.n2637 gnd.n2636 585
R1272 gnd.n2636 gnd.n2635 585
R1273 gnd.n1987 gnd.n1986 585
R1274 gnd.n2634 gnd.n1987 585
R1275 gnd.n2632 gnd.n2631 585
R1276 gnd.n2633 gnd.n2632 585
R1277 gnd.n2630 gnd.n1989 585
R1278 gnd.n1989 gnd.n1988 585
R1279 gnd.n2629 gnd.n2628 585
R1280 gnd.n2628 gnd.n2627 585
R1281 gnd.n1995 gnd.n1994 585
R1282 gnd.n2626 gnd.n1995 585
R1283 gnd.n2624 gnd.n2623 585
R1284 gnd.n2625 gnd.n2624 585
R1285 gnd.n2622 gnd.n1997 585
R1286 gnd.n1997 gnd.n1996 585
R1287 gnd.n2621 gnd.n2620 585
R1288 gnd.n2620 gnd.n2619 585
R1289 gnd.n2003 gnd.n2002 585
R1290 gnd.n2618 gnd.n2003 585
R1291 gnd.n2616 gnd.n2615 585
R1292 gnd.n2617 gnd.n2616 585
R1293 gnd.n2614 gnd.n2005 585
R1294 gnd.n2005 gnd.n2004 585
R1295 gnd.n2613 gnd.n2612 585
R1296 gnd.n2612 gnd.n2611 585
R1297 gnd.n2011 gnd.n2010 585
R1298 gnd.n2610 gnd.n2011 585
R1299 gnd.n2608 gnd.n2607 585
R1300 gnd.n2609 gnd.n2608 585
R1301 gnd.n2606 gnd.n2013 585
R1302 gnd.n2013 gnd.n2012 585
R1303 gnd.n2605 gnd.n2604 585
R1304 gnd.n2604 gnd.n2603 585
R1305 gnd.n2019 gnd.n2018 585
R1306 gnd.n2602 gnd.n2019 585
R1307 gnd.n2600 gnd.n2599 585
R1308 gnd.n2601 gnd.n2600 585
R1309 gnd.n2598 gnd.n2021 585
R1310 gnd.n2021 gnd.n2020 585
R1311 gnd.n2597 gnd.n2596 585
R1312 gnd.n2596 gnd.n2595 585
R1313 gnd.n2027 gnd.n2026 585
R1314 gnd.n2594 gnd.n2027 585
R1315 gnd.n2592 gnd.n2591 585
R1316 gnd.n2593 gnd.n2592 585
R1317 gnd.n2590 gnd.n2029 585
R1318 gnd.n2029 gnd.n2028 585
R1319 gnd.n2589 gnd.n2588 585
R1320 gnd.n2588 gnd.n2587 585
R1321 gnd.n2035 gnd.n2034 585
R1322 gnd.n2586 gnd.n2035 585
R1323 gnd.n2584 gnd.n2583 585
R1324 gnd.n2585 gnd.n2584 585
R1325 gnd.n2582 gnd.n2037 585
R1326 gnd.n2037 gnd.n2036 585
R1327 gnd.n2581 gnd.n2580 585
R1328 gnd.n2580 gnd.n2579 585
R1329 gnd.n2043 gnd.n2042 585
R1330 gnd.n2578 gnd.n2043 585
R1331 gnd.n2576 gnd.n2575 585
R1332 gnd.n2577 gnd.n2576 585
R1333 gnd.n2574 gnd.n2045 585
R1334 gnd.n2045 gnd.n2044 585
R1335 gnd.n2573 gnd.n2572 585
R1336 gnd.n2572 gnd.n2571 585
R1337 gnd.n2051 gnd.n2050 585
R1338 gnd.n2570 gnd.n2051 585
R1339 gnd.n2568 gnd.n2567 585
R1340 gnd.n2569 gnd.n2568 585
R1341 gnd.n2566 gnd.n2053 585
R1342 gnd.n2053 gnd.n2052 585
R1343 gnd.n2565 gnd.n2564 585
R1344 gnd.n2564 gnd.n2563 585
R1345 gnd.n2059 gnd.n2058 585
R1346 gnd.n2562 gnd.n2059 585
R1347 gnd.n2560 gnd.n2559 585
R1348 gnd.n2561 gnd.n2560 585
R1349 gnd.n2558 gnd.n2061 585
R1350 gnd.n2061 gnd.n2060 585
R1351 gnd.n2557 gnd.n2556 585
R1352 gnd.n2556 gnd.n2555 585
R1353 gnd.n2067 gnd.n2066 585
R1354 gnd.n2554 gnd.n2067 585
R1355 gnd.n2552 gnd.n2551 585
R1356 gnd.n2553 gnd.n2552 585
R1357 gnd.n2550 gnd.n2069 585
R1358 gnd.n2069 gnd.n2068 585
R1359 gnd.n2549 gnd.n2548 585
R1360 gnd.n2548 gnd.n2547 585
R1361 gnd.n2075 gnd.n2074 585
R1362 gnd.n2546 gnd.n2075 585
R1363 gnd.n2544 gnd.n2543 585
R1364 gnd.n2545 gnd.n2544 585
R1365 gnd.n2542 gnd.n2077 585
R1366 gnd.n2077 gnd.n2076 585
R1367 gnd.n2541 gnd.n2540 585
R1368 gnd.n2540 gnd.n2539 585
R1369 gnd.n2083 gnd.n2082 585
R1370 gnd.n2538 gnd.n2083 585
R1371 gnd.n2536 gnd.n2535 585
R1372 gnd.n2537 gnd.n2536 585
R1373 gnd.n2534 gnd.n2085 585
R1374 gnd.n2085 gnd.n2084 585
R1375 gnd.n2533 gnd.n2532 585
R1376 gnd.n2532 gnd.n2531 585
R1377 gnd.n2091 gnd.n2090 585
R1378 gnd.n2530 gnd.n2091 585
R1379 gnd.n2528 gnd.n2527 585
R1380 gnd.n2529 gnd.n2528 585
R1381 gnd.n2526 gnd.n2093 585
R1382 gnd.n2093 gnd.n2092 585
R1383 gnd.n2525 gnd.n2524 585
R1384 gnd.n2524 gnd.n2523 585
R1385 gnd.n2099 gnd.n2098 585
R1386 gnd.n2522 gnd.n2099 585
R1387 gnd.n2520 gnd.n2519 585
R1388 gnd.n2521 gnd.n2520 585
R1389 gnd.n2518 gnd.n2101 585
R1390 gnd.n2101 gnd.n2100 585
R1391 gnd.n2517 gnd.n2516 585
R1392 gnd.n2516 gnd.n2515 585
R1393 gnd.n2107 gnd.n2106 585
R1394 gnd.n2514 gnd.n2107 585
R1395 gnd.n2512 gnd.n2511 585
R1396 gnd.n2513 gnd.n2512 585
R1397 gnd.n2510 gnd.n2109 585
R1398 gnd.n2109 gnd.n2108 585
R1399 gnd.n2509 gnd.n2508 585
R1400 gnd.n2508 gnd.n2507 585
R1401 gnd.n2115 gnd.n2114 585
R1402 gnd.n2506 gnd.n2115 585
R1403 gnd.n2504 gnd.n2503 585
R1404 gnd.n2505 gnd.n2504 585
R1405 gnd.n2502 gnd.n2117 585
R1406 gnd.n2117 gnd.n2116 585
R1407 gnd.n2501 gnd.n2500 585
R1408 gnd.n2500 gnd.n2499 585
R1409 gnd.n2123 gnd.n2122 585
R1410 gnd.n2498 gnd.n2123 585
R1411 gnd.n2496 gnd.n2495 585
R1412 gnd.n2497 gnd.n2496 585
R1413 gnd.n2494 gnd.n2125 585
R1414 gnd.n2125 gnd.n2124 585
R1415 gnd.n2493 gnd.n2492 585
R1416 gnd.n2492 gnd.n2491 585
R1417 gnd.n2131 gnd.n2130 585
R1418 gnd.n2490 gnd.n2131 585
R1419 gnd.n2488 gnd.n2487 585
R1420 gnd.n2489 gnd.n2488 585
R1421 gnd.n2486 gnd.n2133 585
R1422 gnd.n2133 gnd.n2132 585
R1423 gnd.n2485 gnd.n2484 585
R1424 gnd.n2484 gnd.n2483 585
R1425 gnd.n2139 gnd.n2138 585
R1426 gnd.n2482 gnd.n2139 585
R1427 gnd.n2480 gnd.n2479 585
R1428 gnd.n2481 gnd.n2480 585
R1429 gnd.n2478 gnd.n2141 585
R1430 gnd.n2141 gnd.n2140 585
R1431 gnd.n337 gnd.n335 585
R1432 gnd.n2306 gnd.n335 585
R1433 gnd.n2310 gnd.n2309 585
R1434 gnd.n2311 gnd.n2310 585
R1435 gnd.n2305 gnd.n2304 585
R1436 gnd.n2312 gnd.n2305 585
R1437 gnd.n2315 gnd.n2314 585
R1438 gnd.n2314 gnd.n2313 585
R1439 gnd.n2316 gnd.n2299 585
R1440 gnd.n2299 gnd.n2298 585
R1441 gnd.n2318 gnd.n2317 585
R1442 gnd.n2319 gnd.n2318 585
R1443 gnd.n2297 gnd.n2296 585
R1444 gnd.n2320 gnd.n2297 585
R1445 gnd.n2323 gnd.n2322 585
R1446 gnd.n2322 gnd.n2321 585
R1447 gnd.n2324 gnd.n2291 585
R1448 gnd.n2291 gnd.n2290 585
R1449 gnd.n2326 gnd.n2325 585
R1450 gnd.n2327 gnd.n2326 585
R1451 gnd.n2289 gnd.n2288 585
R1452 gnd.n2328 gnd.n2289 585
R1453 gnd.n2331 gnd.n2330 585
R1454 gnd.n2330 gnd.n2329 585
R1455 gnd.n2332 gnd.n2283 585
R1456 gnd.n2283 gnd.n2282 585
R1457 gnd.n2334 gnd.n2333 585
R1458 gnd.n2335 gnd.n2334 585
R1459 gnd.n2281 gnd.n2280 585
R1460 gnd.n2336 gnd.n2281 585
R1461 gnd.n2339 gnd.n2338 585
R1462 gnd.n2338 gnd.n2337 585
R1463 gnd.n2340 gnd.n2275 585
R1464 gnd.n2275 gnd.n2274 585
R1465 gnd.n2342 gnd.n2341 585
R1466 gnd.n2343 gnd.n2342 585
R1467 gnd.n2273 gnd.n2272 585
R1468 gnd.n2344 gnd.n2273 585
R1469 gnd.n2347 gnd.n2346 585
R1470 gnd.n2346 gnd.n2345 585
R1471 gnd.n2348 gnd.n2267 585
R1472 gnd.n2267 gnd.n2266 585
R1473 gnd.n2350 gnd.n2349 585
R1474 gnd.n2351 gnd.n2350 585
R1475 gnd.n2265 gnd.n2264 585
R1476 gnd.n2352 gnd.n2265 585
R1477 gnd.n2355 gnd.n2354 585
R1478 gnd.n2354 gnd.n2353 585
R1479 gnd.n2356 gnd.n2259 585
R1480 gnd.n2259 gnd.n2258 585
R1481 gnd.n2358 gnd.n2357 585
R1482 gnd.n2359 gnd.n2358 585
R1483 gnd.n2257 gnd.n2256 585
R1484 gnd.n2360 gnd.n2257 585
R1485 gnd.n2363 gnd.n2362 585
R1486 gnd.n2362 gnd.n2361 585
R1487 gnd.n2364 gnd.n2251 585
R1488 gnd.n2251 gnd.n2250 585
R1489 gnd.n2366 gnd.n2365 585
R1490 gnd.n2367 gnd.n2366 585
R1491 gnd.n2249 gnd.n2248 585
R1492 gnd.n2368 gnd.n2249 585
R1493 gnd.n2371 gnd.n2370 585
R1494 gnd.n2370 gnd.n2369 585
R1495 gnd.n2372 gnd.n2243 585
R1496 gnd.n2243 gnd.n2242 585
R1497 gnd.n2374 gnd.n2373 585
R1498 gnd.n2375 gnd.n2374 585
R1499 gnd.n2241 gnd.n2240 585
R1500 gnd.n2376 gnd.n2241 585
R1501 gnd.n2379 gnd.n2378 585
R1502 gnd.n2378 gnd.n2377 585
R1503 gnd.n2380 gnd.n2235 585
R1504 gnd.n2235 gnd.n2234 585
R1505 gnd.n2382 gnd.n2381 585
R1506 gnd.n2383 gnd.n2382 585
R1507 gnd.n2233 gnd.n2232 585
R1508 gnd.n2384 gnd.n2233 585
R1509 gnd.n2387 gnd.n2386 585
R1510 gnd.n2386 gnd.n2385 585
R1511 gnd.n2388 gnd.n2227 585
R1512 gnd.n2227 gnd.n2226 585
R1513 gnd.n2390 gnd.n2389 585
R1514 gnd.n2391 gnd.n2390 585
R1515 gnd.n2225 gnd.n2224 585
R1516 gnd.n2392 gnd.n2225 585
R1517 gnd.n2395 gnd.n2394 585
R1518 gnd.n2394 gnd.n2393 585
R1519 gnd.n2396 gnd.n2219 585
R1520 gnd.n2219 gnd.n2218 585
R1521 gnd.n2398 gnd.n2397 585
R1522 gnd.n2399 gnd.n2398 585
R1523 gnd.n2217 gnd.n2216 585
R1524 gnd.n2400 gnd.n2217 585
R1525 gnd.n2403 gnd.n2402 585
R1526 gnd.n2402 gnd.n2401 585
R1527 gnd.n2404 gnd.n2211 585
R1528 gnd.n2211 gnd.n2210 585
R1529 gnd.n2406 gnd.n2405 585
R1530 gnd.n2407 gnd.n2406 585
R1531 gnd.n2209 gnd.n2208 585
R1532 gnd.n2408 gnd.n2209 585
R1533 gnd.n2411 gnd.n2410 585
R1534 gnd.n2410 gnd.n2409 585
R1535 gnd.n2412 gnd.n2203 585
R1536 gnd.n2203 gnd.n2202 585
R1537 gnd.n2414 gnd.n2413 585
R1538 gnd.n2415 gnd.n2414 585
R1539 gnd.n2201 gnd.n2200 585
R1540 gnd.n2416 gnd.n2201 585
R1541 gnd.n2419 gnd.n2418 585
R1542 gnd.n2418 gnd.n2417 585
R1543 gnd.n2420 gnd.n2195 585
R1544 gnd.n2195 gnd.n2194 585
R1545 gnd.n2422 gnd.n2421 585
R1546 gnd.n2423 gnd.n2422 585
R1547 gnd.n2193 gnd.n2192 585
R1548 gnd.n2424 gnd.n2193 585
R1549 gnd.n2427 gnd.n2426 585
R1550 gnd.n2426 gnd.n2425 585
R1551 gnd.n2428 gnd.n2187 585
R1552 gnd.n2187 gnd.n2186 585
R1553 gnd.n2430 gnd.n2429 585
R1554 gnd.n2431 gnd.n2430 585
R1555 gnd.n2185 gnd.n2184 585
R1556 gnd.n2432 gnd.n2185 585
R1557 gnd.n2435 gnd.n2434 585
R1558 gnd.n2434 gnd.n2433 585
R1559 gnd.n2436 gnd.n2179 585
R1560 gnd.n2179 gnd.n2178 585
R1561 gnd.n2438 gnd.n2437 585
R1562 gnd.n2439 gnd.n2438 585
R1563 gnd.n2177 gnd.n2176 585
R1564 gnd.n2440 gnd.n2177 585
R1565 gnd.n2443 gnd.n2442 585
R1566 gnd.n2442 gnd.n2441 585
R1567 gnd.n2444 gnd.n2171 585
R1568 gnd.n2171 gnd.n2170 585
R1569 gnd.n2446 gnd.n2445 585
R1570 gnd.n2447 gnd.n2446 585
R1571 gnd.n2169 gnd.n2168 585
R1572 gnd.n2448 gnd.n2169 585
R1573 gnd.n2451 gnd.n2450 585
R1574 gnd.n2450 gnd.n2449 585
R1575 gnd.n2452 gnd.n2163 585
R1576 gnd.n2163 gnd.n2162 585
R1577 gnd.n2454 gnd.n2453 585
R1578 gnd.n2455 gnd.n2454 585
R1579 gnd.n2161 gnd.n2160 585
R1580 gnd.n2456 gnd.n2161 585
R1581 gnd.n2459 gnd.n2458 585
R1582 gnd.n2458 gnd.n2457 585
R1583 gnd.n2460 gnd.n2155 585
R1584 gnd.n2155 gnd.n2154 585
R1585 gnd.n2462 gnd.n2461 585
R1586 gnd.n2463 gnd.n2462 585
R1587 gnd.n2153 gnd.n2152 585
R1588 gnd.n2464 gnd.n2153 585
R1589 gnd.n2467 gnd.n2466 585
R1590 gnd.n2466 gnd.n2465 585
R1591 gnd.n2468 gnd.n2148 585
R1592 gnd.n2148 gnd.n2147 585
R1593 gnd.n2470 gnd.n2469 585
R1594 gnd.n2471 gnd.n2470 585
R1595 gnd.n2146 gnd.n2145 585
R1596 gnd.n2472 gnd.n2146 585
R1597 gnd.n2475 gnd.n2474 585
R1598 gnd.n2474 gnd.n2473 585
R1599 gnd.n5661 gnd.n1178 585
R1600 gnd.n5741 gnd.n1178 585
R1601 gnd.n5663 gnd.n5662 585
R1602 gnd.n5664 gnd.n5663 585
R1603 gnd.n1267 gnd.n1266 585
R1604 gnd.n5152 gnd.n1266 585
R1605 gnd.n5346 gnd.n5345 585
R1606 gnd.n5345 gnd.n5344 585
R1607 gnd.n1270 gnd.n1269 585
R1608 gnd.n5118 gnd.n1270 585
R1609 gnd.n5333 gnd.n5332 585
R1610 gnd.n5334 gnd.n5333 585
R1611 gnd.n1286 gnd.n1285 585
R1612 gnd.n5107 gnd.n1285 585
R1613 gnd.n5328 gnd.n5327 585
R1614 gnd.n5327 gnd.n5326 585
R1615 gnd.n1289 gnd.n1288 585
R1616 gnd.n5103 gnd.n1289 585
R1617 gnd.n5317 gnd.n5316 585
R1618 gnd.n5318 gnd.n5317 585
R1619 gnd.n1303 gnd.n1302 585
R1620 gnd.n5097 gnd.n1302 585
R1621 gnd.n5312 gnd.n5311 585
R1622 gnd.n5311 gnd.n5310 585
R1623 gnd.n1306 gnd.n1305 585
R1624 gnd.n5019 gnd.n1306 585
R1625 gnd.n5301 gnd.n5300 585
R1626 gnd.n5302 gnd.n5301 585
R1627 gnd.n1321 gnd.n1320 585
R1628 gnd.n5023 gnd.n1320 585
R1629 gnd.n5296 gnd.n5295 585
R1630 gnd.n5295 gnd.n5294 585
R1631 gnd.n1324 gnd.n1323 585
R1632 gnd.n5027 gnd.n1324 585
R1633 gnd.n5285 gnd.n5284 585
R1634 gnd.n5286 gnd.n5285 585
R1635 gnd.n1338 gnd.n1337 585
R1636 gnd.n5033 gnd.n1337 585
R1637 gnd.n5280 gnd.n5279 585
R1638 gnd.n5279 gnd.n5278 585
R1639 gnd.n1341 gnd.n1340 585
R1640 gnd.n5007 gnd.n1341 585
R1641 gnd.n5269 gnd.n5268 585
R1642 gnd.n5270 gnd.n5269 585
R1643 gnd.n1356 gnd.n1355 585
R1644 gnd.n5003 gnd.n1355 585
R1645 gnd.n5264 gnd.n5263 585
R1646 gnd.n5263 gnd.n5262 585
R1647 gnd.n1359 gnd.n1358 585
R1648 gnd.n4997 gnd.n1359 585
R1649 gnd.n5253 gnd.n5252 585
R1650 gnd.n5254 gnd.n5253 585
R1651 gnd.n1373 gnd.n1372 585
R1652 gnd.n4993 gnd.n1372 585
R1653 gnd.n5248 gnd.n5247 585
R1654 gnd.n5247 gnd.n5246 585
R1655 gnd.n1376 gnd.n1375 585
R1656 gnd.n5197 gnd.n1376 585
R1657 gnd.n5214 gnd.n5213 585
R1658 gnd.n5219 gnd.n5214 585
R1659 gnd.n1427 gnd.n1426 585
R1660 gnd.n1426 gnd.n1422 585
R1661 gnd.n5209 gnd.n5208 585
R1662 gnd.n5208 gnd.n1412 585
R1663 gnd.n1403 gnd.n1402 585
R1664 gnd.n5227 gnd.n1403 585
R1665 gnd.n5234 gnd.n5233 585
R1666 gnd.n5233 gnd.n5232 585
R1667 gnd.n5235 gnd.n1397 585
R1668 gnd.n1397 gnd.n1395 585
R1669 gnd.n5237 gnd.n5236 585
R1670 gnd.n5238 gnd.n5237 585
R1671 gnd.n1398 gnd.n1396 585
R1672 gnd.n4901 gnd.n1396 585
R1673 gnd.n1471 gnd.n1470 585
R1674 gnd.n1470 gnd.n1443 585
R1675 gnd.n1472 gnd.n1450 585
R1676 gnd.n4888 gnd.n1450 585
R1677 gnd.n4875 gnd.n4874 585
R1678 gnd.n4874 gnd.n4873 585
R1679 gnd.n4876 gnd.n1462 585
R1680 gnd.n1462 gnd.n1460 585
R1681 gnd.n4878 gnd.n4877 585
R1682 gnd.n4879 gnd.n4878 585
R1683 gnd.n1463 gnd.n1461 585
R1684 gnd.n4861 gnd.n1461 585
R1685 gnd.n4833 gnd.n4832 585
R1686 gnd.n4832 gnd.n1478 585
R1687 gnd.n4834 gnd.n1486 585
R1688 gnd.n4848 gnd.n1486 585
R1689 gnd.n4835 gnd.n1496 585
R1690 gnd.n1496 gnd.n1484 585
R1691 gnd.n4837 gnd.n4836 585
R1692 gnd.n4838 gnd.n4837 585
R1693 gnd.n1497 gnd.n1495 585
R1694 gnd.n1504 gnd.n1495 585
R1695 gnd.n4824 gnd.n4823 585
R1696 gnd.n4823 gnd.n4822 585
R1697 gnd.n1500 gnd.n1499 585
R1698 gnd.n1501 gnd.n1500 585
R1699 gnd.n4813 gnd.n4812 585
R1700 gnd.n4814 gnd.n4813 585
R1701 gnd.n1514 gnd.n1513 585
R1702 gnd.n1513 gnd.n1510 585
R1703 gnd.n4808 gnd.n4807 585
R1704 gnd.n4807 gnd.n4806 585
R1705 gnd.n1517 gnd.n1516 585
R1706 gnd.n1518 gnd.n1517 585
R1707 gnd.n4797 gnd.n4796 585
R1708 gnd.n4798 gnd.n4797 585
R1709 gnd.n1529 gnd.n1528 585
R1710 gnd.n1536 gnd.n1528 585
R1711 gnd.n4792 gnd.n4791 585
R1712 gnd.n4791 gnd.n4790 585
R1713 gnd.n1532 gnd.n1531 585
R1714 gnd.n1533 gnd.n1532 585
R1715 gnd.n4781 gnd.n4780 585
R1716 gnd.n4782 gnd.n4781 585
R1717 gnd.n1546 gnd.n1545 585
R1718 gnd.n1545 gnd.n1542 585
R1719 gnd.n4776 gnd.n4775 585
R1720 gnd.n4775 gnd.n4774 585
R1721 gnd.n1549 gnd.n1548 585
R1722 gnd.n1550 gnd.n1549 585
R1723 gnd.n4765 gnd.n4764 585
R1724 gnd.n4766 gnd.n4765 585
R1725 gnd.n1561 gnd.n1560 585
R1726 gnd.n4566 gnd.n1560 585
R1727 gnd.n4760 gnd.n4759 585
R1728 gnd.n4759 gnd.n4758 585
R1729 gnd.n4467 gnd.n1563 585
R1730 gnd.n4470 gnd.n4468 585
R1731 gnd.n4473 gnd.n4472 585
R1732 gnd.n4465 gnd.n4464 585
R1733 gnd.n4478 gnd.n4477 585
R1734 gnd.n4480 gnd.n4463 585
R1735 gnd.n4483 gnd.n4482 585
R1736 gnd.n4461 gnd.n4460 585
R1737 gnd.n4488 gnd.n4487 585
R1738 gnd.n4490 gnd.n4459 585
R1739 gnd.n4493 gnd.n4492 585
R1740 gnd.n4457 gnd.n4456 585
R1741 gnd.n4498 gnd.n4497 585
R1742 gnd.n4500 gnd.n4455 585
R1743 gnd.n4503 gnd.n4502 585
R1744 gnd.n4453 gnd.n4452 585
R1745 gnd.n4508 gnd.n4507 585
R1746 gnd.n4510 gnd.n4451 585
R1747 gnd.n4512 gnd.n4511 585
R1748 gnd.n4511 gnd.n4444 585
R1749 gnd.n5744 gnd.n5743 585
R1750 gnd.n1171 gnd.n1163 585
R1751 gnd.n5751 gnd.n1160 585
R1752 gnd.n5752 gnd.n1159 585
R1753 gnd.n1193 gnd.n1153 585
R1754 gnd.n5759 gnd.n1152 585
R1755 gnd.n5760 gnd.n1151 585
R1756 gnd.n1191 gnd.n1143 585
R1757 gnd.n5767 gnd.n1142 585
R1758 gnd.n5768 gnd.n1141 585
R1759 gnd.n1188 gnd.n1135 585
R1760 gnd.n5775 gnd.n1134 585
R1761 gnd.n5776 gnd.n1133 585
R1762 gnd.n1186 gnd.n1126 585
R1763 gnd.n5783 gnd.n1125 585
R1764 gnd.n5784 gnd.n1124 585
R1765 gnd.n5352 gnd.n1123 585
R1766 gnd.n5355 gnd.n5354 585
R1767 gnd.n5351 gnd.n5350 585
R1768 gnd.n5351 gnd.n1196 585
R1769 gnd.n5742 gnd.n1174 585
R1770 gnd.n5742 gnd.n5741 585
R1771 gnd.n5154 gnd.n1173 585
R1772 gnd.n5664 gnd.n1173 585
R1773 gnd.n5155 gnd.n5153 585
R1774 gnd.n5153 gnd.n5152 585
R1775 gnd.n5120 gnd.n1273 585
R1776 gnd.n5344 gnd.n1273 585
R1777 gnd.n5159 gnd.n5119 585
R1778 gnd.n5119 gnd.n5118 585
R1779 gnd.n5160 gnd.n1283 585
R1780 gnd.n5334 gnd.n1283 585
R1781 gnd.n5161 gnd.n4938 585
R1782 gnd.n5107 gnd.n4938 585
R1783 gnd.n4936 gnd.n1292 585
R1784 gnd.n5326 gnd.n1292 585
R1785 gnd.n5165 gnd.n4935 585
R1786 gnd.n5103 gnd.n4935 585
R1787 gnd.n5166 gnd.n1300 585
R1788 gnd.n5318 gnd.n1300 585
R1789 gnd.n5167 gnd.n4934 585
R1790 gnd.n5097 gnd.n4934 585
R1791 gnd.n4932 gnd.n1309 585
R1792 gnd.n5310 gnd.n1309 585
R1793 gnd.n5171 gnd.n4931 585
R1794 gnd.n5019 gnd.n4931 585
R1795 gnd.n5172 gnd.n1318 585
R1796 gnd.n5302 gnd.n1318 585
R1797 gnd.n5173 gnd.n4930 585
R1798 gnd.n5023 gnd.n4930 585
R1799 gnd.n4928 gnd.n1327 585
R1800 gnd.n5294 gnd.n1327 585
R1801 gnd.n5177 gnd.n4927 585
R1802 gnd.n5027 gnd.n4927 585
R1803 gnd.n5178 gnd.n1335 585
R1804 gnd.n5286 gnd.n1335 585
R1805 gnd.n5179 gnd.n4926 585
R1806 gnd.n5033 gnd.n4926 585
R1807 gnd.n4924 gnd.n1344 585
R1808 gnd.n5278 gnd.n1344 585
R1809 gnd.n5183 gnd.n4923 585
R1810 gnd.n5007 gnd.n4923 585
R1811 gnd.n5184 gnd.n1353 585
R1812 gnd.n5270 gnd.n1353 585
R1813 gnd.n5185 gnd.n4922 585
R1814 gnd.n5003 gnd.n4922 585
R1815 gnd.n4920 gnd.n1362 585
R1816 gnd.n5262 gnd.n1362 585
R1817 gnd.n5189 gnd.n4919 585
R1818 gnd.n4997 gnd.n4919 585
R1819 gnd.n5190 gnd.n1370 585
R1820 gnd.n5254 gnd.n1370 585
R1821 gnd.n5191 gnd.n4918 585
R1822 gnd.n4993 gnd.n4918 585
R1823 gnd.n1436 gnd.n1379 585
R1824 gnd.n5246 gnd.n1379 585
R1825 gnd.n5196 gnd.n5195 585
R1826 gnd.n5197 gnd.n5196 585
R1827 gnd.n1435 gnd.n1424 585
R1828 gnd.n5219 gnd.n1424 585
R1829 gnd.n4914 gnd.n4913 585
R1830 gnd.n4913 gnd.n1422 585
R1831 gnd.n4912 gnd.n4911 585
R1832 gnd.n4912 gnd.n1412 585
R1833 gnd.n4910 gnd.n1411 585
R1834 gnd.n5227 gnd.n1411 585
R1835 gnd.n1438 gnd.n1405 585
R1836 gnd.n5232 gnd.n1405 585
R1837 gnd.n4906 gnd.n4905 585
R1838 gnd.n4905 gnd.n1395 585
R1839 gnd.n4904 gnd.n1394 585
R1840 gnd.n5238 gnd.n1394 585
R1841 gnd.n4903 gnd.n4902 585
R1842 gnd.n4902 gnd.n4901 585
R1843 gnd.n1442 gnd.n1440 585
R1844 gnd.n1443 gnd.n1442 585
R1845 gnd.n4870 gnd.n1449 585
R1846 gnd.n4888 gnd.n1449 585
R1847 gnd.n4872 gnd.n4871 585
R1848 gnd.n4873 gnd.n4872 585
R1849 gnd.n1474 gnd.n1473 585
R1850 gnd.n1473 gnd.n1460 585
R1851 gnd.n4864 gnd.n1459 585
R1852 gnd.n4879 gnd.n1459 585
R1853 gnd.n4863 gnd.n4862 585
R1854 gnd.n4862 gnd.n4861 585
R1855 gnd.n1477 gnd.n1476 585
R1856 gnd.n1478 gnd.n1477 585
R1857 gnd.n4536 gnd.n1485 585
R1858 gnd.n4848 gnd.n1485 585
R1859 gnd.n4538 gnd.n4537 585
R1860 gnd.n4537 gnd.n1484 585
R1861 gnd.n4539 gnd.n1494 585
R1862 gnd.n4838 gnd.n1494 585
R1863 gnd.n4541 gnd.n4540 585
R1864 gnd.n4540 gnd.n1504 585
R1865 gnd.n4542 gnd.n1503 585
R1866 gnd.n4822 gnd.n1503 585
R1867 gnd.n4544 gnd.n4543 585
R1868 gnd.n4543 gnd.n1501 585
R1869 gnd.n4545 gnd.n1512 585
R1870 gnd.n4814 gnd.n1512 585
R1871 gnd.n4547 gnd.n4546 585
R1872 gnd.n4546 gnd.n1510 585
R1873 gnd.n4548 gnd.n1520 585
R1874 gnd.n4806 gnd.n1520 585
R1875 gnd.n4550 gnd.n4549 585
R1876 gnd.n4549 gnd.n1518 585
R1877 gnd.n4551 gnd.n1527 585
R1878 gnd.n4798 gnd.n1527 585
R1879 gnd.n4553 gnd.n4552 585
R1880 gnd.n4552 gnd.n1536 585
R1881 gnd.n4554 gnd.n1535 585
R1882 gnd.n4790 gnd.n1535 585
R1883 gnd.n4556 gnd.n4555 585
R1884 gnd.n4555 gnd.n1533 585
R1885 gnd.n4557 gnd.n1544 585
R1886 gnd.n4782 gnd.n1544 585
R1887 gnd.n4559 gnd.n4558 585
R1888 gnd.n4558 gnd.n1542 585
R1889 gnd.n4560 gnd.n1552 585
R1890 gnd.n4774 gnd.n1552 585
R1891 gnd.n4562 gnd.n4561 585
R1892 gnd.n4561 gnd.n1550 585
R1893 gnd.n4563 gnd.n1559 585
R1894 gnd.n4766 gnd.n1559 585
R1895 gnd.n4565 gnd.n4564 585
R1896 gnd.n4566 gnd.n4565 585
R1897 gnd.n4447 gnd.n4446 585
R1898 gnd.n4758 gnd.n4446 585
R1899 gnd.n7741 gnd.n129 585
R1900 gnd.n7837 gnd.n129 585
R1901 gnd.n7742 gnd.n7679 585
R1902 gnd.n7679 gnd.n126 585
R1903 gnd.n7743 gnd.n207 585
R1904 gnd.n7757 gnd.n207 585
R1905 gnd.n219 gnd.n217 585
R1906 gnd.n217 gnd.n206 585
R1907 gnd.n7748 gnd.n7747 585
R1908 gnd.n7749 gnd.n7748 585
R1909 gnd.n218 gnd.n216 585
R1910 gnd.n216 gnd.n213 585
R1911 gnd.n7675 gnd.n7674 585
R1912 gnd.n7674 gnd.n7673 585
R1913 gnd.n222 gnd.n221 585
R1914 gnd.n7492 gnd.n222 585
R1915 gnd.n7664 gnd.n7663 585
R1916 gnd.n7665 gnd.n7664 585
R1917 gnd.n234 gnd.n233 585
R1918 gnd.n233 gnd.n229 585
R1919 gnd.n7659 gnd.n7658 585
R1920 gnd.n7658 gnd.n7657 585
R1921 gnd.n237 gnd.n236 585
R1922 gnd.n238 gnd.n237 585
R1923 gnd.n7648 gnd.n7647 585
R1924 gnd.n7649 gnd.n7648 585
R1925 gnd.n248 gnd.n247 585
R1926 gnd.n253 gnd.n247 585
R1927 gnd.n7643 gnd.n7642 585
R1928 gnd.n7642 gnd.n7641 585
R1929 gnd.n251 gnd.n250 585
R1930 gnd.n262 gnd.n251 585
R1931 gnd.n7632 gnd.n7631 585
R1932 gnd.n7633 gnd.n7632 585
R1933 gnd.n264 gnd.n263 585
R1934 gnd.n263 gnd.n259 585
R1935 gnd.n7627 gnd.n7626 585
R1936 gnd.n7626 gnd.n7625 585
R1937 gnd.n267 gnd.n266 585
R1938 gnd.n268 gnd.n267 585
R1939 gnd.n7616 gnd.n7615 585
R1940 gnd.n7617 gnd.n7616 585
R1941 gnd.n278 gnd.n277 585
R1942 gnd.n283 gnd.n277 585
R1943 gnd.n7611 gnd.n7610 585
R1944 gnd.n7610 gnd.n7609 585
R1945 gnd.n281 gnd.n280 585
R1946 gnd.n292 gnd.n281 585
R1947 gnd.n7600 gnd.n7599 585
R1948 gnd.n7601 gnd.n7600 585
R1949 gnd.n294 gnd.n293 585
R1950 gnd.n293 gnd.n289 585
R1951 gnd.n7595 gnd.n7594 585
R1952 gnd.n7594 gnd.n7593 585
R1953 gnd.n297 gnd.n296 585
R1954 gnd.n298 gnd.n297 585
R1955 gnd.n7571 gnd.n7570 585
R1956 gnd.n7570 gnd.n7569 585
R1957 gnd.n7572 gnd.n326 585
R1958 gnd.n7565 gnd.n326 585
R1959 gnd.n332 gnd.n324 585
R1960 gnd.n333 gnd.n332 585
R1961 gnd.n7576 gnd.n323 585
R1962 gnd.n7555 gnd.n323 585
R1963 gnd.n7577 gnd.n322 585
R1964 gnd.n343 gnd.n322 585
R1965 gnd.n7578 gnd.n321 585
R1966 gnd.n7549 gnd.n321 585
R1967 gnd.n318 gnd.n316 585
R1968 gnd.n7533 gnd.n316 585
R1969 gnd.n7583 gnd.n7582 585
R1970 gnd.n7584 gnd.n7583 585
R1971 gnd.n317 gnd.n315 585
R1972 gnd.n7539 gnd.n315 585
R1973 gnd.n7430 gnd.n7428 585
R1974 gnd.n7428 gnd.n7427 585
R1975 gnd.n7431 gnd.n365 585
R1976 gnd.n7447 gnd.n365 585
R1977 gnd.n7432 gnd.n7426 585
R1978 gnd.n7426 gnd.n7425 585
R1979 gnd.n380 gnd.n378 585
R1980 gnd.n7409 gnd.n378 585
R1981 gnd.n7437 gnd.n7436 585
R1982 gnd.n7438 gnd.n7437 585
R1983 gnd.n379 gnd.n377 585
R1984 gnd.n7415 gnd.n377 585
R1985 gnd.n7384 gnd.n7383 585
R1986 gnd.n7383 gnd.n7382 585
R1987 gnd.n7385 gnd.n398 585
R1988 gnd.n7401 gnd.n398 585
R1989 gnd.n412 gnd.n410 585
R1990 gnd.n7332 gnd.n410 585
R1991 gnd.n7390 gnd.n7389 585
R1992 gnd.n7391 gnd.n7390 585
R1993 gnd.n411 gnd.n409 585
R1994 gnd.n7341 gnd.n409 585
R1995 gnd.n7308 gnd.n7307 585
R1996 gnd.n7307 gnd.n422 585
R1997 gnd.n7309 gnd.n433 585
R1998 gnd.n7325 gnd.n433 585
R1999 gnd.n447 gnd.n445 585
R2000 gnd.n7145 gnd.n445 585
R2001 gnd.n7314 gnd.n7313 585
R2002 gnd.n7315 gnd.n7314 585
R2003 gnd.n446 gnd.n444 585
R2004 gnd.n7151 gnd.n444 585
R2005 gnd.n7303 gnd.n7302 585
R2006 gnd.n7302 gnd.n7301 585
R2007 gnd.n450 gnd.n449 585
R2008 gnd.n7128 gnd.n450 585
R2009 gnd.n7292 gnd.n7291 585
R2010 gnd.n7293 gnd.n7292 585
R2011 gnd.n464 gnd.n463 585
R2012 gnd.n617 gnd.n463 585
R2013 gnd.n7287 gnd.n7286 585
R2014 gnd.n7286 gnd.n7285 585
R2015 gnd.n467 gnd.n466 585
R2016 gnd.n611 gnd.n467 585
R2017 gnd.n7276 gnd.n7275 585
R2018 gnd.n7277 gnd.n7276 585
R2019 gnd.n482 gnd.n481 585
R2020 gnd.n607 gnd.n481 585
R2021 gnd.n7271 gnd.n7270 585
R2022 gnd.n7270 gnd.n7269 585
R2023 gnd.n485 gnd.n484 585
R2024 gnd.n601 gnd.n485 585
R2025 gnd.n7260 gnd.n7259 585
R2026 gnd.n7261 gnd.n7260 585
R2027 gnd.n500 gnd.n499 585
R2028 gnd.n7176 gnd.n499 585
R2029 gnd.n7255 gnd.n7254 585
R2030 gnd.n503 gnd.n502 585
R2031 gnd.n6728 gnd.n6599 585
R2032 gnd.n6727 gnd.n6600 585
R2033 gnd.n6602 gnd.n6601 585
R2034 gnd.n6720 gnd.n6610 585
R2035 gnd.n6719 gnd.n6611 585
R2036 gnd.n6618 gnd.n6612 585
R2037 gnd.n6712 gnd.n6619 585
R2038 gnd.n6711 gnd.n6620 585
R2039 gnd.n6622 gnd.n6621 585
R2040 gnd.n6704 gnd.n6630 585
R2041 gnd.n6703 gnd.n6631 585
R2042 gnd.n6638 gnd.n6632 585
R2043 gnd.n6696 gnd.n6639 585
R2044 gnd.n6695 gnd.n6640 585
R2045 gnd.n6642 gnd.n6641 585
R2046 gnd.n6688 gnd.n6685 585
R2047 gnd.n6684 gnd.n531 585
R2048 gnd.n7252 gnd.n531 585
R2049 gnd.n7840 gnd.n7839 585
R2050 gnd.n7712 gnd.n124 585
R2051 gnd.n7714 gnd.n7713 585
R2052 gnd.n7710 gnd.n7709 585
R2053 gnd.n7718 gnd.n7708 585
R2054 gnd.n7719 gnd.n7706 585
R2055 gnd.n7720 gnd.n7705 585
R2056 gnd.n7703 gnd.n7701 585
R2057 gnd.n7724 gnd.n7700 585
R2058 gnd.n7725 gnd.n7698 585
R2059 gnd.n7726 gnd.n7697 585
R2060 gnd.n7695 gnd.n7693 585
R2061 gnd.n7730 gnd.n7692 585
R2062 gnd.n7731 gnd.n7690 585
R2063 gnd.n7732 gnd.n7689 585
R2064 gnd.n7687 gnd.n7685 585
R2065 gnd.n7736 gnd.n7684 585
R2066 gnd.n7737 gnd.n7682 585
R2067 gnd.n7738 gnd.n7681 585
R2068 gnd.n7681 gnd.n128 585
R2069 gnd.n7838 gnd.n120 585
R2070 gnd.n7838 gnd.n7837 585
R2071 gnd.n7844 gnd.n119 585
R2072 gnd.n126 gnd.n119 585
R2073 gnd.n7845 gnd.n118 585
R2074 gnd.n7757 gnd.n118 585
R2075 gnd.n7846 gnd.n117 585
R2076 gnd.n206 gnd.n117 585
R2077 gnd.n215 gnd.n115 585
R2078 gnd.n7749 gnd.n215 585
R2079 gnd.n7850 gnd.n114 585
R2080 gnd.n213 gnd.n114 585
R2081 gnd.n7851 gnd.n113 585
R2082 gnd.n7673 gnd.n113 585
R2083 gnd.n7852 gnd.n112 585
R2084 gnd.n7492 gnd.n112 585
R2085 gnd.n231 gnd.n110 585
R2086 gnd.n7665 gnd.n231 585
R2087 gnd.n7856 gnd.n109 585
R2088 gnd.n229 gnd.n109 585
R2089 gnd.n7857 gnd.n108 585
R2090 gnd.n7657 gnd.n108 585
R2091 gnd.n7858 gnd.n107 585
R2092 gnd.n238 gnd.n107 585
R2093 gnd.n246 gnd.n105 585
R2094 gnd.n7649 gnd.n246 585
R2095 gnd.n7862 gnd.n104 585
R2096 gnd.n253 gnd.n104 585
R2097 gnd.n7863 gnd.n103 585
R2098 gnd.n7641 gnd.n103 585
R2099 gnd.n7864 gnd.n102 585
R2100 gnd.n262 gnd.n102 585
R2101 gnd.n261 gnd.n100 585
R2102 gnd.n7633 gnd.n261 585
R2103 gnd.n7868 gnd.n99 585
R2104 gnd.n259 gnd.n99 585
R2105 gnd.n7869 gnd.n98 585
R2106 gnd.n7625 gnd.n98 585
R2107 gnd.n7870 gnd.n97 585
R2108 gnd.n268 gnd.n97 585
R2109 gnd.n276 gnd.n95 585
R2110 gnd.n7617 gnd.n276 585
R2111 gnd.n7874 gnd.n94 585
R2112 gnd.n283 gnd.n94 585
R2113 gnd.n7875 gnd.n93 585
R2114 gnd.n7609 gnd.n93 585
R2115 gnd.n7876 gnd.n92 585
R2116 gnd.n292 gnd.n92 585
R2117 gnd.n291 gnd.n90 585
R2118 gnd.n7601 gnd.n291 585
R2119 gnd.n7880 gnd.n89 585
R2120 gnd.n289 gnd.n89 585
R2121 gnd.n7881 gnd.n88 585
R2122 gnd.n7593 gnd.n88 585
R2123 gnd.n7882 gnd.n87 585
R2124 gnd.n298 gnd.n87 585
R2125 gnd.n328 gnd.n85 585
R2126 gnd.n7569 gnd.n328 585
R2127 gnd.n7886 gnd.n84 585
R2128 gnd.n7565 gnd.n84 585
R2129 gnd.n7887 gnd.n83 585
R2130 gnd.n333 gnd.n83 585
R2131 gnd.n7888 gnd.n82 585
R2132 gnd.n7555 gnd.n82 585
R2133 gnd.n351 gnd.n80 585
R2134 gnd.n351 gnd.n343 585
R2135 gnd.n7547 gnd.n7546 585
R2136 gnd.n7549 gnd.n7547 585
R2137 gnd.n7545 gnd.n350 585
R2138 gnd.n7533 gnd.n350 585
R2139 gnd.n352 gnd.n313 585
R2140 gnd.n7584 gnd.n313 585
R2141 gnd.n7541 gnd.n7540 585
R2142 gnd.n7540 gnd.n7539 585
R2143 gnd.n355 gnd.n354 585
R2144 gnd.n7427 gnd.n355 585
R2145 gnd.n386 gnd.n363 585
R2146 gnd.n7447 gnd.n363 585
R2147 gnd.n7424 gnd.n7423 585
R2148 gnd.n7425 gnd.n7424 585
R2149 gnd.n385 gnd.n384 585
R2150 gnd.n7409 gnd.n384 585
R2151 gnd.n7418 gnd.n375 585
R2152 gnd.n7438 gnd.n375 585
R2153 gnd.n7417 gnd.n7416 585
R2154 gnd.n7416 gnd.n7415 585
R2155 gnd.n389 gnd.n388 585
R2156 gnd.n7382 gnd.n389 585
R2157 gnd.n7334 gnd.n397 585
R2158 gnd.n7401 gnd.n397 585
R2159 gnd.n7335 gnd.n7333 585
R2160 gnd.n7333 gnd.n7332 585
R2161 gnd.n426 gnd.n407 585
R2162 gnd.n7391 gnd.n407 585
R2163 gnd.n7340 gnd.n7339 585
R2164 gnd.n7341 gnd.n7340 585
R2165 gnd.n425 gnd.n424 585
R2166 gnd.n424 gnd.n422 585
R2167 gnd.n7327 gnd.n7326 585
R2168 gnd.n7326 gnd.n7325 585
R2169 gnd.n429 gnd.n428 585
R2170 gnd.n7145 gnd.n429 585
R2171 gnd.n7153 gnd.n442 585
R2172 gnd.n7315 gnd.n442 585
R2173 gnd.n7156 gnd.n7152 585
R2174 gnd.n7152 gnd.n7151 585
R2175 gnd.n7157 gnd.n453 585
R2176 gnd.n7301 gnd.n453 585
R2177 gnd.n7158 gnd.n593 585
R2178 gnd.n7128 gnd.n593 585
R2179 gnd.n591 gnd.n462 585
R2180 gnd.n7293 gnd.n462 585
R2181 gnd.n7162 gnd.n590 585
R2182 gnd.n617 gnd.n590 585
R2183 gnd.n7163 gnd.n470 585
R2184 gnd.n7285 gnd.n470 585
R2185 gnd.n7164 gnd.n589 585
R2186 gnd.n611 gnd.n589 585
R2187 gnd.n587 gnd.n479 585
R2188 gnd.n7277 gnd.n479 585
R2189 gnd.n7168 gnd.n586 585
R2190 gnd.n607 gnd.n586 585
R2191 gnd.n7169 gnd.n488 585
R2192 gnd.n7269 gnd.n488 585
R2193 gnd.n7170 gnd.n585 585
R2194 gnd.n601 gnd.n585 585
R2195 gnd.n582 gnd.n497 585
R2196 gnd.n7261 gnd.n497 585
R2197 gnd.n7175 gnd.n7174 585
R2198 gnd.n7176 gnd.n7175 585
R2199 gnd.n4351 gnd.n4350 585
R2200 gnd.n4352 gnd.n4351 585
R2201 gnd.n1640 gnd.n1639 585
R2202 gnd.n1646 gnd.n1639 585
R2203 gnd.n4326 gnd.n3064 585
R2204 gnd.n3064 gnd.n1645 585
R2205 gnd.n4328 gnd.n4327 585
R2206 gnd.n4329 gnd.n4328 585
R2207 gnd.n3065 gnd.n3063 585
R2208 gnd.n3063 gnd.n1653 585
R2209 gnd.n4060 gnd.n4059 585
R2210 gnd.n4059 gnd.n4058 585
R2211 gnd.n3070 gnd.n3069 585
R2212 gnd.n4029 gnd.n3070 585
R2213 gnd.n4049 gnd.n4048 585
R2214 gnd.n4048 gnd.n4047 585
R2215 gnd.n3077 gnd.n3076 585
R2216 gnd.n4035 gnd.n3077 585
R2217 gnd.n4005 gnd.n3097 585
R2218 gnd.n3097 gnd.n3096 585
R2219 gnd.n4007 gnd.n4006 585
R2220 gnd.n4008 gnd.n4007 585
R2221 gnd.n3098 gnd.n3095 585
R2222 gnd.n3106 gnd.n3095 585
R2223 gnd.n3983 gnd.n3118 585
R2224 gnd.n3118 gnd.n3105 585
R2225 gnd.n3985 gnd.n3984 585
R2226 gnd.n3986 gnd.n3985 585
R2227 gnd.n3119 gnd.n3117 585
R2228 gnd.n3117 gnd.n3113 585
R2229 gnd.n3971 gnd.n3970 585
R2230 gnd.n3970 gnd.n3969 585
R2231 gnd.n3124 gnd.n3123 585
R2232 gnd.n3134 gnd.n3124 585
R2233 gnd.n3960 gnd.n3959 585
R2234 gnd.n3959 gnd.n3958 585
R2235 gnd.n3131 gnd.n3130 585
R2236 gnd.n3946 gnd.n3131 585
R2237 gnd.n3920 gnd.n3152 585
R2238 gnd.n3152 gnd.n3141 585
R2239 gnd.n3922 gnd.n3921 585
R2240 gnd.n3923 gnd.n3922 585
R2241 gnd.n3153 gnd.n3151 585
R2242 gnd.n3161 gnd.n3151 585
R2243 gnd.n3898 gnd.n3173 585
R2244 gnd.n3173 gnd.n3160 585
R2245 gnd.n3900 gnd.n3899 585
R2246 gnd.n3901 gnd.n3900 585
R2247 gnd.n3174 gnd.n3172 585
R2248 gnd.n3172 gnd.n3168 585
R2249 gnd.n3886 gnd.n3885 585
R2250 gnd.n3885 gnd.n3884 585
R2251 gnd.n3179 gnd.n3178 585
R2252 gnd.n3188 gnd.n3179 585
R2253 gnd.n3875 gnd.n3874 585
R2254 gnd.n3874 gnd.n3873 585
R2255 gnd.n3186 gnd.n3185 585
R2256 gnd.n3861 gnd.n3186 585
R2257 gnd.n3299 gnd.n3298 585
R2258 gnd.n3299 gnd.n3195 585
R2259 gnd.n3818 gnd.n3817 585
R2260 gnd.n3817 gnd.n3816 585
R2261 gnd.n3819 gnd.n3293 585
R2262 gnd.n3304 gnd.n3293 585
R2263 gnd.n3821 gnd.n3820 585
R2264 gnd.n3822 gnd.n3821 585
R2265 gnd.n3294 gnd.n3292 585
R2266 gnd.n3317 gnd.n3292 585
R2267 gnd.n3277 gnd.n3276 585
R2268 gnd.n3280 gnd.n3277 585
R2269 gnd.n3832 gnd.n3831 585
R2270 gnd.n3831 gnd.n3830 585
R2271 gnd.n3833 gnd.n3271 585
R2272 gnd.n3792 gnd.n3271 585
R2273 gnd.n3835 gnd.n3834 585
R2274 gnd.n3836 gnd.n3835 585
R2275 gnd.n3272 gnd.n3270 585
R2276 gnd.n3331 gnd.n3270 585
R2277 gnd.n3784 gnd.n3783 585
R2278 gnd.n3783 gnd.n3782 585
R2279 gnd.n3328 gnd.n3327 585
R2280 gnd.n3766 gnd.n3328 585
R2281 gnd.n3753 gnd.n3347 585
R2282 gnd.n3347 gnd.n3346 585
R2283 gnd.n3755 gnd.n3754 585
R2284 gnd.n3756 gnd.n3755 585
R2285 gnd.n3348 gnd.n3345 585
R2286 gnd.n3354 gnd.n3345 585
R2287 gnd.n3734 gnd.n3733 585
R2288 gnd.n3735 gnd.n3734 585
R2289 gnd.n3365 gnd.n3364 585
R2290 gnd.n3364 gnd.n3360 585
R2291 gnd.n3724 gnd.n3723 585
R2292 gnd.n3725 gnd.n3724 585
R2293 gnd.n3375 gnd.n3374 585
R2294 gnd.n3380 gnd.n3374 585
R2295 gnd.n3702 gnd.n3393 585
R2296 gnd.n3393 gnd.n3379 585
R2297 gnd.n3704 gnd.n3703 585
R2298 gnd.n3705 gnd.n3704 585
R2299 gnd.n3394 gnd.n3392 585
R2300 gnd.n3392 gnd.n3388 585
R2301 gnd.n3693 gnd.n3692 585
R2302 gnd.n3694 gnd.n3693 585
R2303 gnd.n3401 gnd.n3400 585
R2304 gnd.n3405 gnd.n3400 585
R2305 gnd.n3670 gnd.n3422 585
R2306 gnd.n3422 gnd.n3404 585
R2307 gnd.n3672 gnd.n3671 585
R2308 gnd.n3673 gnd.n3672 585
R2309 gnd.n3423 gnd.n3421 585
R2310 gnd.n3421 gnd.n3412 585
R2311 gnd.n3665 gnd.n3664 585
R2312 gnd.n3664 gnd.n3663 585
R2313 gnd.n3470 gnd.n3469 585
R2314 gnd.n3471 gnd.n3470 585
R2315 gnd.n3624 gnd.n3623 585
R2316 gnd.n3625 gnd.n3624 585
R2317 gnd.n3480 gnd.n3479 585
R2318 gnd.n3479 gnd.n3478 585
R2319 gnd.n3619 gnd.n3618 585
R2320 gnd.n3618 gnd.n3617 585
R2321 gnd.n3483 gnd.n3482 585
R2322 gnd.n3484 gnd.n3483 585
R2323 gnd.n3608 gnd.n3607 585
R2324 gnd.n3609 gnd.n3608 585
R2325 gnd.n3491 gnd.n3490 585
R2326 gnd.n3600 gnd.n3490 585
R2327 gnd.n3603 gnd.n3602 585
R2328 gnd.n3602 gnd.n3601 585
R2329 gnd.n3494 gnd.n3493 585
R2330 gnd.n3495 gnd.n3494 585
R2331 gnd.n3589 gnd.n3588 585
R2332 gnd.n3587 gnd.n3513 585
R2333 gnd.n3586 gnd.n3512 585
R2334 gnd.n3591 gnd.n3512 585
R2335 gnd.n3585 gnd.n3584 585
R2336 gnd.n3583 gnd.n3582 585
R2337 gnd.n3581 gnd.n3580 585
R2338 gnd.n3579 gnd.n3578 585
R2339 gnd.n3577 gnd.n3576 585
R2340 gnd.n3575 gnd.n3574 585
R2341 gnd.n3573 gnd.n3572 585
R2342 gnd.n3571 gnd.n3570 585
R2343 gnd.n3569 gnd.n3568 585
R2344 gnd.n3567 gnd.n3566 585
R2345 gnd.n3565 gnd.n3564 585
R2346 gnd.n3563 gnd.n3562 585
R2347 gnd.n3561 gnd.n3560 585
R2348 gnd.n3559 gnd.n3558 585
R2349 gnd.n3557 gnd.n3556 585
R2350 gnd.n3555 gnd.n3554 585
R2351 gnd.n3553 gnd.n3552 585
R2352 gnd.n3551 gnd.n3550 585
R2353 gnd.n3549 gnd.n3548 585
R2354 gnd.n3547 gnd.n3546 585
R2355 gnd.n3545 gnd.n3544 585
R2356 gnd.n3543 gnd.n3542 585
R2357 gnd.n3500 gnd.n3499 585
R2358 gnd.n3594 gnd.n3593 585
R2359 gnd.n4355 gnd.n4354 585
R2360 gnd.n4357 gnd.n4356 585
R2361 gnd.n4359 gnd.n4358 585
R2362 gnd.n4361 gnd.n4360 585
R2363 gnd.n4363 gnd.n4362 585
R2364 gnd.n4365 gnd.n4364 585
R2365 gnd.n4367 gnd.n4366 585
R2366 gnd.n4369 gnd.n4368 585
R2367 gnd.n4371 gnd.n4370 585
R2368 gnd.n4373 gnd.n4372 585
R2369 gnd.n4375 gnd.n4374 585
R2370 gnd.n4377 gnd.n4376 585
R2371 gnd.n4379 gnd.n4378 585
R2372 gnd.n4381 gnd.n4380 585
R2373 gnd.n4383 gnd.n4382 585
R2374 gnd.n4385 gnd.n4384 585
R2375 gnd.n4387 gnd.n4386 585
R2376 gnd.n4389 gnd.n4388 585
R2377 gnd.n4391 gnd.n4390 585
R2378 gnd.n4393 gnd.n4392 585
R2379 gnd.n4395 gnd.n4394 585
R2380 gnd.n4397 gnd.n4396 585
R2381 gnd.n4399 gnd.n4398 585
R2382 gnd.n4401 gnd.n4400 585
R2383 gnd.n4403 gnd.n4402 585
R2384 gnd.n4404 gnd.n1607 585
R2385 gnd.n4405 gnd.n1565 585
R2386 gnd.n4443 gnd.n1565 585
R2387 gnd.n4353 gnd.n1637 585
R2388 gnd.n4353 gnd.n4352 585
R2389 gnd.n4022 gnd.n1636 585
R2390 gnd.n1646 gnd.n1636 585
R2391 gnd.n4024 gnd.n4023 585
R2392 gnd.n4023 gnd.n1645 585
R2393 gnd.n4025 gnd.n1655 585
R2394 gnd.n4329 gnd.n1655 585
R2395 gnd.n4027 gnd.n4026 585
R2396 gnd.n4026 gnd.n1653 585
R2397 gnd.n4028 gnd.n3072 585
R2398 gnd.n4058 gnd.n3072 585
R2399 gnd.n4031 gnd.n4030 585
R2400 gnd.n4030 gnd.n4029 585
R2401 gnd.n4032 gnd.n3079 585
R2402 gnd.n4047 gnd.n3079 585
R2403 gnd.n4034 gnd.n4033 585
R2404 gnd.n4035 gnd.n4034 585
R2405 gnd.n3089 gnd.n3088 585
R2406 gnd.n3096 gnd.n3088 585
R2407 gnd.n4010 gnd.n4009 585
R2408 gnd.n4009 gnd.n4008 585
R2409 gnd.n3092 gnd.n3091 585
R2410 gnd.n3106 gnd.n3092 585
R2411 gnd.n3936 gnd.n3935 585
R2412 gnd.n3935 gnd.n3105 585
R2413 gnd.n3937 gnd.n3115 585
R2414 gnd.n3986 gnd.n3115 585
R2415 gnd.n3939 gnd.n3938 585
R2416 gnd.n3938 gnd.n3113 585
R2417 gnd.n3940 gnd.n3126 585
R2418 gnd.n3969 gnd.n3126 585
R2419 gnd.n3942 gnd.n3941 585
R2420 gnd.n3941 gnd.n3134 585
R2421 gnd.n3943 gnd.n3133 585
R2422 gnd.n3958 gnd.n3133 585
R2423 gnd.n3945 gnd.n3944 585
R2424 gnd.n3946 gnd.n3945 585
R2425 gnd.n3145 gnd.n3144 585
R2426 gnd.n3144 gnd.n3141 585
R2427 gnd.n3925 gnd.n3924 585
R2428 gnd.n3924 gnd.n3923 585
R2429 gnd.n3148 gnd.n3147 585
R2430 gnd.n3161 gnd.n3148 585
R2431 gnd.n3849 gnd.n3848 585
R2432 gnd.n3848 gnd.n3160 585
R2433 gnd.n3850 gnd.n3170 585
R2434 gnd.n3901 gnd.n3170 585
R2435 gnd.n3852 gnd.n3851 585
R2436 gnd.n3851 gnd.n3168 585
R2437 gnd.n3853 gnd.n3181 585
R2438 gnd.n3884 gnd.n3181 585
R2439 gnd.n3855 gnd.n3854 585
R2440 gnd.n3854 gnd.n3188 585
R2441 gnd.n3856 gnd.n3187 585
R2442 gnd.n3873 gnd.n3187 585
R2443 gnd.n3858 gnd.n3857 585
R2444 gnd.n3861 gnd.n3858 585
R2445 gnd.n3198 gnd.n3197 585
R2446 gnd.n3197 gnd.n3195 585
R2447 gnd.n3301 gnd.n3300 585
R2448 gnd.n3816 gnd.n3300 585
R2449 gnd.n3303 gnd.n3302 585
R2450 gnd.n3304 gnd.n3303 585
R2451 gnd.n3314 gnd.n3290 585
R2452 gnd.n3822 gnd.n3290 585
R2453 gnd.n3316 gnd.n3315 585
R2454 gnd.n3317 gnd.n3316 585
R2455 gnd.n3313 gnd.n3312 585
R2456 gnd.n3313 gnd.n3280 585
R2457 gnd.n3311 gnd.n3278 585
R2458 gnd.n3830 gnd.n3278 585
R2459 gnd.n3267 gnd.n3265 585
R2460 gnd.n3792 gnd.n3267 585
R2461 gnd.n3838 gnd.n3837 585
R2462 gnd.n3837 gnd.n3836 585
R2463 gnd.n3266 gnd.n3264 585
R2464 gnd.n3331 gnd.n3266 585
R2465 gnd.n3763 gnd.n3330 585
R2466 gnd.n3782 gnd.n3330 585
R2467 gnd.n3765 gnd.n3764 585
R2468 gnd.n3766 gnd.n3765 585
R2469 gnd.n3340 gnd.n3339 585
R2470 gnd.n3346 gnd.n3339 585
R2471 gnd.n3758 gnd.n3757 585
R2472 gnd.n3757 gnd.n3756 585
R2473 gnd.n3343 gnd.n3342 585
R2474 gnd.n3354 gnd.n3343 585
R2475 gnd.n3643 gnd.n3362 585
R2476 gnd.n3735 gnd.n3362 585
R2477 gnd.n3645 gnd.n3644 585
R2478 gnd.n3644 gnd.n3360 585
R2479 gnd.n3646 gnd.n3373 585
R2480 gnd.n3725 gnd.n3373 585
R2481 gnd.n3648 gnd.n3647 585
R2482 gnd.n3648 gnd.n3380 585
R2483 gnd.n3650 gnd.n3649 585
R2484 gnd.n3649 gnd.n3379 585
R2485 gnd.n3651 gnd.n3390 585
R2486 gnd.n3705 gnd.n3390 585
R2487 gnd.n3653 gnd.n3652 585
R2488 gnd.n3652 gnd.n3388 585
R2489 gnd.n3654 gnd.n3399 585
R2490 gnd.n3694 gnd.n3399 585
R2491 gnd.n3656 gnd.n3655 585
R2492 gnd.n3656 gnd.n3405 585
R2493 gnd.n3658 gnd.n3657 585
R2494 gnd.n3657 gnd.n3404 585
R2495 gnd.n3659 gnd.n3420 585
R2496 gnd.n3673 gnd.n3420 585
R2497 gnd.n3660 gnd.n3473 585
R2498 gnd.n3473 gnd.n3412 585
R2499 gnd.n3662 gnd.n3661 585
R2500 gnd.n3663 gnd.n3662 585
R2501 gnd.n3474 gnd.n3472 585
R2502 gnd.n3472 gnd.n3471 585
R2503 gnd.n3627 gnd.n3626 585
R2504 gnd.n3626 gnd.n3625 585
R2505 gnd.n3477 gnd.n3476 585
R2506 gnd.n3478 gnd.n3477 585
R2507 gnd.n3616 gnd.n3615 585
R2508 gnd.n3617 gnd.n3616 585
R2509 gnd.n3486 gnd.n3485 585
R2510 gnd.n3485 gnd.n3484 585
R2511 gnd.n3611 gnd.n3610 585
R2512 gnd.n3610 gnd.n3609 585
R2513 gnd.n3489 gnd.n3488 585
R2514 gnd.n3600 gnd.n3489 585
R2515 gnd.n3599 gnd.n3598 585
R2516 gnd.n3601 gnd.n3599 585
R2517 gnd.n3497 gnd.n3496 585
R2518 gnd.n3496 gnd.n3495 585
R2519 gnd.n4338 gnd.n1587 585
R2520 gnd.n1587 gnd.n1564 585
R2521 gnd.n4339 gnd.n1648 585
R2522 gnd.n1648 gnd.n1638 585
R2523 gnd.n4341 gnd.n4340 585
R2524 gnd.n4342 gnd.n4341 585
R2525 gnd.n1649 gnd.n1647 585
R2526 gnd.n3062 gnd.n1647 585
R2527 gnd.n4332 gnd.n4331 585
R2528 gnd.n4331 gnd.n4330 585
R2529 gnd.n1652 gnd.n1651 585
R2530 gnd.n4057 gnd.n1652 585
R2531 gnd.n4043 gnd.n3081 585
R2532 gnd.n3081 gnd.n3071 585
R2533 gnd.n4045 gnd.n4044 585
R2534 gnd.n4046 gnd.n4045 585
R2535 gnd.n3082 gnd.n3080 585
R2536 gnd.n3080 gnd.n3078 585
R2537 gnd.n4038 gnd.n4037 585
R2538 gnd.n4037 gnd.n4036 585
R2539 gnd.n3085 gnd.n3084 585
R2540 gnd.n3094 gnd.n3085 585
R2541 gnd.n3994 gnd.n3108 585
R2542 gnd.n3108 gnd.n3093 585
R2543 gnd.n3996 gnd.n3995 585
R2544 gnd.n3997 gnd.n3996 585
R2545 gnd.n3109 gnd.n3107 585
R2546 gnd.n3116 gnd.n3107 585
R2547 gnd.n3989 gnd.n3988 585
R2548 gnd.n3988 gnd.n3987 585
R2549 gnd.n3112 gnd.n3111 585
R2550 gnd.n3968 gnd.n3112 585
R2551 gnd.n3954 gnd.n3136 585
R2552 gnd.n3136 gnd.n3125 585
R2553 gnd.n3956 gnd.n3955 585
R2554 gnd.n3957 gnd.n3956 585
R2555 gnd.n3137 gnd.n3135 585
R2556 gnd.n3135 gnd.n3132 585
R2557 gnd.n3949 gnd.n3948 585
R2558 gnd.n3948 gnd.n3947 585
R2559 gnd.n3140 gnd.n3139 585
R2560 gnd.n3150 gnd.n3140 585
R2561 gnd.n3909 gnd.n3163 585
R2562 gnd.n3163 gnd.n3149 585
R2563 gnd.n3911 gnd.n3910 585
R2564 gnd.n3912 gnd.n3911 585
R2565 gnd.n3164 gnd.n3162 585
R2566 gnd.n3171 gnd.n3162 585
R2567 gnd.n3904 gnd.n3903 585
R2568 gnd.n3903 gnd.n3902 585
R2569 gnd.n3167 gnd.n3166 585
R2570 gnd.n3883 gnd.n3167 585
R2571 gnd.n3869 gnd.n3190 585
R2572 gnd.n3190 gnd.n3180 585
R2573 gnd.n3871 gnd.n3870 585
R2574 gnd.n3872 gnd.n3871 585
R2575 gnd.n3191 gnd.n3189 585
R2576 gnd.n3860 gnd.n3189 585
R2577 gnd.n3864 gnd.n3863 585
R2578 gnd.n3863 gnd.n3862 585
R2579 gnd.n3194 gnd.n3193 585
R2580 gnd.n3815 gnd.n3194 585
R2581 gnd.n3308 gnd.n3307 585
R2582 gnd.n3309 gnd.n3308 585
R2583 gnd.n3288 gnd.n3287 585
R2584 gnd.n3291 gnd.n3288 585
R2585 gnd.n3825 gnd.n3824 585
R2586 gnd.n3824 gnd.n3823 585
R2587 gnd.n3826 gnd.n3282 585
R2588 gnd.n3318 gnd.n3282 585
R2589 gnd.n3828 gnd.n3827 585
R2590 gnd.n3829 gnd.n3828 585
R2591 gnd.n3283 gnd.n3281 585
R2592 gnd.n3793 gnd.n3281 585
R2593 gnd.n3777 gnd.n3776 585
R2594 gnd.n3776 gnd.n3269 585
R2595 gnd.n3778 gnd.n3333 585
R2596 gnd.n3333 gnd.n3268 585
R2597 gnd.n3780 gnd.n3779 585
R2598 gnd.n3781 gnd.n3780 585
R2599 gnd.n3334 gnd.n3332 585
R2600 gnd.n3332 gnd.n3329 585
R2601 gnd.n3769 gnd.n3768 585
R2602 gnd.n3768 gnd.n3767 585
R2603 gnd.n3337 gnd.n3336 585
R2604 gnd.n3344 gnd.n3337 585
R2605 gnd.n3743 gnd.n3742 585
R2606 gnd.n3744 gnd.n3743 585
R2607 gnd.n3356 gnd.n3355 585
R2608 gnd.n3363 gnd.n3355 585
R2609 gnd.n3738 gnd.n3737 585
R2610 gnd.n3737 gnd.n3736 585
R2611 gnd.n3359 gnd.n3358 585
R2612 gnd.n3726 gnd.n3359 585
R2613 gnd.n3713 gnd.n3383 585
R2614 gnd.n3383 gnd.n3382 585
R2615 gnd.n3715 gnd.n3714 585
R2616 gnd.n3716 gnd.n3715 585
R2617 gnd.n3384 gnd.n3381 585
R2618 gnd.n3391 gnd.n3381 585
R2619 gnd.n3708 gnd.n3707 585
R2620 gnd.n3707 gnd.n3706 585
R2621 gnd.n3387 gnd.n3386 585
R2622 gnd.n3695 gnd.n3387 585
R2623 gnd.n3682 gnd.n3408 585
R2624 gnd.n3408 gnd.n3407 585
R2625 gnd.n3684 gnd.n3683 585
R2626 gnd.n3685 gnd.n3684 585
R2627 gnd.n3678 gnd.n3406 585
R2628 gnd.n3677 gnd.n3676 585
R2629 gnd.n3411 gnd.n3410 585
R2630 gnd.n3674 gnd.n3411 585
R2631 gnd.n3433 gnd.n3432 585
R2632 gnd.n3436 gnd.n3435 585
R2633 gnd.n3434 gnd.n3429 585
R2634 gnd.n3441 gnd.n3440 585
R2635 gnd.n3443 gnd.n3442 585
R2636 gnd.n3446 gnd.n3445 585
R2637 gnd.n3444 gnd.n3427 585
R2638 gnd.n3451 gnd.n3450 585
R2639 gnd.n3453 gnd.n3452 585
R2640 gnd.n3456 gnd.n3455 585
R2641 gnd.n3454 gnd.n3425 585
R2642 gnd.n3461 gnd.n3460 585
R2643 gnd.n3465 gnd.n3462 585
R2644 gnd.n3466 gnd.n3403 585
R2645 gnd.n4344 gnd.n1602 585
R2646 gnd.n4411 gnd.n4410 585
R2647 gnd.n4413 gnd.n4412 585
R2648 gnd.n4415 gnd.n4414 585
R2649 gnd.n4417 gnd.n4416 585
R2650 gnd.n4419 gnd.n4418 585
R2651 gnd.n4421 gnd.n4420 585
R2652 gnd.n4423 gnd.n4422 585
R2653 gnd.n4425 gnd.n4424 585
R2654 gnd.n4427 gnd.n4426 585
R2655 gnd.n4429 gnd.n4428 585
R2656 gnd.n4431 gnd.n4430 585
R2657 gnd.n4433 gnd.n4432 585
R2658 gnd.n4436 gnd.n4435 585
R2659 gnd.n4434 gnd.n1590 585
R2660 gnd.n4440 gnd.n1588 585
R2661 gnd.n4442 gnd.n4441 585
R2662 gnd.n4443 gnd.n4442 585
R2663 gnd.n4345 gnd.n1643 585
R2664 gnd.n4345 gnd.n1564 585
R2665 gnd.n4347 gnd.n4346 585
R2666 gnd.n4346 gnd.n1638 585
R2667 gnd.n4343 gnd.n1642 585
R2668 gnd.n4343 gnd.n4342 585
R2669 gnd.n4322 gnd.n1644 585
R2670 gnd.n3062 gnd.n1644 585
R2671 gnd.n4321 gnd.n1654 585
R2672 gnd.n4330 gnd.n1654 585
R2673 gnd.n4056 gnd.n3067 585
R2674 gnd.n4057 gnd.n4056 585
R2675 gnd.n4055 gnd.n4054 585
R2676 gnd.n4055 gnd.n3071 585
R2677 gnd.n4053 gnd.n3073 585
R2678 gnd.n4046 gnd.n3073 585
R2679 gnd.n3086 gnd.n3074 585
R2680 gnd.n3086 gnd.n3078 585
R2681 gnd.n4002 gnd.n3087 585
R2682 gnd.n4036 gnd.n3087 585
R2683 gnd.n4001 gnd.n4000 585
R2684 gnd.n4000 gnd.n3094 585
R2685 gnd.n3999 gnd.n3102 585
R2686 gnd.n3999 gnd.n3093 585
R2687 gnd.n3998 gnd.n3104 585
R2688 gnd.n3998 gnd.n3997 585
R2689 gnd.n3977 gnd.n3103 585
R2690 gnd.n3116 gnd.n3103 585
R2691 gnd.n3976 gnd.n3114 585
R2692 gnd.n3987 gnd.n3114 585
R2693 gnd.n3967 gnd.n3121 585
R2694 gnd.n3968 gnd.n3967 585
R2695 gnd.n3966 gnd.n3965 585
R2696 gnd.n3966 gnd.n3125 585
R2697 gnd.n3964 gnd.n3127 585
R2698 gnd.n3957 gnd.n3127 585
R2699 gnd.n3142 gnd.n3128 585
R2700 gnd.n3142 gnd.n3132 585
R2701 gnd.n3917 gnd.n3143 585
R2702 gnd.n3947 gnd.n3143 585
R2703 gnd.n3916 gnd.n3915 585
R2704 gnd.n3915 gnd.n3150 585
R2705 gnd.n3914 gnd.n3157 585
R2706 gnd.n3914 gnd.n3149 585
R2707 gnd.n3913 gnd.n3159 585
R2708 gnd.n3913 gnd.n3912 585
R2709 gnd.n3892 gnd.n3158 585
R2710 gnd.n3171 gnd.n3158 585
R2711 gnd.n3891 gnd.n3169 585
R2712 gnd.n3902 gnd.n3169 585
R2713 gnd.n3882 gnd.n3176 585
R2714 gnd.n3883 gnd.n3882 585
R2715 gnd.n3881 gnd.n3880 585
R2716 gnd.n3881 gnd.n3180 585
R2717 gnd.n3879 gnd.n3182 585
R2718 gnd.n3872 gnd.n3182 585
R2719 gnd.n3859 gnd.n3183 585
R2720 gnd.n3860 gnd.n3859 585
R2721 gnd.n3812 gnd.n3196 585
R2722 gnd.n3862 gnd.n3196 585
R2723 gnd.n3814 gnd.n3813 585
R2724 gnd.n3815 gnd.n3814 585
R2725 gnd.n3807 gnd.n3310 585
R2726 gnd.n3310 gnd.n3309 585
R2727 gnd.n3805 gnd.n3804 585
R2728 gnd.n3804 gnd.n3291 585
R2729 gnd.n3802 gnd.n3289 585
R2730 gnd.n3823 gnd.n3289 585
R2731 gnd.n3320 gnd.n3319 585
R2732 gnd.n3319 gnd.n3318 585
R2733 gnd.n3796 gnd.n3279 585
R2734 gnd.n3829 gnd.n3279 585
R2735 gnd.n3795 gnd.n3794 585
R2736 gnd.n3794 gnd.n3793 585
R2737 gnd.n3791 gnd.n3322 585
R2738 gnd.n3791 gnd.n3269 585
R2739 gnd.n3790 gnd.n3789 585
R2740 gnd.n3790 gnd.n3268 585
R2741 gnd.n3325 gnd.n3324 585
R2742 gnd.n3781 gnd.n3324 585
R2743 gnd.n3749 gnd.n3748 585
R2744 gnd.n3748 gnd.n3329 585
R2745 gnd.n3750 gnd.n3338 585
R2746 gnd.n3767 gnd.n3338 585
R2747 gnd.n3747 gnd.n3746 585
R2748 gnd.n3746 gnd.n3344 585
R2749 gnd.n3745 gnd.n3352 585
R2750 gnd.n3745 gnd.n3744 585
R2751 gnd.n3730 gnd.n3353 585
R2752 gnd.n3363 gnd.n3353 585
R2753 gnd.n3729 gnd.n3361 585
R2754 gnd.n3736 gnd.n3361 585
R2755 gnd.n3728 gnd.n3727 585
R2756 gnd.n3727 gnd.n3726 585
R2757 gnd.n3372 gnd.n3369 585
R2758 gnd.n3382 gnd.n3372 585
R2759 gnd.n3718 gnd.n3717 585
R2760 gnd.n3717 gnd.n3716 585
R2761 gnd.n3378 gnd.n3377 585
R2762 gnd.n3391 gnd.n3378 585
R2763 gnd.n3698 gnd.n3389 585
R2764 gnd.n3706 gnd.n3389 585
R2765 gnd.n3697 gnd.n3696 585
R2766 gnd.n3696 gnd.n3695 585
R2767 gnd.n3398 gnd.n3396 585
R2768 gnd.n3407 gnd.n3398 585
R2769 gnd.n3687 gnd.n3686 585
R2770 gnd.n3686 gnd.n3685 585
R2771 gnd.n5740 gnd.n5739 585
R2772 gnd.n5741 gnd.n5740 585
R2773 gnd.n1181 gnd.n1179 585
R2774 gnd.n5664 gnd.n1179 585
R2775 gnd.n5341 gnd.n1276 585
R2776 gnd.n5152 gnd.n1276 585
R2777 gnd.n5343 gnd.n5342 585
R2778 gnd.n5344 gnd.n5343 585
R2779 gnd.n1277 gnd.n1275 585
R2780 gnd.n5118 gnd.n1275 585
R2781 gnd.n5336 gnd.n5335 585
R2782 gnd.n5335 gnd.n5334 585
R2783 gnd.n1280 gnd.n1279 585
R2784 gnd.n5107 gnd.n1280 585
R2785 gnd.n5325 gnd.n5324 585
R2786 gnd.n5326 gnd.n5325 585
R2787 gnd.n1295 gnd.n1294 585
R2788 gnd.n5103 gnd.n1294 585
R2789 gnd.n5320 gnd.n5319 585
R2790 gnd.n5319 gnd.n5318 585
R2791 gnd.n1298 gnd.n1297 585
R2792 gnd.n5097 gnd.n1298 585
R2793 gnd.n5309 gnd.n5308 585
R2794 gnd.n5310 gnd.n5309 585
R2795 gnd.n1312 gnd.n1311 585
R2796 gnd.n5019 gnd.n1311 585
R2797 gnd.n5304 gnd.n5303 585
R2798 gnd.n5303 gnd.n5302 585
R2799 gnd.n1315 gnd.n1314 585
R2800 gnd.n5023 gnd.n1315 585
R2801 gnd.n5293 gnd.n5292 585
R2802 gnd.n5294 gnd.n5293 585
R2803 gnd.n1330 gnd.n1329 585
R2804 gnd.n5027 gnd.n1329 585
R2805 gnd.n5288 gnd.n5287 585
R2806 gnd.n5287 gnd.n5286 585
R2807 gnd.n1333 gnd.n1332 585
R2808 gnd.n5033 gnd.n1333 585
R2809 gnd.n5277 gnd.n5276 585
R2810 gnd.n5278 gnd.n5277 585
R2811 gnd.n1347 gnd.n1346 585
R2812 gnd.n5007 gnd.n1346 585
R2813 gnd.n5272 gnd.n5271 585
R2814 gnd.n5271 gnd.n5270 585
R2815 gnd.n1350 gnd.n1349 585
R2816 gnd.n5003 gnd.n1350 585
R2817 gnd.n5261 gnd.n5260 585
R2818 gnd.n5262 gnd.n5261 585
R2819 gnd.n1365 gnd.n1364 585
R2820 gnd.n4997 gnd.n1364 585
R2821 gnd.n5256 gnd.n5255 585
R2822 gnd.n5255 gnd.n5254 585
R2823 gnd.n1368 gnd.n1367 585
R2824 gnd.n4993 gnd.n1368 585
R2825 gnd.n5245 gnd.n5244 585
R2826 gnd.n5246 gnd.n5245 585
R2827 gnd.n1382 gnd.n1381 585
R2828 gnd.n5197 gnd.n1381 585
R2829 gnd.n5218 gnd.n5217 585
R2830 gnd.n5219 gnd.n5218 585
R2831 gnd.n5216 gnd.n5215 585
R2832 gnd.n5215 gnd.n1422 585
R2833 gnd.n1408 gnd.n1407 585
R2834 gnd.n1412 gnd.n1407 585
R2835 gnd.n5228 gnd.n1409 585
R2836 gnd.n5228 gnd.n5227 585
R2837 gnd.n5231 gnd.n5230 585
R2838 gnd.n5232 gnd.n5231 585
R2839 gnd.n5229 gnd.n1391 585
R2840 gnd.n1395 gnd.n1391 585
R2841 gnd.n5240 gnd.n5239 585
R2842 gnd.n5239 gnd.n5238 585
R2843 gnd.n5241 gnd.n1390 585
R2844 gnd.n4901 gnd.n1390 585
R2845 gnd.n1452 gnd.n1389 585
R2846 gnd.n1452 gnd.n1443 585
R2847 gnd.n4887 gnd.n4886 585
R2848 gnd.n4888 gnd.n4887 585
R2849 gnd.n4885 gnd.n1451 585
R2850 gnd.n4873 gnd.n1451 585
R2851 gnd.n1457 gnd.n1453 585
R2852 gnd.n1460 gnd.n1457 585
R2853 gnd.n4881 gnd.n4880 585
R2854 gnd.n4880 gnd.n4879 585
R2855 gnd.n1456 gnd.n1455 585
R2856 gnd.n4861 gnd.n1456 585
R2857 gnd.n4845 gnd.n1488 585
R2858 gnd.n1488 gnd.n1478 585
R2859 gnd.n4847 gnd.n4846 585
R2860 gnd.n4848 gnd.n4847 585
R2861 gnd.n1489 gnd.n1487 585
R2862 gnd.n1487 gnd.n1484 585
R2863 gnd.n4840 gnd.n4839 585
R2864 gnd.n4839 gnd.n4838 585
R2865 gnd.n1492 gnd.n1491 585
R2866 gnd.n1504 gnd.n1492 585
R2867 gnd.n4821 gnd.n4820 585
R2868 gnd.n4822 gnd.n4821 585
R2869 gnd.n1506 gnd.n1505 585
R2870 gnd.n1505 gnd.n1501 585
R2871 gnd.n4816 gnd.n4815 585
R2872 gnd.n4815 gnd.n4814 585
R2873 gnd.n1509 gnd.n1508 585
R2874 gnd.n1510 gnd.n1509 585
R2875 gnd.n4805 gnd.n4804 585
R2876 gnd.n4806 gnd.n4805 585
R2877 gnd.n1522 gnd.n1521 585
R2878 gnd.n1521 gnd.n1518 585
R2879 gnd.n4800 gnd.n4799 585
R2880 gnd.n4799 gnd.n4798 585
R2881 gnd.n1525 gnd.n1524 585
R2882 gnd.n1536 gnd.n1525 585
R2883 gnd.n4789 gnd.n4788 585
R2884 gnd.n4790 gnd.n4789 585
R2885 gnd.n1538 gnd.n1537 585
R2886 gnd.n1537 gnd.n1533 585
R2887 gnd.n4784 gnd.n4783 585
R2888 gnd.n4783 gnd.n4782 585
R2889 gnd.n1541 gnd.n1540 585
R2890 gnd.n1542 gnd.n1541 585
R2891 gnd.n4773 gnd.n4772 585
R2892 gnd.n4774 gnd.n4773 585
R2893 gnd.n1554 gnd.n1553 585
R2894 gnd.n1553 gnd.n1550 585
R2895 gnd.n4768 gnd.n4767 585
R2896 gnd.n4767 gnd.n4766 585
R2897 gnd.n1557 gnd.n1556 585
R2898 gnd.n4566 gnd.n1557 585
R2899 gnd.n4757 gnd.n4756 585
R2900 gnd.n4758 gnd.n4757 585
R2901 gnd.n4753 gnd.n4567 585
R2902 gnd.n4752 gnd.n4751 585
R2903 gnd.n4749 gnd.n4569 585
R2904 gnd.n4749 gnd.n4444 585
R2905 gnd.n4748 gnd.n4747 585
R2906 gnd.n4746 gnd.n4745 585
R2907 gnd.n4744 gnd.n4574 585
R2908 gnd.n4742 gnd.n4741 585
R2909 gnd.n4740 gnd.n4575 585
R2910 gnd.n4739 gnd.n4738 585
R2911 gnd.n4736 gnd.n4580 585
R2912 gnd.n4734 gnd.n4733 585
R2913 gnd.n4732 gnd.n4581 585
R2914 gnd.n4731 gnd.n4730 585
R2915 gnd.n4728 gnd.n4586 585
R2916 gnd.n4726 gnd.n4725 585
R2917 gnd.n4724 gnd.n4587 585
R2918 gnd.n4723 gnd.n4722 585
R2919 gnd.n4720 gnd.n4592 585
R2920 gnd.n4718 gnd.n4717 585
R2921 gnd.n4716 gnd.n4593 585
R2922 gnd.n4715 gnd.n4714 585
R2923 gnd.n4712 gnd.n4601 585
R2924 gnd.n4710 gnd.n4709 585
R2925 gnd.n4708 gnd.n4602 585
R2926 gnd.n4707 gnd.n4706 585
R2927 gnd.n4704 gnd.n4607 585
R2928 gnd.n4702 gnd.n4701 585
R2929 gnd.n4700 gnd.n4608 585
R2930 gnd.n4699 gnd.n4698 585
R2931 gnd.n4696 gnd.n4613 585
R2932 gnd.n4694 gnd.n4693 585
R2933 gnd.n4692 gnd.n4614 585
R2934 gnd.n4691 gnd.n4690 585
R2935 gnd.n4688 gnd.n4619 585
R2936 gnd.n4686 gnd.n4685 585
R2937 gnd.n4684 gnd.n4620 585
R2938 gnd.n4683 gnd.n4625 585
R2939 gnd.n4676 gnd.n4628 585
R2940 gnd.n4679 gnd.n4678 585
R2941 gnd.n5671 gnd.n5670 585
R2942 gnd.n5673 gnd.n1259 585
R2943 gnd.n5675 gnd.n5674 585
R2944 gnd.n5676 gnd.n1252 585
R2945 gnd.n5678 gnd.n5677 585
R2946 gnd.n5680 gnd.n1250 585
R2947 gnd.n5682 gnd.n5681 585
R2948 gnd.n5683 gnd.n1245 585
R2949 gnd.n5685 gnd.n5684 585
R2950 gnd.n5687 gnd.n1243 585
R2951 gnd.n5689 gnd.n5688 585
R2952 gnd.n5690 gnd.n1238 585
R2953 gnd.n5692 gnd.n5691 585
R2954 gnd.n5694 gnd.n1236 585
R2955 gnd.n5696 gnd.n5695 585
R2956 gnd.n5697 gnd.n1231 585
R2957 gnd.n5699 gnd.n5698 585
R2958 gnd.n5701 gnd.n1229 585
R2959 gnd.n5703 gnd.n5702 585
R2960 gnd.n5704 gnd.n1223 585
R2961 gnd.n5706 gnd.n5705 585
R2962 gnd.n5710 gnd.n1218 585
R2963 gnd.n5712 gnd.n5711 585
R2964 gnd.n5713 gnd.n1213 585
R2965 gnd.n5715 gnd.n5714 585
R2966 gnd.n5717 gnd.n1211 585
R2967 gnd.n5719 gnd.n5718 585
R2968 gnd.n5720 gnd.n1206 585
R2969 gnd.n5722 gnd.n5721 585
R2970 gnd.n5724 gnd.n1204 585
R2971 gnd.n5726 gnd.n5725 585
R2972 gnd.n5727 gnd.n1198 585
R2973 gnd.n5729 gnd.n5728 585
R2974 gnd.n5731 gnd.n1197 585
R2975 gnd.n5732 gnd.n1184 585
R2976 gnd.n5735 gnd.n5734 585
R2977 gnd.n5736 gnd.n1180 585
R2978 gnd.n1196 gnd.n1180 585
R2979 gnd.n5667 gnd.n1176 585
R2980 gnd.n5741 gnd.n1176 585
R2981 gnd.n5666 gnd.n5665 585
R2982 gnd.n5665 gnd.n5664 585
R2983 gnd.n1264 gnd.n1263 585
R2984 gnd.n5152 gnd.n1264 585
R2985 gnd.n5115 gnd.n1272 585
R2986 gnd.n5344 gnd.n1272 585
R2987 gnd.n5117 gnd.n5116 585
R2988 gnd.n5118 gnd.n5117 585
R2989 gnd.n4939 gnd.n1282 585
R2990 gnd.n5334 gnd.n1282 585
R2991 gnd.n5109 gnd.n5108 585
R2992 gnd.n5108 gnd.n5107 585
R2993 gnd.n5106 gnd.n1291 585
R2994 gnd.n5326 gnd.n1291 585
R2995 gnd.n5105 gnd.n5104 585
R2996 gnd.n5104 gnd.n5103 585
R2997 gnd.n4941 gnd.n1299 585
R2998 gnd.n5318 gnd.n1299 585
R2999 gnd.n5099 gnd.n5098 585
R3000 gnd.n5098 gnd.n5097 585
R3001 gnd.n4943 gnd.n1308 585
R3002 gnd.n5310 gnd.n1308 585
R3003 gnd.n5021 gnd.n5020 585
R3004 gnd.n5020 gnd.n5019 585
R3005 gnd.n5022 gnd.n1317 585
R3006 gnd.n5302 gnd.n1317 585
R3007 gnd.n5025 gnd.n5024 585
R3008 gnd.n5024 gnd.n5023 585
R3009 gnd.n5026 gnd.n1326 585
R3010 gnd.n5294 gnd.n1326 585
R3011 gnd.n5029 gnd.n5028 585
R3012 gnd.n5028 gnd.n5027 585
R3013 gnd.n5030 gnd.n1334 585
R3014 gnd.n5286 gnd.n1334 585
R3015 gnd.n5032 gnd.n5031 585
R3016 gnd.n5033 gnd.n5032 585
R3017 gnd.n4955 gnd.n1343 585
R3018 gnd.n5278 gnd.n1343 585
R3019 gnd.n5009 gnd.n5008 585
R3020 gnd.n5008 gnd.n5007 585
R3021 gnd.n5006 gnd.n1352 585
R3022 gnd.n5270 gnd.n1352 585
R3023 gnd.n5005 gnd.n5004 585
R3024 gnd.n5004 gnd.n5003 585
R3025 gnd.n4957 gnd.n1361 585
R3026 gnd.n5262 gnd.n1361 585
R3027 gnd.n4999 gnd.n4998 585
R3028 gnd.n4998 gnd.n4997 585
R3029 gnd.n4996 gnd.n1369 585
R3030 gnd.n5254 gnd.n1369 585
R3031 gnd.n4995 gnd.n4994 585
R3032 gnd.n4994 gnd.n4993 585
R3033 gnd.n1434 gnd.n1378 585
R3034 gnd.n5246 gnd.n1378 585
R3035 gnd.n5199 gnd.n5198 585
R3036 gnd.n5198 gnd.n5197 585
R3037 gnd.n5200 gnd.n1423 585
R3038 gnd.n5219 gnd.n1423 585
R3039 gnd.n5202 gnd.n5201 585
R3040 gnd.n5202 gnd.n1422 585
R3041 gnd.n5204 gnd.n5203 585
R3042 gnd.n5203 gnd.n1412 585
R3043 gnd.n5205 gnd.n1410 585
R3044 gnd.n5227 gnd.n1410 585
R3045 gnd.n1430 gnd.n1404 585
R3046 gnd.n5232 gnd.n1404 585
R3047 gnd.n4897 gnd.n4896 585
R3048 gnd.n4896 gnd.n1395 585
R3049 gnd.n4898 gnd.n1393 585
R3050 gnd.n5238 gnd.n1393 585
R3051 gnd.n4900 gnd.n4899 585
R3052 gnd.n4901 gnd.n4900 585
R3053 gnd.n1445 gnd.n1444 585
R3054 gnd.n1444 gnd.n1443 585
R3055 gnd.n4890 gnd.n4889 585
R3056 gnd.n4889 gnd.n4888 585
R3057 gnd.n1448 gnd.n1447 585
R3058 gnd.n4873 gnd.n1448 585
R3059 gnd.n4857 gnd.n4856 585
R3060 gnd.n4856 gnd.n1460 585
R3061 gnd.n4858 gnd.n1458 585
R3062 gnd.n4879 gnd.n1458 585
R3063 gnd.n4860 gnd.n4859 585
R3064 gnd.n4861 gnd.n4860 585
R3065 gnd.n1480 gnd.n1479 585
R3066 gnd.n1479 gnd.n1478 585
R3067 gnd.n4850 gnd.n4849 585
R3068 gnd.n4849 gnd.n4848 585
R3069 gnd.n1483 gnd.n1482 585
R3070 gnd.n1484 gnd.n1483 585
R3071 gnd.n4648 gnd.n1493 585
R3072 gnd.n4838 gnd.n1493 585
R3073 gnd.n4650 gnd.n4649 585
R3074 gnd.n4649 gnd.n1504 585
R3075 gnd.n4651 gnd.n1502 585
R3076 gnd.n4822 gnd.n1502 585
R3077 gnd.n4653 gnd.n4652 585
R3078 gnd.n4652 gnd.n1501 585
R3079 gnd.n4654 gnd.n1511 585
R3080 gnd.n4814 gnd.n1511 585
R3081 gnd.n4656 gnd.n4655 585
R3082 gnd.n4655 gnd.n1510 585
R3083 gnd.n4657 gnd.n1519 585
R3084 gnd.n4806 gnd.n1519 585
R3085 gnd.n4659 gnd.n4658 585
R3086 gnd.n4658 gnd.n1518 585
R3087 gnd.n4660 gnd.n1526 585
R3088 gnd.n4798 gnd.n1526 585
R3089 gnd.n4662 gnd.n4661 585
R3090 gnd.n4661 gnd.n1536 585
R3091 gnd.n4663 gnd.n1534 585
R3092 gnd.n4790 gnd.n1534 585
R3093 gnd.n4665 gnd.n4664 585
R3094 gnd.n4664 gnd.n1533 585
R3095 gnd.n4666 gnd.n1543 585
R3096 gnd.n4782 gnd.n1543 585
R3097 gnd.n4668 gnd.n4667 585
R3098 gnd.n4667 gnd.n1542 585
R3099 gnd.n4669 gnd.n1551 585
R3100 gnd.n4774 gnd.n1551 585
R3101 gnd.n4671 gnd.n4670 585
R3102 gnd.n4670 gnd.n1550 585
R3103 gnd.n4672 gnd.n1558 585
R3104 gnd.n4766 gnd.n1558 585
R3105 gnd.n4673 gnd.n4630 585
R3106 gnd.n4630 gnd.n4566 585
R3107 gnd.n4674 gnd.n4445 585
R3108 gnd.n4758 gnd.n4445 585
R3109 gnd.n7836 gnd.n7835 585
R3110 gnd.n7837 gnd.n7836 585
R3111 gnd.n132 gnd.n130 585
R3112 gnd.n130 gnd.n126 585
R3113 gnd.n7756 gnd.n7755 585
R3114 gnd.n7757 gnd.n7756 585
R3115 gnd.n209 gnd.n208 585
R3116 gnd.n208 gnd.n206 585
R3117 gnd.n7751 gnd.n7750 585
R3118 gnd.n7750 gnd.n7749 585
R3119 gnd.n212 gnd.n211 585
R3120 gnd.n213 gnd.n212 585
R3121 gnd.n7672 gnd.n7671 585
R3122 gnd.n7673 gnd.n7672 585
R3123 gnd.n225 gnd.n224 585
R3124 gnd.n7492 gnd.n224 585
R3125 gnd.n7667 gnd.n7666 585
R3126 gnd.n7666 gnd.n7665 585
R3127 gnd.n228 gnd.n227 585
R3128 gnd.n229 gnd.n228 585
R3129 gnd.n7656 gnd.n7655 585
R3130 gnd.n7657 gnd.n7656 585
R3131 gnd.n241 gnd.n240 585
R3132 gnd.n240 gnd.n238 585
R3133 gnd.n7651 gnd.n7650 585
R3134 gnd.n7650 gnd.n7649 585
R3135 gnd.n244 gnd.n243 585
R3136 gnd.n253 gnd.n244 585
R3137 gnd.n7640 gnd.n7639 585
R3138 gnd.n7641 gnd.n7640 585
R3139 gnd.n255 gnd.n254 585
R3140 gnd.n262 gnd.n254 585
R3141 gnd.n7635 gnd.n7634 585
R3142 gnd.n7634 gnd.n7633 585
R3143 gnd.n258 gnd.n257 585
R3144 gnd.n259 gnd.n258 585
R3145 gnd.n7624 gnd.n7623 585
R3146 gnd.n7625 gnd.n7624 585
R3147 gnd.n271 gnd.n270 585
R3148 gnd.n270 gnd.n268 585
R3149 gnd.n7619 gnd.n7618 585
R3150 gnd.n7618 gnd.n7617 585
R3151 gnd.n274 gnd.n273 585
R3152 gnd.n283 gnd.n274 585
R3153 gnd.n7608 gnd.n7607 585
R3154 gnd.n7609 gnd.n7608 585
R3155 gnd.n285 gnd.n284 585
R3156 gnd.n292 gnd.n284 585
R3157 gnd.n7603 gnd.n7602 585
R3158 gnd.n7602 gnd.n7601 585
R3159 gnd.n288 gnd.n287 585
R3160 gnd.n289 gnd.n288 585
R3161 gnd.n7592 gnd.n7591 585
R3162 gnd.n7593 gnd.n7592 585
R3163 gnd.n301 gnd.n300 585
R3164 gnd.n300 gnd.n298 585
R3165 gnd.n7568 gnd.n7567 585
R3166 gnd.n7569 gnd.n7568 585
R3167 gnd.n7566 gnd.n331 585
R3168 gnd.n7566 gnd.n7565 585
R3169 gnd.n330 gnd.n329 585
R3170 gnd.n333 gnd.n329 585
R3171 gnd.n7554 gnd.n7553 585
R3172 gnd.n7555 gnd.n7554 585
R3173 gnd.n7552 gnd.n7551 585
R3174 gnd.n7551 gnd.n343 585
R3175 gnd.n7550 gnd.n347 585
R3176 gnd.n7550 gnd.n7549 585
R3177 gnd.n346 gnd.n310 585
R3178 gnd.n7533 gnd.n310 585
R3179 gnd.n7586 gnd.n7585 585
R3180 gnd.n7585 gnd.n7584 585
R3181 gnd.n7587 gnd.n309 585
R3182 gnd.n7539 gnd.n309 585
R3183 gnd.n367 gnd.n308 585
R3184 gnd.n7427 gnd.n367 585
R3185 gnd.n7446 gnd.n7445 585
R3186 gnd.n7447 gnd.n7446 585
R3187 gnd.n7444 gnd.n366 585
R3188 gnd.n7425 gnd.n366 585
R3189 gnd.n372 gnd.n368 585
R3190 gnd.n7409 gnd.n372 585
R3191 gnd.n7440 gnd.n7439 585
R3192 gnd.n7439 gnd.n7438 585
R3193 gnd.n371 gnd.n370 585
R3194 gnd.n7415 gnd.n371 585
R3195 gnd.n7398 gnd.n400 585
R3196 gnd.n7382 gnd.n400 585
R3197 gnd.n7400 gnd.n7399 585
R3198 gnd.n7401 gnd.n7400 585
R3199 gnd.n401 gnd.n399 585
R3200 gnd.n7332 gnd.n399 585
R3201 gnd.n7393 gnd.n7392 585
R3202 gnd.n7392 gnd.n7391 585
R3203 gnd.n404 gnd.n403 585
R3204 gnd.n7341 gnd.n404 585
R3205 gnd.n7322 gnd.n435 585
R3206 gnd.n435 gnd.n422 585
R3207 gnd.n7324 gnd.n7323 585
R3208 gnd.n7325 gnd.n7324 585
R3209 gnd.n436 gnd.n434 585
R3210 gnd.n7145 gnd.n434 585
R3211 gnd.n7317 gnd.n7316 585
R3212 gnd.n7316 gnd.n7315 585
R3213 gnd.n439 gnd.n438 585
R3214 gnd.n7151 gnd.n439 585
R3215 gnd.n7300 gnd.n7299 585
R3216 gnd.n7301 gnd.n7300 585
R3217 gnd.n456 gnd.n455 585
R3218 gnd.n7128 gnd.n455 585
R3219 gnd.n7295 gnd.n7294 585
R3220 gnd.n7294 gnd.n7293 585
R3221 gnd.n459 gnd.n458 585
R3222 gnd.n617 gnd.n459 585
R3223 gnd.n7284 gnd.n7283 585
R3224 gnd.n7285 gnd.n7284 585
R3225 gnd.n473 gnd.n472 585
R3226 gnd.n611 gnd.n472 585
R3227 gnd.n7279 gnd.n7278 585
R3228 gnd.n7278 gnd.n7277 585
R3229 gnd.n476 gnd.n475 585
R3230 gnd.n607 gnd.n476 585
R3231 gnd.n7268 gnd.n7267 585
R3232 gnd.n7269 gnd.n7268 585
R3233 gnd.n491 gnd.n490 585
R3234 gnd.n601 gnd.n490 585
R3235 gnd.n7263 gnd.n7262 585
R3236 gnd.n7262 gnd.n7261 585
R3237 gnd.n494 gnd.n493 585
R3238 gnd.n7176 gnd.n494 585
R3239 gnd.n7250 gnd.n7249 585
R3240 gnd.n7248 gnd.n534 585
R3241 gnd.n7247 gnd.n533 585
R3242 gnd.n7252 gnd.n533 585
R3243 gnd.n7246 gnd.n7245 585
R3244 gnd.n7244 gnd.n7243 585
R3245 gnd.n7242 gnd.n7241 585
R3246 gnd.n7240 gnd.n7239 585
R3247 gnd.n7238 gnd.n7237 585
R3248 gnd.n7236 gnd.n7235 585
R3249 gnd.n7234 gnd.n7233 585
R3250 gnd.n7232 gnd.n7231 585
R3251 gnd.n7230 gnd.n7229 585
R3252 gnd.n7228 gnd.n7227 585
R3253 gnd.n7226 gnd.n7225 585
R3254 gnd.n7224 gnd.n7223 585
R3255 gnd.n7222 gnd.n7221 585
R3256 gnd.n7219 gnd.n7218 585
R3257 gnd.n7217 gnd.n7216 585
R3258 gnd.n7215 gnd.n7214 585
R3259 gnd.n7213 gnd.n7212 585
R3260 gnd.n7211 gnd.n7210 585
R3261 gnd.n7209 gnd.n7208 585
R3262 gnd.n7207 gnd.n7206 585
R3263 gnd.n7205 gnd.n7204 585
R3264 gnd.n7203 gnd.n7202 585
R3265 gnd.n7201 gnd.n7200 585
R3266 gnd.n7199 gnd.n7198 585
R3267 gnd.n7197 gnd.n7196 585
R3268 gnd.n7195 gnd.n7194 585
R3269 gnd.n7193 gnd.n7192 585
R3270 gnd.n7191 gnd.n7190 585
R3271 gnd.n7189 gnd.n7188 585
R3272 gnd.n7187 gnd.n7186 585
R3273 gnd.n7185 gnd.n7184 585
R3274 gnd.n7183 gnd.n574 585
R3275 gnd.n578 gnd.n575 585
R3276 gnd.n7179 gnd.n7178 585
R3277 gnd.n200 gnd.n199 585
R3278 gnd.n7765 gnd.n195 585
R3279 gnd.n7767 gnd.n7766 585
R3280 gnd.n7769 gnd.n193 585
R3281 gnd.n7771 gnd.n7770 585
R3282 gnd.n7772 gnd.n188 585
R3283 gnd.n7774 gnd.n7773 585
R3284 gnd.n7776 gnd.n186 585
R3285 gnd.n7778 gnd.n7777 585
R3286 gnd.n7779 gnd.n181 585
R3287 gnd.n7781 gnd.n7780 585
R3288 gnd.n7783 gnd.n179 585
R3289 gnd.n7785 gnd.n7784 585
R3290 gnd.n7786 gnd.n174 585
R3291 gnd.n7788 gnd.n7787 585
R3292 gnd.n7790 gnd.n172 585
R3293 gnd.n7792 gnd.n7791 585
R3294 gnd.n7793 gnd.n167 585
R3295 gnd.n7795 gnd.n7794 585
R3296 gnd.n7797 gnd.n165 585
R3297 gnd.n7799 gnd.n7798 585
R3298 gnd.n7803 gnd.n160 585
R3299 gnd.n7805 gnd.n7804 585
R3300 gnd.n7807 gnd.n158 585
R3301 gnd.n7809 gnd.n7808 585
R3302 gnd.n7810 gnd.n153 585
R3303 gnd.n7812 gnd.n7811 585
R3304 gnd.n7814 gnd.n151 585
R3305 gnd.n7816 gnd.n7815 585
R3306 gnd.n7817 gnd.n146 585
R3307 gnd.n7819 gnd.n7818 585
R3308 gnd.n7821 gnd.n144 585
R3309 gnd.n7823 gnd.n7822 585
R3310 gnd.n7824 gnd.n139 585
R3311 gnd.n7826 gnd.n7825 585
R3312 gnd.n7828 gnd.n137 585
R3313 gnd.n7830 gnd.n7829 585
R3314 gnd.n7831 gnd.n135 585
R3315 gnd.n7832 gnd.n131 585
R3316 gnd.n131 gnd.n128 585
R3317 gnd.n7761 gnd.n127 585
R3318 gnd.n7837 gnd.n127 585
R3319 gnd.n7760 gnd.n7759 585
R3320 gnd.n7759 gnd.n126 585
R3321 gnd.n7758 gnd.n204 585
R3322 gnd.n7758 gnd.n7757 585
R3323 gnd.n7487 gnd.n205 585
R3324 gnd.n206 gnd.n205 585
R3325 gnd.n7488 gnd.n214 585
R3326 gnd.n7749 gnd.n214 585
R3327 gnd.n7490 gnd.n7489 585
R3328 gnd.n7489 gnd.n213 585
R3329 gnd.n7491 gnd.n223 585
R3330 gnd.n7673 gnd.n223 585
R3331 gnd.n7494 gnd.n7493 585
R3332 gnd.n7493 gnd.n7492 585
R3333 gnd.n7495 gnd.n230 585
R3334 gnd.n7665 gnd.n230 585
R3335 gnd.n7497 gnd.n7496 585
R3336 gnd.n7496 gnd.n229 585
R3337 gnd.n7498 gnd.n239 585
R3338 gnd.n7657 gnd.n239 585
R3339 gnd.n7500 gnd.n7499 585
R3340 gnd.n7499 gnd.n238 585
R3341 gnd.n7501 gnd.n245 585
R3342 gnd.n7649 gnd.n245 585
R3343 gnd.n7503 gnd.n7502 585
R3344 gnd.n7502 gnd.n253 585
R3345 gnd.n7504 gnd.n252 585
R3346 gnd.n7641 gnd.n252 585
R3347 gnd.n7506 gnd.n7505 585
R3348 gnd.n7505 gnd.n262 585
R3349 gnd.n7507 gnd.n260 585
R3350 gnd.n7633 gnd.n260 585
R3351 gnd.n7509 gnd.n7508 585
R3352 gnd.n7508 gnd.n259 585
R3353 gnd.n7510 gnd.n269 585
R3354 gnd.n7625 gnd.n269 585
R3355 gnd.n7512 gnd.n7511 585
R3356 gnd.n7511 gnd.n268 585
R3357 gnd.n7513 gnd.n275 585
R3358 gnd.n7617 gnd.n275 585
R3359 gnd.n7515 gnd.n7514 585
R3360 gnd.n7514 gnd.n283 585
R3361 gnd.n7516 gnd.n282 585
R3362 gnd.n7609 gnd.n282 585
R3363 gnd.n7518 gnd.n7517 585
R3364 gnd.n7517 gnd.n292 585
R3365 gnd.n7519 gnd.n290 585
R3366 gnd.n7601 gnd.n290 585
R3367 gnd.n7521 gnd.n7520 585
R3368 gnd.n7520 gnd.n289 585
R3369 gnd.n7522 gnd.n299 585
R3370 gnd.n7593 gnd.n299 585
R3371 gnd.n7524 gnd.n7523 585
R3372 gnd.n7523 gnd.n298 585
R3373 gnd.n7525 gnd.n327 585
R3374 gnd.n7569 gnd.n327 585
R3375 gnd.n7526 gnd.n334 585
R3376 gnd.n7565 gnd.n334 585
R3377 gnd.n7528 gnd.n7527 585
R3378 gnd.n7527 gnd.n333 585
R3379 gnd.n7529 gnd.n344 585
R3380 gnd.n7555 gnd.n344 585
R3381 gnd.n7531 gnd.n7530 585
R3382 gnd.n7530 gnd.n343 585
R3383 gnd.n7532 gnd.n349 585
R3384 gnd.n7549 gnd.n349 585
R3385 gnd.n7535 gnd.n7534 585
R3386 gnd.n7534 gnd.n7533 585
R3387 gnd.n7536 gnd.n312 585
R3388 gnd.n7584 gnd.n312 585
R3389 gnd.n7538 gnd.n7537 585
R3390 gnd.n7539 gnd.n7538 585
R3391 gnd.n358 gnd.n357 585
R3392 gnd.n7427 gnd.n357 585
R3393 gnd.n7449 gnd.n7448 585
R3394 gnd.n7448 gnd.n7447 585
R3395 gnd.n361 gnd.n360 585
R3396 gnd.n7425 gnd.n361 585
R3397 gnd.n7411 gnd.n7410 585
R3398 gnd.n7410 gnd.n7409 585
R3399 gnd.n7412 gnd.n374 585
R3400 gnd.n7438 gnd.n374 585
R3401 gnd.n7414 gnd.n7413 585
R3402 gnd.n7415 gnd.n7414 585
R3403 gnd.n392 gnd.n391 585
R3404 gnd.n7382 gnd.n391 585
R3405 gnd.n7403 gnd.n7402 585
R3406 gnd.n7402 gnd.n7401 585
R3407 gnd.n395 gnd.n394 585
R3408 gnd.n7332 gnd.n395 585
R3409 gnd.n7140 gnd.n406 585
R3410 gnd.n7391 gnd.n406 585
R3411 gnd.n7141 gnd.n423 585
R3412 gnd.n7341 gnd.n423 585
R3413 gnd.n7143 gnd.n7142 585
R3414 gnd.n7142 gnd.n422 585
R3415 gnd.n7144 gnd.n431 585
R3416 gnd.n7325 gnd.n431 585
R3417 gnd.n7147 gnd.n7146 585
R3418 gnd.n7146 gnd.n7145 585
R3419 gnd.n7148 gnd.n441 585
R3420 gnd.n7315 gnd.n441 585
R3421 gnd.n7150 gnd.n7149 585
R3422 gnd.n7151 gnd.n7150 585
R3423 gnd.n594 gnd.n452 585
R3424 gnd.n7301 gnd.n452 585
R3425 gnd.n7130 gnd.n7129 585
R3426 gnd.n7129 gnd.n7128 585
R3427 gnd.n620 gnd.n461 585
R3428 gnd.n7293 gnd.n461 585
R3429 gnd.n619 gnd.n618 585
R3430 gnd.n618 gnd.n617 585
R3431 gnd.n596 gnd.n469 585
R3432 gnd.n7285 gnd.n469 585
R3433 gnd.n613 gnd.n612 585
R3434 gnd.n612 gnd.n611 585
R3435 gnd.n610 gnd.n478 585
R3436 gnd.n7277 gnd.n478 585
R3437 gnd.n609 gnd.n608 585
R3438 gnd.n608 gnd.n607 585
R3439 gnd.n598 gnd.n487 585
R3440 gnd.n7269 gnd.n487 585
R3441 gnd.n603 gnd.n602 585
R3442 gnd.n602 gnd.n601 585
R3443 gnd.n600 gnd.n496 585
R3444 gnd.n7261 gnd.n496 585
R3445 gnd.n7177 gnd.n580 585
R3446 gnd.n7177 gnd.n7176 585
R3447 gnd.n6566 gnd.n6129 585
R3448 gnd.n6566 gnd.n6565 585
R3449 gnd.n6568 gnd.n6567 585
R3450 gnd.n6567 gnd.n728 585
R3451 gnd.n6569 gnd.n6127 585
R3452 gnd.n6127 gnd.n726 585
R3453 gnd.n6571 gnd.n6570 585
R3454 gnd.n6572 gnd.n6571 585
R3455 gnd.n6128 gnd.n6126 585
R3456 gnd.n6126 gnd.n735 585
R3457 gnd.n6366 gnd.n6365 585
R3458 gnd.n6367 gnd.n6366 585
R3459 gnd.n6364 gnd.n6137 585
R3460 gnd.n6137 gnd.n6136 585
R3461 gnd.n6363 gnd.n6362 585
R3462 gnd.n6362 gnd.n742 585
R3463 gnd.n6361 gnd.n6138 585
R3464 gnd.n6361 gnd.n6360 585
R3465 gnd.n6347 gnd.n6139 585
R3466 gnd.n6139 gnd.n750 585
R3467 gnd.n6348 gnd.n748 585
R3468 gnd.n6969 gnd.n748 585
R3469 gnd.n6350 gnd.n6349 585
R3470 gnd.n6351 gnd.n6350 585
R3471 gnd.n6346 gnd.n6146 585
R3472 gnd.n6146 gnd.n759 585
R3473 gnd.n6345 gnd.n6344 585
R3474 gnd.n6344 gnd.n757 585
R3475 gnd.n6343 gnd.n6147 585
R3476 gnd.n6343 gnd.n6342 585
R3477 gnd.n6330 gnd.n6148 585
R3478 gnd.n6148 gnd.n767 585
R3479 gnd.n6331 gnd.n6156 585
R3480 gnd.n6156 gnd.n765 585
R3481 gnd.n6333 gnd.n6332 585
R3482 gnd.n6334 gnd.n6333 585
R3483 gnd.n6329 gnd.n6155 585
R3484 gnd.n6155 gnd.n775 585
R3485 gnd.n6328 gnd.n6327 585
R3486 gnd.n6327 gnd.n773 585
R3487 gnd.n6326 gnd.n6157 585
R3488 gnd.n6326 gnd.n6325 585
R3489 gnd.n6312 gnd.n6158 585
R3490 gnd.n6158 gnd.n783 585
R3491 gnd.n6313 gnd.n6166 585
R3492 gnd.n6166 gnd.n781 585
R3493 gnd.n6315 gnd.n6314 585
R3494 gnd.n6316 gnd.n6315 585
R3495 gnd.n6311 gnd.n6165 585
R3496 gnd.n6165 gnd.n791 585
R3497 gnd.n6310 gnd.n6309 585
R3498 gnd.n6309 gnd.n789 585
R3499 gnd.n6308 gnd.n6167 585
R3500 gnd.n6308 gnd.n6307 585
R3501 gnd.n6294 gnd.n6168 585
R3502 gnd.n6168 gnd.n799 585
R3503 gnd.n6295 gnd.n6177 585
R3504 gnd.n6177 gnd.n797 585
R3505 gnd.n6297 gnd.n6296 585
R3506 gnd.n6298 gnd.n6297 585
R3507 gnd.n6293 gnd.n6176 585
R3508 gnd.n6176 gnd.n6175 585
R3509 gnd.n6292 gnd.n6291 585
R3510 gnd.n6291 gnd.n805 585
R3511 gnd.n6290 gnd.n6178 585
R3512 gnd.n6290 gnd.n6289 585
R3513 gnd.n6276 gnd.n6179 585
R3514 gnd.n6179 gnd.n814 585
R3515 gnd.n6277 gnd.n6186 585
R3516 gnd.n6186 gnd.n812 585
R3517 gnd.n6279 gnd.n6278 585
R3518 gnd.n6280 gnd.n6279 585
R3519 gnd.n6275 gnd.n6185 585
R3520 gnd.n6185 gnd.n822 585
R3521 gnd.n6274 gnd.n6273 585
R3522 gnd.n6273 gnd.n820 585
R3523 gnd.n6272 gnd.n6187 585
R3524 gnd.n6272 gnd.n6271 585
R3525 gnd.n6257 gnd.n6188 585
R3526 gnd.n6188 gnd.n830 585
R3527 gnd.n6258 gnd.n6195 585
R3528 gnd.n6195 gnd.n828 585
R3529 gnd.n6260 gnd.n6259 585
R3530 gnd.n6261 gnd.n6260 585
R3531 gnd.n6256 gnd.n6194 585
R3532 gnd.n6194 gnd.n838 585
R3533 gnd.n6255 gnd.n6254 585
R3534 gnd.n6254 gnd.n836 585
R3535 gnd.n6253 gnd.n6196 585
R3536 gnd.n6253 gnd.n6252 585
R3537 gnd.n6238 gnd.n6197 585
R3538 gnd.n6197 gnd.n846 585
R3539 gnd.n6239 gnd.n6204 585
R3540 gnd.n6204 gnd.n844 585
R3541 gnd.n6241 gnd.n6240 585
R3542 gnd.n6242 gnd.n6241 585
R3543 gnd.n6237 gnd.n6203 585
R3544 gnd.n6203 gnd.n854 585
R3545 gnd.n6236 gnd.n6235 585
R3546 gnd.n6235 gnd.n852 585
R3547 gnd.n6234 gnd.n6205 585
R3548 gnd.n6234 gnd.n6233 585
R3549 gnd.n6219 gnd.n6206 585
R3550 gnd.n6206 gnd.n862 585
R3551 gnd.n6220 gnd.n6217 585
R3552 gnd.n6217 gnd.n860 585
R3553 gnd.n6222 gnd.n6221 585
R3554 gnd.n6223 gnd.n6222 585
R3555 gnd.n6218 gnd.n6216 585
R3556 gnd.n6216 gnd.n870 585
R3557 gnd.n898 gnd.n897 585
R3558 gnd.n898 gnd.n868 585
R3559 gnd.n6823 gnd.n6822 585
R3560 gnd.n6822 gnd.n6821 585
R3561 gnd.n6824 gnd.n895 585
R3562 gnd.n895 gnd.n877 585
R3563 gnd.n6826 gnd.n6825 585
R3564 gnd.n6827 gnd.n6826 585
R3565 gnd.n896 gnd.n894 585
R3566 gnd.n894 gnd.n893 585
R3567 gnd.n6051 gnd.n884 585
R3568 gnd.n6833 gnd.n884 585
R3569 gnd.n6052 gnd.n929 585
R3570 gnd.n929 gnd.n883 585
R3571 gnd.n6054 gnd.n6053 585
R3572 gnd.n6055 gnd.n6054 585
R3573 gnd.n6050 gnd.n928 585
R3574 gnd.n6040 gnd.n928 585
R3575 gnd.n6049 gnd.n6048 585
R3576 gnd.n6048 gnd.n909 585
R3577 gnd.n6047 gnd.n930 585
R3578 gnd.n6047 gnd.n6046 585
R3579 gnd.n6026 gnd.n931 585
R3580 gnd.n933 gnd.n931 585
R3581 gnd.n6028 gnd.n6027 585
R3582 gnd.n6027 gnd.n919 585
R3583 gnd.n6029 gnd.n942 585
R3584 gnd.n942 gnd.n917 585
R3585 gnd.n6031 gnd.n6030 585
R3586 gnd.n6032 gnd.n6031 585
R3587 gnd.n6025 gnd.n941 585
R3588 gnd.n941 gnd.n939 585
R3589 gnd.n6024 gnd.n6023 585
R3590 gnd.n6023 gnd.n6022 585
R3591 gnd.n944 gnd.n943 585
R3592 gnd.n5943 gnd.n944 585
R3593 gnd.n5930 gnd.n5929 585
R3594 gnd.n5929 gnd.n955 585
R3595 gnd.n5931 gnd.n5926 585
R3596 gnd.n5926 gnd.n953 585
R3597 gnd.n5933 gnd.n5932 585
R3598 gnd.n5934 gnd.n5933 585
R3599 gnd.n5928 gnd.n5925 585
R3600 gnd.n5925 gnd.n965 585
R3601 gnd.n5927 gnd.n1000 585
R3602 gnd.n1000 gnd.n963 585
R3603 gnd.n5964 gnd.n999 585
R3604 gnd.n5964 gnd.n5963 585
R3605 gnd.n5966 gnd.n5965 585
R3606 gnd.n5965 gnd.n973 585
R3607 gnd.n5967 gnd.n997 585
R3608 gnd.n997 gnd.n971 585
R3609 gnd.n5969 gnd.n5968 585
R3610 gnd.n5970 gnd.n5969 585
R3611 gnd.n998 gnd.n996 585
R3612 gnd.n996 gnd.n981 585
R3613 gnd.n5385 gnd.n5384 585
R3614 gnd.n5385 gnd.n979 585
R3615 gnd.n5389 gnd.n5388 585
R3616 gnd.n5388 gnd.n5387 585
R3617 gnd.n5390 gnd.n987 585
R3618 gnd.n5978 gnd.n987 585
R3619 gnd.n5391 gnd.n5383 585
R3620 gnd.n5383 gnd.n1011 585
R3621 gnd.n5393 gnd.n5392 585
R3622 gnd.n5393 gnd.n1010 585
R3623 gnd.n5614 gnd.n5382 585
R3624 gnd.n5614 gnd.n5613 585
R3625 gnd.n5616 gnd.n5615 585
R3626 gnd.n5615 gnd.n1020 585
R3627 gnd.n5617 gnd.n5380 585
R3628 gnd.n5380 gnd.n1018 585
R3629 gnd.n5619 gnd.n5618 585
R3630 gnd.n5620 gnd.n5619 585
R3631 gnd.n5381 gnd.n5379 585
R3632 gnd.n5379 gnd.n1028 585
R3633 gnd.n5600 gnd.n5599 585
R3634 gnd.n5601 gnd.n5600 585
R3635 gnd.n5598 gnd.n5401 585
R3636 gnd.n5401 gnd.n5400 585
R3637 gnd.n5597 gnd.n5596 585
R3638 gnd.n5596 gnd.n1035 585
R3639 gnd.n5595 gnd.n5594 585
R3640 gnd.n5593 gnd.n5592 585
R3641 gnd.n5591 gnd.n5424 585
R3642 gnd.n5591 gnd.n1042 585
R3643 gnd.n5590 gnd.n5589 585
R3644 gnd.n5588 gnd.n5587 585
R3645 gnd.n5586 gnd.n5426 585
R3646 gnd.n5584 gnd.n5583 585
R3647 gnd.n5582 gnd.n5427 585
R3648 gnd.n5581 gnd.n5580 585
R3649 gnd.n5578 gnd.n5428 585
R3650 gnd.n5576 gnd.n5575 585
R3651 gnd.n5574 gnd.n5429 585
R3652 gnd.n5573 gnd.n5572 585
R3653 gnd.n5570 gnd.n5430 585
R3654 gnd.n5568 gnd.n5567 585
R3655 gnd.n5566 gnd.n5431 585
R3656 gnd.n5565 gnd.n5564 585
R3657 gnd.n5562 gnd.n5432 585
R3658 gnd.n5560 gnd.n5559 585
R3659 gnd.n5558 gnd.n5433 585
R3660 gnd.n5557 gnd.n5556 585
R3661 gnd.n5554 gnd.n5434 585
R3662 gnd.n5552 gnd.n5551 585
R3663 gnd.n5550 gnd.n5435 585
R3664 gnd.n5549 gnd.n5548 585
R3665 gnd.n5546 gnd.n5436 585
R3666 gnd.n5544 gnd.n5543 585
R3667 gnd.n5542 gnd.n5437 585
R3668 gnd.n5541 gnd.n5540 585
R3669 gnd.n5538 gnd.n5537 585
R3670 gnd.n5536 gnd.n5535 585
R3671 gnd.n5534 gnd.n5442 585
R3672 gnd.n5531 gnd.n5530 585
R3673 gnd.n5529 gnd.n5444 585
R3674 gnd.n5527 gnd.n5526 585
R3675 gnd.n5525 gnd.n5445 585
R3676 gnd.n5523 gnd.n5522 585
R3677 gnd.n5520 gnd.n5448 585
R3678 gnd.n5518 gnd.n5517 585
R3679 gnd.n5516 gnd.n5449 585
R3680 gnd.n5515 gnd.n5514 585
R3681 gnd.n5512 gnd.n5450 585
R3682 gnd.n5510 gnd.n5509 585
R3683 gnd.n5508 gnd.n5451 585
R3684 gnd.n5507 gnd.n5506 585
R3685 gnd.n5504 gnd.n5452 585
R3686 gnd.n5502 gnd.n5501 585
R3687 gnd.n5500 gnd.n5453 585
R3688 gnd.n5499 gnd.n5498 585
R3689 gnd.n5496 gnd.n5454 585
R3690 gnd.n5494 gnd.n5493 585
R3691 gnd.n5492 gnd.n5455 585
R3692 gnd.n5491 gnd.n5490 585
R3693 gnd.n5488 gnd.n5456 585
R3694 gnd.n5486 gnd.n5485 585
R3695 gnd.n5484 gnd.n5457 585
R3696 gnd.n5483 gnd.n5482 585
R3697 gnd.n5480 gnd.n5458 585
R3698 gnd.n5478 gnd.n5477 585
R3699 gnd.n5476 gnd.n5459 585
R3700 gnd.n5475 gnd.n5474 585
R3701 gnd.n5472 gnd.n5460 585
R3702 gnd.n5470 gnd.n5469 585
R3703 gnd.n5468 gnd.n5461 585
R3704 gnd.n5467 gnd.n5466 585
R3705 gnd.n6562 gnd.n6132 585
R3706 gnd.n6561 gnd.n6560 585
R3707 gnd.n6558 gnd.n6375 585
R3708 gnd.n6556 gnd.n6555 585
R3709 gnd.n6554 gnd.n6376 585
R3710 gnd.n6553 gnd.n6552 585
R3711 gnd.n6550 gnd.n6377 585
R3712 gnd.n6548 gnd.n6547 585
R3713 gnd.n6546 gnd.n6378 585
R3714 gnd.n6545 gnd.n6544 585
R3715 gnd.n6542 gnd.n6379 585
R3716 gnd.n6540 gnd.n6539 585
R3717 gnd.n6538 gnd.n6380 585
R3718 gnd.n6537 gnd.n6536 585
R3719 gnd.n6534 gnd.n6381 585
R3720 gnd.n6532 gnd.n6531 585
R3721 gnd.n6530 gnd.n6382 585
R3722 gnd.n6529 gnd.n6528 585
R3723 gnd.n6526 gnd.n6383 585
R3724 gnd.n6524 gnd.n6523 585
R3725 gnd.n6522 gnd.n6384 585
R3726 gnd.n6521 gnd.n6520 585
R3727 gnd.n6518 gnd.n6385 585
R3728 gnd.n6516 gnd.n6515 585
R3729 gnd.n6514 gnd.n6386 585
R3730 gnd.n6513 gnd.n6512 585
R3731 gnd.n6510 gnd.n6387 585
R3732 gnd.n6508 gnd.n6507 585
R3733 gnd.n6506 gnd.n6388 585
R3734 gnd.n6504 gnd.n6503 585
R3735 gnd.n6501 gnd.n6391 585
R3736 gnd.n6499 gnd.n6498 585
R3737 gnd.n6497 gnd.n720 585
R3738 gnd.n6494 gnd.n551 585
R3739 gnd.n6493 gnd.n6492 585
R3740 gnd.n6491 gnd.n6490 585
R3741 gnd.n6489 gnd.n6393 585
R3742 gnd.n6487 gnd.n6486 585
R3743 gnd.n6482 gnd.n6394 585
R3744 gnd.n6481 gnd.n6480 585
R3745 gnd.n6478 gnd.n6395 585
R3746 gnd.n6476 gnd.n6475 585
R3747 gnd.n6474 gnd.n6396 585
R3748 gnd.n6473 gnd.n6472 585
R3749 gnd.n6470 gnd.n6397 585
R3750 gnd.n6468 gnd.n6467 585
R3751 gnd.n6466 gnd.n6398 585
R3752 gnd.n6465 gnd.n6464 585
R3753 gnd.n6462 gnd.n6399 585
R3754 gnd.n6460 gnd.n6459 585
R3755 gnd.n6458 gnd.n6400 585
R3756 gnd.n6457 gnd.n6456 585
R3757 gnd.n6454 gnd.n6401 585
R3758 gnd.n6452 gnd.n6451 585
R3759 gnd.n6450 gnd.n6402 585
R3760 gnd.n6449 gnd.n6448 585
R3761 gnd.n6446 gnd.n6403 585
R3762 gnd.n6444 gnd.n6443 585
R3763 gnd.n6442 gnd.n6404 585
R3764 gnd.n6441 gnd.n6440 585
R3765 gnd.n6438 gnd.n6405 585
R3766 gnd.n6436 gnd.n6435 585
R3767 gnd.n6434 gnd.n6406 585
R3768 gnd.n6433 gnd.n6432 585
R3769 gnd.n6430 gnd.n6428 585
R3770 gnd.n6427 gnd.n6130 585
R3771 gnd.n6564 gnd.n6563 585
R3772 gnd.n6565 gnd.n6564 585
R3773 gnd.n6374 gnd.n6131 585
R3774 gnd.n6131 gnd.n728 585
R3775 gnd.n6373 gnd.n6372 585
R3776 gnd.n6372 gnd.n726 585
R3777 gnd.n6371 gnd.n6125 585
R3778 gnd.n6572 gnd.n6125 585
R3779 gnd.n6370 gnd.n6369 585
R3780 gnd.n6369 gnd.n735 585
R3781 gnd.n6368 gnd.n6133 585
R3782 gnd.n6368 gnd.n6367 585
R3783 gnd.n6356 gnd.n6134 585
R3784 gnd.n6136 gnd.n6134 585
R3785 gnd.n6357 gnd.n6142 585
R3786 gnd.n6142 gnd.n742 585
R3787 gnd.n6359 gnd.n6358 585
R3788 gnd.n6360 gnd.n6359 585
R3789 gnd.n6355 gnd.n6141 585
R3790 gnd.n6141 gnd.n750 585
R3791 gnd.n6354 gnd.n751 585
R3792 gnd.n6969 gnd.n751 585
R3793 gnd.n6353 gnd.n6352 585
R3794 gnd.n6352 gnd.n6351 585
R3795 gnd.n6144 gnd.n6143 585
R3796 gnd.n6144 gnd.n759 585
R3797 gnd.n6339 gnd.n6151 585
R3798 gnd.n6151 gnd.n757 585
R3799 gnd.n6341 gnd.n6340 585
R3800 gnd.n6342 gnd.n6341 585
R3801 gnd.n6338 gnd.n6150 585
R3802 gnd.n6150 gnd.n767 585
R3803 gnd.n6337 gnd.n6336 585
R3804 gnd.n6336 gnd.n765 585
R3805 gnd.n6335 gnd.n6152 585
R3806 gnd.n6335 gnd.n6334 585
R3807 gnd.n6321 gnd.n6153 585
R3808 gnd.n6153 gnd.n775 585
R3809 gnd.n6322 gnd.n6161 585
R3810 gnd.n6161 gnd.n773 585
R3811 gnd.n6324 gnd.n6323 585
R3812 gnd.n6325 gnd.n6324 585
R3813 gnd.n6320 gnd.n6160 585
R3814 gnd.n6160 gnd.n783 585
R3815 gnd.n6319 gnd.n6318 585
R3816 gnd.n6318 gnd.n781 585
R3817 gnd.n6317 gnd.n6162 585
R3818 gnd.n6317 gnd.n6316 585
R3819 gnd.n6303 gnd.n6163 585
R3820 gnd.n6163 gnd.n791 585
R3821 gnd.n6304 gnd.n6171 585
R3822 gnd.n6171 gnd.n789 585
R3823 gnd.n6306 gnd.n6305 585
R3824 gnd.n6307 gnd.n6306 585
R3825 gnd.n6302 gnd.n6170 585
R3826 gnd.n6170 gnd.n799 585
R3827 gnd.n6301 gnd.n6300 585
R3828 gnd.n6300 gnd.n797 585
R3829 gnd.n6299 gnd.n6172 585
R3830 gnd.n6299 gnd.n6298 585
R3831 gnd.n6285 gnd.n6173 585
R3832 gnd.n6175 gnd.n6173 585
R3833 gnd.n6286 gnd.n6182 585
R3834 gnd.n6182 gnd.n805 585
R3835 gnd.n6288 gnd.n6287 585
R3836 gnd.n6289 gnd.n6288 585
R3837 gnd.n6284 gnd.n6181 585
R3838 gnd.n6181 gnd.n814 585
R3839 gnd.n6283 gnd.n6282 585
R3840 gnd.n6282 gnd.n812 585
R3841 gnd.n6281 gnd.n6183 585
R3842 gnd.n6281 gnd.n6280 585
R3843 gnd.n6266 gnd.n6184 585
R3844 gnd.n6184 gnd.n822 585
R3845 gnd.n6267 gnd.n6190 585
R3846 gnd.n6190 gnd.n820 585
R3847 gnd.n6269 gnd.n6268 585
R3848 gnd.n6271 gnd.n6269 585
R3849 gnd.n6265 gnd.n6189 585
R3850 gnd.n6189 gnd.n830 585
R3851 gnd.n6264 gnd.n6263 585
R3852 gnd.n6263 gnd.n828 585
R3853 gnd.n6262 gnd.n6191 585
R3854 gnd.n6262 gnd.n6261 585
R3855 gnd.n6247 gnd.n6192 585
R3856 gnd.n6192 gnd.n838 585
R3857 gnd.n6248 gnd.n6199 585
R3858 gnd.n6199 gnd.n836 585
R3859 gnd.n6250 gnd.n6249 585
R3860 gnd.n6252 gnd.n6250 585
R3861 gnd.n6246 gnd.n6198 585
R3862 gnd.n6198 gnd.n846 585
R3863 gnd.n6245 gnd.n6244 585
R3864 gnd.n6244 gnd.n844 585
R3865 gnd.n6243 gnd.n6200 585
R3866 gnd.n6243 gnd.n6242 585
R3867 gnd.n6228 gnd.n6201 585
R3868 gnd.n6201 gnd.n854 585
R3869 gnd.n6229 gnd.n6208 585
R3870 gnd.n6208 gnd.n852 585
R3871 gnd.n6231 gnd.n6230 585
R3872 gnd.n6233 gnd.n6231 585
R3873 gnd.n6227 gnd.n6207 585
R3874 gnd.n6207 gnd.n862 585
R3875 gnd.n6226 gnd.n6225 585
R3876 gnd.n6225 gnd.n860 585
R3877 gnd.n6224 gnd.n6209 585
R3878 gnd.n6224 gnd.n6223 585
R3879 gnd.n6214 gnd.n6213 585
R3880 gnd.n6214 gnd.n870 585
R3881 gnd.n6212 gnd.n6210 585
R3882 gnd.n6210 gnd.n868 585
R3883 gnd.n6211 gnd.n899 585
R3884 gnd.n6821 gnd.n899 585
R3885 gnd.n891 gnd.n890 585
R3886 gnd.n891 gnd.n877 585
R3887 gnd.n6829 gnd.n6828 585
R3888 gnd.n6828 gnd.n6827 585
R3889 gnd.n6830 gnd.n888 585
R3890 gnd.n893 gnd.n888 585
R3891 gnd.n6832 gnd.n6831 585
R3892 gnd.n6833 gnd.n6832 585
R3893 gnd.n889 gnd.n887 585
R3894 gnd.n887 gnd.n883 585
R3895 gnd.n6038 gnd.n927 585
R3896 gnd.n6055 gnd.n927 585
R3897 gnd.n6042 gnd.n6041 585
R3898 gnd.n6041 gnd.n6040 585
R3899 gnd.n6043 gnd.n935 585
R3900 gnd.n935 gnd.n909 585
R3901 gnd.n6045 gnd.n6044 585
R3902 gnd.n6046 gnd.n6045 585
R3903 gnd.n6037 gnd.n934 585
R3904 gnd.n934 gnd.n933 585
R3905 gnd.n6036 gnd.n6035 585
R3906 gnd.n6035 gnd.n919 585
R3907 gnd.n6034 gnd.n936 585
R3908 gnd.n6034 gnd.n917 585
R3909 gnd.n6033 gnd.n938 585
R3910 gnd.n6033 gnd.n6032 585
R3911 gnd.n5939 gnd.n937 585
R3912 gnd.n939 gnd.n937 585
R3913 gnd.n5940 gnd.n945 585
R3914 gnd.n6022 gnd.n945 585
R3915 gnd.n5942 gnd.n5941 585
R3916 gnd.n5943 gnd.n5942 585
R3917 gnd.n5938 gnd.n5914 585
R3918 gnd.n5914 gnd.n955 585
R3919 gnd.n5937 gnd.n5936 585
R3920 gnd.n5936 gnd.n953 585
R3921 gnd.n5935 gnd.n5915 585
R3922 gnd.n5935 gnd.n5934 585
R3923 gnd.n5923 gnd.n5922 585
R3924 gnd.n5923 gnd.n965 585
R3925 gnd.n5921 gnd.n5916 585
R3926 gnd.n5916 gnd.n963 585
R3927 gnd.n5920 gnd.n1001 585
R3928 gnd.n5963 gnd.n1001 585
R3929 gnd.n5919 gnd.n5918 585
R3930 gnd.n5918 gnd.n973 585
R3931 gnd.n5917 gnd.n994 585
R3932 gnd.n994 gnd.n971 585
R3933 gnd.n5971 gnd.n995 585
R3934 gnd.n5971 gnd.n5970 585
R3935 gnd.n5972 gnd.n993 585
R3936 gnd.n5972 gnd.n981 585
R3937 gnd.n5974 gnd.n5973 585
R3938 gnd.n5973 gnd.n979 585
R3939 gnd.n5975 gnd.n991 585
R3940 gnd.n5387 gnd.n991 585
R3941 gnd.n5977 gnd.n5976 585
R3942 gnd.n5978 gnd.n5977 585
R3943 gnd.n992 gnd.n990 585
R3944 gnd.n1011 gnd.n990 585
R3945 gnd.n5609 gnd.n5395 585
R3946 gnd.n5395 gnd.n1010 585
R3947 gnd.n5611 gnd.n5610 585
R3948 gnd.n5613 gnd.n5611 585
R3949 gnd.n5608 gnd.n5394 585
R3950 gnd.n5394 gnd.n1020 585
R3951 gnd.n5607 gnd.n5606 585
R3952 gnd.n5606 gnd.n1018 585
R3953 gnd.n5605 gnd.n5378 585
R3954 gnd.n5620 gnd.n5378 585
R3955 gnd.n5604 gnd.n5603 585
R3956 gnd.n5603 gnd.n1028 585
R3957 gnd.n5602 gnd.n5396 585
R3958 gnd.n5602 gnd.n5601 585
R3959 gnd.n5462 gnd.n5397 585
R3960 gnd.n5400 gnd.n5397 585
R3961 gnd.n5464 gnd.n5463 585
R3962 gnd.n5464 gnd.n1035 585
R3963 gnd.n3057 gnd.n1658 585
R3964 gnd.n1658 gnd.n1392 585
R3965 gnd.n7563 gnd.n7562 585
R3966 gnd.n7564 gnd.n7563 585
R3967 gnd.n7559 gnd.n336 585
R3968 gnd.n345 gnd.n336 585
R3969 gnd.n7558 gnd.n7557 585
R3970 gnd.n7557 gnd.n7556 585
R3971 gnd.n342 gnd.n341 585
R3972 gnd.n7548 gnd.n342 585
R3973 gnd.n7365 gnd.n7364 585
R3974 gnd.n7364 gnd.n348 585
R3975 gnd.n7366 gnd.n7359 585
R3976 gnd.n7359 gnd.n314 585
R3977 gnd.n7368 gnd.n7367 585
R3978 gnd.n7368 gnd.n311 585
R3979 gnd.n7369 gnd.n7358 585
R3980 gnd.n7369 gnd.n356 585
R3981 gnd.n7371 gnd.n7370 585
R3982 gnd.n7370 gnd.n364 585
R3983 gnd.n7372 gnd.n7353 585
R3984 gnd.n7353 gnd.n362 585
R3985 gnd.n7374 gnd.n7373 585
R3986 gnd.n7374 gnd.n383 585
R3987 gnd.n7375 gnd.n7352 585
R3988 gnd.n7375 gnd.n376 585
R3989 gnd.n7377 gnd.n7376 585
R3990 gnd.n7376 gnd.n373 585
R3991 gnd.n7378 gnd.n416 585
R3992 gnd.n416 gnd.n390 585
R3993 gnd.n7380 gnd.n7379 585
R3994 gnd.n7381 gnd.n7380 585
R3995 gnd.n417 gnd.n415 585
R3996 gnd.n415 gnd.n396 585
R3997 gnd.n7346 gnd.n7345 585
R3998 gnd.n7345 gnd.n408 585
R3999 gnd.n7344 gnd.n419 585
R4000 gnd.n7344 gnd.n405 585
R4001 gnd.n7343 gnd.n421 585
R4002 gnd.n7343 gnd.n7342 585
R4003 gnd.n7117 gnd.n420 585
R4004 gnd.n432 gnd.n420 585
R4005 gnd.n7118 gnd.n7111 585
R4006 gnd.n7111 gnd.n430 585
R4007 gnd.n7120 gnd.n7119 585
R4008 gnd.n7120 gnd.n443 585
R4009 gnd.n7121 gnd.n7110 585
R4010 gnd.n7121 gnd.n440 585
R4011 gnd.n7123 gnd.n7122 585
R4012 gnd.n7122 gnd.n454 585
R4013 gnd.n7124 gnd.n622 585
R4014 gnd.n622 gnd.n451 585
R4015 gnd.n7126 gnd.n7125 585
R4016 gnd.n7127 gnd.n7126 585
R4017 gnd.n623 gnd.n621 585
R4018 gnd.n621 gnd.n460 585
R4019 gnd.n7104 gnd.n7103 585
R4020 gnd.n7103 gnd.n471 585
R4021 gnd.n7102 gnd.n625 585
R4022 gnd.n7102 gnd.n468 585
R4023 gnd.n7101 gnd.n7100 585
R4024 gnd.n7101 gnd.n480 585
R4025 gnd.n627 gnd.n626 585
R4026 gnd.n626 gnd.n477 585
R4027 gnd.n7096 gnd.n7095 585
R4028 gnd.n7095 gnd.n489 585
R4029 gnd.n7094 gnd.n629 585
R4030 gnd.n7094 gnd.n486 585
R4031 gnd.n7093 gnd.n7092 585
R4032 gnd.n7093 gnd.n498 585
R4033 gnd.n631 gnd.n630 585
R4034 gnd.n630 gnd.n495 585
R4035 gnd.n7088 gnd.n7087 585
R4036 gnd.n7087 gnd.n581 585
R4037 gnd.n7086 gnd.n633 585
R4038 gnd.n7086 gnd.n532 585
R4039 gnd.n7085 gnd.n7084 585
R4040 gnd.n7085 gnd.n504 585
R4041 gnd.n635 gnd.n634 585
R4042 gnd.n7077 gnd.n634 585
R4043 gnd.n7080 gnd.n7079 585
R4044 gnd.n7079 gnd.n7078 585
R4045 gnd.n638 gnd.n637 585
R4046 gnd.n639 gnd.n638 585
R4047 gnd.n7065 gnd.n664 585
R4048 gnd.n664 gnd.n662 585
R4049 gnd.n7067 gnd.n7066 585
R4050 gnd.n7068 gnd.n7067 585
R4051 gnd.n665 gnd.n663 585
R4052 gnd.n671 gnd.n663 585
R4053 gnd.n7060 gnd.n7059 585
R4054 gnd.n7059 gnd.n7058 585
R4055 gnd.n668 gnd.n667 585
R4056 gnd.n669 gnd.n668 585
R4057 gnd.n7048 gnd.n7047 585
R4058 gnd.n7049 gnd.n7048 585
R4059 gnd.n680 gnd.n679 585
R4060 gnd.n679 gnd.n677 585
R4061 gnd.n7043 gnd.n7042 585
R4062 gnd.n7042 gnd.n7041 585
R4063 gnd.n683 gnd.n682 585
R4064 gnd.n684 gnd.n683 585
R4065 gnd.n7032 gnd.n7031 585
R4066 gnd.n7033 gnd.n7032 585
R4067 gnd.n694 gnd.n693 585
R4068 gnd.n693 gnd.n691 585
R4069 gnd.n7027 gnd.n7026 585
R4070 gnd.n7026 gnd.n7025 585
R4071 gnd.n697 gnd.n696 585
R4072 gnd.n706 gnd.n697 585
R4073 gnd.n7016 gnd.n7015 585
R4074 gnd.n7017 gnd.n7016 585
R4075 gnd.n708 gnd.n707 585
R4076 gnd.n707 gnd.n704 585
R4077 gnd.n7011 gnd.n7010 585
R4078 gnd.n7010 gnd.n7009 585
R4079 gnd.n711 gnd.n710 585
R4080 gnd.n6578 gnd.n711 585
R4081 gnd.n7000 gnd.n6999 585
R4082 gnd.n7001 gnd.n7000 585
R4083 gnd.n722 gnd.n721 585
R4084 gnd.n721 gnd.n718 585
R4085 gnd.n6995 gnd.n6994 585
R4086 gnd.n6994 gnd.n6993 585
R4087 gnd.n725 gnd.n724 585
R4088 gnd.n6573 gnd.n725 585
R4089 gnd.n6984 gnd.n6983 585
R4090 gnd.n6985 gnd.n6984 585
R4091 gnd.n737 gnd.n736 585
R4092 gnd.n6135 gnd.n736 585
R4093 gnd.n6979 gnd.n6978 585
R4094 gnd.n6978 gnd.n6977 585
R4095 gnd.n740 gnd.n739 585
R4096 gnd.n6140 gnd.n740 585
R4097 gnd.n6968 gnd.n6967 585
R4098 gnd.n6969 gnd.n6968 585
R4099 gnd.n753 gnd.n752 585
R4100 gnd.n6145 gnd.n752 585
R4101 gnd.n6963 gnd.n6962 585
R4102 gnd.n6962 gnd.n6961 585
R4103 gnd.n756 gnd.n755 585
R4104 gnd.n6149 gnd.n756 585
R4105 gnd.n6952 gnd.n6951 585
R4106 gnd.n6953 gnd.n6952 585
R4107 gnd.n769 gnd.n768 585
R4108 gnd.n6154 gnd.n768 585
R4109 gnd.n6947 gnd.n6946 585
R4110 gnd.n6946 gnd.n6945 585
R4111 gnd.n772 gnd.n771 585
R4112 gnd.n6159 gnd.n772 585
R4113 gnd.n6936 gnd.n6935 585
R4114 gnd.n6937 gnd.n6936 585
R4115 gnd.n785 gnd.n784 585
R4116 gnd.n6164 gnd.n784 585
R4117 gnd.n6931 gnd.n6930 585
R4118 gnd.n6930 gnd.n6929 585
R4119 gnd.n788 gnd.n787 585
R4120 gnd.n6169 gnd.n788 585
R4121 gnd.n6920 gnd.n6919 585
R4122 gnd.n6921 gnd.n6920 585
R4123 gnd.n801 gnd.n800 585
R4124 gnd.n6174 gnd.n800 585
R4125 gnd.n6915 gnd.n6914 585
R4126 gnd.n6914 gnd.n6913 585
R4127 gnd.n804 gnd.n803 585
R4128 gnd.n6180 gnd.n804 585
R4129 gnd.n6904 gnd.n6903 585
R4130 gnd.n6905 gnd.n6904 585
R4131 gnd.n816 gnd.n815 585
R4132 gnd.n6280 gnd.n815 585
R4133 gnd.n6899 gnd.n6898 585
R4134 gnd.n6898 gnd.n6897 585
R4135 gnd.n819 gnd.n818 585
R4136 gnd.n6270 gnd.n819 585
R4137 gnd.n6888 gnd.n6887 585
R4138 gnd.n6889 gnd.n6888 585
R4139 gnd.n832 gnd.n831 585
R4140 gnd.n6193 gnd.n831 585
R4141 gnd.n6883 gnd.n6882 585
R4142 gnd.n6882 gnd.n6881 585
R4143 gnd.n835 gnd.n834 585
R4144 gnd.n6251 gnd.n835 585
R4145 gnd.n6872 gnd.n6871 585
R4146 gnd.n6873 gnd.n6872 585
R4147 gnd.n848 gnd.n847 585
R4148 gnd.n6202 gnd.n847 585
R4149 gnd.n6867 gnd.n6866 585
R4150 gnd.n6866 gnd.n6865 585
R4151 gnd.n851 gnd.n850 585
R4152 gnd.n6232 gnd.n851 585
R4153 gnd.n6856 gnd.n6855 585
R4154 gnd.n6857 gnd.n6856 585
R4155 gnd.n864 gnd.n863 585
R4156 gnd.n6215 gnd.n863 585
R4157 gnd.n6851 gnd.n6850 585
R4158 gnd.n6850 gnd.n6849 585
R4159 gnd.n867 gnd.n866 585
R4160 gnd.n6820 gnd.n867 585
R4161 gnd.n6840 gnd.n6839 585
R4162 gnd.n6841 gnd.n6840 585
R4163 gnd.n879 gnd.n878 585
R4164 gnd.n892 gnd.n878 585
R4165 gnd.n6835 gnd.n6834 585
R4166 gnd.n6834 gnd.n6833 585
R4167 gnd.n882 gnd.n881 585
R4168 gnd.n6056 gnd.n882 585
R4169 gnd.n6076 gnd.n912 585
R4170 gnd.n6039 gnd.n912 585
R4171 gnd.n6078 gnd.n6077 585
R4172 gnd.n6079 gnd.n6078 585
R4173 gnd.n913 gnd.n911 585
R4174 gnd.n932 gnd.n911 585
R4175 gnd.n6071 gnd.n6070 585
R4176 gnd.n6070 gnd.n6069 585
R4177 gnd.n916 gnd.n915 585
R4178 gnd.n940 gnd.n916 585
R4179 gnd.n6020 gnd.n6019 585
R4180 gnd.n6021 gnd.n6020 585
R4181 gnd.n949 gnd.n948 585
R4182 gnd.n5944 gnd.n948 585
R4183 gnd.n6015 gnd.n6014 585
R4184 gnd.n6014 gnd.n6013 585
R4185 gnd.n952 gnd.n951 585
R4186 gnd.n5924 gnd.n952 585
R4187 gnd.n6001 gnd.n6000 585
R4188 gnd.n6002 gnd.n6001 585
R4189 gnd.n967 gnd.n966 585
R4190 gnd.n5962 gnd.n966 585
R4191 gnd.n5996 gnd.n5995 585
R4192 gnd.n5995 gnd.n5994 585
R4193 gnd.n970 gnd.n969 585
R4194 gnd.n5907 gnd.n970 585
R4195 gnd.n5985 gnd.n5984 585
R4196 gnd.n5986 gnd.n5985 585
R4197 gnd.n983 gnd.n982 585
R4198 gnd.n5386 gnd.n982 585
R4199 gnd.n5980 gnd.n5979 585
R4200 gnd.n5979 gnd.n5978 585
R4201 gnd.n986 gnd.n985 585
R4202 gnd.n5899 gnd.n986 585
R4203 gnd.n5887 gnd.n1022 585
R4204 gnd.n5612 gnd.n1022 585
R4205 gnd.n5889 gnd.n5888 585
R4206 gnd.n5890 gnd.n5889 585
R4207 gnd.n1023 gnd.n1021 585
R4208 gnd.n5621 gnd.n1021 585
R4209 gnd.n5882 gnd.n5881 585
R4210 gnd.n5881 gnd.n5880 585
R4211 gnd.n1026 gnd.n1025 585
R4212 gnd.n5399 gnd.n1026 585
R4213 gnd.n5871 gnd.n5870 585
R4214 gnd.n5872 gnd.n5871 585
R4215 gnd.n1037 gnd.n1036 585
R4216 gnd.n5374 gnd.n1036 585
R4217 gnd.n5866 gnd.n5865 585
R4218 gnd.n5865 gnd.n5864 585
R4219 gnd.n1040 gnd.n1039 585
R4220 gnd.n1050 gnd.n1040 585
R4221 gnd.n5855 gnd.n5854 585
R4222 gnd.n5856 gnd.n5855 585
R4223 gnd.n1052 gnd.n1051 585
R4224 gnd.n1051 gnd.n1048 585
R4225 gnd.n5850 gnd.n5849 585
R4226 gnd.n5849 gnd.n5848 585
R4227 gnd.n1055 gnd.n1054 585
R4228 gnd.n1064 gnd.n1055 585
R4229 gnd.n5839 gnd.n5838 585
R4230 gnd.n5840 gnd.n5839 585
R4231 gnd.n1066 gnd.n1065 585
R4232 gnd.n1065 gnd.n1062 585
R4233 gnd.n5834 gnd.n5833 585
R4234 gnd.n5833 gnd.n5832 585
R4235 gnd.n1069 gnd.n1068 585
R4236 gnd.n1070 gnd.n1069 585
R4237 gnd.n5823 gnd.n5822 585
R4238 gnd.n5824 gnd.n5823 585
R4239 gnd.n1080 gnd.n1079 585
R4240 gnd.n1079 gnd.n1077 585
R4241 gnd.n5818 gnd.n5817 585
R4242 gnd.n5817 gnd.n5816 585
R4243 gnd.n1083 gnd.n1082 585
R4244 gnd.n1084 gnd.n1083 585
R4245 gnd.n5807 gnd.n5806 585
R4246 gnd.n5808 gnd.n5807 585
R4247 gnd.n1093 gnd.n1092 585
R4248 gnd.n1099 gnd.n1092 585
R4249 gnd.n5802 gnd.n5801 585
R4250 gnd.n5801 gnd.n5800 585
R4251 gnd.n1096 gnd.n1095 585
R4252 gnd.n1097 gnd.n1096 585
R4253 gnd.n5071 gnd.n5070 585
R4254 gnd.n5070 gnd.n1104 585
R4255 gnd.n5072 gnd.n5065 585
R4256 gnd.n5074 gnd.n5065 585
R4257 gnd.n5076 gnd.n5073 585
R4258 gnd.n5076 gnd.n5075 585
R4259 gnd.n5078 gnd.n5064 585
R4260 gnd.n5078 gnd.n5077 585
R4261 gnd.n5080 gnd.n5079 585
R4262 gnd.n5079 gnd.n1177 585
R4263 gnd.n5081 gnd.n5059 585
R4264 gnd.n5059 gnd.n1175 585
R4265 gnd.n5083 gnd.n5082 585
R4266 gnd.n5083 gnd.n1265 585
R4267 gnd.n5084 gnd.n5058 585
R4268 gnd.n5084 gnd.n1274 585
R4269 gnd.n5086 gnd.n5085 585
R4270 gnd.n5085 gnd.n1271 585
R4271 gnd.n5087 gnd.n5053 585
R4272 gnd.n5053 gnd.n1284 585
R4273 gnd.n5089 gnd.n5088 585
R4274 gnd.n5089 gnd.n1281 585
R4275 gnd.n5090 gnd.n5052 585
R4276 gnd.n5090 gnd.n1293 585
R4277 gnd.n5092 gnd.n5091 585
R4278 gnd.n5091 gnd.n1290 585
R4279 gnd.n5093 gnd.n4945 585
R4280 gnd.n4945 gnd.n1301 585
R4281 gnd.n5095 gnd.n5094 585
R4282 gnd.n5096 gnd.n5095 585
R4283 gnd.n4946 gnd.n4944 585
R4284 gnd.n4944 gnd.n1310 585
R4285 gnd.n5046 gnd.n5045 585
R4286 gnd.n5045 gnd.n1307 585
R4287 gnd.n5044 gnd.n4948 585
R4288 gnd.n5044 gnd.n1319 585
R4289 gnd.n5043 gnd.n5042 585
R4290 gnd.n5043 gnd.n1316 585
R4291 gnd.n4950 gnd.n4949 585
R4292 gnd.n4949 gnd.n1328 585
R4293 gnd.n5038 gnd.n5037 585
R4294 gnd.n5037 gnd.n1325 585
R4295 gnd.n5036 gnd.n4952 585
R4296 gnd.n5036 gnd.n1336 585
R4297 gnd.n5035 gnd.n4954 585
R4298 gnd.n5035 gnd.n5034 585
R4299 gnd.n4980 gnd.n4953 585
R4300 gnd.n4953 gnd.n1345 585
R4301 gnd.n4982 gnd.n4981 585
R4302 gnd.n4981 gnd.n1342 585
R4303 gnd.n4983 gnd.n4973 585
R4304 gnd.n4973 gnd.n1354 585
R4305 gnd.n4985 gnd.n4984 585
R4306 gnd.n4985 gnd.n1351 585
R4307 gnd.n4986 gnd.n4972 585
R4308 gnd.n4986 gnd.n1363 585
R4309 gnd.n4988 gnd.n4987 585
R4310 gnd.n4987 gnd.n1360 585
R4311 gnd.n4989 gnd.n4962 585
R4312 gnd.n4962 gnd.n1371 585
R4313 gnd.n4991 gnd.n4990 585
R4314 gnd.n4992 gnd.n4991 585
R4315 gnd.n4963 gnd.n4961 585
R4316 gnd.n4961 gnd.n1380 585
R4317 gnd.n4966 gnd.n4965 585
R4318 gnd.n4965 gnd.n1377 585
R4319 gnd.n1420 gnd.n1419 585
R4320 gnd.n1425 gnd.n1420 585
R4321 gnd.n5222 gnd.n5221 585
R4322 gnd.n5221 gnd.n5220 585
R4323 gnd.n5223 gnd.n1414 585
R4324 gnd.n1421 gnd.n1414 585
R4325 gnd.n5225 gnd.n5224 585
R4326 gnd.n5226 gnd.n5225 585
R4327 gnd.n1415 gnd.n1413 585
R4328 gnd.n1413 gnd.n1406 585
R4329 gnd.n3054 gnd.n3053 585
R4330 gnd.n3053 gnd.n3052 585
R4331 gnd.n6734 gnd.n6733 585
R4332 gnd.n6733 gnd.n662 585
R4333 gnd.n6735 gnd.n661 585
R4334 gnd.n7068 gnd.n661 585
R4335 gnd.n6736 gnd.n6594 585
R4336 gnd.n6594 gnd.n671 585
R4337 gnd.n6592 gnd.n670 585
R4338 gnd.n7058 gnd.n670 585
R4339 gnd.n6740 gnd.n6591 585
R4340 gnd.n6591 gnd.n669 585
R4341 gnd.n6741 gnd.n678 585
R4342 gnd.n7049 gnd.n678 585
R4343 gnd.n6742 gnd.n6590 585
R4344 gnd.n6590 gnd.n677 585
R4345 gnd.n6588 gnd.n685 585
R4346 gnd.n7041 gnd.n685 585
R4347 gnd.n6746 gnd.n6587 585
R4348 gnd.n6587 gnd.n684 585
R4349 gnd.n6747 gnd.n692 585
R4350 gnd.n7033 gnd.n692 585
R4351 gnd.n6748 gnd.n6586 585
R4352 gnd.n6586 gnd.n691 585
R4353 gnd.n6584 gnd.n698 585
R4354 gnd.n7025 gnd.n698 585
R4355 gnd.n6752 gnd.n6583 585
R4356 gnd.n6583 gnd.n706 585
R4357 gnd.n6753 gnd.n705 585
R4358 gnd.n7017 gnd.n705 585
R4359 gnd.n6754 gnd.n6582 585
R4360 gnd.n6582 gnd.n704 585
R4361 gnd.n6580 gnd.n712 585
R4362 gnd.n7009 gnd.n712 585
R4363 gnd.n6758 gnd.n6579 585
R4364 gnd.n6579 gnd.n6578 585
R4365 gnd.n6759 gnd.n719 585
R4366 gnd.n7001 gnd.n719 585
R4367 gnd.n6760 gnd.n6577 585
R4368 gnd.n6577 gnd.n718 585
R4369 gnd.n6575 gnd.n727 585
R4370 gnd.n6993 gnd.n727 585
R4371 gnd.n6764 gnd.n6574 585
R4372 gnd.n6574 gnd.n6573 585
R4373 gnd.n6765 gnd.n734 585
R4374 gnd.n6985 gnd.n734 585
R4375 gnd.n6766 gnd.n6124 585
R4376 gnd.n6135 gnd.n6124 585
R4377 gnd.n6122 gnd.n741 585
R4378 gnd.n6977 gnd.n741 585
R4379 gnd.n6770 gnd.n6121 585
R4380 gnd.n6140 gnd.n6121 585
R4381 gnd.n6771 gnd.n749 585
R4382 gnd.n6969 gnd.n749 585
R4383 gnd.n6772 gnd.n6120 585
R4384 gnd.n6145 gnd.n6120 585
R4385 gnd.n6118 gnd.n758 585
R4386 gnd.n6961 gnd.n758 585
R4387 gnd.n6776 gnd.n6117 585
R4388 gnd.n6149 gnd.n6117 585
R4389 gnd.n6777 gnd.n766 585
R4390 gnd.n6953 gnd.n766 585
R4391 gnd.n6778 gnd.n6116 585
R4392 gnd.n6154 gnd.n6116 585
R4393 gnd.n6114 gnd.n774 585
R4394 gnd.n6945 gnd.n774 585
R4395 gnd.n6782 gnd.n6113 585
R4396 gnd.n6159 gnd.n6113 585
R4397 gnd.n6783 gnd.n782 585
R4398 gnd.n6937 gnd.n782 585
R4399 gnd.n6784 gnd.n6112 585
R4400 gnd.n6164 gnd.n6112 585
R4401 gnd.n6110 gnd.n790 585
R4402 gnd.n6929 gnd.n790 585
R4403 gnd.n6788 gnd.n6109 585
R4404 gnd.n6169 gnd.n6109 585
R4405 gnd.n6789 gnd.n798 585
R4406 gnd.n6921 gnd.n798 585
R4407 gnd.n6790 gnd.n6108 585
R4408 gnd.n6174 gnd.n6108 585
R4409 gnd.n6106 gnd.n806 585
R4410 gnd.n6913 gnd.n806 585
R4411 gnd.n6794 gnd.n6105 585
R4412 gnd.n6180 gnd.n6105 585
R4413 gnd.n6795 gnd.n813 585
R4414 gnd.n6905 gnd.n813 585
R4415 gnd.n6796 gnd.n6104 585
R4416 gnd.n6280 gnd.n6104 585
R4417 gnd.n6102 gnd.n821 585
R4418 gnd.n6897 gnd.n821 585
R4419 gnd.n6800 gnd.n6101 585
R4420 gnd.n6270 gnd.n6101 585
R4421 gnd.n6801 gnd.n829 585
R4422 gnd.n6889 gnd.n829 585
R4423 gnd.n6802 gnd.n6100 585
R4424 gnd.n6193 gnd.n6100 585
R4425 gnd.n6098 gnd.n837 585
R4426 gnd.n6881 gnd.n837 585
R4427 gnd.n6806 gnd.n6097 585
R4428 gnd.n6251 gnd.n6097 585
R4429 gnd.n6807 gnd.n845 585
R4430 gnd.n6873 gnd.n845 585
R4431 gnd.n6808 gnd.n6096 585
R4432 gnd.n6202 gnd.n6096 585
R4433 gnd.n6094 gnd.n853 585
R4434 gnd.n6865 gnd.n853 585
R4435 gnd.n6812 gnd.n6093 585
R4436 gnd.n6232 gnd.n6093 585
R4437 gnd.n6813 gnd.n861 585
R4438 gnd.n6857 gnd.n861 585
R4439 gnd.n6814 gnd.n6092 585
R4440 gnd.n6215 gnd.n6092 585
R4441 gnd.n901 gnd.n869 585
R4442 gnd.n6849 gnd.n869 585
R4443 gnd.n6819 gnd.n6818 585
R4444 gnd.n6820 gnd.n6819 585
R4445 gnd.n900 gnd.n876 585
R4446 gnd.n6841 gnd.n876 585
R4447 gnd.n6088 gnd.n6087 585
R4448 gnd.n6087 gnd.n892 585
R4449 gnd.n6086 gnd.n885 585
R4450 gnd.n6833 gnd.n885 585
R4451 gnd.n6085 gnd.n904 585
R4452 gnd.n6056 gnd.n904 585
R4453 gnd.n908 gnd.n903 585
R4454 gnd.n6039 gnd.n908 585
R4455 gnd.n6081 gnd.n6080 585
R4456 gnd.n6080 gnd.n6079 585
R4457 gnd.n907 gnd.n906 585
R4458 gnd.n932 gnd.n907 585
R4459 gnd.n5949 gnd.n918 585
R4460 gnd.n6069 gnd.n918 585
R4461 gnd.n5950 gnd.n5948 585
R4462 gnd.n5948 gnd.n940 585
R4463 gnd.n5946 gnd.n946 585
R4464 gnd.n6021 gnd.n946 585
R4465 gnd.n5954 gnd.n5945 585
R4466 gnd.n5945 gnd.n5944 585
R4467 gnd.n5955 gnd.n954 585
R4468 gnd.n6013 gnd.n954 585
R4469 gnd.n5956 gnd.n5913 585
R4470 gnd.n5924 gnd.n5913 585
R4471 gnd.n1003 gnd.n964 585
R4472 gnd.n6002 gnd.n964 585
R4473 gnd.n5961 gnd.n5960 585
R4474 gnd.n5962 gnd.n5961 585
R4475 gnd.n1002 gnd.n972 585
R4476 gnd.n5994 gnd.n972 585
R4477 gnd.n5909 gnd.n5908 585
R4478 gnd.n5908 gnd.n5907 585
R4479 gnd.n5906 gnd.n980 585
R4480 gnd.n5986 gnd.n980 585
R4481 gnd.n5905 gnd.n1006 585
R4482 gnd.n5386 gnd.n1006 585
R4483 gnd.n1005 gnd.n988 585
R4484 gnd.n5978 gnd.n988 585
R4485 gnd.n5901 gnd.n5900 585
R4486 gnd.n5900 gnd.n5899 585
R4487 gnd.n1009 gnd.n1008 585
R4488 gnd.n5612 gnd.n1009 585
R4489 gnd.n5624 gnd.n1019 585
R4490 gnd.n5890 gnd.n1019 585
R4491 gnd.n5625 gnd.n5622 585
R4492 gnd.n5622 gnd.n5621 585
R4493 gnd.n5626 gnd.n1027 585
R4494 gnd.n5880 gnd.n1027 585
R4495 gnd.n5398 gnd.n5376 585
R4496 gnd.n5399 gnd.n5398 585
R4497 gnd.n5630 gnd.n1034 585
R4498 gnd.n5872 gnd.n1034 585
R4499 gnd.n5631 gnd.n5375 585
R4500 gnd.n5375 gnd.n5374 585
R4501 gnd.n5632 gnd.n1041 585
R4502 gnd.n5864 gnd.n1041 585
R4503 gnd.n5372 gnd.n5371 585
R4504 gnd.n5371 gnd.n1050 585
R4505 gnd.n5636 gnd.n1049 585
R4506 gnd.n5856 gnd.n1049 585
R4507 gnd.n5637 gnd.n5370 585
R4508 gnd.n5370 gnd.n1048 585
R4509 gnd.n5638 gnd.n1056 585
R4510 gnd.n5848 gnd.n1056 585
R4511 gnd.n5368 gnd.n5367 585
R4512 gnd.n5367 gnd.n1064 585
R4513 gnd.n5642 gnd.n1063 585
R4514 gnd.n5840 gnd.n1063 585
R4515 gnd.n5643 gnd.n5366 585
R4516 gnd.n5366 gnd.n1062 585
R4517 gnd.n5644 gnd.n1071 585
R4518 gnd.n5832 gnd.n1071 585
R4519 gnd.n5364 gnd.n5363 585
R4520 gnd.n5363 gnd.n1070 585
R4521 gnd.n5648 gnd.n1078 585
R4522 gnd.n5824 gnd.n1078 585
R4523 gnd.n5649 gnd.n5362 585
R4524 gnd.n5362 gnd.n1077 585
R4525 gnd.n5650 gnd.n1085 585
R4526 gnd.n5816 gnd.n1085 585
R4527 gnd.n5360 gnd.n5359 585
R4528 gnd.n5359 gnd.n1084 585
R4529 gnd.n5654 gnd.n1091 585
R4530 gnd.n5808 gnd.n1091 585
R4531 gnd.n5655 gnd.n5358 585
R4532 gnd.n5358 gnd.n1099 585
R4533 gnd.n5656 gnd.n1098 585
R4534 gnd.n5800 gnd.n1098 585
R4535 gnd.n5789 gnd.n5788 585
R4536 gnd.n5787 gnd.n1118 585
R4537 gnd.n1120 gnd.n1117 585
R4538 gnd.n5791 gnd.n1117 585
R4539 gnd.n5780 gnd.n1128 585
R4540 gnd.n5779 gnd.n1129 585
R4541 gnd.n1131 gnd.n1130 585
R4542 gnd.n5772 gnd.n1137 585
R4543 gnd.n5771 gnd.n1138 585
R4544 gnd.n1145 gnd.n1139 585
R4545 gnd.n5764 gnd.n1146 585
R4546 gnd.n5763 gnd.n1147 585
R4547 gnd.n1149 gnd.n1148 585
R4548 gnd.n5756 gnd.n1155 585
R4549 gnd.n5755 gnd.n1156 585
R4550 gnd.n1165 gnd.n1157 585
R4551 gnd.n5748 gnd.n1166 585
R4552 gnd.n5747 gnd.n1167 585
R4553 gnd.n1169 gnd.n1168 585
R4554 gnd.n5147 gnd.n5122 585
R4555 gnd.n5146 gnd.n5123 585
R4556 gnd.n5145 gnd.n5124 585
R4557 gnd.n5126 gnd.n5125 585
R4558 gnd.n5141 gnd.n5128 585
R4559 gnd.n5140 gnd.n5129 585
R4560 gnd.n5139 gnd.n5130 585
R4561 gnd.n5136 gnd.n5135 585
R4562 gnd.n1103 gnd.n1102 585
R4563 gnd.n5794 gnd.n5793 585
R4564 gnd.n5795 gnd.n1100 585
R4565 gnd.n7071 gnd.n655 585
R4566 gnd.n662 gnd.n655 585
R4567 gnd.n7070 gnd.n7069 585
R4568 gnd.n7069 gnd.n7068 585
R4569 gnd.n660 gnd.n659 585
R4570 gnd.n671 gnd.n660 585
R4571 gnd.n7057 gnd.n7056 585
R4572 gnd.n7058 gnd.n7057 585
R4573 gnd.n673 gnd.n672 585
R4574 gnd.n672 gnd.n669 585
R4575 gnd.n7051 gnd.n7050 585
R4576 gnd.n7050 gnd.n7049 585
R4577 gnd.n676 gnd.n675 585
R4578 gnd.n677 gnd.n676 585
R4579 gnd.n7040 gnd.n7039 585
R4580 gnd.n7041 gnd.n7040 585
R4581 gnd.n687 gnd.n686 585
R4582 gnd.n686 gnd.n684 585
R4583 gnd.n7035 gnd.n7034 585
R4584 gnd.n7034 gnd.n7033 585
R4585 gnd.n690 gnd.n689 585
R4586 gnd.n691 gnd.n690 585
R4587 gnd.n7024 gnd.n7023 585
R4588 gnd.n7025 gnd.n7024 585
R4589 gnd.n700 gnd.n699 585
R4590 gnd.n706 gnd.n699 585
R4591 gnd.n7019 gnd.n7018 585
R4592 gnd.n7018 gnd.n7017 585
R4593 gnd.n703 gnd.n702 585
R4594 gnd.n704 gnd.n703 585
R4595 gnd.n7008 gnd.n7007 585
R4596 gnd.n7009 gnd.n7008 585
R4597 gnd.n714 gnd.n713 585
R4598 gnd.n6578 gnd.n713 585
R4599 gnd.n7003 gnd.n7002 585
R4600 gnd.n7002 gnd.n7001 585
R4601 gnd.n717 gnd.n716 585
R4602 gnd.n718 gnd.n717 585
R4603 gnd.n6992 gnd.n6991 585
R4604 gnd.n6993 gnd.n6992 585
R4605 gnd.n730 gnd.n729 585
R4606 gnd.n6573 gnd.n729 585
R4607 gnd.n6987 gnd.n6986 585
R4608 gnd.n6986 gnd.n6985 585
R4609 gnd.n733 gnd.n732 585
R4610 gnd.n6135 gnd.n733 585
R4611 gnd.n6976 gnd.n6975 585
R4612 gnd.n6977 gnd.n6976 585
R4613 gnd.n744 gnd.n743 585
R4614 gnd.n6140 gnd.n743 585
R4615 gnd.n6971 gnd.n6970 585
R4616 gnd.n6970 gnd.n6969 585
R4617 gnd.n747 gnd.n746 585
R4618 gnd.n6145 gnd.n747 585
R4619 gnd.n6960 gnd.n6959 585
R4620 gnd.n6961 gnd.n6960 585
R4621 gnd.n761 gnd.n760 585
R4622 gnd.n6149 gnd.n760 585
R4623 gnd.n6955 gnd.n6954 585
R4624 gnd.n6954 gnd.n6953 585
R4625 gnd.n764 gnd.n763 585
R4626 gnd.n6154 gnd.n764 585
R4627 gnd.n6944 gnd.n6943 585
R4628 gnd.n6945 gnd.n6944 585
R4629 gnd.n777 gnd.n776 585
R4630 gnd.n6159 gnd.n776 585
R4631 gnd.n6939 gnd.n6938 585
R4632 gnd.n6938 gnd.n6937 585
R4633 gnd.n780 gnd.n779 585
R4634 gnd.n6164 gnd.n780 585
R4635 gnd.n6928 gnd.n6927 585
R4636 gnd.n6929 gnd.n6928 585
R4637 gnd.n793 gnd.n792 585
R4638 gnd.n6169 gnd.n792 585
R4639 gnd.n6923 gnd.n6922 585
R4640 gnd.n6922 gnd.n6921 585
R4641 gnd.n796 gnd.n795 585
R4642 gnd.n6174 gnd.n796 585
R4643 gnd.n6912 gnd.n6911 585
R4644 gnd.n6913 gnd.n6912 585
R4645 gnd.n808 gnd.n807 585
R4646 gnd.n6180 gnd.n807 585
R4647 gnd.n6907 gnd.n6906 585
R4648 gnd.n6906 gnd.n6905 585
R4649 gnd.n811 gnd.n810 585
R4650 gnd.n6280 gnd.n811 585
R4651 gnd.n6896 gnd.n6895 585
R4652 gnd.n6897 gnd.n6896 585
R4653 gnd.n824 gnd.n823 585
R4654 gnd.n6270 gnd.n823 585
R4655 gnd.n6891 gnd.n6890 585
R4656 gnd.n6890 gnd.n6889 585
R4657 gnd.n827 gnd.n826 585
R4658 gnd.n6193 gnd.n827 585
R4659 gnd.n6880 gnd.n6879 585
R4660 gnd.n6881 gnd.n6880 585
R4661 gnd.n840 gnd.n839 585
R4662 gnd.n6251 gnd.n839 585
R4663 gnd.n6875 gnd.n6874 585
R4664 gnd.n6874 gnd.n6873 585
R4665 gnd.n843 gnd.n842 585
R4666 gnd.n6202 gnd.n843 585
R4667 gnd.n6864 gnd.n6863 585
R4668 gnd.n6865 gnd.n6864 585
R4669 gnd.n856 gnd.n855 585
R4670 gnd.n6232 gnd.n855 585
R4671 gnd.n6859 gnd.n6858 585
R4672 gnd.n6858 gnd.n6857 585
R4673 gnd.n859 gnd.n858 585
R4674 gnd.n6215 gnd.n859 585
R4675 gnd.n6848 gnd.n6847 585
R4676 gnd.n6849 gnd.n6848 585
R4677 gnd.n872 gnd.n871 585
R4678 gnd.n6820 gnd.n871 585
R4679 gnd.n6843 gnd.n6842 585
R4680 gnd.n6842 gnd.n6841 585
R4681 gnd.n875 gnd.n874 585
R4682 gnd.n892 gnd.n875 585
R4683 gnd.n6058 gnd.n886 585
R4684 gnd.n6833 gnd.n886 585
R4685 gnd.n6061 gnd.n6057 585
R4686 gnd.n6057 gnd.n6056 585
R4687 gnd.n6062 gnd.n926 585
R4688 gnd.n6039 gnd.n926 585
R4689 gnd.n6063 gnd.n910 585
R4690 gnd.n6079 gnd.n910 585
R4691 gnd.n923 gnd.n921 585
R4692 gnd.n932 gnd.n921 585
R4693 gnd.n6068 gnd.n6067 585
R4694 gnd.n6069 gnd.n6068 585
R4695 gnd.n922 gnd.n920 585
R4696 gnd.n940 gnd.n920 585
R4697 gnd.n6007 gnd.n947 585
R4698 gnd.n6021 gnd.n947 585
R4699 gnd.n959 gnd.n957 585
R4700 gnd.n5944 gnd.n957 585
R4701 gnd.n6012 gnd.n6011 585
R4702 gnd.n6013 gnd.n6012 585
R4703 gnd.n958 gnd.n956 585
R4704 gnd.n5924 gnd.n956 585
R4705 gnd.n6004 gnd.n6003 585
R4706 gnd.n6003 gnd.n6002 585
R4707 gnd.n962 gnd.n961 585
R4708 gnd.n5962 gnd.n962 585
R4709 gnd.n5993 gnd.n5992 585
R4710 gnd.n5994 gnd.n5993 585
R4711 gnd.n975 gnd.n974 585
R4712 gnd.n5907 gnd.n974 585
R4713 gnd.n5988 gnd.n5987 585
R4714 gnd.n5987 gnd.n5986 585
R4715 gnd.n978 gnd.n977 585
R4716 gnd.n5386 gnd.n978 585
R4717 gnd.n1014 gnd.n989 585
R4718 gnd.n5978 gnd.n989 585
R4719 gnd.n5898 gnd.n5897 585
R4720 gnd.n5899 gnd.n5898 585
R4721 gnd.n1013 gnd.n1012 585
R4722 gnd.n5612 gnd.n1012 585
R4723 gnd.n5892 gnd.n5891 585
R4724 gnd.n5891 gnd.n5890 585
R4725 gnd.n1017 gnd.n1016 585
R4726 gnd.n5621 gnd.n1017 585
R4727 gnd.n5879 gnd.n5878 585
R4728 gnd.n5880 gnd.n5879 585
R4729 gnd.n1030 gnd.n1029 585
R4730 gnd.n5399 gnd.n1029 585
R4731 gnd.n5874 gnd.n5873 585
R4732 gnd.n5873 gnd.n5872 585
R4733 gnd.n1033 gnd.n1032 585
R4734 gnd.n5374 gnd.n1033 585
R4735 gnd.n5863 gnd.n5862 585
R4736 gnd.n5864 gnd.n5863 585
R4737 gnd.n1044 gnd.n1043 585
R4738 gnd.n1050 gnd.n1043 585
R4739 gnd.n5858 gnd.n5857 585
R4740 gnd.n5857 gnd.n5856 585
R4741 gnd.n1047 gnd.n1046 585
R4742 gnd.n1048 gnd.n1047 585
R4743 gnd.n5847 gnd.n5846 585
R4744 gnd.n5848 gnd.n5847 585
R4745 gnd.n1058 gnd.n1057 585
R4746 gnd.n1064 gnd.n1057 585
R4747 gnd.n5842 gnd.n5841 585
R4748 gnd.n5841 gnd.n5840 585
R4749 gnd.n1061 gnd.n1060 585
R4750 gnd.n1062 gnd.n1061 585
R4751 gnd.n5831 gnd.n5830 585
R4752 gnd.n5832 gnd.n5831 585
R4753 gnd.n1073 gnd.n1072 585
R4754 gnd.n1072 gnd.n1070 585
R4755 gnd.n5826 gnd.n5825 585
R4756 gnd.n5825 gnd.n5824 585
R4757 gnd.n1076 gnd.n1075 585
R4758 gnd.n1077 gnd.n1076 585
R4759 gnd.n5815 gnd.n5814 585
R4760 gnd.n5816 gnd.n5815 585
R4761 gnd.n1087 gnd.n1086 585
R4762 gnd.n1086 gnd.n1084 585
R4763 gnd.n5810 gnd.n5809 585
R4764 gnd.n5809 gnd.n5808 585
R4765 gnd.n1090 gnd.n1089 585
R4766 gnd.n1099 gnd.n1090 585
R4767 gnd.n5799 gnd.n5798 585
R4768 gnd.n5800 gnd.n5799 585
R4769 gnd.n7075 gnd.n7074 585
R4770 gnd.n7076 gnd.n7075 585
R4771 gnd.n656 gnd.n654 585
R4772 gnd.n6668 gnd.n6667 585
R4773 gnd.n6669 gnd.n6666 585
R4774 gnd.n6661 gnd.n6660 585
R4775 gnd.n6673 gnd.n6659 585
R4776 gnd.n6674 gnd.n6658 585
R4777 gnd.n6675 gnd.n6657 585
R4778 gnd.n6655 gnd.n6654 585
R4779 gnd.n6679 gnd.n6653 585
R4780 gnd.n6680 gnd.n6652 585
R4781 gnd.n6681 gnd.n6651 585
R4782 gnd.n6648 gnd.n6647 585
R4783 gnd.n6691 gnd.n6646 585
R4784 gnd.n6692 gnd.n6645 585
R4785 gnd.n6644 gnd.n6636 585
R4786 gnd.n6699 gnd.n6635 585
R4787 gnd.n6700 gnd.n6634 585
R4788 gnd.n6628 gnd.n6627 585
R4789 gnd.n6707 gnd.n6626 585
R4790 gnd.n6708 gnd.n6625 585
R4791 gnd.n6624 gnd.n6616 585
R4792 gnd.n6715 gnd.n6615 585
R4793 gnd.n6716 gnd.n6614 585
R4794 gnd.n6608 gnd.n6607 585
R4795 gnd.n6723 gnd.n6606 585
R4796 gnd.n6724 gnd.n6605 585
R4797 gnd.n6604 gnd.n6596 585
R4798 gnd.n6732 gnd.n6731 585
R4799 gnd.n6566 gnd.n6130 482.89
R4800 gnd.n6564 gnd.n6132 482.89
R4801 gnd.n5466 gnd.n5464 482.89
R4802 gnd.n5596 gnd.n5595 482.89
R4803 gnd.n5446 gnd.t240 443.966
R4804 gnd.n6389 gnd.t257 443.966
R4805 gnd.n5438 gnd.t289 443.966
R4806 gnd.n6483 gnd.t202 443.966
R4807 gnd.n2844 gnd.n2843 374.827
R4808 gnd.n5131 gnd.t223 371.625
R4809 gnd.n122 gnd.t234 371.625
R4810 gnd.n6686 gnd.t247 371.625
R4811 gnd.n1161 gnd.t274 371.625
R4812 gnd.n554 gnd.t217 371.625
R4813 gnd.n576 gnd.t206 371.625
R4814 gnd.n201 gnd.t267 371.625
R4815 gnd.n7800 gnd.t187 371.625
R4816 gnd.n4594 gnd.t283 371.625
R4817 gnd.n4626 gnd.t260 371.625
R4818 gnd.n4449 gnd.t280 371.625
R4819 gnd.n1257 gnd.t277 371.625
R4820 gnd.n1220 gnd.t195 371.625
R4821 gnd.n6663 gnd.t191 371.625
R4822 gnd.n3463 gnd.t270 323.425
R4823 gnd.n1603 gnd.t213 323.425
R4824 gnd.n4311 gnd.n4285 289.615
R4825 gnd.n4279 gnd.n4253 289.615
R4826 gnd.n4247 gnd.n4221 289.615
R4827 gnd.n4216 gnd.n4190 289.615
R4828 gnd.n4184 gnd.n4158 289.615
R4829 gnd.n4152 gnd.n4126 289.615
R4830 gnd.n4120 gnd.n4094 289.615
R4831 gnd.n4089 gnd.n4063 289.615
R4832 gnd.n3537 gnd.t250 279.217
R4833 gnd.n1629 gnd.t227 279.217
R4834 gnd.n5408 gnd.t266 260.649
R4835 gnd.n6418 gnd.t201 260.649
R4836 gnd.n5423 gnd.n1042 256.663
R4837 gnd.n5425 gnd.n1042 256.663
R4838 gnd.n5585 gnd.n1042 256.663
R4839 gnd.n5579 gnd.n1042 256.663
R4840 gnd.n5577 gnd.n1042 256.663
R4841 gnd.n5571 gnd.n1042 256.663
R4842 gnd.n5569 gnd.n1042 256.663
R4843 gnd.n5563 gnd.n1042 256.663
R4844 gnd.n5561 gnd.n1042 256.663
R4845 gnd.n5555 gnd.n1042 256.663
R4846 gnd.n5553 gnd.n1042 256.663
R4847 gnd.n5547 gnd.n1042 256.663
R4848 gnd.n5545 gnd.n1042 256.663
R4849 gnd.n5539 gnd.n1042 256.663
R4850 gnd.n5441 gnd.n1042 256.663
R4851 gnd.n5533 gnd.n1042 256.663
R4852 gnd.n5532 gnd.n5531 256.663
R4853 gnd.n5443 gnd.n1042 256.663
R4854 gnd.n5528 gnd.n1042 256.663
R4855 gnd.n5521 gnd.n1042 256.663
R4856 gnd.n5519 gnd.n1042 256.663
R4857 gnd.n5513 gnd.n1042 256.663
R4858 gnd.n5511 gnd.n1042 256.663
R4859 gnd.n5505 gnd.n1042 256.663
R4860 gnd.n5503 gnd.n1042 256.663
R4861 gnd.n5497 gnd.n1042 256.663
R4862 gnd.n5495 gnd.n1042 256.663
R4863 gnd.n5489 gnd.n1042 256.663
R4864 gnd.n5487 gnd.n1042 256.663
R4865 gnd.n5481 gnd.n1042 256.663
R4866 gnd.n5479 gnd.n1042 256.663
R4867 gnd.n5473 gnd.n1042 256.663
R4868 gnd.n5471 gnd.n1042 256.663
R4869 gnd.n5465 gnd.n1042 256.663
R4870 gnd.n6559 gnd.n720 256.663
R4871 gnd.n6557 gnd.n720 256.663
R4872 gnd.n6551 gnd.n720 256.663
R4873 gnd.n6549 gnd.n720 256.663
R4874 gnd.n6543 gnd.n720 256.663
R4875 gnd.n6541 gnd.n720 256.663
R4876 gnd.n6535 gnd.n720 256.663
R4877 gnd.n6533 gnd.n720 256.663
R4878 gnd.n6527 gnd.n720 256.663
R4879 gnd.n6525 gnd.n720 256.663
R4880 gnd.n6519 gnd.n720 256.663
R4881 gnd.n6517 gnd.n720 256.663
R4882 gnd.n6511 gnd.n720 256.663
R4883 gnd.n6509 gnd.n720 256.663
R4884 gnd.n6502 gnd.n720 256.663
R4885 gnd.n6500 gnd.n720 256.663
R4886 gnd.n6496 gnd.n551 256.663
R4887 gnd.n6495 gnd.n720 256.663
R4888 gnd.n6392 gnd.n720 256.663
R4889 gnd.n6488 gnd.n720 256.663
R4890 gnd.n6479 gnd.n720 256.663
R4891 gnd.n6477 gnd.n720 256.663
R4892 gnd.n6471 gnd.n720 256.663
R4893 gnd.n6469 gnd.n720 256.663
R4894 gnd.n6463 gnd.n720 256.663
R4895 gnd.n6461 gnd.n720 256.663
R4896 gnd.n6455 gnd.n720 256.663
R4897 gnd.n6453 gnd.n720 256.663
R4898 gnd.n6447 gnd.n720 256.663
R4899 gnd.n6445 gnd.n720 256.663
R4900 gnd.n6439 gnd.n720 256.663
R4901 gnd.n6437 gnd.n720 256.663
R4902 gnd.n6431 gnd.n720 256.663
R4903 gnd.n6429 gnd.n720 256.663
R4904 gnd.n4469 gnd.n4444 242.672
R4905 gnd.n4471 gnd.n4444 242.672
R4906 gnd.n4479 gnd.n4444 242.672
R4907 gnd.n4481 gnd.n4444 242.672
R4908 gnd.n4489 gnd.n4444 242.672
R4909 gnd.n4491 gnd.n4444 242.672
R4910 gnd.n4499 gnd.n4444 242.672
R4911 gnd.n4501 gnd.n4444 242.672
R4912 gnd.n4509 gnd.n4444 242.672
R4913 gnd.n1196 gnd.n1172 242.672
R4914 gnd.n1196 gnd.n1195 242.672
R4915 gnd.n1196 gnd.n1194 242.672
R4916 gnd.n1196 gnd.n1192 242.672
R4917 gnd.n1196 gnd.n1190 242.672
R4918 gnd.n1196 gnd.n1189 242.672
R4919 gnd.n1196 gnd.n1187 242.672
R4920 gnd.n1196 gnd.n1185 242.672
R4921 gnd.n5353 gnd.n1196 242.672
R4922 gnd.n7253 gnd.n7252 242.672
R4923 gnd.n7252 gnd.n523 242.672
R4924 gnd.n7252 gnd.n524 242.672
R4925 gnd.n7252 gnd.n525 242.672
R4926 gnd.n7252 gnd.n526 242.672
R4927 gnd.n7252 gnd.n527 242.672
R4928 gnd.n7252 gnd.n528 242.672
R4929 gnd.n7252 gnd.n529 242.672
R4930 gnd.n7252 gnd.n530 242.672
R4931 gnd.n128 gnd.n125 242.672
R4932 gnd.n7711 gnd.n128 242.672
R4933 gnd.n7707 gnd.n128 242.672
R4934 gnd.n7704 gnd.n128 242.672
R4935 gnd.n7699 gnd.n128 242.672
R4936 gnd.n7696 gnd.n128 242.672
R4937 gnd.n7691 gnd.n128 242.672
R4938 gnd.n7688 gnd.n128 242.672
R4939 gnd.n7683 gnd.n128 242.672
R4940 gnd.n3591 gnd.n3590 242.672
R4941 gnd.n3591 gnd.n3501 242.672
R4942 gnd.n3591 gnd.n3502 242.672
R4943 gnd.n3591 gnd.n3503 242.672
R4944 gnd.n3591 gnd.n3504 242.672
R4945 gnd.n3591 gnd.n3505 242.672
R4946 gnd.n3591 gnd.n3506 242.672
R4947 gnd.n3591 gnd.n3507 242.672
R4948 gnd.n3591 gnd.n3508 242.672
R4949 gnd.n3591 gnd.n3509 242.672
R4950 gnd.n3591 gnd.n3510 242.672
R4951 gnd.n3591 gnd.n3511 242.672
R4952 gnd.n3592 gnd.n3591 242.672
R4953 gnd.n4443 gnd.n1578 242.672
R4954 gnd.n4443 gnd.n1577 242.672
R4955 gnd.n4443 gnd.n1576 242.672
R4956 gnd.n4443 gnd.n1575 242.672
R4957 gnd.n4443 gnd.n1574 242.672
R4958 gnd.n4443 gnd.n1573 242.672
R4959 gnd.n4443 gnd.n1572 242.672
R4960 gnd.n4443 gnd.n1571 242.672
R4961 gnd.n4443 gnd.n1570 242.672
R4962 gnd.n4443 gnd.n1569 242.672
R4963 gnd.n4443 gnd.n1568 242.672
R4964 gnd.n4443 gnd.n1567 242.672
R4965 gnd.n4443 gnd.n1566 242.672
R4966 gnd.n3675 gnd.n3674 242.672
R4967 gnd.n3674 gnd.n3413 242.672
R4968 gnd.n3674 gnd.n3414 242.672
R4969 gnd.n3674 gnd.n3415 242.672
R4970 gnd.n3674 gnd.n3416 242.672
R4971 gnd.n3674 gnd.n3417 242.672
R4972 gnd.n3674 gnd.n3418 242.672
R4973 gnd.n3674 gnd.n3419 242.672
R4974 gnd.n4443 gnd.n1579 242.672
R4975 gnd.n4443 gnd.n1580 242.672
R4976 gnd.n4443 gnd.n1581 242.672
R4977 gnd.n4443 gnd.n1582 242.672
R4978 gnd.n4443 gnd.n1583 242.672
R4979 gnd.n4443 gnd.n1584 242.672
R4980 gnd.n4443 gnd.n1585 242.672
R4981 gnd.n4443 gnd.n1586 242.672
R4982 gnd.n4750 gnd.n4444 242.672
R4983 gnd.n4570 gnd.n4444 242.672
R4984 gnd.n4743 gnd.n4444 242.672
R4985 gnd.n4737 gnd.n4444 242.672
R4986 gnd.n4735 gnd.n4444 242.672
R4987 gnd.n4729 gnd.n4444 242.672
R4988 gnd.n4727 gnd.n4444 242.672
R4989 gnd.n4721 gnd.n4444 242.672
R4990 gnd.n4719 gnd.n4444 242.672
R4991 gnd.n4713 gnd.n4444 242.672
R4992 gnd.n4711 gnd.n4444 242.672
R4993 gnd.n4705 gnd.n4444 242.672
R4994 gnd.n4703 gnd.n4444 242.672
R4995 gnd.n4697 gnd.n4444 242.672
R4996 gnd.n4695 gnd.n4444 242.672
R4997 gnd.n4689 gnd.n4444 242.672
R4998 gnd.n4687 gnd.n4444 242.672
R4999 gnd.n4624 gnd.n4444 242.672
R5000 gnd.n4677 gnd.n4444 242.672
R5001 gnd.n5672 gnd.n1196 242.672
R5002 gnd.n1260 gnd.n1196 242.672
R5003 gnd.n5679 gnd.n1196 242.672
R5004 gnd.n1251 gnd.n1196 242.672
R5005 gnd.n5686 gnd.n1196 242.672
R5006 gnd.n1244 gnd.n1196 242.672
R5007 gnd.n5693 gnd.n1196 242.672
R5008 gnd.n1237 gnd.n1196 242.672
R5009 gnd.n5700 gnd.n1196 242.672
R5010 gnd.n1230 gnd.n1196 242.672
R5011 gnd.n5707 gnd.n1196 242.672
R5012 gnd.n5708 gnd.n1222 242.672
R5013 gnd.n5709 gnd.n1196 242.672
R5014 gnd.n1219 gnd.n1196 242.672
R5015 gnd.n5716 gnd.n1196 242.672
R5016 gnd.n1212 gnd.n1196 242.672
R5017 gnd.n5723 gnd.n1196 242.672
R5018 gnd.n1205 gnd.n1196 242.672
R5019 gnd.n5730 gnd.n1196 242.672
R5020 gnd.n5733 gnd.n1196 242.672
R5021 gnd.n7252 gnd.n7251 242.672
R5022 gnd.n7252 gnd.n505 242.672
R5023 gnd.n7252 gnd.n506 242.672
R5024 gnd.n7252 gnd.n507 242.672
R5025 gnd.n7252 gnd.n508 242.672
R5026 gnd.n7252 gnd.n509 242.672
R5027 gnd.n7252 gnd.n510 242.672
R5028 gnd.n7252 gnd.n511 242.672
R5029 gnd.n7220 gnd.n552 242.672
R5030 gnd.n7252 gnd.n512 242.672
R5031 gnd.n7252 gnd.n513 242.672
R5032 gnd.n7252 gnd.n514 242.672
R5033 gnd.n7252 gnd.n515 242.672
R5034 gnd.n7252 gnd.n516 242.672
R5035 gnd.n7252 gnd.n517 242.672
R5036 gnd.n7252 gnd.n518 242.672
R5037 gnd.n7252 gnd.n519 242.672
R5038 gnd.n7252 gnd.n520 242.672
R5039 gnd.n7252 gnd.n521 242.672
R5040 gnd.n7252 gnd.n522 242.672
R5041 gnd.n198 gnd.n128 242.672
R5042 gnd.n7768 gnd.n128 242.672
R5043 gnd.n194 gnd.n128 242.672
R5044 gnd.n7775 gnd.n128 242.672
R5045 gnd.n187 gnd.n128 242.672
R5046 gnd.n7782 gnd.n128 242.672
R5047 gnd.n180 gnd.n128 242.672
R5048 gnd.n7789 gnd.n128 242.672
R5049 gnd.n173 gnd.n128 242.672
R5050 gnd.n7796 gnd.n128 242.672
R5051 gnd.n166 gnd.n128 242.672
R5052 gnd.n7806 gnd.n128 242.672
R5053 gnd.n159 gnd.n128 242.672
R5054 gnd.n7813 gnd.n128 242.672
R5055 gnd.n152 gnd.n128 242.672
R5056 gnd.n7820 gnd.n128 242.672
R5057 gnd.n145 gnd.n128 242.672
R5058 gnd.n7827 gnd.n128 242.672
R5059 gnd.n138 gnd.n128 242.672
R5060 gnd.n5791 gnd.n5790 242.672
R5061 gnd.n5791 gnd.n1105 242.672
R5062 gnd.n5791 gnd.n1106 242.672
R5063 gnd.n5791 gnd.n1107 242.672
R5064 gnd.n5791 gnd.n1108 242.672
R5065 gnd.n5791 gnd.n1109 242.672
R5066 gnd.n5791 gnd.n1110 242.672
R5067 gnd.n5791 gnd.n1111 242.672
R5068 gnd.n5791 gnd.n1112 242.672
R5069 gnd.n5791 gnd.n1113 242.672
R5070 gnd.n5791 gnd.n1114 242.672
R5071 gnd.n5791 gnd.n1115 242.672
R5072 gnd.n5791 gnd.n1116 242.672
R5073 gnd.n5792 gnd.n5791 242.672
R5074 gnd.n7076 gnd.n653 242.672
R5075 gnd.n7076 gnd.n652 242.672
R5076 gnd.n7076 gnd.n651 242.672
R5077 gnd.n7076 gnd.n650 242.672
R5078 gnd.n7076 gnd.n649 242.672
R5079 gnd.n7076 gnd.n648 242.672
R5080 gnd.n7076 gnd.n647 242.672
R5081 gnd.n7076 gnd.n646 242.672
R5082 gnd.n7076 gnd.n645 242.672
R5083 gnd.n7076 gnd.n644 242.672
R5084 gnd.n7076 gnd.n643 242.672
R5085 gnd.n7076 gnd.n642 242.672
R5086 gnd.n7076 gnd.n641 242.672
R5087 gnd.n7076 gnd.n640 242.672
R5088 gnd.n135 gnd.n131 240.244
R5089 gnd.n7829 gnd.n7828 240.244
R5090 gnd.n7826 gnd.n139 240.244
R5091 gnd.n7822 gnd.n7821 240.244
R5092 gnd.n7819 gnd.n146 240.244
R5093 gnd.n7815 gnd.n7814 240.244
R5094 gnd.n7812 gnd.n153 240.244
R5095 gnd.n7808 gnd.n7807 240.244
R5096 gnd.n7805 gnd.n160 240.244
R5097 gnd.n7798 gnd.n7797 240.244
R5098 gnd.n7795 gnd.n167 240.244
R5099 gnd.n7791 gnd.n7790 240.244
R5100 gnd.n7788 gnd.n174 240.244
R5101 gnd.n7784 gnd.n7783 240.244
R5102 gnd.n7781 gnd.n181 240.244
R5103 gnd.n7777 gnd.n7776 240.244
R5104 gnd.n7774 gnd.n188 240.244
R5105 gnd.n7770 gnd.n7769 240.244
R5106 gnd.n7767 gnd.n195 240.244
R5107 gnd.n7177 gnd.n496 240.244
R5108 gnd.n602 gnd.n496 240.244
R5109 gnd.n602 gnd.n487 240.244
R5110 gnd.n608 gnd.n487 240.244
R5111 gnd.n608 gnd.n478 240.244
R5112 gnd.n612 gnd.n478 240.244
R5113 gnd.n612 gnd.n469 240.244
R5114 gnd.n618 gnd.n469 240.244
R5115 gnd.n618 gnd.n461 240.244
R5116 gnd.n7129 gnd.n461 240.244
R5117 gnd.n7129 gnd.n452 240.244
R5118 gnd.n7150 gnd.n452 240.244
R5119 gnd.n7150 gnd.n441 240.244
R5120 gnd.n7146 gnd.n441 240.244
R5121 gnd.n7146 gnd.n431 240.244
R5122 gnd.n7142 gnd.n431 240.244
R5123 gnd.n7142 gnd.n423 240.244
R5124 gnd.n423 gnd.n406 240.244
R5125 gnd.n406 gnd.n395 240.244
R5126 gnd.n7402 gnd.n395 240.244
R5127 gnd.n7402 gnd.n391 240.244
R5128 gnd.n7414 gnd.n391 240.244
R5129 gnd.n7414 gnd.n374 240.244
R5130 gnd.n7410 gnd.n374 240.244
R5131 gnd.n7410 gnd.n361 240.244
R5132 gnd.n7448 gnd.n361 240.244
R5133 gnd.n7448 gnd.n357 240.244
R5134 gnd.n7538 gnd.n357 240.244
R5135 gnd.n7538 gnd.n312 240.244
R5136 gnd.n7534 gnd.n312 240.244
R5137 gnd.n7534 gnd.n349 240.244
R5138 gnd.n7530 gnd.n349 240.244
R5139 gnd.n7530 gnd.n344 240.244
R5140 gnd.n7527 gnd.n344 240.244
R5141 gnd.n7527 gnd.n334 240.244
R5142 gnd.n334 gnd.n327 240.244
R5143 gnd.n7523 gnd.n327 240.244
R5144 gnd.n7523 gnd.n299 240.244
R5145 gnd.n7520 gnd.n299 240.244
R5146 gnd.n7520 gnd.n290 240.244
R5147 gnd.n7517 gnd.n290 240.244
R5148 gnd.n7517 gnd.n282 240.244
R5149 gnd.n7514 gnd.n282 240.244
R5150 gnd.n7514 gnd.n275 240.244
R5151 gnd.n7511 gnd.n275 240.244
R5152 gnd.n7511 gnd.n269 240.244
R5153 gnd.n7508 gnd.n269 240.244
R5154 gnd.n7508 gnd.n260 240.244
R5155 gnd.n7505 gnd.n260 240.244
R5156 gnd.n7505 gnd.n252 240.244
R5157 gnd.n7502 gnd.n252 240.244
R5158 gnd.n7502 gnd.n245 240.244
R5159 gnd.n7499 gnd.n245 240.244
R5160 gnd.n7499 gnd.n239 240.244
R5161 gnd.n7496 gnd.n239 240.244
R5162 gnd.n7496 gnd.n230 240.244
R5163 gnd.n7493 gnd.n230 240.244
R5164 gnd.n7493 gnd.n223 240.244
R5165 gnd.n7489 gnd.n223 240.244
R5166 gnd.n7489 gnd.n214 240.244
R5167 gnd.n214 gnd.n205 240.244
R5168 gnd.n7758 gnd.n205 240.244
R5169 gnd.n7759 gnd.n7758 240.244
R5170 gnd.n7759 gnd.n127 240.244
R5171 gnd.n534 gnd.n533 240.244
R5172 gnd.n7245 gnd.n533 240.244
R5173 gnd.n7243 gnd.n7242 240.244
R5174 gnd.n7239 gnd.n7238 240.244
R5175 gnd.n7235 gnd.n7234 240.244
R5176 gnd.n7231 gnd.n7230 240.244
R5177 gnd.n7227 gnd.n7226 240.244
R5178 gnd.n7223 gnd.n7222 240.244
R5179 gnd.n7218 gnd.n7217 240.244
R5180 gnd.n7214 gnd.n7213 240.244
R5181 gnd.n7210 gnd.n7209 240.244
R5182 gnd.n7206 gnd.n7205 240.244
R5183 gnd.n7202 gnd.n7201 240.244
R5184 gnd.n7198 gnd.n7197 240.244
R5185 gnd.n7194 gnd.n7193 240.244
R5186 gnd.n7190 gnd.n7189 240.244
R5187 gnd.n7186 gnd.n7185 240.244
R5188 gnd.n575 gnd.n574 240.244
R5189 gnd.n7262 gnd.n494 240.244
R5190 gnd.n7262 gnd.n490 240.244
R5191 gnd.n7268 gnd.n490 240.244
R5192 gnd.n7268 gnd.n476 240.244
R5193 gnd.n7278 gnd.n476 240.244
R5194 gnd.n7278 gnd.n472 240.244
R5195 gnd.n7284 gnd.n472 240.244
R5196 gnd.n7284 gnd.n459 240.244
R5197 gnd.n7294 gnd.n459 240.244
R5198 gnd.n7294 gnd.n455 240.244
R5199 gnd.n7300 gnd.n455 240.244
R5200 gnd.n7300 gnd.n439 240.244
R5201 gnd.n7316 gnd.n439 240.244
R5202 gnd.n7316 gnd.n434 240.244
R5203 gnd.n7324 gnd.n434 240.244
R5204 gnd.n7324 gnd.n435 240.244
R5205 gnd.n435 gnd.n404 240.244
R5206 gnd.n7392 gnd.n404 240.244
R5207 gnd.n7392 gnd.n399 240.244
R5208 gnd.n7400 gnd.n399 240.244
R5209 gnd.n7400 gnd.n400 240.244
R5210 gnd.n400 gnd.n371 240.244
R5211 gnd.n7439 gnd.n371 240.244
R5212 gnd.n7439 gnd.n372 240.244
R5213 gnd.n372 gnd.n366 240.244
R5214 gnd.n7446 gnd.n366 240.244
R5215 gnd.n7446 gnd.n367 240.244
R5216 gnd.n367 gnd.n309 240.244
R5217 gnd.n7585 gnd.n309 240.244
R5218 gnd.n7585 gnd.n310 240.244
R5219 gnd.n7550 gnd.n310 240.244
R5220 gnd.n7551 gnd.n7550 240.244
R5221 gnd.n7554 gnd.n7551 240.244
R5222 gnd.n7554 gnd.n329 240.244
R5223 gnd.n7566 gnd.n329 240.244
R5224 gnd.n7568 gnd.n7566 240.244
R5225 gnd.n7568 gnd.n300 240.244
R5226 gnd.n7592 gnd.n300 240.244
R5227 gnd.n7592 gnd.n288 240.244
R5228 gnd.n7602 gnd.n288 240.244
R5229 gnd.n7602 gnd.n284 240.244
R5230 gnd.n7608 gnd.n284 240.244
R5231 gnd.n7608 gnd.n274 240.244
R5232 gnd.n7618 gnd.n274 240.244
R5233 gnd.n7618 gnd.n270 240.244
R5234 gnd.n7624 gnd.n270 240.244
R5235 gnd.n7624 gnd.n258 240.244
R5236 gnd.n7634 gnd.n258 240.244
R5237 gnd.n7634 gnd.n254 240.244
R5238 gnd.n7640 gnd.n254 240.244
R5239 gnd.n7640 gnd.n244 240.244
R5240 gnd.n7650 gnd.n244 240.244
R5241 gnd.n7650 gnd.n240 240.244
R5242 gnd.n7656 gnd.n240 240.244
R5243 gnd.n7656 gnd.n228 240.244
R5244 gnd.n7666 gnd.n228 240.244
R5245 gnd.n7666 gnd.n224 240.244
R5246 gnd.n7672 gnd.n224 240.244
R5247 gnd.n7672 gnd.n212 240.244
R5248 gnd.n7750 gnd.n212 240.244
R5249 gnd.n7750 gnd.n208 240.244
R5250 gnd.n7756 gnd.n208 240.244
R5251 gnd.n7756 gnd.n130 240.244
R5252 gnd.n7836 gnd.n130 240.244
R5253 gnd.n5734 gnd.n1180 240.244
R5254 gnd.n5732 gnd.n5731 240.244
R5255 gnd.n5729 gnd.n1198 240.244
R5256 gnd.n5725 gnd.n5724 240.244
R5257 gnd.n5722 gnd.n1206 240.244
R5258 gnd.n5718 gnd.n5717 240.244
R5259 gnd.n5715 gnd.n1213 240.244
R5260 gnd.n5711 gnd.n5710 240.244
R5261 gnd.n5706 gnd.n1223 240.244
R5262 gnd.n5702 gnd.n5701 240.244
R5263 gnd.n5699 gnd.n1231 240.244
R5264 gnd.n5695 gnd.n5694 240.244
R5265 gnd.n5692 gnd.n1238 240.244
R5266 gnd.n5688 gnd.n5687 240.244
R5267 gnd.n5685 gnd.n1245 240.244
R5268 gnd.n5681 gnd.n5680 240.244
R5269 gnd.n5678 gnd.n1252 240.244
R5270 gnd.n5674 gnd.n5673 240.244
R5271 gnd.n4630 gnd.n4445 240.244
R5272 gnd.n4630 gnd.n1558 240.244
R5273 gnd.n4670 gnd.n1558 240.244
R5274 gnd.n4670 gnd.n1551 240.244
R5275 gnd.n4667 gnd.n1551 240.244
R5276 gnd.n4667 gnd.n1543 240.244
R5277 gnd.n4664 gnd.n1543 240.244
R5278 gnd.n4664 gnd.n1534 240.244
R5279 gnd.n4661 gnd.n1534 240.244
R5280 gnd.n4661 gnd.n1526 240.244
R5281 gnd.n4658 gnd.n1526 240.244
R5282 gnd.n4658 gnd.n1519 240.244
R5283 gnd.n4655 gnd.n1519 240.244
R5284 gnd.n4655 gnd.n1511 240.244
R5285 gnd.n4652 gnd.n1511 240.244
R5286 gnd.n4652 gnd.n1502 240.244
R5287 gnd.n4649 gnd.n1502 240.244
R5288 gnd.n4649 gnd.n1493 240.244
R5289 gnd.n1493 gnd.n1483 240.244
R5290 gnd.n4849 gnd.n1483 240.244
R5291 gnd.n4849 gnd.n1479 240.244
R5292 gnd.n4860 gnd.n1479 240.244
R5293 gnd.n4860 gnd.n1458 240.244
R5294 gnd.n4856 gnd.n1458 240.244
R5295 gnd.n4856 gnd.n1448 240.244
R5296 gnd.n4889 gnd.n1448 240.244
R5297 gnd.n4889 gnd.n1444 240.244
R5298 gnd.n4900 gnd.n1444 240.244
R5299 gnd.n4900 gnd.n1393 240.244
R5300 gnd.n4896 gnd.n1393 240.244
R5301 gnd.n4896 gnd.n1404 240.244
R5302 gnd.n1410 gnd.n1404 240.244
R5303 gnd.n5203 gnd.n1410 240.244
R5304 gnd.n5203 gnd.n5202 240.244
R5305 gnd.n5202 gnd.n1423 240.244
R5306 gnd.n5198 gnd.n1423 240.244
R5307 gnd.n5198 gnd.n1378 240.244
R5308 gnd.n4994 gnd.n1378 240.244
R5309 gnd.n4994 gnd.n1369 240.244
R5310 gnd.n4998 gnd.n1369 240.244
R5311 gnd.n4998 gnd.n1361 240.244
R5312 gnd.n5004 gnd.n1361 240.244
R5313 gnd.n5004 gnd.n1352 240.244
R5314 gnd.n5008 gnd.n1352 240.244
R5315 gnd.n5008 gnd.n1343 240.244
R5316 gnd.n5032 gnd.n1343 240.244
R5317 gnd.n5032 gnd.n1334 240.244
R5318 gnd.n5028 gnd.n1334 240.244
R5319 gnd.n5028 gnd.n1326 240.244
R5320 gnd.n5024 gnd.n1326 240.244
R5321 gnd.n5024 gnd.n1317 240.244
R5322 gnd.n5020 gnd.n1317 240.244
R5323 gnd.n5020 gnd.n1308 240.244
R5324 gnd.n5098 gnd.n1308 240.244
R5325 gnd.n5098 gnd.n1299 240.244
R5326 gnd.n5104 gnd.n1299 240.244
R5327 gnd.n5104 gnd.n1291 240.244
R5328 gnd.n5108 gnd.n1291 240.244
R5329 gnd.n5108 gnd.n1282 240.244
R5330 gnd.n5117 gnd.n1282 240.244
R5331 gnd.n5117 gnd.n1272 240.244
R5332 gnd.n1272 gnd.n1264 240.244
R5333 gnd.n5665 gnd.n1264 240.244
R5334 gnd.n5665 gnd.n1176 240.244
R5335 gnd.n4751 gnd.n4749 240.244
R5336 gnd.n4749 gnd.n4748 240.244
R5337 gnd.n4745 gnd.n4744 240.244
R5338 gnd.n4742 gnd.n4575 240.244
R5339 gnd.n4738 gnd.n4736 240.244
R5340 gnd.n4734 gnd.n4581 240.244
R5341 gnd.n4730 gnd.n4728 240.244
R5342 gnd.n4726 gnd.n4587 240.244
R5343 gnd.n4722 gnd.n4720 240.244
R5344 gnd.n4718 gnd.n4593 240.244
R5345 gnd.n4714 gnd.n4712 240.244
R5346 gnd.n4710 gnd.n4602 240.244
R5347 gnd.n4706 gnd.n4704 240.244
R5348 gnd.n4702 gnd.n4608 240.244
R5349 gnd.n4698 gnd.n4696 240.244
R5350 gnd.n4694 gnd.n4614 240.244
R5351 gnd.n4690 gnd.n4688 240.244
R5352 gnd.n4686 gnd.n4620 240.244
R5353 gnd.n4676 gnd.n4625 240.244
R5354 gnd.n4757 gnd.n1557 240.244
R5355 gnd.n4767 gnd.n1557 240.244
R5356 gnd.n4767 gnd.n1553 240.244
R5357 gnd.n4773 gnd.n1553 240.244
R5358 gnd.n4773 gnd.n1541 240.244
R5359 gnd.n4783 gnd.n1541 240.244
R5360 gnd.n4783 gnd.n1537 240.244
R5361 gnd.n4789 gnd.n1537 240.244
R5362 gnd.n4789 gnd.n1525 240.244
R5363 gnd.n4799 gnd.n1525 240.244
R5364 gnd.n4799 gnd.n1521 240.244
R5365 gnd.n4805 gnd.n1521 240.244
R5366 gnd.n4805 gnd.n1509 240.244
R5367 gnd.n4815 gnd.n1509 240.244
R5368 gnd.n4815 gnd.n1505 240.244
R5369 gnd.n4821 gnd.n1505 240.244
R5370 gnd.n4821 gnd.n1492 240.244
R5371 gnd.n4839 gnd.n1492 240.244
R5372 gnd.n4839 gnd.n1487 240.244
R5373 gnd.n4847 gnd.n1487 240.244
R5374 gnd.n4847 gnd.n1488 240.244
R5375 gnd.n1488 gnd.n1456 240.244
R5376 gnd.n4880 gnd.n1456 240.244
R5377 gnd.n4880 gnd.n1457 240.244
R5378 gnd.n1457 gnd.n1451 240.244
R5379 gnd.n4887 gnd.n1451 240.244
R5380 gnd.n4887 gnd.n1452 240.244
R5381 gnd.n1452 gnd.n1390 240.244
R5382 gnd.n5239 gnd.n1390 240.244
R5383 gnd.n5239 gnd.n1391 240.244
R5384 gnd.n5231 gnd.n1391 240.244
R5385 gnd.n5231 gnd.n5228 240.244
R5386 gnd.n5228 gnd.n1407 240.244
R5387 gnd.n5215 gnd.n1407 240.244
R5388 gnd.n5218 gnd.n5215 240.244
R5389 gnd.n5218 gnd.n1381 240.244
R5390 gnd.n5245 gnd.n1381 240.244
R5391 gnd.n5245 gnd.n1368 240.244
R5392 gnd.n5255 gnd.n1368 240.244
R5393 gnd.n5255 gnd.n1364 240.244
R5394 gnd.n5261 gnd.n1364 240.244
R5395 gnd.n5261 gnd.n1350 240.244
R5396 gnd.n5271 gnd.n1350 240.244
R5397 gnd.n5271 gnd.n1346 240.244
R5398 gnd.n5277 gnd.n1346 240.244
R5399 gnd.n5277 gnd.n1333 240.244
R5400 gnd.n5287 gnd.n1333 240.244
R5401 gnd.n5287 gnd.n1329 240.244
R5402 gnd.n5293 gnd.n1329 240.244
R5403 gnd.n5293 gnd.n1315 240.244
R5404 gnd.n5303 gnd.n1315 240.244
R5405 gnd.n5303 gnd.n1311 240.244
R5406 gnd.n5309 gnd.n1311 240.244
R5407 gnd.n5309 gnd.n1298 240.244
R5408 gnd.n5319 gnd.n1298 240.244
R5409 gnd.n5319 gnd.n1294 240.244
R5410 gnd.n5325 gnd.n1294 240.244
R5411 gnd.n5325 gnd.n1280 240.244
R5412 gnd.n5335 gnd.n1280 240.244
R5413 gnd.n5335 gnd.n1275 240.244
R5414 gnd.n5343 gnd.n1275 240.244
R5415 gnd.n5343 gnd.n1276 240.244
R5416 gnd.n1276 gnd.n1179 240.244
R5417 gnd.n5740 gnd.n1179 240.244
R5418 gnd.n4442 gnd.n1588 240.244
R5419 gnd.n4435 gnd.n4434 240.244
R5420 gnd.n4432 gnd.n4431 240.244
R5421 gnd.n4428 gnd.n4427 240.244
R5422 gnd.n4424 gnd.n4423 240.244
R5423 gnd.n4420 gnd.n4419 240.244
R5424 gnd.n4416 gnd.n4415 240.244
R5425 gnd.n4412 gnd.n4411 240.244
R5426 gnd.n3686 gnd.n3398 240.244
R5427 gnd.n3696 gnd.n3398 240.244
R5428 gnd.n3696 gnd.n3389 240.244
R5429 gnd.n3389 gnd.n3378 240.244
R5430 gnd.n3717 gnd.n3378 240.244
R5431 gnd.n3717 gnd.n3372 240.244
R5432 gnd.n3727 gnd.n3372 240.244
R5433 gnd.n3727 gnd.n3361 240.244
R5434 gnd.n3361 gnd.n3353 240.244
R5435 gnd.n3745 gnd.n3353 240.244
R5436 gnd.n3746 gnd.n3745 240.244
R5437 gnd.n3746 gnd.n3338 240.244
R5438 gnd.n3748 gnd.n3338 240.244
R5439 gnd.n3748 gnd.n3324 240.244
R5440 gnd.n3790 gnd.n3324 240.244
R5441 gnd.n3791 gnd.n3790 240.244
R5442 gnd.n3794 gnd.n3791 240.244
R5443 gnd.n3794 gnd.n3279 240.244
R5444 gnd.n3319 gnd.n3279 240.244
R5445 gnd.n3319 gnd.n3289 240.244
R5446 gnd.n3804 gnd.n3289 240.244
R5447 gnd.n3804 gnd.n3310 240.244
R5448 gnd.n3814 gnd.n3310 240.244
R5449 gnd.n3814 gnd.n3196 240.244
R5450 gnd.n3859 gnd.n3196 240.244
R5451 gnd.n3859 gnd.n3182 240.244
R5452 gnd.n3881 gnd.n3182 240.244
R5453 gnd.n3882 gnd.n3881 240.244
R5454 gnd.n3882 gnd.n3169 240.244
R5455 gnd.n3169 gnd.n3158 240.244
R5456 gnd.n3913 gnd.n3158 240.244
R5457 gnd.n3914 gnd.n3913 240.244
R5458 gnd.n3915 gnd.n3914 240.244
R5459 gnd.n3915 gnd.n3143 240.244
R5460 gnd.n3143 gnd.n3142 240.244
R5461 gnd.n3142 gnd.n3127 240.244
R5462 gnd.n3966 gnd.n3127 240.244
R5463 gnd.n3967 gnd.n3966 240.244
R5464 gnd.n3967 gnd.n3114 240.244
R5465 gnd.n3114 gnd.n3103 240.244
R5466 gnd.n3998 gnd.n3103 240.244
R5467 gnd.n3999 gnd.n3998 240.244
R5468 gnd.n4000 gnd.n3999 240.244
R5469 gnd.n4000 gnd.n3087 240.244
R5470 gnd.n3087 gnd.n3086 240.244
R5471 gnd.n3086 gnd.n3073 240.244
R5472 gnd.n4055 gnd.n3073 240.244
R5473 gnd.n4056 gnd.n4055 240.244
R5474 gnd.n4056 gnd.n1654 240.244
R5475 gnd.n1654 gnd.n1644 240.244
R5476 gnd.n4343 gnd.n1644 240.244
R5477 gnd.n4346 gnd.n4343 240.244
R5478 gnd.n4346 gnd.n4345 240.244
R5479 gnd.n3676 gnd.n3411 240.244
R5480 gnd.n3432 gnd.n3411 240.244
R5481 gnd.n3435 gnd.n3434 240.244
R5482 gnd.n3442 gnd.n3441 240.244
R5483 gnd.n3445 gnd.n3444 240.244
R5484 gnd.n3452 gnd.n3451 240.244
R5485 gnd.n3455 gnd.n3454 240.244
R5486 gnd.n3462 gnd.n3461 240.244
R5487 gnd.n3684 gnd.n3408 240.244
R5488 gnd.n3408 gnd.n3387 240.244
R5489 gnd.n3707 gnd.n3387 240.244
R5490 gnd.n3707 gnd.n3381 240.244
R5491 gnd.n3715 gnd.n3381 240.244
R5492 gnd.n3715 gnd.n3383 240.244
R5493 gnd.n3383 gnd.n3359 240.244
R5494 gnd.n3737 gnd.n3359 240.244
R5495 gnd.n3737 gnd.n3355 240.244
R5496 gnd.n3743 gnd.n3355 240.244
R5497 gnd.n3743 gnd.n3337 240.244
R5498 gnd.n3768 gnd.n3337 240.244
R5499 gnd.n3768 gnd.n3332 240.244
R5500 gnd.n3780 gnd.n3332 240.244
R5501 gnd.n3780 gnd.n3333 240.244
R5502 gnd.n3776 gnd.n3333 240.244
R5503 gnd.n3776 gnd.n3281 240.244
R5504 gnd.n3828 gnd.n3281 240.244
R5505 gnd.n3828 gnd.n3282 240.244
R5506 gnd.n3824 gnd.n3282 240.244
R5507 gnd.n3824 gnd.n3288 240.244
R5508 gnd.n3308 gnd.n3288 240.244
R5509 gnd.n3308 gnd.n3194 240.244
R5510 gnd.n3863 gnd.n3194 240.244
R5511 gnd.n3863 gnd.n3189 240.244
R5512 gnd.n3871 gnd.n3189 240.244
R5513 gnd.n3871 gnd.n3190 240.244
R5514 gnd.n3190 gnd.n3167 240.244
R5515 gnd.n3903 gnd.n3167 240.244
R5516 gnd.n3903 gnd.n3162 240.244
R5517 gnd.n3911 gnd.n3162 240.244
R5518 gnd.n3911 gnd.n3163 240.244
R5519 gnd.n3163 gnd.n3140 240.244
R5520 gnd.n3948 gnd.n3140 240.244
R5521 gnd.n3948 gnd.n3135 240.244
R5522 gnd.n3956 gnd.n3135 240.244
R5523 gnd.n3956 gnd.n3136 240.244
R5524 gnd.n3136 gnd.n3112 240.244
R5525 gnd.n3988 gnd.n3112 240.244
R5526 gnd.n3988 gnd.n3107 240.244
R5527 gnd.n3996 gnd.n3107 240.244
R5528 gnd.n3996 gnd.n3108 240.244
R5529 gnd.n3108 gnd.n3085 240.244
R5530 gnd.n4037 gnd.n3085 240.244
R5531 gnd.n4037 gnd.n3080 240.244
R5532 gnd.n4045 gnd.n3080 240.244
R5533 gnd.n4045 gnd.n3081 240.244
R5534 gnd.n3081 gnd.n1652 240.244
R5535 gnd.n4331 gnd.n1652 240.244
R5536 gnd.n4331 gnd.n1647 240.244
R5537 gnd.n4341 gnd.n1647 240.244
R5538 gnd.n4341 gnd.n1648 240.244
R5539 gnd.n1648 gnd.n1587 240.244
R5540 gnd.n1607 gnd.n1565 240.244
R5541 gnd.n4402 gnd.n4401 240.244
R5542 gnd.n4398 gnd.n4397 240.244
R5543 gnd.n4394 gnd.n4393 240.244
R5544 gnd.n4390 gnd.n4389 240.244
R5545 gnd.n4386 gnd.n4385 240.244
R5546 gnd.n4382 gnd.n4381 240.244
R5547 gnd.n4378 gnd.n4377 240.244
R5548 gnd.n4374 gnd.n4373 240.244
R5549 gnd.n4370 gnd.n4369 240.244
R5550 gnd.n4366 gnd.n4365 240.244
R5551 gnd.n4362 gnd.n4361 240.244
R5552 gnd.n4358 gnd.n4357 240.244
R5553 gnd.n3599 gnd.n3496 240.244
R5554 gnd.n3599 gnd.n3489 240.244
R5555 gnd.n3610 gnd.n3489 240.244
R5556 gnd.n3610 gnd.n3485 240.244
R5557 gnd.n3616 gnd.n3485 240.244
R5558 gnd.n3616 gnd.n3477 240.244
R5559 gnd.n3626 gnd.n3477 240.244
R5560 gnd.n3626 gnd.n3472 240.244
R5561 gnd.n3662 gnd.n3472 240.244
R5562 gnd.n3662 gnd.n3473 240.244
R5563 gnd.n3473 gnd.n3420 240.244
R5564 gnd.n3657 gnd.n3420 240.244
R5565 gnd.n3657 gnd.n3656 240.244
R5566 gnd.n3656 gnd.n3399 240.244
R5567 gnd.n3652 gnd.n3399 240.244
R5568 gnd.n3652 gnd.n3390 240.244
R5569 gnd.n3649 gnd.n3390 240.244
R5570 gnd.n3649 gnd.n3648 240.244
R5571 gnd.n3648 gnd.n3373 240.244
R5572 gnd.n3644 gnd.n3373 240.244
R5573 gnd.n3644 gnd.n3362 240.244
R5574 gnd.n3362 gnd.n3343 240.244
R5575 gnd.n3757 gnd.n3343 240.244
R5576 gnd.n3757 gnd.n3339 240.244
R5577 gnd.n3765 gnd.n3339 240.244
R5578 gnd.n3765 gnd.n3330 240.244
R5579 gnd.n3330 gnd.n3266 240.244
R5580 gnd.n3837 gnd.n3266 240.244
R5581 gnd.n3837 gnd.n3267 240.244
R5582 gnd.n3278 gnd.n3267 240.244
R5583 gnd.n3313 gnd.n3278 240.244
R5584 gnd.n3316 gnd.n3313 240.244
R5585 gnd.n3316 gnd.n3290 240.244
R5586 gnd.n3303 gnd.n3290 240.244
R5587 gnd.n3303 gnd.n3300 240.244
R5588 gnd.n3300 gnd.n3197 240.244
R5589 gnd.n3858 gnd.n3197 240.244
R5590 gnd.n3858 gnd.n3187 240.244
R5591 gnd.n3854 gnd.n3187 240.244
R5592 gnd.n3854 gnd.n3181 240.244
R5593 gnd.n3851 gnd.n3181 240.244
R5594 gnd.n3851 gnd.n3170 240.244
R5595 gnd.n3848 gnd.n3170 240.244
R5596 gnd.n3848 gnd.n3148 240.244
R5597 gnd.n3924 gnd.n3148 240.244
R5598 gnd.n3924 gnd.n3144 240.244
R5599 gnd.n3945 gnd.n3144 240.244
R5600 gnd.n3945 gnd.n3133 240.244
R5601 gnd.n3941 gnd.n3133 240.244
R5602 gnd.n3941 gnd.n3126 240.244
R5603 gnd.n3938 gnd.n3126 240.244
R5604 gnd.n3938 gnd.n3115 240.244
R5605 gnd.n3935 gnd.n3115 240.244
R5606 gnd.n3935 gnd.n3092 240.244
R5607 gnd.n4009 gnd.n3092 240.244
R5608 gnd.n4009 gnd.n3088 240.244
R5609 gnd.n4034 gnd.n3088 240.244
R5610 gnd.n4034 gnd.n3079 240.244
R5611 gnd.n4030 gnd.n3079 240.244
R5612 gnd.n4030 gnd.n3072 240.244
R5613 gnd.n4026 gnd.n3072 240.244
R5614 gnd.n4026 gnd.n1655 240.244
R5615 gnd.n4023 gnd.n1655 240.244
R5616 gnd.n4023 gnd.n1636 240.244
R5617 gnd.n4353 gnd.n1636 240.244
R5618 gnd.n3513 gnd.n3512 240.244
R5619 gnd.n3584 gnd.n3512 240.244
R5620 gnd.n3582 gnd.n3581 240.244
R5621 gnd.n3578 gnd.n3577 240.244
R5622 gnd.n3574 gnd.n3573 240.244
R5623 gnd.n3570 gnd.n3569 240.244
R5624 gnd.n3566 gnd.n3565 240.244
R5625 gnd.n3562 gnd.n3561 240.244
R5626 gnd.n3558 gnd.n3557 240.244
R5627 gnd.n3554 gnd.n3553 240.244
R5628 gnd.n3550 gnd.n3549 240.244
R5629 gnd.n3546 gnd.n3545 240.244
R5630 gnd.n3542 gnd.n3500 240.244
R5631 gnd.n3602 gnd.n3494 240.244
R5632 gnd.n3602 gnd.n3490 240.244
R5633 gnd.n3608 gnd.n3490 240.244
R5634 gnd.n3608 gnd.n3483 240.244
R5635 gnd.n3618 gnd.n3483 240.244
R5636 gnd.n3618 gnd.n3479 240.244
R5637 gnd.n3624 gnd.n3479 240.244
R5638 gnd.n3624 gnd.n3470 240.244
R5639 gnd.n3664 gnd.n3470 240.244
R5640 gnd.n3664 gnd.n3421 240.244
R5641 gnd.n3672 gnd.n3421 240.244
R5642 gnd.n3672 gnd.n3422 240.244
R5643 gnd.n3422 gnd.n3400 240.244
R5644 gnd.n3693 gnd.n3400 240.244
R5645 gnd.n3693 gnd.n3392 240.244
R5646 gnd.n3704 gnd.n3392 240.244
R5647 gnd.n3704 gnd.n3393 240.244
R5648 gnd.n3393 gnd.n3374 240.244
R5649 gnd.n3724 gnd.n3374 240.244
R5650 gnd.n3724 gnd.n3364 240.244
R5651 gnd.n3734 gnd.n3364 240.244
R5652 gnd.n3734 gnd.n3345 240.244
R5653 gnd.n3755 gnd.n3345 240.244
R5654 gnd.n3755 gnd.n3347 240.244
R5655 gnd.n3347 gnd.n3328 240.244
R5656 gnd.n3783 gnd.n3328 240.244
R5657 gnd.n3783 gnd.n3270 240.244
R5658 gnd.n3835 gnd.n3270 240.244
R5659 gnd.n3835 gnd.n3271 240.244
R5660 gnd.n3831 gnd.n3271 240.244
R5661 gnd.n3831 gnd.n3277 240.244
R5662 gnd.n3292 gnd.n3277 240.244
R5663 gnd.n3821 gnd.n3292 240.244
R5664 gnd.n3821 gnd.n3293 240.244
R5665 gnd.n3817 gnd.n3293 240.244
R5666 gnd.n3817 gnd.n3299 240.244
R5667 gnd.n3299 gnd.n3186 240.244
R5668 gnd.n3874 gnd.n3186 240.244
R5669 gnd.n3874 gnd.n3179 240.244
R5670 gnd.n3885 gnd.n3179 240.244
R5671 gnd.n3885 gnd.n3172 240.244
R5672 gnd.n3900 gnd.n3172 240.244
R5673 gnd.n3900 gnd.n3173 240.244
R5674 gnd.n3173 gnd.n3151 240.244
R5675 gnd.n3922 gnd.n3151 240.244
R5676 gnd.n3922 gnd.n3152 240.244
R5677 gnd.n3152 gnd.n3131 240.244
R5678 gnd.n3959 gnd.n3131 240.244
R5679 gnd.n3959 gnd.n3124 240.244
R5680 gnd.n3970 gnd.n3124 240.244
R5681 gnd.n3970 gnd.n3117 240.244
R5682 gnd.n3985 gnd.n3117 240.244
R5683 gnd.n3985 gnd.n3118 240.244
R5684 gnd.n3118 gnd.n3095 240.244
R5685 gnd.n4007 gnd.n3095 240.244
R5686 gnd.n4007 gnd.n3097 240.244
R5687 gnd.n3097 gnd.n3077 240.244
R5688 gnd.n4048 gnd.n3077 240.244
R5689 gnd.n4048 gnd.n3070 240.244
R5690 gnd.n4059 gnd.n3070 240.244
R5691 gnd.n4059 gnd.n3063 240.244
R5692 gnd.n4328 gnd.n3063 240.244
R5693 gnd.n4328 gnd.n3064 240.244
R5694 gnd.n3064 gnd.n1639 240.244
R5695 gnd.n4351 gnd.n1639 240.244
R5696 gnd.n7682 gnd.n7681 240.244
R5697 gnd.n7687 gnd.n7684 240.244
R5698 gnd.n7690 gnd.n7689 240.244
R5699 gnd.n7695 gnd.n7692 240.244
R5700 gnd.n7698 gnd.n7697 240.244
R5701 gnd.n7703 gnd.n7700 240.244
R5702 gnd.n7706 gnd.n7705 240.244
R5703 gnd.n7710 gnd.n7708 240.244
R5704 gnd.n7713 gnd.n7712 240.244
R5705 gnd.n7175 gnd.n497 240.244
R5706 gnd.n585 gnd.n497 240.244
R5707 gnd.n585 gnd.n488 240.244
R5708 gnd.n586 gnd.n488 240.244
R5709 gnd.n586 gnd.n479 240.244
R5710 gnd.n589 gnd.n479 240.244
R5711 gnd.n589 gnd.n470 240.244
R5712 gnd.n590 gnd.n470 240.244
R5713 gnd.n590 gnd.n462 240.244
R5714 gnd.n593 gnd.n462 240.244
R5715 gnd.n593 gnd.n453 240.244
R5716 gnd.n7152 gnd.n453 240.244
R5717 gnd.n7152 gnd.n442 240.244
R5718 gnd.n442 gnd.n429 240.244
R5719 gnd.n7326 gnd.n429 240.244
R5720 gnd.n7326 gnd.n424 240.244
R5721 gnd.n7340 gnd.n424 240.244
R5722 gnd.n7340 gnd.n407 240.244
R5723 gnd.n7333 gnd.n407 240.244
R5724 gnd.n7333 gnd.n397 240.244
R5725 gnd.n397 gnd.n389 240.244
R5726 gnd.n7416 gnd.n389 240.244
R5727 gnd.n7416 gnd.n375 240.244
R5728 gnd.n384 gnd.n375 240.244
R5729 gnd.n7424 gnd.n384 240.244
R5730 gnd.n7424 gnd.n363 240.244
R5731 gnd.n363 gnd.n355 240.244
R5732 gnd.n7540 gnd.n355 240.244
R5733 gnd.n7540 gnd.n313 240.244
R5734 gnd.n350 gnd.n313 240.244
R5735 gnd.n7547 gnd.n350 240.244
R5736 gnd.n7547 gnd.n351 240.244
R5737 gnd.n351 gnd.n82 240.244
R5738 gnd.n83 gnd.n82 240.244
R5739 gnd.n84 gnd.n83 240.244
R5740 gnd.n328 gnd.n84 240.244
R5741 gnd.n328 gnd.n87 240.244
R5742 gnd.n88 gnd.n87 240.244
R5743 gnd.n89 gnd.n88 240.244
R5744 gnd.n291 gnd.n89 240.244
R5745 gnd.n291 gnd.n92 240.244
R5746 gnd.n93 gnd.n92 240.244
R5747 gnd.n94 gnd.n93 240.244
R5748 gnd.n276 gnd.n94 240.244
R5749 gnd.n276 gnd.n97 240.244
R5750 gnd.n98 gnd.n97 240.244
R5751 gnd.n99 gnd.n98 240.244
R5752 gnd.n261 gnd.n99 240.244
R5753 gnd.n261 gnd.n102 240.244
R5754 gnd.n103 gnd.n102 240.244
R5755 gnd.n104 gnd.n103 240.244
R5756 gnd.n246 gnd.n104 240.244
R5757 gnd.n246 gnd.n107 240.244
R5758 gnd.n108 gnd.n107 240.244
R5759 gnd.n109 gnd.n108 240.244
R5760 gnd.n231 gnd.n109 240.244
R5761 gnd.n231 gnd.n112 240.244
R5762 gnd.n113 gnd.n112 240.244
R5763 gnd.n114 gnd.n113 240.244
R5764 gnd.n215 gnd.n114 240.244
R5765 gnd.n215 gnd.n117 240.244
R5766 gnd.n118 gnd.n117 240.244
R5767 gnd.n119 gnd.n118 240.244
R5768 gnd.n7838 gnd.n119 240.244
R5769 gnd.n6599 gnd.n503 240.244
R5770 gnd.n6601 gnd.n6600 240.244
R5771 gnd.n6611 gnd.n6610 240.244
R5772 gnd.n6619 gnd.n6618 240.244
R5773 gnd.n6621 gnd.n6620 240.244
R5774 gnd.n6631 gnd.n6630 240.244
R5775 gnd.n6639 gnd.n6638 240.244
R5776 gnd.n6641 gnd.n6640 240.244
R5777 gnd.n6685 gnd.n531 240.244
R5778 gnd.n7260 gnd.n499 240.244
R5779 gnd.n7260 gnd.n485 240.244
R5780 gnd.n7270 gnd.n485 240.244
R5781 gnd.n7270 gnd.n481 240.244
R5782 gnd.n7276 gnd.n481 240.244
R5783 gnd.n7276 gnd.n467 240.244
R5784 gnd.n7286 gnd.n467 240.244
R5785 gnd.n7286 gnd.n463 240.244
R5786 gnd.n7292 gnd.n463 240.244
R5787 gnd.n7292 gnd.n450 240.244
R5788 gnd.n7302 gnd.n450 240.244
R5789 gnd.n7302 gnd.n444 240.244
R5790 gnd.n7314 gnd.n444 240.244
R5791 gnd.n7314 gnd.n445 240.244
R5792 gnd.n445 gnd.n433 240.244
R5793 gnd.n7307 gnd.n433 240.244
R5794 gnd.n7307 gnd.n409 240.244
R5795 gnd.n7390 gnd.n409 240.244
R5796 gnd.n7390 gnd.n410 240.244
R5797 gnd.n410 gnd.n398 240.244
R5798 gnd.n7383 gnd.n398 240.244
R5799 gnd.n7383 gnd.n377 240.244
R5800 gnd.n7437 gnd.n377 240.244
R5801 gnd.n7437 gnd.n378 240.244
R5802 gnd.n7426 gnd.n378 240.244
R5803 gnd.n7426 gnd.n365 240.244
R5804 gnd.n7428 gnd.n365 240.244
R5805 gnd.n7428 gnd.n315 240.244
R5806 gnd.n7583 gnd.n315 240.244
R5807 gnd.n7583 gnd.n316 240.244
R5808 gnd.n321 gnd.n316 240.244
R5809 gnd.n322 gnd.n321 240.244
R5810 gnd.n323 gnd.n322 240.244
R5811 gnd.n332 gnd.n323 240.244
R5812 gnd.n332 gnd.n326 240.244
R5813 gnd.n7570 gnd.n326 240.244
R5814 gnd.n7570 gnd.n297 240.244
R5815 gnd.n7594 gnd.n297 240.244
R5816 gnd.n7594 gnd.n293 240.244
R5817 gnd.n7600 gnd.n293 240.244
R5818 gnd.n7600 gnd.n281 240.244
R5819 gnd.n7610 gnd.n281 240.244
R5820 gnd.n7610 gnd.n277 240.244
R5821 gnd.n7616 gnd.n277 240.244
R5822 gnd.n7616 gnd.n267 240.244
R5823 gnd.n7626 gnd.n267 240.244
R5824 gnd.n7626 gnd.n263 240.244
R5825 gnd.n7632 gnd.n263 240.244
R5826 gnd.n7632 gnd.n251 240.244
R5827 gnd.n7642 gnd.n251 240.244
R5828 gnd.n7642 gnd.n247 240.244
R5829 gnd.n7648 gnd.n247 240.244
R5830 gnd.n7648 gnd.n237 240.244
R5831 gnd.n7658 gnd.n237 240.244
R5832 gnd.n7658 gnd.n233 240.244
R5833 gnd.n7664 gnd.n233 240.244
R5834 gnd.n7664 gnd.n222 240.244
R5835 gnd.n7674 gnd.n222 240.244
R5836 gnd.n7674 gnd.n216 240.244
R5837 gnd.n7748 gnd.n216 240.244
R5838 gnd.n7748 gnd.n217 240.244
R5839 gnd.n217 gnd.n207 240.244
R5840 gnd.n7679 gnd.n207 240.244
R5841 gnd.n7679 gnd.n129 240.244
R5842 gnd.n5354 gnd.n5351 240.244
R5843 gnd.n5352 gnd.n1124 240.244
R5844 gnd.n1186 gnd.n1125 240.244
R5845 gnd.n1134 gnd.n1133 240.244
R5846 gnd.n1188 gnd.n1141 240.244
R5847 gnd.n1191 gnd.n1142 240.244
R5848 gnd.n1152 gnd.n1151 240.244
R5849 gnd.n1193 gnd.n1159 240.244
R5850 gnd.n1171 gnd.n1160 240.244
R5851 gnd.n4565 gnd.n4446 240.244
R5852 gnd.n4565 gnd.n1559 240.244
R5853 gnd.n4561 gnd.n1559 240.244
R5854 gnd.n4561 gnd.n1552 240.244
R5855 gnd.n4558 gnd.n1552 240.244
R5856 gnd.n4558 gnd.n1544 240.244
R5857 gnd.n4555 gnd.n1544 240.244
R5858 gnd.n4555 gnd.n1535 240.244
R5859 gnd.n4552 gnd.n1535 240.244
R5860 gnd.n4552 gnd.n1527 240.244
R5861 gnd.n4549 gnd.n1527 240.244
R5862 gnd.n4549 gnd.n1520 240.244
R5863 gnd.n4546 gnd.n1520 240.244
R5864 gnd.n4546 gnd.n1512 240.244
R5865 gnd.n4543 gnd.n1512 240.244
R5866 gnd.n4543 gnd.n1503 240.244
R5867 gnd.n4540 gnd.n1503 240.244
R5868 gnd.n4540 gnd.n1494 240.244
R5869 gnd.n4537 gnd.n1494 240.244
R5870 gnd.n4537 gnd.n1485 240.244
R5871 gnd.n1485 gnd.n1477 240.244
R5872 gnd.n4862 gnd.n1477 240.244
R5873 gnd.n4862 gnd.n1459 240.244
R5874 gnd.n1473 gnd.n1459 240.244
R5875 gnd.n4872 gnd.n1473 240.244
R5876 gnd.n4872 gnd.n1449 240.244
R5877 gnd.n1449 gnd.n1442 240.244
R5878 gnd.n4902 gnd.n1442 240.244
R5879 gnd.n4902 gnd.n1394 240.244
R5880 gnd.n4905 gnd.n1394 240.244
R5881 gnd.n4905 gnd.n1405 240.244
R5882 gnd.n1411 gnd.n1405 240.244
R5883 gnd.n4912 gnd.n1411 240.244
R5884 gnd.n4913 gnd.n4912 240.244
R5885 gnd.n4913 gnd.n1424 240.244
R5886 gnd.n5196 gnd.n1424 240.244
R5887 gnd.n5196 gnd.n1379 240.244
R5888 gnd.n4918 gnd.n1379 240.244
R5889 gnd.n4918 gnd.n1370 240.244
R5890 gnd.n4919 gnd.n1370 240.244
R5891 gnd.n4919 gnd.n1362 240.244
R5892 gnd.n4922 gnd.n1362 240.244
R5893 gnd.n4922 gnd.n1353 240.244
R5894 gnd.n4923 gnd.n1353 240.244
R5895 gnd.n4923 gnd.n1344 240.244
R5896 gnd.n4926 gnd.n1344 240.244
R5897 gnd.n4926 gnd.n1335 240.244
R5898 gnd.n4927 gnd.n1335 240.244
R5899 gnd.n4927 gnd.n1327 240.244
R5900 gnd.n4930 gnd.n1327 240.244
R5901 gnd.n4930 gnd.n1318 240.244
R5902 gnd.n4931 gnd.n1318 240.244
R5903 gnd.n4931 gnd.n1309 240.244
R5904 gnd.n4934 gnd.n1309 240.244
R5905 gnd.n4934 gnd.n1300 240.244
R5906 gnd.n4935 gnd.n1300 240.244
R5907 gnd.n4935 gnd.n1292 240.244
R5908 gnd.n4938 gnd.n1292 240.244
R5909 gnd.n4938 gnd.n1283 240.244
R5910 gnd.n5119 gnd.n1283 240.244
R5911 gnd.n5119 gnd.n1273 240.244
R5912 gnd.n5153 gnd.n1273 240.244
R5913 gnd.n5153 gnd.n1173 240.244
R5914 gnd.n5742 gnd.n1173 240.244
R5915 gnd.n4472 gnd.n4470 240.244
R5916 gnd.n4478 gnd.n4464 240.244
R5917 gnd.n4482 gnd.n4480 240.244
R5918 gnd.n4488 gnd.n4460 240.244
R5919 gnd.n4492 gnd.n4490 240.244
R5920 gnd.n4498 gnd.n4456 240.244
R5921 gnd.n4502 gnd.n4500 240.244
R5922 gnd.n4508 gnd.n4452 240.244
R5923 gnd.n4511 gnd.n4510 240.244
R5924 gnd.n4759 gnd.n1560 240.244
R5925 gnd.n4765 gnd.n1560 240.244
R5926 gnd.n4765 gnd.n1549 240.244
R5927 gnd.n4775 gnd.n1549 240.244
R5928 gnd.n4775 gnd.n1545 240.244
R5929 gnd.n4781 gnd.n1545 240.244
R5930 gnd.n4781 gnd.n1532 240.244
R5931 gnd.n4791 gnd.n1532 240.244
R5932 gnd.n4791 gnd.n1528 240.244
R5933 gnd.n4797 gnd.n1528 240.244
R5934 gnd.n4797 gnd.n1517 240.244
R5935 gnd.n4807 gnd.n1517 240.244
R5936 gnd.n4807 gnd.n1513 240.244
R5937 gnd.n4813 gnd.n1513 240.244
R5938 gnd.n4813 gnd.n1500 240.244
R5939 gnd.n4823 gnd.n1500 240.244
R5940 gnd.n4823 gnd.n1495 240.244
R5941 gnd.n4837 gnd.n1495 240.244
R5942 gnd.n4837 gnd.n1496 240.244
R5943 gnd.n1496 gnd.n1486 240.244
R5944 gnd.n4832 gnd.n1486 240.244
R5945 gnd.n4832 gnd.n1461 240.244
R5946 gnd.n4878 gnd.n1461 240.244
R5947 gnd.n4878 gnd.n1462 240.244
R5948 gnd.n4874 gnd.n1462 240.244
R5949 gnd.n4874 gnd.n1450 240.244
R5950 gnd.n1470 gnd.n1450 240.244
R5951 gnd.n1470 gnd.n1396 240.244
R5952 gnd.n5237 gnd.n1396 240.244
R5953 gnd.n5237 gnd.n1397 240.244
R5954 gnd.n5233 gnd.n1397 240.244
R5955 gnd.n5233 gnd.n1403 240.244
R5956 gnd.n5208 gnd.n1403 240.244
R5957 gnd.n5208 gnd.n1426 240.244
R5958 gnd.n5214 gnd.n1426 240.244
R5959 gnd.n5214 gnd.n1376 240.244
R5960 gnd.n5247 gnd.n1376 240.244
R5961 gnd.n5247 gnd.n1372 240.244
R5962 gnd.n5253 gnd.n1372 240.244
R5963 gnd.n5253 gnd.n1359 240.244
R5964 gnd.n5263 gnd.n1359 240.244
R5965 gnd.n5263 gnd.n1355 240.244
R5966 gnd.n5269 gnd.n1355 240.244
R5967 gnd.n5269 gnd.n1341 240.244
R5968 gnd.n5279 gnd.n1341 240.244
R5969 gnd.n5279 gnd.n1337 240.244
R5970 gnd.n5285 gnd.n1337 240.244
R5971 gnd.n5285 gnd.n1324 240.244
R5972 gnd.n5295 gnd.n1324 240.244
R5973 gnd.n5295 gnd.n1320 240.244
R5974 gnd.n5301 gnd.n1320 240.244
R5975 gnd.n5301 gnd.n1306 240.244
R5976 gnd.n5311 gnd.n1306 240.244
R5977 gnd.n5311 gnd.n1302 240.244
R5978 gnd.n5317 gnd.n1302 240.244
R5979 gnd.n5317 gnd.n1289 240.244
R5980 gnd.n5327 gnd.n1289 240.244
R5981 gnd.n5327 gnd.n1285 240.244
R5982 gnd.n5333 gnd.n1285 240.244
R5983 gnd.n5333 gnd.n1270 240.244
R5984 gnd.n5345 gnd.n1270 240.244
R5985 gnd.n5345 gnd.n1266 240.244
R5986 gnd.n5663 gnd.n1266 240.244
R5987 gnd.n5663 gnd.n1178 240.244
R5988 gnd.n2842 gnd.n1784 240.244
R5989 gnd.n2836 gnd.n1784 240.244
R5990 gnd.n2836 gnd.n1788 240.244
R5991 gnd.n2832 gnd.n1788 240.244
R5992 gnd.n2832 gnd.n1790 240.244
R5993 gnd.n2828 gnd.n1790 240.244
R5994 gnd.n2828 gnd.n1795 240.244
R5995 gnd.n2824 gnd.n1795 240.244
R5996 gnd.n2824 gnd.n1797 240.244
R5997 gnd.n2820 gnd.n1797 240.244
R5998 gnd.n2820 gnd.n1803 240.244
R5999 gnd.n2816 gnd.n1803 240.244
R6000 gnd.n2816 gnd.n1805 240.244
R6001 gnd.n2812 gnd.n1805 240.244
R6002 gnd.n2812 gnd.n1811 240.244
R6003 gnd.n2808 gnd.n1811 240.244
R6004 gnd.n2808 gnd.n1813 240.244
R6005 gnd.n2804 gnd.n1813 240.244
R6006 gnd.n2804 gnd.n1819 240.244
R6007 gnd.n2800 gnd.n1819 240.244
R6008 gnd.n2800 gnd.n1821 240.244
R6009 gnd.n2796 gnd.n1821 240.244
R6010 gnd.n2796 gnd.n1827 240.244
R6011 gnd.n2792 gnd.n1827 240.244
R6012 gnd.n2792 gnd.n1829 240.244
R6013 gnd.n2788 gnd.n1829 240.244
R6014 gnd.n2788 gnd.n1835 240.244
R6015 gnd.n2784 gnd.n1835 240.244
R6016 gnd.n2784 gnd.n1837 240.244
R6017 gnd.n2780 gnd.n1837 240.244
R6018 gnd.n2780 gnd.n1843 240.244
R6019 gnd.n2776 gnd.n1843 240.244
R6020 gnd.n2776 gnd.n1845 240.244
R6021 gnd.n2772 gnd.n1845 240.244
R6022 gnd.n2772 gnd.n1851 240.244
R6023 gnd.n2768 gnd.n1851 240.244
R6024 gnd.n2768 gnd.n1853 240.244
R6025 gnd.n2764 gnd.n1853 240.244
R6026 gnd.n2764 gnd.n1859 240.244
R6027 gnd.n2760 gnd.n1859 240.244
R6028 gnd.n2760 gnd.n1861 240.244
R6029 gnd.n2756 gnd.n1861 240.244
R6030 gnd.n2756 gnd.n1867 240.244
R6031 gnd.n2752 gnd.n1867 240.244
R6032 gnd.n2752 gnd.n1869 240.244
R6033 gnd.n2748 gnd.n1869 240.244
R6034 gnd.n2748 gnd.n1875 240.244
R6035 gnd.n2744 gnd.n1875 240.244
R6036 gnd.n2744 gnd.n1877 240.244
R6037 gnd.n2740 gnd.n1877 240.244
R6038 gnd.n2740 gnd.n1883 240.244
R6039 gnd.n2736 gnd.n1883 240.244
R6040 gnd.n2736 gnd.n1885 240.244
R6041 gnd.n2732 gnd.n1885 240.244
R6042 gnd.n2732 gnd.n1891 240.244
R6043 gnd.n2728 gnd.n1891 240.244
R6044 gnd.n2728 gnd.n1893 240.244
R6045 gnd.n2724 gnd.n1893 240.244
R6046 gnd.n2724 gnd.n1899 240.244
R6047 gnd.n2720 gnd.n1899 240.244
R6048 gnd.n2720 gnd.n1901 240.244
R6049 gnd.n2716 gnd.n1901 240.244
R6050 gnd.n2716 gnd.n1907 240.244
R6051 gnd.n2712 gnd.n1907 240.244
R6052 gnd.n2712 gnd.n1909 240.244
R6053 gnd.n2708 gnd.n1909 240.244
R6054 gnd.n2708 gnd.n1915 240.244
R6055 gnd.n2704 gnd.n1915 240.244
R6056 gnd.n2704 gnd.n1917 240.244
R6057 gnd.n2700 gnd.n1917 240.244
R6058 gnd.n2700 gnd.n1923 240.244
R6059 gnd.n2696 gnd.n1923 240.244
R6060 gnd.n2696 gnd.n1925 240.244
R6061 gnd.n2692 gnd.n1925 240.244
R6062 gnd.n2692 gnd.n1931 240.244
R6063 gnd.n2688 gnd.n1931 240.244
R6064 gnd.n2688 gnd.n1933 240.244
R6065 gnd.n2684 gnd.n1933 240.244
R6066 gnd.n2684 gnd.n1939 240.244
R6067 gnd.n2680 gnd.n1939 240.244
R6068 gnd.n2680 gnd.n1941 240.244
R6069 gnd.n2676 gnd.n1941 240.244
R6070 gnd.n2676 gnd.n1947 240.244
R6071 gnd.n2672 gnd.n1947 240.244
R6072 gnd.n2672 gnd.n1949 240.244
R6073 gnd.n2668 gnd.n1949 240.244
R6074 gnd.n2668 gnd.n1955 240.244
R6075 gnd.n2664 gnd.n1955 240.244
R6076 gnd.n2664 gnd.n1957 240.244
R6077 gnd.n2660 gnd.n1957 240.244
R6078 gnd.n2660 gnd.n1963 240.244
R6079 gnd.n2656 gnd.n1963 240.244
R6080 gnd.n2656 gnd.n1965 240.244
R6081 gnd.n2652 gnd.n1965 240.244
R6082 gnd.n2652 gnd.n1971 240.244
R6083 gnd.n2648 gnd.n1971 240.244
R6084 gnd.n2648 gnd.n1973 240.244
R6085 gnd.n2644 gnd.n1973 240.244
R6086 gnd.n2644 gnd.n1979 240.244
R6087 gnd.n2640 gnd.n1979 240.244
R6088 gnd.n2640 gnd.n1981 240.244
R6089 gnd.n2636 gnd.n1981 240.244
R6090 gnd.n2636 gnd.n1987 240.244
R6091 gnd.n2632 gnd.n1987 240.244
R6092 gnd.n2632 gnd.n1989 240.244
R6093 gnd.n2628 gnd.n1989 240.244
R6094 gnd.n2628 gnd.n1995 240.244
R6095 gnd.n2624 gnd.n1995 240.244
R6096 gnd.n2624 gnd.n1997 240.244
R6097 gnd.n2620 gnd.n1997 240.244
R6098 gnd.n2620 gnd.n2003 240.244
R6099 gnd.n2616 gnd.n2003 240.244
R6100 gnd.n2616 gnd.n2005 240.244
R6101 gnd.n2612 gnd.n2005 240.244
R6102 gnd.n2612 gnd.n2011 240.244
R6103 gnd.n2608 gnd.n2011 240.244
R6104 gnd.n2608 gnd.n2013 240.244
R6105 gnd.n2604 gnd.n2013 240.244
R6106 gnd.n2604 gnd.n2019 240.244
R6107 gnd.n2600 gnd.n2019 240.244
R6108 gnd.n2600 gnd.n2021 240.244
R6109 gnd.n2596 gnd.n2021 240.244
R6110 gnd.n2596 gnd.n2027 240.244
R6111 gnd.n2592 gnd.n2027 240.244
R6112 gnd.n2592 gnd.n2029 240.244
R6113 gnd.n2588 gnd.n2029 240.244
R6114 gnd.n2588 gnd.n2035 240.244
R6115 gnd.n2584 gnd.n2035 240.244
R6116 gnd.n2584 gnd.n2037 240.244
R6117 gnd.n2580 gnd.n2037 240.244
R6118 gnd.n2580 gnd.n2043 240.244
R6119 gnd.n2576 gnd.n2043 240.244
R6120 gnd.n2576 gnd.n2045 240.244
R6121 gnd.n2572 gnd.n2045 240.244
R6122 gnd.n2572 gnd.n2051 240.244
R6123 gnd.n2568 gnd.n2051 240.244
R6124 gnd.n2568 gnd.n2053 240.244
R6125 gnd.n2564 gnd.n2053 240.244
R6126 gnd.n2564 gnd.n2059 240.244
R6127 gnd.n2560 gnd.n2059 240.244
R6128 gnd.n2560 gnd.n2061 240.244
R6129 gnd.n2556 gnd.n2061 240.244
R6130 gnd.n2556 gnd.n2067 240.244
R6131 gnd.n2552 gnd.n2067 240.244
R6132 gnd.n2552 gnd.n2069 240.244
R6133 gnd.n2548 gnd.n2069 240.244
R6134 gnd.n2548 gnd.n2075 240.244
R6135 gnd.n2544 gnd.n2075 240.244
R6136 gnd.n2544 gnd.n2077 240.244
R6137 gnd.n2540 gnd.n2077 240.244
R6138 gnd.n2540 gnd.n2083 240.244
R6139 gnd.n2536 gnd.n2083 240.244
R6140 gnd.n2536 gnd.n2085 240.244
R6141 gnd.n2532 gnd.n2085 240.244
R6142 gnd.n2532 gnd.n2091 240.244
R6143 gnd.n2528 gnd.n2091 240.244
R6144 gnd.n2528 gnd.n2093 240.244
R6145 gnd.n2524 gnd.n2093 240.244
R6146 gnd.n2524 gnd.n2099 240.244
R6147 gnd.n2520 gnd.n2099 240.244
R6148 gnd.n2520 gnd.n2101 240.244
R6149 gnd.n2516 gnd.n2101 240.244
R6150 gnd.n2516 gnd.n2107 240.244
R6151 gnd.n2512 gnd.n2107 240.244
R6152 gnd.n2512 gnd.n2109 240.244
R6153 gnd.n2508 gnd.n2109 240.244
R6154 gnd.n2508 gnd.n2115 240.244
R6155 gnd.n2504 gnd.n2115 240.244
R6156 gnd.n2504 gnd.n2117 240.244
R6157 gnd.n2500 gnd.n2117 240.244
R6158 gnd.n2500 gnd.n2123 240.244
R6159 gnd.n2496 gnd.n2123 240.244
R6160 gnd.n2496 gnd.n2125 240.244
R6161 gnd.n2492 gnd.n2125 240.244
R6162 gnd.n2492 gnd.n2131 240.244
R6163 gnd.n2488 gnd.n2131 240.244
R6164 gnd.n2488 gnd.n2133 240.244
R6165 gnd.n2484 gnd.n2133 240.244
R6166 gnd.n2484 gnd.n2139 240.244
R6167 gnd.n2480 gnd.n2139 240.244
R6168 gnd.n2480 gnd.n2141 240.244
R6169 gnd.n2474 gnd.n2146 240.244
R6170 gnd.n2470 gnd.n2146 240.244
R6171 gnd.n2470 gnd.n2148 240.244
R6172 gnd.n2466 gnd.n2148 240.244
R6173 gnd.n2466 gnd.n2153 240.244
R6174 gnd.n2462 gnd.n2153 240.244
R6175 gnd.n2462 gnd.n2155 240.244
R6176 gnd.n2458 gnd.n2155 240.244
R6177 gnd.n2458 gnd.n2161 240.244
R6178 gnd.n2454 gnd.n2161 240.244
R6179 gnd.n2454 gnd.n2163 240.244
R6180 gnd.n2450 gnd.n2163 240.244
R6181 gnd.n2450 gnd.n2169 240.244
R6182 gnd.n2446 gnd.n2169 240.244
R6183 gnd.n2446 gnd.n2171 240.244
R6184 gnd.n2442 gnd.n2171 240.244
R6185 gnd.n2442 gnd.n2177 240.244
R6186 gnd.n2438 gnd.n2177 240.244
R6187 gnd.n2438 gnd.n2179 240.244
R6188 gnd.n2434 gnd.n2179 240.244
R6189 gnd.n2434 gnd.n2185 240.244
R6190 gnd.n2430 gnd.n2185 240.244
R6191 gnd.n2430 gnd.n2187 240.244
R6192 gnd.n2426 gnd.n2187 240.244
R6193 gnd.n2426 gnd.n2193 240.244
R6194 gnd.n2422 gnd.n2193 240.244
R6195 gnd.n2422 gnd.n2195 240.244
R6196 gnd.n2418 gnd.n2195 240.244
R6197 gnd.n2418 gnd.n2201 240.244
R6198 gnd.n2414 gnd.n2201 240.244
R6199 gnd.n2414 gnd.n2203 240.244
R6200 gnd.n2410 gnd.n2203 240.244
R6201 gnd.n2410 gnd.n2209 240.244
R6202 gnd.n2406 gnd.n2209 240.244
R6203 gnd.n2406 gnd.n2211 240.244
R6204 gnd.n2402 gnd.n2211 240.244
R6205 gnd.n2402 gnd.n2217 240.244
R6206 gnd.n2398 gnd.n2217 240.244
R6207 gnd.n2398 gnd.n2219 240.244
R6208 gnd.n2394 gnd.n2219 240.244
R6209 gnd.n2394 gnd.n2225 240.244
R6210 gnd.n2390 gnd.n2225 240.244
R6211 gnd.n2390 gnd.n2227 240.244
R6212 gnd.n2386 gnd.n2227 240.244
R6213 gnd.n2386 gnd.n2233 240.244
R6214 gnd.n2382 gnd.n2233 240.244
R6215 gnd.n2382 gnd.n2235 240.244
R6216 gnd.n2378 gnd.n2235 240.244
R6217 gnd.n2378 gnd.n2241 240.244
R6218 gnd.n2374 gnd.n2241 240.244
R6219 gnd.n2374 gnd.n2243 240.244
R6220 gnd.n2370 gnd.n2243 240.244
R6221 gnd.n2370 gnd.n2249 240.244
R6222 gnd.n2366 gnd.n2249 240.244
R6223 gnd.n2366 gnd.n2251 240.244
R6224 gnd.n2362 gnd.n2251 240.244
R6225 gnd.n2362 gnd.n2257 240.244
R6226 gnd.n2358 gnd.n2257 240.244
R6227 gnd.n2358 gnd.n2259 240.244
R6228 gnd.n2354 gnd.n2259 240.244
R6229 gnd.n2354 gnd.n2265 240.244
R6230 gnd.n2350 gnd.n2265 240.244
R6231 gnd.n2350 gnd.n2267 240.244
R6232 gnd.n2346 gnd.n2267 240.244
R6233 gnd.n2346 gnd.n2273 240.244
R6234 gnd.n2342 gnd.n2273 240.244
R6235 gnd.n2342 gnd.n2275 240.244
R6236 gnd.n2338 gnd.n2275 240.244
R6237 gnd.n2338 gnd.n2281 240.244
R6238 gnd.n2334 gnd.n2281 240.244
R6239 gnd.n2334 gnd.n2283 240.244
R6240 gnd.n2330 gnd.n2283 240.244
R6241 gnd.n2330 gnd.n2289 240.244
R6242 gnd.n2326 gnd.n2289 240.244
R6243 gnd.n2326 gnd.n2291 240.244
R6244 gnd.n2322 gnd.n2291 240.244
R6245 gnd.n2322 gnd.n2297 240.244
R6246 gnd.n2318 gnd.n2297 240.244
R6247 gnd.n2318 gnd.n2299 240.244
R6248 gnd.n2314 gnd.n2299 240.244
R6249 gnd.n2314 gnd.n2305 240.244
R6250 gnd.n2310 gnd.n2305 240.244
R6251 gnd.n2310 gnd.n335 240.244
R6252 gnd.n7563 gnd.n335 240.244
R6253 gnd.n3053 gnd.n1413 240.244
R6254 gnd.n5225 gnd.n1413 240.244
R6255 gnd.n5225 gnd.n1414 240.244
R6256 gnd.n5221 gnd.n1414 240.244
R6257 gnd.n5221 gnd.n1420 240.244
R6258 gnd.n4965 gnd.n1420 240.244
R6259 gnd.n4965 gnd.n4961 240.244
R6260 gnd.n4991 gnd.n4961 240.244
R6261 gnd.n4991 gnd.n4962 240.244
R6262 gnd.n4987 gnd.n4962 240.244
R6263 gnd.n4987 gnd.n4986 240.244
R6264 gnd.n4986 gnd.n4985 240.244
R6265 gnd.n4985 gnd.n4973 240.244
R6266 gnd.n4981 gnd.n4973 240.244
R6267 gnd.n4981 gnd.n4953 240.244
R6268 gnd.n5035 gnd.n4953 240.244
R6269 gnd.n5036 gnd.n5035 240.244
R6270 gnd.n5037 gnd.n5036 240.244
R6271 gnd.n5037 gnd.n4949 240.244
R6272 gnd.n5043 gnd.n4949 240.244
R6273 gnd.n5044 gnd.n5043 240.244
R6274 gnd.n5045 gnd.n5044 240.244
R6275 gnd.n5045 gnd.n4944 240.244
R6276 gnd.n5095 gnd.n4944 240.244
R6277 gnd.n5095 gnd.n4945 240.244
R6278 gnd.n5091 gnd.n4945 240.244
R6279 gnd.n5091 gnd.n5090 240.244
R6280 gnd.n5090 gnd.n5089 240.244
R6281 gnd.n5089 gnd.n5053 240.244
R6282 gnd.n5085 gnd.n5053 240.244
R6283 gnd.n5085 gnd.n5084 240.244
R6284 gnd.n5084 gnd.n5083 240.244
R6285 gnd.n5083 gnd.n5059 240.244
R6286 gnd.n5079 gnd.n5059 240.244
R6287 gnd.n5079 gnd.n5078 240.244
R6288 gnd.n5078 gnd.n5076 240.244
R6289 gnd.n5076 gnd.n5065 240.244
R6290 gnd.n5070 gnd.n5065 240.244
R6291 gnd.n5070 gnd.n1096 240.244
R6292 gnd.n5801 gnd.n1096 240.244
R6293 gnd.n5801 gnd.n1092 240.244
R6294 gnd.n5807 gnd.n1092 240.244
R6295 gnd.n5807 gnd.n1083 240.244
R6296 gnd.n5817 gnd.n1083 240.244
R6297 gnd.n5817 gnd.n1079 240.244
R6298 gnd.n5823 gnd.n1079 240.244
R6299 gnd.n5823 gnd.n1069 240.244
R6300 gnd.n5833 gnd.n1069 240.244
R6301 gnd.n5833 gnd.n1065 240.244
R6302 gnd.n5839 gnd.n1065 240.244
R6303 gnd.n5839 gnd.n1055 240.244
R6304 gnd.n5849 gnd.n1055 240.244
R6305 gnd.n5849 gnd.n1051 240.244
R6306 gnd.n5855 gnd.n1051 240.244
R6307 gnd.n5855 gnd.n1040 240.244
R6308 gnd.n5865 gnd.n1040 240.244
R6309 gnd.n5865 gnd.n1036 240.244
R6310 gnd.n5871 gnd.n1036 240.244
R6311 gnd.n5871 gnd.n1026 240.244
R6312 gnd.n5881 gnd.n1026 240.244
R6313 gnd.n5881 gnd.n1021 240.244
R6314 gnd.n5889 gnd.n1021 240.244
R6315 gnd.n5889 gnd.n1022 240.244
R6316 gnd.n1022 gnd.n986 240.244
R6317 gnd.n5979 gnd.n986 240.244
R6318 gnd.n5979 gnd.n982 240.244
R6319 gnd.n5985 gnd.n982 240.244
R6320 gnd.n5985 gnd.n970 240.244
R6321 gnd.n5995 gnd.n970 240.244
R6322 gnd.n5995 gnd.n966 240.244
R6323 gnd.n6001 gnd.n966 240.244
R6324 gnd.n6001 gnd.n952 240.244
R6325 gnd.n6014 gnd.n952 240.244
R6326 gnd.n6014 gnd.n948 240.244
R6327 gnd.n6020 gnd.n948 240.244
R6328 gnd.n6020 gnd.n916 240.244
R6329 gnd.n6070 gnd.n916 240.244
R6330 gnd.n6070 gnd.n911 240.244
R6331 gnd.n6078 gnd.n911 240.244
R6332 gnd.n6078 gnd.n912 240.244
R6333 gnd.n912 gnd.n882 240.244
R6334 gnd.n6834 gnd.n882 240.244
R6335 gnd.n6834 gnd.n878 240.244
R6336 gnd.n6840 gnd.n878 240.244
R6337 gnd.n6840 gnd.n867 240.244
R6338 gnd.n6850 gnd.n867 240.244
R6339 gnd.n6850 gnd.n863 240.244
R6340 gnd.n6856 gnd.n863 240.244
R6341 gnd.n6856 gnd.n851 240.244
R6342 gnd.n6866 gnd.n851 240.244
R6343 gnd.n6866 gnd.n847 240.244
R6344 gnd.n6872 gnd.n847 240.244
R6345 gnd.n6872 gnd.n835 240.244
R6346 gnd.n6882 gnd.n835 240.244
R6347 gnd.n6882 gnd.n831 240.244
R6348 gnd.n6888 gnd.n831 240.244
R6349 gnd.n6888 gnd.n819 240.244
R6350 gnd.n6898 gnd.n819 240.244
R6351 gnd.n6898 gnd.n815 240.244
R6352 gnd.n6904 gnd.n815 240.244
R6353 gnd.n6904 gnd.n804 240.244
R6354 gnd.n6914 gnd.n804 240.244
R6355 gnd.n6914 gnd.n800 240.244
R6356 gnd.n6920 gnd.n800 240.244
R6357 gnd.n6920 gnd.n788 240.244
R6358 gnd.n6930 gnd.n788 240.244
R6359 gnd.n6930 gnd.n784 240.244
R6360 gnd.n6936 gnd.n784 240.244
R6361 gnd.n6936 gnd.n772 240.244
R6362 gnd.n6946 gnd.n772 240.244
R6363 gnd.n6946 gnd.n768 240.244
R6364 gnd.n6952 gnd.n768 240.244
R6365 gnd.n6952 gnd.n756 240.244
R6366 gnd.n6962 gnd.n756 240.244
R6367 gnd.n6962 gnd.n752 240.244
R6368 gnd.n6968 gnd.n752 240.244
R6369 gnd.n6968 gnd.n740 240.244
R6370 gnd.n6978 gnd.n740 240.244
R6371 gnd.n6978 gnd.n736 240.244
R6372 gnd.n6984 gnd.n736 240.244
R6373 gnd.n6984 gnd.n725 240.244
R6374 gnd.n6994 gnd.n725 240.244
R6375 gnd.n6994 gnd.n721 240.244
R6376 gnd.n7000 gnd.n721 240.244
R6377 gnd.n7000 gnd.n711 240.244
R6378 gnd.n7010 gnd.n711 240.244
R6379 gnd.n7010 gnd.n707 240.244
R6380 gnd.n7016 gnd.n707 240.244
R6381 gnd.n7016 gnd.n697 240.244
R6382 gnd.n7026 gnd.n697 240.244
R6383 gnd.n7026 gnd.n693 240.244
R6384 gnd.n7032 gnd.n693 240.244
R6385 gnd.n7032 gnd.n683 240.244
R6386 gnd.n7042 gnd.n683 240.244
R6387 gnd.n7042 gnd.n679 240.244
R6388 gnd.n7048 gnd.n679 240.244
R6389 gnd.n7048 gnd.n668 240.244
R6390 gnd.n7059 gnd.n668 240.244
R6391 gnd.n7059 gnd.n663 240.244
R6392 gnd.n7067 gnd.n663 240.244
R6393 gnd.n7067 gnd.n664 240.244
R6394 gnd.n664 gnd.n638 240.244
R6395 gnd.n7079 gnd.n638 240.244
R6396 gnd.n7079 gnd.n634 240.244
R6397 gnd.n7085 gnd.n634 240.244
R6398 gnd.n7086 gnd.n7085 240.244
R6399 gnd.n7087 gnd.n7086 240.244
R6400 gnd.n7087 gnd.n630 240.244
R6401 gnd.n7093 gnd.n630 240.244
R6402 gnd.n7094 gnd.n7093 240.244
R6403 gnd.n7095 gnd.n7094 240.244
R6404 gnd.n7095 gnd.n626 240.244
R6405 gnd.n7101 gnd.n626 240.244
R6406 gnd.n7102 gnd.n7101 240.244
R6407 gnd.n7103 gnd.n7102 240.244
R6408 gnd.n7103 gnd.n621 240.244
R6409 gnd.n7126 gnd.n621 240.244
R6410 gnd.n7126 gnd.n622 240.244
R6411 gnd.n7122 gnd.n622 240.244
R6412 gnd.n7122 gnd.n7121 240.244
R6413 gnd.n7121 gnd.n7120 240.244
R6414 gnd.n7120 gnd.n7111 240.244
R6415 gnd.n7111 gnd.n420 240.244
R6416 gnd.n7343 gnd.n420 240.244
R6417 gnd.n7344 gnd.n7343 240.244
R6418 gnd.n7345 gnd.n7344 240.244
R6419 gnd.n7345 gnd.n415 240.244
R6420 gnd.n7380 gnd.n415 240.244
R6421 gnd.n7380 gnd.n416 240.244
R6422 gnd.n7376 gnd.n416 240.244
R6423 gnd.n7376 gnd.n7375 240.244
R6424 gnd.n7375 gnd.n7374 240.244
R6425 gnd.n7374 gnd.n7353 240.244
R6426 gnd.n7370 gnd.n7353 240.244
R6427 gnd.n7370 gnd.n7369 240.244
R6428 gnd.n7369 gnd.n7368 240.244
R6429 gnd.n7368 gnd.n7359 240.244
R6430 gnd.n7364 gnd.n7359 240.244
R6431 gnd.n7364 gnd.n342 240.244
R6432 gnd.n7557 gnd.n342 240.244
R6433 gnd.n7557 gnd.n336 240.244
R6434 gnd.n2846 gnd.n1782 240.244
R6435 gnd.n2846 gnd.n1778 240.244
R6436 gnd.n2852 gnd.n1778 240.244
R6437 gnd.n2852 gnd.n1776 240.244
R6438 gnd.n2856 gnd.n1776 240.244
R6439 gnd.n2856 gnd.n1772 240.244
R6440 gnd.n2862 gnd.n1772 240.244
R6441 gnd.n2862 gnd.n1770 240.244
R6442 gnd.n2866 gnd.n1770 240.244
R6443 gnd.n2866 gnd.n1766 240.244
R6444 gnd.n2872 gnd.n1766 240.244
R6445 gnd.n2872 gnd.n1764 240.244
R6446 gnd.n2876 gnd.n1764 240.244
R6447 gnd.n2876 gnd.n1760 240.244
R6448 gnd.n2882 gnd.n1760 240.244
R6449 gnd.n2882 gnd.n1758 240.244
R6450 gnd.n2886 gnd.n1758 240.244
R6451 gnd.n2886 gnd.n1754 240.244
R6452 gnd.n2892 gnd.n1754 240.244
R6453 gnd.n2892 gnd.n1752 240.244
R6454 gnd.n2896 gnd.n1752 240.244
R6455 gnd.n2896 gnd.n1748 240.244
R6456 gnd.n2902 gnd.n1748 240.244
R6457 gnd.n2902 gnd.n1746 240.244
R6458 gnd.n2906 gnd.n1746 240.244
R6459 gnd.n2906 gnd.n1742 240.244
R6460 gnd.n2912 gnd.n1742 240.244
R6461 gnd.n2912 gnd.n1740 240.244
R6462 gnd.n2916 gnd.n1740 240.244
R6463 gnd.n2916 gnd.n1736 240.244
R6464 gnd.n2922 gnd.n1736 240.244
R6465 gnd.n2922 gnd.n1734 240.244
R6466 gnd.n2926 gnd.n1734 240.244
R6467 gnd.n2926 gnd.n1730 240.244
R6468 gnd.n2932 gnd.n1730 240.244
R6469 gnd.n2932 gnd.n1728 240.244
R6470 gnd.n2936 gnd.n1728 240.244
R6471 gnd.n2936 gnd.n1724 240.244
R6472 gnd.n2942 gnd.n1724 240.244
R6473 gnd.n2942 gnd.n1722 240.244
R6474 gnd.n2946 gnd.n1722 240.244
R6475 gnd.n2946 gnd.n1718 240.244
R6476 gnd.n2952 gnd.n1718 240.244
R6477 gnd.n2952 gnd.n1716 240.244
R6478 gnd.n2956 gnd.n1716 240.244
R6479 gnd.n2956 gnd.n1712 240.244
R6480 gnd.n2962 gnd.n1712 240.244
R6481 gnd.n2962 gnd.n1710 240.244
R6482 gnd.n2966 gnd.n1710 240.244
R6483 gnd.n2966 gnd.n1706 240.244
R6484 gnd.n2972 gnd.n1706 240.244
R6485 gnd.n2972 gnd.n1704 240.244
R6486 gnd.n2976 gnd.n1704 240.244
R6487 gnd.n2976 gnd.n1700 240.244
R6488 gnd.n2982 gnd.n1700 240.244
R6489 gnd.n2982 gnd.n1698 240.244
R6490 gnd.n2986 gnd.n1698 240.244
R6491 gnd.n2986 gnd.n1694 240.244
R6492 gnd.n2992 gnd.n1694 240.244
R6493 gnd.n2992 gnd.n1692 240.244
R6494 gnd.n2996 gnd.n1692 240.244
R6495 gnd.n2996 gnd.n1688 240.244
R6496 gnd.n3002 gnd.n1688 240.244
R6497 gnd.n3002 gnd.n1686 240.244
R6498 gnd.n3006 gnd.n1686 240.244
R6499 gnd.n3006 gnd.n1682 240.244
R6500 gnd.n3012 gnd.n1682 240.244
R6501 gnd.n3012 gnd.n1680 240.244
R6502 gnd.n3016 gnd.n1680 240.244
R6503 gnd.n3016 gnd.n1676 240.244
R6504 gnd.n3022 gnd.n1676 240.244
R6505 gnd.n3022 gnd.n1674 240.244
R6506 gnd.n3026 gnd.n1674 240.244
R6507 gnd.n3026 gnd.n1670 240.244
R6508 gnd.n3032 gnd.n1670 240.244
R6509 gnd.n3032 gnd.n1668 240.244
R6510 gnd.n3036 gnd.n1668 240.244
R6511 gnd.n3036 gnd.n1664 240.244
R6512 gnd.n3042 gnd.n1664 240.244
R6513 gnd.n3042 gnd.n1662 240.244
R6514 gnd.n3046 gnd.n1662 240.244
R6515 gnd.n3046 gnd.n1657 240.244
R6516 gnd.n3059 gnd.n1657 240.244
R6517 gnd.n3059 gnd.n1658 240.244
R6518 gnd.n5358 gnd.n1098 240.244
R6519 gnd.n5358 gnd.n1091 240.244
R6520 gnd.n5359 gnd.n1091 240.244
R6521 gnd.n5359 gnd.n1085 240.244
R6522 gnd.n5362 gnd.n1085 240.244
R6523 gnd.n5362 gnd.n1078 240.244
R6524 gnd.n5363 gnd.n1078 240.244
R6525 gnd.n5363 gnd.n1071 240.244
R6526 gnd.n5366 gnd.n1071 240.244
R6527 gnd.n5366 gnd.n1063 240.244
R6528 gnd.n5367 gnd.n1063 240.244
R6529 gnd.n5367 gnd.n1056 240.244
R6530 gnd.n5370 gnd.n1056 240.244
R6531 gnd.n5370 gnd.n1049 240.244
R6532 gnd.n5371 gnd.n1049 240.244
R6533 gnd.n5371 gnd.n1041 240.244
R6534 gnd.n5375 gnd.n1041 240.244
R6535 gnd.n5375 gnd.n1034 240.244
R6536 gnd.n5398 gnd.n1034 240.244
R6537 gnd.n5398 gnd.n1027 240.244
R6538 gnd.n5622 gnd.n1027 240.244
R6539 gnd.n5622 gnd.n1019 240.244
R6540 gnd.n1019 gnd.n1009 240.244
R6541 gnd.n5900 gnd.n1009 240.244
R6542 gnd.n5900 gnd.n988 240.244
R6543 gnd.n1006 gnd.n988 240.244
R6544 gnd.n1006 gnd.n980 240.244
R6545 gnd.n5908 gnd.n980 240.244
R6546 gnd.n5908 gnd.n972 240.244
R6547 gnd.n5961 gnd.n972 240.244
R6548 gnd.n5961 gnd.n964 240.244
R6549 gnd.n5913 gnd.n964 240.244
R6550 gnd.n5913 gnd.n954 240.244
R6551 gnd.n5945 gnd.n954 240.244
R6552 gnd.n5945 gnd.n946 240.244
R6553 gnd.n5948 gnd.n946 240.244
R6554 gnd.n5948 gnd.n918 240.244
R6555 gnd.n918 gnd.n907 240.244
R6556 gnd.n6080 gnd.n907 240.244
R6557 gnd.n6080 gnd.n908 240.244
R6558 gnd.n908 gnd.n904 240.244
R6559 gnd.n904 gnd.n885 240.244
R6560 gnd.n6087 gnd.n885 240.244
R6561 gnd.n6087 gnd.n876 240.244
R6562 gnd.n6819 gnd.n876 240.244
R6563 gnd.n6819 gnd.n869 240.244
R6564 gnd.n6092 gnd.n869 240.244
R6565 gnd.n6092 gnd.n861 240.244
R6566 gnd.n6093 gnd.n861 240.244
R6567 gnd.n6093 gnd.n853 240.244
R6568 gnd.n6096 gnd.n853 240.244
R6569 gnd.n6096 gnd.n845 240.244
R6570 gnd.n6097 gnd.n845 240.244
R6571 gnd.n6097 gnd.n837 240.244
R6572 gnd.n6100 gnd.n837 240.244
R6573 gnd.n6100 gnd.n829 240.244
R6574 gnd.n6101 gnd.n829 240.244
R6575 gnd.n6101 gnd.n821 240.244
R6576 gnd.n6104 gnd.n821 240.244
R6577 gnd.n6104 gnd.n813 240.244
R6578 gnd.n6105 gnd.n813 240.244
R6579 gnd.n6105 gnd.n806 240.244
R6580 gnd.n6108 gnd.n806 240.244
R6581 gnd.n6108 gnd.n798 240.244
R6582 gnd.n6109 gnd.n798 240.244
R6583 gnd.n6109 gnd.n790 240.244
R6584 gnd.n6112 gnd.n790 240.244
R6585 gnd.n6112 gnd.n782 240.244
R6586 gnd.n6113 gnd.n782 240.244
R6587 gnd.n6113 gnd.n774 240.244
R6588 gnd.n6116 gnd.n774 240.244
R6589 gnd.n6116 gnd.n766 240.244
R6590 gnd.n6117 gnd.n766 240.244
R6591 gnd.n6117 gnd.n758 240.244
R6592 gnd.n6120 gnd.n758 240.244
R6593 gnd.n6120 gnd.n749 240.244
R6594 gnd.n6121 gnd.n749 240.244
R6595 gnd.n6121 gnd.n741 240.244
R6596 gnd.n6124 gnd.n741 240.244
R6597 gnd.n6124 gnd.n734 240.244
R6598 gnd.n6574 gnd.n734 240.244
R6599 gnd.n6574 gnd.n727 240.244
R6600 gnd.n6577 gnd.n727 240.244
R6601 gnd.n6577 gnd.n719 240.244
R6602 gnd.n6579 gnd.n719 240.244
R6603 gnd.n6579 gnd.n712 240.244
R6604 gnd.n6582 gnd.n712 240.244
R6605 gnd.n6582 gnd.n705 240.244
R6606 gnd.n6583 gnd.n705 240.244
R6607 gnd.n6583 gnd.n698 240.244
R6608 gnd.n6586 gnd.n698 240.244
R6609 gnd.n6586 gnd.n692 240.244
R6610 gnd.n6587 gnd.n692 240.244
R6611 gnd.n6587 gnd.n685 240.244
R6612 gnd.n6590 gnd.n685 240.244
R6613 gnd.n6590 gnd.n678 240.244
R6614 gnd.n6591 gnd.n678 240.244
R6615 gnd.n6591 gnd.n670 240.244
R6616 gnd.n6594 gnd.n670 240.244
R6617 gnd.n6594 gnd.n661 240.244
R6618 gnd.n6733 gnd.n661 240.244
R6619 gnd.n1118 gnd.n1117 240.244
R6620 gnd.n1128 gnd.n1117 240.244
R6621 gnd.n1130 gnd.n1129 240.244
R6622 gnd.n1138 gnd.n1137 240.244
R6623 gnd.n1146 gnd.n1145 240.244
R6624 gnd.n1148 gnd.n1147 240.244
R6625 gnd.n1156 gnd.n1155 240.244
R6626 gnd.n1166 gnd.n1165 240.244
R6627 gnd.n1168 gnd.n1167 240.244
R6628 gnd.n5123 gnd.n5122 240.244
R6629 gnd.n5125 gnd.n5124 240.244
R6630 gnd.n5129 gnd.n5128 240.244
R6631 gnd.n5135 gnd.n5130 240.244
R6632 gnd.n5793 gnd.n1103 240.244
R6633 gnd.n5799 gnd.n1090 240.244
R6634 gnd.n5809 gnd.n1090 240.244
R6635 gnd.n5809 gnd.n1086 240.244
R6636 gnd.n5815 gnd.n1086 240.244
R6637 gnd.n5815 gnd.n1076 240.244
R6638 gnd.n5825 gnd.n1076 240.244
R6639 gnd.n5825 gnd.n1072 240.244
R6640 gnd.n5831 gnd.n1072 240.244
R6641 gnd.n5831 gnd.n1061 240.244
R6642 gnd.n5841 gnd.n1061 240.244
R6643 gnd.n5841 gnd.n1057 240.244
R6644 gnd.n5847 gnd.n1057 240.244
R6645 gnd.n5847 gnd.n1047 240.244
R6646 gnd.n5857 gnd.n1047 240.244
R6647 gnd.n5857 gnd.n1043 240.244
R6648 gnd.n5863 gnd.n1043 240.244
R6649 gnd.n5863 gnd.n1033 240.244
R6650 gnd.n5873 gnd.n1033 240.244
R6651 gnd.n5873 gnd.n1029 240.244
R6652 gnd.n5879 gnd.n1029 240.244
R6653 gnd.n5879 gnd.n1017 240.244
R6654 gnd.n5891 gnd.n1017 240.244
R6655 gnd.n5891 gnd.n1012 240.244
R6656 gnd.n5898 gnd.n1012 240.244
R6657 gnd.n5898 gnd.n989 240.244
R6658 gnd.n989 gnd.n978 240.244
R6659 gnd.n5987 gnd.n978 240.244
R6660 gnd.n5987 gnd.n974 240.244
R6661 gnd.n5993 gnd.n974 240.244
R6662 gnd.n5993 gnd.n962 240.244
R6663 gnd.n6003 gnd.n962 240.244
R6664 gnd.n6003 gnd.n956 240.244
R6665 gnd.n6012 gnd.n956 240.244
R6666 gnd.n6012 gnd.n957 240.244
R6667 gnd.n957 gnd.n947 240.244
R6668 gnd.n947 gnd.n920 240.244
R6669 gnd.n6068 gnd.n920 240.244
R6670 gnd.n6068 gnd.n921 240.244
R6671 gnd.n921 gnd.n910 240.244
R6672 gnd.n926 gnd.n910 240.244
R6673 gnd.n6057 gnd.n926 240.244
R6674 gnd.n6057 gnd.n886 240.244
R6675 gnd.n886 gnd.n875 240.244
R6676 gnd.n6842 gnd.n875 240.244
R6677 gnd.n6842 gnd.n871 240.244
R6678 gnd.n6848 gnd.n871 240.244
R6679 gnd.n6848 gnd.n859 240.244
R6680 gnd.n6858 gnd.n859 240.244
R6681 gnd.n6858 gnd.n855 240.244
R6682 gnd.n6864 gnd.n855 240.244
R6683 gnd.n6864 gnd.n843 240.244
R6684 gnd.n6874 gnd.n843 240.244
R6685 gnd.n6874 gnd.n839 240.244
R6686 gnd.n6880 gnd.n839 240.244
R6687 gnd.n6880 gnd.n827 240.244
R6688 gnd.n6890 gnd.n827 240.244
R6689 gnd.n6890 gnd.n823 240.244
R6690 gnd.n6896 gnd.n823 240.244
R6691 gnd.n6896 gnd.n811 240.244
R6692 gnd.n6906 gnd.n811 240.244
R6693 gnd.n6906 gnd.n807 240.244
R6694 gnd.n6912 gnd.n807 240.244
R6695 gnd.n6912 gnd.n796 240.244
R6696 gnd.n6922 gnd.n796 240.244
R6697 gnd.n6922 gnd.n792 240.244
R6698 gnd.n6928 gnd.n792 240.244
R6699 gnd.n6928 gnd.n780 240.244
R6700 gnd.n6938 gnd.n780 240.244
R6701 gnd.n6938 gnd.n776 240.244
R6702 gnd.n6944 gnd.n776 240.244
R6703 gnd.n6944 gnd.n764 240.244
R6704 gnd.n6954 gnd.n764 240.244
R6705 gnd.n6954 gnd.n760 240.244
R6706 gnd.n6960 gnd.n760 240.244
R6707 gnd.n6960 gnd.n747 240.244
R6708 gnd.n6970 gnd.n747 240.244
R6709 gnd.n6970 gnd.n743 240.244
R6710 gnd.n6976 gnd.n743 240.244
R6711 gnd.n6976 gnd.n733 240.244
R6712 gnd.n6986 gnd.n733 240.244
R6713 gnd.n6986 gnd.n729 240.244
R6714 gnd.n6992 gnd.n729 240.244
R6715 gnd.n6992 gnd.n717 240.244
R6716 gnd.n7002 gnd.n717 240.244
R6717 gnd.n7002 gnd.n713 240.244
R6718 gnd.n7008 gnd.n713 240.244
R6719 gnd.n7008 gnd.n703 240.244
R6720 gnd.n7018 gnd.n703 240.244
R6721 gnd.n7018 gnd.n699 240.244
R6722 gnd.n7024 gnd.n699 240.244
R6723 gnd.n7024 gnd.n690 240.244
R6724 gnd.n7034 gnd.n690 240.244
R6725 gnd.n7034 gnd.n686 240.244
R6726 gnd.n7040 gnd.n686 240.244
R6727 gnd.n7040 gnd.n676 240.244
R6728 gnd.n7050 gnd.n676 240.244
R6729 gnd.n7050 gnd.n672 240.244
R6730 gnd.n7057 gnd.n672 240.244
R6731 gnd.n7057 gnd.n660 240.244
R6732 gnd.n7069 gnd.n660 240.244
R6733 gnd.n7069 gnd.n655 240.244
R6734 gnd.n6605 gnd.n6604 240.244
R6735 gnd.n6607 gnd.n6606 240.244
R6736 gnd.n6615 gnd.n6614 240.244
R6737 gnd.n6625 gnd.n6624 240.244
R6738 gnd.n6627 gnd.n6626 240.244
R6739 gnd.n6635 gnd.n6634 240.244
R6740 gnd.n6645 gnd.n6644 240.244
R6741 gnd.n6647 gnd.n6646 240.244
R6742 gnd.n6652 gnd.n6651 240.244
R6743 gnd.n6654 gnd.n6653 240.244
R6744 gnd.n6658 gnd.n6657 240.244
R6745 gnd.n6660 gnd.n6659 240.244
R6746 gnd.n6667 gnd.n6666 240.244
R6747 gnd.n7075 gnd.n654 240.244
R6748 gnd.n5408 gnd.n5407 240.132
R6749 gnd.n6418 gnd.n6417 240.132
R6750 gnd.n2843 gnd.n1783 225.874
R6751 gnd.n2835 gnd.n1783 225.874
R6752 gnd.n2835 gnd.n2834 225.874
R6753 gnd.n2834 gnd.n2833 225.874
R6754 gnd.n2833 gnd.n1789 225.874
R6755 gnd.n2827 gnd.n1789 225.874
R6756 gnd.n2827 gnd.n2826 225.874
R6757 gnd.n2826 gnd.n2825 225.874
R6758 gnd.n2825 gnd.n1796 225.874
R6759 gnd.n2819 gnd.n1796 225.874
R6760 gnd.n2819 gnd.n2818 225.874
R6761 gnd.n2818 gnd.n2817 225.874
R6762 gnd.n2817 gnd.n1804 225.874
R6763 gnd.n2811 gnd.n1804 225.874
R6764 gnd.n2811 gnd.n2810 225.874
R6765 gnd.n2810 gnd.n2809 225.874
R6766 gnd.n2809 gnd.n1812 225.874
R6767 gnd.n2803 gnd.n1812 225.874
R6768 gnd.n2803 gnd.n2802 225.874
R6769 gnd.n2802 gnd.n2801 225.874
R6770 gnd.n2801 gnd.n1820 225.874
R6771 gnd.n2795 gnd.n1820 225.874
R6772 gnd.n2795 gnd.n2794 225.874
R6773 gnd.n2794 gnd.n2793 225.874
R6774 gnd.n2793 gnd.n1828 225.874
R6775 gnd.n2787 gnd.n1828 225.874
R6776 gnd.n2787 gnd.n2786 225.874
R6777 gnd.n2786 gnd.n2785 225.874
R6778 gnd.n2785 gnd.n1836 225.874
R6779 gnd.n2779 gnd.n1836 225.874
R6780 gnd.n2779 gnd.n2778 225.874
R6781 gnd.n2778 gnd.n2777 225.874
R6782 gnd.n2777 gnd.n1844 225.874
R6783 gnd.n2771 gnd.n1844 225.874
R6784 gnd.n2771 gnd.n2770 225.874
R6785 gnd.n2770 gnd.n2769 225.874
R6786 gnd.n2769 gnd.n1852 225.874
R6787 gnd.n2763 gnd.n1852 225.874
R6788 gnd.n2763 gnd.n2762 225.874
R6789 gnd.n2762 gnd.n2761 225.874
R6790 gnd.n2761 gnd.n1860 225.874
R6791 gnd.n2755 gnd.n1860 225.874
R6792 gnd.n2755 gnd.n2754 225.874
R6793 gnd.n2754 gnd.n2753 225.874
R6794 gnd.n2753 gnd.n1868 225.874
R6795 gnd.n2747 gnd.n1868 225.874
R6796 gnd.n2747 gnd.n2746 225.874
R6797 gnd.n2746 gnd.n2745 225.874
R6798 gnd.n2745 gnd.n1876 225.874
R6799 gnd.n2739 gnd.n1876 225.874
R6800 gnd.n2739 gnd.n2738 225.874
R6801 gnd.n2738 gnd.n2737 225.874
R6802 gnd.n2737 gnd.n1884 225.874
R6803 gnd.n2731 gnd.n1884 225.874
R6804 gnd.n2731 gnd.n2730 225.874
R6805 gnd.n2730 gnd.n2729 225.874
R6806 gnd.n2729 gnd.n1892 225.874
R6807 gnd.n2723 gnd.n1892 225.874
R6808 gnd.n2723 gnd.n2722 225.874
R6809 gnd.n2722 gnd.n2721 225.874
R6810 gnd.n2721 gnd.n1900 225.874
R6811 gnd.n2715 gnd.n1900 225.874
R6812 gnd.n2715 gnd.n2714 225.874
R6813 gnd.n2714 gnd.n2713 225.874
R6814 gnd.n2713 gnd.n1908 225.874
R6815 gnd.n2707 gnd.n1908 225.874
R6816 gnd.n2707 gnd.n2706 225.874
R6817 gnd.n2706 gnd.n2705 225.874
R6818 gnd.n2705 gnd.n1916 225.874
R6819 gnd.n2699 gnd.n1916 225.874
R6820 gnd.n2699 gnd.n2698 225.874
R6821 gnd.n2698 gnd.n2697 225.874
R6822 gnd.n2697 gnd.n1924 225.874
R6823 gnd.n2691 gnd.n1924 225.874
R6824 gnd.n2691 gnd.n2690 225.874
R6825 gnd.n2690 gnd.n2689 225.874
R6826 gnd.n2689 gnd.n1932 225.874
R6827 gnd.n2683 gnd.n1932 225.874
R6828 gnd.n2683 gnd.n2682 225.874
R6829 gnd.n2682 gnd.n2681 225.874
R6830 gnd.n2681 gnd.n1940 225.874
R6831 gnd.n2675 gnd.n1940 225.874
R6832 gnd.n2675 gnd.n2674 225.874
R6833 gnd.n2674 gnd.n2673 225.874
R6834 gnd.n2673 gnd.n1948 225.874
R6835 gnd.n2667 gnd.n1948 225.874
R6836 gnd.n2667 gnd.n2666 225.874
R6837 gnd.n2666 gnd.n2665 225.874
R6838 gnd.n2665 gnd.n1956 225.874
R6839 gnd.n2659 gnd.n1956 225.874
R6840 gnd.n2659 gnd.n2658 225.874
R6841 gnd.n2658 gnd.n2657 225.874
R6842 gnd.n2657 gnd.n1964 225.874
R6843 gnd.n2651 gnd.n1964 225.874
R6844 gnd.n2651 gnd.n2650 225.874
R6845 gnd.n2650 gnd.n2649 225.874
R6846 gnd.n2649 gnd.n1972 225.874
R6847 gnd.n2643 gnd.n1972 225.874
R6848 gnd.n2643 gnd.n2642 225.874
R6849 gnd.n2642 gnd.n2641 225.874
R6850 gnd.n2641 gnd.n1980 225.874
R6851 gnd.n2635 gnd.n1980 225.874
R6852 gnd.n2635 gnd.n2634 225.874
R6853 gnd.n2634 gnd.n2633 225.874
R6854 gnd.n2633 gnd.n1988 225.874
R6855 gnd.n2627 gnd.n1988 225.874
R6856 gnd.n2627 gnd.n2626 225.874
R6857 gnd.n2626 gnd.n2625 225.874
R6858 gnd.n2625 gnd.n1996 225.874
R6859 gnd.n2619 gnd.n1996 225.874
R6860 gnd.n2619 gnd.n2618 225.874
R6861 gnd.n2618 gnd.n2617 225.874
R6862 gnd.n2617 gnd.n2004 225.874
R6863 gnd.n2611 gnd.n2004 225.874
R6864 gnd.n2611 gnd.n2610 225.874
R6865 gnd.n2610 gnd.n2609 225.874
R6866 gnd.n2609 gnd.n2012 225.874
R6867 gnd.n2603 gnd.n2012 225.874
R6868 gnd.n2603 gnd.n2602 225.874
R6869 gnd.n2602 gnd.n2601 225.874
R6870 gnd.n2601 gnd.n2020 225.874
R6871 gnd.n2595 gnd.n2020 225.874
R6872 gnd.n2595 gnd.n2594 225.874
R6873 gnd.n2594 gnd.n2593 225.874
R6874 gnd.n2593 gnd.n2028 225.874
R6875 gnd.n2587 gnd.n2028 225.874
R6876 gnd.n2587 gnd.n2586 225.874
R6877 gnd.n2586 gnd.n2585 225.874
R6878 gnd.n2585 gnd.n2036 225.874
R6879 gnd.n2579 gnd.n2036 225.874
R6880 gnd.n2579 gnd.n2578 225.874
R6881 gnd.n2578 gnd.n2577 225.874
R6882 gnd.n2577 gnd.n2044 225.874
R6883 gnd.n2571 gnd.n2044 225.874
R6884 gnd.n2571 gnd.n2570 225.874
R6885 gnd.n2570 gnd.n2569 225.874
R6886 gnd.n2569 gnd.n2052 225.874
R6887 gnd.n2563 gnd.n2052 225.874
R6888 gnd.n2563 gnd.n2562 225.874
R6889 gnd.n2562 gnd.n2561 225.874
R6890 gnd.n2561 gnd.n2060 225.874
R6891 gnd.n2555 gnd.n2060 225.874
R6892 gnd.n2555 gnd.n2554 225.874
R6893 gnd.n2554 gnd.n2553 225.874
R6894 gnd.n2553 gnd.n2068 225.874
R6895 gnd.n2547 gnd.n2068 225.874
R6896 gnd.n2547 gnd.n2546 225.874
R6897 gnd.n2546 gnd.n2545 225.874
R6898 gnd.n2545 gnd.n2076 225.874
R6899 gnd.n2539 gnd.n2076 225.874
R6900 gnd.n2539 gnd.n2538 225.874
R6901 gnd.n2538 gnd.n2537 225.874
R6902 gnd.n2537 gnd.n2084 225.874
R6903 gnd.n2531 gnd.n2084 225.874
R6904 gnd.n2531 gnd.n2530 225.874
R6905 gnd.n2530 gnd.n2529 225.874
R6906 gnd.n2529 gnd.n2092 225.874
R6907 gnd.n2523 gnd.n2092 225.874
R6908 gnd.n2523 gnd.n2522 225.874
R6909 gnd.n2522 gnd.n2521 225.874
R6910 gnd.n2521 gnd.n2100 225.874
R6911 gnd.n2515 gnd.n2100 225.874
R6912 gnd.n2515 gnd.n2514 225.874
R6913 gnd.n2514 gnd.n2513 225.874
R6914 gnd.n2513 gnd.n2108 225.874
R6915 gnd.n2507 gnd.n2108 225.874
R6916 gnd.n2507 gnd.n2506 225.874
R6917 gnd.n2506 gnd.n2505 225.874
R6918 gnd.n2505 gnd.n2116 225.874
R6919 gnd.n2499 gnd.n2116 225.874
R6920 gnd.n2499 gnd.n2498 225.874
R6921 gnd.n2498 gnd.n2497 225.874
R6922 gnd.n2497 gnd.n2124 225.874
R6923 gnd.n2491 gnd.n2124 225.874
R6924 gnd.n2491 gnd.n2490 225.874
R6925 gnd.n2490 gnd.n2489 225.874
R6926 gnd.n2489 gnd.n2132 225.874
R6927 gnd.n2483 gnd.n2132 225.874
R6928 gnd.n2483 gnd.n2482 225.874
R6929 gnd.n2482 gnd.n2481 225.874
R6930 gnd.n2481 gnd.n2140 225.874
R6931 gnd.n3537 gnd.t253 224.174
R6932 gnd.n1629 gnd.t229 224.174
R6933 gnd.n552 gnd.n511 199.319
R6934 gnd.n552 gnd.n512 199.319
R6935 gnd.n5709 gnd.n5708 199.319
R6936 gnd.n5708 gnd.n5707 199.319
R6937 gnd.n5409 gnd.n5406 186.49
R6938 gnd.n6419 gnd.n6416 186.49
R6939 gnd.n4312 gnd.n4311 185
R6940 gnd.n4310 gnd.n4309 185
R6941 gnd.n4289 gnd.n4288 185
R6942 gnd.n4304 gnd.n4303 185
R6943 gnd.n4302 gnd.n4301 185
R6944 gnd.n4293 gnd.n4292 185
R6945 gnd.n4296 gnd.n4295 185
R6946 gnd.n4280 gnd.n4279 185
R6947 gnd.n4278 gnd.n4277 185
R6948 gnd.n4257 gnd.n4256 185
R6949 gnd.n4272 gnd.n4271 185
R6950 gnd.n4270 gnd.n4269 185
R6951 gnd.n4261 gnd.n4260 185
R6952 gnd.n4264 gnd.n4263 185
R6953 gnd.n4248 gnd.n4247 185
R6954 gnd.n4246 gnd.n4245 185
R6955 gnd.n4225 gnd.n4224 185
R6956 gnd.n4240 gnd.n4239 185
R6957 gnd.n4238 gnd.n4237 185
R6958 gnd.n4229 gnd.n4228 185
R6959 gnd.n4232 gnd.n4231 185
R6960 gnd.n4217 gnd.n4216 185
R6961 gnd.n4215 gnd.n4214 185
R6962 gnd.n4194 gnd.n4193 185
R6963 gnd.n4209 gnd.n4208 185
R6964 gnd.n4207 gnd.n4206 185
R6965 gnd.n4198 gnd.n4197 185
R6966 gnd.n4201 gnd.n4200 185
R6967 gnd.n4185 gnd.n4184 185
R6968 gnd.n4183 gnd.n4182 185
R6969 gnd.n4162 gnd.n4161 185
R6970 gnd.n4177 gnd.n4176 185
R6971 gnd.n4175 gnd.n4174 185
R6972 gnd.n4166 gnd.n4165 185
R6973 gnd.n4169 gnd.n4168 185
R6974 gnd.n4153 gnd.n4152 185
R6975 gnd.n4151 gnd.n4150 185
R6976 gnd.n4130 gnd.n4129 185
R6977 gnd.n4145 gnd.n4144 185
R6978 gnd.n4143 gnd.n4142 185
R6979 gnd.n4134 gnd.n4133 185
R6980 gnd.n4137 gnd.n4136 185
R6981 gnd.n4121 gnd.n4120 185
R6982 gnd.n4119 gnd.n4118 185
R6983 gnd.n4098 gnd.n4097 185
R6984 gnd.n4113 gnd.n4112 185
R6985 gnd.n4111 gnd.n4110 185
R6986 gnd.n4102 gnd.n4101 185
R6987 gnd.n4105 gnd.n4104 185
R6988 gnd.n4090 gnd.n4089 185
R6989 gnd.n4088 gnd.n4087 185
R6990 gnd.n4067 gnd.n4066 185
R6991 gnd.n4082 gnd.n4081 185
R6992 gnd.n4080 gnd.n4079 185
R6993 gnd.n4071 gnd.n4070 185
R6994 gnd.n4074 gnd.n4073 185
R6995 gnd.n3538 gnd.t252 178.987
R6996 gnd.n1630 gnd.t230 178.987
R6997 gnd.n1 gnd.t154 170.774
R6998 gnd.n9 gnd.t363 170.103
R6999 gnd.n8 gnd.t296 170.103
R7000 gnd.n7 gnd.t116 170.103
R7001 gnd.n6 gnd.t2 170.103
R7002 gnd.n5 gnd.t160 170.103
R7003 gnd.n4 gnd.t360 170.103
R7004 gnd.n3 gnd.t4 170.103
R7005 gnd.n2 gnd.t6 170.103
R7006 gnd.n1 gnd.t317 170.103
R7007 gnd.n6432 gnd.n6430 163.367
R7008 gnd.n6436 gnd.n6406 163.367
R7009 gnd.n6440 gnd.n6438 163.367
R7010 gnd.n6444 gnd.n6404 163.367
R7011 gnd.n6448 gnd.n6446 163.367
R7012 gnd.n6452 gnd.n6402 163.367
R7013 gnd.n6456 gnd.n6454 163.367
R7014 gnd.n6460 gnd.n6400 163.367
R7015 gnd.n6464 gnd.n6462 163.367
R7016 gnd.n6468 gnd.n6398 163.367
R7017 gnd.n6472 gnd.n6470 163.367
R7018 gnd.n6476 gnd.n6396 163.367
R7019 gnd.n6480 gnd.n6478 163.367
R7020 gnd.n6487 gnd.n6394 163.367
R7021 gnd.n6490 gnd.n6489 163.367
R7022 gnd.n6494 gnd.n6493 163.367
R7023 gnd.n6499 gnd.n6497 163.367
R7024 gnd.n6503 gnd.n6501 163.367
R7025 gnd.n6508 gnd.n6388 163.367
R7026 gnd.n6512 gnd.n6510 163.367
R7027 gnd.n6516 gnd.n6386 163.367
R7028 gnd.n6520 gnd.n6518 163.367
R7029 gnd.n6524 gnd.n6384 163.367
R7030 gnd.n6528 gnd.n6526 163.367
R7031 gnd.n6532 gnd.n6382 163.367
R7032 gnd.n6536 gnd.n6534 163.367
R7033 gnd.n6540 gnd.n6380 163.367
R7034 gnd.n6544 gnd.n6542 163.367
R7035 gnd.n6548 gnd.n6378 163.367
R7036 gnd.n6552 gnd.n6550 163.367
R7037 gnd.n6556 gnd.n6376 163.367
R7038 gnd.n6560 gnd.n6558 163.367
R7039 gnd.n5464 gnd.n5397 163.367
R7040 gnd.n5602 gnd.n5397 163.367
R7041 gnd.n5603 gnd.n5602 163.367
R7042 gnd.n5603 gnd.n5378 163.367
R7043 gnd.n5606 gnd.n5378 163.367
R7044 gnd.n5606 gnd.n5394 163.367
R7045 gnd.n5611 gnd.n5394 163.367
R7046 gnd.n5611 gnd.n5395 163.367
R7047 gnd.n5395 gnd.n990 163.367
R7048 gnd.n5977 gnd.n990 163.367
R7049 gnd.n5977 gnd.n991 163.367
R7050 gnd.n5973 gnd.n991 163.367
R7051 gnd.n5973 gnd.n5972 163.367
R7052 gnd.n5972 gnd.n5971 163.367
R7053 gnd.n5971 gnd.n994 163.367
R7054 gnd.n5918 gnd.n994 163.367
R7055 gnd.n5918 gnd.n1001 163.367
R7056 gnd.n5916 gnd.n1001 163.367
R7057 gnd.n5923 gnd.n5916 163.367
R7058 gnd.n5935 gnd.n5923 163.367
R7059 gnd.n5936 gnd.n5935 163.367
R7060 gnd.n5936 gnd.n5914 163.367
R7061 gnd.n5942 gnd.n5914 163.367
R7062 gnd.n5942 gnd.n945 163.367
R7063 gnd.n945 gnd.n937 163.367
R7064 gnd.n6033 gnd.n937 163.367
R7065 gnd.n6034 gnd.n6033 163.367
R7066 gnd.n6035 gnd.n6034 163.367
R7067 gnd.n6035 gnd.n934 163.367
R7068 gnd.n6045 gnd.n934 163.367
R7069 gnd.n6045 gnd.n935 163.367
R7070 gnd.n6041 gnd.n935 163.367
R7071 gnd.n6041 gnd.n927 163.367
R7072 gnd.n927 gnd.n887 163.367
R7073 gnd.n6832 gnd.n887 163.367
R7074 gnd.n6832 gnd.n888 163.367
R7075 gnd.n6828 gnd.n888 163.367
R7076 gnd.n6828 gnd.n891 163.367
R7077 gnd.n899 gnd.n891 163.367
R7078 gnd.n6210 gnd.n899 163.367
R7079 gnd.n6214 gnd.n6210 163.367
R7080 gnd.n6224 gnd.n6214 163.367
R7081 gnd.n6225 gnd.n6224 163.367
R7082 gnd.n6225 gnd.n6207 163.367
R7083 gnd.n6231 gnd.n6207 163.367
R7084 gnd.n6231 gnd.n6208 163.367
R7085 gnd.n6208 gnd.n6201 163.367
R7086 gnd.n6243 gnd.n6201 163.367
R7087 gnd.n6244 gnd.n6243 163.367
R7088 gnd.n6244 gnd.n6198 163.367
R7089 gnd.n6250 gnd.n6198 163.367
R7090 gnd.n6250 gnd.n6199 163.367
R7091 gnd.n6199 gnd.n6192 163.367
R7092 gnd.n6262 gnd.n6192 163.367
R7093 gnd.n6263 gnd.n6262 163.367
R7094 gnd.n6263 gnd.n6189 163.367
R7095 gnd.n6269 gnd.n6189 163.367
R7096 gnd.n6269 gnd.n6190 163.367
R7097 gnd.n6190 gnd.n6184 163.367
R7098 gnd.n6281 gnd.n6184 163.367
R7099 gnd.n6282 gnd.n6281 163.367
R7100 gnd.n6282 gnd.n6181 163.367
R7101 gnd.n6288 gnd.n6181 163.367
R7102 gnd.n6288 gnd.n6182 163.367
R7103 gnd.n6182 gnd.n6173 163.367
R7104 gnd.n6299 gnd.n6173 163.367
R7105 gnd.n6300 gnd.n6299 163.367
R7106 gnd.n6300 gnd.n6170 163.367
R7107 gnd.n6306 gnd.n6170 163.367
R7108 gnd.n6306 gnd.n6171 163.367
R7109 gnd.n6171 gnd.n6163 163.367
R7110 gnd.n6317 gnd.n6163 163.367
R7111 gnd.n6318 gnd.n6317 163.367
R7112 gnd.n6318 gnd.n6160 163.367
R7113 gnd.n6324 gnd.n6160 163.367
R7114 gnd.n6324 gnd.n6161 163.367
R7115 gnd.n6161 gnd.n6153 163.367
R7116 gnd.n6335 gnd.n6153 163.367
R7117 gnd.n6336 gnd.n6335 163.367
R7118 gnd.n6336 gnd.n6150 163.367
R7119 gnd.n6341 gnd.n6150 163.367
R7120 gnd.n6341 gnd.n6151 163.367
R7121 gnd.n6151 gnd.n6144 163.367
R7122 gnd.n6352 gnd.n6144 163.367
R7123 gnd.n6352 gnd.n751 163.367
R7124 gnd.n6141 gnd.n751 163.367
R7125 gnd.n6359 gnd.n6141 163.367
R7126 gnd.n6359 gnd.n6142 163.367
R7127 gnd.n6142 gnd.n6134 163.367
R7128 gnd.n6368 gnd.n6134 163.367
R7129 gnd.n6369 gnd.n6368 163.367
R7130 gnd.n6369 gnd.n6125 163.367
R7131 gnd.n6372 gnd.n6125 163.367
R7132 gnd.n6372 gnd.n6131 163.367
R7133 gnd.n6564 gnd.n6131 163.367
R7134 gnd.n5592 gnd.n5591 163.367
R7135 gnd.n5591 gnd.n5590 163.367
R7136 gnd.n5587 gnd.n5586 163.367
R7137 gnd.n5584 gnd.n5427 163.367
R7138 gnd.n5580 gnd.n5578 163.367
R7139 gnd.n5576 gnd.n5429 163.367
R7140 gnd.n5572 gnd.n5570 163.367
R7141 gnd.n5568 gnd.n5431 163.367
R7142 gnd.n5564 gnd.n5562 163.367
R7143 gnd.n5560 gnd.n5433 163.367
R7144 gnd.n5556 gnd.n5554 163.367
R7145 gnd.n5552 gnd.n5435 163.367
R7146 gnd.n5548 gnd.n5546 163.367
R7147 gnd.n5544 gnd.n5437 163.367
R7148 gnd.n5540 gnd.n5538 163.367
R7149 gnd.n5535 gnd.n5534 163.367
R7150 gnd.n5530 gnd.n5529 163.367
R7151 gnd.n5527 gnd.n5445 163.367
R7152 gnd.n5522 gnd.n5520 163.367
R7153 gnd.n5518 gnd.n5449 163.367
R7154 gnd.n5514 gnd.n5512 163.367
R7155 gnd.n5510 gnd.n5451 163.367
R7156 gnd.n5506 gnd.n5504 163.367
R7157 gnd.n5502 gnd.n5453 163.367
R7158 gnd.n5498 gnd.n5496 163.367
R7159 gnd.n5494 gnd.n5455 163.367
R7160 gnd.n5490 gnd.n5488 163.367
R7161 gnd.n5486 gnd.n5457 163.367
R7162 gnd.n5482 gnd.n5480 163.367
R7163 gnd.n5478 gnd.n5459 163.367
R7164 gnd.n5474 gnd.n5472 163.367
R7165 gnd.n5470 gnd.n5461 163.367
R7166 gnd.n5596 gnd.n5401 163.367
R7167 gnd.n5600 gnd.n5401 163.367
R7168 gnd.n5600 gnd.n5379 163.367
R7169 gnd.n5619 gnd.n5379 163.367
R7170 gnd.n5619 gnd.n5380 163.367
R7171 gnd.n5615 gnd.n5380 163.367
R7172 gnd.n5615 gnd.n5614 163.367
R7173 gnd.n5614 gnd.n5393 163.367
R7174 gnd.n5393 gnd.n5383 163.367
R7175 gnd.n5383 gnd.n987 163.367
R7176 gnd.n5388 gnd.n987 163.367
R7177 gnd.n5388 gnd.n5385 163.367
R7178 gnd.n5385 gnd.n996 163.367
R7179 gnd.n5969 gnd.n996 163.367
R7180 gnd.n5969 gnd.n997 163.367
R7181 gnd.n5965 gnd.n997 163.367
R7182 gnd.n5965 gnd.n5964 163.367
R7183 gnd.n5964 gnd.n1000 163.367
R7184 gnd.n5925 gnd.n1000 163.367
R7185 gnd.n5933 gnd.n5925 163.367
R7186 gnd.n5933 gnd.n5926 163.367
R7187 gnd.n5929 gnd.n5926 163.367
R7188 gnd.n5929 gnd.n944 163.367
R7189 gnd.n6023 gnd.n944 163.367
R7190 gnd.n6023 gnd.n941 163.367
R7191 gnd.n6031 gnd.n941 163.367
R7192 gnd.n6031 gnd.n942 163.367
R7193 gnd.n6027 gnd.n942 163.367
R7194 gnd.n6027 gnd.n931 163.367
R7195 gnd.n6047 gnd.n931 163.367
R7196 gnd.n6048 gnd.n6047 163.367
R7197 gnd.n6048 gnd.n928 163.367
R7198 gnd.n6054 gnd.n928 163.367
R7199 gnd.n6054 gnd.n929 163.367
R7200 gnd.n929 gnd.n884 163.367
R7201 gnd.n894 gnd.n884 163.367
R7202 gnd.n6826 gnd.n894 163.367
R7203 gnd.n6826 gnd.n895 163.367
R7204 gnd.n6822 gnd.n895 163.367
R7205 gnd.n6822 gnd.n898 163.367
R7206 gnd.n6216 gnd.n898 163.367
R7207 gnd.n6222 gnd.n6216 163.367
R7208 gnd.n6222 gnd.n6217 163.367
R7209 gnd.n6217 gnd.n6206 163.367
R7210 gnd.n6234 gnd.n6206 163.367
R7211 gnd.n6235 gnd.n6234 163.367
R7212 gnd.n6235 gnd.n6203 163.367
R7213 gnd.n6241 gnd.n6203 163.367
R7214 gnd.n6241 gnd.n6204 163.367
R7215 gnd.n6204 gnd.n6197 163.367
R7216 gnd.n6253 gnd.n6197 163.367
R7217 gnd.n6254 gnd.n6253 163.367
R7218 gnd.n6254 gnd.n6194 163.367
R7219 gnd.n6260 gnd.n6194 163.367
R7220 gnd.n6260 gnd.n6195 163.367
R7221 gnd.n6195 gnd.n6188 163.367
R7222 gnd.n6272 gnd.n6188 163.367
R7223 gnd.n6273 gnd.n6272 163.367
R7224 gnd.n6273 gnd.n6185 163.367
R7225 gnd.n6279 gnd.n6185 163.367
R7226 gnd.n6279 gnd.n6186 163.367
R7227 gnd.n6186 gnd.n6179 163.367
R7228 gnd.n6290 gnd.n6179 163.367
R7229 gnd.n6291 gnd.n6290 163.367
R7230 gnd.n6291 gnd.n6176 163.367
R7231 gnd.n6297 gnd.n6176 163.367
R7232 gnd.n6297 gnd.n6177 163.367
R7233 gnd.n6177 gnd.n6168 163.367
R7234 gnd.n6308 gnd.n6168 163.367
R7235 gnd.n6309 gnd.n6308 163.367
R7236 gnd.n6309 gnd.n6165 163.367
R7237 gnd.n6315 gnd.n6165 163.367
R7238 gnd.n6315 gnd.n6166 163.367
R7239 gnd.n6166 gnd.n6158 163.367
R7240 gnd.n6326 gnd.n6158 163.367
R7241 gnd.n6327 gnd.n6326 163.367
R7242 gnd.n6327 gnd.n6155 163.367
R7243 gnd.n6333 gnd.n6155 163.367
R7244 gnd.n6333 gnd.n6156 163.367
R7245 gnd.n6156 gnd.n6148 163.367
R7246 gnd.n6343 gnd.n6148 163.367
R7247 gnd.n6344 gnd.n6343 163.367
R7248 gnd.n6344 gnd.n6146 163.367
R7249 gnd.n6350 gnd.n6146 163.367
R7250 gnd.n6350 gnd.n748 163.367
R7251 gnd.n6139 gnd.n748 163.367
R7252 gnd.n6361 gnd.n6139 163.367
R7253 gnd.n6362 gnd.n6361 163.367
R7254 gnd.n6362 gnd.n6137 163.367
R7255 gnd.n6366 gnd.n6137 163.367
R7256 gnd.n6366 gnd.n6126 163.367
R7257 gnd.n6571 gnd.n6126 163.367
R7258 gnd.n6571 gnd.n6127 163.367
R7259 gnd.n6567 gnd.n6127 163.367
R7260 gnd.n6567 gnd.n6566 163.367
R7261 gnd.n6425 gnd.n6424 156.462
R7262 gnd.n4252 gnd.n4220 153.042
R7263 gnd.n4316 gnd.n4315 152.079
R7264 gnd.n4284 gnd.n4283 152.079
R7265 gnd.n4252 gnd.n4251 152.079
R7266 gnd.n5414 gnd.n5413 152
R7267 gnd.n5415 gnd.n5404 152
R7268 gnd.n5417 gnd.n5416 152
R7269 gnd.n5419 gnd.n5402 152
R7270 gnd.n5421 gnd.n5420 152
R7271 gnd.n6423 gnd.n6407 152
R7272 gnd.n6415 gnd.n6408 152
R7273 gnd.n6414 gnd.n6413 152
R7274 gnd.n6412 gnd.n6409 152
R7275 gnd.n6410 gnd.t199 150.546
R7276 gnd.t22 gnd.n4294 147.661
R7277 gnd.t293 gnd.n4262 147.661
R7278 gnd.t175 gnd.n4230 147.661
R7279 gnd.t24 gnd.n4199 147.661
R7280 gnd.t353 gnd.n4167 147.661
R7281 gnd.t109 gnd.n4135 147.661
R7282 gnd.t149 gnd.n4103 147.661
R7283 gnd.t151 gnd.n4072 147.661
R7284 gnd.n6496 gnd.n6495 143.351
R7285 gnd.n5533 gnd.n5532 143.351
R7286 gnd.n5532 gnd.n5443 143.351
R7287 gnd.n7220 gnd.n551 138.177
R7288 gnd.n5531 gnd.n1222 138.177
R7289 gnd.n5411 gnd.t244 130.484
R7290 gnd.n5420 gnd.t264 126.766
R7291 gnd.n5418 gnd.t210 126.766
R7292 gnd.n5404 gnd.t254 126.766
R7293 gnd.n5412 gnd.t231 126.766
R7294 gnd.n6411 gnd.t184 126.766
R7295 gnd.n6413 gnd.t286 126.766
R7296 gnd.n6422 gnd.t237 126.766
R7297 gnd.n6424 gnd.t220 126.766
R7298 gnd.n4311 gnd.n4310 104.615
R7299 gnd.n4310 gnd.n4288 104.615
R7300 gnd.n4303 gnd.n4288 104.615
R7301 gnd.n4303 gnd.n4302 104.615
R7302 gnd.n4302 gnd.n4292 104.615
R7303 gnd.n4295 gnd.n4292 104.615
R7304 gnd.n4279 gnd.n4278 104.615
R7305 gnd.n4278 gnd.n4256 104.615
R7306 gnd.n4271 gnd.n4256 104.615
R7307 gnd.n4271 gnd.n4270 104.615
R7308 gnd.n4270 gnd.n4260 104.615
R7309 gnd.n4263 gnd.n4260 104.615
R7310 gnd.n4247 gnd.n4246 104.615
R7311 gnd.n4246 gnd.n4224 104.615
R7312 gnd.n4239 gnd.n4224 104.615
R7313 gnd.n4239 gnd.n4238 104.615
R7314 gnd.n4238 gnd.n4228 104.615
R7315 gnd.n4231 gnd.n4228 104.615
R7316 gnd.n4216 gnd.n4215 104.615
R7317 gnd.n4215 gnd.n4193 104.615
R7318 gnd.n4208 gnd.n4193 104.615
R7319 gnd.n4208 gnd.n4207 104.615
R7320 gnd.n4207 gnd.n4197 104.615
R7321 gnd.n4200 gnd.n4197 104.615
R7322 gnd.n4184 gnd.n4183 104.615
R7323 gnd.n4183 gnd.n4161 104.615
R7324 gnd.n4176 gnd.n4161 104.615
R7325 gnd.n4176 gnd.n4175 104.615
R7326 gnd.n4175 gnd.n4165 104.615
R7327 gnd.n4168 gnd.n4165 104.615
R7328 gnd.n4152 gnd.n4151 104.615
R7329 gnd.n4151 gnd.n4129 104.615
R7330 gnd.n4144 gnd.n4129 104.615
R7331 gnd.n4144 gnd.n4143 104.615
R7332 gnd.n4143 gnd.n4133 104.615
R7333 gnd.n4136 gnd.n4133 104.615
R7334 gnd.n4120 gnd.n4119 104.615
R7335 gnd.n4119 gnd.n4097 104.615
R7336 gnd.n4112 gnd.n4097 104.615
R7337 gnd.n4112 gnd.n4111 104.615
R7338 gnd.n4111 gnd.n4101 104.615
R7339 gnd.n4104 gnd.n4101 104.615
R7340 gnd.n4089 gnd.n4088 104.615
R7341 gnd.n4088 gnd.n4066 104.615
R7342 gnd.n4081 gnd.n4066 104.615
R7343 gnd.n4081 gnd.n4080 104.615
R7344 gnd.n4080 gnd.n4070 104.615
R7345 gnd.n4073 gnd.n4070 104.615
R7346 gnd.n3463 gnd.t273 100.632
R7347 gnd.n1603 gnd.t215 100.632
R7348 gnd.n7829 gnd.n138 99.6594
R7349 gnd.n7827 gnd.n7826 99.6594
R7350 gnd.n7822 gnd.n145 99.6594
R7351 gnd.n7820 gnd.n7819 99.6594
R7352 gnd.n7815 gnd.n152 99.6594
R7353 gnd.n7813 gnd.n7812 99.6594
R7354 gnd.n7808 gnd.n159 99.6594
R7355 gnd.n7806 gnd.n7805 99.6594
R7356 gnd.n7798 gnd.n166 99.6594
R7357 gnd.n7796 gnd.n7795 99.6594
R7358 gnd.n7791 gnd.n173 99.6594
R7359 gnd.n7789 gnd.n7788 99.6594
R7360 gnd.n7784 gnd.n180 99.6594
R7361 gnd.n7782 gnd.n7781 99.6594
R7362 gnd.n7777 gnd.n187 99.6594
R7363 gnd.n7775 gnd.n7774 99.6594
R7364 gnd.n7770 gnd.n194 99.6594
R7365 gnd.n7768 gnd.n7767 99.6594
R7366 gnd.n199 gnd.n198 99.6594
R7367 gnd.n7251 gnd.n7250 99.6594
R7368 gnd.n7245 gnd.n505 99.6594
R7369 gnd.n7242 gnd.n506 99.6594
R7370 gnd.n7238 gnd.n507 99.6594
R7371 gnd.n7234 gnd.n508 99.6594
R7372 gnd.n7230 gnd.n509 99.6594
R7373 gnd.n7226 gnd.n510 99.6594
R7374 gnd.n7222 gnd.n511 99.6594
R7375 gnd.n7217 gnd.n513 99.6594
R7376 gnd.n7213 gnd.n514 99.6594
R7377 gnd.n7209 gnd.n515 99.6594
R7378 gnd.n7205 gnd.n516 99.6594
R7379 gnd.n7201 gnd.n517 99.6594
R7380 gnd.n7197 gnd.n518 99.6594
R7381 gnd.n7193 gnd.n519 99.6594
R7382 gnd.n7189 gnd.n520 99.6594
R7383 gnd.n7185 gnd.n521 99.6594
R7384 gnd.n575 gnd.n522 99.6594
R7385 gnd.n5733 gnd.n5732 99.6594
R7386 gnd.n5730 gnd.n5729 99.6594
R7387 gnd.n5725 gnd.n1205 99.6594
R7388 gnd.n5723 gnd.n5722 99.6594
R7389 gnd.n5718 gnd.n1212 99.6594
R7390 gnd.n5716 gnd.n5715 99.6594
R7391 gnd.n5711 gnd.n1219 99.6594
R7392 gnd.n5707 gnd.n5706 99.6594
R7393 gnd.n5702 gnd.n1230 99.6594
R7394 gnd.n5700 gnd.n5699 99.6594
R7395 gnd.n5695 gnd.n1237 99.6594
R7396 gnd.n5693 gnd.n5692 99.6594
R7397 gnd.n5688 gnd.n1244 99.6594
R7398 gnd.n5686 gnd.n5685 99.6594
R7399 gnd.n5681 gnd.n1251 99.6594
R7400 gnd.n5679 gnd.n5678 99.6594
R7401 gnd.n5674 gnd.n1260 99.6594
R7402 gnd.n5672 gnd.n5671 99.6594
R7403 gnd.n4750 gnd.n4567 99.6594
R7404 gnd.n4748 gnd.n4570 99.6594
R7405 gnd.n4744 gnd.n4743 99.6594
R7406 gnd.n4737 gnd.n4575 99.6594
R7407 gnd.n4736 gnd.n4735 99.6594
R7408 gnd.n4729 gnd.n4581 99.6594
R7409 gnd.n4728 gnd.n4727 99.6594
R7410 gnd.n4721 gnd.n4587 99.6594
R7411 gnd.n4720 gnd.n4719 99.6594
R7412 gnd.n4713 gnd.n4593 99.6594
R7413 gnd.n4712 gnd.n4711 99.6594
R7414 gnd.n4705 gnd.n4602 99.6594
R7415 gnd.n4704 gnd.n4703 99.6594
R7416 gnd.n4697 gnd.n4608 99.6594
R7417 gnd.n4696 gnd.n4695 99.6594
R7418 gnd.n4689 gnd.n4614 99.6594
R7419 gnd.n4688 gnd.n4687 99.6594
R7420 gnd.n4624 gnd.n4620 99.6594
R7421 gnd.n4677 gnd.n4676 99.6594
R7422 gnd.n4434 gnd.n1586 99.6594
R7423 gnd.n4432 gnd.n1585 99.6594
R7424 gnd.n4428 gnd.n1584 99.6594
R7425 gnd.n4424 gnd.n1583 99.6594
R7426 gnd.n4420 gnd.n1582 99.6594
R7427 gnd.n4416 gnd.n1581 99.6594
R7428 gnd.n4412 gnd.n1580 99.6594
R7429 gnd.n4344 gnd.n1579 99.6594
R7430 gnd.n3675 gnd.n3406 99.6594
R7431 gnd.n3432 gnd.n3413 99.6594
R7432 gnd.n3434 gnd.n3414 99.6594
R7433 gnd.n3442 gnd.n3415 99.6594
R7434 gnd.n3444 gnd.n3416 99.6594
R7435 gnd.n3452 gnd.n3417 99.6594
R7436 gnd.n3454 gnd.n3418 99.6594
R7437 gnd.n3462 gnd.n3419 99.6594
R7438 gnd.n4402 gnd.n1566 99.6594
R7439 gnd.n4398 gnd.n1567 99.6594
R7440 gnd.n4394 gnd.n1568 99.6594
R7441 gnd.n4390 gnd.n1569 99.6594
R7442 gnd.n4386 gnd.n1570 99.6594
R7443 gnd.n4382 gnd.n1571 99.6594
R7444 gnd.n4378 gnd.n1572 99.6594
R7445 gnd.n4374 gnd.n1573 99.6594
R7446 gnd.n4370 gnd.n1574 99.6594
R7447 gnd.n4366 gnd.n1575 99.6594
R7448 gnd.n4362 gnd.n1576 99.6594
R7449 gnd.n4358 gnd.n1577 99.6594
R7450 gnd.n4354 gnd.n1578 99.6594
R7451 gnd.n3590 gnd.n3589 99.6594
R7452 gnd.n3584 gnd.n3501 99.6594
R7453 gnd.n3581 gnd.n3502 99.6594
R7454 gnd.n3577 gnd.n3503 99.6594
R7455 gnd.n3573 gnd.n3504 99.6594
R7456 gnd.n3569 gnd.n3505 99.6594
R7457 gnd.n3565 gnd.n3506 99.6594
R7458 gnd.n3561 gnd.n3507 99.6594
R7459 gnd.n3557 gnd.n3508 99.6594
R7460 gnd.n3553 gnd.n3509 99.6594
R7461 gnd.n3549 gnd.n3510 99.6594
R7462 gnd.n3545 gnd.n3511 99.6594
R7463 gnd.n3592 gnd.n3500 99.6594
R7464 gnd.n7684 gnd.n7683 99.6594
R7465 gnd.n7689 gnd.n7688 99.6594
R7466 gnd.n7692 gnd.n7691 99.6594
R7467 gnd.n7697 gnd.n7696 99.6594
R7468 gnd.n7700 gnd.n7699 99.6594
R7469 gnd.n7705 gnd.n7704 99.6594
R7470 gnd.n7708 gnd.n7707 99.6594
R7471 gnd.n7713 gnd.n7711 99.6594
R7472 gnd.n7839 gnd.n125 99.6594
R7473 gnd.n7254 gnd.n7253 99.6594
R7474 gnd.n6599 gnd.n523 99.6594
R7475 gnd.n6601 gnd.n524 99.6594
R7476 gnd.n6611 gnd.n525 99.6594
R7477 gnd.n6619 gnd.n526 99.6594
R7478 gnd.n6621 gnd.n527 99.6594
R7479 gnd.n6631 gnd.n528 99.6594
R7480 gnd.n6639 gnd.n529 99.6594
R7481 gnd.n6641 gnd.n530 99.6594
R7482 gnd.n5353 gnd.n5352 99.6594
R7483 gnd.n1185 gnd.n1125 99.6594
R7484 gnd.n1187 gnd.n1133 99.6594
R7485 gnd.n1189 gnd.n1188 99.6594
R7486 gnd.n1190 gnd.n1142 99.6594
R7487 gnd.n1192 gnd.n1151 99.6594
R7488 gnd.n1194 gnd.n1193 99.6594
R7489 gnd.n1195 gnd.n1160 99.6594
R7490 gnd.n5743 gnd.n1172 99.6594
R7491 gnd.n4469 gnd.n1563 99.6594
R7492 gnd.n4472 gnd.n4471 99.6594
R7493 gnd.n4479 gnd.n4478 99.6594
R7494 gnd.n4482 gnd.n4481 99.6594
R7495 gnd.n4489 gnd.n4488 99.6594
R7496 gnd.n4492 gnd.n4491 99.6594
R7497 gnd.n4499 gnd.n4498 99.6594
R7498 gnd.n4502 gnd.n4501 99.6594
R7499 gnd.n4509 gnd.n4508 99.6594
R7500 gnd.n4470 gnd.n4469 99.6594
R7501 gnd.n4471 gnd.n4464 99.6594
R7502 gnd.n4480 gnd.n4479 99.6594
R7503 gnd.n4481 gnd.n4460 99.6594
R7504 gnd.n4490 gnd.n4489 99.6594
R7505 gnd.n4491 gnd.n4456 99.6594
R7506 gnd.n4500 gnd.n4499 99.6594
R7507 gnd.n4501 gnd.n4452 99.6594
R7508 gnd.n4510 gnd.n4509 99.6594
R7509 gnd.n1172 gnd.n1171 99.6594
R7510 gnd.n1195 gnd.n1159 99.6594
R7511 gnd.n1194 gnd.n1152 99.6594
R7512 gnd.n1192 gnd.n1191 99.6594
R7513 gnd.n1190 gnd.n1141 99.6594
R7514 gnd.n1189 gnd.n1134 99.6594
R7515 gnd.n1187 gnd.n1186 99.6594
R7516 gnd.n1185 gnd.n1124 99.6594
R7517 gnd.n5354 gnd.n5353 99.6594
R7518 gnd.n7253 gnd.n503 99.6594
R7519 gnd.n6600 gnd.n523 99.6594
R7520 gnd.n6610 gnd.n524 99.6594
R7521 gnd.n6618 gnd.n525 99.6594
R7522 gnd.n6620 gnd.n526 99.6594
R7523 gnd.n6630 gnd.n527 99.6594
R7524 gnd.n6638 gnd.n528 99.6594
R7525 gnd.n6640 gnd.n529 99.6594
R7526 gnd.n6685 gnd.n530 99.6594
R7527 gnd.n7712 gnd.n125 99.6594
R7528 gnd.n7711 gnd.n7710 99.6594
R7529 gnd.n7707 gnd.n7706 99.6594
R7530 gnd.n7704 gnd.n7703 99.6594
R7531 gnd.n7699 gnd.n7698 99.6594
R7532 gnd.n7696 gnd.n7695 99.6594
R7533 gnd.n7691 gnd.n7690 99.6594
R7534 gnd.n7688 gnd.n7687 99.6594
R7535 gnd.n7683 gnd.n7682 99.6594
R7536 gnd.n3590 gnd.n3513 99.6594
R7537 gnd.n3582 gnd.n3501 99.6594
R7538 gnd.n3578 gnd.n3502 99.6594
R7539 gnd.n3574 gnd.n3503 99.6594
R7540 gnd.n3570 gnd.n3504 99.6594
R7541 gnd.n3566 gnd.n3505 99.6594
R7542 gnd.n3562 gnd.n3506 99.6594
R7543 gnd.n3558 gnd.n3507 99.6594
R7544 gnd.n3554 gnd.n3508 99.6594
R7545 gnd.n3550 gnd.n3509 99.6594
R7546 gnd.n3546 gnd.n3510 99.6594
R7547 gnd.n3542 gnd.n3511 99.6594
R7548 gnd.n3593 gnd.n3592 99.6594
R7549 gnd.n4357 gnd.n1578 99.6594
R7550 gnd.n4361 gnd.n1577 99.6594
R7551 gnd.n4365 gnd.n1576 99.6594
R7552 gnd.n4369 gnd.n1575 99.6594
R7553 gnd.n4373 gnd.n1574 99.6594
R7554 gnd.n4377 gnd.n1573 99.6594
R7555 gnd.n4381 gnd.n1572 99.6594
R7556 gnd.n4385 gnd.n1571 99.6594
R7557 gnd.n4389 gnd.n1570 99.6594
R7558 gnd.n4393 gnd.n1569 99.6594
R7559 gnd.n4397 gnd.n1568 99.6594
R7560 gnd.n4401 gnd.n1567 99.6594
R7561 gnd.n1607 gnd.n1566 99.6594
R7562 gnd.n3676 gnd.n3675 99.6594
R7563 gnd.n3435 gnd.n3413 99.6594
R7564 gnd.n3441 gnd.n3414 99.6594
R7565 gnd.n3445 gnd.n3415 99.6594
R7566 gnd.n3451 gnd.n3416 99.6594
R7567 gnd.n3455 gnd.n3417 99.6594
R7568 gnd.n3461 gnd.n3418 99.6594
R7569 gnd.n3419 gnd.n3403 99.6594
R7570 gnd.n4411 gnd.n1579 99.6594
R7571 gnd.n4415 gnd.n1580 99.6594
R7572 gnd.n4419 gnd.n1581 99.6594
R7573 gnd.n4423 gnd.n1582 99.6594
R7574 gnd.n4427 gnd.n1583 99.6594
R7575 gnd.n4431 gnd.n1584 99.6594
R7576 gnd.n4435 gnd.n1585 99.6594
R7577 gnd.n1588 gnd.n1586 99.6594
R7578 gnd.n4751 gnd.n4750 99.6594
R7579 gnd.n4745 gnd.n4570 99.6594
R7580 gnd.n4743 gnd.n4742 99.6594
R7581 gnd.n4738 gnd.n4737 99.6594
R7582 gnd.n4735 gnd.n4734 99.6594
R7583 gnd.n4730 gnd.n4729 99.6594
R7584 gnd.n4727 gnd.n4726 99.6594
R7585 gnd.n4722 gnd.n4721 99.6594
R7586 gnd.n4719 gnd.n4718 99.6594
R7587 gnd.n4714 gnd.n4713 99.6594
R7588 gnd.n4711 gnd.n4710 99.6594
R7589 gnd.n4706 gnd.n4705 99.6594
R7590 gnd.n4703 gnd.n4702 99.6594
R7591 gnd.n4698 gnd.n4697 99.6594
R7592 gnd.n4695 gnd.n4694 99.6594
R7593 gnd.n4690 gnd.n4689 99.6594
R7594 gnd.n4687 gnd.n4686 99.6594
R7595 gnd.n4625 gnd.n4624 99.6594
R7596 gnd.n4678 gnd.n4677 99.6594
R7597 gnd.n5673 gnd.n5672 99.6594
R7598 gnd.n1260 gnd.n1252 99.6594
R7599 gnd.n5680 gnd.n5679 99.6594
R7600 gnd.n1251 gnd.n1245 99.6594
R7601 gnd.n5687 gnd.n5686 99.6594
R7602 gnd.n1244 gnd.n1238 99.6594
R7603 gnd.n5694 gnd.n5693 99.6594
R7604 gnd.n1237 gnd.n1231 99.6594
R7605 gnd.n5701 gnd.n5700 99.6594
R7606 gnd.n1230 gnd.n1223 99.6594
R7607 gnd.n5710 gnd.n5709 99.6594
R7608 gnd.n1219 gnd.n1213 99.6594
R7609 gnd.n5717 gnd.n5716 99.6594
R7610 gnd.n1212 gnd.n1206 99.6594
R7611 gnd.n5724 gnd.n5723 99.6594
R7612 gnd.n1205 gnd.n1198 99.6594
R7613 gnd.n5731 gnd.n5730 99.6594
R7614 gnd.n5734 gnd.n5733 99.6594
R7615 gnd.n7251 gnd.n534 99.6594
R7616 gnd.n7243 gnd.n505 99.6594
R7617 gnd.n7239 gnd.n506 99.6594
R7618 gnd.n7235 gnd.n507 99.6594
R7619 gnd.n7231 gnd.n508 99.6594
R7620 gnd.n7227 gnd.n509 99.6594
R7621 gnd.n7223 gnd.n510 99.6594
R7622 gnd.n7218 gnd.n512 99.6594
R7623 gnd.n7214 gnd.n513 99.6594
R7624 gnd.n7210 gnd.n514 99.6594
R7625 gnd.n7206 gnd.n515 99.6594
R7626 gnd.n7202 gnd.n516 99.6594
R7627 gnd.n7198 gnd.n517 99.6594
R7628 gnd.n7194 gnd.n518 99.6594
R7629 gnd.n7190 gnd.n519 99.6594
R7630 gnd.n7186 gnd.n520 99.6594
R7631 gnd.n574 gnd.n521 99.6594
R7632 gnd.n7178 gnd.n522 99.6594
R7633 gnd.n198 gnd.n195 99.6594
R7634 gnd.n7769 gnd.n7768 99.6594
R7635 gnd.n194 gnd.n188 99.6594
R7636 gnd.n7776 gnd.n7775 99.6594
R7637 gnd.n187 gnd.n181 99.6594
R7638 gnd.n7783 gnd.n7782 99.6594
R7639 gnd.n180 gnd.n174 99.6594
R7640 gnd.n7790 gnd.n7789 99.6594
R7641 gnd.n173 gnd.n167 99.6594
R7642 gnd.n7797 gnd.n7796 99.6594
R7643 gnd.n166 gnd.n160 99.6594
R7644 gnd.n7807 gnd.n7806 99.6594
R7645 gnd.n159 gnd.n153 99.6594
R7646 gnd.n7814 gnd.n7813 99.6594
R7647 gnd.n152 gnd.n146 99.6594
R7648 gnd.n7821 gnd.n7820 99.6594
R7649 gnd.n145 gnd.n139 99.6594
R7650 gnd.n7828 gnd.n7827 99.6594
R7651 gnd.n138 gnd.n135 99.6594
R7652 gnd.n5790 gnd.n5789 99.6594
R7653 gnd.n1128 gnd.n1105 99.6594
R7654 gnd.n1130 gnd.n1106 99.6594
R7655 gnd.n1138 gnd.n1107 99.6594
R7656 gnd.n1146 gnd.n1108 99.6594
R7657 gnd.n1148 gnd.n1109 99.6594
R7658 gnd.n1156 gnd.n1110 99.6594
R7659 gnd.n1166 gnd.n1111 99.6594
R7660 gnd.n1168 gnd.n1112 99.6594
R7661 gnd.n5123 gnd.n1113 99.6594
R7662 gnd.n5125 gnd.n1114 99.6594
R7663 gnd.n5129 gnd.n1115 99.6594
R7664 gnd.n5135 gnd.n1116 99.6594
R7665 gnd.n5793 gnd.n5792 99.6594
R7666 gnd.n5790 gnd.n1118 99.6594
R7667 gnd.n1129 gnd.n1105 99.6594
R7668 gnd.n1137 gnd.n1106 99.6594
R7669 gnd.n1145 gnd.n1107 99.6594
R7670 gnd.n1147 gnd.n1108 99.6594
R7671 gnd.n1155 gnd.n1109 99.6594
R7672 gnd.n1165 gnd.n1110 99.6594
R7673 gnd.n1167 gnd.n1111 99.6594
R7674 gnd.n5122 gnd.n1112 99.6594
R7675 gnd.n5124 gnd.n1113 99.6594
R7676 gnd.n5128 gnd.n1114 99.6594
R7677 gnd.n5130 gnd.n1115 99.6594
R7678 gnd.n1116 gnd.n1103 99.6594
R7679 gnd.n5792 gnd.n1100 99.6594
R7680 gnd.n6604 gnd.n640 99.6594
R7681 gnd.n6606 gnd.n641 99.6594
R7682 gnd.n6614 gnd.n642 99.6594
R7683 gnd.n6624 gnd.n643 99.6594
R7684 gnd.n6626 gnd.n644 99.6594
R7685 gnd.n6634 gnd.n645 99.6594
R7686 gnd.n6644 gnd.n646 99.6594
R7687 gnd.n6646 gnd.n647 99.6594
R7688 gnd.n6651 gnd.n648 99.6594
R7689 gnd.n6653 gnd.n649 99.6594
R7690 gnd.n6657 gnd.n650 99.6594
R7691 gnd.n6659 gnd.n651 99.6594
R7692 gnd.n6666 gnd.n652 99.6594
R7693 gnd.n654 gnd.n653 99.6594
R7694 gnd.n6667 gnd.n653 99.6594
R7695 gnd.n6660 gnd.n652 99.6594
R7696 gnd.n6658 gnd.n651 99.6594
R7697 gnd.n6654 gnd.n650 99.6594
R7698 gnd.n6652 gnd.n649 99.6594
R7699 gnd.n6647 gnd.n648 99.6594
R7700 gnd.n6645 gnd.n647 99.6594
R7701 gnd.n6635 gnd.n646 99.6594
R7702 gnd.n6627 gnd.n645 99.6594
R7703 gnd.n6625 gnd.n644 99.6594
R7704 gnd.n6615 gnd.n643 99.6594
R7705 gnd.n6607 gnd.n642 99.6594
R7706 gnd.n6605 gnd.n641 99.6594
R7707 gnd.n6732 gnd.n640 99.6594
R7708 gnd.n5131 gnd.t226 98.63
R7709 gnd.n122 gnd.t235 98.63
R7710 gnd.n6686 gnd.t249 98.63
R7711 gnd.n1161 gnd.t275 98.63
R7712 gnd.n554 gnd.t219 98.63
R7713 gnd.n576 gnd.t209 98.63
R7714 gnd.n201 gnd.t268 98.63
R7715 gnd.n7800 gnd.t189 98.63
R7716 gnd.n4594 gnd.t285 98.63
R7717 gnd.n4626 gnd.t263 98.63
R7718 gnd.n4449 gnd.t282 98.63
R7719 gnd.n1257 gnd.t278 98.63
R7720 gnd.n1220 gnd.t197 98.63
R7721 gnd.n6663 gnd.t193 98.63
R7722 gnd.n2473 gnd.n2472 97.3241
R7723 gnd.n2472 gnd.n2471 97.3241
R7724 gnd.n2471 gnd.n2147 97.3241
R7725 gnd.n2465 gnd.n2147 97.3241
R7726 gnd.n2465 gnd.n2464 97.3241
R7727 gnd.n2464 gnd.n2463 97.3241
R7728 gnd.n2463 gnd.n2154 97.3241
R7729 gnd.n2457 gnd.n2154 97.3241
R7730 gnd.n2457 gnd.n2456 97.3241
R7731 gnd.n2456 gnd.n2455 97.3241
R7732 gnd.n2455 gnd.n2162 97.3241
R7733 gnd.n2449 gnd.n2162 97.3241
R7734 gnd.n2449 gnd.n2448 97.3241
R7735 gnd.n2448 gnd.n2447 97.3241
R7736 gnd.n2447 gnd.n2170 97.3241
R7737 gnd.n2441 gnd.n2170 97.3241
R7738 gnd.n2441 gnd.n2440 97.3241
R7739 gnd.n2440 gnd.n2439 97.3241
R7740 gnd.n2439 gnd.n2178 97.3241
R7741 gnd.n2433 gnd.n2178 97.3241
R7742 gnd.n2433 gnd.n2432 97.3241
R7743 gnd.n2432 gnd.n2431 97.3241
R7744 gnd.n2431 gnd.n2186 97.3241
R7745 gnd.n2425 gnd.n2186 97.3241
R7746 gnd.n2425 gnd.n2424 97.3241
R7747 gnd.n2424 gnd.n2423 97.3241
R7748 gnd.n2423 gnd.n2194 97.3241
R7749 gnd.n2417 gnd.n2194 97.3241
R7750 gnd.n2417 gnd.n2416 97.3241
R7751 gnd.n2416 gnd.n2415 97.3241
R7752 gnd.n2415 gnd.n2202 97.3241
R7753 gnd.n2409 gnd.n2202 97.3241
R7754 gnd.n2409 gnd.n2408 97.3241
R7755 gnd.n2408 gnd.n2407 97.3241
R7756 gnd.n2407 gnd.n2210 97.3241
R7757 gnd.n2401 gnd.n2210 97.3241
R7758 gnd.n2401 gnd.n2400 97.3241
R7759 gnd.n2400 gnd.n2399 97.3241
R7760 gnd.n2399 gnd.n2218 97.3241
R7761 gnd.n2393 gnd.n2218 97.3241
R7762 gnd.n2393 gnd.n2392 97.3241
R7763 gnd.n2392 gnd.n2391 97.3241
R7764 gnd.n2391 gnd.n2226 97.3241
R7765 gnd.n2385 gnd.n2226 97.3241
R7766 gnd.n2385 gnd.n2384 97.3241
R7767 gnd.n2384 gnd.n2383 97.3241
R7768 gnd.n2383 gnd.n2234 97.3241
R7769 gnd.n2377 gnd.n2234 97.3241
R7770 gnd.n2377 gnd.n2376 97.3241
R7771 gnd.n2376 gnd.n2375 97.3241
R7772 gnd.n2375 gnd.n2242 97.3241
R7773 gnd.n2369 gnd.n2242 97.3241
R7774 gnd.n2369 gnd.n2368 97.3241
R7775 gnd.n2368 gnd.n2367 97.3241
R7776 gnd.n2367 gnd.n2250 97.3241
R7777 gnd.n2361 gnd.n2250 97.3241
R7778 gnd.n2361 gnd.n2360 97.3241
R7779 gnd.n2360 gnd.n2359 97.3241
R7780 gnd.n2359 gnd.n2258 97.3241
R7781 gnd.n2353 gnd.n2258 97.3241
R7782 gnd.n2353 gnd.n2352 97.3241
R7783 gnd.n2352 gnd.n2351 97.3241
R7784 gnd.n2351 gnd.n2266 97.3241
R7785 gnd.n2345 gnd.n2266 97.3241
R7786 gnd.n2345 gnd.n2344 97.3241
R7787 gnd.n2344 gnd.n2343 97.3241
R7788 gnd.n2343 gnd.n2274 97.3241
R7789 gnd.n2337 gnd.n2274 97.3241
R7790 gnd.n2337 gnd.n2336 97.3241
R7791 gnd.n2336 gnd.n2335 97.3241
R7792 gnd.n2335 gnd.n2282 97.3241
R7793 gnd.n2329 gnd.n2282 97.3241
R7794 gnd.n2329 gnd.n2328 97.3241
R7795 gnd.n2328 gnd.n2327 97.3241
R7796 gnd.n2327 gnd.n2290 97.3241
R7797 gnd.n2321 gnd.n2290 97.3241
R7798 gnd.n2321 gnd.n2320 97.3241
R7799 gnd.n2320 gnd.n2319 97.3241
R7800 gnd.n2319 gnd.n2298 97.3241
R7801 gnd.n2313 gnd.n2298 97.3241
R7802 gnd.n2313 gnd.n2312 97.3241
R7803 gnd.n2312 gnd.n2311 97.3241
R7804 gnd.n2311 gnd.n2306 97.3241
R7805 gnd.n5446 gnd.t243 92.8196
R7806 gnd.n6389 gnd.t258 92.8196
R7807 gnd.n5438 gnd.t291 92.8118
R7808 gnd.n6483 gnd.t204 92.8118
R7809 gnd.n5411 gnd.n5410 81.8399
R7810 gnd.n3464 gnd.t272 74.8376
R7811 gnd.n1604 gnd.t216 74.8376
R7812 gnd.n5447 gnd.t242 72.8438
R7813 gnd.n6390 gnd.t259 72.8438
R7814 gnd.n5412 gnd.n5405 72.8411
R7815 gnd.n5418 gnd.n5403 72.8411
R7816 gnd.n6422 gnd.n6421 72.8411
R7817 gnd.n5132 gnd.t225 72.836
R7818 gnd.n5439 gnd.t290 72.836
R7819 gnd.n6484 gnd.t205 72.836
R7820 gnd.n123 gnd.t236 72.836
R7821 gnd.n6687 gnd.t248 72.836
R7822 gnd.n1162 gnd.t276 72.836
R7823 gnd.n555 gnd.t218 72.836
R7824 gnd.n577 gnd.t208 72.836
R7825 gnd.n202 gnd.t269 72.836
R7826 gnd.n7801 gnd.t190 72.836
R7827 gnd.n4595 gnd.t284 72.836
R7828 gnd.n4627 gnd.t262 72.836
R7829 gnd.n4450 gnd.t281 72.836
R7830 gnd.n1258 gnd.t279 72.836
R7831 gnd.n1221 gnd.t198 72.836
R7832 gnd.n6664 gnd.t194 72.836
R7833 gnd.n6430 gnd.n6429 71.676
R7834 gnd.n6431 gnd.n6406 71.676
R7835 gnd.n6438 gnd.n6437 71.676
R7836 gnd.n6439 gnd.n6404 71.676
R7837 gnd.n6446 gnd.n6445 71.676
R7838 gnd.n6447 gnd.n6402 71.676
R7839 gnd.n6454 gnd.n6453 71.676
R7840 gnd.n6455 gnd.n6400 71.676
R7841 gnd.n6462 gnd.n6461 71.676
R7842 gnd.n6463 gnd.n6398 71.676
R7843 gnd.n6470 gnd.n6469 71.676
R7844 gnd.n6471 gnd.n6396 71.676
R7845 gnd.n6478 gnd.n6477 71.676
R7846 gnd.n6479 gnd.n6394 71.676
R7847 gnd.n6489 gnd.n6488 71.676
R7848 gnd.n6493 gnd.n6392 71.676
R7849 gnd.n6497 gnd.n6496 71.676
R7850 gnd.n6501 gnd.n6500 71.676
R7851 gnd.n6502 gnd.n6388 71.676
R7852 gnd.n6510 gnd.n6509 71.676
R7853 gnd.n6511 gnd.n6386 71.676
R7854 gnd.n6518 gnd.n6517 71.676
R7855 gnd.n6519 gnd.n6384 71.676
R7856 gnd.n6526 gnd.n6525 71.676
R7857 gnd.n6527 gnd.n6382 71.676
R7858 gnd.n6534 gnd.n6533 71.676
R7859 gnd.n6535 gnd.n6380 71.676
R7860 gnd.n6542 gnd.n6541 71.676
R7861 gnd.n6543 gnd.n6378 71.676
R7862 gnd.n6550 gnd.n6549 71.676
R7863 gnd.n6551 gnd.n6376 71.676
R7864 gnd.n6558 gnd.n6557 71.676
R7865 gnd.n6559 gnd.n6132 71.676
R7866 gnd.n5595 gnd.n5423 71.676
R7867 gnd.n5590 gnd.n5425 71.676
R7868 gnd.n5586 gnd.n5585 71.676
R7869 gnd.n5579 gnd.n5427 71.676
R7870 gnd.n5578 gnd.n5577 71.676
R7871 gnd.n5571 gnd.n5429 71.676
R7872 gnd.n5570 gnd.n5569 71.676
R7873 gnd.n5563 gnd.n5431 71.676
R7874 gnd.n5562 gnd.n5561 71.676
R7875 gnd.n5555 gnd.n5433 71.676
R7876 gnd.n5554 gnd.n5553 71.676
R7877 gnd.n5547 gnd.n5435 71.676
R7878 gnd.n5546 gnd.n5545 71.676
R7879 gnd.n5539 gnd.n5437 71.676
R7880 gnd.n5538 gnd.n5441 71.676
R7881 gnd.n5534 gnd.n5533 71.676
R7882 gnd.n5529 gnd.n5528 71.676
R7883 gnd.n5521 gnd.n5445 71.676
R7884 gnd.n5520 gnd.n5519 71.676
R7885 gnd.n5513 gnd.n5449 71.676
R7886 gnd.n5512 gnd.n5511 71.676
R7887 gnd.n5505 gnd.n5451 71.676
R7888 gnd.n5504 gnd.n5503 71.676
R7889 gnd.n5497 gnd.n5453 71.676
R7890 gnd.n5496 gnd.n5495 71.676
R7891 gnd.n5489 gnd.n5455 71.676
R7892 gnd.n5488 gnd.n5487 71.676
R7893 gnd.n5481 gnd.n5457 71.676
R7894 gnd.n5480 gnd.n5479 71.676
R7895 gnd.n5473 gnd.n5459 71.676
R7896 gnd.n5472 gnd.n5471 71.676
R7897 gnd.n5465 gnd.n5461 71.676
R7898 gnd.n5592 gnd.n5423 71.676
R7899 gnd.n5587 gnd.n5425 71.676
R7900 gnd.n5585 gnd.n5584 71.676
R7901 gnd.n5580 gnd.n5579 71.676
R7902 gnd.n5577 gnd.n5576 71.676
R7903 gnd.n5572 gnd.n5571 71.676
R7904 gnd.n5569 gnd.n5568 71.676
R7905 gnd.n5564 gnd.n5563 71.676
R7906 gnd.n5561 gnd.n5560 71.676
R7907 gnd.n5556 gnd.n5555 71.676
R7908 gnd.n5553 gnd.n5552 71.676
R7909 gnd.n5548 gnd.n5547 71.676
R7910 gnd.n5545 gnd.n5544 71.676
R7911 gnd.n5540 gnd.n5539 71.676
R7912 gnd.n5535 gnd.n5441 71.676
R7913 gnd.n5530 gnd.n5443 71.676
R7914 gnd.n5528 gnd.n5527 71.676
R7915 gnd.n5522 gnd.n5521 71.676
R7916 gnd.n5519 gnd.n5518 71.676
R7917 gnd.n5514 gnd.n5513 71.676
R7918 gnd.n5511 gnd.n5510 71.676
R7919 gnd.n5506 gnd.n5505 71.676
R7920 gnd.n5503 gnd.n5502 71.676
R7921 gnd.n5498 gnd.n5497 71.676
R7922 gnd.n5495 gnd.n5494 71.676
R7923 gnd.n5490 gnd.n5489 71.676
R7924 gnd.n5487 gnd.n5486 71.676
R7925 gnd.n5482 gnd.n5481 71.676
R7926 gnd.n5479 gnd.n5478 71.676
R7927 gnd.n5474 gnd.n5473 71.676
R7928 gnd.n5471 gnd.n5470 71.676
R7929 gnd.n5466 gnd.n5465 71.676
R7930 gnd.n6560 gnd.n6559 71.676
R7931 gnd.n6557 gnd.n6556 71.676
R7932 gnd.n6552 gnd.n6551 71.676
R7933 gnd.n6549 gnd.n6548 71.676
R7934 gnd.n6544 gnd.n6543 71.676
R7935 gnd.n6541 gnd.n6540 71.676
R7936 gnd.n6536 gnd.n6535 71.676
R7937 gnd.n6533 gnd.n6532 71.676
R7938 gnd.n6528 gnd.n6527 71.676
R7939 gnd.n6525 gnd.n6524 71.676
R7940 gnd.n6520 gnd.n6519 71.676
R7941 gnd.n6517 gnd.n6516 71.676
R7942 gnd.n6512 gnd.n6511 71.676
R7943 gnd.n6509 gnd.n6508 71.676
R7944 gnd.n6503 gnd.n6502 71.676
R7945 gnd.n6500 gnd.n6499 71.676
R7946 gnd.n6495 gnd.n6494 71.676
R7947 gnd.n6490 gnd.n6392 71.676
R7948 gnd.n6488 gnd.n6487 71.676
R7949 gnd.n6480 gnd.n6479 71.676
R7950 gnd.n6477 gnd.n6476 71.676
R7951 gnd.n6472 gnd.n6471 71.676
R7952 gnd.n6469 gnd.n6468 71.676
R7953 gnd.n6464 gnd.n6463 71.676
R7954 gnd.n6461 gnd.n6460 71.676
R7955 gnd.n6456 gnd.n6455 71.676
R7956 gnd.n6453 gnd.n6452 71.676
R7957 gnd.n6448 gnd.n6447 71.676
R7958 gnd.n6445 gnd.n6444 71.676
R7959 gnd.n6440 gnd.n6439 71.676
R7960 gnd.n6437 gnd.n6436 71.676
R7961 gnd.n6432 gnd.n6431 71.676
R7962 gnd.n6429 gnd.n6130 71.676
R7963 gnd.n10 gnd.t340 69.1507
R7964 gnd.n18 gnd.t165 68.4792
R7965 gnd.n17 gnd.t328 68.4792
R7966 gnd.n16 gnd.t112 68.4792
R7967 gnd.n15 gnd.t342 68.4792
R7968 gnd.n14 gnd.t101 68.4792
R7969 gnd.n13 gnd.t103 68.4792
R7970 gnd.n12 gnd.t319 68.4792
R7971 gnd.n11 gnd.t344 68.4792
R7972 gnd.n10 gnd.t67 68.4792
R7973 gnd.n3591 gnd.n3495 64.369
R7974 gnd.n5524 gnd.n5447 59.5399
R7975 gnd.n6505 gnd.n6390 59.5399
R7976 gnd.n5440 gnd.n5439 59.5399
R7977 gnd.n6485 gnd.n6484 59.5399
R7978 gnd.n5422 gnd.n5421 59.1804
R7979 gnd.n2306 gnd.n232 58.3947
R7980 gnd.n4443 gnd.n1564 57.3586
R7981 gnd.n3242 gnd.t145 56.607
R7982 gnd.n60 gnd.t93 56.607
R7983 gnd.n3203 gnd.t181 56.407
R7984 gnd.n3222 gnd.t8 56.407
R7985 gnd.n21 gnd.t87 56.407
R7986 gnd.n40 gnd.t127 56.407
R7987 gnd.n3259 gnd.t357 55.8337
R7988 gnd.n3220 gnd.t131 55.8337
R7989 gnd.n3239 gnd.t313 55.8337
R7990 gnd.n77 gnd.t155 55.8337
R7991 gnd.n38 gnd.t89 55.8337
R7992 gnd.n57 gnd.t297 55.8337
R7993 gnd.n5409 gnd.n5408 54.358
R7994 gnd.n6419 gnd.n6418 54.358
R7995 gnd.n3242 gnd.n3241 53.0052
R7996 gnd.n3244 gnd.n3243 53.0052
R7997 gnd.n3246 gnd.n3245 53.0052
R7998 gnd.n3248 gnd.n3247 53.0052
R7999 gnd.n3250 gnd.n3249 53.0052
R8000 gnd.n3252 gnd.n3251 53.0052
R8001 gnd.n3254 gnd.n3253 53.0052
R8002 gnd.n3256 gnd.n3255 53.0052
R8003 gnd.n3258 gnd.n3257 53.0052
R8004 gnd.n3203 gnd.n3202 53.0052
R8005 gnd.n3205 gnd.n3204 53.0052
R8006 gnd.n3207 gnd.n3206 53.0052
R8007 gnd.n3209 gnd.n3208 53.0052
R8008 gnd.n3211 gnd.n3210 53.0052
R8009 gnd.n3213 gnd.n3212 53.0052
R8010 gnd.n3215 gnd.n3214 53.0052
R8011 gnd.n3217 gnd.n3216 53.0052
R8012 gnd.n3219 gnd.n3218 53.0052
R8013 gnd.n3222 gnd.n3221 53.0052
R8014 gnd.n3224 gnd.n3223 53.0052
R8015 gnd.n3226 gnd.n3225 53.0052
R8016 gnd.n3228 gnd.n3227 53.0052
R8017 gnd.n3230 gnd.n3229 53.0052
R8018 gnd.n3232 gnd.n3231 53.0052
R8019 gnd.n3234 gnd.n3233 53.0052
R8020 gnd.n3236 gnd.n3235 53.0052
R8021 gnd.n3238 gnd.n3237 53.0052
R8022 gnd.n76 gnd.n75 53.0052
R8023 gnd.n74 gnd.n73 53.0052
R8024 gnd.n72 gnd.n71 53.0052
R8025 gnd.n70 gnd.n69 53.0052
R8026 gnd.n68 gnd.n67 53.0052
R8027 gnd.n66 gnd.n65 53.0052
R8028 gnd.n64 gnd.n63 53.0052
R8029 gnd.n62 gnd.n61 53.0052
R8030 gnd.n60 gnd.n59 53.0052
R8031 gnd.n37 gnd.n36 53.0052
R8032 gnd.n35 gnd.n34 53.0052
R8033 gnd.n33 gnd.n32 53.0052
R8034 gnd.n31 gnd.n30 53.0052
R8035 gnd.n29 gnd.n28 53.0052
R8036 gnd.n27 gnd.n26 53.0052
R8037 gnd.n25 gnd.n24 53.0052
R8038 gnd.n23 gnd.n22 53.0052
R8039 gnd.n21 gnd.n20 53.0052
R8040 gnd.n56 gnd.n55 53.0052
R8041 gnd.n54 gnd.n53 53.0052
R8042 gnd.n52 gnd.n51 53.0052
R8043 gnd.n50 gnd.n49 53.0052
R8044 gnd.n48 gnd.n47 53.0052
R8045 gnd.n46 gnd.n45 53.0052
R8046 gnd.n44 gnd.n43 53.0052
R8047 gnd.n42 gnd.n41 53.0052
R8048 gnd.n40 gnd.n39 53.0052
R8049 gnd.n6410 gnd.n6409 52.4801
R8050 gnd.n4295 gnd.t22 52.3082
R8051 gnd.n4263 gnd.t293 52.3082
R8052 gnd.n4231 gnd.t175 52.3082
R8053 gnd.n4200 gnd.t24 52.3082
R8054 gnd.n4168 gnd.t353 52.3082
R8055 gnd.n4136 gnd.t109 52.3082
R8056 gnd.n4104 gnd.t149 52.3082
R8057 gnd.n4073 gnd.t151 52.3082
R8058 gnd.n4758 gnd.n4444 51.6227
R8059 gnd.n7837 gnd.n128 51.6227
R8060 gnd.n4125 gnd.n4093 51.4173
R8061 gnd.n4189 gnd.n4188 50.455
R8062 gnd.n4157 gnd.n4156 50.455
R8063 gnd.n4125 gnd.n4124 50.455
R8064 gnd.n3538 gnd.n3537 45.1884
R8065 gnd.n1630 gnd.n1629 45.1884
R8066 gnd.n6426 gnd.n6425 44.3322
R8067 gnd.n5412 gnd.n5411 44.3189
R8068 gnd.n5133 gnd.n5132 42.4732
R8069 gnd.n6665 gnd.n6664 42.4732
R8070 gnd.n3539 gnd.n3538 42.2793
R8071 gnd.n1631 gnd.n1630 42.2793
R8072 gnd.n3465 gnd.n3464 42.2793
R8073 gnd.n4410 gnd.n1604 42.2793
R8074 gnd.n124 gnd.n123 42.2793
R8075 gnd.n6688 gnd.n6687 42.2793
R8076 gnd.n1163 gnd.n1162 42.2793
R8077 gnd.n578 gnd.n577 42.2793
R8078 gnd.n7765 gnd.n202 42.2793
R8079 gnd.n7802 gnd.n7801 42.2793
R8080 gnd.n4596 gnd.n4595 42.2793
R8081 gnd.n4628 gnd.n4627 42.2793
R8082 gnd.n4451 gnd.n4450 42.2793
R8083 gnd.n1259 gnd.n1258 42.2793
R8084 gnd.n5410 gnd.n5409 41.6274
R8085 gnd.n6420 gnd.n6419 41.6274
R8086 gnd.n5419 gnd.n5418 40.8975
R8087 gnd.n6423 gnd.n6422 40.8975
R8088 gnd.n7220 gnd.n555 36.9518
R8089 gnd.n1222 gnd.n1221 36.9518
R8090 gnd.n5418 gnd.n5417 35.055
R8091 gnd.n5413 gnd.n5412 35.055
R8092 gnd.n6412 gnd.n6411 35.055
R8093 gnd.n6422 gnd.n6408 35.055
R8094 gnd.n2845 gnd.n2844 33.6191
R8095 gnd.n2845 gnd.n1777 33.6191
R8096 gnd.n2853 gnd.n1777 33.6191
R8097 gnd.n2854 gnd.n2853 33.6191
R8098 gnd.n2855 gnd.n2854 33.6191
R8099 gnd.n2855 gnd.n1771 33.6191
R8100 gnd.n2863 gnd.n1771 33.6191
R8101 gnd.n2864 gnd.n2863 33.6191
R8102 gnd.n2865 gnd.n2864 33.6191
R8103 gnd.n2865 gnd.n1765 33.6191
R8104 gnd.n2873 gnd.n1765 33.6191
R8105 gnd.n2874 gnd.n2873 33.6191
R8106 gnd.n2875 gnd.n2874 33.6191
R8107 gnd.n2875 gnd.n1759 33.6191
R8108 gnd.n2883 gnd.n1759 33.6191
R8109 gnd.n2884 gnd.n2883 33.6191
R8110 gnd.n2885 gnd.n2884 33.6191
R8111 gnd.n2885 gnd.n1753 33.6191
R8112 gnd.n2893 gnd.n1753 33.6191
R8113 gnd.n2894 gnd.n2893 33.6191
R8114 gnd.n2895 gnd.n2894 33.6191
R8115 gnd.n2895 gnd.n1747 33.6191
R8116 gnd.n2903 gnd.n1747 33.6191
R8117 gnd.n2904 gnd.n2903 33.6191
R8118 gnd.n2905 gnd.n2904 33.6191
R8119 gnd.n2905 gnd.n1741 33.6191
R8120 gnd.n2913 gnd.n1741 33.6191
R8121 gnd.n2914 gnd.n2913 33.6191
R8122 gnd.n2915 gnd.n2914 33.6191
R8123 gnd.n2915 gnd.n1735 33.6191
R8124 gnd.n2923 gnd.n1735 33.6191
R8125 gnd.n2924 gnd.n2923 33.6191
R8126 gnd.n2925 gnd.n2924 33.6191
R8127 gnd.n2925 gnd.n1729 33.6191
R8128 gnd.n2933 gnd.n1729 33.6191
R8129 gnd.n2934 gnd.n2933 33.6191
R8130 gnd.n2935 gnd.n2934 33.6191
R8131 gnd.n2935 gnd.n1723 33.6191
R8132 gnd.n2943 gnd.n1723 33.6191
R8133 gnd.n2944 gnd.n2943 33.6191
R8134 gnd.n2945 gnd.n2944 33.6191
R8135 gnd.n2945 gnd.n1717 33.6191
R8136 gnd.n2953 gnd.n1717 33.6191
R8137 gnd.n2954 gnd.n2953 33.6191
R8138 gnd.n2955 gnd.n2954 33.6191
R8139 gnd.n2955 gnd.n1711 33.6191
R8140 gnd.n2963 gnd.n1711 33.6191
R8141 gnd.n2964 gnd.n2963 33.6191
R8142 gnd.n2965 gnd.n2964 33.6191
R8143 gnd.n2965 gnd.n1705 33.6191
R8144 gnd.n2973 gnd.n1705 33.6191
R8145 gnd.n2974 gnd.n2973 33.6191
R8146 gnd.n2975 gnd.n2974 33.6191
R8147 gnd.n2975 gnd.n1699 33.6191
R8148 gnd.n2983 gnd.n1699 33.6191
R8149 gnd.n2984 gnd.n2983 33.6191
R8150 gnd.n2985 gnd.n2984 33.6191
R8151 gnd.n2985 gnd.n1693 33.6191
R8152 gnd.n2993 gnd.n1693 33.6191
R8153 gnd.n2994 gnd.n2993 33.6191
R8154 gnd.n2995 gnd.n2994 33.6191
R8155 gnd.n2995 gnd.n1687 33.6191
R8156 gnd.n3003 gnd.n1687 33.6191
R8157 gnd.n3004 gnd.n3003 33.6191
R8158 gnd.n3005 gnd.n3004 33.6191
R8159 gnd.n3005 gnd.n1681 33.6191
R8160 gnd.n3013 gnd.n1681 33.6191
R8161 gnd.n3014 gnd.n3013 33.6191
R8162 gnd.n3015 gnd.n3014 33.6191
R8163 gnd.n3015 gnd.n1675 33.6191
R8164 gnd.n3023 gnd.n1675 33.6191
R8165 gnd.n3024 gnd.n3023 33.6191
R8166 gnd.n3025 gnd.n3024 33.6191
R8167 gnd.n3025 gnd.n1669 33.6191
R8168 gnd.n3033 gnd.n1669 33.6191
R8169 gnd.n3034 gnd.n3033 33.6191
R8170 gnd.n3035 gnd.n3034 33.6191
R8171 gnd.n3035 gnd.n1663 33.6191
R8172 gnd.n3043 gnd.n1663 33.6191
R8173 gnd.n3044 gnd.n3043 33.6191
R8174 gnd.n3045 gnd.n3044 33.6191
R8175 gnd.n3045 gnd.n1656 33.6191
R8176 gnd.n3060 gnd.n1656 33.6191
R8177 gnd.n3601 gnd.n3495 31.8661
R8178 gnd.n3601 gnd.n3600 31.8661
R8179 gnd.n3609 gnd.n3484 31.8661
R8180 gnd.n3617 gnd.n3484 31.8661
R8181 gnd.n3617 gnd.n3478 31.8661
R8182 gnd.n3625 gnd.n3478 31.8661
R8183 gnd.n3625 gnd.n3471 31.8661
R8184 gnd.n3663 gnd.n3471 31.8661
R8185 gnd.n3673 gnd.n3404 31.8661
R8186 gnd.n4758 gnd.n4566 31.8661
R8187 gnd.n4766 gnd.n1550 31.8661
R8188 gnd.n4774 gnd.n1550 31.8661
R8189 gnd.n4774 gnd.n1542 31.8661
R8190 gnd.n4782 gnd.n1542 31.8661
R8191 gnd.n4790 gnd.n1533 31.8661
R8192 gnd.n4790 gnd.n1536 31.8661
R8193 gnd.n4798 gnd.n1518 31.8661
R8194 gnd.n4806 gnd.n1518 31.8661
R8195 gnd.n4814 gnd.n1510 31.8661
R8196 gnd.n4822 gnd.n1501 31.8661
R8197 gnd.n4822 gnd.n1504 31.8661
R8198 gnd.n4838 gnd.n1484 31.8661
R8199 gnd.n4848 gnd.n1484 31.8661
R8200 gnd.n4861 gnd.n1478 31.8661
R8201 gnd.n4879 gnd.n1460 31.8661
R8202 gnd.n4873 gnd.n1460 31.8661
R8203 gnd.n4888 gnd.n1443 31.8661
R8204 gnd.n4901 gnd.n1443 31.8661
R8205 gnd.n5238 gnd.n1395 31.8661
R8206 gnd.n5077 gnd.n1177 31.8661
R8207 gnd.n5075 gnd.n5074 31.8661
R8208 gnd.n5074 gnd.n1104 31.8661
R8209 gnd.n5800 gnd.n1097 31.8661
R8210 gnd.n5800 gnd.n1099 31.8661
R8211 gnd.n5808 gnd.n1084 31.8661
R8212 gnd.n5816 gnd.n1084 31.8661
R8213 gnd.n5816 gnd.n1077 31.8661
R8214 gnd.n5824 gnd.n1077 31.8661
R8215 gnd.n5832 gnd.n1070 31.8661
R8216 gnd.n5832 gnd.n1062 31.8661
R8217 gnd.n5840 gnd.n1062 31.8661
R8218 gnd.n5840 gnd.n1064 31.8661
R8219 gnd.n5848 gnd.n1048 31.8661
R8220 gnd.n5856 gnd.n1048 31.8661
R8221 gnd.n5856 gnd.n1050 31.8661
R8222 gnd.n7001 gnd.n718 31.8661
R8223 gnd.n7009 gnd.n704 31.8661
R8224 gnd.n7017 gnd.n704 31.8661
R8225 gnd.n7017 gnd.n706 31.8661
R8226 gnd.n7025 gnd.n691 31.8661
R8227 gnd.n7033 gnd.n691 31.8661
R8228 gnd.n7033 gnd.n684 31.8661
R8229 gnd.n7041 gnd.n684 31.8661
R8230 gnd.n7049 gnd.n677 31.8661
R8231 gnd.n7049 gnd.n669 31.8661
R8232 gnd.n7058 gnd.n669 31.8661
R8233 gnd.n7058 gnd.n671 31.8661
R8234 gnd.n7068 gnd.n662 31.8661
R8235 gnd.n662 gnd.n639 31.8661
R8236 gnd.n7078 gnd.n7077 31.8661
R8237 gnd.n7077 gnd.n504 31.8661
R8238 gnd.n581 gnd.n532 31.8661
R8239 gnd.n7565 gnd.n333 31.8661
R8240 gnd.n7569 gnd.n298 31.8661
R8241 gnd.n7593 gnd.n298 31.8661
R8242 gnd.n7601 gnd.n289 31.8661
R8243 gnd.n7601 gnd.n292 31.8661
R8244 gnd.n7609 gnd.n283 31.8661
R8245 gnd.n7617 gnd.n268 31.8661
R8246 gnd.n7625 gnd.n268 31.8661
R8247 gnd.n7633 gnd.n259 31.8661
R8248 gnd.n7633 gnd.n262 31.8661
R8249 gnd.n7641 gnd.n253 31.8661
R8250 gnd.n7649 gnd.n238 31.8661
R8251 gnd.n7657 gnd.n238 31.8661
R8252 gnd.n7665 gnd.n229 31.8661
R8253 gnd.n7673 gnd.n213 31.8661
R8254 gnd.n7749 gnd.n213 31.8661
R8255 gnd.n7749 gnd.n206 31.8661
R8256 gnd.n7757 gnd.n206 31.8661
R8257 gnd.n7837 gnd.n126 31.8661
R8258 gnd.n6563 gnd.n6562 31.3761
R8259 gnd.n5467 gnd.n5463 31.3761
R8260 gnd.t132 gnd.n1478 30.9101
R8261 gnd.n5864 gnd.n1042 30.9101
R8262 gnd.n283 gnd.t96 30.9101
R8263 gnd.n5374 gnd.t265 30.5915
R8264 gnd.t73 gnd.n1510 30.2728
R8265 gnd.n253 gnd.t9 30.2728
R8266 gnd.n4566 gnd.t261 28.3609
R8267 gnd.t188 gnd.n126 28.3609
R8268 gnd.n1050 gnd.t316 27.0862
R8269 gnd.n7009 gnd.t327 27.0862
R8270 gnd.n6578 gnd.t221 26.1303
R8271 gnd.n5132 gnd.n5131 25.7944
R8272 gnd.n3464 gnd.n3463 25.7944
R8273 gnd.n1604 gnd.n1603 25.7944
R8274 gnd.n123 gnd.n122 25.7944
R8275 gnd.n6687 gnd.n6686 25.7944
R8276 gnd.n1162 gnd.n1161 25.7944
R8277 gnd.n555 gnd.n554 25.7944
R8278 gnd.n577 gnd.n576 25.7944
R8279 gnd.n202 gnd.n201 25.7944
R8280 gnd.n7801 gnd.n7800 25.7944
R8281 gnd.n4595 gnd.n4594 25.7944
R8282 gnd.n4627 gnd.n4626 25.7944
R8283 gnd.n4450 gnd.n4449 25.7944
R8284 gnd.n1258 gnd.n1257 25.7944
R8285 gnd.n1221 gnd.n1220 25.7944
R8286 gnd.n6664 gnd.n6663 25.7944
R8287 gnd.n3685 gnd.n3405 24.8557
R8288 gnd.n3695 gnd.n3388 24.8557
R8289 gnd.n3391 gnd.n3379 24.8557
R8290 gnd.n3716 gnd.n3380 24.8557
R8291 gnd.n3726 gnd.n3360 24.8557
R8292 gnd.n3736 gnd.n3735 24.8557
R8293 gnd.n3346 gnd.n3344 24.8557
R8294 gnd.n3767 gnd.n3766 24.8557
R8295 gnd.n3782 gnd.n3329 24.8557
R8296 gnd.n3836 gnd.n3268 24.8557
R8297 gnd.n3792 gnd.n3269 24.8557
R8298 gnd.n3829 gnd.n3280 24.8557
R8299 gnd.n3318 gnd.n3317 24.8557
R8300 gnd.n3823 gnd.n3822 24.8557
R8301 gnd.n3304 gnd.n3291 24.8557
R8302 gnd.n3862 gnd.n3861 24.8557
R8303 gnd.n3872 gnd.n3188 24.8557
R8304 gnd.n3884 gnd.n3180 24.8557
R8305 gnd.n3883 gnd.n3168 24.8557
R8306 gnd.n3902 gnd.n3901 24.8557
R8307 gnd.n3912 gnd.n3161 24.8557
R8308 gnd.n3923 gnd.n3149 24.8557
R8309 gnd.n3947 gnd.n3946 24.8557
R8310 gnd.n3958 gnd.n3132 24.8557
R8311 gnd.n3957 gnd.n3134 24.8557
R8312 gnd.n3969 gnd.n3125 24.8557
R8313 gnd.n3987 gnd.n3986 24.8557
R8314 gnd.n3116 gnd.n3105 24.8557
R8315 gnd.n4008 gnd.n3093 24.8557
R8316 gnd.n4036 gnd.n4035 24.8557
R8317 gnd.n4047 gnd.n3078 24.8557
R8318 gnd.n4058 gnd.n3071 24.8557
R8319 gnd.n4057 gnd.n1653 24.8557
R8320 gnd.n4330 gnd.n4329 24.8557
R8321 gnd.n4352 gnd.n1638 24.8557
R8322 gnd.n1099 gnd.t224 24.537
R8323 gnd.n5848 gnd.t339 24.537
R8324 gnd.n706 gnd.t362 24.537
R8325 gnd.n7068 gnd.t192 24.537
R8326 gnd.n5227 gnd.n1406 24.2183
R8327 gnd.n5226 gnd.n1412 24.2183
R8328 gnd.n5220 gnd.n5219 24.2183
R8329 gnd.n5246 gnd.n1377 24.2183
R8330 gnd.n4993 gnd.n1380 24.2183
R8331 gnd.n4997 gnd.n1371 24.2183
R8332 gnd.n5262 gnd.n1360 24.2183
R8333 gnd.n5270 gnd.n1351 24.2183
R8334 gnd.n5278 gnd.n1342 24.2183
R8335 gnd.n5033 gnd.n1345 24.2183
R8336 gnd.n5027 gnd.n1336 24.2183
R8337 gnd.n5294 gnd.n1325 24.2183
R8338 gnd.n5302 gnd.n1316 24.2183
R8339 gnd.n5310 gnd.n1307 24.2183
R8340 gnd.n5097 gnd.n1310 24.2183
R8341 gnd.n5103 gnd.n1301 24.2183
R8342 gnd.n5326 gnd.n1290 24.2183
R8343 gnd.n5334 gnd.n1281 24.2183
R8344 gnd.n5118 gnd.n1284 24.2183
R8345 gnd.n5344 gnd.n1271 24.2183
R8346 gnd.n5152 gnd.n1274 24.2183
R8347 gnd.n5664 gnd.n1265 24.2183
R8348 gnd.n5741 gnd.n1175 24.2183
R8349 gnd.n7176 gnd.n495 24.2183
R8350 gnd.n7261 gnd.n498 24.2183
R8351 gnd.n601 gnd.n486 24.2183
R8352 gnd.n7269 gnd.n489 24.2183
R8353 gnd.n607 gnd.n477 24.2183
R8354 gnd.n7277 gnd.n480 24.2183
R8355 gnd.n7285 gnd.n471 24.2183
R8356 gnd.n617 gnd.n460 24.2183
R8357 gnd.n7128 gnd.n451 24.2183
R8358 gnd.n7301 gnd.n454 24.2183
R8359 gnd.n7315 gnd.n443 24.2183
R8360 gnd.n7325 gnd.n432 24.2183
R8361 gnd.n7342 gnd.n422 24.2183
R8362 gnd.n7391 gnd.n408 24.2183
R8363 gnd.n7332 gnd.n396 24.2183
R8364 gnd.n7382 gnd.n390 24.2183
R8365 gnd.n7438 gnd.n376 24.2183
R8366 gnd.n7409 gnd.n383 24.2183
R8367 gnd.n7447 gnd.n364 24.2183
R8368 gnd.n7427 gnd.n356 24.2183
R8369 gnd.n7584 gnd.n314 24.2183
R8370 gnd.n7549 gnd.n7548 24.2183
R8371 gnd.n7556 gnd.n343 24.2183
R8372 gnd.t171 gnd.n1425 23.8997
R8373 gnd.n5791 gnd.n1097 23.8997
R8374 gnd.n7076 gnd.n639 23.8997
R8375 gnd.t59 gnd.n311 23.8997
R8376 gnd.n3706 gnd.t150 23.2624
R8377 gnd.n4782 gnd.t130 23.2624
R8378 gnd.t98 gnd.n1354 23.2624
R8379 gnd.n5107 gnd.t7 23.2624
R8380 gnd.n611 gnd.t86 23.2624
R8381 gnd.n7381 gnd.t27 23.2624
R8382 gnd.n7673 gnd.t88 23.2624
R8383 gnd.n3407 gnd.t271 22.6251
R8384 gnd.n4814 gnd.t77 22.6251
R8385 gnd.n5023 gnd.t36 22.6251
R8386 gnd.t146 gnd.n1319 22.6251
R8387 gnd.t19 gnd.n440 22.6251
R8388 gnd.n7145 gnd.t90 22.6251
R8389 gnd.n7641 gnd.t81 22.6251
R8390 gnd.n4861 gnd.t40 21.9878
R8391 gnd.n5003 gnd.t157 21.9878
R8392 gnd.n7415 gnd.t17 21.9878
R8393 gnd.n7609 gnd.t42 21.9878
R8394 gnd.n5400 gnd.n1035 21.6691
R8395 gnd.n5970 gnd.n981 21.6691
R8396 gnd.n5934 gnd.n965 21.6691
R8397 gnd.n5943 gnd.n955 21.6691
R8398 gnd.n6032 gnd.n939 21.6691
R8399 gnd.n933 gnd.n919 21.6691
R8400 gnd.n6040 gnd.n909 21.6691
R8401 gnd.n6833 gnd.n883 21.6691
R8402 gnd.n6242 gnd.n854 21.6691
R8403 gnd.n6280 gnd.n812 21.6691
R8404 gnd.n6289 gnd.n805 21.6691
R8405 gnd.n6298 gnd.n797 21.6691
R8406 gnd.n6307 gnd.n789 21.6691
R8407 gnd.n6316 gnd.n781 21.6691
R8408 gnd.n6325 gnd.n773 21.6691
R8409 gnd.n6342 gnd.n757 21.6691
R8410 gnd.n6969 gnd.n750 21.6691
R8411 gnd.n6136 gnd.n742 21.6691
R8412 gnd.t23 gnd.n3412 21.3504
R8413 gnd.n1422 gnd.t162 21.3504
R8414 gnd.n7533 gnd.t75 21.3504
R8415 gnd.t232 gnd.n1020 21.0318
R8416 gnd.t48 gnd.n3106 20.7131
R8417 gnd.n4888 gnd.t69 20.7131
R8418 gnd.n7593 gnd.t84 20.7131
R8419 gnd.t123 gnd.n1392 20.3945
R8420 gnd.n5612 gnd.n1010 20.3945
R8421 gnd.n5986 gnd.n979 20.3945
R8422 gnd.n6961 gnd.n759 20.3945
R8423 gnd.n7564 gnd.t63 20.3945
R8424 gnd.n3061 gnd.n3060 20.1716
R8425 gnd.t12 gnd.n3141 20.0758
R8426 gnd.n4838 gnd.t79 20.0758
R8427 gnd.t343 gnd.n973 20.0758
R8428 gnd.t115 gnd.n765 20.0758
R8429 gnd.n7625 gnd.t55 20.0758
R8430 gnd.n5447 gnd.n5446 19.9763
R8431 gnd.n6390 gnd.n6389 19.9763
R8432 gnd.n5439 gnd.n5438 19.9763
R8433 gnd.n6484 gnd.n6483 19.9763
R8434 gnd.n5406 gnd.t233 19.8005
R8435 gnd.n5406 gnd.t246 19.8005
R8436 gnd.n5407 gnd.t212 19.8005
R8437 gnd.n5407 gnd.t256 19.8005
R8438 gnd.n6416 gnd.t239 19.8005
R8439 gnd.n6416 gnd.t222 19.8005
R8440 gnd.n6417 gnd.t186 19.8005
R8441 gnd.n6417 gnd.t288 19.8005
R8442 gnd.n5075 gnd.n1196 19.7572
R8443 gnd.n7252 gnd.n504 19.7572
R8444 gnd.n5403 gnd.n5402 19.5087
R8445 gnd.n5416 gnd.n5403 19.5087
R8446 gnd.n5414 gnd.n5405 19.5087
R8447 gnd.n6421 gnd.n6415 19.5087
R8448 gnd.n3873 gnd.t321 19.4385
R8449 gnd.n4798 gnd.t31 19.4385
R8450 gnd.n5824 gnd.t153 19.4385
R8451 gnd.t164 gnd.n677 19.4385
R8452 gnd.n7657 gnd.t135 19.4385
R8453 gnd.n5798 gnd.n1089 19.3944
R8454 gnd.n5810 gnd.n1089 19.3944
R8455 gnd.n5810 gnd.n1087 19.3944
R8456 gnd.n5814 gnd.n1087 19.3944
R8457 gnd.n5814 gnd.n1075 19.3944
R8458 gnd.n5826 gnd.n1075 19.3944
R8459 gnd.n5826 gnd.n1073 19.3944
R8460 gnd.n5830 gnd.n1073 19.3944
R8461 gnd.n5830 gnd.n1060 19.3944
R8462 gnd.n5842 gnd.n1060 19.3944
R8463 gnd.n5842 gnd.n1058 19.3944
R8464 gnd.n5846 gnd.n1058 19.3944
R8465 gnd.n5846 gnd.n1046 19.3944
R8466 gnd.n5858 gnd.n1046 19.3944
R8467 gnd.n5858 gnd.n1044 19.3944
R8468 gnd.n5862 gnd.n1044 19.3944
R8469 gnd.n5862 gnd.n1032 19.3944
R8470 gnd.n5874 gnd.n1032 19.3944
R8471 gnd.n5874 gnd.n1030 19.3944
R8472 gnd.n5878 gnd.n1030 19.3944
R8473 gnd.n5878 gnd.n1016 19.3944
R8474 gnd.n5892 gnd.n1016 19.3944
R8475 gnd.n5892 gnd.n1013 19.3944
R8476 gnd.n5897 gnd.n1013 19.3944
R8477 gnd.n5897 gnd.n1014 19.3944
R8478 gnd.n1014 gnd.n977 19.3944
R8479 gnd.n5988 gnd.n977 19.3944
R8480 gnd.n5988 gnd.n975 19.3944
R8481 gnd.n5992 gnd.n975 19.3944
R8482 gnd.n5992 gnd.n961 19.3944
R8483 gnd.n6004 gnd.n961 19.3944
R8484 gnd.n6004 gnd.n958 19.3944
R8485 gnd.n6011 gnd.n958 19.3944
R8486 gnd.n6011 gnd.n959 19.3944
R8487 gnd.n6007 gnd.n959 19.3944
R8488 gnd.n6007 gnd.n922 19.3944
R8489 gnd.n6067 gnd.n922 19.3944
R8490 gnd.n6067 gnd.n923 19.3944
R8491 gnd.n6063 gnd.n923 19.3944
R8492 gnd.n6063 gnd.n6062 19.3944
R8493 gnd.n6062 gnd.n6061 19.3944
R8494 gnd.n6061 gnd.n6058 19.3944
R8495 gnd.n6058 gnd.n874 19.3944
R8496 gnd.n6843 gnd.n874 19.3944
R8497 gnd.n6843 gnd.n872 19.3944
R8498 gnd.n6847 gnd.n872 19.3944
R8499 gnd.n6847 gnd.n858 19.3944
R8500 gnd.n6859 gnd.n858 19.3944
R8501 gnd.n6859 gnd.n856 19.3944
R8502 gnd.n6863 gnd.n856 19.3944
R8503 gnd.n6863 gnd.n842 19.3944
R8504 gnd.n6875 gnd.n842 19.3944
R8505 gnd.n6875 gnd.n840 19.3944
R8506 gnd.n6879 gnd.n840 19.3944
R8507 gnd.n6879 gnd.n826 19.3944
R8508 gnd.n6891 gnd.n826 19.3944
R8509 gnd.n6891 gnd.n824 19.3944
R8510 gnd.n6895 gnd.n824 19.3944
R8511 gnd.n6895 gnd.n810 19.3944
R8512 gnd.n6907 gnd.n810 19.3944
R8513 gnd.n6907 gnd.n808 19.3944
R8514 gnd.n6911 gnd.n808 19.3944
R8515 gnd.n6911 gnd.n795 19.3944
R8516 gnd.n6923 gnd.n795 19.3944
R8517 gnd.n6923 gnd.n793 19.3944
R8518 gnd.n6927 gnd.n793 19.3944
R8519 gnd.n6927 gnd.n779 19.3944
R8520 gnd.n6939 gnd.n779 19.3944
R8521 gnd.n6939 gnd.n777 19.3944
R8522 gnd.n6943 gnd.n777 19.3944
R8523 gnd.n6943 gnd.n763 19.3944
R8524 gnd.n6955 gnd.n763 19.3944
R8525 gnd.n6955 gnd.n761 19.3944
R8526 gnd.n6959 gnd.n761 19.3944
R8527 gnd.n6959 gnd.n746 19.3944
R8528 gnd.n6971 gnd.n746 19.3944
R8529 gnd.n6971 gnd.n744 19.3944
R8530 gnd.n6975 gnd.n744 19.3944
R8531 gnd.n6975 gnd.n732 19.3944
R8532 gnd.n6987 gnd.n732 19.3944
R8533 gnd.n6987 gnd.n730 19.3944
R8534 gnd.n6991 gnd.n730 19.3944
R8535 gnd.n6991 gnd.n716 19.3944
R8536 gnd.n7003 gnd.n716 19.3944
R8537 gnd.n7003 gnd.n714 19.3944
R8538 gnd.n7007 gnd.n714 19.3944
R8539 gnd.n7007 gnd.n702 19.3944
R8540 gnd.n7019 gnd.n702 19.3944
R8541 gnd.n7019 gnd.n700 19.3944
R8542 gnd.n7023 gnd.n700 19.3944
R8543 gnd.n7023 gnd.n689 19.3944
R8544 gnd.n7035 gnd.n689 19.3944
R8545 gnd.n7035 gnd.n687 19.3944
R8546 gnd.n7039 gnd.n687 19.3944
R8547 gnd.n7039 gnd.n675 19.3944
R8548 gnd.n7051 gnd.n675 19.3944
R8549 gnd.n7051 gnd.n673 19.3944
R8550 gnd.n7056 gnd.n673 19.3944
R8551 gnd.n7056 gnd.n659 19.3944
R8552 gnd.n7070 gnd.n659 19.3944
R8553 gnd.n7071 gnd.n7070 19.3944
R8554 gnd.n5136 gnd.n1102 19.3944
R8555 gnd.n5794 gnd.n1102 19.3944
R8556 gnd.n5795 gnd.n5794 19.3944
R8557 gnd.n5788 gnd.n5787 19.3944
R8558 gnd.n5787 gnd.n1120 19.3944
R8559 gnd.n5780 gnd.n1120 19.3944
R8560 gnd.n5780 gnd.n5779 19.3944
R8561 gnd.n5779 gnd.n1131 19.3944
R8562 gnd.n5772 gnd.n1131 19.3944
R8563 gnd.n5772 gnd.n5771 19.3944
R8564 gnd.n5771 gnd.n1139 19.3944
R8565 gnd.n5764 gnd.n1139 19.3944
R8566 gnd.n5764 gnd.n5763 19.3944
R8567 gnd.n5763 gnd.n1149 19.3944
R8568 gnd.n5756 gnd.n1149 19.3944
R8569 gnd.n5756 gnd.n5755 19.3944
R8570 gnd.n5755 gnd.n1157 19.3944
R8571 gnd.n5748 gnd.n1157 19.3944
R8572 gnd.n5748 gnd.n5747 19.3944
R8573 gnd.n5747 gnd.n1169 19.3944
R8574 gnd.n5147 gnd.n1169 19.3944
R8575 gnd.n5147 gnd.n5146 19.3944
R8576 gnd.n5146 gnd.n5145 19.3944
R8577 gnd.n5145 gnd.n5126 19.3944
R8578 gnd.n5141 gnd.n5126 19.3944
R8579 gnd.n5141 gnd.n5140 19.3944
R8580 gnd.n5140 gnd.n5139 19.3944
R8581 gnd.n3588 gnd.n3587 19.3944
R8582 gnd.n3587 gnd.n3586 19.3944
R8583 gnd.n3586 gnd.n3585 19.3944
R8584 gnd.n3585 gnd.n3583 19.3944
R8585 gnd.n3583 gnd.n3580 19.3944
R8586 gnd.n3580 gnd.n3579 19.3944
R8587 gnd.n3579 gnd.n3576 19.3944
R8588 gnd.n3576 gnd.n3575 19.3944
R8589 gnd.n3575 gnd.n3572 19.3944
R8590 gnd.n3572 gnd.n3571 19.3944
R8591 gnd.n3571 gnd.n3568 19.3944
R8592 gnd.n3568 gnd.n3567 19.3944
R8593 gnd.n3567 gnd.n3564 19.3944
R8594 gnd.n3564 gnd.n3563 19.3944
R8595 gnd.n3563 gnd.n3560 19.3944
R8596 gnd.n3560 gnd.n3559 19.3944
R8597 gnd.n3559 gnd.n3556 19.3944
R8598 gnd.n3556 gnd.n3555 19.3944
R8599 gnd.n3555 gnd.n3552 19.3944
R8600 gnd.n3552 gnd.n3551 19.3944
R8601 gnd.n3551 gnd.n3548 19.3944
R8602 gnd.n3548 gnd.n3547 19.3944
R8603 gnd.n3544 gnd.n3543 19.3944
R8604 gnd.n3543 gnd.n3499 19.3944
R8605 gnd.n3594 gnd.n3499 19.3944
R8606 gnd.n4360 gnd.n4359 19.3944
R8607 gnd.n4359 gnd.n4356 19.3944
R8608 gnd.n4356 gnd.n4355 19.3944
R8609 gnd.n4405 gnd.n4404 19.3944
R8610 gnd.n4404 gnd.n4403 19.3944
R8611 gnd.n4403 gnd.n4400 19.3944
R8612 gnd.n4400 gnd.n4399 19.3944
R8613 gnd.n4399 gnd.n4396 19.3944
R8614 gnd.n4396 gnd.n4395 19.3944
R8615 gnd.n4395 gnd.n4392 19.3944
R8616 gnd.n4392 gnd.n4391 19.3944
R8617 gnd.n4391 gnd.n4388 19.3944
R8618 gnd.n4388 gnd.n4387 19.3944
R8619 gnd.n4387 gnd.n4384 19.3944
R8620 gnd.n4384 gnd.n4383 19.3944
R8621 gnd.n4383 gnd.n4380 19.3944
R8622 gnd.n4380 gnd.n4379 19.3944
R8623 gnd.n4379 gnd.n4376 19.3944
R8624 gnd.n4376 gnd.n4375 19.3944
R8625 gnd.n4375 gnd.n4372 19.3944
R8626 gnd.n4372 gnd.n4371 19.3944
R8627 gnd.n4371 gnd.n4368 19.3944
R8628 gnd.n4368 gnd.n4367 19.3944
R8629 gnd.n4367 gnd.n4364 19.3944
R8630 gnd.n4364 gnd.n4363 19.3944
R8631 gnd.n3687 gnd.n3396 19.3944
R8632 gnd.n3697 gnd.n3396 19.3944
R8633 gnd.n3698 gnd.n3697 19.3944
R8634 gnd.n3698 gnd.n3377 19.3944
R8635 gnd.n3718 gnd.n3377 19.3944
R8636 gnd.n3718 gnd.n3369 19.3944
R8637 gnd.n3728 gnd.n3369 19.3944
R8638 gnd.n3729 gnd.n3728 19.3944
R8639 gnd.n3730 gnd.n3729 19.3944
R8640 gnd.n3730 gnd.n3352 19.3944
R8641 gnd.n3747 gnd.n3352 19.3944
R8642 gnd.n3750 gnd.n3747 19.3944
R8643 gnd.n3750 gnd.n3749 19.3944
R8644 gnd.n3749 gnd.n3325 19.3944
R8645 gnd.n3789 gnd.n3325 19.3944
R8646 gnd.n3789 gnd.n3322 19.3944
R8647 gnd.n3795 gnd.n3322 19.3944
R8648 gnd.n3796 gnd.n3795 19.3944
R8649 gnd.n3796 gnd.n3320 19.3944
R8650 gnd.n3802 gnd.n3320 19.3944
R8651 gnd.n3805 gnd.n3802 19.3944
R8652 gnd.n3807 gnd.n3805 19.3944
R8653 gnd.n3813 gnd.n3807 19.3944
R8654 gnd.n3813 gnd.n3812 19.3944
R8655 gnd.n3812 gnd.n3183 19.3944
R8656 gnd.n3879 gnd.n3183 19.3944
R8657 gnd.n3880 gnd.n3879 19.3944
R8658 gnd.n3880 gnd.n3176 19.3944
R8659 gnd.n3891 gnd.n3176 19.3944
R8660 gnd.n3892 gnd.n3891 19.3944
R8661 gnd.n3892 gnd.n3159 19.3944
R8662 gnd.n3159 gnd.n3157 19.3944
R8663 gnd.n3916 gnd.n3157 19.3944
R8664 gnd.n3917 gnd.n3916 19.3944
R8665 gnd.n3917 gnd.n3128 19.3944
R8666 gnd.n3964 gnd.n3128 19.3944
R8667 gnd.n3965 gnd.n3964 19.3944
R8668 gnd.n3965 gnd.n3121 19.3944
R8669 gnd.n3976 gnd.n3121 19.3944
R8670 gnd.n3977 gnd.n3976 19.3944
R8671 gnd.n3977 gnd.n3104 19.3944
R8672 gnd.n3104 gnd.n3102 19.3944
R8673 gnd.n4001 gnd.n3102 19.3944
R8674 gnd.n4002 gnd.n4001 19.3944
R8675 gnd.n4002 gnd.n3074 19.3944
R8676 gnd.n4053 gnd.n3074 19.3944
R8677 gnd.n4054 gnd.n4053 19.3944
R8678 gnd.n4054 gnd.n3067 19.3944
R8679 gnd.n4321 gnd.n3067 19.3944
R8680 gnd.n4322 gnd.n4321 19.3944
R8681 gnd.n4322 gnd.n1642 19.3944
R8682 gnd.n4347 gnd.n1642 19.3944
R8683 gnd.n4347 gnd.n1643 19.3944
R8684 gnd.n3678 gnd.n3677 19.3944
R8685 gnd.n3677 gnd.n3410 19.3944
R8686 gnd.n3433 gnd.n3410 19.3944
R8687 gnd.n3436 gnd.n3433 19.3944
R8688 gnd.n3436 gnd.n3429 19.3944
R8689 gnd.n3440 gnd.n3429 19.3944
R8690 gnd.n3443 gnd.n3440 19.3944
R8691 gnd.n3446 gnd.n3443 19.3944
R8692 gnd.n3446 gnd.n3427 19.3944
R8693 gnd.n3450 gnd.n3427 19.3944
R8694 gnd.n3453 gnd.n3450 19.3944
R8695 gnd.n3456 gnd.n3453 19.3944
R8696 gnd.n3456 gnd.n3425 19.3944
R8697 gnd.n3460 gnd.n3425 19.3944
R8698 gnd.n3683 gnd.n3682 19.3944
R8699 gnd.n3682 gnd.n3386 19.3944
R8700 gnd.n3708 gnd.n3386 19.3944
R8701 gnd.n3708 gnd.n3384 19.3944
R8702 gnd.n3714 gnd.n3384 19.3944
R8703 gnd.n3714 gnd.n3713 19.3944
R8704 gnd.n3713 gnd.n3358 19.3944
R8705 gnd.n3738 gnd.n3358 19.3944
R8706 gnd.n3738 gnd.n3356 19.3944
R8707 gnd.n3742 gnd.n3356 19.3944
R8708 gnd.n3742 gnd.n3336 19.3944
R8709 gnd.n3769 gnd.n3336 19.3944
R8710 gnd.n3769 gnd.n3334 19.3944
R8711 gnd.n3779 gnd.n3334 19.3944
R8712 gnd.n3779 gnd.n3778 19.3944
R8713 gnd.n3778 gnd.n3777 19.3944
R8714 gnd.n3777 gnd.n3283 19.3944
R8715 gnd.n3827 gnd.n3283 19.3944
R8716 gnd.n3827 gnd.n3826 19.3944
R8717 gnd.n3826 gnd.n3825 19.3944
R8718 gnd.n3825 gnd.n3287 19.3944
R8719 gnd.n3307 gnd.n3287 19.3944
R8720 gnd.n3307 gnd.n3193 19.3944
R8721 gnd.n3864 gnd.n3193 19.3944
R8722 gnd.n3864 gnd.n3191 19.3944
R8723 gnd.n3870 gnd.n3191 19.3944
R8724 gnd.n3870 gnd.n3869 19.3944
R8725 gnd.n3869 gnd.n3166 19.3944
R8726 gnd.n3904 gnd.n3166 19.3944
R8727 gnd.n3904 gnd.n3164 19.3944
R8728 gnd.n3910 gnd.n3164 19.3944
R8729 gnd.n3910 gnd.n3909 19.3944
R8730 gnd.n3909 gnd.n3139 19.3944
R8731 gnd.n3949 gnd.n3139 19.3944
R8732 gnd.n3949 gnd.n3137 19.3944
R8733 gnd.n3955 gnd.n3137 19.3944
R8734 gnd.n3955 gnd.n3954 19.3944
R8735 gnd.n3954 gnd.n3111 19.3944
R8736 gnd.n3989 gnd.n3111 19.3944
R8737 gnd.n3989 gnd.n3109 19.3944
R8738 gnd.n3995 gnd.n3109 19.3944
R8739 gnd.n3995 gnd.n3994 19.3944
R8740 gnd.n3994 gnd.n3084 19.3944
R8741 gnd.n4038 gnd.n3084 19.3944
R8742 gnd.n4038 gnd.n3082 19.3944
R8743 gnd.n4044 gnd.n3082 19.3944
R8744 gnd.n4044 gnd.n4043 19.3944
R8745 gnd.n4043 gnd.n1651 19.3944
R8746 gnd.n4332 gnd.n1651 19.3944
R8747 gnd.n4332 gnd.n1649 19.3944
R8748 gnd.n4340 gnd.n1649 19.3944
R8749 gnd.n4340 gnd.n4339 19.3944
R8750 gnd.n4339 gnd.n4338 19.3944
R8751 gnd.n4441 gnd.n4440 19.3944
R8752 gnd.n4440 gnd.n1590 19.3944
R8753 gnd.n4436 gnd.n1590 19.3944
R8754 gnd.n4436 gnd.n4433 19.3944
R8755 gnd.n4433 gnd.n4430 19.3944
R8756 gnd.n4430 gnd.n4429 19.3944
R8757 gnd.n4429 gnd.n4426 19.3944
R8758 gnd.n4426 gnd.n4425 19.3944
R8759 gnd.n4425 gnd.n4422 19.3944
R8760 gnd.n4422 gnd.n4421 19.3944
R8761 gnd.n4421 gnd.n4418 19.3944
R8762 gnd.n4418 gnd.n4417 19.3944
R8763 gnd.n4417 gnd.n4414 19.3944
R8764 gnd.n4414 gnd.n4413 19.3944
R8765 gnd.n3598 gnd.n3497 19.3944
R8766 gnd.n3598 gnd.n3488 19.3944
R8767 gnd.n3611 gnd.n3488 19.3944
R8768 gnd.n3611 gnd.n3486 19.3944
R8769 gnd.n3615 gnd.n3486 19.3944
R8770 gnd.n3615 gnd.n3476 19.3944
R8771 gnd.n3627 gnd.n3476 19.3944
R8772 gnd.n3627 gnd.n3474 19.3944
R8773 gnd.n3661 gnd.n3474 19.3944
R8774 gnd.n3661 gnd.n3660 19.3944
R8775 gnd.n3660 gnd.n3659 19.3944
R8776 gnd.n3659 gnd.n3658 19.3944
R8777 gnd.n3658 gnd.n3655 19.3944
R8778 gnd.n3655 gnd.n3654 19.3944
R8779 gnd.n3654 gnd.n3653 19.3944
R8780 gnd.n3653 gnd.n3651 19.3944
R8781 gnd.n3651 gnd.n3650 19.3944
R8782 gnd.n3650 gnd.n3647 19.3944
R8783 gnd.n3647 gnd.n3646 19.3944
R8784 gnd.n3646 gnd.n3645 19.3944
R8785 gnd.n3645 gnd.n3643 19.3944
R8786 gnd.n3643 gnd.n3342 19.3944
R8787 gnd.n3758 gnd.n3342 19.3944
R8788 gnd.n3758 gnd.n3340 19.3944
R8789 gnd.n3764 gnd.n3340 19.3944
R8790 gnd.n3764 gnd.n3763 19.3944
R8791 gnd.n3763 gnd.n3264 19.3944
R8792 gnd.n3838 gnd.n3264 19.3944
R8793 gnd.n3838 gnd.n3265 19.3944
R8794 gnd.n3312 gnd.n3311 19.3944
R8795 gnd.n3315 gnd.n3314 19.3944
R8796 gnd.n3302 gnd.n3301 19.3944
R8797 gnd.n3857 gnd.n3198 19.3944
R8798 gnd.n3857 gnd.n3856 19.3944
R8799 gnd.n3856 gnd.n3855 19.3944
R8800 gnd.n3855 gnd.n3853 19.3944
R8801 gnd.n3853 gnd.n3852 19.3944
R8802 gnd.n3852 gnd.n3850 19.3944
R8803 gnd.n3850 gnd.n3849 19.3944
R8804 gnd.n3849 gnd.n3147 19.3944
R8805 gnd.n3925 gnd.n3147 19.3944
R8806 gnd.n3925 gnd.n3145 19.3944
R8807 gnd.n3944 gnd.n3145 19.3944
R8808 gnd.n3944 gnd.n3943 19.3944
R8809 gnd.n3943 gnd.n3942 19.3944
R8810 gnd.n3942 gnd.n3940 19.3944
R8811 gnd.n3940 gnd.n3939 19.3944
R8812 gnd.n3939 gnd.n3937 19.3944
R8813 gnd.n3937 gnd.n3936 19.3944
R8814 gnd.n3936 gnd.n3091 19.3944
R8815 gnd.n4010 gnd.n3091 19.3944
R8816 gnd.n4010 gnd.n3089 19.3944
R8817 gnd.n4033 gnd.n3089 19.3944
R8818 gnd.n4033 gnd.n4032 19.3944
R8819 gnd.n4032 gnd.n4031 19.3944
R8820 gnd.n4031 gnd.n4028 19.3944
R8821 gnd.n4028 gnd.n4027 19.3944
R8822 gnd.n4027 gnd.n4025 19.3944
R8823 gnd.n4025 gnd.n4024 19.3944
R8824 gnd.n4024 gnd.n4022 19.3944
R8825 gnd.n4022 gnd.n1637 19.3944
R8826 gnd.n3603 gnd.n3493 19.3944
R8827 gnd.n3603 gnd.n3491 19.3944
R8828 gnd.n3607 gnd.n3491 19.3944
R8829 gnd.n3607 gnd.n3482 19.3944
R8830 gnd.n3619 gnd.n3482 19.3944
R8831 gnd.n3619 gnd.n3480 19.3944
R8832 gnd.n3623 gnd.n3480 19.3944
R8833 gnd.n3623 gnd.n3469 19.3944
R8834 gnd.n3665 gnd.n3469 19.3944
R8835 gnd.n3665 gnd.n3423 19.3944
R8836 gnd.n3671 gnd.n3423 19.3944
R8837 gnd.n3671 gnd.n3670 19.3944
R8838 gnd.n3670 gnd.n3401 19.3944
R8839 gnd.n3692 gnd.n3401 19.3944
R8840 gnd.n3692 gnd.n3394 19.3944
R8841 gnd.n3703 gnd.n3394 19.3944
R8842 gnd.n3703 gnd.n3702 19.3944
R8843 gnd.n3702 gnd.n3375 19.3944
R8844 gnd.n3723 gnd.n3375 19.3944
R8845 gnd.n3723 gnd.n3365 19.3944
R8846 gnd.n3733 gnd.n3365 19.3944
R8847 gnd.n3733 gnd.n3348 19.3944
R8848 gnd.n3754 gnd.n3348 19.3944
R8849 gnd.n3754 gnd.n3753 19.3944
R8850 gnd.n3753 gnd.n3327 19.3944
R8851 gnd.n3784 gnd.n3327 19.3944
R8852 gnd.n3784 gnd.n3272 19.3944
R8853 gnd.n3834 gnd.n3272 19.3944
R8854 gnd.n3834 gnd.n3833 19.3944
R8855 gnd.n3833 gnd.n3832 19.3944
R8856 gnd.n3832 gnd.n3276 19.3944
R8857 gnd.n3294 gnd.n3276 19.3944
R8858 gnd.n3820 gnd.n3294 19.3944
R8859 gnd.n3820 gnd.n3819 19.3944
R8860 gnd.n3819 gnd.n3818 19.3944
R8861 gnd.n3818 gnd.n3298 19.3944
R8862 gnd.n3298 gnd.n3185 19.3944
R8863 gnd.n3875 gnd.n3185 19.3944
R8864 gnd.n3875 gnd.n3178 19.3944
R8865 gnd.n3886 gnd.n3178 19.3944
R8866 gnd.n3886 gnd.n3174 19.3944
R8867 gnd.n3899 gnd.n3174 19.3944
R8868 gnd.n3899 gnd.n3898 19.3944
R8869 gnd.n3898 gnd.n3153 19.3944
R8870 gnd.n3921 gnd.n3153 19.3944
R8871 gnd.n3921 gnd.n3920 19.3944
R8872 gnd.n3920 gnd.n3130 19.3944
R8873 gnd.n3960 gnd.n3130 19.3944
R8874 gnd.n3960 gnd.n3123 19.3944
R8875 gnd.n3971 gnd.n3123 19.3944
R8876 gnd.n3971 gnd.n3119 19.3944
R8877 gnd.n3984 gnd.n3119 19.3944
R8878 gnd.n3984 gnd.n3983 19.3944
R8879 gnd.n3983 gnd.n3098 19.3944
R8880 gnd.n4006 gnd.n3098 19.3944
R8881 gnd.n4006 gnd.n4005 19.3944
R8882 gnd.n4005 gnd.n3076 19.3944
R8883 gnd.n4049 gnd.n3076 19.3944
R8884 gnd.n4049 gnd.n3069 19.3944
R8885 gnd.n4060 gnd.n3069 19.3944
R8886 gnd.n4060 gnd.n3065 19.3944
R8887 gnd.n4327 gnd.n3065 19.3944
R8888 gnd.n4327 gnd.n4326 19.3944
R8889 gnd.n4326 gnd.n1640 19.3944
R8890 gnd.n4350 gnd.n1640 19.3944
R8891 gnd.n7174 gnd.n582 19.3944
R8892 gnd.n7170 gnd.n582 19.3944
R8893 gnd.n7170 gnd.n7169 19.3944
R8894 gnd.n7169 gnd.n7168 19.3944
R8895 gnd.n7168 gnd.n587 19.3944
R8896 gnd.n7164 gnd.n587 19.3944
R8897 gnd.n7164 gnd.n7163 19.3944
R8898 gnd.n7163 gnd.n7162 19.3944
R8899 gnd.n7162 gnd.n591 19.3944
R8900 gnd.n7158 gnd.n591 19.3944
R8901 gnd.n7158 gnd.n7157 19.3944
R8902 gnd.n7157 gnd.n7156 19.3944
R8903 gnd.n7156 gnd.n7153 19.3944
R8904 gnd.n7153 gnd.n428 19.3944
R8905 gnd.n7327 gnd.n428 19.3944
R8906 gnd.n7327 gnd.n425 19.3944
R8907 gnd.n7339 gnd.n425 19.3944
R8908 gnd.n7339 gnd.n426 19.3944
R8909 gnd.n7335 gnd.n426 19.3944
R8910 gnd.n7335 gnd.n7334 19.3944
R8911 gnd.n7334 gnd.n388 19.3944
R8912 gnd.n7417 gnd.n388 19.3944
R8913 gnd.n7418 gnd.n7417 19.3944
R8914 gnd.n7418 gnd.n385 19.3944
R8915 gnd.n7423 gnd.n385 19.3944
R8916 gnd.n7423 gnd.n386 19.3944
R8917 gnd.n386 gnd.n354 19.3944
R8918 gnd.n7541 gnd.n354 19.3944
R8919 gnd.n7541 gnd.n352 19.3944
R8920 gnd.n7545 gnd.n352 19.3944
R8921 gnd.n7546 gnd.n7545 19.3944
R8922 gnd.n7546 gnd.n80 19.3944
R8923 gnd.n7888 gnd.n80 19.3944
R8924 gnd.n7888 gnd.n7887 19.3944
R8925 gnd.n7887 gnd.n7886 19.3944
R8926 gnd.n7886 gnd.n85 19.3944
R8927 gnd.n7882 gnd.n85 19.3944
R8928 gnd.n7882 gnd.n7881 19.3944
R8929 gnd.n7881 gnd.n7880 19.3944
R8930 gnd.n7880 gnd.n90 19.3944
R8931 gnd.n7876 gnd.n90 19.3944
R8932 gnd.n7876 gnd.n7875 19.3944
R8933 gnd.n7875 gnd.n7874 19.3944
R8934 gnd.n7874 gnd.n95 19.3944
R8935 gnd.n7870 gnd.n95 19.3944
R8936 gnd.n7870 gnd.n7869 19.3944
R8937 gnd.n7869 gnd.n7868 19.3944
R8938 gnd.n7868 gnd.n100 19.3944
R8939 gnd.n7864 gnd.n100 19.3944
R8940 gnd.n7864 gnd.n7863 19.3944
R8941 gnd.n7863 gnd.n7862 19.3944
R8942 gnd.n7862 gnd.n105 19.3944
R8943 gnd.n7858 gnd.n105 19.3944
R8944 gnd.n7858 gnd.n7857 19.3944
R8945 gnd.n7857 gnd.n7856 19.3944
R8946 gnd.n7856 gnd.n110 19.3944
R8947 gnd.n7852 gnd.n110 19.3944
R8948 gnd.n7852 gnd.n7851 19.3944
R8949 gnd.n7851 gnd.n7850 19.3944
R8950 gnd.n7850 gnd.n115 19.3944
R8951 gnd.n7846 gnd.n115 19.3944
R8952 gnd.n7846 gnd.n7845 19.3944
R8953 gnd.n7845 gnd.n7844 19.3944
R8954 gnd.n7844 gnd.n120 19.3944
R8955 gnd.n7738 gnd.n7737 19.3944
R8956 gnd.n7737 gnd.n7736 19.3944
R8957 gnd.n7736 gnd.n7685 19.3944
R8958 gnd.n7732 gnd.n7685 19.3944
R8959 gnd.n7732 gnd.n7731 19.3944
R8960 gnd.n7731 gnd.n7730 19.3944
R8961 gnd.n7730 gnd.n7693 19.3944
R8962 gnd.n7726 gnd.n7693 19.3944
R8963 gnd.n7726 gnd.n7725 19.3944
R8964 gnd.n7725 gnd.n7724 19.3944
R8965 gnd.n7724 gnd.n7701 19.3944
R8966 gnd.n7720 gnd.n7701 19.3944
R8967 gnd.n7720 gnd.n7719 19.3944
R8968 gnd.n7719 gnd.n7718 19.3944
R8969 gnd.n7718 gnd.n7709 19.3944
R8970 gnd.n7714 gnd.n7709 19.3944
R8971 gnd.n7255 gnd.n502 19.3944
R8972 gnd.n6728 gnd.n502 19.3944
R8973 gnd.n6728 gnd.n6727 19.3944
R8974 gnd.n6727 gnd.n6602 19.3944
R8975 gnd.n6720 gnd.n6602 19.3944
R8976 gnd.n6720 gnd.n6719 19.3944
R8977 gnd.n6719 gnd.n6612 19.3944
R8978 gnd.n6712 gnd.n6612 19.3944
R8979 gnd.n6712 gnd.n6711 19.3944
R8980 gnd.n6711 gnd.n6622 19.3944
R8981 gnd.n6704 gnd.n6622 19.3944
R8982 gnd.n6704 gnd.n6703 19.3944
R8983 gnd.n6703 gnd.n6632 19.3944
R8984 gnd.n6696 gnd.n6632 19.3944
R8985 gnd.n6696 gnd.n6695 19.3944
R8986 gnd.n6695 gnd.n6642 19.3944
R8987 gnd.n7259 gnd.n500 19.3944
R8988 gnd.n7259 gnd.n484 19.3944
R8989 gnd.n7271 gnd.n484 19.3944
R8990 gnd.n7271 gnd.n482 19.3944
R8991 gnd.n7275 gnd.n482 19.3944
R8992 gnd.n7275 gnd.n466 19.3944
R8993 gnd.n7287 gnd.n466 19.3944
R8994 gnd.n7287 gnd.n464 19.3944
R8995 gnd.n7291 gnd.n464 19.3944
R8996 gnd.n7291 gnd.n449 19.3944
R8997 gnd.n7303 gnd.n449 19.3944
R8998 gnd.n7303 gnd.n446 19.3944
R8999 gnd.n7313 gnd.n446 19.3944
R9000 gnd.n7313 gnd.n447 19.3944
R9001 gnd.n7309 gnd.n447 19.3944
R9002 gnd.n7309 gnd.n7308 19.3944
R9003 gnd.n7308 gnd.n411 19.3944
R9004 gnd.n7389 gnd.n411 19.3944
R9005 gnd.n7389 gnd.n412 19.3944
R9006 gnd.n7385 gnd.n412 19.3944
R9007 gnd.n7385 gnd.n7384 19.3944
R9008 gnd.n7384 gnd.n379 19.3944
R9009 gnd.n7436 gnd.n379 19.3944
R9010 gnd.n7436 gnd.n380 19.3944
R9011 gnd.n7432 gnd.n380 19.3944
R9012 gnd.n7432 gnd.n7431 19.3944
R9013 gnd.n7431 gnd.n7430 19.3944
R9014 gnd.n7430 gnd.n317 19.3944
R9015 gnd.n7582 gnd.n317 19.3944
R9016 gnd.n7582 gnd.n318 19.3944
R9017 gnd.n7578 gnd.n318 19.3944
R9018 gnd.n7578 gnd.n7577 19.3944
R9019 gnd.n7577 gnd.n7576 19.3944
R9020 gnd.n7576 gnd.n324 19.3944
R9021 gnd.n7572 gnd.n324 19.3944
R9022 gnd.n7572 gnd.n7571 19.3944
R9023 gnd.n7571 gnd.n296 19.3944
R9024 gnd.n7595 gnd.n296 19.3944
R9025 gnd.n7595 gnd.n294 19.3944
R9026 gnd.n7599 gnd.n294 19.3944
R9027 gnd.n7599 gnd.n280 19.3944
R9028 gnd.n7611 gnd.n280 19.3944
R9029 gnd.n7611 gnd.n278 19.3944
R9030 gnd.n7615 gnd.n278 19.3944
R9031 gnd.n7615 gnd.n266 19.3944
R9032 gnd.n7627 gnd.n266 19.3944
R9033 gnd.n7627 gnd.n264 19.3944
R9034 gnd.n7631 gnd.n264 19.3944
R9035 gnd.n7631 gnd.n250 19.3944
R9036 gnd.n7643 gnd.n250 19.3944
R9037 gnd.n7643 gnd.n248 19.3944
R9038 gnd.n7647 gnd.n248 19.3944
R9039 gnd.n7647 gnd.n236 19.3944
R9040 gnd.n7659 gnd.n236 19.3944
R9041 gnd.n7659 gnd.n234 19.3944
R9042 gnd.n7663 gnd.n234 19.3944
R9043 gnd.n7663 gnd.n221 19.3944
R9044 gnd.n7675 gnd.n221 19.3944
R9045 gnd.n7675 gnd.n218 19.3944
R9046 gnd.n7747 gnd.n218 19.3944
R9047 gnd.n7747 gnd.n219 19.3944
R9048 gnd.n7743 gnd.n219 19.3944
R9049 gnd.n7743 gnd.n7742 19.3944
R9050 gnd.n7742 gnd.n7741 19.3944
R9051 gnd.n5355 gnd.n5350 19.3944
R9052 gnd.n5355 gnd.n1123 19.3944
R9053 gnd.n5784 gnd.n1123 19.3944
R9054 gnd.n5784 gnd.n5783 19.3944
R9055 gnd.n5783 gnd.n1126 19.3944
R9056 gnd.n5776 gnd.n1126 19.3944
R9057 gnd.n5776 gnd.n5775 19.3944
R9058 gnd.n5775 gnd.n1135 19.3944
R9059 gnd.n5768 gnd.n1135 19.3944
R9060 gnd.n5768 gnd.n5767 19.3944
R9061 gnd.n5767 gnd.n1143 19.3944
R9062 gnd.n5760 gnd.n1143 19.3944
R9063 gnd.n5760 gnd.n5759 19.3944
R9064 gnd.n5759 gnd.n1153 19.3944
R9065 gnd.n5752 gnd.n1153 19.3944
R9066 gnd.n5752 gnd.n5751 19.3944
R9067 gnd.n3054 gnd.n1415 19.3944
R9068 gnd.n5224 gnd.n1415 19.3944
R9069 gnd.n5224 gnd.n5223 19.3944
R9070 gnd.n5223 gnd.n5222 19.3944
R9071 gnd.n5222 gnd.n1419 19.3944
R9072 gnd.n4966 gnd.n1419 19.3944
R9073 gnd.n4966 gnd.n4963 19.3944
R9074 gnd.n4990 gnd.n4963 19.3944
R9075 gnd.n4990 gnd.n4989 19.3944
R9076 gnd.n4989 gnd.n4988 19.3944
R9077 gnd.n4988 gnd.n4972 19.3944
R9078 gnd.n4984 gnd.n4972 19.3944
R9079 gnd.n4984 gnd.n4983 19.3944
R9080 gnd.n4983 gnd.n4982 19.3944
R9081 gnd.n4982 gnd.n4980 19.3944
R9082 gnd.n4980 gnd.n4954 19.3944
R9083 gnd.n4954 gnd.n4952 19.3944
R9084 gnd.n5038 gnd.n4952 19.3944
R9085 gnd.n5038 gnd.n4950 19.3944
R9086 gnd.n5042 gnd.n4950 19.3944
R9087 gnd.n5042 gnd.n4948 19.3944
R9088 gnd.n5046 gnd.n4948 19.3944
R9089 gnd.n5046 gnd.n4946 19.3944
R9090 gnd.n5094 gnd.n4946 19.3944
R9091 gnd.n5094 gnd.n5093 19.3944
R9092 gnd.n5093 gnd.n5092 19.3944
R9093 gnd.n5092 gnd.n5052 19.3944
R9094 gnd.n5088 gnd.n5052 19.3944
R9095 gnd.n5088 gnd.n5087 19.3944
R9096 gnd.n5087 gnd.n5086 19.3944
R9097 gnd.n5086 gnd.n5058 19.3944
R9098 gnd.n5082 gnd.n5058 19.3944
R9099 gnd.n5082 gnd.n5081 19.3944
R9100 gnd.n5081 gnd.n5080 19.3944
R9101 gnd.n5080 gnd.n5064 19.3944
R9102 gnd.n5073 gnd.n5064 19.3944
R9103 gnd.n5073 gnd.n5072 19.3944
R9104 gnd.n5072 gnd.n5071 19.3944
R9105 gnd.n5071 gnd.n1095 19.3944
R9106 gnd.n5802 gnd.n1095 19.3944
R9107 gnd.n5802 gnd.n1093 19.3944
R9108 gnd.n5806 gnd.n1093 19.3944
R9109 gnd.n5806 gnd.n1082 19.3944
R9110 gnd.n5818 gnd.n1082 19.3944
R9111 gnd.n5818 gnd.n1080 19.3944
R9112 gnd.n5822 gnd.n1080 19.3944
R9113 gnd.n5822 gnd.n1068 19.3944
R9114 gnd.n5834 gnd.n1068 19.3944
R9115 gnd.n5834 gnd.n1066 19.3944
R9116 gnd.n5838 gnd.n1066 19.3944
R9117 gnd.n5838 gnd.n1054 19.3944
R9118 gnd.n5850 gnd.n1054 19.3944
R9119 gnd.n5850 gnd.n1052 19.3944
R9120 gnd.n5854 gnd.n1052 19.3944
R9121 gnd.n5854 gnd.n1039 19.3944
R9122 gnd.n5866 gnd.n1039 19.3944
R9123 gnd.n5866 gnd.n1037 19.3944
R9124 gnd.n5870 gnd.n1037 19.3944
R9125 gnd.n5870 gnd.n1025 19.3944
R9126 gnd.n5882 gnd.n1025 19.3944
R9127 gnd.n5882 gnd.n1023 19.3944
R9128 gnd.n5888 gnd.n1023 19.3944
R9129 gnd.n5888 gnd.n5887 19.3944
R9130 gnd.n5887 gnd.n985 19.3944
R9131 gnd.n5980 gnd.n985 19.3944
R9132 gnd.n5980 gnd.n983 19.3944
R9133 gnd.n5984 gnd.n983 19.3944
R9134 gnd.n5984 gnd.n969 19.3944
R9135 gnd.n5996 gnd.n969 19.3944
R9136 gnd.n5996 gnd.n967 19.3944
R9137 gnd.n6000 gnd.n967 19.3944
R9138 gnd.n6000 gnd.n951 19.3944
R9139 gnd.n6015 gnd.n951 19.3944
R9140 gnd.n6015 gnd.n949 19.3944
R9141 gnd.n6019 gnd.n949 19.3944
R9142 gnd.n6019 gnd.n915 19.3944
R9143 gnd.n6071 gnd.n915 19.3944
R9144 gnd.n6071 gnd.n913 19.3944
R9145 gnd.n6077 gnd.n913 19.3944
R9146 gnd.n6077 gnd.n6076 19.3944
R9147 gnd.n6076 gnd.n881 19.3944
R9148 gnd.n6835 gnd.n881 19.3944
R9149 gnd.n6835 gnd.n879 19.3944
R9150 gnd.n6839 gnd.n879 19.3944
R9151 gnd.n6839 gnd.n866 19.3944
R9152 gnd.n6851 gnd.n866 19.3944
R9153 gnd.n6851 gnd.n864 19.3944
R9154 gnd.n6855 gnd.n864 19.3944
R9155 gnd.n6855 gnd.n850 19.3944
R9156 gnd.n6867 gnd.n850 19.3944
R9157 gnd.n6867 gnd.n848 19.3944
R9158 gnd.n6871 gnd.n848 19.3944
R9159 gnd.n6871 gnd.n834 19.3944
R9160 gnd.n6883 gnd.n834 19.3944
R9161 gnd.n6883 gnd.n832 19.3944
R9162 gnd.n6887 gnd.n832 19.3944
R9163 gnd.n6887 gnd.n818 19.3944
R9164 gnd.n6899 gnd.n818 19.3944
R9165 gnd.n6899 gnd.n816 19.3944
R9166 gnd.n6903 gnd.n816 19.3944
R9167 gnd.n6903 gnd.n803 19.3944
R9168 gnd.n6915 gnd.n803 19.3944
R9169 gnd.n6915 gnd.n801 19.3944
R9170 gnd.n6919 gnd.n801 19.3944
R9171 gnd.n6919 gnd.n787 19.3944
R9172 gnd.n6931 gnd.n787 19.3944
R9173 gnd.n6931 gnd.n785 19.3944
R9174 gnd.n6935 gnd.n785 19.3944
R9175 gnd.n6935 gnd.n771 19.3944
R9176 gnd.n6947 gnd.n771 19.3944
R9177 gnd.n6947 gnd.n769 19.3944
R9178 gnd.n6951 gnd.n769 19.3944
R9179 gnd.n6951 gnd.n755 19.3944
R9180 gnd.n6963 gnd.n755 19.3944
R9181 gnd.n6963 gnd.n753 19.3944
R9182 gnd.n6967 gnd.n753 19.3944
R9183 gnd.n6967 gnd.n739 19.3944
R9184 gnd.n6979 gnd.n739 19.3944
R9185 gnd.n6979 gnd.n737 19.3944
R9186 gnd.n6983 gnd.n737 19.3944
R9187 gnd.n6983 gnd.n724 19.3944
R9188 gnd.n6995 gnd.n724 19.3944
R9189 gnd.n6995 gnd.n722 19.3944
R9190 gnd.n6999 gnd.n722 19.3944
R9191 gnd.n6999 gnd.n710 19.3944
R9192 gnd.n7011 gnd.n710 19.3944
R9193 gnd.n7011 gnd.n708 19.3944
R9194 gnd.n7015 gnd.n708 19.3944
R9195 gnd.n7015 gnd.n696 19.3944
R9196 gnd.n7027 gnd.n696 19.3944
R9197 gnd.n7027 gnd.n694 19.3944
R9198 gnd.n7031 gnd.n694 19.3944
R9199 gnd.n7031 gnd.n682 19.3944
R9200 gnd.n7043 gnd.n682 19.3944
R9201 gnd.n7043 gnd.n680 19.3944
R9202 gnd.n7047 gnd.n680 19.3944
R9203 gnd.n7047 gnd.n667 19.3944
R9204 gnd.n7060 gnd.n667 19.3944
R9205 gnd.n7060 gnd.n665 19.3944
R9206 gnd.n7066 gnd.n665 19.3944
R9207 gnd.n7066 gnd.n7065 19.3944
R9208 gnd.n7065 gnd.n637 19.3944
R9209 gnd.n7080 gnd.n637 19.3944
R9210 gnd.n7080 gnd.n635 19.3944
R9211 gnd.n7084 gnd.n635 19.3944
R9212 gnd.n7084 gnd.n633 19.3944
R9213 gnd.n7088 gnd.n633 19.3944
R9214 gnd.n7088 gnd.n631 19.3944
R9215 gnd.n7092 gnd.n631 19.3944
R9216 gnd.n7092 gnd.n629 19.3944
R9217 gnd.n7096 gnd.n629 19.3944
R9218 gnd.n7096 gnd.n627 19.3944
R9219 gnd.n7100 gnd.n627 19.3944
R9220 gnd.n7100 gnd.n625 19.3944
R9221 gnd.n7104 gnd.n625 19.3944
R9222 gnd.n7104 gnd.n623 19.3944
R9223 gnd.n7125 gnd.n623 19.3944
R9224 gnd.n7125 gnd.n7124 19.3944
R9225 gnd.n7124 gnd.n7123 19.3944
R9226 gnd.n7123 gnd.n7110 19.3944
R9227 gnd.n7119 gnd.n7110 19.3944
R9228 gnd.n7119 gnd.n7118 19.3944
R9229 gnd.n7118 gnd.n7117 19.3944
R9230 gnd.n7117 gnd.n421 19.3944
R9231 gnd.n421 gnd.n419 19.3944
R9232 gnd.n7346 gnd.n419 19.3944
R9233 gnd.n7346 gnd.n417 19.3944
R9234 gnd.n7379 gnd.n417 19.3944
R9235 gnd.n7379 gnd.n7378 19.3944
R9236 gnd.n7378 gnd.n7377 19.3944
R9237 gnd.n7377 gnd.n7352 19.3944
R9238 gnd.n7373 gnd.n7352 19.3944
R9239 gnd.n7373 gnd.n7372 19.3944
R9240 gnd.n7372 gnd.n7371 19.3944
R9241 gnd.n7371 gnd.n7358 19.3944
R9242 gnd.n7367 gnd.n7358 19.3944
R9243 gnd.n7367 gnd.n7366 19.3944
R9244 gnd.n7366 gnd.n7365 19.3944
R9245 gnd.n7365 gnd.n341 19.3944
R9246 gnd.n7558 gnd.n341 19.3944
R9247 gnd.n7559 gnd.n7558 19.3944
R9248 gnd.n2475 gnd.n2145 19.3944
R9249 gnd.n2469 gnd.n2145 19.3944
R9250 gnd.n2469 gnd.n2468 19.3944
R9251 gnd.n2468 gnd.n2467 19.3944
R9252 gnd.n2467 gnd.n2152 19.3944
R9253 gnd.n2461 gnd.n2152 19.3944
R9254 gnd.n2461 gnd.n2460 19.3944
R9255 gnd.n2460 gnd.n2459 19.3944
R9256 gnd.n2459 gnd.n2160 19.3944
R9257 gnd.n2453 gnd.n2160 19.3944
R9258 gnd.n2453 gnd.n2452 19.3944
R9259 gnd.n2452 gnd.n2451 19.3944
R9260 gnd.n2451 gnd.n2168 19.3944
R9261 gnd.n2445 gnd.n2168 19.3944
R9262 gnd.n2445 gnd.n2444 19.3944
R9263 gnd.n2444 gnd.n2443 19.3944
R9264 gnd.n2443 gnd.n2176 19.3944
R9265 gnd.n2437 gnd.n2176 19.3944
R9266 gnd.n2437 gnd.n2436 19.3944
R9267 gnd.n2436 gnd.n2435 19.3944
R9268 gnd.n2435 gnd.n2184 19.3944
R9269 gnd.n2429 gnd.n2184 19.3944
R9270 gnd.n2429 gnd.n2428 19.3944
R9271 gnd.n2428 gnd.n2427 19.3944
R9272 gnd.n2427 gnd.n2192 19.3944
R9273 gnd.n2421 gnd.n2192 19.3944
R9274 gnd.n2421 gnd.n2420 19.3944
R9275 gnd.n2420 gnd.n2419 19.3944
R9276 gnd.n2419 gnd.n2200 19.3944
R9277 gnd.n2413 gnd.n2200 19.3944
R9278 gnd.n2413 gnd.n2412 19.3944
R9279 gnd.n2412 gnd.n2411 19.3944
R9280 gnd.n2411 gnd.n2208 19.3944
R9281 gnd.n2405 gnd.n2208 19.3944
R9282 gnd.n2405 gnd.n2404 19.3944
R9283 gnd.n2404 gnd.n2403 19.3944
R9284 gnd.n2403 gnd.n2216 19.3944
R9285 gnd.n2397 gnd.n2216 19.3944
R9286 gnd.n2397 gnd.n2396 19.3944
R9287 gnd.n2396 gnd.n2395 19.3944
R9288 gnd.n2395 gnd.n2224 19.3944
R9289 gnd.n2389 gnd.n2224 19.3944
R9290 gnd.n2389 gnd.n2388 19.3944
R9291 gnd.n2388 gnd.n2387 19.3944
R9292 gnd.n2387 gnd.n2232 19.3944
R9293 gnd.n2381 gnd.n2232 19.3944
R9294 gnd.n2381 gnd.n2380 19.3944
R9295 gnd.n2380 gnd.n2379 19.3944
R9296 gnd.n2379 gnd.n2240 19.3944
R9297 gnd.n2373 gnd.n2240 19.3944
R9298 gnd.n2373 gnd.n2372 19.3944
R9299 gnd.n2372 gnd.n2371 19.3944
R9300 gnd.n2371 gnd.n2248 19.3944
R9301 gnd.n2365 gnd.n2248 19.3944
R9302 gnd.n2365 gnd.n2364 19.3944
R9303 gnd.n2364 gnd.n2363 19.3944
R9304 gnd.n2363 gnd.n2256 19.3944
R9305 gnd.n2357 gnd.n2256 19.3944
R9306 gnd.n2357 gnd.n2356 19.3944
R9307 gnd.n2356 gnd.n2355 19.3944
R9308 gnd.n2355 gnd.n2264 19.3944
R9309 gnd.n2349 gnd.n2264 19.3944
R9310 gnd.n2349 gnd.n2348 19.3944
R9311 gnd.n2348 gnd.n2347 19.3944
R9312 gnd.n2347 gnd.n2272 19.3944
R9313 gnd.n2341 gnd.n2272 19.3944
R9314 gnd.n2341 gnd.n2340 19.3944
R9315 gnd.n2340 gnd.n2339 19.3944
R9316 gnd.n2339 gnd.n2280 19.3944
R9317 gnd.n2333 gnd.n2280 19.3944
R9318 gnd.n2333 gnd.n2332 19.3944
R9319 gnd.n2332 gnd.n2331 19.3944
R9320 gnd.n2331 gnd.n2288 19.3944
R9321 gnd.n2325 gnd.n2288 19.3944
R9322 gnd.n2325 gnd.n2324 19.3944
R9323 gnd.n2324 gnd.n2323 19.3944
R9324 gnd.n2323 gnd.n2296 19.3944
R9325 gnd.n2317 gnd.n2296 19.3944
R9326 gnd.n2317 gnd.n2316 19.3944
R9327 gnd.n2316 gnd.n2315 19.3944
R9328 gnd.n2315 gnd.n2304 19.3944
R9329 gnd.n2309 gnd.n2304 19.3944
R9330 gnd.n2309 gnd.n337 19.3944
R9331 gnd.n7562 gnd.n337 19.3944
R9332 gnd.n2841 gnd.n1785 19.3944
R9333 gnd.n2837 gnd.n1785 19.3944
R9334 gnd.n2837 gnd.n1787 19.3944
R9335 gnd.n2831 gnd.n1787 19.3944
R9336 gnd.n2831 gnd.n2830 19.3944
R9337 gnd.n2830 gnd.n2829 19.3944
R9338 gnd.n2829 gnd.n1794 19.3944
R9339 gnd.n2823 gnd.n1794 19.3944
R9340 gnd.n2823 gnd.n2822 19.3944
R9341 gnd.n2822 gnd.n2821 19.3944
R9342 gnd.n2821 gnd.n1802 19.3944
R9343 gnd.n2815 gnd.n1802 19.3944
R9344 gnd.n2815 gnd.n2814 19.3944
R9345 gnd.n2814 gnd.n2813 19.3944
R9346 gnd.n2813 gnd.n1810 19.3944
R9347 gnd.n2807 gnd.n1810 19.3944
R9348 gnd.n2807 gnd.n2806 19.3944
R9349 gnd.n2806 gnd.n2805 19.3944
R9350 gnd.n2805 gnd.n1818 19.3944
R9351 gnd.n2799 gnd.n1818 19.3944
R9352 gnd.n2799 gnd.n2798 19.3944
R9353 gnd.n2798 gnd.n2797 19.3944
R9354 gnd.n2797 gnd.n1826 19.3944
R9355 gnd.n2791 gnd.n1826 19.3944
R9356 gnd.n2791 gnd.n2790 19.3944
R9357 gnd.n2790 gnd.n2789 19.3944
R9358 gnd.n2789 gnd.n1834 19.3944
R9359 gnd.n2783 gnd.n1834 19.3944
R9360 gnd.n2783 gnd.n2782 19.3944
R9361 gnd.n2782 gnd.n2781 19.3944
R9362 gnd.n2781 gnd.n1842 19.3944
R9363 gnd.n2775 gnd.n1842 19.3944
R9364 gnd.n2775 gnd.n2774 19.3944
R9365 gnd.n2774 gnd.n2773 19.3944
R9366 gnd.n2773 gnd.n1850 19.3944
R9367 gnd.n2767 gnd.n1850 19.3944
R9368 gnd.n2767 gnd.n2766 19.3944
R9369 gnd.n2766 gnd.n2765 19.3944
R9370 gnd.n2765 gnd.n1858 19.3944
R9371 gnd.n2759 gnd.n1858 19.3944
R9372 gnd.n2759 gnd.n2758 19.3944
R9373 gnd.n2758 gnd.n2757 19.3944
R9374 gnd.n2757 gnd.n1866 19.3944
R9375 gnd.n2751 gnd.n1866 19.3944
R9376 gnd.n2751 gnd.n2750 19.3944
R9377 gnd.n2750 gnd.n2749 19.3944
R9378 gnd.n2749 gnd.n1874 19.3944
R9379 gnd.n2743 gnd.n1874 19.3944
R9380 gnd.n2743 gnd.n2742 19.3944
R9381 gnd.n2742 gnd.n2741 19.3944
R9382 gnd.n2741 gnd.n1882 19.3944
R9383 gnd.n2735 gnd.n1882 19.3944
R9384 gnd.n2735 gnd.n2734 19.3944
R9385 gnd.n2734 gnd.n2733 19.3944
R9386 gnd.n2733 gnd.n1890 19.3944
R9387 gnd.n2727 gnd.n1890 19.3944
R9388 gnd.n2727 gnd.n2726 19.3944
R9389 gnd.n2726 gnd.n2725 19.3944
R9390 gnd.n2725 gnd.n1898 19.3944
R9391 gnd.n2719 gnd.n1898 19.3944
R9392 gnd.n2719 gnd.n2718 19.3944
R9393 gnd.n2718 gnd.n2717 19.3944
R9394 gnd.n2717 gnd.n1906 19.3944
R9395 gnd.n2711 gnd.n1906 19.3944
R9396 gnd.n2711 gnd.n2710 19.3944
R9397 gnd.n2710 gnd.n2709 19.3944
R9398 gnd.n2709 gnd.n1914 19.3944
R9399 gnd.n2703 gnd.n1914 19.3944
R9400 gnd.n2703 gnd.n2702 19.3944
R9401 gnd.n2702 gnd.n2701 19.3944
R9402 gnd.n2701 gnd.n1922 19.3944
R9403 gnd.n2695 gnd.n1922 19.3944
R9404 gnd.n2695 gnd.n2694 19.3944
R9405 gnd.n2694 gnd.n2693 19.3944
R9406 gnd.n2693 gnd.n1930 19.3944
R9407 gnd.n2687 gnd.n1930 19.3944
R9408 gnd.n2687 gnd.n2686 19.3944
R9409 gnd.n2686 gnd.n2685 19.3944
R9410 gnd.n2685 gnd.n1938 19.3944
R9411 gnd.n2679 gnd.n1938 19.3944
R9412 gnd.n2679 gnd.n2678 19.3944
R9413 gnd.n2678 gnd.n2677 19.3944
R9414 gnd.n2677 gnd.n1946 19.3944
R9415 gnd.n2671 gnd.n1946 19.3944
R9416 gnd.n2671 gnd.n2670 19.3944
R9417 gnd.n2670 gnd.n2669 19.3944
R9418 gnd.n2669 gnd.n1954 19.3944
R9419 gnd.n2663 gnd.n1954 19.3944
R9420 gnd.n2663 gnd.n2662 19.3944
R9421 gnd.n2662 gnd.n2661 19.3944
R9422 gnd.n2661 gnd.n1962 19.3944
R9423 gnd.n2655 gnd.n1962 19.3944
R9424 gnd.n2655 gnd.n2654 19.3944
R9425 gnd.n2654 gnd.n2653 19.3944
R9426 gnd.n2653 gnd.n1970 19.3944
R9427 gnd.n2647 gnd.n1970 19.3944
R9428 gnd.n2647 gnd.n2646 19.3944
R9429 gnd.n2646 gnd.n2645 19.3944
R9430 gnd.n2645 gnd.n1978 19.3944
R9431 gnd.n2639 gnd.n1978 19.3944
R9432 gnd.n2639 gnd.n2638 19.3944
R9433 gnd.n2638 gnd.n2637 19.3944
R9434 gnd.n2637 gnd.n1986 19.3944
R9435 gnd.n2631 gnd.n1986 19.3944
R9436 gnd.n2631 gnd.n2630 19.3944
R9437 gnd.n2630 gnd.n2629 19.3944
R9438 gnd.n2629 gnd.n1994 19.3944
R9439 gnd.n2623 gnd.n1994 19.3944
R9440 gnd.n2623 gnd.n2622 19.3944
R9441 gnd.n2622 gnd.n2621 19.3944
R9442 gnd.n2621 gnd.n2002 19.3944
R9443 gnd.n2615 gnd.n2002 19.3944
R9444 gnd.n2615 gnd.n2614 19.3944
R9445 gnd.n2614 gnd.n2613 19.3944
R9446 gnd.n2613 gnd.n2010 19.3944
R9447 gnd.n2607 gnd.n2010 19.3944
R9448 gnd.n2607 gnd.n2606 19.3944
R9449 gnd.n2606 gnd.n2605 19.3944
R9450 gnd.n2605 gnd.n2018 19.3944
R9451 gnd.n2599 gnd.n2018 19.3944
R9452 gnd.n2599 gnd.n2598 19.3944
R9453 gnd.n2598 gnd.n2597 19.3944
R9454 gnd.n2597 gnd.n2026 19.3944
R9455 gnd.n2591 gnd.n2026 19.3944
R9456 gnd.n2591 gnd.n2590 19.3944
R9457 gnd.n2590 gnd.n2589 19.3944
R9458 gnd.n2589 gnd.n2034 19.3944
R9459 gnd.n2583 gnd.n2034 19.3944
R9460 gnd.n2583 gnd.n2582 19.3944
R9461 gnd.n2582 gnd.n2581 19.3944
R9462 gnd.n2581 gnd.n2042 19.3944
R9463 gnd.n2575 gnd.n2042 19.3944
R9464 gnd.n2575 gnd.n2574 19.3944
R9465 gnd.n2574 gnd.n2573 19.3944
R9466 gnd.n2573 gnd.n2050 19.3944
R9467 gnd.n2567 gnd.n2050 19.3944
R9468 gnd.n2567 gnd.n2566 19.3944
R9469 gnd.n2566 gnd.n2565 19.3944
R9470 gnd.n2565 gnd.n2058 19.3944
R9471 gnd.n2559 gnd.n2058 19.3944
R9472 gnd.n2559 gnd.n2558 19.3944
R9473 gnd.n2558 gnd.n2557 19.3944
R9474 gnd.n2557 gnd.n2066 19.3944
R9475 gnd.n2551 gnd.n2066 19.3944
R9476 gnd.n2551 gnd.n2550 19.3944
R9477 gnd.n2550 gnd.n2549 19.3944
R9478 gnd.n2549 gnd.n2074 19.3944
R9479 gnd.n2543 gnd.n2074 19.3944
R9480 gnd.n2543 gnd.n2542 19.3944
R9481 gnd.n2542 gnd.n2541 19.3944
R9482 gnd.n2541 gnd.n2082 19.3944
R9483 gnd.n2535 gnd.n2082 19.3944
R9484 gnd.n2535 gnd.n2534 19.3944
R9485 gnd.n2534 gnd.n2533 19.3944
R9486 gnd.n2533 gnd.n2090 19.3944
R9487 gnd.n2527 gnd.n2090 19.3944
R9488 gnd.n2527 gnd.n2526 19.3944
R9489 gnd.n2526 gnd.n2525 19.3944
R9490 gnd.n2525 gnd.n2098 19.3944
R9491 gnd.n2519 gnd.n2098 19.3944
R9492 gnd.n2519 gnd.n2518 19.3944
R9493 gnd.n2518 gnd.n2517 19.3944
R9494 gnd.n2517 gnd.n2106 19.3944
R9495 gnd.n2511 gnd.n2106 19.3944
R9496 gnd.n2511 gnd.n2510 19.3944
R9497 gnd.n2510 gnd.n2509 19.3944
R9498 gnd.n2509 gnd.n2114 19.3944
R9499 gnd.n2503 gnd.n2114 19.3944
R9500 gnd.n2503 gnd.n2502 19.3944
R9501 gnd.n2502 gnd.n2501 19.3944
R9502 gnd.n2501 gnd.n2122 19.3944
R9503 gnd.n2495 gnd.n2122 19.3944
R9504 gnd.n2495 gnd.n2494 19.3944
R9505 gnd.n2494 gnd.n2493 19.3944
R9506 gnd.n2493 gnd.n2130 19.3944
R9507 gnd.n2487 gnd.n2130 19.3944
R9508 gnd.n2487 gnd.n2486 19.3944
R9509 gnd.n2486 gnd.n2485 19.3944
R9510 gnd.n2485 gnd.n2138 19.3944
R9511 gnd.n2479 gnd.n2138 19.3944
R9512 gnd.n2479 gnd.n2478 19.3944
R9513 gnd.n7249 gnd.n7248 19.3944
R9514 gnd.n7248 gnd.n7247 19.3944
R9515 gnd.n7247 gnd.n7246 19.3944
R9516 gnd.n7246 gnd.n7244 19.3944
R9517 gnd.n7244 gnd.n7241 19.3944
R9518 gnd.n7241 gnd.n7240 19.3944
R9519 gnd.n7240 gnd.n7237 19.3944
R9520 gnd.n7237 gnd.n7236 19.3944
R9521 gnd.n7236 gnd.n7233 19.3944
R9522 gnd.n7233 gnd.n7232 19.3944
R9523 gnd.n7232 gnd.n7229 19.3944
R9524 gnd.n7229 gnd.n7228 19.3944
R9525 gnd.n7228 gnd.n7225 19.3944
R9526 gnd.n7225 gnd.n7224 19.3944
R9527 gnd.n7224 gnd.n7221 19.3944
R9528 gnd.n7219 gnd.n7216 19.3944
R9529 gnd.n7216 gnd.n7215 19.3944
R9530 gnd.n7215 gnd.n7212 19.3944
R9531 gnd.n7212 gnd.n7211 19.3944
R9532 gnd.n7211 gnd.n7208 19.3944
R9533 gnd.n7208 gnd.n7207 19.3944
R9534 gnd.n7207 gnd.n7204 19.3944
R9535 gnd.n7204 gnd.n7203 19.3944
R9536 gnd.n7203 gnd.n7200 19.3944
R9537 gnd.n7200 gnd.n7199 19.3944
R9538 gnd.n7199 gnd.n7196 19.3944
R9539 gnd.n7196 gnd.n7195 19.3944
R9540 gnd.n7195 gnd.n7192 19.3944
R9541 gnd.n7192 gnd.n7191 19.3944
R9542 gnd.n7191 gnd.n7188 19.3944
R9543 gnd.n7188 gnd.n7187 19.3944
R9544 gnd.n7187 gnd.n7184 19.3944
R9545 gnd.n7184 gnd.n7183 19.3944
R9546 gnd.n600 gnd.n580 19.3944
R9547 gnd.n603 gnd.n600 19.3944
R9548 gnd.n603 gnd.n598 19.3944
R9549 gnd.n609 gnd.n598 19.3944
R9550 gnd.n610 gnd.n609 19.3944
R9551 gnd.n613 gnd.n610 19.3944
R9552 gnd.n613 gnd.n596 19.3944
R9553 gnd.n619 gnd.n596 19.3944
R9554 gnd.n620 gnd.n619 19.3944
R9555 gnd.n7130 gnd.n620 19.3944
R9556 gnd.n7130 gnd.n594 19.3944
R9557 gnd.n7149 gnd.n594 19.3944
R9558 gnd.n7149 gnd.n7148 19.3944
R9559 gnd.n7148 gnd.n7147 19.3944
R9560 gnd.n7147 gnd.n7144 19.3944
R9561 gnd.n7144 gnd.n7143 19.3944
R9562 gnd.n7143 gnd.n7141 19.3944
R9563 gnd.n7141 gnd.n7140 19.3944
R9564 gnd.n7140 gnd.n394 19.3944
R9565 gnd.n7403 gnd.n394 19.3944
R9566 gnd.n7403 gnd.n392 19.3944
R9567 gnd.n7413 gnd.n392 19.3944
R9568 gnd.n7413 gnd.n7412 19.3944
R9569 gnd.n7412 gnd.n7411 19.3944
R9570 gnd.n7411 gnd.n360 19.3944
R9571 gnd.n7449 gnd.n360 19.3944
R9572 gnd.n7449 gnd.n358 19.3944
R9573 gnd.n7537 gnd.n358 19.3944
R9574 gnd.n7537 gnd.n7536 19.3944
R9575 gnd.n7536 gnd.n7535 19.3944
R9576 gnd.n7535 gnd.n7532 19.3944
R9577 gnd.n7532 gnd.n7531 19.3944
R9578 gnd.n7531 gnd.n7529 19.3944
R9579 gnd.n7529 gnd.n7528 19.3944
R9580 gnd.n7528 gnd.n7526 19.3944
R9581 gnd.n7526 gnd.n7525 19.3944
R9582 gnd.n7525 gnd.n7524 19.3944
R9583 gnd.n7524 gnd.n7522 19.3944
R9584 gnd.n7522 gnd.n7521 19.3944
R9585 gnd.n7521 gnd.n7519 19.3944
R9586 gnd.n7519 gnd.n7518 19.3944
R9587 gnd.n7518 gnd.n7516 19.3944
R9588 gnd.n7516 gnd.n7515 19.3944
R9589 gnd.n7515 gnd.n7513 19.3944
R9590 gnd.n7513 gnd.n7512 19.3944
R9591 gnd.n7512 gnd.n7510 19.3944
R9592 gnd.n7510 gnd.n7509 19.3944
R9593 gnd.n7509 gnd.n7507 19.3944
R9594 gnd.n7507 gnd.n7506 19.3944
R9595 gnd.n7506 gnd.n7504 19.3944
R9596 gnd.n7504 gnd.n7503 19.3944
R9597 gnd.n7503 gnd.n7501 19.3944
R9598 gnd.n7501 gnd.n7500 19.3944
R9599 gnd.n7500 gnd.n7498 19.3944
R9600 gnd.n7498 gnd.n7497 19.3944
R9601 gnd.n7497 gnd.n7495 19.3944
R9602 gnd.n7495 gnd.n7494 19.3944
R9603 gnd.n7494 gnd.n7491 19.3944
R9604 gnd.n7491 gnd.n7490 19.3944
R9605 gnd.n7490 gnd.n7488 19.3944
R9606 gnd.n7488 gnd.n7487 19.3944
R9607 gnd.n7487 gnd.n204 19.3944
R9608 gnd.n7760 gnd.n204 19.3944
R9609 gnd.n7761 gnd.n7760 19.3944
R9610 gnd.n7799 gnd.n165 19.3944
R9611 gnd.n7794 gnd.n165 19.3944
R9612 gnd.n7794 gnd.n7793 19.3944
R9613 gnd.n7793 gnd.n7792 19.3944
R9614 gnd.n7792 gnd.n172 19.3944
R9615 gnd.n7787 gnd.n172 19.3944
R9616 gnd.n7787 gnd.n7786 19.3944
R9617 gnd.n7786 gnd.n7785 19.3944
R9618 gnd.n7785 gnd.n179 19.3944
R9619 gnd.n7780 gnd.n179 19.3944
R9620 gnd.n7780 gnd.n7779 19.3944
R9621 gnd.n7779 gnd.n7778 19.3944
R9622 gnd.n7778 gnd.n186 19.3944
R9623 gnd.n7773 gnd.n186 19.3944
R9624 gnd.n7773 gnd.n7772 19.3944
R9625 gnd.n7772 gnd.n7771 19.3944
R9626 gnd.n7771 gnd.n193 19.3944
R9627 gnd.n7766 gnd.n193 19.3944
R9628 gnd.n7832 gnd.n7831 19.3944
R9629 gnd.n7831 gnd.n7830 19.3944
R9630 gnd.n7830 gnd.n137 19.3944
R9631 gnd.n7825 gnd.n137 19.3944
R9632 gnd.n7825 gnd.n7824 19.3944
R9633 gnd.n7824 gnd.n7823 19.3944
R9634 gnd.n7823 gnd.n144 19.3944
R9635 gnd.n7818 gnd.n144 19.3944
R9636 gnd.n7818 gnd.n7817 19.3944
R9637 gnd.n7817 gnd.n7816 19.3944
R9638 gnd.n7816 gnd.n151 19.3944
R9639 gnd.n7811 gnd.n151 19.3944
R9640 gnd.n7811 gnd.n7810 19.3944
R9641 gnd.n7810 gnd.n7809 19.3944
R9642 gnd.n7809 gnd.n158 19.3944
R9643 gnd.n7804 gnd.n158 19.3944
R9644 gnd.n7804 gnd.n7803 19.3944
R9645 gnd.n7263 gnd.n493 19.3944
R9646 gnd.n7263 gnd.n491 19.3944
R9647 gnd.n7267 gnd.n491 19.3944
R9648 gnd.n7267 gnd.n475 19.3944
R9649 gnd.n7279 gnd.n475 19.3944
R9650 gnd.n7279 gnd.n473 19.3944
R9651 gnd.n7283 gnd.n473 19.3944
R9652 gnd.n7283 gnd.n458 19.3944
R9653 gnd.n7295 gnd.n458 19.3944
R9654 gnd.n7295 gnd.n456 19.3944
R9655 gnd.n7299 gnd.n456 19.3944
R9656 gnd.n7299 gnd.n438 19.3944
R9657 gnd.n7317 gnd.n438 19.3944
R9658 gnd.n7317 gnd.n436 19.3944
R9659 gnd.n7323 gnd.n436 19.3944
R9660 gnd.n7323 gnd.n7322 19.3944
R9661 gnd.n7322 gnd.n403 19.3944
R9662 gnd.n7393 gnd.n403 19.3944
R9663 gnd.n7393 gnd.n401 19.3944
R9664 gnd.n7399 gnd.n401 19.3944
R9665 gnd.n7399 gnd.n7398 19.3944
R9666 gnd.n7398 gnd.n370 19.3944
R9667 gnd.n7440 gnd.n370 19.3944
R9668 gnd.n7440 gnd.n368 19.3944
R9669 gnd.n7444 gnd.n368 19.3944
R9670 gnd.n7445 gnd.n7444 19.3944
R9671 gnd.n7445 gnd.n308 19.3944
R9672 gnd.n7587 gnd.n7586 19.3944
R9673 gnd.n347 gnd.n346 19.3944
R9674 gnd.n7553 gnd.n7552 19.3944
R9675 gnd.n331 gnd.n330 19.3944
R9676 gnd.n7567 gnd.n301 19.3944
R9677 gnd.n7591 gnd.n301 19.3944
R9678 gnd.n7591 gnd.n287 19.3944
R9679 gnd.n7603 gnd.n287 19.3944
R9680 gnd.n7603 gnd.n285 19.3944
R9681 gnd.n7607 gnd.n285 19.3944
R9682 gnd.n7607 gnd.n273 19.3944
R9683 gnd.n7619 gnd.n273 19.3944
R9684 gnd.n7619 gnd.n271 19.3944
R9685 gnd.n7623 gnd.n271 19.3944
R9686 gnd.n7623 gnd.n257 19.3944
R9687 gnd.n7635 gnd.n257 19.3944
R9688 gnd.n7635 gnd.n255 19.3944
R9689 gnd.n7639 gnd.n255 19.3944
R9690 gnd.n7639 gnd.n243 19.3944
R9691 gnd.n7651 gnd.n243 19.3944
R9692 gnd.n7651 gnd.n241 19.3944
R9693 gnd.n7655 gnd.n241 19.3944
R9694 gnd.n7655 gnd.n227 19.3944
R9695 gnd.n7667 gnd.n227 19.3944
R9696 gnd.n7667 gnd.n225 19.3944
R9697 gnd.n7671 gnd.n225 19.3944
R9698 gnd.n7671 gnd.n211 19.3944
R9699 gnd.n7751 gnd.n211 19.3944
R9700 gnd.n7751 gnd.n209 19.3944
R9701 gnd.n7755 gnd.n209 19.3944
R9702 gnd.n7755 gnd.n132 19.3944
R9703 gnd.n7835 gnd.n132 19.3944
R9704 gnd.n4753 gnd.n4752 19.3944
R9705 gnd.n4752 gnd.n4569 19.3944
R9706 gnd.n4747 gnd.n4569 19.3944
R9707 gnd.n4747 gnd.n4746 19.3944
R9708 gnd.n4746 gnd.n4574 19.3944
R9709 gnd.n4741 gnd.n4574 19.3944
R9710 gnd.n4741 gnd.n4740 19.3944
R9711 gnd.n4740 gnd.n4739 19.3944
R9712 gnd.n4739 gnd.n4580 19.3944
R9713 gnd.n4733 gnd.n4580 19.3944
R9714 gnd.n4733 gnd.n4732 19.3944
R9715 gnd.n4732 gnd.n4731 19.3944
R9716 gnd.n4731 gnd.n4586 19.3944
R9717 gnd.n4725 gnd.n4586 19.3944
R9718 gnd.n4725 gnd.n4724 19.3944
R9719 gnd.n4724 gnd.n4723 19.3944
R9720 gnd.n4723 gnd.n4592 19.3944
R9721 gnd.n4717 gnd.n4716 19.3944
R9722 gnd.n4716 gnd.n4715 19.3944
R9723 gnd.n4715 gnd.n4601 19.3944
R9724 gnd.n4709 gnd.n4601 19.3944
R9725 gnd.n4709 gnd.n4708 19.3944
R9726 gnd.n4708 gnd.n4707 19.3944
R9727 gnd.n4707 gnd.n4607 19.3944
R9728 gnd.n4701 gnd.n4607 19.3944
R9729 gnd.n4701 gnd.n4700 19.3944
R9730 gnd.n4700 gnd.n4699 19.3944
R9731 gnd.n4699 gnd.n4613 19.3944
R9732 gnd.n4693 gnd.n4613 19.3944
R9733 gnd.n4693 gnd.n4692 19.3944
R9734 gnd.n4692 gnd.n4691 19.3944
R9735 gnd.n4691 gnd.n4619 19.3944
R9736 gnd.n4685 gnd.n4619 19.3944
R9737 gnd.n4685 gnd.n4684 19.3944
R9738 gnd.n4684 gnd.n4683 19.3944
R9739 gnd.n4760 gnd.n1561 19.3944
R9740 gnd.n4764 gnd.n1561 19.3944
R9741 gnd.n4764 gnd.n1548 19.3944
R9742 gnd.n4776 gnd.n1548 19.3944
R9743 gnd.n4776 gnd.n1546 19.3944
R9744 gnd.n4780 gnd.n1546 19.3944
R9745 gnd.n4780 gnd.n1531 19.3944
R9746 gnd.n4792 gnd.n1531 19.3944
R9747 gnd.n4792 gnd.n1529 19.3944
R9748 gnd.n4796 gnd.n1529 19.3944
R9749 gnd.n4796 gnd.n1516 19.3944
R9750 gnd.n4808 gnd.n1516 19.3944
R9751 gnd.n4808 gnd.n1514 19.3944
R9752 gnd.n4812 gnd.n1514 19.3944
R9753 gnd.n4812 gnd.n1499 19.3944
R9754 gnd.n4824 gnd.n1499 19.3944
R9755 gnd.n4824 gnd.n1497 19.3944
R9756 gnd.n4836 gnd.n1497 19.3944
R9757 gnd.n4836 gnd.n4835 19.3944
R9758 gnd.n4835 gnd.n4834 19.3944
R9759 gnd.n4834 gnd.n4833 19.3944
R9760 gnd.n4833 gnd.n1463 19.3944
R9761 gnd.n4877 gnd.n1463 19.3944
R9762 gnd.n4877 gnd.n4876 19.3944
R9763 gnd.n4876 gnd.n4875 19.3944
R9764 gnd.n4875 gnd.n1472 19.3944
R9765 gnd.n1472 gnd.n1471 19.3944
R9766 gnd.n1471 gnd.n1398 19.3944
R9767 gnd.n5236 gnd.n1398 19.3944
R9768 gnd.n5236 gnd.n5235 19.3944
R9769 gnd.n5235 gnd.n5234 19.3944
R9770 gnd.n5234 gnd.n1402 19.3944
R9771 gnd.n5209 gnd.n1402 19.3944
R9772 gnd.n5209 gnd.n1427 19.3944
R9773 gnd.n5213 gnd.n1427 19.3944
R9774 gnd.n5213 gnd.n1375 19.3944
R9775 gnd.n5248 gnd.n1375 19.3944
R9776 gnd.n5248 gnd.n1373 19.3944
R9777 gnd.n5252 gnd.n1373 19.3944
R9778 gnd.n5252 gnd.n1358 19.3944
R9779 gnd.n5264 gnd.n1358 19.3944
R9780 gnd.n5264 gnd.n1356 19.3944
R9781 gnd.n5268 gnd.n1356 19.3944
R9782 gnd.n5268 gnd.n1340 19.3944
R9783 gnd.n5280 gnd.n1340 19.3944
R9784 gnd.n5280 gnd.n1338 19.3944
R9785 gnd.n5284 gnd.n1338 19.3944
R9786 gnd.n5284 gnd.n1323 19.3944
R9787 gnd.n5296 gnd.n1323 19.3944
R9788 gnd.n5296 gnd.n1321 19.3944
R9789 gnd.n5300 gnd.n1321 19.3944
R9790 gnd.n5300 gnd.n1305 19.3944
R9791 gnd.n5312 gnd.n1305 19.3944
R9792 gnd.n5312 gnd.n1303 19.3944
R9793 gnd.n5316 gnd.n1303 19.3944
R9794 gnd.n5316 gnd.n1288 19.3944
R9795 gnd.n5328 gnd.n1288 19.3944
R9796 gnd.n5328 gnd.n1286 19.3944
R9797 gnd.n5332 gnd.n1286 19.3944
R9798 gnd.n5332 gnd.n1269 19.3944
R9799 gnd.n5346 gnd.n1269 19.3944
R9800 gnd.n5346 gnd.n1267 19.3944
R9801 gnd.n5662 gnd.n1267 19.3944
R9802 gnd.n5662 gnd.n5661 19.3944
R9803 gnd.n4468 gnd.n4467 19.3944
R9804 gnd.n4473 gnd.n4468 19.3944
R9805 gnd.n4473 gnd.n4465 19.3944
R9806 gnd.n4477 gnd.n4465 19.3944
R9807 gnd.n4477 gnd.n4463 19.3944
R9808 gnd.n4483 gnd.n4463 19.3944
R9809 gnd.n4483 gnd.n4461 19.3944
R9810 gnd.n4487 gnd.n4461 19.3944
R9811 gnd.n4487 gnd.n4459 19.3944
R9812 gnd.n4493 gnd.n4459 19.3944
R9813 gnd.n4493 gnd.n4457 19.3944
R9814 gnd.n4497 gnd.n4457 19.3944
R9815 gnd.n4497 gnd.n4455 19.3944
R9816 gnd.n4503 gnd.n4455 19.3944
R9817 gnd.n4503 gnd.n4453 19.3944
R9818 gnd.n4507 gnd.n4453 19.3944
R9819 gnd.n4564 gnd.n4447 19.3944
R9820 gnd.n4564 gnd.n4563 19.3944
R9821 gnd.n4563 gnd.n4562 19.3944
R9822 gnd.n4562 gnd.n4560 19.3944
R9823 gnd.n4560 gnd.n4559 19.3944
R9824 gnd.n4559 gnd.n4557 19.3944
R9825 gnd.n4557 gnd.n4556 19.3944
R9826 gnd.n4556 gnd.n4554 19.3944
R9827 gnd.n4554 gnd.n4553 19.3944
R9828 gnd.n4553 gnd.n4551 19.3944
R9829 gnd.n4551 gnd.n4550 19.3944
R9830 gnd.n4550 gnd.n4548 19.3944
R9831 gnd.n4548 gnd.n4547 19.3944
R9832 gnd.n4547 gnd.n4545 19.3944
R9833 gnd.n4545 gnd.n4544 19.3944
R9834 gnd.n4544 gnd.n4542 19.3944
R9835 gnd.n4542 gnd.n4541 19.3944
R9836 gnd.n4541 gnd.n4539 19.3944
R9837 gnd.n4539 gnd.n4538 19.3944
R9838 gnd.n4538 gnd.n4536 19.3944
R9839 gnd.n4536 gnd.n1476 19.3944
R9840 gnd.n4863 gnd.n1476 19.3944
R9841 gnd.n4864 gnd.n4863 19.3944
R9842 gnd.n4864 gnd.n1474 19.3944
R9843 gnd.n4871 gnd.n1474 19.3944
R9844 gnd.n4871 gnd.n4870 19.3944
R9845 gnd.n4870 gnd.n1440 19.3944
R9846 gnd.n4903 gnd.n1440 19.3944
R9847 gnd.n4904 gnd.n4903 19.3944
R9848 gnd.n4906 gnd.n4904 19.3944
R9849 gnd.n4906 gnd.n1438 19.3944
R9850 gnd.n4910 gnd.n1438 19.3944
R9851 gnd.n4911 gnd.n4910 19.3944
R9852 gnd.n4914 gnd.n4911 19.3944
R9853 gnd.n4914 gnd.n1435 19.3944
R9854 gnd.n5195 gnd.n1435 19.3944
R9855 gnd.n5195 gnd.n1436 19.3944
R9856 gnd.n5191 gnd.n1436 19.3944
R9857 gnd.n5191 gnd.n5190 19.3944
R9858 gnd.n5190 gnd.n5189 19.3944
R9859 gnd.n5189 gnd.n4920 19.3944
R9860 gnd.n5185 gnd.n4920 19.3944
R9861 gnd.n5185 gnd.n5184 19.3944
R9862 gnd.n5184 gnd.n5183 19.3944
R9863 gnd.n5183 gnd.n4924 19.3944
R9864 gnd.n5179 gnd.n4924 19.3944
R9865 gnd.n5179 gnd.n5178 19.3944
R9866 gnd.n5178 gnd.n5177 19.3944
R9867 gnd.n5177 gnd.n4928 19.3944
R9868 gnd.n5173 gnd.n4928 19.3944
R9869 gnd.n5173 gnd.n5172 19.3944
R9870 gnd.n5172 gnd.n5171 19.3944
R9871 gnd.n5171 gnd.n4932 19.3944
R9872 gnd.n5167 gnd.n4932 19.3944
R9873 gnd.n5167 gnd.n5166 19.3944
R9874 gnd.n5166 gnd.n5165 19.3944
R9875 gnd.n5165 gnd.n4936 19.3944
R9876 gnd.n5161 gnd.n4936 19.3944
R9877 gnd.n5161 gnd.n5160 19.3944
R9878 gnd.n5160 gnd.n5159 19.3944
R9879 gnd.n5159 gnd.n5120 19.3944
R9880 gnd.n5155 gnd.n5120 19.3944
R9881 gnd.n5155 gnd.n5154 19.3944
R9882 gnd.n5154 gnd.n1174 19.3944
R9883 gnd.n4674 gnd.n4673 19.3944
R9884 gnd.n4673 gnd.n4672 19.3944
R9885 gnd.n4672 gnd.n4671 19.3944
R9886 gnd.n4671 gnd.n4669 19.3944
R9887 gnd.n4669 gnd.n4668 19.3944
R9888 gnd.n4668 gnd.n4666 19.3944
R9889 gnd.n4666 gnd.n4665 19.3944
R9890 gnd.n4665 gnd.n4663 19.3944
R9891 gnd.n4663 gnd.n4662 19.3944
R9892 gnd.n4662 gnd.n4660 19.3944
R9893 gnd.n4660 gnd.n4659 19.3944
R9894 gnd.n4659 gnd.n4657 19.3944
R9895 gnd.n4657 gnd.n4656 19.3944
R9896 gnd.n4656 gnd.n4654 19.3944
R9897 gnd.n4654 gnd.n4653 19.3944
R9898 gnd.n4653 gnd.n4651 19.3944
R9899 gnd.n4651 gnd.n4650 19.3944
R9900 gnd.n4650 gnd.n4648 19.3944
R9901 gnd.n4648 gnd.n1482 19.3944
R9902 gnd.n4850 gnd.n1482 19.3944
R9903 gnd.n4850 gnd.n1480 19.3944
R9904 gnd.n4859 gnd.n1480 19.3944
R9905 gnd.n4859 gnd.n4858 19.3944
R9906 gnd.n4858 gnd.n4857 19.3944
R9907 gnd.n4857 gnd.n1447 19.3944
R9908 gnd.n4890 gnd.n1447 19.3944
R9909 gnd.n4890 gnd.n1445 19.3944
R9910 gnd.n4899 gnd.n1445 19.3944
R9911 gnd.n4899 gnd.n4898 19.3944
R9912 gnd.n4898 gnd.n4897 19.3944
R9913 gnd.n4897 gnd.n1430 19.3944
R9914 gnd.n5205 gnd.n1430 19.3944
R9915 gnd.n5205 gnd.n5204 19.3944
R9916 gnd.n5204 gnd.n5201 19.3944
R9917 gnd.n5201 gnd.n5200 19.3944
R9918 gnd.n5200 gnd.n5199 19.3944
R9919 gnd.n5199 gnd.n1434 19.3944
R9920 gnd.n4995 gnd.n1434 19.3944
R9921 gnd.n4996 gnd.n4995 19.3944
R9922 gnd.n4999 gnd.n4996 19.3944
R9923 gnd.n4999 gnd.n4957 19.3944
R9924 gnd.n5005 gnd.n4957 19.3944
R9925 gnd.n5006 gnd.n5005 19.3944
R9926 gnd.n5009 gnd.n5006 19.3944
R9927 gnd.n5009 gnd.n4955 19.3944
R9928 gnd.n5031 gnd.n4955 19.3944
R9929 gnd.n5031 gnd.n5030 19.3944
R9930 gnd.n5030 gnd.n5029 19.3944
R9931 gnd.n5029 gnd.n5026 19.3944
R9932 gnd.n5026 gnd.n5025 19.3944
R9933 gnd.n5025 gnd.n5022 19.3944
R9934 gnd.n5022 gnd.n5021 19.3944
R9935 gnd.n5021 gnd.n4943 19.3944
R9936 gnd.n5099 gnd.n4943 19.3944
R9937 gnd.n5099 gnd.n4941 19.3944
R9938 gnd.n5105 gnd.n4941 19.3944
R9939 gnd.n5106 gnd.n5105 19.3944
R9940 gnd.n5109 gnd.n5106 19.3944
R9941 gnd.n5109 gnd.n4939 19.3944
R9942 gnd.n5116 gnd.n4939 19.3944
R9943 gnd.n5116 gnd.n5115 19.3944
R9944 gnd.n5115 gnd.n1263 19.3944
R9945 gnd.n5666 gnd.n1263 19.3944
R9946 gnd.n5667 gnd.n5666 19.3944
R9947 gnd.n5705 gnd.n5704 19.3944
R9948 gnd.n5704 gnd.n5703 19.3944
R9949 gnd.n5703 gnd.n1229 19.3944
R9950 gnd.n5698 gnd.n1229 19.3944
R9951 gnd.n5698 gnd.n5697 19.3944
R9952 gnd.n5697 gnd.n5696 19.3944
R9953 gnd.n5696 gnd.n1236 19.3944
R9954 gnd.n5691 gnd.n1236 19.3944
R9955 gnd.n5691 gnd.n5690 19.3944
R9956 gnd.n5690 gnd.n5689 19.3944
R9957 gnd.n5689 gnd.n1243 19.3944
R9958 gnd.n5684 gnd.n1243 19.3944
R9959 gnd.n5684 gnd.n5683 19.3944
R9960 gnd.n5683 gnd.n5682 19.3944
R9961 gnd.n5682 gnd.n1250 19.3944
R9962 gnd.n5677 gnd.n1250 19.3944
R9963 gnd.n5677 gnd.n5676 19.3944
R9964 gnd.n5676 gnd.n5675 19.3944
R9965 gnd.n5736 gnd.n5735 19.3944
R9966 gnd.n5735 gnd.n1184 19.3944
R9967 gnd.n1197 gnd.n1184 19.3944
R9968 gnd.n5728 gnd.n1197 19.3944
R9969 gnd.n5728 gnd.n5727 19.3944
R9970 gnd.n5727 gnd.n5726 19.3944
R9971 gnd.n5726 gnd.n1204 19.3944
R9972 gnd.n5721 gnd.n1204 19.3944
R9973 gnd.n5721 gnd.n5720 19.3944
R9974 gnd.n5720 gnd.n5719 19.3944
R9975 gnd.n5719 gnd.n1211 19.3944
R9976 gnd.n5714 gnd.n1211 19.3944
R9977 gnd.n5714 gnd.n5713 19.3944
R9978 gnd.n5713 gnd.n5712 19.3944
R9979 gnd.n5712 gnd.n1218 19.3944
R9980 gnd.n4756 gnd.n1556 19.3944
R9981 gnd.n4768 gnd.n1556 19.3944
R9982 gnd.n4768 gnd.n1554 19.3944
R9983 gnd.n4772 gnd.n1554 19.3944
R9984 gnd.n4772 gnd.n1540 19.3944
R9985 gnd.n4784 gnd.n1540 19.3944
R9986 gnd.n4784 gnd.n1538 19.3944
R9987 gnd.n4788 gnd.n1538 19.3944
R9988 gnd.n4788 gnd.n1524 19.3944
R9989 gnd.n4800 gnd.n1524 19.3944
R9990 gnd.n4800 gnd.n1522 19.3944
R9991 gnd.n4804 gnd.n1522 19.3944
R9992 gnd.n4804 gnd.n1508 19.3944
R9993 gnd.n4816 gnd.n1508 19.3944
R9994 gnd.n4816 gnd.n1506 19.3944
R9995 gnd.n4820 gnd.n1506 19.3944
R9996 gnd.n4820 gnd.n1491 19.3944
R9997 gnd.n4840 gnd.n1491 19.3944
R9998 gnd.n4840 gnd.n1489 19.3944
R9999 gnd.n4846 gnd.n1489 19.3944
R10000 gnd.n4846 gnd.n4845 19.3944
R10001 gnd.n4845 gnd.n1455 19.3944
R10002 gnd.n4881 gnd.n1455 19.3944
R10003 gnd.n4881 gnd.n1453 19.3944
R10004 gnd.n4885 gnd.n1453 19.3944
R10005 gnd.n4886 gnd.n4885 19.3944
R10006 gnd.n4886 gnd.n1389 19.3944
R10007 gnd.n5241 gnd.n5240 19.3944
R10008 gnd.n5230 gnd.n5229 19.3944
R10009 gnd.n1409 gnd.n1408 19.3944
R10010 gnd.n5217 gnd.n5216 19.3944
R10011 gnd.n5244 gnd.n1382 19.3944
R10012 gnd.n5244 gnd.n1367 19.3944
R10013 gnd.n5256 gnd.n1367 19.3944
R10014 gnd.n5256 gnd.n1365 19.3944
R10015 gnd.n5260 gnd.n1365 19.3944
R10016 gnd.n5260 gnd.n1349 19.3944
R10017 gnd.n5272 gnd.n1349 19.3944
R10018 gnd.n5272 gnd.n1347 19.3944
R10019 gnd.n5276 gnd.n1347 19.3944
R10020 gnd.n5276 gnd.n1332 19.3944
R10021 gnd.n5288 gnd.n1332 19.3944
R10022 gnd.n5288 gnd.n1330 19.3944
R10023 gnd.n5292 gnd.n1330 19.3944
R10024 gnd.n5292 gnd.n1314 19.3944
R10025 gnd.n5304 gnd.n1314 19.3944
R10026 gnd.n5304 gnd.n1312 19.3944
R10027 gnd.n5308 gnd.n1312 19.3944
R10028 gnd.n5308 gnd.n1297 19.3944
R10029 gnd.n5320 gnd.n1297 19.3944
R10030 gnd.n5320 gnd.n1295 19.3944
R10031 gnd.n5324 gnd.n1295 19.3944
R10032 gnd.n5324 gnd.n1279 19.3944
R10033 gnd.n5336 gnd.n1279 19.3944
R10034 gnd.n5336 gnd.n1277 19.3944
R10035 gnd.n5342 gnd.n1277 19.3944
R10036 gnd.n5342 gnd.n5341 19.3944
R10037 gnd.n5341 gnd.n1181 19.3944
R10038 gnd.n5739 gnd.n1181 19.3944
R10039 gnd.n2847 gnd.n1781 19.3944
R10040 gnd.n2847 gnd.n1779 19.3944
R10041 gnd.n2851 gnd.n1779 19.3944
R10042 gnd.n2851 gnd.n1775 19.3944
R10043 gnd.n2857 gnd.n1775 19.3944
R10044 gnd.n2857 gnd.n1773 19.3944
R10045 gnd.n2861 gnd.n1773 19.3944
R10046 gnd.n2861 gnd.n1769 19.3944
R10047 gnd.n2867 gnd.n1769 19.3944
R10048 gnd.n2867 gnd.n1767 19.3944
R10049 gnd.n2871 gnd.n1767 19.3944
R10050 gnd.n2871 gnd.n1763 19.3944
R10051 gnd.n2877 gnd.n1763 19.3944
R10052 gnd.n2877 gnd.n1761 19.3944
R10053 gnd.n2881 gnd.n1761 19.3944
R10054 gnd.n2881 gnd.n1757 19.3944
R10055 gnd.n2887 gnd.n1757 19.3944
R10056 gnd.n2887 gnd.n1755 19.3944
R10057 gnd.n2891 gnd.n1755 19.3944
R10058 gnd.n2891 gnd.n1751 19.3944
R10059 gnd.n2897 gnd.n1751 19.3944
R10060 gnd.n2897 gnd.n1749 19.3944
R10061 gnd.n2901 gnd.n1749 19.3944
R10062 gnd.n2901 gnd.n1745 19.3944
R10063 gnd.n2907 gnd.n1745 19.3944
R10064 gnd.n2907 gnd.n1743 19.3944
R10065 gnd.n2911 gnd.n1743 19.3944
R10066 gnd.n2911 gnd.n1739 19.3944
R10067 gnd.n2917 gnd.n1739 19.3944
R10068 gnd.n2917 gnd.n1737 19.3944
R10069 gnd.n2921 gnd.n1737 19.3944
R10070 gnd.n2921 gnd.n1733 19.3944
R10071 gnd.n2927 gnd.n1733 19.3944
R10072 gnd.n2927 gnd.n1731 19.3944
R10073 gnd.n2931 gnd.n1731 19.3944
R10074 gnd.n2931 gnd.n1727 19.3944
R10075 gnd.n2937 gnd.n1727 19.3944
R10076 gnd.n2937 gnd.n1725 19.3944
R10077 gnd.n2941 gnd.n1725 19.3944
R10078 gnd.n2941 gnd.n1721 19.3944
R10079 gnd.n2947 gnd.n1721 19.3944
R10080 gnd.n2947 gnd.n1719 19.3944
R10081 gnd.n2951 gnd.n1719 19.3944
R10082 gnd.n2951 gnd.n1715 19.3944
R10083 gnd.n2957 gnd.n1715 19.3944
R10084 gnd.n2957 gnd.n1713 19.3944
R10085 gnd.n2961 gnd.n1713 19.3944
R10086 gnd.n2961 gnd.n1709 19.3944
R10087 gnd.n2967 gnd.n1709 19.3944
R10088 gnd.n2967 gnd.n1707 19.3944
R10089 gnd.n2971 gnd.n1707 19.3944
R10090 gnd.n2971 gnd.n1703 19.3944
R10091 gnd.n2977 gnd.n1703 19.3944
R10092 gnd.n2977 gnd.n1701 19.3944
R10093 gnd.n2981 gnd.n1701 19.3944
R10094 gnd.n2981 gnd.n1697 19.3944
R10095 gnd.n2987 gnd.n1697 19.3944
R10096 gnd.n2987 gnd.n1695 19.3944
R10097 gnd.n2991 gnd.n1695 19.3944
R10098 gnd.n2991 gnd.n1691 19.3944
R10099 gnd.n2997 gnd.n1691 19.3944
R10100 gnd.n2997 gnd.n1689 19.3944
R10101 gnd.n3001 gnd.n1689 19.3944
R10102 gnd.n3001 gnd.n1685 19.3944
R10103 gnd.n3007 gnd.n1685 19.3944
R10104 gnd.n3007 gnd.n1683 19.3944
R10105 gnd.n3011 gnd.n1683 19.3944
R10106 gnd.n3011 gnd.n1679 19.3944
R10107 gnd.n3017 gnd.n1679 19.3944
R10108 gnd.n3017 gnd.n1677 19.3944
R10109 gnd.n3021 gnd.n1677 19.3944
R10110 gnd.n3021 gnd.n1673 19.3944
R10111 gnd.n3027 gnd.n1673 19.3944
R10112 gnd.n3027 gnd.n1671 19.3944
R10113 gnd.n3031 gnd.n1671 19.3944
R10114 gnd.n3031 gnd.n1667 19.3944
R10115 gnd.n3037 gnd.n1667 19.3944
R10116 gnd.n3037 gnd.n1665 19.3944
R10117 gnd.n3041 gnd.n1665 19.3944
R10118 gnd.n3041 gnd.n1661 19.3944
R10119 gnd.n3047 gnd.n1661 19.3944
R10120 gnd.n3047 gnd.n1659 19.3944
R10121 gnd.n3058 gnd.n1659 19.3944
R10122 gnd.n3058 gnd.n3057 19.3944
R10123 gnd.n5656 gnd.n5655 19.3944
R10124 gnd.n5655 gnd.n5654 19.3944
R10125 gnd.n5654 gnd.n5360 19.3944
R10126 gnd.n5650 gnd.n5360 19.3944
R10127 gnd.n5650 gnd.n5649 19.3944
R10128 gnd.n5649 gnd.n5648 19.3944
R10129 gnd.n5648 gnd.n5364 19.3944
R10130 gnd.n5644 gnd.n5364 19.3944
R10131 gnd.n5644 gnd.n5643 19.3944
R10132 gnd.n5643 gnd.n5642 19.3944
R10133 gnd.n5642 gnd.n5368 19.3944
R10134 gnd.n5638 gnd.n5368 19.3944
R10135 gnd.n5638 gnd.n5637 19.3944
R10136 gnd.n5637 gnd.n5636 19.3944
R10137 gnd.n5636 gnd.n5372 19.3944
R10138 gnd.n5632 gnd.n5372 19.3944
R10139 gnd.n5632 gnd.n5631 19.3944
R10140 gnd.n5631 gnd.n5630 19.3944
R10141 gnd.n5630 gnd.n5376 19.3944
R10142 gnd.n5626 gnd.n5376 19.3944
R10143 gnd.n5626 gnd.n5625 19.3944
R10144 gnd.n5625 gnd.n5624 19.3944
R10145 gnd.n5624 gnd.n1008 19.3944
R10146 gnd.n5901 gnd.n1008 19.3944
R10147 gnd.n5901 gnd.n1005 19.3944
R10148 gnd.n5905 gnd.n1005 19.3944
R10149 gnd.n5906 gnd.n5905 19.3944
R10150 gnd.n5909 gnd.n5906 19.3944
R10151 gnd.n5909 gnd.n1002 19.3944
R10152 gnd.n5960 gnd.n1002 19.3944
R10153 gnd.n5960 gnd.n1003 19.3944
R10154 gnd.n5956 gnd.n1003 19.3944
R10155 gnd.n5956 gnd.n5955 19.3944
R10156 gnd.n5955 gnd.n5954 19.3944
R10157 gnd.n5954 gnd.n5946 19.3944
R10158 gnd.n5950 gnd.n5946 19.3944
R10159 gnd.n5950 gnd.n5949 19.3944
R10160 gnd.n5949 gnd.n906 19.3944
R10161 gnd.n6081 gnd.n906 19.3944
R10162 gnd.n6081 gnd.n903 19.3944
R10163 gnd.n6085 gnd.n903 19.3944
R10164 gnd.n6086 gnd.n6085 19.3944
R10165 gnd.n6088 gnd.n6086 19.3944
R10166 gnd.n6088 gnd.n900 19.3944
R10167 gnd.n6818 gnd.n900 19.3944
R10168 gnd.n6818 gnd.n901 19.3944
R10169 gnd.n6814 gnd.n901 19.3944
R10170 gnd.n6814 gnd.n6813 19.3944
R10171 gnd.n6813 gnd.n6812 19.3944
R10172 gnd.n6812 gnd.n6094 19.3944
R10173 gnd.n6808 gnd.n6094 19.3944
R10174 gnd.n6808 gnd.n6807 19.3944
R10175 gnd.n6807 gnd.n6806 19.3944
R10176 gnd.n6806 gnd.n6098 19.3944
R10177 gnd.n6802 gnd.n6098 19.3944
R10178 gnd.n6802 gnd.n6801 19.3944
R10179 gnd.n6801 gnd.n6800 19.3944
R10180 gnd.n6800 gnd.n6102 19.3944
R10181 gnd.n6796 gnd.n6102 19.3944
R10182 gnd.n6796 gnd.n6795 19.3944
R10183 gnd.n6795 gnd.n6794 19.3944
R10184 gnd.n6794 gnd.n6106 19.3944
R10185 gnd.n6790 gnd.n6106 19.3944
R10186 gnd.n6790 gnd.n6789 19.3944
R10187 gnd.n6789 gnd.n6788 19.3944
R10188 gnd.n6788 gnd.n6110 19.3944
R10189 gnd.n6784 gnd.n6110 19.3944
R10190 gnd.n6784 gnd.n6783 19.3944
R10191 gnd.n6783 gnd.n6782 19.3944
R10192 gnd.n6782 gnd.n6114 19.3944
R10193 gnd.n6778 gnd.n6114 19.3944
R10194 gnd.n6778 gnd.n6777 19.3944
R10195 gnd.n6777 gnd.n6776 19.3944
R10196 gnd.n6776 gnd.n6118 19.3944
R10197 gnd.n6772 gnd.n6118 19.3944
R10198 gnd.n6772 gnd.n6771 19.3944
R10199 gnd.n6771 gnd.n6770 19.3944
R10200 gnd.n6770 gnd.n6122 19.3944
R10201 gnd.n6766 gnd.n6122 19.3944
R10202 gnd.n6766 gnd.n6765 19.3944
R10203 gnd.n6765 gnd.n6764 19.3944
R10204 gnd.n6764 gnd.n6575 19.3944
R10205 gnd.n6760 gnd.n6575 19.3944
R10206 gnd.n6760 gnd.n6759 19.3944
R10207 gnd.n6759 gnd.n6758 19.3944
R10208 gnd.n6758 gnd.n6580 19.3944
R10209 gnd.n6754 gnd.n6580 19.3944
R10210 gnd.n6754 gnd.n6753 19.3944
R10211 gnd.n6753 gnd.n6752 19.3944
R10212 gnd.n6752 gnd.n6584 19.3944
R10213 gnd.n6748 gnd.n6584 19.3944
R10214 gnd.n6748 gnd.n6747 19.3944
R10215 gnd.n6747 gnd.n6746 19.3944
R10216 gnd.n6746 gnd.n6588 19.3944
R10217 gnd.n6742 gnd.n6588 19.3944
R10218 gnd.n6742 gnd.n6741 19.3944
R10219 gnd.n6741 gnd.n6740 19.3944
R10220 gnd.n6740 gnd.n6592 19.3944
R10221 gnd.n6736 gnd.n6592 19.3944
R10222 gnd.n6736 gnd.n6735 19.3944
R10223 gnd.n6735 gnd.n6734 19.3944
R10224 gnd.n6669 gnd.n6668 19.3944
R10225 gnd.n6668 gnd.n656 19.3944
R10226 gnd.n7074 gnd.n656 19.3944
R10227 gnd.n6731 gnd.n6596 19.3944
R10228 gnd.n6724 gnd.n6596 19.3944
R10229 gnd.n6724 gnd.n6723 19.3944
R10230 gnd.n6723 gnd.n6608 19.3944
R10231 gnd.n6716 gnd.n6608 19.3944
R10232 gnd.n6716 gnd.n6715 19.3944
R10233 gnd.n6715 gnd.n6616 19.3944
R10234 gnd.n6708 gnd.n6616 19.3944
R10235 gnd.n6708 gnd.n6707 19.3944
R10236 gnd.n6707 gnd.n6628 19.3944
R10237 gnd.n6700 gnd.n6628 19.3944
R10238 gnd.n6700 gnd.n6699 19.3944
R10239 gnd.n6699 gnd.n6636 19.3944
R10240 gnd.n6692 gnd.n6636 19.3944
R10241 gnd.n6692 gnd.n6691 19.3944
R10242 gnd.n6691 gnd.n6648 19.3944
R10243 gnd.n6681 gnd.n6648 19.3944
R10244 gnd.n6681 gnd.n6680 19.3944
R10245 gnd.n6680 gnd.n6679 19.3944
R10246 gnd.n6679 gnd.n6655 19.3944
R10247 gnd.n6675 gnd.n6655 19.3944
R10248 gnd.n6675 gnd.n6674 19.3944
R10249 gnd.n6674 gnd.n6673 19.3944
R10250 gnd.n6673 gnd.n6661 19.3944
R10251 gnd.n5597 gnd.n5422 19.2005
R10252 gnd.n6426 gnd.n6129 19.2005
R10253 gnd.n5994 gnd.n971 19.1199
R10254 gnd.n6849 gnd.n868 19.1199
R10255 gnd.n6193 gnd.n828 19.1199
R10256 gnd.n6953 gnd.n767 19.1199
R10257 gnd.n3830 gnd.t50 18.8012
R10258 gnd.n3815 gnd.t292 18.8012
R10259 gnd.n5387 gnd.t5 18.8012
R10260 gnd.n6351 gnd.t111 18.8012
R10261 gnd.n3674 gnd.n3673 18.4825
R10262 gnd.n7221 gnd.n7220 18.4247
R10263 gnd.n1222 gnd.n1218 18.4247
R10264 gnd.n7714 gnd.n124 18.2308
R10265 gnd.n6688 gnd.n6642 18.2308
R10266 gnd.n5751 gnd.n1163 18.2308
R10267 gnd.n4507 gnd.n4451 18.2308
R10268 gnd.t49 gnd.n3354 18.1639
R10269 gnd.n5601 gnd.n5399 17.8452
R10270 gnd.n6002 gnd.n963 17.8452
R10271 gnd.n6857 gnd.n860 17.8452
R10272 gnd.n6251 gnd.n836 17.8452
R10273 gnd.n6945 gnd.n775 17.8452
R10274 gnd.n6993 gnd.n726 17.8452
R10275 gnd.n3382 gnd.t15 17.5266
R10276 gnd.n7665 gnd.n232 17.5266
R10277 gnd.t167 gnd.n917 17.2079
R10278 gnd.t166 gnd.n799 17.2079
R10279 gnd.n3781 gnd.t322 16.8893
R10280 gnd.n6013 gnd.n953 16.5706
R10281 gnd.n6046 gnd.t338 16.5706
R10282 gnd.n6865 gnd.n852 16.5706
R10283 gnd.n6202 gnd.n844 16.5706
R10284 gnd.n6175 gnd.t336 16.5706
R10285 gnd.n6937 gnd.n783 16.5706
R10286 gnd.n3609 gnd.t251 16.2519
R10287 gnd.n3309 gnd.t45 16.2519
R10288 gnd.n6055 gnd.t113 15.9333
R10289 gnd.t118 gnd.n814 15.9333
R10290 gnd.n4296 gnd.n4294 15.6674
R10291 gnd.n4264 gnd.n4262 15.6674
R10292 gnd.n4232 gnd.n4230 15.6674
R10293 gnd.n4201 gnd.n4199 15.6674
R10294 gnd.n4169 gnd.n4167 15.6674
R10295 gnd.n4137 gnd.n4135 15.6674
R10296 gnd.n4105 gnd.n4103 15.6674
R10297 gnd.n4074 gnd.n4072 15.6674
R10298 gnd.n3600 gnd.t251 15.6146
R10299 gnd.t214 gnd.n1646 15.6146
R10300 gnd.n5924 gnd.n953 15.296
R10301 gnd.n6022 gnd.n6021 15.296
R10302 gnd.n893 gnd.t65 15.296
R10303 gnd.n6232 gnd.n852 15.296
R10304 gnd.n6873 gnd.n844 15.296
R10305 gnd.t330 gnd.n822 15.296
R10306 gnd.n6929 gnd.n791 15.296
R10307 gnd.n6159 gnd.n783 15.296
R10308 gnd.n6985 gnd.t203 15.296
R10309 gnd.n6411 gnd.n6410 15.0827
R10310 gnd.n5410 gnd.n5405 15.0481
R10311 gnd.n6421 gnd.n6420 15.0481
R10312 gnd.n3968 gnd.t13 14.9773
R10313 gnd.n6821 gnd.t331 14.6587
R10314 gnd.t329 gnd.n830 14.6587
R10315 gnd.n6977 gnd.t200 14.6587
R10316 gnd.t352 gnd.n3094 14.34
R10317 gnd.n4046 gnd.t33 14.34
R10318 gnd.n5620 gnd.t66 14.34
R10319 gnd.t295 gnd.n735 14.34
R10320 gnd.n7492 gnd.n232 14.34
R10321 gnd.n5962 gnd.n963 14.0214
R10322 gnd.n6069 gnd.n917 14.0214
R10323 gnd.n6223 gnd.t294 14.0214
R10324 gnd.n6215 gnd.n860 14.0214
R10325 gnd.n6881 gnd.n836 14.0214
R10326 gnd.t25 gnd.n838 14.0214
R10327 gnd.n6921 gnd.n799 14.0214
R10328 gnd.n6154 gnd.n775 14.0214
R10329 gnd.n6573 gnd.n726 14.0214
R10330 gnd.n3756 gnd.t174 13.7027
R10331 gnd.n3052 gnd.t51 13.7027
R10332 gnd.n6841 gnd.t359 13.7027
R10333 gnd.n6270 gnd.t100 13.7027
R10334 gnd.t143 gnd.n345 13.7027
R10335 gnd.n3466 gnd.n3465 13.5763
R10336 gnd.n4410 gnd.n1602 13.5763
R10337 gnd.n7183 gnd.n578 13.5763
R10338 gnd.n7766 gnd.n7765 13.5763
R10339 gnd.n4683 gnd.n4628 13.5763
R10340 gnd.n5675 gnd.n1259 13.5763
R10341 gnd.n3674 gnd.n3412 13.384
R10342 gnd.n6233 gnd.t332 13.384
R10343 gnd.t114 gnd.n846 13.384
R10344 gnd.n5421 gnd.n5402 13.1884
R10345 gnd.n5416 gnd.n5415 13.1884
R10346 gnd.n5415 gnd.n5414 13.1884
R10347 gnd.n6414 gnd.n6409 13.1884
R10348 gnd.n6415 gnd.n6414 13.1884
R10349 gnd.n5417 gnd.n5404 13.146
R10350 gnd.n5413 gnd.n5404 13.146
R10351 gnd.n6413 gnd.n6412 13.146
R10352 gnd.n6413 gnd.n6408 13.146
R10353 gnd.n4992 gnd.t128 13.0654
R10354 gnd.t53 gnd.n362 13.0654
R10355 gnd.n4297 gnd.n4293 12.8005
R10356 gnd.n4265 gnd.n4261 12.8005
R10357 gnd.n4233 gnd.n4229 12.8005
R10358 gnd.n4202 gnd.n4198 12.8005
R10359 gnd.n4170 gnd.n4166 12.8005
R10360 gnd.n4138 gnd.n4134 12.8005
R10361 gnd.n4106 gnd.n4102 12.8005
R10362 gnd.n4075 gnd.n4071 12.8005
R10363 gnd.n5890 gnd.n1018 12.7467
R10364 gnd.n5978 gnd.t245 12.7467
R10365 gnd.n5907 gnd.n971 12.7467
R10366 gnd.n6820 gnd.n868 12.7467
R10367 gnd.n6889 gnd.n828 12.7467
R10368 gnd.n6149 gnd.n767 12.7467
R10369 gnd.t238 gnd.n728 12.7467
R10370 gnd.n1536 gnd.t31 12.4281
R10371 gnd.n5034 gnd.t29 12.4281
R10372 gnd.n5318 gnd.t125 12.4281
R10373 gnd.t153 gnd.n1070 12.4281
R10374 gnd.n7041 gnd.t164 12.4281
R10375 gnd.n7293 gnd.t38 12.4281
R10376 gnd.t57 gnd.n405 12.4281
R10377 gnd.t135 gnd.n229 12.4281
R10378 gnd.n3465 gnd.n3460 12.4126
R10379 gnd.n4413 gnd.n4410 12.4126
R10380 gnd.n7179 gnd.n578 12.4126
R10381 gnd.n7765 gnd.n200 12.4126
R10382 gnd.n4679 gnd.n4628 12.4126
R10383 gnd.n5670 gnd.n1259 12.4126
R10384 gnd.n5594 gnd.n5422 12.1761
R10385 gnd.n6427 gnd.n6426 12.1761
R10386 gnd.n5077 gnd.n1196 12.1094
R10387 gnd.n5880 gnd.t211 12.1094
R10388 gnd.n7252 gnd.n532 12.1094
R10389 gnd.n4301 gnd.n4300 12.0247
R10390 gnd.n4269 gnd.n4268 12.0247
R10391 gnd.n4237 gnd.n4236 12.0247
R10392 gnd.n4206 gnd.n4205 12.0247
R10393 gnd.n4174 gnd.n4173 12.0247
R10394 gnd.n4142 gnd.n4141 12.0247
R10395 gnd.n4110 gnd.n4109 12.0247
R10396 gnd.n4079 gnd.n4078 12.0247
R10397 gnd.n1504 gnd.t79 11.7908
R10398 gnd.n5286 gnd.t29 11.7908
R10399 gnd.n5096 gnd.t125 11.7908
R10400 gnd.n7127 gnd.t38 11.7908
R10401 gnd.n7341 gnd.t57 11.7908
R10402 gnd.t55 gnd.n259 11.7908
R10403 gnd.n5899 gnd.n1010 11.4721
R10404 gnd.n5386 gnd.n979 11.4721
R10405 gnd.n6056 gnd.n6055 11.4721
R10406 gnd.n6827 gnd.n892 11.4721
R10407 gnd.n6897 gnd.n820 11.4721
R10408 gnd.n6905 gnd.n814 11.4721
R10409 gnd.n6145 gnd.n759 11.4721
R10410 gnd.n6360 gnd.n6140 11.4721
R10411 gnd.n4304 gnd.n4291 11.249
R10412 gnd.n4272 gnd.n4259 11.249
R10413 gnd.n4240 gnd.n4227 11.249
R10414 gnd.n4209 gnd.n4196 11.249
R10415 gnd.n4177 gnd.n4164 11.249
R10416 gnd.n4145 gnd.n4132 11.249
R10417 gnd.n4113 gnd.n4100 11.249
R10418 gnd.n4082 gnd.n4069 11.249
R10419 gnd.n3744 gnd.t174 11.1535
R10420 gnd.n4873 gnd.t69 11.1535
R10421 gnd.n5238 gnd.n1392 11.1535
R10422 gnd.n5254 gnd.t128 11.1535
R10423 gnd.n6046 gnd.t318 11.1535
R10424 gnd.n6175 gnd.t1 11.1535
R10425 gnd.n7425 gnd.t53 11.1535
R10426 gnd.n7565 gnd.n7564 11.1535
R10427 gnd.t84 gnd.n289 11.1535
R10428 gnd.n6498 gnd.n6391 10.6151
R10429 gnd.n6504 gnd.n6391 10.6151
R10430 gnd.n6507 gnd.n6506 10.6151
R10431 gnd.n6507 gnd.n6387 10.6151
R10432 gnd.n6513 gnd.n6387 10.6151
R10433 gnd.n6514 gnd.n6513 10.6151
R10434 gnd.n6515 gnd.n6514 10.6151
R10435 gnd.n6515 gnd.n6385 10.6151
R10436 gnd.n6521 gnd.n6385 10.6151
R10437 gnd.n6522 gnd.n6521 10.6151
R10438 gnd.n6523 gnd.n6522 10.6151
R10439 gnd.n6523 gnd.n6383 10.6151
R10440 gnd.n6529 gnd.n6383 10.6151
R10441 gnd.n6530 gnd.n6529 10.6151
R10442 gnd.n6531 gnd.n6530 10.6151
R10443 gnd.n6531 gnd.n6381 10.6151
R10444 gnd.n6537 gnd.n6381 10.6151
R10445 gnd.n6538 gnd.n6537 10.6151
R10446 gnd.n6539 gnd.n6538 10.6151
R10447 gnd.n6539 gnd.n6379 10.6151
R10448 gnd.n6545 gnd.n6379 10.6151
R10449 gnd.n6546 gnd.n6545 10.6151
R10450 gnd.n6547 gnd.n6546 10.6151
R10451 gnd.n6547 gnd.n6377 10.6151
R10452 gnd.n6553 gnd.n6377 10.6151
R10453 gnd.n6554 gnd.n6553 10.6151
R10454 gnd.n6555 gnd.n6554 10.6151
R10455 gnd.n6555 gnd.n6375 10.6151
R10456 gnd.n6561 gnd.n6375 10.6151
R10457 gnd.n6562 gnd.n6561 10.6151
R10458 gnd.n5463 gnd.n5462 10.6151
R10459 gnd.n5462 gnd.n5396 10.6151
R10460 gnd.n5604 gnd.n5396 10.6151
R10461 gnd.n5605 gnd.n5604 10.6151
R10462 gnd.n5607 gnd.n5605 10.6151
R10463 gnd.n5608 gnd.n5607 10.6151
R10464 gnd.n5610 gnd.n5608 10.6151
R10465 gnd.n5610 gnd.n5609 10.6151
R10466 gnd.n5609 gnd.n992 10.6151
R10467 gnd.n5976 gnd.n992 10.6151
R10468 gnd.n5976 gnd.n5975 10.6151
R10469 gnd.n5975 gnd.n5974 10.6151
R10470 gnd.n5974 gnd.n993 10.6151
R10471 gnd.n995 gnd.n993 10.6151
R10472 gnd.n5917 gnd.n995 10.6151
R10473 gnd.n5919 gnd.n5917 10.6151
R10474 gnd.n5920 gnd.n5919 10.6151
R10475 gnd.n5921 gnd.n5920 10.6151
R10476 gnd.n5922 gnd.n5921 10.6151
R10477 gnd.n5922 gnd.n5915 10.6151
R10478 gnd.n5937 gnd.n5915 10.6151
R10479 gnd.n5938 gnd.n5937 10.6151
R10480 gnd.n5941 gnd.n5938 10.6151
R10481 gnd.n5941 gnd.n5940 10.6151
R10482 gnd.n5940 gnd.n5939 10.6151
R10483 gnd.n5939 gnd.n938 10.6151
R10484 gnd.n938 gnd.n936 10.6151
R10485 gnd.n6036 gnd.n936 10.6151
R10486 gnd.n6037 gnd.n6036 10.6151
R10487 gnd.n6044 gnd.n6037 10.6151
R10488 gnd.n6044 gnd.n6043 10.6151
R10489 gnd.n6043 gnd.n6042 10.6151
R10490 gnd.n6042 gnd.n6038 10.6151
R10491 gnd.n6038 gnd.n889 10.6151
R10492 gnd.n6831 gnd.n889 10.6151
R10493 gnd.n6831 gnd.n6830 10.6151
R10494 gnd.n6830 gnd.n6829 10.6151
R10495 gnd.n6829 gnd.n890 10.6151
R10496 gnd.n6211 gnd.n890 10.6151
R10497 gnd.n6212 gnd.n6211 10.6151
R10498 gnd.n6213 gnd.n6212 10.6151
R10499 gnd.n6213 gnd.n6209 10.6151
R10500 gnd.n6226 gnd.n6209 10.6151
R10501 gnd.n6227 gnd.n6226 10.6151
R10502 gnd.n6230 gnd.n6227 10.6151
R10503 gnd.n6230 gnd.n6229 10.6151
R10504 gnd.n6229 gnd.n6228 10.6151
R10505 gnd.n6228 gnd.n6200 10.6151
R10506 gnd.n6245 gnd.n6200 10.6151
R10507 gnd.n6246 gnd.n6245 10.6151
R10508 gnd.n6249 gnd.n6246 10.6151
R10509 gnd.n6249 gnd.n6248 10.6151
R10510 gnd.n6248 gnd.n6247 10.6151
R10511 gnd.n6247 gnd.n6191 10.6151
R10512 gnd.n6264 gnd.n6191 10.6151
R10513 gnd.n6265 gnd.n6264 10.6151
R10514 gnd.n6268 gnd.n6265 10.6151
R10515 gnd.n6268 gnd.n6267 10.6151
R10516 gnd.n6267 gnd.n6266 10.6151
R10517 gnd.n6266 gnd.n6183 10.6151
R10518 gnd.n6283 gnd.n6183 10.6151
R10519 gnd.n6284 gnd.n6283 10.6151
R10520 gnd.n6287 gnd.n6284 10.6151
R10521 gnd.n6287 gnd.n6286 10.6151
R10522 gnd.n6286 gnd.n6285 10.6151
R10523 gnd.n6285 gnd.n6172 10.6151
R10524 gnd.n6301 gnd.n6172 10.6151
R10525 gnd.n6302 gnd.n6301 10.6151
R10526 gnd.n6305 gnd.n6302 10.6151
R10527 gnd.n6305 gnd.n6304 10.6151
R10528 gnd.n6304 gnd.n6303 10.6151
R10529 gnd.n6303 gnd.n6162 10.6151
R10530 gnd.n6319 gnd.n6162 10.6151
R10531 gnd.n6320 gnd.n6319 10.6151
R10532 gnd.n6323 gnd.n6320 10.6151
R10533 gnd.n6323 gnd.n6322 10.6151
R10534 gnd.n6322 gnd.n6321 10.6151
R10535 gnd.n6321 gnd.n6152 10.6151
R10536 gnd.n6337 gnd.n6152 10.6151
R10537 gnd.n6338 gnd.n6337 10.6151
R10538 gnd.n6340 gnd.n6338 10.6151
R10539 gnd.n6340 gnd.n6339 10.6151
R10540 gnd.n6339 gnd.n6143 10.6151
R10541 gnd.n6353 gnd.n6143 10.6151
R10542 gnd.n6354 gnd.n6353 10.6151
R10543 gnd.n6355 gnd.n6354 10.6151
R10544 gnd.n6358 gnd.n6355 10.6151
R10545 gnd.n6358 gnd.n6357 10.6151
R10546 gnd.n6357 gnd.n6356 10.6151
R10547 gnd.n6356 gnd.n6133 10.6151
R10548 gnd.n6370 gnd.n6133 10.6151
R10549 gnd.n6371 gnd.n6370 10.6151
R10550 gnd.n6373 gnd.n6371 10.6151
R10551 gnd.n6374 gnd.n6373 10.6151
R10552 gnd.n6563 gnd.n6374 10.6151
R10553 gnd.n5526 gnd.n5444 10.6151
R10554 gnd.n5526 gnd.n5525 10.6151
R10555 gnd.n5523 gnd.n5448 10.6151
R10556 gnd.n5517 gnd.n5448 10.6151
R10557 gnd.n5517 gnd.n5516 10.6151
R10558 gnd.n5516 gnd.n5515 10.6151
R10559 gnd.n5515 gnd.n5450 10.6151
R10560 gnd.n5509 gnd.n5450 10.6151
R10561 gnd.n5509 gnd.n5508 10.6151
R10562 gnd.n5508 gnd.n5507 10.6151
R10563 gnd.n5507 gnd.n5452 10.6151
R10564 gnd.n5501 gnd.n5452 10.6151
R10565 gnd.n5501 gnd.n5500 10.6151
R10566 gnd.n5500 gnd.n5499 10.6151
R10567 gnd.n5499 gnd.n5454 10.6151
R10568 gnd.n5493 gnd.n5454 10.6151
R10569 gnd.n5493 gnd.n5492 10.6151
R10570 gnd.n5492 gnd.n5491 10.6151
R10571 gnd.n5491 gnd.n5456 10.6151
R10572 gnd.n5485 gnd.n5456 10.6151
R10573 gnd.n5485 gnd.n5484 10.6151
R10574 gnd.n5484 gnd.n5483 10.6151
R10575 gnd.n5483 gnd.n5458 10.6151
R10576 gnd.n5477 gnd.n5458 10.6151
R10577 gnd.n5477 gnd.n5476 10.6151
R10578 gnd.n5476 gnd.n5475 10.6151
R10579 gnd.n5475 gnd.n5460 10.6151
R10580 gnd.n5469 gnd.n5460 10.6151
R10581 gnd.n5469 gnd.n5468 10.6151
R10582 gnd.n5468 gnd.n5467 10.6151
R10583 gnd.n5594 gnd.n5593 10.6151
R10584 gnd.n5593 gnd.n5424 10.6151
R10585 gnd.n5589 gnd.n5424 10.6151
R10586 gnd.n5589 gnd.n5588 10.6151
R10587 gnd.n5588 gnd.n5426 10.6151
R10588 gnd.n5583 gnd.n5426 10.6151
R10589 gnd.n5583 gnd.n5582 10.6151
R10590 gnd.n5582 gnd.n5581 10.6151
R10591 gnd.n5581 gnd.n5428 10.6151
R10592 gnd.n5575 gnd.n5428 10.6151
R10593 gnd.n5575 gnd.n5574 10.6151
R10594 gnd.n5574 gnd.n5573 10.6151
R10595 gnd.n5573 gnd.n5430 10.6151
R10596 gnd.n5567 gnd.n5430 10.6151
R10597 gnd.n5567 gnd.n5566 10.6151
R10598 gnd.n5566 gnd.n5565 10.6151
R10599 gnd.n5565 gnd.n5432 10.6151
R10600 gnd.n5559 gnd.n5432 10.6151
R10601 gnd.n5559 gnd.n5558 10.6151
R10602 gnd.n5558 gnd.n5557 10.6151
R10603 gnd.n5557 gnd.n5434 10.6151
R10604 gnd.n5551 gnd.n5434 10.6151
R10605 gnd.n5551 gnd.n5550 10.6151
R10606 gnd.n5550 gnd.n5549 10.6151
R10607 gnd.n5549 gnd.n5436 10.6151
R10608 gnd.n5543 gnd.n5436 10.6151
R10609 gnd.n5543 gnd.n5542 10.6151
R10610 gnd.n5542 gnd.n5541 10.6151
R10611 gnd.n5537 gnd.n5536 10.6151
R10612 gnd.n5536 gnd.n5442 10.6151
R10613 gnd.n6428 gnd.n6427 10.6151
R10614 gnd.n6433 gnd.n6428 10.6151
R10615 gnd.n6434 gnd.n6433 10.6151
R10616 gnd.n6435 gnd.n6434 10.6151
R10617 gnd.n6435 gnd.n6405 10.6151
R10618 gnd.n6441 gnd.n6405 10.6151
R10619 gnd.n6442 gnd.n6441 10.6151
R10620 gnd.n6443 gnd.n6442 10.6151
R10621 gnd.n6443 gnd.n6403 10.6151
R10622 gnd.n6449 gnd.n6403 10.6151
R10623 gnd.n6450 gnd.n6449 10.6151
R10624 gnd.n6451 gnd.n6450 10.6151
R10625 gnd.n6451 gnd.n6401 10.6151
R10626 gnd.n6457 gnd.n6401 10.6151
R10627 gnd.n6458 gnd.n6457 10.6151
R10628 gnd.n6459 gnd.n6458 10.6151
R10629 gnd.n6459 gnd.n6399 10.6151
R10630 gnd.n6465 gnd.n6399 10.6151
R10631 gnd.n6466 gnd.n6465 10.6151
R10632 gnd.n6467 gnd.n6466 10.6151
R10633 gnd.n6467 gnd.n6397 10.6151
R10634 gnd.n6473 gnd.n6397 10.6151
R10635 gnd.n6474 gnd.n6473 10.6151
R10636 gnd.n6475 gnd.n6474 10.6151
R10637 gnd.n6475 gnd.n6395 10.6151
R10638 gnd.n6481 gnd.n6395 10.6151
R10639 gnd.n6482 gnd.n6481 10.6151
R10640 gnd.n6486 gnd.n6482 10.6151
R10641 gnd.n6491 gnd.n6393 10.6151
R10642 gnd.n6492 gnd.n6491 10.6151
R10643 gnd.n5598 gnd.n5597 10.6151
R10644 gnd.n5599 gnd.n5598 10.6151
R10645 gnd.n5599 gnd.n5381 10.6151
R10646 gnd.n5618 gnd.n5381 10.6151
R10647 gnd.n5618 gnd.n5617 10.6151
R10648 gnd.n5617 gnd.n5616 10.6151
R10649 gnd.n5616 gnd.n5382 10.6151
R10650 gnd.n5392 gnd.n5382 10.6151
R10651 gnd.n5392 gnd.n5391 10.6151
R10652 gnd.n5391 gnd.n5390 10.6151
R10653 gnd.n5390 gnd.n5389 10.6151
R10654 gnd.n5389 gnd.n5384 10.6151
R10655 gnd.n5384 gnd.n998 10.6151
R10656 gnd.n5968 gnd.n998 10.6151
R10657 gnd.n5968 gnd.n5967 10.6151
R10658 gnd.n5967 gnd.n5966 10.6151
R10659 gnd.n5966 gnd.n999 10.6151
R10660 gnd.n5927 gnd.n999 10.6151
R10661 gnd.n5928 gnd.n5927 10.6151
R10662 gnd.n5932 gnd.n5928 10.6151
R10663 gnd.n5932 gnd.n5931 10.6151
R10664 gnd.n5931 gnd.n5930 10.6151
R10665 gnd.n5930 gnd.n943 10.6151
R10666 gnd.n6024 gnd.n943 10.6151
R10667 gnd.n6025 gnd.n6024 10.6151
R10668 gnd.n6030 gnd.n6025 10.6151
R10669 gnd.n6030 gnd.n6029 10.6151
R10670 gnd.n6029 gnd.n6028 10.6151
R10671 gnd.n6028 gnd.n6026 10.6151
R10672 gnd.n6026 gnd.n930 10.6151
R10673 gnd.n6049 gnd.n930 10.6151
R10674 gnd.n6050 gnd.n6049 10.6151
R10675 gnd.n6053 gnd.n6050 10.6151
R10676 gnd.n6053 gnd.n6052 10.6151
R10677 gnd.n6052 gnd.n6051 10.6151
R10678 gnd.n6051 gnd.n896 10.6151
R10679 gnd.n6825 gnd.n896 10.6151
R10680 gnd.n6825 gnd.n6824 10.6151
R10681 gnd.n6824 gnd.n6823 10.6151
R10682 gnd.n6823 gnd.n897 10.6151
R10683 gnd.n6218 gnd.n897 10.6151
R10684 gnd.n6221 gnd.n6218 10.6151
R10685 gnd.n6221 gnd.n6220 10.6151
R10686 gnd.n6220 gnd.n6219 10.6151
R10687 gnd.n6219 gnd.n6205 10.6151
R10688 gnd.n6236 gnd.n6205 10.6151
R10689 gnd.n6237 gnd.n6236 10.6151
R10690 gnd.n6240 gnd.n6237 10.6151
R10691 gnd.n6240 gnd.n6239 10.6151
R10692 gnd.n6239 gnd.n6238 10.6151
R10693 gnd.n6238 gnd.n6196 10.6151
R10694 gnd.n6255 gnd.n6196 10.6151
R10695 gnd.n6256 gnd.n6255 10.6151
R10696 gnd.n6259 gnd.n6256 10.6151
R10697 gnd.n6259 gnd.n6258 10.6151
R10698 gnd.n6258 gnd.n6257 10.6151
R10699 gnd.n6257 gnd.n6187 10.6151
R10700 gnd.n6274 gnd.n6187 10.6151
R10701 gnd.n6275 gnd.n6274 10.6151
R10702 gnd.n6278 gnd.n6275 10.6151
R10703 gnd.n6278 gnd.n6277 10.6151
R10704 gnd.n6277 gnd.n6276 10.6151
R10705 gnd.n6276 gnd.n6178 10.6151
R10706 gnd.n6292 gnd.n6178 10.6151
R10707 gnd.n6293 gnd.n6292 10.6151
R10708 gnd.n6296 gnd.n6293 10.6151
R10709 gnd.n6296 gnd.n6295 10.6151
R10710 gnd.n6295 gnd.n6294 10.6151
R10711 gnd.n6294 gnd.n6167 10.6151
R10712 gnd.n6310 gnd.n6167 10.6151
R10713 gnd.n6311 gnd.n6310 10.6151
R10714 gnd.n6314 gnd.n6311 10.6151
R10715 gnd.n6314 gnd.n6313 10.6151
R10716 gnd.n6313 gnd.n6312 10.6151
R10717 gnd.n6312 gnd.n6157 10.6151
R10718 gnd.n6328 gnd.n6157 10.6151
R10719 gnd.n6329 gnd.n6328 10.6151
R10720 gnd.n6332 gnd.n6329 10.6151
R10721 gnd.n6332 gnd.n6331 10.6151
R10722 gnd.n6331 gnd.n6330 10.6151
R10723 gnd.n6330 gnd.n6147 10.6151
R10724 gnd.n6345 gnd.n6147 10.6151
R10725 gnd.n6346 gnd.n6345 10.6151
R10726 gnd.n6349 gnd.n6346 10.6151
R10727 gnd.n6349 gnd.n6348 10.6151
R10728 gnd.n6348 gnd.n6347 10.6151
R10729 gnd.n6347 gnd.n6138 10.6151
R10730 gnd.n6363 gnd.n6138 10.6151
R10731 gnd.n6364 gnd.n6363 10.6151
R10732 gnd.n6365 gnd.n6364 10.6151
R10733 gnd.n6365 gnd.n6128 10.6151
R10734 gnd.n6570 gnd.n6128 10.6151
R10735 gnd.n6570 gnd.n6569 10.6151
R10736 gnd.n6569 gnd.n6568 10.6151
R10737 gnd.n6568 gnd.n6129 10.6151
R10738 gnd.n3663 gnd.t23 10.5161
R10739 gnd.n3096 gnd.t352 10.5161
R10740 gnd.n4029 gnd.t33 10.5161
R10741 gnd.n5232 gnd.t51 10.5161
R10742 gnd.n5944 gnd.t3 10.5161
R10743 gnd.n6164 gnd.t341 10.5161
R10744 gnd.n7555 gnd.t143 10.5161
R10745 gnd.n4305 gnd.n4289 10.4732
R10746 gnd.n4273 gnd.n4257 10.4732
R10747 gnd.n4241 gnd.n4225 10.4732
R10748 gnd.n4210 gnd.n4194 10.4732
R10749 gnd.n4178 gnd.n4162 10.4732
R10750 gnd.n4146 gnd.n4130 10.4732
R10751 gnd.n4114 gnd.n4098 10.4732
R10752 gnd.n4083 gnd.n4067 10.4732
R10753 gnd.n5899 gnd.n1011 10.1975
R10754 gnd.n6056 gnd.n883 10.1975
R10755 gnd.n893 gnd.n892 10.1975
R10756 gnd.n6897 gnd.n822 10.1975
R10757 gnd.n6905 gnd.n812 10.1975
R10758 gnd.n6140 gnd.n750 10.1975
R10759 gnd.t13 gnd.n3113 9.87883
R10760 gnd.n4879 gnd.t40 9.87883
R10761 gnd.n292 gnd.t42 9.87883
R10762 gnd.n7891 gnd.n78 9.81789
R10763 gnd.n4309 gnd.n4308 9.69747
R10764 gnd.n4277 gnd.n4276 9.69747
R10765 gnd.n4245 gnd.n4244 9.69747
R10766 gnd.n4214 gnd.n4213 9.69747
R10767 gnd.n4182 gnd.n4181 9.69747
R10768 gnd.n4150 gnd.n4149 9.69747
R10769 gnd.n4118 gnd.n4117 9.69747
R10770 gnd.n4087 gnd.n4086 9.69747
R10771 gnd.n5659 gnd.n5350 9.45751
R10772 gnd.n7256 gnd.n7255 9.45599
R10773 gnd.n4315 gnd.n4314 9.45567
R10774 gnd.n4283 gnd.n4282 9.45567
R10775 gnd.n4251 gnd.n4250 9.45567
R10776 gnd.n4220 gnd.n4219 9.45567
R10777 gnd.n4188 gnd.n4187 9.45567
R10778 gnd.n4156 gnd.n4155 9.45567
R10779 gnd.n4124 gnd.n4123 9.45567
R10780 gnd.n4093 gnd.n4092 9.45567
R10781 gnd.n3261 gnd.n3260 9.39724
R10782 gnd.n4314 gnd.n4313 9.3005
R10783 gnd.n4287 gnd.n4286 9.3005
R10784 gnd.n4308 gnd.n4307 9.3005
R10785 gnd.n4306 gnd.n4305 9.3005
R10786 gnd.n4291 gnd.n4290 9.3005
R10787 gnd.n4300 gnd.n4299 9.3005
R10788 gnd.n4298 gnd.n4297 9.3005
R10789 gnd.n4282 gnd.n4281 9.3005
R10790 gnd.n4255 gnd.n4254 9.3005
R10791 gnd.n4276 gnd.n4275 9.3005
R10792 gnd.n4274 gnd.n4273 9.3005
R10793 gnd.n4259 gnd.n4258 9.3005
R10794 gnd.n4268 gnd.n4267 9.3005
R10795 gnd.n4266 gnd.n4265 9.3005
R10796 gnd.n4250 gnd.n4249 9.3005
R10797 gnd.n4223 gnd.n4222 9.3005
R10798 gnd.n4244 gnd.n4243 9.3005
R10799 gnd.n4242 gnd.n4241 9.3005
R10800 gnd.n4227 gnd.n4226 9.3005
R10801 gnd.n4236 gnd.n4235 9.3005
R10802 gnd.n4234 gnd.n4233 9.3005
R10803 gnd.n4219 gnd.n4218 9.3005
R10804 gnd.n4192 gnd.n4191 9.3005
R10805 gnd.n4213 gnd.n4212 9.3005
R10806 gnd.n4211 gnd.n4210 9.3005
R10807 gnd.n4196 gnd.n4195 9.3005
R10808 gnd.n4205 gnd.n4204 9.3005
R10809 gnd.n4203 gnd.n4202 9.3005
R10810 gnd.n4187 gnd.n4186 9.3005
R10811 gnd.n4160 gnd.n4159 9.3005
R10812 gnd.n4181 gnd.n4180 9.3005
R10813 gnd.n4179 gnd.n4178 9.3005
R10814 gnd.n4164 gnd.n4163 9.3005
R10815 gnd.n4173 gnd.n4172 9.3005
R10816 gnd.n4171 gnd.n4170 9.3005
R10817 gnd.n4155 gnd.n4154 9.3005
R10818 gnd.n4128 gnd.n4127 9.3005
R10819 gnd.n4149 gnd.n4148 9.3005
R10820 gnd.n4147 gnd.n4146 9.3005
R10821 gnd.n4132 gnd.n4131 9.3005
R10822 gnd.n4141 gnd.n4140 9.3005
R10823 gnd.n4139 gnd.n4138 9.3005
R10824 gnd.n4123 gnd.n4122 9.3005
R10825 gnd.n4096 gnd.n4095 9.3005
R10826 gnd.n4117 gnd.n4116 9.3005
R10827 gnd.n4115 gnd.n4114 9.3005
R10828 gnd.n4100 gnd.n4099 9.3005
R10829 gnd.n4109 gnd.n4108 9.3005
R10830 gnd.n4107 gnd.n4106 9.3005
R10831 gnd.n4092 gnd.n4091 9.3005
R10832 gnd.n4065 gnd.n4064 9.3005
R10833 gnd.n4086 gnd.n4085 9.3005
R10834 gnd.n4084 gnd.n4083 9.3005
R10835 gnd.n4069 gnd.n4068 9.3005
R10836 gnd.n4078 gnd.n4077 9.3005
R10837 gnd.n4076 gnd.n4075 9.3005
R10838 gnd.n4440 gnd.n4439 9.3005
R10839 gnd.n4438 gnd.n1590 9.3005
R10840 gnd.n4437 gnd.n4436 9.3005
R10841 gnd.n4433 gnd.n1591 9.3005
R10842 gnd.n4430 gnd.n1592 9.3005
R10843 gnd.n4429 gnd.n1593 9.3005
R10844 gnd.n4426 gnd.n1594 9.3005
R10845 gnd.n4425 gnd.n1595 9.3005
R10846 gnd.n4422 gnd.n1596 9.3005
R10847 gnd.n4421 gnd.n1597 9.3005
R10848 gnd.n4418 gnd.n1598 9.3005
R10849 gnd.n4417 gnd.n1599 9.3005
R10850 gnd.n4414 gnd.n1600 9.3005
R10851 gnd.n4413 gnd.n1601 9.3005
R10852 gnd.n4410 gnd.n4409 9.3005
R10853 gnd.n4408 gnd.n1602 9.3005
R10854 gnd.n4441 gnd.n1589 9.3005
R10855 gnd.n3682 gnd.n3681 9.3005
R10856 gnd.n3386 gnd.n3385 9.3005
R10857 gnd.n3709 gnd.n3708 9.3005
R10858 gnd.n3710 gnd.n3384 9.3005
R10859 gnd.n3714 gnd.n3711 9.3005
R10860 gnd.n3713 gnd.n3712 9.3005
R10861 gnd.n3358 gnd.n3357 9.3005
R10862 gnd.n3739 gnd.n3738 9.3005
R10863 gnd.n3740 gnd.n3356 9.3005
R10864 gnd.n3742 gnd.n3741 9.3005
R10865 gnd.n3336 gnd.n3335 9.3005
R10866 gnd.n3770 gnd.n3769 9.3005
R10867 gnd.n3771 gnd.n3334 9.3005
R10868 gnd.n3779 gnd.n3772 9.3005
R10869 gnd.n3778 gnd.n3773 9.3005
R10870 gnd.n3777 gnd.n3775 9.3005
R10871 gnd.n3774 gnd.n3283 9.3005
R10872 gnd.n3827 gnd.n3284 9.3005
R10873 gnd.n3826 gnd.n3285 9.3005
R10874 gnd.n3825 gnd.n3286 9.3005
R10875 gnd.n3305 gnd.n3287 9.3005
R10876 gnd.n3307 gnd.n3306 9.3005
R10877 gnd.n3193 gnd.n3192 9.3005
R10878 gnd.n3865 gnd.n3864 9.3005
R10879 gnd.n3866 gnd.n3191 9.3005
R10880 gnd.n3870 gnd.n3867 9.3005
R10881 gnd.n3869 gnd.n3868 9.3005
R10882 gnd.n3166 gnd.n3165 9.3005
R10883 gnd.n3905 gnd.n3904 9.3005
R10884 gnd.n3906 gnd.n3164 9.3005
R10885 gnd.n3910 gnd.n3907 9.3005
R10886 gnd.n3909 gnd.n3908 9.3005
R10887 gnd.n3139 gnd.n3138 9.3005
R10888 gnd.n3950 gnd.n3949 9.3005
R10889 gnd.n3951 gnd.n3137 9.3005
R10890 gnd.n3955 gnd.n3952 9.3005
R10891 gnd.n3954 gnd.n3953 9.3005
R10892 gnd.n3111 gnd.n3110 9.3005
R10893 gnd.n3990 gnd.n3989 9.3005
R10894 gnd.n3991 gnd.n3109 9.3005
R10895 gnd.n3995 gnd.n3992 9.3005
R10896 gnd.n3994 gnd.n3993 9.3005
R10897 gnd.n3084 gnd.n3083 9.3005
R10898 gnd.n4039 gnd.n4038 9.3005
R10899 gnd.n4040 gnd.n3082 9.3005
R10900 gnd.n4044 gnd.n4041 9.3005
R10901 gnd.n4043 gnd.n4042 9.3005
R10902 gnd.n1651 gnd.n1650 9.3005
R10903 gnd.n4333 gnd.n4332 9.3005
R10904 gnd.n4334 gnd.n1649 9.3005
R10905 gnd.n4340 gnd.n4335 9.3005
R10906 gnd.n4339 gnd.n4336 9.3005
R10907 gnd.n4338 gnd.n4337 9.3005
R10908 gnd.n3683 gnd.n3680 9.3005
R10909 gnd.n3465 gnd.n3424 9.3005
R10910 gnd.n3460 gnd.n3459 9.3005
R10911 gnd.n3458 gnd.n3425 9.3005
R10912 gnd.n3457 gnd.n3456 9.3005
R10913 gnd.n3453 gnd.n3426 9.3005
R10914 gnd.n3450 gnd.n3449 9.3005
R10915 gnd.n3448 gnd.n3427 9.3005
R10916 gnd.n3447 gnd.n3446 9.3005
R10917 gnd.n3443 gnd.n3428 9.3005
R10918 gnd.n3440 gnd.n3439 9.3005
R10919 gnd.n3438 gnd.n3429 9.3005
R10920 gnd.n3437 gnd.n3436 9.3005
R10921 gnd.n3433 gnd.n3431 9.3005
R10922 gnd.n3430 gnd.n3410 9.3005
R10923 gnd.n3677 gnd.n3409 9.3005
R10924 gnd.n3679 gnd.n3678 9.3005
R10925 gnd.n3467 gnd.n3466 9.3005
R10926 gnd.n3690 gnd.n3396 9.3005
R10927 gnd.n3697 gnd.n3397 9.3005
R10928 gnd.n3699 gnd.n3698 9.3005
R10929 gnd.n3700 gnd.n3377 9.3005
R10930 gnd.n3719 gnd.n3718 9.3005
R10931 gnd.n3721 gnd.n3369 9.3005
R10932 gnd.n3728 gnd.n3371 9.3005
R10933 gnd.n3729 gnd.n3366 9.3005
R10934 gnd.n3731 gnd.n3730 9.3005
R10935 gnd.n3367 gnd.n3352 9.3005
R10936 gnd.n3747 gnd.n3350 9.3005
R10937 gnd.n3751 gnd.n3750 9.3005
R10938 gnd.n3749 gnd.n3326 9.3005
R10939 gnd.n3786 gnd.n3325 9.3005
R10940 gnd.n3789 gnd.n3788 9.3005
R10941 gnd.n3322 gnd.n3321 9.3005
R10942 gnd.n3795 gnd.n3323 9.3005
R10943 gnd.n3797 gnd.n3796 9.3005
R10944 gnd.n3799 gnd.n3320 9.3005
R10945 gnd.n3802 gnd.n3801 9.3005
R10946 gnd.n3805 gnd.n3803 9.3005
R10947 gnd.n3807 gnd.n3806 9.3005
R10948 gnd.n3813 gnd.n3808 9.3005
R10949 gnd.n3812 gnd.n3811 9.3005
R10950 gnd.n3184 gnd.n3183 9.3005
R10951 gnd.n3879 gnd.n3878 9.3005
R10952 gnd.n3880 gnd.n3177 9.3005
R10953 gnd.n3888 gnd.n3176 9.3005
R10954 gnd.n3891 gnd.n3890 9.3005
R10955 gnd.n3893 gnd.n3892 9.3005
R10956 gnd.n3896 gnd.n3159 9.3005
R10957 gnd.n3894 gnd.n3157 9.3005
R10958 gnd.n3916 gnd.n3155 9.3005
R10959 gnd.n3918 gnd.n3917 9.3005
R10960 gnd.n3129 gnd.n3128 9.3005
R10961 gnd.n3964 gnd.n3963 9.3005
R10962 gnd.n3965 gnd.n3122 9.3005
R10963 gnd.n3973 gnd.n3121 9.3005
R10964 gnd.n3976 gnd.n3975 9.3005
R10965 gnd.n3978 gnd.n3977 9.3005
R10966 gnd.n3981 gnd.n3104 9.3005
R10967 gnd.n3979 gnd.n3102 9.3005
R10968 gnd.n4001 gnd.n3100 9.3005
R10969 gnd.n4003 gnd.n4002 9.3005
R10970 gnd.n3075 gnd.n3074 9.3005
R10971 gnd.n4053 gnd.n4052 9.3005
R10972 gnd.n4054 gnd.n3068 9.3005
R10973 gnd.n4062 gnd.n3067 9.3005
R10974 gnd.n4321 gnd.n4320 9.3005
R10975 gnd.n4323 gnd.n4322 9.3005
R10976 gnd.n4324 gnd.n1642 9.3005
R10977 gnd.n4348 gnd.n4347 9.3005
R10978 gnd.n1643 gnd.n1605 9.3005
R10979 gnd.n3688 gnd.n3687 9.3005
R10980 gnd.n4404 gnd.n1606 9.3005
R10981 gnd.n4403 gnd.n1608 9.3005
R10982 gnd.n4400 gnd.n1609 9.3005
R10983 gnd.n4399 gnd.n1610 9.3005
R10984 gnd.n4396 gnd.n1611 9.3005
R10985 gnd.n4395 gnd.n1612 9.3005
R10986 gnd.n4392 gnd.n1613 9.3005
R10987 gnd.n4391 gnd.n1614 9.3005
R10988 gnd.n4388 gnd.n1615 9.3005
R10989 gnd.n4387 gnd.n1616 9.3005
R10990 gnd.n4384 gnd.n1617 9.3005
R10991 gnd.n4383 gnd.n1618 9.3005
R10992 gnd.n4380 gnd.n1619 9.3005
R10993 gnd.n4379 gnd.n1620 9.3005
R10994 gnd.n4376 gnd.n1621 9.3005
R10995 gnd.n4375 gnd.n1622 9.3005
R10996 gnd.n4372 gnd.n1623 9.3005
R10997 gnd.n4371 gnd.n1624 9.3005
R10998 gnd.n4368 gnd.n1625 9.3005
R10999 gnd.n4367 gnd.n1626 9.3005
R11000 gnd.n4364 gnd.n1627 9.3005
R11001 gnd.n4363 gnd.n1628 9.3005
R11002 gnd.n4360 gnd.n1632 9.3005
R11003 gnd.n4359 gnd.n1633 9.3005
R11004 gnd.n4356 gnd.n1634 9.3005
R11005 gnd.n4355 gnd.n1635 9.3005
R11006 gnd.n4406 gnd.n4405 9.3005
R11007 gnd.n3857 gnd.n3841 9.3005
R11008 gnd.n3856 gnd.n3842 9.3005
R11009 gnd.n3855 gnd.n3843 9.3005
R11010 gnd.n3853 gnd.n3844 9.3005
R11011 gnd.n3852 gnd.n3845 9.3005
R11012 gnd.n3850 gnd.n3846 9.3005
R11013 gnd.n3849 gnd.n3847 9.3005
R11014 gnd.n3147 gnd.n3146 9.3005
R11015 gnd.n3926 gnd.n3925 9.3005
R11016 gnd.n3927 gnd.n3145 9.3005
R11017 gnd.n3944 gnd.n3928 9.3005
R11018 gnd.n3943 gnd.n3929 9.3005
R11019 gnd.n3942 gnd.n3930 9.3005
R11020 gnd.n3940 gnd.n3931 9.3005
R11021 gnd.n3939 gnd.n3932 9.3005
R11022 gnd.n3937 gnd.n3933 9.3005
R11023 gnd.n3936 gnd.n3934 9.3005
R11024 gnd.n3091 gnd.n3090 9.3005
R11025 gnd.n4011 gnd.n4010 9.3005
R11026 gnd.n4012 gnd.n3089 9.3005
R11027 gnd.n4033 gnd.n4013 9.3005
R11028 gnd.n4032 gnd.n4014 9.3005
R11029 gnd.n4031 gnd.n4015 9.3005
R11030 gnd.n4028 gnd.n4016 9.3005
R11031 gnd.n4027 gnd.n4017 9.3005
R11032 gnd.n4025 gnd.n4018 9.3005
R11033 gnd.n4024 gnd.n4019 9.3005
R11034 gnd.n4022 gnd.n4021 9.3005
R11035 gnd.n4020 gnd.n1637 9.3005
R11036 gnd.n3598 gnd.n3597 9.3005
R11037 gnd.n3488 gnd.n3487 9.3005
R11038 gnd.n3612 gnd.n3611 9.3005
R11039 gnd.n3613 gnd.n3486 9.3005
R11040 gnd.n3615 gnd.n3614 9.3005
R11041 gnd.n3476 gnd.n3475 9.3005
R11042 gnd.n3628 gnd.n3627 9.3005
R11043 gnd.n3629 gnd.n3474 9.3005
R11044 gnd.n3661 gnd.n3630 9.3005
R11045 gnd.n3660 gnd.n3631 9.3005
R11046 gnd.n3659 gnd.n3632 9.3005
R11047 gnd.n3658 gnd.n3633 9.3005
R11048 gnd.n3655 gnd.n3634 9.3005
R11049 gnd.n3654 gnd.n3635 9.3005
R11050 gnd.n3653 gnd.n3636 9.3005
R11051 gnd.n3651 gnd.n3637 9.3005
R11052 gnd.n3650 gnd.n3638 9.3005
R11053 gnd.n3647 gnd.n3639 9.3005
R11054 gnd.n3646 gnd.n3640 9.3005
R11055 gnd.n3645 gnd.n3641 9.3005
R11056 gnd.n3643 gnd.n3642 9.3005
R11057 gnd.n3342 gnd.n3341 9.3005
R11058 gnd.n3759 gnd.n3758 9.3005
R11059 gnd.n3760 gnd.n3340 9.3005
R11060 gnd.n3764 gnd.n3761 9.3005
R11061 gnd.n3763 gnd.n3762 9.3005
R11062 gnd.n3264 gnd.n3263 9.3005
R11063 gnd.n3839 gnd.n3838 9.3005
R11064 gnd.n3596 gnd.n3497 9.3005
R11065 gnd.n3499 gnd.n3498 9.3005
R11066 gnd.n3543 gnd.n3541 9.3005
R11067 gnd.n3544 gnd.n3540 9.3005
R11068 gnd.n3547 gnd.n3536 9.3005
R11069 gnd.n3548 gnd.n3535 9.3005
R11070 gnd.n3551 gnd.n3534 9.3005
R11071 gnd.n3552 gnd.n3533 9.3005
R11072 gnd.n3555 gnd.n3532 9.3005
R11073 gnd.n3556 gnd.n3531 9.3005
R11074 gnd.n3559 gnd.n3530 9.3005
R11075 gnd.n3560 gnd.n3529 9.3005
R11076 gnd.n3563 gnd.n3528 9.3005
R11077 gnd.n3564 gnd.n3527 9.3005
R11078 gnd.n3567 gnd.n3526 9.3005
R11079 gnd.n3568 gnd.n3525 9.3005
R11080 gnd.n3571 gnd.n3524 9.3005
R11081 gnd.n3572 gnd.n3523 9.3005
R11082 gnd.n3575 gnd.n3522 9.3005
R11083 gnd.n3576 gnd.n3521 9.3005
R11084 gnd.n3579 gnd.n3520 9.3005
R11085 gnd.n3580 gnd.n3519 9.3005
R11086 gnd.n3583 gnd.n3518 9.3005
R11087 gnd.n3585 gnd.n3517 9.3005
R11088 gnd.n3586 gnd.n3516 9.3005
R11089 gnd.n3587 gnd.n3515 9.3005
R11090 gnd.n3588 gnd.n3514 9.3005
R11091 gnd.n3595 gnd.n3594 9.3005
R11092 gnd.n3604 gnd.n3603 9.3005
R11093 gnd.n3605 gnd.n3491 9.3005
R11094 gnd.n3607 gnd.n3606 9.3005
R11095 gnd.n3482 gnd.n3481 9.3005
R11096 gnd.n3620 gnd.n3619 9.3005
R11097 gnd.n3621 gnd.n3480 9.3005
R11098 gnd.n3623 gnd.n3622 9.3005
R11099 gnd.n3469 gnd.n3468 9.3005
R11100 gnd.n3666 gnd.n3665 9.3005
R11101 gnd.n3667 gnd.n3423 9.3005
R11102 gnd.n3671 gnd.n3669 9.3005
R11103 gnd.n3670 gnd.n3402 9.3005
R11104 gnd.n3689 gnd.n3401 9.3005
R11105 gnd.n3692 gnd.n3691 9.3005
R11106 gnd.n3395 gnd.n3394 9.3005
R11107 gnd.n3703 gnd.n3701 9.3005
R11108 gnd.n3702 gnd.n3376 9.3005
R11109 gnd.n3720 gnd.n3375 9.3005
R11110 gnd.n3723 gnd.n3722 9.3005
R11111 gnd.n3370 gnd.n3365 9.3005
R11112 gnd.n3733 gnd.n3732 9.3005
R11113 gnd.n3368 gnd.n3348 9.3005
R11114 gnd.n3754 gnd.n3349 9.3005
R11115 gnd.n3753 gnd.n3752 9.3005
R11116 gnd.n3351 gnd.n3327 9.3005
R11117 gnd.n3785 gnd.n3784 9.3005
R11118 gnd.n3787 gnd.n3272 9.3005
R11119 gnd.n3834 gnd.n3273 9.3005
R11120 gnd.n3833 gnd.n3274 9.3005
R11121 gnd.n3832 gnd.n3275 9.3005
R11122 gnd.n3798 gnd.n3276 9.3005
R11123 gnd.n3800 gnd.n3294 9.3005
R11124 gnd.n3820 gnd.n3295 9.3005
R11125 gnd.n3819 gnd.n3296 9.3005
R11126 gnd.n3818 gnd.n3297 9.3005
R11127 gnd.n3809 gnd.n3298 9.3005
R11128 gnd.n3810 gnd.n3185 9.3005
R11129 gnd.n3876 gnd.n3875 9.3005
R11130 gnd.n3877 gnd.n3178 9.3005
R11131 gnd.n3887 gnd.n3886 9.3005
R11132 gnd.n3889 gnd.n3174 9.3005
R11133 gnd.n3899 gnd.n3175 9.3005
R11134 gnd.n3898 gnd.n3897 9.3005
R11135 gnd.n3895 gnd.n3153 9.3005
R11136 gnd.n3921 gnd.n3154 9.3005
R11137 gnd.n3920 gnd.n3919 9.3005
R11138 gnd.n3156 gnd.n3130 9.3005
R11139 gnd.n3961 gnd.n3960 9.3005
R11140 gnd.n3962 gnd.n3123 9.3005
R11141 gnd.n3972 gnd.n3971 9.3005
R11142 gnd.n3974 gnd.n3119 9.3005
R11143 gnd.n3984 gnd.n3120 9.3005
R11144 gnd.n3983 gnd.n3982 9.3005
R11145 gnd.n3980 gnd.n3098 9.3005
R11146 gnd.n4006 gnd.n3099 9.3005
R11147 gnd.n4005 gnd.n4004 9.3005
R11148 gnd.n3101 gnd.n3076 9.3005
R11149 gnd.n4050 gnd.n4049 9.3005
R11150 gnd.n4051 gnd.n3069 9.3005
R11151 gnd.n4061 gnd.n4060 9.3005
R11152 gnd.n4319 gnd.n3065 9.3005
R11153 gnd.n4327 gnd.n3066 9.3005
R11154 gnd.n4326 gnd.n4325 9.3005
R11155 gnd.n1641 gnd.n1640 9.3005
R11156 gnd.n4350 gnd.n4349 9.3005
R11157 gnd.n3493 gnd.n3492 9.3005
R11158 gnd.n2841 gnd.n2840 9.3005
R11159 gnd.n2839 gnd.n1785 9.3005
R11160 gnd.n2838 gnd.n2837 9.3005
R11161 gnd.n1787 gnd.n1786 9.3005
R11162 gnd.n2831 gnd.n1791 9.3005
R11163 gnd.n2830 gnd.n1792 9.3005
R11164 gnd.n2829 gnd.n1793 9.3005
R11165 gnd.n1798 gnd.n1794 9.3005
R11166 gnd.n2823 gnd.n1799 9.3005
R11167 gnd.n2822 gnd.n1800 9.3005
R11168 gnd.n2821 gnd.n1801 9.3005
R11169 gnd.n1806 gnd.n1802 9.3005
R11170 gnd.n2815 gnd.n1807 9.3005
R11171 gnd.n2814 gnd.n1808 9.3005
R11172 gnd.n2813 gnd.n1809 9.3005
R11173 gnd.n1814 gnd.n1810 9.3005
R11174 gnd.n2807 gnd.n1815 9.3005
R11175 gnd.n2806 gnd.n1816 9.3005
R11176 gnd.n2805 gnd.n1817 9.3005
R11177 gnd.n1822 gnd.n1818 9.3005
R11178 gnd.n2799 gnd.n1823 9.3005
R11179 gnd.n2798 gnd.n1824 9.3005
R11180 gnd.n2797 gnd.n1825 9.3005
R11181 gnd.n1830 gnd.n1826 9.3005
R11182 gnd.n2791 gnd.n1831 9.3005
R11183 gnd.n2790 gnd.n1832 9.3005
R11184 gnd.n2789 gnd.n1833 9.3005
R11185 gnd.n1838 gnd.n1834 9.3005
R11186 gnd.n2783 gnd.n1839 9.3005
R11187 gnd.n2782 gnd.n1840 9.3005
R11188 gnd.n2781 gnd.n1841 9.3005
R11189 gnd.n1846 gnd.n1842 9.3005
R11190 gnd.n2775 gnd.n1847 9.3005
R11191 gnd.n2774 gnd.n1848 9.3005
R11192 gnd.n2773 gnd.n1849 9.3005
R11193 gnd.n1854 gnd.n1850 9.3005
R11194 gnd.n2767 gnd.n1855 9.3005
R11195 gnd.n2766 gnd.n1856 9.3005
R11196 gnd.n2765 gnd.n1857 9.3005
R11197 gnd.n1862 gnd.n1858 9.3005
R11198 gnd.n2759 gnd.n1863 9.3005
R11199 gnd.n2758 gnd.n1864 9.3005
R11200 gnd.n2757 gnd.n1865 9.3005
R11201 gnd.n1870 gnd.n1866 9.3005
R11202 gnd.n2751 gnd.n1871 9.3005
R11203 gnd.n2750 gnd.n1872 9.3005
R11204 gnd.n2749 gnd.n1873 9.3005
R11205 gnd.n1878 gnd.n1874 9.3005
R11206 gnd.n2743 gnd.n1879 9.3005
R11207 gnd.n2742 gnd.n1880 9.3005
R11208 gnd.n2741 gnd.n1881 9.3005
R11209 gnd.n1886 gnd.n1882 9.3005
R11210 gnd.n2735 gnd.n1887 9.3005
R11211 gnd.n2734 gnd.n1888 9.3005
R11212 gnd.n2733 gnd.n1889 9.3005
R11213 gnd.n1894 gnd.n1890 9.3005
R11214 gnd.n2727 gnd.n1895 9.3005
R11215 gnd.n2726 gnd.n1896 9.3005
R11216 gnd.n2725 gnd.n1897 9.3005
R11217 gnd.n1902 gnd.n1898 9.3005
R11218 gnd.n2719 gnd.n1903 9.3005
R11219 gnd.n2718 gnd.n1904 9.3005
R11220 gnd.n2717 gnd.n1905 9.3005
R11221 gnd.n1910 gnd.n1906 9.3005
R11222 gnd.n2711 gnd.n1911 9.3005
R11223 gnd.n2710 gnd.n1912 9.3005
R11224 gnd.n2709 gnd.n1913 9.3005
R11225 gnd.n1918 gnd.n1914 9.3005
R11226 gnd.n2703 gnd.n1919 9.3005
R11227 gnd.n2702 gnd.n1920 9.3005
R11228 gnd.n2701 gnd.n1921 9.3005
R11229 gnd.n1926 gnd.n1922 9.3005
R11230 gnd.n2695 gnd.n1927 9.3005
R11231 gnd.n2694 gnd.n1928 9.3005
R11232 gnd.n2693 gnd.n1929 9.3005
R11233 gnd.n1934 gnd.n1930 9.3005
R11234 gnd.n2687 gnd.n1935 9.3005
R11235 gnd.n2686 gnd.n1936 9.3005
R11236 gnd.n2685 gnd.n1937 9.3005
R11237 gnd.n1942 gnd.n1938 9.3005
R11238 gnd.n2679 gnd.n1943 9.3005
R11239 gnd.n2678 gnd.n1944 9.3005
R11240 gnd.n2677 gnd.n1945 9.3005
R11241 gnd.n1950 gnd.n1946 9.3005
R11242 gnd.n2671 gnd.n1951 9.3005
R11243 gnd.n2670 gnd.n1952 9.3005
R11244 gnd.n2669 gnd.n1953 9.3005
R11245 gnd.n1958 gnd.n1954 9.3005
R11246 gnd.n2663 gnd.n1959 9.3005
R11247 gnd.n2662 gnd.n1960 9.3005
R11248 gnd.n2661 gnd.n1961 9.3005
R11249 gnd.n1966 gnd.n1962 9.3005
R11250 gnd.n2655 gnd.n1967 9.3005
R11251 gnd.n2654 gnd.n1968 9.3005
R11252 gnd.n2653 gnd.n1969 9.3005
R11253 gnd.n1974 gnd.n1970 9.3005
R11254 gnd.n2647 gnd.n1975 9.3005
R11255 gnd.n2646 gnd.n1976 9.3005
R11256 gnd.n2645 gnd.n1977 9.3005
R11257 gnd.n1982 gnd.n1978 9.3005
R11258 gnd.n2639 gnd.n1983 9.3005
R11259 gnd.n2638 gnd.n1984 9.3005
R11260 gnd.n2637 gnd.n1985 9.3005
R11261 gnd.n1990 gnd.n1986 9.3005
R11262 gnd.n2631 gnd.n1991 9.3005
R11263 gnd.n2630 gnd.n1992 9.3005
R11264 gnd.n2629 gnd.n1993 9.3005
R11265 gnd.n1998 gnd.n1994 9.3005
R11266 gnd.n2623 gnd.n1999 9.3005
R11267 gnd.n2622 gnd.n2000 9.3005
R11268 gnd.n2621 gnd.n2001 9.3005
R11269 gnd.n2006 gnd.n2002 9.3005
R11270 gnd.n2615 gnd.n2007 9.3005
R11271 gnd.n2614 gnd.n2008 9.3005
R11272 gnd.n2613 gnd.n2009 9.3005
R11273 gnd.n2014 gnd.n2010 9.3005
R11274 gnd.n2607 gnd.n2015 9.3005
R11275 gnd.n2606 gnd.n2016 9.3005
R11276 gnd.n2605 gnd.n2017 9.3005
R11277 gnd.n2022 gnd.n2018 9.3005
R11278 gnd.n2599 gnd.n2023 9.3005
R11279 gnd.n2598 gnd.n2024 9.3005
R11280 gnd.n2597 gnd.n2025 9.3005
R11281 gnd.n2030 gnd.n2026 9.3005
R11282 gnd.n2591 gnd.n2031 9.3005
R11283 gnd.n2590 gnd.n2032 9.3005
R11284 gnd.n2589 gnd.n2033 9.3005
R11285 gnd.n2038 gnd.n2034 9.3005
R11286 gnd.n2583 gnd.n2039 9.3005
R11287 gnd.n2582 gnd.n2040 9.3005
R11288 gnd.n2581 gnd.n2041 9.3005
R11289 gnd.n2046 gnd.n2042 9.3005
R11290 gnd.n2575 gnd.n2047 9.3005
R11291 gnd.n2574 gnd.n2048 9.3005
R11292 gnd.n2573 gnd.n2049 9.3005
R11293 gnd.n2054 gnd.n2050 9.3005
R11294 gnd.n2567 gnd.n2055 9.3005
R11295 gnd.n2566 gnd.n2056 9.3005
R11296 gnd.n2565 gnd.n2057 9.3005
R11297 gnd.n2062 gnd.n2058 9.3005
R11298 gnd.n2559 gnd.n2063 9.3005
R11299 gnd.n2558 gnd.n2064 9.3005
R11300 gnd.n2557 gnd.n2065 9.3005
R11301 gnd.n2070 gnd.n2066 9.3005
R11302 gnd.n2551 gnd.n2071 9.3005
R11303 gnd.n2550 gnd.n2072 9.3005
R11304 gnd.n2549 gnd.n2073 9.3005
R11305 gnd.n2078 gnd.n2074 9.3005
R11306 gnd.n2543 gnd.n2079 9.3005
R11307 gnd.n2542 gnd.n2080 9.3005
R11308 gnd.n2541 gnd.n2081 9.3005
R11309 gnd.n2086 gnd.n2082 9.3005
R11310 gnd.n2535 gnd.n2087 9.3005
R11311 gnd.n2534 gnd.n2088 9.3005
R11312 gnd.n2533 gnd.n2089 9.3005
R11313 gnd.n2094 gnd.n2090 9.3005
R11314 gnd.n2527 gnd.n2095 9.3005
R11315 gnd.n2526 gnd.n2096 9.3005
R11316 gnd.n2525 gnd.n2097 9.3005
R11317 gnd.n2102 gnd.n2098 9.3005
R11318 gnd.n2519 gnd.n2103 9.3005
R11319 gnd.n2518 gnd.n2104 9.3005
R11320 gnd.n2517 gnd.n2105 9.3005
R11321 gnd.n2110 gnd.n2106 9.3005
R11322 gnd.n2511 gnd.n2111 9.3005
R11323 gnd.n2510 gnd.n2112 9.3005
R11324 gnd.n2509 gnd.n2113 9.3005
R11325 gnd.n2118 gnd.n2114 9.3005
R11326 gnd.n2503 gnd.n2119 9.3005
R11327 gnd.n2502 gnd.n2120 9.3005
R11328 gnd.n2501 gnd.n2121 9.3005
R11329 gnd.n2126 gnd.n2122 9.3005
R11330 gnd.n2495 gnd.n2127 9.3005
R11331 gnd.n2494 gnd.n2128 9.3005
R11332 gnd.n2493 gnd.n2129 9.3005
R11333 gnd.n2134 gnd.n2130 9.3005
R11334 gnd.n2487 gnd.n2135 9.3005
R11335 gnd.n2486 gnd.n2136 9.3005
R11336 gnd.n2485 gnd.n2137 9.3005
R11337 gnd.n2142 gnd.n2138 9.3005
R11338 gnd.n2479 gnd.n2143 9.3005
R11339 gnd.n2478 gnd.n2477 9.3005
R11340 gnd.n2145 gnd.n2144 9.3005
R11341 gnd.n2469 gnd.n2149 9.3005
R11342 gnd.n2468 gnd.n2150 9.3005
R11343 gnd.n2467 gnd.n2151 9.3005
R11344 gnd.n2156 gnd.n2152 9.3005
R11345 gnd.n2461 gnd.n2157 9.3005
R11346 gnd.n2460 gnd.n2158 9.3005
R11347 gnd.n2459 gnd.n2159 9.3005
R11348 gnd.n2164 gnd.n2160 9.3005
R11349 gnd.n2453 gnd.n2165 9.3005
R11350 gnd.n2452 gnd.n2166 9.3005
R11351 gnd.n2451 gnd.n2167 9.3005
R11352 gnd.n2172 gnd.n2168 9.3005
R11353 gnd.n2445 gnd.n2173 9.3005
R11354 gnd.n2444 gnd.n2174 9.3005
R11355 gnd.n2443 gnd.n2175 9.3005
R11356 gnd.n2180 gnd.n2176 9.3005
R11357 gnd.n2437 gnd.n2181 9.3005
R11358 gnd.n2436 gnd.n2182 9.3005
R11359 gnd.n2435 gnd.n2183 9.3005
R11360 gnd.n2188 gnd.n2184 9.3005
R11361 gnd.n2429 gnd.n2189 9.3005
R11362 gnd.n2428 gnd.n2190 9.3005
R11363 gnd.n2427 gnd.n2191 9.3005
R11364 gnd.n2196 gnd.n2192 9.3005
R11365 gnd.n2421 gnd.n2197 9.3005
R11366 gnd.n2420 gnd.n2198 9.3005
R11367 gnd.n2419 gnd.n2199 9.3005
R11368 gnd.n2204 gnd.n2200 9.3005
R11369 gnd.n2413 gnd.n2205 9.3005
R11370 gnd.n2412 gnd.n2206 9.3005
R11371 gnd.n2411 gnd.n2207 9.3005
R11372 gnd.n2212 gnd.n2208 9.3005
R11373 gnd.n2405 gnd.n2213 9.3005
R11374 gnd.n2404 gnd.n2214 9.3005
R11375 gnd.n2403 gnd.n2215 9.3005
R11376 gnd.n2220 gnd.n2216 9.3005
R11377 gnd.n2397 gnd.n2221 9.3005
R11378 gnd.n2396 gnd.n2222 9.3005
R11379 gnd.n2395 gnd.n2223 9.3005
R11380 gnd.n2228 gnd.n2224 9.3005
R11381 gnd.n2389 gnd.n2229 9.3005
R11382 gnd.n2388 gnd.n2230 9.3005
R11383 gnd.n2387 gnd.n2231 9.3005
R11384 gnd.n2236 gnd.n2232 9.3005
R11385 gnd.n2381 gnd.n2237 9.3005
R11386 gnd.n2380 gnd.n2238 9.3005
R11387 gnd.n2379 gnd.n2239 9.3005
R11388 gnd.n2244 gnd.n2240 9.3005
R11389 gnd.n2373 gnd.n2245 9.3005
R11390 gnd.n2372 gnd.n2246 9.3005
R11391 gnd.n2371 gnd.n2247 9.3005
R11392 gnd.n2252 gnd.n2248 9.3005
R11393 gnd.n2365 gnd.n2253 9.3005
R11394 gnd.n2364 gnd.n2254 9.3005
R11395 gnd.n2363 gnd.n2255 9.3005
R11396 gnd.n2260 gnd.n2256 9.3005
R11397 gnd.n2357 gnd.n2261 9.3005
R11398 gnd.n2356 gnd.n2262 9.3005
R11399 gnd.n2355 gnd.n2263 9.3005
R11400 gnd.n2268 gnd.n2264 9.3005
R11401 gnd.n2349 gnd.n2269 9.3005
R11402 gnd.n2348 gnd.n2270 9.3005
R11403 gnd.n2347 gnd.n2271 9.3005
R11404 gnd.n2276 gnd.n2272 9.3005
R11405 gnd.n2341 gnd.n2277 9.3005
R11406 gnd.n2340 gnd.n2278 9.3005
R11407 gnd.n2339 gnd.n2279 9.3005
R11408 gnd.n2284 gnd.n2280 9.3005
R11409 gnd.n2333 gnd.n2285 9.3005
R11410 gnd.n2332 gnd.n2286 9.3005
R11411 gnd.n2331 gnd.n2287 9.3005
R11412 gnd.n2292 gnd.n2288 9.3005
R11413 gnd.n2325 gnd.n2293 9.3005
R11414 gnd.n2324 gnd.n2294 9.3005
R11415 gnd.n2323 gnd.n2295 9.3005
R11416 gnd.n2300 gnd.n2296 9.3005
R11417 gnd.n2317 gnd.n2301 9.3005
R11418 gnd.n2316 gnd.n2302 9.3005
R11419 gnd.n2315 gnd.n2303 9.3005
R11420 gnd.n2307 gnd.n2304 9.3005
R11421 gnd.n2309 gnd.n2308 9.3005
R11422 gnd.n338 gnd.n337 9.3005
R11423 gnd.n7562 gnd.n7561 9.3005
R11424 gnd.n2476 gnd.n2475 9.3005
R11425 gnd.n7831 gnd.n134 9.3005
R11426 gnd.n7830 gnd.n136 9.3005
R11427 gnd.n140 gnd.n137 9.3005
R11428 gnd.n7825 gnd.n141 9.3005
R11429 gnd.n7824 gnd.n142 9.3005
R11430 gnd.n7823 gnd.n143 9.3005
R11431 gnd.n147 gnd.n144 9.3005
R11432 gnd.n7818 gnd.n148 9.3005
R11433 gnd.n7817 gnd.n149 9.3005
R11434 gnd.n7816 gnd.n150 9.3005
R11435 gnd.n154 gnd.n151 9.3005
R11436 gnd.n7811 gnd.n155 9.3005
R11437 gnd.n7810 gnd.n156 9.3005
R11438 gnd.n7809 gnd.n157 9.3005
R11439 gnd.n161 gnd.n158 9.3005
R11440 gnd.n7804 gnd.n162 9.3005
R11441 gnd.n7803 gnd.n163 9.3005
R11442 gnd.n7799 gnd.n164 9.3005
R11443 gnd.n168 gnd.n165 9.3005
R11444 gnd.n7794 gnd.n169 9.3005
R11445 gnd.n7793 gnd.n170 9.3005
R11446 gnd.n7792 gnd.n171 9.3005
R11447 gnd.n175 gnd.n172 9.3005
R11448 gnd.n7787 gnd.n176 9.3005
R11449 gnd.n7786 gnd.n177 9.3005
R11450 gnd.n7785 gnd.n178 9.3005
R11451 gnd.n182 gnd.n179 9.3005
R11452 gnd.n7780 gnd.n183 9.3005
R11453 gnd.n7779 gnd.n184 9.3005
R11454 gnd.n7778 gnd.n185 9.3005
R11455 gnd.n189 gnd.n186 9.3005
R11456 gnd.n7773 gnd.n190 9.3005
R11457 gnd.n7772 gnd.n191 9.3005
R11458 gnd.n7771 gnd.n192 9.3005
R11459 gnd.n196 gnd.n193 9.3005
R11460 gnd.n7766 gnd.n197 9.3005
R11461 gnd.n7765 gnd.n7764 9.3005
R11462 gnd.n7763 gnd.n200 9.3005
R11463 gnd.n7833 gnd.n7832 9.3005
R11464 gnd.n600 gnd.n599 9.3005
R11465 gnd.n604 gnd.n603 9.3005
R11466 gnd.n605 gnd.n598 9.3005
R11467 gnd.n609 gnd.n606 9.3005
R11468 gnd.n610 gnd.n597 9.3005
R11469 gnd.n614 gnd.n613 9.3005
R11470 gnd.n615 gnd.n596 9.3005
R11471 gnd.n619 gnd.n616 9.3005
R11472 gnd.n620 gnd.n595 9.3005
R11473 gnd.n7131 gnd.n7130 9.3005
R11474 gnd.n7132 gnd.n594 9.3005
R11475 gnd.n7149 gnd.n7133 9.3005
R11476 gnd.n7148 gnd.n7134 9.3005
R11477 gnd.n7147 gnd.n7135 9.3005
R11478 gnd.n7144 gnd.n7136 9.3005
R11479 gnd.n7143 gnd.n7137 9.3005
R11480 gnd.n7141 gnd.n7138 9.3005
R11481 gnd.n7140 gnd.n7139 9.3005
R11482 gnd.n394 gnd.n393 9.3005
R11483 gnd.n7404 gnd.n7403 9.3005
R11484 gnd.n7405 gnd.n392 9.3005
R11485 gnd.n7413 gnd.n7406 9.3005
R11486 gnd.n7412 gnd.n7407 9.3005
R11487 gnd.n7411 gnd.n7408 9.3005
R11488 gnd.n360 gnd.n359 9.3005
R11489 gnd.n7450 gnd.n7449 9.3005
R11490 gnd.n7451 gnd.n358 9.3005
R11491 gnd.n7537 gnd.n7452 9.3005
R11492 gnd.n7536 gnd.n7453 9.3005
R11493 gnd.n7535 gnd.n7454 9.3005
R11494 gnd.n7532 gnd.n7455 9.3005
R11495 gnd.n7531 gnd.n7456 9.3005
R11496 gnd.n7529 gnd.n7457 9.3005
R11497 gnd.n7528 gnd.n7458 9.3005
R11498 gnd.n7526 gnd.n7459 9.3005
R11499 gnd.n7525 gnd.n7460 9.3005
R11500 gnd.n7524 gnd.n7461 9.3005
R11501 gnd.n7522 gnd.n7462 9.3005
R11502 gnd.n7521 gnd.n7463 9.3005
R11503 gnd.n7519 gnd.n7464 9.3005
R11504 gnd.n7518 gnd.n7465 9.3005
R11505 gnd.n7516 gnd.n7466 9.3005
R11506 gnd.n7515 gnd.n7467 9.3005
R11507 gnd.n7513 gnd.n7468 9.3005
R11508 gnd.n7512 gnd.n7469 9.3005
R11509 gnd.n7510 gnd.n7470 9.3005
R11510 gnd.n7509 gnd.n7471 9.3005
R11511 gnd.n7507 gnd.n7472 9.3005
R11512 gnd.n7506 gnd.n7473 9.3005
R11513 gnd.n7504 gnd.n7474 9.3005
R11514 gnd.n7503 gnd.n7475 9.3005
R11515 gnd.n7501 gnd.n7476 9.3005
R11516 gnd.n7500 gnd.n7477 9.3005
R11517 gnd.n7498 gnd.n7478 9.3005
R11518 gnd.n7497 gnd.n7479 9.3005
R11519 gnd.n7495 gnd.n7480 9.3005
R11520 gnd.n7494 gnd.n7481 9.3005
R11521 gnd.n7491 gnd.n7482 9.3005
R11522 gnd.n7490 gnd.n7483 9.3005
R11523 gnd.n7488 gnd.n7484 9.3005
R11524 gnd.n7487 gnd.n7486 9.3005
R11525 gnd.n7485 gnd.n204 9.3005
R11526 gnd.n7760 gnd.n203 9.3005
R11527 gnd.n7762 gnd.n7761 9.3005
R11528 gnd.n580 gnd.n579 9.3005
R11529 gnd.n7183 gnd.n7182 9.3005
R11530 gnd.n7184 gnd.n573 9.3005
R11531 gnd.n7187 gnd.n572 9.3005
R11532 gnd.n7188 gnd.n571 9.3005
R11533 gnd.n7191 gnd.n570 9.3005
R11534 gnd.n7192 gnd.n569 9.3005
R11535 gnd.n7195 gnd.n568 9.3005
R11536 gnd.n7196 gnd.n567 9.3005
R11537 gnd.n7199 gnd.n566 9.3005
R11538 gnd.n7200 gnd.n565 9.3005
R11539 gnd.n7203 gnd.n564 9.3005
R11540 gnd.n7204 gnd.n563 9.3005
R11541 gnd.n7207 gnd.n562 9.3005
R11542 gnd.n7208 gnd.n561 9.3005
R11543 gnd.n7211 gnd.n560 9.3005
R11544 gnd.n7212 gnd.n559 9.3005
R11545 gnd.n7215 gnd.n558 9.3005
R11546 gnd.n7216 gnd.n557 9.3005
R11547 gnd.n7219 gnd.n556 9.3005
R11548 gnd.n7221 gnd.n550 9.3005
R11549 gnd.n7224 gnd.n549 9.3005
R11550 gnd.n7225 gnd.n548 9.3005
R11551 gnd.n7228 gnd.n547 9.3005
R11552 gnd.n7229 gnd.n546 9.3005
R11553 gnd.n7232 gnd.n545 9.3005
R11554 gnd.n7233 gnd.n544 9.3005
R11555 gnd.n7236 gnd.n543 9.3005
R11556 gnd.n7237 gnd.n542 9.3005
R11557 gnd.n7240 gnd.n541 9.3005
R11558 gnd.n7241 gnd.n540 9.3005
R11559 gnd.n7244 gnd.n539 9.3005
R11560 gnd.n7246 gnd.n538 9.3005
R11561 gnd.n7247 gnd.n537 9.3005
R11562 gnd.n7248 gnd.n536 9.3005
R11563 gnd.n7249 gnd.n535 9.3005
R11564 gnd.n7181 gnd.n578 9.3005
R11565 gnd.n7180 gnd.n7179 9.3005
R11566 gnd.n7264 gnd.n7263 9.3005
R11567 gnd.n7265 gnd.n491 9.3005
R11568 gnd.n7267 gnd.n7266 9.3005
R11569 gnd.n475 gnd.n474 9.3005
R11570 gnd.n7280 gnd.n7279 9.3005
R11571 gnd.n7281 gnd.n473 9.3005
R11572 gnd.n7283 gnd.n7282 9.3005
R11573 gnd.n458 gnd.n457 9.3005
R11574 gnd.n7296 gnd.n7295 9.3005
R11575 gnd.n7297 gnd.n456 9.3005
R11576 gnd.n7299 gnd.n7298 9.3005
R11577 gnd.n438 gnd.n437 9.3005
R11578 gnd.n7318 gnd.n7317 9.3005
R11579 gnd.n7319 gnd.n436 9.3005
R11580 gnd.n7323 gnd.n7320 9.3005
R11581 gnd.n7322 gnd.n7321 9.3005
R11582 gnd.n403 gnd.n402 9.3005
R11583 gnd.n7394 gnd.n7393 9.3005
R11584 gnd.n7395 gnd.n401 9.3005
R11585 gnd.n7399 gnd.n7396 9.3005
R11586 gnd.n7398 gnd.n7397 9.3005
R11587 gnd.n370 gnd.n369 9.3005
R11588 gnd.n7441 gnd.n7440 9.3005
R11589 gnd.n7442 gnd.n368 9.3005
R11590 gnd.n7444 gnd.n7443 9.3005
R11591 gnd.n7445 gnd.n302 9.3005
R11592 gnd.n7591 gnd.n7590 9.3005
R11593 gnd.n287 gnd.n286 9.3005
R11594 gnd.n7604 gnd.n7603 9.3005
R11595 gnd.n7605 gnd.n285 9.3005
R11596 gnd.n7607 gnd.n7606 9.3005
R11597 gnd.n273 gnd.n272 9.3005
R11598 gnd.n7620 gnd.n7619 9.3005
R11599 gnd.n7621 gnd.n271 9.3005
R11600 gnd.n7623 gnd.n7622 9.3005
R11601 gnd.n257 gnd.n256 9.3005
R11602 gnd.n7636 gnd.n7635 9.3005
R11603 gnd.n7637 gnd.n255 9.3005
R11604 gnd.n7639 gnd.n7638 9.3005
R11605 gnd.n243 gnd.n242 9.3005
R11606 gnd.n7652 gnd.n7651 9.3005
R11607 gnd.n7653 gnd.n241 9.3005
R11608 gnd.n7655 gnd.n7654 9.3005
R11609 gnd.n227 gnd.n226 9.3005
R11610 gnd.n7668 gnd.n7667 9.3005
R11611 gnd.n7669 gnd.n225 9.3005
R11612 gnd.n7671 gnd.n7670 9.3005
R11613 gnd.n211 gnd.n210 9.3005
R11614 gnd.n7752 gnd.n7751 9.3005
R11615 gnd.n7753 gnd.n209 9.3005
R11616 gnd.n7755 gnd.n7754 9.3005
R11617 gnd.n133 gnd.n132 9.3005
R11618 gnd.n7835 gnd.n7834 9.3005
R11619 gnd.n493 gnd.n492 9.3005
R11620 gnd.n7589 gnd.n301 9.3005
R11621 gnd.n7360 gnd.n7358 9.3005
R11622 gnd.n7367 gnd.n7361 9.3005
R11623 gnd.n7366 gnd.n7362 9.3005
R11624 gnd.n7365 gnd.n7363 9.3005
R11625 gnd.n341 gnd.n340 9.3005
R11626 gnd.n7558 gnd.n339 9.3005
R11627 gnd.n7560 gnd.n7559 9.3005
R11628 gnd.n4968 gnd.n4963 9.3005
R11629 gnd.n4990 gnd.n4969 9.3005
R11630 gnd.n4989 gnd.n4970 9.3005
R11631 gnd.n4988 gnd.n4971 9.3005
R11632 gnd.n4974 gnd.n4972 9.3005
R11633 gnd.n4984 gnd.n4975 9.3005
R11634 gnd.n4983 gnd.n4976 9.3005
R11635 gnd.n4982 gnd.n4977 9.3005
R11636 gnd.n4980 gnd.n4979 9.3005
R11637 gnd.n4978 gnd.n4954 9.3005
R11638 gnd.n4952 gnd.n4951 9.3005
R11639 gnd.n5039 gnd.n5038 9.3005
R11640 gnd.n5040 gnd.n4950 9.3005
R11641 gnd.n5042 gnd.n5041 9.3005
R11642 gnd.n4948 gnd.n4947 9.3005
R11643 gnd.n5047 gnd.n5046 9.3005
R11644 gnd.n5048 gnd.n4946 9.3005
R11645 gnd.n5094 gnd.n5049 9.3005
R11646 gnd.n5093 gnd.n5050 9.3005
R11647 gnd.n5092 gnd.n5051 9.3005
R11648 gnd.n5054 gnd.n5052 9.3005
R11649 gnd.n5088 gnd.n5055 9.3005
R11650 gnd.n5087 gnd.n5056 9.3005
R11651 gnd.n5086 gnd.n5057 9.3005
R11652 gnd.n5060 gnd.n5058 9.3005
R11653 gnd.n5082 gnd.n5061 9.3005
R11654 gnd.n5081 gnd.n5062 9.3005
R11655 gnd.n5080 gnd.n5063 9.3005
R11656 gnd.n5066 gnd.n5064 9.3005
R11657 gnd.n5073 gnd.n5067 9.3005
R11658 gnd.n5072 gnd.n5068 9.3005
R11659 gnd.n5071 gnd.n5069 9.3005
R11660 gnd.n1095 gnd.n1094 9.3005
R11661 gnd.n5803 gnd.n5802 9.3005
R11662 gnd.n5804 gnd.n1093 9.3005
R11663 gnd.n5806 gnd.n5805 9.3005
R11664 gnd.n1082 gnd.n1081 9.3005
R11665 gnd.n5819 gnd.n5818 9.3005
R11666 gnd.n5820 gnd.n1080 9.3005
R11667 gnd.n5822 gnd.n5821 9.3005
R11668 gnd.n1068 gnd.n1067 9.3005
R11669 gnd.n5835 gnd.n5834 9.3005
R11670 gnd.n5836 gnd.n1066 9.3005
R11671 gnd.n5838 gnd.n5837 9.3005
R11672 gnd.n1054 gnd.n1053 9.3005
R11673 gnd.n5851 gnd.n5850 9.3005
R11674 gnd.n5852 gnd.n1052 9.3005
R11675 gnd.n5854 gnd.n5853 9.3005
R11676 gnd.n1039 gnd.n1038 9.3005
R11677 gnd.n5867 gnd.n5866 9.3005
R11678 gnd.n5868 gnd.n1037 9.3005
R11679 gnd.n5870 gnd.n5869 9.3005
R11680 gnd.n1025 gnd.n1024 9.3005
R11681 gnd.n5883 gnd.n5882 9.3005
R11682 gnd.n5884 gnd.n1023 9.3005
R11683 gnd.n5888 gnd.n5885 9.3005
R11684 gnd.n5887 gnd.n5886 9.3005
R11685 gnd.n985 gnd.n984 9.3005
R11686 gnd.n5981 gnd.n5980 9.3005
R11687 gnd.n5982 gnd.n983 9.3005
R11688 gnd.n5984 gnd.n5983 9.3005
R11689 gnd.n969 gnd.n968 9.3005
R11690 gnd.n5997 gnd.n5996 9.3005
R11691 gnd.n5998 gnd.n967 9.3005
R11692 gnd.n6000 gnd.n5999 9.3005
R11693 gnd.n951 gnd.n950 9.3005
R11694 gnd.n6016 gnd.n6015 9.3005
R11695 gnd.n6017 gnd.n949 9.3005
R11696 gnd.n6019 gnd.n6018 9.3005
R11697 gnd.n915 gnd.n914 9.3005
R11698 gnd.n6072 gnd.n6071 9.3005
R11699 gnd.n6073 gnd.n913 9.3005
R11700 gnd.n6077 gnd.n6074 9.3005
R11701 gnd.n6076 gnd.n6075 9.3005
R11702 gnd.n881 gnd.n880 9.3005
R11703 gnd.n6836 gnd.n6835 9.3005
R11704 gnd.n6837 gnd.n879 9.3005
R11705 gnd.n6839 gnd.n6838 9.3005
R11706 gnd.n866 gnd.n865 9.3005
R11707 gnd.n6852 gnd.n6851 9.3005
R11708 gnd.n6853 gnd.n864 9.3005
R11709 gnd.n6855 gnd.n6854 9.3005
R11710 gnd.n850 gnd.n849 9.3005
R11711 gnd.n6868 gnd.n6867 9.3005
R11712 gnd.n6869 gnd.n848 9.3005
R11713 gnd.n6871 gnd.n6870 9.3005
R11714 gnd.n834 gnd.n833 9.3005
R11715 gnd.n6884 gnd.n6883 9.3005
R11716 gnd.n6885 gnd.n832 9.3005
R11717 gnd.n6887 gnd.n6886 9.3005
R11718 gnd.n818 gnd.n817 9.3005
R11719 gnd.n6900 gnd.n6899 9.3005
R11720 gnd.n6901 gnd.n816 9.3005
R11721 gnd.n6903 gnd.n6902 9.3005
R11722 gnd.n803 gnd.n802 9.3005
R11723 gnd.n6916 gnd.n6915 9.3005
R11724 gnd.n6917 gnd.n801 9.3005
R11725 gnd.n6919 gnd.n6918 9.3005
R11726 gnd.n787 gnd.n786 9.3005
R11727 gnd.n6932 gnd.n6931 9.3005
R11728 gnd.n6933 gnd.n785 9.3005
R11729 gnd.n6935 gnd.n6934 9.3005
R11730 gnd.n771 gnd.n770 9.3005
R11731 gnd.n6948 gnd.n6947 9.3005
R11732 gnd.n6949 gnd.n769 9.3005
R11733 gnd.n6951 gnd.n6950 9.3005
R11734 gnd.n755 gnd.n754 9.3005
R11735 gnd.n6964 gnd.n6963 9.3005
R11736 gnd.n6965 gnd.n753 9.3005
R11737 gnd.n6967 gnd.n6966 9.3005
R11738 gnd.n739 gnd.n738 9.3005
R11739 gnd.n6980 gnd.n6979 9.3005
R11740 gnd.n6981 gnd.n737 9.3005
R11741 gnd.n6983 gnd.n6982 9.3005
R11742 gnd.n724 gnd.n723 9.3005
R11743 gnd.n6996 gnd.n6995 9.3005
R11744 gnd.n6997 gnd.n722 9.3005
R11745 gnd.n6999 gnd.n6998 9.3005
R11746 gnd.n710 gnd.n709 9.3005
R11747 gnd.n7012 gnd.n7011 9.3005
R11748 gnd.n7013 gnd.n708 9.3005
R11749 gnd.n7015 gnd.n7014 9.3005
R11750 gnd.n696 gnd.n695 9.3005
R11751 gnd.n7028 gnd.n7027 9.3005
R11752 gnd.n7029 gnd.n694 9.3005
R11753 gnd.n7031 gnd.n7030 9.3005
R11754 gnd.n682 gnd.n681 9.3005
R11755 gnd.n7044 gnd.n7043 9.3005
R11756 gnd.n7045 gnd.n680 9.3005
R11757 gnd.n7047 gnd.n7046 9.3005
R11758 gnd.n667 gnd.n666 9.3005
R11759 gnd.n7061 gnd.n7060 9.3005
R11760 gnd.n7062 gnd.n665 9.3005
R11761 gnd.n7066 gnd.n7063 9.3005
R11762 gnd.n7065 gnd.n7064 9.3005
R11763 gnd.n637 gnd.n636 9.3005
R11764 gnd.n7081 gnd.n7080 9.3005
R11765 gnd.n7082 gnd.n635 9.3005
R11766 gnd.n7084 gnd.n7083 9.3005
R11767 gnd.n633 gnd.n632 9.3005
R11768 gnd.n7089 gnd.n7088 9.3005
R11769 gnd.n7090 gnd.n631 9.3005
R11770 gnd.n7092 gnd.n7091 9.3005
R11771 gnd.n629 gnd.n628 9.3005
R11772 gnd.n7097 gnd.n7096 9.3005
R11773 gnd.n7098 gnd.n627 9.3005
R11774 gnd.n7100 gnd.n7099 9.3005
R11775 gnd.n625 gnd.n624 9.3005
R11776 gnd.n7105 gnd.n7104 9.3005
R11777 gnd.n7106 gnd.n623 9.3005
R11778 gnd.n7125 gnd.n7107 9.3005
R11779 gnd.n7124 gnd.n7108 9.3005
R11780 gnd.n7123 gnd.n7109 9.3005
R11781 gnd.n7112 gnd.n7110 9.3005
R11782 gnd.n7119 gnd.n7113 9.3005
R11783 gnd.n7118 gnd.n7114 9.3005
R11784 gnd.n7117 gnd.n7116 9.3005
R11785 gnd.n7115 gnd.n421 9.3005
R11786 gnd.n419 gnd.n418 9.3005
R11787 gnd.n7347 gnd.n7346 9.3005
R11788 gnd.n7348 gnd.n417 9.3005
R11789 gnd.n7379 gnd.n7349 9.3005
R11790 gnd.n7378 gnd.n7350 9.3005
R11791 gnd.n7377 gnd.n7351 9.3005
R11792 gnd.n7354 gnd.n7352 9.3005
R11793 gnd.n7373 gnd.n7355 9.3005
R11794 gnd.n7372 gnd.n7356 9.3005
R11795 gnd.n7371 gnd.n7357 9.3005
R11796 gnd.n4910 gnd.n4909 9.3005
R11797 gnd.n4564 gnd.n4515 9.3005
R11798 gnd.n4563 gnd.n4516 9.3005
R11799 gnd.n4562 gnd.n4517 9.3005
R11800 gnd.n4560 gnd.n4518 9.3005
R11801 gnd.n4559 gnd.n4519 9.3005
R11802 gnd.n4557 gnd.n4520 9.3005
R11803 gnd.n4556 gnd.n4521 9.3005
R11804 gnd.n4554 gnd.n4522 9.3005
R11805 gnd.n4553 gnd.n4523 9.3005
R11806 gnd.n4551 gnd.n4524 9.3005
R11807 gnd.n4550 gnd.n4525 9.3005
R11808 gnd.n4548 gnd.n4526 9.3005
R11809 gnd.n4547 gnd.n4527 9.3005
R11810 gnd.n4545 gnd.n4528 9.3005
R11811 gnd.n4544 gnd.n4529 9.3005
R11812 gnd.n4542 gnd.n4530 9.3005
R11813 gnd.n4541 gnd.n4531 9.3005
R11814 gnd.n4539 gnd.n4532 9.3005
R11815 gnd.n4538 gnd.n4533 9.3005
R11816 gnd.n4536 gnd.n4535 9.3005
R11817 gnd.n4534 gnd.n1476 9.3005
R11818 gnd.n4863 gnd.n1475 9.3005
R11819 gnd.n4865 gnd.n4864 9.3005
R11820 gnd.n4866 gnd.n1474 9.3005
R11821 gnd.n4871 gnd.n4867 9.3005
R11822 gnd.n4870 gnd.n4869 9.3005
R11823 gnd.n4868 gnd.n1440 9.3005
R11824 gnd.n4903 gnd.n1441 9.3005
R11825 gnd.n4904 gnd.n1439 9.3005
R11826 gnd.n4907 gnd.n4906 9.3005
R11827 gnd.n4908 gnd.n1438 9.3005
R11828 gnd.n4514 gnd.n4447 9.3005
R11829 gnd.n4507 gnd.n4506 9.3005
R11830 gnd.n4505 gnd.n4453 9.3005
R11831 gnd.n4504 gnd.n4503 9.3005
R11832 gnd.n4455 gnd.n4454 9.3005
R11833 gnd.n4497 gnd.n4496 9.3005
R11834 gnd.n4495 gnd.n4457 9.3005
R11835 gnd.n4494 gnd.n4493 9.3005
R11836 gnd.n4459 gnd.n4458 9.3005
R11837 gnd.n4487 gnd.n4486 9.3005
R11838 gnd.n4485 gnd.n4461 9.3005
R11839 gnd.n4484 gnd.n4483 9.3005
R11840 gnd.n4463 gnd.n4462 9.3005
R11841 gnd.n4477 gnd.n4476 9.3005
R11842 gnd.n4475 gnd.n4465 9.3005
R11843 gnd.n4474 gnd.n4473 9.3005
R11844 gnd.n4468 gnd.n4466 9.3005
R11845 gnd.n4467 gnd.n1562 9.3005
R11846 gnd.n4451 gnd.n4448 9.3005
R11847 gnd.n4513 gnd.n4512 9.3005
R11848 gnd.n4762 gnd.n1561 9.3005
R11849 gnd.n4764 gnd.n4763 9.3005
R11850 gnd.n1548 gnd.n1547 9.3005
R11851 gnd.n4777 gnd.n4776 9.3005
R11852 gnd.n4778 gnd.n1546 9.3005
R11853 gnd.n4780 gnd.n4779 9.3005
R11854 gnd.n1531 gnd.n1530 9.3005
R11855 gnd.n4793 gnd.n4792 9.3005
R11856 gnd.n4794 gnd.n1529 9.3005
R11857 gnd.n4796 gnd.n4795 9.3005
R11858 gnd.n1516 gnd.n1515 9.3005
R11859 gnd.n4809 gnd.n4808 9.3005
R11860 gnd.n4810 gnd.n1514 9.3005
R11861 gnd.n4812 gnd.n4811 9.3005
R11862 gnd.n1499 gnd.n1498 9.3005
R11863 gnd.n4825 gnd.n4824 9.3005
R11864 gnd.n4826 gnd.n1497 9.3005
R11865 gnd.n4836 gnd.n4827 9.3005
R11866 gnd.n4835 gnd.n4828 9.3005
R11867 gnd.n4834 gnd.n4829 9.3005
R11868 gnd.n4833 gnd.n4831 9.3005
R11869 gnd.n4830 gnd.n1463 9.3005
R11870 gnd.n4877 gnd.n1464 9.3005
R11871 gnd.n4876 gnd.n1465 9.3005
R11872 gnd.n4875 gnd.n1466 9.3005
R11873 gnd.n1472 gnd.n1467 9.3005
R11874 gnd.n1471 gnd.n1469 9.3005
R11875 gnd.n1468 gnd.n1398 9.3005
R11876 gnd.n5236 gnd.n1399 9.3005
R11877 gnd.n5235 gnd.n1400 9.3005
R11878 gnd.n5234 gnd.n1401 9.3005
R11879 gnd.n5207 gnd.n1402 9.3005
R11880 gnd.n5210 gnd.n5209 9.3005
R11881 gnd.n5211 gnd.n1427 9.3005
R11882 gnd.n5213 gnd.n5212 9.3005
R11883 gnd.n1375 gnd.n1374 9.3005
R11884 gnd.n5249 gnd.n5248 9.3005
R11885 gnd.n5250 gnd.n1373 9.3005
R11886 gnd.n5252 gnd.n5251 9.3005
R11887 gnd.n1358 gnd.n1357 9.3005
R11888 gnd.n5265 gnd.n5264 9.3005
R11889 gnd.n5266 gnd.n1356 9.3005
R11890 gnd.n5268 gnd.n5267 9.3005
R11891 gnd.n1340 gnd.n1339 9.3005
R11892 gnd.n5281 gnd.n5280 9.3005
R11893 gnd.n5282 gnd.n1338 9.3005
R11894 gnd.n5284 gnd.n5283 9.3005
R11895 gnd.n1323 gnd.n1322 9.3005
R11896 gnd.n5297 gnd.n5296 9.3005
R11897 gnd.n5298 gnd.n1321 9.3005
R11898 gnd.n5300 gnd.n5299 9.3005
R11899 gnd.n1305 gnd.n1304 9.3005
R11900 gnd.n5313 gnd.n5312 9.3005
R11901 gnd.n5314 gnd.n1303 9.3005
R11902 gnd.n5316 gnd.n5315 9.3005
R11903 gnd.n1288 gnd.n1287 9.3005
R11904 gnd.n5329 gnd.n5328 9.3005
R11905 gnd.n5330 gnd.n1286 9.3005
R11906 gnd.n5332 gnd.n5331 9.3005
R11907 gnd.n1269 gnd.n1268 9.3005
R11908 gnd.n5347 gnd.n5346 9.3005
R11909 gnd.n5348 gnd.n1267 9.3005
R11910 gnd.n5662 gnd.n5349 9.3005
R11911 gnd.n5661 gnd.n5660 9.3005
R11912 gnd.n4761 gnd.n4760 9.3005
R11913 gnd.n1224 gnd.n1218 9.3005
R11914 gnd.n5712 gnd.n1217 9.3005
R11915 gnd.n5713 gnd.n1216 9.3005
R11916 gnd.n5714 gnd.n1215 9.3005
R11917 gnd.n1214 gnd.n1211 9.3005
R11918 gnd.n5719 gnd.n1210 9.3005
R11919 gnd.n5720 gnd.n1209 9.3005
R11920 gnd.n5721 gnd.n1208 9.3005
R11921 gnd.n1207 gnd.n1204 9.3005
R11922 gnd.n5726 gnd.n1203 9.3005
R11923 gnd.n5727 gnd.n1202 9.3005
R11924 gnd.n5728 gnd.n1201 9.3005
R11925 gnd.n1200 gnd.n1197 9.3005
R11926 gnd.n1199 gnd.n1184 9.3005
R11927 gnd.n5735 gnd.n1183 9.3005
R11928 gnd.n5737 gnd.n5736 9.3005
R11929 gnd.n5704 gnd.n1227 9.3005
R11930 gnd.n5703 gnd.n1228 9.3005
R11931 gnd.n1232 gnd.n1229 9.3005
R11932 gnd.n5698 gnd.n1233 9.3005
R11933 gnd.n5697 gnd.n1234 9.3005
R11934 gnd.n5696 gnd.n1235 9.3005
R11935 gnd.n1239 gnd.n1236 9.3005
R11936 gnd.n5691 gnd.n1240 9.3005
R11937 gnd.n5690 gnd.n1241 9.3005
R11938 gnd.n5689 gnd.n1242 9.3005
R11939 gnd.n1246 gnd.n1243 9.3005
R11940 gnd.n5684 gnd.n1247 9.3005
R11941 gnd.n5683 gnd.n1248 9.3005
R11942 gnd.n5682 gnd.n1249 9.3005
R11943 gnd.n1253 gnd.n1250 9.3005
R11944 gnd.n5677 gnd.n1254 9.3005
R11945 gnd.n5676 gnd.n1255 9.3005
R11946 gnd.n5675 gnd.n1256 9.3005
R11947 gnd.n1261 gnd.n1259 9.3005
R11948 gnd.n5670 gnd.n5669 9.3005
R11949 gnd.n5705 gnd.n1226 9.3005
R11950 gnd.n4673 gnd.n4629 9.3005
R11951 gnd.n4672 gnd.n4631 9.3005
R11952 gnd.n4671 gnd.n4632 9.3005
R11953 gnd.n4669 gnd.n4633 9.3005
R11954 gnd.n4668 gnd.n4634 9.3005
R11955 gnd.n4666 gnd.n4635 9.3005
R11956 gnd.n4665 gnd.n4636 9.3005
R11957 gnd.n4663 gnd.n4637 9.3005
R11958 gnd.n4662 gnd.n4638 9.3005
R11959 gnd.n4660 gnd.n4639 9.3005
R11960 gnd.n4659 gnd.n4640 9.3005
R11961 gnd.n4657 gnd.n4641 9.3005
R11962 gnd.n4656 gnd.n4642 9.3005
R11963 gnd.n4654 gnd.n4643 9.3005
R11964 gnd.n4653 gnd.n4644 9.3005
R11965 gnd.n4651 gnd.n4645 9.3005
R11966 gnd.n4650 gnd.n4646 9.3005
R11967 gnd.n4648 gnd.n4647 9.3005
R11968 gnd.n1482 gnd.n1481 9.3005
R11969 gnd.n4851 gnd.n4850 9.3005
R11970 gnd.n4852 gnd.n1480 9.3005
R11971 gnd.n4859 gnd.n4853 9.3005
R11972 gnd.n4858 gnd.n4854 9.3005
R11973 gnd.n4857 gnd.n4855 9.3005
R11974 gnd.n1447 gnd.n1446 9.3005
R11975 gnd.n4891 gnd.n4890 9.3005
R11976 gnd.n4892 gnd.n1445 9.3005
R11977 gnd.n4899 gnd.n4893 9.3005
R11978 gnd.n4898 gnd.n4894 9.3005
R11979 gnd.n4897 gnd.n4895 9.3005
R11980 gnd.n1430 gnd.n1428 9.3005
R11981 gnd.n5206 gnd.n5205 9.3005
R11982 gnd.n5204 gnd.n1429 9.3005
R11983 gnd.n5201 gnd.n1431 9.3005
R11984 gnd.n5200 gnd.n1432 9.3005
R11985 gnd.n5199 gnd.n1433 9.3005
R11986 gnd.n4959 gnd.n1434 9.3005
R11987 gnd.n4995 gnd.n4960 9.3005
R11988 gnd.n4996 gnd.n4958 9.3005
R11989 gnd.n5000 gnd.n4999 9.3005
R11990 gnd.n5001 gnd.n4957 9.3005
R11991 gnd.n5005 gnd.n5002 9.3005
R11992 gnd.n5006 gnd.n4956 9.3005
R11993 gnd.n5010 gnd.n5009 9.3005
R11994 gnd.n5011 gnd.n4955 9.3005
R11995 gnd.n5031 gnd.n5012 9.3005
R11996 gnd.n5030 gnd.n5013 9.3005
R11997 gnd.n5029 gnd.n5014 9.3005
R11998 gnd.n5026 gnd.n5015 9.3005
R11999 gnd.n5025 gnd.n5016 9.3005
R12000 gnd.n5022 gnd.n5017 9.3005
R12001 gnd.n5021 gnd.n5018 9.3005
R12002 gnd.n4943 gnd.n4942 9.3005
R12003 gnd.n5100 gnd.n5099 9.3005
R12004 gnd.n5101 gnd.n4941 9.3005
R12005 gnd.n5105 gnd.n5102 9.3005
R12006 gnd.n5106 gnd.n4940 9.3005
R12007 gnd.n5110 gnd.n5109 9.3005
R12008 gnd.n5111 gnd.n4939 9.3005
R12009 gnd.n5116 gnd.n5112 9.3005
R12010 gnd.n5115 gnd.n5114 9.3005
R12011 gnd.n5113 gnd.n1263 9.3005
R12012 gnd.n5666 gnd.n1262 9.3005
R12013 gnd.n5668 gnd.n5667 9.3005
R12014 gnd.n4675 gnd.n4674 9.3005
R12015 gnd.n4683 gnd.n4682 9.3005
R12016 gnd.n4684 gnd.n4623 9.3005
R12017 gnd.n4685 gnd.n4622 9.3005
R12018 gnd.n4621 gnd.n4619 9.3005
R12019 gnd.n4691 gnd.n4618 9.3005
R12020 gnd.n4692 gnd.n4617 9.3005
R12021 gnd.n4693 gnd.n4616 9.3005
R12022 gnd.n4615 gnd.n4613 9.3005
R12023 gnd.n4699 gnd.n4612 9.3005
R12024 gnd.n4700 gnd.n4611 9.3005
R12025 gnd.n4701 gnd.n4610 9.3005
R12026 gnd.n4609 gnd.n4607 9.3005
R12027 gnd.n4707 gnd.n4606 9.3005
R12028 gnd.n4708 gnd.n4605 9.3005
R12029 gnd.n4709 gnd.n4604 9.3005
R12030 gnd.n4603 gnd.n4601 9.3005
R12031 gnd.n4715 gnd.n4600 9.3005
R12032 gnd.n4716 gnd.n4599 9.3005
R12033 gnd.n4717 gnd.n4598 9.3005
R12034 gnd.n4597 gnd.n4592 9.3005
R12035 gnd.n4723 gnd.n4591 9.3005
R12036 gnd.n4724 gnd.n4590 9.3005
R12037 gnd.n4725 gnd.n4589 9.3005
R12038 gnd.n4588 gnd.n4586 9.3005
R12039 gnd.n4731 gnd.n4585 9.3005
R12040 gnd.n4732 gnd.n4584 9.3005
R12041 gnd.n4733 gnd.n4583 9.3005
R12042 gnd.n4582 gnd.n4580 9.3005
R12043 gnd.n4739 gnd.n4579 9.3005
R12044 gnd.n4740 gnd.n4578 9.3005
R12045 gnd.n4741 gnd.n4577 9.3005
R12046 gnd.n4576 gnd.n4574 9.3005
R12047 gnd.n4746 gnd.n4573 9.3005
R12048 gnd.n4747 gnd.n4572 9.3005
R12049 gnd.n4571 gnd.n4569 9.3005
R12050 gnd.n4752 gnd.n4568 9.3005
R12051 gnd.n4754 gnd.n4753 9.3005
R12052 gnd.n4681 gnd.n4628 9.3005
R12053 gnd.n4680 gnd.n4679 9.3005
R12054 gnd.n1556 gnd.n1555 9.3005
R12055 gnd.n4769 gnd.n4768 9.3005
R12056 gnd.n4770 gnd.n1554 9.3005
R12057 gnd.n4772 gnd.n4771 9.3005
R12058 gnd.n1540 gnd.n1539 9.3005
R12059 gnd.n4785 gnd.n4784 9.3005
R12060 gnd.n4786 gnd.n1538 9.3005
R12061 gnd.n4788 gnd.n4787 9.3005
R12062 gnd.n1524 gnd.n1523 9.3005
R12063 gnd.n4801 gnd.n4800 9.3005
R12064 gnd.n4802 gnd.n1522 9.3005
R12065 gnd.n4804 gnd.n4803 9.3005
R12066 gnd.n1508 gnd.n1507 9.3005
R12067 gnd.n4817 gnd.n4816 9.3005
R12068 gnd.n4818 gnd.n1506 9.3005
R12069 gnd.n4820 gnd.n4819 9.3005
R12070 gnd.n1491 gnd.n1490 9.3005
R12071 gnd.n4841 gnd.n4840 9.3005
R12072 gnd.n4842 gnd.n1489 9.3005
R12073 gnd.n4846 gnd.n4843 9.3005
R12074 gnd.n4845 gnd.n4844 9.3005
R12075 gnd.n1455 gnd.n1454 9.3005
R12076 gnd.n4882 gnd.n4881 9.3005
R12077 gnd.n4883 gnd.n1453 9.3005
R12078 gnd.n4885 gnd.n4884 9.3005
R12079 gnd.n4886 gnd.n1383 9.3005
R12080 gnd.n1367 gnd.n1366 9.3005
R12081 gnd.n5257 gnd.n5256 9.3005
R12082 gnd.n5258 gnd.n1365 9.3005
R12083 gnd.n5260 gnd.n5259 9.3005
R12084 gnd.n1349 gnd.n1348 9.3005
R12085 gnd.n5273 gnd.n5272 9.3005
R12086 gnd.n5274 gnd.n1347 9.3005
R12087 gnd.n5276 gnd.n5275 9.3005
R12088 gnd.n1332 gnd.n1331 9.3005
R12089 gnd.n5289 gnd.n5288 9.3005
R12090 gnd.n5290 gnd.n1330 9.3005
R12091 gnd.n5292 gnd.n5291 9.3005
R12092 gnd.n1314 gnd.n1313 9.3005
R12093 gnd.n5305 gnd.n5304 9.3005
R12094 gnd.n5306 gnd.n1312 9.3005
R12095 gnd.n5308 gnd.n5307 9.3005
R12096 gnd.n1297 gnd.n1296 9.3005
R12097 gnd.n5321 gnd.n5320 9.3005
R12098 gnd.n5322 gnd.n1295 9.3005
R12099 gnd.n5324 gnd.n5323 9.3005
R12100 gnd.n1279 gnd.n1278 9.3005
R12101 gnd.n5337 gnd.n5336 9.3005
R12102 gnd.n5338 gnd.n1277 9.3005
R12103 gnd.n5342 gnd.n5339 9.3005
R12104 gnd.n5341 gnd.n5340 9.3005
R12105 gnd.n1182 gnd.n1181 9.3005
R12106 gnd.n5739 gnd.n5738 9.3005
R12107 gnd.n4756 gnd.n4755 9.3005
R12108 gnd.n5244 gnd.n5243 9.3005
R12109 gnd.n3051 gnd.n1415 9.3005
R12110 gnd.n5224 gnd.n1416 9.3005
R12111 gnd.n5223 gnd.n1417 9.3005
R12112 gnd.n5222 gnd.n1418 9.3005
R12113 gnd.n4964 gnd.n1419 9.3005
R12114 gnd.n4967 gnd.n4966 9.3005
R12115 gnd.n3055 gnd.n3054 9.3005
R12116 gnd.n3058 gnd.n3050 9.3005
R12117 gnd.n3049 gnd.n1659 9.3005
R12118 gnd.n3048 gnd.n3047 9.3005
R12119 gnd.n1661 gnd.n1660 9.3005
R12120 gnd.n3041 gnd.n3040 9.3005
R12121 gnd.n3039 gnd.n1665 9.3005
R12122 gnd.n3038 gnd.n3037 9.3005
R12123 gnd.n1667 gnd.n1666 9.3005
R12124 gnd.n3031 gnd.n3030 9.3005
R12125 gnd.n3029 gnd.n1671 9.3005
R12126 gnd.n3028 gnd.n3027 9.3005
R12127 gnd.n1673 gnd.n1672 9.3005
R12128 gnd.n3021 gnd.n3020 9.3005
R12129 gnd.n3019 gnd.n1677 9.3005
R12130 gnd.n3018 gnd.n3017 9.3005
R12131 gnd.n1679 gnd.n1678 9.3005
R12132 gnd.n3011 gnd.n3010 9.3005
R12133 gnd.n3009 gnd.n1683 9.3005
R12134 gnd.n3008 gnd.n3007 9.3005
R12135 gnd.n1685 gnd.n1684 9.3005
R12136 gnd.n3001 gnd.n3000 9.3005
R12137 gnd.n2999 gnd.n1689 9.3005
R12138 gnd.n2998 gnd.n2997 9.3005
R12139 gnd.n1691 gnd.n1690 9.3005
R12140 gnd.n2991 gnd.n2990 9.3005
R12141 gnd.n2989 gnd.n1695 9.3005
R12142 gnd.n2988 gnd.n2987 9.3005
R12143 gnd.n1697 gnd.n1696 9.3005
R12144 gnd.n2981 gnd.n2980 9.3005
R12145 gnd.n2979 gnd.n1701 9.3005
R12146 gnd.n2978 gnd.n2977 9.3005
R12147 gnd.n1703 gnd.n1702 9.3005
R12148 gnd.n2971 gnd.n2970 9.3005
R12149 gnd.n2969 gnd.n1707 9.3005
R12150 gnd.n2968 gnd.n2967 9.3005
R12151 gnd.n1709 gnd.n1708 9.3005
R12152 gnd.n2961 gnd.n2960 9.3005
R12153 gnd.n2959 gnd.n1713 9.3005
R12154 gnd.n2958 gnd.n2957 9.3005
R12155 gnd.n1715 gnd.n1714 9.3005
R12156 gnd.n2951 gnd.n2950 9.3005
R12157 gnd.n2949 gnd.n1719 9.3005
R12158 gnd.n2948 gnd.n2947 9.3005
R12159 gnd.n1721 gnd.n1720 9.3005
R12160 gnd.n2941 gnd.n2940 9.3005
R12161 gnd.n2939 gnd.n1725 9.3005
R12162 gnd.n2938 gnd.n2937 9.3005
R12163 gnd.n1727 gnd.n1726 9.3005
R12164 gnd.n2931 gnd.n2930 9.3005
R12165 gnd.n2929 gnd.n1731 9.3005
R12166 gnd.n2928 gnd.n2927 9.3005
R12167 gnd.n1733 gnd.n1732 9.3005
R12168 gnd.n2921 gnd.n2920 9.3005
R12169 gnd.n2919 gnd.n1737 9.3005
R12170 gnd.n2918 gnd.n2917 9.3005
R12171 gnd.n1739 gnd.n1738 9.3005
R12172 gnd.n2911 gnd.n2910 9.3005
R12173 gnd.n2909 gnd.n1743 9.3005
R12174 gnd.n2908 gnd.n2907 9.3005
R12175 gnd.n1745 gnd.n1744 9.3005
R12176 gnd.n2901 gnd.n2900 9.3005
R12177 gnd.n2899 gnd.n1749 9.3005
R12178 gnd.n2898 gnd.n2897 9.3005
R12179 gnd.n1751 gnd.n1750 9.3005
R12180 gnd.n2891 gnd.n2890 9.3005
R12181 gnd.n2889 gnd.n1755 9.3005
R12182 gnd.n2888 gnd.n2887 9.3005
R12183 gnd.n1757 gnd.n1756 9.3005
R12184 gnd.n2881 gnd.n2880 9.3005
R12185 gnd.n2879 gnd.n1761 9.3005
R12186 gnd.n2878 gnd.n2877 9.3005
R12187 gnd.n1763 gnd.n1762 9.3005
R12188 gnd.n2871 gnd.n2870 9.3005
R12189 gnd.n2869 gnd.n1767 9.3005
R12190 gnd.n2868 gnd.n2867 9.3005
R12191 gnd.n1769 gnd.n1768 9.3005
R12192 gnd.n2861 gnd.n2860 9.3005
R12193 gnd.n2859 gnd.n1773 9.3005
R12194 gnd.n2858 gnd.n2857 9.3005
R12195 gnd.n1775 gnd.n1774 9.3005
R12196 gnd.n2851 gnd.n2850 9.3005
R12197 gnd.n2849 gnd.n1779 9.3005
R12198 gnd.n2848 gnd.n2847 9.3005
R12199 gnd.n1781 gnd.n1780 9.3005
R12200 gnd.n3057 gnd.n3056 9.3005
R12201 gnd.n6598 gnd.n6596 9.3005
R12202 gnd.n6725 gnd.n6724 9.3005
R12203 gnd.n6723 gnd.n6722 9.3005
R12204 gnd.n6609 gnd.n6608 9.3005
R12205 gnd.n6717 gnd.n6716 9.3005
R12206 gnd.n6715 gnd.n6714 9.3005
R12207 gnd.n6617 gnd.n6616 9.3005
R12208 gnd.n6709 gnd.n6708 9.3005
R12209 gnd.n6707 gnd.n6706 9.3005
R12210 gnd.n6629 gnd.n6628 9.3005
R12211 gnd.n6701 gnd.n6700 9.3005
R12212 gnd.n6699 gnd.n6698 9.3005
R12213 gnd.n6637 gnd.n6636 9.3005
R12214 gnd.n6693 gnd.n6692 9.3005
R12215 gnd.n6691 gnd.n6690 9.3005
R12216 gnd.n6649 gnd.n6648 9.3005
R12217 gnd.n6682 gnd.n6681 9.3005
R12218 gnd.n6680 gnd.n6650 9.3005
R12219 gnd.n6731 gnd.n6730 9.3005
R12220 gnd.n6643 gnd.n6642 9.3005
R12221 gnd.n6695 gnd.n6694 9.3005
R12222 gnd.n6697 gnd.n6696 9.3005
R12223 gnd.n6633 gnd.n6632 9.3005
R12224 gnd.n6703 gnd.n6702 9.3005
R12225 gnd.n6705 gnd.n6704 9.3005
R12226 gnd.n6623 gnd.n6622 9.3005
R12227 gnd.n6711 gnd.n6710 9.3005
R12228 gnd.n6713 gnd.n6712 9.3005
R12229 gnd.n6613 gnd.n6612 9.3005
R12230 gnd.n6719 gnd.n6718 9.3005
R12231 gnd.n6721 gnd.n6720 9.3005
R12232 gnd.n6603 gnd.n6602 9.3005
R12233 gnd.n6727 gnd.n6726 9.3005
R12234 gnd.n6729 gnd.n6728 9.3005
R12235 gnd.n6597 gnd.n502 9.3005
R12236 gnd.n6689 gnd.n6688 9.3005
R12237 gnd.n6684 gnd.n6683 9.3005
R12238 gnd.n6679 gnd.n6678 9.3005
R12239 gnd.n6677 gnd.n6655 9.3005
R12240 gnd.n6676 gnd.n6675 9.3005
R12241 gnd.n6674 gnd.n6656 9.3005
R12242 gnd.n6673 gnd.n6672 9.3005
R12243 gnd.n6671 gnd.n6661 9.3005
R12244 gnd.n6670 gnd.n6669 9.3005
R12245 gnd.n6668 gnd.n6662 9.3005
R12246 gnd.n657 gnd.n656 9.3005
R12247 gnd.n7074 gnd.n7073 9.3005
R12248 gnd.n1089 gnd.n1088 9.3005
R12249 gnd.n5811 gnd.n5810 9.3005
R12250 gnd.n5812 gnd.n1087 9.3005
R12251 gnd.n5814 gnd.n5813 9.3005
R12252 gnd.n1075 gnd.n1074 9.3005
R12253 gnd.n5827 gnd.n5826 9.3005
R12254 gnd.n5828 gnd.n1073 9.3005
R12255 gnd.n5830 gnd.n5829 9.3005
R12256 gnd.n1060 gnd.n1059 9.3005
R12257 gnd.n5843 gnd.n5842 9.3005
R12258 gnd.n5844 gnd.n1058 9.3005
R12259 gnd.n5846 gnd.n5845 9.3005
R12260 gnd.n1046 gnd.n1045 9.3005
R12261 gnd.n5859 gnd.n5858 9.3005
R12262 gnd.n5860 gnd.n1044 9.3005
R12263 gnd.n5862 gnd.n5861 9.3005
R12264 gnd.n1032 gnd.n1031 9.3005
R12265 gnd.n5875 gnd.n5874 9.3005
R12266 gnd.n5876 gnd.n1030 9.3005
R12267 gnd.n5878 gnd.n5877 9.3005
R12268 gnd.n1016 gnd.n1015 9.3005
R12269 gnd.n5893 gnd.n5892 9.3005
R12270 gnd.n5894 gnd.n1013 9.3005
R12271 gnd.n5897 gnd.n5896 9.3005
R12272 gnd.n5895 gnd.n1014 9.3005
R12273 gnd.n977 gnd.n976 9.3005
R12274 gnd.n5989 gnd.n5988 9.3005
R12275 gnd.n5990 gnd.n975 9.3005
R12276 gnd.n5992 gnd.n5991 9.3005
R12277 gnd.n961 gnd.n960 9.3005
R12278 gnd.n6005 gnd.n6004 9.3005
R12279 gnd.n6006 gnd.n958 9.3005
R12280 gnd.n6011 gnd.n6010 9.3005
R12281 gnd.n6009 gnd.n959 9.3005
R12282 gnd.n6008 gnd.n6007 9.3005
R12283 gnd.n924 gnd.n922 9.3005
R12284 gnd.n6067 gnd.n6066 9.3005
R12285 gnd.n6065 gnd.n923 9.3005
R12286 gnd.n6064 gnd.n6063 9.3005
R12287 gnd.n6062 gnd.n925 9.3005
R12288 gnd.n6061 gnd.n6060 9.3005
R12289 gnd.n6059 gnd.n6058 9.3005
R12290 gnd.n874 gnd.n873 9.3005
R12291 gnd.n6844 gnd.n6843 9.3005
R12292 gnd.n6845 gnd.n872 9.3005
R12293 gnd.n6847 gnd.n6846 9.3005
R12294 gnd.n858 gnd.n857 9.3005
R12295 gnd.n6860 gnd.n6859 9.3005
R12296 gnd.n6861 gnd.n856 9.3005
R12297 gnd.n6863 gnd.n6862 9.3005
R12298 gnd.n842 gnd.n841 9.3005
R12299 gnd.n6876 gnd.n6875 9.3005
R12300 gnd.n6877 gnd.n840 9.3005
R12301 gnd.n6879 gnd.n6878 9.3005
R12302 gnd.n826 gnd.n825 9.3005
R12303 gnd.n6892 gnd.n6891 9.3005
R12304 gnd.n6893 gnd.n824 9.3005
R12305 gnd.n6895 gnd.n6894 9.3005
R12306 gnd.n810 gnd.n809 9.3005
R12307 gnd.n6908 gnd.n6907 9.3005
R12308 gnd.n6909 gnd.n808 9.3005
R12309 gnd.n6911 gnd.n6910 9.3005
R12310 gnd.n795 gnd.n794 9.3005
R12311 gnd.n6924 gnd.n6923 9.3005
R12312 gnd.n6925 gnd.n793 9.3005
R12313 gnd.n6927 gnd.n6926 9.3005
R12314 gnd.n779 gnd.n778 9.3005
R12315 gnd.n6940 gnd.n6939 9.3005
R12316 gnd.n6941 gnd.n777 9.3005
R12317 gnd.n6943 gnd.n6942 9.3005
R12318 gnd.n763 gnd.n762 9.3005
R12319 gnd.n6956 gnd.n6955 9.3005
R12320 gnd.n6957 gnd.n761 9.3005
R12321 gnd.n6959 gnd.n6958 9.3005
R12322 gnd.n746 gnd.n745 9.3005
R12323 gnd.n6972 gnd.n6971 9.3005
R12324 gnd.n6973 gnd.n744 9.3005
R12325 gnd.n6975 gnd.n6974 9.3005
R12326 gnd.n732 gnd.n731 9.3005
R12327 gnd.n6988 gnd.n6987 9.3005
R12328 gnd.n6989 gnd.n730 9.3005
R12329 gnd.n6991 gnd.n6990 9.3005
R12330 gnd.n716 gnd.n715 9.3005
R12331 gnd.n7004 gnd.n7003 9.3005
R12332 gnd.n7005 gnd.n714 9.3005
R12333 gnd.n7007 gnd.n7006 9.3005
R12334 gnd.n702 gnd.n701 9.3005
R12335 gnd.n7020 gnd.n7019 9.3005
R12336 gnd.n7021 gnd.n700 9.3005
R12337 gnd.n7023 gnd.n7022 9.3005
R12338 gnd.n689 gnd.n688 9.3005
R12339 gnd.n7036 gnd.n7035 9.3005
R12340 gnd.n7037 gnd.n687 9.3005
R12341 gnd.n7039 gnd.n7038 9.3005
R12342 gnd.n675 gnd.n674 9.3005
R12343 gnd.n7052 gnd.n7051 9.3005
R12344 gnd.n7053 gnd.n673 9.3005
R12345 gnd.n7056 gnd.n7055 9.3005
R12346 gnd.n7054 gnd.n659 9.3005
R12347 gnd.n7070 gnd.n658 9.3005
R12348 gnd.n7072 gnd.n7071 9.3005
R12349 gnd.n5798 gnd.n5797 9.3005
R12350 gnd.n5794 gnd.n1101 9.3005
R12351 gnd.n5134 gnd.n1102 9.3005
R12352 gnd.n5137 gnd.n5136 9.3005
R12353 gnd.n5139 gnd.n5138 9.3005
R12354 gnd.n5140 gnd.n5127 9.3005
R12355 gnd.n5142 gnd.n5141 9.3005
R12356 gnd.n5143 gnd.n5126 9.3005
R12357 gnd.n5145 gnd.n5144 9.3005
R12358 gnd.n5146 gnd.n5121 9.3005
R12359 gnd.n5796 gnd.n5795 9.3005
R12360 gnd.n4911 gnd.n1437 9.3005
R12361 gnd.n4915 gnd.n4914 9.3005
R12362 gnd.n4916 gnd.n1435 9.3005
R12363 gnd.n5195 gnd.n5194 9.3005
R12364 gnd.n5193 gnd.n1436 9.3005
R12365 gnd.n5192 gnd.n5191 9.3005
R12366 gnd.n5190 gnd.n4917 9.3005
R12367 gnd.n5189 gnd.n5188 9.3005
R12368 gnd.n5187 gnd.n4920 9.3005
R12369 gnd.n5186 gnd.n5185 9.3005
R12370 gnd.n5184 gnd.n4921 9.3005
R12371 gnd.n5183 gnd.n5182 9.3005
R12372 gnd.n5181 gnd.n4924 9.3005
R12373 gnd.n5180 gnd.n5179 9.3005
R12374 gnd.n5178 gnd.n4925 9.3005
R12375 gnd.n5177 gnd.n5176 9.3005
R12376 gnd.n5175 gnd.n4928 9.3005
R12377 gnd.n5174 gnd.n5173 9.3005
R12378 gnd.n5172 gnd.n4929 9.3005
R12379 gnd.n5171 gnd.n5170 9.3005
R12380 gnd.n5169 gnd.n4932 9.3005
R12381 gnd.n5168 gnd.n5167 9.3005
R12382 gnd.n5166 gnd.n4933 9.3005
R12383 gnd.n5165 gnd.n5164 9.3005
R12384 gnd.n5163 gnd.n4936 9.3005
R12385 gnd.n5162 gnd.n5161 9.3005
R12386 gnd.n5160 gnd.n4937 9.3005
R12387 gnd.n5159 gnd.n5158 9.3005
R12388 gnd.n5157 gnd.n5120 9.3005
R12389 gnd.n5156 gnd.n5155 9.3005
R12390 gnd.n5154 gnd.n5151 9.3005
R12391 gnd.n5150 gnd.n1174 9.3005
R12392 gnd.n5148 gnd.n5147 9.3005
R12393 gnd.n1170 gnd.n1169 9.3005
R12394 gnd.n5747 gnd.n5746 9.3005
R12395 gnd.n5749 gnd.n5748 9.3005
R12396 gnd.n1158 gnd.n1157 9.3005
R12397 gnd.n5755 gnd.n5754 9.3005
R12398 gnd.n5757 gnd.n5756 9.3005
R12399 gnd.n1150 gnd.n1149 9.3005
R12400 gnd.n5763 gnd.n5762 9.3005
R12401 gnd.n5765 gnd.n5764 9.3005
R12402 gnd.n1140 gnd.n1139 9.3005
R12403 gnd.n5771 gnd.n5770 9.3005
R12404 gnd.n5773 gnd.n5772 9.3005
R12405 gnd.n1132 gnd.n1131 9.3005
R12406 gnd.n5779 gnd.n5778 9.3005
R12407 gnd.n5781 gnd.n5780 9.3005
R12408 gnd.n1122 gnd.n1120 9.3005
R12409 gnd.n5787 gnd.n5786 9.3005
R12410 gnd.n5788 gnd.n1119 9.3005
R12411 gnd.n5356 gnd.n5355 9.3005
R12412 gnd.n1123 gnd.n1121 9.3005
R12413 gnd.n5785 gnd.n5784 9.3005
R12414 gnd.n5783 gnd.n5782 9.3005
R12415 gnd.n1127 gnd.n1126 9.3005
R12416 gnd.n5777 gnd.n5776 9.3005
R12417 gnd.n5775 gnd.n5774 9.3005
R12418 gnd.n1136 gnd.n1135 9.3005
R12419 gnd.n5769 gnd.n5768 9.3005
R12420 gnd.n5767 gnd.n5766 9.3005
R12421 gnd.n1144 gnd.n1143 9.3005
R12422 gnd.n5761 gnd.n5760 9.3005
R12423 gnd.n5759 gnd.n5758 9.3005
R12424 gnd.n1154 gnd.n1153 9.3005
R12425 gnd.n5753 gnd.n5752 9.3005
R12426 gnd.n5751 gnd.n5750 9.3005
R12427 gnd.n1164 gnd.n1163 9.3005
R12428 gnd.n5745 gnd.n5744 9.3005
R12429 gnd.n5655 gnd.n5357 9.3005
R12430 gnd.n5654 gnd.n5653 9.3005
R12431 gnd.n5652 gnd.n5360 9.3005
R12432 gnd.n5651 gnd.n5650 9.3005
R12433 gnd.n5649 gnd.n5361 9.3005
R12434 gnd.n5648 gnd.n5647 9.3005
R12435 gnd.n5646 gnd.n5364 9.3005
R12436 gnd.n5645 gnd.n5644 9.3005
R12437 gnd.n5643 gnd.n5365 9.3005
R12438 gnd.n5642 gnd.n5641 9.3005
R12439 gnd.n5640 gnd.n5368 9.3005
R12440 gnd.n5639 gnd.n5638 9.3005
R12441 gnd.n5637 gnd.n5369 9.3005
R12442 gnd.n5636 gnd.n5635 9.3005
R12443 gnd.n5634 gnd.n5372 9.3005
R12444 gnd.n5633 gnd.n5632 9.3005
R12445 gnd.n5631 gnd.n5373 9.3005
R12446 gnd.n5630 gnd.n5629 9.3005
R12447 gnd.n5628 gnd.n5376 9.3005
R12448 gnd.n5627 gnd.n5626 9.3005
R12449 gnd.n5625 gnd.n5377 9.3005
R12450 gnd.n5624 gnd.n5623 9.3005
R12451 gnd.n1008 gnd.n1007 9.3005
R12452 gnd.n5902 gnd.n5901 9.3005
R12453 gnd.n5903 gnd.n1005 9.3005
R12454 gnd.n5905 gnd.n5904 9.3005
R12455 gnd.n5906 gnd.n1004 9.3005
R12456 gnd.n5910 gnd.n5909 9.3005
R12457 gnd.n5911 gnd.n1002 9.3005
R12458 gnd.n5960 gnd.n5959 9.3005
R12459 gnd.n5958 gnd.n1003 9.3005
R12460 gnd.n5957 gnd.n5956 9.3005
R12461 gnd.n5955 gnd.n5912 9.3005
R12462 gnd.n5954 gnd.n5953 9.3005
R12463 gnd.n5952 gnd.n5946 9.3005
R12464 gnd.n5951 gnd.n5950 9.3005
R12465 gnd.n5949 gnd.n5947 9.3005
R12466 gnd.n906 gnd.n905 9.3005
R12467 gnd.n6082 gnd.n6081 9.3005
R12468 gnd.n6083 gnd.n903 9.3005
R12469 gnd.n6085 gnd.n6084 9.3005
R12470 gnd.n6086 gnd.n902 9.3005
R12471 gnd.n6089 gnd.n6088 9.3005
R12472 gnd.n6090 gnd.n900 9.3005
R12473 gnd.n6818 gnd.n6817 9.3005
R12474 gnd.n6816 gnd.n901 9.3005
R12475 gnd.n6815 gnd.n6814 9.3005
R12476 gnd.n6813 gnd.n6091 9.3005
R12477 gnd.n6812 gnd.n6811 9.3005
R12478 gnd.n6810 gnd.n6094 9.3005
R12479 gnd.n6809 gnd.n6808 9.3005
R12480 gnd.n6807 gnd.n6095 9.3005
R12481 gnd.n6806 gnd.n6805 9.3005
R12482 gnd.n6804 gnd.n6098 9.3005
R12483 gnd.n6803 gnd.n6802 9.3005
R12484 gnd.n6801 gnd.n6099 9.3005
R12485 gnd.n6800 gnd.n6799 9.3005
R12486 gnd.n6798 gnd.n6102 9.3005
R12487 gnd.n6797 gnd.n6796 9.3005
R12488 gnd.n6795 gnd.n6103 9.3005
R12489 gnd.n6794 gnd.n6793 9.3005
R12490 gnd.n6792 gnd.n6106 9.3005
R12491 gnd.n6791 gnd.n6790 9.3005
R12492 gnd.n6789 gnd.n6107 9.3005
R12493 gnd.n6788 gnd.n6787 9.3005
R12494 gnd.n6786 gnd.n6110 9.3005
R12495 gnd.n6785 gnd.n6784 9.3005
R12496 gnd.n6783 gnd.n6111 9.3005
R12497 gnd.n6782 gnd.n6781 9.3005
R12498 gnd.n6780 gnd.n6114 9.3005
R12499 gnd.n6779 gnd.n6778 9.3005
R12500 gnd.n6777 gnd.n6115 9.3005
R12501 gnd.n6776 gnd.n6775 9.3005
R12502 gnd.n6774 gnd.n6118 9.3005
R12503 gnd.n6773 gnd.n6772 9.3005
R12504 gnd.n6771 gnd.n6119 9.3005
R12505 gnd.n6770 gnd.n6769 9.3005
R12506 gnd.n6768 gnd.n6122 9.3005
R12507 gnd.n6767 gnd.n6766 9.3005
R12508 gnd.n6765 gnd.n6123 9.3005
R12509 gnd.n6764 gnd.n6763 9.3005
R12510 gnd.n6762 gnd.n6575 9.3005
R12511 gnd.n6761 gnd.n6760 9.3005
R12512 gnd.n6759 gnd.n6576 9.3005
R12513 gnd.n6758 gnd.n6757 9.3005
R12514 gnd.n6756 gnd.n6580 9.3005
R12515 gnd.n6755 gnd.n6754 9.3005
R12516 gnd.n6753 gnd.n6581 9.3005
R12517 gnd.n6752 gnd.n6751 9.3005
R12518 gnd.n6750 gnd.n6584 9.3005
R12519 gnd.n6749 gnd.n6748 9.3005
R12520 gnd.n6747 gnd.n6585 9.3005
R12521 gnd.n6746 gnd.n6745 9.3005
R12522 gnd.n6744 gnd.n6588 9.3005
R12523 gnd.n6743 gnd.n6742 9.3005
R12524 gnd.n6741 gnd.n6589 9.3005
R12525 gnd.n6740 gnd.n6739 9.3005
R12526 gnd.n6738 gnd.n6592 9.3005
R12527 gnd.n6737 gnd.n6736 9.3005
R12528 gnd.n6735 gnd.n6593 9.3005
R12529 gnd.n6734 gnd.n6595 9.3005
R12530 gnd.n5657 gnd.n5656 9.3005
R12531 gnd.n7259 gnd.n7258 9.3005
R12532 gnd.n484 gnd.n483 9.3005
R12533 gnd.n7272 gnd.n7271 9.3005
R12534 gnd.n7273 gnd.n482 9.3005
R12535 gnd.n7275 gnd.n7274 9.3005
R12536 gnd.n466 gnd.n465 9.3005
R12537 gnd.n7288 gnd.n7287 9.3005
R12538 gnd.n7289 gnd.n464 9.3005
R12539 gnd.n7291 gnd.n7290 9.3005
R12540 gnd.n449 gnd.n448 9.3005
R12541 gnd.n7304 gnd.n7303 9.3005
R12542 gnd.n7305 gnd.n446 9.3005
R12543 gnd.n7313 gnd.n7312 9.3005
R12544 gnd.n7311 gnd.n447 9.3005
R12545 gnd.n7310 gnd.n7309 9.3005
R12546 gnd.n7308 gnd.n7306 9.3005
R12547 gnd.n413 gnd.n411 9.3005
R12548 gnd.n7389 gnd.n7388 9.3005
R12549 gnd.n7387 gnd.n412 9.3005
R12550 gnd.n7386 gnd.n7385 9.3005
R12551 gnd.n7384 gnd.n414 9.3005
R12552 gnd.n381 gnd.n379 9.3005
R12553 gnd.n7436 gnd.n7435 9.3005
R12554 gnd.n7434 gnd.n380 9.3005
R12555 gnd.n7433 gnd.n7432 9.3005
R12556 gnd.n7431 gnd.n382 9.3005
R12557 gnd.n7430 gnd.n7429 9.3005
R12558 gnd.n319 gnd.n317 9.3005
R12559 gnd.n7582 gnd.n7581 9.3005
R12560 gnd.n7580 gnd.n318 9.3005
R12561 gnd.n7579 gnd.n7578 9.3005
R12562 gnd.n7577 gnd.n320 9.3005
R12563 gnd.n7576 gnd.n7575 9.3005
R12564 gnd.n7574 gnd.n324 9.3005
R12565 gnd.n7573 gnd.n7572 9.3005
R12566 gnd.n7571 gnd.n325 9.3005
R12567 gnd.n296 gnd.n295 9.3005
R12568 gnd.n7596 gnd.n7595 9.3005
R12569 gnd.n7597 gnd.n294 9.3005
R12570 gnd.n7599 gnd.n7598 9.3005
R12571 gnd.n280 gnd.n279 9.3005
R12572 gnd.n7612 gnd.n7611 9.3005
R12573 gnd.n7613 gnd.n278 9.3005
R12574 gnd.n7615 gnd.n7614 9.3005
R12575 gnd.n266 gnd.n265 9.3005
R12576 gnd.n7628 gnd.n7627 9.3005
R12577 gnd.n7629 gnd.n264 9.3005
R12578 gnd.n7631 gnd.n7630 9.3005
R12579 gnd.n250 gnd.n249 9.3005
R12580 gnd.n7644 gnd.n7643 9.3005
R12581 gnd.n7645 gnd.n248 9.3005
R12582 gnd.n7647 gnd.n7646 9.3005
R12583 gnd.n236 gnd.n235 9.3005
R12584 gnd.n7660 gnd.n7659 9.3005
R12585 gnd.n7661 gnd.n234 9.3005
R12586 gnd.n7663 gnd.n7662 9.3005
R12587 gnd.n221 gnd.n220 9.3005
R12588 gnd.n7676 gnd.n7675 9.3005
R12589 gnd.n7677 gnd.n218 9.3005
R12590 gnd.n7747 gnd.n7746 9.3005
R12591 gnd.n7745 gnd.n219 9.3005
R12592 gnd.n7744 gnd.n7743 9.3005
R12593 gnd.n7742 gnd.n7678 9.3005
R12594 gnd.n7741 gnd.n7740 9.3005
R12595 gnd.n7257 gnd.n500 9.3005
R12596 gnd.n7737 gnd.n7680 9.3005
R12597 gnd.n7736 gnd.n7735 9.3005
R12598 gnd.n7734 gnd.n7685 9.3005
R12599 gnd.n7733 gnd.n7732 9.3005
R12600 gnd.n7731 gnd.n7686 9.3005
R12601 gnd.n7730 gnd.n7729 9.3005
R12602 gnd.n7728 gnd.n7693 9.3005
R12603 gnd.n7727 gnd.n7726 9.3005
R12604 gnd.n7725 gnd.n7694 9.3005
R12605 gnd.n7724 gnd.n7723 9.3005
R12606 gnd.n7722 gnd.n7701 9.3005
R12607 gnd.n7721 gnd.n7720 9.3005
R12608 gnd.n7719 gnd.n7702 9.3005
R12609 gnd.n7718 gnd.n7717 9.3005
R12610 gnd.n7716 gnd.n7709 9.3005
R12611 gnd.n7715 gnd.n7714 9.3005
R12612 gnd.n124 gnd.n121 9.3005
R12613 gnd.n7841 gnd.n7840 9.3005
R12614 gnd.n7739 gnd.n7738 9.3005
R12615 gnd.n7172 gnd.n582 9.3005
R12616 gnd.n7171 gnd.n7170 9.3005
R12617 gnd.n7169 gnd.n584 9.3005
R12618 gnd.n7168 gnd.n7167 9.3005
R12619 gnd.n7166 gnd.n587 9.3005
R12620 gnd.n7165 gnd.n7164 9.3005
R12621 gnd.n7163 gnd.n588 9.3005
R12622 gnd.n7162 gnd.n7161 9.3005
R12623 gnd.n7160 gnd.n591 9.3005
R12624 gnd.n7159 gnd.n7158 9.3005
R12625 gnd.n7157 gnd.n592 9.3005
R12626 gnd.n7156 gnd.n7155 9.3005
R12627 gnd.n7154 gnd.n7153 9.3005
R12628 gnd.n428 gnd.n427 9.3005
R12629 gnd.n7328 gnd.n7327 9.3005
R12630 gnd.n7329 gnd.n425 9.3005
R12631 gnd.n7339 gnd.n7338 9.3005
R12632 gnd.n7337 gnd.n426 9.3005
R12633 gnd.n7336 gnd.n7335 9.3005
R12634 gnd.n7334 gnd.n7331 9.3005
R12635 gnd.n7330 gnd.n388 9.3005
R12636 gnd.n7417 gnd.n387 9.3005
R12637 gnd.n7419 gnd.n7418 9.3005
R12638 gnd.n7420 gnd.n385 9.3005
R12639 gnd.n7423 gnd.n7422 9.3005
R12640 gnd.n7421 gnd.n386 9.3005
R12641 gnd.n354 gnd.n353 9.3005
R12642 gnd.n7542 gnd.n7541 9.3005
R12643 gnd.n7543 gnd.n352 9.3005
R12644 gnd.n7545 gnd.n7544 9.3005
R12645 gnd.n7546 gnd.n79 9.3005
R12646 gnd.n7890 gnd.n80 9.3005
R12647 gnd.n7889 gnd.n7888 9.3005
R12648 gnd.n7887 gnd.n81 9.3005
R12649 gnd.n7886 gnd.n7885 9.3005
R12650 gnd.n7884 gnd.n85 9.3005
R12651 gnd.n7883 gnd.n7882 9.3005
R12652 gnd.n7881 gnd.n86 9.3005
R12653 gnd.n7880 gnd.n7879 9.3005
R12654 gnd.n7878 gnd.n90 9.3005
R12655 gnd.n7877 gnd.n7876 9.3005
R12656 gnd.n7875 gnd.n91 9.3005
R12657 gnd.n7874 gnd.n7873 9.3005
R12658 gnd.n7872 gnd.n95 9.3005
R12659 gnd.n7871 gnd.n7870 9.3005
R12660 gnd.n7869 gnd.n96 9.3005
R12661 gnd.n7868 gnd.n7867 9.3005
R12662 gnd.n7866 gnd.n100 9.3005
R12663 gnd.n7865 gnd.n7864 9.3005
R12664 gnd.n7863 gnd.n101 9.3005
R12665 gnd.n7862 gnd.n7861 9.3005
R12666 gnd.n7860 gnd.n105 9.3005
R12667 gnd.n7859 gnd.n7858 9.3005
R12668 gnd.n7857 gnd.n106 9.3005
R12669 gnd.n7856 gnd.n7855 9.3005
R12670 gnd.n7854 gnd.n110 9.3005
R12671 gnd.n7853 gnd.n7852 9.3005
R12672 gnd.n7851 gnd.n111 9.3005
R12673 gnd.n7850 gnd.n7849 9.3005
R12674 gnd.n7848 gnd.n115 9.3005
R12675 gnd.n7847 gnd.n7846 9.3005
R12676 gnd.n7845 gnd.n116 9.3005
R12677 gnd.n7844 gnd.n7843 9.3005
R12678 gnd.n7842 gnd.n120 9.3005
R12679 gnd.n7174 gnd.n7173 9.3005
R12680 gnd.t11 gnd.n3160 9.24152
R12681 gnd.n3062 gnd.t228 9.24152
R12682 gnd.n4342 gnd.t214 9.24152
R12683 gnd.t77 gnd.n1501 9.24152
R12684 gnd.n262 gnd.t81 9.24152
R12685 gnd.t108 gnd.t11 8.92286
R12686 gnd.n5621 gnd.t255 8.92286
R12687 gnd.n5890 gnd.n1020 8.92286
R12688 gnd.n1011 gnd.t245 8.92286
R12689 gnd.t68 gnd.n5386 8.92286
R12690 gnd.n6079 gnd.n909 8.92286
R12691 gnd.n6821 gnd.n6820 8.92286
R12692 gnd.n6889 gnd.n830 8.92286
R12693 gnd.n6913 gnd.n805 8.92286
R12694 gnd.t337 gnd.n6145 8.92286
R12695 gnd.n6136 gnd.n6135 8.92286
R12696 gnd.n6565 gnd.t238 8.92286
R12697 gnd.n4312 gnd.n4287 8.92171
R12698 gnd.n4280 gnd.n4255 8.92171
R12699 gnd.n4248 gnd.n4223 8.92171
R12700 gnd.n4217 gnd.n4192 8.92171
R12701 gnd.n4185 gnd.n4160 8.92171
R12702 gnd.n4153 gnd.n4128 8.92171
R12703 gnd.n4121 gnd.n4096 8.92171
R12704 gnd.n4090 gnd.n4065 8.92171
R12705 gnd.n6425 gnd.n6407 8.72777
R12706 gnd.n3816 gnd.t45 8.60421
R12707 gnd.t130 gnd.n1533 8.60421
R12708 gnd.n7492 gnd.t88 8.60421
R12709 gnd.n3240 gnd.n3220 8.43467
R12710 gnd.n58 gnd.n38 8.43467
R12711 gnd.n4909 gnd.n0 8.41456
R12712 gnd.n7891 gnd.n7890 8.41456
R12713 gnd.n4313 gnd.n4285 8.14595
R12714 gnd.n4281 gnd.n4253 8.14595
R12715 gnd.n4249 gnd.n4221 8.14595
R12716 gnd.n4218 gnd.n4190 8.14595
R12717 gnd.n4186 gnd.n4158 8.14595
R12718 gnd.n4154 gnd.n4126 8.14595
R12719 gnd.n4122 gnd.n4094 8.14595
R12720 gnd.n4091 gnd.n4063 8.14595
R12721 gnd.n4318 gnd.n4317 7.97301
R12722 gnd.t322 gnd.n3331 7.9669
R12723 gnd.n3061 gnd.n1645 7.9669
R12724 gnd.n5791 gnd.n1104 7.9669
R12725 gnd.n7078 gnd.n7076 7.9669
R12726 gnd.n7840 gnd.n124 7.75808
R12727 gnd.n6688 gnd.n6684 7.75808
R12728 gnd.n5744 gnd.n1163 7.75808
R12729 gnd.n4512 gnd.n4451 7.75808
R12730 gnd.t228 gnd.n3061 7.64824
R12731 gnd.n3052 gnd.n1395 7.64824
R12732 gnd.n5232 gnd.n1406 7.64824
R12733 gnd.n5227 gnd.n5226 7.64824
R12734 gnd.n1421 gnd.n1412 7.64824
R12735 gnd.n5220 gnd.n1422 7.64824
R12736 gnd.n5219 gnd.n1425 7.64824
R12737 gnd.n5197 gnd.n1377 7.64824
R12738 gnd.n5246 gnd.n1380 7.64824
R12739 gnd.n4993 gnd.n4992 7.64824
R12740 gnd.n5254 gnd.n1371 7.64824
R12741 gnd.n4997 gnd.n1360 7.64824
R12742 gnd.n5262 gnd.n1363 7.64824
R12743 gnd.n5003 gnd.n1351 7.64824
R12744 gnd.n5270 gnd.n1354 7.64824
R12745 gnd.n5007 gnd.n1342 7.64824
R12746 gnd.n5278 gnd.n1345 7.64824
R12747 gnd.n5034 gnd.n5033 7.64824
R12748 gnd.n5286 gnd.n1336 7.64824
R12749 gnd.n5027 gnd.n1325 7.64824
R12750 gnd.n5294 gnd.n1328 7.64824
R12751 gnd.n5023 gnd.n1316 7.64824
R12752 gnd.n5302 gnd.n1319 7.64824
R12753 gnd.n5019 gnd.n1307 7.64824
R12754 gnd.n5310 gnd.n1310 7.64824
R12755 gnd.n5097 gnd.n5096 7.64824
R12756 gnd.n5318 gnd.n1301 7.64824
R12757 gnd.n5103 gnd.n1290 7.64824
R12758 gnd.n5326 gnd.n1293 7.64824
R12759 gnd.n5107 gnd.n1281 7.64824
R12760 gnd.n5334 gnd.n1284 7.64824
R12761 gnd.n5118 gnd.n1271 7.64824
R12762 gnd.n5344 gnd.n1274 7.64824
R12763 gnd.n5664 gnd.n1175 7.64824
R12764 gnd.n5741 gnd.n1177 7.64824
R12765 gnd.n5880 gnd.n1028 7.64824
R12766 gnd.n6069 gnd.n919 7.64824
R12767 gnd.t294 gnd.n870 7.64824
R12768 gnd.n6223 gnd.n6215 7.64824
R12769 gnd.n6881 gnd.n838 7.64824
R12770 gnd.n6261 gnd.t25 7.64824
R12771 gnd.n6921 gnd.n797 7.64824
R12772 gnd.n7176 gnd.n581 7.64824
R12773 gnd.n7261 gnd.n495 7.64824
R12774 gnd.n7269 gnd.n486 7.64824
R12775 gnd.n607 gnd.n489 7.64824
R12776 gnd.n7277 gnd.n477 7.64824
R12777 gnd.n611 gnd.n480 7.64824
R12778 gnd.n7285 gnd.n468 7.64824
R12779 gnd.n617 gnd.n471 7.64824
R12780 gnd.n7293 gnd.n460 7.64824
R12781 gnd.n7128 gnd.n7127 7.64824
R12782 gnd.n7301 gnd.n451 7.64824
R12783 gnd.n7151 gnd.n454 7.64824
R12784 gnd.n7315 gnd.n440 7.64824
R12785 gnd.n7145 gnd.n443 7.64824
R12786 gnd.n7325 gnd.n430 7.64824
R12787 gnd.n432 gnd.n422 7.64824
R12788 gnd.n7342 gnd.n7341 7.64824
R12789 gnd.n7391 gnd.n405 7.64824
R12790 gnd.n7332 gnd.n408 7.64824
R12791 gnd.n7401 gnd.n396 7.64824
R12792 gnd.n7382 gnd.n7381 7.64824
R12793 gnd.n7415 gnd.n390 7.64824
R12794 gnd.n7438 gnd.n373 7.64824
R12795 gnd.n7409 gnd.n376 7.64824
R12796 gnd.n7425 gnd.n383 7.64824
R12797 gnd.n7447 gnd.n362 7.64824
R12798 gnd.n7427 gnd.n364 7.64824
R12799 gnd.n7539 gnd.n356 7.64824
R12800 gnd.n7584 gnd.n311 7.64824
R12801 gnd.n7533 gnd.n314 7.64824
R12802 gnd.n7549 gnd.n348 7.64824
R12803 gnd.n7548 gnd.n343 7.64824
R12804 gnd.n7556 gnd.n7555 7.64824
R12805 gnd.n345 gnd.n333 7.64824
R12806 gnd.n3725 gnd.t15 7.32958
R12807 gnd.n5808 gnd.t224 7.32958
R12808 gnd.n1064 gnd.t339 7.32958
R12809 gnd.t66 gnd.n1028 7.32958
R12810 gnd.n6572 gnd.t295 7.32958
R12811 gnd.n7025 gnd.t362 7.32958
R12812 gnd.n671 gnd.t192 7.32958
R12813 gnd.n5420 gnd.n5419 7.30353
R12814 gnd.n6424 gnd.n6423 7.30353
R12815 gnd.n3685 gnd.n3404 7.01093
R12816 gnd.n3407 gnd.n3405 7.01093
R12817 gnd.n3695 gnd.n3694 7.01093
R12818 gnd.n3706 gnd.n3388 7.01093
R12819 gnd.n3705 gnd.n3391 7.01093
R12820 gnd.n3716 gnd.n3379 7.01093
R12821 gnd.n3382 gnd.n3380 7.01093
R12822 gnd.n3726 gnd.n3725 7.01093
R12823 gnd.n3736 gnd.n3360 7.01093
R12824 gnd.n3735 gnd.n3363 7.01093
R12825 gnd.n3744 gnd.n3354 7.01093
R12826 gnd.n3756 gnd.n3344 7.01093
R12827 gnd.n3766 gnd.n3329 7.01093
R12828 gnd.n3782 gnd.n3781 7.01093
R12829 gnd.n3331 gnd.n3268 7.01093
R12830 gnd.n3836 gnd.n3269 7.01093
R12831 gnd.n3830 gnd.n3829 7.01093
R12832 gnd.n3318 gnd.n3280 7.01093
R12833 gnd.n3822 gnd.n3291 7.01093
R12834 gnd.n3309 gnd.n3304 7.01093
R12835 gnd.n3816 gnd.n3815 7.01093
R12836 gnd.n3862 gnd.n3195 7.01093
R12837 gnd.n3861 gnd.n3860 7.01093
R12838 gnd.n3873 gnd.n3872 7.01093
R12839 gnd.n3188 gnd.n3180 7.01093
R12840 gnd.n3902 gnd.n3168 7.01093
R12841 gnd.n3901 gnd.n3171 7.01093
R12842 gnd.n3912 gnd.n3160 7.01093
R12843 gnd.n3161 gnd.n3149 7.01093
R12844 gnd.n3923 gnd.n3150 7.01093
R12845 gnd.n3947 gnd.n3141 7.01093
R12846 gnd.n3946 gnd.n3132 7.01093
R12847 gnd.n3969 gnd.n3968 7.01093
R12848 gnd.n3987 gnd.n3113 7.01093
R12849 gnd.n3986 gnd.n3116 7.01093
R12850 gnd.n3997 gnd.n3105 7.01093
R12851 gnd.n3106 gnd.n3093 7.01093
R12852 gnd.n4008 gnd.n3094 7.01093
R12853 gnd.n4035 gnd.n3078 7.01093
R12854 gnd.n4047 gnd.n4046 7.01093
R12855 gnd.n4029 gnd.n3071 7.01093
R12856 gnd.n4058 gnd.n4057 7.01093
R12857 gnd.n4330 gnd.n1653 7.01093
R12858 gnd.n4329 gnd.n3062 7.01093
R12859 gnd.n4342 gnd.n1645 7.01093
R12860 gnd.n1646 gnd.n1638 7.01093
R12861 gnd.n4352 gnd.n1564 7.01093
R12862 gnd.n5907 gnd.t152 7.01093
R12863 gnd.t331 gnd.n877 7.01093
R12864 gnd.n6271 gnd.t329 7.01093
R12865 gnd.t335 gnd.n6149 7.01093
R12866 gnd.n3363 gnd.t49 6.69227
R12867 gnd.n3171 gnd.t108 6.69227
R12868 gnd.n4036 gnd.t46 6.69227
R12869 gnd.n6827 gnd.t359 6.69227
R12870 gnd.t100 gnd.n820 6.69227
R12871 gnd.n6505 gnd.n6504 6.5566
R12872 gnd.n5525 gnd.n5524 6.5566
R12873 gnd.n5537 gnd.n5440 6.5566
R12874 gnd.n6485 gnd.n6393 6.5566
R12875 gnd.n5872 gnd.n1035 6.37362
R12876 gnd.t255 gnd.t241 6.37362
R12877 gnd.n6021 gnd.n939 6.37362
R12878 gnd.n6833 gnd.t65 6.37362
R12879 gnd.n6233 gnd.n6232 6.37362
R12880 gnd.n6873 gnd.n846 6.37362
R12881 gnd.n6280 gnd.t330 6.37362
R12882 gnd.n6929 gnd.n789 6.37362
R12883 gnd.n6135 gnd.t185 6.37362
R12884 gnd.n6367 gnd.t185 6.37362
R12885 gnd.n6565 gnd.n718 6.37362
R12886 gnd.n5136 gnd.n5133 6.20656
R12887 gnd.n7802 gnd.n7799 6.20656
R12888 gnd.n4717 gnd.n4596 6.20656
R12889 gnd.n6669 gnd.n6665 6.20656
R12890 gnd.t148 gnd.n3792 6.05496
R12891 gnd.n3793 gnd.t50 6.05496
R12892 gnd.t292 gnd.n3195 6.05496
R12893 gnd.t34 gnd.n3957 6.05496
R12894 gnd.n6022 gnd.t3 6.05496
R12895 gnd.t332 gnd.t102 6.05496
R12896 gnd.t159 gnd.t114 6.05496
R12897 gnd.t341 gnd.n791 6.05496
R12898 gnd.n4315 gnd.n4285 5.81868
R12899 gnd.n4283 gnd.n4253 5.81868
R12900 gnd.n4251 gnd.n4221 5.81868
R12901 gnd.n4220 gnd.n4190 5.81868
R12902 gnd.n4188 gnd.n4158 5.81868
R12903 gnd.n4156 gnd.n4126 5.81868
R12904 gnd.n4124 gnd.n4094 5.81868
R12905 gnd.n4093 gnd.n4063 5.81868
R12906 gnd.n6360 gnd.t200 5.73631
R12907 gnd.n6498 gnd.n551 5.62001
R12908 gnd.n5531 gnd.n5444 5.62001
R12909 gnd.n5531 gnd.n5442 5.62001
R12910 gnd.n6492 gnd.n551 5.62001
R12911 gnd.n3544 gnd.n3539 5.4308
R12912 gnd.n4360 gnd.n1631 5.4308
R12913 gnd.n3860 gnd.t321 5.41765
R12914 gnd.t16 gnd.n3883 5.41765
R12915 gnd.t21 gnd.n3125 5.41765
R12916 gnd.t26 gnd.n5962 5.09899
R12917 gnd.n6013 gnd.n955 5.09899
R12918 gnd.n6865 gnd.n854 5.09899
R12919 gnd.n6242 gnd.n6202 5.09899
R12920 gnd.n6937 gnd.n781 5.09899
R12921 gnd.t110 gnd.n6154 5.09899
R12922 gnd.n4313 gnd.n4312 5.04292
R12923 gnd.n4281 gnd.n4280 5.04292
R12924 gnd.n4249 gnd.n4248 5.04292
R12925 gnd.n4218 gnd.n4217 5.04292
R12926 gnd.n4186 gnd.n4185 5.04292
R12927 gnd.n4154 gnd.n4153 5.04292
R12928 gnd.n4122 gnd.n4121 5.04292
R12929 gnd.n4091 gnd.n4090 5.04292
R12930 gnd.n3260 gnd.n3259 4.82753
R12931 gnd.n78 gnd.n77 4.82753
R12932 gnd.n3823 gnd.t14 4.78034
R12933 gnd.n3150 gnd.t12 4.78034
R12934 gnd.n5864 gnd.t316 4.78034
R12935 gnd.t221 gnd.n720 4.78034
R12936 gnd.n6578 gnd.t327 4.78034
R12937 gnd.n3265 gnd.n3262 4.74817
R12938 gnd.n3315 gnd.n3201 4.74817
R12939 gnd.n3302 gnd.n3200 4.74817
R12940 gnd.n3199 gnd.n3198 4.74817
R12941 gnd.n3311 gnd.n3262 4.74817
R12942 gnd.n3312 gnd.n3201 4.74817
R12943 gnd.n3314 gnd.n3200 4.74817
R12944 gnd.n3301 gnd.n3199 4.74817
R12945 gnd.n7588 gnd.n7587 4.74817
R12946 gnd.n346 gnd.n307 4.74817
R12947 gnd.n7552 gnd.n306 4.74817
R12948 gnd.n330 gnd.n305 4.74817
R12949 gnd.n7567 gnd.n304 4.74817
R12950 gnd.n7588 gnd.n308 4.74817
R12951 gnd.n7586 gnd.n307 4.74817
R12952 gnd.n347 gnd.n306 4.74817
R12953 gnd.n7553 gnd.n305 4.74817
R12954 gnd.n331 gnd.n304 4.74817
R12955 gnd.n5242 gnd.n5241 4.74817
R12956 gnd.n5229 gnd.n1388 4.74817
R12957 gnd.n1409 gnd.n1387 4.74817
R12958 gnd.n5216 gnd.n1386 4.74817
R12959 gnd.n1385 gnd.n1382 4.74817
R12960 gnd.n5242 gnd.n1389 4.74817
R12961 gnd.n5240 gnd.n1388 4.74817
R12962 gnd.n5230 gnd.n1387 4.74817
R12963 gnd.n1408 gnd.n1386 4.74817
R12964 gnd.n5217 gnd.n1385 4.74817
R12965 gnd.n3240 gnd.n3239 4.7074
R12966 gnd.n58 gnd.n57 4.7074
R12967 gnd.n3260 gnd.n3240 4.65959
R12968 gnd.n78 gnd.n58 4.65959
R12969 gnd.n7220 gnd.n553 4.6132
R12970 gnd.n1225 gnd.n1222 4.6132
R12971 gnd.n6039 gnd.t113 4.46168
R12972 gnd.n6180 gnd.t118 4.46168
R12973 gnd.n6573 gnd.t287 4.46168
R12974 gnd.n6420 gnd.n6407 4.46111
R12975 gnd.n4298 gnd.n4294 4.38594
R12976 gnd.n4266 gnd.n4262 4.38594
R12977 gnd.n4234 gnd.n4230 4.38594
R12978 gnd.n4203 gnd.n4199 4.38594
R12979 gnd.n4171 gnd.n4167 4.38594
R12980 gnd.n4139 gnd.n4135 4.38594
R12981 gnd.n4107 gnd.n4103 4.38594
R12982 gnd.n4076 gnd.n4072 4.38594
R12983 gnd.n4309 gnd.n4287 4.26717
R12984 gnd.n4277 gnd.n4255 4.26717
R12985 gnd.n4245 gnd.n4223 4.26717
R12986 gnd.n4214 gnd.n4192 4.26717
R12987 gnd.n4182 gnd.n4160 4.26717
R12988 gnd.n4150 gnd.n4128 4.26717
R12989 gnd.n4118 gnd.n4096 4.26717
R12990 gnd.n4087 gnd.n4065 4.26717
R12991 gnd.n3767 gnd.t47 4.14303
R12992 gnd.n3997 gnd.t48 4.14303
R12993 gnd.t196 gnd.n1265 4.14303
R12994 gnd.t207 gnd.n498 4.14303
R12995 gnd.n4317 gnd.n4316 4.08274
R12996 gnd.n6506 gnd.n6505 4.05904
R12997 gnd.n5524 gnd.n5523 4.05904
R12998 gnd.n5541 gnd.n5440 4.05904
R12999 gnd.n6486 gnd.n6485 4.05904
R13000 gnd.n19 gnd.n9 3.99943
R13001 gnd.n5400 gnd.n5399 3.82437
R13002 gnd.t241 gnd.n1018 3.82437
R13003 gnd.n6002 gnd.n965 3.82437
R13004 gnd.t117 gnd.n5943 3.82437
R13005 gnd.n6032 gnd.n940 3.82437
R13006 gnd.n6857 gnd.n862 3.82437
R13007 gnd.n6252 gnd.n6251 3.82437
R13008 gnd.n6307 gnd.n6169 3.82437
R13009 gnd.n6316 gnd.t333 3.82437
R13010 gnd.n6945 gnd.n773 3.82437
R13011 gnd.n6367 gnd.t203 3.82437
R13012 gnd.n6993 gnd.n728 3.82437
R13013 gnd.n4317 gnd.n4189 3.70378
R13014 gnd.n3840 gnd.n3261 3.65935
R13015 gnd.n19 gnd.n18 3.60163
R13016 gnd.n4766 gnd.t261 3.50571
R13017 gnd.n5152 gnd.t196 3.50571
R13018 gnd.n601 gnd.t207 3.50571
R13019 gnd.n7757 gnd.t188 3.50571
R13020 gnd.n4308 gnd.n4289 3.49141
R13021 gnd.n4276 gnd.n4257 3.49141
R13022 gnd.n4244 gnd.n4225 3.49141
R13023 gnd.n4213 gnd.n4194 3.49141
R13024 gnd.n4181 gnd.n4162 3.49141
R13025 gnd.n4149 gnd.n4130 3.49141
R13026 gnd.n4117 gnd.n4098 3.49141
R13027 gnd.n4086 gnd.n4067 3.49141
R13028 gnd.n5934 gnd.t0 3.18706
R13029 gnd.t0 gnd.n5924 3.18706
R13030 gnd.t334 gnd.n6159 3.18706
R13031 gnd.n6325 gnd.t334 3.18706
R13032 gnd.t287 gnd.n6572 3.18706
R13033 gnd.n3346 gnd.t47 2.8684
R13034 gnd.t162 gnd.n1421 2.8684
R13035 gnd.n5978 gnd.t5 2.8684
R13036 gnd.n6969 gnd.t111 2.8684
R13037 gnd.t75 gnd.n348 2.8684
R13038 gnd.n3241 gnd.t147 2.82907
R13039 gnd.n3241 gnd.t183 2.82907
R13040 gnd.n3243 gnd.t95 2.82907
R13041 gnd.n3243 gnd.t37 2.82907
R13042 gnd.n3245 gnd.t182 2.82907
R13043 gnd.n3245 gnd.t99 2.82907
R13044 gnd.n3247 gnd.t172 2.82907
R13045 gnd.n3247 gnd.t142 2.82907
R13046 gnd.n3249 gnd.t94 2.82907
R13047 gnd.n3249 gnd.t163 2.82907
R13048 gnd.n3251 gnd.t161 2.82907
R13049 gnd.n3251 gnd.t361 2.82907
R13050 gnd.n3253 gnd.t309 2.82907
R13051 gnd.n3253 gnd.t41 2.82907
R13052 gnd.n3255 gnd.t310 2.82907
R13053 gnd.n3255 gnd.t308 2.82907
R13054 gnd.n3257 gnd.t311 2.82907
R13055 gnd.n3257 gnd.t74 2.82907
R13056 gnd.n3202 gnd.t348 2.82907
R13057 gnd.n3202 gnd.t126 2.82907
R13058 gnd.n3204 gnd.t30 2.82907
R13059 gnd.n3204 gnd.t299 2.82907
R13060 gnd.n3206 gnd.t158 2.82907
R13061 gnd.n3206 gnd.t176 2.82907
R13062 gnd.n3208 gnd.t320 2.82907
R13063 gnd.n3208 gnd.t303 2.82907
R13064 gnd.n3210 gnd.t120 2.82907
R13065 gnd.n3210 gnd.t345 2.82907
R13066 gnd.n3212 gnd.t70 2.82907
R13067 gnd.n3212 gnd.t355 2.82907
R13068 gnd.n3214 gnd.t138 2.82907
R13069 gnd.n3214 gnd.t168 2.82907
R13070 gnd.n3216 gnd.t78 2.82907
R13071 gnd.n3216 gnd.t302 2.82907
R13072 gnd.n3218 gnd.t137 2.82907
R13073 gnd.n3218 gnd.t105 2.82907
R13074 gnd.n3221 gnd.t323 2.82907
R13075 gnd.n3221 gnd.t349 2.82907
R13076 gnd.n3223 gnd.t177 2.82907
R13077 gnd.n3223 gnd.t62 2.82907
R13078 gnd.n3225 gnd.t307 2.82907
R13079 gnd.n3225 gnd.t156 2.82907
R13080 gnd.n3227 gnd.t350 2.82907
R13081 gnd.n3227 gnd.t129 2.82907
R13082 gnd.n3229 gnd.t52 2.82907
R13083 gnd.n3229 gnd.t324 2.82907
R13084 gnd.n3231 gnd.t354 2.82907
R13085 gnd.n3231 gnd.t124 2.82907
R13086 gnd.n3233 gnd.t133 2.82907
R13087 gnd.n3233 gnd.t347 2.82907
R13088 gnd.n3235 gnd.t169 2.82907
R13089 gnd.n3235 gnd.t80 2.82907
R13090 gnd.n3237 gnd.t32 2.82907
R13091 gnd.n3237 gnd.t122 2.82907
R13092 gnd.n75 gnd.t358 2.82907
R13093 gnd.n75 gnd.t315 2.82907
R13094 gnd.n73 gnd.t56 2.82907
R13095 gnd.n73 gnd.t170 2.82907
R13096 gnd.n71 gnd.t141 2.82907
R13097 gnd.n71 gnd.t97 2.82907
R13098 gnd.n69 gnd.t64 2.82907
R13099 gnd.n69 gnd.t326 2.82907
R13100 gnd.n67 gnd.t76 2.82907
R13101 gnd.n67 gnd.t144 2.82907
R13102 gnd.n65 gnd.t106 2.82907
R13103 gnd.n65 gnd.t107 2.82907
R13104 gnd.n63 gnd.t35 2.82907
R13105 gnd.n63 gnd.t18 2.82907
R13106 gnd.n61 gnd.t173 2.82907
R13107 gnd.n61 gnd.t58 2.82907
R13108 gnd.n59 gnd.t39 2.82907
R13109 gnd.n59 gnd.t356 2.82907
R13110 gnd.n36 gnd.t10 2.82907
R13111 gnd.n36 gnd.t140 2.82907
R13112 gnd.n34 gnd.t92 2.82907
R13113 gnd.n34 gnd.t82 2.82907
R13114 gnd.n32 gnd.t71 2.82907
R13115 gnd.n32 gnd.t305 2.82907
R13116 gnd.n30 gnd.t300 2.82907
R13117 gnd.n30 gnd.t85 2.82907
R13118 gnd.n28 gnd.t178 2.82907
R13119 gnd.n28 gnd.t346 2.82907
R13120 gnd.n26 gnd.t54 2.82907
R13121 gnd.n26 gnd.t60 2.82907
R13122 gnd.n24 gnd.t44 2.82907
R13123 gnd.n24 gnd.t139 2.82907
R13124 gnd.n22 gnd.t91 2.82907
R13125 gnd.n22 gnd.t61 2.82907
R13126 gnd.n20 gnd.t72 2.82907
R13127 gnd.n20 gnd.t20 2.82907
R13128 gnd.n55 gnd.t104 2.82907
R13129 gnd.n55 gnd.t136 2.82907
R13130 gnd.n53 gnd.t83 2.82907
R13131 gnd.n53 gnd.t351 2.82907
R13132 gnd.n51 gnd.t43 2.82907
R13133 gnd.n51 gnd.t298 2.82907
R13134 gnd.n49 gnd.t180 2.82907
R13135 gnd.n49 gnd.t314 2.82907
R13136 gnd.n47 gnd.t119 2.82907
R13137 gnd.n47 gnd.t306 2.82907
R13138 gnd.n45 gnd.t304 2.82907
R13139 gnd.n45 gnd.t325 2.82907
R13140 gnd.n43 gnd.t28 2.82907
R13141 gnd.n43 gnd.t134 2.82907
R13142 gnd.n41 gnd.t301 2.82907
R13143 gnd.n41 gnd.t312 2.82907
R13144 gnd.n39 gnd.t179 2.82907
R13145 gnd.n39 gnd.t121 2.82907
R13146 gnd.n4305 gnd.n4304 2.71565
R13147 gnd.n4273 gnd.n4272 2.71565
R13148 gnd.n4241 gnd.n4240 2.71565
R13149 gnd.n4210 gnd.n4209 2.71565
R13150 gnd.n4178 gnd.n4177 2.71565
R13151 gnd.n4146 gnd.n4145 2.71565
R13152 gnd.n4114 gnd.n4113 2.71565
R13153 gnd.n4083 gnd.n4082 2.71565
R13154 gnd.n5621 gnd.n5620 2.54975
R13155 gnd.n5994 gnd.n973 2.54975
R13156 gnd.n5963 gnd.t26 2.54975
R13157 gnd.n933 gnd.n932 2.54975
R13158 gnd.n932 gnd.t338 2.54975
R13159 gnd.n6849 gnd.n870 2.54975
R13160 gnd.n6261 gnd.n6193 2.54975
R13161 gnd.t336 gnd.n6174 2.54975
R13162 gnd.n6298 gnd.n6174 2.54975
R13163 gnd.n6334 gnd.t110 2.54975
R13164 gnd.n6953 gnd.n765 2.54975
R13165 gnd.n6985 gnd.n735 2.54975
R13166 gnd.n3840 gnd.n3262 2.27742
R13167 gnd.n3840 gnd.n3201 2.27742
R13168 gnd.n3840 gnd.n3200 2.27742
R13169 gnd.n3840 gnd.n3199 2.27742
R13170 gnd.n7589 gnd.n7588 2.27742
R13171 gnd.n7589 gnd.n307 2.27742
R13172 gnd.n7589 gnd.n306 2.27742
R13173 gnd.n7589 gnd.n305 2.27742
R13174 gnd.n7589 gnd.n304 2.27742
R13175 gnd.n5243 gnd.n5242 2.27742
R13176 gnd.n5243 gnd.n1388 2.27742
R13177 gnd.n5243 gnd.n1387 2.27742
R13178 gnd.n5243 gnd.n1386 2.27742
R13179 gnd.n5243 gnd.n1385 2.27742
R13180 gnd.n3694 gnd.t271 2.23109
R13181 gnd.n3317 gnd.t14 2.23109
R13182 gnd.t157 gnd.n1363 2.23109
R13183 gnd.t102 gnd.n862 2.23109
R13184 gnd.n6252 gnd.t159 2.23109
R13185 gnd.t17 gnd.n373 2.23109
R13186 gnd.n4301 gnd.n4291 1.93989
R13187 gnd.n4269 gnd.n4259 1.93989
R13188 gnd.n4237 gnd.n4227 1.93989
R13189 gnd.n4206 gnd.n4196 1.93989
R13190 gnd.n4174 gnd.n4164 1.93989
R13191 gnd.n4142 gnd.n4132 1.93989
R13192 gnd.n4110 gnd.n4100 1.93989
R13193 gnd.n4079 gnd.n4069 1.93989
R13194 gnd.n5601 gnd.t211 1.91244
R13195 gnd.n5970 gnd.t152 1.91244
R13196 gnd.n6342 gnd.t335 1.91244
R13197 gnd.t150 gnd.n3705 1.59378
R13198 gnd.n3884 gnd.t16 1.59378
R13199 gnd.n3134 gnd.t21 1.59378
R13200 gnd.n4806 gnd.t73 1.59378
R13201 gnd.t36 gnd.n1328 1.59378
R13202 gnd.n5019 gnd.t146 1.59378
R13203 gnd.n5963 gnd.t343 1.59378
R13204 gnd.n6079 gnd.t318 1.59378
R13205 gnd.n6913 gnd.t1 1.59378
R13206 gnd.n6334 gnd.t115 1.59378
R13207 gnd.n7151 gnd.t19 1.59378
R13208 gnd.t90 gnd.n430 1.59378
R13209 gnd.n7649 gnd.t9 1.59378
R13210 gnd.n5872 gnd.t265 1.27512
R13211 gnd.n5613 gnd.n5612 1.27512
R13212 gnd.n5387 gnd.t68 1.27512
R13213 gnd.n5986 gnd.n981 1.27512
R13214 gnd.n5944 gnd.t117 1.27512
R13215 gnd.n6040 gnd.n6039 1.27512
R13216 gnd.n6841 gnd.n877 1.27512
R13217 gnd.n6271 gnd.n6270 1.27512
R13218 gnd.n6289 gnd.n6180 1.27512
R13219 gnd.t333 gnd.n6164 1.27512
R13220 gnd.n6961 gnd.n757 1.27512
R13221 gnd.n6351 gnd.t337 1.27512
R13222 gnd.n6977 gnd.n742 1.27512
R13223 gnd.n3547 gnd.n3539 1.16414
R13224 gnd.n4363 gnd.n1631 1.16414
R13225 gnd.n4300 gnd.n4293 1.16414
R13226 gnd.n4268 gnd.n4261 1.16414
R13227 gnd.n4236 gnd.n4229 1.16414
R13228 gnd.n4205 gnd.n4198 1.16414
R13229 gnd.n4173 gnd.n4166 1.16414
R13230 gnd.n4141 gnd.n4134 1.16414
R13231 gnd.n4109 gnd.n4102 1.16414
R13232 gnd.n4078 gnd.n4071 1.16414
R13233 gnd.n7220 gnd.n7219 0.970197
R13234 gnd.n5705 gnd.n1222 0.970197
R13235 gnd.n4284 gnd.n4252 0.962709
R13236 gnd.n4316 gnd.n4284 0.962709
R13237 gnd.n4157 gnd.n4125 0.962709
R13238 gnd.n4189 gnd.n4157 0.962709
R13239 gnd.n3793 gnd.t148 0.956468
R13240 gnd.n3958 gnd.t34 0.956468
R13241 gnd.n4848 gnd.t132 0.956468
R13242 gnd.n5007 gnd.t98 0.956468
R13243 gnd.t7 gnd.n1293 0.956468
R13244 gnd.n5374 gnd.n1042 0.956468
R13245 gnd.n7001 gnd.n720 0.956468
R13246 gnd.t86 gnd.n468 0.956468
R13247 gnd.n7401 gnd.t27 0.956468
R13248 gnd.n7617 gnd.t96 0.956468
R13249 gnd.n3252 gnd.n3250 0.773756
R13250 gnd.n70 gnd.n68 0.773756
R13251 gnd.n3259 gnd.n3258 0.773756
R13252 gnd.n3258 gnd.n3256 0.773756
R13253 gnd.n3256 gnd.n3254 0.773756
R13254 gnd.n3254 gnd.n3252 0.773756
R13255 gnd.n3250 gnd.n3248 0.773756
R13256 gnd.n3248 gnd.n3246 0.773756
R13257 gnd.n3246 gnd.n3244 0.773756
R13258 gnd.n3244 gnd.n3242 0.773756
R13259 gnd.n62 gnd.n60 0.773756
R13260 gnd.n64 gnd.n62 0.773756
R13261 gnd.n66 gnd.n64 0.773756
R13262 gnd.n68 gnd.n66 0.773756
R13263 gnd.n72 gnd.n70 0.773756
R13264 gnd.n74 gnd.n72 0.773756
R13265 gnd.n76 gnd.n74 0.773756
R13266 gnd.n77 gnd.n76 0.773756
R13267 gnd gnd.n0 0.70738
R13268 gnd.n2 gnd.n1 0.672012
R13269 gnd.n3 gnd.n2 0.672012
R13270 gnd.n4 gnd.n3 0.672012
R13271 gnd.n5 gnd.n4 0.672012
R13272 gnd.n6 gnd.n5 0.672012
R13273 gnd.n7 gnd.n6 0.672012
R13274 gnd.n8 gnd.n7 0.672012
R13275 gnd.n9 gnd.n8 0.672012
R13276 gnd.n11 gnd.n10 0.672012
R13277 gnd.n12 gnd.n11 0.672012
R13278 gnd.n13 gnd.n12 0.672012
R13279 gnd.n14 gnd.n13 0.672012
R13280 gnd.n15 gnd.n14 0.672012
R13281 gnd.n16 gnd.n15 0.672012
R13282 gnd.n17 gnd.n16 0.672012
R13283 gnd.n18 gnd.n17 0.672012
R13284 gnd.n5613 gnd.t232 0.637812
R13285 gnd.n940 gnd.t167 0.637812
R13286 gnd.n6169 gnd.t166 0.637812
R13287 gnd.n7892 gnd.n7891 0.637193
R13288 gnd.n3220 gnd.n3219 0.573776
R13289 gnd.n3219 gnd.n3217 0.573776
R13290 gnd.n3217 gnd.n3215 0.573776
R13291 gnd.n3215 gnd.n3213 0.573776
R13292 gnd.n3213 gnd.n3211 0.573776
R13293 gnd.n3211 gnd.n3209 0.573776
R13294 gnd.n3209 gnd.n3207 0.573776
R13295 gnd.n3207 gnd.n3205 0.573776
R13296 gnd.n3205 gnd.n3203 0.573776
R13297 gnd.n3239 gnd.n3238 0.573776
R13298 gnd.n3238 gnd.n3236 0.573776
R13299 gnd.n3236 gnd.n3234 0.573776
R13300 gnd.n3234 gnd.n3232 0.573776
R13301 gnd.n3232 gnd.n3230 0.573776
R13302 gnd.n3230 gnd.n3228 0.573776
R13303 gnd.n3228 gnd.n3226 0.573776
R13304 gnd.n3226 gnd.n3224 0.573776
R13305 gnd.n3224 gnd.n3222 0.573776
R13306 gnd.n23 gnd.n21 0.573776
R13307 gnd.n25 gnd.n23 0.573776
R13308 gnd.n27 gnd.n25 0.573776
R13309 gnd.n29 gnd.n27 0.573776
R13310 gnd.n31 gnd.n29 0.573776
R13311 gnd.n33 gnd.n31 0.573776
R13312 gnd.n35 gnd.n33 0.573776
R13313 gnd.n37 gnd.n35 0.573776
R13314 gnd.n38 gnd.n37 0.573776
R13315 gnd.n42 gnd.n40 0.573776
R13316 gnd.n44 gnd.n42 0.573776
R13317 gnd.n46 gnd.n44 0.573776
R13318 gnd.n48 gnd.n46 0.573776
R13319 gnd.n50 gnd.n48 0.573776
R13320 gnd.n52 gnd.n50 0.573776
R13321 gnd.n54 gnd.n52 0.573776
R13322 gnd.n56 gnd.n54 0.573776
R13323 gnd.n57 gnd.n56 0.573776
R13324 gnd.n7589 gnd.n303 0.5435
R13325 gnd.n5243 gnd.n1384 0.5435
R13326 gnd.n4020 gnd.n1635 0.486781
R13327 gnd.n6595 gnd.n501 0.486781
R13328 gnd.n3596 gnd.n3595 0.48678
R13329 gnd.n5658 gnd.n5657 0.485256
R13330 gnd.n4337 gnd.n1589 0.480683
R13331 gnd.n3680 gnd.n3679 0.480683
R13332 gnd.n4514 gnd.n4513 0.477634
R13333 gnd.n4761 gnd.n1562 0.477634
R13334 gnd.n7740 gnd.n7739 0.477634
R13335 gnd.n7842 gnd.n7841 0.477634
R13336 gnd.n7834 gnd.n7833 0.465439
R13337 gnd.n7763 gnd.n7762 0.465439
R13338 gnd.n7180 gnd.n579 0.465439
R13339 gnd.n535 gnd.n492 0.465439
R13340 gnd.n5738 gnd.n5737 0.465439
R13341 gnd.n5669 gnd.n5668 0.465439
R13342 gnd.n4680 gnd.n4675 0.465439
R13343 gnd.n4755 gnd.n4754 0.465439
R13344 gnd.n7073 gnd.n7072 0.451719
R13345 gnd.n5797 gnd.n5796 0.451719
R13346 gnd.n2840 gnd.n1780 0.425805
R13347 gnd.n2477 gnd.n2476 0.425805
R13348 gnd.n7561 gnd.n7560 0.425805
R13349 gnd.n3056 gnd.n3055 0.425805
R13350 gnd.n5139 gnd.n5133 0.388379
R13351 gnd.n4297 gnd.n4296 0.388379
R13352 gnd.n4265 gnd.n4264 0.388379
R13353 gnd.n4233 gnd.n4232 0.388379
R13354 gnd.n4202 gnd.n4201 0.388379
R13355 gnd.n4170 gnd.n4169 0.388379
R13356 gnd.n4138 gnd.n4137 0.388379
R13357 gnd.n4106 gnd.n4105 0.388379
R13358 gnd.n4075 gnd.n4074 0.388379
R13359 gnd.n7803 gnd.n7802 0.388379
R13360 gnd.n4596 gnd.n4592 0.388379
R13361 gnd.n6665 gnd.n6661 0.388379
R13362 gnd.n5660 gnd.n5659 0.378829
R13363 gnd.n7257 gnd.n7256 0.377553
R13364 gnd.n7892 gnd.n19 0.374463
R13365 gnd gnd.n7892 0.367492
R13366 gnd.n3096 gnd.t46 0.319156
R13367 gnd.n4901 gnd.t123 0.319156
R13368 gnd.n5197 gnd.t171 0.319156
R13369 gnd.n7539 gnd.t59 0.319156
R13370 gnd.n7569 gnd.t63 0.319156
R13371 gnd.n3514 gnd.n3492 0.311721
R13372 gnd.n4408 gnd.n4407 0.268793
R13373 gnd.n5150 gnd.n5149 0.247451
R13374 gnd.n7173 gnd.n583 0.247451
R13375 gnd.n4407 gnd.n4406 0.241354
R13376 gnd.n553 gnd.n550 0.229039
R13377 gnd.n556 gnd.n553 0.229039
R13378 gnd.n1225 gnd.n1224 0.229039
R13379 gnd.n1226 gnd.n1225 0.229039
R13380 gnd.n3261 gnd.n0 0.210825
R13381 gnd.n3668 gnd.n3467 0.206293
R13382 gnd.n4314 gnd.n4286 0.155672
R13383 gnd.n4307 gnd.n4286 0.155672
R13384 gnd.n4307 gnd.n4306 0.155672
R13385 gnd.n4306 gnd.n4290 0.155672
R13386 gnd.n4299 gnd.n4290 0.155672
R13387 gnd.n4299 gnd.n4298 0.155672
R13388 gnd.n4282 gnd.n4254 0.155672
R13389 gnd.n4275 gnd.n4254 0.155672
R13390 gnd.n4275 gnd.n4274 0.155672
R13391 gnd.n4274 gnd.n4258 0.155672
R13392 gnd.n4267 gnd.n4258 0.155672
R13393 gnd.n4267 gnd.n4266 0.155672
R13394 gnd.n4250 gnd.n4222 0.155672
R13395 gnd.n4243 gnd.n4222 0.155672
R13396 gnd.n4243 gnd.n4242 0.155672
R13397 gnd.n4242 gnd.n4226 0.155672
R13398 gnd.n4235 gnd.n4226 0.155672
R13399 gnd.n4235 gnd.n4234 0.155672
R13400 gnd.n4219 gnd.n4191 0.155672
R13401 gnd.n4212 gnd.n4191 0.155672
R13402 gnd.n4212 gnd.n4211 0.155672
R13403 gnd.n4211 gnd.n4195 0.155672
R13404 gnd.n4204 gnd.n4195 0.155672
R13405 gnd.n4204 gnd.n4203 0.155672
R13406 gnd.n4187 gnd.n4159 0.155672
R13407 gnd.n4180 gnd.n4159 0.155672
R13408 gnd.n4180 gnd.n4179 0.155672
R13409 gnd.n4179 gnd.n4163 0.155672
R13410 gnd.n4172 gnd.n4163 0.155672
R13411 gnd.n4172 gnd.n4171 0.155672
R13412 gnd.n4155 gnd.n4127 0.155672
R13413 gnd.n4148 gnd.n4127 0.155672
R13414 gnd.n4148 gnd.n4147 0.155672
R13415 gnd.n4147 gnd.n4131 0.155672
R13416 gnd.n4140 gnd.n4131 0.155672
R13417 gnd.n4140 gnd.n4139 0.155672
R13418 gnd.n4123 gnd.n4095 0.155672
R13419 gnd.n4116 gnd.n4095 0.155672
R13420 gnd.n4116 gnd.n4115 0.155672
R13421 gnd.n4115 gnd.n4099 0.155672
R13422 gnd.n4108 gnd.n4099 0.155672
R13423 gnd.n4108 gnd.n4107 0.155672
R13424 gnd.n4092 gnd.n4064 0.155672
R13425 gnd.n4085 gnd.n4064 0.155672
R13426 gnd.n4085 gnd.n4084 0.155672
R13427 gnd.n4084 gnd.n4068 0.155672
R13428 gnd.n4077 gnd.n4068 0.155672
R13429 gnd.n4077 gnd.n4076 0.155672
R13430 gnd.n4439 gnd.n1589 0.152939
R13431 gnd.n4439 gnd.n4438 0.152939
R13432 gnd.n4438 gnd.n4437 0.152939
R13433 gnd.n4437 gnd.n1591 0.152939
R13434 gnd.n1592 gnd.n1591 0.152939
R13435 gnd.n1593 gnd.n1592 0.152939
R13436 gnd.n1594 gnd.n1593 0.152939
R13437 gnd.n1595 gnd.n1594 0.152939
R13438 gnd.n1596 gnd.n1595 0.152939
R13439 gnd.n1597 gnd.n1596 0.152939
R13440 gnd.n1598 gnd.n1597 0.152939
R13441 gnd.n1599 gnd.n1598 0.152939
R13442 gnd.n1600 gnd.n1599 0.152939
R13443 gnd.n1601 gnd.n1600 0.152939
R13444 gnd.n4409 gnd.n1601 0.152939
R13445 gnd.n4409 gnd.n4408 0.152939
R13446 gnd.n3681 gnd.n3680 0.152939
R13447 gnd.n3681 gnd.n3385 0.152939
R13448 gnd.n3709 gnd.n3385 0.152939
R13449 gnd.n3710 gnd.n3709 0.152939
R13450 gnd.n3711 gnd.n3710 0.152939
R13451 gnd.n3712 gnd.n3711 0.152939
R13452 gnd.n3712 gnd.n3357 0.152939
R13453 gnd.n3739 gnd.n3357 0.152939
R13454 gnd.n3740 gnd.n3739 0.152939
R13455 gnd.n3741 gnd.n3740 0.152939
R13456 gnd.n3741 gnd.n3335 0.152939
R13457 gnd.n3770 gnd.n3335 0.152939
R13458 gnd.n3771 gnd.n3770 0.152939
R13459 gnd.n3772 gnd.n3771 0.152939
R13460 gnd.n3773 gnd.n3772 0.152939
R13461 gnd.n3775 gnd.n3773 0.152939
R13462 gnd.n3775 gnd.n3774 0.152939
R13463 gnd.n3774 gnd.n3284 0.152939
R13464 gnd.n3285 gnd.n3284 0.152939
R13465 gnd.n3286 gnd.n3285 0.152939
R13466 gnd.n3305 gnd.n3286 0.152939
R13467 gnd.n3306 gnd.n3305 0.152939
R13468 gnd.n3306 gnd.n3192 0.152939
R13469 gnd.n3865 gnd.n3192 0.152939
R13470 gnd.n3866 gnd.n3865 0.152939
R13471 gnd.n3867 gnd.n3866 0.152939
R13472 gnd.n3868 gnd.n3867 0.152939
R13473 gnd.n3868 gnd.n3165 0.152939
R13474 gnd.n3905 gnd.n3165 0.152939
R13475 gnd.n3906 gnd.n3905 0.152939
R13476 gnd.n3907 gnd.n3906 0.152939
R13477 gnd.n3908 gnd.n3907 0.152939
R13478 gnd.n3908 gnd.n3138 0.152939
R13479 gnd.n3950 gnd.n3138 0.152939
R13480 gnd.n3951 gnd.n3950 0.152939
R13481 gnd.n3952 gnd.n3951 0.152939
R13482 gnd.n3953 gnd.n3952 0.152939
R13483 gnd.n3953 gnd.n3110 0.152939
R13484 gnd.n3990 gnd.n3110 0.152939
R13485 gnd.n3991 gnd.n3990 0.152939
R13486 gnd.n3992 gnd.n3991 0.152939
R13487 gnd.n3993 gnd.n3992 0.152939
R13488 gnd.n3993 gnd.n3083 0.152939
R13489 gnd.n4039 gnd.n3083 0.152939
R13490 gnd.n4040 gnd.n4039 0.152939
R13491 gnd.n4041 gnd.n4040 0.152939
R13492 gnd.n4042 gnd.n4041 0.152939
R13493 gnd.n4042 gnd.n1650 0.152939
R13494 gnd.n4333 gnd.n1650 0.152939
R13495 gnd.n4334 gnd.n4333 0.152939
R13496 gnd.n4335 gnd.n4334 0.152939
R13497 gnd.n4336 gnd.n4335 0.152939
R13498 gnd.n4337 gnd.n4336 0.152939
R13499 gnd.n3679 gnd.n3409 0.152939
R13500 gnd.n3430 gnd.n3409 0.152939
R13501 gnd.n3431 gnd.n3430 0.152939
R13502 gnd.n3437 gnd.n3431 0.152939
R13503 gnd.n3438 gnd.n3437 0.152939
R13504 gnd.n3439 gnd.n3438 0.152939
R13505 gnd.n3439 gnd.n3428 0.152939
R13506 gnd.n3447 gnd.n3428 0.152939
R13507 gnd.n3448 gnd.n3447 0.152939
R13508 gnd.n3449 gnd.n3448 0.152939
R13509 gnd.n3449 gnd.n3426 0.152939
R13510 gnd.n3457 gnd.n3426 0.152939
R13511 gnd.n3458 gnd.n3457 0.152939
R13512 gnd.n3459 gnd.n3458 0.152939
R13513 gnd.n3459 gnd.n3424 0.152939
R13514 gnd.n3467 gnd.n3424 0.152939
R13515 gnd.n4406 gnd.n1606 0.152939
R13516 gnd.n1608 gnd.n1606 0.152939
R13517 gnd.n1609 gnd.n1608 0.152939
R13518 gnd.n1610 gnd.n1609 0.152939
R13519 gnd.n1611 gnd.n1610 0.152939
R13520 gnd.n1612 gnd.n1611 0.152939
R13521 gnd.n1613 gnd.n1612 0.152939
R13522 gnd.n1614 gnd.n1613 0.152939
R13523 gnd.n1615 gnd.n1614 0.152939
R13524 gnd.n1616 gnd.n1615 0.152939
R13525 gnd.n1617 gnd.n1616 0.152939
R13526 gnd.n1618 gnd.n1617 0.152939
R13527 gnd.n1619 gnd.n1618 0.152939
R13528 gnd.n1620 gnd.n1619 0.152939
R13529 gnd.n1621 gnd.n1620 0.152939
R13530 gnd.n1622 gnd.n1621 0.152939
R13531 gnd.n1623 gnd.n1622 0.152939
R13532 gnd.n1624 gnd.n1623 0.152939
R13533 gnd.n1625 gnd.n1624 0.152939
R13534 gnd.n1626 gnd.n1625 0.152939
R13535 gnd.n1627 gnd.n1626 0.152939
R13536 gnd.n1628 gnd.n1627 0.152939
R13537 gnd.n1632 gnd.n1628 0.152939
R13538 gnd.n1633 gnd.n1632 0.152939
R13539 gnd.n1634 gnd.n1633 0.152939
R13540 gnd.n1635 gnd.n1634 0.152939
R13541 gnd.n3842 gnd.n3841 0.152939
R13542 gnd.n3843 gnd.n3842 0.152939
R13543 gnd.n3844 gnd.n3843 0.152939
R13544 gnd.n3845 gnd.n3844 0.152939
R13545 gnd.n3846 gnd.n3845 0.152939
R13546 gnd.n3847 gnd.n3846 0.152939
R13547 gnd.n3847 gnd.n3146 0.152939
R13548 gnd.n3926 gnd.n3146 0.152939
R13549 gnd.n3927 gnd.n3926 0.152939
R13550 gnd.n3928 gnd.n3927 0.152939
R13551 gnd.n3929 gnd.n3928 0.152939
R13552 gnd.n3930 gnd.n3929 0.152939
R13553 gnd.n3931 gnd.n3930 0.152939
R13554 gnd.n3932 gnd.n3931 0.152939
R13555 gnd.n3933 gnd.n3932 0.152939
R13556 gnd.n3934 gnd.n3933 0.152939
R13557 gnd.n3934 gnd.n3090 0.152939
R13558 gnd.n4011 gnd.n3090 0.152939
R13559 gnd.n4012 gnd.n4011 0.152939
R13560 gnd.n4013 gnd.n4012 0.152939
R13561 gnd.n4014 gnd.n4013 0.152939
R13562 gnd.n4015 gnd.n4014 0.152939
R13563 gnd.n4016 gnd.n4015 0.152939
R13564 gnd.n4017 gnd.n4016 0.152939
R13565 gnd.n4018 gnd.n4017 0.152939
R13566 gnd.n4019 gnd.n4018 0.152939
R13567 gnd.n4021 gnd.n4019 0.152939
R13568 gnd.n4021 gnd.n4020 0.152939
R13569 gnd.n3597 gnd.n3596 0.152939
R13570 gnd.n3597 gnd.n3487 0.152939
R13571 gnd.n3612 gnd.n3487 0.152939
R13572 gnd.n3613 gnd.n3612 0.152939
R13573 gnd.n3614 gnd.n3613 0.152939
R13574 gnd.n3614 gnd.n3475 0.152939
R13575 gnd.n3628 gnd.n3475 0.152939
R13576 gnd.n3629 gnd.n3628 0.152939
R13577 gnd.n3630 gnd.n3629 0.152939
R13578 gnd.n3631 gnd.n3630 0.152939
R13579 gnd.n3632 gnd.n3631 0.152939
R13580 gnd.n3633 gnd.n3632 0.152939
R13581 gnd.n3634 gnd.n3633 0.152939
R13582 gnd.n3635 gnd.n3634 0.152939
R13583 gnd.n3636 gnd.n3635 0.152939
R13584 gnd.n3637 gnd.n3636 0.152939
R13585 gnd.n3638 gnd.n3637 0.152939
R13586 gnd.n3639 gnd.n3638 0.152939
R13587 gnd.n3640 gnd.n3639 0.152939
R13588 gnd.n3641 gnd.n3640 0.152939
R13589 gnd.n3642 gnd.n3641 0.152939
R13590 gnd.n3642 gnd.n3341 0.152939
R13591 gnd.n3759 gnd.n3341 0.152939
R13592 gnd.n3760 gnd.n3759 0.152939
R13593 gnd.n3761 gnd.n3760 0.152939
R13594 gnd.n3762 gnd.n3761 0.152939
R13595 gnd.n3762 gnd.n3263 0.152939
R13596 gnd.n3839 gnd.n3263 0.152939
R13597 gnd.n3515 gnd.n3514 0.152939
R13598 gnd.n3516 gnd.n3515 0.152939
R13599 gnd.n3517 gnd.n3516 0.152939
R13600 gnd.n3518 gnd.n3517 0.152939
R13601 gnd.n3519 gnd.n3518 0.152939
R13602 gnd.n3520 gnd.n3519 0.152939
R13603 gnd.n3521 gnd.n3520 0.152939
R13604 gnd.n3522 gnd.n3521 0.152939
R13605 gnd.n3523 gnd.n3522 0.152939
R13606 gnd.n3524 gnd.n3523 0.152939
R13607 gnd.n3525 gnd.n3524 0.152939
R13608 gnd.n3526 gnd.n3525 0.152939
R13609 gnd.n3527 gnd.n3526 0.152939
R13610 gnd.n3528 gnd.n3527 0.152939
R13611 gnd.n3529 gnd.n3528 0.152939
R13612 gnd.n3530 gnd.n3529 0.152939
R13613 gnd.n3531 gnd.n3530 0.152939
R13614 gnd.n3532 gnd.n3531 0.152939
R13615 gnd.n3533 gnd.n3532 0.152939
R13616 gnd.n3534 gnd.n3533 0.152939
R13617 gnd.n3535 gnd.n3534 0.152939
R13618 gnd.n3536 gnd.n3535 0.152939
R13619 gnd.n3540 gnd.n3536 0.152939
R13620 gnd.n3541 gnd.n3540 0.152939
R13621 gnd.n3541 gnd.n3498 0.152939
R13622 gnd.n3595 gnd.n3498 0.152939
R13623 gnd.n2840 gnd.n2839 0.152939
R13624 gnd.n2839 gnd.n2838 0.152939
R13625 gnd.n2838 gnd.n1786 0.152939
R13626 gnd.n1791 gnd.n1786 0.152939
R13627 gnd.n1792 gnd.n1791 0.152939
R13628 gnd.n1793 gnd.n1792 0.152939
R13629 gnd.n1798 gnd.n1793 0.152939
R13630 gnd.n1799 gnd.n1798 0.152939
R13631 gnd.n1800 gnd.n1799 0.152939
R13632 gnd.n1801 gnd.n1800 0.152939
R13633 gnd.n1806 gnd.n1801 0.152939
R13634 gnd.n1807 gnd.n1806 0.152939
R13635 gnd.n1808 gnd.n1807 0.152939
R13636 gnd.n1809 gnd.n1808 0.152939
R13637 gnd.n1814 gnd.n1809 0.152939
R13638 gnd.n1815 gnd.n1814 0.152939
R13639 gnd.n1816 gnd.n1815 0.152939
R13640 gnd.n1817 gnd.n1816 0.152939
R13641 gnd.n1822 gnd.n1817 0.152939
R13642 gnd.n1823 gnd.n1822 0.152939
R13643 gnd.n1824 gnd.n1823 0.152939
R13644 gnd.n1825 gnd.n1824 0.152939
R13645 gnd.n1830 gnd.n1825 0.152939
R13646 gnd.n1831 gnd.n1830 0.152939
R13647 gnd.n1832 gnd.n1831 0.152939
R13648 gnd.n1833 gnd.n1832 0.152939
R13649 gnd.n1838 gnd.n1833 0.152939
R13650 gnd.n1839 gnd.n1838 0.152939
R13651 gnd.n1840 gnd.n1839 0.152939
R13652 gnd.n1841 gnd.n1840 0.152939
R13653 gnd.n1846 gnd.n1841 0.152939
R13654 gnd.n1847 gnd.n1846 0.152939
R13655 gnd.n1848 gnd.n1847 0.152939
R13656 gnd.n1849 gnd.n1848 0.152939
R13657 gnd.n1854 gnd.n1849 0.152939
R13658 gnd.n1855 gnd.n1854 0.152939
R13659 gnd.n1856 gnd.n1855 0.152939
R13660 gnd.n1857 gnd.n1856 0.152939
R13661 gnd.n1862 gnd.n1857 0.152939
R13662 gnd.n1863 gnd.n1862 0.152939
R13663 gnd.n1864 gnd.n1863 0.152939
R13664 gnd.n1865 gnd.n1864 0.152939
R13665 gnd.n1870 gnd.n1865 0.152939
R13666 gnd.n1871 gnd.n1870 0.152939
R13667 gnd.n1872 gnd.n1871 0.152939
R13668 gnd.n1873 gnd.n1872 0.152939
R13669 gnd.n1878 gnd.n1873 0.152939
R13670 gnd.n1879 gnd.n1878 0.152939
R13671 gnd.n1880 gnd.n1879 0.152939
R13672 gnd.n1881 gnd.n1880 0.152939
R13673 gnd.n1886 gnd.n1881 0.152939
R13674 gnd.n1887 gnd.n1886 0.152939
R13675 gnd.n1888 gnd.n1887 0.152939
R13676 gnd.n1889 gnd.n1888 0.152939
R13677 gnd.n1894 gnd.n1889 0.152939
R13678 gnd.n1895 gnd.n1894 0.152939
R13679 gnd.n1896 gnd.n1895 0.152939
R13680 gnd.n1897 gnd.n1896 0.152939
R13681 gnd.n1902 gnd.n1897 0.152939
R13682 gnd.n1903 gnd.n1902 0.152939
R13683 gnd.n1904 gnd.n1903 0.152939
R13684 gnd.n1905 gnd.n1904 0.152939
R13685 gnd.n1910 gnd.n1905 0.152939
R13686 gnd.n1911 gnd.n1910 0.152939
R13687 gnd.n1912 gnd.n1911 0.152939
R13688 gnd.n1913 gnd.n1912 0.152939
R13689 gnd.n1918 gnd.n1913 0.152939
R13690 gnd.n1919 gnd.n1918 0.152939
R13691 gnd.n1920 gnd.n1919 0.152939
R13692 gnd.n1921 gnd.n1920 0.152939
R13693 gnd.n1926 gnd.n1921 0.152939
R13694 gnd.n1927 gnd.n1926 0.152939
R13695 gnd.n1928 gnd.n1927 0.152939
R13696 gnd.n1929 gnd.n1928 0.152939
R13697 gnd.n1934 gnd.n1929 0.152939
R13698 gnd.n1935 gnd.n1934 0.152939
R13699 gnd.n1936 gnd.n1935 0.152939
R13700 gnd.n1937 gnd.n1936 0.152939
R13701 gnd.n1942 gnd.n1937 0.152939
R13702 gnd.n1943 gnd.n1942 0.152939
R13703 gnd.n1944 gnd.n1943 0.152939
R13704 gnd.n1945 gnd.n1944 0.152939
R13705 gnd.n1950 gnd.n1945 0.152939
R13706 gnd.n1951 gnd.n1950 0.152939
R13707 gnd.n1952 gnd.n1951 0.152939
R13708 gnd.n1953 gnd.n1952 0.152939
R13709 gnd.n1958 gnd.n1953 0.152939
R13710 gnd.n1959 gnd.n1958 0.152939
R13711 gnd.n1960 gnd.n1959 0.152939
R13712 gnd.n1961 gnd.n1960 0.152939
R13713 gnd.n1966 gnd.n1961 0.152939
R13714 gnd.n1967 gnd.n1966 0.152939
R13715 gnd.n1968 gnd.n1967 0.152939
R13716 gnd.n1969 gnd.n1968 0.152939
R13717 gnd.n1974 gnd.n1969 0.152939
R13718 gnd.n1975 gnd.n1974 0.152939
R13719 gnd.n1976 gnd.n1975 0.152939
R13720 gnd.n1977 gnd.n1976 0.152939
R13721 gnd.n1982 gnd.n1977 0.152939
R13722 gnd.n1983 gnd.n1982 0.152939
R13723 gnd.n1984 gnd.n1983 0.152939
R13724 gnd.n1985 gnd.n1984 0.152939
R13725 gnd.n1990 gnd.n1985 0.152939
R13726 gnd.n1991 gnd.n1990 0.152939
R13727 gnd.n1992 gnd.n1991 0.152939
R13728 gnd.n1993 gnd.n1992 0.152939
R13729 gnd.n1998 gnd.n1993 0.152939
R13730 gnd.n1999 gnd.n1998 0.152939
R13731 gnd.n2000 gnd.n1999 0.152939
R13732 gnd.n2001 gnd.n2000 0.152939
R13733 gnd.n2006 gnd.n2001 0.152939
R13734 gnd.n2007 gnd.n2006 0.152939
R13735 gnd.n2008 gnd.n2007 0.152939
R13736 gnd.n2009 gnd.n2008 0.152939
R13737 gnd.n2014 gnd.n2009 0.152939
R13738 gnd.n2015 gnd.n2014 0.152939
R13739 gnd.n2016 gnd.n2015 0.152939
R13740 gnd.n2017 gnd.n2016 0.152939
R13741 gnd.n2022 gnd.n2017 0.152939
R13742 gnd.n2023 gnd.n2022 0.152939
R13743 gnd.n2024 gnd.n2023 0.152939
R13744 gnd.n2025 gnd.n2024 0.152939
R13745 gnd.n2030 gnd.n2025 0.152939
R13746 gnd.n2031 gnd.n2030 0.152939
R13747 gnd.n2032 gnd.n2031 0.152939
R13748 gnd.n2033 gnd.n2032 0.152939
R13749 gnd.n2038 gnd.n2033 0.152939
R13750 gnd.n2039 gnd.n2038 0.152939
R13751 gnd.n2040 gnd.n2039 0.152939
R13752 gnd.n2041 gnd.n2040 0.152939
R13753 gnd.n2046 gnd.n2041 0.152939
R13754 gnd.n2047 gnd.n2046 0.152939
R13755 gnd.n2048 gnd.n2047 0.152939
R13756 gnd.n2049 gnd.n2048 0.152939
R13757 gnd.n2054 gnd.n2049 0.152939
R13758 gnd.n2055 gnd.n2054 0.152939
R13759 gnd.n2056 gnd.n2055 0.152939
R13760 gnd.n2057 gnd.n2056 0.152939
R13761 gnd.n2062 gnd.n2057 0.152939
R13762 gnd.n2063 gnd.n2062 0.152939
R13763 gnd.n2064 gnd.n2063 0.152939
R13764 gnd.n2065 gnd.n2064 0.152939
R13765 gnd.n2070 gnd.n2065 0.152939
R13766 gnd.n2071 gnd.n2070 0.152939
R13767 gnd.n2072 gnd.n2071 0.152939
R13768 gnd.n2073 gnd.n2072 0.152939
R13769 gnd.n2078 gnd.n2073 0.152939
R13770 gnd.n2079 gnd.n2078 0.152939
R13771 gnd.n2080 gnd.n2079 0.152939
R13772 gnd.n2081 gnd.n2080 0.152939
R13773 gnd.n2086 gnd.n2081 0.152939
R13774 gnd.n2087 gnd.n2086 0.152939
R13775 gnd.n2088 gnd.n2087 0.152939
R13776 gnd.n2089 gnd.n2088 0.152939
R13777 gnd.n2094 gnd.n2089 0.152939
R13778 gnd.n2095 gnd.n2094 0.152939
R13779 gnd.n2096 gnd.n2095 0.152939
R13780 gnd.n2097 gnd.n2096 0.152939
R13781 gnd.n2102 gnd.n2097 0.152939
R13782 gnd.n2103 gnd.n2102 0.152939
R13783 gnd.n2104 gnd.n2103 0.152939
R13784 gnd.n2105 gnd.n2104 0.152939
R13785 gnd.n2110 gnd.n2105 0.152939
R13786 gnd.n2111 gnd.n2110 0.152939
R13787 gnd.n2112 gnd.n2111 0.152939
R13788 gnd.n2113 gnd.n2112 0.152939
R13789 gnd.n2118 gnd.n2113 0.152939
R13790 gnd.n2119 gnd.n2118 0.152939
R13791 gnd.n2120 gnd.n2119 0.152939
R13792 gnd.n2121 gnd.n2120 0.152939
R13793 gnd.n2126 gnd.n2121 0.152939
R13794 gnd.n2127 gnd.n2126 0.152939
R13795 gnd.n2128 gnd.n2127 0.152939
R13796 gnd.n2129 gnd.n2128 0.152939
R13797 gnd.n2134 gnd.n2129 0.152939
R13798 gnd.n2135 gnd.n2134 0.152939
R13799 gnd.n2136 gnd.n2135 0.152939
R13800 gnd.n2137 gnd.n2136 0.152939
R13801 gnd.n2142 gnd.n2137 0.152939
R13802 gnd.n2143 gnd.n2142 0.152939
R13803 gnd.n2477 gnd.n2143 0.152939
R13804 gnd.n2476 gnd.n2144 0.152939
R13805 gnd.n2149 gnd.n2144 0.152939
R13806 gnd.n2150 gnd.n2149 0.152939
R13807 gnd.n2151 gnd.n2150 0.152939
R13808 gnd.n2156 gnd.n2151 0.152939
R13809 gnd.n2157 gnd.n2156 0.152939
R13810 gnd.n2158 gnd.n2157 0.152939
R13811 gnd.n2159 gnd.n2158 0.152939
R13812 gnd.n2164 gnd.n2159 0.152939
R13813 gnd.n2165 gnd.n2164 0.152939
R13814 gnd.n2166 gnd.n2165 0.152939
R13815 gnd.n2167 gnd.n2166 0.152939
R13816 gnd.n2172 gnd.n2167 0.152939
R13817 gnd.n2173 gnd.n2172 0.152939
R13818 gnd.n2174 gnd.n2173 0.152939
R13819 gnd.n2175 gnd.n2174 0.152939
R13820 gnd.n2180 gnd.n2175 0.152939
R13821 gnd.n2181 gnd.n2180 0.152939
R13822 gnd.n2182 gnd.n2181 0.152939
R13823 gnd.n2183 gnd.n2182 0.152939
R13824 gnd.n2188 gnd.n2183 0.152939
R13825 gnd.n2189 gnd.n2188 0.152939
R13826 gnd.n2190 gnd.n2189 0.152939
R13827 gnd.n2191 gnd.n2190 0.152939
R13828 gnd.n2196 gnd.n2191 0.152939
R13829 gnd.n2197 gnd.n2196 0.152939
R13830 gnd.n2198 gnd.n2197 0.152939
R13831 gnd.n2199 gnd.n2198 0.152939
R13832 gnd.n2204 gnd.n2199 0.152939
R13833 gnd.n2205 gnd.n2204 0.152939
R13834 gnd.n2206 gnd.n2205 0.152939
R13835 gnd.n2207 gnd.n2206 0.152939
R13836 gnd.n2212 gnd.n2207 0.152939
R13837 gnd.n2213 gnd.n2212 0.152939
R13838 gnd.n2214 gnd.n2213 0.152939
R13839 gnd.n2215 gnd.n2214 0.152939
R13840 gnd.n2220 gnd.n2215 0.152939
R13841 gnd.n2221 gnd.n2220 0.152939
R13842 gnd.n2222 gnd.n2221 0.152939
R13843 gnd.n2223 gnd.n2222 0.152939
R13844 gnd.n2228 gnd.n2223 0.152939
R13845 gnd.n2229 gnd.n2228 0.152939
R13846 gnd.n2230 gnd.n2229 0.152939
R13847 gnd.n2231 gnd.n2230 0.152939
R13848 gnd.n2236 gnd.n2231 0.152939
R13849 gnd.n2237 gnd.n2236 0.152939
R13850 gnd.n2238 gnd.n2237 0.152939
R13851 gnd.n2239 gnd.n2238 0.152939
R13852 gnd.n2244 gnd.n2239 0.152939
R13853 gnd.n2245 gnd.n2244 0.152939
R13854 gnd.n2246 gnd.n2245 0.152939
R13855 gnd.n2247 gnd.n2246 0.152939
R13856 gnd.n2252 gnd.n2247 0.152939
R13857 gnd.n2253 gnd.n2252 0.152939
R13858 gnd.n2254 gnd.n2253 0.152939
R13859 gnd.n2255 gnd.n2254 0.152939
R13860 gnd.n2260 gnd.n2255 0.152939
R13861 gnd.n2261 gnd.n2260 0.152939
R13862 gnd.n2262 gnd.n2261 0.152939
R13863 gnd.n2263 gnd.n2262 0.152939
R13864 gnd.n2268 gnd.n2263 0.152939
R13865 gnd.n2269 gnd.n2268 0.152939
R13866 gnd.n2270 gnd.n2269 0.152939
R13867 gnd.n2271 gnd.n2270 0.152939
R13868 gnd.n2276 gnd.n2271 0.152939
R13869 gnd.n2277 gnd.n2276 0.152939
R13870 gnd.n2278 gnd.n2277 0.152939
R13871 gnd.n2279 gnd.n2278 0.152939
R13872 gnd.n2284 gnd.n2279 0.152939
R13873 gnd.n2285 gnd.n2284 0.152939
R13874 gnd.n2286 gnd.n2285 0.152939
R13875 gnd.n2287 gnd.n2286 0.152939
R13876 gnd.n2292 gnd.n2287 0.152939
R13877 gnd.n2293 gnd.n2292 0.152939
R13878 gnd.n2294 gnd.n2293 0.152939
R13879 gnd.n2295 gnd.n2294 0.152939
R13880 gnd.n2300 gnd.n2295 0.152939
R13881 gnd.n2301 gnd.n2300 0.152939
R13882 gnd.n2302 gnd.n2301 0.152939
R13883 gnd.n2303 gnd.n2302 0.152939
R13884 gnd.n2307 gnd.n2303 0.152939
R13885 gnd.n2308 gnd.n2307 0.152939
R13886 gnd.n2308 gnd.n338 0.152939
R13887 gnd.n7561 gnd.n338 0.152939
R13888 gnd.n7590 gnd.n7589 0.152939
R13889 gnd.n7590 gnd.n286 0.152939
R13890 gnd.n7604 gnd.n286 0.152939
R13891 gnd.n7605 gnd.n7604 0.152939
R13892 gnd.n7606 gnd.n7605 0.152939
R13893 gnd.n7606 gnd.n272 0.152939
R13894 gnd.n7620 gnd.n272 0.152939
R13895 gnd.n7621 gnd.n7620 0.152939
R13896 gnd.n7622 gnd.n7621 0.152939
R13897 gnd.n7622 gnd.n256 0.152939
R13898 gnd.n7636 gnd.n256 0.152939
R13899 gnd.n7637 gnd.n7636 0.152939
R13900 gnd.n7638 gnd.n7637 0.152939
R13901 gnd.n7638 gnd.n242 0.152939
R13902 gnd.n7652 gnd.n242 0.152939
R13903 gnd.n7653 gnd.n7652 0.152939
R13904 gnd.n7654 gnd.n7653 0.152939
R13905 gnd.n7654 gnd.n226 0.152939
R13906 gnd.n7668 gnd.n226 0.152939
R13907 gnd.n7669 gnd.n7668 0.152939
R13908 gnd.n7670 gnd.n7669 0.152939
R13909 gnd.n7670 gnd.n210 0.152939
R13910 gnd.n7752 gnd.n210 0.152939
R13911 gnd.n7753 gnd.n7752 0.152939
R13912 gnd.n7754 gnd.n7753 0.152939
R13913 gnd.n7754 gnd.n133 0.152939
R13914 gnd.n7834 gnd.n133 0.152939
R13915 gnd.n7833 gnd.n134 0.152939
R13916 gnd.n136 gnd.n134 0.152939
R13917 gnd.n140 gnd.n136 0.152939
R13918 gnd.n141 gnd.n140 0.152939
R13919 gnd.n142 gnd.n141 0.152939
R13920 gnd.n143 gnd.n142 0.152939
R13921 gnd.n147 gnd.n143 0.152939
R13922 gnd.n148 gnd.n147 0.152939
R13923 gnd.n149 gnd.n148 0.152939
R13924 gnd.n150 gnd.n149 0.152939
R13925 gnd.n154 gnd.n150 0.152939
R13926 gnd.n155 gnd.n154 0.152939
R13927 gnd.n156 gnd.n155 0.152939
R13928 gnd.n157 gnd.n156 0.152939
R13929 gnd.n161 gnd.n157 0.152939
R13930 gnd.n162 gnd.n161 0.152939
R13931 gnd.n163 gnd.n162 0.152939
R13932 gnd.n164 gnd.n163 0.152939
R13933 gnd.n168 gnd.n164 0.152939
R13934 gnd.n169 gnd.n168 0.152939
R13935 gnd.n170 gnd.n169 0.152939
R13936 gnd.n171 gnd.n170 0.152939
R13937 gnd.n175 gnd.n171 0.152939
R13938 gnd.n176 gnd.n175 0.152939
R13939 gnd.n177 gnd.n176 0.152939
R13940 gnd.n178 gnd.n177 0.152939
R13941 gnd.n182 gnd.n178 0.152939
R13942 gnd.n183 gnd.n182 0.152939
R13943 gnd.n184 gnd.n183 0.152939
R13944 gnd.n185 gnd.n184 0.152939
R13945 gnd.n189 gnd.n185 0.152939
R13946 gnd.n190 gnd.n189 0.152939
R13947 gnd.n191 gnd.n190 0.152939
R13948 gnd.n192 gnd.n191 0.152939
R13949 gnd.n196 gnd.n192 0.152939
R13950 gnd.n197 gnd.n196 0.152939
R13951 gnd.n7764 gnd.n197 0.152939
R13952 gnd.n7764 gnd.n7763 0.152939
R13953 gnd.n599 gnd.n579 0.152939
R13954 gnd.n604 gnd.n599 0.152939
R13955 gnd.n605 gnd.n604 0.152939
R13956 gnd.n606 gnd.n605 0.152939
R13957 gnd.n606 gnd.n597 0.152939
R13958 gnd.n614 gnd.n597 0.152939
R13959 gnd.n615 gnd.n614 0.152939
R13960 gnd.n616 gnd.n615 0.152939
R13961 gnd.n616 gnd.n595 0.152939
R13962 gnd.n7131 gnd.n595 0.152939
R13963 gnd.n7132 gnd.n7131 0.152939
R13964 gnd.n7133 gnd.n7132 0.152939
R13965 gnd.n7134 gnd.n7133 0.152939
R13966 gnd.n7135 gnd.n7134 0.152939
R13967 gnd.n7136 gnd.n7135 0.152939
R13968 gnd.n7137 gnd.n7136 0.152939
R13969 gnd.n7138 gnd.n7137 0.152939
R13970 gnd.n7139 gnd.n7138 0.152939
R13971 gnd.n7139 gnd.n393 0.152939
R13972 gnd.n7404 gnd.n393 0.152939
R13973 gnd.n7405 gnd.n7404 0.152939
R13974 gnd.n7406 gnd.n7405 0.152939
R13975 gnd.n7407 gnd.n7406 0.152939
R13976 gnd.n7408 gnd.n7407 0.152939
R13977 gnd.n7408 gnd.n359 0.152939
R13978 gnd.n7450 gnd.n359 0.152939
R13979 gnd.n7451 gnd.n7450 0.152939
R13980 gnd.n7452 gnd.n7451 0.152939
R13981 gnd.n7453 gnd.n7452 0.152939
R13982 gnd.n7454 gnd.n7453 0.152939
R13983 gnd.n7455 gnd.n7454 0.152939
R13984 gnd.n7456 gnd.n7455 0.152939
R13985 gnd.n7457 gnd.n7456 0.152939
R13986 gnd.n7458 gnd.n7457 0.152939
R13987 gnd.n7459 gnd.n7458 0.152939
R13988 gnd.n7460 gnd.n7459 0.152939
R13989 gnd.n7461 gnd.n7460 0.152939
R13990 gnd.n7462 gnd.n7461 0.152939
R13991 gnd.n7463 gnd.n7462 0.152939
R13992 gnd.n7464 gnd.n7463 0.152939
R13993 gnd.n7465 gnd.n7464 0.152939
R13994 gnd.n7466 gnd.n7465 0.152939
R13995 gnd.n7467 gnd.n7466 0.152939
R13996 gnd.n7468 gnd.n7467 0.152939
R13997 gnd.n7469 gnd.n7468 0.152939
R13998 gnd.n7470 gnd.n7469 0.152939
R13999 gnd.n7471 gnd.n7470 0.152939
R14000 gnd.n7472 gnd.n7471 0.152939
R14001 gnd.n7473 gnd.n7472 0.152939
R14002 gnd.n7474 gnd.n7473 0.152939
R14003 gnd.n7475 gnd.n7474 0.152939
R14004 gnd.n7476 gnd.n7475 0.152939
R14005 gnd.n7477 gnd.n7476 0.152939
R14006 gnd.n7478 gnd.n7477 0.152939
R14007 gnd.n7479 gnd.n7478 0.152939
R14008 gnd.n7480 gnd.n7479 0.152939
R14009 gnd.n7481 gnd.n7480 0.152939
R14010 gnd.n7482 gnd.n7481 0.152939
R14011 gnd.n7483 gnd.n7482 0.152939
R14012 gnd.n7484 gnd.n7483 0.152939
R14013 gnd.n7486 gnd.n7484 0.152939
R14014 gnd.n7486 gnd.n7485 0.152939
R14015 gnd.n7485 gnd.n203 0.152939
R14016 gnd.n7762 gnd.n203 0.152939
R14017 gnd.n536 gnd.n535 0.152939
R14018 gnd.n537 gnd.n536 0.152939
R14019 gnd.n538 gnd.n537 0.152939
R14020 gnd.n539 gnd.n538 0.152939
R14021 gnd.n540 gnd.n539 0.152939
R14022 gnd.n541 gnd.n540 0.152939
R14023 gnd.n542 gnd.n541 0.152939
R14024 gnd.n543 gnd.n542 0.152939
R14025 gnd.n544 gnd.n543 0.152939
R14026 gnd.n545 gnd.n544 0.152939
R14027 gnd.n546 gnd.n545 0.152939
R14028 gnd.n547 gnd.n546 0.152939
R14029 gnd.n548 gnd.n547 0.152939
R14030 gnd.n549 gnd.n548 0.152939
R14031 gnd.n550 gnd.n549 0.152939
R14032 gnd.n557 gnd.n556 0.152939
R14033 gnd.n558 gnd.n557 0.152939
R14034 gnd.n559 gnd.n558 0.152939
R14035 gnd.n560 gnd.n559 0.152939
R14036 gnd.n561 gnd.n560 0.152939
R14037 gnd.n562 gnd.n561 0.152939
R14038 gnd.n563 gnd.n562 0.152939
R14039 gnd.n564 gnd.n563 0.152939
R14040 gnd.n565 gnd.n564 0.152939
R14041 gnd.n566 gnd.n565 0.152939
R14042 gnd.n567 gnd.n566 0.152939
R14043 gnd.n568 gnd.n567 0.152939
R14044 gnd.n569 gnd.n568 0.152939
R14045 gnd.n570 gnd.n569 0.152939
R14046 gnd.n571 gnd.n570 0.152939
R14047 gnd.n572 gnd.n571 0.152939
R14048 gnd.n573 gnd.n572 0.152939
R14049 gnd.n7182 gnd.n573 0.152939
R14050 gnd.n7182 gnd.n7181 0.152939
R14051 gnd.n7181 gnd.n7180 0.152939
R14052 gnd.n7264 gnd.n492 0.152939
R14053 gnd.n7265 gnd.n7264 0.152939
R14054 gnd.n7266 gnd.n7265 0.152939
R14055 gnd.n7266 gnd.n474 0.152939
R14056 gnd.n7280 gnd.n474 0.152939
R14057 gnd.n7281 gnd.n7280 0.152939
R14058 gnd.n7282 gnd.n7281 0.152939
R14059 gnd.n7282 gnd.n457 0.152939
R14060 gnd.n7296 gnd.n457 0.152939
R14061 gnd.n7297 gnd.n7296 0.152939
R14062 gnd.n7298 gnd.n7297 0.152939
R14063 gnd.n7298 gnd.n437 0.152939
R14064 gnd.n7318 gnd.n437 0.152939
R14065 gnd.n7319 gnd.n7318 0.152939
R14066 gnd.n7320 gnd.n7319 0.152939
R14067 gnd.n7321 gnd.n7320 0.152939
R14068 gnd.n7321 gnd.n402 0.152939
R14069 gnd.n7394 gnd.n402 0.152939
R14070 gnd.n7395 gnd.n7394 0.152939
R14071 gnd.n7396 gnd.n7395 0.152939
R14072 gnd.n7397 gnd.n7396 0.152939
R14073 gnd.n7397 gnd.n369 0.152939
R14074 gnd.n7441 gnd.n369 0.152939
R14075 gnd.n7442 gnd.n7441 0.152939
R14076 gnd.n7443 gnd.n7442 0.152939
R14077 gnd.n7443 gnd.n302 0.152939
R14078 gnd.n7589 gnd.n302 0.152939
R14079 gnd.n7360 gnd.n7357 0.152939
R14080 gnd.n7361 gnd.n7360 0.152939
R14081 gnd.n7362 gnd.n7361 0.152939
R14082 gnd.n7363 gnd.n7362 0.152939
R14083 gnd.n340 gnd.n339 0.152939
R14084 gnd.n7560 gnd.n339 0.152939
R14085 gnd.n4968 gnd.n4967 0.152939
R14086 gnd.n4969 gnd.n4968 0.152939
R14087 gnd.n4970 gnd.n4969 0.152939
R14088 gnd.n4971 gnd.n4970 0.152939
R14089 gnd.n4974 gnd.n4971 0.152939
R14090 gnd.n4975 gnd.n4974 0.152939
R14091 gnd.n4976 gnd.n4975 0.152939
R14092 gnd.n4977 gnd.n4976 0.152939
R14093 gnd.n4979 gnd.n4977 0.152939
R14094 gnd.n4979 gnd.n4978 0.152939
R14095 gnd.n4978 gnd.n4951 0.152939
R14096 gnd.n5039 gnd.n4951 0.152939
R14097 gnd.n5040 gnd.n5039 0.152939
R14098 gnd.n5041 gnd.n5040 0.152939
R14099 gnd.n5041 gnd.n4947 0.152939
R14100 gnd.n5047 gnd.n4947 0.152939
R14101 gnd.n5048 gnd.n5047 0.152939
R14102 gnd.n5049 gnd.n5048 0.152939
R14103 gnd.n5050 gnd.n5049 0.152939
R14104 gnd.n5051 gnd.n5050 0.152939
R14105 gnd.n5054 gnd.n5051 0.152939
R14106 gnd.n5055 gnd.n5054 0.152939
R14107 gnd.n5056 gnd.n5055 0.152939
R14108 gnd.n5057 gnd.n5056 0.152939
R14109 gnd.n5060 gnd.n5057 0.152939
R14110 gnd.n5061 gnd.n5060 0.152939
R14111 gnd.n5062 gnd.n5061 0.152939
R14112 gnd.n5063 gnd.n5062 0.152939
R14113 gnd.n5066 gnd.n5063 0.152939
R14114 gnd.n5067 gnd.n5066 0.152939
R14115 gnd.n5068 gnd.n5067 0.152939
R14116 gnd.n5069 gnd.n5068 0.152939
R14117 gnd.n5069 gnd.n1094 0.152939
R14118 gnd.n5803 gnd.n1094 0.152939
R14119 gnd.n5804 gnd.n5803 0.152939
R14120 gnd.n5805 gnd.n5804 0.152939
R14121 gnd.n5805 gnd.n1081 0.152939
R14122 gnd.n5819 gnd.n1081 0.152939
R14123 gnd.n5820 gnd.n5819 0.152939
R14124 gnd.n5821 gnd.n5820 0.152939
R14125 gnd.n5821 gnd.n1067 0.152939
R14126 gnd.n5835 gnd.n1067 0.152939
R14127 gnd.n5836 gnd.n5835 0.152939
R14128 gnd.n5837 gnd.n5836 0.152939
R14129 gnd.n5837 gnd.n1053 0.152939
R14130 gnd.n5851 gnd.n1053 0.152939
R14131 gnd.n5852 gnd.n5851 0.152939
R14132 gnd.n5853 gnd.n5852 0.152939
R14133 gnd.n5853 gnd.n1038 0.152939
R14134 gnd.n5867 gnd.n1038 0.152939
R14135 gnd.n5868 gnd.n5867 0.152939
R14136 gnd.n5869 gnd.n5868 0.152939
R14137 gnd.n5869 gnd.n1024 0.152939
R14138 gnd.n5883 gnd.n1024 0.152939
R14139 gnd.n5884 gnd.n5883 0.152939
R14140 gnd.n5885 gnd.n5884 0.152939
R14141 gnd.n5886 gnd.n5885 0.152939
R14142 gnd.n5886 gnd.n984 0.152939
R14143 gnd.n5981 gnd.n984 0.152939
R14144 gnd.n5982 gnd.n5981 0.152939
R14145 gnd.n5983 gnd.n5982 0.152939
R14146 gnd.n5983 gnd.n968 0.152939
R14147 gnd.n5997 gnd.n968 0.152939
R14148 gnd.n5998 gnd.n5997 0.152939
R14149 gnd.n5999 gnd.n5998 0.152939
R14150 gnd.n5999 gnd.n950 0.152939
R14151 gnd.n6016 gnd.n950 0.152939
R14152 gnd.n6017 gnd.n6016 0.152939
R14153 gnd.n6018 gnd.n6017 0.152939
R14154 gnd.n6018 gnd.n914 0.152939
R14155 gnd.n6072 gnd.n914 0.152939
R14156 gnd.n6073 gnd.n6072 0.152939
R14157 gnd.n6074 gnd.n6073 0.152939
R14158 gnd.n6075 gnd.n6074 0.152939
R14159 gnd.n6075 gnd.n880 0.152939
R14160 gnd.n6836 gnd.n880 0.152939
R14161 gnd.n6837 gnd.n6836 0.152939
R14162 gnd.n6838 gnd.n6837 0.152939
R14163 gnd.n6838 gnd.n865 0.152939
R14164 gnd.n6852 gnd.n865 0.152939
R14165 gnd.n6853 gnd.n6852 0.152939
R14166 gnd.n6854 gnd.n6853 0.152939
R14167 gnd.n6854 gnd.n849 0.152939
R14168 gnd.n6868 gnd.n849 0.152939
R14169 gnd.n6869 gnd.n6868 0.152939
R14170 gnd.n6870 gnd.n6869 0.152939
R14171 gnd.n6870 gnd.n833 0.152939
R14172 gnd.n6884 gnd.n833 0.152939
R14173 gnd.n6885 gnd.n6884 0.152939
R14174 gnd.n6886 gnd.n6885 0.152939
R14175 gnd.n6886 gnd.n817 0.152939
R14176 gnd.n6900 gnd.n817 0.152939
R14177 gnd.n6901 gnd.n6900 0.152939
R14178 gnd.n6902 gnd.n6901 0.152939
R14179 gnd.n6902 gnd.n802 0.152939
R14180 gnd.n6916 gnd.n802 0.152939
R14181 gnd.n6917 gnd.n6916 0.152939
R14182 gnd.n6918 gnd.n6917 0.152939
R14183 gnd.n6918 gnd.n786 0.152939
R14184 gnd.n6932 gnd.n786 0.152939
R14185 gnd.n6933 gnd.n6932 0.152939
R14186 gnd.n6934 gnd.n6933 0.152939
R14187 gnd.n6934 gnd.n770 0.152939
R14188 gnd.n6948 gnd.n770 0.152939
R14189 gnd.n6949 gnd.n6948 0.152939
R14190 gnd.n6950 gnd.n6949 0.152939
R14191 gnd.n6950 gnd.n754 0.152939
R14192 gnd.n6964 gnd.n754 0.152939
R14193 gnd.n6965 gnd.n6964 0.152939
R14194 gnd.n6966 gnd.n6965 0.152939
R14195 gnd.n6966 gnd.n738 0.152939
R14196 gnd.n6980 gnd.n738 0.152939
R14197 gnd.n6981 gnd.n6980 0.152939
R14198 gnd.n6982 gnd.n6981 0.152939
R14199 gnd.n6982 gnd.n723 0.152939
R14200 gnd.n6996 gnd.n723 0.152939
R14201 gnd.n6997 gnd.n6996 0.152939
R14202 gnd.n6998 gnd.n6997 0.152939
R14203 gnd.n6998 gnd.n709 0.152939
R14204 gnd.n7012 gnd.n709 0.152939
R14205 gnd.n7013 gnd.n7012 0.152939
R14206 gnd.n7014 gnd.n7013 0.152939
R14207 gnd.n7014 gnd.n695 0.152939
R14208 gnd.n7028 gnd.n695 0.152939
R14209 gnd.n7029 gnd.n7028 0.152939
R14210 gnd.n7030 gnd.n7029 0.152939
R14211 gnd.n7030 gnd.n681 0.152939
R14212 gnd.n7044 gnd.n681 0.152939
R14213 gnd.n7045 gnd.n7044 0.152939
R14214 gnd.n7046 gnd.n7045 0.152939
R14215 gnd.n7046 gnd.n666 0.152939
R14216 gnd.n7061 gnd.n666 0.152939
R14217 gnd.n7062 gnd.n7061 0.152939
R14218 gnd.n7063 gnd.n7062 0.152939
R14219 gnd.n7064 gnd.n7063 0.152939
R14220 gnd.n7064 gnd.n636 0.152939
R14221 gnd.n7081 gnd.n636 0.152939
R14222 gnd.n7082 gnd.n7081 0.152939
R14223 gnd.n7083 gnd.n7082 0.152939
R14224 gnd.n7083 gnd.n632 0.152939
R14225 gnd.n7089 gnd.n632 0.152939
R14226 gnd.n7090 gnd.n7089 0.152939
R14227 gnd.n7091 gnd.n7090 0.152939
R14228 gnd.n7091 gnd.n628 0.152939
R14229 gnd.n7097 gnd.n628 0.152939
R14230 gnd.n7098 gnd.n7097 0.152939
R14231 gnd.n7099 gnd.n7098 0.152939
R14232 gnd.n7099 gnd.n624 0.152939
R14233 gnd.n7105 gnd.n624 0.152939
R14234 gnd.n7106 gnd.n7105 0.152939
R14235 gnd.n7107 gnd.n7106 0.152939
R14236 gnd.n7108 gnd.n7107 0.152939
R14237 gnd.n7109 gnd.n7108 0.152939
R14238 gnd.n7112 gnd.n7109 0.152939
R14239 gnd.n7113 gnd.n7112 0.152939
R14240 gnd.n7114 gnd.n7113 0.152939
R14241 gnd.n7116 gnd.n7114 0.152939
R14242 gnd.n7116 gnd.n7115 0.152939
R14243 gnd.n7115 gnd.n418 0.152939
R14244 gnd.n7347 gnd.n418 0.152939
R14245 gnd.n7348 gnd.n7347 0.152939
R14246 gnd.n7349 gnd.n7348 0.152939
R14247 gnd.n7350 gnd.n7349 0.152939
R14248 gnd.n7351 gnd.n7350 0.152939
R14249 gnd.n7354 gnd.n7351 0.152939
R14250 gnd.n7355 gnd.n7354 0.152939
R14251 gnd.n7356 gnd.n7355 0.152939
R14252 gnd.n7357 gnd.n7356 0.152939
R14253 gnd.n4515 gnd.n4514 0.152939
R14254 gnd.n4516 gnd.n4515 0.152939
R14255 gnd.n4517 gnd.n4516 0.152939
R14256 gnd.n4518 gnd.n4517 0.152939
R14257 gnd.n4519 gnd.n4518 0.152939
R14258 gnd.n4520 gnd.n4519 0.152939
R14259 gnd.n4521 gnd.n4520 0.152939
R14260 gnd.n4522 gnd.n4521 0.152939
R14261 gnd.n4523 gnd.n4522 0.152939
R14262 gnd.n4524 gnd.n4523 0.152939
R14263 gnd.n4525 gnd.n4524 0.152939
R14264 gnd.n4526 gnd.n4525 0.152939
R14265 gnd.n4527 gnd.n4526 0.152939
R14266 gnd.n4528 gnd.n4527 0.152939
R14267 gnd.n4529 gnd.n4528 0.152939
R14268 gnd.n4530 gnd.n4529 0.152939
R14269 gnd.n4531 gnd.n4530 0.152939
R14270 gnd.n4532 gnd.n4531 0.152939
R14271 gnd.n4533 gnd.n4532 0.152939
R14272 gnd.n4535 gnd.n4533 0.152939
R14273 gnd.n4535 gnd.n4534 0.152939
R14274 gnd.n4534 gnd.n1475 0.152939
R14275 gnd.n4865 gnd.n1475 0.152939
R14276 gnd.n4866 gnd.n4865 0.152939
R14277 gnd.n4867 gnd.n4866 0.152939
R14278 gnd.n4869 gnd.n4867 0.152939
R14279 gnd.n4869 gnd.n4868 0.152939
R14280 gnd.n4868 gnd.n1441 0.152939
R14281 gnd.n1441 gnd.n1439 0.152939
R14282 gnd.n4907 gnd.n1439 0.152939
R14283 gnd.n4908 gnd.n4907 0.152939
R14284 gnd.n4466 gnd.n1562 0.152939
R14285 gnd.n4474 gnd.n4466 0.152939
R14286 gnd.n4475 gnd.n4474 0.152939
R14287 gnd.n4476 gnd.n4475 0.152939
R14288 gnd.n4476 gnd.n4462 0.152939
R14289 gnd.n4484 gnd.n4462 0.152939
R14290 gnd.n4485 gnd.n4484 0.152939
R14291 gnd.n4486 gnd.n4485 0.152939
R14292 gnd.n4486 gnd.n4458 0.152939
R14293 gnd.n4494 gnd.n4458 0.152939
R14294 gnd.n4495 gnd.n4494 0.152939
R14295 gnd.n4496 gnd.n4495 0.152939
R14296 gnd.n4496 gnd.n4454 0.152939
R14297 gnd.n4504 gnd.n4454 0.152939
R14298 gnd.n4505 gnd.n4504 0.152939
R14299 gnd.n4506 gnd.n4505 0.152939
R14300 gnd.n4506 gnd.n4448 0.152939
R14301 gnd.n4513 gnd.n4448 0.152939
R14302 gnd.n4762 gnd.n4761 0.152939
R14303 gnd.n4763 gnd.n4762 0.152939
R14304 gnd.n4763 gnd.n1547 0.152939
R14305 gnd.n4777 gnd.n1547 0.152939
R14306 gnd.n4778 gnd.n4777 0.152939
R14307 gnd.n4779 gnd.n4778 0.152939
R14308 gnd.n4779 gnd.n1530 0.152939
R14309 gnd.n4793 gnd.n1530 0.152939
R14310 gnd.n4794 gnd.n4793 0.152939
R14311 gnd.n4795 gnd.n4794 0.152939
R14312 gnd.n4795 gnd.n1515 0.152939
R14313 gnd.n4809 gnd.n1515 0.152939
R14314 gnd.n4810 gnd.n4809 0.152939
R14315 gnd.n4811 gnd.n4810 0.152939
R14316 gnd.n4811 gnd.n1498 0.152939
R14317 gnd.n4825 gnd.n1498 0.152939
R14318 gnd.n4826 gnd.n4825 0.152939
R14319 gnd.n4827 gnd.n4826 0.152939
R14320 gnd.n4828 gnd.n4827 0.152939
R14321 gnd.n4829 gnd.n4828 0.152939
R14322 gnd.n4831 gnd.n4829 0.152939
R14323 gnd.n4831 gnd.n4830 0.152939
R14324 gnd.n4830 gnd.n1464 0.152939
R14325 gnd.n1465 gnd.n1464 0.152939
R14326 gnd.n1466 gnd.n1465 0.152939
R14327 gnd.n1467 gnd.n1466 0.152939
R14328 gnd.n1469 gnd.n1467 0.152939
R14329 gnd.n1469 gnd.n1468 0.152939
R14330 gnd.n1468 gnd.n1399 0.152939
R14331 gnd.n1400 gnd.n1399 0.152939
R14332 gnd.n1401 gnd.n1400 0.152939
R14333 gnd.n5207 gnd.n1401 0.152939
R14334 gnd.n5210 gnd.n5207 0.152939
R14335 gnd.n5211 gnd.n5210 0.152939
R14336 gnd.n5212 gnd.n5211 0.152939
R14337 gnd.n5212 gnd.n1374 0.152939
R14338 gnd.n5249 gnd.n1374 0.152939
R14339 gnd.n5250 gnd.n5249 0.152939
R14340 gnd.n5251 gnd.n5250 0.152939
R14341 gnd.n5251 gnd.n1357 0.152939
R14342 gnd.n5265 gnd.n1357 0.152939
R14343 gnd.n5266 gnd.n5265 0.152939
R14344 gnd.n5267 gnd.n5266 0.152939
R14345 gnd.n5267 gnd.n1339 0.152939
R14346 gnd.n5281 gnd.n1339 0.152939
R14347 gnd.n5282 gnd.n5281 0.152939
R14348 gnd.n5283 gnd.n5282 0.152939
R14349 gnd.n5283 gnd.n1322 0.152939
R14350 gnd.n5297 gnd.n1322 0.152939
R14351 gnd.n5298 gnd.n5297 0.152939
R14352 gnd.n5299 gnd.n5298 0.152939
R14353 gnd.n5299 gnd.n1304 0.152939
R14354 gnd.n5313 gnd.n1304 0.152939
R14355 gnd.n5314 gnd.n5313 0.152939
R14356 gnd.n5315 gnd.n5314 0.152939
R14357 gnd.n5315 gnd.n1287 0.152939
R14358 gnd.n5329 gnd.n1287 0.152939
R14359 gnd.n5330 gnd.n5329 0.152939
R14360 gnd.n5331 gnd.n5330 0.152939
R14361 gnd.n5331 gnd.n1268 0.152939
R14362 gnd.n5347 gnd.n1268 0.152939
R14363 gnd.n5348 gnd.n5347 0.152939
R14364 gnd.n5349 gnd.n5348 0.152939
R14365 gnd.n5660 gnd.n5349 0.152939
R14366 gnd.n5243 gnd.n1366 0.152939
R14367 gnd.n5257 gnd.n1366 0.152939
R14368 gnd.n5258 gnd.n5257 0.152939
R14369 gnd.n5259 gnd.n5258 0.152939
R14370 gnd.n5259 gnd.n1348 0.152939
R14371 gnd.n5273 gnd.n1348 0.152939
R14372 gnd.n5274 gnd.n5273 0.152939
R14373 gnd.n5275 gnd.n5274 0.152939
R14374 gnd.n5275 gnd.n1331 0.152939
R14375 gnd.n5289 gnd.n1331 0.152939
R14376 gnd.n5290 gnd.n5289 0.152939
R14377 gnd.n5291 gnd.n5290 0.152939
R14378 gnd.n5291 gnd.n1313 0.152939
R14379 gnd.n5305 gnd.n1313 0.152939
R14380 gnd.n5306 gnd.n5305 0.152939
R14381 gnd.n5307 gnd.n5306 0.152939
R14382 gnd.n5307 gnd.n1296 0.152939
R14383 gnd.n5321 gnd.n1296 0.152939
R14384 gnd.n5322 gnd.n5321 0.152939
R14385 gnd.n5323 gnd.n5322 0.152939
R14386 gnd.n5323 gnd.n1278 0.152939
R14387 gnd.n5337 gnd.n1278 0.152939
R14388 gnd.n5338 gnd.n5337 0.152939
R14389 gnd.n5339 gnd.n5338 0.152939
R14390 gnd.n5340 gnd.n5339 0.152939
R14391 gnd.n5340 gnd.n1182 0.152939
R14392 gnd.n5738 gnd.n1182 0.152939
R14393 gnd.n5737 gnd.n1183 0.152939
R14394 gnd.n1199 gnd.n1183 0.152939
R14395 gnd.n1200 gnd.n1199 0.152939
R14396 gnd.n1201 gnd.n1200 0.152939
R14397 gnd.n1202 gnd.n1201 0.152939
R14398 gnd.n1203 gnd.n1202 0.152939
R14399 gnd.n1207 gnd.n1203 0.152939
R14400 gnd.n1208 gnd.n1207 0.152939
R14401 gnd.n1209 gnd.n1208 0.152939
R14402 gnd.n1210 gnd.n1209 0.152939
R14403 gnd.n1214 gnd.n1210 0.152939
R14404 gnd.n1215 gnd.n1214 0.152939
R14405 gnd.n1216 gnd.n1215 0.152939
R14406 gnd.n1217 gnd.n1216 0.152939
R14407 gnd.n1224 gnd.n1217 0.152939
R14408 gnd.n1227 gnd.n1226 0.152939
R14409 gnd.n1228 gnd.n1227 0.152939
R14410 gnd.n1232 gnd.n1228 0.152939
R14411 gnd.n1233 gnd.n1232 0.152939
R14412 gnd.n1234 gnd.n1233 0.152939
R14413 gnd.n1235 gnd.n1234 0.152939
R14414 gnd.n1239 gnd.n1235 0.152939
R14415 gnd.n1240 gnd.n1239 0.152939
R14416 gnd.n1241 gnd.n1240 0.152939
R14417 gnd.n1242 gnd.n1241 0.152939
R14418 gnd.n1246 gnd.n1242 0.152939
R14419 gnd.n1247 gnd.n1246 0.152939
R14420 gnd.n1248 gnd.n1247 0.152939
R14421 gnd.n1249 gnd.n1248 0.152939
R14422 gnd.n1253 gnd.n1249 0.152939
R14423 gnd.n1254 gnd.n1253 0.152939
R14424 gnd.n1255 gnd.n1254 0.152939
R14425 gnd.n1256 gnd.n1255 0.152939
R14426 gnd.n1261 gnd.n1256 0.152939
R14427 gnd.n5669 gnd.n1261 0.152939
R14428 gnd.n4675 gnd.n4629 0.152939
R14429 gnd.n4631 gnd.n4629 0.152939
R14430 gnd.n4632 gnd.n4631 0.152939
R14431 gnd.n4633 gnd.n4632 0.152939
R14432 gnd.n4634 gnd.n4633 0.152939
R14433 gnd.n4635 gnd.n4634 0.152939
R14434 gnd.n4636 gnd.n4635 0.152939
R14435 gnd.n4637 gnd.n4636 0.152939
R14436 gnd.n4638 gnd.n4637 0.152939
R14437 gnd.n4639 gnd.n4638 0.152939
R14438 gnd.n4640 gnd.n4639 0.152939
R14439 gnd.n4641 gnd.n4640 0.152939
R14440 gnd.n4642 gnd.n4641 0.152939
R14441 gnd.n4643 gnd.n4642 0.152939
R14442 gnd.n4644 gnd.n4643 0.152939
R14443 gnd.n4645 gnd.n4644 0.152939
R14444 gnd.n4646 gnd.n4645 0.152939
R14445 gnd.n4647 gnd.n4646 0.152939
R14446 gnd.n4647 gnd.n1481 0.152939
R14447 gnd.n4851 gnd.n1481 0.152939
R14448 gnd.n4852 gnd.n4851 0.152939
R14449 gnd.n4853 gnd.n4852 0.152939
R14450 gnd.n4854 gnd.n4853 0.152939
R14451 gnd.n4855 gnd.n4854 0.152939
R14452 gnd.n4855 gnd.n1446 0.152939
R14453 gnd.n4891 gnd.n1446 0.152939
R14454 gnd.n4892 gnd.n4891 0.152939
R14455 gnd.n4893 gnd.n4892 0.152939
R14456 gnd.n4894 gnd.n4893 0.152939
R14457 gnd.n4895 gnd.n4894 0.152939
R14458 gnd.n4895 gnd.n1428 0.152939
R14459 gnd.n5206 gnd.n1428 0.152939
R14460 gnd.n5206 gnd.n1429 0.152939
R14461 gnd.n1431 gnd.n1429 0.152939
R14462 gnd.n1432 gnd.n1431 0.152939
R14463 gnd.n1433 gnd.n1432 0.152939
R14464 gnd.n4959 gnd.n1433 0.152939
R14465 gnd.n4960 gnd.n4959 0.152939
R14466 gnd.n4960 gnd.n4958 0.152939
R14467 gnd.n5000 gnd.n4958 0.152939
R14468 gnd.n5001 gnd.n5000 0.152939
R14469 gnd.n5002 gnd.n5001 0.152939
R14470 gnd.n5002 gnd.n4956 0.152939
R14471 gnd.n5010 gnd.n4956 0.152939
R14472 gnd.n5011 gnd.n5010 0.152939
R14473 gnd.n5012 gnd.n5011 0.152939
R14474 gnd.n5013 gnd.n5012 0.152939
R14475 gnd.n5014 gnd.n5013 0.152939
R14476 gnd.n5015 gnd.n5014 0.152939
R14477 gnd.n5016 gnd.n5015 0.152939
R14478 gnd.n5017 gnd.n5016 0.152939
R14479 gnd.n5018 gnd.n5017 0.152939
R14480 gnd.n5018 gnd.n4942 0.152939
R14481 gnd.n5100 gnd.n4942 0.152939
R14482 gnd.n5101 gnd.n5100 0.152939
R14483 gnd.n5102 gnd.n5101 0.152939
R14484 gnd.n5102 gnd.n4940 0.152939
R14485 gnd.n5110 gnd.n4940 0.152939
R14486 gnd.n5111 gnd.n5110 0.152939
R14487 gnd.n5112 gnd.n5111 0.152939
R14488 gnd.n5114 gnd.n5112 0.152939
R14489 gnd.n5114 gnd.n5113 0.152939
R14490 gnd.n5113 gnd.n1262 0.152939
R14491 gnd.n5668 gnd.n1262 0.152939
R14492 gnd.n4754 gnd.n4568 0.152939
R14493 gnd.n4571 gnd.n4568 0.152939
R14494 gnd.n4572 gnd.n4571 0.152939
R14495 gnd.n4573 gnd.n4572 0.152939
R14496 gnd.n4576 gnd.n4573 0.152939
R14497 gnd.n4577 gnd.n4576 0.152939
R14498 gnd.n4578 gnd.n4577 0.152939
R14499 gnd.n4579 gnd.n4578 0.152939
R14500 gnd.n4582 gnd.n4579 0.152939
R14501 gnd.n4583 gnd.n4582 0.152939
R14502 gnd.n4584 gnd.n4583 0.152939
R14503 gnd.n4585 gnd.n4584 0.152939
R14504 gnd.n4588 gnd.n4585 0.152939
R14505 gnd.n4589 gnd.n4588 0.152939
R14506 gnd.n4590 gnd.n4589 0.152939
R14507 gnd.n4591 gnd.n4590 0.152939
R14508 gnd.n4597 gnd.n4591 0.152939
R14509 gnd.n4598 gnd.n4597 0.152939
R14510 gnd.n4599 gnd.n4598 0.152939
R14511 gnd.n4600 gnd.n4599 0.152939
R14512 gnd.n4603 gnd.n4600 0.152939
R14513 gnd.n4604 gnd.n4603 0.152939
R14514 gnd.n4605 gnd.n4604 0.152939
R14515 gnd.n4606 gnd.n4605 0.152939
R14516 gnd.n4609 gnd.n4606 0.152939
R14517 gnd.n4610 gnd.n4609 0.152939
R14518 gnd.n4611 gnd.n4610 0.152939
R14519 gnd.n4612 gnd.n4611 0.152939
R14520 gnd.n4615 gnd.n4612 0.152939
R14521 gnd.n4616 gnd.n4615 0.152939
R14522 gnd.n4617 gnd.n4616 0.152939
R14523 gnd.n4618 gnd.n4617 0.152939
R14524 gnd.n4621 gnd.n4618 0.152939
R14525 gnd.n4622 gnd.n4621 0.152939
R14526 gnd.n4623 gnd.n4622 0.152939
R14527 gnd.n4682 gnd.n4623 0.152939
R14528 gnd.n4682 gnd.n4681 0.152939
R14529 gnd.n4681 gnd.n4680 0.152939
R14530 gnd.n4755 gnd.n1555 0.152939
R14531 gnd.n4769 gnd.n1555 0.152939
R14532 gnd.n4770 gnd.n4769 0.152939
R14533 gnd.n4771 gnd.n4770 0.152939
R14534 gnd.n4771 gnd.n1539 0.152939
R14535 gnd.n4785 gnd.n1539 0.152939
R14536 gnd.n4786 gnd.n4785 0.152939
R14537 gnd.n4787 gnd.n4786 0.152939
R14538 gnd.n4787 gnd.n1523 0.152939
R14539 gnd.n4801 gnd.n1523 0.152939
R14540 gnd.n4802 gnd.n4801 0.152939
R14541 gnd.n4803 gnd.n4802 0.152939
R14542 gnd.n4803 gnd.n1507 0.152939
R14543 gnd.n4817 gnd.n1507 0.152939
R14544 gnd.n4818 gnd.n4817 0.152939
R14545 gnd.n4819 gnd.n4818 0.152939
R14546 gnd.n4819 gnd.n1490 0.152939
R14547 gnd.n4841 gnd.n1490 0.152939
R14548 gnd.n4842 gnd.n4841 0.152939
R14549 gnd.n4843 gnd.n4842 0.152939
R14550 gnd.n4844 gnd.n4843 0.152939
R14551 gnd.n4844 gnd.n1454 0.152939
R14552 gnd.n4882 gnd.n1454 0.152939
R14553 gnd.n4883 gnd.n4882 0.152939
R14554 gnd.n4884 gnd.n4883 0.152939
R14555 gnd.n4884 gnd.n1383 0.152939
R14556 gnd.n5243 gnd.n1383 0.152939
R14557 gnd.n3055 gnd.n3051 0.152939
R14558 gnd.n3051 gnd.n1416 0.152939
R14559 gnd.n1418 gnd.n1417 0.152939
R14560 gnd.n4964 gnd.n1418 0.152939
R14561 gnd.n4967 gnd.n4964 0.152939
R14562 gnd.n2848 gnd.n1780 0.152939
R14563 gnd.n2849 gnd.n2848 0.152939
R14564 gnd.n2850 gnd.n2849 0.152939
R14565 gnd.n2850 gnd.n1774 0.152939
R14566 gnd.n2858 gnd.n1774 0.152939
R14567 gnd.n2859 gnd.n2858 0.152939
R14568 gnd.n2860 gnd.n2859 0.152939
R14569 gnd.n2860 gnd.n1768 0.152939
R14570 gnd.n2868 gnd.n1768 0.152939
R14571 gnd.n2869 gnd.n2868 0.152939
R14572 gnd.n2870 gnd.n2869 0.152939
R14573 gnd.n2870 gnd.n1762 0.152939
R14574 gnd.n2878 gnd.n1762 0.152939
R14575 gnd.n2879 gnd.n2878 0.152939
R14576 gnd.n2880 gnd.n2879 0.152939
R14577 gnd.n2880 gnd.n1756 0.152939
R14578 gnd.n2888 gnd.n1756 0.152939
R14579 gnd.n2889 gnd.n2888 0.152939
R14580 gnd.n2890 gnd.n2889 0.152939
R14581 gnd.n2890 gnd.n1750 0.152939
R14582 gnd.n2898 gnd.n1750 0.152939
R14583 gnd.n2899 gnd.n2898 0.152939
R14584 gnd.n2900 gnd.n2899 0.152939
R14585 gnd.n2900 gnd.n1744 0.152939
R14586 gnd.n2908 gnd.n1744 0.152939
R14587 gnd.n2909 gnd.n2908 0.152939
R14588 gnd.n2910 gnd.n2909 0.152939
R14589 gnd.n2910 gnd.n1738 0.152939
R14590 gnd.n2918 gnd.n1738 0.152939
R14591 gnd.n2919 gnd.n2918 0.152939
R14592 gnd.n2920 gnd.n2919 0.152939
R14593 gnd.n2920 gnd.n1732 0.152939
R14594 gnd.n2928 gnd.n1732 0.152939
R14595 gnd.n2929 gnd.n2928 0.152939
R14596 gnd.n2930 gnd.n2929 0.152939
R14597 gnd.n2930 gnd.n1726 0.152939
R14598 gnd.n2938 gnd.n1726 0.152939
R14599 gnd.n2939 gnd.n2938 0.152939
R14600 gnd.n2940 gnd.n2939 0.152939
R14601 gnd.n2940 gnd.n1720 0.152939
R14602 gnd.n2948 gnd.n1720 0.152939
R14603 gnd.n2949 gnd.n2948 0.152939
R14604 gnd.n2950 gnd.n2949 0.152939
R14605 gnd.n2950 gnd.n1714 0.152939
R14606 gnd.n2958 gnd.n1714 0.152939
R14607 gnd.n2959 gnd.n2958 0.152939
R14608 gnd.n2960 gnd.n2959 0.152939
R14609 gnd.n2960 gnd.n1708 0.152939
R14610 gnd.n2968 gnd.n1708 0.152939
R14611 gnd.n2969 gnd.n2968 0.152939
R14612 gnd.n2970 gnd.n2969 0.152939
R14613 gnd.n2970 gnd.n1702 0.152939
R14614 gnd.n2978 gnd.n1702 0.152939
R14615 gnd.n2979 gnd.n2978 0.152939
R14616 gnd.n2980 gnd.n2979 0.152939
R14617 gnd.n2980 gnd.n1696 0.152939
R14618 gnd.n2988 gnd.n1696 0.152939
R14619 gnd.n2989 gnd.n2988 0.152939
R14620 gnd.n2990 gnd.n2989 0.152939
R14621 gnd.n2990 gnd.n1690 0.152939
R14622 gnd.n2998 gnd.n1690 0.152939
R14623 gnd.n2999 gnd.n2998 0.152939
R14624 gnd.n3000 gnd.n2999 0.152939
R14625 gnd.n3000 gnd.n1684 0.152939
R14626 gnd.n3008 gnd.n1684 0.152939
R14627 gnd.n3009 gnd.n3008 0.152939
R14628 gnd.n3010 gnd.n3009 0.152939
R14629 gnd.n3010 gnd.n1678 0.152939
R14630 gnd.n3018 gnd.n1678 0.152939
R14631 gnd.n3019 gnd.n3018 0.152939
R14632 gnd.n3020 gnd.n3019 0.152939
R14633 gnd.n3020 gnd.n1672 0.152939
R14634 gnd.n3028 gnd.n1672 0.152939
R14635 gnd.n3029 gnd.n3028 0.152939
R14636 gnd.n3030 gnd.n3029 0.152939
R14637 gnd.n3030 gnd.n1666 0.152939
R14638 gnd.n3038 gnd.n1666 0.152939
R14639 gnd.n3039 gnd.n3038 0.152939
R14640 gnd.n3040 gnd.n3039 0.152939
R14641 gnd.n3040 gnd.n1660 0.152939
R14642 gnd.n3048 gnd.n1660 0.152939
R14643 gnd.n3049 gnd.n3048 0.152939
R14644 gnd.n3050 gnd.n3049 0.152939
R14645 gnd.n3056 gnd.n3050 0.152939
R14646 gnd.n6678 gnd.n6677 0.152939
R14647 gnd.n6677 gnd.n6676 0.152939
R14648 gnd.n6676 gnd.n6656 0.152939
R14649 gnd.n6672 gnd.n6656 0.152939
R14650 gnd.n6672 gnd.n6671 0.152939
R14651 gnd.n6671 gnd.n6670 0.152939
R14652 gnd.n6670 gnd.n6662 0.152939
R14653 gnd.n6662 gnd.n657 0.152939
R14654 gnd.n7073 gnd.n657 0.152939
R14655 gnd.n5797 gnd.n1088 0.152939
R14656 gnd.n5811 gnd.n1088 0.152939
R14657 gnd.n5812 gnd.n5811 0.152939
R14658 gnd.n5813 gnd.n5812 0.152939
R14659 gnd.n5813 gnd.n1074 0.152939
R14660 gnd.n5827 gnd.n1074 0.152939
R14661 gnd.n5828 gnd.n5827 0.152939
R14662 gnd.n5829 gnd.n5828 0.152939
R14663 gnd.n5829 gnd.n1059 0.152939
R14664 gnd.n5843 gnd.n1059 0.152939
R14665 gnd.n5844 gnd.n5843 0.152939
R14666 gnd.n5845 gnd.n5844 0.152939
R14667 gnd.n5845 gnd.n1045 0.152939
R14668 gnd.n5859 gnd.n1045 0.152939
R14669 gnd.n5860 gnd.n5859 0.152939
R14670 gnd.n5861 gnd.n5860 0.152939
R14671 gnd.n5861 gnd.n1031 0.152939
R14672 gnd.n5875 gnd.n1031 0.152939
R14673 gnd.n5876 gnd.n5875 0.152939
R14674 gnd.n5877 gnd.n5876 0.152939
R14675 gnd.n5877 gnd.n1015 0.152939
R14676 gnd.n5893 gnd.n1015 0.152939
R14677 gnd.n5894 gnd.n5893 0.152939
R14678 gnd.n5896 gnd.n5894 0.152939
R14679 gnd.n5896 gnd.n5895 0.152939
R14680 gnd.n5895 gnd.n976 0.152939
R14681 gnd.n5989 gnd.n976 0.152939
R14682 gnd.n5990 gnd.n5989 0.152939
R14683 gnd.n5991 gnd.n5990 0.152939
R14684 gnd.n5991 gnd.n960 0.152939
R14685 gnd.n6005 gnd.n960 0.152939
R14686 gnd.n6006 gnd.n6005 0.152939
R14687 gnd.n6010 gnd.n6006 0.152939
R14688 gnd.n6010 gnd.n6009 0.152939
R14689 gnd.n6009 gnd.n6008 0.152939
R14690 gnd.n6008 gnd.n924 0.152939
R14691 gnd.n6066 gnd.n924 0.152939
R14692 gnd.n6066 gnd.n6065 0.152939
R14693 gnd.n6065 gnd.n6064 0.152939
R14694 gnd.n6064 gnd.n925 0.152939
R14695 gnd.n6060 gnd.n925 0.152939
R14696 gnd.n6060 gnd.n6059 0.152939
R14697 gnd.n6059 gnd.n873 0.152939
R14698 gnd.n6844 gnd.n873 0.152939
R14699 gnd.n6845 gnd.n6844 0.152939
R14700 gnd.n6846 gnd.n6845 0.152939
R14701 gnd.n6846 gnd.n857 0.152939
R14702 gnd.n6860 gnd.n857 0.152939
R14703 gnd.n6861 gnd.n6860 0.152939
R14704 gnd.n6862 gnd.n6861 0.152939
R14705 gnd.n6862 gnd.n841 0.152939
R14706 gnd.n6876 gnd.n841 0.152939
R14707 gnd.n6877 gnd.n6876 0.152939
R14708 gnd.n6878 gnd.n6877 0.152939
R14709 gnd.n6878 gnd.n825 0.152939
R14710 gnd.n6892 gnd.n825 0.152939
R14711 gnd.n6893 gnd.n6892 0.152939
R14712 gnd.n6894 gnd.n6893 0.152939
R14713 gnd.n6894 gnd.n809 0.152939
R14714 gnd.n6908 gnd.n809 0.152939
R14715 gnd.n6909 gnd.n6908 0.152939
R14716 gnd.n6910 gnd.n6909 0.152939
R14717 gnd.n6910 gnd.n794 0.152939
R14718 gnd.n6924 gnd.n794 0.152939
R14719 gnd.n6925 gnd.n6924 0.152939
R14720 gnd.n6926 gnd.n6925 0.152939
R14721 gnd.n6926 gnd.n778 0.152939
R14722 gnd.n6940 gnd.n778 0.152939
R14723 gnd.n6941 gnd.n6940 0.152939
R14724 gnd.n6942 gnd.n6941 0.152939
R14725 gnd.n6942 gnd.n762 0.152939
R14726 gnd.n6956 gnd.n762 0.152939
R14727 gnd.n6957 gnd.n6956 0.152939
R14728 gnd.n6958 gnd.n6957 0.152939
R14729 gnd.n6958 gnd.n745 0.152939
R14730 gnd.n6972 gnd.n745 0.152939
R14731 gnd.n6973 gnd.n6972 0.152939
R14732 gnd.n6974 gnd.n6973 0.152939
R14733 gnd.n6974 gnd.n731 0.152939
R14734 gnd.n6988 gnd.n731 0.152939
R14735 gnd.n6989 gnd.n6988 0.152939
R14736 gnd.n6990 gnd.n6989 0.152939
R14737 gnd.n6990 gnd.n715 0.152939
R14738 gnd.n7004 gnd.n715 0.152939
R14739 gnd.n7005 gnd.n7004 0.152939
R14740 gnd.n7006 gnd.n7005 0.152939
R14741 gnd.n7006 gnd.n701 0.152939
R14742 gnd.n7020 gnd.n701 0.152939
R14743 gnd.n7021 gnd.n7020 0.152939
R14744 gnd.n7022 gnd.n7021 0.152939
R14745 gnd.n7022 gnd.n688 0.152939
R14746 gnd.n7036 gnd.n688 0.152939
R14747 gnd.n7037 gnd.n7036 0.152939
R14748 gnd.n7038 gnd.n7037 0.152939
R14749 gnd.n7038 gnd.n674 0.152939
R14750 gnd.n7052 gnd.n674 0.152939
R14751 gnd.n7053 gnd.n7052 0.152939
R14752 gnd.n7055 gnd.n7053 0.152939
R14753 gnd.n7055 gnd.n7054 0.152939
R14754 gnd.n7054 gnd.n658 0.152939
R14755 gnd.n7072 gnd.n658 0.152939
R14756 gnd.n5144 gnd.n5121 0.152939
R14757 gnd.n5144 gnd.n5143 0.152939
R14758 gnd.n5143 gnd.n5142 0.152939
R14759 gnd.n5142 gnd.n5127 0.152939
R14760 gnd.n5138 gnd.n5127 0.152939
R14761 gnd.n5138 gnd.n5137 0.152939
R14762 gnd.n5137 gnd.n5134 0.152939
R14763 gnd.n5134 gnd.n1101 0.152939
R14764 gnd.n5796 gnd.n1101 0.152939
R14765 gnd.n4915 gnd.n1437 0.152939
R14766 gnd.n4916 gnd.n4915 0.152939
R14767 gnd.n5194 gnd.n4916 0.152939
R14768 gnd.n5194 gnd.n5193 0.152939
R14769 gnd.n5193 gnd.n5192 0.152939
R14770 gnd.n5192 gnd.n4917 0.152939
R14771 gnd.n5188 gnd.n4917 0.152939
R14772 gnd.n5188 gnd.n5187 0.152939
R14773 gnd.n5187 gnd.n5186 0.152939
R14774 gnd.n5186 gnd.n4921 0.152939
R14775 gnd.n5182 gnd.n4921 0.152939
R14776 gnd.n5182 gnd.n5181 0.152939
R14777 gnd.n5181 gnd.n5180 0.152939
R14778 gnd.n5180 gnd.n4925 0.152939
R14779 gnd.n5176 gnd.n4925 0.152939
R14780 gnd.n5176 gnd.n5175 0.152939
R14781 gnd.n5175 gnd.n5174 0.152939
R14782 gnd.n5174 gnd.n4929 0.152939
R14783 gnd.n5170 gnd.n4929 0.152939
R14784 gnd.n5170 gnd.n5169 0.152939
R14785 gnd.n5169 gnd.n5168 0.152939
R14786 gnd.n5168 gnd.n4933 0.152939
R14787 gnd.n5164 gnd.n4933 0.152939
R14788 gnd.n5164 gnd.n5163 0.152939
R14789 gnd.n5163 gnd.n5162 0.152939
R14790 gnd.n5162 gnd.n4937 0.152939
R14791 gnd.n5158 gnd.n4937 0.152939
R14792 gnd.n5158 gnd.n5157 0.152939
R14793 gnd.n5157 gnd.n5156 0.152939
R14794 gnd.n5156 gnd.n5151 0.152939
R14795 gnd.n5151 gnd.n5150 0.152939
R14796 gnd.n5657 gnd.n5357 0.152939
R14797 gnd.n5653 gnd.n5357 0.152939
R14798 gnd.n5653 gnd.n5652 0.152939
R14799 gnd.n5652 gnd.n5651 0.152939
R14800 gnd.n5651 gnd.n5361 0.152939
R14801 gnd.n5647 gnd.n5361 0.152939
R14802 gnd.n5647 gnd.n5646 0.152939
R14803 gnd.n5646 gnd.n5645 0.152939
R14804 gnd.n5645 gnd.n5365 0.152939
R14805 gnd.n5641 gnd.n5365 0.152939
R14806 gnd.n5641 gnd.n5640 0.152939
R14807 gnd.n5640 gnd.n5639 0.152939
R14808 gnd.n5639 gnd.n5369 0.152939
R14809 gnd.n5635 gnd.n5369 0.152939
R14810 gnd.n5635 gnd.n5634 0.152939
R14811 gnd.n5634 gnd.n5633 0.152939
R14812 gnd.n5633 gnd.n5373 0.152939
R14813 gnd.n5629 gnd.n5373 0.152939
R14814 gnd.n5629 gnd.n5628 0.152939
R14815 gnd.n5628 gnd.n5627 0.152939
R14816 gnd.n5627 gnd.n5377 0.152939
R14817 gnd.n5623 gnd.n5377 0.152939
R14818 gnd.n5623 gnd.n1007 0.152939
R14819 gnd.n5902 gnd.n1007 0.152939
R14820 gnd.n5903 gnd.n5902 0.152939
R14821 gnd.n5904 gnd.n5903 0.152939
R14822 gnd.n5904 gnd.n1004 0.152939
R14823 gnd.n5910 gnd.n1004 0.152939
R14824 gnd.n5911 gnd.n5910 0.152939
R14825 gnd.n5959 gnd.n5911 0.152939
R14826 gnd.n5959 gnd.n5958 0.152939
R14827 gnd.n5958 gnd.n5957 0.152939
R14828 gnd.n5957 gnd.n5912 0.152939
R14829 gnd.n5953 gnd.n5912 0.152939
R14830 gnd.n5953 gnd.n5952 0.152939
R14831 gnd.n5952 gnd.n5951 0.152939
R14832 gnd.n5951 gnd.n5947 0.152939
R14833 gnd.n5947 gnd.n905 0.152939
R14834 gnd.n6082 gnd.n905 0.152939
R14835 gnd.n6083 gnd.n6082 0.152939
R14836 gnd.n6084 gnd.n6083 0.152939
R14837 gnd.n6084 gnd.n902 0.152939
R14838 gnd.n6089 gnd.n902 0.152939
R14839 gnd.n6090 gnd.n6089 0.152939
R14840 gnd.n6817 gnd.n6090 0.152939
R14841 gnd.n6817 gnd.n6816 0.152939
R14842 gnd.n6816 gnd.n6815 0.152939
R14843 gnd.n6815 gnd.n6091 0.152939
R14844 gnd.n6811 gnd.n6091 0.152939
R14845 gnd.n6811 gnd.n6810 0.152939
R14846 gnd.n6810 gnd.n6809 0.152939
R14847 gnd.n6809 gnd.n6095 0.152939
R14848 gnd.n6805 gnd.n6095 0.152939
R14849 gnd.n6805 gnd.n6804 0.152939
R14850 gnd.n6804 gnd.n6803 0.152939
R14851 gnd.n6803 gnd.n6099 0.152939
R14852 gnd.n6799 gnd.n6099 0.152939
R14853 gnd.n6799 gnd.n6798 0.152939
R14854 gnd.n6798 gnd.n6797 0.152939
R14855 gnd.n6797 gnd.n6103 0.152939
R14856 gnd.n6793 gnd.n6103 0.152939
R14857 gnd.n6793 gnd.n6792 0.152939
R14858 gnd.n6792 gnd.n6791 0.152939
R14859 gnd.n6791 gnd.n6107 0.152939
R14860 gnd.n6787 gnd.n6107 0.152939
R14861 gnd.n6787 gnd.n6786 0.152939
R14862 gnd.n6786 gnd.n6785 0.152939
R14863 gnd.n6785 gnd.n6111 0.152939
R14864 gnd.n6781 gnd.n6111 0.152939
R14865 gnd.n6781 gnd.n6780 0.152939
R14866 gnd.n6780 gnd.n6779 0.152939
R14867 gnd.n6779 gnd.n6115 0.152939
R14868 gnd.n6775 gnd.n6115 0.152939
R14869 gnd.n6775 gnd.n6774 0.152939
R14870 gnd.n6774 gnd.n6773 0.152939
R14871 gnd.n6773 gnd.n6119 0.152939
R14872 gnd.n6769 gnd.n6119 0.152939
R14873 gnd.n6769 gnd.n6768 0.152939
R14874 gnd.n6768 gnd.n6767 0.152939
R14875 gnd.n6767 gnd.n6123 0.152939
R14876 gnd.n6763 gnd.n6123 0.152939
R14877 gnd.n6763 gnd.n6762 0.152939
R14878 gnd.n6762 gnd.n6761 0.152939
R14879 gnd.n6761 gnd.n6576 0.152939
R14880 gnd.n6757 gnd.n6576 0.152939
R14881 gnd.n6757 gnd.n6756 0.152939
R14882 gnd.n6756 gnd.n6755 0.152939
R14883 gnd.n6755 gnd.n6581 0.152939
R14884 gnd.n6751 gnd.n6581 0.152939
R14885 gnd.n6751 gnd.n6750 0.152939
R14886 gnd.n6750 gnd.n6749 0.152939
R14887 gnd.n6749 gnd.n6585 0.152939
R14888 gnd.n6745 gnd.n6585 0.152939
R14889 gnd.n6745 gnd.n6744 0.152939
R14890 gnd.n6744 gnd.n6743 0.152939
R14891 gnd.n6743 gnd.n6589 0.152939
R14892 gnd.n6739 gnd.n6589 0.152939
R14893 gnd.n6739 gnd.n6738 0.152939
R14894 gnd.n6738 gnd.n6737 0.152939
R14895 gnd.n6737 gnd.n6593 0.152939
R14896 gnd.n6595 gnd.n6593 0.152939
R14897 gnd.n7258 gnd.n7257 0.152939
R14898 gnd.n7258 gnd.n483 0.152939
R14899 gnd.n7272 gnd.n483 0.152939
R14900 gnd.n7273 gnd.n7272 0.152939
R14901 gnd.n7274 gnd.n7273 0.152939
R14902 gnd.n7274 gnd.n465 0.152939
R14903 gnd.n7288 gnd.n465 0.152939
R14904 gnd.n7289 gnd.n7288 0.152939
R14905 gnd.n7290 gnd.n7289 0.152939
R14906 gnd.n7290 gnd.n448 0.152939
R14907 gnd.n7304 gnd.n448 0.152939
R14908 gnd.n7305 gnd.n7304 0.152939
R14909 gnd.n7312 gnd.n7305 0.152939
R14910 gnd.n7312 gnd.n7311 0.152939
R14911 gnd.n7311 gnd.n7310 0.152939
R14912 gnd.n7310 gnd.n7306 0.152939
R14913 gnd.n7306 gnd.n413 0.152939
R14914 gnd.n7388 gnd.n413 0.152939
R14915 gnd.n7388 gnd.n7387 0.152939
R14916 gnd.n7387 gnd.n7386 0.152939
R14917 gnd.n7386 gnd.n414 0.152939
R14918 gnd.n414 gnd.n381 0.152939
R14919 gnd.n7435 gnd.n381 0.152939
R14920 gnd.n7435 gnd.n7434 0.152939
R14921 gnd.n7434 gnd.n7433 0.152939
R14922 gnd.n7433 gnd.n382 0.152939
R14923 gnd.n7429 gnd.n382 0.152939
R14924 gnd.n7429 gnd.n319 0.152939
R14925 gnd.n7581 gnd.n319 0.152939
R14926 gnd.n7581 gnd.n7580 0.152939
R14927 gnd.n7580 gnd.n7579 0.152939
R14928 gnd.n7579 gnd.n320 0.152939
R14929 gnd.n7575 gnd.n320 0.152939
R14930 gnd.n7575 gnd.n7574 0.152939
R14931 gnd.n7574 gnd.n7573 0.152939
R14932 gnd.n7573 gnd.n325 0.152939
R14933 gnd.n325 gnd.n295 0.152939
R14934 gnd.n7596 gnd.n295 0.152939
R14935 gnd.n7597 gnd.n7596 0.152939
R14936 gnd.n7598 gnd.n7597 0.152939
R14937 gnd.n7598 gnd.n279 0.152939
R14938 gnd.n7612 gnd.n279 0.152939
R14939 gnd.n7613 gnd.n7612 0.152939
R14940 gnd.n7614 gnd.n7613 0.152939
R14941 gnd.n7614 gnd.n265 0.152939
R14942 gnd.n7628 gnd.n265 0.152939
R14943 gnd.n7629 gnd.n7628 0.152939
R14944 gnd.n7630 gnd.n7629 0.152939
R14945 gnd.n7630 gnd.n249 0.152939
R14946 gnd.n7644 gnd.n249 0.152939
R14947 gnd.n7645 gnd.n7644 0.152939
R14948 gnd.n7646 gnd.n7645 0.152939
R14949 gnd.n7646 gnd.n235 0.152939
R14950 gnd.n7660 gnd.n235 0.152939
R14951 gnd.n7661 gnd.n7660 0.152939
R14952 gnd.n7662 gnd.n7661 0.152939
R14953 gnd.n7662 gnd.n220 0.152939
R14954 gnd.n7676 gnd.n220 0.152939
R14955 gnd.n7677 gnd.n7676 0.152939
R14956 gnd.n7746 gnd.n7677 0.152939
R14957 gnd.n7746 gnd.n7745 0.152939
R14958 gnd.n7745 gnd.n7744 0.152939
R14959 gnd.n7744 gnd.n7678 0.152939
R14960 gnd.n7740 gnd.n7678 0.152939
R14961 gnd.n7739 gnd.n7680 0.152939
R14962 gnd.n7735 gnd.n7680 0.152939
R14963 gnd.n7735 gnd.n7734 0.152939
R14964 gnd.n7734 gnd.n7733 0.152939
R14965 gnd.n7733 gnd.n7686 0.152939
R14966 gnd.n7729 gnd.n7686 0.152939
R14967 gnd.n7729 gnd.n7728 0.152939
R14968 gnd.n7728 gnd.n7727 0.152939
R14969 gnd.n7727 gnd.n7694 0.152939
R14970 gnd.n7723 gnd.n7694 0.152939
R14971 gnd.n7723 gnd.n7722 0.152939
R14972 gnd.n7722 gnd.n7721 0.152939
R14973 gnd.n7721 gnd.n7702 0.152939
R14974 gnd.n7717 gnd.n7702 0.152939
R14975 gnd.n7717 gnd.n7716 0.152939
R14976 gnd.n7716 gnd.n7715 0.152939
R14977 gnd.n7715 gnd.n121 0.152939
R14978 gnd.n7841 gnd.n121 0.152939
R14979 gnd.n7173 gnd.n7172 0.152939
R14980 gnd.n7172 gnd.n7171 0.152939
R14981 gnd.n7171 gnd.n584 0.152939
R14982 gnd.n7167 gnd.n584 0.152939
R14983 gnd.n7167 gnd.n7166 0.152939
R14984 gnd.n7166 gnd.n7165 0.152939
R14985 gnd.n7165 gnd.n588 0.152939
R14986 gnd.n7161 gnd.n588 0.152939
R14987 gnd.n7161 gnd.n7160 0.152939
R14988 gnd.n7160 gnd.n7159 0.152939
R14989 gnd.n7159 gnd.n592 0.152939
R14990 gnd.n7155 gnd.n592 0.152939
R14991 gnd.n7155 gnd.n7154 0.152939
R14992 gnd.n7154 gnd.n427 0.152939
R14993 gnd.n7328 gnd.n427 0.152939
R14994 gnd.n7329 gnd.n7328 0.152939
R14995 gnd.n7338 gnd.n7329 0.152939
R14996 gnd.n7338 gnd.n7337 0.152939
R14997 gnd.n7337 gnd.n7336 0.152939
R14998 gnd.n7336 gnd.n7331 0.152939
R14999 gnd.n7331 gnd.n7330 0.152939
R15000 gnd.n7330 gnd.n387 0.152939
R15001 gnd.n7419 gnd.n387 0.152939
R15002 gnd.n7420 gnd.n7419 0.152939
R15003 gnd.n7422 gnd.n7420 0.152939
R15004 gnd.n7422 gnd.n7421 0.152939
R15005 gnd.n7421 gnd.n353 0.152939
R15006 gnd.n7542 gnd.n353 0.152939
R15007 gnd.n7543 gnd.n7542 0.152939
R15008 gnd.n7544 gnd.n7543 0.152939
R15009 gnd.n7544 gnd.n79 0.152939
R15010 gnd.n7890 gnd.n79 0.152939
R15011 gnd.n7890 gnd.n7889 0.152939
R15012 gnd.n7889 gnd.n81 0.152939
R15013 gnd.n7885 gnd.n81 0.152939
R15014 gnd.n7885 gnd.n7884 0.152939
R15015 gnd.n7884 gnd.n7883 0.152939
R15016 gnd.n7883 gnd.n86 0.152939
R15017 gnd.n7879 gnd.n86 0.152939
R15018 gnd.n7879 gnd.n7878 0.152939
R15019 gnd.n7878 gnd.n7877 0.152939
R15020 gnd.n7877 gnd.n91 0.152939
R15021 gnd.n7873 gnd.n91 0.152939
R15022 gnd.n7873 gnd.n7872 0.152939
R15023 gnd.n7872 gnd.n7871 0.152939
R15024 gnd.n7871 gnd.n96 0.152939
R15025 gnd.n7867 gnd.n96 0.152939
R15026 gnd.n7867 gnd.n7866 0.152939
R15027 gnd.n7866 gnd.n7865 0.152939
R15028 gnd.n7865 gnd.n101 0.152939
R15029 gnd.n7861 gnd.n101 0.152939
R15030 gnd.n7861 gnd.n7860 0.152939
R15031 gnd.n7860 gnd.n7859 0.152939
R15032 gnd.n7859 gnd.n106 0.152939
R15033 gnd.n7855 gnd.n106 0.152939
R15034 gnd.n7855 gnd.n7854 0.152939
R15035 gnd.n7854 gnd.n7853 0.152939
R15036 gnd.n7853 gnd.n111 0.152939
R15037 gnd.n7849 gnd.n111 0.152939
R15038 gnd.n7849 gnd.n7848 0.152939
R15039 gnd.n7848 gnd.n7847 0.152939
R15040 gnd.n7847 gnd.n116 0.152939
R15041 gnd.n7843 gnd.n116 0.152939
R15042 gnd.n7843 gnd.n7842 0.152939
R15043 gnd.n6678 gnd.n583 0.151415
R15044 gnd.n5149 gnd.n5121 0.151415
R15045 gnd.n4909 gnd.n4908 0.145814
R15046 gnd.n4909 gnd.n1437 0.145814
R15047 gnd.n7363 gnd.n303 0.0950122
R15048 gnd.n1417 gnd.n1384 0.0950122
R15049 gnd.n3841 gnd.n3840 0.0767195
R15050 gnd.n3840 gnd.n3839 0.0767195
R15051 gnd.n5659 gnd.n5658 0.063
R15052 gnd.n7256 gnd.n501 0.063
R15053 gnd.n340 gnd.n303 0.0584268
R15054 gnd.n1416 gnd.n1384 0.0584268
R15055 gnd.n4407 gnd.n1605 0.0477147
R15056 gnd.n3604 gnd.n3492 0.0442063
R15057 gnd.n3605 gnd.n3604 0.0442063
R15058 gnd.n3606 gnd.n3605 0.0442063
R15059 gnd.n3606 gnd.n3481 0.0442063
R15060 gnd.n3620 gnd.n3481 0.0442063
R15061 gnd.n3621 gnd.n3620 0.0442063
R15062 gnd.n3622 gnd.n3621 0.0442063
R15063 gnd.n3622 gnd.n3468 0.0442063
R15064 gnd.n3666 gnd.n3468 0.0442063
R15065 gnd.n3667 gnd.n3666 0.0442063
R15066 gnd.n3669 gnd.n3402 0.0344674
R15067 gnd.n6682 gnd.n6650 0.0343753
R15068 gnd.n5148 gnd.n1170 0.0343753
R15069 gnd.n3689 gnd.n3688 0.0269946
R15070 gnd.n3691 gnd.n3690 0.0269946
R15071 gnd.n3397 gnd.n3395 0.0269946
R15072 gnd.n3701 gnd.n3699 0.0269946
R15073 gnd.n3700 gnd.n3376 0.0269946
R15074 gnd.n3720 gnd.n3719 0.0269946
R15075 gnd.n3722 gnd.n3721 0.0269946
R15076 gnd.n3371 gnd.n3370 0.0269946
R15077 gnd.n3732 gnd.n3366 0.0269946
R15078 gnd.n3731 gnd.n3368 0.0269946
R15079 gnd.n3367 gnd.n3349 0.0269946
R15080 gnd.n3752 gnd.n3350 0.0269946
R15081 gnd.n3751 gnd.n3351 0.0269946
R15082 gnd.n3785 gnd.n3326 0.0269946
R15083 gnd.n3787 gnd.n3786 0.0269946
R15084 gnd.n3788 gnd.n3273 0.0269946
R15085 gnd.n3321 gnd.n3274 0.0269946
R15086 gnd.n3323 gnd.n3275 0.0269946
R15087 gnd.n3798 gnd.n3797 0.0269946
R15088 gnd.n3800 gnd.n3799 0.0269946
R15089 gnd.n3801 gnd.n3295 0.0269946
R15090 gnd.n3803 gnd.n3296 0.0269946
R15091 gnd.n3806 gnd.n3297 0.0269946
R15092 gnd.n3809 gnd.n3808 0.0269946
R15093 gnd.n3811 gnd.n3810 0.0269946
R15094 gnd.n3876 gnd.n3184 0.0269946
R15095 gnd.n3878 gnd.n3877 0.0269946
R15096 gnd.n3887 gnd.n3177 0.0269946
R15097 gnd.n3889 gnd.n3888 0.0269946
R15098 gnd.n3890 gnd.n3175 0.0269946
R15099 gnd.n3897 gnd.n3893 0.0269946
R15100 gnd.n3896 gnd.n3895 0.0269946
R15101 gnd.n3894 gnd.n3154 0.0269946
R15102 gnd.n3919 gnd.n3155 0.0269946
R15103 gnd.n3918 gnd.n3156 0.0269946
R15104 gnd.n3961 gnd.n3129 0.0269946
R15105 gnd.n3963 gnd.n3962 0.0269946
R15106 gnd.n3972 gnd.n3122 0.0269946
R15107 gnd.n3974 gnd.n3973 0.0269946
R15108 gnd.n3975 gnd.n3120 0.0269946
R15109 gnd.n3982 gnd.n3978 0.0269946
R15110 gnd.n3981 gnd.n3980 0.0269946
R15111 gnd.n3979 gnd.n3099 0.0269946
R15112 gnd.n4004 gnd.n3100 0.0269946
R15113 gnd.n4003 gnd.n3101 0.0269946
R15114 gnd.n4050 gnd.n3075 0.0269946
R15115 gnd.n4052 gnd.n4051 0.0269946
R15116 gnd.n4061 gnd.n3068 0.0269946
R15117 gnd.n4320 gnd.n3066 0.0269946
R15118 gnd.n4325 gnd.n4323 0.0269946
R15119 gnd.n4324 gnd.n1641 0.0269946
R15120 gnd.n4349 gnd.n4348 0.0269946
R15121 gnd.n6597 gnd.n501 0.0245515
R15122 gnd.n5658 gnd.n5356 0.0245515
R15123 gnd.n3669 gnd.n3668 0.0202011
R15124 gnd.n6730 gnd.n6597 0.0174377
R15125 gnd.n6730 gnd.n6729 0.0174377
R15126 gnd.n6729 gnd.n6598 0.0174377
R15127 gnd.n6726 gnd.n6598 0.0174377
R15128 gnd.n6726 gnd.n6725 0.0174377
R15129 gnd.n6725 gnd.n6603 0.0174377
R15130 gnd.n6722 gnd.n6603 0.0174377
R15131 gnd.n6722 gnd.n6721 0.0174377
R15132 gnd.n6721 gnd.n6609 0.0174377
R15133 gnd.n6718 gnd.n6609 0.0174377
R15134 gnd.n6718 gnd.n6717 0.0174377
R15135 gnd.n6717 gnd.n6613 0.0174377
R15136 gnd.n6714 gnd.n6613 0.0174377
R15137 gnd.n6714 gnd.n6713 0.0174377
R15138 gnd.n6713 gnd.n6617 0.0174377
R15139 gnd.n6710 gnd.n6617 0.0174377
R15140 gnd.n6710 gnd.n6709 0.0174377
R15141 gnd.n6709 gnd.n6623 0.0174377
R15142 gnd.n6706 gnd.n6623 0.0174377
R15143 gnd.n6706 gnd.n6705 0.0174377
R15144 gnd.n6705 gnd.n6629 0.0174377
R15145 gnd.n6702 gnd.n6629 0.0174377
R15146 gnd.n6702 gnd.n6701 0.0174377
R15147 gnd.n6701 gnd.n6633 0.0174377
R15148 gnd.n6698 gnd.n6633 0.0174377
R15149 gnd.n6698 gnd.n6697 0.0174377
R15150 gnd.n6697 gnd.n6637 0.0174377
R15151 gnd.n6694 gnd.n6637 0.0174377
R15152 gnd.n6694 gnd.n6693 0.0174377
R15153 gnd.n6693 gnd.n6643 0.0174377
R15154 gnd.n6690 gnd.n6643 0.0174377
R15155 gnd.n6690 gnd.n6689 0.0174377
R15156 gnd.n6689 gnd.n6649 0.0174377
R15157 gnd.n6683 gnd.n6649 0.0174377
R15158 gnd.n6683 gnd.n6682 0.0174377
R15159 gnd.n5356 gnd.n1119 0.0174377
R15160 gnd.n1121 gnd.n1119 0.0174377
R15161 gnd.n5786 gnd.n1121 0.0174377
R15162 gnd.n5786 gnd.n5785 0.0174377
R15163 gnd.n5785 gnd.n1122 0.0174377
R15164 gnd.n5782 gnd.n1122 0.0174377
R15165 gnd.n5782 gnd.n5781 0.0174377
R15166 gnd.n5781 gnd.n1127 0.0174377
R15167 gnd.n5778 gnd.n1127 0.0174377
R15168 gnd.n5778 gnd.n5777 0.0174377
R15169 gnd.n5777 gnd.n1132 0.0174377
R15170 gnd.n5774 gnd.n1132 0.0174377
R15171 gnd.n5774 gnd.n5773 0.0174377
R15172 gnd.n5773 gnd.n1136 0.0174377
R15173 gnd.n5770 gnd.n1136 0.0174377
R15174 gnd.n5770 gnd.n5769 0.0174377
R15175 gnd.n5769 gnd.n1140 0.0174377
R15176 gnd.n5766 gnd.n1140 0.0174377
R15177 gnd.n5766 gnd.n5765 0.0174377
R15178 gnd.n5765 gnd.n1144 0.0174377
R15179 gnd.n5762 gnd.n1144 0.0174377
R15180 gnd.n5762 gnd.n5761 0.0174377
R15181 gnd.n5761 gnd.n1150 0.0174377
R15182 gnd.n5758 gnd.n1150 0.0174377
R15183 gnd.n5758 gnd.n5757 0.0174377
R15184 gnd.n5757 gnd.n1154 0.0174377
R15185 gnd.n5754 gnd.n1154 0.0174377
R15186 gnd.n5754 gnd.n5753 0.0174377
R15187 gnd.n5753 gnd.n1158 0.0174377
R15188 gnd.n5750 gnd.n1158 0.0174377
R15189 gnd.n5750 gnd.n5749 0.0174377
R15190 gnd.n5749 gnd.n1164 0.0174377
R15191 gnd.n5746 gnd.n1164 0.0174377
R15192 gnd.n5746 gnd.n5745 0.0174377
R15193 gnd.n5745 gnd.n1170 0.0174377
R15194 gnd.n3668 gnd.n3667 0.0148637
R15195 gnd.n4318 gnd.n4062 0.0144266
R15196 gnd.n4319 gnd.n4318 0.0130679
R15197 gnd.n3688 gnd.n3402 0.00797283
R15198 gnd.n3690 gnd.n3689 0.00797283
R15199 gnd.n3691 gnd.n3397 0.00797283
R15200 gnd.n3699 gnd.n3395 0.00797283
R15201 gnd.n3701 gnd.n3700 0.00797283
R15202 gnd.n3719 gnd.n3376 0.00797283
R15203 gnd.n3721 gnd.n3720 0.00797283
R15204 gnd.n3722 gnd.n3371 0.00797283
R15205 gnd.n3370 gnd.n3366 0.00797283
R15206 gnd.n3732 gnd.n3731 0.00797283
R15207 gnd.n3368 gnd.n3367 0.00797283
R15208 gnd.n3350 gnd.n3349 0.00797283
R15209 gnd.n3752 gnd.n3751 0.00797283
R15210 gnd.n3351 gnd.n3326 0.00797283
R15211 gnd.n3786 gnd.n3785 0.00797283
R15212 gnd.n3788 gnd.n3787 0.00797283
R15213 gnd.n3321 gnd.n3273 0.00797283
R15214 gnd.n3323 gnd.n3274 0.00797283
R15215 gnd.n3797 gnd.n3275 0.00797283
R15216 gnd.n3799 gnd.n3798 0.00797283
R15217 gnd.n3801 gnd.n3800 0.00797283
R15218 gnd.n3803 gnd.n3295 0.00797283
R15219 gnd.n3806 gnd.n3296 0.00797283
R15220 gnd.n3808 gnd.n3297 0.00797283
R15221 gnd.n3811 gnd.n3809 0.00797283
R15222 gnd.n3810 gnd.n3184 0.00797283
R15223 gnd.n3878 gnd.n3876 0.00797283
R15224 gnd.n3877 gnd.n3177 0.00797283
R15225 gnd.n3888 gnd.n3887 0.00797283
R15226 gnd.n3890 gnd.n3889 0.00797283
R15227 gnd.n3893 gnd.n3175 0.00797283
R15228 gnd.n3897 gnd.n3896 0.00797283
R15229 gnd.n3895 gnd.n3894 0.00797283
R15230 gnd.n3155 gnd.n3154 0.00797283
R15231 gnd.n3919 gnd.n3918 0.00797283
R15232 gnd.n3156 gnd.n3129 0.00797283
R15233 gnd.n3963 gnd.n3961 0.00797283
R15234 gnd.n3962 gnd.n3122 0.00797283
R15235 gnd.n3973 gnd.n3972 0.00797283
R15236 gnd.n3975 gnd.n3974 0.00797283
R15237 gnd.n3978 gnd.n3120 0.00797283
R15238 gnd.n3982 gnd.n3981 0.00797283
R15239 gnd.n3980 gnd.n3979 0.00797283
R15240 gnd.n3100 gnd.n3099 0.00797283
R15241 gnd.n4004 gnd.n4003 0.00797283
R15242 gnd.n3101 gnd.n3075 0.00797283
R15243 gnd.n4052 gnd.n4050 0.00797283
R15244 gnd.n4051 gnd.n3068 0.00797283
R15245 gnd.n4062 gnd.n4061 0.00797283
R15246 gnd.n4320 gnd.n4319 0.00797283
R15247 gnd.n4323 gnd.n3066 0.00797283
R15248 gnd.n4325 gnd.n4324 0.00797283
R15249 gnd.n4348 gnd.n1641 0.00797283
R15250 gnd.n4349 gnd.n1605 0.00797283
R15251 gnd.n7456 gnd.n320 0.00433921
R15252 gnd.n5207 gnd.n5206 0.00433921
R15253 gnd.n6650 gnd.n583 0.000838753
R15254 gnd.n5149 gnd.n5148 0.000838753
R15255 vdd.n315 vdd.n279 756.745
R15256 vdd.n260 vdd.n224 756.745
R15257 vdd.n217 vdd.n181 756.745
R15258 vdd.n162 vdd.n126 756.745
R15259 vdd.n120 vdd.n84 756.745
R15260 vdd.n65 vdd.n29 756.745
R15261 vdd.n1764 vdd.n1728 756.745
R15262 vdd.n1819 vdd.n1783 756.745
R15263 vdd.n1666 vdd.n1630 756.745
R15264 vdd.n1721 vdd.n1685 756.745
R15265 vdd.n1569 vdd.n1533 756.745
R15266 vdd.n1624 vdd.n1588 756.745
R15267 vdd.n1107 vdd.t152 640.208
R15268 vdd.n968 vdd.t190 640.208
R15269 vdd.n1101 vdd.t217 640.208
R15270 vdd.n959 vdd.t214 640.208
R15271 vdd.n856 vdd.t163 640.208
R15272 vdd.n2678 vdd.t208 640.208
R15273 vdd.n804 vdd.t184 640.208
R15274 vdd.n2747 vdd.t194 640.208
R15275 vdd.n768 vdd.t148 640.208
R15276 vdd.n1029 vdd.t204 640.208
R15277 vdd.n1228 vdd.t177 592.009
R15278 vdd.n1384 vdd.t201 592.009
R15279 vdd.n1420 vdd.t211 592.009
R15280 vdd.n2117 vdd.t170 592.009
R15281 vdd.n1967 vdd.t187 592.009
R15282 vdd.n1927 vdd.t198 592.009
R15283 vdd.n405 vdd.t174 592.009
R15284 vdd.n419 vdd.t159 592.009
R15285 vdd.n431 vdd.t181 592.009
R15286 vdd.n723 vdd.t144 592.009
R15287 vdd.n686 vdd.t156 592.009
R15288 vdd.n3195 vdd.t167 592.009
R15289 vdd.n316 vdd.n315 585
R15290 vdd.n314 vdd.n281 585
R15291 vdd.n313 vdd.n312 585
R15292 vdd.n284 vdd.n282 585
R15293 vdd.n307 vdd.n306 585
R15294 vdd.n305 vdd.n304 585
R15295 vdd.n288 vdd.n287 585
R15296 vdd.n299 vdd.n298 585
R15297 vdd.n297 vdd.n296 585
R15298 vdd.n292 vdd.n291 585
R15299 vdd.n261 vdd.n260 585
R15300 vdd.n259 vdd.n226 585
R15301 vdd.n258 vdd.n257 585
R15302 vdd.n229 vdd.n227 585
R15303 vdd.n252 vdd.n251 585
R15304 vdd.n250 vdd.n249 585
R15305 vdd.n233 vdd.n232 585
R15306 vdd.n244 vdd.n243 585
R15307 vdd.n242 vdd.n241 585
R15308 vdd.n237 vdd.n236 585
R15309 vdd.n218 vdd.n217 585
R15310 vdd.n216 vdd.n183 585
R15311 vdd.n215 vdd.n214 585
R15312 vdd.n186 vdd.n184 585
R15313 vdd.n209 vdd.n208 585
R15314 vdd.n207 vdd.n206 585
R15315 vdd.n190 vdd.n189 585
R15316 vdd.n201 vdd.n200 585
R15317 vdd.n199 vdd.n198 585
R15318 vdd.n194 vdd.n193 585
R15319 vdd.n163 vdd.n162 585
R15320 vdd.n161 vdd.n128 585
R15321 vdd.n160 vdd.n159 585
R15322 vdd.n131 vdd.n129 585
R15323 vdd.n154 vdd.n153 585
R15324 vdd.n152 vdd.n151 585
R15325 vdd.n135 vdd.n134 585
R15326 vdd.n146 vdd.n145 585
R15327 vdd.n144 vdd.n143 585
R15328 vdd.n139 vdd.n138 585
R15329 vdd.n121 vdd.n120 585
R15330 vdd.n119 vdd.n86 585
R15331 vdd.n118 vdd.n117 585
R15332 vdd.n89 vdd.n87 585
R15333 vdd.n112 vdd.n111 585
R15334 vdd.n110 vdd.n109 585
R15335 vdd.n93 vdd.n92 585
R15336 vdd.n104 vdd.n103 585
R15337 vdd.n102 vdd.n101 585
R15338 vdd.n97 vdd.n96 585
R15339 vdd.n66 vdd.n65 585
R15340 vdd.n64 vdd.n31 585
R15341 vdd.n63 vdd.n62 585
R15342 vdd.n34 vdd.n32 585
R15343 vdd.n57 vdd.n56 585
R15344 vdd.n55 vdd.n54 585
R15345 vdd.n38 vdd.n37 585
R15346 vdd.n49 vdd.n48 585
R15347 vdd.n47 vdd.n46 585
R15348 vdd.n42 vdd.n41 585
R15349 vdd.n1765 vdd.n1764 585
R15350 vdd.n1763 vdd.n1730 585
R15351 vdd.n1762 vdd.n1761 585
R15352 vdd.n1733 vdd.n1731 585
R15353 vdd.n1756 vdd.n1755 585
R15354 vdd.n1754 vdd.n1753 585
R15355 vdd.n1737 vdd.n1736 585
R15356 vdd.n1748 vdd.n1747 585
R15357 vdd.n1746 vdd.n1745 585
R15358 vdd.n1741 vdd.n1740 585
R15359 vdd.n1820 vdd.n1819 585
R15360 vdd.n1818 vdd.n1785 585
R15361 vdd.n1817 vdd.n1816 585
R15362 vdd.n1788 vdd.n1786 585
R15363 vdd.n1811 vdd.n1810 585
R15364 vdd.n1809 vdd.n1808 585
R15365 vdd.n1792 vdd.n1791 585
R15366 vdd.n1803 vdd.n1802 585
R15367 vdd.n1801 vdd.n1800 585
R15368 vdd.n1796 vdd.n1795 585
R15369 vdd.n1667 vdd.n1666 585
R15370 vdd.n1665 vdd.n1632 585
R15371 vdd.n1664 vdd.n1663 585
R15372 vdd.n1635 vdd.n1633 585
R15373 vdd.n1658 vdd.n1657 585
R15374 vdd.n1656 vdd.n1655 585
R15375 vdd.n1639 vdd.n1638 585
R15376 vdd.n1650 vdd.n1649 585
R15377 vdd.n1648 vdd.n1647 585
R15378 vdd.n1643 vdd.n1642 585
R15379 vdd.n1722 vdd.n1721 585
R15380 vdd.n1720 vdd.n1687 585
R15381 vdd.n1719 vdd.n1718 585
R15382 vdd.n1690 vdd.n1688 585
R15383 vdd.n1713 vdd.n1712 585
R15384 vdd.n1711 vdd.n1710 585
R15385 vdd.n1694 vdd.n1693 585
R15386 vdd.n1705 vdd.n1704 585
R15387 vdd.n1703 vdd.n1702 585
R15388 vdd.n1698 vdd.n1697 585
R15389 vdd.n1570 vdd.n1569 585
R15390 vdd.n1568 vdd.n1535 585
R15391 vdd.n1567 vdd.n1566 585
R15392 vdd.n1538 vdd.n1536 585
R15393 vdd.n1561 vdd.n1560 585
R15394 vdd.n1559 vdd.n1558 585
R15395 vdd.n1542 vdd.n1541 585
R15396 vdd.n1553 vdd.n1552 585
R15397 vdd.n1551 vdd.n1550 585
R15398 vdd.n1546 vdd.n1545 585
R15399 vdd.n1625 vdd.n1624 585
R15400 vdd.n1623 vdd.n1590 585
R15401 vdd.n1622 vdd.n1621 585
R15402 vdd.n1593 vdd.n1591 585
R15403 vdd.n1616 vdd.n1615 585
R15404 vdd.n1614 vdd.n1613 585
R15405 vdd.n1597 vdd.n1596 585
R15406 vdd.n1608 vdd.n1607 585
R15407 vdd.n1606 vdd.n1605 585
R15408 vdd.n1601 vdd.n1600 585
R15409 vdd.n445 vdd.n370 462.44
R15410 vdd.n3433 vdd.n372 462.44
R15411 vdd.n3328 vdd.n657 462.44
R15412 vdd.n3326 vdd.n660 462.44
R15413 vdd.n2112 vdd.n1127 462.44
R15414 vdd.n2115 vdd.n2114 462.44
R15415 vdd.n1455 vdd.n1225 462.44
R15416 vdd.n1452 vdd.n1223 462.44
R15417 vdd.n293 vdd.t30 329.043
R15418 vdd.n238 vdd.t80 329.043
R15419 vdd.n195 vdd.t137 329.043
R15420 vdd.n140 vdd.t64 329.043
R15421 vdd.n98 vdd.t59 329.043
R15422 vdd.n43 vdd.t118 329.043
R15423 vdd.n1742 vdd.t138 329.043
R15424 vdd.n1797 vdd.t78 329.043
R15425 vdd.n1644 vdd.t130 329.043
R15426 vdd.n1699 vdd.t60 329.043
R15427 vdd.n1547 vdd.t96 329.043
R15428 vdd.n1602 vdd.t14 329.043
R15429 vdd.n1228 vdd.t180 319.788
R15430 vdd.n1384 vdd.t203 319.788
R15431 vdd.n1420 vdd.t213 319.788
R15432 vdd.n2117 vdd.t172 319.788
R15433 vdd.n1967 vdd.t188 319.788
R15434 vdd.n1927 vdd.t199 319.788
R15435 vdd.n405 vdd.t175 319.788
R15436 vdd.n419 vdd.t161 319.788
R15437 vdd.n431 vdd.t182 319.788
R15438 vdd.n723 vdd.t147 319.788
R15439 vdd.n686 vdd.t158 319.788
R15440 vdd.n3195 vdd.t169 319.788
R15441 vdd.n1229 vdd.t179 303.69
R15442 vdd.n1385 vdd.t202 303.69
R15443 vdd.n1421 vdd.t212 303.69
R15444 vdd.n2118 vdd.t173 303.69
R15445 vdd.n1968 vdd.t189 303.69
R15446 vdd.n1928 vdd.t200 303.69
R15447 vdd.n406 vdd.t176 303.69
R15448 vdd.n420 vdd.t162 303.69
R15449 vdd.n432 vdd.t183 303.69
R15450 vdd.n724 vdd.t146 303.69
R15451 vdd.n687 vdd.t157 303.69
R15452 vdd.n3196 vdd.t168 303.69
R15453 vdd.n2933 vdd.n918 285.366
R15454 vdd.n3157 vdd.n778 285.366
R15455 vdd.n3094 vdd.n775 285.366
R15456 vdd.n2812 vdd.n915 285.366
R15457 vdd.n2642 vdd.n956 285.366
R15458 vdd.n2573 vdd.n2572 285.366
R15459 vdd.n2313 vdd.n1082 285.366
R15460 vdd.n2383 vdd.n1084 285.366
R15461 vdd.n3073 vdd.n776 285.366
R15462 vdd.n3160 vdd.n3159 285.366
R15463 vdd.n2926 vdd.n916 285.366
R15464 vdd.n2935 vdd.n914 285.366
R15465 vdd.n2570 vdd.n966 285.366
R15466 vdd.n964 vdd.n938 285.366
R15467 vdd.n2199 vdd.n1083 285.366
R15468 vdd.n2385 vdd.n1080 285.366
R15469 vdd.n1125 vdd.n1081 216.982
R15470 vdd.n756 vdd.n658 216.982
R15471 vdd.n3075 vdd.n776 185
R15472 vdd.n3158 vdd.n776 185
R15473 vdd.n3077 vdd.n3076 185
R15474 vdd.n3076 vdd.n774 185
R15475 vdd.n3078 vdd.n810 185
R15476 vdd.n3088 vdd.n810 185
R15477 vdd.n3079 vdd.n819 185
R15478 vdd.n819 vdd.n817 185
R15479 vdd.n3081 vdd.n3080 185
R15480 vdd.n3082 vdd.n3081 185
R15481 vdd.n3034 vdd.n818 185
R15482 vdd.n818 vdd.n814 185
R15483 vdd.n3033 vdd.n3032 185
R15484 vdd.n3032 vdd.n3031 185
R15485 vdd.n821 vdd.n820 185
R15486 vdd.n822 vdd.n821 185
R15487 vdd.n3024 vdd.n3023 185
R15488 vdd.n3025 vdd.n3024 185
R15489 vdd.n3022 vdd.n830 185
R15490 vdd.n835 vdd.n830 185
R15491 vdd.n3021 vdd.n3020 185
R15492 vdd.n3020 vdd.n3019 185
R15493 vdd.n832 vdd.n831 185
R15494 vdd.n841 vdd.n832 185
R15495 vdd.n3012 vdd.n3011 185
R15496 vdd.n3013 vdd.n3012 185
R15497 vdd.n3010 vdd.n842 185
R15498 vdd.n848 vdd.n842 185
R15499 vdd.n3009 vdd.n3008 185
R15500 vdd.n3008 vdd.n3007 185
R15501 vdd.n844 vdd.n843 185
R15502 vdd.n845 vdd.n844 185
R15503 vdd.n3000 vdd.n2999 185
R15504 vdd.n3001 vdd.n3000 185
R15505 vdd.n2998 vdd.n855 185
R15506 vdd.n855 vdd.n852 185
R15507 vdd.n2996 vdd.n2995 185
R15508 vdd.n2995 vdd.n2994 185
R15509 vdd.n858 vdd.n857 185
R15510 vdd.n859 vdd.n858 185
R15511 vdd.n2987 vdd.n2986 185
R15512 vdd.n2988 vdd.n2987 185
R15513 vdd.n2985 vdd.n867 185
R15514 vdd.n872 vdd.n867 185
R15515 vdd.n2984 vdd.n2983 185
R15516 vdd.n2983 vdd.n2982 185
R15517 vdd.n869 vdd.n868 185
R15518 vdd.n2894 vdd.n869 185
R15519 vdd.n2975 vdd.n2974 185
R15520 vdd.n2976 vdd.n2975 185
R15521 vdd.n2973 vdd.n879 185
R15522 vdd.n879 vdd.n876 185
R15523 vdd.n2972 vdd.n2971 185
R15524 vdd.n2971 vdd.n2970 185
R15525 vdd.n881 vdd.n880 185
R15526 vdd.n882 vdd.n881 185
R15527 vdd.n2963 vdd.n2962 185
R15528 vdd.n2964 vdd.n2963 185
R15529 vdd.n2961 vdd.n890 185
R15530 vdd.n2906 vdd.n890 185
R15531 vdd.n2960 vdd.n2959 185
R15532 vdd.n2959 vdd.n2958 185
R15533 vdd.n892 vdd.n891 185
R15534 vdd.n901 vdd.n892 185
R15535 vdd.n2951 vdd.n2950 185
R15536 vdd.n2952 vdd.n2951 185
R15537 vdd.n2949 vdd.n902 185
R15538 vdd.n902 vdd.n898 185
R15539 vdd.n2948 vdd.n2947 185
R15540 vdd.n2947 vdd.n2946 185
R15541 vdd.n904 vdd.n903 185
R15542 vdd.n2918 vdd.n904 185
R15543 vdd.n2939 vdd.n2938 185
R15544 vdd.n2940 vdd.n2939 185
R15545 vdd.n2937 vdd.n912 185
R15546 vdd.n917 vdd.n912 185
R15547 vdd.n2936 vdd.n2935 185
R15548 vdd.n2935 vdd.n2934 185
R15549 vdd.n914 vdd.n913 185
R15550 vdd.n2682 vdd.n2681 185
R15551 vdd.n2684 vdd.n2683 185
R15552 vdd.n2686 vdd.n2685 185
R15553 vdd.n2688 vdd.n2687 185
R15554 vdd.n2690 vdd.n2689 185
R15555 vdd.n2692 vdd.n2691 185
R15556 vdd.n2694 vdd.n2693 185
R15557 vdd.n2696 vdd.n2695 185
R15558 vdd.n2698 vdd.n2697 185
R15559 vdd.n2700 vdd.n2699 185
R15560 vdd.n2702 vdd.n2701 185
R15561 vdd.n2704 vdd.n2703 185
R15562 vdd.n2706 vdd.n2705 185
R15563 vdd.n2708 vdd.n2707 185
R15564 vdd.n2710 vdd.n2709 185
R15565 vdd.n2712 vdd.n2711 185
R15566 vdd.n2714 vdd.n2713 185
R15567 vdd.n2716 vdd.n2715 185
R15568 vdd.n2718 vdd.n2717 185
R15569 vdd.n2720 vdd.n2719 185
R15570 vdd.n2722 vdd.n2721 185
R15571 vdd.n2724 vdd.n2723 185
R15572 vdd.n2726 vdd.n2725 185
R15573 vdd.n2728 vdd.n2727 185
R15574 vdd.n2730 vdd.n2729 185
R15575 vdd.n2732 vdd.n2731 185
R15576 vdd.n2734 vdd.n2733 185
R15577 vdd.n2736 vdd.n2735 185
R15578 vdd.n2738 vdd.n2737 185
R15579 vdd.n2740 vdd.n2739 185
R15580 vdd.n2742 vdd.n2741 185
R15581 vdd.n2744 vdd.n2743 185
R15582 vdd.n2745 vdd.n2677 185
R15583 vdd.n2926 vdd.n2925 185
R15584 vdd.n2927 vdd.n2926 185
R15585 vdd.n3161 vdd.n3160 185
R15586 vdd.n3162 vdd.n767 185
R15587 vdd.n3164 vdd.n3163 185
R15588 vdd.n3166 vdd.n765 185
R15589 vdd.n3168 vdd.n3167 185
R15590 vdd.n3169 vdd.n764 185
R15591 vdd.n3171 vdd.n3170 185
R15592 vdd.n3173 vdd.n762 185
R15593 vdd.n3175 vdd.n3174 185
R15594 vdd.n3176 vdd.n761 185
R15595 vdd.n3178 vdd.n3177 185
R15596 vdd.n3180 vdd.n759 185
R15597 vdd.n3182 vdd.n3181 185
R15598 vdd.n3183 vdd.n758 185
R15599 vdd.n3185 vdd.n3184 185
R15600 vdd.n3187 vdd.n757 185
R15601 vdd.n3188 vdd.n754 185
R15602 vdd.n3191 vdd.n3190 185
R15603 vdd.n755 vdd.n753 185
R15604 vdd.n3047 vdd.n3046 185
R15605 vdd.n3049 vdd.n3048 185
R15606 vdd.n3051 vdd.n3043 185
R15607 vdd.n3053 vdd.n3052 185
R15608 vdd.n3054 vdd.n3042 185
R15609 vdd.n3056 vdd.n3055 185
R15610 vdd.n3058 vdd.n3040 185
R15611 vdd.n3060 vdd.n3059 185
R15612 vdd.n3061 vdd.n3039 185
R15613 vdd.n3063 vdd.n3062 185
R15614 vdd.n3065 vdd.n3037 185
R15615 vdd.n3067 vdd.n3066 185
R15616 vdd.n3068 vdd.n3036 185
R15617 vdd.n3070 vdd.n3069 185
R15618 vdd.n3072 vdd.n3035 185
R15619 vdd.n3074 vdd.n3073 185
R15620 vdd.n3073 vdd.n756 185
R15621 vdd.n3159 vdd.n771 185
R15622 vdd.n3159 vdd.n3158 185
R15623 vdd.n2825 vdd.n773 185
R15624 vdd.n774 vdd.n773 185
R15625 vdd.n2826 vdd.n809 185
R15626 vdd.n3088 vdd.n809 185
R15627 vdd.n2828 vdd.n2827 185
R15628 vdd.n2827 vdd.n817 185
R15629 vdd.n2829 vdd.n816 185
R15630 vdd.n3082 vdd.n816 185
R15631 vdd.n2831 vdd.n2830 185
R15632 vdd.n2830 vdd.n814 185
R15633 vdd.n2832 vdd.n824 185
R15634 vdd.n3031 vdd.n824 185
R15635 vdd.n2834 vdd.n2833 185
R15636 vdd.n2833 vdd.n822 185
R15637 vdd.n2835 vdd.n829 185
R15638 vdd.n3025 vdd.n829 185
R15639 vdd.n2837 vdd.n2836 185
R15640 vdd.n2836 vdd.n835 185
R15641 vdd.n2838 vdd.n834 185
R15642 vdd.n3019 vdd.n834 185
R15643 vdd.n2840 vdd.n2839 185
R15644 vdd.n2839 vdd.n841 185
R15645 vdd.n2841 vdd.n840 185
R15646 vdd.n3013 vdd.n840 185
R15647 vdd.n2843 vdd.n2842 185
R15648 vdd.n2842 vdd.n848 185
R15649 vdd.n2844 vdd.n847 185
R15650 vdd.n3007 vdd.n847 185
R15651 vdd.n2846 vdd.n2845 185
R15652 vdd.n2845 vdd.n845 185
R15653 vdd.n2847 vdd.n854 185
R15654 vdd.n3001 vdd.n854 185
R15655 vdd.n2849 vdd.n2848 185
R15656 vdd.n2848 vdd.n852 185
R15657 vdd.n2850 vdd.n861 185
R15658 vdd.n2994 vdd.n861 185
R15659 vdd.n2852 vdd.n2851 185
R15660 vdd.n2851 vdd.n859 185
R15661 vdd.n2853 vdd.n866 185
R15662 vdd.n2988 vdd.n866 185
R15663 vdd.n2855 vdd.n2854 185
R15664 vdd.n2854 vdd.n872 185
R15665 vdd.n2856 vdd.n871 185
R15666 vdd.n2982 vdd.n871 185
R15667 vdd.n2896 vdd.n2895 185
R15668 vdd.n2895 vdd.n2894 185
R15669 vdd.n2897 vdd.n878 185
R15670 vdd.n2976 vdd.n878 185
R15671 vdd.n2899 vdd.n2898 185
R15672 vdd.n2898 vdd.n876 185
R15673 vdd.n2900 vdd.n884 185
R15674 vdd.n2970 vdd.n884 185
R15675 vdd.n2902 vdd.n2901 185
R15676 vdd.n2901 vdd.n882 185
R15677 vdd.n2903 vdd.n889 185
R15678 vdd.n2964 vdd.n889 185
R15679 vdd.n2905 vdd.n2904 185
R15680 vdd.n2906 vdd.n2905 185
R15681 vdd.n2824 vdd.n894 185
R15682 vdd.n2958 vdd.n894 185
R15683 vdd.n2823 vdd.n2822 185
R15684 vdd.n2822 vdd.n901 185
R15685 vdd.n2821 vdd.n900 185
R15686 vdd.n2952 vdd.n900 185
R15687 vdd.n2820 vdd.n2819 185
R15688 vdd.n2819 vdd.n898 185
R15689 vdd.n2746 vdd.n906 185
R15690 vdd.n2946 vdd.n906 185
R15691 vdd.n2920 vdd.n2919 185
R15692 vdd.n2919 vdd.n2918 185
R15693 vdd.n2921 vdd.n911 185
R15694 vdd.n2940 vdd.n911 185
R15695 vdd.n2923 vdd.n2922 185
R15696 vdd.n2922 vdd.n917 185
R15697 vdd.n2924 vdd.n916 185
R15698 vdd.n2934 vdd.n916 185
R15699 vdd.n2112 vdd.n2111 185
R15700 vdd.n2113 vdd.n2112 185
R15701 vdd.n1128 vdd.n1126 185
R15702 vdd.n1126 vdd.n1124 185
R15703 vdd.n1894 vdd.n1893 185
R15704 vdd.n1893 vdd.n1892 185
R15705 vdd.n1131 vdd.n1130 185
R15706 vdd.n1132 vdd.n1131 185
R15707 vdd.n1881 vdd.n1880 185
R15708 vdd.n1882 vdd.n1881 185
R15709 vdd.n1140 vdd.n1139 185
R15710 vdd.n1873 vdd.n1139 185
R15711 vdd.n1876 vdd.n1875 185
R15712 vdd.n1875 vdd.n1874 185
R15713 vdd.n1143 vdd.n1142 185
R15714 vdd.n1149 vdd.n1143 185
R15715 vdd.n1864 vdd.n1863 185
R15716 vdd.n1865 vdd.n1864 185
R15717 vdd.n1151 vdd.n1150 185
R15718 vdd.n1856 vdd.n1150 185
R15719 vdd.n1859 vdd.n1858 185
R15720 vdd.n1858 vdd.n1857 185
R15721 vdd.n1154 vdd.n1153 185
R15722 vdd.n1155 vdd.n1154 185
R15723 vdd.n1847 vdd.n1846 185
R15724 vdd.n1848 vdd.n1847 185
R15725 vdd.n1163 vdd.n1162 185
R15726 vdd.n1162 vdd.n1161 185
R15727 vdd.n1842 vdd.n1841 185
R15728 vdd.n1841 vdd.n1840 185
R15729 vdd.n1166 vdd.n1165 185
R15730 vdd.n1172 vdd.n1166 185
R15731 vdd.n1831 vdd.n1830 185
R15732 vdd.n1832 vdd.n1831 185
R15733 vdd.n1174 vdd.n1173 185
R15734 vdd.n1528 vdd.n1173 185
R15735 vdd.n1531 vdd.n1530 185
R15736 vdd.n1530 vdd.n1529 185
R15737 vdd.n1177 vdd.n1176 185
R15738 vdd.n1184 vdd.n1177 185
R15739 vdd.n1519 vdd.n1518 185
R15740 vdd.n1520 vdd.n1519 185
R15741 vdd.n1186 vdd.n1185 185
R15742 vdd.n1185 vdd.n1183 185
R15743 vdd.n1514 vdd.n1513 185
R15744 vdd.n1513 vdd.n1512 185
R15745 vdd.n1189 vdd.n1188 185
R15746 vdd.n1190 vdd.n1189 185
R15747 vdd.n1503 vdd.n1502 185
R15748 vdd.n1504 vdd.n1503 185
R15749 vdd.n1197 vdd.n1196 185
R15750 vdd.n1495 vdd.n1196 185
R15751 vdd.n1498 vdd.n1497 185
R15752 vdd.n1497 vdd.n1496 185
R15753 vdd.n1200 vdd.n1199 185
R15754 vdd.n1206 vdd.n1200 185
R15755 vdd.n1486 vdd.n1485 185
R15756 vdd.n1487 vdd.n1486 185
R15757 vdd.n1208 vdd.n1207 185
R15758 vdd.n1478 vdd.n1207 185
R15759 vdd.n1481 vdd.n1480 185
R15760 vdd.n1480 vdd.n1479 185
R15761 vdd.n1211 vdd.n1210 185
R15762 vdd.n1212 vdd.n1211 185
R15763 vdd.n1469 vdd.n1468 185
R15764 vdd.n1470 vdd.n1469 185
R15765 vdd.n1220 vdd.n1219 185
R15766 vdd.n1219 vdd.n1218 185
R15767 vdd.n1464 vdd.n1463 185
R15768 vdd.n1463 vdd.n1462 185
R15769 vdd.n1223 vdd.n1222 185
R15770 vdd.n1224 vdd.n1223 185
R15771 vdd.n1452 vdd.n1451 185
R15772 vdd.n1450 vdd.n1263 185
R15773 vdd.n1265 vdd.n1262 185
R15774 vdd.n1454 vdd.n1262 185
R15775 vdd.n1446 vdd.n1267 185
R15776 vdd.n1445 vdd.n1268 185
R15777 vdd.n1444 vdd.n1269 185
R15778 vdd.n1272 vdd.n1270 185
R15779 vdd.n1440 vdd.n1273 185
R15780 vdd.n1439 vdd.n1274 185
R15781 vdd.n1438 vdd.n1275 185
R15782 vdd.n1278 vdd.n1276 185
R15783 vdd.n1434 vdd.n1279 185
R15784 vdd.n1433 vdd.n1280 185
R15785 vdd.n1432 vdd.n1281 185
R15786 vdd.n1284 vdd.n1282 185
R15787 vdd.n1428 vdd.n1285 185
R15788 vdd.n1427 vdd.n1286 185
R15789 vdd.n1426 vdd.n1287 185
R15790 vdd.n1418 vdd.n1288 185
R15791 vdd.n1422 vdd.n1419 185
R15792 vdd.n1417 vdd.n1290 185
R15793 vdd.n1416 vdd.n1291 185
R15794 vdd.n1294 vdd.n1292 185
R15795 vdd.n1412 vdd.n1295 185
R15796 vdd.n1411 vdd.n1296 185
R15797 vdd.n1410 vdd.n1297 185
R15798 vdd.n1300 vdd.n1298 185
R15799 vdd.n1406 vdd.n1301 185
R15800 vdd.n1405 vdd.n1302 185
R15801 vdd.n1404 vdd.n1303 185
R15802 vdd.n1306 vdd.n1304 185
R15803 vdd.n1400 vdd.n1307 185
R15804 vdd.n1399 vdd.n1308 185
R15805 vdd.n1398 vdd.n1309 185
R15806 vdd.n1312 vdd.n1310 185
R15807 vdd.n1394 vdd.n1313 185
R15808 vdd.n1393 vdd.n1314 185
R15809 vdd.n1392 vdd.n1315 185
R15810 vdd.n1318 vdd.n1316 185
R15811 vdd.n1388 vdd.n1319 185
R15812 vdd.n1387 vdd.n1320 185
R15813 vdd.n1386 vdd.n1383 185
R15814 vdd.n1323 vdd.n1321 185
R15815 vdd.n1379 vdd.n1324 185
R15816 vdd.n1378 vdd.n1325 185
R15817 vdd.n1377 vdd.n1326 185
R15818 vdd.n1329 vdd.n1327 185
R15819 vdd.n1373 vdd.n1330 185
R15820 vdd.n1372 vdd.n1331 185
R15821 vdd.n1371 vdd.n1332 185
R15822 vdd.n1335 vdd.n1333 185
R15823 vdd.n1367 vdd.n1336 185
R15824 vdd.n1366 vdd.n1337 185
R15825 vdd.n1365 vdd.n1338 185
R15826 vdd.n1341 vdd.n1339 185
R15827 vdd.n1361 vdd.n1342 185
R15828 vdd.n1360 vdd.n1343 185
R15829 vdd.n1359 vdd.n1344 185
R15830 vdd.n1347 vdd.n1345 185
R15831 vdd.n1355 vdd.n1348 185
R15832 vdd.n1354 vdd.n1349 185
R15833 vdd.n1353 vdd.n1350 185
R15834 vdd.n1351 vdd.n1231 185
R15835 vdd.n1456 vdd.n1455 185
R15836 vdd.n1455 vdd.n1454 185
R15837 vdd.n2116 vdd.n2115 185
R15838 vdd.n2120 vdd.n1120 185
R15839 vdd.n1996 vdd.n1119 185
R15840 vdd.n1999 vdd.n1998 185
R15841 vdd.n2001 vdd.n2000 185
R15842 vdd.n2004 vdd.n2003 185
R15843 vdd.n2006 vdd.n2005 185
R15844 vdd.n2008 vdd.n1994 185
R15845 vdd.n2010 vdd.n2009 185
R15846 vdd.n2011 vdd.n1988 185
R15847 vdd.n2013 vdd.n2012 185
R15848 vdd.n2015 vdd.n1986 185
R15849 vdd.n2017 vdd.n2016 185
R15850 vdd.n2018 vdd.n1981 185
R15851 vdd.n2020 vdd.n2019 185
R15852 vdd.n2022 vdd.n1979 185
R15853 vdd.n2024 vdd.n2023 185
R15854 vdd.n2025 vdd.n1975 185
R15855 vdd.n2027 vdd.n2026 185
R15856 vdd.n2029 vdd.n1972 185
R15857 vdd.n2031 vdd.n2030 185
R15858 vdd.n1973 vdd.n1966 185
R15859 vdd.n2035 vdd.n1970 185
R15860 vdd.n2036 vdd.n1962 185
R15861 vdd.n2038 vdd.n2037 185
R15862 vdd.n2040 vdd.n1960 185
R15863 vdd.n2042 vdd.n2041 185
R15864 vdd.n2043 vdd.n1955 185
R15865 vdd.n2045 vdd.n2044 185
R15866 vdd.n2047 vdd.n1953 185
R15867 vdd.n2049 vdd.n2048 185
R15868 vdd.n2050 vdd.n1948 185
R15869 vdd.n2052 vdd.n2051 185
R15870 vdd.n2054 vdd.n1946 185
R15871 vdd.n2056 vdd.n2055 185
R15872 vdd.n2057 vdd.n1941 185
R15873 vdd.n2059 vdd.n2058 185
R15874 vdd.n2061 vdd.n1939 185
R15875 vdd.n2063 vdd.n2062 185
R15876 vdd.n2064 vdd.n1935 185
R15877 vdd.n2066 vdd.n2065 185
R15878 vdd.n2068 vdd.n1932 185
R15879 vdd.n2070 vdd.n2069 185
R15880 vdd.n1933 vdd.n1926 185
R15881 vdd.n2074 vdd.n1930 185
R15882 vdd.n2075 vdd.n1922 185
R15883 vdd.n2077 vdd.n2076 185
R15884 vdd.n2079 vdd.n1920 185
R15885 vdd.n2081 vdd.n2080 185
R15886 vdd.n2082 vdd.n1915 185
R15887 vdd.n2084 vdd.n2083 185
R15888 vdd.n2086 vdd.n1913 185
R15889 vdd.n2088 vdd.n2087 185
R15890 vdd.n2089 vdd.n1908 185
R15891 vdd.n2091 vdd.n2090 185
R15892 vdd.n2093 vdd.n1907 185
R15893 vdd.n2094 vdd.n1904 185
R15894 vdd.n2097 vdd.n2096 185
R15895 vdd.n1906 vdd.n1902 185
R15896 vdd.n2101 vdd.n1900 185
R15897 vdd.n2103 vdd.n2102 185
R15898 vdd.n2105 vdd.n1898 185
R15899 vdd.n2107 vdd.n2106 185
R15900 vdd.n2108 vdd.n1127 185
R15901 vdd.n2114 vdd.n1123 185
R15902 vdd.n2114 vdd.n2113 185
R15903 vdd.n1135 vdd.n1122 185
R15904 vdd.n1124 vdd.n1122 185
R15905 vdd.n1891 vdd.n1890 185
R15906 vdd.n1892 vdd.n1891 185
R15907 vdd.n1134 vdd.n1133 185
R15908 vdd.n1133 vdd.n1132 185
R15909 vdd.n1884 vdd.n1883 185
R15910 vdd.n1883 vdd.n1882 185
R15911 vdd.n1138 vdd.n1137 185
R15912 vdd.n1873 vdd.n1138 185
R15913 vdd.n1872 vdd.n1871 185
R15914 vdd.n1874 vdd.n1872 185
R15915 vdd.n1145 vdd.n1144 185
R15916 vdd.n1149 vdd.n1144 185
R15917 vdd.n1867 vdd.n1866 185
R15918 vdd.n1866 vdd.n1865 185
R15919 vdd.n1148 vdd.n1147 185
R15920 vdd.n1856 vdd.n1148 185
R15921 vdd.n1855 vdd.n1854 185
R15922 vdd.n1857 vdd.n1855 185
R15923 vdd.n1157 vdd.n1156 185
R15924 vdd.n1156 vdd.n1155 185
R15925 vdd.n1850 vdd.n1849 185
R15926 vdd.n1849 vdd.n1848 185
R15927 vdd.n1160 vdd.n1159 185
R15928 vdd.n1161 vdd.n1160 185
R15929 vdd.n1839 vdd.n1838 185
R15930 vdd.n1840 vdd.n1839 185
R15931 vdd.n1168 vdd.n1167 185
R15932 vdd.n1172 vdd.n1167 185
R15933 vdd.n1834 vdd.n1833 185
R15934 vdd.n1833 vdd.n1832 185
R15935 vdd.n1171 vdd.n1170 185
R15936 vdd.n1528 vdd.n1171 185
R15937 vdd.n1527 vdd.n1526 185
R15938 vdd.n1529 vdd.n1527 185
R15939 vdd.n1179 vdd.n1178 185
R15940 vdd.n1184 vdd.n1178 185
R15941 vdd.n1522 vdd.n1521 185
R15942 vdd.n1521 vdd.n1520 185
R15943 vdd.n1182 vdd.n1181 185
R15944 vdd.n1183 vdd.n1182 185
R15945 vdd.n1511 vdd.n1510 185
R15946 vdd.n1512 vdd.n1511 185
R15947 vdd.n1192 vdd.n1191 185
R15948 vdd.n1191 vdd.n1190 185
R15949 vdd.n1506 vdd.n1505 185
R15950 vdd.n1505 vdd.n1504 185
R15951 vdd.n1195 vdd.n1194 185
R15952 vdd.n1495 vdd.n1195 185
R15953 vdd.n1494 vdd.n1493 185
R15954 vdd.n1496 vdd.n1494 185
R15955 vdd.n1202 vdd.n1201 185
R15956 vdd.n1206 vdd.n1201 185
R15957 vdd.n1489 vdd.n1488 185
R15958 vdd.n1488 vdd.n1487 185
R15959 vdd.n1205 vdd.n1204 185
R15960 vdd.n1478 vdd.n1205 185
R15961 vdd.n1477 vdd.n1476 185
R15962 vdd.n1479 vdd.n1477 185
R15963 vdd.n1214 vdd.n1213 185
R15964 vdd.n1213 vdd.n1212 185
R15965 vdd.n1472 vdd.n1471 185
R15966 vdd.n1471 vdd.n1470 185
R15967 vdd.n1217 vdd.n1216 185
R15968 vdd.n1218 vdd.n1217 185
R15969 vdd.n1461 vdd.n1460 185
R15970 vdd.n1462 vdd.n1461 185
R15971 vdd.n1226 vdd.n1225 185
R15972 vdd.n1225 vdd.n1224 185
R15973 vdd.n958 vdd.n956 185
R15974 vdd.n2571 vdd.n956 185
R15975 vdd.n2493 vdd.n976 185
R15976 vdd.n976 vdd.n963 185
R15977 vdd.n2495 vdd.n2494 185
R15978 vdd.n2496 vdd.n2495 185
R15979 vdd.n2492 vdd.n975 185
R15980 vdd.n2251 vdd.n975 185
R15981 vdd.n2491 vdd.n2490 185
R15982 vdd.n2490 vdd.n2489 185
R15983 vdd.n978 vdd.n977 185
R15984 vdd.n979 vdd.n978 185
R15985 vdd.n2480 vdd.n2479 185
R15986 vdd.n2481 vdd.n2480 185
R15987 vdd.n2478 vdd.n989 185
R15988 vdd.n989 vdd.n986 185
R15989 vdd.n2477 vdd.n2476 185
R15990 vdd.n2476 vdd.n2475 185
R15991 vdd.n991 vdd.n990 185
R15992 vdd.n2263 vdd.n991 185
R15993 vdd.n2468 vdd.n2467 185
R15994 vdd.n2469 vdd.n2468 185
R15995 vdd.n2466 vdd.n999 185
R15996 vdd.n1004 vdd.n999 185
R15997 vdd.n2465 vdd.n2464 185
R15998 vdd.n2464 vdd.n2463 185
R15999 vdd.n1001 vdd.n1000 185
R16000 vdd.n1010 vdd.n1001 185
R16001 vdd.n2456 vdd.n2455 185
R16002 vdd.n2457 vdd.n2456 185
R16003 vdd.n2454 vdd.n1011 185
R16004 vdd.n2275 vdd.n1011 185
R16005 vdd.n2453 vdd.n2452 185
R16006 vdd.n2452 vdd.n2451 185
R16007 vdd.n1013 vdd.n1012 185
R16008 vdd.n1014 vdd.n1013 185
R16009 vdd.n2444 vdd.n2443 185
R16010 vdd.n2445 vdd.n2444 185
R16011 vdd.n2442 vdd.n1023 185
R16012 vdd.n1023 vdd.n1020 185
R16013 vdd.n2441 vdd.n2440 185
R16014 vdd.n2440 vdd.n2439 185
R16015 vdd.n1025 vdd.n1024 185
R16016 vdd.n1034 vdd.n1025 185
R16017 vdd.n2431 vdd.n2430 185
R16018 vdd.n2432 vdd.n2431 185
R16019 vdd.n2429 vdd.n1035 185
R16020 vdd.n1041 vdd.n1035 185
R16021 vdd.n2428 vdd.n2427 185
R16022 vdd.n2427 vdd.n2426 185
R16023 vdd.n1037 vdd.n1036 185
R16024 vdd.n1038 vdd.n1037 185
R16025 vdd.n2419 vdd.n2418 185
R16026 vdd.n2420 vdd.n2419 185
R16027 vdd.n2417 vdd.n1048 185
R16028 vdd.n1048 vdd.n1045 185
R16029 vdd.n2416 vdd.n2415 185
R16030 vdd.n2415 vdd.n2414 185
R16031 vdd.n1050 vdd.n1049 185
R16032 vdd.n1051 vdd.n1050 185
R16033 vdd.n2407 vdd.n2406 185
R16034 vdd.n2408 vdd.n2407 185
R16035 vdd.n2405 vdd.n1060 185
R16036 vdd.n1060 vdd.n1057 185
R16037 vdd.n2404 vdd.n2403 185
R16038 vdd.n2403 vdd.n2402 185
R16039 vdd.n1062 vdd.n1061 185
R16040 vdd.n1063 vdd.n1062 185
R16041 vdd.n2395 vdd.n2394 185
R16042 vdd.n2396 vdd.n2395 185
R16043 vdd.n2393 vdd.n1072 185
R16044 vdd.n1072 vdd.n1069 185
R16045 vdd.n2392 vdd.n2391 185
R16046 vdd.n2391 vdd.n2390 185
R16047 vdd.n1074 vdd.n1073 185
R16048 vdd.n1075 vdd.n1074 185
R16049 vdd.n2383 vdd.n2382 185
R16050 vdd.n2384 vdd.n2383 185
R16051 vdd.n2381 vdd.n1084 185
R16052 vdd.n2380 vdd.n2379 185
R16053 vdd.n2377 vdd.n1085 185
R16054 vdd.n2377 vdd.n1081 185
R16055 vdd.n2376 vdd.n2375 185
R16056 vdd.n2374 vdd.n2373 185
R16057 vdd.n2372 vdd.n1087 185
R16058 vdd.n2370 vdd.n2369 185
R16059 vdd.n2368 vdd.n1088 185
R16060 vdd.n2367 vdd.n2366 185
R16061 vdd.n2364 vdd.n1089 185
R16062 vdd.n2362 vdd.n2361 185
R16063 vdd.n2360 vdd.n1090 185
R16064 vdd.n2359 vdd.n2358 185
R16065 vdd.n2356 vdd.n1091 185
R16066 vdd.n2354 vdd.n2353 185
R16067 vdd.n2352 vdd.n1092 185
R16068 vdd.n2351 vdd.n2350 185
R16069 vdd.n2348 vdd.n1093 185
R16070 vdd.n2346 vdd.n2345 185
R16071 vdd.n2344 vdd.n1094 185
R16072 vdd.n2343 vdd.n2342 185
R16073 vdd.n2340 vdd.n1095 185
R16074 vdd.n2338 vdd.n2337 185
R16075 vdd.n2336 vdd.n1096 185
R16076 vdd.n2335 vdd.n2334 185
R16077 vdd.n2332 vdd.n1097 185
R16078 vdd.n2330 vdd.n2329 185
R16079 vdd.n2328 vdd.n1098 185
R16080 vdd.n2327 vdd.n2326 185
R16081 vdd.n2324 vdd.n1099 185
R16082 vdd.n2322 vdd.n2321 185
R16083 vdd.n2320 vdd.n1100 185
R16084 vdd.n2318 vdd.n2317 185
R16085 vdd.n2315 vdd.n1103 185
R16086 vdd.n2313 vdd.n2312 185
R16087 vdd.n2574 vdd.n2573 185
R16088 vdd.n2576 vdd.n2575 185
R16089 vdd.n2578 vdd.n2577 185
R16090 vdd.n2581 vdd.n2580 185
R16091 vdd.n2583 vdd.n2582 185
R16092 vdd.n2585 vdd.n2584 185
R16093 vdd.n2587 vdd.n2586 185
R16094 vdd.n2589 vdd.n2588 185
R16095 vdd.n2591 vdd.n2590 185
R16096 vdd.n2593 vdd.n2592 185
R16097 vdd.n2595 vdd.n2594 185
R16098 vdd.n2597 vdd.n2596 185
R16099 vdd.n2599 vdd.n2598 185
R16100 vdd.n2601 vdd.n2600 185
R16101 vdd.n2603 vdd.n2602 185
R16102 vdd.n2605 vdd.n2604 185
R16103 vdd.n2607 vdd.n2606 185
R16104 vdd.n2609 vdd.n2608 185
R16105 vdd.n2611 vdd.n2610 185
R16106 vdd.n2613 vdd.n2612 185
R16107 vdd.n2615 vdd.n2614 185
R16108 vdd.n2617 vdd.n2616 185
R16109 vdd.n2619 vdd.n2618 185
R16110 vdd.n2621 vdd.n2620 185
R16111 vdd.n2623 vdd.n2622 185
R16112 vdd.n2625 vdd.n2624 185
R16113 vdd.n2627 vdd.n2626 185
R16114 vdd.n2629 vdd.n2628 185
R16115 vdd.n2631 vdd.n2630 185
R16116 vdd.n2633 vdd.n2632 185
R16117 vdd.n2635 vdd.n2634 185
R16118 vdd.n2637 vdd.n2636 185
R16119 vdd.n2639 vdd.n2638 185
R16120 vdd.n2640 vdd.n957 185
R16121 vdd.n2642 vdd.n2641 185
R16122 vdd.n2643 vdd.n2642 185
R16123 vdd.n2572 vdd.n961 185
R16124 vdd.n2572 vdd.n2571 185
R16125 vdd.n2249 vdd.n962 185
R16126 vdd.n963 vdd.n962 185
R16127 vdd.n2250 vdd.n973 185
R16128 vdd.n2496 vdd.n973 185
R16129 vdd.n2253 vdd.n2252 185
R16130 vdd.n2252 vdd.n2251 185
R16131 vdd.n2254 vdd.n980 185
R16132 vdd.n2489 vdd.n980 185
R16133 vdd.n2256 vdd.n2255 185
R16134 vdd.n2255 vdd.n979 185
R16135 vdd.n2257 vdd.n987 185
R16136 vdd.n2481 vdd.n987 185
R16137 vdd.n2259 vdd.n2258 185
R16138 vdd.n2258 vdd.n986 185
R16139 vdd.n2260 vdd.n992 185
R16140 vdd.n2475 vdd.n992 185
R16141 vdd.n2262 vdd.n2261 185
R16142 vdd.n2263 vdd.n2262 185
R16143 vdd.n2248 vdd.n997 185
R16144 vdd.n2469 vdd.n997 185
R16145 vdd.n2247 vdd.n2246 185
R16146 vdd.n2246 vdd.n1004 185
R16147 vdd.n2245 vdd.n1002 185
R16148 vdd.n2463 vdd.n1002 185
R16149 vdd.n2244 vdd.n2243 185
R16150 vdd.n2243 vdd.n1010 185
R16151 vdd.n1104 vdd.n1008 185
R16152 vdd.n2457 vdd.n1008 185
R16153 vdd.n2277 vdd.n2276 185
R16154 vdd.n2276 vdd.n2275 185
R16155 vdd.n2278 vdd.n1015 185
R16156 vdd.n2451 vdd.n1015 185
R16157 vdd.n2280 vdd.n2279 185
R16158 vdd.n2279 vdd.n1014 185
R16159 vdd.n2281 vdd.n1021 185
R16160 vdd.n2445 vdd.n1021 185
R16161 vdd.n2283 vdd.n2282 185
R16162 vdd.n2282 vdd.n1020 185
R16163 vdd.n2284 vdd.n1026 185
R16164 vdd.n2439 vdd.n1026 185
R16165 vdd.n2286 vdd.n2285 185
R16166 vdd.n2285 vdd.n1034 185
R16167 vdd.n2287 vdd.n1032 185
R16168 vdd.n2432 vdd.n1032 185
R16169 vdd.n2289 vdd.n2288 185
R16170 vdd.n2288 vdd.n1041 185
R16171 vdd.n2290 vdd.n1039 185
R16172 vdd.n2426 vdd.n1039 185
R16173 vdd.n2292 vdd.n2291 185
R16174 vdd.n2291 vdd.n1038 185
R16175 vdd.n2293 vdd.n1046 185
R16176 vdd.n2420 vdd.n1046 185
R16177 vdd.n2295 vdd.n2294 185
R16178 vdd.n2294 vdd.n1045 185
R16179 vdd.n2296 vdd.n1052 185
R16180 vdd.n2414 vdd.n1052 185
R16181 vdd.n2298 vdd.n2297 185
R16182 vdd.n2297 vdd.n1051 185
R16183 vdd.n2299 vdd.n1058 185
R16184 vdd.n2408 vdd.n1058 185
R16185 vdd.n2301 vdd.n2300 185
R16186 vdd.n2300 vdd.n1057 185
R16187 vdd.n2302 vdd.n1064 185
R16188 vdd.n2402 vdd.n1064 185
R16189 vdd.n2304 vdd.n2303 185
R16190 vdd.n2303 vdd.n1063 185
R16191 vdd.n2305 vdd.n1070 185
R16192 vdd.n2396 vdd.n1070 185
R16193 vdd.n2307 vdd.n2306 185
R16194 vdd.n2306 vdd.n1069 185
R16195 vdd.n2308 vdd.n1076 185
R16196 vdd.n2390 vdd.n1076 185
R16197 vdd.n2310 vdd.n2309 185
R16198 vdd.n2309 vdd.n1075 185
R16199 vdd.n2311 vdd.n1082 185
R16200 vdd.n2384 vdd.n1082 185
R16201 vdd.n370 vdd.n369 185
R16202 vdd.n3436 vdd.n370 185
R16203 vdd.n3439 vdd.n3438 185
R16204 vdd.n3438 vdd.n3437 185
R16205 vdd.n3440 vdd.n364 185
R16206 vdd.n364 vdd.n363 185
R16207 vdd.n3442 vdd.n3441 185
R16208 vdd.n3443 vdd.n3442 185
R16209 vdd.n359 vdd.n358 185
R16210 vdd.n3444 vdd.n359 185
R16211 vdd.n3447 vdd.n3446 185
R16212 vdd.n3446 vdd.n3445 185
R16213 vdd.n3448 vdd.n353 185
R16214 vdd.n3418 vdd.n353 185
R16215 vdd.n3450 vdd.n3449 185
R16216 vdd.n3451 vdd.n3450 185
R16217 vdd.n348 vdd.n347 185
R16218 vdd.n3452 vdd.n348 185
R16219 vdd.n3455 vdd.n3454 185
R16220 vdd.n3454 vdd.n3453 185
R16221 vdd.n3456 vdd.n342 185
R16222 vdd.n349 vdd.n342 185
R16223 vdd.n3458 vdd.n3457 185
R16224 vdd.n3459 vdd.n3458 185
R16225 vdd.n338 vdd.n337 185
R16226 vdd.n3460 vdd.n338 185
R16227 vdd.n3463 vdd.n3462 185
R16228 vdd.n3462 vdd.n3461 185
R16229 vdd.n3464 vdd.n333 185
R16230 vdd.n333 vdd.n332 185
R16231 vdd.n3466 vdd.n3465 185
R16232 vdd.n3467 vdd.n3466 185
R16233 vdd.n327 vdd.n325 185
R16234 vdd.n3468 vdd.n327 185
R16235 vdd.n3471 vdd.n3470 185
R16236 vdd.n3470 vdd.n3469 185
R16237 vdd.n326 vdd.n324 185
R16238 vdd.n328 vdd.n326 185
R16239 vdd.n3394 vdd.n3393 185
R16240 vdd.n3395 vdd.n3394 185
R16241 vdd.n615 vdd.n614 185
R16242 vdd.n614 vdd.n613 185
R16243 vdd.n3389 vdd.n3388 185
R16244 vdd.n3388 vdd.n3387 185
R16245 vdd.n618 vdd.n617 185
R16246 vdd.n624 vdd.n618 185
R16247 vdd.n3375 vdd.n3374 185
R16248 vdd.n3376 vdd.n3375 185
R16249 vdd.n626 vdd.n625 185
R16250 vdd.n3367 vdd.n625 185
R16251 vdd.n3370 vdd.n3369 185
R16252 vdd.n3369 vdd.n3368 185
R16253 vdd.n629 vdd.n628 185
R16254 vdd.n636 vdd.n629 185
R16255 vdd.n3358 vdd.n3357 185
R16256 vdd.n3359 vdd.n3358 185
R16257 vdd.n638 vdd.n637 185
R16258 vdd.n637 vdd.n635 185
R16259 vdd.n3353 vdd.n3352 185
R16260 vdd.n3352 vdd.n3351 185
R16261 vdd.n641 vdd.n640 185
R16262 vdd.n642 vdd.n641 185
R16263 vdd.n3342 vdd.n3341 185
R16264 vdd.n3343 vdd.n3342 185
R16265 vdd.n650 vdd.n649 185
R16266 vdd.n649 vdd.n648 185
R16267 vdd.n3337 vdd.n3336 185
R16268 vdd.n3336 vdd.n3335 185
R16269 vdd.n653 vdd.n652 185
R16270 vdd.n659 vdd.n653 185
R16271 vdd.n3326 vdd.n3325 185
R16272 vdd.n3327 vdd.n3326 185
R16273 vdd.n3322 vdd.n660 185
R16274 vdd.n3321 vdd.n3320 185
R16275 vdd.n3318 vdd.n662 185
R16276 vdd.n3318 vdd.n658 185
R16277 vdd.n3317 vdd.n3316 185
R16278 vdd.n3315 vdd.n3314 185
R16279 vdd.n3313 vdd.n3312 185
R16280 vdd.n3311 vdd.n3310 185
R16281 vdd.n3309 vdd.n668 185
R16282 vdd.n3307 vdd.n3306 185
R16283 vdd.n3305 vdd.n669 185
R16284 vdd.n3304 vdd.n3303 185
R16285 vdd.n3301 vdd.n674 185
R16286 vdd.n3299 vdd.n3298 185
R16287 vdd.n3297 vdd.n675 185
R16288 vdd.n3296 vdd.n3295 185
R16289 vdd.n3293 vdd.n680 185
R16290 vdd.n3291 vdd.n3290 185
R16291 vdd.n3289 vdd.n681 185
R16292 vdd.n3288 vdd.n3287 185
R16293 vdd.n3285 vdd.n688 185
R16294 vdd.n3283 vdd.n3282 185
R16295 vdd.n3281 vdd.n689 185
R16296 vdd.n3280 vdd.n3279 185
R16297 vdd.n3277 vdd.n694 185
R16298 vdd.n3275 vdd.n3274 185
R16299 vdd.n3273 vdd.n695 185
R16300 vdd.n3272 vdd.n3271 185
R16301 vdd.n3269 vdd.n700 185
R16302 vdd.n3267 vdd.n3266 185
R16303 vdd.n3265 vdd.n701 185
R16304 vdd.n3264 vdd.n3263 185
R16305 vdd.n3261 vdd.n706 185
R16306 vdd.n3259 vdd.n3258 185
R16307 vdd.n3257 vdd.n707 185
R16308 vdd.n3256 vdd.n3255 185
R16309 vdd.n3253 vdd.n712 185
R16310 vdd.n3251 vdd.n3250 185
R16311 vdd.n3249 vdd.n713 185
R16312 vdd.n3248 vdd.n3247 185
R16313 vdd.n3245 vdd.n718 185
R16314 vdd.n3243 vdd.n3242 185
R16315 vdd.n3241 vdd.n719 185
R16316 vdd.n728 vdd.n722 185
R16317 vdd.n3237 vdd.n3236 185
R16318 vdd.n3234 vdd.n726 185
R16319 vdd.n3233 vdd.n3232 185
R16320 vdd.n3231 vdd.n3230 185
R16321 vdd.n3229 vdd.n732 185
R16322 vdd.n3227 vdd.n3226 185
R16323 vdd.n3225 vdd.n733 185
R16324 vdd.n3224 vdd.n3223 185
R16325 vdd.n3221 vdd.n738 185
R16326 vdd.n3219 vdd.n3218 185
R16327 vdd.n3217 vdd.n739 185
R16328 vdd.n3216 vdd.n3215 185
R16329 vdd.n3213 vdd.n744 185
R16330 vdd.n3211 vdd.n3210 185
R16331 vdd.n3209 vdd.n745 185
R16332 vdd.n3208 vdd.n3207 185
R16333 vdd.n3205 vdd.n3204 185
R16334 vdd.n3203 vdd.n3202 185
R16335 vdd.n3201 vdd.n3200 185
R16336 vdd.n3199 vdd.n3198 185
R16337 vdd.n3194 vdd.n657 185
R16338 vdd.n658 vdd.n657 185
R16339 vdd.n3433 vdd.n3432 185
R16340 vdd.n599 vdd.n404 185
R16341 vdd.n598 vdd.n597 185
R16342 vdd.n596 vdd.n595 185
R16343 vdd.n594 vdd.n409 185
R16344 vdd.n590 vdd.n589 185
R16345 vdd.n588 vdd.n587 185
R16346 vdd.n586 vdd.n585 185
R16347 vdd.n584 vdd.n411 185
R16348 vdd.n580 vdd.n579 185
R16349 vdd.n578 vdd.n577 185
R16350 vdd.n576 vdd.n575 185
R16351 vdd.n574 vdd.n413 185
R16352 vdd.n570 vdd.n569 185
R16353 vdd.n568 vdd.n567 185
R16354 vdd.n566 vdd.n565 185
R16355 vdd.n564 vdd.n415 185
R16356 vdd.n560 vdd.n559 185
R16357 vdd.n558 vdd.n557 185
R16358 vdd.n556 vdd.n555 185
R16359 vdd.n554 vdd.n417 185
R16360 vdd.n550 vdd.n549 185
R16361 vdd.n548 vdd.n547 185
R16362 vdd.n546 vdd.n545 185
R16363 vdd.n544 vdd.n421 185
R16364 vdd.n540 vdd.n539 185
R16365 vdd.n538 vdd.n537 185
R16366 vdd.n536 vdd.n535 185
R16367 vdd.n534 vdd.n423 185
R16368 vdd.n530 vdd.n529 185
R16369 vdd.n528 vdd.n527 185
R16370 vdd.n526 vdd.n525 185
R16371 vdd.n524 vdd.n425 185
R16372 vdd.n520 vdd.n519 185
R16373 vdd.n518 vdd.n517 185
R16374 vdd.n516 vdd.n515 185
R16375 vdd.n514 vdd.n427 185
R16376 vdd.n510 vdd.n509 185
R16377 vdd.n508 vdd.n507 185
R16378 vdd.n506 vdd.n505 185
R16379 vdd.n504 vdd.n429 185
R16380 vdd.n500 vdd.n499 185
R16381 vdd.n498 vdd.n497 185
R16382 vdd.n496 vdd.n495 185
R16383 vdd.n494 vdd.n433 185
R16384 vdd.n490 vdd.n489 185
R16385 vdd.n488 vdd.n487 185
R16386 vdd.n486 vdd.n485 185
R16387 vdd.n484 vdd.n435 185
R16388 vdd.n480 vdd.n479 185
R16389 vdd.n478 vdd.n477 185
R16390 vdd.n476 vdd.n475 185
R16391 vdd.n474 vdd.n437 185
R16392 vdd.n470 vdd.n469 185
R16393 vdd.n468 vdd.n467 185
R16394 vdd.n466 vdd.n465 185
R16395 vdd.n464 vdd.n439 185
R16396 vdd.n460 vdd.n459 185
R16397 vdd.n458 vdd.n457 185
R16398 vdd.n456 vdd.n455 185
R16399 vdd.n454 vdd.n441 185
R16400 vdd.n450 vdd.n449 185
R16401 vdd.n448 vdd.n447 185
R16402 vdd.n446 vdd.n445 185
R16403 vdd.n3429 vdd.n372 185
R16404 vdd.n3436 vdd.n372 185
R16405 vdd.n3428 vdd.n371 185
R16406 vdd.n3437 vdd.n371 185
R16407 vdd.n3427 vdd.n3426 185
R16408 vdd.n3426 vdd.n363 185
R16409 vdd.n602 vdd.n362 185
R16410 vdd.n3443 vdd.n362 185
R16411 vdd.n3422 vdd.n361 185
R16412 vdd.n3444 vdd.n361 185
R16413 vdd.n3421 vdd.n360 185
R16414 vdd.n3445 vdd.n360 185
R16415 vdd.n3420 vdd.n3419 185
R16416 vdd.n3419 vdd.n3418 185
R16417 vdd.n604 vdd.n352 185
R16418 vdd.n3451 vdd.n352 185
R16419 vdd.n3414 vdd.n351 185
R16420 vdd.n3452 vdd.n351 185
R16421 vdd.n3413 vdd.n350 185
R16422 vdd.n3453 vdd.n350 185
R16423 vdd.n3412 vdd.n3411 185
R16424 vdd.n3411 vdd.n349 185
R16425 vdd.n606 vdd.n341 185
R16426 vdd.n3459 vdd.n341 185
R16427 vdd.n3407 vdd.n340 185
R16428 vdd.n3460 vdd.n340 185
R16429 vdd.n3406 vdd.n339 185
R16430 vdd.n3461 vdd.n339 185
R16431 vdd.n3405 vdd.n3404 185
R16432 vdd.n3404 vdd.n332 185
R16433 vdd.n608 vdd.n331 185
R16434 vdd.n3467 vdd.n331 185
R16435 vdd.n3400 vdd.n330 185
R16436 vdd.n3468 vdd.n330 185
R16437 vdd.n3399 vdd.n329 185
R16438 vdd.n3469 vdd.n329 185
R16439 vdd.n3398 vdd.n3397 185
R16440 vdd.n3397 vdd.n328 185
R16441 vdd.n3396 vdd.n610 185
R16442 vdd.n3396 vdd.n3395 185
R16443 vdd.n3384 vdd.n612 185
R16444 vdd.n613 vdd.n612 185
R16445 vdd.n3386 vdd.n3385 185
R16446 vdd.n3387 vdd.n3386 185
R16447 vdd.n620 vdd.n619 185
R16448 vdd.n624 vdd.n619 185
R16449 vdd.n3378 vdd.n3377 185
R16450 vdd.n3377 vdd.n3376 185
R16451 vdd.n623 vdd.n622 185
R16452 vdd.n3367 vdd.n623 185
R16453 vdd.n3366 vdd.n3365 185
R16454 vdd.n3368 vdd.n3366 185
R16455 vdd.n631 vdd.n630 185
R16456 vdd.n636 vdd.n630 185
R16457 vdd.n3361 vdd.n3360 185
R16458 vdd.n3360 vdd.n3359 185
R16459 vdd.n634 vdd.n633 185
R16460 vdd.n635 vdd.n634 185
R16461 vdd.n3350 vdd.n3349 185
R16462 vdd.n3351 vdd.n3350 185
R16463 vdd.n644 vdd.n643 185
R16464 vdd.n643 vdd.n642 185
R16465 vdd.n3345 vdd.n3344 185
R16466 vdd.n3344 vdd.n3343 185
R16467 vdd.n647 vdd.n646 185
R16468 vdd.n648 vdd.n647 185
R16469 vdd.n3334 vdd.n3333 185
R16470 vdd.n3335 vdd.n3334 185
R16471 vdd.n655 vdd.n654 185
R16472 vdd.n659 vdd.n654 185
R16473 vdd.n3329 vdd.n3328 185
R16474 vdd.n3328 vdd.n3327 185
R16475 vdd.n2931 vdd.n918 185
R16476 vdd.n2930 vdd.n2929 185
R16477 vdd.n920 vdd.n919 185
R16478 vdd.n2927 vdd.n920 185
R16479 vdd.n2750 vdd.n2749 185
R16480 vdd.n2752 vdd.n2751 185
R16481 vdd.n2754 vdd.n2753 185
R16482 vdd.n2756 vdd.n2755 185
R16483 vdd.n2758 vdd.n2757 185
R16484 vdd.n2760 vdd.n2759 185
R16485 vdd.n2762 vdd.n2761 185
R16486 vdd.n2764 vdd.n2763 185
R16487 vdd.n2766 vdd.n2765 185
R16488 vdd.n2768 vdd.n2767 185
R16489 vdd.n2770 vdd.n2769 185
R16490 vdd.n2772 vdd.n2771 185
R16491 vdd.n2774 vdd.n2773 185
R16492 vdd.n2776 vdd.n2775 185
R16493 vdd.n2778 vdd.n2777 185
R16494 vdd.n2780 vdd.n2779 185
R16495 vdd.n2782 vdd.n2781 185
R16496 vdd.n2784 vdd.n2783 185
R16497 vdd.n2786 vdd.n2785 185
R16498 vdd.n2788 vdd.n2787 185
R16499 vdd.n2790 vdd.n2789 185
R16500 vdd.n2792 vdd.n2791 185
R16501 vdd.n2794 vdd.n2793 185
R16502 vdd.n2796 vdd.n2795 185
R16503 vdd.n2798 vdd.n2797 185
R16504 vdd.n2800 vdd.n2799 185
R16505 vdd.n2802 vdd.n2801 185
R16506 vdd.n2804 vdd.n2803 185
R16507 vdd.n2806 vdd.n2805 185
R16508 vdd.n2809 vdd.n2808 185
R16509 vdd.n2811 vdd.n2810 185
R16510 vdd.n2813 vdd.n2812 185
R16511 vdd.n3095 vdd.n3094 185
R16512 vdd.n3096 vdd.n803 185
R16513 vdd.n3098 vdd.n3097 185
R16514 vdd.n3100 vdd.n801 185
R16515 vdd.n3102 vdd.n3101 185
R16516 vdd.n3103 vdd.n800 185
R16517 vdd.n3105 vdd.n3104 185
R16518 vdd.n3107 vdd.n798 185
R16519 vdd.n3109 vdd.n3108 185
R16520 vdd.n3110 vdd.n797 185
R16521 vdd.n3112 vdd.n3111 185
R16522 vdd.n3114 vdd.n795 185
R16523 vdd.n3116 vdd.n3115 185
R16524 vdd.n3117 vdd.n794 185
R16525 vdd.n3119 vdd.n3118 185
R16526 vdd.n3121 vdd.n792 185
R16527 vdd.n3123 vdd.n3122 185
R16528 vdd.n3125 vdd.n791 185
R16529 vdd.n3127 vdd.n3126 185
R16530 vdd.n3129 vdd.n789 185
R16531 vdd.n3131 vdd.n3130 185
R16532 vdd.n3132 vdd.n788 185
R16533 vdd.n3134 vdd.n3133 185
R16534 vdd.n3136 vdd.n786 185
R16535 vdd.n3138 vdd.n3137 185
R16536 vdd.n3139 vdd.n785 185
R16537 vdd.n3141 vdd.n3140 185
R16538 vdd.n3143 vdd.n783 185
R16539 vdd.n3145 vdd.n3144 185
R16540 vdd.n3146 vdd.n782 185
R16541 vdd.n3148 vdd.n3147 185
R16542 vdd.n3150 vdd.n781 185
R16543 vdd.n3151 vdd.n780 185
R16544 vdd.n3154 vdd.n3153 185
R16545 vdd.n3155 vdd.n778 185
R16546 vdd.n778 vdd.n756 185
R16547 vdd.n3092 vdd.n775 185
R16548 vdd.n3158 vdd.n775 185
R16549 vdd.n3091 vdd.n3090 185
R16550 vdd.n3090 vdd.n774 185
R16551 vdd.n3089 vdd.n807 185
R16552 vdd.n3089 vdd.n3088 185
R16553 vdd.n2863 vdd.n808 185
R16554 vdd.n817 vdd.n808 185
R16555 vdd.n2864 vdd.n815 185
R16556 vdd.n3082 vdd.n815 185
R16557 vdd.n2866 vdd.n2865 185
R16558 vdd.n2865 vdd.n814 185
R16559 vdd.n2867 vdd.n823 185
R16560 vdd.n3031 vdd.n823 185
R16561 vdd.n2869 vdd.n2868 185
R16562 vdd.n2868 vdd.n822 185
R16563 vdd.n2870 vdd.n828 185
R16564 vdd.n3025 vdd.n828 185
R16565 vdd.n2872 vdd.n2871 185
R16566 vdd.n2871 vdd.n835 185
R16567 vdd.n2873 vdd.n833 185
R16568 vdd.n3019 vdd.n833 185
R16569 vdd.n2875 vdd.n2874 185
R16570 vdd.n2874 vdd.n841 185
R16571 vdd.n2876 vdd.n839 185
R16572 vdd.n3013 vdd.n839 185
R16573 vdd.n2878 vdd.n2877 185
R16574 vdd.n2877 vdd.n848 185
R16575 vdd.n2879 vdd.n846 185
R16576 vdd.n3007 vdd.n846 185
R16577 vdd.n2881 vdd.n2880 185
R16578 vdd.n2880 vdd.n845 185
R16579 vdd.n2882 vdd.n853 185
R16580 vdd.n3001 vdd.n853 185
R16581 vdd.n2884 vdd.n2883 185
R16582 vdd.n2883 vdd.n852 185
R16583 vdd.n2885 vdd.n860 185
R16584 vdd.n2994 vdd.n860 185
R16585 vdd.n2887 vdd.n2886 185
R16586 vdd.n2886 vdd.n859 185
R16587 vdd.n2888 vdd.n865 185
R16588 vdd.n2988 vdd.n865 185
R16589 vdd.n2890 vdd.n2889 185
R16590 vdd.n2889 vdd.n872 185
R16591 vdd.n2891 vdd.n870 185
R16592 vdd.n2982 vdd.n870 185
R16593 vdd.n2893 vdd.n2892 185
R16594 vdd.n2894 vdd.n2893 185
R16595 vdd.n2862 vdd.n877 185
R16596 vdd.n2976 vdd.n877 185
R16597 vdd.n2861 vdd.n2860 185
R16598 vdd.n2860 vdd.n876 185
R16599 vdd.n2859 vdd.n883 185
R16600 vdd.n2970 vdd.n883 185
R16601 vdd.n2858 vdd.n2857 185
R16602 vdd.n2857 vdd.n882 185
R16603 vdd.n2818 vdd.n888 185
R16604 vdd.n2964 vdd.n888 185
R16605 vdd.n2908 vdd.n2907 185
R16606 vdd.n2907 vdd.n2906 185
R16607 vdd.n2909 vdd.n893 185
R16608 vdd.n2958 vdd.n893 185
R16609 vdd.n2911 vdd.n2910 185
R16610 vdd.n2910 vdd.n901 185
R16611 vdd.n2912 vdd.n899 185
R16612 vdd.n2952 vdd.n899 185
R16613 vdd.n2914 vdd.n2913 185
R16614 vdd.n2913 vdd.n898 185
R16615 vdd.n2915 vdd.n905 185
R16616 vdd.n2946 vdd.n905 185
R16617 vdd.n2917 vdd.n2916 185
R16618 vdd.n2918 vdd.n2917 185
R16619 vdd.n2817 vdd.n910 185
R16620 vdd.n2940 vdd.n910 185
R16621 vdd.n2816 vdd.n2815 185
R16622 vdd.n2815 vdd.n917 185
R16623 vdd.n2814 vdd.n915 185
R16624 vdd.n2934 vdd.n915 185
R16625 vdd.n2933 vdd.n2932 185
R16626 vdd.n2934 vdd.n2933 185
R16627 vdd.n909 vdd.n908 185
R16628 vdd.n917 vdd.n909 185
R16629 vdd.n2942 vdd.n2941 185
R16630 vdd.n2941 vdd.n2940 185
R16631 vdd.n2943 vdd.n907 185
R16632 vdd.n2918 vdd.n907 185
R16633 vdd.n2945 vdd.n2944 185
R16634 vdd.n2946 vdd.n2945 185
R16635 vdd.n897 vdd.n896 185
R16636 vdd.n898 vdd.n897 185
R16637 vdd.n2954 vdd.n2953 185
R16638 vdd.n2953 vdd.n2952 185
R16639 vdd.n2955 vdd.n895 185
R16640 vdd.n901 vdd.n895 185
R16641 vdd.n2957 vdd.n2956 185
R16642 vdd.n2958 vdd.n2957 185
R16643 vdd.n887 vdd.n886 185
R16644 vdd.n2906 vdd.n887 185
R16645 vdd.n2966 vdd.n2965 185
R16646 vdd.n2965 vdd.n2964 185
R16647 vdd.n2967 vdd.n885 185
R16648 vdd.n885 vdd.n882 185
R16649 vdd.n2969 vdd.n2968 185
R16650 vdd.n2970 vdd.n2969 185
R16651 vdd.n875 vdd.n874 185
R16652 vdd.n876 vdd.n875 185
R16653 vdd.n2978 vdd.n2977 185
R16654 vdd.n2977 vdd.n2976 185
R16655 vdd.n2979 vdd.n873 185
R16656 vdd.n2894 vdd.n873 185
R16657 vdd.n2981 vdd.n2980 185
R16658 vdd.n2982 vdd.n2981 185
R16659 vdd.n864 vdd.n863 185
R16660 vdd.n872 vdd.n864 185
R16661 vdd.n2990 vdd.n2989 185
R16662 vdd.n2989 vdd.n2988 185
R16663 vdd.n2991 vdd.n862 185
R16664 vdd.n862 vdd.n859 185
R16665 vdd.n2993 vdd.n2992 185
R16666 vdd.n2994 vdd.n2993 185
R16667 vdd.n851 vdd.n850 185
R16668 vdd.n852 vdd.n851 185
R16669 vdd.n3003 vdd.n3002 185
R16670 vdd.n3002 vdd.n3001 185
R16671 vdd.n3004 vdd.n849 185
R16672 vdd.n849 vdd.n845 185
R16673 vdd.n3006 vdd.n3005 185
R16674 vdd.n3007 vdd.n3006 185
R16675 vdd.n838 vdd.n837 185
R16676 vdd.n848 vdd.n838 185
R16677 vdd.n3015 vdd.n3014 185
R16678 vdd.n3014 vdd.n3013 185
R16679 vdd.n3016 vdd.n836 185
R16680 vdd.n841 vdd.n836 185
R16681 vdd.n3018 vdd.n3017 185
R16682 vdd.n3019 vdd.n3018 185
R16683 vdd.n827 vdd.n826 185
R16684 vdd.n835 vdd.n827 185
R16685 vdd.n3027 vdd.n3026 185
R16686 vdd.n3026 vdd.n3025 185
R16687 vdd.n3028 vdd.n825 185
R16688 vdd.n825 vdd.n822 185
R16689 vdd.n3030 vdd.n3029 185
R16690 vdd.n3031 vdd.n3030 185
R16691 vdd.n813 vdd.n812 185
R16692 vdd.n814 vdd.n813 185
R16693 vdd.n3084 vdd.n3083 185
R16694 vdd.n3083 vdd.n3082 185
R16695 vdd.n3085 vdd.n811 185
R16696 vdd.n817 vdd.n811 185
R16697 vdd.n3087 vdd.n3086 185
R16698 vdd.n3088 vdd.n3087 185
R16699 vdd.n779 vdd.n777 185
R16700 vdd.n777 vdd.n774 185
R16701 vdd.n3157 vdd.n3156 185
R16702 vdd.n3158 vdd.n3157 185
R16703 vdd.n2570 vdd.n2569 185
R16704 vdd.n2571 vdd.n2570 185
R16705 vdd.n967 vdd.n965 185
R16706 vdd.n965 vdd.n963 185
R16707 vdd.n2485 vdd.n974 185
R16708 vdd.n2496 vdd.n974 185
R16709 vdd.n2486 vdd.n983 185
R16710 vdd.n2251 vdd.n983 185
R16711 vdd.n2488 vdd.n2487 185
R16712 vdd.n2489 vdd.n2488 185
R16713 vdd.n2484 vdd.n982 185
R16714 vdd.n982 vdd.n979 185
R16715 vdd.n2483 vdd.n2482 185
R16716 vdd.n2482 vdd.n2481 185
R16717 vdd.n985 vdd.n984 185
R16718 vdd.n986 vdd.n985 185
R16719 vdd.n2474 vdd.n2473 185
R16720 vdd.n2475 vdd.n2474 185
R16721 vdd.n2472 vdd.n994 185
R16722 vdd.n2263 vdd.n994 185
R16723 vdd.n2471 vdd.n2470 185
R16724 vdd.n2470 vdd.n2469 185
R16725 vdd.n996 vdd.n995 185
R16726 vdd.n1004 vdd.n996 185
R16727 vdd.n2462 vdd.n2461 185
R16728 vdd.n2463 vdd.n2462 185
R16729 vdd.n2460 vdd.n1005 185
R16730 vdd.n1010 vdd.n1005 185
R16731 vdd.n2459 vdd.n2458 185
R16732 vdd.n2458 vdd.n2457 185
R16733 vdd.n1007 vdd.n1006 185
R16734 vdd.n2275 vdd.n1007 185
R16735 vdd.n2450 vdd.n2449 185
R16736 vdd.n2451 vdd.n2450 185
R16737 vdd.n2448 vdd.n1017 185
R16738 vdd.n1017 vdd.n1014 185
R16739 vdd.n2447 vdd.n2446 185
R16740 vdd.n2446 vdd.n2445 185
R16741 vdd.n1019 vdd.n1018 185
R16742 vdd.n1020 vdd.n1019 185
R16743 vdd.n2438 vdd.n2437 185
R16744 vdd.n2439 vdd.n2438 185
R16745 vdd.n2435 vdd.n1028 185
R16746 vdd.n1034 vdd.n1028 185
R16747 vdd.n2434 vdd.n2433 185
R16748 vdd.n2433 vdd.n2432 185
R16749 vdd.n1031 vdd.n1030 185
R16750 vdd.n1041 vdd.n1031 185
R16751 vdd.n2425 vdd.n2424 185
R16752 vdd.n2426 vdd.n2425 185
R16753 vdd.n2423 vdd.n1042 185
R16754 vdd.n1042 vdd.n1038 185
R16755 vdd.n2422 vdd.n2421 185
R16756 vdd.n2421 vdd.n2420 185
R16757 vdd.n1044 vdd.n1043 185
R16758 vdd.n1045 vdd.n1044 185
R16759 vdd.n2413 vdd.n2412 185
R16760 vdd.n2414 vdd.n2413 185
R16761 vdd.n2411 vdd.n1054 185
R16762 vdd.n1054 vdd.n1051 185
R16763 vdd.n2410 vdd.n2409 185
R16764 vdd.n2409 vdd.n2408 185
R16765 vdd.n1056 vdd.n1055 185
R16766 vdd.n1057 vdd.n1056 185
R16767 vdd.n2401 vdd.n2400 185
R16768 vdd.n2402 vdd.n2401 185
R16769 vdd.n2399 vdd.n1066 185
R16770 vdd.n1066 vdd.n1063 185
R16771 vdd.n2398 vdd.n2397 185
R16772 vdd.n2397 vdd.n2396 185
R16773 vdd.n1068 vdd.n1067 185
R16774 vdd.n1069 vdd.n1068 185
R16775 vdd.n2389 vdd.n2388 185
R16776 vdd.n2390 vdd.n2389 185
R16777 vdd.n2387 vdd.n1078 185
R16778 vdd.n1078 vdd.n1075 185
R16779 vdd.n2386 vdd.n2385 185
R16780 vdd.n2385 vdd.n2384 185
R16781 vdd.n2501 vdd.n938 185
R16782 vdd.n2643 vdd.n938 185
R16783 vdd.n2503 vdd.n2502 185
R16784 vdd.n2505 vdd.n2504 185
R16785 vdd.n2507 vdd.n2506 185
R16786 vdd.n2509 vdd.n2508 185
R16787 vdd.n2511 vdd.n2510 185
R16788 vdd.n2513 vdd.n2512 185
R16789 vdd.n2515 vdd.n2514 185
R16790 vdd.n2517 vdd.n2516 185
R16791 vdd.n2519 vdd.n2518 185
R16792 vdd.n2521 vdd.n2520 185
R16793 vdd.n2523 vdd.n2522 185
R16794 vdd.n2525 vdd.n2524 185
R16795 vdd.n2527 vdd.n2526 185
R16796 vdd.n2529 vdd.n2528 185
R16797 vdd.n2531 vdd.n2530 185
R16798 vdd.n2533 vdd.n2532 185
R16799 vdd.n2535 vdd.n2534 185
R16800 vdd.n2537 vdd.n2536 185
R16801 vdd.n2539 vdd.n2538 185
R16802 vdd.n2541 vdd.n2540 185
R16803 vdd.n2543 vdd.n2542 185
R16804 vdd.n2545 vdd.n2544 185
R16805 vdd.n2547 vdd.n2546 185
R16806 vdd.n2549 vdd.n2548 185
R16807 vdd.n2551 vdd.n2550 185
R16808 vdd.n2553 vdd.n2552 185
R16809 vdd.n2555 vdd.n2554 185
R16810 vdd.n2557 vdd.n2556 185
R16811 vdd.n2559 vdd.n2558 185
R16812 vdd.n2561 vdd.n2560 185
R16813 vdd.n2563 vdd.n2562 185
R16814 vdd.n2565 vdd.n2564 185
R16815 vdd.n2567 vdd.n2566 185
R16816 vdd.n2568 vdd.n966 185
R16817 vdd.n2500 vdd.n964 185
R16818 vdd.n2571 vdd.n964 185
R16819 vdd.n2499 vdd.n2498 185
R16820 vdd.n2498 vdd.n963 185
R16821 vdd.n2497 vdd.n971 185
R16822 vdd.n2497 vdd.n2496 185
R16823 vdd.n2235 vdd.n972 185
R16824 vdd.n2251 vdd.n972 185
R16825 vdd.n2236 vdd.n981 185
R16826 vdd.n2489 vdd.n981 185
R16827 vdd.n2238 vdd.n2237 185
R16828 vdd.n2237 vdd.n979 185
R16829 vdd.n2239 vdd.n988 185
R16830 vdd.n2481 vdd.n988 185
R16831 vdd.n2241 vdd.n2240 185
R16832 vdd.n2240 vdd.n986 185
R16833 vdd.n2242 vdd.n993 185
R16834 vdd.n2475 vdd.n993 185
R16835 vdd.n2265 vdd.n2264 185
R16836 vdd.n2264 vdd.n2263 185
R16837 vdd.n2266 vdd.n998 185
R16838 vdd.n2469 vdd.n998 185
R16839 vdd.n2268 vdd.n2267 185
R16840 vdd.n2267 vdd.n1004 185
R16841 vdd.n2269 vdd.n1003 185
R16842 vdd.n2463 vdd.n1003 185
R16843 vdd.n2271 vdd.n2270 185
R16844 vdd.n2270 vdd.n1010 185
R16845 vdd.n2272 vdd.n1009 185
R16846 vdd.n2457 vdd.n1009 185
R16847 vdd.n2274 vdd.n2273 185
R16848 vdd.n2275 vdd.n2274 185
R16849 vdd.n2234 vdd.n1016 185
R16850 vdd.n2451 vdd.n1016 185
R16851 vdd.n2233 vdd.n2232 185
R16852 vdd.n2232 vdd.n1014 185
R16853 vdd.n2231 vdd.n1022 185
R16854 vdd.n2445 vdd.n1022 185
R16855 vdd.n2230 vdd.n2229 185
R16856 vdd.n2229 vdd.n1020 185
R16857 vdd.n2228 vdd.n1027 185
R16858 vdd.n2439 vdd.n1027 185
R16859 vdd.n2227 vdd.n2226 185
R16860 vdd.n2226 vdd.n1034 185
R16861 vdd.n2225 vdd.n1033 185
R16862 vdd.n2432 vdd.n1033 185
R16863 vdd.n2224 vdd.n2223 185
R16864 vdd.n2223 vdd.n1041 185
R16865 vdd.n2222 vdd.n1040 185
R16866 vdd.n2426 vdd.n1040 185
R16867 vdd.n2221 vdd.n2220 185
R16868 vdd.n2220 vdd.n1038 185
R16869 vdd.n2219 vdd.n1047 185
R16870 vdd.n2420 vdd.n1047 185
R16871 vdd.n2218 vdd.n2217 185
R16872 vdd.n2217 vdd.n1045 185
R16873 vdd.n2216 vdd.n1053 185
R16874 vdd.n2414 vdd.n1053 185
R16875 vdd.n2215 vdd.n2214 185
R16876 vdd.n2214 vdd.n1051 185
R16877 vdd.n2213 vdd.n1059 185
R16878 vdd.n2408 vdd.n1059 185
R16879 vdd.n2212 vdd.n2211 185
R16880 vdd.n2211 vdd.n1057 185
R16881 vdd.n2210 vdd.n1065 185
R16882 vdd.n2402 vdd.n1065 185
R16883 vdd.n2209 vdd.n2208 185
R16884 vdd.n2208 vdd.n1063 185
R16885 vdd.n2207 vdd.n1071 185
R16886 vdd.n2396 vdd.n1071 185
R16887 vdd.n2206 vdd.n2205 185
R16888 vdd.n2205 vdd.n1069 185
R16889 vdd.n2204 vdd.n1077 185
R16890 vdd.n2390 vdd.n1077 185
R16891 vdd.n2203 vdd.n2202 185
R16892 vdd.n2202 vdd.n1075 185
R16893 vdd.n2201 vdd.n1083 185
R16894 vdd.n2384 vdd.n1083 185
R16895 vdd.n1080 vdd.n1079 185
R16896 vdd.n2133 vdd.n2131 185
R16897 vdd.n2136 vdd.n2135 185
R16898 vdd.n2137 vdd.n2130 185
R16899 vdd.n2139 vdd.n2138 185
R16900 vdd.n2141 vdd.n2129 185
R16901 vdd.n2144 vdd.n2143 185
R16902 vdd.n2145 vdd.n2128 185
R16903 vdd.n2147 vdd.n2146 185
R16904 vdd.n2149 vdd.n2127 185
R16905 vdd.n2152 vdd.n2151 185
R16906 vdd.n2153 vdd.n2126 185
R16907 vdd.n2155 vdd.n2154 185
R16908 vdd.n2157 vdd.n2125 185
R16909 vdd.n2160 vdd.n2159 185
R16910 vdd.n2161 vdd.n2124 185
R16911 vdd.n2163 vdd.n2162 185
R16912 vdd.n2165 vdd.n2123 185
R16913 vdd.n2168 vdd.n2167 185
R16914 vdd.n2169 vdd.n1114 185
R16915 vdd.n2171 vdd.n2170 185
R16916 vdd.n2173 vdd.n1113 185
R16917 vdd.n2176 vdd.n2175 185
R16918 vdd.n2177 vdd.n1112 185
R16919 vdd.n2179 vdd.n2178 185
R16920 vdd.n2181 vdd.n1111 185
R16921 vdd.n2184 vdd.n2183 185
R16922 vdd.n2185 vdd.n1110 185
R16923 vdd.n2187 vdd.n2186 185
R16924 vdd.n2189 vdd.n1109 185
R16925 vdd.n2192 vdd.n2191 185
R16926 vdd.n2193 vdd.n1106 185
R16927 vdd.n2196 vdd.n2195 185
R16928 vdd.n2198 vdd.n1105 185
R16929 vdd.n2200 vdd.n2199 185
R16930 vdd.n2199 vdd.n1081 185
R16931 vdd.n315 vdd.n314 171.744
R16932 vdd.n314 vdd.n313 171.744
R16933 vdd.n313 vdd.n282 171.744
R16934 vdd.n306 vdd.n282 171.744
R16935 vdd.n306 vdd.n305 171.744
R16936 vdd.n305 vdd.n287 171.744
R16937 vdd.n298 vdd.n287 171.744
R16938 vdd.n298 vdd.n297 171.744
R16939 vdd.n297 vdd.n291 171.744
R16940 vdd.n260 vdd.n259 171.744
R16941 vdd.n259 vdd.n258 171.744
R16942 vdd.n258 vdd.n227 171.744
R16943 vdd.n251 vdd.n227 171.744
R16944 vdd.n251 vdd.n250 171.744
R16945 vdd.n250 vdd.n232 171.744
R16946 vdd.n243 vdd.n232 171.744
R16947 vdd.n243 vdd.n242 171.744
R16948 vdd.n242 vdd.n236 171.744
R16949 vdd.n217 vdd.n216 171.744
R16950 vdd.n216 vdd.n215 171.744
R16951 vdd.n215 vdd.n184 171.744
R16952 vdd.n208 vdd.n184 171.744
R16953 vdd.n208 vdd.n207 171.744
R16954 vdd.n207 vdd.n189 171.744
R16955 vdd.n200 vdd.n189 171.744
R16956 vdd.n200 vdd.n199 171.744
R16957 vdd.n199 vdd.n193 171.744
R16958 vdd.n162 vdd.n161 171.744
R16959 vdd.n161 vdd.n160 171.744
R16960 vdd.n160 vdd.n129 171.744
R16961 vdd.n153 vdd.n129 171.744
R16962 vdd.n153 vdd.n152 171.744
R16963 vdd.n152 vdd.n134 171.744
R16964 vdd.n145 vdd.n134 171.744
R16965 vdd.n145 vdd.n144 171.744
R16966 vdd.n144 vdd.n138 171.744
R16967 vdd.n120 vdd.n119 171.744
R16968 vdd.n119 vdd.n118 171.744
R16969 vdd.n118 vdd.n87 171.744
R16970 vdd.n111 vdd.n87 171.744
R16971 vdd.n111 vdd.n110 171.744
R16972 vdd.n110 vdd.n92 171.744
R16973 vdd.n103 vdd.n92 171.744
R16974 vdd.n103 vdd.n102 171.744
R16975 vdd.n102 vdd.n96 171.744
R16976 vdd.n65 vdd.n64 171.744
R16977 vdd.n64 vdd.n63 171.744
R16978 vdd.n63 vdd.n32 171.744
R16979 vdd.n56 vdd.n32 171.744
R16980 vdd.n56 vdd.n55 171.744
R16981 vdd.n55 vdd.n37 171.744
R16982 vdd.n48 vdd.n37 171.744
R16983 vdd.n48 vdd.n47 171.744
R16984 vdd.n47 vdd.n41 171.744
R16985 vdd.n1764 vdd.n1763 171.744
R16986 vdd.n1763 vdd.n1762 171.744
R16987 vdd.n1762 vdd.n1731 171.744
R16988 vdd.n1755 vdd.n1731 171.744
R16989 vdd.n1755 vdd.n1754 171.744
R16990 vdd.n1754 vdd.n1736 171.744
R16991 vdd.n1747 vdd.n1736 171.744
R16992 vdd.n1747 vdd.n1746 171.744
R16993 vdd.n1746 vdd.n1740 171.744
R16994 vdd.n1819 vdd.n1818 171.744
R16995 vdd.n1818 vdd.n1817 171.744
R16996 vdd.n1817 vdd.n1786 171.744
R16997 vdd.n1810 vdd.n1786 171.744
R16998 vdd.n1810 vdd.n1809 171.744
R16999 vdd.n1809 vdd.n1791 171.744
R17000 vdd.n1802 vdd.n1791 171.744
R17001 vdd.n1802 vdd.n1801 171.744
R17002 vdd.n1801 vdd.n1795 171.744
R17003 vdd.n1666 vdd.n1665 171.744
R17004 vdd.n1665 vdd.n1664 171.744
R17005 vdd.n1664 vdd.n1633 171.744
R17006 vdd.n1657 vdd.n1633 171.744
R17007 vdd.n1657 vdd.n1656 171.744
R17008 vdd.n1656 vdd.n1638 171.744
R17009 vdd.n1649 vdd.n1638 171.744
R17010 vdd.n1649 vdd.n1648 171.744
R17011 vdd.n1648 vdd.n1642 171.744
R17012 vdd.n1721 vdd.n1720 171.744
R17013 vdd.n1720 vdd.n1719 171.744
R17014 vdd.n1719 vdd.n1688 171.744
R17015 vdd.n1712 vdd.n1688 171.744
R17016 vdd.n1712 vdd.n1711 171.744
R17017 vdd.n1711 vdd.n1693 171.744
R17018 vdd.n1704 vdd.n1693 171.744
R17019 vdd.n1704 vdd.n1703 171.744
R17020 vdd.n1703 vdd.n1697 171.744
R17021 vdd.n1569 vdd.n1568 171.744
R17022 vdd.n1568 vdd.n1567 171.744
R17023 vdd.n1567 vdd.n1536 171.744
R17024 vdd.n1560 vdd.n1536 171.744
R17025 vdd.n1560 vdd.n1559 171.744
R17026 vdd.n1559 vdd.n1541 171.744
R17027 vdd.n1552 vdd.n1541 171.744
R17028 vdd.n1552 vdd.n1551 171.744
R17029 vdd.n1551 vdd.n1545 171.744
R17030 vdd.n1624 vdd.n1623 171.744
R17031 vdd.n1623 vdd.n1622 171.744
R17032 vdd.n1622 vdd.n1591 171.744
R17033 vdd.n1615 vdd.n1591 171.744
R17034 vdd.n1615 vdd.n1614 171.744
R17035 vdd.n1614 vdd.n1596 171.744
R17036 vdd.n1607 vdd.n1596 171.744
R17037 vdd.n1607 vdd.n1606 171.744
R17038 vdd.n1606 vdd.n1600 171.744
R17039 vdd.n449 vdd.n448 146.341
R17040 vdd.n455 vdd.n454 146.341
R17041 vdd.n459 vdd.n458 146.341
R17042 vdd.n465 vdd.n464 146.341
R17043 vdd.n469 vdd.n468 146.341
R17044 vdd.n475 vdd.n474 146.341
R17045 vdd.n479 vdd.n478 146.341
R17046 vdd.n485 vdd.n484 146.341
R17047 vdd.n489 vdd.n488 146.341
R17048 vdd.n495 vdd.n494 146.341
R17049 vdd.n499 vdd.n498 146.341
R17050 vdd.n505 vdd.n504 146.341
R17051 vdd.n509 vdd.n508 146.341
R17052 vdd.n515 vdd.n514 146.341
R17053 vdd.n519 vdd.n518 146.341
R17054 vdd.n525 vdd.n524 146.341
R17055 vdd.n529 vdd.n528 146.341
R17056 vdd.n535 vdd.n534 146.341
R17057 vdd.n539 vdd.n538 146.341
R17058 vdd.n545 vdd.n544 146.341
R17059 vdd.n549 vdd.n548 146.341
R17060 vdd.n555 vdd.n554 146.341
R17061 vdd.n559 vdd.n558 146.341
R17062 vdd.n565 vdd.n564 146.341
R17063 vdd.n569 vdd.n568 146.341
R17064 vdd.n575 vdd.n574 146.341
R17065 vdd.n579 vdd.n578 146.341
R17066 vdd.n585 vdd.n584 146.341
R17067 vdd.n589 vdd.n588 146.341
R17068 vdd.n595 vdd.n594 146.341
R17069 vdd.n597 vdd.n404 146.341
R17070 vdd.n3328 vdd.n654 146.341
R17071 vdd.n3334 vdd.n654 146.341
R17072 vdd.n3334 vdd.n647 146.341
R17073 vdd.n3344 vdd.n647 146.341
R17074 vdd.n3344 vdd.n643 146.341
R17075 vdd.n3350 vdd.n643 146.341
R17076 vdd.n3350 vdd.n634 146.341
R17077 vdd.n3360 vdd.n634 146.341
R17078 vdd.n3360 vdd.n630 146.341
R17079 vdd.n3366 vdd.n630 146.341
R17080 vdd.n3366 vdd.n623 146.341
R17081 vdd.n3377 vdd.n623 146.341
R17082 vdd.n3377 vdd.n619 146.341
R17083 vdd.n3386 vdd.n619 146.341
R17084 vdd.n3386 vdd.n612 146.341
R17085 vdd.n3396 vdd.n612 146.341
R17086 vdd.n3397 vdd.n3396 146.341
R17087 vdd.n3397 vdd.n329 146.341
R17088 vdd.n330 vdd.n329 146.341
R17089 vdd.n331 vdd.n330 146.341
R17090 vdd.n3404 vdd.n331 146.341
R17091 vdd.n3404 vdd.n339 146.341
R17092 vdd.n340 vdd.n339 146.341
R17093 vdd.n341 vdd.n340 146.341
R17094 vdd.n3411 vdd.n341 146.341
R17095 vdd.n3411 vdd.n350 146.341
R17096 vdd.n351 vdd.n350 146.341
R17097 vdd.n352 vdd.n351 146.341
R17098 vdd.n3419 vdd.n352 146.341
R17099 vdd.n3419 vdd.n360 146.341
R17100 vdd.n361 vdd.n360 146.341
R17101 vdd.n362 vdd.n361 146.341
R17102 vdd.n3426 vdd.n362 146.341
R17103 vdd.n3426 vdd.n371 146.341
R17104 vdd.n372 vdd.n371 146.341
R17105 vdd.n3320 vdd.n3318 146.341
R17106 vdd.n3318 vdd.n3317 146.341
R17107 vdd.n3314 vdd.n3313 146.341
R17108 vdd.n3310 vdd.n3309 146.341
R17109 vdd.n3307 vdd.n669 146.341
R17110 vdd.n3303 vdd.n3301 146.341
R17111 vdd.n3299 vdd.n675 146.341
R17112 vdd.n3295 vdd.n3293 146.341
R17113 vdd.n3291 vdd.n681 146.341
R17114 vdd.n3287 vdd.n3285 146.341
R17115 vdd.n3283 vdd.n689 146.341
R17116 vdd.n3279 vdd.n3277 146.341
R17117 vdd.n3275 vdd.n695 146.341
R17118 vdd.n3271 vdd.n3269 146.341
R17119 vdd.n3267 vdd.n701 146.341
R17120 vdd.n3263 vdd.n3261 146.341
R17121 vdd.n3259 vdd.n707 146.341
R17122 vdd.n3255 vdd.n3253 146.341
R17123 vdd.n3251 vdd.n713 146.341
R17124 vdd.n3247 vdd.n3245 146.341
R17125 vdd.n3243 vdd.n719 146.341
R17126 vdd.n3236 vdd.n728 146.341
R17127 vdd.n3234 vdd.n3233 146.341
R17128 vdd.n3230 vdd.n3229 146.341
R17129 vdd.n3227 vdd.n733 146.341
R17130 vdd.n3223 vdd.n3221 146.341
R17131 vdd.n3219 vdd.n739 146.341
R17132 vdd.n3215 vdd.n3213 146.341
R17133 vdd.n3211 vdd.n745 146.341
R17134 vdd.n3207 vdd.n3205 146.341
R17135 vdd.n3202 vdd.n3201 146.341
R17136 vdd.n3198 vdd.n657 146.341
R17137 vdd.n3326 vdd.n653 146.341
R17138 vdd.n3336 vdd.n653 146.341
R17139 vdd.n3336 vdd.n649 146.341
R17140 vdd.n3342 vdd.n649 146.341
R17141 vdd.n3342 vdd.n641 146.341
R17142 vdd.n3352 vdd.n641 146.341
R17143 vdd.n3352 vdd.n637 146.341
R17144 vdd.n3358 vdd.n637 146.341
R17145 vdd.n3358 vdd.n629 146.341
R17146 vdd.n3369 vdd.n629 146.341
R17147 vdd.n3369 vdd.n625 146.341
R17148 vdd.n3375 vdd.n625 146.341
R17149 vdd.n3375 vdd.n618 146.341
R17150 vdd.n3388 vdd.n618 146.341
R17151 vdd.n3388 vdd.n614 146.341
R17152 vdd.n3394 vdd.n614 146.341
R17153 vdd.n3394 vdd.n326 146.341
R17154 vdd.n3470 vdd.n326 146.341
R17155 vdd.n3470 vdd.n327 146.341
R17156 vdd.n3466 vdd.n327 146.341
R17157 vdd.n3466 vdd.n333 146.341
R17158 vdd.n3462 vdd.n333 146.341
R17159 vdd.n3462 vdd.n338 146.341
R17160 vdd.n3458 vdd.n338 146.341
R17161 vdd.n3458 vdd.n342 146.341
R17162 vdd.n3454 vdd.n342 146.341
R17163 vdd.n3454 vdd.n348 146.341
R17164 vdd.n3450 vdd.n348 146.341
R17165 vdd.n3450 vdd.n353 146.341
R17166 vdd.n3446 vdd.n353 146.341
R17167 vdd.n3446 vdd.n359 146.341
R17168 vdd.n3442 vdd.n359 146.341
R17169 vdd.n3442 vdd.n364 146.341
R17170 vdd.n3438 vdd.n364 146.341
R17171 vdd.n3438 vdd.n370 146.341
R17172 vdd.n2106 vdd.n2105 146.341
R17173 vdd.n2103 vdd.n1900 146.341
R17174 vdd.n2096 vdd.n1906 146.341
R17175 vdd.n2094 vdd.n2093 146.341
R17176 vdd.n2091 vdd.n1908 146.341
R17177 vdd.n2087 vdd.n2086 146.341
R17178 vdd.n2084 vdd.n1915 146.341
R17179 vdd.n2080 vdd.n2079 146.341
R17180 vdd.n2077 vdd.n1922 146.341
R17181 vdd.n1933 vdd.n1930 146.341
R17182 vdd.n2069 vdd.n2068 146.341
R17183 vdd.n2066 vdd.n1935 146.341
R17184 vdd.n2062 vdd.n2061 146.341
R17185 vdd.n2059 vdd.n1941 146.341
R17186 vdd.n2055 vdd.n2054 146.341
R17187 vdd.n2052 vdd.n1948 146.341
R17188 vdd.n2048 vdd.n2047 146.341
R17189 vdd.n2045 vdd.n1955 146.341
R17190 vdd.n2041 vdd.n2040 146.341
R17191 vdd.n2038 vdd.n1962 146.341
R17192 vdd.n1973 vdd.n1970 146.341
R17193 vdd.n2030 vdd.n2029 146.341
R17194 vdd.n2027 vdd.n1975 146.341
R17195 vdd.n2023 vdd.n2022 146.341
R17196 vdd.n2020 vdd.n1981 146.341
R17197 vdd.n2016 vdd.n2015 146.341
R17198 vdd.n2013 vdd.n1988 146.341
R17199 vdd.n2009 vdd.n2008 146.341
R17200 vdd.n2006 vdd.n2003 146.341
R17201 vdd.n2001 vdd.n1998 146.341
R17202 vdd.n1996 vdd.n1120 146.341
R17203 vdd.n1461 vdd.n1225 146.341
R17204 vdd.n1461 vdd.n1217 146.341
R17205 vdd.n1471 vdd.n1217 146.341
R17206 vdd.n1471 vdd.n1213 146.341
R17207 vdd.n1477 vdd.n1213 146.341
R17208 vdd.n1477 vdd.n1205 146.341
R17209 vdd.n1488 vdd.n1205 146.341
R17210 vdd.n1488 vdd.n1201 146.341
R17211 vdd.n1494 vdd.n1201 146.341
R17212 vdd.n1494 vdd.n1195 146.341
R17213 vdd.n1505 vdd.n1195 146.341
R17214 vdd.n1505 vdd.n1191 146.341
R17215 vdd.n1511 vdd.n1191 146.341
R17216 vdd.n1511 vdd.n1182 146.341
R17217 vdd.n1521 vdd.n1182 146.341
R17218 vdd.n1521 vdd.n1178 146.341
R17219 vdd.n1527 vdd.n1178 146.341
R17220 vdd.n1527 vdd.n1171 146.341
R17221 vdd.n1833 vdd.n1171 146.341
R17222 vdd.n1833 vdd.n1167 146.341
R17223 vdd.n1839 vdd.n1167 146.341
R17224 vdd.n1839 vdd.n1160 146.341
R17225 vdd.n1849 vdd.n1160 146.341
R17226 vdd.n1849 vdd.n1156 146.341
R17227 vdd.n1855 vdd.n1156 146.341
R17228 vdd.n1855 vdd.n1148 146.341
R17229 vdd.n1866 vdd.n1148 146.341
R17230 vdd.n1866 vdd.n1144 146.341
R17231 vdd.n1872 vdd.n1144 146.341
R17232 vdd.n1872 vdd.n1138 146.341
R17233 vdd.n1883 vdd.n1138 146.341
R17234 vdd.n1883 vdd.n1133 146.341
R17235 vdd.n1891 vdd.n1133 146.341
R17236 vdd.n1891 vdd.n1122 146.341
R17237 vdd.n2114 vdd.n1122 146.341
R17238 vdd.n1263 vdd.n1262 146.341
R17239 vdd.n1267 vdd.n1262 146.341
R17240 vdd.n1269 vdd.n1268 146.341
R17241 vdd.n1273 vdd.n1272 146.341
R17242 vdd.n1275 vdd.n1274 146.341
R17243 vdd.n1279 vdd.n1278 146.341
R17244 vdd.n1281 vdd.n1280 146.341
R17245 vdd.n1285 vdd.n1284 146.341
R17246 vdd.n1287 vdd.n1286 146.341
R17247 vdd.n1419 vdd.n1418 146.341
R17248 vdd.n1291 vdd.n1290 146.341
R17249 vdd.n1295 vdd.n1294 146.341
R17250 vdd.n1297 vdd.n1296 146.341
R17251 vdd.n1301 vdd.n1300 146.341
R17252 vdd.n1303 vdd.n1302 146.341
R17253 vdd.n1307 vdd.n1306 146.341
R17254 vdd.n1309 vdd.n1308 146.341
R17255 vdd.n1313 vdd.n1312 146.341
R17256 vdd.n1315 vdd.n1314 146.341
R17257 vdd.n1319 vdd.n1318 146.341
R17258 vdd.n1383 vdd.n1320 146.341
R17259 vdd.n1324 vdd.n1323 146.341
R17260 vdd.n1326 vdd.n1325 146.341
R17261 vdd.n1330 vdd.n1329 146.341
R17262 vdd.n1332 vdd.n1331 146.341
R17263 vdd.n1336 vdd.n1335 146.341
R17264 vdd.n1338 vdd.n1337 146.341
R17265 vdd.n1342 vdd.n1341 146.341
R17266 vdd.n1344 vdd.n1343 146.341
R17267 vdd.n1348 vdd.n1347 146.341
R17268 vdd.n1350 vdd.n1349 146.341
R17269 vdd.n1455 vdd.n1231 146.341
R17270 vdd.n1463 vdd.n1223 146.341
R17271 vdd.n1463 vdd.n1219 146.341
R17272 vdd.n1469 vdd.n1219 146.341
R17273 vdd.n1469 vdd.n1211 146.341
R17274 vdd.n1480 vdd.n1211 146.341
R17275 vdd.n1480 vdd.n1207 146.341
R17276 vdd.n1486 vdd.n1207 146.341
R17277 vdd.n1486 vdd.n1200 146.341
R17278 vdd.n1497 vdd.n1200 146.341
R17279 vdd.n1497 vdd.n1196 146.341
R17280 vdd.n1503 vdd.n1196 146.341
R17281 vdd.n1503 vdd.n1189 146.341
R17282 vdd.n1513 vdd.n1189 146.341
R17283 vdd.n1513 vdd.n1185 146.341
R17284 vdd.n1519 vdd.n1185 146.341
R17285 vdd.n1519 vdd.n1177 146.341
R17286 vdd.n1530 vdd.n1177 146.341
R17287 vdd.n1530 vdd.n1173 146.341
R17288 vdd.n1831 vdd.n1173 146.341
R17289 vdd.n1831 vdd.n1166 146.341
R17290 vdd.n1841 vdd.n1166 146.341
R17291 vdd.n1841 vdd.n1162 146.341
R17292 vdd.n1847 vdd.n1162 146.341
R17293 vdd.n1847 vdd.n1154 146.341
R17294 vdd.n1858 vdd.n1154 146.341
R17295 vdd.n1858 vdd.n1150 146.341
R17296 vdd.n1864 vdd.n1150 146.341
R17297 vdd.n1864 vdd.n1143 146.341
R17298 vdd.n1875 vdd.n1143 146.341
R17299 vdd.n1875 vdd.n1139 146.341
R17300 vdd.n1881 vdd.n1139 146.341
R17301 vdd.n1881 vdd.n1131 146.341
R17302 vdd.n1893 vdd.n1131 146.341
R17303 vdd.n1893 vdd.n1126 146.341
R17304 vdd.n2112 vdd.n1126 146.341
R17305 vdd.n1107 vdd.t155 127.284
R17306 vdd.n968 vdd.t192 127.284
R17307 vdd.n1101 vdd.t219 127.284
R17308 vdd.n959 vdd.t215 127.284
R17309 vdd.n856 vdd.t165 127.284
R17310 vdd.n856 vdd.t166 127.284
R17311 vdd.n2678 vdd.t210 127.284
R17312 vdd.n804 vdd.t185 127.284
R17313 vdd.n2747 vdd.t197 127.284
R17314 vdd.n768 vdd.t150 127.284
R17315 vdd.n1029 vdd.t206 127.284
R17316 vdd.n1029 vdd.t207 127.284
R17317 vdd.n22 vdd.n20 117.314
R17318 vdd.n17 vdd.n15 117.314
R17319 vdd.n27 vdd.n26 116.927
R17320 vdd.n24 vdd.n23 116.927
R17321 vdd.n22 vdd.n21 116.927
R17322 vdd.n17 vdd.n16 116.927
R17323 vdd.n19 vdd.n18 116.927
R17324 vdd.n27 vdd.n25 116.927
R17325 vdd.n1108 vdd.t154 111.188
R17326 vdd.n969 vdd.t193 111.188
R17327 vdd.n1102 vdd.t218 111.188
R17328 vdd.n960 vdd.t216 111.188
R17329 vdd.n2679 vdd.t209 111.188
R17330 vdd.n805 vdd.t186 111.188
R17331 vdd.n2748 vdd.t196 111.188
R17332 vdd.n769 vdd.t151 111.188
R17333 vdd.n2933 vdd.n909 99.5127
R17334 vdd.n2941 vdd.n909 99.5127
R17335 vdd.n2941 vdd.n907 99.5127
R17336 vdd.n2945 vdd.n907 99.5127
R17337 vdd.n2945 vdd.n897 99.5127
R17338 vdd.n2953 vdd.n897 99.5127
R17339 vdd.n2953 vdd.n895 99.5127
R17340 vdd.n2957 vdd.n895 99.5127
R17341 vdd.n2957 vdd.n887 99.5127
R17342 vdd.n2965 vdd.n887 99.5127
R17343 vdd.n2965 vdd.n885 99.5127
R17344 vdd.n2969 vdd.n885 99.5127
R17345 vdd.n2969 vdd.n875 99.5127
R17346 vdd.n2977 vdd.n875 99.5127
R17347 vdd.n2977 vdd.n873 99.5127
R17348 vdd.n2981 vdd.n873 99.5127
R17349 vdd.n2981 vdd.n864 99.5127
R17350 vdd.n2989 vdd.n864 99.5127
R17351 vdd.n2989 vdd.n862 99.5127
R17352 vdd.n2993 vdd.n862 99.5127
R17353 vdd.n2993 vdd.n851 99.5127
R17354 vdd.n3002 vdd.n851 99.5127
R17355 vdd.n3002 vdd.n849 99.5127
R17356 vdd.n3006 vdd.n849 99.5127
R17357 vdd.n3006 vdd.n838 99.5127
R17358 vdd.n3014 vdd.n838 99.5127
R17359 vdd.n3014 vdd.n836 99.5127
R17360 vdd.n3018 vdd.n836 99.5127
R17361 vdd.n3018 vdd.n827 99.5127
R17362 vdd.n3026 vdd.n827 99.5127
R17363 vdd.n3026 vdd.n825 99.5127
R17364 vdd.n3030 vdd.n825 99.5127
R17365 vdd.n3030 vdd.n813 99.5127
R17366 vdd.n3083 vdd.n813 99.5127
R17367 vdd.n3083 vdd.n811 99.5127
R17368 vdd.n3087 vdd.n811 99.5127
R17369 vdd.n3087 vdd.n777 99.5127
R17370 vdd.n3157 vdd.n777 99.5127
R17371 vdd.n3153 vdd.n778 99.5127
R17372 vdd.n3151 vdd.n3150 99.5127
R17373 vdd.n3148 vdd.n782 99.5127
R17374 vdd.n3144 vdd.n3143 99.5127
R17375 vdd.n3141 vdd.n785 99.5127
R17376 vdd.n3137 vdd.n3136 99.5127
R17377 vdd.n3134 vdd.n788 99.5127
R17378 vdd.n3130 vdd.n3129 99.5127
R17379 vdd.n3127 vdd.n791 99.5127
R17380 vdd.n3122 vdd.n3121 99.5127
R17381 vdd.n3119 vdd.n794 99.5127
R17382 vdd.n3115 vdd.n3114 99.5127
R17383 vdd.n3112 vdd.n797 99.5127
R17384 vdd.n3108 vdd.n3107 99.5127
R17385 vdd.n3105 vdd.n800 99.5127
R17386 vdd.n3101 vdd.n3100 99.5127
R17387 vdd.n3098 vdd.n803 99.5127
R17388 vdd.n2815 vdd.n915 99.5127
R17389 vdd.n2815 vdd.n910 99.5127
R17390 vdd.n2917 vdd.n910 99.5127
R17391 vdd.n2917 vdd.n905 99.5127
R17392 vdd.n2913 vdd.n905 99.5127
R17393 vdd.n2913 vdd.n899 99.5127
R17394 vdd.n2910 vdd.n899 99.5127
R17395 vdd.n2910 vdd.n893 99.5127
R17396 vdd.n2907 vdd.n893 99.5127
R17397 vdd.n2907 vdd.n888 99.5127
R17398 vdd.n2857 vdd.n888 99.5127
R17399 vdd.n2857 vdd.n883 99.5127
R17400 vdd.n2860 vdd.n883 99.5127
R17401 vdd.n2860 vdd.n877 99.5127
R17402 vdd.n2893 vdd.n877 99.5127
R17403 vdd.n2893 vdd.n870 99.5127
R17404 vdd.n2889 vdd.n870 99.5127
R17405 vdd.n2889 vdd.n865 99.5127
R17406 vdd.n2886 vdd.n865 99.5127
R17407 vdd.n2886 vdd.n860 99.5127
R17408 vdd.n2883 vdd.n860 99.5127
R17409 vdd.n2883 vdd.n853 99.5127
R17410 vdd.n2880 vdd.n853 99.5127
R17411 vdd.n2880 vdd.n846 99.5127
R17412 vdd.n2877 vdd.n846 99.5127
R17413 vdd.n2877 vdd.n839 99.5127
R17414 vdd.n2874 vdd.n839 99.5127
R17415 vdd.n2874 vdd.n833 99.5127
R17416 vdd.n2871 vdd.n833 99.5127
R17417 vdd.n2871 vdd.n828 99.5127
R17418 vdd.n2868 vdd.n828 99.5127
R17419 vdd.n2868 vdd.n823 99.5127
R17420 vdd.n2865 vdd.n823 99.5127
R17421 vdd.n2865 vdd.n815 99.5127
R17422 vdd.n815 vdd.n808 99.5127
R17423 vdd.n3089 vdd.n808 99.5127
R17424 vdd.n3090 vdd.n3089 99.5127
R17425 vdd.n3090 vdd.n775 99.5127
R17426 vdd.n2929 vdd.n920 99.5127
R17427 vdd.n2749 vdd.n920 99.5127
R17428 vdd.n2753 vdd.n2752 99.5127
R17429 vdd.n2757 vdd.n2756 99.5127
R17430 vdd.n2761 vdd.n2760 99.5127
R17431 vdd.n2765 vdd.n2764 99.5127
R17432 vdd.n2769 vdd.n2768 99.5127
R17433 vdd.n2773 vdd.n2772 99.5127
R17434 vdd.n2777 vdd.n2776 99.5127
R17435 vdd.n2781 vdd.n2780 99.5127
R17436 vdd.n2785 vdd.n2784 99.5127
R17437 vdd.n2789 vdd.n2788 99.5127
R17438 vdd.n2793 vdd.n2792 99.5127
R17439 vdd.n2797 vdd.n2796 99.5127
R17440 vdd.n2801 vdd.n2800 99.5127
R17441 vdd.n2805 vdd.n2804 99.5127
R17442 vdd.n2810 vdd.n2809 99.5127
R17443 vdd.n2642 vdd.n957 99.5127
R17444 vdd.n2638 vdd.n2637 99.5127
R17445 vdd.n2634 vdd.n2633 99.5127
R17446 vdd.n2630 vdd.n2629 99.5127
R17447 vdd.n2626 vdd.n2625 99.5127
R17448 vdd.n2622 vdd.n2621 99.5127
R17449 vdd.n2618 vdd.n2617 99.5127
R17450 vdd.n2614 vdd.n2613 99.5127
R17451 vdd.n2610 vdd.n2609 99.5127
R17452 vdd.n2606 vdd.n2605 99.5127
R17453 vdd.n2602 vdd.n2601 99.5127
R17454 vdd.n2598 vdd.n2597 99.5127
R17455 vdd.n2594 vdd.n2593 99.5127
R17456 vdd.n2590 vdd.n2589 99.5127
R17457 vdd.n2586 vdd.n2585 99.5127
R17458 vdd.n2582 vdd.n2581 99.5127
R17459 vdd.n2577 vdd.n2576 99.5127
R17460 vdd.n2309 vdd.n1082 99.5127
R17461 vdd.n2309 vdd.n1076 99.5127
R17462 vdd.n2306 vdd.n1076 99.5127
R17463 vdd.n2306 vdd.n1070 99.5127
R17464 vdd.n2303 vdd.n1070 99.5127
R17465 vdd.n2303 vdd.n1064 99.5127
R17466 vdd.n2300 vdd.n1064 99.5127
R17467 vdd.n2300 vdd.n1058 99.5127
R17468 vdd.n2297 vdd.n1058 99.5127
R17469 vdd.n2297 vdd.n1052 99.5127
R17470 vdd.n2294 vdd.n1052 99.5127
R17471 vdd.n2294 vdd.n1046 99.5127
R17472 vdd.n2291 vdd.n1046 99.5127
R17473 vdd.n2291 vdd.n1039 99.5127
R17474 vdd.n2288 vdd.n1039 99.5127
R17475 vdd.n2288 vdd.n1032 99.5127
R17476 vdd.n2285 vdd.n1032 99.5127
R17477 vdd.n2285 vdd.n1026 99.5127
R17478 vdd.n2282 vdd.n1026 99.5127
R17479 vdd.n2282 vdd.n1021 99.5127
R17480 vdd.n2279 vdd.n1021 99.5127
R17481 vdd.n2279 vdd.n1015 99.5127
R17482 vdd.n2276 vdd.n1015 99.5127
R17483 vdd.n2276 vdd.n1008 99.5127
R17484 vdd.n2243 vdd.n1008 99.5127
R17485 vdd.n2243 vdd.n1002 99.5127
R17486 vdd.n2246 vdd.n1002 99.5127
R17487 vdd.n2246 vdd.n997 99.5127
R17488 vdd.n2262 vdd.n997 99.5127
R17489 vdd.n2262 vdd.n992 99.5127
R17490 vdd.n2258 vdd.n992 99.5127
R17491 vdd.n2258 vdd.n987 99.5127
R17492 vdd.n2255 vdd.n987 99.5127
R17493 vdd.n2255 vdd.n980 99.5127
R17494 vdd.n2252 vdd.n980 99.5127
R17495 vdd.n2252 vdd.n973 99.5127
R17496 vdd.n973 vdd.n962 99.5127
R17497 vdd.n2572 vdd.n962 99.5127
R17498 vdd.n2379 vdd.n2377 99.5127
R17499 vdd.n2377 vdd.n2376 99.5127
R17500 vdd.n2373 vdd.n2372 99.5127
R17501 vdd.n2370 vdd.n1088 99.5127
R17502 vdd.n2366 vdd.n2364 99.5127
R17503 vdd.n2362 vdd.n1090 99.5127
R17504 vdd.n2358 vdd.n2356 99.5127
R17505 vdd.n2354 vdd.n1092 99.5127
R17506 vdd.n2350 vdd.n2348 99.5127
R17507 vdd.n2346 vdd.n1094 99.5127
R17508 vdd.n2342 vdd.n2340 99.5127
R17509 vdd.n2338 vdd.n1096 99.5127
R17510 vdd.n2334 vdd.n2332 99.5127
R17511 vdd.n2330 vdd.n1098 99.5127
R17512 vdd.n2326 vdd.n2324 99.5127
R17513 vdd.n2322 vdd.n1100 99.5127
R17514 vdd.n2317 vdd.n2315 99.5127
R17515 vdd.n2383 vdd.n1074 99.5127
R17516 vdd.n2391 vdd.n1074 99.5127
R17517 vdd.n2391 vdd.n1072 99.5127
R17518 vdd.n2395 vdd.n1072 99.5127
R17519 vdd.n2395 vdd.n1062 99.5127
R17520 vdd.n2403 vdd.n1062 99.5127
R17521 vdd.n2403 vdd.n1060 99.5127
R17522 vdd.n2407 vdd.n1060 99.5127
R17523 vdd.n2407 vdd.n1050 99.5127
R17524 vdd.n2415 vdd.n1050 99.5127
R17525 vdd.n2415 vdd.n1048 99.5127
R17526 vdd.n2419 vdd.n1048 99.5127
R17527 vdd.n2419 vdd.n1037 99.5127
R17528 vdd.n2427 vdd.n1037 99.5127
R17529 vdd.n2427 vdd.n1035 99.5127
R17530 vdd.n2431 vdd.n1035 99.5127
R17531 vdd.n2431 vdd.n1025 99.5127
R17532 vdd.n2440 vdd.n1025 99.5127
R17533 vdd.n2440 vdd.n1023 99.5127
R17534 vdd.n2444 vdd.n1023 99.5127
R17535 vdd.n2444 vdd.n1013 99.5127
R17536 vdd.n2452 vdd.n1013 99.5127
R17537 vdd.n2452 vdd.n1011 99.5127
R17538 vdd.n2456 vdd.n1011 99.5127
R17539 vdd.n2456 vdd.n1001 99.5127
R17540 vdd.n2464 vdd.n1001 99.5127
R17541 vdd.n2464 vdd.n999 99.5127
R17542 vdd.n2468 vdd.n999 99.5127
R17543 vdd.n2468 vdd.n991 99.5127
R17544 vdd.n2476 vdd.n991 99.5127
R17545 vdd.n2476 vdd.n989 99.5127
R17546 vdd.n2480 vdd.n989 99.5127
R17547 vdd.n2480 vdd.n978 99.5127
R17548 vdd.n2490 vdd.n978 99.5127
R17549 vdd.n2490 vdd.n975 99.5127
R17550 vdd.n2495 vdd.n975 99.5127
R17551 vdd.n2495 vdd.n976 99.5127
R17552 vdd.n976 vdd.n956 99.5127
R17553 vdd.n3073 vdd.n3072 99.5127
R17554 vdd.n3070 vdd.n3036 99.5127
R17555 vdd.n3066 vdd.n3065 99.5127
R17556 vdd.n3063 vdd.n3039 99.5127
R17557 vdd.n3059 vdd.n3058 99.5127
R17558 vdd.n3056 vdd.n3042 99.5127
R17559 vdd.n3052 vdd.n3051 99.5127
R17560 vdd.n3049 vdd.n3046 99.5127
R17561 vdd.n3190 vdd.n755 99.5127
R17562 vdd.n3188 vdd.n3187 99.5127
R17563 vdd.n3185 vdd.n758 99.5127
R17564 vdd.n3181 vdd.n3180 99.5127
R17565 vdd.n3178 vdd.n761 99.5127
R17566 vdd.n3174 vdd.n3173 99.5127
R17567 vdd.n3171 vdd.n764 99.5127
R17568 vdd.n3167 vdd.n3166 99.5127
R17569 vdd.n3164 vdd.n767 99.5127
R17570 vdd.n2922 vdd.n916 99.5127
R17571 vdd.n2922 vdd.n911 99.5127
R17572 vdd.n2919 vdd.n911 99.5127
R17573 vdd.n2919 vdd.n906 99.5127
R17574 vdd.n2819 vdd.n906 99.5127
R17575 vdd.n2819 vdd.n900 99.5127
R17576 vdd.n2822 vdd.n900 99.5127
R17577 vdd.n2822 vdd.n894 99.5127
R17578 vdd.n2905 vdd.n894 99.5127
R17579 vdd.n2905 vdd.n889 99.5127
R17580 vdd.n2901 vdd.n889 99.5127
R17581 vdd.n2901 vdd.n884 99.5127
R17582 vdd.n2898 vdd.n884 99.5127
R17583 vdd.n2898 vdd.n878 99.5127
R17584 vdd.n2895 vdd.n878 99.5127
R17585 vdd.n2895 vdd.n871 99.5127
R17586 vdd.n2854 vdd.n871 99.5127
R17587 vdd.n2854 vdd.n866 99.5127
R17588 vdd.n2851 vdd.n866 99.5127
R17589 vdd.n2851 vdd.n861 99.5127
R17590 vdd.n2848 vdd.n861 99.5127
R17591 vdd.n2848 vdd.n854 99.5127
R17592 vdd.n2845 vdd.n854 99.5127
R17593 vdd.n2845 vdd.n847 99.5127
R17594 vdd.n2842 vdd.n847 99.5127
R17595 vdd.n2842 vdd.n840 99.5127
R17596 vdd.n2839 vdd.n840 99.5127
R17597 vdd.n2839 vdd.n834 99.5127
R17598 vdd.n2836 vdd.n834 99.5127
R17599 vdd.n2836 vdd.n829 99.5127
R17600 vdd.n2833 vdd.n829 99.5127
R17601 vdd.n2833 vdd.n824 99.5127
R17602 vdd.n2830 vdd.n824 99.5127
R17603 vdd.n2830 vdd.n816 99.5127
R17604 vdd.n2827 vdd.n816 99.5127
R17605 vdd.n2827 vdd.n809 99.5127
R17606 vdd.n809 vdd.n773 99.5127
R17607 vdd.n3159 vdd.n773 99.5127
R17608 vdd.n2683 vdd.n2682 99.5127
R17609 vdd.n2687 vdd.n2686 99.5127
R17610 vdd.n2691 vdd.n2690 99.5127
R17611 vdd.n2695 vdd.n2694 99.5127
R17612 vdd.n2699 vdd.n2698 99.5127
R17613 vdd.n2703 vdd.n2702 99.5127
R17614 vdd.n2707 vdd.n2706 99.5127
R17615 vdd.n2711 vdd.n2710 99.5127
R17616 vdd.n2715 vdd.n2714 99.5127
R17617 vdd.n2719 vdd.n2718 99.5127
R17618 vdd.n2723 vdd.n2722 99.5127
R17619 vdd.n2727 vdd.n2726 99.5127
R17620 vdd.n2731 vdd.n2730 99.5127
R17621 vdd.n2735 vdd.n2734 99.5127
R17622 vdd.n2739 vdd.n2738 99.5127
R17623 vdd.n2743 vdd.n2742 99.5127
R17624 vdd.n2926 vdd.n2677 99.5127
R17625 vdd.n2935 vdd.n912 99.5127
R17626 vdd.n2939 vdd.n912 99.5127
R17627 vdd.n2939 vdd.n904 99.5127
R17628 vdd.n2947 vdd.n904 99.5127
R17629 vdd.n2947 vdd.n902 99.5127
R17630 vdd.n2951 vdd.n902 99.5127
R17631 vdd.n2951 vdd.n892 99.5127
R17632 vdd.n2959 vdd.n892 99.5127
R17633 vdd.n2959 vdd.n890 99.5127
R17634 vdd.n2963 vdd.n890 99.5127
R17635 vdd.n2963 vdd.n881 99.5127
R17636 vdd.n2971 vdd.n881 99.5127
R17637 vdd.n2971 vdd.n879 99.5127
R17638 vdd.n2975 vdd.n879 99.5127
R17639 vdd.n2975 vdd.n869 99.5127
R17640 vdd.n2983 vdd.n869 99.5127
R17641 vdd.n2983 vdd.n867 99.5127
R17642 vdd.n2987 vdd.n867 99.5127
R17643 vdd.n2987 vdd.n858 99.5127
R17644 vdd.n2995 vdd.n858 99.5127
R17645 vdd.n2995 vdd.n855 99.5127
R17646 vdd.n3000 vdd.n855 99.5127
R17647 vdd.n3000 vdd.n844 99.5127
R17648 vdd.n3008 vdd.n844 99.5127
R17649 vdd.n3008 vdd.n842 99.5127
R17650 vdd.n3012 vdd.n842 99.5127
R17651 vdd.n3012 vdd.n832 99.5127
R17652 vdd.n3020 vdd.n832 99.5127
R17653 vdd.n3020 vdd.n830 99.5127
R17654 vdd.n3024 vdd.n830 99.5127
R17655 vdd.n3024 vdd.n821 99.5127
R17656 vdd.n3032 vdd.n821 99.5127
R17657 vdd.n3032 vdd.n818 99.5127
R17658 vdd.n3081 vdd.n818 99.5127
R17659 vdd.n3081 vdd.n819 99.5127
R17660 vdd.n819 vdd.n810 99.5127
R17661 vdd.n3076 vdd.n810 99.5127
R17662 vdd.n3076 vdd.n776 99.5127
R17663 vdd.n2566 vdd.n2565 99.5127
R17664 vdd.n2562 vdd.n2561 99.5127
R17665 vdd.n2558 vdd.n2557 99.5127
R17666 vdd.n2554 vdd.n2553 99.5127
R17667 vdd.n2550 vdd.n2549 99.5127
R17668 vdd.n2546 vdd.n2545 99.5127
R17669 vdd.n2542 vdd.n2541 99.5127
R17670 vdd.n2538 vdd.n2537 99.5127
R17671 vdd.n2534 vdd.n2533 99.5127
R17672 vdd.n2530 vdd.n2529 99.5127
R17673 vdd.n2526 vdd.n2525 99.5127
R17674 vdd.n2522 vdd.n2521 99.5127
R17675 vdd.n2518 vdd.n2517 99.5127
R17676 vdd.n2514 vdd.n2513 99.5127
R17677 vdd.n2510 vdd.n2509 99.5127
R17678 vdd.n2506 vdd.n2505 99.5127
R17679 vdd.n2502 vdd.n938 99.5127
R17680 vdd.n2202 vdd.n1083 99.5127
R17681 vdd.n2202 vdd.n1077 99.5127
R17682 vdd.n2205 vdd.n1077 99.5127
R17683 vdd.n2205 vdd.n1071 99.5127
R17684 vdd.n2208 vdd.n1071 99.5127
R17685 vdd.n2208 vdd.n1065 99.5127
R17686 vdd.n2211 vdd.n1065 99.5127
R17687 vdd.n2211 vdd.n1059 99.5127
R17688 vdd.n2214 vdd.n1059 99.5127
R17689 vdd.n2214 vdd.n1053 99.5127
R17690 vdd.n2217 vdd.n1053 99.5127
R17691 vdd.n2217 vdd.n1047 99.5127
R17692 vdd.n2220 vdd.n1047 99.5127
R17693 vdd.n2220 vdd.n1040 99.5127
R17694 vdd.n2223 vdd.n1040 99.5127
R17695 vdd.n2223 vdd.n1033 99.5127
R17696 vdd.n2226 vdd.n1033 99.5127
R17697 vdd.n2226 vdd.n1027 99.5127
R17698 vdd.n2229 vdd.n1027 99.5127
R17699 vdd.n2229 vdd.n1022 99.5127
R17700 vdd.n2232 vdd.n1022 99.5127
R17701 vdd.n2232 vdd.n1016 99.5127
R17702 vdd.n2274 vdd.n1016 99.5127
R17703 vdd.n2274 vdd.n1009 99.5127
R17704 vdd.n2270 vdd.n1009 99.5127
R17705 vdd.n2270 vdd.n1003 99.5127
R17706 vdd.n2267 vdd.n1003 99.5127
R17707 vdd.n2267 vdd.n998 99.5127
R17708 vdd.n2264 vdd.n998 99.5127
R17709 vdd.n2264 vdd.n993 99.5127
R17710 vdd.n2240 vdd.n993 99.5127
R17711 vdd.n2240 vdd.n988 99.5127
R17712 vdd.n2237 vdd.n988 99.5127
R17713 vdd.n2237 vdd.n981 99.5127
R17714 vdd.n981 vdd.n972 99.5127
R17715 vdd.n2497 vdd.n972 99.5127
R17716 vdd.n2498 vdd.n2497 99.5127
R17717 vdd.n2498 vdd.n964 99.5127
R17718 vdd.n2135 vdd.n2133 99.5127
R17719 vdd.n2139 vdd.n2130 99.5127
R17720 vdd.n2143 vdd.n2141 99.5127
R17721 vdd.n2147 vdd.n2128 99.5127
R17722 vdd.n2151 vdd.n2149 99.5127
R17723 vdd.n2155 vdd.n2126 99.5127
R17724 vdd.n2159 vdd.n2157 99.5127
R17725 vdd.n2163 vdd.n2124 99.5127
R17726 vdd.n2167 vdd.n2165 99.5127
R17727 vdd.n2171 vdd.n1114 99.5127
R17728 vdd.n2175 vdd.n2173 99.5127
R17729 vdd.n2179 vdd.n1112 99.5127
R17730 vdd.n2183 vdd.n2181 99.5127
R17731 vdd.n2187 vdd.n1110 99.5127
R17732 vdd.n2191 vdd.n2189 99.5127
R17733 vdd.n2196 vdd.n1106 99.5127
R17734 vdd.n2199 vdd.n2198 99.5127
R17735 vdd.n2385 vdd.n1078 99.5127
R17736 vdd.n2389 vdd.n1078 99.5127
R17737 vdd.n2389 vdd.n1068 99.5127
R17738 vdd.n2397 vdd.n1068 99.5127
R17739 vdd.n2397 vdd.n1066 99.5127
R17740 vdd.n2401 vdd.n1066 99.5127
R17741 vdd.n2401 vdd.n1056 99.5127
R17742 vdd.n2409 vdd.n1056 99.5127
R17743 vdd.n2409 vdd.n1054 99.5127
R17744 vdd.n2413 vdd.n1054 99.5127
R17745 vdd.n2413 vdd.n1044 99.5127
R17746 vdd.n2421 vdd.n1044 99.5127
R17747 vdd.n2421 vdd.n1042 99.5127
R17748 vdd.n2425 vdd.n1042 99.5127
R17749 vdd.n2425 vdd.n1031 99.5127
R17750 vdd.n2433 vdd.n1031 99.5127
R17751 vdd.n2433 vdd.n1028 99.5127
R17752 vdd.n2438 vdd.n1028 99.5127
R17753 vdd.n2438 vdd.n1019 99.5127
R17754 vdd.n2446 vdd.n1019 99.5127
R17755 vdd.n2446 vdd.n1017 99.5127
R17756 vdd.n2450 vdd.n1017 99.5127
R17757 vdd.n2450 vdd.n1007 99.5127
R17758 vdd.n2458 vdd.n1007 99.5127
R17759 vdd.n2458 vdd.n1005 99.5127
R17760 vdd.n2462 vdd.n1005 99.5127
R17761 vdd.n2462 vdd.n996 99.5127
R17762 vdd.n2470 vdd.n996 99.5127
R17763 vdd.n2470 vdd.n994 99.5127
R17764 vdd.n2474 vdd.n994 99.5127
R17765 vdd.n2474 vdd.n985 99.5127
R17766 vdd.n2482 vdd.n985 99.5127
R17767 vdd.n2482 vdd.n982 99.5127
R17768 vdd.n2488 vdd.n982 99.5127
R17769 vdd.n2488 vdd.n983 99.5127
R17770 vdd.n983 vdd.n974 99.5127
R17771 vdd.n974 vdd.n965 99.5127
R17772 vdd.n2570 vdd.n965 99.5127
R17773 vdd.n9 vdd.n7 98.9633
R17774 vdd.n2 vdd.n0 98.9633
R17775 vdd.n9 vdd.n8 98.6055
R17776 vdd.n11 vdd.n10 98.6055
R17777 vdd.n13 vdd.n12 98.6055
R17778 vdd.n6 vdd.n5 98.6055
R17779 vdd.n4 vdd.n3 98.6055
R17780 vdd.n2 vdd.n1 98.6055
R17781 vdd.t30 vdd.n291 85.8723
R17782 vdd.t80 vdd.n236 85.8723
R17783 vdd.t137 vdd.n193 85.8723
R17784 vdd.t64 vdd.n138 85.8723
R17785 vdd.t59 vdd.n96 85.8723
R17786 vdd.t118 vdd.n41 85.8723
R17787 vdd.t138 vdd.n1740 85.8723
R17788 vdd.t78 vdd.n1795 85.8723
R17789 vdd.t130 vdd.n1642 85.8723
R17790 vdd.t60 vdd.n1697 85.8723
R17791 vdd.t96 vdd.n1545 85.8723
R17792 vdd.t14 vdd.n1600 85.8723
R17793 vdd.n2997 vdd.n856 78.546
R17794 vdd.n2436 vdd.n1029 78.546
R17795 vdd.n278 vdd.n277 75.1835
R17796 vdd.n276 vdd.n275 75.1835
R17797 vdd.n274 vdd.n273 75.1835
R17798 vdd.n272 vdd.n271 75.1835
R17799 vdd.n270 vdd.n269 75.1835
R17800 vdd.n268 vdd.n267 75.1835
R17801 vdd.n266 vdd.n265 75.1835
R17802 vdd.n180 vdd.n179 75.1835
R17803 vdd.n178 vdd.n177 75.1835
R17804 vdd.n176 vdd.n175 75.1835
R17805 vdd.n174 vdd.n173 75.1835
R17806 vdd.n172 vdd.n171 75.1835
R17807 vdd.n170 vdd.n169 75.1835
R17808 vdd.n168 vdd.n167 75.1835
R17809 vdd.n83 vdd.n82 75.1835
R17810 vdd.n81 vdd.n80 75.1835
R17811 vdd.n79 vdd.n78 75.1835
R17812 vdd.n77 vdd.n76 75.1835
R17813 vdd.n75 vdd.n74 75.1835
R17814 vdd.n73 vdd.n72 75.1835
R17815 vdd.n71 vdd.n70 75.1835
R17816 vdd.n1770 vdd.n1769 75.1835
R17817 vdd.n1772 vdd.n1771 75.1835
R17818 vdd.n1774 vdd.n1773 75.1835
R17819 vdd.n1776 vdd.n1775 75.1835
R17820 vdd.n1778 vdd.n1777 75.1835
R17821 vdd.n1780 vdd.n1779 75.1835
R17822 vdd.n1782 vdd.n1781 75.1835
R17823 vdd.n1672 vdd.n1671 75.1835
R17824 vdd.n1674 vdd.n1673 75.1835
R17825 vdd.n1676 vdd.n1675 75.1835
R17826 vdd.n1678 vdd.n1677 75.1835
R17827 vdd.n1680 vdd.n1679 75.1835
R17828 vdd.n1682 vdd.n1681 75.1835
R17829 vdd.n1684 vdd.n1683 75.1835
R17830 vdd.n1575 vdd.n1574 75.1835
R17831 vdd.n1577 vdd.n1576 75.1835
R17832 vdd.n1579 vdd.n1578 75.1835
R17833 vdd.n1581 vdd.n1580 75.1835
R17834 vdd.n1583 vdd.n1582 75.1835
R17835 vdd.n1585 vdd.n1584 75.1835
R17836 vdd.n1587 vdd.n1586 75.1835
R17837 vdd.n2927 vdd.n2660 72.8958
R17838 vdd.n2927 vdd.n2661 72.8958
R17839 vdd.n2927 vdd.n2662 72.8958
R17840 vdd.n2927 vdd.n2663 72.8958
R17841 vdd.n2927 vdd.n2664 72.8958
R17842 vdd.n2927 vdd.n2665 72.8958
R17843 vdd.n2927 vdd.n2666 72.8958
R17844 vdd.n2927 vdd.n2667 72.8958
R17845 vdd.n2927 vdd.n2668 72.8958
R17846 vdd.n2927 vdd.n2669 72.8958
R17847 vdd.n2927 vdd.n2670 72.8958
R17848 vdd.n2927 vdd.n2671 72.8958
R17849 vdd.n2927 vdd.n2672 72.8958
R17850 vdd.n2927 vdd.n2673 72.8958
R17851 vdd.n2927 vdd.n2674 72.8958
R17852 vdd.n2927 vdd.n2675 72.8958
R17853 vdd.n2927 vdd.n2676 72.8958
R17854 vdd.n772 vdd.n756 72.8958
R17855 vdd.n3165 vdd.n756 72.8958
R17856 vdd.n766 vdd.n756 72.8958
R17857 vdd.n3172 vdd.n756 72.8958
R17858 vdd.n763 vdd.n756 72.8958
R17859 vdd.n3179 vdd.n756 72.8958
R17860 vdd.n760 vdd.n756 72.8958
R17861 vdd.n3186 vdd.n756 72.8958
R17862 vdd.n3189 vdd.n756 72.8958
R17863 vdd.n3045 vdd.n756 72.8958
R17864 vdd.n3050 vdd.n756 72.8958
R17865 vdd.n3044 vdd.n756 72.8958
R17866 vdd.n3057 vdd.n756 72.8958
R17867 vdd.n3041 vdd.n756 72.8958
R17868 vdd.n3064 vdd.n756 72.8958
R17869 vdd.n3038 vdd.n756 72.8958
R17870 vdd.n3071 vdd.n756 72.8958
R17871 vdd.n2378 vdd.n1081 72.8958
R17872 vdd.n1086 vdd.n1081 72.8958
R17873 vdd.n2371 vdd.n1081 72.8958
R17874 vdd.n2365 vdd.n1081 72.8958
R17875 vdd.n2363 vdd.n1081 72.8958
R17876 vdd.n2357 vdd.n1081 72.8958
R17877 vdd.n2355 vdd.n1081 72.8958
R17878 vdd.n2349 vdd.n1081 72.8958
R17879 vdd.n2347 vdd.n1081 72.8958
R17880 vdd.n2341 vdd.n1081 72.8958
R17881 vdd.n2339 vdd.n1081 72.8958
R17882 vdd.n2333 vdd.n1081 72.8958
R17883 vdd.n2331 vdd.n1081 72.8958
R17884 vdd.n2325 vdd.n1081 72.8958
R17885 vdd.n2323 vdd.n1081 72.8958
R17886 vdd.n2316 vdd.n1081 72.8958
R17887 vdd.n2314 vdd.n1081 72.8958
R17888 vdd.n2643 vdd.n939 72.8958
R17889 vdd.n2643 vdd.n940 72.8958
R17890 vdd.n2643 vdd.n941 72.8958
R17891 vdd.n2643 vdd.n942 72.8958
R17892 vdd.n2643 vdd.n943 72.8958
R17893 vdd.n2643 vdd.n944 72.8958
R17894 vdd.n2643 vdd.n945 72.8958
R17895 vdd.n2643 vdd.n946 72.8958
R17896 vdd.n2643 vdd.n947 72.8958
R17897 vdd.n2643 vdd.n948 72.8958
R17898 vdd.n2643 vdd.n949 72.8958
R17899 vdd.n2643 vdd.n950 72.8958
R17900 vdd.n2643 vdd.n951 72.8958
R17901 vdd.n2643 vdd.n952 72.8958
R17902 vdd.n2643 vdd.n953 72.8958
R17903 vdd.n2643 vdd.n954 72.8958
R17904 vdd.n2643 vdd.n955 72.8958
R17905 vdd.n2928 vdd.n2927 72.8958
R17906 vdd.n2927 vdd.n2644 72.8958
R17907 vdd.n2927 vdd.n2645 72.8958
R17908 vdd.n2927 vdd.n2646 72.8958
R17909 vdd.n2927 vdd.n2647 72.8958
R17910 vdd.n2927 vdd.n2648 72.8958
R17911 vdd.n2927 vdd.n2649 72.8958
R17912 vdd.n2927 vdd.n2650 72.8958
R17913 vdd.n2927 vdd.n2651 72.8958
R17914 vdd.n2927 vdd.n2652 72.8958
R17915 vdd.n2927 vdd.n2653 72.8958
R17916 vdd.n2927 vdd.n2654 72.8958
R17917 vdd.n2927 vdd.n2655 72.8958
R17918 vdd.n2927 vdd.n2656 72.8958
R17919 vdd.n2927 vdd.n2657 72.8958
R17920 vdd.n2927 vdd.n2658 72.8958
R17921 vdd.n2927 vdd.n2659 72.8958
R17922 vdd.n3093 vdd.n756 72.8958
R17923 vdd.n3099 vdd.n756 72.8958
R17924 vdd.n802 vdd.n756 72.8958
R17925 vdd.n3106 vdd.n756 72.8958
R17926 vdd.n799 vdd.n756 72.8958
R17927 vdd.n3113 vdd.n756 72.8958
R17928 vdd.n796 vdd.n756 72.8958
R17929 vdd.n3120 vdd.n756 72.8958
R17930 vdd.n793 vdd.n756 72.8958
R17931 vdd.n3128 vdd.n756 72.8958
R17932 vdd.n790 vdd.n756 72.8958
R17933 vdd.n3135 vdd.n756 72.8958
R17934 vdd.n787 vdd.n756 72.8958
R17935 vdd.n3142 vdd.n756 72.8958
R17936 vdd.n784 vdd.n756 72.8958
R17937 vdd.n3149 vdd.n756 72.8958
R17938 vdd.n3152 vdd.n756 72.8958
R17939 vdd.n2643 vdd.n937 72.8958
R17940 vdd.n2643 vdd.n936 72.8958
R17941 vdd.n2643 vdd.n935 72.8958
R17942 vdd.n2643 vdd.n934 72.8958
R17943 vdd.n2643 vdd.n933 72.8958
R17944 vdd.n2643 vdd.n932 72.8958
R17945 vdd.n2643 vdd.n931 72.8958
R17946 vdd.n2643 vdd.n930 72.8958
R17947 vdd.n2643 vdd.n929 72.8958
R17948 vdd.n2643 vdd.n928 72.8958
R17949 vdd.n2643 vdd.n927 72.8958
R17950 vdd.n2643 vdd.n926 72.8958
R17951 vdd.n2643 vdd.n925 72.8958
R17952 vdd.n2643 vdd.n924 72.8958
R17953 vdd.n2643 vdd.n923 72.8958
R17954 vdd.n2643 vdd.n922 72.8958
R17955 vdd.n2643 vdd.n921 72.8958
R17956 vdd.n2132 vdd.n1081 72.8958
R17957 vdd.n2134 vdd.n1081 72.8958
R17958 vdd.n2140 vdd.n1081 72.8958
R17959 vdd.n2142 vdd.n1081 72.8958
R17960 vdd.n2148 vdd.n1081 72.8958
R17961 vdd.n2150 vdd.n1081 72.8958
R17962 vdd.n2156 vdd.n1081 72.8958
R17963 vdd.n2158 vdd.n1081 72.8958
R17964 vdd.n2164 vdd.n1081 72.8958
R17965 vdd.n2166 vdd.n1081 72.8958
R17966 vdd.n2172 vdd.n1081 72.8958
R17967 vdd.n2174 vdd.n1081 72.8958
R17968 vdd.n2180 vdd.n1081 72.8958
R17969 vdd.n2182 vdd.n1081 72.8958
R17970 vdd.n2188 vdd.n1081 72.8958
R17971 vdd.n2190 vdd.n1081 72.8958
R17972 vdd.n2197 vdd.n1081 72.8958
R17973 vdd.n1454 vdd.n1453 66.2847
R17974 vdd.n1454 vdd.n1232 66.2847
R17975 vdd.n1454 vdd.n1233 66.2847
R17976 vdd.n1454 vdd.n1234 66.2847
R17977 vdd.n1454 vdd.n1235 66.2847
R17978 vdd.n1454 vdd.n1236 66.2847
R17979 vdd.n1454 vdd.n1237 66.2847
R17980 vdd.n1454 vdd.n1238 66.2847
R17981 vdd.n1454 vdd.n1239 66.2847
R17982 vdd.n1454 vdd.n1240 66.2847
R17983 vdd.n1454 vdd.n1241 66.2847
R17984 vdd.n1454 vdd.n1242 66.2847
R17985 vdd.n1454 vdd.n1243 66.2847
R17986 vdd.n1454 vdd.n1244 66.2847
R17987 vdd.n1454 vdd.n1245 66.2847
R17988 vdd.n1454 vdd.n1246 66.2847
R17989 vdd.n1454 vdd.n1247 66.2847
R17990 vdd.n1454 vdd.n1248 66.2847
R17991 vdd.n1454 vdd.n1249 66.2847
R17992 vdd.n1454 vdd.n1250 66.2847
R17993 vdd.n1454 vdd.n1251 66.2847
R17994 vdd.n1454 vdd.n1252 66.2847
R17995 vdd.n1454 vdd.n1253 66.2847
R17996 vdd.n1454 vdd.n1254 66.2847
R17997 vdd.n1454 vdd.n1255 66.2847
R17998 vdd.n1454 vdd.n1256 66.2847
R17999 vdd.n1454 vdd.n1257 66.2847
R18000 vdd.n1454 vdd.n1258 66.2847
R18001 vdd.n1454 vdd.n1259 66.2847
R18002 vdd.n1454 vdd.n1260 66.2847
R18003 vdd.n1454 vdd.n1261 66.2847
R18004 vdd.n1125 vdd.n1121 66.2847
R18005 vdd.n1997 vdd.n1125 66.2847
R18006 vdd.n2002 vdd.n1125 66.2847
R18007 vdd.n2007 vdd.n1125 66.2847
R18008 vdd.n1995 vdd.n1125 66.2847
R18009 vdd.n2014 vdd.n1125 66.2847
R18010 vdd.n1987 vdd.n1125 66.2847
R18011 vdd.n2021 vdd.n1125 66.2847
R18012 vdd.n1980 vdd.n1125 66.2847
R18013 vdd.n2028 vdd.n1125 66.2847
R18014 vdd.n1974 vdd.n1125 66.2847
R18015 vdd.n1969 vdd.n1125 66.2847
R18016 vdd.n2039 vdd.n1125 66.2847
R18017 vdd.n1961 vdd.n1125 66.2847
R18018 vdd.n2046 vdd.n1125 66.2847
R18019 vdd.n1954 vdd.n1125 66.2847
R18020 vdd.n2053 vdd.n1125 66.2847
R18021 vdd.n1947 vdd.n1125 66.2847
R18022 vdd.n2060 vdd.n1125 66.2847
R18023 vdd.n1940 vdd.n1125 66.2847
R18024 vdd.n2067 vdd.n1125 66.2847
R18025 vdd.n1934 vdd.n1125 66.2847
R18026 vdd.n1929 vdd.n1125 66.2847
R18027 vdd.n2078 vdd.n1125 66.2847
R18028 vdd.n1921 vdd.n1125 66.2847
R18029 vdd.n2085 vdd.n1125 66.2847
R18030 vdd.n1914 vdd.n1125 66.2847
R18031 vdd.n2092 vdd.n1125 66.2847
R18032 vdd.n2095 vdd.n1125 66.2847
R18033 vdd.n1905 vdd.n1125 66.2847
R18034 vdd.n2104 vdd.n1125 66.2847
R18035 vdd.n1899 vdd.n1125 66.2847
R18036 vdd.n3319 vdd.n658 66.2847
R18037 vdd.n663 vdd.n658 66.2847
R18038 vdd.n666 vdd.n658 66.2847
R18039 vdd.n3308 vdd.n658 66.2847
R18040 vdd.n3302 vdd.n658 66.2847
R18041 vdd.n3300 vdd.n658 66.2847
R18042 vdd.n3294 vdd.n658 66.2847
R18043 vdd.n3292 vdd.n658 66.2847
R18044 vdd.n3286 vdd.n658 66.2847
R18045 vdd.n3284 vdd.n658 66.2847
R18046 vdd.n3278 vdd.n658 66.2847
R18047 vdd.n3276 vdd.n658 66.2847
R18048 vdd.n3270 vdd.n658 66.2847
R18049 vdd.n3268 vdd.n658 66.2847
R18050 vdd.n3262 vdd.n658 66.2847
R18051 vdd.n3260 vdd.n658 66.2847
R18052 vdd.n3254 vdd.n658 66.2847
R18053 vdd.n3252 vdd.n658 66.2847
R18054 vdd.n3246 vdd.n658 66.2847
R18055 vdd.n3244 vdd.n658 66.2847
R18056 vdd.n727 vdd.n658 66.2847
R18057 vdd.n3235 vdd.n658 66.2847
R18058 vdd.n729 vdd.n658 66.2847
R18059 vdd.n3228 vdd.n658 66.2847
R18060 vdd.n3222 vdd.n658 66.2847
R18061 vdd.n3220 vdd.n658 66.2847
R18062 vdd.n3214 vdd.n658 66.2847
R18063 vdd.n3212 vdd.n658 66.2847
R18064 vdd.n3206 vdd.n658 66.2847
R18065 vdd.n750 vdd.n658 66.2847
R18066 vdd.n752 vdd.n658 66.2847
R18067 vdd.n3435 vdd.n3434 66.2847
R18068 vdd.n3435 vdd.n403 66.2847
R18069 vdd.n3435 vdd.n402 66.2847
R18070 vdd.n3435 vdd.n401 66.2847
R18071 vdd.n3435 vdd.n400 66.2847
R18072 vdd.n3435 vdd.n399 66.2847
R18073 vdd.n3435 vdd.n398 66.2847
R18074 vdd.n3435 vdd.n397 66.2847
R18075 vdd.n3435 vdd.n396 66.2847
R18076 vdd.n3435 vdd.n395 66.2847
R18077 vdd.n3435 vdd.n394 66.2847
R18078 vdd.n3435 vdd.n393 66.2847
R18079 vdd.n3435 vdd.n392 66.2847
R18080 vdd.n3435 vdd.n391 66.2847
R18081 vdd.n3435 vdd.n390 66.2847
R18082 vdd.n3435 vdd.n389 66.2847
R18083 vdd.n3435 vdd.n388 66.2847
R18084 vdd.n3435 vdd.n387 66.2847
R18085 vdd.n3435 vdd.n386 66.2847
R18086 vdd.n3435 vdd.n385 66.2847
R18087 vdd.n3435 vdd.n384 66.2847
R18088 vdd.n3435 vdd.n383 66.2847
R18089 vdd.n3435 vdd.n382 66.2847
R18090 vdd.n3435 vdd.n381 66.2847
R18091 vdd.n3435 vdd.n380 66.2847
R18092 vdd.n3435 vdd.n379 66.2847
R18093 vdd.n3435 vdd.n378 66.2847
R18094 vdd.n3435 vdd.n377 66.2847
R18095 vdd.n3435 vdd.n376 66.2847
R18096 vdd.n3435 vdd.n375 66.2847
R18097 vdd.n3435 vdd.n374 66.2847
R18098 vdd.n3435 vdd.n373 66.2847
R18099 vdd.n448 vdd.n373 52.4337
R18100 vdd.n454 vdd.n374 52.4337
R18101 vdd.n458 vdd.n375 52.4337
R18102 vdd.n464 vdd.n376 52.4337
R18103 vdd.n468 vdd.n377 52.4337
R18104 vdd.n474 vdd.n378 52.4337
R18105 vdd.n478 vdd.n379 52.4337
R18106 vdd.n484 vdd.n380 52.4337
R18107 vdd.n488 vdd.n381 52.4337
R18108 vdd.n494 vdd.n382 52.4337
R18109 vdd.n498 vdd.n383 52.4337
R18110 vdd.n504 vdd.n384 52.4337
R18111 vdd.n508 vdd.n385 52.4337
R18112 vdd.n514 vdd.n386 52.4337
R18113 vdd.n518 vdd.n387 52.4337
R18114 vdd.n524 vdd.n388 52.4337
R18115 vdd.n528 vdd.n389 52.4337
R18116 vdd.n534 vdd.n390 52.4337
R18117 vdd.n538 vdd.n391 52.4337
R18118 vdd.n544 vdd.n392 52.4337
R18119 vdd.n548 vdd.n393 52.4337
R18120 vdd.n554 vdd.n394 52.4337
R18121 vdd.n558 vdd.n395 52.4337
R18122 vdd.n564 vdd.n396 52.4337
R18123 vdd.n568 vdd.n397 52.4337
R18124 vdd.n574 vdd.n398 52.4337
R18125 vdd.n578 vdd.n399 52.4337
R18126 vdd.n584 vdd.n400 52.4337
R18127 vdd.n588 vdd.n401 52.4337
R18128 vdd.n594 vdd.n402 52.4337
R18129 vdd.n597 vdd.n403 52.4337
R18130 vdd.n3434 vdd.n3433 52.4337
R18131 vdd.n3319 vdd.n660 52.4337
R18132 vdd.n3317 vdd.n663 52.4337
R18133 vdd.n3313 vdd.n666 52.4337
R18134 vdd.n3309 vdd.n3308 52.4337
R18135 vdd.n3302 vdd.n669 52.4337
R18136 vdd.n3301 vdd.n3300 52.4337
R18137 vdd.n3294 vdd.n675 52.4337
R18138 vdd.n3293 vdd.n3292 52.4337
R18139 vdd.n3286 vdd.n681 52.4337
R18140 vdd.n3285 vdd.n3284 52.4337
R18141 vdd.n3278 vdd.n689 52.4337
R18142 vdd.n3277 vdd.n3276 52.4337
R18143 vdd.n3270 vdd.n695 52.4337
R18144 vdd.n3269 vdd.n3268 52.4337
R18145 vdd.n3262 vdd.n701 52.4337
R18146 vdd.n3261 vdd.n3260 52.4337
R18147 vdd.n3254 vdd.n707 52.4337
R18148 vdd.n3253 vdd.n3252 52.4337
R18149 vdd.n3246 vdd.n713 52.4337
R18150 vdd.n3245 vdd.n3244 52.4337
R18151 vdd.n727 vdd.n719 52.4337
R18152 vdd.n3236 vdd.n3235 52.4337
R18153 vdd.n3233 vdd.n729 52.4337
R18154 vdd.n3229 vdd.n3228 52.4337
R18155 vdd.n3222 vdd.n733 52.4337
R18156 vdd.n3221 vdd.n3220 52.4337
R18157 vdd.n3214 vdd.n739 52.4337
R18158 vdd.n3213 vdd.n3212 52.4337
R18159 vdd.n3206 vdd.n745 52.4337
R18160 vdd.n3205 vdd.n750 52.4337
R18161 vdd.n3201 vdd.n752 52.4337
R18162 vdd.n2106 vdd.n1899 52.4337
R18163 vdd.n2104 vdd.n2103 52.4337
R18164 vdd.n1906 vdd.n1905 52.4337
R18165 vdd.n2095 vdd.n2094 52.4337
R18166 vdd.n2092 vdd.n2091 52.4337
R18167 vdd.n2087 vdd.n1914 52.4337
R18168 vdd.n2085 vdd.n2084 52.4337
R18169 vdd.n2080 vdd.n1921 52.4337
R18170 vdd.n2078 vdd.n2077 52.4337
R18171 vdd.n1930 vdd.n1929 52.4337
R18172 vdd.n2069 vdd.n1934 52.4337
R18173 vdd.n2067 vdd.n2066 52.4337
R18174 vdd.n2062 vdd.n1940 52.4337
R18175 vdd.n2060 vdd.n2059 52.4337
R18176 vdd.n2055 vdd.n1947 52.4337
R18177 vdd.n2053 vdd.n2052 52.4337
R18178 vdd.n2048 vdd.n1954 52.4337
R18179 vdd.n2046 vdd.n2045 52.4337
R18180 vdd.n2041 vdd.n1961 52.4337
R18181 vdd.n2039 vdd.n2038 52.4337
R18182 vdd.n1970 vdd.n1969 52.4337
R18183 vdd.n2030 vdd.n1974 52.4337
R18184 vdd.n2028 vdd.n2027 52.4337
R18185 vdd.n2023 vdd.n1980 52.4337
R18186 vdd.n2021 vdd.n2020 52.4337
R18187 vdd.n2016 vdd.n1987 52.4337
R18188 vdd.n2014 vdd.n2013 52.4337
R18189 vdd.n2009 vdd.n1995 52.4337
R18190 vdd.n2007 vdd.n2006 52.4337
R18191 vdd.n2002 vdd.n2001 52.4337
R18192 vdd.n1997 vdd.n1996 52.4337
R18193 vdd.n2115 vdd.n1121 52.4337
R18194 vdd.n1453 vdd.n1452 52.4337
R18195 vdd.n1267 vdd.n1232 52.4337
R18196 vdd.n1269 vdd.n1233 52.4337
R18197 vdd.n1273 vdd.n1234 52.4337
R18198 vdd.n1275 vdd.n1235 52.4337
R18199 vdd.n1279 vdd.n1236 52.4337
R18200 vdd.n1281 vdd.n1237 52.4337
R18201 vdd.n1285 vdd.n1238 52.4337
R18202 vdd.n1287 vdd.n1239 52.4337
R18203 vdd.n1419 vdd.n1240 52.4337
R18204 vdd.n1291 vdd.n1241 52.4337
R18205 vdd.n1295 vdd.n1242 52.4337
R18206 vdd.n1297 vdd.n1243 52.4337
R18207 vdd.n1301 vdd.n1244 52.4337
R18208 vdd.n1303 vdd.n1245 52.4337
R18209 vdd.n1307 vdd.n1246 52.4337
R18210 vdd.n1309 vdd.n1247 52.4337
R18211 vdd.n1313 vdd.n1248 52.4337
R18212 vdd.n1315 vdd.n1249 52.4337
R18213 vdd.n1319 vdd.n1250 52.4337
R18214 vdd.n1383 vdd.n1251 52.4337
R18215 vdd.n1324 vdd.n1252 52.4337
R18216 vdd.n1326 vdd.n1253 52.4337
R18217 vdd.n1330 vdd.n1254 52.4337
R18218 vdd.n1332 vdd.n1255 52.4337
R18219 vdd.n1336 vdd.n1256 52.4337
R18220 vdd.n1338 vdd.n1257 52.4337
R18221 vdd.n1342 vdd.n1258 52.4337
R18222 vdd.n1344 vdd.n1259 52.4337
R18223 vdd.n1348 vdd.n1260 52.4337
R18224 vdd.n1350 vdd.n1261 52.4337
R18225 vdd.n1453 vdd.n1263 52.4337
R18226 vdd.n1268 vdd.n1232 52.4337
R18227 vdd.n1272 vdd.n1233 52.4337
R18228 vdd.n1274 vdd.n1234 52.4337
R18229 vdd.n1278 vdd.n1235 52.4337
R18230 vdd.n1280 vdd.n1236 52.4337
R18231 vdd.n1284 vdd.n1237 52.4337
R18232 vdd.n1286 vdd.n1238 52.4337
R18233 vdd.n1418 vdd.n1239 52.4337
R18234 vdd.n1290 vdd.n1240 52.4337
R18235 vdd.n1294 vdd.n1241 52.4337
R18236 vdd.n1296 vdd.n1242 52.4337
R18237 vdd.n1300 vdd.n1243 52.4337
R18238 vdd.n1302 vdd.n1244 52.4337
R18239 vdd.n1306 vdd.n1245 52.4337
R18240 vdd.n1308 vdd.n1246 52.4337
R18241 vdd.n1312 vdd.n1247 52.4337
R18242 vdd.n1314 vdd.n1248 52.4337
R18243 vdd.n1318 vdd.n1249 52.4337
R18244 vdd.n1320 vdd.n1250 52.4337
R18245 vdd.n1323 vdd.n1251 52.4337
R18246 vdd.n1325 vdd.n1252 52.4337
R18247 vdd.n1329 vdd.n1253 52.4337
R18248 vdd.n1331 vdd.n1254 52.4337
R18249 vdd.n1335 vdd.n1255 52.4337
R18250 vdd.n1337 vdd.n1256 52.4337
R18251 vdd.n1341 vdd.n1257 52.4337
R18252 vdd.n1343 vdd.n1258 52.4337
R18253 vdd.n1347 vdd.n1259 52.4337
R18254 vdd.n1349 vdd.n1260 52.4337
R18255 vdd.n1261 vdd.n1231 52.4337
R18256 vdd.n1121 vdd.n1120 52.4337
R18257 vdd.n1998 vdd.n1997 52.4337
R18258 vdd.n2003 vdd.n2002 52.4337
R18259 vdd.n2008 vdd.n2007 52.4337
R18260 vdd.n1995 vdd.n1988 52.4337
R18261 vdd.n2015 vdd.n2014 52.4337
R18262 vdd.n1987 vdd.n1981 52.4337
R18263 vdd.n2022 vdd.n2021 52.4337
R18264 vdd.n1980 vdd.n1975 52.4337
R18265 vdd.n2029 vdd.n2028 52.4337
R18266 vdd.n1974 vdd.n1973 52.4337
R18267 vdd.n1969 vdd.n1962 52.4337
R18268 vdd.n2040 vdd.n2039 52.4337
R18269 vdd.n1961 vdd.n1955 52.4337
R18270 vdd.n2047 vdd.n2046 52.4337
R18271 vdd.n1954 vdd.n1948 52.4337
R18272 vdd.n2054 vdd.n2053 52.4337
R18273 vdd.n1947 vdd.n1941 52.4337
R18274 vdd.n2061 vdd.n2060 52.4337
R18275 vdd.n1940 vdd.n1935 52.4337
R18276 vdd.n2068 vdd.n2067 52.4337
R18277 vdd.n1934 vdd.n1933 52.4337
R18278 vdd.n1929 vdd.n1922 52.4337
R18279 vdd.n2079 vdd.n2078 52.4337
R18280 vdd.n1921 vdd.n1915 52.4337
R18281 vdd.n2086 vdd.n2085 52.4337
R18282 vdd.n1914 vdd.n1908 52.4337
R18283 vdd.n2093 vdd.n2092 52.4337
R18284 vdd.n2096 vdd.n2095 52.4337
R18285 vdd.n1905 vdd.n1900 52.4337
R18286 vdd.n2105 vdd.n2104 52.4337
R18287 vdd.n1899 vdd.n1127 52.4337
R18288 vdd.n3320 vdd.n3319 52.4337
R18289 vdd.n3314 vdd.n663 52.4337
R18290 vdd.n3310 vdd.n666 52.4337
R18291 vdd.n3308 vdd.n3307 52.4337
R18292 vdd.n3303 vdd.n3302 52.4337
R18293 vdd.n3300 vdd.n3299 52.4337
R18294 vdd.n3295 vdd.n3294 52.4337
R18295 vdd.n3292 vdd.n3291 52.4337
R18296 vdd.n3287 vdd.n3286 52.4337
R18297 vdd.n3284 vdd.n3283 52.4337
R18298 vdd.n3279 vdd.n3278 52.4337
R18299 vdd.n3276 vdd.n3275 52.4337
R18300 vdd.n3271 vdd.n3270 52.4337
R18301 vdd.n3268 vdd.n3267 52.4337
R18302 vdd.n3263 vdd.n3262 52.4337
R18303 vdd.n3260 vdd.n3259 52.4337
R18304 vdd.n3255 vdd.n3254 52.4337
R18305 vdd.n3252 vdd.n3251 52.4337
R18306 vdd.n3247 vdd.n3246 52.4337
R18307 vdd.n3244 vdd.n3243 52.4337
R18308 vdd.n728 vdd.n727 52.4337
R18309 vdd.n3235 vdd.n3234 52.4337
R18310 vdd.n3230 vdd.n729 52.4337
R18311 vdd.n3228 vdd.n3227 52.4337
R18312 vdd.n3223 vdd.n3222 52.4337
R18313 vdd.n3220 vdd.n3219 52.4337
R18314 vdd.n3215 vdd.n3214 52.4337
R18315 vdd.n3212 vdd.n3211 52.4337
R18316 vdd.n3207 vdd.n3206 52.4337
R18317 vdd.n3202 vdd.n750 52.4337
R18318 vdd.n3198 vdd.n752 52.4337
R18319 vdd.n3434 vdd.n404 52.4337
R18320 vdd.n595 vdd.n403 52.4337
R18321 vdd.n589 vdd.n402 52.4337
R18322 vdd.n585 vdd.n401 52.4337
R18323 vdd.n579 vdd.n400 52.4337
R18324 vdd.n575 vdd.n399 52.4337
R18325 vdd.n569 vdd.n398 52.4337
R18326 vdd.n565 vdd.n397 52.4337
R18327 vdd.n559 vdd.n396 52.4337
R18328 vdd.n555 vdd.n395 52.4337
R18329 vdd.n549 vdd.n394 52.4337
R18330 vdd.n545 vdd.n393 52.4337
R18331 vdd.n539 vdd.n392 52.4337
R18332 vdd.n535 vdd.n391 52.4337
R18333 vdd.n529 vdd.n390 52.4337
R18334 vdd.n525 vdd.n389 52.4337
R18335 vdd.n519 vdd.n388 52.4337
R18336 vdd.n515 vdd.n387 52.4337
R18337 vdd.n509 vdd.n386 52.4337
R18338 vdd.n505 vdd.n385 52.4337
R18339 vdd.n499 vdd.n384 52.4337
R18340 vdd.n495 vdd.n383 52.4337
R18341 vdd.n489 vdd.n382 52.4337
R18342 vdd.n485 vdd.n381 52.4337
R18343 vdd.n479 vdd.n380 52.4337
R18344 vdd.n475 vdd.n379 52.4337
R18345 vdd.n469 vdd.n378 52.4337
R18346 vdd.n465 vdd.n377 52.4337
R18347 vdd.n459 vdd.n376 52.4337
R18348 vdd.n455 vdd.n375 52.4337
R18349 vdd.n449 vdd.n374 52.4337
R18350 vdd.n445 vdd.n373 52.4337
R18351 vdd.t250 vdd.t233 51.4683
R18352 vdd.n266 vdd.n264 42.0461
R18353 vdd.n168 vdd.n166 42.0461
R18354 vdd.n71 vdd.n69 42.0461
R18355 vdd.n1770 vdd.n1768 42.0461
R18356 vdd.n1672 vdd.n1670 42.0461
R18357 vdd.n1575 vdd.n1573 42.0461
R18358 vdd.n320 vdd.n319 41.6884
R18359 vdd.n222 vdd.n221 41.6884
R18360 vdd.n125 vdd.n124 41.6884
R18361 vdd.n1824 vdd.n1823 41.6884
R18362 vdd.n1726 vdd.n1725 41.6884
R18363 vdd.n1629 vdd.n1628 41.6884
R18364 vdd.n1230 vdd.n1229 41.1157
R18365 vdd.n1386 vdd.n1385 41.1157
R18366 vdd.n1422 vdd.n1421 41.1157
R18367 vdd.n407 vdd.n406 41.1157
R18368 vdd.n547 vdd.n420 41.1157
R18369 vdd.n433 vdd.n432 41.1157
R18370 vdd.n3152 vdd.n3151 39.2114
R18371 vdd.n3149 vdd.n3148 39.2114
R18372 vdd.n3144 vdd.n784 39.2114
R18373 vdd.n3142 vdd.n3141 39.2114
R18374 vdd.n3137 vdd.n787 39.2114
R18375 vdd.n3135 vdd.n3134 39.2114
R18376 vdd.n3130 vdd.n790 39.2114
R18377 vdd.n3128 vdd.n3127 39.2114
R18378 vdd.n3122 vdd.n793 39.2114
R18379 vdd.n3120 vdd.n3119 39.2114
R18380 vdd.n3115 vdd.n796 39.2114
R18381 vdd.n3113 vdd.n3112 39.2114
R18382 vdd.n3108 vdd.n799 39.2114
R18383 vdd.n3106 vdd.n3105 39.2114
R18384 vdd.n3101 vdd.n802 39.2114
R18385 vdd.n3099 vdd.n3098 39.2114
R18386 vdd.n3094 vdd.n3093 39.2114
R18387 vdd.n2928 vdd.n918 39.2114
R18388 vdd.n2749 vdd.n2644 39.2114
R18389 vdd.n2753 vdd.n2645 39.2114
R18390 vdd.n2757 vdd.n2646 39.2114
R18391 vdd.n2761 vdd.n2647 39.2114
R18392 vdd.n2765 vdd.n2648 39.2114
R18393 vdd.n2769 vdd.n2649 39.2114
R18394 vdd.n2773 vdd.n2650 39.2114
R18395 vdd.n2777 vdd.n2651 39.2114
R18396 vdd.n2781 vdd.n2652 39.2114
R18397 vdd.n2785 vdd.n2653 39.2114
R18398 vdd.n2789 vdd.n2654 39.2114
R18399 vdd.n2793 vdd.n2655 39.2114
R18400 vdd.n2797 vdd.n2656 39.2114
R18401 vdd.n2801 vdd.n2657 39.2114
R18402 vdd.n2805 vdd.n2658 39.2114
R18403 vdd.n2810 vdd.n2659 39.2114
R18404 vdd.n2638 vdd.n955 39.2114
R18405 vdd.n2634 vdd.n954 39.2114
R18406 vdd.n2630 vdd.n953 39.2114
R18407 vdd.n2626 vdd.n952 39.2114
R18408 vdd.n2622 vdd.n951 39.2114
R18409 vdd.n2618 vdd.n950 39.2114
R18410 vdd.n2614 vdd.n949 39.2114
R18411 vdd.n2610 vdd.n948 39.2114
R18412 vdd.n2606 vdd.n947 39.2114
R18413 vdd.n2602 vdd.n946 39.2114
R18414 vdd.n2598 vdd.n945 39.2114
R18415 vdd.n2594 vdd.n944 39.2114
R18416 vdd.n2590 vdd.n943 39.2114
R18417 vdd.n2586 vdd.n942 39.2114
R18418 vdd.n2582 vdd.n941 39.2114
R18419 vdd.n2577 vdd.n940 39.2114
R18420 vdd.n2573 vdd.n939 39.2114
R18421 vdd.n2378 vdd.n1084 39.2114
R18422 vdd.n2376 vdd.n1086 39.2114
R18423 vdd.n2372 vdd.n2371 39.2114
R18424 vdd.n2365 vdd.n1088 39.2114
R18425 vdd.n2364 vdd.n2363 39.2114
R18426 vdd.n2357 vdd.n1090 39.2114
R18427 vdd.n2356 vdd.n2355 39.2114
R18428 vdd.n2349 vdd.n1092 39.2114
R18429 vdd.n2348 vdd.n2347 39.2114
R18430 vdd.n2341 vdd.n1094 39.2114
R18431 vdd.n2340 vdd.n2339 39.2114
R18432 vdd.n2333 vdd.n1096 39.2114
R18433 vdd.n2332 vdd.n2331 39.2114
R18434 vdd.n2325 vdd.n1098 39.2114
R18435 vdd.n2324 vdd.n2323 39.2114
R18436 vdd.n2316 vdd.n1100 39.2114
R18437 vdd.n2315 vdd.n2314 39.2114
R18438 vdd.n3071 vdd.n3070 39.2114
R18439 vdd.n3066 vdd.n3038 39.2114
R18440 vdd.n3064 vdd.n3063 39.2114
R18441 vdd.n3059 vdd.n3041 39.2114
R18442 vdd.n3057 vdd.n3056 39.2114
R18443 vdd.n3052 vdd.n3044 39.2114
R18444 vdd.n3050 vdd.n3049 39.2114
R18445 vdd.n3045 vdd.n755 39.2114
R18446 vdd.n3189 vdd.n3188 39.2114
R18447 vdd.n3186 vdd.n3185 39.2114
R18448 vdd.n3181 vdd.n760 39.2114
R18449 vdd.n3179 vdd.n3178 39.2114
R18450 vdd.n3174 vdd.n763 39.2114
R18451 vdd.n3172 vdd.n3171 39.2114
R18452 vdd.n3167 vdd.n766 39.2114
R18453 vdd.n3165 vdd.n3164 39.2114
R18454 vdd.n3160 vdd.n772 39.2114
R18455 vdd.n2660 vdd.n914 39.2114
R18456 vdd.n2683 vdd.n2661 39.2114
R18457 vdd.n2687 vdd.n2662 39.2114
R18458 vdd.n2691 vdd.n2663 39.2114
R18459 vdd.n2695 vdd.n2664 39.2114
R18460 vdd.n2699 vdd.n2665 39.2114
R18461 vdd.n2703 vdd.n2666 39.2114
R18462 vdd.n2707 vdd.n2667 39.2114
R18463 vdd.n2711 vdd.n2668 39.2114
R18464 vdd.n2715 vdd.n2669 39.2114
R18465 vdd.n2719 vdd.n2670 39.2114
R18466 vdd.n2723 vdd.n2671 39.2114
R18467 vdd.n2727 vdd.n2672 39.2114
R18468 vdd.n2731 vdd.n2673 39.2114
R18469 vdd.n2735 vdd.n2674 39.2114
R18470 vdd.n2739 vdd.n2675 39.2114
R18471 vdd.n2743 vdd.n2676 39.2114
R18472 vdd.n2682 vdd.n2660 39.2114
R18473 vdd.n2686 vdd.n2661 39.2114
R18474 vdd.n2690 vdd.n2662 39.2114
R18475 vdd.n2694 vdd.n2663 39.2114
R18476 vdd.n2698 vdd.n2664 39.2114
R18477 vdd.n2702 vdd.n2665 39.2114
R18478 vdd.n2706 vdd.n2666 39.2114
R18479 vdd.n2710 vdd.n2667 39.2114
R18480 vdd.n2714 vdd.n2668 39.2114
R18481 vdd.n2718 vdd.n2669 39.2114
R18482 vdd.n2722 vdd.n2670 39.2114
R18483 vdd.n2726 vdd.n2671 39.2114
R18484 vdd.n2730 vdd.n2672 39.2114
R18485 vdd.n2734 vdd.n2673 39.2114
R18486 vdd.n2738 vdd.n2674 39.2114
R18487 vdd.n2742 vdd.n2675 39.2114
R18488 vdd.n2677 vdd.n2676 39.2114
R18489 vdd.n772 vdd.n767 39.2114
R18490 vdd.n3166 vdd.n3165 39.2114
R18491 vdd.n766 vdd.n764 39.2114
R18492 vdd.n3173 vdd.n3172 39.2114
R18493 vdd.n763 vdd.n761 39.2114
R18494 vdd.n3180 vdd.n3179 39.2114
R18495 vdd.n760 vdd.n758 39.2114
R18496 vdd.n3187 vdd.n3186 39.2114
R18497 vdd.n3190 vdd.n3189 39.2114
R18498 vdd.n3046 vdd.n3045 39.2114
R18499 vdd.n3051 vdd.n3050 39.2114
R18500 vdd.n3044 vdd.n3042 39.2114
R18501 vdd.n3058 vdd.n3057 39.2114
R18502 vdd.n3041 vdd.n3039 39.2114
R18503 vdd.n3065 vdd.n3064 39.2114
R18504 vdd.n3038 vdd.n3036 39.2114
R18505 vdd.n3072 vdd.n3071 39.2114
R18506 vdd.n2379 vdd.n2378 39.2114
R18507 vdd.n2373 vdd.n1086 39.2114
R18508 vdd.n2371 vdd.n2370 39.2114
R18509 vdd.n2366 vdd.n2365 39.2114
R18510 vdd.n2363 vdd.n2362 39.2114
R18511 vdd.n2358 vdd.n2357 39.2114
R18512 vdd.n2355 vdd.n2354 39.2114
R18513 vdd.n2350 vdd.n2349 39.2114
R18514 vdd.n2347 vdd.n2346 39.2114
R18515 vdd.n2342 vdd.n2341 39.2114
R18516 vdd.n2339 vdd.n2338 39.2114
R18517 vdd.n2334 vdd.n2333 39.2114
R18518 vdd.n2331 vdd.n2330 39.2114
R18519 vdd.n2326 vdd.n2325 39.2114
R18520 vdd.n2323 vdd.n2322 39.2114
R18521 vdd.n2317 vdd.n2316 39.2114
R18522 vdd.n2314 vdd.n2313 39.2114
R18523 vdd.n2576 vdd.n939 39.2114
R18524 vdd.n2581 vdd.n940 39.2114
R18525 vdd.n2585 vdd.n941 39.2114
R18526 vdd.n2589 vdd.n942 39.2114
R18527 vdd.n2593 vdd.n943 39.2114
R18528 vdd.n2597 vdd.n944 39.2114
R18529 vdd.n2601 vdd.n945 39.2114
R18530 vdd.n2605 vdd.n946 39.2114
R18531 vdd.n2609 vdd.n947 39.2114
R18532 vdd.n2613 vdd.n948 39.2114
R18533 vdd.n2617 vdd.n949 39.2114
R18534 vdd.n2621 vdd.n950 39.2114
R18535 vdd.n2625 vdd.n951 39.2114
R18536 vdd.n2629 vdd.n952 39.2114
R18537 vdd.n2633 vdd.n953 39.2114
R18538 vdd.n2637 vdd.n954 39.2114
R18539 vdd.n957 vdd.n955 39.2114
R18540 vdd.n2929 vdd.n2928 39.2114
R18541 vdd.n2752 vdd.n2644 39.2114
R18542 vdd.n2756 vdd.n2645 39.2114
R18543 vdd.n2760 vdd.n2646 39.2114
R18544 vdd.n2764 vdd.n2647 39.2114
R18545 vdd.n2768 vdd.n2648 39.2114
R18546 vdd.n2772 vdd.n2649 39.2114
R18547 vdd.n2776 vdd.n2650 39.2114
R18548 vdd.n2780 vdd.n2651 39.2114
R18549 vdd.n2784 vdd.n2652 39.2114
R18550 vdd.n2788 vdd.n2653 39.2114
R18551 vdd.n2792 vdd.n2654 39.2114
R18552 vdd.n2796 vdd.n2655 39.2114
R18553 vdd.n2800 vdd.n2656 39.2114
R18554 vdd.n2804 vdd.n2657 39.2114
R18555 vdd.n2809 vdd.n2658 39.2114
R18556 vdd.n2812 vdd.n2659 39.2114
R18557 vdd.n3093 vdd.n803 39.2114
R18558 vdd.n3100 vdd.n3099 39.2114
R18559 vdd.n802 vdd.n800 39.2114
R18560 vdd.n3107 vdd.n3106 39.2114
R18561 vdd.n799 vdd.n797 39.2114
R18562 vdd.n3114 vdd.n3113 39.2114
R18563 vdd.n796 vdd.n794 39.2114
R18564 vdd.n3121 vdd.n3120 39.2114
R18565 vdd.n793 vdd.n791 39.2114
R18566 vdd.n3129 vdd.n3128 39.2114
R18567 vdd.n790 vdd.n788 39.2114
R18568 vdd.n3136 vdd.n3135 39.2114
R18569 vdd.n787 vdd.n785 39.2114
R18570 vdd.n3143 vdd.n3142 39.2114
R18571 vdd.n784 vdd.n782 39.2114
R18572 vdd.n3150 vdd.n3149 39.2114
R18573 vdd.n3153 vdd.n3152 39.2114
R18574 vdd.n966 vdd.n921 39.2114
R18575 vdd.n2565 vdd.n922 39.2114
R18576 vdd.n2561 vdd.n923 39.2114
R18577 vdd.n2557 vdd.n924 39.2114
R18578 vdd.n2553 vdd.n925 39.2114
R18579 vdd.n2549 vdd.n926 39.2114
R18580 vdd.n2545 vdd.n927 39.2114
R18581 vdd.n2541 vdd.n928 39.2114
R18582 vdd.n2537 vdd.n929 39.2114
R18583 vdd.n2533 vdd.n930 39.2114
R18584 vdd.n2529 vdd.n931 39.2114
R18585 vdd.n2525 vdd.n932 39.2114
R18586 vdd.n2521 vdd.n933 39.2114
R18587 vdd.n2517 vdd.n934 39.2114
R18588 vdd.n2513 vdd.n935 39.2114
R18589 vdd.n2509 vdd.n936 39.2114
R18590 vdd.n2505 vdd.n937 39.2114
R18591 vdd.n2132 vdd.n1080 39.2114
R18592 vdd.n2135 vdd.n2134 39.2114
R18593 vdd.n2140 vdd.n2139 39.2114
R18594 vdd.n2143 vdd.n2142 39.2114
R18595 vdd.n2148 vdd.n2147 39.2114
R18596 vdd.n2151 vdd.n2150 39.2114
R18597 vdd.n2156 vdd.n2155 39.2114
R18598 vdd.n2159 vdd.n2158 39.2114
R18599 vdd.n2164 vdd.n2163 39.2114
R18600 vdd.n2167 vdd.n2166 39.2114
R18601 vdd.n2172 vdd.n2171 39.2114
R18602 vdd.n2175 vdd.n2174 39.2114
R18603 vdd.n2180 vdd.n2179 39.2114
R18604 vdd.n2183 vdd.n2182 39.2114
R18605 vdd.n2188 vdd.n2187 39.2114
R18606 vdd.n2191 vdd.n2190 39.2114
R18607 vdd.n2197 vdd.n2196 39.2114
R18608 vdd.n2502 vdd.n937 39.2114
R18609 vdd.n2506 vdd.n936 39.2114
R18610 vdd.n2510 vdd.n935 39.2114
R18611 vdd.n2514 vdd.n934 39.2114
R18612 vdd.n2518 vdd.n933 39.2114
R18613 vdd.n2522 vdd.n932 39.2114
R18614 vdd.n2526 vdd.n931 39.2114
R18615 vdd.n2530 vdd.n930 39.2114
R18616 vdd.n2534 vdd.n929 39.2114
R18617 vdd.n2538 vdd.n928 39.2114
R18618 vdd.n2542 vdd.n927 39.2114
R18619 vdd.n2546 vdd.n926 39.2114
R18620 vdd.n2550 vdd.n925 39.2114
R18621 vdd.n2554 vdd.n924 39.2114
R18622 vdd.n2558 vdd.n923 39.2114
R18623 vdd.n2562 vdd.n922 39.2114
R18624 vdd.n2566 vdd.n921 39.2114
R18625 vdd.n2133 vdd.n2132 39.2114
R18626 vdd.n2134 vdd.n2130 39.2114
R18627 vdd.n2141 vdd.n2140 39.2114
R18628 vdd.n2142 vdd.n2128 39.2114
R18629 vdd.n2149 vdd.n2148 39.2114
R18630 vdd.n2150 vdd.n2126 39.2114
R18631 vdd.n2157 vdd.n2156 39.2114
R18632 vdd.n2158 vdd.n2124 39.2114
R18633 vdd.n2165 vdd.n2164 39.2114
R18634 vdd.n2166 vdd.n1114 39.2114
R18635 vdd.n2173 vdd.n2172 39.2114
R18636 vdd.n2174 vdd.n1112 39.2114
R18637 vdd.n2181 vdd.n2180 39.2114
R18638 vdd.n2182 vdd.n1110 39.2114
R18639 vdd.n2189 vdd.n2188 39.2114
R18640 vdd.n2190 vdd.n1106 39.2114
R18641 vdd.n2198 vdd.n2197 39.2114
R18642 vdd.n2119 vdd.n2118 37.2369
R18643 vdd.n2035 vdd.n1968 37.2369
R18644 vdd.n2074 vdd.n1928 37.2369
R18645 vdd.n3241 vdd.n724 37.2369
R18646 vdd.n688 vdd.n687 37.2369
R18647 vdd.n3197 vdd.n3196 37.2369
R18648 vdd.n2194 vdd.n1108 30.449
R18649 vdd.n970 vdd.n969 30.449
R18650 vdd.n2319 vdd.n1102 30.449
R18651 vdd.n2579 vdd.n960 30.449
R18652 vdd.n2680 vdd.n2679 30.449
R18653 vdd.n806 vdd.n805 30.449
R18654 vdd.n2807 vdd.n2748 30.449
R18655 vdd.n770 vdd.n769 30.449
R18656 vdd.n2382 vdd.n2381 30.4395
R18657 vdd.n2641 vdd.n958 30.4395
R18658 vdd.n2574 vdd.n961 30.4395
R18659 vdd.n2312 vdd.n2311 30.4395
R18660 vdd.n2814 vdd.n2813 30.4395
R18661 vdd.n3095 vdd.n3092 30.4395
R18662 vdd.n2932 vdd.n2931 30.4395
R18663 vdd.n3156 vdd.n3155 30.4395
R18664 vdd.n3075 vdd.n3074 30.4395
R18665 vdd.n3161 vdd.n771 30.4395
R18666 vdd.n2925 vdd.n2924 30.4395
R18667 vdd.n2936 vdd.n913 30.4395
R18668 vdd.n2386 vdd.n1079 30.4395
R18669 vdd.n2569 vdd.n2568 30.4395
R18670 vdd.n2501 vdd.n2500 30.4395
R18671 vdd.n2201 vdd.n2200 30.4395
R18672 vdd.n1460 vdd.n1226 19.3944
R18673 vdd.n1460 vdd.n1216 19.3944
R18674 vdd.n1472 vdd.n1216 19.3944
R18675 vdd.n1472 vdd.n1214 19.3944
R18676 vdd.n1476 vdd.n1214 19.3944
R18677 vdd.n1476 vdd.n1204 19.3944
R18678 vdd.n1489 vdd.n1204 19.3944
R18679 vdd.n1489 vdd.n1202 19.3944
R18680 vdd.n1493 vdd.n1202 19.3944
R18681 vdd.n1493 vdd.n1194 19.3944
R18682 vdd.n1506 vdd.n1194 19.3944
R18683 vdd.n1506 vdd.n1192 19.3944
R18684 vdd.n1510 vdd.n1192 19.3944
R18685 vdd.n1510 vdd.n1181 19.3944
R18686 vdd.n1522 vdd.n1181 19.3944
R18687 vdd.n1522 vdd.n1179 19.3944
R18688 vdd.n1526 vdd.n1179 19.3944
R18689 vdd.n1526 vdd.n1170 19.3944
R18690 vdd.n1834 vdd.n1170 19.3944
R18691 vdd.n1834 vdd.n1168 19.3944
R18692 vdd.n1838 vdd.n1168 19.3944
R18693 vdd.n1838 vdd.n1159 19.3944
R18694 vdd.n1850 vdd.n1159 19.3944
R18695 vdd.n1850 vdd.n1157 19.3944
R18696 vdd.n1854 vdd.n1157 19.3944
R18697 vdd.n1854 vdd.n1147 19.3944
R18698 vdd.n1867 vdd.n1147 19.3944
R18699 vdd.n1867 vdd.n1145 19.3944
R18700 vdd.n1871 vdd.n1145 19.3944
R18701 vdd.n1871 vdd.n1137 19.3944
R18702 vdd.n1884 vdd.n1137 19.3944
R18703 vdd.n1884 vdd.n1134 19.3944
R18704 vdd.n1890 vdd.n1134 19.3944
R18705 vdd.n1890 vdd.n1135 19.3944
R18706 vdd.n1135 vdd.n1123 19.3944
R18707 vdd.n1379 vdd.n1321 19.3944
R18708 vdd.n1379 vdd.n1378 19.3944
R18709 vdd.n1378 vdd.n1377 19.3944
R18710 vdd.n1377 vdd.n1327 19.3944
R18711 vdd.n1373 vdd.n1327 19.3944
R18712 vdd.n1373 vdd.n1372 19.3944
R18713 vdd.n1372 vdd.n1371 19.3944
R18714 vdd.n1371 vdd.n1333 19.3944
R18715 vdd.n1367 vdd.n1333 19.3944
R18716 vdd.n1367 vdd.n1366 19.3944
R18717 vdd.n1366 vdd.n1365 19.3944
R18718 vdd.n1365 vdd.n1339 19.3944
R18719 vdd.n1361 vdd.n1339 19.3944
R18720 vdd.n1361 vdd.n1360 19.3944
R18721 vdd.n1360 vdd.n1359 19.3944
R18722 vdd.n1359 vdd.n1345 19.3944
R18723 vdd.n1355 vdd.n1345 19.3944
R18724 vdd.n1355 vdd.n1354 19.3944
R18725 vdd.n1354 vdd.n1353 19.3944
R18726 vdd.n1353 vdd.n1351 19.3944
R18727 vdd.n1417 vdd.n1416 19.3944
R18728 vdd.n1416 vdd.n1292 19.3944
R18729 vdd.n1412 vdd.n1292 19.3944
R18730 vdd.n1412 vdd.n1411 19.3944
R18731 vdd.n1411 vdd.n1410 19.3944
R18732 vdd.n1410 vdd.n1298 19.3944
R18733 vdd.n1406 vdd.n1298 19.3944
R18734 vdd.n1406 vdd.n1405 19.3944
R18735 vdd.n1405 vdd.n1404 19.3944
R18736 vdd.n1404 vdd.n1304 19.3944
R18737 vdd.n1400 vdd.n1304 19.3944
R18738 vdd.n1400 vdd.n1399 19.3944
R18739 vdd.n1399 vdd.n1398 19.3944
R18740 vdd.n1398 vdd.n1310 19.3944
R18741 vdd.n1394 vdd.n1310 19.3944
R18742 vdd.n1394 vdd.n1393 19.3944
R18743 vdd.n1393 vdd.n1392 19.3944
R18744 vdd.n1392 vdd.n1316 19.3944
R18745 vdd.n1388 vdd.n1316 19.3944
R18746 vdd.n1388 vdd.n1387 19.3944
R18747 vdd.n1451 vdd.n1450 19.3944
R18748 vdd.n1450 vdd.n1265 19.3944
R18749 vdd.n1446 vdd.n1265 19.3944
R18750 vdd.n1446 vdd.n1445 19.3944
R18751 vdd.n1445 vdd.n1444 19.3944
R18752 vdd.n1444 vdd.n1270 19.3944
R18753 vdd.n1440 vdd.n1270 19.3944
R18754 vdd.n1440 vdd.n1439 19.3944
R18755 vdd.n1439 vdd.n1438 19.3944
R18756 vdd.n1438 vdd.n1276 19.3944
R18757 vdd.n1434 vdd.n1276 19.3944
R18758 vdd.n1434 vdd.n1433 19.3944
R18759 vdd.n1433 vdd.n1432 19.3944
R18760 vdd.n1432 vdd.n1282 19.3944
R18761 vdd.n1428 vdd.n1282 19.3944
R18762 vdd.n1428 vdd.n1427 19.3944
R18763 vdd.n1427 vdd.n1426 19.3944
R18764 vdd.n1426 vdd.n1288 19.3944
R18765 vdd.n2031 vdd.n1966 19.3944
R18766 vdd.n2031 vdd.n1972 19.3944
R18767 vdd.n2026 vdd.n1972 19.3944
R18768 vdd.n2026 vdd.n2025 19.3944
R18769 vdd.n2025 vdd.n2024 19.3944
R18770 vdd.n2024 vdd.n1979 19.3944
R18771 vdd.n2019 vdd.n1979 19.3944
R18772 vdd.n2019 vdd.n2018 19.3944
R18773 vdd.n2018 vdd.n2017 19.3944
R18774 vdd.n2017 vdd.n1986 19.3944
R18775 vdd.n2012 vdd.n1986 19.3944
R18776 vdd.n2012 vdd.n2011 19.3944
R18777 vdd.n2011 vdd.n2010 19.3944
R18778 vdd.n2010 vdd.n1994 19.3944
R18779 vdd.n2005 vdd.n1994 19.3944
R18780 vdd.n2005 vdd.n2004 19.3944
R18781 vdd.n2000 vdd.n1999 19.3944
R18782 vdd.n2120 vdd.n1119 19.3944
R18783 vdd.n2070 vdd.n1926 19.3944
R18784 vdd.n2070 vdd.n1932 19.3944
R18785 vdd.n2065 vdd.n1932 19.3944
R18786 vdd.n2065 vdd.n2064 19.3944
R18787 vdd.n2064 vdd.n2063 19.3944
R18788 vdd.n2063 vdd.n1939 19.3944
R18789 vdd.n2058 vdd.n1939 19.3944
R18790 vdd.n2058 vdd.n2057 19.3944
R18791 vdd.n2057 vdd.n2056 19.3944
R18792 vdd.n2056 vdd.n1946 19.3944
R18793 vdd.n2051 vdd.n1946 19.3944
R18794 vdd.n2051 vdd.n2050 19.3944
R18795 vdd.n2050 vdd.n2049 19.3944
R18796 vdd.n2049 vdd.n1953 19.3944
R18797 vdd.n2044 vdd.n1953 19.3944
R18798 vdd.n2044 vdd.n2043 19.3944
R18799 vdd.n2043 vdd.n2042 19.3944
R18800 vdd.n2042 vdd.n1960 19.3944
R18801 vdd.n2037 vdd.n1960 19.3944
R18802 vdd.n2037 vdd.n2036 19.3944
R18803 vdd.n2108 vdd.n2107 19.3944
R18804 vdd.n2107 vdd.n1898 19.3944
R18805 vdd.n2102 vdd.n2101 19.3944
R18806 vdd.n2097 vdd.n1902 19.3944
R18807 vdd.n2097 vdd.n1904 19.3944
R18808 vdd.n1907 vdd.n1904 19.3944
R18809 vdd.n2090 vdd.n1907 19.3944
R18810 vdd.n2090 vdd.n2089 19.3944
R18811 vdd.n2089 vdd.n2088 19.3944
R18812 vdd.n2088 vdd.n1913 19.3944
R18813 vdd.n2083 vdd.n1913 19.3944
R18814 vdd.n2083 vdd.n2082 19.3944
R18815 vdd.n2082 vdd.n2081 19.3944
R18816 vdd.n2081 vdd.n1920 19.3944
R18817 vdd.n2076 vdd.n1920 19.3944
R18818 vdd.n2076 vdd.n2075 19.3944
R18819 vdd.n1464 vdd.n1222 19.3944
R18820 vdd.n1464 vdd.n1220 19.3944
R18821 vdd.n1468 vdd.n1220 19.3944
R18822 vdd.n1468 vdd.n1210 19.3944
R18823 vdd.n1481 vdd.n1210 19.3944
R18824 vdd.n1481 vdd.n1208 19.3944
R18825 vdd.n1485 vdd.n1208 19.3944
R18826 vdd.n1485 vdd.n1199 19.3944
R18827 vdd.n1498 vdd.n1199 19.3944
R18828 vdd.n1498 vdd.n1197 19.3944
R18829 vdd.n1502 vdd.n1197 19.3944
R18830 vdd.n1502 vdd.n1188 19.3944
R18831 vdd.n1514 vdd.n1188 19.3944
R18832 vdd.n1514 vdd.n1186 19.3944
R18833 vdd.n1518 vdd.n1186 19.3944
R18834 vdd.n1518 vdd.n1176 19.3944
R18835 vdd.n1531 vdd.n1176 19.3944
R18836 vdd.n1531 vdd.n1174 19.3944
R18837 vdd.n1830 vdd.n1174 19.3944
R18838 vdd.n1830 vdd.n1165 19.3944
R18839 vdd.n1842 vdd.n1165 19.3944
R18840 vdd.n1842 vdd.n1163 19.3944
R18841 vdd.n1846 vdd.n1163 19.3944
R18842 vdd.n1846 vdd.n1153 19.3944
R18843 vdd.n1859 vdd.n1153 19.3944
R18844 vdd.n1859 vdd.n1151 19.3944
R18845 vdd.n1863 vdd.n1151 19.3944
R18846 vdd.n1863 vdd.n1142 19.3944
R18847 vdd.n1876 vdd.n1142 19.3944
R18848 vdd.n1876 vdd.n1140 19.3944
R18849 vdd.n1880 vdd.n1140 19.3944
R18850 vdd.n1880 vdd.n1130 19.3944
R18851 vdd.n1894 vdd.n1130 19.3944
R18852 vdd.n1894 vdd.n1128 19.3944
R18853 vdd.n2111 vdd.n1128 19.3944
R18854 vdd.n3329 vdd.n655 19.3944
R18855 vdd.n3333 vdd.n655 19.3944
R18856 vdd.n3333 vdd.n646 19.3944
R18857 vdd.n3345 vdd.n646 19.3944
R18858 vdd.n3345 vdd.n644 19.3944
R18859 vdd.n3349 vdd.n644 19.3944
R18860 vdd.n3349 vdd.n633 19.3944
R18861 vdd.n3361 vdd.n633 19.3944
R18862 vdd.n3361 vdd.n631 19.3944
R18863 vdd.n3365 vdd.n631 19.3944
R18864 vdd.n3365 vdd.n622 19.3944
R18865 vdd.n3378 vdd.n622 19.3944
R18866 vdd.n3378 vdd.n620 19.3944
R18867 vdd.n3385 vdd.n620 19.3944
R18868 vdd.n3385 vdd.n3384 19.3944
R18869 vdd.n3384 vdd.n610 19.3944
R18870 vdd.n3398 vdd.n610 19.3944
R18871 vdd.n3399 vdd.n3398 19.3944
R18872 vdd.n3400 vdd.n3399 19.3944
R18873 vdd.n3400 vdd.n608 19.3944
R18874 vdd.n3405 vdd.n608 19.3944
R18875 vdd.n3406 vdd.n3405 19.3944
R18876 vdd.n3407 vdd.n3406 19.3944
R18877 vdd.n3407 vdd.n606 19.3944
R18878 vdd.n3412 vdd.n606 19.3944
R18879 vdd.n3413 vdd.n3412 19.3944
R18880 vdd.n3414 vdd.n3413 19.3944
R18881 vdd.n3414 vdd.n604 19.3944
R18882 vdd.n3420 vdd.n604 19.3944
R18883 vdd.n3421 vdd.n3420 19.3944
R18884 vdd.n3422 vdd.n3421 19.3944
R18885 vdd.n3422 vdd.n602 19.3944
R18886 vdd.n3427 vdd.n602 19.3944
R18887 vdd.n3428 vdd.n3427 19.3944
R18888 vdd.n3429 vdd.n3428 19.3944
R18889 vdd.n550 vdd.n417 19.3944
R18890 vdd.n556 vdd.n417 19.3944
R18891 vdd.n557 vdd.n556 19.3944
R18892 vdd.n560 vdd.n557 19.3944
R18893 vdd.n560 vdd.n415 19.3944
R18894 vdd.n566 vdd.n415 19.3944
R18895 vdd.n567 vdd.n566 19.3944
R18896 vdd.n570 vdd.n567 19.3944
R18897 vdd.n570 vdd.n413 19.3944
R18898 vdd.n576 vdd.n413 19.3944
R18899 vdd.n577 vdd.n576 19.3944
R18900 vdd.n580 vdd.n577 19.3944
R18901 vdd.n580 vdd.n411 19.3944
R18902 vdd.n586 vdd.n411 19.3944
R18903 vdd.n587 vdd.n586 19.3944
R18904 vdd.n590 vdd.n587 19.3944
R18905 vdd.n590 vdd.n409 19.3944
R18906 vdd.n596 vdd.n409 19.3944
R18907 vdd.n598 vdd.n596 19.3944
R18908 vdd.n599 vdd.n598 19.3944
R18909 vdd.n497 vdd.n496 19.3944
R18910 vdd.n500 vdd.n497 19.3944
R18911 vdd.n500 vdd.n429 19.3944
R18912 vdd.n506 vdd.n429 19.3944
R18913 vdd.n507 vdd.n506 19.3944
R18914 vdd.n510 vdd.n507 19.3944
R18915 vdd.n510 vdd.n427 19.3944
R18916 vdd.n516 vdd.n427 19.3944
R18917 vdd.n517 vdd.n516 19.3944
R18918 vdd.n520 vdd.n517 19.3944
R18919 vdd.n520 vdd.n425 19.3944
R18920 vdd.n526 vdd.n425 19.3944
R18921 vdd.n527 vdd.n526 19.3944
R18922 vdd.n530 vdd.n527 19.3944
R18923 vdd.n530 vdd.n423 19.3944
R18924 vdd.n536 vdd.n423 19.3944
R18925 vdd.n537 vdd.n536 19.3944
R18926 vdd.n540 vdd.n537 19.3944
R18927 vdd.n540 vdd.n421 19.3944
R18928 vdd.n546 vdd.n421 19.3944
R18929 vdd.n447 vdd.n446 19.3944
R18930 vdd.n450 vdd.n447 19.3944
R18931 vdd.n450 vdd.n441 19.3944
R18932 vdd.n456 vdd.n441 19.3944
R18933 vdd.n457 vdd.n456 19.3944
R18934 vdd.n460 vdd.n457 19.3944
R18935 vdd.n460 vdd.n439 19.3944
R18936 vdd.n466 vdd.n439 19.3944
R18937 vdd.n467 vdd.n466 19.3944
R18938 vdd.n470 vdd.n467 19.3944
R18939 vdd.n470 vdd.n437 19.3944
R18940 vdd.n476 vdd.n437 19.3944
R18941 vdd.n477 vdd.n476 19.3944
R18942 vdd.n480 vdd.n477 19.3944
R18943 vdd.n480 vdd.n435 19.3944
R18944 vdd.n486 vdd.n435 19.3944
R18945 vdd.n487 vdd.n486 19.3944
R18946 vdd.n490 vdd.n487 19.3944
R18947 vdd.n3325 vdd.n652 19.3944
R18948 vdd.n3337 vdd.n652 19.3944
R18949 vdd.n3337 vdd.n650 19.3944
R18950 vdd.n3341 vdd.n650 19.3944
R18951 vdd.n3341 vdd.n640 19.3944
R18952 vdd.n3353 vdd.n640 19.3944
R18953 vdd.n3353 vdd.n638 19.3944
R18954 vdd.n3357 vdd.n638 19.3944
R18955 vdd.n3357 vdd.n628 19.3944
R18956 vdd.n3370 vdd.n628 19.3944
R18957 vdd.n3370 vdd.n626 19.3944
R18958 vdd.n3374 vdd.n626 19.3944
R18959 vdd.n3374 vdd.n617 19.3944
R18960 vdd.n3389 vdd.n617 19.3944
R18961 vdd.n3389 vdd.n615 19.3944
R18962 vdd.n3393 vdd.n615 19.3944
R18963 vdd.n3393 vdd.n324 19.3944
R18964 vdd.n3471 vdd.n324 19.3944
R18965 vdd.n3471 vdd.n325 19.3944
R18966 vdd.n3465 vdd.n325 19.3944
R18967 vdd.n3465 vdd.n3464 19.3944
R18968 vdd.n3464 vdd.n3463 19.3944
R18969 vdd.n3463 vdd.n337 19.3944
R18970 vdd.n3457 vdd.n337 19.3944
R18971 vdd.n3457 vdd.n3456 19.3944
R18972 vdd.n3456 vdd.n3455 19.3944
R18973 vdd.n3455 vdd.n347 19.3944
R18974 vdd.n3449 vdd.n347 19.3944
R18975 vdd.n3449 vdd.n3448 19.3944
R18976 vdd.n3448 vdd.n3447 19.3944
R18977 vdd.n3447 vdd.n358 19.3944
R18978 vdd.n3441 vdd.n358 19.3944
R18979 vdd.n3441 vdd.n3440 19.3944
R18980 vdd.n3440 vdd.n3439 19.3944
R18981 vdd.n3439 vdd.n369 19.3944
R18982 vdd.n3282 vdd.n3281 19.3944
R18983 vdd.n3281 vdd.n3280 19.3944
R18984 vdd.n3280 vdd.n694 19.3944
R18985 vdd.n3274 vdd.n694 19.3944
R18986 vdd.n3274 vdd.n3273 19.3944
R18987 vdd.n3273 vdd.n3272 19.3944
R18988 vdd.n3272 vdd.n700 19.3944
R18989 vdd.n3266 vdd.n700 19.3944
R18990 vdd.n3266 vdd.n3265 19.3944
R18991 vdd.n3265 vdd.n3264 19.3944
R18992 vdd.n3264 vdd.n706 19.3944
R18993 vdd.n3258 vdd.n706 19.3944
R18994 vdd.n3258 vdd.n3257 19.3944
R18995 vdd.n3257 vdd.n3256 19.3944
R18996 vdd.n3256 vdd.n712 19.3944
R18997 vdd.n3250 vdd.n712 19.3944
R18998 vdd.n3250 vdd.n3249 19.3944
R18999 vdd.n3249 vdd.n3248 19.3944
R19000 vdd.n3248 vdd.n718 19.3944
R19001 vdd.n3242 vdd.n718 19.3944
R19002 vdd.n3322 vdd.n3321 19.3944
R19003 vdd.n3321 vdd.n662 19.3944
R19004 vdd.n3316 vdd.n3315 19.3944
R19005 vdd.n3312 vdd.n3311 19.3944
R19006 vdd.n3311 vdd.n668 19.3944
R19007 vdd.n3306 vdd.n668 19.3944
R19008 vdd.n3306 vdd.n3305 19.3944
R19009 vdd.n3305 vdd.n3304 19.3944
R19010 vdd.n3304 vdd.n674 19.3944
R19011 vdd.n3298 vdd.n674 19.3944
R19012 vdd.n3298 vdd.n3297 19.3944
R19013 vdd.n3297 vdd.n3296 19.3944
R19014 vdd.n3296 vdd.n680 19.3944
R19015 vdd.n3290 vdd.n680 19.3944
R19016 vdd.n3290 vdd.n3289 19.3944
R19017 vdd.n3289 vdd.n3288 19.3944
R19018 vdd.n3237 vdd.n722 19.3944
R19019 vdd.n3237 vdd.n726 19.3944
R19020 vdd.n3232 vdd.n726 19.3944
R19021 vdd.n3232 vdd.n3231 19.3944
R19022 vdd.n3231 vdd.n732 19.3944
R19023 vdd.n3226 vdd.n732 19.3944
R19024 vdd.n3226 vdd.n3225 19.3944
R19025 vdd.n3225 vdd.n3224 19.3944
R19026 vdd.n3224 vdd.n738 19.3944
R19027 vdd.n3218 vdd.n738 19.3944
R19028 vdd.n3218 vdd.n3217 19.3944
R19029 vdd.n3217 vdd.n3216 19.3944
R19030 vdd.n3216 vdd.n744 19.3944
R19031 vdd.n3210 vdd.n744 19.3944
R19032 vdd.n3210 vdd.n3209 19.3944
R19033 vdd.n3209 vdd.n3208 19.3944
R19034 vdd.n3204 vdd.n3203 19.3944
R19035 vdd.n3200 vdd.n3199 19.3944
R19036 vdd.n1386 vdd.n1321 19.0066
R19037 vdd.n2035 vdd.n1966 19.0066
R19038 vdd.n550 vdd.n547 19.0066
R19039 vdd.n3241 vdd.n722 19.0066
R19040 vdd.n1454 vdd.n1224 18.5924
R19041 vdd.n2113 vdd.n1125 18.5924
R19042 vdd.n3327 vdd.n658 18.5924
R19043 vdd.n3436 vdd.n3435 18.5924
R19044 vdd.n1108 vdd.n1107 16.0975
R19045 vdd.n969 vdd.n968 16.0975
R19046 vdd.n1229 vdd.n1228 16.0975
R19047 vdd.n1385 vdd.n1384 16.0975
R19048 vdd.n1421 vdd.n1420 16.0975
R19049 vdd.n2118 vdd.n2117 16.0975
R19050 vdd.n1968 vdd.n1967 16.0975
R19051 vdd.n1928 vdd.n1927 16.0975
R19052 vdd.n1102 vdd.n1101 16.0975
R19053 vdd.n960 vdd.n959 16.0975
R19054 vdd.n2679 vdd.n2678 16.0975
R19055 vdd.n406 vdd.n405 16.0975
R19056 vdd.n420 vdd.n419 16.0975
R19057 vdd.n432 vdd.n431 16.0975
R19058 vdd.n724 vdd.n723 16.0975
R19059 vdd.n687 vdd.n686 16.0975
R19060 vdd.n805 vdd.n804 16.0975
R19061 vdd.n2748 vdd.n2747 16.0975
R19062 vdd.n3196 vdd.n3195 16.0975
R19063 vdd.n769 vdd.n768 16.0975
R19064 vdd.t233 vdd.n2643 15.4182
R19065 vdd.n2927 vdd.t250 15.4182
R19066 vdd.n28 vdd.n27 15.0023
R19067 vdd.n2384 vdd.n1081 13.6043
R19068 vdd.n3158 vdd.n756 13.6043
R19069 vdd.n316 vdd.n281 13.1884
R19070 vdd.n261 vdd.n226 13.1884
R19071 vdd.n218 vdd.n183 13.1884
R19072 vdd.n163 vdd.n128 13.1884
R19073 vdd.n121 vdd.n86 13.1884
R19074 vdd.n66 vdd.n31 13.1884
R19075 vdd.n1765 vdd.n1730 13.1884
R19076 vdd.n1820 vdd.n1785 13.1884
R19077 vdd.n1667 vdd.n1632 13.1884
R19078 vdd.n1722 vdd.n1687 13.1884
R19079 vdd.n1570 vdd.n1535 13.1884
R19080 vdd.n1625 vdd.n1590 13.1884
R19081 vdd.n1422 vdd.n1417 12.9944
R19082 vdd.n1422 vdd.n1288 12.9944
R19083 vdd.n2074 vdd.n1926 12.9944
R19084 vdd.n2075 vdd.n2074 12.9944
R19085 vdd.n496 vdd.n433 12.9944
R19086 vdd.n490 vdd.n433 12.9944
R19087 vdd.n3282 vdd.n688 12.9944
R19088 vdd.n3288 vdd.n688 12.9944
R19089 vdd.n317 vdd.n279 12.8005
R19090 vdd.n312 vdd.n283 12.8005
R19091 vdd.n262 vdd.n224 12.8005
R19092 vdd.n257 vdd.n228 12.8005
R19093 vdd.n219 vdd.n181 12.8005
R19094 vdd.n214 vdd.n185 12.8005
R19095 vdd.n164 vdd.n126 12.8005
R19096 vdd.n159 vdd.n130 12.8005
R19097 vdd.n122 vdd.n84 12.8005
R19098 vdd.n117 vdd.n88 12.8005
R19099 vdd.n67 vdd.n29 12.8005
R19100 vdd.n62 vdd.n33 12.8005
R19101 vdd.n1766 vdd.n1728 12.8005
R19102 vdd.n1761 vdd.n1732 12.8005
R19103 vdd.n1821 vdd.n1783 12.8005
R19104 vdd.n1816 vdd.n1787 12.8005
R19105 vdd.n1668 vdd.n1630 12.8005
R19106 vdd.n1663 vdd.n1634 12.8005
R19107 vdd.n1723 vdd.n1685 12.8005
R19108 vdd.n1718 vdd.n1689 12.8005
R19109 vdd.n1571 vdd.n1533 12.8005
R19110 vdd.n1566 vdd.n1537 12.8005
R19111 vdd.n1626 vdd.n1588 12.8005
R19112 vdd.n1621 vdd.n1592 12.8005
R19113 vdd.n311 vdd.n284 12.0247
R19114 vdd.n256 vdd.n229 12.0247
R19115 vdd.n213 vdd.n186 12.0247
R19116 vdd.n158 vdd.n131 12.0247
R19117 vdd.n116 vdd.n89 12.0247
R19118 vdd.n61 vdd.n34 12.0247
R19119 vdd.n1760 vdd.n1733 12.0247
R19120 vdd.n1815 vdd.n1788 12.0247
R19121 vdd.n1662 vdd.n1635 12.0247
R19122 vdd.n1717 vdd.n1690 12.0247
R19123 vdd.n1565 vdd.n1538 12.0247
R19124 vdd.n1620 vdd.n1593 12.0247
R19125 vdd.n1462 vdd.n1224 11.337
R19126 vdd.n1470 vdd.n1218 11.337
R19127 vdd.n1470 vdd.n1212 11.337
R19128 vdd.n1479 vdd.n1212 11.337
R19129 vdd.n1487 vdd.n1206 11.337
R19130 vdd.n1496 vdd.n1495 11.337
R19131 vdd.n1512 vdd.n1190 11.337
R19132 vdd.n1520 vdd.n1183 11.337
R19133 vdd.n1529 vdd.n1528 11.337
R19134 vdd.n1832 vdd.n1172 11.337
R19135 vdd.n1848 vdd.n1161 11.337
R19136 vdd.n1857 vdd.n1155 11.337
R19137 vdd.n1865 vdd.n1149 11.337
R19138 vdd.n1874 vdd.n1873 11.337
R19139 vdd.n1882 vdd.n1132 11.337
R19140 vdd.n1892 vdd.n1132 11.337
R19141 vdd.n2113 vdd.n1124 11.337
R19142 vdd.n3327 vdd.n659 11.337
R19143 vdd.n3335 vdd.n648 11.337
R19144 vdd.n3343 vdd.n648 11.337
R19145 vdd.n3351 vdd.n642 11.337
R19146 vdd.n3359 vdd.n635 11.337
R19147 vdd.n3368 vdd.n3367 11.337
R19148 vdd.n3376 vdd.n624 11.337
R19149 vdd.n3395 vdd.n613 11.337
R19150 vdd.n3469 vdd.n328 11.337
R19151 vdd.n3467 vdd.n332 11.337
R19152 vdd.n3461 vdd.n3460 11.337
R19153 vdd.n3453 vdd.n349 11.337
R19154 vdd.n3452 vdd.n3451 11.337
R19155 vdd.n3445 vdd.n3444 11.337
R19156 vdd.n3444 vdd.n3443 11.337
R19157 vdd.n3443 vdd.n363 11.337
R19158 vdd.n3437 vdd.n3436 11.337
R19159 vdd.n308 vdd.n307 11.249
R19160 vdd.n253 vdd.n252 11.249
R19161 vdd.n210 vdd.n209 11.249
R19162 vdd.n155 vdd.n154 11.249
R19163 vdd.n113 vdd.n112 11.249
R19164 vdd.n58 vdd.n57 11.249
R19165 vdd.n1757 vdd.n1756 11.249
R19166 vdd.n1812 vdd.n1811 11.249
R19167 vdd.n1659 vdd.n1658 11.249
R19168 vdd.n1714 vdd.n1713 11.249
R19169 vdd.n1562 vdd.n1561 11.249
R19170 vdd.n1617 vdd.n1616 11.249
R19171 vdd.n1882 vdd.t95 10.7702
R19172 vdd.n3343 vdd.t63 10.7702
R19173 vdd.n293 vdd.n292 10.7238
R19174 vdd.n238 vdd.n237 10.7238
R19175 vdd.n195 vdd.n194 10.7238
R19176 vdd.n140 vdd.n139 10.7238
R19177 vdd.n98 vdd.n97 10.7238
R19178 vdd.n43 vdd.n42 10.7238
R19179 vdd.n1742 vdd.n1741 10.7238
R19180 vdd.n1797 vdd.n1796 10.7238
R19181 vdd.n1644 vdd.n1643 10.7238
R19182 vdd.n1699 vdd.n1698 10.7238
R19183 vdd.n1547 vdd.n1546 10.7238
R19184 vdd.n1602 vdd.n1601 10.7238
R19185 vdd.n2382 vdd.n1073 10.6151
R19186 vdd.n2392 vdd.n1073 10.6151
R19187 vdd.n2393 vdd.n2392 10.6151
R19188 vdd.n2394 vdd.n2393 10.6151
R19189 vdd.n2394 vdd.n1061 10.6151
R19190 vdd.n2404 vdd.n1061 10.6151
R19191 vdd.n2405 vdd.n2404 10.6151
R19192 vdd.n2406 vdd.n2405 10.6151
R19193 vdd.n2406 vdd.n1049 10.6151
R19194 vdd.n2416 vdd.n1049 10.6151
R19195 vdd.n2417 vdd.n2416 10.6151
R19196 vdd.n2418 vdd.n2417 10.6151
R19197 vdd.n2418 vdd.n1036 10.6151
R19198 vdd.n2428 vdd.n1036 10.6151
R19199 vdd.n2429 vdd.n2428 10.6151
R19200 vdd.n2430 vdd.n2429 10.6151
R19201 vdd.n2430 vdd.n1024 10.6151
R19202 vdd.n2441 vdd.n1024 10.6151
R19203 vdd.n2442 vdd.n2441 10.6151
R19204 vdd.n2443 vdd.n2442 10.6151
R19205 vdd.n2443 vdd.n1012 10.6151
R19206 vdd.n2453 vdd.n1012 10.6151
R19207 vdd.n2454 vdd.n2453 10.6151
R19208 vdd.n2455 vdd.n2454 10.6151
R19209 vdd.n2455 vdd.n1000 10.6151
R19210 vdd.n2465 vdd.n1000 10.6151
R19211 vdd.n2466 vdd.n2465 10.6151
R19212 vdd.n2467 vdd.n2466 10.6151
R19213 vdd.n2467 vdd.n990 10.6151
R19214 vdd.n2477 vdd.n990 10.6151
R19215 vdd.n2478 vdd.n2477 10.6151
R19216 vdd.n2479 vdd.n2478 10.6151
R19217 vdd.n2479 vdd.n977 10.6151
R19218 vdd.n2491 vdd.n977 10.6151
R19219 vdd.n2492 vdd.n2491 10.6151
R19220 vdd.n2494 vdd.n2492 10.6151
R19221 vdd.n2494 vdd.n2493 10.6151
R19222 vdd.n2493 vdd.n958 10.6151
R19223 vdd.n2641 vdd.n2640 10.6151
R19224 vdd.n2640 vdd.n2639 10.6151
R19225 vdd.n2639 vdd.n2636 10.6151
R19226 vdd.n2636 vdd.n2635 10.6151
R19227 vdd.n2635 vdd.n2632 10.6151
R19228 vdd.n2632 vdd.n2631 10.6151
R19229 vdd.n2631 vdd.n2628 10.6151
R19230 vdd.n2628 vdd.n2627 10.6151
R19231 vdd.n2627 vdd.n2624 10.6151
R19232 vdd.n2624 vdd.n2623 10.6151
R19233 vdd.n2623 vdd.n2620 10.6151
R19234 vdd.n2620 vdd.n2619 10.6151
R19235 vdd.n2619 vdd.n2616 10.6151
R19236 vdd.n2616 vdd.n2615 10.6151
R19237 vdd.n2615 vdd.n2612 10.6151
R19238 vdd.n2612 vdd.n2611 10.6151
R19239 vdd.n2611 vdd.n2608 10.6151
R19240 vdd.n2608 vdd.n2607 10.6151
R19241 vdd.n2607 vdd.n2604 10.6151
R19242 vdd.n2604 vdd.n2603 10.6151
R19243 vdd.n2603 vdd.n2600 10.6151
R19244 vdd.n2600 vdd.n2599 10.6151
R19245 vdd.n2599 vdd.n2596 10.6151
R19246 vdd.n2596 vdd.n2595 10.6151
R19247 vdd.n2595 vdd.n2592 10.6151
R19248 vdd.n2592 vdd.n2591 10.6151
R19249 vdd.n2591 vdd.n2588 10.6151
R19250 vdd.n2588 vdd.n2587 10.6151
R19251 vdd.n2587 vdd.n2584 10.6151
R19252 vdd.n2584 vdd.n2583 10.6151
R19253 vdd.n2583 vdd.n2580 10.6151
R19254 vdd.n2578 vdd.n2575 10.6151
R19255 vdd.n2575 vdd.n2574 10.6151
R19256 vdd.n2311 vdd.n2310 10.6151
R19257 vdd.n2310 vdd.n2308 10.6151
R19258 vdd.n2308 vdd.n2307 10.6151
R19259 vdd.n2307 vdd.n2305 10.6151
R19260 vdd.n2305 vdd.n2304 10.6151
R19261 vdd.n2304 vdd.n2302 10.6151
R19262 vdd.n2302 vdd.n2301 10.6151
R19263 vdd.n2301 vdd.n2299 10.6151
R19264 vdd.n2299 vdd.n2298 10.6151
R19265 vdd.n2298 vdd.n2296 10.6151
R19266 vdd.n2296 vdd.n2295 10.6151
R19267 vdd.n2295 vdd.n2293 10.6151
R19268 vdd.n2293 vdd.n2292 10.6151
R19269 vdd.n2292 vdd.n2290 10.6151
R19270 vdd.n2290 vdd.n2289 10.6151
R19271 vdd.n2289 vdd.n2287 10.6151
R19272 vdd.n2287 vdd.n2286 10.6151
R19273 vdd.n2286 vdd.n2284 10.6151
R19274 vdd.n2284 vdd.n2283 10.6151
R19275 vdd.n2283 vdd.n2281 10.6151
R19276 vdd.n2281 vdd.n2280 10.6151
R19277 vdd.n2280 vdd.n2278 10.6151
R19278 vdd.n2278 vdd.n2277 10.6151
R19279 vdd.n2277 vdd.n1104 10.6151
R19280 vdd.n2244 vdd.n1104 10.6151
R19281 vdd.n2245 vdd.n2244 10.6151
R19282 vdd.n2247 vdd.n2245 10.6151
R19283 vdd.n2248 vdd.n2247 10.6151
R19284 vdd.n2261 vdd.n2248 10.6151
R19285 vdd.n2261 vdd.n2260 10.6151
R19286 vdd.n2260 vdd.n2259 10.6151
R19287 vdd.n2259 vdd.n2257 10.6151
R19288 vdd.n2257 vdd.n2256 10.6151
R19289 vdd.n2256 vdd.n2254 10.6151
R19290 vdd.n2254 vdd.n2253 10.6151
R19291 vdd.n2253 vdd.n2250 10.6151
R19292 vdd.n2250 vdd.n2249 10.6151
R19293 vdd.n2249 vdd.n961 10.6151
R19294 vdd.n2381 vdd.n2380 10.6151
R19295 vdd.n2380 vdd.n1085 10.6151
R19296 vdd.n2375 vdd.n1085 10.6151
R19297 vdd.n2375 vdd.n2374 10.6151
R19298 vdd.n2374 vdd.n1087 10.6151
R19299 vdd.n2369 vdd.n1087 10.6151
R19300 vdd.n2369 vdd.n2368 10.6151
R19301 vdd.n2368 vdd.n2367 10.6151
R19302 vdd.n2367 vdd.n1089 10.6151
R19303 vdd.n2361 vdd.n1089 10.6151
R19304 vdd.n2361 vdd.n2360 10.6151
R19305 vdd.n2360 vdd.n2359 10.6151
R19306 vdd.n2359 vdd.n1091 10.6151
R19307 vdd.n2353 vdd.n1091 10.6151
R19308 vdd.n2353 vdd.n2352 10.6151
R19309 vdd.n2352 vdd.n2351 10.6151
R19310 vdd.n2351 vdd.n1093 10.6151
R19311 vdd.n2345 vdd.n1093 10.6151
R19312 vdd.n2345 vdd.n2344 10.6151
R19313 vdd.n2344 vdd.n2343 10.6151
R19314 vdd.n2343 vdd.n1095 10.6151
R19315 vdd.n2337 vdd.n1095 10.6151
R19316 vdd.n2337 vdd.n2336 10.6151
R19317 vdd.n2336 vdd.n2335 10.6151
R19318 vdd.n2335 vdd.n1097 10.6151
R19319 vdd.n2329 vdd.n1097 10.6151
R19320 vdd.n2329 vdd.n2328 10.6151
R19321 vdd.n2328 vdd.n2327 10.6151
R19322 vdd.n2327 vdd.n1099 10.6151
R19323 vdd.n2321 vdd.n1099 10.6151
R19324 vdd.n2321 vdd.n2320 10.6151
R19325 vdd.n2318 vdd.n1103 10.6151
R19326 vdd.n2312 vdd.n1103 10.6151
R19327 vdd.n2816 vdd.n2814 10.6151
R19328 vdd.n2817 vdd.n2816 10.6151
R19329 vdd.n2916 vdd.n2817 10.6151
R19330 vdd.n2916 vdd.n2915 10.6151
R19331 vdd.n2915 vdd.n2914 10.6151
R19332 vdd.n2914 vdd.n2912 10.6151
R19333 vdd.n2912 vdd.n2911 10.6151
R19334 vdd.n2911 vdd.n2909 10.6151
R19335 vdd.n2909 vdd.n2908 10.6151
R19336 vdd.n2908 vdd.n2818 10.6151
R19337 vdd.n2858 vdd.n2818 10.6151
R19338 vdd.n2859 vdd.n2858 10.6151
R19339 vdd.n2861 vdd.n2859 10.6151
R19340 vdd.n2862 vdd.n2861 10.6151
R19341 vdd.n2892 vdd.n2862 10.6151
R19342 vdd.n2892 vdd.n2891 10.6151
R19343 vdd.n2891 vdd.n2890 10.6151
R19344 vdd.n2890 vdd.n2888 10.6151
R19345 vdd.n2888 vdd.n2887 10.6151
R19346 vdd.n2887 vdd.n2885 10.6151
R19347 vdd.n2885 vdd.n2884 10.6151
R19348 vdd.n2884 vdd.n2882 10.6151
R19349 vdd.n2882 vdd.n2881 10.6151
R19350 vdd.n2881 vdd.n2879 10.6151
R19351 vdd.n2879 vdd.n2878 10.6151
R19352 vdd.n2878 vdd.n2876 10.6151
R19353 vdd.n2876 vdd.n2875 10.6151
R19354 vdd.n2875 vdd.n2873 10.6151
R19355 vdd.n2873 vdd.n2872 10.6151
R19356 vdd.n2872 vdd.n2870 10.6151
R19357 vdd.n2870 vdd.n2869 10.6151
R19358 vdd.n2869 vdd.n2867 10.6151
R19359 vdd.n2867 vdd.n2866 10.6151
R19360 vdd.n2866 vdd.n2864 10.6151
R19361 vdd.n2864 vdd.n2863 10.6151
R19362 vdd.n2863 vdd.n807 10.6151
R19363 vdd.n3091 vdd.n807 10.6151
R19364 vdd.n3092 vdd.n3091 10.6151
R19365 vdd.n2931 vdd.n2930 10.6151
R19366 vdd.n2930 vdd.n919 10.6151
R19367 vdd.n2750 vdd.n919 10.6151
R19368 vdd.n2751 vdd.n2750 10.6151
R19369 vdd.n2754 vdd.n2751 10.6151
R19370 vdd.n2755 vdd.n2754 10.6151
R19371 vdd.n2758 vdd.n2755 10.6151
R19372 vdd.n2759 vdd.n2758 10.6151
R19373 vdd.n2762 vdd.n2759 10.6151
R19374 vdd.n2763 vdd.n2762 10.6151
R19375 vdd.n2766 vdd.n2763 10.6151
R19376 vdd.n2767 vdd.n2766 10.6151
R19377 vdd.n2770 vdd.n2767 10.6151
R19378 vdd.n2771 vdd.n2770 10.6151
R19379 vdd.n2774 vdd.n2771 10.6151
R19380 vdd.n2775 vdd.n2774 10.6151
R19381 vdd.n2778 vdd.n2775 10.6151
R19382 vdd.n2779 vdd.n2778 10.6151
R19383 vdd.n2782 vdd.n2779 10.6151
R19384 vdd.n2783 vdd.n2782 10.6151
R19385 vdd.n2786 vdd.n2783 10.6151
R19386 vdd.n2787 vdd.n2786 10.6151
R19387 vdd.n2790 vdd.n2787 10.6151
R19388 vdd.n2791 vdd.n2790 10.6151
R19389 vdd.n2794 vdd.n2791 10.6151
R19390 vdd.n2795 vdd.n2794 10.6151
R19391 vdd.n2798 vdd.n2795 10.6151
R19392 vdd.n2799 vdd.n2798 10.6151
R19393 vdd.n2802 vdd.n2799 10.6151
R19394 vdd.n2803 vdd.n2802 10.6151
R19395 vdd.n2806 vdd.n2803 10.6151
R19396 vdd.n2811 vdd.n2808 10.6151
R19397 vdd.n2813 vdd.n2811 10.6151
R19398 vdd.n2932 vdd.n908 10.6151
R19399 vdd.n2942 vdd.n908 10.6151
R19400 vdd.n2943 vdd.n2942 10.6151
R19401 vdd.n2944 vdd.n2943 10.6151
R19402 vdd.n2944 vdd.n896 10.6151
R19403 vdd.n2954 vdd.n896 10.6151
R19404 vdd.n2955 vdd.n2954 10.6151
R19405 vdd.n2956 vdd.n2955 10.6151
R19406 vdd.n2956 vdd.n886 10.6151
R19407 vdd.n2966 vdd.n886 10.6151
R19408 vdd.n2967 vdd.n2966 10.6151
R19409 vdd.n2968 vdd.n2967 10.6151
R19410 vdd.n2968 vdd.n874 10.6151
R19411 vdd.n2978 vdd.n874 10.6151
R19412 vdd.n2979 vdd.n2978 10.6151
R19413 vdd.n2980 vdd.n2979 10.6151
R19414 vdd.n2980 vdd.n863 10.6151
R19415 vdd.n2990 vdd.n863 10.6151
R19416 vdd.n2991 vdd.n2990 10.6151
R19417 vdd.n2992 vdd.n2991 10.6151
R19418 vdd.n2992 vdd.n850 10.6151
R19419 vdd.n3003 vdd.n850 10.6151
R19420 vdd.n3004 vdd.n3003 10.6151
R19421 vdd.n3005 vdd.n3004 10.6151
R19422 vdd.n3005 vdd.n837 10.6151
R19423 vdd.n3015 vdd.n837 10.6151
R19424 vdd.n3016 vdd.n3015 10.6151
R19425 vdd.n3017 vdd.n3016 10.6151
R19426 vdd.n3017 vdd.n826 10.6151
R19427 vdd.n3027 vdd.n826 10.6151
R19428 vdd.n3028 vdd.n3027 10.6151
R19429 vdd.n3029 vdd.n3028 10.6151
R19430 vdd.n3029 vdd.n812 10.6151
R19431 vdd.n3084 vdd.n812 10.6151
R19432 vdd.n3085 vdd.n3084 10.6151
R19433 vdd.n3086 vdd.n3085 10.6151
R19434 vdd.n3086 vdd.n779 10.6151
R19435 vdd.n3156 vdd.n779 10.6151
R19436 vdd.n3155 vdd.n3154 10.6151
R19437 vdd.n3154 vdd.n780 10.6151
R19438 vdd.n781 vdd.n780 10.6151
R19439 vdd.n3147 vdd.n781 10.6151
R19440 vdd.n3147 vdd.n3146 10.6151
R19441 vdd.n3146 vdd.n3145 10.6151
R19442 vdd.n3145 vdd.n783 10.6151
R19443 vdd.n3140 vdd.n783 10.6151
R19444 vdd.n3140 vdd.n3139 10.6151
R19445 vdd.n3139 vdd.n3138 10.6151
R19446 vdd.n3138 vdd.n786 10.6151
R19447 vdd.n3133 vdd.n786 10.6151
R19448 vdd.n3133 vdd.n3132 10.6151
R19449 vdd.n3132 vdd.n3131 10.6151
R19450 vdd.n3131 vdd.n789 10.6151
R19451 vdd.n3126 vdd.n789 10.6151
R19452 vdd.n3126 vdd.n3125 10.6151
R19453 vdd.n3125 vdd.n3123 10.6151
R19454 vdd.n3123 vdd.n792 10.6151
R19455 vdd.n3118 vdd.n792 10.6151
R19456 vdd.n3118 vdd.n3117 10.6151
R19457 vdd.n3117 vdd.n3116 10.6151
R19458 vdd.n3116 vdd.n795 10.6151
R19459 vdd.n3111 vdd.n795 10.6151
R19460 vdd.n3111 vdd.n3110 10.6151
R19461 vdd.n3110 vdd.n3109 10.6151
R19462 vdd.n3109 vdd.n798 10.6151
R19463 vdd.n3104 vdd.n798 10.6151
R19464 vdd.n3104 vdd.n3103 10.6151
R19465 vdd.n3103 vdd.n3102 10.6151
R19466 vdd.n3102 vdd.n801 10.6151
R19467 vdd.n3097 vdd.n3096 10.6151
R19468 vdd.n3096 vdd.n3095 10.6151
R19469 vdd.n3074 vdd.n3035 10.6151
R19470 vdd.n3069 vdd.n3035 10.6151
R19471 vdd.n3069 vdd.n3068 10.6151
R19472 vdd.n3068 vdd.n3067 10.6151
R19473 vdd.n3067 vdd.n3037 10.6151
R19474 vdd.n3062 vdd.n3037 10.6151
R19475 vdd.n3062 vdd.n3061 10.6151
R19476 vdd.n3061 vdd.n3060 10.6151
R19477 vdd.n3060 vdd.n3040 10.6151
R19478 vdd.n3055 vdd.n3040 10.6151
R19479 vdd.n3055 vdd.n3054 10.6151
R19480 vdd.n3054 vdd.n3053 10.6151
R19481 vdd.n3053 vdd.n3043 10.6151
R19482 vdd.n3048 vdd.n3043 10.6151
R19483 vdd.n3048 vdd.n3047 10.6151
R19484 vdd.n3047 vdd.n753 10.6151
R19485 vdd.n3191 vdd.n753 10.6151
R19486 vdd.n3191 vdd.n754 10.6151
R19487 vdd.n757 vdd.n754 10.6151
R19488 vdd.n3184 vdd.n757 10.6151
R19489 vdd.n3184 vdd.n3183 10.6151
R19490 vdd.n3183 vdd.n3182 10.6151
R19491 vdd.n3182 vdd.n759 10.6151
R19492 vdd.n3177 vdd.n759 10.6151
R19493 vdd.n3177 vdd.n3176 10.6151
R19494 vdd.n3176 vdd.n3175 10.6151
R19495 vdd.n3175 vdd.n762 10.6151
R19496 vdd.n3170 vdd.n762 10.6151
R19497 vdd.n3170 vdd.n3169 10.6151
R19498 vdd.n3169 vdd.n3168 10.6151
R19499 vdd.n3168 vdd.n765 10.6151
R19500 vdd.n3163 vdd.n3162 10.6151
R19501 vdd.n3162 vdd.n3161 10.6151
R19502 vdd.n2924 vdd.n2923 10.6151
R19503 vdd.n2923 vdd.n2921 10.6151
R19504 vdd.n2921 vdd.n2920 10.6151
R19505 vdd.n2920 vdd.n2746 10.6151
R19506 vdd.n2820 vdd.n2746 10.6151
R19507 vdd.n2821 vdd.n2820 10.6151
R19508 vdd.n2823 vdd.n2821 10.6151
R19509 vdd.n2824 vdd.n2823 10.6151
R19510 vdd.n2904 vdd.n2824 10.6151
R19511 vdd.n2904 vdd.n2903 10.6151
R19512 vdd.n2903 vdd.n2902 10.6151
R19513 vdd.n2902 vdd.n2900 10.6151
R19514 vdd.n2900 vdd.n2899 10.6151
R19515 vdd.n2899 vdd.n2897 10.6151
R19516 vdd.n2897 vdd.n2896 10.6151
R19517 vdd.n2896 vdd.n2856 10.6151
R19518 vdd.n2856 vdd.n2855 10.6151
R19519 vdd.n2855 vdd.n2853 10.6151
R19520 vdd.n2853 vdd.n2852 10.6151
R19521 vdd.n2852 vdd.n2850 10.6151
R19522 vdd.n2850 vdd.n2849 10.6151
R19523 vdd.n2849 vdd.n2847 10.6151
R19524 vdd.n2847 vdd.n2846 10.6151
R19525 vdd.n2846 vdd.n2844 10.6151
R19526 vdd.n2844 vdd.n2843 10.6151
R19527 vdd.n2843 vdd.n2841 10.6151
R19528 vdd.n2841 vdd.n2840 10.6151
R19529 vdd.n2840 vdd.n2838 10.6151
R19530 vdd.n2838 vdd.n2837 10.6151
R19531 vdd.n2837 vdd.n2835 10.6151
R19532 vdd.n2835 vdd.n2834 10.6151
R19533 vdd.n2834 vdd.n2832 10.6151
R19534 vdd.n2832 vdd.n2831 10.6151
R19535 vdd.n2831 vdd.n2829 10.6151
R19536 vdd.n2829 vdd.n2828 10.6151
R19537 vdd.n2828 vdd.n2826 10.6151
R19538 vdd.n2826 vdd.n2825 10.6151
R19539 vdd.n2825 vdd.n771 10.6151
R19540 vdd.n2681 vdd.n913 10.6151
R19541 vdd.n2684 vdd.n2681 10.6151
R19542 vdd.n2685 vdd.n2684 10.6151
R19543 vdd.n2688 vdd.n2685 10.6151
R19544 vdd.n2689 vdd.n2688 10.6151
R19545 vdd.n2692 vdd.n2689 10.6151
R19546 vdd.n2693 vdd.n2692 10.6151
R19547 vdd.n2696 vdd.n2693 10.6151
R19548 vdd.n2697 vdd.n2696 10.6151
R19549 vdd.n2700 vdd.n2697 10.6151
R19550 vdd.n2701 vdd.n2700 10.6151
R19551 vdd.n2704 vdd.n2701 10.6151
R19552 vdd.n2705 vdd.n2704 10.6151
R19553 vdd.n2708 vdd.n2705 10.6151
R19554 vdd.n2709 vdd.n2708 10.6151
R19555 vdd.n2712 vdd.n2709 10.6151
R19556 vdd.n2713 vdd.n2712 10.6151
R19557 vdd.n2716 vdd.n2713 10.6151
R19558 vdd.n2717 vdd.n2716 10.6151
R19559 vdd.n2720 vdd.n2717 10.6151
R19560 vdd.n2721 vdd.n2720 10.6151
R19561 vdd.n2724 vdd.n2721 10.6151
R19562 vdd.n2725 vdd.n2724 10.6151
R19563 vdd.n2728 vdd.n2725 10.6151
R19564 vdd.n2729 vdd.n2728 10.6151
R19565 vdd.n2732 vdd.n2729 10.6151
R19566 vdd.n2733 vdd.n2732 10.6151
R19567 vdd.n2736 vdd.n2733 10.6151
R19568 vdd.n2737 vdd.n2736 10.6151
R19569 vdd.n2740 vdd.n2737 10.6151
R19570 vdd.n2741 vdd.n2740 10.6151
R19571 vdd.n2745 vdd.n2744 10.6151
R19572 vdd.n2925 vdd.n2745 10.6151
R19573 vdd.n2937 vdd.n2936 10.6151
R19574 vdd.n2938 vdd.n2937 10.6151
R19575 vdd.n2938 vdd.n903 10.6151
R19576 vdd.n2948 vdd.n903 10.6151
R19577 vdd.n2949 vdd.n2948 10.6151
R19578 vdd.n2950 vdd.n2949 10.6151
R19579 vdd.n2950 vdd.n891 10.6151
R19580 vdd.n2960 vdd.n891 10.6151
R19581 vdd.n2961 vdd.n2960 10.6151
R19582 vdd.n2962 vdd.n2961 10.6151
R19583 vdd.n2962 vdd.n880 10.6151
R19584 vdd.n2972 vdd.n880 10.6151
R19585 vdd.n2973 vdd.n2972 10.6151
R19586 vdd.n2974 vdd.n2973 10.6151
R19587 vdd.n2974 vdd.n868 10.6151
R19588 vdd.n2984 vdd.n868 10.6151
R19589 vdd.n2985 vdd.n2984 10.6151
R19590 vdd.n2986 vdd.n2985 10.6151
R19591 vdd.n2986 vdd.n857 10.6151
R19592 vdd.n2996 vdd.n857 10.6151
R19593 vdd.n2999 vdd.n2998 10.6151
R19594 vdd.n2999 vdd.n843 10.6151
R19595 vdd.n3009 vdd.n843 10.6151
R19596 vdd.n3010 vdd.n3009 10.6151
R19597 vdd.n3011 vdd.n3010 10.6151
R19598 vdd.n3011 vdd.n831 10.6151
R19599 vdd.n3021 vdd.n831 10.6151
R19600 vdd.n3022 vdd.n3021 10.6151
R19601 vdd.n3023 vdd.n3022 10.6151
R19602 vdd.n3023 vdd.n820 10.6151
R19603 vdd.n3033 vdd.n820 10.6151
R19604 vdd.n3034 vdd.n3033 10.6151
R19605 vdd.n3080 vdd.n3034 10.6151
R19606 vdd.n3080 vdd.n3079 10.6151
R19607 vdd.n3079 vdd.n3078 10.6151
R19608 vdd.n3078 vdd.n3077 10.6151
R19609 vdd.n3077 vdd.n3075 10.6151
R19610 vdd.n2387 vdd.n2386 10.6151
R19611 vdd.n2388 vdd.n2387 10.6151
R19612 vdd.n2388 vdd.n1067 10.6151
R19613 vdd.n2398 vdd.n1067 10.6151
R19614 vdd.n2399 vdd.n2398 10.6151
R19615 vdd.n2400 vdd.n2399 10.6151
R19616 vdd.n2400 vdd.n1055 10.6151
R19617 vdd.n2410 vdd.n1055 10.6151
R19618 vdd.n2411 vdd.n2410 10.6151
R19619 vdd.n2412 vdd.n2411 10.6151
R19620 vdd.n2412 vdd.n1043 10.6151
R19621 vdd.n2422 vdd.n1043 10.6151
R19622 vdd.n2423 vdd.n2422 10.6151
R19623 vdd.n2424 vdd.n2423 10.6151
R19624 vdd.n2424 vdd.n1030 10.6151
R19625 vdd.n2434 vdd.n1030 10.6151
R19626 vdd.n2435 vdd.n2434 10.6151
R19627 vdd.n2437 vdd.n1018 10.6151
R19628 vdd.n2447 vdd.n1018 10.6151
R19629 vdd.n2448 vdd.n2447 10.6151
R19630 vdd.n2449 vdd.n2448 10.6151
R19631 vdd.n2449 vdd.n1006 10.6151
R19632 vdd.n2459 vdd.n1006 10.6151
R19633 vdd.n2460 vdd.n2459 10.6151
R19634 vdd.n2461 vdd.n2460 10.6151
R19635 vdd.n2461 vdd.n995 10.6151
R19636 vdd.n2471 vdd.n995 10.6151
R19637 vdd.n2472 vdd.n2471 10.6151
R19638 vdd.n2473 vdd.n2472 10.6151
R19639 vdd.n2473 vdd.n984 10.6151
R19640 vdd.n2483 vdd.n984 10.6151
R19641 vdd.n2484 vdd.n2483 10.6151
R19642 vdd.n2487 vdd.n2484 10.6151
R19643 vdd.n2487 vdd.n2486 10.6151
R19644 vdd.n2486 vdd.n2485 10.6151
R19645 vdd.n2485 vdd.n967 10.6151
R19646 vdd.n2569 vdd.n967 10.6151
R19647 vdd.n2568 vdd.n2567 10.6151
R19648 vdd.n2567 vdd.n2564 10.6151
R19649 vdd.n2564 vdd.n2563 10.6151
R19650 vdd.n2563 vdd.n2560 10.6151
R19651 vdd.n2560 vdd.n2559 10.6151
R19652 vdd.n2559 vdd.n2556 10.6151
R19653 vdd.n2556 vdd.n2555 10.6151
R19654 vdd.n2555 vdd.n2552 10.6151
R19655 vdd.n2552 vdd.n2551 10.6151
R19656 vdd.n2551 vdd.n2548 10.6151
R19657 vdd.n2548 vdd.n2547 10.6151
R19658 vdd.n2547 vdd.n2544 10.6151
R19659 vdd.n2544 vdd.n2543 10.6151
R19660 vdd.n2543 vdd.n2540 10.6151
R19661 vdd.n2540 vdd.n2539 10.6151
R19662 vdd.n2539 vdd.n2536 10.6151
R19663 vdd.n2536 vdd.n2535 10.6151
R19664 vdd.n2535 vdd.n2532 10.6151
R19665 vdd.n2532 vdd.n2531 10.6151
R19666 vdd.n2531 vdd.n2528 10.6151
R19667 vdd.n2528 vdd.n2527 10.6151
R19668 vdd.n2527 vdd.n2524 10.6151
R19669 vdd.n2524 vdd.n2523 10.6151
R19670 vdd.n2523 vdd.n2520 10.6151
R19671 vdd.n2520 vdd.n2519 10.6151
R19672 vdd.n2519 vdd.n2516 10.6151
R19673 vdd.n2516 vdd.n2515 10.6151
R19674 vdd.n2515 vdd.n2512 10.6151
R19675 vdd.n2512 vdd.n2511 10.6151
R19676 vdd.n2511 vdd.n2508 10.6151
R19677 vdd.n2508 vdd.n2507 10.6151
R19678 vdd.n2504 vdd.n2503 10.6151
R19679 vdd.n2503 vdd.n2501 10.6151
R19680 vdd.n2203 vdd.n2201 10.6151
R19681 vdd.n2204 vdd.n2203 10.6151
R19682 vdd.n2206 vdd.n2204 10.6151
R19683 vdd.n2207 vdd.n2206 10.6151
R19684 vdd.n2209 vdd.n2207 10.6151
R19685 vdd.n2210 vdd.n2209 10.6151
R19686 vdd.n2212 vdd.n2210 10.6151
R19687 vdd.n2213 vdd.n2212 10.6151
R19688 vdd.n2215 vdd.n2213 10.6151
R19689 vdd.n2216 vdd.n2215 10.6151
R19690 vdd.n2218 vdd.n2216 10.6151
R19691 vdd.n2219 vdd.n2218 10.6151
R19692 vdd.n2221 vdd.n2219 10.6151
R19693 vdd.n2222 vdd.n2221 10.6151
R19694 vdd.n2224 vdd.n2222 10.6151
R19695 vdd.n2225 vdd.n2224 10.6151
R19696 vdd.n2227 vdd.n2225 10.6151
R19697 vdd.n2228 vdd.n2227 10.6151
R19698 vdd.n2230 vdd.n2228 10.6151
R19699 vdd.n2231 vdd.n2230 10.6151
R19700 vdd.n2233 vdd.n2231 10.6151
R19701 vdd.n2234 vdd.n2233 10.6151
R19702 vdd.n2273 vdd.n2234 10.6151
R19703 vdd.n2273 vdd.n2272 10.6151
R19704 vdd.n2272 vdd.n2271 10.6151
R19705 vdd.n2271 vdd.n2269 10.6151
R19706 vdd.n2269 vdd.n2268 10.6151
R19707 vdd.n2268 vdd.n2266 10.6151
R19708 vdd.n2266 vdd.n2265 10.6151
R19709 vdd.n2265 vdd.n2242 10.6151
R19710 vdd.n2242 vdd.n2241 10.6151
R19711 vdd.n2241 vdd.n2239 10.6151
R19712 vdd.n2239 vdd.n2238 10.6151
R19713 vdd.n2238 vdd.n2236 10.6151
R19714 vdd.n2236 vdd.n2235 10.6151
R19715 vdd.n2235 vdd.n971 10.6151
R19716 vdd.n2499 vdd.n971 10.6151
R19717 vdd.n2500 vdd.n2499 10.6151
R19718 vdd.n2131 vdd.n1079 10.6151
R19719 vdd.n2136 vdd.n2131 10.6151
R19720 vdd.n2137 vdd.n2136 10.6151
R19721 vdd.n2138 vdd.n2137 10.6151
R19722 vdd.n2138 vdd.n2129 10.6151
R19723 vdd.n2144 vdd.n2129 10.6151
R19724 vdd.n2145 vdd.n2144 10.6151
R19725 vdd.n2146 vdd.n2145 10.6151
R19726 vdd.n2146 vdd.n2127 10.6151
R19727 vdd.n2152 vdd.n2127 10.6151
R19728 vdd.n2153 vdd.n2152 10.6151
R19729 vdd.n2154 vdd.n2153 10.6151
R19730 vdd.n2154 vdd.n2125 10.6151
R19731 vdd.n2160 vdd.n2125 10.6151
R19732 vdd.n2161 vdd.n2160 10.6151
R19733 vdd.n2162 vdd.n2161 10.6151
R19734 vdd.n2162 vdd.n2123 10.6151
R19735 vdd.n2168 vdd.n2123 10.6151
R19736 vdd.n2169 vdd.n2168 10.6151
R19737 vdd.n2170 vdd.n2169 10.6151
R19738 vdd.n2170 vdd.n1113 10.6151
R19739 vdd.n2176 vdd.n1113 10.6151
R19740 vdd.n2177 vdd.n2176 10.6151
R19741 vdd.n2178 vdd.n2177 10.6151
R19742 vdd.n2178 vdd.n1111 10.6151
R19743 vdd.n2184 vdd.n1111 10.6151
R19744 vdd.n2185 vdd.n2184 10.6151
R19745 vdd.n2186 vdd.n2185 10.6151
R19746 vdd.n2186 vdd.n1109 10.6151
R19747 vdd.n2192 vdd.n1109 10.6151
R19748 vdd.n2193 vdd.n2192 10.6151
R19749 vdd.n2195 vdd.n1105 10.6151
R19750 vdd.n2200 vdd.n1105 10.6151
R19751 vdd.t36 vdd.n1856 10.5435
R19752 vdd.n636 vdd.t33 10.5435
R19753 vdd.n304 vdd.n286 10.4732
R19754 vdd.n249 vdd.n231 10.4732
R19755 vdd.n206 vdd.n188 10.4732
R19756 vdd.n151 vdd.n133 10.4732
R19757 vdd.n109 vdd.n91 10.4732
R19758 vdd.n54 vdd.n36 10.4732
R19759 vdd.n1753 vdd.n1735 10.4732
R19760 vdd.n1808 vdd.n1790 10.4732
R19761 vdd.n1655 vdd.n1637 10.4732
R19762 vdd.n1710 vdd.n1692 10.4732
R19763 vdd.n1558 vdd.n1540 10.4732
R19764 vdd.n1613 vdd.n1595 10.4732
R19765 vdd.n1840 vdd.t93 10.3167
R19766 vdd.n3387 vdd.t31 10.3167
R19767 vdd.n2571 vdd.t242 10.2034
R19768 vdd.n2934 vdd.t230 10.2034
R19769 vdd.t48 vdd.n1184 10.09
R19770 vdd.n1892 vdd.t171 10.09
R19771 vdd.n3335 vdd.t145 10.09
R19772 vdd.n3468 vdd.t27 10.09
R19773 vdd.n2099 vdd.n1093 9.88581
R19774 vdd.n3125 vdd.n3124 9.88581
R19775 vdd.n3192 vdd.n3191 9.88581
R19776 vdd.n2123 vdd.n2122 9.88581
R19777 vdd.n1504 vdd.t69 9.86327
R19778 vdd.n3459 vdd.t17 9.86327
R19779 vdd.n303 vdd.n288 9.69747
R19780 vdd.n248 vdd.n233 9.69747
R19781 vdd.n205 vdd.n190 9.69747
R19782 vdd.n150 vdd.n135 9.69747
R19783 vdd.n108 vdd.n93 9.69747
R19784 vdd.n53 vdd.n38 9.69747
R19785 vdd.n1752 vdd.n1737 9.69747
R19786 vdd.n1807 vdd.n1792 9.69747
R19787 vdd.n1654 vdd.n1639 9.69747
R19788 vdd.n1709 vdd.n1694 9.69747
R19789 vdd.n1557 vdd.n1542 9.69747
R19790 vdd.n1612 vdd.n1597 9.69747
R19791 vdd.t13 vdd.n1478 9.63654
R19792 vdd.n3418 vdd.t29 9.63654
R19793 vdd.n319 vdd.n318 9.45567
R19794 vdd.n264 vdd.n263 9.45567
R19795 vdd.n221 vdd.n220 9.45567
R19796 vdd.n166 vdd.n165 9.45567
R19797 vdd.n124 vdd.n123 9.45567
R19798 vdd.n69 vdd.n68 9.45567
R19799 vdd.n1768 vdd.n1767 9.45567
R19800 vdd.n1823 vdd.n1822 9.45567
R19801 vdd.n1670 vdd.n1669 9.45567
R19802 vdd.n1725 vdd.n1724 9.45567
R19803 vdd.n1573 vdd.n1572 9.45567
R19804 vdd.n1628 vdd.n1627 9.45567
R19805 vdd.n2072 vdd.n1926 9.3005
R19806 vdd.n2071 vdd.n2070 9.3005
R19807 vdd.n1932 vdd.n1931 9.3005
R19808 vdd.n2065 vdd.n1936 9.3005
R19809 vdd.n2064 vdd.n1937 9.3005
R19810 vdd.n2063 vdd.n1938 9.3005
R19811 vdd.n1942 vdd.n1939 9.3005
R19812 vdd.n2058 vdd.n1943 9.3005
R19813 vdd.n2057 vdd.n1944 9.3005
R19814 vdd.n2056 vdd.n1945 9.3005
R19815 vdd.n1949 vdd.n1946 9.3005
R19816 vdd.n2051 vdd.n1950 9.3005
R19817 vdd.n2050 vdd.n1951 9.3005
R19818 vdd.n2049 vdd.n1952 9.3005
R19819 vdd.n1956 vdd.n1953 9.3005
R19820 vdd.n2044 vdd.n1957 9.3005
R19821 vdd.n2043 vdd.n1958 9.3005
R19822 vdd.n2042 vdd.n1959 9.3005
R19823 vdd.n1963 vdd.n1960 9.3005
R19824 vdd.n2037 vdd.n1964 9.3005
R19825 vdd.n2036 vdd.n1965 9.3005
R19826 vdd.n2035 vdd.n2034 9.3005
R19827 vdd.n2033 vdd.n1966 9.3005
R19828 vdd.n2032 vdd.n2031 9.3005
R19829 vdd.n1972 vdd.n1971 9.3005
R19830 vdd.n2026 vdd.n1976 9.3005
R19831 vdd.n2025 vdd.n1977 9.3005
R19832 vdd.n2024 vdd.n1978 9.3005
R19833 vdd.n1982 vdd.n1979 9.3005
R19834 vdd.n2019 vdd.n1983 9.3005
R19835 vdd.n2018 vdd.n1984 9.3005
R19836 vdd.n2017 vdd.n1985 9.3005
R19837 vdd.n1989 vdd.n1986 9.3005
R19838 vdd.n2012 vdd.n1990 9.3005
R19839 vdd.n2011 vdd.n1991 9.3005
R19840 vdd.n2010 vdd.n1992 9.3005
R19841 vdd.n1994 vdd.n1993 9.3005
R19842 vdd.n2005 vdd.n1115 9.3005
R19843 vdd.n2074 vdd.n2073 9.3005
R19844 vdd.n2098 vdd.n2097 9.3005
R19845 vdd.n1904 vdd.n1903 9.3005
R19846 vdd.n1909 vdd.n1907 9.3005
R19847 vdd.n2090 vdd.n1910 9.3005
R19848 vdd.n2089 vdd.n1911 9.3005
R19849 vdd.n2088 vdd.n1912 9.3005
R19850 vdd.n1916 vdd.n1913 9.3005
R19851 vdd.n2083 vdd.n1917 9.3005
R19852 vdd.n2082 vdd.n1918 9.3005
R19853 vdd.n2081 vdd.n1919 9.3005
R19854 vdd.n1923 vdd.n1920 9.3005
R19855 vdd.n2076 vdd.n1924 9.3005
R19856 vdd.n2075 vdd.n1925 9.3005
R19857 vdd.n2107 vdd.n1897 9.3005
R19858 vdd.n2109 vdd.n2108 9.3005
R19859 vdd.n1828 vdd.n1174 9.3005
R19860 vdd.n1830 vdd.n1829 9.3005
R19861 vdd.n1165 vdd.n1164 9.3005
R19862 vdd.n1843 vdd.n1842 9.3005
R19863 vdd.n1844 vdd.n1163 9.3005
R19864 vdd.n1846 vdd.n1845 9.3005
R19865 vdd.n1153 vdd.n1152 9.3005
R19866 vdd.n1860 vdd.n1859 9.3005
R19867 vdd.n1861 vdd.n1151 9.3005
R19868 vdd.n1863 vdd.n1862 9.3005
R19869 vdd.n1142 vdd.n1141 9.3005
R19870 vdd.n1877 vdd.n1876 9.3005
R19871 vdd.n1878 vdd.n1140 9.3005
R19872 vdd.n1880 vdd.n1879 9.3005
R19873 vdd.n1130 vdd.n1129 9.3005
R19874 vdd.n1895 vdd.n1894 9.3005
R19875 vdd.n1896 vdd.n1128 9.3005
R19876 vdd.n2111 vdd.n2110 9.3005
R19877 vdd.n295 vdd.n294 9.3005
R19878 vdd.n290 vdd.n289 9.3005
R19879 vdd.n301 vdd.n300 9.3005
R19880 vdd.n303 vdd.n302 9.3005
R19881 vdd.n286 vdd.n285 9.3005
R19882 vdd.n309 vdd.n308 9.3005
R19883 vdd.n311 vdd.n310 9.3005
R19884 vdd.n283 vdd.n280 9.3005
R19885 vdd.n318 vdd.n317 9.3005
R19886 vdd.n240 vdd.n239 9.3005
R19887 vdd.n235 vdd.n234 9.3005
R19888 vdd.n246 vdd.n245 9.3005
R19889 vdd.n248 vdd.n247 9.3005
R19890 vdd.n231 vdd.n230 9.3005
R19891 vdd.n254 vdd.n253 9.3005
R19892 vdd.n256 vdd.n255 9.3005
R19893 vdd.n228 vdd.n225 9.3005
R19894 vdd.n263 vdd.n262 9.3005
R19895 vdd.n197 vdd.n196 9.3005
R19896 vdd.n192 vdd.n191 9.3005
R19897 vdd.n203 vdd.n202 9.3005
R19898 vdd.n205 vdd.n204 9.3005
R19899 vdd.n188 vdd.n187 9.3005
R19900 vdd.n211 vdd.n210 9.3005
R19901 vdd.n213 vdd.n212 9.3005
R19902 vdd.n185 vdd.n182 9.3005
R19903 vdd.n220 vdd.n219 9.3005
R19904 vdd.n142 vdd.n141 9.3005
R19905 vdd.n137 vdd.n136 9.3005
R19906 vdd.n148 vdd.n147 9.3005
R19907 vdd.n150 vdd.n149 9.3005
R19908 vdd.n133 vdd.n132 9.3005
R19909 vdd.n156 vdd.n155 9.3005
R19910 vdd.n158 vdd.n157 9.3005
R19911 vdd.n130 vdd.n127 9.3005
R19912 vdd.n165 vdd.n164 9.3005
R19913 vdd.n100 vdd.n99 9.3005
R19914 vdd.n95 vdd.n94 9.3005
R19915 vdd.n106 vdd.n105 9.3005
R19916 vdd.n108 vdd.n107 9.3005
R19917 vdd.n91 vdd.n90 9.3005
R19918 vdd.n114 vdd.n113 9.3005
R19919 vdd.n116 vdd.n115 9.3005
R19920 vdd.n88 vdd.n85 9.3005
R19921 vdd.n123 vdd.n122 9.3005
R19922 vdd.n45 vdd.n44 9.3005
R19923 vdd.n40 vdd.n39 9.3005
R19924 vdd.n51 vdd.n50 9.3005
R19925 vdd.n53 vdd.n52 9.3005
R19926 vdd.n36 vdd.n35 9.3005
R19927 vdd.n59 vdd.n58 9.3005
R19928 vdd.n61 vdd.n60 9.3005
R19929 vdd.n33 vdd.n30 9.3005
R19930 vdd.n68 vdd.n67 9.3005
R19931 vdd.n3241 vdd.n3240 9.3005
R19932 vdd.n3242 vdd.n721 9.3005
R19933 vdd.n720 vdd.n718 9.3005
R19934 vdd.n3248 vdd.n717 9.3005
R19935 vdd.n3249 vdd.n716 9.3005
R19936 vdd.n3250 vdd.n715 9.3005
R19937 vdd.n714 vdd.n712 9.3005
R19938 vdd.n3256 vdd.n711 9.3005
R19939 vdd.n3257 vdd.n710 9.3005
R19940 vdd.n3258 vdd.n709 9.3005
R19941 vdd.n708 vdd.n706 9.3005
R19942 vdd.n3264 vdd.n705 9.3005
R19943 vdd.n3265 vdd.n704 9.3005
R19944 vdd.n3266 vdd.n703 9.3005
R19945 vdd.n702 vdd.n700 9.3005
R19946 vdd.n3272 vdd.n699 9.3005
R19947 vdd.n3273 vdd.n698 9.3005
R19948 vdd.n3274 vdd.n697 9.3005
R19949 vdd.n696 vdd.n694 9.3005
R19950 vdd.n3280 vdd.n693 9.3005
R19951 vdd.n3281 vdd.n692 9.3005
R19952 vdd.n3282 vdd.n691 9.3005
R19953 vdd.n690 vdd.n688 9.3005
R19954 vdd.n3288 vdd.n685 9.3005
R19955 vdd.n3289 vdd.n684 9.3005
R19956 vdd.n3290 vdd.n683 9.3005
R19957 vdd.n682 vdd.n680 9.3005
R19958 vdd.n3296 vdd.n679 9.3005
R19959 vdd.n3297 vdd.n678 9.3005
R19960 vdd.n3298 vdd.n677 9.3005
R19961 vdd.n676 vdd.n674 9.3005
R19962 vdd.n3304 vdd.n673 9.3005
R19963 vdd.n3305 vdd.n672 9.3005
R19964 vdd.n3306 vdd.n671 9.3005
R19965 vdd.n670 vdd.n668 9.3005
R19966 vdd.n3311 vdd.n667 9.3005
R19967 vdd.n3321 vdd.n661 9.3005
R19968 vdd.n3323 vdd.n3322 9.3005
R19969 vdd.n652 vdd.n651 9.3005
R19970 vdd.n3338 vdd.n3337 9.3005
R19971 vdd.n3339 vdd.n650 9.3005
R19972 vdd.n3341 vdd.n3340 9.3005
R19973 vdd.n640 vdd.n639 9.3005
R19974 vdd.n3354 vdd.n3353 9.3005
R19975 vdd.n3355 vdd.n638 9.3005
R19976 vdd.n3357 vdd.n3356 9.3005
R19977 vdd.n628 vdd.n627 9.3005
R19978 vdd.n3371 vdd.n3370 9.3005
R19979 vdd.n3372 vdd.n626 9.3005
R19980 vdd.n3374 vdd.n3373 9.3005
R19981 vdd.n617 vdd.n616 9.3005
R19982 vdd.n3390 vdd.n3389 9.3005
R19983 vdd.n3391 vdd.n615 9.3005
R19984 vdd.n3393 vdd.n3392 9.3005
R19985 vdd.n324 vdd.n322 9.3005
R19986 vdd.n3325 vdd.n3324 9.3005
R19987 vdd.n3472 vdd.n3471 9.3005
R19988 vdd.n325 vdd.n323 9.3005
R19989 vdd.n3465 vdd.n334 9.3005
R19990 vdd.n3464 vdd.n335 9.3005
R19991 vdd.n3463 vdd.n336 9.3005
R19992 vdd.n343 vdd.n337 9.3005
R19993 vdd.n3457 vdd.n344 9.3005
R19994 vdd.n3456 vdd.n345 9.3005
R19995 vdd.n3455 vdd.n346 9.3005
R19996 vdd.n354 vdd.n347 9.3005
R19997 vdd.n3449 vdd.n355 9.3005
R19998 vdd.n3448 vdd.n356 9.3005
R19999 vdd.n3447 vdd.n357 9.3005
R20000 vdd.n365 vdd.n358 9.3005
R20001 vdd.n3441 vdd.n366 9.3005
R20002 vdd.n3440 vdd.n367 9.3005
R20003 vdd.n3439 vdd.n368 9.3005
R20004 vdd.n443 vdd.n369 9.3005
R20005 vdd.n447 vdd.n442 9.3005
R20006 vdd.n451 vdd.n450 9.3005
R20007 vdd.n452 vdd.n441 9.3005
R20008 vdd.n456 vdd.n453 9.3005
R20009 vdd.n457 vdd.n440 9.3005
R20010 vdd.n461 vdd.n460 9.3005
R20011 vdd.n462 vdd.n439 9.3005
R20012 vdd.n466 vdd.n463 9.3005
R20013 vdd.n467 vdd.n438 9.3005
R20014 vdd.n471 vdd.n470 9.3005
R20015 vdd.n472 vdd.n437 9.3005
R20016 vdd.n476 vdd.n473 9.3005
R20017 vdd.n477 vdd.n436 9.3005
R20018 vdd.n481 vdd.n480 9.3005
R20019 vdd.n482 vdd.n435 9.3005
R20020 vdd.n486 vdd.n483 9.3005
R20021 vdd.n487 vdd.n434 9.3005
R20022 vdd.n491 vdd.n490 9.3005
R20023 vdd.n492 vdd.n433 9.3005
R20024 vdd.n496 vdd.n493 9.3005
R20025 vdd.n497 vdd.n430 9.3005
R20026 vdd.n501 vdd.n500 9.3005
R20027 vdd.n502 vdd.n429 9.3005
R20028 vdd.n506 vdd.n503 9.3005
R20029 vdd.n507 vdd.n428 9.3005
R20030 vdd.n511 vdd.n510 9.3005
R20031 vdd.n512 vdd.n427 9.3005
R20032 vdd.n516 vdd.n513 9.3005
R20033 vdd.n517 vdd.n426 9.3005
R20034 vdd.n521 vdd.n520 9.3005
R20035 vdd.n522 vdd.n425 9.3005
R20036 vdd.n526 vdd.n523 9.3005
R20037 vdd.n527 vdd.n424 9.3005
R20038 vdd.n531 vdd.n530 9.3005
R20039 vdd.n532 vdd.n423 9.3005
R20040 vdd.n536 vdd.n533 9.3005
R20041 vdd.n537 vdd.n422 9.3005
R20042 vdd.n541 vdd.n540 9.3005
R20043 vdd.n542 vdd.n421 9.3005
R20044 vdd.n546 vdd.n543 9.3005
R20045 vdd.n547 vdd.n418 9.3005
R20046 vdd.n551 vdd.n550 9.3005
R20047 vdd.n552 vdd.n417 9.3005
R20048 vdd.n556 vdd.n553 9.3005
R20049 vdd.n557 vdd.n416 9.3005
R20050 vdd.n561 vdd.n560 9.3005
R20051 vdd.n562 vdd.n415 9.3005
R20052 vdd.n566 vdd.n563 9.3005
R20053 vdd.n567 vdd.n414 9.3005
R20054 vdd.n571 vdd.n570 9.3005
R20055 vdd.n572 vdd.n413 9.3005
R20056 vdd.n576 vdd.n573 9.3005
R20057 vdd.n577 vdd.n412 9.3005
R20058 vdd.n581 vdd.n580 9.3005
R20059 vdd.n582 vdd.n411 9.3005
R20060 vdd.n586 vdd.n583 9.3005
R20061 vdd.n587 vdd.n410 9.3005
R20062 vdd.n591 vdd.n590 9.3005
R20063 vdd.n592 vdd.n409 9.3005
R20064 vdd.n596 vdd.n593 9.3005
R20065 vdd.n598 vdd.n408 9.3005
R20066 vdd.n600 vdd.n599 9.3005
R20067 vdd.n3432 vdd.n3431 9.3005
R20068 vdd.n446 vdd.n444 9.3005
R20069 vdd.n3331 vdd.n655 9.3005
R20070 vdd.n3333 vdd.n3332 9.3005
R20071 vdd.n646 vdd.n645 9.3005
R20072 vdd.n3346 vdd.n3345 9.3005
R20073 vdd.n3347 vdd.n644 9.3005
R20074 vdd.n3349 vdd.n3348 9.3005
R20075 vdd.n633 vdd.n632 9.3005
R20076 vdd.n3362 vdd.n3361 9.3005
R20077 vdd.n3363 vdd.n631 9.3005
R20078 vdd.n3365 vdd.n3364 9.3005
R20079 vdd.n622 vdd.n621 9.3005
R20080 vdd.n3379 vdd.n3378 9.3005
R20081 vdd.n3380 vdd.n620 9.3005
R20082 vdd.n3385 vdd.n3381 9.3005
R20083 vdd.n3384 vdd.n3383 9.3005
R20084 vdd.n3382 vdd.n610 9.3005
R20085 vdd.n3398 vdd.n611 9.3005
R20086 vdd.n3399 vdd.n609 9.3005
R20087 vdd.n3401 vdd.n3400 9.3005
R20088 vdd.n3402 vdd.n608 9.3005
R20089 vdd.n3405 vdd.n3403 9.3005
R20090 vdd.n3406 vdd.n607 9.3005
R20091 vdd.n3408 vdd.n3407 9.3005
R20092 vdd.n3409 vdd.n606 9.3005
R20093 vdd.n3412 vdd.n3410 9.3005
R20094 vdd.n3413 vdd.n605 9.3005
R20095 vdd.n3415 vdd.n3414 9.3005
R20096 vdd.n3416 vdd.n604 9.3005
R20097 vdd.n3420 vdd.n3417 9.3005
R20098 vdd.n3421 vdd.n603 9.3005
R20099 vdd.n3423 vdd.n3422 9.3005
R20100 vdd.n3424 vdd.n602 9.3005
R20101 vdd.n3427 vdd.n3425 9.3005
R20102 vdd.n3428 vdd.n601 9.3005
R20103 vdd.n3430 vdd.n3429 9.3005
R20104 vdd.n3330 vdd.n3329 9.3005
R20105 vdd.n3194 vdd.n656 9.3005
R20106 vdd.n3199 vdd.n3193 9.3005
R20107 vdd.n3209 vdd.n748 9.3005
R20108 vdd.n3210 vdd.n747 9.3005
R20109 vdd.n746 vdd.n744 9.3005
R20110 vdd.n3216 vdd.n743 9.3005
R20111 vdd.n3217 vdd.n742 9.3005
R20112 vdd.n3218 vdd.n741 9.3005
R20113 vdd.n740 vdd.n738 9.3005
R20114 vdd.n3224 vdd.n737 9.3005
R20115 vdd.n3225 vdd.n736 9.3005
R20116 vdd.n3226 vdd.n735 9.3005
R20117 vdd.n734 vdd.n732 9.3005
R20118 vdd.n3231 vdd.n731 9.3005
R20119 vdd.n3232 vdd.n730 9.3005
R20120 vdd.n726 vdd.n725 9.3005
R20121 vdd.n3238 vdd.n3237 9.3005
R20122 vdd.n3239 vdd.n722 9.3005
R20123 vdd.n2121 vdd.n2120 9.3005
R20124 vdd.n2116 vdd.n1118 9.3005
R20125 vdd.n1460 vdd.n1459 9.3005
R20126 vdd.n1216 vdd.n1215 9.3005
R20127 vdd.n1473 vdd.n1472 9.3005
R20128 vdd.n1474 vdd.n1214 9.3005
R20129 vdd.n1476 vdd.n1475 9.3005
R20130 vdd.n1204 vdd.n1203 9.3005
R20131 vdd.n1490 vdd.n1489 9.3005
R20132 vdd.n1491 vdd.n1202 9.3005
R20133 vdd.n1493 vdd.n1492 9.3005
R20134 vdd.n1194 vdd.n1193 9.3005
R20135 vdd.n1507 vdd.n1506 9.3005
R20136 vdd.n1508 vdd.n1192 9.3005
R20137 vdd.n1510 vdd.n1509 9.3005
R20138 vdd.n1181 vdd.n1180 9.3005
R20139 vdd.n1523 vdd.n1522 9.3005
R20140 vdd.n1524 vdd.n1179 9.3005
R20141 vdd.n1526 vdd.n1525 9.3005
R20142 vdd.n1170 vdd.n1169 9.3005
R20143 vdd.n1835 vdd.n1834 9.3005
R20144 vdd.n1836 vdd.n1168 9.3005
R20145 vdd.n1838 vdd.n1837 9.3005
R20146 vdd.n1159 vdd.n1158 9.3005
R20147 vdd.n1851 vdd.n1850 9.3005
R20148 vdd.n1852 vdd.n1157 9.3005
R20149 vdd.n1854 vdd.n1853 9.3005
R20150 vdd.n1147 vdd.n1146 9.3005
R20151 vdd.n1868 vdd.n1867 9.3005
R20152 vdd.n1869 vdd.n1145 9.3005
R20153 vdd.n1871 vdd.n1870 9.3005
R20154 vdd.n1137 vdd.n1136 9.3005
R20155 vdd.n1885 vdd.n1884 9.3005
R20156 vdd.n1886 vdd.n1134 9.3005
R20157 vdd.n1890 vdd.n1889 9.3005
R20158 vdd.n1888 vdd.n1135 9.3005
R20159 vdd.n1887 vdd.n1123 9.3005
R20160 vdd.n1458 vdd.n1226 9.3005
R20161 vdd.n1351 vdd.n1227 9.3005
R20162 vdd.n1353 vdd.n1352 9.3005
R20163 vdd.n1354 vdd.n1346 9.3005
R20164 vdd.n1356 vdd.n1355 9.3005
R20165 vdd.n1357 vdd.n1345 9.3005
R20166 vdd.n1359 vdd.n1358 9.3005
R20167 vdd.n1360 vdd.n1340 9.3005
R20168 vdd.n1362 vdd.n1361 9.3005
R20169 vdd.n1363 vdd.n1339 9.3005
R20170 vdd.n1365 vdd.n1364 9.3005
R20171 vdd.n1366 vdd.n1334 9.3005
R20172 vdd.n1368 vdd.n1367 9.3005
R20173 vdd.n1369 vdd.n1333 9.3005
R20174 vdd.n1371 vdd.n1370 9.3005
R20175 vdd.n1372 vdd.n1328 9.3005
R20176 vdd.n1374 vdd.n1373 9.3005
R20177 vdd.n1375 vdd.n1327 9.3005
R20178 vdd.n1377 vdd.n1376 9.3005
R20179 vdd.n1378 vdd.n1322 9.3005
R20180 vdd.n1380 vdd.n1379 9.3005
R20181 vdd.n1381 vdd.n1321 9.3005
R20182 vdd.n1386 vdd.n1382 9.3005
R20183 vdd.n1387 vdd.n1317 9.3005
R20184 vdd.n1389 vdd.n1388 9.3005
R20185 vdd.n1390 vdd.n1316 9.3005
R20186 vdd.n1392 vdd.n1391 9.3005
R20187 vdd.n1393 vdd.n1311 9.3005
R20188 vdd.n1395 vdd.n1394 9.3005
R20189 vdd.n1396 vdd.n1310 9.3005
R20190 vdd.n1398 vdd.n1397 9.3005
R20191 vdd.n1399 vdd.n1305 9.3005
R20192 vdd.n1401 vdd.n1400 9.3005
R20193 vdd.n1402 vdd.n1304 9.3005
R20194 vdd.n1404 vdd.n1403 9.3005
R20195 vdd.n1405 vdd.n1299 9.3005
R20196 vdd.n1407 vdd.n1406 9.3005
R20197 vdd.n1408 vdd.n1298 9.3005
R20198 vdd.n1410 vdd.n1409 9.3005
R20199 vdd.n1411 vdd.n1293 9.3005
R20200 vdd.n1413 vdd.n1412 9.3005
R20201 vdd.n1414 vdd.n1292 9.3005
R20202 vdd.n1416 vdd.n1415 9.3005
R20203 vdd.n1417 vdd.n1289 9.3005
R20204 vdd.n1423 vdd.n1422 9.3005
R20205 vdd.n1424 vdd.n1288 9.3005
R20206 vdd.n1426 vdd.n1425 9.3005
R20207 vdd.n1427 vdd.n1283 9.3005
R20208 vdd.n1429 vdd.n1428 9.3005
R20209 vdd.n1430 vdd.n1282 9.3005
R20210 vdd.n1432 vdd.n1431 9.3005
R20211 vdd.n1433 vdd.n1277 9.3005
R20212 vdd.n1435 vdd.n1434 9.3005
R20213 vdd.n1436 vdd.n1276 9.3005
R20214 vdd.n1438 vdd.n1437 9.3005
R20215 vdd.n1439 vdd.n1271 9.3005
R20216 vdd.n1441 vdd.n1440 9.3005
R20217 vdd.n1442 vdd.n1270 9.3005
R20218 vdd.n1444 vdd.n1443 9.3005
R20219 vdd.n1445 vdd.n1266 9.3005
R20220 vdd.n1447 vdd.n1446 9.3005
R20221 vdd.n1448 vdd.n1265 9.3005
R20222 vdd.n1450 vdd.n1449 9.3005
R20223 vdd.n1451 vdd.n1264 9.3005
R20224 vdd.n1457 vdd.n1456 9.3005
R20225 vdd.n1465 vdd.n1464 9.3005
R20226 vdd.n1466 vdd.n1220 9.3005
R20227 vdd.n1468 vdd.n1467 9.3005
R20228 vdd.n1210 vdd.n1209 9.3005
R20229 vdd.n1482 vdd.n1481 9.3005
R20230 vdd.n1483 vdd.n1208 9.3005
R20231 vdd.n1485 vdd.n1484 9.3005
R20232 vdd.n1199 vdd.n1198 9.3005
R20233 vdd.n1499 vdd.n1498 9.3005
R20234 vdd.n1500 vdd.n1197 9.3005
R20235 vdd.n1502 vdd.n1501 9.3005
R20236 vdd.n1188 vdd.n1187 9.3005
R20237 vdd.n1515 vdd.n1514 9.3005
R20238 vdd.n1516 vdd.n1186 9.3005
R20239 vdd.n1518 vdd.n1517 9.3005
R20240 vdd.n1176 vdd.n1175 9.3005
R20241 vdd.n1532 vdd.n1531 9.3005
R20242 vdd.n1222 vdd.n1221 9.3005
R20243 vdd.n1744 vdd.n1743 9.3005
R20244 vdd.n1739 vdd.n1738 9.3005
R20245 vdd.n1750 vdd.n1749 9.3005
R20246 vdd.n1752 vdd.n1751 9.3005
R20247 vdd.n1735 vdd.n1734 9.3005
R20248 vdd.n1758 vdd.n1757 9.3005
R20249 vdd.n1760 vdd.n1759 9.3005
R20250 vdd.n1732 vdd.n1729 9.3005
R20251 vdd.n1767 vdd.n1766 9.3005
R20252 vdd.n1799 vdd.n1798 9.3005
R20253 vdd.n1794 vdd.n1793 9.3005
R20254 vdd.n1805 vdd.n1804 9.3005
R20255 vdd.n1807 vdd.n1806 9.3005
R20256 vdd.n1790 vdd.n1789 9.3005
R20257 vdd.n1813 vdd.n1812 9.3005
R20258 vdd.n1815 vdd.n1814 9.3005
R20259 vdd.n1787 vdd.n1784 9.3005
R20260 vdd.n1822 vdd.n1821 9.3005
R20261 vdd.n1646 vdd.n1645 9.3005
R20262 vdd.n1641 vdd.n1640 9.3005
R20263 vdd.n1652 vdd.n1651 9.3005
R20264 vdd.n1654 vdd.n1653 9.3005
R20265 vdd.n1637 vdd.n1636 9.3005
R20266 vdd.n1660 vdd.n1659 9.3005
R20267 vdd.n1662 vdd.n1661 9.3005
R20268 vdd.n1634 vdd.n1631 9.3005
R20269 vdd.n1669 vdd.n1668 9.3005
R20270 vdd.n1701 vdd.n1700 9.3005
R20271 vdd.n1696 vdd.n1695 9.3005
R20272 vdd.n1707 vdd.n1706 9.3005
R20273 vdd.n1709 vdd.n1708 9.3005
R20274 vdd.n1692 vdd.n1691 9.3005
R20275 vdd.n1715 vdd.n1714 9.3005
R20276 vdd.n1717 vdd.n1716 9.3005
R20277 vdd.n1689 vdd.n1686 9.3005
R20278 vdd.n1724 vdd.n1723 9.3005
R20279 vdd.n1549 vdd.n1548 9.3005
R20280 vdd.n1544 vdd.n1543 9.3005
R20281 vdd.n1555 vdd.n1554 9.3005
R20282 vdd.n1557 vdd.n1556 9.3005
R20283 vdd.n1540 vdd.n1539 9.3005
R20284 vdd.n1563 vdd.n1562 9.3005
R20285 vdd.n1565 vdd.n1564 9.3005
R20286 vdd.n1537 vdd.n1534 9.3005
R20287 vdd.n1572 vdd.n1571 9.3005
R20288 vdd.n1604 vdd.n1603 9.3005
R20289 vdd.n1599 vdd.n1598 9.3005
R20290 vdd.n1610 vdd.n1609 9.3005
R20291 vdd.n1612 vdd.n1611 9.3005
R20292 vdd.n1595 vdd.n1594 9.3005
R20293 vdd.n1618 vdd.n1617 9.3005
R20294 vdd.n1620 vdd.n1619 9.3005
R20295 vdd.n1592 vdd.n1589 9.3005
R20296 vdd.n1627 vdd.n1626 9.3005
R20297 vdd.n1478 vdd.t11 9.18308
R20298 vdd.n3418 vdd.t108 9.18308
R20299 vdd.n1504 vdd.t19 8.95635
R20300 vdd.t72 vdd.n3459 8.95635
R20301 vdd.n300 vdd.n299 8.92171
R20302 vdd.n245 vdd.n244 8.92171
R20303 vdd.n202 vdd.n201 8.92171
R20304 vdd.n147 vdd.n146 8.92171
R20305 vdd.n105 vdd.n104 8.92171
R20306 vdd.n50 vdd.n49 8.92171
R20307 vdd.n1749 vdd.n1748 8.92171
R20308 vdd.n1804 vdd.n1803 8.92171
R20309 vdd.n1651 vdd.n1650 8.92171
R20310 vdd.n1706 vdd.n1705 8.92171
R20311 vdd.n1554 vdd.n1553 8.92171
R20312 vdd.n1609 vdd.n1608 8.92171
R20313 vdd.n223 vdd.n125 8.81535
R20314 vdd.n1727 vdd.n1629 8.81535
R20315 vdd.n1184 vdd.t46 8.72962
R20316 vdd.t104 vdd.n3468 8.72962
R20317 vdd.n1840 vdd.t91 8.50289
R20318 vdd.n3387 vdd.t57 8.50289
R20319 vdd.n28 vdd.n14 8.42249
R20320 vdd.n1856 vdd.t67 8.27616
R20321 vdd.t54 vdd.n636 8.27616
R20322 vdd.n3474 vdd.n3473 8.16225
R20323 vdd.n1827 vdd.n1826 8.16225
R20324 vdd.n296 vdd.n290 8.14595
R20325 vdd.n241 vdd.n235 8.14595
R20326 vdd.n198 vdd.n192 8.14595
R20327 vdd.n143 vdd.n137 8.14595
R20328 vdd.n101 vdd.n95 8.14595
R20329 vdd.n46 vdd.n40 8.14595
R20330 vdd.n1745 vdd.n1739 8.14595
R20331 vdd.n1800 vdd.n1794 8.14595
R20332 vdd.n1647 vdd.n1641 8.14595
R20333 vdd.n1702 vdd.n1696 8.14595
R20334 vdd.n1550 vdd.n1544 8.14595
R20335 vdd.n1605 vdd.n1599 8.14595
R20336 vdd.t178 vdd.n1218 7.8227
R20337 vdd.t160 vdd.n363 7.8227
R20338 vdd.n2384 vdd.n1075 7.70933
R20339 vdd.n2390 vdd.n1075 7.70933
R20340 vdd.n2396 vdd.n1069 7.70933
R20341 vdd.n2396 vdd.n1063 7.70933
R20342 vdd.n2402 vdd.n1063 7.70933
R20343 vdd.n2402 vdd.n1057 7.70933
R20344 vdd.n2408 vdd.n1057 7.70933
R20345 vdd.n2414 vdd.n1051 7.70933
R20346 vdd.n2420 vdd.n1045 7.70933
R20347 vdd.n2426 vdd.n1038 7.70933
R20348 vdd.n2426 vdd.n1041 7.70933
R20349 vdd.n2432 vdd.n1034 7.70933
R20350 vdd.n2439 vdd.n1020 7.70933
R20351 vdd.n2445 vdd.n1020 7.70933
R20352 vdd.n2451 vdd.n1014 7.70933
R20353 vdd.n2457 vdd.n1010 7.70933
R20354 vdd.n2463 vdd.n1004 7.70933
R20355 vdd.n2481 vdd.n986 7.70933
R20356 vdd.n2481 vdd.n979 7.70933
R20357 vdd.n2489 vdd.n979 7.70933
R20358 vdd.n2571 vdd.n963 7.70933
R20359 vdd.n2934 vdd.n917 7.70933
R20360 vdd.n2946 vdd.n898 7.70933
R20361 vdd.n2952 vdd.n898 7.70933
R20362 vdd.n2952 vdd.n901 7.70933
R20363 vdd.n2970 vdd.n882 7.70933
R20364 vdd.n2976 vdd.n876 7.70933
R20365 vdd.n2982 vdd.n872 7.70933
R20366 vdd.n2988 vdd.n859 7.70933
R20367 vdd.n2994 vdd.n859 7.70933
R20368 vdd.n3001 vdd.n852 7.70933
R20369 vdd.n3007 vdd.n845 7.70933
R20370 vdd.n3007 vdd.n848 7.70933
R20371 vdd.n3013 vdd.n841 7.70933
R20372 vdd.n3019 vdd.n835 7.70933
R20373 vdd.n3025 vdd.n822 7.70933
R20374 vdd.n3031 vdd.n822 7.70933
R20375 vdd.n3031 vdd.n814 7.70933
R20376 vdd.n3082 vdd.n814 7.70933
R20377 vdd.n3082 vdd.n817 7.70933
R20378 vdd.n3088 vdd.n774 7.70933
R20379 vdd.n3158 vdd.n774 7.70933
R20380 vdd.t253 vdd.n1051 7.59597
R20381 vdd.n2263 vdd.t269 7.59597
R20382 vdd.n2906 vdd.t223 7.59597
R20383 vdd.n835 vdd.t252 7.59597
R20384 vdd.n295 vdd.n292 7.3702
R20385 vdd.n240 vdd.n237 7.3702
R20386 vdd.n197 vdd.n194 7.3702
R20387 vdd.n142 vdd.n139 7.3702
R20388 vdd.n100 vdd.n97 7.3702
R20389 vdd.n45 vdd.n42 7.3702
R20390 vdd.n1744 vdd.n1741 7.3702
R20391 vdd.n1799 vdd.n1796 7.3702
R20392 vdd.n1646 vdd.n1643 7.3702
R20393 vdd.n1701 vdd.n1698 7.3702
R20394 vdd.n1549 vdd.n1546 7.3702
R20395 vdd.n1604 vdd.n1601 7.3702
R20396 vdd.n1387 vdd.n1386 6.98232
R20397 vdd.n2036 vdd.n2035 6.98232
R20398 vdd.n547 vdd.n546 6.98232
R20399 vdd.n3242 vdd.n3241 6.98232
R20400 vdd.n1874 vdd.t25 6.91577
R20401 vdd.n2420 vdd.t260 6.91577
R20402 vdd.n3013 vdd.t268 6.91577
R20403 vdd.n3351 vdd.t21 6.91577
R20404 vdd.n2998 vdd.n2997 6.86879
R20405 vdd.n2436 vdd.n2435 6.86879
R20406 vdd.n2496 vdd.t240 6.80241
R20407 vdd.n2940 vdd.t238 6.80241
R20408 vdd.t50 vdd.n1155 6.68904
R20409 vdd.n3367 vdd.t84 6.68904
R20410 vdd.n1832 vdd.t23 6.46231
R20411 vdd.n3395 vdd.t38 6.46231
R20412 vdd.n2263 vdd.t246 6.34895
R20413 vdd.n2906 vdd.t244 6.34895
R20414 vdd.n3474 vdd.n321 6.32949
R20415 vdd.n1826 vdd.n1825 6.32949
R20416 vdd.t15 vdd.n1183 6.23558
R20417 vdd.t82 vdd.n332 6.23558
R20418 vdd.n1496 vdd.t89 6.00885
R20419 vdd.t249 vdd.n1014 6.00885
R20420 vdd.n872 vdd.t263 6.00885
R20421 vdd.n3453 vdd.t61 6.00885
R20422 vdd.n296 vdd.n295 5.81868
R20423 vdd.n241 vdd.n240 5.81868
R20424 vdd.n198 vdd.n197 5.81868
R20425 vdd.n143 vdd.n142 5.81868
R20426 vdd.n101 vdd.n100 5.81868
R20427 vdd.n46 vdd.n45 5.81868
R20428 vdd.n1745 vdd.n1744 5.81868
R20429 vdd.n1800 vdd.n1799 5.81868
R20430 vdd.n1647 vdd.n1646 5.81868
R20431 vdd.n1702 vdd.n1701 5.81868
R20432 vdd.n1550 vdd.n1549 5.81868
R20433 vdd.n1605 vdd.n1604 5.81868
R20434 vdd.n2579 vdd.n2578 5.77611
R20435 vdd.n2319 vdd.n2318 5.77611
R20436 vdd.n2808 vdd.n2807 5.77611
R20437 vdd.n3097 vdd.n806 5.77611
R20438 vdd.n3163 vdd.n770 5.77611
R20439 vdd.n2744 vdd.n2680 5.77611
R20440 vdd.n2504 vdd.n970 5.77611
R20441 vdd.n2195 vdd.n2194 5.77611
R20442 vdd.n1456 vdd.n1230 5.62474
R20443 vdd.n2119 vdd.n2116 5.62474
R20444 vdd.n3432 vdd.n407 5.62474
R20445 vdd.n3197 vdd.n3194 5.62474
R20446 vdd.n2457 vdd.t255 5.44203
R20447 vdd.n2976 vdd.t266 5.44203
R20448 vdd.n1206 vdd.t89 5.32866
R20449 vdd.t61 vdd.n3452 5.32866
R20450 vdd.n1512 vdd.t15 5.10193
R20451 vdd.n2432 vdd.t259 5.10193
R20452 vdd.n2451 vdd.t141 5.10193
R20453 vdd.n2982 vdd.t254 5.10193
R20454 vdd.n3001 vdd.t220 5.10193
R20455 vdd.n3461 vdd.t82 5.10193
R20456 vdd.n299 vdd.n290 5.04292
R20457 vdd.n244 vdd.n235 5.04292
R20458 vdd.n201 vdd.n192 5.04292
R20459 vdd.n146 vdd.n137 5.04292
R20460 vdd.n104 vdd.n95 5.04292
R20461 vdd.n49 vdd.n40 5.04292
R20462 vdd.n1748 vdd.n1739 5.04292
R20463 vdd.n1803 vdd.n1794 5.04292
R20464 vdd.n1650 vdd.n1641 5.04292
R20465 vdd.n1705 vdd.n1696 5.04292
R20466 vdd.n1553 vdd.n1544 5.04292
R20467 vdd.n1608 vdd.n1599 5.04292
R20468 vdd.n1034 vdd.t205 4.98857
R20469 vdd.t164 vdd.n852 4.98857
R20470 vdd.n1528 vdd.t23 4.8752
R20471 vdd.t153 vdd.n1069 4.8752
R20472 vdd.t257 vdd.t9 4.8752
R20473 vdd.n2251 vdd.t191 4.8752
R20474 vdd.n2918 vdd.t195 4.8752
R20475 vdd.t139 vdd.t232 4.8752
R20476 vdd.n817 vdd.t149 4.8752
R20477 vdd.t38 vdd.n328 4.8752
R20478 vdd.n2580 vdd.n2579 4.83952
R20479 vdd.n2320 vdd.n2319 4.83952
R20480 vdd.n2807 vdd.n2806 4.83952
R20481 vdd.n806 vdd.n801 4.83952
R20482 vdd.n770 vdd.n765 4.83952
R20483 vdd.n2741 vdd.n2680 4.83952
R20484 vdd.n2507 vdd.n970 4.83952
R20485 vdd.n2194 vdd.n2193 4.83952
R20486 vdd.n2475 vdd.t235 4.76184
R20487 vdd.n2958 vdd.t6 4.76184
R20488 vdd.n2004 vdd.n1116 4.74817
R20489 vdd.n1999 vdd.n1117 4.74817
R20490 vdd.n1901 vdd.n1898 4.74817
R20491 vdd.n2100 vdd.n1902 4.74817
R20492 vdd.n2102 vdd.n1901 4.74817
R20493 vdd.n2101 vdd.n2100 4.74817
R20494 vdd.n664 vdd.n662 4.74817
R20495 vdd.n3312 vdd.n665 4.74817
R20496 vdd.n3315 vdd.n665 4.74817
R20497 vdd.n3316 vdd.n664 4.74817
R20498 vdd.n3204 vdd.n749 4.74817
R20499 vdd.n3200 vdd.n751 4.74817
R20500 vdd.n3203 vdd.n751 4.74817
R20501 vdd.n3208 vdd.n749 4.74817
R20502 vdd.n2000 vdd.n1116 4.74817
R20503 vdd.n1119 vdd.n1117 4.74817
R20504 vdd.n321 vdd.n320 4.7074
R20505 vdd.n223 vdd.n222 4.7074
R20506 vdd.n1825 vdd.n1824 4.7074
R20507 vdd.n1727 vdd.n1726 4.7074
R20508 vdd.n1848 vdd.t50 4.64847
R20509 vdd.n3376 vdd.t84 4.64847
R20510 vdd.n1149 vdd.t25 4.42174
R20511 vdd.t21 vdd.n635 4.42174
R20512 vdd.n2251 vdd.t264 4.30838
R20513 vdd.n2918 vdd.t221 4.30838
R20514 vdd.n300 vdd.n288 4.26717
R20515 vdd.n245 vdd.n233 4.26717
R20516 vdd.n202 vdd.n190 4.26717
R20517 vdd.n147 vdd.n135 4.26717
R20518 vdd.n105 vdd.n93 4.26717
R20519 vdd.n50 vdd.n38 4.26717
R20520 vdd.n1749 vdd.n1737 4.26717
R20521 vdd.n1804 vdd.n1792 4.26717
R20522 vdd.n1651 vdd.n1639 4.26717
R20523 vdd.n1706 vdd.n1694 4.26717
R20524 vdd.n1554 vdd.n1542 4.26717
R20525 vdd.n1609 vdd.n1597 4.26717
R20526 vdd.t261 vdd.n1045 4.19501
R20527 vdd.n1004 vdd.t8 4.19501
R20528 vdd.t258 vdd.n882 4.19501
R20529 vdd.n841 vdd.t237 4.19501
R20530 vdd.n321 vdd.n223 4.10845
R20531 vdd.n1825 vdd.n1727 4.10845
R20532 vdd.n277 vdd.t79 4.06363
R20533 vdd.n277 vdd.t119 4.06363
R20534 vdd.n275 vdd.t122 4.06363
R20535 vdd.n275 vdd.t18 4.06363
R20536 vdd.n273 vdd.t45 4.06363
R20537 vdd.n273 vdd.t98 4.06363
R20538 vdd.n271 vdd.t121 4.06363
R20539 vdd.n271 vdd.t131 4.06363
R20540 vdd.n269 vdd.t134 4.06363
R20541 vdd.n269 vdd.t52 4.06363
R20542 vdd.n267 vdd.t77 4.06363
R20543 vdd.n267 vdd.t133 4.06363
R20544 vdd.n265 vdd.t135 4.06363
R20545 vdd.n265 vdd.t76 4.06363
R20546 vdd.n179 vdd.t62 4.06363
R20547 vdd.n179 vdd.t109 4.06363
R20548 vdd.n177 vdd.t110 4.06363
R20549 vdd.n177 vdd.t132 4.06363
R20550 vdd.n175 vdd.t28 4.06363
R20551 vdd.n175 vdd.t83 4.06363
R20552 vdd.n173 vdd.t113 4.06363
R20553 vdd.n173 vdd.t123 4.06363
R20554 vdd.n171 vdd.t126 4.06363
R20555 vdd.n171 vdd.t32 4.06363
R20556 vdd.n169 vdd.t56 4.06363
R20557 vdd.n169 vdd.t114 4.06363
R20558 vdd.n167 vdd.t127 4.06363
R20559 vdd.n167 vdd.t55 4.06363
R20560 vdd.n82 vdd.t88 4.06363
R20561 vdd.n82 vdd.t111 4.06363
R20562 vdd.n80 vdd.t73 4.06363
R20563 vdd.n80 vdd.t128 4.06363
R20564 vdd.n78 vdd.t44 4.06363
R20565 vdd.n78 vdd.t120 4.06363
R20566 vdd.n76 vdd.t39 4.06363
R20567 vdd.n76 vdd.t105 4.06363
R20568 vdd.n74 vdd.t58 4.06363
R20569 vdd.n74 vdd.t124 4.06363
R20570 vdd.n72 vdd.t34 4.06363
R20571 vdd.n72 vdd.t85 4.06363
R20572 vdd.n70 vdd.t22 4.06363
R20573 vdd.n70 vdd.t65 4.06363
R20574 vdd.n1769 vdd.t115 4.06363
R20575 vdd.n1769 vdd.t75 4.06363
R20576 vdd.n1771 vdd.t71 4.06363
R20577 vdd.n1771 vdd.t116 4.06363
R20578 vdd.n1773 vdd.t101 4.06363
R20579 vdd.n1773 vdd.t100 4.06363
R20580 vdd.n1775 vdd.t66 4.06363
R20581 vdd.n1775 vdd.t43 4.06363
R20582 vdd.n1777 vdd.t41 4.06363
R20583 vdd.n1777 vdd.t99 4.06363
R20584 vdd.n1779 vdd.t81 4.06363
R20585 vdd.n1779 vdd.t42 4.06363
R20586 vdd.n1781 vdd.t35 4.06363
R20587 vdd.n1781 vdd.t117 4.06363
R20588 vdd.n1671 vdd.t102 4.06363
R20589 vdd.n1671 vdd.t53 4.06363
R20590 vdd.n1673 vdd.t51 4.06363
R20591 vdd.n1673 vdd.t103 4.06363
R20592 vdd.n1675 vdd.t94 4.06363
R20593 vdd.n1675 vdd.t92 4.06363
R20594 vdd.n1677 vdd.t47 4.06363
R20595 vdd.n1677 vdd.t24 4.06363
R20596 vdd.n1679 vdd.t16 4.06363
R20597 vdd.n1679 vdd.t87 4.06363
R20598 vdd.n1681 vdd.t70 4.06363
R20599 vdd.n1681 vdd.t20 4.06363
R20600 vdd.n1683 vdd.t12 4.06363
R20601 vdd.n1683 vdd.t107 4.06363
R20602 vdd.n1574 vdd.t68 4.06363
R20603 vdd.n1574 vdd.t26 4.06363
R20604 vdd.n1576 vdd.t86 4.06363
R20605 vdd.n1576 vdd.t37 4.06363
R20606 vdd.n1578 vdd.t125 4.06363
R20607 vdd.n1578 vdd.t136 4.06363
R20608 vdd.n1580 vdd.t106 4.06363
R20609 vdd.n1580 vdd.t40 4.06363
R20610 vdd.n1582 vdd.t97 4.06363
R20611 vdd.n1582 vdd.t49 4.06363
R20612 vdd.n1584 vdd.t129 4.06363
R20613 vdd.n1584 vdd.t74 4.06363
R20614 vdd.n1586 vdd.t112 4.06363
R20615 vdd.n1586 vdd.t90 4.06363
R20616 vdd.n26 vdd.t5 3.9605
R20617 vdd.n26 vdd.t0 3.9605
R20618 vdd.n23 vdd.t229 3.9605
R20619 vdd.n23 vdd.t3 3.9605
R20620 vdd.n21 vdd.t226 3.9605
R20621 vdd.n21 vdd.t271 3.9605
R20622 vdd.n20 vdd.t4 3.9605
R20623 vdd.n20 vdd.t228 3.9605
R20624 vdd.n15 vdd.t225 3.9605
R20625 vdd.n15 vdd.t142 3.9605
R20626 vdd.n16 vdd.t2 3.9605
R20627 vdd.n16 vdd.t227 3.9605
R20628 vdd.n18 vdd.t1 3.9605
R20629 vdd.n18 vdd.t143 3.9605
R20630 vdd.n25 vdd.t224 3.9605
R20631 vdd.n25 vdd.t270 3.9605
R20632 vdd.n2997 vdd.n2996 3.74684
R20633 vdd.n2437 vdd.n2436 3.74684
R20634 vdd.n7 vdd.t140 3.61217
R20635 vdd.n7 vdd.t267 3.61217
R20636 vdd.n8 vdd.t7 3.61217
R20637 vdd.n8 vdd.t245 3.61217
R20638 vdd.n10 vdd.t239 3.61217
R20639 vdd.n10 vdd.t222 3.61217
R20640 vdd.n12 vdd.t251 3.61217
R20641 vdd.n12 vdd.t231 3.61217
R20642 vdd.n5 vdd.t243 3.61217
R20643 vdd.n5 vdd.t234 3.61217
R20644 vdd.n3 vdd.t265 3.61217
R20645 vdd.n3 vdd.t241 3.61217
R20646 vdd.n1 vdd.t247 3.61217
R20647 vdd.n1 vdd.t236 3.61217
R20648 vdd.n0 vdd.t256 3.61217
R20649 vdd.n0 vdd.t10 3.61217
R20650 vdd.n1462 vdd.t178 3.51482
R20651 vdd.n2414 vdd.t261 3.51482
R20652 vdd.n2469 vdd.t8 3.51482
R20653 vdd.n2964 vdd.t258 3.51482
R20654 vdd.n3019 vdd.t237 3.51482
R20655 vdd.n3437 vdd.t160 3.51482
R20656 vdd.n304 vdd.n303 3.49141
R20657 vdd.n249 vdd.n248 3.49141
R20658 vdd.n206 vdd.n205 3.49141
R20659 vdd.n151 vdd.n150 3.49141
R20660 vdd.n109 vdd.n108 3.49141
R20661 vdd.n54 vdd.n53 3.49141
R20662 vdd.n1753 vdd.n1752 3.49141
R20663 vdd.n1808 vdd.n1807 3.49141
R20664 vdd.n1655 vdd.n1654 3.49141
R20665 vdd.n1710 vdd.n1709 3.49141
R20666 vdd.n1558 vdd.n1557 3.49141
R20667 vdd.n1613 vdd.n1612 3.49141
R20668 vdd.n2489 vdd.t264 3.40145
R20669 vdd.n2643 vdd.t242 3.40145
R20670 vdd.n2927 vdd.t230 3.40145
R20671 vdd.n2946 vdd.t221 3.40145
R20672 vdd.n1865 vdd.t67 3.06136
R20673 vdd.n3359 vdd.t54 3.06136
R20674 vdd.t235 vdd.n986 2.94799
R20675 vdd.n901 vdd.t6 2.94799
R20676 vdd.t91 vdd.n1161 2.83463
R20677 vdd.n2390 vdd.t153 2.83463
R20678 vdd.n2496 vdd.t191 2.83463
R20679 vdd.n2940 vdd.t195 2.83463
R20680 vdd.n3088 vdd.t149 2.83463
R20681 vdd.n624 vdd.t57 2.83463
R20682 vdd.n307 vdd.n286 2.71565
R20683 vdd.n252 vdd.n231 2.71565
R20684 vdd.n209 vdd.n188 2.71565
R20685 vdd.n154 vdd.n133 2.71565
R20686 vdd.n112 vdd.n91 2.71565
R20687 vdd.n57 vdd.n36 2.71565
R20688 vdd.n1756 vdd.n1735 2.71565
R20689 vdd.n1811 vdd.n1790 2.71565
R20690 vdd.n1658 vdd.n1637 2.71565
R20691 vdd.n1713 vdd.n1692 2.71565
R20692 vdd.n1561 vdd.n1540 2.71565
R20693 vdd.n1616 vdd.n1595 2.71565
R20694 vdd.n1529 vdd.t46 2.6079
R20695 vdd.n1041 vdd.t259 2.6079
R20696 vdd.n2275 vdd.t141 2.6079
R20697 vdd.n2894 vdd.t254 2.6079
R20698 vdd.t220 vdd.n845 2.6079
R20699 vdd.n3469 vdd.t104 2.6079
R20700 vdd.n294 vdd.n293 2.4129
R20701 vdd.n239 vdd.n238 2.4129
R20702 vdd.n196 vdd.n195 2.4129
R20703 vdd.n141 vdd.n140 2.4129
R20704 vdd.n99 vdd.n98 2.4129
R20705 vdd.n44 vdd.n43 2.4129
R20706 vdd.n1743 vdd.n1742 2.4129
R20707 vdd.n1798 vdd.n1797 2.4129
R20708 vdd.n1645 vdd.n1644 2.4129
R20709 vdd.n1700 vdd.n1699 2.4129
R20710 vdd.n1548 vdd.n1547 2.4129
R20711 vdd.n1603 vdd.n1602 2.4129
R20712 vdd.t19 vdd.n1190 2.38117
R20713 vdd.n3460 vdd.t72 2.38117
R20714 vdd.n2099 vdd.n1901 2.27742
R20715 vdd.n2100 vdd.n2099 2.27742
R20716 vdd.n3124 vdd.n665 2.27742
R20717 vdd.n3124 vdd.n664 2.27742
R20718 vdd.n3192 vdd.n751 2.27742
R20719 vdd.n3192 vdd.n749 2.27742
R20720 vdd.n2122 vdd.n1116 2.27742
R20721 vdd.n2122 vdd.n1117 2.27742
R20722 vdd.n2275 vdd.t255 2.2678
R20723 vdd.n2894 vdd.t266 2.2678
R20724 vdd.n1487 vdd.t11 2.15444
R20725 vdd.n3451 vdd.t108 2.15444
R20726 vdd.n2463 vdd.t9 2.04107
R20727 vdd.n2970 vdd.t139 2.04107
R20728 vdd.n308 vdd.n284 1.93989
R20729 vdd.n253 vdd.n229 1.93989
R20730 vdd.n210 vdd.n186 1.93989
R20731 vdd.n155 vdd.n131 1.93989
R20732 vdd.n113 vdd.n89 1.93989
R20733 vdd.n58 vdd.n34 1.93989
R20734 vdd.n1757 vdd.n1733 1.93989
R20735 vdd.n1812 vdd.n1788 1.93989
R20736 vdd.n1659 vdd.n1635 1.93989
R20737 vdd.n1714 vdd.n1690 1.93989
R20738 vdd.n1562 vdd.n1538 1.93989
R20739 vdd.n1617 vdd.n1593 1.93989
R20740 vdd.n1479 vdd.t13 1.70098
R20741 vdd.n2439 vdd.t248 1.70098
R20742 vdd.n2445 vdd.t249 1.70098
R20743 vdd.n2988 vdd.t263 1.70098
R20744 vdd.n2994 vdd.t262 1.70098
R20745 vdd.n3445 vdd.t29 1.70098
R20746 vdd.n1495 vdd.t69 1.47425
R20747 vdd.n349 vdd.t17 1.47425
R20748 vdd.n2469 vdd.t246 1.36088
R20749 vdd.n2964 vdd.t244 1.36088
R20750 vdd.n1520 vdd.t48 1.24752
R20751 vdd.t171 vdd.n1124 1.24752
R20752 vdd.n659 vdd.t145 1.24752
R20753 vdd.t27 vdd.n3467 1.24752
R20754 vdd.n319 vdd.n279 1.16414
R20755 vdd.n312 vdd.n311 1.16414
R20756 vdd.n264 vdd.n224 1.16414
R20757 vdd.n257 vdd.n256 1.16414
R20758 vdd.n221 vdd.n181 1.16414
R20759 vdd.n214 vdd.n213 1.16414
R20760 vdd.n166 vdd.n126 1.16414
R20761 vdd.n159 vdd.n158 1.16414
R20762 vdd.n124 vdd.n84 1.16414
R20763 vdd.n117 vdd.n116 1.16414
R20764 vdd.n69 vdd.n29 1.16414
R20765 vdd.n62 vdd.n61 1.16414
R20766 vdd.n1768 vdd.n1728 1.16414
R20767 vdd.n1761 vdd.n1760 1.16414
R20768 vdd.n1823 vdd.n1783 1.16414
R20769 vdd.n1816 vdd.n1815 1.16414
R20770 vdd.n1670 vdd.n1630 1.16414
R20771 vdd.n1663 vdd.n1662 1.16414
R20772 vdd.n1725 vdd.n1685 1.16414
R20773 vdd.n1718 vdd.n1717 1.16414
R20774 vdd.n1573 vdd.n1533 1.16414
R20775 vdd.n1566 vdd.n1565 1.16414
R20776 vdd.n1628 vdd.n1588 1.16414
R20777 vdd.n1621 vdd.n1620 1.16414
R20778 vdd.n1826 vdd.n28 1.06035
R20779 vdd vdd.n3474 1.05252
R20780 vdd.n1172 vdd.t93 1.02079
R20781 vdd.t205 vdd.t248 1.02079
R20782 vdd.t262 vdd.t164 1.02079
R20783 vdd.t31 vdd.n613 1.02079
R20784 vdd.n1351 vdd.n1230 0.970197
R20785 vdd.n2120 vdd.n2119 0.970197
R20786 vdd.n599 vdd.n407 0.970197
R20787 vdd.n3199 vdd.n3197 0.970197
R20788 vdd.t240 vdd.n963 0.907421
R20789 vdd.n917 vdd.t238 0.907421
R20790 vdd.n1857 vdd.t36 0.794056
R20791 vdd.t260 vdd.n1038 0.794056
R20792 vdd.n1010 vdd.t257 0.794056
R20793 vdd.t232 vdd.n876 0.794056
R20794 vdd.n848 vdd.t268 0.794056
R20795 vdd.n3368 vdd.t33 0.794056
R20796 vdd.n1873 vdd.t95 0.567326
R20797 vdd.t63 vdd.n642 0.567326
R20798 vdd.n2110 vdd.n2109 0.482207
R20799 vdd.n3324 vdd.n3323 0.482207
R20800 vdd.n444 vdd.n443 0.482207
R20801 vdd.n3431 vdd.n3430 0.482207
R20802 vdd.n3330 vdd.n656 0.482207
R20803 vdd.n1887 vdd.n1118 0.482207
R20804 vdd.n1458 vdd.n1457 0.482207
R20805 vdd.n1264 vdd.n1221 0.482207
R20806 vdd.n4 vdd.n2 0.459552
R20807 vdd.n11 vdd.n9 0.459552
R20808 vdd.n317 vdd.n316 0.388379
R20809 vdd.n283 vdd.n281 0.388379
R20810 vdd.n262 vdd.n261 0.388379
R20811 vdd.n228 vdd.n226 0.388379
R20812 vdd.n219 vdd.n218 0.388379
R20813 vdd.n185 vdd.n183 0.388379
R20814 vdd.n164 vdd.n163 0.388379
R20815 vdd.n130 vdd.n128 0.388379
R20816 vdd.n122 vdd.n121 0.388379
R20817 vdd.n88 vdd.n86 0.388379
R20818 vdd.n67 vdd.n66 0.388379
R20819 vdd.n33 vdd.n31 0.388379
R20820 vdd.n1766 vdd.n1765 0.388379
R20821 vdd.n1732 vdd.n1730 0.388379
R20822 vdd.n1821 vdd.n1820 0.388379
R20823 vdd.n1787 vdd.n1785 0.388379
R20824 vdd.n1668 vdd.n1667 0.388379
R20825 vdd.n1634 vdd.n1632 0.388379
R20826 vdd.n1723 vdd.n1722 0.388379
R20827 vdd.n1689 vdd.n1687 0.388379
R20828 vdd.n1571 vdd.n1570 0.388379
R20829 vdd.n1537 vdd.n1535 0.388379
R20830 vdd.n1626 vdd.n1625 0.388379
R20831 vdd.n1592 vdd.n1590 0.388379
R20832 vdd.n19 vdd.n17 0.387128
R20833 vdd.n24 vdd.n22 0.387128
R20834 vdd.n6 vdd.n4 0.358259
R20835 vdd.n13 vdd.n11 0.358259
R20836 vdd.n268 vdd.n266 0.358259
R20837 vdd.n270 vdd.n268 0.358259
R20838 vdd.n272 vdd.n270 0.358259
R20839 vdd.n274 vdd.n272 0.358259
R20840 vdd.n276 vdd.n274 0.358259
R20841 vdd.n278 vdd.n276 0.358259
R20842 vdd.n320 vdd.n278 0.358259
R20843 vdd.n170 vdd.n168 0.358259
R20844 vdd.n172 vdd.n170 0.358259
R20845 vdd.n174 vdd.n172 0.358259
R20846 vdd.n176 vdd.n174 0.358259
R20847 vdd.n178 vdd.n176 0.358259
R20848 vdd.n180 vdd.n178 0.358259
R20849 vdd.n222 vdd.n180 0.358259
R20850 vdd.n73 vdd.n71 0.358259
R20851 vdd.n75 vdd.n73 0.358259
R20852 vdd.n77 vdd.n75 0.358259
R20853 vdd.n79 vdd.n77 0.358259
R20854 vdd.n81 vdd.n79 0.358259
R20855 vdd.n83 vdd.n81 0.358259
R20856 vdd.n125 vdd.n83 0.358259
R20857 vdd.n1824 vdd.n1782 0.358259
R20858 vdd.n1782 vdd.n1780 0.358259
R20859 vdd.n1780 vdd.n1778 0.358259
R20860 vdd.n1778 vdd.n1776 0.358259
R20861 vdd.n1776 vdd.n1774 0.358259
R20862 vdd.n1774 vdd.n1772 0.358259
R20863 vdd.n1772 vdd.n1770 0.358259
R20864 vdd.n1726 vdd.n1684 0.358259
R20865 vdd.n1684 vdd.n1682 0.358259
R20866 vdd.n1682 vdd.n1680 0.358259
R20867 vdd.n1680 vdd.n1678 0.358259
R20868 vdd.n1678 vdd.n1676 0.358259
R20869 vdd.n1676 vdd.n1674 0.358259
R20870 vdd.n1674 vdd.n1672 0.358259
R20871 vdd.n1629 vdd.n1587 0.358259
R20872 vdd.n1587 vdd.n1585 0.358259
R20873 vdd.n1585 vdd.n1583 0.358259
R20874 vdd.n1583 vdd.n1581 0.358259
R20875 vdd.n1581 vdd.n1579 0.358259
R20876 vdd.n1579 vdd.n1577 0.358259
R20877 vdd.n1577 vdd.n1575 0.358259
R20878 vdd.n14 vdd.n6 0.334552
R20879 vdd.n14 vdd.n13 0.334552
R20880 vdd.n27 vdd.n19 0.21707
R20881 vdd.n27 vdd.n24 0.21707
R20882 vdd.n318 vdd.n280 0.155672
R20883 vdd.n310 vdd.n280 0.155672
R20884 vdd.n310 vdd.n309 0.155672
R20885 vdd.n309 vdd.n285 0.155672
R20886 vdd.n302 vdd.n285 0.155672
R20887 vdd.n302 vdd.n301 0.155672
R20888 vdd.n301 vdd.n289 0.155672
R20889 vdd.n294 vdd.n289 0.155672
R20890 vdd.n263 vdd.n225 0.155672
R20891 vdd.n255 vdd.n225 0.155672
R20892 vdd.n255 vdd.n254 0.155672
R20893 vdd.n254 vdd.n230 0.155672
R20894 vdd.n247 vdd.n230 0.155672
R20895 vdd.n247 vdd.n246 0.155672
R20896 vdd.n246 vdd.n234 0.155672
R20897 vdd.n239 vdd.n234 0.155672
R20898 vdd.n220 vdd.n182 0.155672
R20899 vdd.n212 vdd.n182 0.155672
R20900 vdd.n212 vdd.n211 0.155672
R20901 vdd.n211 vdd.n187 0.155672
R20902 vdd.n204 vdd.n187 0.155672
R20903 vdd.n204 vdd.n203 0.155672
R20904 vdd.n203 vdd.n191 0.155672
R20905 vdd.n196 vdd.n191 0.155672
R20906 vdd.n165 vdd.n127 0.155672
R20907 vdd.n157 vdd.n127 0.155672
R20908 vdd.n157 vdd.n156 0.155672
R20909 vdd.n156 vdd.n132 0.155672
R20910 vdd.n149 vdd.n132 0.155672
R20911 vdd.n149 vdd.n148 0.155672
R20912 vdd.n148 vdd.n136 0.155672
R20913 vdd.n141 vdd.n136 0.155672
R20914 vdd.n123 vdd.n85 0.155672
R20915 vdd.n115 vdd.n85 0.155672
R20916 vdd.n115 vdd.n114 0.155672
R20917 vdd.n114 vdd.n90 0.155672
R20918 vdd.n107 vdd.n90 0.155672
R20919 vdd.n107 vdd.n106 0.155672
R20920 vdd.n106 vdd.n94 0.155672
R20921 vdd.n99 vdd.n94 0.155672
R20922 vdd.n68 vdd.n30 0.155672
R20923 vdd.n60 vdd.n30 0.155672
R20924 vdd.n60 vdd.n59 0.155672
R20925 vdd.n59 vdd.n35 0.155672
R20926 vdd.n52 vdd.n35 0.155672
R20927 vdd.n52 vdd.n51 0.155672
R20928 vdd.n51 vdd.n39 0.155672
R20929 vdd.n44 vdd.n39 0.155672
R20930 vdd.n1767 vdd.n1729 0.155672
R20931 vdd.n1759 vdd.n1729 0.155672
R20932 vdd.n1759 vdd.n1758 0.155672
R20933 vdd.n1758 vdd.n1734 0.155672
R20934 vdd.n1751 vdd.n1734 0.155672
R20935 vdd.n1751 vdd.n1750 0.155672
R20936 vdd.n1750 vdd.n1738 0.155672
R20937 vdd.n1743 vdd.n1738 0.155672
R20938 vdd.n1822 vdd.n1784 0.155672
R20939 vdd.n1814 vdd.n1784 0.155672
R20940 vdd.n1814 vdd.n1813 0.155672
R20941 vdd.n1813 vdd.n1789 0.155672
R20942 vdd.n1806 vdd.n1789 0.155672
R20943 vdd.n1806 vdd.n1805 0.155672
R20944 vdd.n1805 vdd.n1793 0.155672
R20945 vdd.n1798 vdd.n1793 0.155672
R20946 vdd.n1669 vdd.n1631 0.155672
R20947 vdd.n1661 vdd.n1631 0.155672
R20948 vdd.n1661 vdd.n1660 0.155672
R20949 vdd.n1660 vdd.n1636 0.155672
R20950 vdd.n1653 vdd.n1636 0.155672
R20951 vdd.n1653 vdd.n1652 0.155672
R20952 vdd.n1652 vdd.n1640 0.155672
R20953 vdd.n1645 vdd.n1640 0.155672
R20954 vdd.n1724 vdd.n1686 0.155672
R20955 vdd.n1716 vdd.n1686 0.155672
R20956 vdd.n1716 vdd.n1715 0.155672
R20957 vdd.n1715 vdd.n1691 0.155672
R20958 vdd.n1708 vdd.n1691 0.155672
R20959 vdd.n1708 vdd.n1707 0.155672
R20960 vdd.n1707 vdd.n1695 0.155672
R20961 vdd.n1700 vdd.n1695 0.155672
R20962 vdd.n1572 vdd.n1534 0.155672
R20963 vdd.n1564 vdd.n1534 0.155672
R20964 vdd.n1564 vdd.n1563 0.155672
R20965 vdd.n1563 vdd.n1539 0.155672
R20966 vdd.n1556 vdd.n1539 0.155672
R20967 vdd.n1556 vdd.n1555 0.155672
R20968 vdd.n1555 vdd.n1543 0.155672
R20969 vdd.n1548 vdd.n1543 0.155672
R20970 vdd.n1627 vdd.n1589 0.155672
R20971 vdd.n1619 vdd.n1589 0.155672
R20972 vdd.n1619 vdd.n1618 0.155672
R20973 vdd.n1618 vdd.n1594 0.155672
R20974 vdd.n1611 vdd.n1594 0.155672
R20975 vdd.n1611 vdd.n1610 0.155672
R20976 vdd.n1610 vdd.n1598 0.155672
R20977 vdd.n1603 vdd.n1598 0.155672
R20978 vdd.n2098 vdd.n1903 0.152939
R20979 vdd.n1909 vdd.n1903 0.152939
R20980 vdd.n1910 vdd.n1909 0.152939
R20981 vdd.n1911 vdd.n1910 0.152939
R20982 vdd.n1912 vdd.n1911 0.152939
R20983 vdd.n1916 vdd.n1912 0.152939
R20984 vdd.n1917 vdd.n1916 0.152939
R20985 vdd.n1918 vdd.n1917 0.152939
R20986 vdd.n1919 vdd.n1918 0.152939
R20987 vdd.n1923 vdd.n1919 0.152939
R20988 vdd.n1924 vdd.n1923 0.152939
R20989 vdd.n1925 vdd.n1924 0.152939
R20990 vdd.n2073 vdd.n1925 0.152939
R20991 vdd.n2073 vdd.n2072 0.152939
R20992 vdd.n2072 vdd.n2071 0.152939
R20993 vdd.n2071 vdd.n1931 0.152939
R20994 vdd.n1936 vdd.n1931 0.152939
R20995 vdd.n1937 vdd.n1936 0.152939
R20996 vdd.n1938 vdd.n1937 0.152939
R20997 vdd.n1942 vdd.n1938 0.152939
R20998 vdd.n1943 vdd.n1942 0.152939
R20999 vdd.n1944 vdd.n1943 0.152939
R21000 vdd.n1945 vdd.n1944 0.152939
R21001 vdd.n1949 vdd.n1945 0.152939
R21002 vdd.n1950 vdd.n1949 0.152939
R21003 vdd.n1951 vdd.n1950 0.152939
R21004 vdd.n1952 vdd.n1951 0.152939
R21005 vdd.n1956 vdd.n1952 0.152939
R21006 vdd.n1957 vdd.n1956 0.152939
R21007 vdd.n1958 vdd.n1957 0.152939
R21008 vdd.n1959 vdd.n1958 0.152939
R21009 vdd.n1963 vdd.n1959 0.152939
R21010 vdd.n1964 vdd.n1963 0.152939
R21011 vdd.n1965 vdd.n1964 0.152939
R21012 vdd.n2034 vdd.n1965 0.152939
R21013 vdd.n2034 vdd.n2033 0.152939
R21014 vdd.n2033 vdd.n2032 0.152939
R21015 vdd.n2032 vdd.n1971 0.152939
R21016 vdd.n1976 vdd.n1971 0.152939
R21017 vdd.n1977 vdd.n1976 0.152939
R21018 vdd.n1978 vdd.n1977 0.152939
R21019 vdd.n1982 vdd.n1978 0.152939
R21020 vdd.n1983 vdd.n1982 0.152939
R21021 vdd.n1984 vdd.n1983 0.152939
R21022 vdd.n1985 vdd.n1984 0.152939
R21023 vdd.n1989 vdd.n1985 0.152939
R21024 vdd.n1990 vdd.n1989 0.152939
R21025 vdd.n1991 vdd.n1990 0.152939
R21026 vdd.n1992 vdd.n1991 0.152939
R21027 vdd.n1993 vdd.n1992 0.152939
R21028 vdd.n1993 vdd.n1115 0.152939
R21029 vdd.n2109 vdd.n1897 0.152939
R21030 vdd.n1829 vdd.n1828 0.152939
R21031 vdd.n1829 vdd.n1164 0.152939
R21032 vdd.n1843 vdd.n1164 0.152939
R21033 vdd.n1844 vdd.n1843 0.152939
R21034 vdd.n1845 vdd.n1844 0.152939
R21035 vdd.n1845 vdd.n1152 0.152939
R21036 vdd.n1860 vdd.n1152 0.152939
R21037 vdd.n1861 vdd.n1860 0.152939
R21038 vdd.n1862 vdd.n1861 0.152939
R21039 vdd.n1862 vdd.n1141 0.152939
R21040 vdd.n1877 vdd.n1141 0.152939
R21041 vdd.n1878 vdd.n1877 0.152939
R21042 vdd.n1879 vdd.n1878 0.152939
R21043 vdd.n1879 vdd.n1129 0.152939
R21044 vdd.n1895 vdd.n1129 0.152939
R21045 vdd.n1896 vdd.n1895 0.152939
R21046 vdd.n2110 vdd.n1896 0.152939
R21047 vdd.n670 vdd.n667 0.152939
R21048 vdd.n671 vdd.n670 0.152939
R21049 vdd.n672 vdd.n671 0.152939
R21050 vdd.n673 vdd.n672 0.152939
R21051 vdd.n676 vdd.n673 0.152939
R21052 vdd.n677 vdd.n676 0.152939
R21053 vdd.n678 vdd.n677 0.152939
R21054 vdd.n679 vdd.n678 0.152939
R21055 vdd.n682 vdd.n679 0.152939
R21056 vdd.n683 vdd.n682 0.152939
R21057 vdd.n684 vdd.n683 0.152939
R21058 vdd.n685 vdd.n684 0.152939
R21059 vdd.n690 vdd.n685 0.152939
R21060 vdd.n691 vdd.n690 0.152939
R21061 vdd.n692 vdd.n691 0.152939
R21062 vdd.n693 vdd.n692 0.152939
R21063 vdd.n696 vdd.n693 0.152939
R21064 vdd.n697 vdd.n696 0.152939
R21065 vdd.n698 vdd.n697 0.152939
R21066 vdd.n699 vdd.n698 0.152939
R21067 vdd.n702 vdd.n699 0.152939
R21068 vdd.n703 vdd.n702 0.152939
R21069 vdd.n704 vdd.n703 0.152939
R21070 vdd.n705 vdd.n704 0.152939
R21071 vdd.n708 vdd.n705 0.152939
R21072 vdd.n709 vdd.n708 0.152939
R21073 vdd.n710 vdd.n709 0.152939
R21074 vdd.n711 vdd.n710 0.152939
R21075 vdd.n714 vdd.n711 0.152939
R21076 vdd.n715 vdd.n714 0.152939
R21077 vdd.n716 vdd.n715 0.152939
R21078 vdd.n717 vdd.n716 0.152939
R21079 vdd.n720 vdd.n717 0.152939
R21080 vdd.n721 vdd.n720 0.152939
R21081 vdd.n3240 vdd.n721 0.152939
R21082 vdd.n3240 vdd.n3239 0.152939
R21083 vdd.n3239 vdd.n3238 0.152939
R21084 vdd.n3238 vdd.n725 0.152939
R21085 vdd.n730 vdd.n725 0.152939
R21086 vdd.n731 vdd.n730 0.152939
R21087 vdd.n734 vdd.n731 0.152939
R21088 vdd.n735 vdd.n734 0.152939
R21089 vdd.n736 vdd.n735 0.152939
R21090 vdd.n737 vdd.n736 0.152939
R21091 vdd.n740 vdd.n737 0.152939
R21092 vdd.n741 vdd.n740 0.152939
R21093 vdd.n742 vdd.n741 0.152939
R21094 vdd.n743 vdd.n742 0.152939
R21095 vdd.n746 vdd.n743 0.152939
R21096 vdd.n747 vdd.n746 0.152939
R21097 vdd.n748 vdd.n747 0.152939
R21098 vdd.n3323 vdd.n661 0.152939
R21099 vdd.n3324 vdd.n651 0.152939
R21100 vdd.n3338 vdd.n651 0.152939
R21101 vdd.n3339 vdd.n3338 0.152939
R21102 vdd.n3340 vdd.n3339 0.152939
R21103 vdd.n3340 vdd.n639 0.152939
R21104 vdd.n3354 vdd.n639 0.152939
R21105 vdd.n3355 vdd.n3354 0.152939
R21106 vdd.n3356 vdd.n3355 0.152939
R21107 vdd.n3356 vdd.n627 0.152939
R21108 vdd.n3371 vdd.n627 0.152939
R21109 vdd.n3372 vdd.n3371 0.152939
R21110 vdd.n3373 vdd.n3372 0.152939
R21111 vdd.n3373 vdd.n616 0.152939
R21112 vdd.n3390 vdd.n616 0.152939
R21113 vdd.n3391 vdd.n3390 0.152939
R21114 vdd.n3392 vdd.n3391 0.152939
R21115 vdd.n3392 vdd.n322 0.152939
R21116 vdd.n3472 vdd.n323 0.152939
R21117 vdd.n334 vdd.n323 0.152939
R21118 vdd.n335 vdd.n334 0.152939
R21119 vdd.n336 vdd.n335 0.152939
R21120 vdd.n343 vdd.n336 0.152939
R21121 vdd.n344 vdd.n343 0.152939
R21122 vdd.n345 vdd.n344 0.152939
R21123 vdd.n346 vdd.n345 0.152939
R21124 vdd.n354 vdd.n346 0.152939
R21125 vdd.n355 vdd.n354 0.152939
R21126 vdd.n356 vdd.n355 0.152939
R21127 vdd.n357 vdd.n356 0.152939
R21128 vdd.n365 vdd.n357 0.152939
R21129 vdd.n366 vdd.n365 0.152939
R21130 vdd.n367 vdd.n366 0.152939
R21131 vdd.n368 vdd.n367 0.152939
R21132 vdd.n443 vdd.n368 0.152939
R21133 vdd.n444 vdd.n442 0.152939
R21134 vdd.n451 vdd.n442 0.152939
R21135 vdd.n452 vdd.n451 0.152939
R21136 vdd.n453 vdd.n452 0.152939
R21137 vdd.n453 vdd.n440 0.152939
R21138 vdd.n461 vdd.n440 0.152939
R21139 vdd.n462 vdd.n461 0.152939
R21140 vdd.n463 vdd.n462 0.152939
R21141 vdd.n463 vdd.n438 0.152939
R21142 vdd.n471 vdd.n438 0.152939
R21143 vdd.n472 vdd.n471 0.152939
R21144 vdd.n473 vdd.n472 0.152939
R21145 vdd.n473 vdd.n436 0.152939
R21146 vdd.n481 vdd.n436 0.152939
R21147 vdd.n482 vdd.n481 0.152939
R21148 vdd.n483 vdd.n482 0.152939
R21149 vdd.n483 vdd.n434 0.152939
R21150 vdd.n491 vdd.n434 0.152939
R21151 vdd.n492 vdd.n491 0.152939
R21152 vdd.n493 vdd.n492 0.152939
R21153 vdd.n493 vdd.n430 0.152939
R21154 vdd.n501 vdd.n430 0.152939
R21155 vdd.n502 vdd.n501 0.152939
R21156 vdd.n503 vdd.n502 0.152939
R21157 vdd.n503 vdd.n428 0.152939
R21158 vdd.n511 vdd.n428 0.152939
R21159 vdd.n512 vdd.n511 0.152939
R21160 vdd.n513 vdd.n512 0.152939
R21161 vdd.n513 vdd.n426 0.152939
R21162 vdd.n521 vdd.n426 0.152939
R21163 vdd.n522 vdd.n521 0.152939
R21164 vdd.n523 vdd.n522 0.152939
R21165 vdd.n523 vdd.n424 0.152939
R21166 vdd.n531 vdd.n424 0.152939
R21167 vdd.n532 vdd.n531 0.152939
R21168 vdd.n533 vdd.n532 0.152939
R21169 vdd.n533 vdd.n422 0.152939
R21170 vdd.n541 vdd.n422 0.152939
R21171 vdd.n542 vdd.n541 0.152939
R21172 vdd.n543 vdd.n542 0.152939
R21173 vdd.n543 vdd.n418 0.152939
R21174 vdd.n551 vdd.n418 0.152939
R21175 vdd.n552 vdd.n551 0.152939
R21176 vdd.n553 vdd.n552 0.152939
R21177 vdd.n553 vdd.n416 0.152939
R21178 vdd.n561 vdd.n416 0.152939
R21179 vdd.n562 vdd.n561 0.152939
R21180 vdd.n563 vdd.n562 0.152939
R21181 vdd.n563 vdd.n414 0.152939
R21182 vdd.n571 vdd.n414 0.152939
R21183 vdd.n572 vdd.n571 0.152939
R21184 vdd.n573 vdd.n572 0.152939
R21185 vdd.n573 vdd.n412 0.152939
R21186 vdd.n581 vdd.n412 0.152939
R21187 vdd.n582 vdd.n581 0.152939
R21188 vdd.n583 vdd.n582 0.152939
R21189 vdd.n583 vdd.n410 0.152939
R21190 vdd.n591 vdd.n410 0.152939
R21191 vdd.n592 vdd.n591 0.152939
R21192 vdd.n593 vdd.n592 0.152939
R21193 vdd.n593 vdd.n408 0.152939
R21194 vdd.n600 vdd.n408 0.152939
R21195 vdd.n3431 vdd.n600 0.152939
R21196 vdd.n3331 vdd.n3330 0.152939
R21197 vdd.n3332 vdd.n3331 0.152939
R21198 vdd.n3332 vdd.n645 0.152939
R21199 vdd.n3346 vdd.n645 0.152939
R21200 vdd.n3347 vdd.n3346 0.152939
R21201 vdd.n3348 vdd.n3347 0.152939
R21202 vdd.n3348 vdd.n632 0.152939
R21203 vdd.n3362 vdd.n632 0.152939
R21204 vdd.n3363 vdd.n3362 0.152939
R21205 vdd.n3364 vdd.n3363 0.152939
R21206 vdd.n3364 vdd.n621 0.152939
R21207 vdd.n3379 vdd.n621 0.152939
R21208 vdd.n3380 vdd.n3379 0.152939
R21209 vdd.n3381 vdd.n3380 0.152939
R21210 vdd.n3383 vdd.n3381 0.152939
R21211 vdd.n3383 vdd.n3382 0.152939
R21212 vdd.n3382 vdd.n611 0.152939
R21213 vdd.n611 vdd.n609 0.152939
R21214 vdd.n3401 vdd.n609 0.152939
R21215 vdd.n3402 vdd.n3401 0.152939
R21216 vdd.n3403 vdd.n3402 0.152939
R21217 vdd.n3403 vdd.n607 0.152939
R21218 vdd.n3408 vdd.n607 0.152939
R21219 vdd.n3409 vdd.n3408 0.152939
R21220 vdd.n3410 vdd.n3409 0.152939
R21221 vdd.n3410 vdd.n605 0.152939
R21222 vdd.n3415 vdd.n605 0.152939
R21223 vdd.n3416 vdd.n3415 0.152939
R21224 vdd.n3417 vdd.n3416 0.152939
R21225 vdd.n3417 vdd.n603 0.152939
R21226 vdd.n3423 vdd.n603 0.152939
R21227 vdd.n3424 vdd.n3423 0.152939
R21228 vdd.n3425 vdd.n3424 0.152939
R21229 vdd.n3425 vdd.n601 0.152939
R21230 vdd.n3430 vdd.n601 0.152939
R21231 vdd.n3193 vdd.n656 0.152939
R21232 vdd.n2121 vdd.n1118 0.152939
R21233 vdd.n1459 vdd.n1458 0.152939
R21234 vdd.n1459 vdd.n1215 0.152939
R21235 vdd.n1473 vdd.n1215 0.152939
R21236 vdd.n1474 vdd.n1473 0.152939
R21237 vdd.n1475 vdd.n1474 0.152939
R21238 vdd.n1475 vdd.n1203 0.152939
R21239 vdd.n1490 vdd.n1203 0.152939
R21240 vdd.n1491 vdd.n1490 0.152939
R21241 vdd.n1492 vdd.n1491 0.152939
R21242 vdd.n1492 vdd.n1193 0.152939
R21243 vdd.n1507 vdd.n1193 0.152939
R21244 vdd.n1508 vdd.n1507 0.152939
R21245 vdd.n1509 vdd.n1508 0.152939
R21246 vdd.n1509 vdd.n1180 0.152939
R21247 vdd.n1523 vdd.n1180 0.152939
R21248 vdd.n1524 vdd.n1523 0.152939
R21249 vdd.n1525 vdd.n1524 0.152939
R21250 vdd.n1525 vdd.n1169 0.152939
R21251 vdd.n1835 vdd.n1169 0.152939
R21252 vdd.n1836 vdd.n1835 0.152939
R21253 vdd.n1837 vdd.n1836 0.152939
R21254 vdd.n1837 vdd.n1158 0.152939
R21255 vdd.n1851 vdd.n1158 0.152939
R21256 vdd.n1852 vdd.n1851 0.152939
R21257 vdd.n1853 vdd.n1852 0.152939
R21258 vdd.n1853 vdd.n1146 0.152939
R21259 vdd.n1868 vdd.n1146 0.152939
R21260 vdd.n1869 vdd.n1868 0.152939
R21261 vdd.n1870 vdd.n1869 0.152939
R21262 vdd.n1870 vdd.n1136 0.152939
R21263 vdd.n1885 vdd.n1136 0.152939
R21264 vdd.n1886 vdd.n1885 0.152939
R21265 vdd.n1889 vdd.n1886 0.152939
R21266 vdd.n1889 vdd.n1888 0.152939
R21267 vdd.n1888 vdd.n1887 0.152939
R21268 vdd.n1449 vdd.n1264 0.152939
R21269 vdd.n1449 vdd.n1448 0.152939
R21270 vdd.n1448 vdd.n1447 0.152939
R21271 vdd.n1447 vdd.n1266 0.152939
R21272 vdd.n1443 vdd.n1266 0.152939
R21273 vdd.n1443 vdd.n1442 0.152939
R21274 vdd.n1442 vdd.n1441 0.152939
R21275 vdd.n1441 vdd.n1271 0.152939
R21276 vdd.n1437 vdd.n1271 0.152939
R21277 vdd.n1437 vdd.n1436 0.152939
R21278 vdd.n1436 vdd.n1435 0.152939
R21279 vdd.n1435 vdd.n1277 0.152939
R21280 vdd.n1431 vdd.n1277 0.152939
R21281 vdd.n1431 vdd.n1430 0.152939
R21282 vdd.n1430 vdd.n1429 0.152939
R21283 vdd.n1429 vdd.n1283 0.152939
R21284 vdd.n1425 vdd.n1283 0.152939
R21285 vdd.n1425 vdd.n1424 0.152939
R21286 vdd.n1424 vdd.n1423 0.152939
R21287 vdd.n1423 vdd.n1289 0.152939
R21288 vdd.n1415 vdd.n1289 0.152939
R21289 vdd.n1415 vdd.n1414 0.152939
R21290 vdd.n1414 vdd.n1413 0.152939
R21291 vdd.n1413 vdd.n1293 0.152939
R21292 vdd.n1409 vdd.n1293 0.152939
R21293 vdd.n1409 vdd.n1408 0.152939
R21294 vdd.n1408 vdd.n1407 0.152939
R21295 vdd.n1407 vdd.n1299 0.152939
R21296 vdd.n1403 vdd.n1299 0.152939
R21297 vdd.n1403 vdd.n1402 0.152939
R21298 vdd.n1402 vdd.n1401 0.152939
R21299 vdd.n1401 vdd.n1305 0.152939
R21300 vdd.n1397 vdd.n1305 0.152939
R21301 vdd.n1397 vdd.n1396 0.152939
R21302 vdd.n1396 vdd.n1395 0.152939
R21303 vdd.n1395 vdd.n1311 0.152939
R21304 vdd.n1391 vdd.n1311 0.152939
R21305 vdd.n1391 vdd.n1390 0.152939
R21306 vdd.n1390 vdd.n1389 0.152939
R21307 vdd.n1389 vdd.n1317 0.152939
R21308 vdd.n1382 vdd.n1317 0.152939
R21309 vdd.n1382 vdd.n1381 0.152939
R21310 vdd.n1381 vdd.n1380 0.152939
R21311 vdd.n1380 vdd.n1322 0.152939
R21312 vdd.n1376 vdd.n1322 0.152939
R21313 vdd.n1376 vdd.n1375 0.152939
R21314 vdd.n1375 vdd.n1374 0.152939
R21315 vdd.n1374 vdd.n1328 0.152939
R21316 vdd.n1370 vdd.n1328 0.152939
R21317 vdd.n1370 vdd.n1369 0.152939
R21318 vdd.n1369 vdd.n1368 0.152939
R21319 vdd.n1368 vdd.n1334 0.152939
R21320 vdd.n1364 vdd.n1334 0.152939
R21321 vdd.n1364 vdd.n1363 0.152939
R21322 vdd.n1363 vdd.n1362 0.152939
R21323 vdd.n1362 vdd.n1340 0.152939
R21324 vdd.n1358 vdd.n1340 0.152939
R21325 vdd.n1358 vdd.n1357 0.152939
R21326 vdd.n1357 vdd.n1356 0.152939
R21327 vdd.n1356 vdd.n1346 0.152939
R21328 vdd.n1352 vdd.n1346 0.152939
R21329 vdd.n1352 vdd.n1227 0.152939
R21330 vdd.n1457 vdd.n1227 0.152939
R21331 vdd.n1465 vdd.n1221 0.152939
R21332 vdd.n1466 vdd.n1465 0.152939
R21333 vdd.n1467 vdd.n1466 0.152939
R21334 vdd.n1467 vdd.n1209 0.152939
R21335 vdd.n1482 vdd.n1209 0.152939
R21336 vdd.n1483 vdd.n1482 0.152939
R21337 vdd.n1484 vdd.n1483 0.152939
R21338 vdd.n1484 vdd.n1198 0.152939
R21339 vdd.n1499 vdd.n1198 0.152939
R21340 vdd.n1500 vdd.n1499 0.152939
R21341 vdd.n1501 vdd.n1500 0.152939
R21342 vdd.n1501 vdd.n1187 0.152939
R21343 vdd.n1515 vdd.n1187 0.152939
R21344 vdd.n1516 vdd.n1515 0.152939
R21345 vdd.n1517 vdd.n1516 0.152939
R21346 vdd.n1517 vdd.n1175 0.152939
R21347 vdd.n1532 vdd.n1175 0.152939
R21348 vdd.n2408 vdd.t253 0.113865
R21349 vdd.n2475 vdd.t269 0.113865
R21350 vdd.n2958 vdd.t223 0.113865
R21351 vdd.n3025 vdd.t252 0.113865
R21352 vdd.n2099 vdd.n1897 0.110256
R21353 vdd.n3124 vdd.n661 0.110256
R21354 vdd.n3193 vdd.n3192 0.110256
R21355 vdd.n2122 vdd.n2121 0.110256
R21356 vdd.n1828 vdd.n1827 0.0695946
R21357 vdd.n3473 vdd.n322 0.0695946
R21358 vdd.n3473 vdd.n3472 0.0695946
R21359 vdd.n1827 vdd.n1532 0.0695946
R21360 vdd.n2099 vdd.n2098 0.0431829
R21361 vdd.n2122 vdd.n1115 0.0431829
R21362 vdd.n3124 vdd.n667 0.0431829
R21363 vdd.n3192 vdd.n748 0.0431829
R21364 vdd vdd.n28 0.00833333
R21365 CSoutput.n19 CSoutput.t180 184.661
R21366 CSoutput.n78 CSoutput.n77 165.8
R21367 CSoutput.n76 CSoutput.n0 165.8
R21368 CSoutput.n75 CSoutput.n74 165.8
R21369 CSoutput.n73 CSoutput.n72 165.8
R21370 CSoutput.n71 CSoutput.n2 165.8
R21371 CSoutput.n69 CSoutput.n68 165.8
R21372 CSoutput.n67 CSoutput.n3 165.8
R21373 CSoutput.n66 CSoutput.n65 165.8
R21374 CSoutput.n63 CSoutput.n4 165.8
R21375 CSoutput.n61 CSoutput.n60 165.8
R21376 CSoutput.n59 CSoutput.n5 165.8
R21377 CSoutput.n58 CSoutput.n57 165.8
R21378 CSoutput.n55 CSoutput.n6 165.8
R21379 CSoutput.n54 CSoutput.n53 165.8
R21380 CSoutput.n52 CSoutput.n51 165.8
R21381 CSoutput.n50 CSoutput.n8 165.8
R21382 CSoutput.n48 CSoutput.n47 165.8
R21383 CSoutput.n46 CSoutput.n9 165.8
R21384 CSoutput.n45 CSoutput.n44 165.8
R21385 CSoutput.n42 CSoutput.n10 165.8
R21386 CSoutput.n41 CSoutput.n40 165.8
R21387 CSoutput.n39 CSoutput.n38 165.8
R21388 CSoutput.n37 CSoutput.n12 165.8
R21389 CSoutput.n35 CSoutput.n34 165.8
R21390 CSoutput.n33 CSoutput.n13 165.8
R21391 CSoutput.n32 CSoutput.n31 165.8
R21392 CSoutput.n29 CSoutput.n14 165.8
R21393 CSoutput.n28 CSoutput.n27 165.8
R21394 CSoutput.n26 CSoutput.n25 165.8
R21395 CSoutput.n24 CSoutput.n16 165.8
R21396 CSoutput.n22 CSoutput.n21 165.8
R21397 CSoutput.n20 CSoutput.n17 165.8
R21398 CSoutput.n77 CSoutput.t183 162.194
R21399 CSoutput.n18 CSoutput.t177 120.501
R21400 CSoutput.n23 CSoutput.t194 120.501
R21401 CSoutput.n15 CSoutput.t189 120.501
R21402 CSoutput.n30 CSoutput.t178 120.501
R21403 CSoutput.n36 CSoutput.t179 120.501
R21404 CSoutput.n11 CSoutput.t191 120.501
R21405 CSoutput.n43 CSoutput.t188 120.501
R21406 CSoutput.n49 CSoutput.t182 120.501
R21407 CSoutput.n7 CSoutput.t195 120.501
R21408 CSoutput.n56 CSoutput.t196 120.501
R21409 CSoutput.n62 CSoutput.t185 120.501
R21410 CSoutput.n64 CSoutput.t197 120.501
R21411 CSoutput.n70 CSoutput.t176 120.501
R21412 CSoutput.n1 CSoutput.t193 120.501
R21413 CSoutput.n310 CSoutput.n308 103.469
R21414 CSoutput.n294 CSoutput.n292 103.469
R21415 CSoutput.n279 CSoutput.n277 103.469
R21416 CSoutput.n112 CSoutput.n110 103.469
R21417 CSoutput.n96 CSoutput.n94 103.469
R21418 CSoutput.n81 CSoutput.n79 103.469
R21419 CSoutput.n320 CSoutput.n319 103.111
R21420 CSoutput.n318 CSoutput.n317 103.111
R21421 CSoutput.n316 CSoutput.n315 103.111
R21422 CSoutput.n314 CSoutput.n313 103.111
R21423 CSoutput.n312 CSoutput.n311 103.111
R21424 CSoutput.n310 CSoutput.n309 103.111
R21425 CSoutput.n306 CSoutput.n305 103.111
R21426 CSoutput.n304 CSoutput.n303 103.111
R21427 CSoutput.n302 CSoutput.n301 103.111
R21428 CSoutput.n300 CSoutput.n299 103.111
R21429 CSoutput.n298 CSoutput.n297 103.111
R21430 CSoutput.n296 CSoutput.n295 103.111
R21431 CSoutput.n294 CSoutput.n293 103.111
R21432 CSoutput.n291 CSoutput.n290 103.111
R21433 CSoutput.n289 CSoutput.n288 103.111
R21434 CSoutput.n287 CSoutput.n286 103.111
R21435 CSoutput.n285 CSoutput.n284 103.111
R21436 CSoutput.n283 CSoutput.n282 103.111
R21437 CSoutput.n281 CSoutput.n280 103.111
R21438 CSoutput.n279 CSoutput.n278 103.111
R21439 CSoutput.n112 CSoutput.n111 103.111
R21440 CSoutput.n114 CSoutput.n113 103.111
R21441 CSoutput.n116 CSoutput.n115 103.111
R21442 CSoutput.n118 CSoutput.n117 103.111
R21443 CSoutput.n120 CSoutput.n119 103.111
R21444 CSoutput.n122 CSoutput.n121 103.111
R21445 CSoutput.n124 CSoutput.n123 103.111
R21446 CSoutput.n96 CSoutput.n95 103.111
R21447 CSoutput.n98 CSoutput.n97 103.111
R21448 CSoutput.n100 CSoutput.n99 103.111
R21449 CSoutput.n102 CSoutput.n101 103.111
R21450 CSoutput.n104 CSoutput.n103 103.111
R21451 CSoutput.n106 CSoutput.n105 103.111
R21452 CSoutput.n108 CSoutput.n107 103.111
R21453 CSoutput.n81 CSoutput.n80 103.111
R21454 CSoutput.n83 CSoutput.n82 103.111
R21455 CSoutput.n85 CSoutput.n84 103.111
R21456 CSoutput.n87 CSoutput.n86 103.111
R21457 CSoutput.n89 CSoutput.n88 103.111
R21458 CSoutput.n91 CSoutput.n90 103.111
R21459 CSoutput.n93 CSoutput.n92 103.111
R21460 CSoutput.n322 CSoutput.n321 103.111
R21461 CSoutput.n346 CSoutput.n344 81.5057
R21462 CSoutput.n327 CSoutput.n325 81.5057
R21463 CSoutput.n386 CSoutput.n384 81.5057
R21464 CSoutput.n367 CSoutput.n365 81.5057
R21465 CSoutput.n362 CSoutput.n361 80.9324
R21466 CSoutput.n360 CSoutput.n359 80.9324
R21467 CSoutput.n358 CSoutput.n357 80.9324
R21468 CSoutput.n356 CSoutput.n355 80.9324
R21469 CSoutput.n354 CSoutput.n353 80.9324
R21470 CSoutput.n352 CSoutput.n351 80.9324
R21471 CSoutput.n350 CSoutput.n349 80.9324
R21472 CSoutput.n348 CSoutput.n347 80.9324
R21473 CSoutput.n346 CSoutput.n345 80.9324
R21474 CSoutput.n343 CSoutput.n342 80.9324
R21475 CSoutput.n341 CSoutput.n340 80.9324
R21476 CSoutput.n339 CSoutput.n338 80.9324
R21477 CSoutput.n337 CSoutput.n336 80.9324
R21478 CSoutput.n335 CSoutput.n334 80.9324
R21479 CSoutput.n333 CSoutput.n332 80.9324
R21480 CSoutput.n331 CSoutput.n330 80.9324
R21481 CSoutput.n329 CSoutput.n328 80.9324
R21482 CSoutput.n327 CSoutput.n326 80.9324
R21483 CSoutput.n386 CSoutput.n385 80.9324
R21484 CSoutput.n388 CSoutput.n387 80.9324
R21485 CSoutput.n390 CSoutput.n389 80.9324
R21486 CSoutput.n392 CSoutput.n391 80.9324
R21487 CSoutput.n394 CSoutput.n393 80.9324
R21488 CSoutput.n396 CSoutput.n395 80.9324
R21489 CSoutput.n398 CSoutput.n397 80.9324
R21490 CSoutput.n400 CSoutput.n399 80.9324
R21491 CSoutput.n402 CSoutput.n401 80.9324
R21492 CSoutput.n367 CSoutput.n366 80.9324
R21493 CSoutput.n369 CSoutput.n368 80.9324
R21494 CSoutput.n371 CSoutput.n370 80.9324
R21495 CSoutput.n373 CSoutput.n372 80.9324
R21496 CSoutput.n375 CSoutput.n374 80.9324
R21497 CSoutput.n377 CSoutput.n376 80.9324
R21498 CSoutput.n379 CSoutput.n378 80.9324
R21499 CSoutput.n381 CSoutput.n380 80.9324
R21500 CSoutput.n383 CSoutput.n382 80.9324
R21501 CSoutput.n25 CSoutput.n24 48.1486
R21502 CSoutput.n69 CSoutput.n3 48.1486
R21503 CSoutput.n38 CSoutput.n37 48.1486
R21504 CSoutput.n42 CSoutput.n41 48.1486
R21505 CSoutput.n51 CSoutput.n50 48.1486
R21506 CSoutput.n55 CSoutput.n54 48.1486
R21507 CSoutput.n22 CSoutput.n17 46.462
R21508 CSoutput.n72 CSoutput.n71 46.462
R21509 CSoutput.n20 CSoutput.n19 44.9055
R21510 CSoutput.n29 CSoutput.n28 43.7635
R21511 CSoutput.n65 CSoutput.n63 43.7635
R21512 CSoutput.n35 CSoutput.n13 41.7396
R21513 CSoutput.n57 CSoutput.n5 41.7396
R21514 CSoutput.n44 CSoutput.n9 37.0171
R21515 CSoutput.n48 CSoutput.n9 37.0171
R21516 CSoutput.n76 CSoutput.n75 34.9932
R21517 CSoutput.n31 CSoutput.n13 32.2947
R21518 CSoutput.n61 CSoutput.n5 32.2947
R21519 CSoutput.n30 CSoutput.n29 29.6014
R21520 CSoutput.n63 CSoutput.n62 29.6014
R21521 CSoutput.n19 CSoutput.n18 28.4085
R21522 CSoutput.n18 CSoutput.n17 25.1176
R21523 CSoutput.n72 CSoutput.n1 25.1176
R21524 CSoutput.n43 CSoutput.n42 22.0922
R21525 CSoutput.n50 CSoutput.n49 22.0922
R21526 CSoutput.n77 CSoutput.n76 21.8586
R21527 CSoutput.n37 CSoutput.n36 18.9681
R21528 CSoutput.n56 CSoutput.n55 18.9681
R21529 CSoutput.n25 CSoutput.n15 17.6292
R21530 CSoutput.n64 CSoutput.n3 17.6292
R21531 CSoutput.n24 CSoutput.n23 15.844
R21532 CSoutput.n70 CSoutput.n69 15.844
R21533 CSoutput.n38 CSoutput.n11 14.5051
R21534 CSoutput.n54 CSoutput.n7 14.5051
R21535 CSoutput.n405 CSoutput.n78 11.6139
R21536 CSoutput.n41 CSoutput.n11 11.3811
R21537 CSoutput.n51 CSoutput.n7 11.3811
R21538 CSoutput.n23 CSoutput.n22 10.0422
R21539 CSoutput.n71 CSoutput.n70 10.0422
R21540 CSoutput.n307 CSoutput.n291 9.25285
R21541 CSoutput.n109 CSoutput.n93 9.25285
R21542 CSoutput.n364 CSoutput.n324 8.99065
R21543 CSoutput.n363 CSoutput.n343 8.97993
R21544 CSoutput.n403 CSoutput.n383 8.97993
R21545 CSoutput.n28 CSoutput.n15 8.25698
R21546 CSoutput.n65 CSoutput.n64 8.25698
R21547 CSoutput.n364 CSoutput.n363 7.89345
R21548 CSoutput.n404 CSoutput.n403 7.89345
R21549 CSoutput.n324 CSoutput.n323 7.12641
R21550 CSoutput.n126 CSoutput.n125 7.12641
R21551 CSoutput.n36 CSoutput.n35 6.91809
R21552 CSoutput.n57 CSoutput.n56 6.91809
R21553 CSoutput.n405 CSoutput.n126 5.39821
R21554 CSoutput.n363 CSoutput.n362 5.25266
R21555 CSoutput.n403 CSoutput.n402 5.25266
R21556 CSoutput.n323 CSoutput.n322 5.1449
R21557 CSoutput.n307 CSoutput.n306 5.1449
R21558 CSoutput.n125 CSoutput.n124 5.1449
R21559 CSoutput.n109 CSoutput.n108 5.1449
R21560 CSoutput.n217 CSoutput.n170 4.5005
R21561 CSoutput.n186 CSoutput.n170 4.5005
R21562 CSoutput.n181 CSoutput.n165 4.5005
R21563 CSoutput.n181 CSoutput.n167 4.5005
R21564 CSoutput.n181 CSoutput.n164 4.5005
R21565 CSoutput.n181 CSoutput.n168 4.5005
R21566 CSoutput.n181 CSoutput.n163 4.5005
R21567 CSoutput.n181 CSoutput.t184 4.5005
R21568 CSoutput.n181 CSoutput.n162 4.5005
R21569 CSoutput.n181 CSoutput.n169 4.5005
R21570 CSoutput.n181 CSoutput.n170 4.5005
R21571 CSoutput.n179 CSoutput.n165 4.5005
R21572 CSoutput.n179 CSoutput.n167 4.5005
R21573 CSoutput.n179 CSoutput.n164 4.5005
R21574 CSoutput.n179 CSoutput.n168 4.5005
R21575 CSoutput.n179 CSoutput.n163 4.5005
R21576 CSoutput.n179 CSoutput.t184 4.5005
R21577 CSoutput.n179 CSoutput.n162 4.5005
R21578 CSoutput.n179 CSoutput.n169 4.5005
R21579 CSoutput.n179 CSoutput.n170 4.5005
R21580 CSoutput.n178 CSoutput.n165 4.5005
R21581 CSoutput.n178 CSoutput.n167 4.5005
R21582 CSoutput.n178 CSoutput.n164 4.5005
R21583 CSoutput.n178 CSoutput.n168 4.5005
R21584 CSoutput.n178 CSoutput.n163 4.5005
R21585 CSoutput.n178 CSoutput.t184 4.5005
R21586 CSoutput.n178 CSoutput.n162 4.5005
R21587 CSoutput.n178 CSoutput.n169 4.5005
R21588 CSoutput.n178 CSoutput.n170 4.5005
R21589 CSoutput.n263 CSoutput.n165 4.5005
R21590 CSoutput.n263 CSoutput.n167 4.5005
R21591 CSoutput.n263 CSoutput.n164 4.5005
R21592 CSoutput.n263 CSoutput.n168 4.5005
R21593 CSoutput.n263 CSoutput.n163 4.5005
R21594 CSoutput.n263 CSoutput.t184 4.5005
R21595 CSoutput.n263 CSoutput.n162 4.5005
R21596 CSoutput.n263 CSoutput.n169 4.5005
R21597 CSoutput.n263 CSoutput.n170 4.5005
R21598 CSoutput.n261 CSoutput.n165 4.5005
R21599 CSoutput.n261 CSoutput.n167 4.5005
R21600 CSoutput.n261 CSoutput.n164 4.5005
R21601 CSoutput.n261 CSoutput.n168 4.5005
R21602 CSoutput.n261 CSoutput.n163 4.5005
R21603 CSoutput.n261 CSoutput.t184 4.5005
R21604 CSoutput.n261 CSoutput.n162 4.5005
R21605 CSoutput.n261 CSoutput.n169 4.5005
R21606 CSoutput.n259 CSoutput.n165 4.5005
R21607 CSoutput.n259 CSoutput.n167 4.5005
R21608 CSoutput.n259 CSoutput.n164 4.5005
R21609 CSoutput.n259 CSoutput.n168 4.5005
R21610 CSoutput.n259 CSoutput.n163 4.5005
R21611 CSoutput.n259 CSoutput.t184 4.5005
R21612 CSoutput.n259 CSoutput.n162 4.5005
R21613 CSoutput.n259 CSoutput.n169 4.5005
R21614 CSoutput.n189 CSoutput.n165 4.5005
R21615 CSoutput.n189 CSoutput.n167 4.5005
R21616 CSoutput.n189 CSoutput.n164 4.5005
R21617 CSoutput.n189 CSoutput.n168 4.5005
R21618 CSoutput.n189 CSoutput.n163 4.5005
R21619 CSoutput.n189 CSoutput.t184 4.5005
R21620 CSoutput.n189 CSoutput.n162 4.5005
R21621 CSoutput.n189 CSoutput.n169 4.5005
R21622 CSoutput.n189 CSoutput.n170 4.5005
R21623 CSoutput.n188 CSoutput.n165 4.5005
R21624 CSoutput.n188 CSoutput.n167 4.5005
R21625 CSoutput.n188 CSoutput.n164 4.5005
R21626 CSoutput.n188 CSoutput.n168 4.5005
R21627 CSoutput.n188 CSoutput.n163 4.5005
R21628 CSoutput.n188 CSoutput.t184 4.5005
R21629 CSoutput.n188 CSoutput.n162 4.5005
R21630 CSoutput.n188 CSoutput.n169 4.5005
R21631 CSoutput.n188 CSoutput.n170 4.5005
R21632 CSoutput.n192 CSoutput.n165 4.5005
R21633 CSoutput.n192 CSoutput.n167 4.5005
R21634 CSoutput.n192 CSoutput.n164 4.5005
R21635 CSoutput.n192 CSoutput.n168 4.5005
R21636 CSoutput.n192 CSoutput.n163 4.5005
R21637 CSoutput.n192 CSoutput.t184 4.5005
R21638 CSoutput.n192 CSoutput.n162 4.5005
R21639 CSoutput.n192 CSoutput.n169 4.5005
R21640 CSoutput.n192 CSoutput.n170 4.5005
R21641 CSoutput.n191 CSoutput.n165 4.5005
R21642 CSoutput.n191 CSoutput.n167 4.5005
R21643 CSoutput.n191 CSoutput.n164 4.5005
R21644 CSoutput.n191 CSoutput.n168 4.5005
R21645 CSoutput.n191 CSoutput.n163 4.5005
R21646 CSoutput.n191 CSoutput.t184 4.5005
R21647 CSoutput.n191 CSoutput.n162 4.5005
R21648 CSoutput.n191 CSoutput.n169 4.5005
R21649 CSoutput.n191 CSoutput.n170 4.5005
R21650 CSoutput.n174 CSoutput.n165 4.5005
R21651 CSoutput.n174 CSoutput.n167 4.5005
R21652 CSoutput.n174 CSoutput.n164 4.5005
R21653 CSoutput.n174 CSoutput.n168 4.5005
R21654 CSoutput.n174 CSoutput.n163 4.5005
R21655 CSoutput.n174 CSoutput.t184 4.5005
R21656 CSoutput.n174 CSoutput.n162 4.5005
R21657 CSoutput.n174 CSoutput.n169 4.5005
R21658 CSoutput.n174 CSoutput.n170 4.5005
R21659 CSoutput.n266 CSoutput.n165 4.5005
R21660 CSoutput.n266 CSoutput.n167 4.5005
R21661 CSoutput.n266 CSoutput.n164 4.5005
R21662 CSoutput.n266 CSoutput.n168 4.5005
R21663 CSoutput.n266 CSoutput.n163 4.5005
R21664 CSoutput.n266 CSoutput.t184 4.5005
R21665 CSoutput.n266 CSoutput.n162 4.5005
R21666 CSoutput.n266 CSoutput.n169 4.5005
R21667 CSoutput.n266 CSoutput.n170 4.5005
R21668 CSoutput.n253 CSoutput.n224 4.5005
R21669 CSoutput.n253 CSoutput.n230 4.5005
R21670 CSoutput.n211 CSoutput.n200 4.5005
R21671 CSoutput.n211 CSoutput.n202 4.5005
R21672 CSoutput.n211 CSoutput.n199 4.5005
R21673 CSoutput.n211 CSoutput.n203 4.5005
R21674 CSoutput.n211 CSoutput.n198 4.5005
R21675 CSoutput.n211 CSoutput.t186 4.5005
R21676 CSoutput.n211 CSoutput.n197 4.5005
R21677 CSoutput.n211 CSoutput.n204 4.5005
R21678 CSoutput.n253 CSoutput.n211 4.5005
R21679 CSoutput.n232 CSoutput.n200 4.5005
R21680 CSoutput.n232 CSoutput.n202 4.5005
R21681 CSoutput.n232 CSoutput.n199 4.5005
R21682 CSoutput.n232 CSoutput.n203 4.5005
R21683 CSoutput.n232 CSoutput.n198 4.5005
R21684 CSoutput.n232 CSoutput.t186 4.5005
R21685 CSoutput.n232 CSoutput.n197 4.5005
R21686 CSoutput.n232 CSoutput.n204 4.5005
R21687 CSoutput.n253 CSoutput.n232 4.5005
R21688 CSoutput.n210 CSoutput.n200 4.5005
R21689 CSoutput.n210 CSoutput.n202 4.5005
R21690 CSoutput.n210 CSoutput.n199 4.5005
R21691 CSoutput.n210 CSoutput.n203 4.5005
R21692 CSoutput.n210 CSoutput.n198 4.5005
R21693 CSoutput.n210 CSoutput.t186 4.5005
R21694 CSoutput.n210 CSoutput.n197 4.5005
R21695 CSoutput.n210 CSoutput.n204 4.5005
R21696 CSoutput.n253 CSoutput.n210 4.5005
R21697 CSoutput.n234 CSoutput.n200 4.5005
R21698 CSoutput.n234 CSoutput.n202 4.5005
R21699 CSoutput.n234 CSoutput.n199 4.5005
R21700 CSoutput.n234 CSoutput.n203 4.5005
R21701 CSoutput.n234 CSoutput.n198 4.5005
R21702 CSoutput.n234 CSoutput.t186 4.5005
R21703 CSoutput.n234 CSoutput.n197 4.5005
R21704 CSoutput.n234 CSoutput.n204 4.5005
R21705 CSoutput.n253 CSoutput.n234 4.5005
R21706 CSoutput.n200 CSoutput.n195 4.5005
R21707 CSoutput.n202 CSoutput.n195 4.5005
R21708 CSoutput.n199 CSoutput.n195 4.5005
R21709 CSoutput.n203 CSoutput.n195 4.5005
R21710 CSoutput.n198 CSoutput.n195 4.5005
R21711 CSoutput.t186 CSoutput.n195 4.5005
R21712 CSoutput.n197 CSoutput.n195 4.5005
R21713 CSoutput.n204 CSoutput.n195 4.5005
R21714 CSoutput.n256 CSoutput.n200 4.5005
R21715 CSoutput.n256 CSoutput.n202 4.5005
R21716 CSoutput.n256 CSoutput.n199 4.5005
R21717 CSoutput.n256 CSoutput.n203 4.5005
R21718 CSoutput.n256 CSoutput.n198 4.5005
R21719 CSoutput.n256 CSoutput.t186 4.5005
R21720 CSoutput.n256 CSoutput.n197 4.5005
R21721 CSoutput.n256 CSoutput.n204 4.5005
R21722 CSoutput.n254 CSoutput.n200 4.5005
R21723 CSoutput.n254 CSoutput.n202 4.5005
R21724 CSoutput.n254 CSoutput.n199 4.5005
R21725 CSoutput.n254 CSoutput.n203 4.5005
R21726 CSoutput.n254 CSoutput.n198 4.5005
R21727 CSoutput.n254 CSoutput.t186 4.5005
R21728 CSoutput.n254 CSoutput.n197 4.5005
R21729 CSoutput.n254 CSoutput.n204 4.5005
R21730 CSoutput.n254 CSoutput.n253 4.5005
R21731 CSoutput.n236 CSoutput.n200 4.5005
R21732 CSoutput.n236 CSoutput.n202 4.5005
R21733 CSoutput.n236 CSoutput.n199 4.5005
R21734 CSoutput.n236 CSoutput.n203 4.5005
R21735 CSoutput.n236 CSoutput.n198 4.5005
R21736 CSoutput.n236 CSoutput.t186 4.5005
R21737 CSoutput.n236 CSoutput.n197 4.5005
R21738 CSoutput.n236 CSoutput.n204 4.5005
R21739 CSoutput.n253 CSoutput.n236 4.5005
R21740 CSoutput.n208 CSoutput.n200 4.5005
R21741 CSoutput.n208 CSoutput.n202 4.5005
R21742 CSoutput.n208 CSoutput.n199 4.5005
R21743 CSoutput.n208 CSoutput.n203 4.5005
R21744 CSoutput.n208 CSoutput.n198 4.5005
R21745 CSoutput.n208 CSoutput.t186 4.5005
R21746 CSoutput.n208 CSoutput.n197 4.5005
R21747 CSoutput.n208 CSoutput.n204 4.5005
R21748 CSoutput.n253 CSoutput.n208 4.5005
R21749 CSoutput.n238 CSoutput.n200 4.5005
R21750 CSoutput.n238 CSoutput.n202 4.5005
R21751 CSoutput.n238 CSoutput.n199 4.5005
R21752 CSoutput.n238 CSoutput.n203 4.5005
R21753 CSoutput.n238 CSoutput.n198 4.5005
R21754 CSoutput.n238 CSoutput.t186 4.5005
R21755 CSoutput.n238 CSoutput.n197 4.5005
R21756 CSoutput.n238 CSoutput.n204 4.5005
R21757 CSoutput.n253 CSoutput.n238 4.5005
R21758 CSoutput.n207 CSoutput.n200 4.5005
R21759 CSoutput.n207 CSoutput.n202 4.5005
R21760 CSoutput.n207 CSoutput.n199 4.5005
R21761 CSoutput.n207 CSoutput.n203 4.5005
R21762 CSoutput.n207 CSoutput.n198 4.5005
R21763 CSoutput.n207 CSoutput.t186 4.5005
R21764 CSoutput.n207 CSoutput.n197 4.5005
R21765 CSoutput.n207 CSoutput.n204 4.5005
R21766 CSoutput.n253 CSoutput.n207 4.5005
R21767 CSoutput.n252 CSoutput.n200 4.5005
R21768 CSoutput.n252 CSoutput.n202 4.5005
R21769 CSoutput.n252 CSoutput.n199 4.5005
R21770 CSoutput.n252 CSoutput.n203 4.5005
R21771 CSoutput.n252 CSoutput.n198 4.5005
R21772 CSoutput.n252 CSoutput.t186 4.5005
R21773 CSoutput.n252 CSoutput.n197 4.5005
R21774 CSoutput.n252 CSoutput.n204 4.5005
R21775 CSoutput.n253 CSoutput.n252 4.5005
R21776 CSoutput.n251 CSoutput.n136 4.5005
R21777 CSoutput.n152 CSoutput.n136 4.5005
R21778 CSoutput.n147 CSoutput.n131 4.5005
R21779 CSoutput.n147 CSoutput.n133 4.5005
R21780 CSoutput.n147 CSoutput.n130 4.5005
R21781 CSoutput.n147 CSoutput.n134 4.5005
R21782 CSoutput.n147 CSoutput.n129 4.5005
R21783 CSoutput.n147 CSoutput.t187 4.5005
R21784 CSoutput.n147 CSoutput.n128 4.5005
R21785 CSoutput.n147 CSoutput.n135 4.5005
R21786 CSoutput.n147 CSoutput.n136 4.5005
R21787 CSoutput.n145 CSoutput.n131 4.5005
R21788 CSoutput.n145 CSoutput.n133 4.5005
R21789 CSoutput.n145 CSoutput.n130 4.5005
R21790 CSoutput.n145 CSoutput.n134 4.5005
R21791 CSoutput.n145 CSoutput.n129 4.5005
R21792 CSoutput.n145 CSoutput.t187 4.5005
R21793 CSoutput.n145 CSoutput.n128 4.5005
R21794 CSoutput.n145 CSoutput.n135 4.5005
R21795 CSoutput.n145 CSoutput.n136 4.5005
R21796 CSoutput.n144 CSoutput.n131 4.5005
R21797 CSoutput.n144 CSoutput.n133 4.5005
R21798 CSoutput.n144 CSoutput.n130 4.5005
R21799 CSoutput.n144 CSoutput.n134 4.5005
R21800 CSoutput.n144 CSoutput.n129 4.5005
R21801 CSoutput.n144 CSoutput.t187 4.5005
R21802 CSoutput.n144 CSoutput.n128 4.5005
R21803 CSoutput.n144 CSoutput.n135 4.5005
R21804 CSoutput.n144 CSoutput.n136 4.5005
R21805 CSoutput.n273 CSoutput.n131 4.5005
R21806 CSoutput.n273 CSoutput.n133 4.5005
R21807 CSoutput.n273 CSoutput.n130 4.5005
R21808 CSoutput.n273 CSoutput.n134 4.5005
R21809 CSoutput.n273 CSoutput.n129 4.5005
R21810 CSoutput.n273 CSoutput.t187 4.5005
R21811 CSoutput.n273 CSoutput.n128 4.5005
R21812 CSoutput.n273 CSoutput.n135 4.5005
R21813 CSoutput.n273 CSoutput.n136 4.5005
R21814 CSoutput.n271 CSoutput.n131 4.5005
R21815 CSoutput.n271 CSoutput.n133 4.5005
R21816 CSoutput.n271 CSoutput.n130 4.5005
R21817 CSoutput.n271 CSoutput.n134 4.5005
R21818 CSoutput.n271 CSoutput.n129 4.5005
R21819 CSoutput.n271 CSoutput.t187 4.5005
R21820 CSoutput.n271 CSoutput.n128 4.5005
R21821 CSoutput.n271 CSoutput.n135 4.5005
R21822 CSoutput.n269 CSoutput.n131 4.5005
R21823 CSoutput.n269 CSoutput.n133 4.5005
R21824 CSoutput.n269 CSoutput.n130 4.5005
R21825 CSoutput.n269 CSoutput.n134 4.5005
R21826 CSoutput.n269 CSoutput.n129 4.5005
R21827 CSoutput.n269 CSoutput.t187 4.5005
R21828 CSoutput.n269 CSoutput.n128 4.5005
R21829 CSoutput.n269 CSoutput.n135 4.5005
R21830 CSoutput.n155 CSoutput.n131 4.5005
R21831 CSoutput.n155 CSoutput.n133 4.5005
R21832 CSoutput.n155 CSoutput.n130 4.5005
R21833 CSoutput.n155 CSoutput.n134 4.5005
R21834 CSoutput.n155 CSoutput.n129 4.5005
R21835 CSoutput.n155 CSoutput.t187 4.5005
R21836 CSoutput.n155 CSoutput.n128 4.5005
R21837 CSoutput.n155 CSoutput.n135 4.5005
R21838 CSoutput.n155 CSoutput.n136 4.5005
R21839 CSoutput.n154 CSoutput.n131 4.5005
R21840 CSoutput.n154 CSoutput.n133 4.5005
R21841 CSoutput.n154 CSoutput.n130 4.5005
R21842 CSoutput.n154 CSoutput.n134 4.5005
R21843 CSoutput.n154 CSoutput.n129 4.5005
R21844 CSoutput.n154 CSoutput.t187 4.5005
R21845 CSoutput.n154 CSoutput.n128 4.5005
R21846 CSoutput.n154 CSoutput.n135 4.5005
R21847 CSoutput.n154 CSoutput.n136 4.5005
R21848 CSoutput.n158 CSoutput.n131 4.5005
R21849 CSoutput.n158 CSoutput.n133 4.5005
R21850 CSoutput.n158 CSoutput.n130 4.5005
R21851 CSoutput.n158 CSoutput.n134 4.5005
R21852 CSoutput.n158 CSoutput.n129 4.5005
R21853 CSoutput.n158 CSoutput.t187 4.5005
R21854 CSoutput.n158 CSoutput.n128 4.5005
R21855 CSoutput.n158 CSoutput.n135 4.5005
R21856 CSoutput.n158 CSoutput.n136 4.5005
R21857 CSoutput.n157 CSoutput.n131 4.5005
R21858 CSoutput.n157 CSoutput.n133 4.5005
R21859 CSoutput.n157 CSoutput.n130 4.5005
R21860 CSoutput.n157 CSoutput.n134 4.5005
R21861 CSoutput.n157 CSoutput.n129 4.5005
R21862 CSoutput.n157 CSoutput.t187 4.5005
R21863 CSoutput.n157 CSoutput.n128 4.5005
R21864 CSoutput.n157 CSoutput.n135 4.5005
R21865 CSoutput.n157 CSoutput.n136 4.5005
R21866 CSoutput.n140 CSoutput.n131 4.5005
R21867 CSoutput.n140 CSoutput.n133 4.5005
R21868 CSoutput.n140 CSoutput.n130 4.5005
R21869 CSoutput.n140 CSoutput.n134 4.5005
R21870 CSoutput.n140 CSoutput.n129 4.5005
R21871 CSoutput.n140 CSoutput.t187 4.5005
R21872 CSoutput.n140 CSoutput.n128 4.5005
R21873 CSoutput.n140 CSoutput.n135 4.5005
R21874 CSoutput.n140 CSoutput.n136 4.5005
R21875 CSoutput.n276 CSoutput.n131 4.5005
R21876 CSoutput.n276 CSoutput.n133 4.5005
R21877 CSoutput.n276 CSoutput.n130 4.5005
R21878 CSoutput.n276 CSoutput.n134 4.5005
R21879 CSoutput.n276 CSoutput.n129 4.5005
R21880 CSoutput.n276 CSoutput.t187 4.5005
R21881 CSoutput.n276 CSoutput.n128 4.5005
R21882 CSoutput.n276 CSoutput.n135 4.5005
R21883 CSoutput.n276 CSoutput.n136 4.5005
R21884 CSoutput.n323 CSoutput.n307 4.10845
R21885 CSoutput.n125 CSoutput.n109 4.10845
R21886 CSoutput.n321 CSoutput.t77 4.06363
R21887 CSoutput.n321 CSoutput.t10 4.06363
R21888 CSoutput.n319 CSoutput.t4 4.06363
R21889 CSoutput.n319 CSoutput.t46 4.06363
R21890 CSoutput.n317 CSoutput.t59 4.06363
R21891 CSoutput.n317 CSoutput.t79 4.06363
R21892 CSoutput.n315 CSoutput.t90 4.06363
R21893 CSoutput.n315 CSoutput.t21 4.06363
R21894 CSoutput.n313 CSoutput.t25 4.06363
R21895 CSoutput.n313 CSoutput.t80 4.06363
R21896 CSoutput.n311 CSoutput.t92 4.06363
R21897 CSoutput.n311 CSoutput.t93 4.06363
R21898 CSoutput.n309 CSoutput.t43 4.06363
R21899 CSoutput.n309 CSoutput.t44 4.06363
R21900 CSoutput.n308 CSoutput.t47 4.06363
R21901 CSoutput.n308 CSoutput.t94 4.06363
R21902 CSoutput.n305 CSoutput.t68 4.06363
R21903 CSoutput.n305 CSoutput.t95 4.06363
R21904 CSoutput.n303 CSoutput.t91 4.06363
R21905 CSoutput.n303 CSoutput.t33 4.06363
R21906 CSoutput.n301 CSoutput.t49 4.06363
R21907 CSoutput.n301 CSoutput.t69 4.06363
R21908 CSoutput.n299 CSoutput.t81 4.06363
R21909 CSoutput.n299 CSoutput.t9 4.06363
R21910 CSoutput.n297 CSoutput.t11 4.06363
R21911 CSoutput.n297 CSoutput.t72 4.06363
R21912 CSoutput.n295 CSoutput.t84 4.06363
R21913 CSoutput.n295 CSoutput.t85 4.06363
R21914 CSoutput.n293 CSoutput.t27 4.06363
R21915 CSoutput.n293 CSoutput.t28 4.06363
R21916 CSoutput.n292 CSoutput.t34 4.06363
R21917 CSoutput.n292 CSoutput.t86 4.06363
R21918 CSoutput.n290 CSoutput.t70 4.06363
R21919 CSoutput.n290 CSoutput.t31 4.06363
R21920 CSoutput.n288 CSoutput.t87 4.06363
R21921 CSoutput.n288 CSoutput.t53 4.06363
R21922 CSoutput.n286 CSoutput.t78 4.06363
R21923 CSoutput.n286 CSoutput.t40 4.06363
R21924 CSoutput.n284 CSoutput.t65 4.06363
R21925 CSoutput.n284 CSoutput.t20 4.06363
R21926 CSoutput.n282 CSoutput.t82 4.06363
R21927 CSoutput.n282 CSoutput.t15 4.06363
R21928 CSoutput.n280 CSoutput.t50 4.06363
R21929 CSoutput.n280 CSoutput.t29 4.06363
R21930 CSoutput.n278 CSoutput.t35 4.06363
R21931 CSoutput.n278 CSoutput.t12 4.06363
R21932 CSoutput.n277 CSoutput.t76 4.06363
R21933 CSoutput.n277 CSoutput.t6 4.06363
R21934 CSoutput.n110 CSoutput.t42 4.06363
R21935 CSoutput.n110 CSoutput.t97 4.06363
R21936 CSoutput.n111 CSoutput.t74 4.06363
R21937 CSoutput.n111 CSoutput.t73 4.06363
R21938 CSoutput.n113 CSoutput.t61 4.06363
R21939 CSoutput.n113 CSoutput.t39 4.06363
R21940 CSoutput.n115 CSoutput.t19 4.06363
R21941 CSoutput.n115 CSoutput.t62 4.06363
R21942 CSoutput.n117 CSoutput.t60 4.06363
R21943 CSoutput.n117 CSoutput.t36 4.06363
R21944 CSoutput.n119 CSoutput.t18 4.06363
R21945 CSoutput.n119 CSoutput.t17 4.06363
R21946 CSoutput.n121 CSoutput.t75 4.06363
R21947 CSoutput.n121 CSoutput.t48 4.06363
R21948 CSoutput.n123 CSoutput.t45 4.06363
R21949 CSoutput.n123 CSoutput.t13 4.06363
R21950 CSoutput.n94 CSoutput.t26 4.06363
R21951 CSoutput.n94 CSoutput.t89 4.06363
R21952 CSoutput.n95 CSoutput.t64 4.06363
R21953 CSoutput.n95 CSoutput.t63 4.06363
R21954 CSoutput.n97 CSoutput.t55 4.06363
R21955 CSoutput.n97 CSoutput.t24 4.06363
R21956 CSoutput.n99 CSoutput.t7 4.06363
R21957 CSoutput.n99 CSoutput.t56 4.06363
R21958 CSoutput.n101 CSoutput.t52 4.06363
R21959 CSoutput.n101 CSoutput.t22 4.06363
R21960 CSoutput.n103 CSoutput.t5 4.06363
R21961 CSoutput.n103 CSoutput.t3 4.06363
R21962 CSoutput.n105 CSoutput.t67 4.06363
R21963 CSoutput.n105 CSoutput.t38 4.06363
R21964 CSoutput.n107 CSoutput.t32 4.06363
R21965 CSoutput.n107 CSoutput.t2 4.06363
R21966 CSoutput.n79 CSoutput.t8 4.06363
R21967 CSoutput.n79 CSoutput.t57 4.06363
R21968 CSoutput.n80 CSoutput.t14 4.06363
R21969 CSoutput.n80 CSoutput.t37 4.06363
R21970 CSoutput.n82 CSoutput.t96 4.06363
R21971 CSoutput.n82 CSoutput.t51 4.06363
R21972 CSoutput.n84 CSoutput.t16 4.06363
R21973 CSoutput.n84 CSoutput.t83 4.06363
R21974 CSoutput.n86 CSoutput.t23 4.06363
R21975 CSoutput.n86 CSoutput.t66 4.06363
R21976 CSoutput.n88 CSoutput.t41 4.06363
R21977 CSoutput.n88 CSoutput.t58 4.06363
R21978 CSoutput.n90 CSoutput.t54 4.06363
R21979 CSoutput.n90 CSoutput.t88 4.06363
R21980 CSoutput.n92 CSoutput.t30 4.06363
R21981 CSoutput.n92 CSoutput.t71 4.06363
R21982 CSoutput.n44 CSoutput.n43 3.79402
R21983 CSoutput.n49 CSoutput.n48 3.79402
R21984 CSoutput.n404 CSoutput.n364 3.71319
R21985 CSoutput.n405 CSoutput.n404 3.57343
R21986 CSoutput.n361 CSoutput.t138 2.82907
R21987 CSoutput.n361 CSoutput.t118 2.82907
R21988 CSoutput.n359 CSoutput.t114 2.82907
R21989 CSoutput.n359 CSoutput.t1 2.82907
R21990 CSoutput.n357 CSoutput.t157 2.82907
R21991 CSoutput.n357 CSoutput.t120 2.82907
R21992 CSoutput.n355 CSoutput.t116 2.82907
R21993 CSoutput.n355 CSoutput.t110 2.82907
R21994 CSoutput.n353 CSoutput.t168 2.82907
R21995 CSoutput.n353 CSoutput.t152 2.82907
R21996 CSoutput.n351 CSoutput.t106 2.82907
R21997 CSoutput.n351 CSoutput.t145 2.82907
R21998 CSoutput.n349 CSoutput.t137 2.82907
R21999 CSoutput.n349 CSoutput.t105 2.82907
R22000 CSoutput.n347 CSoutput.t107 2.82907
R22001 CSoutput.n347 CSoutput.t103 2.82907
R22002 CSoutput.n345 CSoutput.t98 2.82907
R22003 CSoutput.n345 CSoutput.t119 2.82907
R22004 CSoutput.n344 CSoutput.t117 2.82907
R22005 CSoutput.n344 CSoutput.t111 2.82907
R22006 CSoutput.n342 CSoutput.t134 2.82907
R22007 CSoutput.n342 CSoutput.t149 2.82907
R22008 CSoutput.n340 CSoutput.t173 2.82907
R22009 CSoutput.n340 CSoutput.t121 2.82907
R22010 CSoutput.n338 CSoutput.t150 2.82907
R22011 CSoutput.n338 CSoutput.t115 2.82907
R22012 CSoutput.n336 CSoutput.t162 2.82907
R22013 CSoutput.n336 CSoutput.t102 2.82907
R22014 CSoutput.n334 CSoutput.t158 2.82907
R22015 CSoutput.n334 CSoutput.t147 2.82907
R22016 CSoutput.n332 CSoutput.t166 2.82907
R22017 CSoutput.n332 CSoutput.t123 2.82907
R22018 CSoutput.n330 CSoutput.t133 2.82907
R22019 CSoutput.n330 CSoutput.t156 2.82907
R22020 CSoutput.n328 CSoutput.t160 2.82907
R22021 CSoutput.n328 CSoutput.t99 2.82907
R22022 CSoutput.n326 CSoutput.t125 2.82907
R22023 CSoutput.n326 CSoutput.t153 2.82907
R22024 CSoutput.n325 CSoutput.t129 2.82907
R22025 CSoutput.n325 CSoutput.t146 2.82907
R22026 CSoutput.n384 CSoutput.t128 2.82907
R22027 CSoutput.n384 CSoutput.t148 2.82907
R22028 CSoutput.n385 CSoutput.t151 2.82907
R22029 CSoutput.n385 CSoutput.t170 2.82907
R22030 CSoutput.n387 CSoutput.t143 2.82907
R22031 CSoutput.n387 CSoutput.t100 2.82907
R22032 CSoutput.n389 CSoutput.t155 2.82907
R22033 CSoutput.n389 CSoutput.t140 2.82907
R22034 CSoutput.n391 CSoutput.t167 2.82907
R22035 CSoutput.n391 CSoutput.t163 2.82907
R22036 CSoutput.n393 CSoutput.t175 2.82907
R22037 CSoutput.n393 CSoutput.t124 2.82907
R22038 CSoutput.n395 CSoutput.t141 2.82907
R22039 CSoutput.n395 CSoutput.t109 2.82907
R22040 CSoutput.n397 CSoutput.t154 2.82907
R22041 CSoutput.n397 CSoutput.t136 2.82907
R22042 CSoutput.n399 CSoutput.t122 2.82907
R22043 CSoutput.n399 CSoutput.t112 2.82907
R22044 CSoutput.n401 CSoutput.t131 2.82907
R22045 CSoutput.n401 CSoutput.t135 2.82907
R22046 CSoutput.n365 CSoutput.t171 2.82907
R22047 CSoutput.n365 CSoutput.t0 2.82907
R22048 CSoutput.n366 CSoutput.t108 2.82907
R22049 CSoutput.n366 CSoutput.t164 2.82907
R22050 CSoutput.n368 CSoutput.t139 2.82907
R22051 CSoutput.n368 CSoutput.t144 2.82907
R22052 CSoutput.n370 CSoutput.t130 2.82907
R22053 CSoutput.n370 CSoutput.t159 2.82907
R22054 CSoutput.n372 CSoutput.t165 2.82907
R22055 CSoutput.n372 CSoutput.t172 2.82907
R22056 CSoutput.n374 CSoutput.t127 2.82907
R22057 CSoutput.n374 CSoutput.t104 2.82907
R22058 CSoutput.n376 CSoutput.t169 2.82907
R22059 CSoutput.n376 CSoutput.t174 2.82907
R22060 CSoutput.n378 CSoutput.t113 2.82907
R22061 CSoutput.n378 CSoutput.t132 2.82907
R22062 CSoutput.n380 CSoutput.t126 2.82907
R22063 CSoutput.n380 CSoutput.t142 2.82907
R22064 CSoutput.n382 CSoutput.t161 2.82907
R22065 CSoutput.n382 CSoutput.t101 2.82907
R22066 CSoutput.n324 CSoutput.n126 2.78353
R22067 CSoutput.n75 CSoutput.n1 2.45513
R22068 CSoutput.n217 CSoutput.n215 2.251
R22069 CSoutput.n217 CSoutput.n214 2.251
R22070 CSoutput.n217 CSoutput.n213 2.251
R22071 CSoutput.n217 CSoutput.n212 2.251
R22072 CSoutput.n186 CSoutput.n185 2.251
R22073 CSoutput.n186 CSoutput.n184 2.251
R22074 CSoutput.n186 CSoutput.n183 2.251
R22075 CSoutput.n186 CSoutput.n182 2.251
R22076 CSoutput.n259 CSoutput.n258 2.251
R22077 CSoutput.n224 CSoutput.n222 2.251
R22078 CSoutput.n224 CSoutput.n221 2.251
R22079 CSoutput.n224 CSoutput.n220 2.251
R22080 CSoutput.n242 CSoutput.n224 2.251
R22081 CSoutput.n230 CSoutput.n229 2.251
R22082 CSoutput.n230 CSoutput.n228 2.251
R22083 CSoutput.n230 CSoutput.n227 2.251
R22084 CSoutput.n230 CSoutput.n226 2.251
R22085 CSoutput.n256 CSoutput.n196 2.251
R22086 CSoutput.n251 CSoutput.n249 2.251
R22087 CSoutput.n251 CSoutput.n248 2.251
R22088 CSoutput.n251 CSoutput.n247 2.251
R22089 CSoutput.n251 CSoutput.n246 2.251
R22090 CSoutput.n152 CSoutput.n151 2.251
R22091 CSoutput.n152 CSoutput.n150 2.251
R22092 CSoutput.n152 CSoutput.n149 2.251
R22093 CSoutput.n152 CSoutput.n148 2.251
R22094 CSoutput.n269 CSoutput.n268 2.251
R22095 CSoutput.n186 CSoutput.n166 2.2505
R22096 CSoutput.n181 CSoutput.n166 2.2505
R22097 CSoutput.n179 CSoutput.n166 2.2505
R22098 CSoutput.n178 CSoutput.n166 2.2505
R22099 CSoutput.n263 CSoutput.n166 2.2505
R22100 CSoutput.n261 CSoutput.n166 2.2505
R22101 CSoutput.n259 CSoutput.n166 2.2505
R22102 CSoutput.n189 CSoutput.n166 2.2505
R22103 CSoutput.n188 CSoutput.n166 2.2505
R22104 CSoutput.n192 CSoutput.n166 2.2505
R22105 CSoutput.n191 CSoutput.n166 2.2505
R22106 CSoutput.n174 CSoutput.n166 2.2505
R22107 CSoutput.n266 CSoutput.n166 2.2505
R22108 CSoutput.n266 CSoutput.n265 2.2505
R22109 CSoutput.n230 CSoutput.n201 2.2505
R22110 CSoutput.n211 CSoutput.n201 2.2505
R22111 CSoutput.n232 CSoutput.n201 2.2505
R22112 CSoutput.n210 CSoutput.n201 2.2505
R22113 CSoutput.n234 CSoutput.n201 2.2505
R22114 CSoutput.n201 CSoutput.n195 2.2505
R22115 CSoutput.n256 CSoutput.n201 2.2505
R22116 CSoutput.n254 CSoutput.n201 2.2505
R22117 CSoutput.n236 CSoutput.n201 2.2505
R22118 CSoutput.n208 CSoutput.n201 2.2505
R22119 CSoutput.n238 CSoutput.n201 2.2505
R22120 CSoutput.n207 CSoutput.n201 2.2505
R22121 CSoutput.n252 CSoutput.n201 2.2505
R22122 CSoutput.n252 CSoutput.n205 2.2505
R22123 CSoutput.n152 CSoutput.n132 2.2505
R22124 CSoutput.n147 CSoutput.n132 2.2505
R22125 CSoutput.n145 CSoutput.n132 2.2505
R22126 CSoutput.n144 CSoutput.n132 2.2505
R22127 CSoutput.n273 CSoutput.n132 2.2505
R22128 CSoutput.n271 CSoutput.n132 2.2505
R22129 CSoutput.n269 CSoutput.n132 2.2505
R22130 CSoutput.n155 CSoutput.n132 2.2505
R22131 CSoutput.n154 CSoutput.n132 2.2505
R22132 CSoutput.n158 CSoutput.n132 2.2505
R22133 CSoutput.n157 CSoutput.n132 2.2505
R22134 CSoutput.n140 CSoutput.n132 2.2505
R22135 CSoutput.n276 CSoutput.n132 2.2505
R22136 CSoutput.n276 CSoutput.n275 2.2505
R22137 CSoutput.n194 CSoutput.n187 2.25024
R22138 CSoutput.n194 CSoutput.n180 2.25024
R22139 CSoutput.n262 CSoutput.n194 2.25024
R22140 CSoutput.n194 CSoutput.n190 2.25024
R22141 CSoutput.n194 CSoutput.n193 2.25024
R22142 CSoutput.n194 CSoutput.n161 2.25024
R22143 CSoutput.n244 CSoutput.n241 2.25024
R22144 CSoutput.n244 CSoutput.n240 2.25024
R22145 CSoutput.n244 CSoutput.n239 2.25024
R22146 CSoutput.n244 CSoutput.n206 2.25024
R22147 CSoutput.n244 CSoutput.n243 2.25024
R22148 CSoutput.n245 CSoutput.n244 2.25024
R22149 CSoutput.n160 CSoutput.n153 2.25024
R22150 CSoutput.n160 CSoutput.n146 2.25024
R22151 CSoutput.n272 CSoutput.n160 2.25024
R22152 CSoutput.n160 CSoutput.n156 2.25024
R22153 CSoutput.n160 CSoutput.n159 2.25024
R22154 CSoutput.n160 CSoutput.n127 2.25024
R22155 CSoutput.n261 CSoutput.n171 1.50111
R22156 CSoutput.n209 CSoutput.n195 1.50111
R22157 CSoutput.n271 CSoutput.n137 1.50111
R22158 CSoutput.n217 CSoutput.n216 1.501
R22159 CSoutput.n224 CSoutput.n223 1.501
R22160 CSoutput.n251 CSoutput.n250 1.501
R22161 CSoutput.n265 CSoutput.n176 1.12536
R22162 CSoutput.n265 CSoutput.n177 1.12536
R22163 CSoutput.n265 CSoutput.n264 1.12536
R22164 CSoutput.n225 CSoutput.n205 1.12536
R22165 CSoutput.n231 CSoutput.n205 1.12536
R22166 CSoutput.n233 CSoutput.n205 1.12536
R22167 CSoutput.n275 CSoutput.n142 1.12536
R22168 CSoutput.n275 CSoutput.n143 1.12536
R22169 CSoutput.n275 CSoutput.n274 1.12536
R22170 CSoutput.n265 CSoutput.n172 1.12536
R22171 CSoutput.n265 CSoutput.n173 1.12536
R22172 CSoutput.n265 CSoutput.n175 1.12536
R22173 CSoutput.n255 CSoutput.n205 1.12536
R22174 CSoutput.n235 CSoutput.n205 1.12536
R22175 CSoutput.n237 CSoutput.n205 1.12536
R22176 CSoutput.n275 CSoutput.n138 1.12536
R22177 CSoutput.n275 CSoutput.n139 1.12536
R22178 CSoutput.n275 CSoutput.n141 1.12536
R22179 CSoutput.n31 CSoutput.n30 0.669944
R22180 CSoutput.n62 CSoutput.n61 0.669944
R22181 CSoutput.n348 CSoutput.n346 0.573776
R22182 CSoutput.n350 CSoutput.n348 0.573776
R22183 CSoutput.n352 CSoutput.n350 0.573776
R22184 CSoutput.n354 CSoutput.n352 0.573776
R22185 CSoutput.n356 CSoutput.n354 0.573776
R22186 CSoutput.n358 CSoutput.n356 0.573776
R22187 CSoutput.n360 CSoutput.n358 0.573776
R22188 CSoutput.n362 CSoutput.n360 0.573776
R22189 CSoutput.n329 CSoutput.n327 0.573776
R22190 CSoutput.n331 CSoutput.n329 0.573776
R22191 CSoutput.n333 CSoutput.n331 0.573776
R22192 CSoutput.n335 CSoutput.n333 0.573776
R22193 CSoutput.n337 CSoutput.n335 0.573776
R22194 CSoutput.n339 CSoutput.n337 0.573776
R22195 CSoutput.n341 CSoutput.n339 0.573776
R22196 CSoutput.n343 CSoutput.n341 0.573776
R22197 CSoutput.n402 CSoutput.n400 0.573776
R22198 CSoutput.n400 CSoutput.n398 0.573776
R22199 CSoutput.n398 CSoutput.n396 0.573776
R22200 CSoutput.n396 CSoutput.n394 0.573776
R22201 CSoutput.n394 CSoutput.n392 0.573776
R22202 CSoutput.n392 CSoutput.n390 0.573776
R22203 CSoutput.n390 CSoutput.n388 0.573776
R22204 CSoutput.n388 CSoutput.n386 0.573776
R22205 CSoutput.n383 CSoutput.n381 0.573776
R22206 CSoutput.n381 CSoutput.n379 0.573776
R22207 CSoutput.n379 CSoutput.n377 0.573776
R22208 CSoutput.n377 CSoutput.n375 0.573776
R22209 CSoutput.n375 CSoutput.n373 0.573776
R22210 CSoutput.n373 CSoutput.n371 0.573776
R22211 CSoutput.n371 CSoutput.n369 0.573776
R22212 CSoutput.n369 CSoutput.n367 0.573776
R22213 CSoutput.n405 CSoutput.n276 0.53442
R22214 CSoutput.n312 CSoutput.n310 0.358259
R22215 CSoutput.n314 CSoutput.n312 0.358259
R22216 CSoutput.n316 CSoutput.n314 0.358259
R22217 CSoutput.n318 CSoutput.n316 0.358259
R22218 CSoutput.n320 CSoutput.n318 0.358259
R22219 CSoutput.n322 CSoutput.n320 0.358259
R22220 CSoutput.n296 CSoutput.n294 0.358259
R22221 CSoutput.n298 CSoutput.n296 0.358259
R22222 CSoutput.n300 CSoutput.n298 0.358259
R22223 CSoutput.n302 CSoutput.n300 0.358259
R22224 CSoutput.n304 CSoutput.n302 0.358259
R22225 CSoutput.n306 CSoutput.n304 0.358259
R22226 CSoutput.n281 CSoutput.n279 0.358259
R22227 CSoutput.n283 CSoutput.n281 0.358259
R22228 CSoutput.n285 CSoutput.n283 0.358259
R22229 CSoutput.n287 CSoutput.n285 0.358259
R22230 CSoutput.n289 CSoutput.n287 0.358259
R22231 CSoutput.n291 CSoutput.n289 0.358259
R22232 CSoutput.n124 CSoutput.n122 0.358259
R22233 CSoutput.n122 CSoutput.n120 0.358259
R22234 CSoutput.n120 CSoutput.n118 0.358259
R22235 CSoutput.n118 CSoutput.n116 0.358259
R22236 CSoutput.n116 CSoutput.n114 0.358259
R22237 CSoutput.n114 CSoutput.n112 0.358259
R22238 CSoutput.n108 CSoutput.n106 0.358259
R22239 CSoutput.n106 CSoutput.n104 0.358259
R22240 CSoutput.n104 CSoutput.n102 0.358259
R22241 CSoutput.n102 CSoutput.n100 0.358259
R22242 CSoutput.n100 CSoutput.n98 0.358259
R22243 CSoutput.n98 CSoutput.n96 0.358259
R22244 CSoutput.n93 CSoutput.n91 0.358259
R22245 CSoutput.n91 CSoutput.n89 0.358259
R22246 CSoutput.n89 CSoutput.n87 0.358259
R22247 CSoutput.n87 CSoutput.n85 0.358259
R22248 CSoutput.n85 CSoutput.n83 0.358259
R22249 CSoutput.n83 CSoutput.n81 0.358259
R22250 CSoutput.n21 CSoutput.n20 0.169105
R22251 CSoutput.n21 CSoutput.n16 0.169105
R22252 CSoutput.n26 CSoutput.n16 0.169105
R22253 CSoutput.n27 CSoutput.n26 0.169105
R22254 CSoutput.n27 CSoutput.n14 0.169105
R22255 CSoutput.n32 CSoutput.n14 0.169105
R22256 CSoutput.n33 CSoutput.n32 0.169105
R22257 CSoutput.n34 CSoutput.n33 0.169105
R22258 CSoutput.n34 CSoutput.n12 0.169105
R22259 CSoutput.n39 CSoutput.n12 0.169105
R22260 CSoutput.n40 CSoutput.n39 0.169105
R22261 CSoutput.n40 CSoutput.n10 0.169105
R22262 CSoutput.n45 CSoutput.n10 0.169105
R22263 CSoutput.n46 CSoutput.n45 0.169105
R22264 CSoutput.n47 CSoutput.n46 0.169105
R22265 CSoutput.n47 CSoutput.n8 0.169105
R22266 CSoutput.n52 CSoutput.n8 0.169105
R22267 CSoutput.n53 CSoutput.n52 0.169105
R22268 CSoutput.n53 CSoutput.n6 0.169105
R22269 CSoutput.n58 CSoutput.n6 0.169105
R22270 CSoutput.n59 CSoutput.n58 0.169105
R22271 CSoutput.n60 CSoutput.n59 0.169105
R22272 CSoutput.n60 CSoutput.n4 0.169105
R22273 CSoutput.n66 CSoutput.n4 0.169105
R22274 CSoutput.n67 CSoutput.n66 0.169105
R22275 CSoutput.n68 CSoutput.n67 0.169105
R22276 CSoutput.n68 CSoutput.n2 0.169105
R22277 CSoutput.n73 CSoutput.n2 0.169105
R22278 CSoutput.n74 CSoutput.n73 0.169105
R22279 CSoutput.n74 CSoutput.n0 0.169105
R22280 CSoutput.n78 CSoutput.n0 0.169105
R22281 CSoutput.n219 CSoutput.n218 0.0910737
R22282 CSoutput.n270 CSoutput.n267 0.0723685
R22283 CSoutput.n224 CSoutput.n219 0.0522944
R22284 CSoutput.n267 CSoutput.n266 0.0499135
R22285 CSoutput.n218 CSoutput.n217 0.0499135
R22286 CSoutput.n252 CSoutput.n251 0.0464294
R22287 CSoutput.n260 CSoutput.n257 0.0391444
R22288 CSoutput.n219 CSoutput.t192 0.023435
R22289 CSoutput.n267 CSoutput.t181 0.02262
R22290 CSoutput.n218 CSoutput.t190 0.02262
R22291 CSoutput CSoutput.n405 0.0052
R22292 CSoutput.n189 CSoutput.n172 0.00365111
R22293 CSoutput.n192 CSoutput.n173 0.00365111
R22294 CSoutput.n175 CSoutput.n174 0.00365111
R22295 CSoutput.n217 CSoutput.n176 0.00365111
R22296 CSoutput.n181 CSoutput.n177 0.00365111
R22297 CSoutput.n264 CSoutput.n178 0.00365111
R22298 CSoutput.n255 CSoutput.n254 0.00365111
R22299 CSoutput.n235 CSoutput.n208 0.00365111
R22300 CSoutput.n237 CSoutput.n207 0.00365111
R22301 CSoutput.n225 CSoutput.n224 0.00365111
R22302 CSoutput.n231 CSoutput.n211 0.00365111
R22303 CSoutput.n233 CSoutput.n210 0.00365111
R22304 CSoutput.n155 CSoutput.n138 0.00365111
R22305 CSoutput.n158 CSoutput.n139 0.00365111
R22306 CSoutput.n141 CSoutput.n140 0.00365111
R22307 CSoutput.n251 CSoutput.n142 0.00365111
R22308 CSoutput.n147 CSoutput.n143 0.00365111
R22309 CSoutput.n274 CSoutput.n144 0.00365111
R22310 CSoutput.n186 CSoutput.n176 0.00340054
R22311 CSoutput.n179 CSoutput.n177 0.00340054
R22312 CSoutput.n264 CSoutput.n263 0.00340054
R22313 CSoutput.n259 CSoutput.n172 0.00340054
R22314 CSoutput.n188 CSoutput.n173 0.00340054
R22315 CSoutput.n191 CSoutput.n175 0.00340054
R22316 CSoutput.n230 CSoutput.n225 0.00340054
R22317 CSoutput.n232 CSoutput.n231 0.00340054
R22318 CSoutput.n234 CSoutput.n233 0.00340054
R22319 CSoutput.n256 CSoutput.n255 0.00340054
R22320 CSoutput.n236 CSoutput.n235 0.00340054
R22321 CSoutput.n238 CSoutput.n237 0.00340054
R22322 CSoutput.n152 CSoutput.n142 0.00340054
R22323 CSoutput.n145 CSoutput.n143 0.00340054
R22324 CSoutput.n274 CSoutput.n273 0.00340054
R22325 CSoutput.n269 CSoutput.n138 0.00340054
R22326 CSoutput.n154 CSoutput.n139 0.00340054
R22327 CSoutput.n157 CSoutput.n141 0.00340054
R22328 CSoutput.n187 CSoutput.n181 0.00252698
R22329 CSoutput.n180 CSoutput.n178 0.00252698
R22330 CSoutput.n262 CSoutput.n261 0.00252698
R22331 CSoutput.n190 CSoutput.n188 0.00252698
R22332 CSoutput.n193 CSoutput.n191 0.00252698
R22333 CSoutput.n266 CSoutput.n161 0.00252698
R22334 CSoutput.n187 CSoutput.n186 0.00252698
R22335 CSoutput.n180 CSoutput.n179 0.00252698
R22336 CSoutput.n263 CSoutput.n262 0.00252698
R22337 CSoutput.n190 CSoutput.n189 0.00252698
R22338 CSoutput.n193 CSoutput.n192 0.00252698
R22339 CSoutput.n174 CSoutput.n161 0.00252698
R22340 CSoutput.n241 CSoutput.n211 0.00252698
R22341 CSoutput.n240 CSoutput.n210 0.00252698
R22342 CSoutput.n239 CSoutput.n195 0.00252698
R22343 CSoutput.n236 CSoutput.n206 0.00252698
R22344 CSoutput.n243 CSoutput.n238 0.00252698
R22345 CSoutput.n252 CSoutput.n245 0.00252698
R22346 CSoutput.n241 CSoutput.n230 0.00252698
R22347 CSoutput.n240 CSoutput.n232 0.00252698
R22348 CSoutput.n239 CSoutput.n234 0.00252698
R22349 CSoutput.n254 CSoutput.n206 0.00252698
R22350 CSoutput.n243 CSoutput.n208 0.00252698
R22351 CSoutput.n245 CSoutput.n207 0.00252698
R22352 CSoutput.n153 CSoutput.n147 0.00252698
R22353 CSoutput.n146 CSoutput.n144 0.00252698
R22354 CSoutput.n272 CSoutput.n271 0.00252698
R22355 CSoutput.n156 CSoutput.n154 0.00252698
R22356 CSoutput.n159 CSoutput.n157 0.00252698
R22357 CSoutput.n276 CSoutput.n127 0.00252698
R22358 CSoutput.n153 CSoutput.n152 0.00252698
R22359 CSoutput.n146 CSoutput.n145 0.00252698
R22360 CSoutput.n273 CSoutput.n272 0.00252698
R22361 CSoutput.n156 CSoutput.n155 0.00252698
R22362 CSoutput.n159 CSoutput.n158 0.00252698
R22363 CSoutput.n140 CSoutput.n127 0.00252698
R22364 CSoutput.n261 CSoutput.n260 0.0020275
R22365 CSoutput.n260 CSoutput.n259 0.0020275
R22366 CSoutput.n257 CSoutput.n195 0.0020275
R22367 CSoutput.n257 CSoutput.n256 0.0020275
R22368 CSoutput.n271 CSoutput.n270 0.0020275
R22369 CSoutput.n270 CSoutput.n269 0.0020275
R22370 CSoutput.n171 CSoutput.n170 0.00166668
R22371 CSoutput.n253 CSoutput.n209 0.00166668
R22372 CSoutput.n137 CSoutput.n136 0.00166668
R22373 CSoutput.n275 CSoutput.n137 0.00133328
R22374 CSoutput.n209 CSoutput.n205 0.00133328
R22375 CSoutput.n265 CSoutput.n171 0.00133328
R22376 CSoutput.n268 CSoutput.n160 0.001
R22377 CSoutput.n246 CSoutput.n160 0.001
R22378 CSoutput.n148 CSoutput.n128 0.001
R22379 CSoutput.n247 CSoutput.n128 0.001
R22380 CSoutput.n149 CSoutput.n129 0.001
R22381 CSoutput.n248 CSoutput.n129 0.001
R22382 CSoutput.n150 CSoutput.n130 0.001
R22383 CSoutput.n249 CSoutput.n130 0.001
R22384 CSoutput.n151 CSoutput.n131 0.001
R22385 CSoutput.n250 CSoutput.n131 0.001
R22386 CSoutput.n244 CSoutput.n196 0.001
R22387 CSoutput.n244 CSoutput.n242 0.001
R22388 CSoutput.n226 CSoutput.n197 0.001
R22389 CSoutput.n220 CSoutput.n197 0.001
R22390 CSoutput.n227 CSoutput.n198 0.001
R22391 CSoutput.n221 CSoutput.n198 0.001
R22392 CSoutput.n228 CSoutput.n199 0.001
R22393 CSoutput.n222 CSoutput.n199 0.001
R22394 CSoutput.n229 CSoutput.n200 0.001
R22395 CSoutput.n223 CSoutput.n200 0.001
R22396 CSoutput.n258 CSoutput.n194 0.001
R22397 CSoutput.n212 CSoutput.n194 0.001
R22398 CSoutput.n182 CSoutput.n162 0.001
R22399 CSoutput.n213 CSoutput.n162 0.001
R22400 CSoutput.n183 CSoutput.n163 0.001
R22401 CSoutput.n214 CSoutput.n163 0.001
R22402 CSoutput.n184 CSoutput.n164 0.001
R22403 CSoutput.n215 CSoutput.n164 0.001
R22404 CSoutput.n185 CSoutput.n165 0.001
R22405 CSoutput.n216 CSoutput.n165 0.001
R22406 CSoutput.n216 CSoutput.n166 0.001
R22407 CSoutput.n215 CSoutput.n167 0.001
R22408 CSoutput.n214 CSoutput.n168 0.001
R22409 CSoutput.n213 CSoutput.t184 0.001
R22410 CSoutput.n212 CSoutput.n169 0.001
R22411 CSoutput.n185 CSoutput.n167 0.001
R22412 CSoutput.n184 CSoutput.n168 0.001
R22413 CSoutput.n183 CSoutput.t184 0.001
R22414 CSoutput.n182 CSoutput.n169 0.001
R22415 CSoutput.n258 CSoutput.n170 0.001
R22416 CSoutput.n223 CSoutput.n201 0.001
R22417 CSoutput.n222 CSoutput.n202 0.001
R22418 CSoutput.n221 CSoutput.n203 0.001
R22419 CSoutput.n220 CSoutput.t186 0.001
R22420 CSoutput.n242 CSoutput.n204 0.001
R22421 CSoutput.n229 CSoutput.n202 0.001
R22422 CSoutput.n228 CSoutput.n203 0.001
R22423 CSoutput.n227 CSoutput.t186 0.001
R22424 CSoutput.n226 CSoutput.n204 0.001
R22425 CSoutput.n253 CSoutput.n196 0.001
R22426 CSoutput.n250 CSoutput.n132 0.001
R22427 CSoutput.n249 CSoutput.n133 0.001
R22428 CSoutput.n248 CSoutput.n134 0.001
R22429 CSoutput.n247 CSoutput.t187 0.001
R22430 CSoutput.n246 CSoutput.n135 0.001
R22431 CSoutput.n151 CSoutput.n133 0.001
R22432 CSoutput.n150 CSoutput.n134 0.001
R22433 CSoutput.n149 CSoutput.t187 0.001
R22434 CSoutput.n148 CSoutput.n135 0.001
R22435 CSoutput.n268 CSoutput.n136 0.001
R22436 a_n2650_13878.n110 a_n2650_13878.t84 512.366
R22437 a_n2650_13878.n100 a_n2650_13878.t74 512.366
R22438 a_n2650_13878.n111 a_n2650_13878.t64 512.366
R22439 a_n2650_13878.n108 a_n2650_13878.t92 512.366
R22440 a_n2650_13878.n101 a_n2650_13878.t81 512.366
R22441 a_n2650_13878.n109 a_n2650_13878.t80 512.366
R22442 a_n2650_13878.n106 a_n2650_13878.t88 512.366
R22443 a_n2650_13878.n102 a_n2650_13878.t72 512.366
R22444 a_n2650_13878.n107 a_n2650_13878.t73 512.366
R22445 a_n2650_13878.n104 a_n2650_13878.t75 512.366
R22446 a_n2650_13878.n103 a_n2650_13878.t86 512.366
R22447 a_n2650_13878.n105 a_n2650_13878.t99 512.366
R22448 a_n2650_13878.n118 a_n2650_13878.t98 512.366
R22449 a_n2650_13878.n117 a_n2650_13878.t77 512.366
R22450 a_n2650_13878.n74 a_n2650_13878.t82 512.366
R22451 a_n2650_13878.n116 a_n2650_13878.t71 512.366
R22452 a_n2650_13878.n115 a_n2650_13878.t87 512.366
R22453 a_n2650_13878.n75 a_n2650_13878.t95 512.366
R22454 a_n2650_13878.n114 a_n2650_13878.t96 512.366
R22455 a_n2650_13878.n113 a_n2650_13878.t66 512.366
R22456 a_n2650_13878.n76 a_n2650_13878.t79 512.366
R22457 a_n2650_13878.n41 a_n2650_13878.t17 533.335
R22458 a_n2650_13878.n119 a_n2650_13878.t33 512.366
R22459 a_n2650_13878.n132 a_n2650_13878.t37 512.366
R22460 a_n2650_13878.n137 a_n2650_13878.t29 512.366
R22461 a_n2650_13878.n136 a_n2650_13878.t7 512.366
R22462 a_n2650_13878.n72 a_n2650_13878.t25 512.366
R22463 a_n2650_13878.n135 a_n2650_13878.t27 512.366
R22464 a_n2650_13878.n134 a_n2650_13878.t13 512.366
R22465 a_n2650_13878.n73 a_n2650_13878.t3 512.366
R22466 a_n2650_13878.n133 a_n2650_13878.t9 512.366
R22467 a_n2650_13878.n92 a_n2650_13878.t35 512.366
R22468 a_n2650_13878.n93 a_n2650_13878.t11 512.366
R22469 a_n2650_13878.n82 a_n2650_13878.t19 512.366
R22470 a_n2650_13878.n94 a_n2650_13878.t23 512.366
R22471 a_n2650_13878.n95 a_n2650_13878.t41 512.366
R22472 a_n2650_13878.n96 a_n2650_13878.t5 512.366
R22473 a_n2650_13878.n97 a_n2650_13878.t21 512.366
R22474 a_n2650_13878.n81 a_n2650_13878.t15 512.366
R22475 a_n2650_13878.n98 a_n2650_13878.t39 512.366
R22476 a_n2650_13878.n85 a_n2650_13878.t70 512.366
R22477 a_n2650_13878.n86 a_n2650_13878.t93 512.366
R22478 a_n2650_13878.n84 a_n2650_13878.t94 512.366
R22479 a_n2650_13878.n87 a_n2650_13878.t68 512.366
R22480 a_n2650_13878.n88 a_n2650_13878.t90 512.366
R22481 a_n2650_13878.n89 a_n2650_13878.t91 512.366
R22482 a_n2650_13878.n90 a_n2650_13878.t65 512.366
R22483 a_n2650_13878.n83 a_n2650_13878.t76 512.366
R22484 a_n2650_13878.n91 a_n2650_13878.t85 512.366
R22485 a_n2650_13878.n5 a_n2650_13878.n70 70.1674
R22486 a_n2650_13878.n7 a_n2650_13878.n68 70.1674
R22487 a_n2650_13878.n9 a_n2650_13878.n66 70.1674
R22488 a_n2650_13878.n12 a_n2650_13878.n64 70.1674
R22489 a_n2650_13878.n23 a_n2650_13878.n48 70.1674
R22490 a_n2650_13878.n40 a_n2650_13878.n27 80.4688
R22491 a_n2650_13878.n40 a_n2650_13878.n133 0.365327
R22492 a_n2650_13878.n27 a_n2650_13878.n39 75.0448
R22493 a_n2650_13878.n38 a_n2650_13878.n26 70.1674
R22494 a_n2650_13878.n135 a_n2650_13878.n38 20.9683
R22495 a_n2650_13878.n26 a_n2650_13878.n37 70.3058
R22496 a_n2650_13878.n37 a_n2650_13878.n72 20.6913
R22497 a_n2650_13878.n36 a_n2650_13878.n28 75.3623
R22498 a_n2650_13878.n136 a_n2650_13878.n36 10.5784
R22499 a_n2650_13878.n28 a_n2650_13878.n137 161.3
R22500 a_n2650_13878.n132 a_n2650_13878.n71 11.843
R22501 a_n2650_13878.n41 a_n2650_13878.n35 70.1674
R22502 a_n2650_13878.n41 a_n2650_13878.n119 20.9683
R22503 a_n2650_13878.n27 a_n2650_13878.n71 74.73
R22504 a_n2650_13878.n48 a_n2650_13878.n76 20.9683
R22505 a_n2650_13878.n47 a_n2650_13878.n23 74.73
R22506 a_n2650_13878.n113 a_n2650_13878.n47 11.843
R22507 a_n2650_13878.n46 a_n2650_13878.n22 80.4688
R22508 a_n2650_13878.n46 a_n2650_13878.n114 0.365327
R22509 a_n2650_13878.n22 a_n2650_13878.n45 75.0448
R22510 a_n2650_13878.n44 a_n2650_13878.n24 70.1674
R22511 a_n2650_13878.n116 a_n2650_13878.n44 20.9683
R22512 a_n2650_13878.n24 a_n2650_13878.n43 70.3058
R22513 a_n2650_13878.n43 a_n2650_13878.n74 20.6913
R22514 a_n2650_13878.n42 a_n2650_13878.n25 75.3623
R22515 a_n2650_13878.n117 a_n2650_13878.n42 10.5784
R22516 a_n2650_13878.n25 a_n2650_13878.n118 161.3
R22517 a_n2650_13878.n15 a_n2650_13878.n62 70.1674
R22518 a_n2650_13878.n19 a_n2650_13878.n55 70.1674
R22519 a_n2650_13878.n91 a_n2650_13878.n55 20.9683
R22520 a_n2650_13878.n54 a_n2650_13878.n19 74.73
R22521 a_n2650_13878.n54 a_n2650_13878.n83 11.843
R22522 a_n2650_13878.n18 a_n2650_13878.n53 80.4688
R22523 a_n2650_13878.n90 a_n2650_13878.n53 0.365327
R22524 a_n2650_13878.n52 a_n2650_13878.n18 75.0448
R22525 a_n2650_13878.n20 a_n2650_13878.n51 70.1674
R22526 a_n2650_13878.n87 a_n2650_13878.n51 20.9683
R22527 a_n2650_13878.n50 a_n2650_13878.n20 70.3058
R22528 a_n2650_13878.n50 a_n2650_13878.n84 20.6913
R22529 a_n2650_13878.n21 a_n2650_13878.n49 75.3623
R22530 a_n2650_13878.n86 a_n2650_13878.n49 10.5784
R22531 a_n2650_13878.n85 a_n2650_13878.n21 161.3
R22532 a_n2650_13878.n98 a_n2650_13878.n62 20.9683
R22533 a_n2650_13878.n61 a_n2650_13878.n15 74.73
R22534 a_n2650_13878.n61 a_n2650_13878.n81 11.843
R22535 a_n2650_13878.n14 a_n2650_13878.n60 80.4688
R22536 a_n2650_13878.n97 a_n2650_13878.n60 0.365327
R22537 a_n2650_13878.n59 a_n2650_13878.n14 75.0448
R22538 a_n2650_13878.n16 a_n2650_13878.n58 70.1674
R22539 a_n2650_13878.n94 a_n2650_13878.n58 20.9683
R22540 a_n2650_13878.n57 a_n2650_13878.n16 70.3058
R22541 a_n2650_13878.n57 a_n2650_13878.n82 20.6913
R22542 a_n2650_13878.n17 a_n2650_13878.n56 75.3623
R22543 a_n2650_13878.n93 a_n2650_13878.n56 10.5784
R22544 a_n2650_13878.n92 a_n2650_13878.n17 161.3
R22545 a_n2650_13878.n105 a_n2650_13878.n64 20.9683
R22546 a_n2650_13878.n63 a_n2650_13878.n13 75.0448
R22547 a_n2650_13878.n63 a_n2650_13878.n103 11.2134
R22548 a_n2650_13878.n13 a_n2650_13878.n104 161.3
R22549 a_n2650_13878.n107 a_n2650_13878.n66 20.9683
R22550 a_n2650_13878.n65 a_n2650_13878.n10 75.0448
R22551 a_n2650_13878.n65 a_n2650_13878.n102 11.2134
R22552 a_n2650_13878.n10 a_n2650_13878.n106 161.3
R22553 a_n2650_13878.n109 a_n2650_13878.n68 20.9683
R22554 a_n2650_13878.n67 a_n2650_13878.n8 75.0448
R22555 a_n2650_13878.n67 a_n2650_13878.n101 11.2134
R22556 a_n2650_13878.n8 a_n2650_13878.n108 161.3
R22557 a_n2650_13878.n111 a_n2650_13878.n70 20.9683
R22558 a_n2650_13878.n69 a_n2650_13878.n6 75.0448
R22559 a_n2650_13878.n69 a_n2650_13878.n100 11.2134
R22560 a_n2650_13878.n6 a_n2650_13878.n110 161.3
R22561 a_n2650_13878.n3 a_n2650_13878.n129 81.3764
R22562 a_n2650_13878.n4 a_n2650_13878.n123 81.3764
R22563 a_n2650_13878.n0 a_n2650_13878.n120 81.3764
R22564 a_n2650_13878.n3 a_n2650_13878.n130 80.9324
R22565 a_n2650_13878.n2 a_n2650_13878.n131 80.9324
R22566 a_n2650_13878.n2 a_n2650_13878.n128 80.9324
R22567 a_n2650_13878.n2 a_n2650_13878.n127 80.9324
R22568 a_n2650_13878.n1 a_n2650_13878.n126 80.9324
R22569 a_n2650_13878.n4 a_n2650_13878.n124 80.9324
R22570 a_n2650_13878.n0 a_n2650_13878.n125 80.9324
R22571 a_n2650_13878.n0 a_n2650_13878.n122 80.9324
R22572 a_n2650_13878.n0 a_n2650_13878.n121 80.9324
R22573 a_n2650_13878.n34 a_n2650_13878.t18 74.6477
R22574 a_n2650_13878.n29 a_n2650_13878.t36 74.6477
R22575 a_n2650_13878.n32 a_n2650_13878.t30 74.2899
R22576 a_n2650_13878.n31 a_n2650_13878.t32 74.2897
R22577 a_n2650_13878.n34 a_n2650_13878.n141 70.6783
R22578 a_n2650_13878.n33 a_n2650_13878.n140 70.6783
R22579 a_n2650_13878.n33 a_n2650_13878.n139 70.6783
R22580 a_n2650_13878.n31 a_n2650_13878.n80 70.6783
R22581 a_n2650_13878.n30 a_n2650_13878.n79 70.6783
R22582 a_n2650_13878.n30 a_n2650_13878.n78 70.6783
R22583 a_n2650_13878.n29 a_n2650_13878.n77 70.6783
R22584 a_n2650_13878.n142 a_n2650_13878.n34 70.6782
R22585 a_n2650_13878.n110 a_n2650_13878.n100 48.2005
R22586 a_n2650_13878.t89 a_n2650_13878.n70 533.335
R22587 a_n2650_13878.n108 a_n2650_13878.n101 48.2005
R22588 a_n2650_13878.t97 a_n2650_13878.n68 533.335
R22589 a_n2650_13878.n106 a_n2650_13878.n102 48.2005
R22590 a_n2650_13878.t83 a_n2650_13878.n66 533.335
R22591 a_n2650_13878.n104 a_n2650_13878.n103 48.2005
R22592 a_n2650_13878.t78 a_n2650_13878.n64 533.335
R22593 a_n2650_13878.n118 a_n2650_13878.n117 48.2005
R22594 a_n2650_13878.n44 a_n2650_13878.n115 20.9683
R22595 a_n2650_13878.n114 a_n2650_13878.n75 48.2005
R22596 a_n2650_13878.t69 a_n2650_13878.n48 533.335
R22597 a_n2650_13878.n137 a_n2650_13878.n136 48.2005
R22598 a_n2650_13878.n38 a_n2650_13878.n134 20.9683
R22599 a_n2650_13878.n133 a_n2650_13878.n73 48.2005
R22600 a_n2650_13878.n93 a_n2650_13878.n92 48.2005
R22601 a_n2650_13878.n95 a_n2650_13878.n58 20.9683
R22602 a_n2650_13878.n97 a_n2650_13878.n96 48.2005
R22603 a_n2650_13878.t31 a_n2650_13878.n62 533.335
R22604 a_n2650_13878.n86 a_n2650_13878.n85 48.2005
R22605 a_n2650_13878.n88 a_n2650_13878.n51 20.9683
R22606 a_n2650_13878.n90 a_n2650_13878.n89 48.2005
R22607 a_n2650_13878.t67 a_n2650_13878.n55 533.335
R22608 a_n2650_13878.n116 a_n2650_13878.n43 21.4216
R22609 a_n2650_13878.n135 a_n2650_13878.n37 21.4216
R22610 a_n2650_13878.n94 a_n2650_13878.n57 21.4216
R22611 a_n2650_13878.n87 a_n2650_13878.n50 21.4216
R22612 a_n2650_13878.n1 a_n2650_13878.n0 32.6799
R22613 a_n2650_13878.n47 a_n2650_13878.n76 34.4824
R22614 a_n2650_13878.n71 a_n2650_13878.n119 34.4824
R22615 a_n2650_13878.n98 a_n2650_13878.n61 34.4824
R22616 a_n2650_13878.n91 a_n2650_13878.n54 34.4824
R22617 a_n2650_13878.n111 a_n2650_13878.n69 35.3134
R22618 a_n2650_13878.n109 a_n2650_13878.n67 35.3134
R22619 a_n2650_13878.n107 a_n2650_13878.n65 35.3134
R22620 a_n2650_13878.n105 a_n2650_13878.n63 35.3134
R22621 a_n2650_13878.n115 a_n2650_13878.n45 35.3134
R22622 a_n2650_13878.n45 a_n2650_13878.n75 11.2134
R22623 a_n2650_13878.n134 a_n2650_13878.n39 35.3134
R22624 a_n2650_13878.n39 a_n2650_13878.n73 11.2134
R22625 a_n2650_13878.n95 a_n2650_13878.n59 35.3134
R22626 a_n2650_13878.n96 a_n2650_13878.n59 11.2134
R22627 a_n2650_13878.n88 a_n2650_13878.n52 35.3134
R22628 a_n2650_13878.n89 a_n2650_13878.n52 11.2134
R22629 a_n2650_13878.n27 a_n2650_13878.n2 23.891
R22630 a_n2650_13878.n42 a_n2650_13878.n74 36.139
R22631 a_n2650_13878.n36 a_n2650_13878.n72 36.139
R22632 a_n2650_13878.n82 a_n2650_13878.n56 36.139
R22633 a_n2650_13878.n84 a_n2650_13878.n49 36.139
R22634 a_n2650_13878.n21 a_n2650_13878.n11 13.3641
R22635 a_n2650_13878.n23 a_n2650_13878.n112 13.1596
R22636 a_n2650_13878.n138 a_n2650_13878.n28 11.8547
R22637 a_n2650_13878.n99 a_n2650_13878.n31 10.2167
R22638 a_n2650_13878.n112 a_n2650_13878.n5 9.99103
R22639 a_n2650_13878.n13 a_n2650_13878.n11 9.99103
R22640 a_n2650_13878.n99 a_n2650_13878.n15 8.01944
R22641 a_n2650_13878.n32 a_n2650_13878.n138 6.37334
R22642 a_n2650_13878.n112 a_n2650_13878.n99 5.3452
R22643 a_n2650_13878.n35 a_n2650_13878.n25 4.07247
R22644 a_n2650_13878.n17 a_n2650_13878.n19 4.07247
R22645 a_n2650_13878.n141 a_n2650_13878.t38 3.61217
R22646 a_n2650_13878.n141 a_n2650_13878.t34 3.61217
R22647 a_n2650_13878.n140 a_n2650_13878.t28 3.61217
R22648 a_n2650_13878.n140 a_n2650_13878.t14 3.61217
R22649 a_n2650_13878.n139 a_n2650_13878.t8 3.61217
R22650 a_n2650_13878.n139 a_n2650_13878.t26 3.61217
R22651 a_n2650_13878.n80 a_n2650_13878.t16 3.61217
R22652 a_n2650_13878.n80 a_n2650_13878.t40 3.61217
R22653 a_n2650_13878.n79 a_n2650_13878.t6 3.61217
R22654 a_n2650_13878.n79 a_n2650_13878.t22 3.61217
R22655 a_n2650_13878.n78 a_n2650_13878.t24 3.61217
R22656 a_n2650_13878.n78 a_n2650_13878.t42 3.61217
R22657 a_n2650_13878.n77 a_n2650_13878.t12 3.61217
R22658 a_n2650_13878.n77 a_n2650_13878.t20 3.61217
R22659 a_n2650_13878.t4 a_n2650_13878.n142 3.61217
R22660 a_n2650_13878.n142 a_n2650_13878.t10 3.61217
R22661 a_n2650_13878.n129 a_n2650_13878.t53 2.82907
R22662 a_n2650_13878.n129 a_n2650_13878.t54 2.82907
R22663 a_n2650_13878.n130 a_n2650_13878.t43 2.82907
R22664 a_n2650_13878.n130 a_n2650_13878.t63 2.82907
R22665 a_n2650_13878.n131 a_n2650_13878.t61 2.82907
R22666 a_n2650_13878.n131 a_n2650_13878.t46 2.82907
R22667 a_n2650_13878.n128 a_n2650_13878.t48 2.82907
R22668 a_n2650_13878.n128 a_n2650_13878.t52 2.82907
R22669 a_n2650_13878.n127 a_n2650_13878.t2 2.82907
R22670 a_n2650_13878.n127 a_n2650_13878.t0 2.82907
R22671 a_n2650_13878.n126 a_n2650_13878.t44 2.82907
R22672 a_n2650_13878.n126 a_n2650_13878.t50 2.82907
R22673 a_n2650_13878.n123 a_n2650_13878.t59 2.82907
R22674 a_n2650_13878.n123 a_n2650_13878.t62 2.82907
R22675 a_n2650_13878.n124 a_n2650_13878.t58 2.82907
R22676 a_n2650_13878.n124 a_n2650_13878.t45 2.82907
R22677 a_n2650_13878.n125 a_n2650_13878.t51 2.82907
R22678 a_n2650_13878.n125 a_n2650_13878.t55 2.82907
R22679 a_n2650_13878.n122 a_n2650_13878.t49 2.82907
R22680 a_n2650_13878.n122 a_n2650_13878.t56 2.82907
R22681 a_n2650_13878.n121 a_n2650_13878.t57 2.82907
R22682 a_n2650_13878.n121 a_n2650_13878.t60 2.82907
R22683 a_n2650_13878.n120 a_n2650_13878.t47 2.82907
R22684 a_n2650_13878.n120 a_n2650_13878.t1 2.82907
R22685 a_n2650_13878.n138 a_n2650_13878.n11 1.30542
R22686 a_n2650_13878.n8 a_n2650_13878.n9 1.04595
R22687 a_n2650_13878.n46 a_n2650_13878.n113 47.835
R22688 a_n2650_13878.n40 a_n2650_13878.n132 47.835
R22689 a_n2650_13878.n81 a_n2650_13878.n60 47.835
R22690 a_n2650_13878.n83 a_n2650_13878.n53 47.835
R22691 a_n2650_13878.n0 a_n2650_13878.n4 1.3324
R22692 a_n2650_13878.n23 a_n2650_13878.n22 1.13686
R22693 a_n2650_13878.n19 a_n2650_13878.n18 1.13686
R22694 a_n2650_13878.n15 a_n2650_13878.n14 1.13686
R22695 a_n2650_13878.n27 a_n2650_13878.n35 1.09898
R22696 a_n2650_13878.n2 a_n2650_13878.n3 0.888431
R22697 a_n2650_13878.n2 a_n2650_13878.n1 0.888431
R22698 a_n2650_13878.n28 a_n2650_13878.n26 0.758076
R22699 a_n2650_13878.n27 a_n2650_13878.n26 0.758076
R22700 a_n2650_13878.n25 a_n2650_13878.n24 0.758076
R22701 a_n2650_13878.n22 a_n2650_13878.n24 0.758076
R22702 a_n2650_13878.n20 a_n2650_13878.n21 0.758076
R22703 a_n2650_13878.n18 a_n2650_13878.n20 0.758076
R22704 a_n2650_13878.n16 a_n2650_13878.n17 0.758076
R22705 a_n2650_13878.n14 a_n2650_13878.n16 0.758076
R22706 a_n2650_13878.n13 a_n2650_13878.n12 0.758076
R22707 a_n2650_13878.n10 a_n2650_13878.n9 0.758076
R22708 a_n2650_13878.n8 a_n2650_13878.n7 0.758076
R22709 a_n2650_13878.n6 a_n2650_13878.n5 0.758076
R22710 a_n2650_13878.n34 a_n2650_13878.n33 0.716017
R22711 a_n2650_13878.n33 a_n2650_13878.n32 0.716017
R22712 a_n2650_13878.n31 a_n2650_13878.n30 0.716017
R22713 a_n2650_13878.n30 a_n2650_13878.n29 0.716017
R22714 a_n2650_13878.n10 a_n2650_13878.n12 0.67853
R22715 a_n2650_13878.n6 a_n2650_13878.n7 0.67853
R22716 a_n2472_13878.n2 a_n2472_13878.n0 98.9633
R22717 a_n2472_13878.n5 a_n2472_13878.n3 98.7517
R22718 a_n2472_13878.n23 a_n2472_13878.n22 98.6055
R22719 a_n2472_13878.n2 a_n2472_13878.n1 98.6055
R22720 a_n2472_13878.n11 a_n2472_13878.n10 98.6055
R22721 a_n2472_13878.n9 a_n2472_13878.n8 98.6055
R22722 a_n2472_13878.n7 a_n2472_13878.n6 98.6055
R22723 a_n2472_13878.n5 a_n2472_13878.n4 98.6055
R22724 a_n2472_13878.n25 a_n2472_13878.n24 98.6054
R22725 a_n2472_13878.n21 a_n2472_13878.n20 98.6054
R22726 a_n2472_13878.n13 a_n2472_13878.t1 74.6477
R22727 a_n2472_13878.n18 a_n2472_13878.t2 74.2899
R22728 a_n2472_13878.n15 a_n2472_13878.t3 74.2899
R22729 a_n2472_13878.n14 a_n2472_13878.t0 74.2899
R22730 a_n2472_13878.n17 a_n2472_13878.n16 70.6783
R22731 a_n2472_13878.n13 a_n2472_13878.n12 70.6783
R22732 a_n2472_13878.n19 a_n2472_13878.n11 15.0004
R22733 a_n2472_13878.n21 a_n2472_13878.n19 12.2917
R22734 a_n2472_13878.n19 a_n2472_13878.n18 7.67184
R22735 a_n2472_13878.n20 a_n2472_13878.t24 3.61217
R22736 a_n2472_13878.n20 a_n2472_13878.t13 3.61217
R22737 a_n2472_13878.n22 a_n2472_13878.t16 3.61217
R22738 a_n2472_13878.n22 a_n2472_13878.t17 3.61217
R22739 a_n2472_13878.n1 a_n2472_13878.t8 3.61217
R22740 a_n2472_13878.n1 a_n2472_13878.t18 3.61217
R22741 a_n2472_13878.n0 a_n2472_13878.t21 3.61217
R22742 a_n2472_13878.n0 a_n2472_13878.t27 3.61217
R22743 a_n2472_13878.n16 a_n2472_13878.t6 3.61217
R22744 a_n2472_13878.n16 a_n2472_13878.t7 3.61217
R22745 a_n2472_13878.n12 a_n2472_13878.t4 3.61217
R22746 a_n2472_13878.n12 a_n2472_13878.t5 3.61217
R22747 a_n2472_13878.n10 a_n2472_13878.t19 3.61217
R22748 a_n2472_13878.n10 a_n2472_13878.t9 3.61217
R22749 a_n2472_13878.n8 a_n2472_13878.t22 3.61217
R22750 a_n2472_13878.n8 a_n2472_13878.t11 3.61217
R22751 a_n2472_13878.n6 a_n2472_13878.t10 3.61217
R22752 a_n2472_13878.n6 a_n2472_13878.t12 3.61217
R22753 a_n2472_13878.n4 a_n2472_13878.t20 3.61217
R22754 a_n2472_13878.n4 a_n2472_13878.t14 3.61217
R22755 a_n2472_13878.n3 a_n2472_13878.t23 3.61217
R22756 a_n2472_13878.n3 a_n2472_13878.t15 3.61217
R22757 a_n2472_13878.n25 a_n2472_13878.t25 3.61217
R22758 a_n2472_13878.t26 a_n2472_13878.n25 3.61217
R22759 a_n2472_13878.n14 a_n2472_13878.n13 0.358259
R22760 a_n2472_13878.n17 a_n2472_13878.n15 0.358259
R22761 a_n2472_13878.n18 a_n2472_13878.n17 0.358259
R22762 a_n2472_13878.n24 a_n2472_13878.n2 0.358259
R22763 a_n2472_13878.n24 a_n2472_13878.n23 0.358259
R22764 a_n2472_13878.n23 a_n2472_13878.n21 0.358259
R22765 a_n2472_13878.n7 a_n2472_13878.n5 0.146627
R22766 a_n2472_13878.n9 a_n2472_13878.n7 0.146627
R22767 a_n2472_13878.n11 a_n2472_13878.n9 0.146627
R22768 a_n2472_13878.n15 a_n2472_13878.n14 0.101793
R22769 outputibias.n27 outputibias.n1 289.615
R22770 outputibias.n58 outputibias.n32 289.615
R22771 outputibias.n90 outputibias.n64 289.615
R22772 outputibias.n122 outputibias.n96 289.615
R22773 outputibias.n28 outputibias.n27 185
R22774 outputibias.n26 outputibias.n25 185
R22775 outputibias.n5 outputibias.n4 185
R22776 outputibias.n20 outputibias.n19 185
R22777 outputibias.n18 outputibias.n17 185
R22778 outputibias.n9 outputibias.n8 185
R22779 outputibias.n12 outputibias.n11 185
R22780 outputibias.n59 outputibias.n58 185
R22781 outputibias.n57 outputibias.n56 185
R22782 outputibias.n36 outputibias.n35 185
R22783 outputibias.n51 outputibias.n50 185
R22784 outputibias.n49 outputibias.n48 185
R22785 outputibias.n40 outputibias.n39 185
R22786 outputibias.n43 outputibias.n42 185
R22787 outputibias.n91 outputibias.n90 185
R22788 outputibias.n89 outputibias.n88 185
R22789 outputibias.n68 outputibias.n67 185
R22790 outputibias.n83 outputibias.n82 185
R22791 outputibias.n81 outputibias.n80 185
R22792 outputibias.n72 outputibias.n71 185
R22793 outputibias.n75 outputibias.n74 185
R22794 outputibias.n123 outputibias.n122 185
R22795 outputibias.n121 outputibias.n120 185
R22796 outputibias.n100 outputibias.n99 185
R22797 outputibias.n115 outputibias.n114 185
R22798 outputibias.n113 outputibias.n112 185
R22799 outputibias.n104 outputibias.n103 185
R22800 outputibias.n107 outputibias.n106 185
R22801 outputibias.n0 outputibias.t8 178.945
R22802 outputibias.n133 outputibias.t9 177.018
R22803 outputibias.n132 outputibias.t11 177.018
R22804 outputibias.n0 outputibias.t10 177.018
R22805 outputibias.t5 outputibias.n10 147.661
R22806 outputibias.t3 outputibias.n41 147.661
R22807 outputibias.t1 outputibias.n73 147.661
R22808 outputibias.t7 outputibias.n105 147.661
R22809 outputibias.n128 outputibias.t4 132.363
R22810 outputibias.n128 outputibias.t2 130.436
R22811 outputibias.n129 outputibias.t0 130.436
R22812 outputibias.n130 outputibias.t6 130.436
R22813 outputibias.n27 outputibias.n26 104.615
R22814 outputibias.n26 outputibias.n4 104.615
R22815 outputibias.n19 outputibias.n4 104.615
R22816 outputibias.n19 outputibias.n18 104.615
R22817 outputibias.n18 outputibias.n8 104.615
R22818 outputibias.n11 outputibias.n8 104.615
R22819 outputibias.n58 outputibias.n57 104.615
R22820 outputibias.n57 outputibias.n35 104.615
R22821 outputibias.n50 outputibias.n35 104.615
R22822 outputibias.n50 outputibias.n49 104.615
R22823 outputibias.n49 outputibias.n39 104.615
R22824 outputibias.n42 outputibias.n39 104.615
R22825 outputibias.n90 outputibias.n89 104.615
R22826 outputibias.n89 outputibias.n67 104.615
R22827 outputibias.n82 outputibias.n67 104.615
R22828 outputibias.n82 outputibias.n81 104.615
R22829 outputibias.n81 outputibias.n71 104.615
R22830 outputibias.n74 outputibias.n71 104.615
R22831 outputibias.n122 outputibias.n121 104.615
R22832 outputibias.n121 outputibias.n99 104.615
R22833 outputibias.n114 outputibias.n99 104.615
R22834 outputibias.n114 outputibias.n113 104.615
R22835 outputibias.n113 outputibias.n103 104.615
R22836 outputibias.n106 outputibias.n103 104.615
R22837 outputibias.n63 outputibias.n31 95.6354
R22838 outputibias.n63 outputibias.n62 94.6732
R22839 outputibias.n95 outputibias.n94 94.6732
R22840 outputibias.n127 outputibias.n126 94.6732
R22841 outputibias.n11 outputibias.t5 52.3082
R22842 outputibias.n42 outputibias.t3 52.3082
R22843 outputibias.n74 outputibias.t1 52.3082
R22844 outputibias.n106 outputibias.t7 52.3082
R22845 outputibias.n12 outputibias.n10 15.6674
R22846 outputibias.n43 outputibias.n41 15.6674
R22847 outputibias.n75 outputibias.n73 15.6674
R22848 outputibias.n107 outputibias.n105 15.6674
R22849 outputibias.n13 outputibias.n9 12.8005
R22850 outputibias.n44 outputibias.n40 12.8005
R22851 outputibias.n76 outputibias.n72 12.8005
R22852 outputibias.n108 outputibias.n104 12.8005
R22853 outputibias.n17 outputibias.n16 12.0247
R22854 outputibias.n48 outputibias.n47 12.0247
R22855 outputibias.n80 outputibias.n79 12.0247
R22856 outputibias.n112 outputibias.n111 12.0247
R22857 outputibias.n20 outputibias.n7 11.249
R22858 outputibias.n51 outputibias.n38 11.249
R22859 outputibias.n83 outputibias.n70 11.249
R22860 outputibias.n115 outputibias.n102 11.249
R22861 outputibias.n21 outputibias.n5 10.4732
R22862 outputibias.n52 outputibias.n36 10.4732
R22863 outputibias.n84 outputibias.n68 10.4732
R22864 outputibias.n116 outputibias.n100 10.4732
R22865 outputibias.n25 outputibias.n24 9.69747
R22866 outputibias.n56 outputibias.n55 9.69747
R22867 outputibias.n88 outputibias.n87 9.69747
R22868 outputibias.n120 outputibias.n119 9.69747
R22869 outputibias.n31 outputibias.n30 9.45567
R22870 outputibias.n62 outputibias.n61 9.45567
R22871 outputibias.n94 outputibias.n93 9.45567
R22872 outputibias.n126 outputibias.n125 9.45567
R22873 outputibias.n30 outputibias.n29 9.3005
R22874 outputibias.n3 outputibias.n2 9.3005
R22875 outputibias.n24 outputibias.n23 9.3005
R22876 outputibias.n22 outputibias.n21 9.3005
R22877 outputibias.n7 outputibias.n6 9.3005
R22878 outputibias.n16 outputibias.n15 9.3005
R22879 outputibias.n14 outputibias.n13 9.3005
R22880 outputibias.n61 outputibias.n60 9.3005
R22881 outputibias.n34 outputibias.n33 9.3005
R22882 outputibias.n55 outputibias.n54 9.3005
R22883 outputibias.n53 outputibias.n52 9.3005
R22884 outputibias.n38 outputibias.n37 9.3005
R22885 outputibias.n47 outputibias.n46 9.3005
R22886 outputibias.n45 outputibias.n44 9.3005
R22887 outputibias.n93 outputibias.n92 9.3005
R22888 outputibias.n66 outputibias.n65 9.3005
R22889 outputibias.n87 outputibias.n86 9.3005
R22890 outputibias.n85 outputibias.n84 9.3005
R22891 outputibias.n70 outputibias.n69 9.3005
R22892 outputibias.n79 outputibias.n78 9.3005
R22893 outputibias.n77 outputibias.n76 9.3005
R22894 outputibias.n125 outputibias.n124 9.3005
R22895 outputibias.n98 outputibias.n97 9.3005
R22896 outputibias.n119 outputibias.n118 9.3005
R22897 outputibias.n117 outputibias.n116 9.3005
R22898 outputibias.n102 outputibias.n101 9.3005
R22899 outputibias.n111 outputibias.n110 9.3005
R22900 outputibias.n109 outputibias.n108 9.3005
R22901 outputibias.n28 outputibias.n3 8.92171
R22902 outputibias.n59 outputibias.n34 8.92171
R22903 outputibias.n91 outputibias.n66 8.92171
R22904 outputibias.n123 outputibias.n98 8.92171
R22905 outputibias.n29 outputibias.n1 8.14595
R22906 outputibias.n60 outputibias.n32 8.14595
R22907 outputibias.n92 outputibias.n64 8.14595
R22908 outputibias.n124 outputibias.n96 8.14595
R22909 outputibias.n31 outputibias.n1 5.81868
R22910 outputibias.n62 outputibias.n32 5.81868
R22911 outputibias.n94 outputibias.n64 5.81868
R22912 outputibias.n126 outputibias.n96 5.81868
R22913 outputibias.n131 outputibias.n130 5.20947
R22914 outputibias.n29 outputibias.n28 5.04292
R22915 outputibias.n60 outputibias.n59 5.04292
R22916 outputibias.n92 outputibias.n91 5.04292
R22917 outputibias.n124 outputibias.n123 5.04292
R22918 outputibias.n131 outputibias.n127 4.42209
R22919 outputibias.n14 outputibias.n10 4.38594
R22920 outputibias.n45 outputibias.n41 4.38594
R22921 outputibias.n77 outputibias.n73 4.38594
R22922 outputibias.n109 outputibias.n105 4.38594
R22923 outputibias.n132 outputibias.n131 4.28454
R22924 outputibias.n25 outputibias.n3 4.26717
R22925 outputibias.n56 outputibias.n34 4.26717
R22926 outputibias.n88 outputibias.n66 4.26717
R22927 outputibias.n120 outputibias.n98 4.26717
R22928 outputibias.n24 outputibias.n5 3.49141
R22929 outputibias.n55 outputibias.n36 3.49141
R22930 outputibias.n87 outputibias.n68 3.49141
R22931 outputibias.n119 outputibias.n100 3.49141
R22932 outputibias.n21 outputibias.n20 2.71565
R22933 outputibias.n52 outputibias.n51 2.71565
R22934 outputibias.n84 outputibias.n83 2.71565
R22935 outputibias.n116 outputibias.n115 2.71565
R22936 outputibias.n17 outputibias.n7 1.93989
R22937 outputibias.n48 outputibias.n38 1.93989
R22938 outputibias.n80 outputibias.n70 1.93989
R22939 outputibias.n112 outputibias.n102 1.93989
R22940 outputibias.n130 outputibias.n129 1.9266
R22941 outputibias.n129 outputibias.n128 1.9266
R22942 outputibias.n133 outputibias.n132 1.92658
R22943 outputibias.n134 outputibias.n133 1.29913
R22944 outputibias.n16 outputibias.n9 1.16414
R22945 outputibias.n47 outputibias.n40 1.16414
R22946 outputibias.n79 outputibias.n72 1.16414
R22947 outputibias.n111 outputibias.n104 1.16414
R22948 outputibias.n127 outputibias.n95 0.962709
R22949 outputibias.n95 outputibias.n63 0.962709
R22950 outputibias.n13 outputibias.n12 0.388379
R22951 outputibias.n44 outputibias.n43 0.388379
R22952 outputibias.n76 outputibias.n75 0.388379
R22953 outputibias.n108 outputibias.n107 0.388379
R22954 outputibias.n134 outputibias.n0 0.337251
R22955 outputibias outputibias.n134 0.302375
R22956 outputibias.n30 outputibias.n2 0.155672
R22957 outputibias.n23 outputibias.n2 0.155672
R22958 outputibias.n23 outputibias.n22 0.155672
R22959 outputibias.n22 outputibias.n6 0.155672
R22960 outputibias.n15 outputibias.n6 0.155672
R22961 outputibias.n15 outputibias.n14 0.155672
R22962 outputibias.n61 outputibias.n33 0.155672
R22963 outputibias.n54 outputibias.n33 0.155672
R22964 outputibias.n54 outputibias.n53 0.155672
R22965 outputibias.n53 outputibias.n37 0.155672
R22966 outputibias.n46 outputibias.n37 0.155672
R22967 outputibias.n46 outputibias.n45 0.155672
R22968 outputibias.n93 outputibias.n65 0.155672
R22969 outputibias.n86 outputibias.n65 0.155672
R22970 outputibias.n86 outputibias.n85 0.155672
R22971 outputibias.n85 outputibias.n69 0.155672
R22972 outputibias.n78 outputibias.n69 0.155672
R22973 outputibias.n78 outputibias.n77 0.155672
R22974 outputibias.n125 outputibias.n97 0.155672
R22975 outputibias.n118 outputibias.n97 0.155672
R22976 outputibias.n118 outputibias.n117 0.155672
R22977 outputibias.n117 outputibias.n101 0.155672
R22978 outputibias.n110 outputibias.n101 0.155672
R22979 outputibias.n110 outputibias.n109 0.155672
R22980 minus.n53 minus.t28 323.478
R22981 minus.n11 minus.t8 323.478
R22982 minus.n82 minus.t13 297.12
R22983 minus.n80 minus.t15 297.12
R22984 minus.n44 minus.t5 297.12
R22985 minus.n74 minus.t6 297.12
R22986 minus.n46 minus.t26 297.12
R22987 minus.n68 minus.t21 297.12
R22988 minus.n48 minus.t23 297.12
R22989 minus.n62 minus.t16 297.12
R22990 minus.n50 minus.t17 297.12
R22991 minus.n56 minus.t9 297.12
R22992 minus.n52 minus.t27 297.12
R22993 minus.n10 minus.t7 297.12
R22994 minus.n14 minus.t11 297.12
R22995 minus.n16 minus.t10 297.12
R22996 minus.n20 minus.t12 297.12
R22997 minus.n22 minus.t20 297.12
R22998 minus.n26 minus.t18 297.12
R22999 minus.n28 minus.t25 297.12
R23000 minus.n32 minus.t24 297.12
R23001 minus.n34 minus.t14 297.12
R23002 minus.n38 minus.t22 297.12
R23003 minus.n40 minus.t19 297.12
R23004 minus.n88 minus.t2 243.255
R23005 minus.n87 minus.n85 224.169
R23006 minus.n87 minus.n86 223.454
R23007 minus.n55 minus.n54 161.3
R23008 minus.n56 minus.n51 161.3
R23009 minus.n58 minus.n57 161.3
R23010 minus.n59 minus.n50 161.3
R23011 minus.n61 minus.n60 161.3
R23012 minus.n62 minus.n49 161.3
R23013 minus.n64 minus.n63 161.3
R23014 minus.n65 minus.n48 161.3
R23015 minus.n67 minus.n66 161.3
R23016 minus.n68 minus.n47 161.3
R23017 minus.n70 minus.n69 161.3
R23018 minus.n71 minus.n46 161.3
R23019 minus.n73 minus.n72 161.3
R23020 minus.n74 minus.n45 161.3
R23021 minus.n76 minus.n75 161.3
R23022 minus.n77 minus.n44 161.3
R23023 minus.n79 minus.n78 161.3
R23024 minus.n80 minus.n43 161.3
R23025 minus.n81 minus.n42 161.3
R23026 minus.n83 minus.n82 161.3
R23027 minus.n41 minus.n40 161.3
R23028 minus.n39 minus.n0 161.3
R23029 minus.n38 minus.n37 161.3
R23030 minus.n36 minus.n1 161.3
R23031 minus.n35 minus.n34 161.3
R23032 minus.n33 minus.n2 161.3
R23033 minus.n32 minus.n31 161.3
R23034 minus.n30 minus.n3 161.3
R23035 minus.n29 minus.n28 161.3
R23036 minus.n27 minus.n4 161.3
R23037 minus.n26 minus.n25 161.3
R23038 minus.n24 minus.n5 161.3
R23039 minus.n23 minus.n22 161.3
R23040 minus.n21 minus.n6 161.3
R23041 minus.n20 minus.n19 161.3
R23042 minus.n18 minus.n7 161.3
R23043 minus.n17 minus.n16 161.3
R23044 minus.n15 minus.n8 161.3
R23045 minus.n14 minus.n13 161.3
R23046 minus.n12 minus.n9 161.3
R23047 minus.n82 minus.n81 46.0096
R23048 minus.n40 minus.n39 46.0096
R23049 minus.n12 minus.n11 45.0871
R23050 minus.n54 minus.n53 45.0871
R23051 minus.n80 minus.n79 41.6278
R23052 minus.n55 minus.n52 41.6278
R23053 minus.n10 minus.n9 41.6278
R23054 minus.n38 minus.n1 41.6278
R23055 minus.n75 minus.n44 37.246
R23056 minus.n57 minus.n56 37.246
R23057 minus.n15 minus.n14 37.246
R23058 minus.n34 minus.n33 37.246
R23059 minus.n84 minus.n83 33.3925
R23060 minus.n74 minus.n73 32.8641
R23061 minus.n61 minus.n50 32.8641
R23062 minus.n16 minus.n7 32.8641
R23063 minus.n32 minus.n3 32.8641
R23064 minus.n69 minus.n46 28.4823
R23065 minus.n63 minus.n62 28.4823
R23066 minus.n21 minus.n20 28.4823
R23067 minus.n28 minus.n27 28.4823
R23068 minus.n68 minus.n67 24.1005
R23069 minus.n67 minus.n48 24.1005
R23070 minus.n22 minus.n5 24.1005
R23071 minus.n26 minus.n5 24.1005
R23072 minus.n86 minus.t4 19.8005
R23073 minus.n86 minus.t3 19.8005
R23074 minus.n85 minus.t1 19.8005
R23075 minus.n85 minus.t0 19.8005
R23076 minus.n69 minus.n68 19.7187
R23077 minus.n63 minus.n48 19.7187
R23078 minus.n22 minus.n21 19.7187
R23079 minus.n27 minus.n26 19.7187
R23080 minus.n73 minus.n46 15.3369
R23081 minus.n62 minus.n61 15.3369
R23082 minus.n20 minus.n7 15.3369
R23083 minus.n28 minus.n3 15.3369
R23084 minus.n53 minus.n52 14.1472
R23085 minus.n11 minus.n10 14.1472
R23086 minus.n84 minus.n41 12.0933
R23087 minus minus.n89 12.0331
R23088 minus.n75 minus.n74 10.955
R23089 minus.n57 minus.n50 10.955
R23090 minus.n16 minus.n15 10.955
R23091 minus.n33 minus.n32 10.955
R23092 minus.n79 minus.n44 6.57323
R23093 minus.n56 minus.n55 6.57323
R23094 minus.n14 minus.n9 6.57323
R23095 minus.n34 minus.n1 6.57323
R23096 minus.n89 minus.n88 4.80222
R23097 minus.n81 minus.n80 2.19141
R23098 minus.n39 minus.n38 2.19141
R23099 minus.n89 minus.n84 0.972091
R23100 minus.n88 minus.n87 0.716017
R23101 minus.n83 minus.n42 0.189894
R23102 minus.n43 minus.n42 0.189894
R23103 minus.n78 minus.n43 0.189894
R23104 minus.n78 minus.n77 0.189894
R23105 minus.n77 minus.n76 0.189894
R23106 minus.n76 minus.n45 0.189894
R23107 minus.n72 minus.n45 0.189894
R23108 minus.n72 minus.n71 0.189894
R23109 minus.n71 minus.n70 0.189894
R23110 minus.n70 minus.n47 0.189894
R23111 minus.n66 minus.n47 0.189894
R23112 minus.n66 minus.n65 0.189894
R23113 minus.n65 minus.n64 0.189894
R23114 minus.n64 minus.n49 0.189894
R23115 minus.n60 minus.n49 0.189894
R23116 minus.n60 minus.n59 0.189894
R23117 minus.n59 minus.n58 0.189894
R23118 minus.n58 minus.n51 0.189894
R23119 minus.n54 minus.n51 0.189894
R23120 minus.n13 minus.n12 0.189894
R23121 minus.n13 minus.n8 0.189894
R23122 minus.n17 minus.n8 0.189894
R23123 minus.n18 minus.n17 0.189894
R23124 minus.n19 minus.n18 0.189894
R23125 minus.n19 minus.n6 0.189894
R23126 minus.n23 minus.n6 0.189894
R23127 minus.n24 minus.n23 0.189894
R23128 minus.n25 minus.n24 0.189894
R23129 minus.n25 minus.n4 0.189894
R23130 minus.n29 minus.n4 0.189894
R23131 minus.n30 minus.n29 0.189894
R23132 minus.n31 minus.n30 0.189894
R23133 minus.n31 minus.n2 0.189894
R23134 minus.n35 minus.n2 0.189894
R23135 minus.n36 minus.n35 0.189894
R23136 minus.n37 minus.n36 0.189894
R23137 minus.n37 minus.n0 0.189894
R23138 minus.n41 minus.n0 0.189894
R23139 diffpairibias.n0 diffpairibias.t27 436.822
R23140 diffpairibias.n27 diffpairibias.t24 435.479
R23141 diffpairibias.n26 diffpairibias.t21 435.479
R23142 diffpairibias.n25 diffpairibias.t22 435.479
R23143 diffpairibias.n24 diffpairibias.t26 435.479
R23144 diffpairibias.n23 diffpairibias.t20 435.479
R23145 diffpairibias.n0 diffpairibias.t23 435.479
R23146 diffpairibias.n1 diffpairibias.t28 435.479
R23147 diffpairibias.n2 diffpairibias.t25 435.479
R23148 diffpairibias.n3 diffpairibias.t29 435.479
R23149 diffpairibias.n13 diffpairibias.t14 377.536
R23150 diffpairibias.n13 diffpairibias.t0 376.193
R23151 diffpairibias.n14 diffpairibias.t10 376.193
R23152 diffpairibias.n15 diffpairibias.t12 376.193
R23153 diffpairibias.n16 diffpairibias.t6 376.193
R23154 diffpairibias.n17 diffpairibias.t2 376.193
R23155 diffpairibias.n18 diffpairibias.t16 376.193
R23156 diffpairibias.n19 diffpairibias.t4 376.193
R23157 diffpairibias.n20 diffpairibias.t18 376.193
R23158 diffpairibias.n21 diffpairibias.t8 376.193
R23159 diffpairibias.n4 diffpairibias.t15 113.368
R23160 diffpairibias.n4 diffpairibias.t1 112.698
R23161 diffpairibias.n5 diffpairibias.t11 112.698
R23162 diffpairibias.n6 diffpairibias.t13 112.698
R23163 diffpairibias.n7 diffpairibias.t7 112.698
R23164 diffpairibias.n8 diffpairibias.t3 112.698
R23165 diffpairibias.n9 diffpairibias.t17 112.698
R23166 diffpairibias.n10 diffpairibias.t5 112.698
R23167 diffpairibias.n11 diffpairibias.t19 112.698
R23168 diffpairibias.n12 diffpairibias.t9 112.698
R23169 diffpairibias.n22 diffpairibias.n21 4.77242
R23170 diffpairibias.n22 diffpairibias.n12 4.30807
R23171 diffpairibias.n23 diffpairibias.n22 4.13945
R23172 diffpairibias.n21 diffpairibias.n20 1.34352
R23173 diffpairibias.n20 diffpairibias.n19 1.34352
R23174 diffpairibias.n19 diffpairibias.n18 1.34352
R23175 diffpairibias.n18 diffpairibias.n17 1.34352
R23176 diffpairibias.n17 diffpairibias.n16 1.34352
R23177 diffpairibias.n16 diffpairibias.n15 1.34352
R23178 diffpairibias.n15 diffpairibias.n14 1.34352
R23179 diffpairibias.n14 diffpairibias.n13 1.34352
R23180 diffpairibias.n3 diffpairibias.n2 1.34352
R23181 diffpairibias.n2 diffpairibias.n1 1.34352
R23182 diffpairibias.n1 diffpairibias.n0 1.34352
R23183 diffpairibias.n24 diffpairibias.n23 1.34352
R23184 diffpairibias.n25 diffpairibias.n24 1.34352
R23185 diffpairibias.n26 diffpairibias.n25 1.34352
R23186 diffpairibias.n27 diffpairibias.n26 1.34352
R23187 diffpairibias.n28 diffpairibias.n27 0.862419
R23188 diffpairibias diffpairibias.n28 0.684875
R23189 diffpairibias.n12 diffpairibias.n11 0.672012
R23190 diffpairibias.n11 diffpairibias.n10 0.672012
R23191 diffpairibias.n10 diffpairibias.n9 0.672012
R23192 diffpairibias.n9 diffpairibias.n8 0.672012
R23193 diffpairibias.n8 diffpairibias.n7 0.672012
R23194 diffpairibias.n7 diffpairibias.n6 0.672012
R23195 diffpairibias.n6 diffpairibias.n5 0.672012
R23196 diffpairibias.n5 diffpairibias.n4 0.672012
R23197 diffpairibias.n28 diffpairibias.n3 0.190907
R23198 commonsourceibias.n281 commonsourceibias.t101 222.032
R23199 commonsourceibias.n44 commonsourceibias.t78 222.032
R23200 commonsourceibias.n166 commonsourceibias.t117 222.032
R23201 commonsourceibias.n643 commonsourceibias.t106 222.032
R23202 commonsourceibias.n413 commonsourceibias.t28 222.032
R23203 commonsourceibias.n529 commonsourceibias.t123 222.032
R23204 commonsourceibias.n364 commonsourceibias.t100 207.983
R23205 commonsourceibias.n127 commonsourceibias.t74 207.983
R23206 commonsourceibias.n249 commonsourceibias.t115 207.983
R23207 commonsourceibias.n731 commonsourceibias.t122 207.983
R23208 commonsourceibias.n501 commonsourceibias.t14 207.983
R23209 commonsourceibias.n616 commonsourceibias.t140 207.983
R23210 commonsourceibias.n280 commonsourceibias.t87 168.701
R23211 commonsourceibias.n286 commonsourceibias.t129 168.701
R23212 commonsourceibias.n292 commonsourceibias.t110 168.701
R23213 commonsourceibias.n276 commonsourceibias.t93 168.701
R23214 commonsourceibias.n300 commonsourceibias.t95 168.701
R23215 commonsourceibias.n306 commonsourceibias.t121 168.701
R23216 commonsourceibias.n271 commonsourceibias.t102 168.701
R23217 commonsourceibias.n314 commonsourceibias.t108 168.701
R23218 commonsourceibias.n320 commonsourceibias.t159 168.701
R23219 commonsourceibias.n266 commonsourceibias.t138 168.701
R23220 commonsourceibias.n328 commonsourceibias.t118 168.701
R23221 commonsourceibias.n334 commonsourceibias.t83 168.701
R23222 commonsourceibias.n261 commonsourceibias.t86 168.701
R23223 commonsourceibias.n342 commonsourceibias.t128 168.701
R23224 commonsourceibias.n348 commonsourceibias.t109 168.701
R23225 commonsourceibias.n256 commonsourceibias.t92 168.701
R23226 commonsourceibias.n356 commonsourceibias.t137 168.701
R23227 commonsourceibias.n362 commonsourceibias.t119 168.701
R23228 commonsourceibias.n125 commonsourceibias.t20 168.701
R23229 commonsourceibias.n119 commonsourceibias.t50 168.701
R23230 commonsourceibias.n19 commonsourceibias.t8 168.701
R23231 commonsourceibias.n111 commonsourceibias.t36 168.701
R23232 commonsourceibias.n105 commonsourceibias.t76 168.701
R23233 commonsourceibias.n24 commonsourceibias.t24 168.701
R23234 commonsourceibias.n97 commonsourceibias.t34 168.701
R23235 commonsourceibias.n91 commonsourceibias.t10 168.701
R23236 commonsourceibias.n29 commonsourceibias.t40 168.701
R23237 commonsourceibias.n83 commonsourceibias.t56 168.701
R23238 commonsourceibias.n77 commonsourceibias.t26 168.701
R23239 commonsourceibias.n34 commonsourceibias.t38 168.701
R23240 commonsourceibias.n69 commonsourceibias.t70 168.701
R23241 commonsourceibias.n63 commonsourceibias.t18 168.701
R23242 commonsourceibias.n39 commonsourceibias.t22 168.701
R23243 commonsourceibias.n55 commonsourceibias.t54 168.701
R23244 commonsourceibias.n49 commonsourceibias.t4 168.701
R23245 commonsourceibias.n43 commonsourceibias.t46 168.701
R23246 commonsourceibias.n247 commonsourceibias.t136 168.701
R23247 commonsourceibias.n241 commonsourceibias.t151 168.701
R23248 commonsourceibias.n5 commonsourceibias.t105 168.701
R23249 commonsourceibias.n233 commonsourceibias.t126 168.701
R23250 commonsourceibias.n227 commonsourceibias.t144 168.701
R23251 commonsourceibias.n10 commonsourceibias.t98 168.701
R23252 commonsourceibias.n219 commonsourceibias.t94 168.701
R23253 commonsourceibias.n213 commonsourceibias.t135 168.701
R23254 commonsourceibias.n150 commonsourceibias.t153 168.701
R23255 commonsourceibias.n151 commonsourceibias.t88 168.701
R23256 commonsourceibias.n153 commonsourceibias.t125 168.701
R23257 commonsourceibias.n155 commonsourceibias.t120 168.701
R23258 commonsourceibias.n191 commonsourceibias.t139 168.701
R23259 commonsourceibias.n185 commonsourceibias.t112 168.701
R23260 commonsourceibias.n161 commonsourceibias.t107 168.701
R23261 commonsourceibias.n177 commonsourceibias.t127 168.701
R23262 commonsourceibias.n171 commonsourceibias.t146 168.701
R23263 commonsourceibias.n165 commonsourceibias.t99 168.701
R23264 commonsourceibias.n642 commonsourceibias.t90 168.701
R23265 commonsourceibias.n648 commonsourceibias.t134 168.701
R23266 commonsourceibias.n654 commonsourceibias.t116 168.701
R23267 commonsourceibias.n656 commonsourceibias.t96 168.701
R23268 commonsourceibias.n663 commonsourceibias.t91 168.701
R23269 commonsourceibias.n669 commonsourceibias.t145 168.701
R23270 commonsourceibias.n671 commonsourceibias.t124 168.701
R23271 commonsourceibias.n678 commonsourceibias.t131 168.701
R23272 commonsourceibias.n684 commonsourceibias.t152 168.701
R23273 commonsourceibias.n686 commonsourceibias.t157 168.701
R23274 commonsourceibias.n693 commonsourceibias.t141 168.701
R23275 commonsourceibias.n699 commonsourceibias.t97 168.701
R23276 commonsourceibias.n701 commonsourceibias.t81 168.701
R23277 commonsourceibias.n708 commonsourceibias.t149 168.701
R23278 commonsourceibias.n714 commonsourceibias.t132 168.701
R23279 commonsourceibias.n716 commonsourceibias.t111 168.701
R23280 commonsourceibias.n723 commonsourceibias.t156 168.701
R23281 commonsourceibias.n729 commonsourceibias.t142 168.701
R23282 commonsourceibias.n412 commonsourceibias.t2 168.701
R23283 commonsourceibias.n418 commonsourceibias.t48 168.701
R23284 commonsourceibias.n424 commonsourceibias.t12 168.701
R23285 commonsourceibias.n426 commonsourceibias.t68 168.701
R23286 commonsourceibias.n433 commonsourceibias.t66 168.701
R23287 commonsourceibias.n439 commonsourceibias.t6 168.701
R23288 commonsourceibias.n441 commonsourceibias.t62 168.701
R23289 commonsourceibias.n448 commonsourceibias.t52 168.701
R23290 commonsourceibias.n454 commonsourceibias.t72 168.701
R23291 commonsourceibias.n456 commonsourceibias.t64 168.701
R23292 commonsourceibias.n463 commonsourceibias.t32 168.701
R23293 commonsourceibias.n469 commonsourceibias.t58 168.701
R23294 commonsourceibias.n471 commonsourceibias.t44 168.701
R23295 commonsourceibias.n478 commonsourceibias.t16 168.701
R23296 commonsourceibias.n484 commonsourceibias.t60 168.701
R23297 commonsourceibias.n486 commonsourceibias.t30 168.701
R23298 commonsourceibias.n493 commonsourceibias.t0 168.701
R23299 commonsourceibias.n499 commonsourceibias.t42 168.701
R23300 commonsourceibias.n614 commonsourceibias.t155 168.701
R23301 commonsourceibias.n608 commonsourceibias.t84 168.701
R23302 commonsourceibias.n601 commonsourceibias.t130 168.701
R23303 commonsourceibias.n599 commonsourceibias.t148 168.701
R23304 commonsourceibias.n593 commonsourceibias.t80 168.701
R23305 commonsourceibias.n586 commonsourceibias.t89 168.701
R23306 commonsourceibias.n584 commonsourceibias.t113 168.701
R23307 commonsourceibias.n578 commonsourceibias.t154 168.701
R23308 commonsourceibias.n571 commonsourceibias.t85 168.701
R23309 commonsourceibias.n528 commonsourceibias.t103 168.701
R23310 commonsourceibias.n534 commonsourceibias.t150 168.701
R23311 commonsourceibias.n540 commonsourceibias.t133 168.701
R23312 commonsourceibias.n542 commonsourceibias.t114 168.701
R23313 commonsourceibias.n549 commonsourceibias.t104 168.701
R23314 commonsourceibias.n555 commonsourceibias.t158 168.701
R23315 commonsourceibias.n519 commonsourceibias.t143 168.701
R23316 commonsourceibias.n517 commonsourceibias.t147 168.701
R23317 commonsourceibias.n515 commonsourceibias.t82 168.701
R23318 commonsourceibias.n363 commonsourceibias.n251 161.3
R23319 commonsourceibias.n361 commonsourceibias.n360 161.3
R23320 commonsourceibias.n359 commonsourceibias.n252 161.3
R23321 commonsourceibias.n358 commonsourceibias.n357 161.3
R23322 commonsourceibias.n355 commonsourceibias.n253 161.3
R23323 commonsourceibias.n354 commonsourceibias.n353 161.3
R23324 commonsourceibias.n352 commonsourceibias.n254 161.3
R23325 commonsourceibias.n351 commonsourceibias.n350 161.3
R23326 commonsourceibias.n349 commonsourceibias.n255 161.3
R23327 commonsourceibias.n347 commonsourceibias.n346 161.3
R23328 commonsourceibias.n345 commonsourceibias.n257 161.3
R23329 commonsourceibias.n344 commonsourceibias.n343 161.3
R23330 commonsourceibias.n341 commonsourceibias.n258 161.3
R23331 commonsourceibias.n340 commonsourceibias.n339 161.3
R23332 commonsourceibias.n338 commonsourceibias.n259 161.3
R23333 commonsourceibias.n337 commonsourceibias.n336 161.3
R23334 commonsourceibias.n335 commonsourceibias.n260 161.3
R23335 commonsourceibias.n333 commonsourceibias.n332 161.3
R23336 commonsourceibias.n331 commonsourceibias.n262 161.3
R23337 commonsourceibias.n330 commonsourceibias.n329 161.3
R23338 commonsourceibias.n327 commonsourceibias.n263 161.3
R23339 commonsourceibias.n326 commonsourceibias.n325 161.3
R23340 commonsourceibias.n324 commonsourceibias.n264 161.3
R23341 commonsourceibias.n323 commonsourceibias.n322 161.3
R23342 commonsourceibias.n321 commonsourceibias.n265 161.3
R23343 commonsourceibias.n319 commonsourceibias.n318 161.3
R23344 commonsourceibias.n317 commonsourceibias.n267 161.3
R23345 commonsourceibias.n316 commonsourceibias.n315 161.3
R23346 commonsourceibias.n313 commonsourceibias.n268 161.3
R23347 commonsourceibias.n312 commonsourceibias.n311 161.3
R23348 commonsourceibias.n310 commonsourceibias.n269 161.3
R23349 commonsourceibias.n309 commonsourceibias.n308 161.3
R23350 commonsourceibias.n307 commonsourceibias.n270 161.3
R23351 commonsourceibias.n305 commonsourceibias.n304 161.3
R23352 commonsourceibias.n303 commonsourceibias.n272 161.3
R23353 commonsourceibias.n302 commonsourceibias.n301 161.3
R23354 commonsourceibias.n299 commonsourceibias.n273 161.3
R23355 commonsourceibias.n298 commonsourceibias.n297 161.3
R23356 commonsourceibias.n296 commonsourceibias.n274 161.3
R23357 commonsourceibias.n295 commonsourceibias.n294 161.3
R23358 commonsourceibias.n293 commonsourceibias.n275 161.3
R23359 commonsourceibias.n291 commonsourceibias.n290 161.3
R23360 commonsourceibias.n289 commonsourceibias.n277 161.3
R23361 commonsourceibias.n288 commonsourceibias.n287 161.3
R23362 commonsourceibias.n285 commonsourceibias.n278 161.3
R23363 commonsourceibias.n284 commonsourceibias.n283 161.3
R23364 commonsourceibias.n282 commonsourceibias.n279 161.3
R23365 commonsourceibias.n45 commonsourceibias.n42 161.3
R23366 commonsourceibias.n47 commonsourceibias.n46 161.3
R23367 commonsourceibias.n48 commonsourceibias.n41 161.3
R23368 commonsourceibias.n51 commonsourceibias.n50 161.3
R23369 commonsourceibias.n52 commonsourceibias.n40 161.3
R23370 commonsourceibias.n54 commonsourceibias.n53 161.3
R23371 commonsourceibias.n56 commonsourceibias.n38 161.3
R23372 commonsourceibias.n58 commonsourceibias.n57 161.3
R23373 commonsourceibias.n59 commonsourceibias.n37 161.3
R23374 commonsourceibias.n61 commonsourceibias.n60 161.3
R23375 commonsourceibias.n62 commonsourceibias.n36 161.3
R23376 commonsourceibias.n65 commonsourceibias.n64 161.3
R23377 commonsourceibias.n66 commonsourceibias.n35 161.3
R23378 commonsourceibias.n68 commonsourceibias.n67 161.3
R23379 commonsourceibias.n70 commonsourceibias.n33 161.3
R23380 commonsourceibias.n72 commonsourceibias.n71 161.3
R23381 commonsourceibias.n73 commonsourceibias.n32 161.3
R23382 commonsourceibias.n75 commonsourceibias.n74 161.3
R23383 commonsourceibias.n76 commonsourceibias.n31 161.3
R23384 commonsourceibias.n79 commonsourceibias.n78 161.3
R23385 commonsourceibias.n80 commonsourceibias.n30 161.3
R23386 commonsourceibias.n82 commonsourceibias.n81 161.3
R23387 commonsourceibias.n84 commonsourceibias.n28 161.3
R23388 commonsourceibias.n86 commonsourceibias.n85 161.3
R23389 commonsourceibias.n87 commonsourceibias.n27 161.3
R23390 commonsourceibias.n89 commonsourceibias.n88 161.3
R23391 commonsourceibias.n90 commonsourceibias.n26 161.3
R23392 commonsourceibias.n93 commonsourceibias.n92 161.3
R23393 commonsourceibias.n94 commonsourceibias.n25 161.3
R23394 commonsourceibias.n96 commonsourceibias.n95 161.3
R23395 commonsourceibias.n98 commonsourceibias.n23 161.3
R23396 commonsourceibias.n100 commonsourceibias.n99 161.3
R23397 commonsourceibias.n101 commonsourceibias.n22 161.3
R23398 commonsourceibias.n103 commonsourceibias.n102 161.3
R23399 commonsourceibias.n104 commonsourceibias.n21 161.3
R23400 commonsourceibias.n107 commonsourceibias.n106 161.3
R23401 commonsourceibias.n108 commonsourceibias.n20 161.3
R23402 commonsourceibias.n110 commonsourceibias.n109 161.3
R23403 commonsourceibias.n112 commonsourceibias.n18 161.3
R23404 commonsourceibias.n114 commonsourceibias.n113 161.3
R23405 commonsourceibias.n115 commonsourceibias.n17 161.3
R23406 commonsourceibias.n117 commonsourceibias.n116 161.3
R23407 commonsourceibias.n118 commonsourceibias.n16 161.3
R23408 commonsourceibias.n121 commonsourceibias.n120 161.3
R23409 commonsourceibias.n122 commonsourceibias.n15 161.3
R23410 commonsourceibias.n124 commonsourceibias.n123 161.3
R23411 commonsourceibias.n126 commonsourceibias.n14 161.3
R23412 commonsourceibias.n167 commonsourceibias.n164 161.3
R23413 commonsourceibias.n169 commonsourceibias.n168 161.3
R23414 commonsourceibias.n170 commonsourceibias.n163 161.3
R23415 commonsourceibias.n173 commonsourceibias.n172 161.3
R23416 commonsourceibias.n174 commonsourceibias.n162 161.3
R23417 commonsourceibias.n176 commonsourceibias.n175 161.3
R23418 commonsourceibias.n178 commonsourceibias.n160 161.3
R23419 commonsourceibias.n180 commonsourceibias.n179 161.3
R23420 commonsourceibias.n181 commonsourceibias.n159 161.3
R23421 commonsourceibias.n183 commonsourceibias.n182 161.3
R23422 commonsourceibias.n184 commonsourceibias.n158 161.3
R23423 commonsourceibias.n187 commonsourceibias.n186 161.3
R23424 commonsourceibias.n188 commonsourceibias.n157 161.3
R23425 commonsourceibias.n190 commonsourceibias.n189 161.3
R23426 commonsourceibias.n192 commonsourceibias.n156 161.3
R23427 commonsourceibias.n194 commonsourceibias.n193 161.3
R23428 commonsourceibias.n196 commonsourceibias.n195 161.3
R23429 commonsourceibias.n197 commonsourceibias.n154 161.3
R23430 commonsourceibias.n199 commonsourceibias.n198 161.3
R23431 commonsourceibias.n201 commonsourceibias.n200 161.3
R23432 commonsourceibias.n202 commonsourceibias.n152 161.3
R23433 commonsourceibias.n204 commonsourceibias.n203 161.3
R23434 commonsourceibias.n206 commonsourceibias.n205 161.3
R23435 commonsourceibias.n208 commonsourceibias.n207 161.3
R23436 commonsourceibias.n209 commonsourceibias.n13 161.3
R23437 commonsourceibias.n211 commonsourceibias.n210 161.3
R23438 commonsourceibias.n212 commonsourceibias.n12 161.3
R23439 commonsourceibias.n215 commonsourceibias.n214 161.3
R23440 commonsourceibias.n216 commonsourceibias.n11 161.3
R23441 commonsourceibias.n218 commonsourceibias.n217 161.3
R23442 commonsourceibias.n220 commonsourceibias.n9 161.3
R23443 commonsourceibias.n222 commonsourceibias.n221 161.3
R23444 commonsourceibias.n223 commonsourceibias.n8 161.3
R23445 commonsourceibias.n225 commonsourceibias.n224 161.3
R23446 commonsourceibias.n226 commonsourceibias.n7 161.3
R23447 commonsourceibias.n229 commonsourceibias.n228 161.3
R23448 commonsourceibias.n230 commonsourceibias.n6 161.3
R23449 commonsourceibias.n232 commonsourceibias.n231 161.3
R23450 commonsourceibias.n234 commonsourceibias.n4 161.3
R23451 commonsourceibias.n236 commonsourceibias.n235 161.3
R23452 commonsourceibias.n237 commonsourceibias.n3 161.3
R23453 commonsourceibias.n239 commonsourceibias.n238 161.3
R23454 commonsourceibias.n240 commonsourceibias.n2 161.3
R23455 commonsourceibias.n243 commonsourceibias.n242 161.3
R23456 commonsourceibias.n244 commonsourceibias.n1 161.3
R23457 commonsourceibias.n246 commonsourceibias.n245 161.3
R23458 commonsourceibias.n248 commonsourceibias.n0 161.3
R23459 commonsourceibias.n730 commonsourceibias.n618 161.3
R23460 commonsourceibias.n728 commonsourceibias.n727 161.3
R23461 commonsourceibias.n726 commonsourceibias.n619 161.3
R23462 commonsourceibias.n725 commonsourceibias.n724 161.3
R23463 commonsourceibias.n722 commonsourceibias.n620 161.3
R23464 commonsourceibias.n721 commonsourceibias.n720 161.3
R23465 commonsourceibias.n719 commonsourceibias.n621 161.3
R23466 commonsourceibias.n718 commonsourceibias.n717 161.3
R23467 commonsourceibias.n715 commonsourceibias.n622 161.3
R23468 commonsourceibias.n713 commonsourceibias.n712 161.3
R23469 commonsourceibias.n711 commonsourceibias.n623 161.3
R23470 commonsourceibias.n710 commonsourceibias.n709 161.3
R23471 commonsourceibias.n707 commonsourceibias.n624 161.3
R23472 commonsourceibias.n706 commonsourceibias.n705 161.3
R23473 commonsourceibias.n704 commonsourceibias.n625 161.3
R23474 commonsourceibias.n703 commonsourceibias.n702 161.3
R23475 commonsourceibias.n700 commonsourceibias.n626 161.3
R23476 commonsourceibias.n698 commonsourceibias.n697 161.3
R23477 commonsourceibias.n696 commonsourceibias.n627 161.3
R23478 commonsourceibias.n695 commonsourceibias.n694 161.3
R23479 commonsourceibias.n692 commonsourceibias.n628 161.3
R23480 commonsourceibias.n691 commonsourceibias.n690 161.3
R23481 commonsourceibias.n689 commonsourceibias.n629 161.3
R23482 commonsourceibias.n688 commonsourceibias.n687 161.3
R23483 commonsourceibias.n685 commonsourceibias.n630 161.3
R23484 commonsourceibias.n683 commonsourceibias.n682 161.3
R23485 commonsourceibias.n681 commonsourceibias.n631 161.3
R23486 commonsourceibias.n680 commonsourceibias.n679 161.3
R23487 commonsourceibias.n677 commonsourceibias.n632 161.3
R23488 commonsourceibias.n676 commonsourceibias.n675 161.3
R23489 commonsourceibias.n674 commonsourceibias.n633 161.3
R23490 commonsourceibias.n673 commonsourceibias.n672 161.3
R23491 commonsourceibias.n670 commonsourceibias.n634 161.3
R23492 commonsourceibias.n668 commonsourceibias.n667 161.3
R23493 commonsourceibias.n666 commonsourceibias.n635 161.3
R23494 commonsourceibias.n665 commonsourceibias.n664 161.3
R23495 commonsourceibias.n662 commonsourceibias.n636 161.3
R23496 commonsourceibias.n661 commonsourceibias.n660 161.3
R23497 commonsourceibias.n659 commonsourceibias.n637 161.3
R23498 commonsourceibias.n658 commonsourceibias.n657 161.3
R23499 commonsourceibias.n655 commonsourceibias.n638 161.3
R23500 commonsourceibias.n653 commonsourceibias.n652 161.3
R23501 commonsourceibias.n651 commonsourceibias.n639 161.3
R23502 commonsourceibias.n650 commonsourceibias.n649 161.3
R23503 commonsourceibias.n647 commonsourceibias.n640 161.3
R23504 commonsourceibias.n646 commonsourceibias.n645 161.3
R23505 commonsourceibias.n644 commonsourceibias.n641 161.3
R23506 commonsourceibias.n500 commonsourceibias.n388 161.3
R23507 commonsourceibias.n498 commonsourceibias.n497 161.3
R23508 commonsourceibias.n496 commonsourceibias.n389 161.3
R23509 commonsourceibias.n495 commonsourceibias.n494 161.3
R23510 commonsourceibias.n492 commonsourceibias.n390 161.3
R23511 commonsourceibias.n491 commonsourceibias.n490 161.3
R23512 commonsourceibias.n489 commonsourceibias.n391 161.3
R23513 commonsourceibias.n488 commonsourceibias.n487 161.3
R23514 commonsourceibias.n485 commonsourceibias.n392 161.3
R23515 commonsourceibias.n483 commonsourceibias.n482 161.3
R23516 commonsourceibias.n481 commonsourceibias.n393 161.3
R23517 commonsourceibias.n480 commonsourceibias.n479 161.3
R23518 commonsourceibias.n477 commonsourceibias.n394 161.3
R23519 commonsourceibias.n476 commonsourceibias.n475 161.3
R23520 commonsourceibias.n474 commonsourceibias.n395 161.3
R23521 commonsourceibias.n473 commonsourceibias.n472 161.3
R23522 commonsourceibias.n470 commonsourceibias.n396 161.3
R23523 commonsourceibias.n468 commonsourceibias.n467 161.3
R23524 commonsourceibias.n466 commonsourceibias.n397 161.3
R23525 commonsourceibias.n465 commonsourceibias.n464 161.3
R23526 commonsourceibias.n462 commonsourceibias.n398 161.3
R23527 commonsourceibias.n461 commonsourceibias.n460 161.3
R23528 commonsourceibias.n459 commonsourceibias.n399 161.3
R23529 commonsourceibias.n458 commonsourceibias.n457 161.3
R23530 commonsourceibias.n455 commonsourceibias.n400 161.3
R23531 commonsourceibias.n453 commonsourceibias.n452 161.3
R23532 commonsourceibias.n451 commonsourceibias.n401 161.3
R23533 commonsourceibias.n450 commonsourceibias.n449 161.3
R23534 commonsourceibias.n447 commonsourceibias.n402 161.3
R23535 commonsourceibias.n446 commonsourceibias.n445 161.3
R23536 commonsourceibias.n444 commonsourceibias.n403 161.3
R23537 commonsourceibias.n443 commonsourceibias.n442 161.3
R23538 commonsourceibias.n440 commonsourceibias.n404 161.3
R23539 commonsourceibias.n438 commonsourceibias.n437 161.3
R23540 commonsourceibias.n436 commonsourceibias.n405 161.3
R23541 commonsourceibias.n435 commonsourceibias.n434 161.3
R23542 commonsourceibias.n432 commonsourceibias.n406 161.3
R23543 commonsourceibias.n431 commonsourceibias.n430 161.3
R23544 commonsourceibias.n429 commonsourceibias.n407 161.3
R23545 commonsourceibias.n428 commonsourceibias.n427 161.3
R23546 commonsourceibias.n425 commonsourceibias.n408 161.3
R23547 commonsourceibias.n423 commonsourceibias.n422 161.3
R23548 commonsourceibias.n421 commonsourceibias.n409 161.3
R23549 commonsourceibias.n420 commonsourceibias.n419 161.3
R23550 commonsourceibias.n417 commonsourceibias.n410 161.3
R23551 commonsourceibias.n416 commonsourceibias.n415 161.3
R23552 commonsourceibias.n414 commonsourceibias.n411 161.3
R23553 commonsourceibias.n570 commonsourceibias.n569 161.3
R23554 commonsourceibias.n568 commonsourceibias.n567 161.3
R23555 commonsourceibias.n566 commonsourceibias.n516 161.3
R23556 commonsourceibias.n565 commonsourceibias.n564 161.3
R23557 commonsourceibias.n563 commonsourceibias.n562 161.3
R23558 commonsourceibias.n561 commonsourceibias.n518 161.3
R23559 commonsourceibias.n560 commonsourceibias.n559 161.3
R23560 commonsourceibias.n558 commonsourceibias.n557 161.3
R23561 commonsourceibias.n556 commonsourceibias.n520 161.3
R23562 commonsourceibias.n554 commonsourceibias.n553 161.3
R23563 commonsourceibias.n552 commonsourceibias.n521 161.3
R23564 commonsourceibias.n551 commonsourceibias.n550 161.3
R23565 commonsourceibias.n548 commonsourceibias.n522 161.3
R23566 commonsourceibias.n547 commonsourceibias.n546 161.3
R23567 commonsourceibias.n545 commonsourceibias.n523 161.3
R23568 commonsourceibias.n544 commonsourceibias.n543 161.3
R23569 commonsourceibias.n541 commonsourceibias.n524 161.3
R23570 commonsourceibias.n539 commonsourceibias.n538 161.3
R23571 commonsourceibias.n537 commonsourceibias.n525 161.3
R23572 commonsourceibias.n536 commonsourceibias.n535 161.3
R23573 commonsourceibias.n533 commonsourceibias.n526 161.3
R23574 commonsourceibias.n532 commonsourceibias.n531 161.3
R23575 commonsourceibias.n530 commonsourceibias.n527 161.3
R23576 commonsourceibias.n615 commonsourceibias.n367 161.3
R23577 commonsourceibias.n613 commonsourceibias.n612 161.3
R23578 commonsourceibias.n611 commonsourceibias.n368 161.3
R23579 commonsourceibias.n610 commonsourceibias.n609 161.3
R23580 commonsourceibias.n607 commonsourceibias.n369 161.3
R23581 commonsourceibias.n606 commonsourceibias.n605 161.3
R23582 commonsourceibias.n604 commonsourceibias.n370 161.3
R23583 commonsourceibias.n603 commonsourceibias.n602 161.3
R23584 commonsourceibias.n600 commonsourceibias.n371 161.3
R23585 commonsourceibias.n598 commonsourceibias.n597 161.3
R23586 commonsourceibias.n596 commonsourceibias.n372 161.3
R23587 commonsourceibias.n595 commonsourceibias.n594 161.3
R23588 commonsourceibias.n592 commonsourceibias.n373 161.3
R23589 commonsourceibias.n591 commonsourceibias.n590 161.3
R23590 commonsourceibias.n589 commonsourceibias.n374 161.3
R23591 commonsourceibias.n588 commonsourceibias.n587 161.3
R23592 commonsourceibias.n585 commonsourceibias.n375 161.3
R23593 commonsourceibias.n583 commonsourceibias.n582 161.3
R23594 commonsourceibias.n581 commonsourceibias.n376 161.3
R23595 commonsourceibias.n580 commonsourceibias.n579 161.3
R23596 commonsourceibias.n577 commonsourceibias.n377 161.3
R23597 commonsourceibias.n576 commonsourceibias.n575 161.3
R23598 commonsourceibias.n574 commonsourceibias.n378 161.3
R23599 commonsourceibias.n573 commonsourceibias.n572 161.3
R23600 commonsourceibias.n141 commonsourceibias.n139 81.5057
R23601 commonsourceibias.n381 commonsourceibias.n379 81.5057
R23602 commonsourceibias.n141 commonsourceibias.n140 80.9324
R23603 commonsourceibias.n143 commonsourceibias.n142 80.9324
R23604 commonsourceibias.n145 commonsourceibias.n144 80.9324
R23605 commonsourceibias.n147 commonsourceibias.n146 80.9324
R23606 commonsourceibias.n138 commonsourceibias.n137 80.9324
R23607 commonsourceibias.n136 commonsourceibias.n135 80.9324
R23608 commonsourceibias.n134 commonsourceibias.n133 80.9324
R23609 commonsourceibias.n132 commonsourceibias.n131 80.9324
R23610 commonsourceibias.n130 commonsourceibias.n129 80.9324
R23611 commonsourceibias.n504 commonsourceibias.n503 80.9324
R23612 commonsourceibias.n506 commonsourceibias.n505 80.9324
R23613 commonsourceibias.n508 commonsourceibias.n507 80.9324
R23614 commonsourceibias.n510 commonsourceibias.n509 80.9324
R23615 commonsourceibias.n512 commonsourceibias.n511 80.9324
R23616 commonsourceibias.n387 commonsourceibias.n386 80.9324
R23617 commonsourceibias.n385 commonsourceibias.n384 80.9324
R23618 commonsourceibias.n383 commonsourceibias.n382 80.9324
R23619 commonsourceibias.n381 commonsourceibias.n380 80.9324
R23620 commonsourceibias.n365 commonsourceibias.n364 80.6037
R23621 commonsourceibias.n128 commonsourceibias.n127 80.6037
R23622 commonsourceibias.n250 commonsourceibias.n249 80.6037
R23623 commonsourceibias.n732 commonsourceibias.n731 80.6037
R23624 commonsourceibias.n502 commonsourceibias.n501 80.6037
R23625 commonsourceibias.n617 commonsourceibias.n616 80.6037
R23626 commonsourceibias.n322 commonsourceibias.n321 56.5617
R23627 commonsourceibias.n336 commonsourceibias.n335 56.5617
R23628 commonsourceibias.n85 commonsourceibias.n84 56.5617
R23629 commonsourceibias.n71 commonsourceibias.n70 56.5617
R23630 commonsourceibias.n207 commonsourceibias.n206 56.5617
R23631 commonsourceibias.n193 commonsourceibias.n192 56.5617
R23632 commonsourceibias.n687 commonsourceibias.n685 56.5617
R23633 commonsourceibias.n702 commonsourceibias.n700 56.5617
R23634 commonsourceibias.n457 commonsourceibias.n455 56.5617
R23635 commonsourceibias.n472 commonsourceibias.n470 56.5617
R23636 commonsourceibias.n572 commonsourceibias.n570 56.5617
R23637 commonsourceibias.n294 commonsourceibias.n293 56.5617
R23638 commonsourceibias.n308 commonsourceibias.n307 56.5617
R23639 commonsourceibias.n350 commonsourceibias.n349 56.5617
R23640 commonsourceibias.n113 commonsourceibias.n112 56.5617
R23641 commonsourceibias.n99 commonsourceibias.n98 56.5617
R23642 commonsourceibias.n57 commonsourceibias.n56 56.5617
R23643 commonsourceibias.n235 commonsourceibias.n234 56.5617
R23644 commonsourceibias.n221 commonsourceibias.n220 56.5617
R23645 commonsourceibias.n179 commonsourceibias.n178 56.5617
R23646 commonsourceibias.n657 commonsourceibias.n655 56.5617
R23647 commonsourceibias.n672 commonsourceibias.n670 56.5617
R23648 commonsourceibias.n717 commonsourceibias.n715 56.5617
R23649 commonsourceibias.n427 commonsourceibias.n425 56.5617
R23650 commonsourceibias.n442 commonsourceibias.n440 56.5617
R23651 commonsourceibias.n487 commonsourceibias.n485 56.5617
R23652 commonsourceibias.n602 commonsourceibias.n600 56.5617
R23653 commonsourceibias.n587 commonsourceibias.n585 56.5617
R23654 commonsourceibias.n543 commonsourceibias.n541 56.5617
R23655 commonsourceibias.n557 commonsourceibias.n556 56.5617
R23656 commonsourceibias.n285 commonsourceibias.n284 51.2335
R23657 commonsourceibias.n357 commonsourceibias.n252 51.2335
R23658 commonsourceibias.n120 commonsourceibias.n15 51.2335
R23659 commonsourceibias.n48 commonsourceibias.n47 51.2335
R23660 commonsourceibias.n242 commonsourceibias.n1 51.2335
R23661 commonsourceibias.n170 commonsourceibias.n169 51.2335
R23662 commonsourceibias.n647 commonsourceibias.n646 51.2335
R23663 commonsourceibias.n724 commonsourceibias.n619 51.2335
R23664 commonsourceibias.n417 commonsourceibias.n416 51.2335
R23665 commonsourceibias.n494 commonsourceibias.n389 51.2335
R23666 commonsourceibias.n609 commonsourceibias.n368 51.2335
R23667 commonsourceibias.n533 commonsourceibias.n532 51.2335
R23668 commonsourceibias.n364 commonsourceibias.n363 50.9056
R23669 commonsourceibias.n127 commonsourceibias.n126 50.9056
R23670 commonsourceibias.n249 commonsourceibias.n248 50.9056
R23671 commonsourceibias.n731 commonsourceibias.n730 50.9056
R23672 commonsourceibias.n501 commonsourceibias.n500 50.9056
R23673 commonsourceibias.n616 commonsourceibias.n615 50.9056
R23674 commonsourceibias.n299 commonsourceibias.n298 50.2647
R23675 commonsourceibias.n343 commonsourceibias.n257 50.2647
R23676 commonsourceibias.n106 commonsourceibias.n20 50.2647
R23677 commonsourceibias.n62 commonsourceibias.n61 50.2647
R23678 commonsourceibias.n228 commonsourceibias.n6 50.2647
R23679 commonsourceibias.n184 commonsourceibias.n183 50.2647
R23680 commonsourceibias.n662 commonsourceibias.n661 50.2647
R23681 commonsourceibias.n709 commonsourceibias.n623 50.2647
R23682 commonsourceibias.n432 commonsourceibias.n431 50.2647
R23683 commonsourceibias.n479 commonsourceibias.n393 50.2647
R23684 commonsourceibias.n594 commonsourceibias.n372 50.2647
R23685 commonsourceibias.n548 commonsourceibias.n547 50.2647
R23686 commonsourceibias.n281 commonsourceibias.n280 49.9027
R23687 commonsourceibias.n44 commonsourceibias.n43 49.9027
R23688 commonsourceibias.n166 commonsourceibias.n165 49.9027
R23689 commonsourceibias.n643 commonsourceibias.n642 49.9027
R23690 commonsourceibias.n413 commonsourceibias.n412 49.9027
R23691 commonsourceibias.n529 commonsourceibias.n528 49.9027
R23692 commonsourceibias.n313 commonsourceibias.n312 49.296
R23693 commonsourceibias.n329 commonsourceibias.n262 49.296
R23694 commonsourceibias.n92 commonsourceibias.n25 49.296
R23695 commonsourceibias.n76 commonsourceibias.n75 49.296
R23696 commonsourceibias.n214 commonsourceibias.n11 49.296
R23697 commonsourceibias.n198 commonsourceibias.n197 49.296
R23698 commonsourceibias.n677 commonsourceibias.n676 49.296
R23699 commonsourceibias.n694 commonsourceibias.n627 49.296
R23700 commonsourceibias.n447 commonsourceibias.n446 49.296
R23701 commonsourceibias.n464 commonsourceibias.n397 49.296
R23702 commonsourceibias.n579 commonsourceibias.n376 49.296
R23703 commonsourceibias.n562 commonsourceibias.n561 49.296
R23704 commonsourceibias.n315 commonsourceibias.n267 48.3272
R23705 commonsourceibias.n327 commonsourceibias.n326 48.3272
R23706 commonsourceibias.n90 commonsourceibias.n89 48.3272
R23707 commonsourceibias.n78 commonsourceibias.n30 48.3272
R23708 commonsourceibias.n212 commonsourceibias.n211 48.3272
R23709 commonsourceibias.n202 commonsourceibias.n201 48.3272
R23710 commonsourceibias.n679 commonsourceibias.n631 48.3272
R23711 commonsourceibias.n692 commonsourceibias.n691 48.3272
R23712 commonsourceibias.n449 commonsourceibias.n401 48.3272
R23713 commonsourceibias.n462 commonsourceibias.n461 48.3272
R23714 commonsourceibias.n577 commonsourceibias.n576 48.3272
R23715 commonsourceibias.n566 commonsourceibias.n565 48.3272
R23716 commonsourceibias.n301 commonsourceibias.n272 47.3584
R23717 commonsourceibias.n341 commonsourceibias.n340 47.3584
R23718 commonsourceibias.n104 commonsourceibias.n103 47.3584
R23719 commonsourceibias.n64 commonsourceibias.n35 47.3584
R23720 commonsourceibias.n226 commonsourceibias.n225 47.3584
R23721 commonsourceibias.n186 commonsourceibias.n157 47.3584
R23722 commonsourceibias.n664 commonsourceibias.n635 47.3584
R23723 commonsourceibias.n707 commonsourceibias.n706 47.3584
R23724 commonsourceibias.n434 commonsourceibias.n405 47.3584
R23725 commonsourceibias.n477 commonsourceibias.n476 47.3584
R23726 commonsourceibias.n592 commonsourceibias.n591 47.3584
R23727 commonsourceibias.n550 commonsourceibias.n521 47.3584
R23728 commonsourceibias.n287 commonsourceibias.n277 46.3896
R23729 commonsourceibias.n355 commonsourceibias.n354 46.3896
R23730 commonsourceibias.n118 commonsourceibias.n117 46.3896
R23731 commonsourceibias.n50 commonsourceibias.n40 46.3896
R23732 commonsourceibias.n240 commonsourceibias.n239 46.3896
R23733 commonsourceibias.n172 commonsourceibias.n162 46.3896
R23734 commonsourceibias.n649 commonsourceibias.n639 46.3896
R23735 commonsourceibias.n722 commonsourceibias.n721 46.3896
R23736 commonsourceibias.n419 commonsourceibias.n409 46.3896
R23737 commonsourceibias.n492 commonsourceibias.n491 46.3896
R23738 commonsourceibias.n607 commonsourceibias.n606 46.3896
R23739 commonsourceibias.n535 commonsourceibias.n525 46.3896
R23740 commonsourceibias.n282 commonsourceibias.n281 44.7059
R23741 commonsourceibias.n644 commonsourceibias.n643 44.7059
R23742 commonsourceibias.n414 commonsourceibias.n413 44.7059
R23743 commonsourceibias.n530 commonsourceibias.n529 44.7059
R23744 commonsourceibias.n45 commonsourceibias.n44 44.7059
R23745 commonsourceibias.n167 commonsourceibias.n166 44.7059
R23746 commonsourceibias.n291 commonsourceibias.n277 34.7644
R23747 commonsourceibias.n354 commonsourceibias.n254 34.7644
R23748 commonsourceibias.n117 commonsourceibias.n17 34.7644
R23749 commonsourceibias.n54 commonsourceibias.n40 34.7644
R23750 commonsourceibias.n239 commonsourceibias.n3 34.7644
R23751 commonsourceibias.n176 commonsourceibias.n162 34.7644
R23752 commonsourceibias.n653 commonsourceibias.n639 34.7644
R23753 commonsourceibias.n721 commonsourceibias.n621 34.7644
R23754 commonsourceibias.n423 commonsourceibias.n409 34.7644
R23755 commonsourceibias.n491 commonsourceibias.n391 34.7644
R23756 commonsourceibias.n606 commonsourceibias.n370 34.7644
R23757 commonsourceibias.n539 commonsourceibias.n525 34.7644
R23758 commonsourceibias.n305 commonsourceibias.n272 33.7956
R23759 commonsourceibias.n340 commonsourceibias.n259 33.7956
R23760 commonsourceibias.n103 commonsourceibias.n22 33.7956
R23761 commonsourceibias.n68 commonsourceibias.n35 33.7956
R23762 commonsourceibias.n225 commonsourceibias.n8 33.7956
R23763 commonsourceibias.n190 commonsourceibias.n157 33.7956
R23764 commonsourceibias.n668 commonsourceibias.n635 33.7956
R23765 commonsourceibias.n706 commonsourceibias.n625 33.7956
R23766 commonsourceibias.n438 commonsourceibias.n405 33.7956
R23767 commonsourceibias.n476 commonsourceibias.n395 33.7956
R23768 commonsourceibias.n591 commonsourceibias.n374 33.7956
R23769 commonsourceibias.n554 commonsourceibias.n521 33.7956
R23770 commonsourceibias.n319 commonsourceibias.n267 32.8269
R23771 commonsourceibias.n326 commonsourceibias.n264 32.8269
R23772 commonsourceibias.n89 commonsourceibias.n27 32.8269
R23773 commonsourceibias.n82 commonsourceibias.n30 32.8269
R23774 commonsourceibias.n211 commonsourceibias.n13 32.8269
R23775 commonsourceibias.n203 commonsourceibias.n202 32.8269
R23776 commonsourceibias.n683 commonsourceibias.n631 32.8269
R23777 commonsourceibias.n691 commonsourceibias.n629 32.8269
R23778 commonsourceibias.n453 commonsourceibias.n401 32.8269
R23779 commonsourceibias.n461 commonsourceibias.n399 32.8269
R23780 commonsourceibias.n576 commonsourceibias.n378 32.8269
R23781 commonsourceibias.n567 commonsourceibias.n566 32.8269
R23782 commonsourceibias.n312 commonsourceibias.n269 31.8581
R23783 commonsourceibias.n333 commonsourceibias.n262 31.8581
R23784 commonsourceibias.n96 commonsourceibias.n25 31.8581
R23785 commonsourceibias.n75 commonsourceibias.n32 31.8581
R23786 commonsourceibias.n218 commonsourceibias.n11 31.8581
R23787 commonsourceibias.n197 commonsourceibias.n196 31.8581
R23788 commonsourceibias.n676 commonsourceibias.n633 31.8581
R23789 commonsourceibias.n698 commonsourceibias.n627 31.8581
R23790 commonsourceibias.n446 commonsourceibias.n403 31.8581
R23791 commonsourceibias.n468 commonsourceibias.n397 31.8581
R23792 commonsourceibias.n583 commonsourceibias.n376 31.8581
R23793 commonsourceibias.n561 commonsourceibias.n560 31.8581
R23794 commonsourceibias.n298 commonsourceibias.n274 30.8893
R23795 commonsourceibias.n347 commonsourceibias.n257 30.8893
R23796 commonsourceibias.n110 commonsourceibias.n20 30.8893
R23797 commonsourceibias.n61 commonsourceibias.n37 30.8893
R23798 commonsourceibias.n232 commonsourceibias.n6 30.8893
R23799 commonsourceibias.n183 commonsourceibias.n159 30.8893
R23800 commonsourceibias.n661 commonsourceibias.n637 30.8893
R23801 commonsourceibias.n713 commonsourceibias.n623 30.8893
R23802 commonsourceibias.n431 commonsourceibias.n407 30.8893
R23803 commonsourceibias.n483 commonsourceibias.n393 30.8893
R23804 commonsourceibias.n598 commonsourceibias.n372 30.8893
R23805 commonsourceibias.n547 commonsourceibias.n523 30.8893
R23806 commonsourceibias.n284 commonsourceibias.n279 29.9206
R23807 commonsourceibias.n361 commonsourceibias.n252 29.9206
R23808 commonsourceibias.n124 commonsourceibias.n15 29.9206
R23809 commonsourceibias.n47 commonsourceibias.n42 29.9206
R23810 commonsourceibias.n246 commonsourceibias.n1 29.9206
R23811 commonsourceibias.n169 commonsourceibias.n164 29.9206
R23812 commonsourceibias.n646 commonsourceibias.n641 29.9206
R23813 commonsourceibias.n728 commonsourceibias.n619 29.9206
R23814 commonsourceibias.n416 commonsourceibias.n411 29.9206
R23815 commonsourceibias.n498 commonsourceibias.n389 29.9206
R23816 commonsourceibias.n613 commonsourceibias.n368 29.9206
R23817 commonsourceibias.n532 commonsourceibias.n527 29.9206
R23818 commonsourceibias.n363 commonsourceibias.n362 21.8872
R23819 commonsourceibias.n126 commonsourceibias.n125 21.8872
R23820 commonsourceibias.n248 commonsourceibias.n247 21.8872
R23821 commonsourceibias.n730 commonsourceibias.n729 21.8872
R23822 commonsourceibias.n500 commonsourceibias.n499 21.8872
R23823 commonsourceibias.n615 commonsourceibias.n614 21.8872
R23824 commonsourceibias.n294 commonsourceibias.n276 21.3954
R23825 commonsourceibias.n349 commonsourceibias.n348 21.3954
R23826 commonsourceibias.n112 commonsourceibias.n111 21.3954
R23827 commonsourceibias.n57 commonsourceibias.n39 21.3954
R23828 commonsourceibias.n234 commonsourceibias.n233 21.3954
R23829 commonsourceibias.n179 commonsourceibias.n161 21.3954
R23830 commonsourceibias.n657 commonsourceibias.n656 21.3954
R23831 commonsourceibias.n715 commonsourceibias.n714 21.3954
R23832 commonsourceibias.n427 commonsourceibias.n426 21.3954
R23833 commonsourceibias.n485 commonsourceibias.n484 21.3954
R23834 commonsourceibias.n600 commonsourceibias.n599 21.3954
R23835 commonsourceibias.n543 commonsourceibias.n542 21.3954
R23836 commonsourceibias.n308 commonsourceibias.n271 20.9036
R23837 commonsourceibias.n335 commonsourceibias.n334 20.9036
R23838 commonsourceibias.n98 commonsourceibias.n97 20.9036
R23839 commonsourceibias.n71 commonsourceibias.n34 20.9036
R23840 commonsourceibias.n220 commonsourceibias.n219 20.9036
R23841 commonsourceibias.n193 commonsourceibias.n155 20.9036
R23842 commonsourceibias.n672 commonsourceibias.n671 20.9036
R23843 commonsourceibias.n700 commonsourceibias.n699 20.9036
R23844 commonsourceibias.n442 commonsourceibias.n441 20.9036
R23845 commonsourceibias.n470 commonsourceibias.n469 20.9036
R23846 commonsourceibias.n585 commonsourceibias.n584 20.9036
R23847 commonsourceibias.n557 commonsourceibias.n519 20.9036
R23848 commonsourceibias.n321 commonsourceibias.n320 20.4117
R23849 commonsourceibias.n322 commonsourceibias.n266 20.4117
R23850 commonsourceibias.n85 commonsourceibias.n29 20.4117
R23851 commonsourceibias.n84 commonsourceibias.n83 20.4117
R23852 commonsourceibias.n207 commonsourceibias.n150 20.4117
R23853 commonsourceibias.n206 commonsourceibias.n151 20.4117
R23854 commonsourceibias.n685 commonsourceibias.n684 20.4117
R23855 commonsourceibias.n687 commonsourceibias.n686 20.4117
R23856 commonsourceibias.n455 commonsourceibias.n454 20.4117
R23857 commonsourceibias.n457 commonsourceibias.n456 20.4117
R23858 commonsourceibias.n572 commonsourceibias.n571 20.4117
R23859 commonsourceibias.n570 commonsourceibias.n515 20.4117
R23860 commonsourceibias.n307 commonsourceibias.n306 19.9199
R23861 commonsourceibias.n336 commonsourceibias.n261 19.9199
R23862 commonsourceibias.n99 commonsourceibias.n24 19.9199
R23863 commonsourceibias.n70 commonsourceibias.n69 19.9199
R23864 commonsourceibias.n221 commonsourceibias.n10 19.9199
R23865 commonsourceibias.n192 commonsourceibias.n191 19.9199
R23866 commonsourceibias.n670 commonsourceibias.n669 19.9199
R23867 commonsourceibias.n702 commonsourceibias.n701 19.9199
R23868 commonsourceibias.n440 commonsourceibias.n439 19.9199
R23869 commonsourceibias.n472 commonsourceibias.n471 19.9199
R23870 commonsourceibias.n587 commonsourceibias.n586 19.9199
R23871 commonsourceibias.n556 commonsourceibias.n555 19.9199
R23872 commonsourceibias.n293 commonsourceibias.n292 19.4281
R23873 commonsourceibias.n350 commonsourceibias.n256 19.4281
R23874 commonsourceibias.n113 commonsourceibias.n19 19.4281
R23875 commonsourceibias.n56 commonsourceibias.n55 19.4281
R23876 commonsourceibias.n235 commonsourceibias.n5 19.4281
R23877 commonsourceibias.n178 commonsourceibias.n177 19.4281
R23878 commonsourceibias.n655 commonsourceibias.n654 19.4281
R23879 commonsourceibias.n717 commonsourceibias.n716 19.4281
R23880 commonsourceibias.n425 commonsourceibias.n424 19.4281
R23881 commonsourceibias.n487 commonsourceibias.n486 19.4281
R23882 commonsourceibias.n602 commonsourceibias.n601 19.4281
R23883 commonsourceibias.n541 commonsourceibias.n540 19.4281
R23884 commonsourceibias.n286 commonsourceibias.n285 13.526
R23885 commonsourceibias.n357 commonsourceibias.n356 13.526
R23886 commonsourceibias.n120 commonsourceibias.n119 13.526
R23887 commonsourceibias.n49 commonsourceibias.n48 13.526
R23888 commonsourceibias.n242 commonsourceibias.n241 13.526
R23889 commonsourceibias.n171 commonsourceibias.n170 13.526
R23890 commonsourceibias.n648 commonsourceibias.n647 13.526
R23891 commonsourceibias.n724 commonsourceibias.n723 13.526
R23892 commonsourceibias.n418 commonsourceibias.n417 13.526
R23893 commonsourceibias.n494 commonsourceibias.n493 13.526
R23894 commonsourceibias.n609 commonsourceibias.n608 13.526
R23895 commonsourceibias.n534 commonsourceibias.n533 13.526
R23896 commonsourceibias.n130 commonsourceibias.n128 13.2322
R23897 commonsourceibias.n504 commonsourceibias.n502 13.2322
R23898 commonsourceibias.n300 commonsourceibias.n299 13.0342
R23899 commonsourceibias.n343 commonsourceibias.n342 13.0342
R23900 commonsourceibias.n106 commonsourceibias.n105 13.0342
R23901 commonsourceibias.n63 commonsourceibias.n62 13.0342
R23902 commonsourceibias.n228 commonsourceibias.n227 13.0342
R23903 commonsourceibias.n185 commonsourceibias.n184 13.0342
R23904 commonsourceibias.n663 commonsourceibias.n662 13.0342
R23905 commonsourceibias.n709 commonsourceibias.n708 13.0342
R23906 commonsourceibias.n433 commonsourceibias.n432 13.0342
R23907 commonsourceibias.n479 commonsourceibias.n478 13.0342
R23908 commonsourceibias.n594 commonsourceibias.n593 13.0342
R23909 commonsourceibias.n549 commonsourceibias.n548 13.0342
R23910 commonsourceibias.n314 commonsourceibias.n313 12.5423
R23911 commonsourceibias.n329 commonsourceibias.n328 12.5423
R23912 commonsourceibias.n92 commonsourceibias.n91 12.5423
R23913 commonsourceibias.n77 commonsourceibias.n76 12.5423
R23914 commonsourceibias.n214 commonsourceibias.n213 12.5423
R23915 commonsourceibias.n198 commonsourceibias.n153 12.5423
R23916 commonsourceibias.n678 commonsourceibias.n677 12.5423
R23917 commonsourceibias.n694 commonsourceibias.n693 12.5423
R23918 commonsourceibias.n448 commonsourceibias.n447 12.5423
R23919 commonsourceibias.n464 commonsourceibias.n463 12.5423
R23920 commonsourceibias.n579 commonsourceibias.n578 12.5423
R23921 commonsourceibias.n562 commonsourceibias.n517 12.5423
R23922 commonsourceibias.n734 commonsourceibias.n366 12.2777
R23923 commonsourceibias.n315 commonsourceibias.n314 12.0505
R23924 commonsourceibias.n328 commonsourceibias.n327 12.0505
R23925 commonsourceibias.n91 commonsourceibias.n90 12.0505
R23926 commonsourceibias.n78 commonsourceibias.n77 12.0505
R23927 commonsourceibias.n213 commonsourceibias.n212 12.0505
R23928 commonsourceibias.n201 commonsourceibias.n153 12.0505
R23929 commonsourceibias.n679 commonsourceibias.n678 12.0505
R23930 commonsourceibias.n693 commonsourceibias.n692 12.0505
R23931 commonsourceibias.n449 commonsourceibias.n448 12.0505
R23932 commonsourceibias.n463 commonsourceibias.n462 12.0505
R23933 commonsourceibias.n578 commonsourceibias.n577 12.0505
R23934 commonsourceibias.n565 commonsourceibias.n517 12.0505
R23935 commonsourceibias.n301 commonsourceibias.n300 11.5587
R23936 commonsourceibias.n342 commonsourceibias.n341 11.5587
R23937 commonsourceibias.n105 commonsourceibias.n104 11.5587
R23938 commonsourceibias.n64 commonsourceibias.n63 11.5587
R23939 commonsourceibias.n227 commonsourceibias.n226 11.5587
R23940 commonsourceibias.n186 commonsourceibias.n185 11.5587
R23941 commonsourceibias.n664 commonsourceibias.n663 11.5587
R23942 commonsourceibias.n708 commonsourceibias.n707 11.5587
R23943 commonsourceibias.n434 commonsourceibias.n433 11.5587
R23944 commonsourceibias.n478 commonsourceibias.n477 11.5587
R23945 commonsourceibias.n593 commonsourceibias.n592 11.5587
R23946 commonsourceibias.n550 commonsourceibias.n549 11.5587
R23947 commonsourceibias.n287 commonsourceibias.n286 11.0668
R23948 commonsourceibias.n356 commonsourceibias.n355 11.0668
R23949 commonsourceibias.n119 commonsourceibias.n118 11.0668
R23950 commonsourceibias.n50 commonsourceibias.n49 11.0668
R23951 commonsourceibias.n241 commonsourceibias.n240 11.0668
R23952 commonsourceibias.n172 commonsourceibias.n171 11.0668
R23953 commonsourceibias.n649 commonsourceibias.n648 11.0668
R23954 commonsourceibias.n723 commonsourceibias.n722 11.0668
R23955 commonsourceibias.n419 commonsourceibias.n418 11.0668
R23956 commonsourceibias.n493 commonsourceibias.n492 11.0668
R23957 commonsourceibias.n608 commonsourceibias.n607 11.0668
R23958 commonsourceibias.n535 commonsourceibias.n534 11.0668
R23959 commonsourceibias.n734 commonsourceibias.n733 10.3347
R23960 commonsourceibias.n149 commonsourceibias.n148 9.50363
R23961 commonsourceibias.n514 commonsourceibias.n513 9.50363
R23962 commonsourceibias.n366 commonsourceibias.n250 8.75852
R23963 commonsourceibias.n733 commonsourceibias.n617 8.75852
R23964 commonsourceibias.n292 commonsourceibias.n291 5.16479
R23965 commonsourceibias.n256 commonsourceibias.n254 5.16479
R23966 commonsourceibias.n19 commonsourceibias.n17 5.16479
R23967 commonsourceibias.n55 commonsourceibias.n54 5.16479
R23968 commonsourceibias.n5 commonsourceibias.n3 5.16479
R23969 commonsourceibias.n177 commonsourceibias.n176 5.16479
R23970 commonsourceibias.n654 commonsourceibias.n653 5.16479
R23971 commonsourceibias.n716 commonsourceibias.n621 5.16479
R23972 commonsourceibias.n424 commonsourceibias.n423 5.16479
R23973 commonsourceibias.n486 commonsourceibias.n391 5.16479
R23974 commonsourceibias.n601 commonsourceibias.n370 5.16479
R23975 commonsourceibias.n540 commonsourceibias.n539 5.16479
R23976 commonsourceibias.n366 commonsourceibias.n365 5.03125
R23977 commonsourceibias.n733 commonsourceibias.n732 5.03125
R23978 commonsourceibias.n306 commonsourceibias.n305 4.67295
R23979 commonsourceibias.n261 commonsourceibias.n259 4.67295
R23980 commonsourceibias.n24 commonsourceibias.n22 4.67295
R23981 commonsourceibias.n69 commonsourceibias.n68 4.67295
R23982 commonsourceibias.n10 commonsourceibias.n8 4.67295
R23983 commonsourceibias.n191 commonsourceibias.n190 4.67295
R23984 commonsourceibias.n669 commonsourceibias.n668 4.67295
R23985 commonsourceibias.n701 commonsourceibias.n625 4.67295
R23986 commonsourceibias.n439 commonsourceibias.n438 4.67295
R23987 commonsourceibias.n471 commonsourceibias.n395 4.67295
R23988 commonsourceibias.n586 commonsourceibias.n374 4.67295
R23989 commonsourceibias.n555 commonsourceibias.n554 4.67295
R23990 commonsourceibias commonsourceibias.n734 4.20978
R23991 commonsourceibias.n320 commonsourceibias.n319 4.18111
R23992 commonsourceibias.n266 commonsourceibias.n264 4.18111
R23993 commonsourceibias.n29 commonsourceibias.n27 4.18111
R23994 commonsourceibias.n83 commonsourceibias.n82 4.18111
R23995 commonsourceibias.n150 commonsourceibias.n13 4.18111
R23996 commonsourceibias.n203 commonsourceibias.n151 4.18111
R23997 commonsourceibias.n684 commonsourceibias.n683 4.18111
R23998 commonsourceibias.n686 commonsourceibias.n629 4.18111
R23999 commonsourceibias.n454 commonsourceibias.n453 4.18111
R24000 commonsourceibias.n456 commonsourceibias.n399 4.18111
R24001 commonsourceibias.n571 commonsourceibias.n378 4.18111
R24002 commonsourceibias.n567 commonsourceibias.n515 4.18111
R24003 commonsourceibias.n271 commonsourceibias.n269 3.68928
R24004 commonsourceibias.n334 commonsourceibias.n333 3.68928
R24005 commonsourceibias.n97 commonsourceibias.n96 3.68928
R24006 commonsourceibias.n34 commonsourceibias.n32 3.68928
R24007 commonsourceibias.n219 commonsourceibias.n218 3.68928
R24008 commonsourceibias.n196 commonsourceibias.n155 3.68928
R24009 commonsourceibias.n671 commonsourceibias.n633 3.68928
R24010 commonsourceibias.n699 commonsourceibias.n698 3.68928
R24011 commonsourceibias.n441 commonsourceibias.n403 3.68928
R24012 commonsourceibias.n469 commonsourceibias.n468 3.68928
R24013 commonsourceibias.n584 commonsourceibias.n583 3.68928
R24014 commonsourceibias.n560 commonsourceibias.n519 3.68928
R24015 commonsourceibias.n276 commonsourceibias.n274 3.19744
R24016 commonsourceibias.n348 commonsourceibias.n347 3.19744
R24017 commonsourceibias.n111 commonsourceibias.n110 3.19744
R24018 commonsourceibias.n39 commonsourceibias.n37 3.19744
R24019 commonsourceibias.n233 commonsourceibias.n232 3.19744
R24020 commonsourceibias.n161 commonsourceibias.n159 3.19744
R24021 commonsourceibias.n656 commonsourceibias.n637 3.19744
R24022 commonsourceibias.n714 commonsourceibias.n713 3.19744
R24023 commonsourceibias.n426 commonsourceibias.n407 3.19744
R24024 commonsourceibias.n484 commonsourceibias.n483 3.19744
R24025 commonsourceibias.n599 commonsourceibias.n598 3.19744
R24026 commonsourceibias.n542 commonsourceibias.n523 3.19744
R24027 commonsourceibias.n139 commonsourceibias.t47 2.82907
R24028 commonsourceibias.n139 commonsourceibias.t79 2.82907
R24029 commonsourceibias.n140 commonsourceibias.t55 2.82907
R24030 commonsourceibias.n140 commonsourceibias.t5 2.82907
R24031 commonsourceibias.n142 commonsourceibias.t19 2.82907
R24032 commonsourceibias.n142 commonsourceibias.t23 2.82907
R24033 commonsourceibias.n144 commonsourceibias.t39 2.82907
R24034 commonsourceibias.n144 commonsourceibias.t71 2.82907
R24035 commonsourceibias.n146 commonsourceibias.t57 2.82907
R24036 commonsourceibias.n146 commonsourceibias.t27 2.82907
R24037 commonsourceibias.n137 commonsourceibias.t11 2.82907
R24038 commonsourceibias.n137 commonsourceibias.t41 2.82907
R24039 commonsourceibias.n135 commonsourceibias.t25 2.82907
R24040 commonsourceibias.n135 commonsourceibias.t35 2.82907
R24041 commonsourceibias.n133 commonsourceibias.t37 2.82907
R24042 commonsourceibias.n133 commonsourceibias.t77 2.82907
R24043 commonsourceibias.n131 commonsourceibias.t51 2.82907
R24044 commonsourceibias.n131 commonsourceibias.t9 2.82907
R24045 commonsourceibias.n129 commonsourceibias.t75 2.82907
R24046 commonsourceibias.n129 commonsourceibias.t21 2.82907
R24047 commonsourceibias.n503 commonsourceibias.t43 2.82907
R24048 commonsourceibias.n503 commonsourceibias.t15 2.82907
R24049 commonsourceibias.n505 commonsourceibias.t31 2.82907
R24050 commonsourceibias.n505 commonsourceibias.t1 2.82907
R24051 commonsourceibias.n507 commonsourceibias.t17 2.82907
R24052 commonsourceibias.n507 commonsourceibias.t61 2.82907
R24053 commonsourceibias.n509 commonsourceibias.t59 2.82907
R24054 commonsourceibias.n509 commonsourceibias.t45 2.82907
R24055 commonsourceibias.n511 commonsourceibias.t65 2.82907
R24056 commonsourceibias.n511 commonsourceibias.t33 2.82907
R24057 commonsourceibias.n386 commonsourceibias.t53 2.82907
R24058 commonsourceibias.n386 commonsourceibias.t73 2.82907
R24059 commonsourceibias.n384 commonsourceibias.t7 2.82907
R24060 commonsourceibias.n384 commonsourceibias.t63 2.82907
R24061 commonsourceibias.n382 commonsourceibias.t69 2.82907
R24062 commonsourceibias.n382 commonsourceibias.t67 2.82907
R24063 commonsourceibias.n380 commonsourceibias.t49 2.82907
R24064 commonsourceibias.n380 commonsourceibias.t13 2.82907
R24065 commonsourceibias.n379 commonsourceibias.t29 2.82907
R24066 commonsourceibias.n379 commonsourceibias.t3 2.82907
R24067 commonsourceibias.n280 commonsourceibias.n279 2.7056
R24068 commonsourceibias.n362 commonsourceibias.n361 2.7056
R24069 commonsourceibias.n125 commonsourceibias.n124 2.7056
R24070 commonsourceibias.n43 commonsourceibias.n42 2.7056
R24071 commonsourceibias.n247 commonsourceibias.n246 2.7056
R24072 commonsourceibias.n165 commonsourceibias.n164 2.7056
R24073 commonsourceibias.n642 commonsourceibias.n641 2.7056
R24074 commonsourceibias.n729 commonsourceibias.n728 2.7056
R24075 commonsourceibias.n412 commonsourceibias.n411 2.7056
R24076 commonsourceibias.n499 commonsourceibias.n498 2.7056
R24077 commonsourceibias.n614 commonsourceibias.n613 2.7056
R24078 commonsourceibias.n528 commonsourceibias.n527 2.7056
R24079 commonsourceibias.n132 commonsourceibias.n130 0.573776
R24080 commonsourceibias.n134 commonsourceibias.n132 0.573776
R24081 commonsourceibias.n136 commonsourceibias.n134 0.573776
R24082 commonsourceibias.n138 commonsourceibias.n136 0.573776
R24083 commonsourceibias.n147 commonsourceibias.n145 0.573776
R24084 commonsourceibias.n145 commonsourceibias.n143 0.573776
R24085 commonsourceibias.n143 commonsourceibias.n141 0.573776
R24086 commonsourceibias.n383 commonsourceibias.n381 0.573776
R24087 commonsourceibias.n385 commonsourceibias.n383 0.573776
R24088 commonsourceibias.n387 commonsourceibias.n385 0.573776
R24089 commonsourceibias.n512 commonsourceibias.n510 0.573776
R24090 commonsourceibias.n510 commonsourceibias.n508 0.573776
R24091 commonsourceibias.n508 commonsourceibias.n506 0.573776
R24092 commonsourceibias.n506 commonsourceibias.n504 0.573776
R24093 commonsourceibias.n148 commonsourceibias.n138 0.287138
R24094 commonsourceibias.n148 commonsourceibias.n147 0.287138
R24095 commonsourceibias.n513 commonsourceibias.n387 0.287138
R24096 commonsourceibias.n513 commonsourceibias.n512 0.287138
R24097 commonsourceibias.n365 commonsourceibias.n251 0.285035
R24098 commonsourceibias.n128 commonsourceibias.n14 0.285035
R24099 commonsourceibias.n250 commonsourceibias.n0 0.285035
R24100 commonsourceibias.n732 commonsourceibias.n618 0.285035
R24101 commonsourceibias.n502 commonsourceibias.n388 0.285035
R24102 commonsourceibias.n617 commonsourceibias.n367 0.285035
R24103 commonsourceibias.n360 commonsourceibias.n251 0.189894
R24104 commonsourceibias.n360 commonsourceibias.n359 0.189894
R24105 commonsourceibias.n359 commonsourceibias.n358 0.189894
R24106 commonsourceibias.n358 commonsourceibias.n253 0.189894
R24107 commonsourceibias.n353 commonsourceibias.n253 0.189894
R24108 commonsourceibias.n353 commonsourceibias.n352 0.189894
R24109 commonsourceibias.n352 commonsourceibias.n351 0.189894
R24110 commonsourceibias.n351 commonsourceibias.n255 0.189894
R24111 commonsourceibias.n346 commonsourceibias.n255 0.189894
R24112 commonsourceibias.n346 commonsourceibias.n345 0.189894
R24113 commonsourceibias.n345 commonsourceibias.n344 0.189894
R24114 commonsourceibias.n344 commonsourceibias.n258 0.189894
R24115 commonsourceibias.n339 commonsourceibias.n258 0.189894
R24116 commonsourceibias.n339 commonsourceibias.n338 0.189894
R24117 commonsourceibias.n338 commonsourceibias.n337 0.189894
R24118 commonsourceibias.n337 commonsourceibias.n260 0.189894
R24119 commonsourceibias.n332 commonsourceibias.n260 0.189894
R24120 commonsourceibias.n332 commonsourceibias.n331 0.189894
R24121 commonsourceibias.n331 commonsourceibias.n330 0.189894
R24122 commonsourceibias.n330 commonsourceibias.n263 0.189894
R24123 commonsourceibias.n325 commonsourceibias.n263 0.189894
R24124 commonsourceibias.n325 commonsourceibias.n324 0.189894
R24125 commonsourceibias.n324 commonsourceibias.n323 0.189894
R24126 commonsourceibias.n323 commonsourceibias.n265 0.189894
R24127 commonsourceibias.n318 commonsourceibias.n265 0.189894
R24128 commonsourceibias.n318 commonsourceibias.n317 0.189894
R24129 commonsourceibias.n317 commonsourceibias.n316 0.189894
R24130 commonsourceibias.n316 commonsourceibias.n268 0.189894
R24131 commonsourceibias.n311 commonsourceibias.n268 0.189894
R24132 commonsourceibias.n311 commonsourceibias.n310 0.189894
R24133 commonsourceibias.n310 commonsourceibias.n309 0.189894
R24134 commonsourceibias.n309 commonsourceibias.n270 0.189894
R24135 commonsourceibias.n304 commonsourceibias.n270 0.189894
R24136 commonsourceibias.n304 commonsourceibias.n303 0.189894
R24137 commonsourceibias.n303 commonsourceibias.n302 0.189894
R24138 commonsourceibias.n302 commonsourceibias.n273 0.189894
R24139 commonsourceibias.n297 commonsourceibias.n273 0.189894
R24140 commonsourceibias.n297 commonsourceibias.n296 0.189894
R24141 commonsourceibias.n296 commonsourceibias.n295 0.189894
R24142 commonsourceibias.n295 commonsourceibias.n275 0.189894
R24143 commonsourceibias.n290 commonsourceibias.n275 0.189894
R24144 commonsourceibias.n290 commonsourceibias.n289 0.189894
R24145 commonsourceibias.n289 commonsourceibias.n288 0.189894
R24146 commonsourceibias.n288 commonsourceibias.n278 0.189894
R24147 commonsourceibias.n283 commonsourceibias.n278 0.189894
R24148 commonsourceibias.n283 commonsourceibias.n282 0.189894
R24149 commonsourceibias.n123 commonsourceibias.n14 0.189894
R24150 commonsourceibias.n123 commonsourceibias.n122 0.189894
R24151 commonsourceibias.n122 commonsourceibias.n121 0.189894
R24152 commonsourceibias.n121 commonsourceibias.n16 0.189894
R24153 commonsourceibias.n116 commonsourceibias.n16 0.189894
R24154 commonsourceibias.n116 commonsourceibias.n115 0.189894
R24155 commonsourceibias.n115 commonsourceibias.n114 0.189894
R24156 commonsourceibias.n114 commonsourceibias.n18 0.189894
R24157 commonsourceibias.n109 commonsourceibias.n18 0.189894
R24158 commonsourceibias.n109 commonsourceibias.n108 0.189894
R24159 commonsourceibias.n108 commonsourceibias.n107 0.189894
R24160 commonsourceibias.n107 commonsourceibias.n21 0.189894
R24161 commonsourceibias.n102 commonsourceibias.n21 0.189894
R24162 commonsourceibias.n102 commonsourceibias.n101 0.189894
R24163 commonsourceibias.n101 commonsourceibias.n100 0.189894
R24164 commonsourceibias.n100 commonsourceibias.n23 0.189894
R24165 commonsourceibias.n95 commonsourceibias.n23 0.189894
R24166 commonsourceibias.n95 commonsourceibias.n94 0.189894
R24167 commonsourceibias.n94 commonsourceibias.n93 0.189894
R24168 commonsourceibias.n93 commonsourceibias.n26 0.189894
R24169 commonsourceibias.n88 commonsourceibias.n26 0.189894
R24170 commonsourceibias.n88 commonsourceibias.n87 0.189894
R24171 commonsourceibias.n87 commonsourceibias.n86 0.189894
R24172 commonsourceibias.n86 commonsourceibias.n28 0.189894
R24173 commonsourceibias.n81 commonsourceibias.n28 0.189894
R24174 commonsourceibias.n81 commonsourceibias.n80 0.189894
R24175 commonsourceibias.n80 commonsourceibias.n79 0.189894
R24176 commonsourceibias.n79 commonsourceibias.n31 0.189894
R24177 commonsourceibias.n74 commonsourceibias.n31 0.189894
R24178 commonsourceibias.n74 commonsourceibias.n73 0.189894
R24179 commonsourceibias.n73 commonsourceibias.n72 0.189894
R24180 commonsourceibias.n72 commonsourceibias.n33 0.189894
R24181 commonsourceibias.n67 commonsourceibias.n33 0.189894
R24182 commonsourceibias.n67 commonsourceibias.n66 0.189894
R24183 commonsourceibias.n66 commonsourceibias.n65 0.189894
R24184 commonsourceibias.n65 commonsourceibias.n36 0.189894
R24185 commonsourceibias.n60 commonsourceibias.n36 0.189894
R24186 commonsourceibias.n60 commonsourceibias.n59 0.189894
R24187 commonsourceibias.n59 commonsourceibias.n58 0.189894
R24188 commonsourceibias.n58 commonsourceibias.n38 0.189894
R24189 commonsourceibias.n53 commonsourceibias.n38 0.189894
R24190 commonsourceibias.n53 commonsourceibias.n52 0.189894
R24191 commonsourceibias.n52 commonsourceibias.n51 0.189894
R24192 commonsourceibias.n51 commonsourceibias.n41 0.189894
R24193 commonsourceibias.n46 commonsourceibias.n41 0.189894
R24194 commonsourceibias.n46 commonsourceibias.n45 0.189894
R24195 commonsourceibias.n205 commonsourceibias.n204 0.189894
R24196 commonsourceibias.n204 commonsourceibias.n152 0.189894
R24197 commonsourceibias.n200 commonsourceibias.n152 0.189894
R24198 commonsourceibias.n200 commonsourceibias.n199 0.189894
R24199 commonsourceibias.n199 commonsourceibias.n154 0.189894
R24200 commonsourceibias.n195 commonsourceibias.n154 0.189894
R24201 commonsourceibias.n195 commonsourceibias.n194 0.189894
R24202 commonsourceibias.n194 commonsourceibias.n156 0.189894
R24203 commonsourceibias.n189 commonsourceibias.n156 0.189894
R24204 commonsourceibias.n189 commonsourceibias.n188 0.189894
R24205 commonsourceibias.n188 commonsourceibias.n187 0.189894
R24206 commonsourceibias.n187 commonsourceibias.n158 0.189894
R24207 commonsourceibias.n182 commonsourceibias.n158 0.189894
R24208 commonsourceibias.n182 commonsourceibias.n181 0.189894
R24209 commonsourceibias.n181 commonsourceibias.n180 0.189894
R24210 commonsourceibias.n180 commonsourceibias.n160 0.189894
R24211 commonsourceibias.n175 commonsourceibias.n160 0.189894
R24212 commonsourceibias.n175 commonsourceibias.n174 0.189894
R24213 commonsourceibias.n174 commonsourceibias.n173 0.189894
R24214 commonsourceibias.n173 commonsourceibias.n163 0.189894
R24215 commonsourceibias.n168 commonsourceibias.n163 0.189894
R24216 commonsourceibias.n168 commonsourceibias.n167 0.189894
R24217 commonsourceibias.n245 commonsourceibias.n0 0.189894
R24218 commonsourceibias.n245 commonsourceibias.n244 0.189894
R24219 commonsourceibias.n244 commonsourceibias.n243 0.189894
R24220 commonsourceibias.n243 commonsourceibias.n2 0.189894
R24221 commonsourceibias.n238 commonsourceibias.n2 0.189894
R24222 commonsourceibias.n238 commonsourceibias.n237 0.189894
R24223 commonsourceibias.n237 commonsourceibias.n236 0.189894
R24224 commonsourceibias.n236 commonsourceibias.n4 0.189894
R24225 commonsourceibias.n231 commonsourceibias.n4 0.189894
R24226 commonsourceibias.n231 commonsourceibias.n230 0.189894
R24227 commonsourceibias.n230 commonsourceibias.n229 0.189894
R24228 commonsourceibias.n229 commonsourceibias.n7 0.189894
R24229 commonsourceibias.n224 commonsourceibias.n7 0.189894
R24230 commonsourceibias.n224 commonsourceibias.n223 0.189894
R24231 commonsourceibias.n223 commonsourceibias.n222 0.189894
R24232 commonsourceibias.n222 commonsourceibias.n9 0.189894
R24233 commonsourceibias.n217 commonsourceibias.n9 0.189894
R24234 commonsourceibias.n217 commonsourceibias.n216 0.189894
R24235 commonsourceibias.n216 commonsourceibias.n215 0.189894
R24236 commonsourceibias.n215 commonsourceibias.n12 0.189894
R24237 commonsourceibias.n210 commonsourceibias.n12 0.189894
R24238 commonsourceibias.n210 commonsourceibias.n209 0.189894
R24239 commonsourceibias.n209 commonsourceibias.n208 0.189894
R24240 commonsourceibias.n645 commonsourceibias.n644 0.189894
R24241 commonsourceibias.n645 commonsourceibias.n640 0.189894
R24242 commonsourceibias.n650 commonsourceibias.n640 0.189894
R24243 commonsourceibias.n651 commonsourceibias.n650 0.189894
R24244 commonsourceibias.n652 commonsourceibias.n651 0.189894
R24245 commonsourceibias.n652 commonsourceibias.n638 0.189894
R24246 commonsourceibias.n658 commonsourceibias.n638 0.189894
R24247 commonsourceibias.n659 commonsourceibias.n658 0.189894
R24248 commonsourceibias.n660 commonsourceibias.n659 0.189894
R24249 commonsourceibias.n660 commonsourceibias.n636 0.189894
R24250 commonsourceibias.n665 commonsourceibias.n636 0.189894
R24251 commonsourceibias.n666 commonsourceibias.n665 0.189894
R24252 commonsourceibias.n667 commonsourceibias.n666 0.189894
R24253 commonsourceibias.n667 commonsourceibias.n634 0.189894
R24254 commonsourceibias.n673 commonsourceibias.n634 0.189894
R24255 commonsourceibias.n674 commonsourceibias.n673 0.189894
R24256 commonsourceibias.n675 commonsourceibias.n674 0.189894
R24257 commonsourceibias.n675 commonsourceibias.n632 0.189894
R24258 commonsourceibias.n680 commonsourceibias.n632 0.189894
R24259 commonsourceibias.n681 commonsourceibias.n680 0.189894
R24260 commonsourceibias.n682 commonsourceibias.n681 0.189894
R24261 commonsourceibias.n682 commonsourceibias.n630 0.189894
R24262 commonsourceibias.n688 commonsourceibias.n630 0.189894
R24263 commonsourceibias.n689 commonsourceibias.n688 0.189894
R24264 commonsourceibias.n690 commonsourceibias.n689 0.189894
R24265 commonsourceibias.n690 commonsourceibias.n628 0.189894
R24266 commonsourceibias.n695 commonsourceibias.n628 0.189894
R24267 commonsourceibias.n696 commonsourceibias.n695 0.189894
R24268 commonsourceibias.n697 commonsourceibias.n696 0.189894
R24269 commonsourceibias.n697 commonsourceibias.n626 0.189894
R24270 commonsourceibias.n703 commonsourceibias.n626 0.189894
R24271 commonsourceibias.n704 commonsourceibias.n703 0.189894
R24272 commonsourceibias.n705 commonsourceibias.n704 0.189894
R24273 commonsourceibias.n705 commonsourceibias.n624 0.189894
R24274 commonsourceibias.n710 commonsourceibias.n624 0.189894
R24275 commonsourceibias.n711 commonsourceibias.n710 0.189894
R24276 commonsourceibias.n712 commonsourceibias.n711 0.189894
R24277 commonsourceibias.n712 commonsourceibias.n622 0.189894
R24278 commonsourceibias.n718 commonsourceibias.n622 0.189894
R24279 commonsourceibias.n719 commonsourceibias.n718 0.189894
R24280 commonsourceibias.n720 commonsourceibias.n719 0.189894
R24281 commonsourceibias.n720 commonsourceibias.n620 0.189894
R24282 commonsourceibias.n725 commonsourceibias.n620 0.189894
R24283 commonsourceibias.n726 commonsourceibias.n725 0.189894
R24284 commonsourceibias.n727 commonsourceibias.n726 0.189894
R24285 commonsourceibias.n727 commonsourceibias.n618 0.189894
R24286 commonsourceibias.n415 commonsourceibias.n414 0.189894
R24287 commonsourceibias.n415 commonsourceibias.n410 0.189894
R24288 commonsourceibias.n420 commonsourceibias.n410 0.189894
R24289 commonsourceibias.n421 commonsourceibias.n420 0.189894
R24290 commonsourceibias.n422 commonsourceibias.n421 0.189894
R24291 commonsourceibias.n422 commonsourceibias.n408 0.189894
R24292 commonsourceibias.n428 commonsourceibias.n408 0.189894
R24293 commonsourceibias.n429 commonsourceibias.n428 0.189894
R24294 commonsourceibias.n430 commonsourceibias.n429 0.189894
R24295 commonsourceibias.n430 commonsourceibias.n406 0.189894
R24296 commonsourceibias.n435 commonsourceibias.n406 0.189894
R24297 commonsourceibias.n436 commonsourceibias.n435 0.189894
R24298 commonsourceibias.n437 commonsourceibias.n436 0.189894
R24299 commonsourceibias.n437 commonsourceibias.n404 0.189894
R24300 commonsourceibias.n443 commonsourceibias.n404 0.189894
R24301 commonsourceibias.n444 commonsourceibias.n443 0.189894
R24302 commonsourceibias.n445 commonsourceibias.n444 0.189894
R24303 commonsourceibias.n445 commonsourceibias.n402 0.189894
R24304 commonsourceibias.n450 commonsourceibias.n402 0.189894
R24305 commonsourceibias.n451 commonsourceibias.n450 0.189894
R24306 commonsourceibias.n452 commonsourceibias.n451 0.189894
R24307 commonsourceibias.n452 commonsourceibias.n400 0.189894
R24308 commonsourceibias.n458 commonsourceibias.n400 0.189894
R24309 commonsourceibias.n459 commonsourceibias.n458 0.189894
R24310 commonsourceibias.n460 commonsourceibias.n459 0.189894
R24311 commonsourceibias.n460 commonsourceibias.n398 0.189894
R24312 commonsourceibias.n465 commonsourceibias.n398 0.189894
R24313 commonsourceibias.n466 commonsourceibias.n465 0.189894
R24314 commonsourceibias.n467 commonsourceibias.n466 0.189894
R24315 commonsourceibias.n467 commonsourceibias.n396 0.189894
R24316 commonsourceibias.n473 commonsourceibias.n396 0.189894
R24317 commonsourceibias.n474 commonsourceibias.n473 0.189894
R24318 commonsourceibias.n475 commonsourceibias.n474 0.189894
R24319 commonsourceibias.n475 commonsourceibias.n394 0.189894
R24320 commonsourceibias.n480 commonsourceibias.n394 0.189894
R24321 commonsourceibias.n481 commonsourceibias.n480 0.189894
R24322 commonsourceibias.n482 commonsourceibias.n481 0.189894
R24323 commonsourceibias.n482 commonsourceibias.n392 0.189894
R24324 commonsourceibias.n488 commonsourceibias.n392 0.189894
R24325 commonsourceibias.n489 commonsourceibias.n488 0.189894
R24326 commonsourceibias.n490 commonsourceibias.n489 0.189894
R24327 commonsourceibias.n490 commonsourceibias.n390 0.189894
R24328 commonsourceibias.n495 commonsourceibias.n390 0.189894
R24329 commonsourceibias.n496 commonsourceibias.n495 0.189894
R24330 commonsourceibias.n497 commonsourceibias.n496 0.189894
R24331 commonsourceibias.n497 commonsourceibias.n388 0.189894
R24332 commonsourceibias.n531 commonsourceibias.n530 0.189894
R24333 commonsourceibias.n531 commonsourceibias.n526 0.189894
R24334 commonsourceibias.n536 commonsourceibias.n526 0.189894
R24335 commonsourceibias.n537 commonsourceibias.n536 0.189894
R24336 commonsourceibias.n538 commonsourceibias.n537 0.189894
R24337 commonsourceibias.n538 commonsourceibias.n524 0.189894
R24338 commonsourceibias.n544 commonsourceibias.n524 0.189894
R24339 commonsourceibias.n545 commonsourceibias.n544 0.189894
R24340 commonsourceibias.n546 commonsourceibias.n545 0.189894
R24341 commonsourceibias.n546 commonsourceibias.n522 0.189894
R24342 commonsourceibias.n551 commonsourceibias.n522 0.189894
R24343 commonsourceibias.n552 commonsourceibias.n551 0.189894
R24344 commonsourceibias.n553 commonsourceibias.n552 0.189894
R24345 commonsourceibias.n553 commonsourceibias.n520 0.189894
R24346 commonsourceibias.n558 commonsourceibias.n520 0.189894
R24347 commonsourceibias.n559 commonsourceibias.n558 0.189894
R24348 commonsourceibias.n559 commonsourceibias.n518 0.189894
R24349 commonsourceibias.n563 commonsourceibias.n518 0.189894
R24350 commonsourceibias.n564 commonsourceibias.n563 0.189894
R24351 commonsourceibias.n564 commonsourceibias.n516 0.189894
R24352 commonsourceibias.n568 commonsourceibias.n516 0.189894
R24353 commonsourceibias.n569 commonsourceibias.n568 0.189894
R24354 commonsourceibias.n574 commonsourceibias.n573 0.189894
R24355 commonsourceibias.n575 commonsourceibias.n574 0.189894
R24356 commonsourceibias.n575 commonsourceibias.n377 0.189894
R24357 commonsourceibias.n580 commonsourceibias.n377 0.189894
R24358 commonsourceibias.n581 commonsourceibias.n580 0.189894
R24359 commonsourceibias.n582 commonsourceibias.n581 0.189894
R24360 commonsourceibias.n582 commonsourceibias.n375 0.189894
R24361 commonsourceibias.n588 commonsourceibias.n375 0.189894
R24362 commonsourceibias.n589 commonsourceibias.n588 0.189894
R24363 commonsourceibias.n590 commonsourceibias.n589 0.189894
R24364 commonsourceibias.n590 commonsourceibias.n373 0.189894
R24365 commonsourceibias.n595 commonsourceibias.n373 0.189894
R24366 commonsourceibias.n596 commonsourceibias.n595 0.189894
R24367 commonsourceibias.n597 commonsourceibias.n596 0.189894
R24368 commonsourceibias.n597 commonsourceibias.n371 0.189894
R24369 commonsourceibias.n603 commonsourceibias.n371 0.189894
R24370 commonsourceibias.n604 commonsourceibias.n603 0.189894
R24371 commonsourceibias.n605 commonsourceibias.n604 0.189894
R24372 commonsourceibias.n605 commonsourceibias.n369 0.189894
R24373 commonsourceibias.n610 commonsourceibias.n369 0.189894
R24374 commonsourceibias.n611 commonsourceibias.n610 0.189894
R24375 commonsourceibias.n612 commonsourceibias.n611 0.189894
R24376 commonsourceibias.n612 commonsourceibias.n367 0.189894
R24377 commonsourceibias.n205 commonsourceibias.n149 0.0762576
R24378 commonsourceibias.n208 commonsourceibias.n149 0.0762576
R24379 commonsourceibias.n569 commonsourceibias.n514 0.0762576
R24380 commonsourceibias.n573 commonsourceibias.n514 0.0762576
R24381 a_n2650_8322.n10 a_n2650_8322.t29 74.6477
R24382 a_n2650_8322.n1 a_n2650_8322.t21 74.6477
R24383 a_n2650_8322.n24 a_n2650_8322.t23 74.6474
R24384 a_n2650_8322.n18 a_n2650_8322.t20 74.2899
R24385 a_n2650_8322.n11 a_n2650_8322.t27 74.2899
R24386 a_n2650_8322.n12 a_n2650_8322.t30 74.2899
R24387 a_n2650_8322.n15 a_n2650_8322.t31 74.2899
R24388 a_n2650_8322.n8 a_n2650_8322.t6 74.2899
R24389 a_n2650_8322.n24 a_n2650_8322.n23 70.6783
R24390 a_n2650_8322.n22 a_n2650_8322.n21 70.6783
R24391 a_n2650_8322.n20 a_n2650_8322.n19 70.6783
R24392 a_n2650_8322.n10 a_n2650_8322.n9 70.6783
R24393 a_n2650_8322.n14 a_n2650_8322.n13 70.6783
R24394 a_n2650_8322.n1 a_n2650_8322.n0 70.6783
R24395 a_n2650_8322.n3 a_n2650_8322.n2 70.6783
R24396 a_n2650_8322.n5 a_n2650_8322.n4 70.6783
R24397 a_n2650_8322.n7 a_n2650_8322.n6 70.6783
R24398 a_n2650_8322.n26 a_n2650_8322.n25 70.6782
R24399 a_n2650_8322.n16 a_n2650_8322.n8 24.1867
R24400 a_n2650_8322.n17 a_n2650_8322.t0 10.0676
R24401 a_n2650_8322.n16 a_n2650_8322.n15 7.67184
R24402 a_n2650_8322.n18 a_n2650_8322.n17 6.55222
R24403 a_n2650_8322.n17 a_n2650_8322.n16 5.3452
R24404 a_n2650_8322.n23 a_n2650_8322.t18 3.61217
R24405 a_n2650_8322.n23 a_n2650_8322.t14 3.61217
R24406 a_n2650_8322.n21 a_n2650_8322.t22 3.61217
R24407 a_n2650_8322.n21 a_n2650_8322.t12 3.61217
R24408 a_n2650_8322.n19 a_n2650_8322.t10 3.61217
R24409 a_n2650_8322.n19 a_n2650_8322.t9 3.61217
R24410 a_n2650_8322.n9 a_n2650_8322.t33 3.61217
R24411 a_n2650_8322.n9 a_n2650_8322.t32 3.61217
R24412 a_n2650_8322.n13 a_n2650_8322.t28 3.61217
R24413 a_n2650_8322.n13 a_n2650_8322.t26 3.61217
R24414 a_n2650_8322.n0 a_n2650_8322.t24 3.61217
R24415 a_n2650_8322.n0 a_n2650_8322.t16 3.61217
R24416 a_n2650_8322.n2 a_n2650_8322.t8 3.61217
R24417 a_n2650_8322.n2 a_n2650_8322.t7 3.61217
R24418 a_n2650_8322.n4 a_n2650_8322.t19 3.61217
R24419 a_n2650_8322.n4 a_n2650_8322.t13 3.61217
R24420 a_n2650_8322.n6 a_n2650_8322.t17 3.61217
R24421 a_n2650_8322.n6 a_n2650_8322.t15 3.61217
R24422 a_n2650_8322.n26 a_n2650_8322.t11 3.61217
R24423 a_n2650_8322.t25 a_n2650_8322.n26 3.61217
R24424 a_n2650_8322.n15 a_n2650_8322.n14 0.358259
R24425 a_n2650_8322.n14 a_n2650_8322.n12 0.358259
R24426 a_n2650_8322.n11 a_n2650_8322.n10 0.358259
R24427 a_n2650_8322.n8 a_n2650_8322.n7 0.358259
R24428 a_n2650_8322.n7 a_n2650_8322.n5 0.358259
R24429 a_n2650_8322.n5 a_n2650_8322.n3 0.358259
R24430 a_n2650_8322.n3 a_n2650_8322.n1 0.358259
R24431 a_n2650_8322.n20 a_n2650_8322.n18 0.358259
R24432 a_n2650_8322.n22 a_n2650_8322.n20 0.358259
R24433 a_n2650_8322.n25 a_n2650_8322.n22 0.358259
R24434 a_n2650_8322.n25 a_n2650_8322.n24 0.358259
R24435 a_n2650_8322.n12 a_n2650_8322.n11 0.101793
R24436 a_n2650_8322.t5 a_n2650_8322.t2 0.0788333
R24437 a_n2650_8322.t4 a_n2650_8322.t3 0.0788333
R24438 a_n2650_8322.t0 a_n2650_8322.t1 0.0788333
R24439 a_n2650_8322.t4 a_n2650_8322.t5 0.0318333
R24440 a_n2650_8322.t0 a_n2650_8322.t3 0.0318333
R24441 a_n2650_8322.t2 a_n2650_8322.t3 0.0318333
R24442 a_n2650_8322.t1 a_n2650_8322.t4 0.0318333
R24443 output.n41 output.n15 289.615
R24444 output.n72 output.n46 289.615
R24445 output.n104 output.n78 289.615
R24446 output.n136 output.n110 289.615
R24447 output.n77 output.n45 197.26
R24448 output.n77 output.n76 196.298
R24449 output.n109 output.n108 196.298
R24450 output.n141 output.n140 196.298
R24451 output.n42 output.n41 185
R24452 output.n40 output.n39 185
R24453 output.n19 output.n18 185
R24454 output.n34 output.n33 185
R24455 output.n32 output.n31 185
R24456 output.n23 output.n22 185
R24457 output.n26 output.n25 185
R24458 output.n73 output.n72 185
R24459 output.n71 output.n70 185
R24460 output.n50 output.n49 185
R24461 output.n65 output.n64 185
R24462 output.n63 output.n62 185
R24463 output.n54 output.n53 185
R24464 output.n57 output.n56 185
R24465 output.n105 output.n104 185
R24466 output.n103 output.n102 185
R24467 output.n82 output.n81 185
R24468 output.n97 output.n96 185
R24469 output.n95 output.n94 185
R24470 output.n86 output.n85 185
R24471 output.n89 output.n88 185
R24472 output.n137 output.n136 185
R24473 output.n135 output.n134 185
R24474 output.n114 output.n113 185
R24475 output.n129 output.n128 185
R24476 output.n127 output.n126 185
R24477 output.n118 output.n117 185
R24478 output.n121 output.n120 185
R24479 output.t19 output.n24 147.661
R24480 output.t17 output.n55 147.661
R24481 output.t18 output.n87 147.661
R24482 output.t16 output.n119 147.661
R24483 output.n41 output.n40 104.615
R24484 output.n40 output.n18 104.615
R24485 output.n33 output.n18 104.615
R24486 output.n33 output.n32 104.615
R24487 output.n32 output.n22 104.615
R24488 output.n25 output.n22 104.615
R24489 output.n72 output.n71 104.615
R24490 output.n71 output.n49 104.615
R24491 output.n64 output.n49 104.615
R24492 output.n64 output.n63 104.615
R24493 output.n63 output.n53 104.615
R24494 output.n56 output.n53 104.615
R24495 output.n104 output.n103 104.615
R24496 output.n103 output.n81 104.615
R24497 output.n96 output.n81 104.615
R24498 output.n96 output.n95 104.615
R24499 output.n95 output.n85 104.615
R24500 output.n88 output.n85 104.615
R24501 output.n136 output.n135 104.615
R24502 output.n135 output.n113 104.615
R24503 output.n128 output.n113 104.615
R24504 output.n128 output.n127 104.615
R24505 output.n127 output.n117 104.615
R24506 output.n120 output.n117 104.615
R24507 output.n1 output.t9 77.056
R24508 output.n14 output.t11 76.6694
R24509 output.n1 output.n0 72.7095
R24510 output.n3 output.n2 72.7095
R24511 output.n5 output.n4 72.7095
R24512 output.n7 output.n6 72.7095
R24513 output.n9 output.n8 72.7095
R24514 output.n11 output.n10 72.7095
R24515 output.n13 output.n12 72.7095
R24516 output.n25 output.t19 52.3082
R24517 output.n56 output.t17 52.3082
R24518 output.n88 output.t18 52.3082
R24519 output.n120 output.t16 52.3082
R24520 output.n26 output.n24 15.6674
R24521 output.n57 output.n55 15.6674
R24522 output.n89 output.n87 15.6674
R24523 output.n121 output.n119 15.6674
R24524 output.n27 output.n23 12.8005
R24525 output.n58 output.n54 12.8005
R24526 output.n90 output.n86 12.8005
R24527 output.n122 output.n118 12.8005
R24528 output.n31 output.n30 12.0247
R24529 output.n62 output.n61 12.0247
R24530 output.n94 output.n93 12.0247
R24531 output.n126 output.n125 12.0247
R24532 output.n34 output.n21 11.249
R24533 output.n65 output.n52 11.249
R24534 output.n97 output.n84 11.249
R24535 output.n129 output.n116 11.249
R24536 output.n35 output.n19 10.4732
R24537 output.n66 output.n50 10.4732
R24538 output.n98 output.n82 10.4732
R24539 output.n130 output.n114 10.4732
R24540 output.n39 output.n38 9.69747
R24541 output.n70 output.n69 9.69747
R24542 output.n102 output.n101 9.69747
R24543 output.n134 output.n133 9.69747
R24544 output.n45 output.n44 9.45567
R24545 output.n76 output.n75 9.45567
R24546 output.n108 output.n107 9.45567
R24547 output.n140 output.n139 9.45567
R24548 output.n44 output.n43 9.3005
R24549 output.n17 output.n16 9.3005
R24550 output.n38 output.n37 9.3005
R24551 output.n36 output.n35 9.3005
R24552 output.n21 output.n20 9.3005
R24553 output.n30 output.n29 9.3005
R24554 output.n28 output.n27 9.3005
R24555 output.n75 output.n74 9.3005
R24556 output.n48 output.n47 9.3005
R24557 output.n69 output.n68 9.3005
R24558 output.n67 output.n66 9.3005
R24559 output.n52 output.n51 9.3005
R24560 output.n61 output.n60 9.3005
R24561 output.n59 output.n58 9.3005
R24562 output.n107 output.n106 9.3005
R24563 output.n80 output.n79 9.3005
R24564 output.n101 output.n100 9.3005
R24565 output.n99 output.n98 9.3005
R24566 output.n84 output.n83 9.3005
R24567 output.n93 output.n92 9.3005
R24568 output.n91 output.n90 9.3005
R24569 output.n139 output.n138 9.3005
R24570 output.n112 output.n111 9.3005
R24571 output.n133 output.n132 9.3005
R24572 output.n131 output.n130 9.3005
R24573 output.n116 output.n115 9.3005
R24574 output.n125 output.n124 9.3005
R24575 output.n123 output.n122 9.3005
R24576 output.n42 output.n17 8.92171
R24577 output.n73 output.n48 8.92171
R24578 output.n105 output.n80 8.92171
R24579 output.n137 output.n112 8.92171
R24580 output output.n141 8.15037
R24581 output.n43 output.n15 8.14595
R24582 output.n74 output.n46 8.14595
R24583 output.n106 output.n78 8.14595
R24584 output.n138 output.n110 8.14595
R24585 output.n45 output.n15 5.81868
R24586 output.n76 output.n46 5.81868
R24587 output.n108 output.n78 5.81868
R24588 output.n140 output.n110 5.81868
R24589 output.n43 output.n42 5.04292
R24590 output.n74 output.n73 5.04292
R24591 output.n106 output.n105 5.04292
R24592 output.n138 output.n137 5.04292
R24593 output.n28 output.n24 4.38594
R24594 output.n59 output.n55 4.38594
R24595 output.n91 output.n87 4.38594
R24596 output.n123 output.n119 4.38594
R24597 output.n39 output.n17 4.26717
R24598 output.n70 output.n48 4.26717
R24599 output.n102 output.n80 4.26717
R24600 output.n134 output.n112 4.26717
R24601 output.n0 output.t15 3.9605
R24602 output.n0 output.t4 3.9605
R24603 output.n2 output.t8 3.9605
R24604 output.n2 output.t0 3.9605
R24605 output.n4 output.t2 3.9605
R24606 output.n4 output.t1 3.9605
R24607 output.n6 output.t7 3.9605
R24608 output.n6 output.t10 3.9605
R24609 output.n8 output.t12 3.9605
R24610 output.n8 output.t5 3.9605
R24611 output.n10 output.t6 3.9605
R24612 output.n10 output.t13 3.9605
R24613 output.n12 output.t14 3.9605
R24614 output.n12 output.t3 3.9605
R24615 output.n38 output.n19 3.49141
R24616 output.n69 output.n50 3.49141
R24617 output.n101 output.n82 3.49141
R24618 output.n133 output.n114 3.49141
R24619 output.n35 output.n34 2.71565
R24620 output.n66 output.n65 2.71565
R24621 output.n98 output.n97 2.71565
R24622 output.n130 output.n129 2.71565
R24623 output.n31 output.n21 1.93989
R24624 output.n62 output.n52 1.93989
R24625 output.n94 output.n84 1.93989
R24626 output.n126 output.n116 1.93989
R24627 output.n30 output.n23 1.16414
R24628 output.n61 output.n54 1.16414
R24629 output.n93 output.n86 1.16414
R24630 output.n125 output.n118 1.16414
R24631 output.n141 output.n109 0.962709
R24632 output.n109 output.n77 0.962709
R24633 output.n27 output.n26 0.388379
R24634 output.n58 output.n57 0.388379
R24635 output.n90 output.n89 0.388379
R24636 output.n122 output.n121 0.388379
R24637 output.n14 output.n13 0.387128
R24638 output.n13 output.n11 0.387128
R24639 output.n11 output.n9 0.387128
R24640 output.n9 output.n7 0.387128
R24641 output.n7 output.n5 0.387128
R24642 output.n5 output.n3 0.387128
R24643 output.n3 output.n1 0.387128
R24644 output.n44 output.n16 0.155672
R24645 output.n37 output.n16 0.155672
R24646 output.n37 output.n36 0.155672
R24647 output.n36 output.n20 0.155672
R24648 output.n29 output.n20 0.155672
R24649 output.n29 output.n28 0.155672
R24650 output.n75 output.n47 0.155672
R24651 output.n68 output.n47 0.155672
R24652 output.n68 output.n67 0.155672
R24653 output.n67 output.n51 0.155672
R24654 output.n60 output.n51 0.155672
R24655 output.n60 output.n59 0.155672
R24656 output.n107 output.n79 0.155672
R24657 output.n100 output.n79 0.155672
R24658 output.n100 output.n99 0.155672
R24659 output.n99 output.n83 0.155672
R24660 output.n92 output.n83 0.155672
R24661 output.n92 output.n91 0.155672
R24662 output.n139 output.n111 0.155672
R24663 output.n132 output.n111 0.155672
R24664 output.n132 output.n131 0.155672
R24665 output.n131 output.n115 0.155672
R24666 output.n124 output.n115 0.155672
R24667 output.n124 output.n123 0.155672
R24668 output output.n14 0.126227
C0 output outputibias 2.34152f
C1 vdd output 7.23429f
C2 CSoutput output 6.13571f
C3 CSoutput outputibias 0.032386f
C4 vdd CSoutput 0.116919p
C5 minus diffpairibias 4.33e-19
C6 commonsourceibias output 0.006808f
C7 CSoutput minus 3.17016f
C8 vdd plus 0.091781f
C9 commonsourceibias outputibias 0.003832f
C10 plus diffpairibias 4.56e-19
C11 vdd commonsourceibias 0.004218f
C12 CSoutput plus 0.91196f
C13 commonsourceibias diffpairibias 0.052527f
C14 CSoutput commonsourceibias 45.462303f
C15 minus plus 10.303599f
C16 minus commonsourceibias 0.337549f
C17 plus commonsourceibias 0.283677f
C18 diffpairibias gnd 59.99123f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.181996p
C22 plus gnd 37.7259f
C23 minus gnd 31.29437f
C24 CSoutput gnd 0.115456p
C25 vdd gnd 0.478096p
C26 output.t9 gnd 0.464308f
C27 output.t15 gnd 0.044422f
C28 output.t4 gnd 0.044422f
C29 output.n0 gnd 0.364624f
C30 output.n1 gnd 0.614102f
C31 output.t8 gnd 0.044422f
C32 output.t0 gnd 0.044422f
C33 output.n2 gnd 0.364624f
C34 output.n3 gnd 0.350265f
C35 output.t2 gnd 0.044422f
C36 output.t1 gnd 0.044422f
C37 output.n4 gnd 0.364624f
C38 output.n5 gnd 0.350265f
C39 output.t7 gnd 0.044422f
C40 output.t10 gnd 0.044422f
C41 output.n6 gnd 0.364624f
C42 output.n7 gnd 0.350265f
C43 output.t12 gnd 0.044422f
C44 output.t5 gnd 0.044422f
C45 output.n8 gnd 0.364624f
C46 output.n9 gnd 0.350265f
C47 output.t6 gnd 0.044422f
C48 output.t13 gnd 0.044422f
C49 output.n10 gnd 0.364624f
C50 output.n11 gnd 0.350265f
C51 output.t14 gnd 0.044422f
C52 output.t3 gnd 0.044422f
C53 output.n12 gnd 0.364624f
C54 output.n13 gnd 0.350265f
C55 output.t11 gnd 0.462979f
C56 output.n14 gnd 0.28994f
C57 output.n15 gnd 0.015803f
C58 output.n16 gnd 0.011243f
C59 output.n17 gnd 0.006041f
C60 output.n18 gnd 0.01428f
C61 output.n19 gnd 0.006397f
C62 output.n20 gnd 0.011243f
C63 output.n21 gnd 0.006041f
C64 output.n22 gnd 0.01428f
C65 output.n23 gnd 0.006397f
C66 output.n24 gnd 0.048111f
C67 output.t19 gnd 0.023274f
C68 output.n25 gnd 0.01071f
C69 output.n26 gnd 0.008435f
C70 output.n27 gnd 0.006041f
C71 output.n28 gnd 0.267512f
C72 output.n29 gnd 0.011243f
C73 output.n30 gnd 0.006041f
C74 output.n31 gnd 0.006397f
C75 output.n32 gnd 0.01428f
C76 output.n33 gnd 0.01428f
C77 output.n34 gnd 0.006397f
C78 output.n35 gnd 0.006041f
C79 output.n36 gnd 0.011243f
C80 output.n37 gnd 0.011243f
C81 output.n38 gnd 0.006041f
C82 output.n39 gnd 0.006397f
C83 output.n40 gnd 0.01428f
C84 output.n41 gnd 0.030913f
C85 output.n42 gnd 0.006397f
C86 output.n43 gnd 0.006041f
C87 output.n44 gnd 0.025987f
C88 output.n45 gnd 0.097665f
C89 output.n46 gnd 0.015803f
C90 output.n47 gnd 0.011243f
C91 output.n48 gnd 0.006041f
C92 output.n49 gnd 0.01428f
C93 output.n50 gnd 0.006397f
C94 output.n51 gnd 0.011243f
C95 output.n52 gnd 0.006041f
C96 output.n53 gnd 0.01428f
C97 output.n54 gnd 0.006397f
C98 output.n55 gnd 0.048111f
C99 output.t17 gnd 0.023274f
C100 output.n56 gnd 0.01071f
C101 output.n57 gnd 0.008435f
C102 output.n58 gnd 0.006041f
C103 output.n59 gnd 0.267512f
C104 output.n60 gnd 0.011243f
C105 output.n61 gnd 0.006041f
C106 output.n62 gnd 0.006397f
C107 output.n63 gnd 0.01428f
C108 output.n64 gnd 0.01428f
C109 output.n65 gnd 0.006397f
C110 output.n66 gnd 0.006041f
C111 output.n67 gnd 0.011243f
C112 output.n68 gnd 0.011243f
C113 output.n69 gnd 0.006041f
C114 output.n70 gnd 0.006397f
C115 output.n71 gnd 0.01428f
C116 output.n72 gnd 0.030913f
C117 output.n73 gnd 0.006397f
C118 output.n74 gnd 0.006041f
C119 output.n75 gnd 0.025987f
C120 output.n76 gnd 0.09306f
C121 output.n77 gnd 1.65264f
C122 output.n78 gnd 0.015803f
C123 output.n79 gnd 0.011243f
C124 output.n80 gnd 0.006041f
C125 output.n81 gnd 0.01428f
C126 output.n82 gnd 0.006397f
C127 output.n83 gnd 0.011243f
C128 output.n84 gnd 0.006041f
C129 output.n85 gnd 0.01428f
C130 output.n86 gnd 0.006397f
C131 output.n87 gnd 0.048111f
C132 output.t18 gnd 0.023274f
C133 output.n88 gnd 0.01071f
C134 output.n89 gnd 0.008435f
C135 output.n90 gnd 0.006041f
C136 output.n91 gnd 0.267512f
C137 output.n92 gnd 0.011243f
C138 output.n93 gnd 0.006041f
C139 output.n94 gnd 0.006397f
C140 output.n95 gnd 0.01428f
C141 output.n96 gnd 0.01428f
C142 output.n97 gnd 0.006397f
C143 output.n98 gnd 0.006041f
C144 output.n99 gnd 0.011243f
C145 output.n100 gnd 0.011243f
C146 output.n101 gnd 0.006041f
C147 output.n102 gnd 0.006397f
C148 output.n103 gnd 0.01428f
C149 output.n104 gnd 0.030913f
C150 output.n105 gnd 0.006397f
C151 output.n106 gnd 0.006041f
C152 output.n107 gnd 0.025987f
C153 output.n108 gnd 0.09306f
C154 output.n109 gnd 0.713089f
C155 output.n110 gnd 0.015803f
C156 output.n111 gnd 0.011243f
C157 output.n112 gnd 0.006041f
C158 output.n113 gnd 0.01428f
C159 output.n114 gnd 0.006397f
C160 output.n115 gnd 0.011243f
C161 output.n116 gnd 0.006041f
C162 output.n117 gnd 0.01428f
C163 output.n118 gnd 0.006397f
C164 output.n119 gnd 0.048111f
C165 output.t16 gnd 0.023274f
C166 output.n120 gnd 0.01071f
C167 output.n121 gnd 0.008435f
C168 output.n122 gnd 0.006041f
C169 output.n123 gnd 0.267512f
C170 output.n124 gnd 0.011243f
C171 output.n125 gnd 0.006041f
C172 output.n126 gnd 0.006397f
C173 output.n127 gnd 0.01428f
C174 output.n128 gnd 0.01428f
C175 output.n129 gnd 0.006397f
C176 output.n130 gnd 0.006041f
C177 output.n131 gnd 0.011243f
C178 output.n132 gnd 0.011243f
C179 output.n133 gnd 0.006041f
C180 output.n134 gnd 0.006397f
C181 output.n135 gnd 0.01428f
C182 output.n136 gnd 0.030913f
C183 output.n137 gnd 0.006397f
C184 output.n138 gnd 0.006041f
C185 output.n139 gnd 0.025987f
C186 output.n140 gnd 0.09306f
C187 output.n141 gnd 1.67353f
C188 a_n2650_8322.t11 gnd 0.097961f
C189 a_n2650_8322.t3 gnd 20.3228f
C190 a_n2650_8322.t2 gnd 20.180302f
C191 a_n2650_8322.t5 gnd 20.180302f
C192 a_n2650_8322.t4 gnd 20.3228f
C193 a_n2650_8322.t1 gnd 20.180302f
C194 a_n2650_8322.t0 gnd 30.033998f
C195 a_n2650_8322.t21 gnd 0.917252f
C196 a_n2650_8322.t24 gnd 0.097961f
C197 a_n2650_8322.t16 gnd 0.097961f
C198 a_n2650_8322.n0 gnd 0.690034f
C199 a_n2650_8322.n1 gnd 0.771011f
C200 a_n2650_8322.t8 gnd 0.097961f
C201 a_n2650_8322.t7 gnd 0.097961f
C202 a_n2650_8322.n2 gnd 0.690034f
C203 a_n2650_8322.n3 gnd 0.391741f
C204 a_n2650_8322.t19 gnd 0.097961f
C205 a_n2650_8322.t13 gnd 0.097961f
C206 a_n2650_8322.n4 gnd 0.690034f
C207 a_n2650_8322.n5 gnd 0.391741f
C208 a_n2650_8322.t17 gnd 0.097961f
C209 a_n2650_8322.t15 gnd 0.097961f
C210 a_n2650_8322.n6 gnd 0.690034f
C211 a_n2650_8322.n7 gnd 0.391741f
C212 a_n2650_8322.t6 gnd 0.915426f
C213 a_n2650_8322.n8 gnd 1.70828f
C214 a_n2650_8322.t29 gnd 0.917252f
C215 a_n2650_8322.t33 gnd 0.097961f
C216 a_n2650_8322.t32 gnd 0.097961f
C217 a_n2650_8322.n9 gnd 0.690034f
C218 a_n2650_8322.n10 gnd 0.771011f
C219 a_n2650_8322.t27 gnd 0.915426f
C220 a_n2650_8322.n11 gnd 0.387983f
C221 a_n2650_8322.t30 gnd 0.915426f
C222 a_n2650_8322.n12 gnd 0.387983f
C223 a_n2650_8322.t28 gnd 0.097961f
C224 a_n2650_8322.t26 gnd 0.097961f
C225 a_n2650_8322.n13 gnd 0.690034f
C226 a_n2650_8322.n14 gnd 0.391741f
C227 a_n2650_8322.t31 gnd 0.915426f
C228 a_n2650_8322.n15 gnd 1.27292f
C229 a_n2650_8322.n16 gnd 2.07982f
C230 a_n2650_8322.n17 gnd 3.90316f
C231 a_n2650_8322.t20 gnd 0.915426f
C232 a_n2650_8322.n18 gnd 0.995719f
C233 a_n2650_8322.t10 gnd 0.097961f
C234 a_n2650_8322.t9 gnd 0.097961f
C235 a_n2650_8322.n19 gnd 0.690034f
C236 a_n2650_8322.n20 gnd 0.391741f
C237 a_n2650_8322.t22 gnd 0.097961f
C238 a_n2650_8322.t12 gnd 0.097961f
C239 a_n2650_8322.n21 gnd 0.690034f
C240 a_n2650_8322.n22 gnd 0.391741f
C241 a_n2650_8322.t23 gnd 0.91725f
C242 a_n2650_8322.t18 gnd 0.097961f
C243 a_n2650_8322.t14 gnd 0.097961f
C244 a_n2650_8322.n23 gnd 0.690034f
C245 a_n2650_8322.n24 gnd 0.771013f
C246 a_n2650_8322.n25 gnd 0.391739f
C247 a_n2650_8322.n26 gnd 0.690035f
C248 a_n2650_8322.t25 gnd 0.097961f
C249 commonsourceibias.n0 gnd 0.010724f
C250 commonsourceibias.t115 gnd 0.162395f
C251 commonsourceibias.t136 gnd 0.150157f
C252 commonsourceibias.n1 gnd 0.007823f
C253 commonsourceibias.n2 gnd 0.008037f
C254 commonsourceibias.t151 gnd 0.150157f
C255 commonsourceibias.n3 gnd 0.01034f
C256 commonsourceibias.n4 gnd 0.008037f
C257 commonsourceibias.t105 gnd 0.150157f
C258 commonsourceibias.n5 gnd 0.059912f
C259 commonsourceibias.t126 gnd 0.150157f
C260 commonsourceibias.n6 gnd 0.007578f
C261 commonsourceibias.n7 gnd 0.008037f
C262 commonsourceibias.t144 gnd 0.150157f
C263 commonsourceibias.n8 gnd 0.010186f
C264 commonsourceibias.n9 gnd 0.008037f
C265 commonsourceibias.t98 gnd 0.150157f
C266 commonsourceibias.n10 gnd 0.059912f
C267 commonsourceibias.t94 gnd 0.150157f
C268 commonsourceibias.n11 gnd 0.007361f
C269 commonsourceibias.n12 gnd 0.008037f
C270 commonsourceibias.t135 gnd 0.150157f
C271 commonsourceibias.n13 gnd 0.010015f
C272 commonsourceibias.n14 gnd 0.010724f
C273 commonsourceibias.t74 gnd 0.162395f
C274 commonsourceibias.t20 gnd 0.150157f
C275 commonsourceibias.n15 gnd 0.007823f
C276 commonsourceibias.n16 gnd 0.008037f
C277 commonsourceibias.t50 gnd 0.150157f
C278 commonsourceibias.n17 gnd 0.01034f
C279 commonsourceibias.n18 gnd 0.008037f
C280 commonsourceibias.t8 gnd 0.150157f
C281 commonsourceibias.n19 gnd 0.059912f
C282 commonsourceibias.t36 gnd 0.150157f
C283 commonsourceibias.n20 gnd 0.007578f
C284 commonsourceibias.n21 gnd 0.008037f
C285 commonsourceibias.t76 gnd 0.150157f
C286 commonsourceibias.n22 gnd 0.010186f
C287 commonsourceibias.n23 gnd 0.008037f
C288 commonsourceibias.t24 gnd 0.150157f
C289 commonsourceibias.n24 gnd 0.059912f
C290 commonsourceibias.t34 gnd 0.150157f
C291 commonsourceibias.n25 gnd 0.007361f
C292 commonsourceibias.n26 gnd 0.008037f
C293 commonsourceibias.t10 gnd 0.150157f
C294 commonsourceibias.n27 gnd 0.010015f
C295 commonsourceibias.n28 gnd 0.008037f
C296 commonsourceibias.t40 gnd 0.150157f
C297 commonsourceibias.n29 gnd 0.059912f
C298 commonsourceibias.t56 gnd 0.150157f
C299 commonsourceibias.n30 gnd 0.007172f
C300 commonsourceibias.n31 gnd 0.008037f
C301 commonsourceibias.t26 gnd 0.150157f
C302 commonsourceibias.n32 gnd 0.009825f
C303 commonsourceibias.n33 gnd 0.008037f
C304 commonsourceibias.t38 gnd 0.150157f
C305 commonsourceibias.n34 gnd 0.059912f
C306 commonsourceibias.t70 gnd 0.150157f
C307 commonsourceibias.n35 gnd 0.007008f
C308 commonsourceibias.n36 gnd 0.008037f
C309 commonsourceibias.t18 gnd 0.150157f
C310 commonsourceibias.n37 gnd 0.009613f
C311 commonsourceibias.n38 gnd 0.008037f
C312 commonsourceibias.t22 gnd 0.150157f
C313 commonsourceibias.n39 gnd 0.059912f
C314 commonsourceibias.t54 gnd 0.150157f
C315 commonsourceibias.n40 gnd 0.006868f
C316 commonsourceibias.n41 gnd 0.008037f
C317 commonsourceibias.t4 gnd 0.150157f
C318 commonsourceibias.n42 gnd 0.009378f
C319 commonsourceibias.t78 gnd 0.166947f
C320 commonsourceibias.t46 gnd 0.150157f
C321 commonsourceibias.n43 gnd 0.065449f
C322 commonsourceibias.n44 gnd 0.071822f
C323 commonsourceibias.n45 gnd 0.033327f
C324 commonsourceibias.n46 gnd 0.008037f
C325 commonsourceibias.n47 gnd 0.007823f
C326 commonsourceibias.n48 gnd 0.01121f
C327 commonsourceibias.n49 gnd 0.059912f
C328 commonsourceibias.n50 gnd 0.011203f
C329 commonsourceibias.n51 gnd 0.008037f
C330 commonsourceibias.n52 gnd 0.008037f
C331 commonsourceibias.n53 gnd 0.008037f
C332 commonsourceibias.n54 gnd 0.01034f
C333 commonsourceibias.n55 gnd 0.059912f
C334 commonsourceibias.n56 gnd 0.010583f
C335 commonsourceibias.n57 gnd 0.010282f
C336 commonsourceibias.n58 gnd 0.008037f
C337 commonsourceibias.n59 gnd 0.008037f
C338 commonsourceibias.n60 gnd 0.008037f
C339 commonsourceibias.n61 gnd 0.007578f
C340 commonsourceibias.n62 gnd 0.01122f
C341 commonsourceibias.n63 gnd 0.059912f
C342 commonsourceibias.n64 gnd 0.011217f
C343 commonsourceibias.n65 gnd 0.008037f
C344 commonsourceibias.n66 gnd 0.008037f
C345 commonsourceibias.n67 gnd 0.008037f
C346 commonsourceibias.n68 gnd 0.010186f
C347 commonsourceibias.n69 gnd 0.059912f
C348 commonsourceibias.n70 gnd 0.010507f
C349 commonsourceibias.n71 gnd 0.010357f
C350 commonsourceibias.n72 gnd 0.008037f
C351 commonsourceibias.n73 gnd 0.008037f
C352 commonsourceibias.n74 gnd 0.008037f
C353 commonsourceibias.n75 gnd 0.007361f
C354 commonsourceibias.n76 gnd 0.011225f
C355 commonsourceibias.n77 gnd 0.059912f
C356 commonsourceibias.n78 gnd 0.011224f
C357 commonsourceibias.n79 gnd 0.008037f
C358 commonsourceibias.n80 gnd 0.008037f
C359 commonsourceibias.n81 gnd 0.008037f
C360 commonsourceibias.n82 gnd 0.010015f
C361 commonsourceibias.n83 gnd 0.059912f
C362 commonsourceibias.n84 gnd 0.010432f
C363 commonsourceibias.n85 gnd 0.010432f
C364 commonsourceibias.n86 gnd 0.008037f
C365 commonsourceibias.n87 gnd 0.008037f
C366 commonsourceibias.n88 gnd 0.008037f
C367 commonsourceibias.n89 gnd 0.007172f
C368 commonsourceibias.n90 gnd 0.011224f
C369 commonsourceibias.n91 gnd 0.059912f
C370 commonsourceibias.n92 gnd 0.011225f
C371 commonsourceibias.n93 gnd 0.008037f
C372 commonsourceibias.n94 gnd 0.008037f
C373 commonsourceibias.n95 gnd 0.008037f
C374 commonsourceibias.n96 gnd 0.009825f
C375 commonsourceibias.n97 gnd 0.059912f
C376 commonsourceibias.n98 gnd 0.010357f
C377 commonsourceibias.n99 gnd 0.010507f
C378 commonsourceibias.n100 gnd 0.008037f
C379 commonsourceibias.n101 gnd 0.008037f
C380 commonsourceibias.n102 gnd 0.008037f
C381 commonsourceibias.n103 gnd 0.007008f
C382 commonsourceibias.n104 gnd 0.011217f
C383 commonsourceibias.n105 gnd 0.059912f
C384 commonsourceibias.n106 gnd 0.01122f
C385 commonsourceibias.n107 gnd 0.008037f
C386 commonsourceibias.n108 gnd 0.008037f
C387 commonsourceibias.n109 gnd 0.008037f
C388 commonsourceibias.n110 gnd 0.009613f
C389 commonsourceibias.n111 gnd 0.059912f
C390 commonsourceibias.n112 gnd 0.010282f
C391 commonsourceibias.n113 gnd 0.010583f
C392 commonsourceibias.n114 gnd 0.008037f
C393 commonsourceibias.n115 gnd 0.008037f
C394 commonsourceibias.n116 gnd 0.008037f
C395 commonsourceibias.n117 gnd 0.006868f
C396 commonsourceibias.n118 gnd 0.011203f
C397 commonsourceibias.n119 gnd 0.059912f
C398 commonsourceibias.n120 gnd 0.01121f
C399 commonsourceibias.n121 gnd 0.008037f
C400 commonsourceibias.n122 gnd 0.008037f
C401 commonsourceibias.n123 gnd 0.008037f
C402 commonsourceibias.n124 gnd 0.009378f
C403 commonsourceibias.n125 gnd 0.059912f
C404 commonsourceibias.n126 gnd 0.009861f
C405 commonsourceibias.n127 gnd 0.07189f
C406 commonsourceibias.n128 gnd 0.080075f
C407 commonsourceibias.t75 gnd 0.017343f
C408 commonsourceibias.t21 gnd 0.017343f
C409 commonsourceibias.n129 gnd 0.15325f
C410 commonsourceibias.n130 gnd 0.132562f
C411 commonsourceibias.t51 gnd 0.017343f
C412 commonsourceibias.t9 gnd 0.017343f
C413 commonsourceibias.n131 gnd 0.15325f
C414 commonsourceibias.n132 gnd 0.070394f
C415 commonsourceibias.t37 gnd 0.017343f
C416 commonsourceibias.t77 gnd 0.017343f
C417 commonsourceibias.n133 gnd 0.15325f
C418 commonsourceibias.n134 gnd 0.070394f
C419 commonsourceibias.t25 gnd 0.017343f
C420 commonsourceibias.t35 gnd 0.017343f
C421 commonsourceibias.n135 gnd 0.15325f
C422 commonsourceibias.n136 gnd 0.070394f
C423 commonsourceibias.t11 gnd 0.017343f
C424 commonsourceibias.t41 gnd 0.017343f
C425 commonsourceibias.n137 gnd 0.15325f
C426 commonsourceibias.n138 gnd 0.058811f
C427 commonsourceibias.t47 gnd 0.017343f
C428 commonsourceibias.t79 gnd 0.017343f
C429 commonsourceibias.n139 gnd 0.153763f
C430 commonsourceibias.t55 gnd 0.017343f
C431 commonsourceibias.t5 gnd 0.017343f
C432 commonsourceibias.n140 gnd 0.15325f
C433 commonsourceibias.n141 gnd 0.1428f
C434 commonsourceibias.t19 gnd 0.017343f
C435 commonsourceibias.t23 gnd 0.017343f
C436 commonsourceibias.n142 gnd 0.15325f
C437 commonsourceibias.n143 gnd 0.070394f
C438 commonsourceibias.t39 gnd 0.017343f
C439 commonsourceibias.t71 gnd 0.017343f
C440 commonsourceibias.n144 gnd 0.15325f
C441 commonsourceibias.n145 gnd 0.070394f
C442 commonsourceibias.t57 gnd 0.017343f
C443 commonsourceibias.t27 gnd 0.017343f
C444 commonsourceibias.n146 gnd 0.15325f
C445 commonsourceibias.n147 gnd 0.058811f
C446 commonsourceibias.n148 gnd 0.071213f
C447 commonsourceibias.n149 gnd 0.052016f
C448 commonsourceibias.t153 gnd 0.150157f
C449 commonsourceibias.n150 gnd 0.059912f
C450 commonsourceibias.t88 gnd 0.150157f
C451 commonsourceibias.n151 gnd 0.059912f
C452 commonsourceibias.n152 gnd 0.008037f
C453 commonsourceibias.t125 gnd 0.150157f
C454 commonsourceibias.n153 gnd 0.059912f
C455 commonsourceibias.n154 gnd 0.008037f
C456 commonsourceibias.t120 gnd 0.150157f
C457 commonsourceibias.n155 gnd 0.059912f
C458 commonsourceibias.n156 gnd 0.008037f
C459 commonsourceibias.t139 gnd 0.150157f
C460 commonsourceibias.n157 gnd 0.007008f
C461 commonsourceibias.n158 gnd 0.008037f
C462 commonsourceibias.t112 gnd 0.150157f
C463 commonsourceibias.n159 gnd 0.009613f
C464 commonsourceibias.n160 gnd 0.008037f
C465 commonsourceibias.t107 gnd 0.150157f
C466 commonsourceibias.n161 gnd 0.059912f
C467 commonsourceibias.t127 gnd 0.150157f
C468 commonsourceibias.n162 gnd 0.006868f
C469 commonsourceibias.n163 gnd 0.008037f
C470 commonsourceibias.t146 gnd 0.150157f
C471 commonsourceibias.n164 gnd 0.009378f
C472 commonsourceibias.t117 gnd 0.166947f
C473 commonsourceibias.t99 gnd 0.150157f
C474 commonsourceibias.n165 gnd 0.065449f
C475 commonsourceibias.n166 gnd 0.071822f
C476 commonsourceibias.n167 gnd 0.033327f
C477 commonsourceibias.n168 gnd 0.008037f
C478 commonsourceibias.n169 gnd 0.007823f
C479 commonsourceibias.n170 gnd 0.01121f
C480 commonsourceibias.n171 gnd 0.059912f
C481 commonsourceibias.n172 gnd 0.011203f
C482 commonsourceibias.n173 gnd 0.008037f
C483 commonsourceibias.n174 gnd 0.008037f
C484 commonsourceibias.n175 gnd 0.008037f
C485 commonsourceibias.n176 gnd 0.01034f
C486 commonsourceibias.n177 gnd 0.059912f
C487 commonsourceibias.n178 gnd 0.010583f
C488 commonsourceibias.n179 gnd 0.010282f
C489 commonsourceibias.n180 gnd 0.008037f
C490 commonsourceibias.n181 gnd 0.008037f
C491 commonsourceibias.n182 gnd 0.008037f
C492 commonsourceibias.n183 gnd 0.007578f
C493 commonsourceibias.n184 gnd 0.01122f
C494 commonsourceibias.n185 gnd 0.059912f
C495 commonsourceibias.n186 gnd 0.011217f
C496 commonsourceibias.n187 gnd 0.008037f
C497 commonsourceibias.n188 gnd 0.008037f
C498 commonsourceibias.n189 gnd 0.008037f
C499 commonsourceibias.n190 gnd 0.010186f
C500 commonsourceibias.n191 gnd 0.059912f
C501 commonsourceibias.n192 gnd 0.010507f
C502 commonsourceibias.n193 gnd 0.010357f
C503 commonsourceibias.n194 gnd 0.008037f
C504 commonsourceibias.n195 gnd 0.008037f
C505 commonsourceibias.n196 gnd 0.009825f
C506 commonsourceibias.n197 gnd 0.007361f
C507 commonsourceibias.n198 gnd 0.011225f
C508 commonsourceibias.n199 gnd 0.008037f
C509 commonsourceibias.n200 gnd 0.008037f
C510 commonsourceibias.n201 gnd 0.011224f
C511 commonsourceibias.n202 gnd 0.007172f
C512 commonsourceibias.n203 gnd 0.010015f
C513 commonsourceibias.n204 gnd 0.008037f
C514 commonsourceibias.n205 gnd 0.007021f
C515 commonsourceibias.n206 gnd 0.010432f
C516 commonsourceibias.n207 gnd 0.010432f
C517 commonsourceibias.n208 gnd 0.007021f
C518 commonsourceibias.n209 gnd 0.008037f
C519 commonsourceibias.n210 gnd 0.008037f
C520 commonsourceibias.n211 gnd 0.007172f
C521 commonsourceibias.n212 gnd 0.011224f
C522 commonsourceibias.n213 gnd 0.059912f
C523 commonsourceibias.n214 gnd 0.011225f
C524 commonsourceibias.n215 gnd 0.008037f
C525 commonsourceibias.n216 gnd 0.008037f
C526 commonsourceibias.n217 gnd 0.008037f
C527 commonsourceibias.n218 gnd 0.009825f
C528 commonsourceibias.n219 gnd 0.059912f
C529 commonsourceibias.n220 gnd 0.010357f
C530 commonsourceibias.n221 gnd 0.010507f
C531 commonsourceibias.n222 gnd 0.008037f
C532 commonsourceibias.n223 gnd 0.008037f
C533 commonsourceibias.n224 gnd 0.008037f
C534 commonsourceibias.n225 gnd 0.007008f
C535 commonsourceibias.n226 gnd 0.011217f
C536 commonsourceibias.n227 gnd 0.059912f
C537 commonsourceibias.n228 gnd 0.01122f
C538 commonsourceibias.n229 gnd 0.008037f
C539 commonsourceibias.n230 gnd 0.008037f
C540 commonsourceibias.n231 gnd 0.008037f
C541 commonsourceibias.n232 gnd 0.009613f
C542 commonsourceibias.n233 gnd 0.059912f
C543 commonsourceibias.n234 gnd 0.010282f
C544 commonsourceibias.n235 gnd 0.010583f
C545 commonsourceibias.n236 gnd 0.008037f
C546 commonsourceibias.n237 gnd 0.008037f
C547 commonsourceibias.n238 gnd 0.008037f
C548 commonsourceibias.n239 gnd 0.006868f
C549 commonsourceibias.n240 gnd 0.011203f
C550 commonsourceibias.n241 gnd 0.059912f
C551 commonsourceibias.n242 gnd 0.01121f
C552 commonsourceibias.n243 gnd 0.008037f
C553 commonsourceibias.n244 gnd 0.008037f
C554 commonsourceibias.n245 gnd 0.008037f
C555 commonsourceibias.n246 gnd 0.009378f
C556 commonsourceibias.n247 gnd 0.059912f
C557 commonsourceibias.n248 gnd 0.009861f
C558 commonsourceibias.n249 gnd 0.07189f
C559 commonsourceibias.n250 gnd 0.04697f
C560 commonsourceibias.n251 gnd 0.010724f
C561 commonsourceibias.t119 gnd 0.150157f
C562 commonsourceibias.n252 gnd 0.007823f
C563 commonsourceibias.n253 gnd 0.008037f
C564 commonsourceibias.t137 gnd 0.150157f
C565 commonsourceibias.n254 gnd 0.01034f
C566 commonsourceibias.n255 gnd 0.008037f
C567 commonsourceibias.t92 gnd 0.150157f
C568 commonsourceibias.n256 gnd 0.059912f
C569 commonsourceibias.t109 gnd 0.150157f
C570 commonsourceibias.n257 gnd 0.007578f
C571 commonsourceibias.n258 gnd 0.008037f
C572 commonsourceibias.t128 gnd 0.150157f
C573 commonsourceibias.n259 gnd 0.010186f
C574 commonsourceibias.n260 gnd 0.008037f
C575 commonsourceibias.t86 gnd 0.150157f
C576 commonsourceibias.n261 gnd 0.059912f
C577 commonsourceibias.t83 gnd 0.150157f
C578 commonsourceibias.n262 gnd 0.007361f
C579 commonsourceibias.n263 gnd 0.008037f
C580 commonsourceibias.t118 gnd 0.150157f
C581 commonsourceibias.n264 gnd 0.010015f
C582 commonsourceibias.n265 gnd 0.008037f
C583 commonsourceibias.t138 gnd 0.150157f
C584 commonsourceibias.n266 gnd 0.059912f
C585 commonsourceibias.t159 gnd 0.150157f
C586 commonsourceibias.n267 gnd 0.007172f
C587 commonsourceibias.n268 gnd 0.008037f
C588 commonsourceibias.t108 gnd 0.150157f
C589 commonsourceibias.n269 gnd 0.009825f
C590 commonsourceibias.n270 gnd 0.008037f
C591 commonsourceibias.t102 gnd 0.150157f
C592 commonsourceibias.n271 gnd 0.059912f
C593 commonsourceibias.t121 gnd 0.150157f
C594 commonsourceibias.n272 gnd 0.007008f
C595 commonsourceibias.n273 gnd 0.008037f
C596 commonsourceibias.t95 gnd 0.150157f
C597 commonsourceibias.n274 gnd 0.009613f
C598 commonsourceibias.n275 gnd 0.008037f
C599 commonsourceibias.t93 gnd 0.150157f
C600 commonsourceibias.n276 gnd 0.059912f
C601 commonsourceibias.t110 gnd 0.150157f
C602 commonsourceibias.n277 gnd 0.006868f
C603 commonsourceibias.n278 gnd 0.008037f
C604 commonsourceibias.t129 gnd 0.150157f
C605 commonsourceibias.n279 gnd 0.009378f
C606 commonsourceibias.t101 gnd 0.166947f
C607 commonsourceibias.t87 gnd 0.150157f
C608 commonsourceibias.n280 gnd 0.065449f
C609 commonsourceibias.n281 gnd 0.071822f
C610 commonsourceibias.n282 gnd 0.033327f
C611 commonsourceibias.n283 gnd 0.008037f
C612 commonsourceibias.n284 gnd 0.007823f
C613 commonsourceibias.n285 gnd 0.01121f
C614 commonsourceibias.n286 gnd 0.059912f
C615 commonsourceibias.n287 gnd 0.011203f
C616 commonsourceibias.n288 gnd 0.008037f
C617 commonsourceibias.n289 gnd 0.008037f
C618 commonsourceibias.n290 gnd 0.008037f
C619 commonsourceibias.n291 gnd 0.01034f
C620 commonsourceibias.n292 gnd 0.059912f
C621 commonsourceibias.n293 gnd 0.010583f
C622 commonsourceibias.n294 gnd 0.010282f
C623 commonsourceibias.n295 gnd 0.008037f
C624 commonsourceibias.n296 gnd 0.008037f
C625 commonsourceibias.n297 gnd 0.008037f
C626 commonsourceibias.n298 gnd 0.007578f
C627 commonsourceibias.n299 gnd 0.01122f
C628 commonsourceibias.n300 gnd 0.059912f
C629 commonsourceibias.n301 gnd 0.011217f
C630 commonsourceibias.n302 gnd 0.008037f
C631 commonsourceibias.n303 gnd 0.008037f
C632 commonsourceibias.n304 gnd 0.008037f
C633 commonsourceibias.n305 gnd 0.010186f
C634 commonsourceibias.n306 gnd 0.059912f
C635 commonsourceibias.n307 gnd 0.010507f
C636 commonsourceibias.n308 gnd 0.010357f
C637 commonsourceibias.n309 gnd 0.008037f
C638 commonsourceibias.n310 gnd 0.008037f
C639 commonsourceibias.n311 gnd 0.008037f
C640 commonsourceibias.n312 gnd 0.007361f
C641 commonsourceibias.n313 gnd 0.011225f
C642 commonsourceibias.n314 gnd 0.059912f
C643 commonsourceibias.n315 gnd 0.011224f
C644 commonsourceibias.n316 gnd 0.008037f
C645 commonsourceibias.n317 gnd 0.008037f
C646 commonsourceibias.n318 gnd 0.008037f
C647 commonsourceibias.n319 gnd 0.010015f
C648 commonsourceibias.n320 gnd 0.059912f
C649 commonsourceibias.n321 gnd 0.010432f
C650 commonsourceibias.n322 gnd 0.010432f
C651 commonsourceibias.n323 gnd 0.008037f
C652 commonsourceibias.n324 gnd 0.008037f
C653 commonsourceibias.n325 gnd 0.008037f
C654 commonsourceibias.n326 gnd 0.007172f
C655 commonsourceibias.n327 gnd 0.011224f
C656 commonsourceibias.n328 gnd 0.059912f
C657 commonsourceibias.n329 gnd 0.011225f
C658 commonsourceibias.n330 gnd 0.008037f
C659 commonsourceibias.n331 gnd 0.008037f
C660 commonsourceibias.n332 gnd 0.008037f
C661 commonsourceibias.n333 gnd 0.009825f
C662 commonsourceibias.n334 gnd 0.059912f
C663 commonsourceibias.n335 gnd 0.010357f
C664 commonsourceibias.n336 gnd 0.010507f
C665 commonsourceibias.n337 gnd 0.008037f
C666 commonsourceibias.n338 gnd 0.008037f
C667 commonsourceibias.n339 gnd 0.008037f
C668 commonsourceibias.n340 gnd 0.007008f
C669 commonsourceibias.n341 gnd 0.011217f
C670 commonsourceibias.n342 gnd 0.059912f
C671 commonsourceibias.n343 gnd 0.01122f
C672 commonsourceibias.n344 gnd 0.008037f
C673 commonsourceibias.n345 gnd 0.008037f
C674 commonsourceibias.n346 gnd 0.008037f
C675 commonsourceibias.n347 gnd 0.009613f
C676 commonsourceibias.n348 gnd 0.059912f
C677 commonsourceibias.n349 gnd 0.010282f
C678 commonsourceibias.n350 gnd 0.010583f
C679 commonsourceibias.n351 gnd 0.008037f
C680 commonsourceibias.n352 gnd 0.008037f
C681 commonsourceibias.n353 gnd 0.008037f
C682 commonsourceibias.n354 gnd 0.006868f
C683 commonsourceibias.n355 gnd 0.011203f
C684 commonsourceibias.n356 gnd 0.059912f
C685 commonsourceibias.n357 gnd 0.01121f
C686 commonsourceibias.n358 gnd 0.008037f
C687 commonsourceibias.n359 gnd 0.008037f
C688 commonsourceibias.n360 gnd 0.008037f
C689 commonsourceibias.n361 gnd 0.009378f
C690 commonsourceibias.n362 gnd 0.059912f
C691 commonsourceibias.n363 gnd 0.009861f
C692 commonsourceibias.t100 gnd 0.162395f
C693 commonsourceibias.n364 gnd 0.07189f
C694 commonsourceibias.n365 gnd 0.025003f
C695 commonsourceibias.n366 gnd 0.464917f
C696 commonsourceibias.n367 gnd 0.010724f
C697 commonsourceibias.t140 gnd 0.162395f
C698 commonsourceibias.t155 gnd 0.150157f
C699 commonsourceibias.n368 gnd 0.007823f
C700 commonsourceibias.n369 gnd 0.008037f
C701 commonsourceibias.t84 gnd 0.150157f
C702 commonsourceibias.n370 gnd 0.01034f
C703 commonsourceibias.n371 gnd 0.008037f
C704 commonsourceibias.t148 gnd 0.150157f
C705 commonsourceibias.n372 gnd 0.007578f
C706 commonsourceibias.n373 gnd 0.008037f
C707 commonsourceibias.t80 gnd 0.150157f
C708 commonsourceibias.n374 gnd 0.010186f
C709 commonsourceibias.n375 gnd 0.008037f
C710 commonsourceibias.t113 gnd 0.150157f
C711 commonsourceibias.n376 gnd 0.007361f
C712 commonsourceibias.n377 gnd 0.008037f
C713 commonsourceibias.t154 gnd 0.150157f
C714 commonsourceibias.n378 gnd 0.010015f
C715 commonsourceibias.t29 gnd 0.017343f
C716 commonsourceibias.t3 gnd 0.017343f
C717 commonsourceibias.n379 gnd 0.153763f
C718 commonsourceibias.t49 gnd 0.017343f
C719 commonsourceibias.t13 gnd 0.017343f
C720 commonsourceibias.n380 gnd 0.15325f
C721 commonsourceibias.n381 gnd 0.1428f
C722 commonsourceibias.t69 gnd 0.017343f
C723 commonsourceibias.t67 gnd 0.017343f
C724 commonsourceibias.n382 gnd 0.15325f
C725 commonsourceibias.n383 gnd 0.070394f
C726 commonsourceibias.t7 gnd 0.017343f
C727 commonsourceibias.t63 gnd 0.017343f
C728 commonsourceibias.n384 gnd 0.15325f
C729 commonsourceibias.n385 gnd 0.070394f
C730 commonsourceibias.t53 gnd 0.017343f
C731 commonsourceibias.t73 gnd 0.017343f
C732 commonsourceibias.n386 gnd 0.15325f
C733 commonsourceibias.n387 gnd 0.058811f
C734 commonsourceibias.n388 gnd 0.010724f
C735 commonsourceibias.t42 gnd 0.150157f
C736 commonsourceibias.n389 gnd 0.007823f
C737 commonsourceibias.n390 gnd 0.008037f
C738 commonsourceibias.t0 gnd 0.150157f
C739 commonsourceibias.n391 gnd 0.01034f
C740 commonsourceibias.n392 gnd 0.008037f
C741 commonsourceibias.t60 gnd 0.150157f
C742 commonsourceibias.n393 gnd 0.007578f
C743 commonsourceibias.n394 gnd 0.008037f
C744 commonsourceibias.t16 gnd 0.150157f
C745 commonsourceibias.n395 gnd 0.010186f
C746 commonsourceibias.n396 gnd 0.008037f
C747 commonsourceibias.t58 gnd 0.150157f
C748 commonsourceibias.n397 gnd 0.007361f
C749 commonsourceibias.n398 gnd 0.008037f
C750 commonsourceibias.t32 gnd 0.150157f
C751 commonsourceibias.n399 gnd 0.010015f
C752 commonsourceibias.n400 gnd 0.008037f
C753 commonsourceibias.t72 gnd 0.150157f
C754 commonsourceibias.n401 gnd 0.007172f
C755 commonsourceibias.n402 gnd 0.008037f
C756 commonsourceibias.t52 gnd 0.150157f
C757 commonsourceibias.n403 gnd 0.009825f
C758 commonsourceibias.n404 gnd 0.008037f
C759 commonsourceibias.t6 gnd 0.150157f
C760 commonsourceibias.n405 gnd 0.007008f
C761 commonsourceibias.n406 gnd 0.008037f
C762 commonsourceibias.t66 gnd 0.150157f
C763 commonsourceibias.n407 gnd 0.009613f
C764 commonsourceibias.n408 gnd 0.008037f
C765 commonsourceibias.t12 gnd 0.150157f
C766 commonsourceibias.n409 gnd 0.006868f
C767 commonsourceibias.n410 gnd 0.008037f
C768 commonsourceibias.t48 gnd 0.150157f
C769 commonsourceibias.n411 gnd 0.009378f
C770 commonsourceibias.t28 gnd 0.166947f
C771 commonsourceibias.t2 gnd 0.150157f
C772 commonsourceibias.n412 gnd 0.065449f
C773 commonsourceibias.n413 gnd 0.071822f
C774 commonsourceibias.n414 gnd 0.033327f
C775 commonsourceibias.n415 gnd 0.008037f
C776 commonsourceibias.n416 gnd 0.007823f
C777 commonsourceibias.n417 gnd 0.01121f
C778 commonsourceibias.n418 gnd 0.059912f
C779 commonsourceibias.n419 gnd 0.011203f
C780 commonsourceibias.n420 gnd 0.008037f
C781 commonsourceibias.n421 gnd 0.008037f
C782 commonsourceibias.n422 gnd 0.008037f
C783 commonsourceibias.n423 gnd 0.01034f
C784 commonsourceibias.n424 gnd 0.059912f
C785 commonsourceibias.n425 gnd 0.010583f
C786 commonsourceibias.t68 gnd 0.150157f
C787 commonsourceibias.n426 gnd 0.059912f
C788 commonsourceibias.n427 gnd 0.010282f
C789 commonsourceibias.n428 gnd 0.008037f
C790 commonsourceibias.n429 gnd 0.008037f
C791 commonsourceibias.n430 gnd 0.008037f
C792 commonsourceibias.n431 gnd 0.007578f
C793 commonsourceibias.n432 gnd 0.01122f
C794 commonsourceibias.n433 gnd 0.059912f
C795 commonsourceibias.n434 gnd 0.011217f
C796 commonsourceibias.n435 gnd 0.008037f
C797 commonsourceibias.n436 gnd 0.008037f
C798 commonsourceibias.n437 gnd 0.008037f
C799 commonsourceibias.n438 gnd 0.010186f
C800 commonsourceibias.n439 gnd 0.059912f
C801 commonsourceibias.n440 gnd 0.010507f
C802 commonsourceibias.t62 gnd 0.150157f
C803 commonsourceibias.n441 gnd 0.059912f
C804 commonsourceibias.n442 gnd 0.010357f
C805 commonsourceibias.n443 gnd 0.008037f
C806 commonsourceibias.n444 gnd 0.008037f
C807 commonsourceibias.n445 gnd 0.008037f
C808 commonsourceibias.n446 gnd 0.007361f
C809 commonsourceibias.n447 gnd 0.011225f
C810 commonsourceibias.n448 gnd 0.059912f
C811 commonsourceibias.n449 gnd 0.011224f
C812 commonsourceibias.n450 gnd 0.008037f
C813 commonsourceibias.n451 gnd 0.008037f
C814 commonsourceibias.n452 gnd 0.008037f
C815 commonsourceibias.n453 gnd 0.010015f
C816 commonsourceibias.n454 gnd 0.059912f
C817 commonsourceibias.n455 gnd 0.010432f
C818 commonsourceibias.t64 gnd 0.150157f
C819 commonsourceibias.n456 gnd 0.059912f
C820 commonsourceibias.n457 gnd 0.010432f
C821 commonsourceibias.n458 gnd 0.008037f
C822 commonsourceibias.n459 gnd 0.008037f
C823 commonsourceibias.n460 gnd 0.008037f
C824 commonsourceibias.n461 gnd 0.007172f
C825 commonsourceibias.n462 gnd 0.011224f
C826 commonsourceibias.n463 gnd 0.059912f
C827 commonsourceibias.n464 gnd 0.011225f
C828 commonsourceibias.n465 gnd 0.008037f
C829 commonsourceibias.n466 gnd 0.008037f
C830 commonsourceibias.n467 gnd 0.008037f
C831 commonsourceibias.n468 gnd 0.009825f
C832 commonsourceibias.n469 gnd 0.059912f
C833 commonsourceibias.n470 gnd 0.010357f
C834 commonsourceibias.t44 gnd 0.150157f
C835 commonsourceibias.n471 gnd 0.059912f
C836 commonsourceibias.n472 gnd 0.010507f
C837 commonsourceibias.n473 gnd 0.008037f
C838 commonsourceibias.n474 gnd 0.008037f
C839 commonsourceibias.n475 gnd 0.008037f
C840 commonsourceibias.n476 gnd 0.007008f
C841 commonsourceibias.n477 gnd 0.011217f
C842 commonsourceibias.n478 gnd 0.059912f
C843 commonsourceibias.n479 gnd 0.01122f
C844 commonsourceibias.n480 gnd 0.008037f
C845 commonsourceibias.n481 gnd 0.008037f
C846 commonsourceibias.n482 gnd 0.008037f
C847 commonsourceibias.n483 gnd 0.009613f
C848 commonsourceibias.n484 gnd 0.059912f
C849 commonsourceibias.n485 gnd 0.010282f
C850 commonsourceibias.t30 gnd 0.150157f
C851 commonsourceibias.n486 gnd 0.059912f
C852 commonsourceibias.n487 gnd 0.010583f
C853 commonsourceibias.n488 gnd 0.008037f
C854 commonsourceibias.n489 gnd 0.008037f
C855 commonsourceibias.n490 gnd 0.008037f
C856 commonsourceibias.n491 gnd 0.006868f
C857 commonsourceibias.n492 gnd 0.011203f
C858 commonsourceibias.n493 gnd 0.059912f
C859 commonsourceibias.n494 gnd 0.01121f
C860 commonsourceibias.n495 gnd 0.008037f
C861 commonsourceibias.n496 gnd 0.008037f
C862 commonsourceibias.n497 gnd 0.008037f
C863 commonsourceibias.n498 gnd 0.009378f
C864 commonsourceibias.n499 gnd 0.059912f
C865 commonsourceibias.n500 gnd 0.009861f
C866 commonsourceibias.t14 gnd 0.162395f
C867 commonsourceibias.n501 gnd 0.07189f
C868 commonsourceibias.n502 gnd 0.080075f
C869 commonsourceibias.t43 gnd 0.017343f
C870 commonsourceibias.t15 gnd 0.017343f
C871 commonsourceibias.n503 gnd 0.15325f
C872 commonsourceibias.n504 gnd 0.132562f
C873 commonsourceibias.t31 gnd 0.017343f
C874 commonsourceibias.t1 gnd 0.017343f
C875 commonsourceibias.n505 gnd 0.15325f
C876 commonsourceibias.n506 gnd 0.070394f
C877 commonsourceibias.t17 gnd 0.017343f
C878 commonsourceibias.t61 gnd 0.017343f
C879 commonsourceibias.n507 gnd 0.15325f
C880 commonsourceibias.n508 gnd 0.070394f
C881 commonsourceibias.t59 gnd 0.017343f
C882 commonsourceibias.t45 gnd 0.017343f
C883 commonsourceibias.n509 gnd 0.15325f
C884 commonsourceibias.n510 gnd 0.070394f
C885 commonsourceibias.t65 gnd 0.017343f
C886 commonsourceibias.t33 gnd 0.017343f
C887 commonsourceibias.n511 gnd 0.15325f
C888 commonsourceibias.n512 gnd 0.058811f
C889 commonsourceibias.n513 gnd 0.071213f
C890 commonsourceibias.n514 gnd 0.052016f
C891 commonsourceibias.t82 gnd 0.150157f
C892 commonsourceibias.n515 gnd 0.059912f
C893 commonsourceibias.n516 gnd 0.008037f
C894 commonsourceibias.t147 gnd 0.150157f
C895 commonsourceibias.n517 gnd 0.059912f
C896 commonsourceibias.n518 gnd 0.008037f
C897 commonsourceibias.t143 gnd 0.150157f
C898 commonsourceibias.n519 gnd 0.059912f
C899 commonsourceibias.n520 gnd 0.008037f
C900 commonsourceibias.t158 gnd 0.150157f
C901 commonsourceibias.n521 gnd 0.007008f
C902 commonsourceibias.n522 gnd 0.008037f
C903 commonsourceibias.t104 gnd 0.150157f
C904 commonsourceibias.n523 gnd 0.009613f
C905 commonsourceibias.n524 gnd 0.008037f
C906 commonsourceibias.t133 gnd 0.150157f
C907 commonsourceibias.n525 gnd 0.006868f
C908 commonsourceibias.n526 gnd 0.008037f
C909 commonsourceibias.t150 gnd 0.150157f
C910 commonsourceibias.n527 gnd 0.009378f
C911 commonsourceibias.t123 gnd 0.166947f
C912 commonsourceibias.t103 gnd 0.150157f
C913 commonsourceibias.n528 gnd 0.065449f
C914 commonsourceibias.n529 gnd 0.071822f
C915 commonsourceibias.n530 gnd 0.033327f
C916 commonsourceibias.n531 gnd 0.008037f
C917 commonsourceibias.n532 gnd 0.007823f
C918 commonsourceibias.n533 gnd 0.01121f
C919 commonsourceibias.n534 gnd 0.059912f
C920 commonsourceibias.n535 gnd 0.011203f
C921 commonsourceibias.n536 gnd 0.008037f
C922 commonsourceibias.n537 gnd 0.008037f
C923 commonsourceibias.n538 gnd 0.008037f
C924 commonsourceibias.n539 gnd 0.01034f
C925 commonsourceibias.n540 gnd 0.059912f
C926 commonsourceibias.n541 gnd 0.010583f
C927 commonsourceibias.t114 gnd 0.150157f
C928 commonsourceibias.n542 gnd 0.059912f
C929 commonsourceibias.n543 gnd 0.010282f
C930 commonsourceibias.n544 gnd 0.008037f
C931 commonsourceibias.n545 gnd 0.008037f
C932 commonsourceibias.n546 gnd 0.008037f
C933 commonsourceibias.n547 gnd 0.007578f
C934 commonsourceibias.n548 gnd 0.01122f
C935 commonsourceibias.n549 gnd 0.059912f
C936 commonsourceibias.n550 gnd 0.011217f
C937 commonsourceibias.n551 gnd 0.008037f
C938 commonsourceibias.n552 gnd 0.008037f
C939 commonsourceibias.n553 gnd 0.008037f
C940 commonsourceibias.n554 gnd 0.010186f
C941 commonsourceibias.n555 gnd 0.059912f
C942 commonsourceibias.n556 gnd 0.010507f
C943 commonsourceibias.n557 gnd 0.010357f
C944 commonsourceibias.n558 gnd 0.008037f
C945 commonsourceibias.n559 gnd 0.008037f
C946 commonsourceibias.n560 gnd 0.009825f
C947 commonsourceibias.n561 gnd 0.007361f
C948 commonsourceibias.n562 gnd 0.011225f
C949 commonsourceibias.n563 gnd 0.008037f
C950 commonsourceibias.n564 gnd 0.008037f
C951 commonsourceibias.n565 gnd 0.011224f
C952 commonsourceibias.n566 gnd 0.007172f
C953 commonsourceibias.n567 gnd 0.010015f
C954 commonsourceibias.n568 gnd 0.008037f
C955 commonsourceibias.n569 gnd 0.007021f
C956 commonsourceibias.n570 gnd 0.010432f
C957 commonsourceibias.t85 gnd 0.150157f
C958 commonsourceibias.n571 gnd 0.059912f
C959 commonsourceibias.n572 gnd 0.010432f
C960 commonsourceibias.n573 gnd 0.007021f
C961 commonsourceibias.n574 gnd 0.008037f
C962 commonsourceibias.n575 gnd 0.008037f
C963 commonsourceibias.n576 gnd 0.007172f
C964 commonsourceibias.n577 gnd 0.011224f
C965 commonsourceibias.n578 gnd 0.059912f
C966 commonsourceibias.n579 gnd 0.011225f
C967 commonsourceibias.n580 gnd 0.008037f
C968 commonsourceibias.n581 gnd 0.008037f
C969 commonsourceibias.n582 gnd 0.008037f
C970 commonsourceibias.n583 gnd 0.009825f
C971 commonsourceibias.n584 gnd 0.059912f
C972 commonsourceibias.n585 gnd 0.010357f
C973 commonsourceibias.t89 gnd 0.150157f
C974 commonsourceibias.n586 gnd 0.059912f
C975 commonsourceibias.n587 gnd 0.010507f
C976 commonsourceibias.n588 gnd 0.008037f
C977 commonsourceibias.n589 gnd 0.008037f
C978 commonsourceibias.n590 gnd 0.008037f
C979 commonsourceibias.n591 gnd 0.007008f
C980 commonsourceibias.n592 gnd 0.011217f
C981 commonsourceibias.n593 gnd 0.059912f
C982 commonsourceibias.n594 gnd 0.01122f
C983 commonsourceibias.n595 gnd 0.008037f
C984 commonsourceibias.n596 gnd 0.008037f
C985 commonsourceibias.n597 gnd 0.008037f
C986 commonsourceibias.n598 gnd 0.009613f
C987 commonsourceibias.n599 gnd 0.059912f
C988 commonsourceibias.n600 gnd 0.010282f
C989 commonsourceibias.t130 gnd 0.150157f
C990 commonsourceibias.n601 gnd 0.059912f
C991 commonsourceibias.n602 gnd 0.010583f
C992 commonsourceibias.n603 gnd 0.008037f
C993 commonsourceibias.n604 gnd 0.008037f
C994 commonsourceibias.n605 gnd 0.008037f
C995 commonsourceibias.n606 gnd 0.006868f
C996 commonsourceibias.n607 gnd 0.011203f
C997 commonsourceibias.n608 gnd 0.059912f
C998 commonsourceibias.n609 gnd 0.01121f
C999 commonsourceibias.n610 gnd 0.008037f
C1000 commonsourceibias.n611 gnd 0.008037f
C1001 commonsourceibias.n612 gnd 0.008037f
C1002 commonsourceibias.n613 gnd 0.009378f
C1003 commonsourceibias.n614 gnd 0.059912f
C1004 commonsourceibias.n615 gnd 0.009861f
C1005 commonsourceibias.n616 gnd 0.07189f
C1006 commonsourceibias.n617 gnd 0.04697f
C1007 commonsourceibias.n618 gnd 0.010724f
C1008 commonsourceibias.t142 gnd 0.150157f
C1009 commonsourceibias.n619 gnd 0.007823f
C1010 commonsourceibias.n620 gnd 0.008037f
C1011 commonsourceibias.t156 gnd 0.150157f
C1012 commonsourceibias.n621 gnd 0.01034f
C1013 commonsourceibias.n622 gnd 0.008037f
C1014 commonsourceibias.t132 gnd 0.150157f
C1015 commonsourceibias.n623 gnd 0.007578f
C1016 commonsourceibias.n624 gnd 0.008037f
C1017 commonsourceibias.t149 gnd 0.150157f
C1018 commonsourceibias.n625 gnd 0.010186f
C1019 commonsourceibias.n626 gnd 0.008037f
C1020 commonsourceibias.t97 gnd 0.150157f
C1021 commonsourceibias.n627 gnd 0.007361f
C1022 commonsourceibias.n628 gnd 0.008037f
C1023 commonsourceibias.t141 gnd 0.150157f
C1024 commonsourceibias.n629 gnd 0.010015f
C1025 commonsourceibias.n630 gnd 0.008037f
C1026 commonsourceibias.t152 gnd 0.150157f
C1027 commonsourceibias.n631 gnd 0.007172f
C1028 commonsourceibias.n632 gnd 0.008037f
C1029 commonsourceibias.t131 gnd 0.150157f
C1030 commonsourceibias.n633 gnd 0.009825f
C1031 commonsourceibias.n634 gnd 0.008037f
C1032 commonsourceibias.t145 gnd 0.150157f
C1033 commonsourceibias.n635 gnd 0.007008f
C1034 commonsourceibias.n636 gnd 0.008037f
C1035 commonsourceibias.t91 gnd 0.150157f
C1036 commonsourceibias.n637 gnd 0.009613f
C1037 commonsourceibias.n638 gnd 0.008037f
C1038 commonsourceibias.t116 gnd 0.150157f
C1039 commonsourceibias.n639 gnd 0.006868f
C1040 commonsourceibias.n640 gnd 0.008037f
C1041 commonsourceibias.t134 gnd 0.150157f
C1042 commonsourceibias.n641 gnd 0.009378f
C1043 commonsourceibias.t106 gnd 0.166947f
C1044 commonsourceibias.t90 gnd 0.150157f
C1045 commonsourceibias.n642 gnd 0.065449f
C1046 commonsourceibias.n643 gnd 0.071822f
C1047 commonsourceibias.n644 gnd 0.033327f
C1048 commonsourceibias.n645 gnd 0.008037f
C1049 commonsourceibias.n646 gnd 0.007823f
C1050 commonsourceibias.n647 gnd 0.01121f
C1051 commonsourceibias.n648 gnd 0.059912f
C1052 commonsourceibias.n649 gnd 0.011203f
C1053 commonsourceibias.n650 gnd 0.008037f
C1054 commonsourceibias.n651 gnd 0.008037f
C1055 commonsourceibias.n652 gnd 0.008037f
C1056 commonsourceibias.n653 gnd 0.01034f
C1057 commonsourceibias.n654 gnd 0.059912f
C1058 commonsourceibias.n655 gnd 0.010583f
C1059 commonsourceibias.t96 gnd 0.150157f
C1060 commonsourceibias.n656 gnd 0.059912f
C1061 commonsourceibias.n657 gnd 0.010282f
C1062 commonsourceibias.n658 gnd 0.008037f
C1063 commonsourceibias.n659 gnd 0.008037f
C1064 commonsourceibias.n660 gnd 0.008037f
C1065 commonsourceibias.n661 gnd 0.007578f
C1066 commonsourceibias.n662 gnd 0.01122f
C1067 commonsourceibias.n663 gnd 0.059912f
C1068 commonsourceibias.n664 gnd 0.011217f
C1069 commonsourceibias.n665 gnd 0.008037f
C1070 commonsourceibias.n666 gnd 0.008037f
C1071 commonsourceibias.n667 gnd 0.008037f
C1072 commonsourceibias.n668 gnd 0.010186f
C1073 commonsourceibias.n669 gnd 0.059912f
C1074 commonsourceibias.n670 gnd 0.010507f
C1075 commonsourceibias.t124 gnd 0.150157f
C1076 commonsourceibias.n671 gnd 0.059912f
C1077 commonsourceibias.n672 gnd 0.010357f
C1078 commonsourceibias.n673 gnd 0.008037f
C1079 commonsourceibias.n674 gnd 0.008037f
C1080 commonsourceibias.n675 gnd 0.008037f
C1081 commonsourceibias.n676 gnd 0.007361f
C1082 commonsourceibias.n677 gnd 0.011225f
C1083 commonsourceibias.n678 gnd 0.059912f
C1084 commonsourceibias.n679 gnd 0.011224f
C1085 commonsourceibias.n680 gnd 0.008037f
C1086 commonsourceibias.n681 gnd 0.008037f
C1087 commonsourceibias.n682 gnd 0.008037f
C1088 commonsourceibias.n683 gnd 0.010015f
C1089 commonsourceibias.n684 gnd 0.059912f
C1090 commonsourceibias.n685 gnd 0.010432f
C1091 commonsourceibias.t157 gnd 0.150157f
C1092 commonsourceibias.n686 gnd 0.059912f
C1093 commonsourceibias.n687 gnd 0.010432f
C1094 commonsourceibias.n688 gnd 0.008037f
C1095 commonsourceibias.n689 gnd 0.008037f
C1096 commonsourceibias.n690 gnd 0.008037f
C1097 commonsourceibias.n691 gnd 0.007172f
C1098 commonsourceibias.n692 gnd 0.011224f
C1099 commonsourceibias.n693 gnd 0.059912f
C1100 commonsourceibias.n694 gnd 0.011225f
C1101 commonsourceibias.n695 gnd 0.008037f
C1102 commonsourceibias.n696 gnd 0.008037f
C1103 commonsourceibias.n697 gnd 0.008037f
C1104 commonsourceibias.n698 gnd 0.009825f
C1105 commonsourceibias.n699 gnd 0.059912f
C1106 commonsourceibias.n700 gnd 0.010357f
C1107 commonsourceibias.t81 gnd 0.150157f
C1108 commonsourceibias.n701 gnd 0.059912f
C1109 commonsourceibias.n702 gnd 0.010507f
C1110 commonsourceibias.n703 gnd 0.008037f
C1111 commonsourceibias.n704 gnd 0.008037f
C1112 commonsourceibias.n705 gnd 0.008037f
C1113 commonsourceibias.n706 gnd 0.007008f
C1114 commonsourceibias.n707 gnd 0.011217f
C1115 commonsourceibias.n708 gnd 0.059912f
C1116 commonsourceibias.n709 gnd 0.01122f
C1117 commonsourceibias.n710 gnd 0.008037f
C1118 commonsourceibias.n711 gnd 0.008037f
C1119 commonsourceibias.n712 gnd 0.008037f
C1120 commonsourceibias.n713 gnd 0.009613f
C1121 commonsourceibias.n714 gnd 0.059912f
C1122 commonsourceibias.n715 gnd 0.010282f
C1123 commonsourceibias.t111 gnd 0.150157f
C1124 commonsourceibias.n716 gnd 0.059912f
C1125 commonsourceibias.n717 gnd 0.010583f
C1126 commonsourceibias.n718 gnd 0.008037f
C1127 commonsourceibias.n719 gnd 0.008037f
C1128 commonsourceibias.n720 gnd 0.008037f
C1129 commonsourceibias.n721 gnd 0.006868f
C1130 commonsourceibias.n722 gnd 0.011203f
C1131 commonsourceibias.n723 gnd 0.059912f
C1132 commonsourceibias.n724 gnd 0.01121f
C1133 commonsourceibias.n725 gnd 0.008037f
C1134 commonsourceibias.n726 gnd 0.008037f
C1135 commonsourceibias.n727 gnd 0.008037f
C1136 commonsourceibias.n728 gnd 0.009378f
C1137 commonsourceibias.n729 gnd 0.059912f
C1138 commonsourceibias.n730 gnd 0.009861f
C1139 commonsourceibias.t122 gnd 0.162395f
C1140 commonsourceibias.n731 gnd 0.07189f
C1141 commonsourceibias.n732 gnd 0.025003f
C1142 commonsourceibias.n733 gnd 0.221951f
C1143 commonsourceibias.n734 gnd 4.85761f
C1144 diffpairibias.t27 gnd 0.090128f
C1145 diffpairibias.t23 gnd 0.08996f
C1146 diffpairibias.n0 gnd 0.105991f
C1147 diffpairibias.t28 gnd 0.08996f
C1148 diffpairibias.n1 gnd 0.051736f
C1149 diffpairibias.t25 gnd 0.08996f
C1150 diffpairibias.n2 gnd 0.051736f
C1151 diffpairibias.t29 gnd 0.08996f
C1152 diffpairibias.n3 gnd 0.041084f
C1153 diffpairibias.t15 gnd 0.086371f
C1154 diffpairibias.t1 gnd 0.085993f
C1155 diffpairibias.n4 gnd 0.13579f
C1156 diffpairibias.t11 gnd 0.085993f
C1157 diffpairibias.n5 gnd 0.072463f
C1158 diffpairibias.t13 gnd 0.085993f
C1159 diffpairibias.n6 gnd 0.072463f
C1160 diffpairibias.t7 gnd 0.085993f
C1161 diffpairibias.n7 gnd 0.072463f
C1162 diffpairibias.t3 gnd 0.085993f
C1163 diffpairibias.n8 gnd 0.072463f
C1164 diffpairibias.t17 gnd 0.085993f
C1165 diffpairibias.n9 gnd 0.072463f
C1166 diffpairibias.t5 gnd 0.085993f
C1167 diffpairibias.n10 gnd 0.072463f
C1168 diffpairibias.t19 gnd 0.085993f
C1169 diffpairibias.n11 gnd 0.072463f
C1170 diffpairibias.t9 gnd 0.085993f
C1171 diffpairibias.n12 gnd 0.102883f
C1172 diffpairibias.t14 gnd 0.086899f
C1173 diffpairibias.t0 gnd 0.086748f
C1174 diffpairibias.n13 gnd 0.094648f
C1175 diffpairibias.t10 gnd 0.086748f
C1176 diffpairibias.n14 gnd 0.052262f
C1177 diffpairibias.t12 gnd 0.086748f
C1178 diffpairibias.n15 gnd 0.052262f
C1179 diffpairibias.t6 gnd 0.086748f
C1180 diffpairibias.n16 gnd 0.052262f
C1181 diffpairibias.t2 gnd 0.086748f
C1182 diffpairibias.n17 gnd 0.052262f
C1183 diffpairibias.t16 gnd 0.086748f
C1184 diffpairibias.n18 gnd 0.052262f
C1185 diffpairibias.t4 gnd 0.086748f
C1186 diffpairibias.n19 gnd 0.052262f
C1187 diffpairibias.t18 gnd 0.086748f
C1188 diffpairibias.n20 gnd 0.052262f
C1189 diffpairibias.t8 gnd 0.086748f
C1190 diffpairibias.n21 gnd 0.061849f
C1191 diffpairibias.n22 gnd 0.233513f
C1192 diffpairibias.t20 gnd 0.08996f
C1193 diffpairibias.n23 gnd 0.051747f
C1194 diffpairibias.t26 gnd 0.08996f
C1195 diffpairibias.n24 gnd 0.051736f
C1196 diffpairibias.t22 gnd 0.08996f
C1197 diffpairibias.n25 gnd 0.051736f
C1198 diffpairibias.t21 gnd 0.08996f
C1199 diffpairibias.n26 gnd 0.051736f
C1200 diffpairibias.t24 gnd 0.08996f
C1201 diffpairibias.n27 gnd 0.04729f
C1202 diffpairibias.n28 gnd 0.047711f
C1203 minus.n0 gnd 0.031253f
C1204 minus.n1 gnd 0.007092f
C1205 minus.n2 gnd 0.031253f
C1206 minus.n3 gnd 0.007092f
C1207 minus.n4 gnd 0.031253f
C1208 minus.n5 gnd 0.007092f
C1209 minus.n6 gnd 0.031253f
C1210 minus.n7 gnd 0.007092f
C1211 minus.n8 gnd 0.031253f
C1212 minus.n9 gnd 0.007092f
C1213 minus.t8 gnd 0.458091f
C1214 minus.t7 gnd 0.442045f
C1215 minus.n10 gnd 0.202766f
C1216 minus.n11 gnd 0.181989f
C1217 minus.n12 gnd 0.134546f
C1218 minus.n13 gnd 0.031253f
C1219 minus.t11 gnd 0.442045f
C1220 minus.n14 gnd 0.196371f
C1221 minus.n15 gnd 0.007092f
C1222 minus.t10 gnd 0.442045f
C1223 minus.n16 gnd 0.196371f
C1224 minus.n17 gnd 0.031253f
C1225 minus.n18 gnd 0.031253f
C1226 minus.n19 gnd 0.031253f
C1227 minus.t12 gnd 0.442045f
C1228 minus.n20 gnd 0.196371f
C1229 minus.n21 gnd 0.007092f
C1230 minus.t20 gnd 0.442045f
C1231 minus.n22 gnd 0.196371f
C1232 minus.n23 gnd 0.031253f
C1233 minus.n24 gnd 0.031253f
C1234 minus.n25 gnd 0.031253f
C1235 minus.t18 gnd 0.442045f
C1236 minus.n26 gnd 0.196371f
C1237 minus.n27 gnd 0.007092f
C1238 minus.t25 gnd 0.442045f
C1239 minus.n28 gnd 0.196371f
C1240 minus.n29 gnd 0.031253f
C1241 minus.n30 gnd 0.031253f
C1242 minus.n31 gnd 0.031253f
C1243 minus.t24 gnd 0.442045f
C1244 minus.n32 gnd 0.196371f
C1245 minus.n33 gnd 0.007092f
C1246 minus.t14 gnd 0.442045f
C1247 minus.n34 gnd 0.196371f
C1248 minus.n35 gnd 0.031253f
C1249 minus.n36 gnd 0.031253f
C1250 minus.n37 gnd 0.031253f
C1251 minus.t22 gnd 0.442045f
C1252 minus.n38 gnd 0.196371f
C1253 minus.n39 gnd 0.007092f
C1254 minus.t19 gnd 0.442045f
C1255 minus.n40 gnd 0.19666f
C1256 minus.n41 gnd 0.361941f
C1257 minus.n42 gnd 0.031253f
C1258 minus.t13 gnd 0.442045f
C1259 minus.t15 gnd 0.442045f
C1260 minus.n43 gnd 0.031253f
C1261 minus.t5 gnd 0.442045f
C1262 minus.n44 gnd 0.196371f
C1263 minus.n45 gnd 0.031253f
C1264 minus.t6 gnd 0.442045f
C1265 minus.t26 gnd 0.442045f
C1266 minus.n46 gnd 0.196371f
C1267 minus.n47 gnd 0.031253f
C1268 minus.t21 gnd 0.442045f
C1269 minus.t23 gnd 0.442045f
C1270 minus.n48 gnd 0.196371f
C1271 minus.n49 gnd 0.031253f
C1272 minus.t16 gnd 0.442045f
C1273 minus.t17 gnd 0.442045f
C1274 minus.n50 gnd 0.196371f
C1275 minus.n51 gnd 0.031253f
C1276 minus.t9 gnd 0.442045f
C1277 minus.t27 gnd 0.442045f
C1278 minus.n52 gnd 0.202766f
C1279 minus.t28 gnd 0.458091f
C1280 minus.n53 gnd 0.181989f
C1281 minus.n54 gnd 0.134546f
C1282 minus.n55 gnd 0.007092f
C1283 minus.n56 gnd 0.196371f
C1284 minus.n57 gnd 0.007092f
C1285 minus.n58 gnd 0.031253f
C1286 minus.n59 gnd 0.031253f
C1287 minus.n60 gnd 0.031253f
C1288 minus.n61 gnd 0.007092f
C1289 minus.n62 gnd 0.196371f
C1290 minus.n63 gnd 0.007092f
C1291 minus.n64 gnd 0.031253f
C1292 minus.n65 gnd 0.031253f
C1293 minus.n66 gnd 0.031253f
C1294 minus.n67 gnd 0.007092f
C1295 minus.n68 gnd 0.196371f
C1296 minus.n69 gnd 0.007092f
C1297 minus.n70 gnd 0.031253f
C1298 minus.n71 gnd 0.031253f
C1299 minus.n72 gnd 0.031253f
C1300 minus.n73 gnd 0.007092f
C1301 minus.n74 gnd 0.196371f
C1302 minus.n75 gnd 0.007092f
C1303 minus.n76 gnd 0.031253f
C1304 minus.n77 gnd 0.031253f
C1305 minus.n78 gnd 0.031253f
C1306 minus.n79 gnd 0.007092f
C1307 minus.n80 gnd 0.196371f
C1308 minus.n81 gnd 0.007092f
C1309 minus.n82 gnd 0.19666f
C1310 minus.n83 gnd 1.04701f
C1311 minus.n84 gnd 1.56003f
C1312 minus.t1 gnd 0.009634f
C1313 minus.t0 gnd 0.009634f
C1314 minus.n85 gnd 0.03168f
C1315 minus.t4 gnd 0.009634f
C1316 minus.t3 gnd 0.009634f
C1317 minus.n86 gnd 0.031246f
C1318 minus.n87 gnd 0.266671f
C1319 minus.t2 gnd 0.053624f
C1320 minus.n88 gnd 0.14552f
C1321 minus.n89 gnd 2.31716f
C1322 outputibias.t10 gnd 0.11477f
C1323 outputibias.t8 gnd 0.115567f
C1324 outputibias.n0 gnd 0.130108f
C1325 outputibias.n1 gnd 0.001372f
C1326 outputibias.n2 gnd 9.76e-19
C1327 outputibias.n3 gnd 5.24e-19
C1328 outputibias.n4 gnd 0.001239f
C1329 outputibias.n5 gnd 5.55e-19
C1330 outputibias.n6 gnd 9.76e-19
C1331 outputibias.n7 gnd 5.24e-19
C1332 outputibias.n8 gnd 0.001239f
C1333 outputibias.n9 gnd 5.55e-19
C1334 outputibias.n10 gnd 0.004176f
C1335 outputibias.t5 gnd 0.00202f
C1336 outputibias.n11 gnd 9.3e-19
C1337 outputibias.n12 gnd 7.32e-19
C1338 outputibias.n13 gnd 5.24e-19
C1339 outputibias.n14 gnd 0.02322f
C1340 outputibias.n15 gnd 9.76e-19
C1341 outputibias.n16 gnd 5.24e-19
C1342 outputibias.n17 gnd 5.55e-19
C1343 outputibias.n18 gnd 0.001239f
C1344 outputibias.n19 gnd 0.001239f
C1345 outputibias.n20 gnd 5.55e-19
C1346 outputibias.n21 gnd 5.24e-19
C1347 outputibias.n22 gnd 9.76e-19
C1348 outputibias.n23 gnd 9.76e-19
C1349 outputibias.n24 gnd 5.24e-19
C1350 outputibias.n25 gnd 5.55e-19
C1351 outputibias.n26 gnd 0.001239f
C1352 outputibias.n27 gnd 0.002683f
C1353 outputibias.n28 gnd 5.55e-19
C1354 outputibias.n29 gnd 5.24e-19
C1355 outputibias.n30 gnd 0.002256f
C1356 outputibias.n31 gnd 0.005781f
C1357 outputibias.n32 gnd 0.001372f
C1358 outputibias.n33 gnd 9.76e-19
C1359 outputibias.n34 gnd 5.24e-19
C1360 outputibias.n35 gnd 0.001239f
C1361 outputibias.n36 gnd 5.55e-19
C1362 outputibias.n37 gnd 9.76e-19
C1363 outputibias.n38 gnd 5.24e-19
C1364 outputibias.n39 gnd 0.001239f
C1365 outputibias.n40 gnd 5.55e-19
C1366 outputibias.n41 gnd 0.004176f
C1367 outputibias.t3 gnd 0.00202f
C1368 outputibias.n42 gnd 9.3e-19
C1369 outputibias.n43 gnd 7.32e-19
C1370 outputibias.n44 gnd 5.24e-19
C1371 outputibias.n45 gnd 0.02322f
C1372 outputibias.n46 gnd 9.76e-19
C1373 outputibias.n47 gnd 5.24e-19
C1374 outputibias.n48 gnd 5.55e-19
C1375 outputibias.n49 gnd 0.001239f
C1376 outputibias.n50 gnd 0.001239f
C1377 outputibias.n51 gnd 5.55e-19
C1378 outputibias.n52 gnd 5.24e-19
C1379 outputibias.n53 gnd 9.76e-19
C1380 outputibias.n54 gnd 9.76e-19
C1381 outputibias.n55 gnd 5.24e-19
C1382 outputibias.n56 gnd 5.55e-19
C1383 outputibias.n57 gnd 0.001239f
C1384 outputibias.n58 gnd 0.002683f
C1385 outputibias.n59 gnd 5.55e-19
C1386 outputibias.n60 gnd 5.24e-19
C1387 outputibias.n61 gnd 0.002256f
C1388 outputibias.n62 gnd 0.005197f
C1389 outputibias.n63 gnd 0.121892f
C1390 outputibias.n64 gnd 0.001372f
C1391 outputibias.n65 gnd 9.76e-19
C1392 outputibias.n66 gnd 5.24e-19
C1393 outputibias.n67 gnd 0.001239f
C1394 outputibias.n68 gnd 5.55e-19
C1395 outputibias.n69 gnd 9.76e-19
C1396 outputibias.n70 gnd 5.24e-19
C1397 outputibias.n71 gnd 0.001239f
C1398 outputibias.n72 gnd 5.55e-19
C1399 outputibias.n73 gnd 0.004176f
C1400 outputibias.t1 gnd 0.00202f
C1401 outputibias.n74 gnd 9.3e-19
C1402 outputibias.n75 gnd 7.32e-19
C1403 outputibias.n76 gnd 5.24e-19
C1404 outputibias.n77 gnd 0.02322f
C1405 outputibias.n78 gnd 9.76e-19
C1406 outputibias.n79 gnd 5.24e-19
C1407 outputibias.n80 gnd 5.55e-19
C1408 outputibias.n81 gnd 0.001239f
C1409 outputibias.n82 gnd 0.001239f
C1410 outputibias.n83 gnd 5.55e-19
C1411 outputibias.n84 gnd 5.24e-19
C1412 outputibias.n85 gnd 9.76e-19
C1413 outputibias.n86 gnd 9.76e-19
C1414 outputibias.n87 gnd 5.24e-19
C1415 outputibias.n88 gnd 5.55e-19
C1416 outputibias.n89 gnd 0.001239f
C1417 outputibias.n90 gnd 0.002683f
C1418 outputibias.n91 gnd 5.55e-19
C1419 outputibias.n92 gnd 5.24e-19
C1420 outputibias.n93 gnd 0.002256f
C1421 outputibias.n94 gnd 0.005197f
C1422 outputibias.n95 gnd 0.064513f
C1423 outputibias.n96 gnd 0.001372f
C1424 outputibias.n97 gnd 9.76e-19
C1425 outputibias.n98 gnd 5.24e-19
C1426 outputibias.n99 gnd 0.001239f
C1427 outputibias.n100 gnd 5.55e-19
C1428 outputibias.n101 gnd 9.76e-19
C1429 outputibias.n102 gnd 5.24e-19
C1430 outputibias.n103 gnd 0.001239f
C1431 outputibias.n104 gnd 5.55e-19
C1432 outputibias.n105 gnd 0.004176f
C1433 outputibias.t7 gnd 0.00202f
C1434 outputibias.n106 gnd 9.3e-19
C1435 outputibias.n107 gnd 7.32e-19
C1436 outputibias.n108 gnd 5.24e-19
C1437 outputibias.n109 gnd 0.02322f
C1438 outputibias.n110 gnd 9.76e-19
C1439 outputibias.n111 gnd 5.24e-19
C1440 outputibias.n112 gnd 5.55e-19
C1441 outputibias.n113 gnd 0.001239f
C1442 outputibias.n114 gnd 0.001239f
C1443 outputibias.n115 gnd 5.55e-19
C1444 outputibias.n116 gnd 5.24e-19
C1445 outputibias.n117 gnd 9.76e-19
C1446 outputibias.n118 gnd 9.76e-19
C1447 outputibias.n119 gnd 5.24e-19
C1448 outputibias.n120 gnd 5.55e-19
C1449 outputibias.n121 gnd 0.001239f
C1450 outputibias.n122 gnd 0.002683f
C1451 outputibias.n123 gnd 5.55e-19
C1452 outputibias.n124 gnd 5.24e-19
C1453 outputibias.n125 gnd 0.002256f
C1454 outputibias.n126 gnd 0.005197f
C1455 outputibias.n127 gnd 0.084814f
C1456 outputibias.t6 gnd 0.108319f
C1457 outputibias.t0 gnd 0.108319f
C1458 outputibias.t2 gnd 0.108319f
C1459 outputibias.t4 gnd 0.109238f
C1460 outputibias.n128 gnd 0.134674f
C1461 outputibias.n129 gnd 0.07244f
C1462 outputibias.n130 gnd 0.079818f
C1463 outputibias.n131 gnd 0.164901f
C1464 outputibias.t11 gnd 0.11477f
C1465 outputibias.n132 gnd 0.067481f
C1466 outputibias.t9 gnd 0.11477f
C1467 outputibias.n133 gnd 0.065115f
C1468 outputibias.n134 gnd 0.029159f
C1469 a_n2472_13878.t25 gnd 0.187389f
C1470 a_n2472_13878.t21 gnd 0.187389f
C1471 a_n2472_13878.t27 gnd 0.187389f
C1472 a_n2472_13878.n0 gnd 1.47796f
C1473 a_n2472_13878.t8 gnd 0.187389f
C1474 a_n2472_13878.t18 gnd 0.187389f
C1475 a_n2472_13878.n1 gnd 1.47552f
C1476 a_n2472_13878.n2 gnd 1.32632f
C1477 a_n2472_13878.t23 gnd 0.187389f
C1478 a_n2472_13878.t15 gnd 0.187389f
C1479 a_n2472_13878.n3 gnd 1.47709f
C1480 a_n2472_13878.t20 gnd 0.187389f
C1481 a_n2472_13878.t14 gnd 0.187389f
C1482 a_n2472_13878.n4 gnd 1.47552f
C1483 a_n2472_13878.n5 gnd 2.06176f
C1484 a_n2472_13878.t10 gnd 0.187389f
C1485 a_n2472_13878.t12 gnd 0.187389f
C1486 a_n2472_13878.n6 gnd 1.47552f
C1487 a_n2472_13878.n7 gnd 1.00568f
C1488 a_n2472_13878.t22 gnd 0.187389f
C1489 a_n2472_13878.t11 gnd 0.187389f
C1490 a_n2472_13878.n8 gnd 1.47552f
C1491 a_n2472_13878.n9 gnd 1.00568f
C1492 a_n2472_13878.t19 gnd 0.187389f
C1493 a_n2472_13878.t9 gnd 0.187389f
C1494 a_n2472_13878.n10 gnd 1.47552f
C1495 a_n2472_13878.n11 gnd 4.40118f
C1496 a_n2472_13878.t1 gnd 1.75461f
C1497 a_n2472_13878.t4 gnd 0.187389f
C1498 a_n2472_13878.t5 gnd 0.187389f
C1499 a_n2472_13878.n12 gnd 1.31997f
C1500 a_n2472_13878.n13 gnd 1.47487f
C1501 a_n2472_13878.t0 gnd 1.75112f
C1502 a_n2472_13878.n14 gnd 0.742173f
C1503 a_n2472_13878.t3 gnd 1.75112f
C1504 a_n2472_13878.n15 gnd 0.742173f
C1505 a_n2472_13878.t6 gnd 0.187389f
C1506 a_n2472_13878.t7 gnd 0.187389f
C1507 a_n2472_13878.n16 gnd 1.31997f
C1508 a_n2472_13878.n17 gnd 0.749361f
C1509 a_n2472_13878.t2 gnd 1.75112f
C1510 a_n2472_13878.n18 gnd 2.43496f
C1511 a_n2472_13878.n19 gnd 3.22551f
C1512 a_n2472_13878.t24 gnd 0.187389f
C1513 a_n2472_13878.t13 gnd 0.187389f
C1514 a_n2472_13878.n20 gnd 1.47552f
C1515 a_n2472_13878.n21 gnd 2.21835f
C1516 a_n2472_13878.t16 gnd 0.187389f
C1517 a_n2472_13878.t17 gnd 0.187389f
C1518 a_n2472_13878.n22 gnd 1.47552f
C1519 a_n2472_13878.n23 gnd 0.653766f
C1520 a_n2472_13878.n24 gnd 0.653763f
C1521 a_n2472_13878.n25 gnd 1.47553f
C1522 a_n2472_13878.t26 gnd 0.187389f
C1523 a_n2650_13878.n0 gnd 3.91621f
C1524 a_n2650_13878.n1 gnd 2.8797f
C1525 a_n2650_13878.n2 gnd 3.85455f
C1526 a_n2650_13878.n3 gnd 0.812882f
C1527 a_n2650_13878.n4 gnd 0.812884f
C1528 a_n2650_13878.n5 gnd 0.796044f
C1529 a_n2650_13878.n6 gnd 0.203125f
C1530 a_n2650_13878.n7 gnd 0.149605f
C1531 a_n2650_13878.n8 gnd 0.235132f
C1532 a_n2650_13878.n9 gnd 0.181613f
C1533 a_n2650_13878.n10 gnd 0.203125f
C1534 a_n2650_13878.n11 gnd 1.22992f
C1535 a_n2650_13878.n12 gnd 0.149605f
C1536 a_n2650_13878.n13 gnd 0.849564f
C1537 a_n2650_13878.n14 gnd 0.214078f
C1538 a_n2650_13878.n15 gnd 0.690816f
C1539 a_n2650_13878.n16 gnd 0.214078f
C1540 a_n2650_13878.n17 gnd 0.498779f
C1541 a_n2650_13878.n18 gnd 0.214078f
C1542 a_n2650_13878.n19 gnd 0.552299f
C1543 a_n2650_13878.n20 gnd 0.214078f
C1544 a_n2650_13878.n21 gnd 0.886227f
C1545 a_n2650_13878.n22 gnd 0.214078f
C1546 a_n2650_13878.n23 gnd 0.926981f
C1547 a_n2650_13878.n24 gnd 0.214078f
C1548 a_n2650_13878.n25 gnd 0.498779f
C1549 a_n2650_13878.n26 gnd 0.214078f
C1550 a_n2650_13878.n27 gnd 2.96592f
C1551 a_n2650_13878.n28 gnd 0.796127f
C1552 a_n2650_13878.n29 gnd 1.16869f
C1553 a_n2650_13878.n30 gnd 1.18759f
C1554 a_n2650_13878.n31 gnd 2.2186f
C1555 a_n2650_13878.n32 gnd 1.43374f
C1556 a_n2650_13878.n33 gnd 1.18759f
C1557 a_n2650_13878.n34 gnd 1.76248f
C1558 a_n2650_13878.n35 gnd 0.44526f
C1559 a_n2650_13878.n36 gnd 0.00859f
C1560 a_n2650_13878.n37 gnd 4.14e-19
C1561 a_n2650_13878.n39 gnd 0.008288f
C1562 a_n2650_13878.n40 gnd 0.012052f
C1563 a_n2650_13878.n41 gnd 0.282797f
C1564 a_n2650_13878.n42 gnd 0.00859f
C1565 a_n2650_13878.n43 gnd 4.14e-19
C1566 a_n2650_13878.n45 gnd 0.008288f
C1567 a_n2650_13878.n46 gnd 0.012052f
C1568 a_n2650_13878.n47 gnd 0.007974f
C1569 a_n2650_13878.n48 gnd 0.282797f
C1570 a_n2650_13878.n49 gnd 0.00859f
C1571 a_n2650_13878.n50 gnd 4.14e-19
C1572 a_n2650_13878.n52 gnd 0.008288f
C1573 a_n2650_13878.n53 gnd 0.012052f
C1574 a_n2650_13878.n54 gnd 0.007974f
C1575 a_n2650_13878.n55 gnd 0.282797f
C1576 a_n2650_13878.n56 gnd 0.00859f
C1577 a_n2650_13878.n57 gnd 4.14e-19
C1578 a_n2650_13878.n59 gnd 0.008288f
C1579 a_n2650_13878.n60 gnd 0.012052f
C1580 a_n2650_13878.n61 gnd 0.007974f
C1581 a_n2650_13878.n62 gnd 0.282797f
C1582 a_n2650_13878.n63 gnd 0.008288f
C1583 a_n2650_13878.n64 gnd 0.282797f
C1584 a_n2650_13878.n65 gnd 0.008288f
C1585 a_n2650_13878.n66 gnd 0.282797f
C1586 a_n2650_13878.n67 gnd 0.008288f
C1587 a_n2650_13878.n68 gnd 0.282797f
C1588 a_n2650_13878.n69 gnd 0.008288f
C1589 a_n2650_13878.n70 gnd 0.282797f
C1590 a_n2650_13878.n71 gnd 0.007974f
C1591 a_n2650_13878.t10 gnd 0.148487f
C1592 a_n2650_13878.t29 gnd 0.69069f
C1593 a_n2650_13878.t7 gnd 0.69069f
C1594 a_n2650_13878.t25 gnd 0.69069f
C1595 a_n2650_13878.n72 gnd 0.303534f
C1596 a_n2650_13878.t27 gnd 0.69069f
C1597 a_n2650_13878.t13 gnd 0.69069f
C1598 a_n2650_13878.t3 gnd 0.69069f
C1599 a_n2650_13878.n73 gnd 0.299815f
C1600 a_n2650_13878.t9 gnd 0.69069f
C1601 a_n2650_13878.t37 gnd 0.69069f
C1602 a_n2650_13878.t98 gnd 0.69069f
C1603 a_n2650_13878.t77 gnd 0.69069f
C1604 a_n2650_13878.t82 gnd 0.69069f
C1605 a_n2650_13878.n74 gnd 0.303534f
C1606 a_n2650_13878.t71 gnd 0.69069f
C1607 a_n2650_13878.t87 gnd 0.69069f
C1608 a_n2650_13878.t95 gnd 0.69069f
C1609 a_n2650_13878.n75 gnd 0.299815f
C1610 a_n2650_13878.t96 gnd 0.69069f
C1611 a_n2650_13878.t66 gnd 0.69069f
C1612 a_n2650_13878.t79 gnd 0.69069f
C1613 a_n2650_13878.n76 gnd 0.303656f
C1614 a_n2650_13878.t36 gnd 1.39036f
C1615 a_n2650_13878.t12 gnd 0.148487f
C1616 a_n2650_13878.t20 gnd 0.148487f
C1617 a_n2650_13878.n77 gnd 1.04594f
C1618 a_n2650_13878.t24 gnd 0.148487f
C1619 a_n2650_13878.t42 gnd 0.148487f
C1620 a_n2650_13878.n78 gnd 1.04594f
C1621 a_n2650_13878.t6 gnd 0.148487f
C1622 a_n2650_13878.t22 gnd 0.148487f
C1623 a_n2650_13878.n79 gnd 1.04594f
C1624 a_n2650_13878.t16 gnd 0.148487f
C1625 a_n2650_13878.t40 gnd 0.148487f
C1626 a_n2650_13878.n80 gnd 1.04594f
C1627 a_n2650_13878.t32 gnd 1.38758f
C1628 a_n2650_13878.t15 gnd 0.69069f
C1629 a_n2650_13878.n81 gnd 0.300072f
C1630 a_n2650_13878.t5 gnd 0.69069f
C1631 a_n2650_13878.t19 gnd 0.69069f
C1632 a_n2650_13878.n82 gnd 0.303534f
C1633 a_n2650_13878.t35 gnd 0.69069f
C1634 a_n2650_13878.t76 gnd 0.69069f
C1635 a_n2650_13878.n83 gnd 0.300072f
C1636 a_n2650_13878.t91 gnd 0.69069f
C1637 a_n2650_13878.t94 gnd 0.69069f
C1638 a_n2650_13878.n84 gnd 0.303534f
C1639 a_n2650_13878.t70 gnd 0.69069f
C1640 a_n2650_13878.n85 gnd 0.29437f
C1641 a_n2650_13878.t93 gnd 0.69069f
C1642 a_n2650_13878.n86 gnd 0.299485f
C1643 a_n2650_13878.t68 gnd 0.69069f
C1644 a_n2650_13878.n87 gnd 0.306266f
C1645 a_n2650_13878.t90 gnd 0.69069f
C1646 a_n2650_13878.n88 gnd 0.303671f
C1647 a_n2650_13878.n89 gnd 0.299815f
C1648 a_n2650_13878.t65 gnd 0.69069f
C1649 a_n2650_13878.n90 gnd 0.294535f
C1650 a_n2650_13878.t85 gnd 0.69069f
C1651 a_n2650_13878.n91 gnd 0.303656f
C1652 a_n2650_13878.t67 gnd 0.702263f
C1653 a_n2650_13878.n92 gnd 0.29437f
C1654 a_n2650_13878.t11 gnd 0.69069f
C1655 a_n2650_13878.n93 gnd 0.299485f
C1656 a_n2650_13878.t23 gnd 0.69069f
C1657 a_n2650_13878.n94 gnd 0.306266f
C1658 a_n2650_13878.t41 gnd 0.69069f
C1659 a_n2650_13878.n95 gnd 0.303671f
C1660 a_n2650_13878.n96 gnd 0.299815f
C1661 a_n2650_13878.t21 gnd 0.69069f
C1662 a_n2650_13878.n97 gnd 0.294535f
C1663 a_n2650_13878.t39 gnd 0.69069f
C1664 a_n2650_13878.n98 gnd 0.303656f
C1665 a_n2650_13878.t31 gnd 0.702263f
C1666 a_n2650_13878.n99 gnd 1.26233f
C1667 a_n2650_13878.t74 gnd 0.69069f
C1668 a_n2650_13878.n100 gnd 0.299815f
C1669 a_n2650_13878.t81 gnd 0.69069f
C1670 a_n2650_13878.n101 gnd 0.299815f
C1671 a_n2650_13878.t72 gnd 0.69069f
C1672 a_n2650_13878.n102 gnd 0.299815f
C1673 a_n2650_13878.t86 gnd 0.69069f
C1674 a_n2650_13878.n103 gnd 0.299815f
C1675 a_n2650_13878.t75 gnd 0.69069f
C1676 a_n2650_13878.n104 gnd 0.29437f
C1677 a_n2650_13878.t99 gnd 0.69069f
C1678 a_n2650_13878.n105 gnd 0.303671f
C1679 a_n2650_13878.t78 gnd 0.702263f
C1680 a_n2650_13878.t88 gnd 0.69069f
C1681 a_n2650_13878.n106 gnd 0.29437f
C1682 a_n2650_13878.t73 gnd 0.69069f
C1683 a_n2650_13878.n107 gnd 0.303671f
C1684 a_n2650_13878.t83 gnd 0.702263f
C1685 a_n2650_13878.t92 gnd 0.69069f
C1686 a_n2650_13878.n108 gnd 0.29437f
C1687 a_n2650_13878.t80 gnd 0.69069f
C1688 a_n2650_13878.n109 gnd 0.303671f
C1689 a_n2650_13878.t97 gnd 0.702263f
C1690 a_n2650_13878.t84 gnd 0.69069f
C1691 a_n2650_13878.n110 gnd 0.29437f
C1692 a_n2650_13878.t64 gnd 0.69069f
C1693 a_n2650_13878.n111 gnd 0.303671f
C1694 a_n2650_13878.t89 gnd 0.702263f
C1695 a_n2650_13878.n112 gnd 1.55896f
C1696 a_n2650_13878.t69 gnd 0.702263f
C1697 a_n2650_13878.n113 gnd 0.300072f
C1698 a_n2650_13878.n114 gnd 0.294535f
C1699 a_n2650_13878.n115 gnd 0.303671f
C1700 a_n2650_13878.n116 gnd 0.306266f
C1701 a_n2650_13878.n117 gnd 0.299485f
C1702 a_n2650_13878.n118 gnd 0.29437f
C1703 a_n2650_13878.t17 gnd 0.702263f
C1704 a_n2650_13878.t33 gnd 0.69069f
C1705 a_n2650_13878.n119 gnd 0.303656f
C1706 a_n2650_13878.t47 gnd 0.11549f
C1707 a_n2650_13878.t1 gnd 0.11549f
C1708 a_n2650_13878.n120 gnd 1.02278f
C1709 a_n2650_13878.t57 gnd 0.11549f
C1710 a_n2650_13878.t60 gnd 0.11549f
C1711 a_n2650_13878.n121 gnd 1.02051f
C1712 a_n2650_13878.t49 gnd 0.11549f
C1713 a_n2650_13878.t56 gnd 0.11549f
C1714 a_n2650_13878.n122 gnd 1.02051f
C1715 a_n2650_13878.t59 gnd 0.11549f
C1716 a_n2650_13878.t62 gnd 0.11549f
C1717 a_n2650_13878.n123 gnd 1.02278f
C1718 a_n2650_13878.t58 gnd 0.11549f
C1719 a_n2650_13878.t45 gnd 0.11549f
C1720 a_n2650_13878.n124 gnd 1.02051f
C1721 a_n2650_13878.t51 gnd 0.11549f
C1722 a_n2650_13878.t55 gnd 0.11549f
C1723 a_n2650_13878.n125 gnd 1.02051f
C1724 a_n2650_13878.t44 gnd 0.11549f
C1725 a_n2650_13878.t50 gnd 0.11549f
C1726 a_n2650_13878.n126 gnd 1.02051f
C1727 a_n2650_13878.t2 gnd 0.11549f
C1728 a_n2650_13878.t0 gnd 0.11549f
C1729 a_n2650_13878.n127 gnd 1.02051f
C1730 a_n2650_13878.t48 gnd 0.11549f
C1731 a_n2650_13878.t52 gnd 0.11549f
C1732 a_n2650_13878.n128 gnd 1.02051f
C1733 a_n2650_13878.t53 gnd 0.11549f
C1734 a_n2650_13878.t54 gnd 0.11549f
C1735 a_n2650_13878.n129 gnd 1.02278f
C1736 a_n2650_13878.t43 gnd 0.11549f
C1737 a_n2650_13878.t63 gnd 0.11549f
C1738 a_n2650_13878.n130 gnd 1.02051f
C1739 a_n2650_13878.t61 gnd 0.11549f
C1740 a_n2650_13878.t46 gnd 0.11549f
C1741 a_n2650_13878.n131 gnd 1.02051f
C1742 a_n2650_13878.n132 gnd 0.300072f
C1743 a_n2650_13878.n133 gnd 0.294535f
C1744 a_n2650_13878.n134 gnd 0.303671f
C1745 a_n2650_13878.n135 gnd 0.306266f
C1746 a_n2650_13878.n136 gnd 0.299485f
C1747 a_n2650_13878.n137 gnd 0.29437f
C1748 a_n2650_13878.n138 gnd 0.933405f
C1749 a_n2650_13878.t30 gnd 1.38759f
C1750 a_n2650_13878.t8 gnd 0.148487f
C1751 a_n2650_13878.t26 gnd 0.148487f
C1752 a_n2650_13878.n139 gnd 1.04594f
C1753 a_n2650_13878.t28 gnd 0.148487f
C1754 a_n2650_13878.t14 gnd 0.148487f
C1755 a_n2650_13878.n140 gnd 1.04594f
C1756 a_n2650_13878.t18 gnd 1.39036f
C1757 a_n2650_13878.t38 gnd 0.148487f
C1758 a_n2650_13878.t34 gnd 0.148487f
C1759 a_n2650_13878.n141 gnd 1.04594f
C1760 a_n2650_13878.n142 gnd 1.04595f
C1761 a_n2650_13878.t4 gnd 0.148487f
C1762 CSoutput.n0 gnd 0.044617f
C1763 CSoutput.t193 gnd 0.295134f
C1764 CSoutput.n1 gnd 0.133268f
C1765 CSoutput.n2 gnd 0.044617f
C1766 CSoutput.t176 gnd 0.295134f
C1767 CSoutput.n3 gnd 0.035363f
C1768 CSoutput.n4 gnd 0.044617f
C1769 CSoutput.t185 gnd 0.295134f
C1770 CSoutput.n5 gnd 0.030494f
C1771 CSoutput.n6 gnd 0.044617f
C1772 CSoutput.t196 gnd 0.295134f
C1773 CSoutput.t195 gnd 0.295134f
C1774 CSoutput.n7 gnd 0.131815f
C1775 CSoutput.n8 gnd 0.044617f
C1776 CSoutput.t182 gnd 0.295134f
C1777 CSoutput.n9 gnd 0.029074f
C1778 CSoutput.n10 gnd 0.044617f
C1779 CSoutput.t188 gnd 0.295134f
C1780 CSoutput.t191 gnd 0.295134f
C1781 CSoutput.n11 gnd 0.131815f
C1782 CSoutput.n12 gnd 0.044617f
C1783 CSoutput.t179 gnd 0.295134f
C1784 CSoutput.n13 gnd 0.030494f
C1785 CSoutput.n14 gnd 0.044617f
C1786 CSoutput.t178 gnd 0.295134f
C1787 CSoutput.t189 gnd 0.295134f
C1788 CSoutput.n15 gnd 0.131815f
C1789 CSoutput.n16 gnd 0.044617f
C1790 CSoutput.t194 gnd 0.295134f
C1791 CSoutput.n17 gnd 0.032569f
C1792 CSoutput.t180 gnd 0.352693f
C1793 CSoutput.t177 gnd 0.295134f
C1794 CSoutput.n18 gnd 0.168277f
C1795 CSoutput.n19 gnd 0.163287f
C1796 CSoutput.n20 gnd 0.189432f
C1797 CSoutput.n21 gnd 0.044617f
C1798 CSoutput.n22 gnd 0.037238f
C1799 CSoutput.n23 gnd 0.131815f
C1800 CSoutput.n24 gnd 0.035896f
C1801 CSoutput.n25 gnd 0.035363f
C1802 CSoutput.n26 gnd 0.044617f
C1803 CSoutput.n27 gnd 0.044617f
C1804 CSoutput.n28 gnd 0.036952f
C1805 CSoutput.n29 gnd 0.031373f
C1806 CSoutput.n30 gnd 0.13475f
C1807 CSoutput.n31 gnd 0.031805f
C1808 CSoutput.n32 gnd 0.044617f
C1809 CSoutput.n33 gnd 0.044617f
C1810 CSoutput.n34 gnd 0.044617f
C1811 CSoutput.n35 gnd 0.036558f
C1812 CSoutput.n36 gnd 0.131815f
C1813 CSoutput.n37 gnd 0.034963f
C1814 CSoutput.n38 gnd 0.036297f
C1815 CSoutput.n39 gnd 0.044617f
C1816 CSoutput.n40 gnd 0.044617f
C1817 CSoutput.n41 gnd 0.03723f
C1818 CSoutput.n42 gnd 0.034029f
C1819 CSoutput.n43 gnd 0.131815f
C1820 CSoutput.n44 gnd 0.034891f
C1821 CSoutput.n45 gnd 0.044617f
C1822 CSoutput.n46 gnd 0.044617f
C1823 CSoutput.n47 gnd 0.044617f
C1824 CSoutput.n48 gnd 0.034891f
C1825 CSoutput.n49 gnd 0.131815f
C1826 CSoutput.n50 gnd 0.034029f
C1827 CSoutput.n51 gnd 0.03723f
C1828 CSoutput.n52 gnd 0.044617f
C1829 CSoutput.n53 gnd 0.044617f
C1830 CSoutput.n54 gnd 0.036297f
C1831 CSoutput.n55 gnd 0.034963f
C1832 CSoutput.n56 gnd 0.131815f
C1833 CSoutput.n57 gnd 0.036558f
C1834 CSoutput.n58 gnd 0.044617f
C1835 CSoutput.n59 gnd 0.044617f
C1836 CSoutput.n60 gnd 0.044617f
C1837 CSoutput.n61 gnd 0.031805f
C1838 CSoutput.n62 gnd 0.13475f
C1839 CSoutput.n63 gnd 0.031373f
C1840 CSoutput.t197 gnd 0.295134f
C1841 CSoutput.n64 gnd 0.131815f
C1842 CSoutput.n65 gnd 0.036952f
C1843 CSoutput.n66 gnd 0.044617f
C1844 CSoutput.n67 gnd 0.044617f
C1845 CSoutput.n68 gnd 0.044617f
C1846 CSoutput.n69 gnd 0.035896f
C1847 CSoutput.n70 gnd 0.131815f
C1848 CSoutput.n71 gnd 0.037238f
C1849 CSoutput.n72 gnd 0.032569f
C1850 CSoutput.n73 gnd 0.044617f
C1851 CSoutput.n74 gnd 0.044617f
C1852 CSoutput.n75 gnd 0.033776f
C1853 CSoutput.n76 gnd 0.02006f
C1854 CSoutput.t183 gnd 0.331604f
C1855 CSoutput.n77 gnd 0.164727f
C1856 CSoutput.n78 gnd 0.704854f
C1857 CSoutput.t8 gnd 0.055654f
C1858 CSoutput.t57 gnd 0.055654f
C1859 CSoutput.n79 gnd 0.43089f
C1860 CSoutput.t14 gnd 0.055654f
C1861 CSoutput.t37 gnd 0.055654f
C1862 CSoutput.n80 gnd 0.430122f
C1863 CSoutput.n81 gnd 0.436573f
C1864 CSoutput.t96 gnd 0.055654f
C1865 CSoutput.t51 gnd 0.055654f
C1866 CSoutput.n82 gnd 0.430122f
C1867 CSoutput.n83 gnd 0.215125f
C1868 CSoutput.t16 gnd 0.055654f
C1869 CSoutput.t83 gnd 0.055654f
C1870 CSoutput.n84 gnd 0.430122f
C1871 CSoutput.n85 gnd 0.215125f
C1872 CSoutput.t23 gnd 0.055654f
C1873 CSoutput.t66 gnd 0.055654f
C1874 CSoutput.n86 gnd 0.430122f
C1875 CSoutput.n87 gnd 0.215125f
C1876 CSoutput.t41 gnd 0.055654f
C1877 CSoutput.t58 gnd 0.055654f
C1878 CSoutput.n88 gnd 0.430122f
C1879 CSoutput.n89 gnd 0.215125f
C1880 CSoutput.t54 gnd 0.055654f
C1881 CSoutput.t88 gnd 0.055654f
C1882 CSoutput.n90 gnd 0.430122f
C1883 CSoutput.n91 gnd 0.215125f
C1884 CSoutput.t30 gnd 0.055654f
C1885 CSoutput.t71 gnd 0.055654f
C1886 CSoutput.n92 gnd 0.430122f
C1887 CSoutput.n93 gnd 0.394489f
C1888 CSoutput.t26 gnd 0.055654f
C1889 CSoutput.t89 gnd 0.055654f
C1890 CSoutput.n94 gnd 0.43089f
C1891 CSoutput.t64 gnd 0.055654f
C1892 CSoutput.t63 gnd 0.055654f
C1893 CSoutput.n95 gnd 0.430122f
C1894 CSoutput.n96 gnd 0.436573f
C1895 CSoutput.t55 gnd 0.055654f
C1896 CSoutput.t24 gnd 0.055654f
C1897 CSoutput.n97 gnd 0.430122f
C1898 CSoutput.n98 gnd 0.215125f
C1899 CSoutput.t7 gnd 0.055654f
C1900 CSoutput.t56 gnd 0.055654f
C1901 CSoutput.n99 gnd 0.430122f
C1902 CSoutput.n100 gnd 0.215125f
C1903 CSoutput.t52 gnd 0.055654f
C1904 CSoutput.t22 gnd 0.055654f
C1905 CSoutput.n101 gnd 0.430122f
C1906 CSoutput.n102 gnd 0.215125f
C1907 CSoutput.t5 gnd 0.055654f
C1908 CSoutput.t3 gnd 0.055654f
C1909 CSoutput.n103 gnd 0.430122f
C1910 CSoutput.n104 gnd 0.215125f
C1911 CSoutput.t67 gnd 0.055654f
C1912 CSoutput.t38 gnd 0.055654f
C1913 CSoutput.n105 gnd 0.430122f
C1914 CSoutput.n106 gnd 0.215125f
C1915 CSoutput.t32 gnd 0.055654f
C1916 CSoutput.t2 gnd 0.055654f
C1917 CSoutput.n107 gnd 0.430122f
C1918 CSoutput.n108 gnd 0.320805f
C1919 CSoutput.n109 gnd 0.404533f
C1920 CSoutput.t42 gnd 0.055654f
C1921 CSoutput.t97 gnd 0.055654f
C1922 CSoutput.n110 gnd 0.43089f
C1923 CSoutput.t74 gnd 0.055654f
C1924 CSoutput.t73 gnd 0.055654f
C1925 CSoutput.n111 gnd 0.430122f
C1926 CSoutput.n112 gnd 0.436573f
C1927 CSoutput.t61 gnd 0.055654f
C1928 CSoutput.t39 gnd 0.055654f
C1929 CSoutput.n113 gnd 0.430122f
C1930 CSoutput.n114 gnd 0.215125f
C1931 CSoutput.t19 gnd 0.055654f
C1932 CSoutput.t62 gnd 0.055654f
C1933 CSoutput.n115 gnd 0.430122f
C1934 CSoutput.n116 gnd 0.215125f
C1935 CSoutput.t60 gnd 0.055654f
C1936 CSoutput.t36 gnd 0.055654f
C1937 CSoutput.n117 gnd 0.430122f
C1938 CSoutput.n118 gnd 0.215125f
C1939 CSoutput.t18 gnd 0.055654f
C1940 CSoutput.t17 gnd 0.055654f
C1941 CSoutput.n119 gnd 0.430122f
C1942 CSoutput.n120 gnd 0.215125f
C1943 CSoutput.t75 gnd 0.055654f
C1944 CSoutput.t48 gnd 0.055654f
C1945 CSoutput.n121 gnd 0.430122f
C1946 CSoutput.n122 gnd 0.215125f
C1947 CSoutput.t45 gnd 0.055654f
C1948 CSoutput.t13 gnd 0.055654f
C1949 CSoutput.n123 gnd 0.430122f
C1950 CSoutput.n124 gnd 0.320805f
C1951 CSoutput.n125 gnd 0.452165f
C1952 CSoutput.n126 gnd 9.49187f
C1953 CSoutput.n128 gnd 0.789272f
C1954 CSoutput.n129 gnd 0.591954f
C1955 CSoutput.n130 gnd 0.789272f
C1956 CSoutput.n131 gnd 0.789272f
C1957 CSoutput.n132 gnd 2.12496f
C1958 CSoutput.n133 gnd 0.789272f
C1959 CSoutput.n134 gnd 0.789272f
C1960 CSoutput.t187 gnd 0.98659f
C1961 CSoutput.n135 gnd 0.789272f
C1962 CSoutput.n136 gnd 0.789272f
C1963 CSoutput.n140 gnd 0.789272f
C1964 CSoutput.n144 gnd 0.789272f
C1965 CSoutput.n145 gnd 0.789272f
C1966 CSoutput.n147 gnd 0.789272f
C1967 CSoutput.n152 gnd 0.789272f
C1968 CSoutput.n154 gnd 0.789272f
C1969 CSoutput.n155 gnd 0.789272f
C1970 CSoutput.n157 gnd 0.789272f
C1971 CSoutput.n158 gnd 0.789272f
C1972 CSoutput.n160 gnd 0.789272f
C1973 CSoutput.t181 gnd 13.1886f
C1974 CSoutput.n162 gnd 0.789272f
C1975 CSoutput.n163 gnd 0.591954f
C1976 CSoutput.n164 gnd 0.789272f
C1977 CSoutput.n165 gnd 0.789272f
C1978 CSoutput.n166 gnd 2.12496f
C1979 CSoutput.n167 gnd 0.789272f
C1980 CSoutput.n168 gnd 0.789272f
C1981 CSoutput.t184 gnd 0.98659f
C1982 CSoutput.n169 gnd 0.789272f
C1983 CSoutput.n170 gnd 0.789272f
C1984 CSoutput.n174 gnd 0.789272f
C1985 CSoutput.n178 gnd 0.789272f
C1986 CSoutput.n179 gnd 0.789272f
C1987 CSoutput.n181 gnd 0.789272f
C1988 CSoutput.n186 gnd 0.789272f
C1989 CSoutput.n188 gnd 0.789272f
C1990 CSoutput.n189 gnd 0.789272f
C1991 CSoutput.n191 gnd 0.789272f
C1992 CSoutput.n192 gnd 0.789272f
C1993 CSoutput.n194 gnd 0.789272f
C1994 CSoutput.n195 gnd 0.591954f
C1995 CSoutput.n197 gnd 0.789272f
C1996 CSoutput.n198 gnd 0.591954f
C1997 CSoutput.n199 gnd 0.789272f
C1998 CSoutput.n200 gnd 0.789272f
C1999 CSoutput.n201 gnd 2.12496f
C2000 CSoutput.n202 gnd 0.789272f
C2001 CSoutput.n203 gnd 0.789272f
C2002 CSoutput.t186 gnd 0.98659f
C2003 CSoutput.n204 gnd 0.789272f
C2004 CSoutput.n205 gnd 2.12496f
C2005 CSoutput.n207 gnd 0.789272f
C2006 CSoutput.n208 gnd 0.789272f
C2007 CSoutput.n210 gnd 0.789272f
C2008 CSoutput.n211 gnd 0.789272f
C2009 CSoutput.t192 gnd 12.973701f
C2010 CSoutput.t190 gnd 13.1886f
C2011 CSoutput.n217 gnd 2.47606f
C2012 CSoutput.n218 gnd 10.086599f
C2013 CSoutput.n219 gnd 10.5086f
C2014 CSoutput.n224 gnd 2.68224f
C2015 CSoutput.n230 gnd 0.789272f
C2016 CSoutput.n232 gnd 0.789272f
C2017 CSoutput.n234 gnd 0.789272f
C2018 CSoutput.n236 gnd 0.789272f
C2019 CSoutput.n238 gnd 0.789272f
C2020 CSoutput.n244 gnd 0.789272f
C2021 CSoutput.n251 gnd 1.44801f
C2022 CSoutput.n252 gnd 1.44801f
C2023 CSoutput.n253 gnd 0.789272f
C2024 CSoutput.n254 gnd 0.789272f
C2025 CSoutput.n256 gnd 0.591954f
C2026 CSoutput.n257 gnd 0.506956f
C2027 CSoutput.n259 gnd 0.591954f
C2028 CSoutput.n260 gnd 0.506956f
C2029 CSoutput.n261 gnd 0.591954f
C2030 CSoutput.n263 gnd 0.789272f
C2031 CSoutput.n265 gnd 2.12496f
C2032 CSoutput.n266 gnd 2.47606f
C2033 CSoutput.n267 gnd 9.27706f
C2034 CSoutput.n269 gnd 0.591954f
C2035 CSoutput.n270 gnd 1.52313f
C2036 CSoutput.n271 gnd 0.591954f
C2037 CSoutput.n273 gnd 0.789272f
C2038 CSoutput.n275 gnd 2.12496f
C2039 CSoutput.n276 gnd 4.62851f
C2040 CSoutput.t76 gnd 0.055654f
C2041 CSoutput.t6 gnd 0.055654f
C2042 CSoutput.n277 gnd 0.43089f
C2043 CSoutput.t35 gnd 0.055654f
C2044 CSoutput.t12 gnd 0.055654f
C2045 CSoutput.n278 gnd 0.430122f
C2046 CSoutput.n279 gnd 0.436573f
C2047 CSoutput.t50 gnd 0.055654f
C2048 CSoutput.t29 gnd 0.055654f
C2049 CSoutput.n280 gnd 0.430122f
C2050 CSoutput.n281 gnd 0.215125f
C2051 CSoutput.t82 gnd 0.055654f
C2052 CSoutput.t15 gnd 0.055654f
C2053 CSoutput.n282 gnd 0.430122f
C2054 CSoutput.n283 gnd 0.215125f
C2055 CSoutput.t65 gnd 0.055654f
C2056 CSoutput.t20 gnd 0.055654f
C2057 CSoutput.n284 gnd 0.430122f
C2058 CSoutput.n285 gnd 0.215125f
C2059 CSoutput.t78 gnd 0.055654f
C2060 CSoutput.t40 gnd 0.055654f
C2061 CSoutput.n286 gnd 0.430122f
C2062 CSoutput.n287 gnd 0.215125f
C2063 CSoutput.t87 gnd 0.055654f
C2064 CSoutput.t53 gnd 0.055654f
C2065 CSoutput.n288 gnd 0.430122f
C2066 CSoutput.n289 gnd 0.215125f
C2067 CSoutput.t70 gnd 0.055654f
C2068 CSoutput.t31 gnd 0.055654f
C2069 CSoutput.n290 gnd 0.430122f
C2070 CSoutput.n291 gnd 0.394489f
C2071 CSoutput.t34 gnd 0.055654f
C2072 CSoutput.t86 gnd 0.055654f
C2073 CSoutput.n292 gnd 0.43089f
C2074 CSoutput.t27 gnd 0.055654f
C2075 CSoutput.t28 gnd 0.055654f
C2076 CSoutput.n293 gnd 0.430122f
C2077 CSoutput.n294 gnd 0.436573f
C2078 CSoutput.t84 gnd 0.055654f
C2079 CSoutput.t85 gnd 0.055654f
C2080 CSoutput.n295 gnd 0.430122f
C2081 CSoutput.n296 gnd 0.215125f
C2082 CSoutput.t11 gnd 0.055654f
C2083 CSoutput.t72 gnd 0.055654f
C2084 CSoutput.n297 gnd 0.430122f
C2085 CSoutput.n298 gnd 0.215125f
C2086 CSoutput.t81 gnd 0.055654f
C2087 CSoutput.t9 gnd 0.055654f
C2088 CSoutput.n299 gnd 0.430122f
C2089 CSoutput.n300 gnd 0.215125f
C2090 CSoutput.t49 gnd 0.055654f
C2091 CSoutput.t69 gnd 0.055654f
C2092 CSoutput.n301 gnd 0.430122f
C2093 CSoutput.n302 gnd 0.215125f
C2094 CSoutput.t91 gnd 0.055654f
C2095 CSoutput.t33 gnd 0.055654f
C2096 CSoutput.n303 gnd 0.430122f
C2097 CSoutput.n304 gnd 0.215125f
C2098 CSoutput.t68 gnd 0.055654f
C2099 CSoutput.t95 gnd 0.055654f
C2100 CSoutput.n305 gnd 0.430122f
C2101 CSoutput.n306 gnd 0.320805f
C2102 CSoutput.n307 gnd 0.404533f
C2103 CSoutput.t47 gnd 0.055654f
C2104 CSoutput.t94 gnd 0.055654f
C2105 CSoutput.n308 gnd 0.43089f
C2106 CSoutput.t43 gnd 0.055654f
C2107 CSoutput.t44 gnd 0.055654f
C2108 CSoutput.n309 gnd 0.430122f
C2109 CSoutput.n310 gnd 0.436573f
C2110 CSoutput.t92 gnd 0.055654f
C2111 CSoutput.t93 gnd 0.055654f
C2112 CSoutput.n311 gnd 0.430122f
C2113 CSoutput.n312 gnd 0.215125f
C2114 CSoutput.t25 gnd 0.055654f
C2115 CSoutput.t80 gnd 0.055654f
C2116 CSoutput.n313 gnd 0.430122f
C2117 CSoutput.n314 gnd 0.215125f
C2118 CSoutput.t90 gnd 0.055654f
C2119 CSoutput.t21 gnd 0.055654f
C2120 CSoutput.n315 gnd 0.430122f
C2121 CSoutput.n316 gnd 0.215125f
C2122 CSoutput.t59 gnd 0.055654f
C2123 CSoutput.t79 gnd 0.055654f
C2124 CSoutput.n317 gnd 0.430122f
C2125 CSoutput.n318 gnd 0.215125f
C2126 CSoutput.t4 gnd 0.055654f
C2127 CSoutput.t46 gnd 0.055654f
C2128 CSoutput.n319 gnd 0.430122f
C2129 CSoutput.n320 gnd 0.215125f
C2130 CSoutput.t77 gnd 0.055654f
C2131 CSoutput.t10 gnd 0.055654f
C2132 CSoutput.n321 gnd 0.43012f
C2133 CSoutput.n322 gnd 0.320807f
C2134 CSoutput.n323 gnd 0.452165f
C2135 CSoutput.n324 gnd 13.0472f
C2136 CSoutput.t129 gnd 0.048697f
C2137 CSoutput.t146 gnd 0.048697f
C2138 CSoutput.n325 gnd 0.431745f
C2139 CSoutput.t125 gnd 0.048697f
C2140 CSoutput.t153 gnd 0.048697f
C2141 CSoutput.n326 gnd 0.430304f
C2142 CSoutput.n327 gnd 0.400963f
C2143 CSoutput.t160 gnd 0.048697f
C2144 CSoutput.t99 gnd 0.048697f
C2145 CSoutput.n328 gnd 0.430304f
C2146 CSoutput.n329 gnd 0.197656f
C2147 CSoutput.t133 gnd 0.048697f
C2148 CSoutput.t156 gnd 0.048697f
C2149 CSoutput.n330 gnd 0.430304f
C2150 CSoutput.n331 gnd 0.197656f
C2151 CSoutput.t166 gnd 0.048697f
C2152 CSoutput.t123 gnd 0.048697f
C2153 CSoutput.n332 gnd 0.430304f
C2154 CSoutput.n333 gnd 0.197656f
C2155 CSoutput.t158 gnd 0.048697f
C2156 CSoutput.t147 gnd 0.048697f
C2157 CSoutput.n334 gnd 0.430304f
C2158 CSoutput.n335 gnd 0.197656f
C2159 CSoutput.t162 gnd 0.048697f
C2160 CSoutput.t102 gnd 0.048697f
C2161 CSoutput.n336 gnd 0.430304f
C2162 CSoutput.n337 gnd 0.197656f
C2163 CSoutput.t150 gnd 0.048697f
C2164 CSoutput.t115 gnd 0.048697f
C2165 CSoutput.n338 gnd 0.430304f
C2166 CSoutput.n339 gnd 0.197656f
C2167 CSoutput.t173 gnd 0.048697f
C2168 CSoutput.t121 gnd 0.048697f
C2169 CSoutput.n340 gnd 0.430304f
C2170 CSoutput.n341 gnd 0.197656f
C2171 CSoutput.t134 gnd 0.048697f
C2172 CSoutput.t149 gnd 0.048697f
C2173 CSoutput.n342 gnd 0.430304f
C2174 CSoutput.n343 gnd 0.364518f
C2175 CSoutput.t117 gnd 0.048697f
C2176 CSoutput.t111 gnd 0.048697f
C2177 CSoutput.n344 gnd 0.431745f
C2178 CSoutput.t98 gnd 0.048697f
C2179 CSoutput.t119 gnd 0.048697f
C2180 CSoutput.n345 gnd 0.430304f
C2181 CSoutput.n346 gnd 0.400963f
C2182 CSoutput.t107 gnd 0.048697f
C2183 CSoutput.t103 gnd 0.048697f
C2184 CSoutput.n347 gnd 0.430304f
C2185 CSoutput.n348 gnd 0.197656f
C2186 CSoutput.t137 gnd 0.048697f
C2187 CSoutput.t105 gnd 0.048697f
C2188 CSoutput.n349 gnd 0.430304f
C2189 CSoutput.n350 gnd 0.197656f
C2190 CSoutput.t106 gnd 0.048697f
C2191 CSoutput.t145 gnd 0.048697f
C2192 CSoutput.n351 gnd 0.430304f
C2193 CSoutput.n352 gnd 0.197656f
C2194 CSoutput.t168 gnd 0.048697f
C2195 CSoutput.t152 gnd 0.048697f
C2196 CSoutput.n353 gnd 0.430304f
C2197 CSoutput.n354 gnd 0.197656f
C2198 CSoutput.t116 gnd 0.048697f
C2199 CSoutput.t110 gnd 0.048697f
C2200 CSoutput.n355 gnd 0.430304f
C2201 CSoutput.n356 gnd 0.197656f
C2202 CSoutput.t157 gnd 0.048697f
C2203 CSoutput.t120 gnd 0.048697f
C2204 CSoutput.n357 gnd 0.430304f
C2205 CSoutput.n358 gnd 0.197656f
C2206 CSoutput.t114 gnd 0.048697f
C2207 CSoutput.t1 gnd 0.048697f
C2208 CSoutput.n359 gnd 0.430304f
C2209 CSoutput.n360 gnd 0.197656f
C2210 CSoutput.t138 gnd 0.048697f
C2211 CSoutput.t118 gnd 0.048697f
C2212 CSoutput.n361 gnd 0.430304f
C2213 CSoutput.n362 gnd 0.300084f
C2214 CSoutput.n363 gnd 0.557579f
C2215 CSoutput.n364 gnd 13.7679f
C2216 CSoutput.t171 gnd 0.048697f
C2217 CSoutput.t0 gnd 0.048697f
C2218 CSoutput.n365 gnd 0.431745f
C2219 CSoutput.t108 gnd 0.048697f
C2220 CSoutput.t164 gnd 0.048697f
C2221 CSoutput.n366 gnd 0.430304f
C2222 CSoutput.n367 gnd 0.400963f
C2223 CSoutput.t139 gnd 0.048697f
C2224 CSoutput.t144 gnd 0.048697f
C2225 CSoutput.n368 gnd 0.430304f
C2226 CSoutput.n369 gnd 0.197656f
C2227 CSoutput.t130 gnd 0.048697f
C2228 CSoutput.t159 gnd 0.048697f
C2229 CSoutput.n370 gnd 0.430304f
C2230 CSoutput.n371 gnd 0.197656f
C2231 CSoutput.t165 gnd 0.048697f
C2232 CSoutput.t172 gnd 0.048697f
C2233 CSoutput.n372 gnd 0.430304f
C2234 CSoutput.n373 gnd 0.197656f
C2235 CSoutput.t127 gnd 0.048697f
C2236 CSoutput.t104 gnd 0.048697f
C2237 CSoutput.n374 gnd 0.430304f
C2238 CSoutput.n375 gnd 0.197656f
C2239 CSoutput.t169 gnd 0.048697f
C2240 CSoutput.t174 gnd 0.048697f
C2241 CSoutput.n376 gnd 0.430304f
C2242 CSoutput.n377 gnd 0.197656f
C2243 CSoutput.t113 gnd 0.048697f
C2244 CSoutput.t132 gnd 0.048697f
C2245 CSoutput.n378 gnd 0.430304f
C2246 CSoutput.n379 gnd 0.197656f
C2247 CSoutput.t126 gnd 0.048697f
C2248 CSoutput.t142 gnd 0.048697f
C2249 CSoutput.n380 gnd 0.430304f
C2250 CSoutput.n381 gnd 0.197656f
C2251 CSoutput.t161 gnd 0.048697f
C2252 CSoutput.t101 gnd 0.048697f
C2253 CSoutput.n382 gnd 0.430304f
C2254 CSoutput.n383 gnd 0.364518f
C2255 CSoutput.t128 gnd 0.048697f
C2256 CSoutput.t148 gnd 0.048697f
C2257 CSoutput.n384 gnd 0.431745f
C2258 CSoutput.t151 gnd 0.048697f
C2259 CSoutput.t170 gnd 0.048697f
C2260 CSoutput.n385 gnd 0.430304f
C2261 CSoutput.n386 gnd 0.400963f
C2262 CSoutput.t143 gnd 0.048697f
C2263 CSoutput.t100 gnd 0.048697f
C2264 CSoutput.n387 gnd 0.430304f
C2265 CSoutput.n388 gnd 0.197656f
C2266 CSoutput.t155 gnd 0.048697f
C2267 CSoutput.t140 gnd 0.048697f
C2268 CSoutput.n389 gnd 0.430304f
C2269 CSoutput.n390 gnd 0.197656f
C2270 CSoutput.t167 gnd 0.048697f
C2271 CSoutput.t163 gnd 0.048697f
C2272 CSoutput.n391 gnd 0.430304f
C2273 CSoutput.n392 gnd 0.197656f
C2274 CSoutput.t175 gnd 0.048697f
C2275 CSoutput.t124 gnd 0.048697f
C2276 CSoutput.n393 gnd 0.430304f
C2277 CSoutput.n394 gnd 0.197656f
C2278 CSoutput.t141 gnd 0.048697f
C2279 CSoutput.t109 gnd 0.048697f
C2280 CSoutput.n395 gnd 0.430304f
C2281 CSoutput.n396 gnd 0.197656f
C2282 CSoutput.t154 gnd 0.048697f
C2283 CSoutput.t136 gnd 0.048697f
C2284 CSoutput.n397 gnd 0.430304f
C2285 CSoutput.n398 gnd 0.197656f
C2286 CSoutput.t122 gnd 0.048697f
C2287 CSoutput.t112 gnd 0.048697f
C2288 CSoutput.n399 gnd 0.430304f
C2289 CSoutput.n400 gnd 0.197656f
C2290 CSoutput.t131 gnd 0.048697f
C2291 CSoutput.t135 gnd 0.048697f
C2292 CSoutput.n401 gnd 0.430304f
C2293 CSoutput.n402 gnd 0.300084f
C2294 CSoutput.n403 gnd 0.557579f
C2295 CSoutput.n404 gnd 8.42525f
C2296 CSoutput.n405 gnd 14.470299f
C2297 vdd.t256 gnd 0.03582f
C2298 vdd.t10 gnd 0.03582f
C2299 vdd.n0 gnd 0.28252f
C2300 vdd.t247 gnd 0.03582f
C2301 vdd.t236 gnd 0.03582f
C2302 vdd.n1 gnd 0.282053f
C2303 vdd.n2 gnd 0.260107f
C2304 vdd.t265 gnd 0.03582f
C2305 vdd.t241 gnd 0.03582f
C2306 vdd.n3 gnd 0.282053f
C2307 vdd.n4 gnd 0.131546f
C2308 vdd.t243 gnd 0.03582f
C2309 vdd.t234 gnd 0.03582f
C2310 vdd.n5 gnd 0.282053f
C2311 vdd.n6 gnd 0.123431f
C2312 vdd.t140 gnd 0.03582f
C2313 vdd.t267 gnd 0.03582f
C2314 vdd.n7 gnd 0.28252f
C2315 vdd.t7 gnd 0.03582f
C2316 vdd.t245 gnd 0.03582f
C2317 vdd.n8 gnd 0.282053f
C2318 vdd.n9 gnd 0.260107f
C2319 vdd.t239 gnd 0.03582f
C2320 vdd.t222 gnd 0.03582f
C2321 vdd.n10 gnd 0.282053f
C2322 vdd.n11 gnd 0.131546f
C2323 vdd.t251 gnd 0.03582f
C2324 vdd.t231 gnd 0.03582f
C2325 vdd.n12 gnd 0.282053f
C2326 vdd.n13 gnd 0.123431f
C2327 vdd.n14 gnd 0.087264f
C2328 vdd.t225 gnd 0.0199f
C2329 vdd.t142 gnd 0.0199f
C2330 vdd.n15 gnd 0.183172f
C2331 vdd.t2 gnd 0.0199f
C2332 vdd.t227 gnd 0.0199f
C2333 vdd.n16 gnd 0.182636f
C2334 vdd.n17 gnd 0.317844f
C2335 vdd.t1 gnd 0.0199f
C2336 vdd.t143 gnd 0.0199f
C2337 vdd.n18 gnd 0.182636f
C2338 vdd.n19 gnd 0.131496f
C2339 vdd.t4 gnd 0.0199f
C2340 vdd.t228 gnd 0.0199f
C2341 vdd.n20 gnd 0.183172f
C2342 vdd.t226 gnd 0.0199f
C2343 vdd.t271 gnd 0.0199f
C2344 vdd.n21 gnd 0.182636f
C2345 vdd.n22 gnd 0.317844f
C2346 vdd.t229 gnd 0.0199f
C2347 vdd.t3 gnd 0.0199f
C2348 vdd.n23 gnd 0.182636f
C2349 vdd.n24 gnd 0.131496f
C2350 vdd.t224 gnd 0.0199f
C2351 vdd.t270 gnd 0.0199f
C2352 vdd.n25 gnd 0.182636f
C2353 vdd.t5 gnd 0.0199f
C2354 vdd.t0 gnd 0.0199f
C2355 vdd.n26 gnd 0.182636f
C2356 vdd.n27 gnd 21.4496f
C2357 vdd.n28 gnd 8.322969f
C2358 vdd.n29 gnd 0.005428f
C2359 vdd.n30 gnd 0.005037f
C2360 vdd.n31 gnd 0.002786f
C2361 vdd.n32 gnd 0.006397f
C2362 vdd.n33 gnd 0.002706f
C2363 vdd.n34 gnd 0.002866f
C2364 vdd.n35 gnd 0.005037f
C2365 vdd.n36 gnd 0.002706f
C2366 vdd.n37 gnd 0.006397f
C2367 vdd.n38 gnd 0.002866f
C2368 vdd.n39 gnd 0.005037f
C2369 vdd.n40 gnd 0.002706f
C2370 vdd.n41 gnd 0.004798f
C2371 vdd.n42 gnd 0.004812f
C2372 vdd.t118 gnd 0.013743f
C2373 vdd.n43 gnd 0.030579f
C2374 vdd.n44 gnd 0.159139f
C2375 vdd.n45 gnd 0.002706f
C2376 vdd.n46 gnd 0.002866f
C2377 vdd.n47 gnd 0.006397f
C2378 vdd.n48 gnd 0.006397f
C2379 vdd.n49 gnd 0.002866f
C2380 vdd.n50 gnd 0.002706f
C2381 vdd.n51 gnd 0.005037f
C2382 vdd.n52 gnd 0.005037f
C2383 vdd.n53 gnd 0.002706f
C2384 vdd.n54 gnd 0.002866f
C2385 vdd.n55 gnd 0.006397f
C2386 vdd.n56 gnd 0.006397f
C2387 vdd.n57 gnd 0.002866f
C2388 vdd.n58 gnd 0.002706f
C2389 vdd.n59 gnd 0.005037f
C2390 vdd.n60 gnd 0.005037f
C2391 vdd.n61 gnd 0.002706f
C2392 vdd.n62 gnd 0.002866f
C2393 vdd.n63 gnd 0.006397f
C2394 vdd.n64 gnd 0.006397f
C2395 vdd.n65 gnd 0.015124f
C2396 vdd.n66 gnd 0.002786f
C2397 vdd.n67 gnd 0.002706f
C2398 vdd.n68 gnd 0.013018f
C2399 vdd.n69 gnd 0.009088f
C2400 vdd.t22 gnd 0.03184f
C2401 vdd.t65 gnd 0.03184f
C2402 vdd.n70 gnd 0.218827f
C2403 vdd.n71 gnd 0.172074f
C2404 vdd.t34 gnd 0.03184f
C2405 vdd.t85 gnd 0.03184f
C2406 vdd.n72 gnd 0.218827f
C2407 vdd.n73 gnd 0.138863f
C2408 vdd.t58 gnd 0.03184f
C2409 vdd.t124 gnd 0.03184f
C2410 vdd.n74 gnd 0.218827f
C2411 vdd.n75 gnd 0.138863f
C2412 vdd.t39 gnd 0.03184f
C2413 vdd.t105 gnd 0.03184f
C2414 vdd.n76 gnd 0.218827f
C2415 vdd.n77 gnd 0.138863f
C2416 vdd.t44 gnd 0.03184f
C2417 vdd.t120 gnd 0.03184f
C2418 vdd.n78 gnd 0.218827f
C2419 vdd.n79 gnd 0.138863f
C2420 vdd.t73 gnd 0.03184f
C2421 vdd.t128 gnd 0.03184f
C2422 vdd.n80 gnd 0.218827f
C2423 vdd.n81 gnd 0.138863f
C2424 vdd.t88 gnd 0.03184f
C2425 vdd.t111 gnd 0.03184f
C2426 vdd.n82 gnd 0.218827f
C2427 vdd.n83 gnd 0.138863f
C2428 vdd.n84 gnd 0.005428f
C2429 vdd.n85 gnd 0.005037f
C2430 vdd.n86 gnd 0.002786f
C2431 vdd.n87 gnd 0.006397f
C2432 vdd.n88 gnd 0.002706f
C2433 vdd.n89 gnd 0.002866f
C2434 vdd.n90 gnd 0.005037f
C2435 vdd.n91 gnd 0.002706f
C2436 vdd.n92 gnd 0.006397f
C2437 vdd.n93 gnd 0.002866f
C2438 vdd.n94 gnd 0.005037f
C2439 vdd.n95 gnd 0.002706f
C2440 vdd.n96 gnd 0.004798f
C2441 vdd.n97 gnd 0.004812f
C2442 vdd.t59 gnd 0.013743f
C2443 vdd.n98 gnd 0.030579f
C2444 vdd.n99 gnd 0.159139f
C2445 vdd.n100 gnd 0.002706f
C2446 vdd.n101 gnd 0.002866f
C2447 vdd.n102 gnd 0.006397f
C2448 vdd.n103 gnd 0.006397f
C2449 vdd.n104 gnd 0.002866f
C2450 vdd.n105 gnd 0.002706f
C2451 vdd.n106 gnd 0.005037f
C2452 vdd.n107 gnd 0.005037f
C2453 vdd.n108 gnd 0.002706f
C2454 vdd.n109 gnd 0.002866f
C2455 vdd.n110 gnd 0.006397f
C2456 vdd.n111 gnd 0.006397f
C2457 vdd.n112 gnd 0.002866f
C2458 vdd.n113 gnd 0.002706f
C2459 vdd.n114 gnd 0.005037f
C2460 vdd.n115 gnd 0.005037f
C2461 vdd.n116 gnd 0.002706f
C2462 vdd.n117 gnd 0.002866f
C2463 vdd.n118 gnd 0.006397f
C2464 vdd.n119 gnd 0.006397f
C2465 vdd.n120 gnd 0.015124f
C2466 vdd.n121 gnd 0.002786f
C2467 vdd.n122 gnd 0.002706f
C2468 vdd.n123 gnd 0.013018f
C2469 vdd.n124 gnd 0.008803f
C2470 vdd.n125 gnd 0.103315f
C2471 vdd.n126 gnd 0.005428f
C2472 vdd.n127 gnd 0.005037f
C2473 vdd.n128 gnd 0.002786f
C2474 vdd.n129 gnd 0.006397f
C2475 vdd.n130 gnd 0.002706f
C2476 vdd.n131 gnd 0.002866f
C2477 vdd.n132 gnd 0.005037f
C2478 vdd.n133 gnd 0.002706f
C2479 vdd.n134 gnd 0.006397f
C2480 vdd.n135 gnd 0.002866f
C2481 vdd.n136 gnd 0.005037f
C2482 vdd.n137 gnd 0.002706f
C2483 vdd.n138 gnd 0.004798f
C2484 vdd.n139 gnd 0.004812f
C2485 vdd.t64 gnd 0.013743f
C2486 vdd.n140 gnd 0.030579f
C2487 vdd.n141 gnd 0.159139f
C2488 vdd.n142 gnd 0.002706f
C2489 vdd.n143 gnd 0.002866f
C2490 vdd.n144 gnd 0.006397f
C2491 vdd.n145 gnd 0.006397f
C2492 vdd.n146 gnd 0.002866f
C2493 vdd.n147 gnd 0.002706f
C2494 vdd.n148 gnd 0.005037f
C2495 vdd.n149 gnd 0.005037f
C2496 vdd.n150 gnd 0.002706f
C2497 vdd.n151 gnd 0.002866f
C2498 vdd.n152 gnd 0.006397f
C2499 vdd.n153 gnd 0.006397f
C2500 vdd.n154 gnd 0.002866f
C2501 vdd.n155 gnd 0.002706f
C2502 vdd.n156 gnd 0.005037f
C2503 vdd.n157 gnd 0.005037f
C2504 vdd.n158 gnd 0.002706f
C2505 vdd.n159 gnd 0.002866f
C2506 vdd.n160 gnd 0.006397f
C2507 vdd.n161 gnd 0.006397f
C2508 vdd.n162 gnd 0.015124f
C2509 vdd.n163 gnd 0.002786f
C2510 vdd.n164 gnd 0.002706f
C2511 vdd.n165 gnd 0.013018f
C2512 vdd.n166 gnd 0.009088f
C2513 vdd.t127 gnd 0.03184f
C2514 vdd.t55 gnd 0.03184f
C2515 vdd.n167 gnd 0.218827f
C2516 vdd.n168 gnd 0.172074f
C2517 vdd.t56 gnd 0.03184f
C2518 vdd.t114 gnd 0.03184f
C2519 vdd.n169 gnd 0.218827f
C2520 vdd.n170 gnd 0.138863f
C2521 vdd.t126 gnd 0.03184f
C2522 vdd.t32 gnd 0.03184f
C2523 vdd.n171 gnd 0.218827f
C2524 vdd.n172 gnd 0.138863f
C2525 vdd.t113 gnd 0.03184f
C2526 vdd.t123 gnd 0.03184f
C2527 vdd.n173 gnd 0.218827f
C2528 vdd.n174 gnd 0.138863f
C2529 vdd.t28 gnd 0.03184f
C2530 vdd.t83 gnd 0.03184f
C2531 vdd.n175 gnd 0.218827f
C2532 vdd.n176 gnd 0.138863f
C2533 vdd.t110 gnd 0.03184f
C2534 vdd.t132 gnd 0.03184f
C2535 vdd.n177 gnd 0.218827f
C2536 vdd.n178 gnd 0.138863f
C2537 vdd.t62 gnd 0.03184f
C2538 vdd.t109 gnd 0.03184f
C2539 vdd.n179 gnd 0.218827f
C2540 vdd.n180 gnd 0.138863f
C2541 vdd.n181 gnd 0.005428f
C2542 vdd.n182 gnd 0.005037f
C2543 vdd.n183 gnd 0.002786f
C2544 vdd.n184 gnd 0.006397f
C2545 vdd.n185 gnd 0.002706f
C2546 vdd.n186 gnd 0.002866f
C2547 vdd.n187 gnd 0.005037f
C2548 vdd.n188 gnd 0.002706f
C2549 vdd.n189 gnd 0.006397f
C2550 vdd.n190 gnd 0.002866f
C2551 vdd.n191 gnd 0.005037f
C2552 vdd.n192 gnd 0.002706f
C2553 vdd.n193 gnd 0.004798f
C2554 vdd.n194 gnd 0.004812f
C2555 vdd.t137 gnd 0.013743f
C2556 vdd.n195 gnd 0.030579f
C2557 vdd.n196 gnd 0.159139f
C2558 vdd.n197 gnd 0.002706f
C2559 vdd.n198 gnd 0.002866f
C2560 vdd.n199 gnd 0.006397f
C2561 vdd.n200 gnd 0.006397f
C2562 vdd.n201 gnd 0.002866f
C2563 vdd.n202 gnd 0.002706f
C2564 vdd.n203 gnd 0.005037f
C2565 vdd.n204 gnd 0.005037f
C2566 vdd.n205 gnd 0.002706f
C2567 vdd.n206 gnd 0.002866f
C2568 vdd.n207 gnd 0.006397f
C2569 vdd.n208 gnd 0.006397f
C2570 vdd.n209 gnd 0.002866f
C2571 vdd.n210 gnd 0.002706f
C2572 vdd.n211 gnd 0.005037f
C2573 vdd.n212 gnd 0.005037f
C2574 vdd.n213 gnd 0.002706f
C2575 vdd.n214 gnd 0.002866f
C2576 vdd.n215 gnd 0.006397f
C2577 vdd.n216 gnd 0.006397f
C2578 vdd.n217 gnd 0.015124f
C2579 vdd.n218 gnd 0.002786f
C2580 vdd.n219 gnd 0.002706f
C2581 vdd.n220 gnd 0.013018f
C2582 vdd.n221 gnd 0.008803f
C2583 vdd.n222 gnd 0.061462f
C2584 vdd.n223 gnd 0.221463f
C2585 vdd.n224 gnd 0.005428f
C2586 vdd.n225 gnd 0.005037f
C2587 vdd.n226 gnd 0.002786f
C2588 vdd.n227 gnd 0.006397f
C2589 vdd.n228 gnd 0.002706f
C2590 vdd.n229 gnd 0.002866f
C2591 vdd.n230 gnd 0.005037f
C2592 vdd.n231 gnd 0.002706f
C2593 vdd.n232 gnd 0.006397f
C2594 vdd.n233 gnd 0.002866f
C2595 vdd.n234 gnd 0.005037f
C2596 vdd.n235 gnd 0.002706f
C2597 vdd.n236 gnd 0.004798f
C2598 vdd.n237 gnd 0.004812f
C2599 vdd.t80 gnd 0.013743f
C2600 vdd.n238 gnd 0.030579f
C2601 vdd.n239 gnd 0.159139f
C2602 vdd.n240 gnd 0.002706f
C2603 vdd.n241 gnd 0.002866f
C2604 vdd.n242 gnd 0.006397f
C2605 vdd.n243 gnd 0.006397f
C2606 vdd.n244 gnd 0.002866f
C2607 vdd.n245 gnd 0.002706f
C2608 vdd.n246 gnd 0.005037f
C2609 vdd.n247 gnd 0.005037f
C2610 vdd.n248 gnd 0.002706f
C2611 vdd.n249 gnd 0.002866f
C2612 vdd.n250 gnd 0.006397f
C2613 vdd.n251 gnd 0.006397f
C2614 vdd.n252 gnd 0.002866f
C2615 vdd.n253 gnd 0.002706f
C2616 vdd.n254 gnd 0.005037f
C2617 vdd.n255 gnd 0.005037f
C2618 vdd.n256 gnd 0.002706f
C2619 vdd.n257 gnd 0.002866f
C2620 vdd.n258 gnd 0.006397f
C2621 vdd.n259 gnd 0.006397f
C2622 vdd.n260 gnd 0.015124f
C2623 vdd.n261 gnd 0.002786f
C2624 vdd.n262 gnd 0.002706f
C2625 vdd.n263 gnd 0.013018f
C2626 vdd.n264 gnd 0.009088f
C2627 vdd.t135 gnd 0.03184f
C2628 vdd.t76 gnd 0.03184f
C2629 vdd.n265 gnd 0.218827f
C2630 vdd.n266 gnd 0.172074f
C2631 vdd.t77 gnd 0.03184f
C2632 vdd.t133 gnd 0.03184f
C2633 vdd.n267 gnd 0.218827f
C2634 vdd.n268 gnd 0.138863f
C2635 vdd.t134 gnd 0.03184f
C2636 vdd.t52 gnd 0.03184f
C2637 vdd.n269 gnd 0.218827f
C2638 vdd.n270 gnd 0.138863f
C2639 vdd.t121 gnd 0.03184f
C2640 vdd.t131 gnd 0.03184f
C2641 vdd.n271 gnd 0.218827f
C2642 vdd.n272 gnd 0.138863f
C2643 vdd.t45 gnd 0.03184f
C2644 vdd.t98 gnd 0.03184f
C2645 vdd.n273 gnd 0.218827f
C2646 vdd.n274 gnd 0.138863f
C2647 vdd.t122 gnd 0.03184f
C2648 vdd.t18 gnd 0.03184f
C2649 vdd.n275 gnd 0.218827f
C2650 vdd.n276 gnd 0.138863f
C2651 vdd.t79 gnd 0.03184f
C2652 vdd.t119 gnd 0.03184f
C2653 vdd.n277 gnd 0.218827f
C2654 vdd.n278 gnd 0.138863f
C2655 vdd.n279 gnd 0.005428f
C2656 vdd.n280 gnd 0.005037f
C2657 vdd.n281 gnd 0.002786f
C2658 vdd.n282 gnd 0.006397f
C2659 vdd.n283 gnd 0.002706f
C2660 vdd.n284 gnd 0.002866f
C2661 vdd.n285 gnd 0.005037f
C2662 vdd.n286 gnd 0.002706f
C2663 vdd.n287 gnd 0.006397f
C2664 vdd.n288 gnd 0.002866f
C2665 vdd.n289 gnd 0.005037f
C2666 vdd.n290 gnd 0.002706f
C2667 vdd.n291 gnd 0.004798f
C2668 vdd.n292 gnd 0.004812f
C2669 vdd.t30 gnd 0.013743f
C2670 vdd.n293 gnd 0.030579f
C2671 vdd.n294 gnd 0.159139f
C2672 vdd.n295 gnd 0.002706f
C2673 vdd.n296 gnd 0.002866f
C2674 vdd.n297 gnd 0.006397f
C2675 vdd.n298 gnd 0.006397f
C2676 vdd.n299 gnd 0.002866f
C2677 vdd.n300 gnd 0.002706f
C2678 vdd.n301 gnd 0.005037f
C2679 vdd.n302 gnd 0.005037f
C2680 vdd.n303 gnd 0.002706f
C2681 vdd.n304 gnd 0.002866f
C2682 vdd.n305 gnd 0.006397f
C2683 vdd.n306 gnd 0.006397f
C2684 vdd.n307 gnd 0.002866f
C2685 vdd.n308 gnd 0.002706f
C2686 vdd.n309 gnd 0.005037f
C2687 vdd.n310 gnd 0.005037f
C2688 vdd.n311 gnd 0.002706f
C2689 vdd.n312 gnd 0.002866f
C2690 vdd.n313 gnd 0.006397f
C2691 vdd.n314 gnd 0.006397f
C2692 vdd.n315 gnd 0.015124f
C2693 vdd.n316 gnd 0.002786f
C2694 vdd.n317 gnd 0.002706f
C2695 vdd.n318 gnd 0.013018f
C2696 vdd.n319 gnd 0.008803f
C2697 vdd.n320 gnd 0.061462f
C2698 vdd.n321 gnd 0.248009f
C2699 vdd.n322 gnd 0.007601f
C2700 vdd.n323 gnd 0.00989f
C2701 vdd.n324 gnd 0.00796f
C2702 vdd.n325 gnd 0.00796f
C2703 vdd.n326 gnd 0.00989f
C2704 vdd.n327 gnd 0.00989f
C2705 vdd.n328 gnd 0.722639f
C2706 vdd.n329 gnd 0.00989f
C2707 vdd.n330 gnd 0.00989f
C2708 vdd.n331 gnd 0.00989f
C2709 vdd.n332 gnd 0.78328f
C2710 vdd.n333 gnd 0.00989f
C2711 vdd.n334 gnd 0.00989f
C2712 vdd.n335 gnd 0.00989f
C2713 vdd.n336 gnd 0.00989f
C2714 vdd.n337 gnd 0.00796f
C2715 vdd.n338 gnd 0.00989f
C2716 vdd.t82 gnd 0.505342f
C2717 vdd.n339 gnd 0.00989f
C2718 vdd.n340 gnd 0.00989f
C2719 vdd.n341 gnd 0.00989f
C2720 vdd.t17 gnd 0.505342f
C2721 vdd.n342 gnd 0.00989f
C2722 vdd.n343 gnd 0.00989f
C2723 vdd.n344 gnd 0.00989f
C2724 vdd.n345 gnd 0.00989f
C2725 vdd.n346 gnd 0.00989f
C2726 vdd.n347 gnd 0.00796f
C2727 vdd.n348 gnd 0.00989f
C2728 vdd.n349 gnd 0.571036f
C2729 vdd.n350 gnd 0.00989f
C2730 vdd.n351 gnd 0.00989f
C2731 vdd.n352 gnd 0.00989f
C2732 vdd.t108 gnd 0.505342f
C2733 vdd.n353 gnd 0.00989f
C2734 vdd.n354 gnd 0.00989f
C2735 vdd.n355 gnd 0.00989f
C2736 vdd.n356 gnd 0.00989f
C2737 vdd.n357 gnd 0.00989f
C2738 vdd.n358 gnd 0.00796f
C2739 vdd.n359 gnd 0.00989f
C2740 vdd.t29 gnd 0.505342f
C2741 vdd.n360 gnd 0.00989f
C2742 vdd.n361 gnd 0.00989f
C2743 vdd.n362 gnd 0.00989f
C2744 vdd.n363 gnd 0.854028f
C2745 vdd.n364 gnd 0.00989f
C2746 vdd.n365 gnd 0.00989f
C2747 vdd.n366 gnd 0.00989f
C2748 vdd.n367 gnd 0.00989f
C2749 vdd.n368 gnd 0.00989f
C2750 vdd.n369 gnd 0.006607f
C2751 vdd.n370 gnd 0.022521f
C2752 vdd.t160 gnd 0.505342f
C2753 vdd.n371 gnd 0.00989f
C2754 vdd.n372 gnd 0.022521f
C2755 vdd.n404 gnd 0.00989f
C2756 vdd.t176 gnd 0.12167f
C2757 vdd.t175 gnd 0.130031f
C2758 vdd.t174 gnd 0.158899f
C2759 vdd.n405 gnd 0.203686f
C2760 vdd.n406 gnd 0.171929f
C2761 vdd.n407 gnd 0.013055f
C2762 vdd.n408 gnd 0.00989f
C2763 vdd.n409 gnd 0.00796f
C2764 vdd.n410 gnd 0.00989f
C2765 vdd.n411 gnd 0.00796f
C2766 vdd.n412 gnd 0.00989f
C2767 vdd.n413 gnd 0.00796f
C2768 vdd.n414 gnd 0.00989f
C2769 vdd.n415 gnd 0.00796f
C2770 vdd.n416 gnd 0.00989f
C2771 vdd.n417 gnd 0.00796f
C2772 vdd.n418 gnd 0.00989f
C2773 vdd.t162 gnd 0.12167f
C2774 vdd.t161 gnd 0.130031f
C2775 vdd.t159 gnd 0.158899f
C2776 vdd.n419 gnd 0.203686f
C2777 vdd.n420 gnd 0.171929f
C2778 vdd.n421 gnd 0.00796f
C2779 vdd.n422 gnd 0.00989f
C2780 vdd.n423 gnd 0.00796f
C2781 vdd.n424 gnd 0.00989f
C2782 vdd.n425 gnd 0.00796f
C2783 vdd.n426 gnd 0.00989f
C2784 vdd.n427 gnd 0.00796f
C2785 vdd.n428 gnd 0.00989f
C2786 vdd.n429 gnd 0.00796f
C2787 vdd.n430 gnd 0.00989f
C2788 vdd.t183 gnd 0.12167f
C2789 vdd.t182 gnd 0.130031f
C2790 vdd.t181 gnd 0.158899f
C2791 vdd.n431 gnd 0.203686f
C2792 vdd.n432 gnd 0.171929f
C2793 vdd.n433 gnd 0.017035f
C2794 vdd.n434 gnd 0.00989f
C2795 vdd.n435 gnd 0.00796f
C2796 vdd.n436 gnd 0.00989f
C2797 vdd.n437 gnd 0.00796f
C2798 vdd.n438 gnd 0.00989f
C2799 vdd.n439 gnd 0.00796f
C2800 vdd.n440 gnd 0.00989f
C2801 vdd.n441 gnd 0.00796f
C2802 vdd.n442 gnd 0.00989f
C2803 vdd.n443 gnd 0.022521f
C2804 vdd.n444 gnd 0.022675f
C2805 vdd.n445 gnd 0.022675f
C2806 vdd.n446 gnd 0.006607f
C2807 vdd.n447 gnd 0.00796f
C2808 vdd.n448 gnd 0.00989f
C2809 vdd.n449 gnd 0.00989f
C2810 vdd.n450 gnd 0.00796f
C2811 vdd.n451 gnd 0.00989f
C2812 vdd.n452 gnd 0.00989f
C2813 vdd.n453 gnd 0.00989f
C2814 vdd.n454 gnd 0.00989f
C2815 vdd.n455 gnd 0.00989f
C2816 vdd.n456 gnd 0.00796f
C2817 vdd.n457 gnd 0.00796f
C2818 vdd.n458 gnd 0.00989f
C2819 vdd.n459 gnd 0.00989f
C2820 vdd.n460 gnd 0.00796f
C2821 vdd.n461 gnd 0.00989f
C2822 vdd.n462 gnd 0.00989f
C2823 vdd.n463 gnd 0.00989f
C2824 vdd.n464 gnd 0.00989f
C2825 vdd.n465 gnd 0.00989f
C2826 vdd.n466 gnd 0.00796f
C2827 vdd.n467 gnd 0.00796f
C2828 vdd.n468 gnd 0.00989f
C2829 vdd.n469 gnd 0.00989f
C2830 vdd.n470 gnd 0.00796f
C2831 vdd.n471 gnd 0.00989f
C2832 vdd.n472 gnd 0.00989f
C2833 vdd.n473 gnd 0.00989f
C2834 vdd.n474 gnd 0.00989f
C2835 vdd.n475 gnd 0.00989f
C2836 vdd.n476 gnd 0.00796f
C2837 vdd.n477 gnd 0.00796f
C2838 vdd.n478 gnd 0.00989f
C2839 vdd.n479 gnd 0.00989f
C2840 vdd.n480 gnd 0.00796f
C2841 vdd.n481 gnd 0.00989f
C2842 vdd.n482 gnd 0.00989f
C2843 vdd.n483 gnd 0.00989f
C2844 vdd.n484 gnd 0.00989f
C2845 vdd.n485 gnd 0.00989f
C2846 vdd.n486 gnd 0.00796f
C2847 vdd.n487 gnd 0.00796f
C2848 vdd.n488 gnd 0.00989f
C2849 vdd.n489 gnd 0.00989f
C2850 vdd.n490 gnd 0.006647f
C2851 vdd.n491 gnd 0.00989f
C2852 vdd.n492 gnd 0.00989f
C2853 vdd.n493 gnd 0.00989f
C2854 vdd.n494 gnd 0.00989f
C2855 vdd.n495 gnd 0.00989f
C2856 vdd.n496 gnd 0.006647f
C2857 vdd.n497 gnd 0.00796f
C2858 vdd.n498 gnd 0.00989f
C2859 vdd.n499 gnd 0.00989f
C2860 vdd.n500 gnd 0.00796f
C2861 vdd.n501 gnd 0.00989f
C2862 vdd.n502 gnd 0.00989f
C2863 vdd.n503 gnd 0.00989f
C2864 vdd.n504 gnd 0.00989f
C2865 vdd.n505 gnd 0.00989f
C2866 vdd.n506 gnd 0.00796f
C2867 vdd.n507 gnd 0.00796f
C2868 vdd.n508 gnd 0.00989f
C2869 vdd.n509 gnd 0.00989f
C2870 vdd.n510 gnd 0.00796f
C2871 vdd.n511 gnd 0.00989f
C2872 vdd.n512 gnd 0.00989f
C2873 vdd.n513 gnd 0.00989f
C2874 vdd.n514 gnd 0.00989f
C2875 vdd.n515 gnd 0.00989f
C2876 vdd.n516 gnd 0.00796f
C2877 vdd.n517 gnd 0.00796f
C2878 vdd.n518 gnd 0.00989f
C2879 vdd.n519 gnd 0.00989f
C2880 vdd.n520 gnd 0.00796f
C2881 vdd.n521 gnd 0.00989f
C2882 vdd.n522 gnd 0.00989f
C2883 vdd.n523 gnd 0.00989f
C2884 vdd.n524 gnd 0.00989f
C2885 vdd.n525 gnd 0.00989f
C2886 vdd.n526 gnd 0.00796f
C2887 vdd.n527 gnd 0.00796f
C2888 vdd.n528 gnd 0.00989f
C2889 vdd.n529 gnd 0.00989f
C2890 vdd.n530 gnd 0.00796f
C2891 vdd.n531 gnd 0.00989f
C2892 vdd.n532 gnd 0.00989f
C2893 vdd.n533 gnd 0.00989f
C2894 vdd.n534 gnd 0.00989f
C2895 vdd.n535 gnd 0.00989f
C2896 vdd.n536 gnd 0.00796f
C2897 vdd.n537 gnd 0.00796f
C2898 vdd.n538 gnd 0.00989f
C2899 vdd.n539 gnd 0.00989f
C2900 vdd.n540 gnd 0.00796f
C2901 vdd.n541 gnd 0.00989f
C2902 vdd.n542 gnd 0.00989f
C2903 vdd.n543 gnd 0.00989f
C2904 vdd.n544 gnd 0.00989f
C2905 vdd.n545 gnd 0.00989f
C2906 vdd.n546 gnd 0.005413f
C2907 vdd.n547 gnd 0.017035f
C2908 vdd.n548 gnd 0.00989f
C2909 vdd.n549 gnd 0.00989f
C2910 vdd.n550 gnd 0.00788f
C2911 vdd.n551 gnd 0.00989f
C2912 vdd.n552 gnd 0.00989f
C2913 vdd.n553 gnd 0.00989f
C2914 vdd.n554 gnd 0.00989f
C2915 vdd.n555 gnd 0.00989f
C2916 vdd.n556 gnd 0.00796f
C2917 vdd.n557 gnd 0.00796f
C2918 vdd.n558 gnd 0.00989f
C2919 vdd.n559 gnd 0.00989f
C2920 vdd.n560 gnd 0.00796f
C2921 vdd.n561 gnd 0.00989f
C2922 vdd.n562 gnd 0.00989f
C2923 vdd.n563 gnd 0.00989f
C2924 vdd.n564 gnd 0.00989f
C2925 vdd.n565 gnd 0.00989f
C2926 vdd.n566 gnd 0.00796f
C2927 vdd.n567 gnd 0.00796f
C2928 vdd.n568 gnd 0.00989f
C2929 vdd.n569 gnd 0.00989f
C2930 vdd.n570 gnd 0.00796f
C2931 vdd.n571 gnd 0.00989f
C2932 vdd.n572 gnd 0.00989f
C2933 vdd.n573 gnd 0.00989f
C2934 vdd.n574 gnd 0.00989f
C2935 vdd.n575 gnd 0.00989f
C2936 vdd.n576 gnd 0.00796f
C2937 vdd.n577 gnd 0.00796f
C2938 vdd.n578 gnd 0.00989f
C2939 vdd.n579 gnd 0.00989f
C2940 vdd.n580 gnd 0.00796f
C2941 vdd.n581 gnd 0.00989f
C2942 vdd.n582 gnd 0.00989f
C2943 vdd.n583 gnd 0.00989f
C2944 vdd.n584 gnd 0.00989f
C2945 vdd.n585 gnd 0.00989f
C2946 vdd.n586 gnd 0.00796f
C2947 vdd.n587 gnd 0.00796f
C2948 vdd.n588 gnd 0.00989f
C2949 vdd.n589 gnd 0.00989f
C2950 vdd.n590 gnd 0.00796f
C2951 vdd.n591 gnd 0.00989f
C2952 vdd.n592 gnd 0.00989f
C2953 vdd.n593 gnd 0.00989f
C2954 vdd.n594 gnd 0.00989f
C2955 vdd.n595 gnd 0.00989f
C2956 vdd.n596 gnd 0.00796f
C2957 vdd.n597 gnd 0.00989f
C2958 vdd.n598 gnd 0.00796f
C2959 vdd.n599 gnd 0.004179f
C2960 vdd.n600 gnd 0.00989f
C2961 vdd.n601 gnd 0.00989f
C2962 vdd.n602 gnd 0.00796f
C2963 vdd.n603 gnd 0.00989f
C2964 vdd.n604 gnd 0.00796f
C2965 vdd.n605 gnd 0.00989f
C2966 vdd.n606 gnd 0.00796f
C2967 vdd.n607 gnd 0.00989f
C2968 vdd.n608 gnd 0.00796f
C2969 vdd.n609 gnd 0.00989f
C2970 vdd.n610 gnd 0.00796f
C2971 vdd.n611 gnd 0.00989f
C2972 vdd.n612 gnd 0.00989f
C2973 vdd.n613 gnd 0.550823f
C2974 vdd.t38 gnd 0.505342f
C2975 vdd.n614 gnd 0.00989f
C2976 vdd.n615 gnd 0.00796f
C2977 vdd.n616 gnd 0.00989f
C2978 vdd.n617 gnd 0.00796f
C2979 vdd.n618 gnd 0.00989f
C2980 vdd.t57 gnd 0.505342f
C2981 vdd.n619 gnd 0.00989f
C2982 vdd.n620 gnd 0.00796f
C2983 vdd.n621 gnd 0.00989f
C2984 vdd.n622 gnd 0.00796f
C2985 vdd.n623 gnd 0.00989f
C2986 vdd.t84 gnd 0.505342f
C2987 vdd.n624 gnd 0.631677f
C2988 vdd.n625 gnd 0.00989f
C2989 vdd.n626 gnd 0.00796f
C2990 vdd.n627 gnd 0.00989f
C2991 vdd.n628 gnd 0.00796f
C2992 vdd.n629 gnd 0.00989f
C2993 vdd.t33 gnd 0.505342f
C2994 vdd.n630 gnd 0.00989f
C2995 vdd.n631 gnd 0.00796f
C2996 vdd.n632 gnd 0.00989f
C2997 vdd.n633 gnd 0.00796f
C2998 vdd.n634 gnd 0.00989f
C2999 vdd.n635 gnd 0.702425f
C3000 vdd.n636 gnd 0.838868f
C3001 vdd.t54 gnd 0.505342f
C3002 vdd.n637 gnd 0.00989f
C3003 vdd.n638 gnd 0.00796f
C3004 vdd.n639 gnd 0.00989f
C3005 vdd.n640 gnd 0.00796f
C3006 vdd.n641 gnd 0.00989f
C3007 vdd.n642 gnd 0.530609f
C3008 vdd.n643 gnd 0.00989f
C3009 vdd.n644 gnd 0.00796f
C3010 vdd.n645 gnd 0.00989f
C3011 vdd.n646 gnd 0.00796f
C3012 vdd.n647 gnd 0.00989f
C3013 vdd.n648 gnd 1.01068f
C3014 vdd.t63 gnd 0.505342f
C3015 vdd.n649 gnd 0.00989f
C3016 vdd.n650 gnd 0.00796f
C3017 vdd.n651 gnd 0.00989f
C3018 vdd.n652 gnd 0.00796f
C3019 vdd.n653 gnd 0.00989f
C3020 vdd.t145 gnd 0.505342f
C3021 vdd.n654 gnd 0.00989f
C3022 vdd.n655 gnd 0.00796f
C3023 vdd.n656 gnd 0.022675f
C3024 vdd.n657 gnd 0.022675f
C3025 vdd.n658 gnd 10.501f
C3026 vdd.n659 gnd 0.56093f
C3027 vdd.n660 gnd 0.022675f
C3028 vdd.n661 gnd 0.008505f
C3029 vdd.n662 gnd 0.00796f
C3030 vdd.n667 gnd 0.006329f
C3031 vdd.n668 gnd 0.00796f
C3032 vdd.n669 gnd 0.00989f
C3033 vdd.n670 gnd 0.00989f
C3034 vdd.n671 gnd 0.00989f
C3035 vdd.n672 gnd 0.00989f
C3036 vdd.n673 gnd 0.00989f
C3037 vdd.n674 gnd 0.00796f
C3038 vdd.n675 gnd 0.00989f
C3039 vdd.n676 gnd 0.00989f
C3040 vdd.n677 gnd 0.00989f
C3041 vdd.n678 gnd 0.00989f
C3042 vdd.n679 gnd 0.00989f
C3043 vdd.n680 gnd 0.00796f
C3044 vdd.n681 gnd 0.00989f
C3045 vdd.n682 gnd 0.00989f
C3046 vdd.n683 gnd 0.00989f
C3047 vdd.n684 gnd 0.00989f
C3048 vdd.n685 gnd 0.00989f
C3049 vdd.t157 gnd 0.12167f
C3050 vdd.t158 gnd 0.130031f
C3051 vdd.t156 gnd 0.158899f
C3052 vdd.n686 gnd 0.203686f
C3053 vdd.n687 gnd 0.171133f
C3054 vdd.n688 gnd 0.016238f
C3055 vdd.n689 gnd 0.00989f
C3056 vdd.n690 gnd 0.00989f
C3057 vdd.n691 gnd 0.00989f
C3058 vdd.n692 gnd 0.00989f
C3059 vdd.n693 gnd 0.00989f
C3060 vdd.n694 gnd 0.00796f
C3061 vdd.n695 gnd 0.00989f
C3062 vdd.n696 gnd 0.00989f
C3063 vdd.n697 gnd 0.00989f
C3064 vdd.n698 gnd 0.00989f
C3065 vdd.n699 gnd 0.00989f
C3066 vdd.n700 gnd 0.00796f
C3067 vdd.n701 gnd 0.00989f
C3068 vdd.n702 gnd 0.00989f
C3069 vdd.n703 gnd 0.00989f
C3070 vdd.n704 gnd 0.00989f
C3071 vdd.n705 gnd 0.00989f
C3072 vdd.n706 gnd 0.00796f
C3073 vdd.n707 gnd 0.00989f
C3074 vdd.n708 gnd 0.00989f
C3075 vdd.n709 gnd 0.00989f
C3076 vdd.n710 gnd 0.00989f
C3077 vdd.n711 gnd 0.00989f
C3078 vdd.n712 gnd 0.00796f
C3079 vdd.n713 gnd 0.00989f
C3080 vdd.n714 gnd 0.00989f
C3081 vdd.n715 gnd 0.00989f
C3082 vdd.n716 gnd 0.00989f
C3083 vdd.n717 gnd 0.00989f
C3084 vdd.n718 gnd 0.00796f
C3085 vdd.n719 gnd 0.00989f
C3086 vdd.n720 gnd 0.00989f
C3087 vdd.n721 gnd 0.00989f
C3088 vdd.n722 gnd 0.00788f
C3089 vdd.t146 gnd 0.12167f
C3090 vdd.t147 gnd 0.130031f
C3091 vdd.t144 gnd 0.158899f
C3092 vdd.n723 gnd 0.203686f
C3093 vdd.n724 gnd 0.171133f
C3094 vdd.n725 gnd 0.00989f
C3095 vdd.n726 gnd 0.00796f
C3096 vdd.n728 gnd 0.00989f
C3097 vdd.n730 gnd 0.00989f
C3098 vdd.n731 gnd 0.00989f
C3099 vdd.n732 gnd 0.00796f
C3100 vdd.n733 gnd 0.00989f
C3101 vdd.n734 gnd 0.00989f
C3102 vdd.n735 gnd 0.00989f
C3103 vdd.n736 gnd 0.00989f
C3104 vdd.n737 gnd 0.00989f
C3105 vdd.n738 gnd 0.00796f
C3106 vdd.n739 gnd 0.00989f
C3107 vdd.n740 gnd 0.00989f
C3108 vdd.n741 gnd 0.00989f
C3109 vdd.n742 gnd 0.00989f
C3110 vdd.n743 gnd 0.00989f
C3111 vdd.n744 gnd 0.00796f
C3112 vdd.n745 gnd 0.00989f
C3113 vdd.n746 gnd 0.00989f
C3114 vdd.n747 gnd 0.00989f
C3115 vdd.n748 gnd 0.006329f
C3116 vdd.n753 gnd 0.006725f
C3117 vdd.n754 gnd 0.006725f
C3118 vdd.n755 gnd 0.006725f
C3119 vdd.n756 gnd 10.2787f
C3120 vdd.n757 gnd 0.006725f
C3121 vdd.n758 gnd 0.006725f
C3122 vdd.n759 gnd 0.006725f
C3123 vdd.n761 gnd 0.006725f
C3124 vdd.n762 gnd 0.006725f
C3125 vdd.n764 gnd 0.006725f
C3126 vdd.n765 gnd 0.004895f
C3127 vdd.n767 gnd 0.006725f
C3128 vdd.t151 gnd 0.271757f
C3129 vdd.t150 gnd 0.278177f
C3130 vdd.t148 gnd 0.177413f
C3131 vdd.n768 gnd 0.095882f
C3132 vdd.n769 gnd 0.054387f
C3133 vdd.n770 gnd 0.009611f
C3134 vdd.n771 gnd 0.015417f
C3135 vdd.n773 gnd 0.006725f
C3136 vdd.n774 gnd 0.687265f
C3137 vdd.n775 gnd 0.014565f
C3138 vdd.n776 gnd 0.014565f
C3139 vdd.n777 gnd 0.006725f
C3140 vdd.n778 gnd 0.0155f
C3141 vdd.n779 gnd 0.006725f
C3142 vdd.n780 gnd 0.006725f
C3143 vdd.n781 gnd 0.006725f
C3144 vdd.n782 gnd 0.006725f
C3145 vdd.n783 gnd 0.006725f
C3146 vdd.n785 gnd 0.006725f
C3147 vdd.n786 gnd 0.006725f
C3148 vdd.n788 gnd 0.006725f
C3149 vdd.n789 gnd 0.006725f
C3150 vdd.n791 gnd 0.006725f
C3151 vdd.n792 gnd 0.006725f
C3152 vdd.n794 gnd 0.006725f
C3153 vdd.n795 gnd 0.006725f
C3154 vdd.n797 gnd 0.006725f
C3155 vdd.n798 gnd 0.006725f
C3156 vdd.n800 gnd 0.006725f
C3157 vdd.n801 gnd 0.004895f
C3158 vdd.n803 gnd 0.006725f
C3159 vdd.t186 gnd 0.271757f
C3160 vdd.t185 gnd 0.278177f
C3161 vdd.t184 gnd 0.177413f
C3162 vdd.n804 gnd 0.095882f
C3163 vdd.n805 gnd 0.054387f
C3164 vdd.n806 gnd 0.009611f
C3165 vdd.n807 gnd 0.006725f
C3166 vdd.n808 gnd 0.006725f
C3167 vdd.t149 gnd 0.343633f
C3168 vdd.n809 gnd 0.006725f
C3169 vdd.n810 gnd 0.006725f
C3170 vdd.n811 gnd 0.006725f
C3171 vdd.n812 gnd 0.006725f
C3172 vdd.n813 gnd 0.006725f
C3173 vdd.n814 gnd 0.687265f
C3174 vdd.n815 gnd 0.006725f
C3175 vdd.n816 gnd 0.006725f
C3176 vdd.n817 gnd 0.56093f
C3177 vdd.n818 gnd 0.006725f
C3178 vdd.n819 gnd 0.006725f
C3179 vdd.n820 gnd 0.006725f
C3180 vdd.n821 gnd 0.006725f
C3181 vdd.n822 gnd 0.687265f
C3182 vdd.n823 gnd 0.006725f
C3183 vdd.n824 gnd 0.006725f
C3184 vdd.n825 gnd 0.006725f
C3185 vdd.n826 gnd 0.006725f
C3186 vdd.n827 gnd 0.006725f
C3187 vdd.t252 gnd 0.343633f
C3188 vdd.n828 gnd 0.006725f
C3189 vdd.n829 gnd 0.006725f
C3190 vdd.n830 gnd 0.006725f
C3191 vdd.n831 gnd 0.006725f
C3192 vdd.n832 gnd 0.006725f
C3193 vdd.t237 gnd 0.343633f
C3194 vdd.n833 gnd 0.006725f
C3195 vdd.n834 gnd 0.006725f
C3196 vdd.n835 gnd 0.682212f
C3197 vdd.n836 gnd 0.006725f
C3198 vdd.n837 gnd 0.006725f
C3199 vdd.n838 gnd 0.006725f
C3200 vdd.t268 gnd 0.343633f
C3201 vdd.n839 gnd 0.006725f
C3202 vdd.n840 gnd 0.006725f
C3203 vdd.n841 gnd 0.530609f
C3204 vdd.n842 gnd 0.006725f
C3205 vdd.n843 gnd 0.006725f
C3206 vdd.n844 gnd 0.006725f
C3207 vdd.n845 gnd 0.459861f
C3208 vdd.n846 gnd 0.006725f
C3209 vdd.n847 gnd 0.006725f
C3210 vdd.n848 gnd 0.379006f
C3211 vdd.n849 gnd 0.006725f
C3212 vdd.n850 gnd 0.006725f
C3213 vdd.n851 gnd 0.006725f
C3214 vdd.n852 gnd 0.565983f
C3215 vdd.n853 gnd 0.006725f
C3216 vdd.n854 gnd 0.006725f
C3217 vdd.t220 gnd 0.343633f
C3218 vdd.n855 gnd 0.006725f
C3219 vdd.t165 gnd 0.278177f
C3220 vdd.t163 gnd 0.177413f
C3221 vdd.t166 gnd 0.278177f
C3222 vdd.n856 gnd 0.156347f
C3223 vdd.n857 gnd 0.006725f
C3224 vdd.n858 gnd 0.006725f
C3225 vdd.n859 gnd 0.687265f
C3226 vdd.n860 gnd 0.006725f
C3227 vdd.n861 gnd 0.006725f
C3228 vdd.t164 gnd 0.267831f
C3229 vdd.t262 gnd 0.121282f
C3230 vdd.n862 gnd 0.006725f
C3231 vdd.n863 gnd 0.006725f
C3232 vdd.n864 gnd 0.006725f
C3233 vdd.t263 gnd 0.343633f
C3234 vdd.n865 gnd 0.006725f
C3235 vdd.n866 gnd 0.006725f
C3236 vdd.n867 gnd 0.006725f
C3237 vdd.n868 gnd 0.006725f
C3238 vdd.n869 gnd 0.006725f
C3239 vdd.t254 gnd 0.343633f
C3240 vdd.n870 gnd 0.006725f
C3241 vdd.n871 gnd 0.006725f
C3242 vdd.n872 gnd 0.611464f
C3243 vdd.n873 gnd 0.006725f
C3244 vdd.n874 gnd 0.006725f
C3245 vdd.n875 gnd 0.006725f
C3246 vdd.n876 gnd 0.379006f
C3247 vdd.n877 gnd 0.006725f
C3248 vdd.n878 gnd 0.006725f
C3249 vdd.t266 gnd 0.343633f
C3250 vdd.n879 gnd 0.006725f
C3251 vdd.n880 gnd 0.006725f
C3252 vdd.n881 gnd 0.006725f
C3253 vdd.n882 gnd 0.530609f
C3254 vdd.n883 gnd 0.006725f
C3255 vdd.n884 gnd 0.006725f
C3256 vdd.t232 gnd 0.252671f
C3257 vdd.t139 gnd 0.308259f
C3258 vdd.n885 gnd 0.006725f
C3259 vdd.n886 gnd 0.006725f
C3260 vdd.n887 gnd 0.006725f
C3261 vdd.t244 gnd 0.343633f
C3262 vdd.n888 gnd 0.006725f
C3263 vdd.n889 gnd 0.006725f
C3264 vdd.t258 gnd 0.343633f
C3265 vdd.n890 gnd 0.006725f
C3266 vdd.n891 gnd 0.006725f
C3267 vdd.n892 gnd 0.006725f
C3268 vdd.t6 gnd 0.343633f
C3269 vdd.n893 gnd 0.006725f
C3270 vdd.n894 gnd 0.006725f
C3271 vdd.t223 gnd 0.343633f
C3272 vdd.n895 gnd 0.006725f
C3273 vdd.n896 gnd 0.006725f
C3274 vdd.n897 gnd 0.006725f
C3275 vdd.n898 gnd 0.687265f
C3276 vdd.n899 gnd 0.006725f
C3277 vdd.n900 gnd 0.006725f
C3278 vdd.n901 gnd 0.475021f
C3279 vdd.n902 gnd 0.006725f
C3280 vdd.n903 gnd 0.006725f
C3281 vdd.n904 gnd 0.006725f
C3282 vdd.t221 gnd 0.343633f
C3283 vdd.n905 gnd 0.006725f
C3284 vdd.n906 gnd 0.006725f
C3285 vdd.n907 gnd 0.006725f
C3286 vdd.n908 gnd 0.006725f
C3287 vdd.n909 gnd 0.006725f
C3288 vdd.t238 gnd 0.343633f
C3289 vdd.n910 gnd 0.006725f
C3290 vdd.n911 gnd 0.006725f
C3291 vdd.t195 gnd 0.343633f
C3292 vdd.n912 gnd 0.006725f
C3293 vdd.n913 gnd 0.0155f
C3294 vdd.n914 gnd 0.0155f
C3295 vdd.t230 gnd 0.60641f
C3296 vdd.n915 gnd 0.014565f
C3297 vdd.n916 gnd 0.014565f
C3298 vdd.n917 gnd 0.38406f
C3299 vdd.n918 gnd 0.0155f
C3300 vdd.n919 gnd 0.006725f
C3301 vdd.n920 gnd 0.006725f
C3302 vdd.t242 gnd 0.60641f
C3303 vdd.n938 gnd 0.0155f
C3304 vdd.n956 gnd 0.014565f
C3305 vdd.n957 gnd 0.006725f
C3306 vdd.n958 gnd 0.014565f
C3307 vdd.t216 gnd 0.271757f
C3308 vdd.t215 gnd 0.278177f
C3309 vdd.t214 gnd 0.177413f
C3310 vdd.n959 gnd 0.095882f
C3311 vdd.n960 gnd 0.054387f
C3312 vdd.n961 gnd 0.015417f
C3313 vdd.n962 gnd 0.006725f
C3314 vdd.n963 gnd 0.38406f
C3315 vdd.n964 gnd 0.014565f
C3316 vdd.n965 gnd 0.006725f
C3317 vdd.n966 gnd 0.0155f
C3318 vdd.n967 gnd 0.006725f
C3319 vdd.t193 gnd 0.271757f
C3320 vdd.t192 gnd 0.278177f
C3321 vdd.t190 gnd 0.177413f
C3322 vdd.n968 gnd 0.095882f
C3323 vdd.n969 gnd 0.054387f
C3324 vdd.n970 gnd 0.009611f
C3325 vdd.n971 gnd 0.006725f
C3326 vdd.n972 gnd 0.006725f
C3327 vdd.t191 gnd 0.343633f
C3328 vdd.n973 gnd 0.006725f
C3329 vdd.t240 gnd 0.343633f
C3330 vdd.n974 gnd 0.006725f
C3331 vdd.n975 gnd 0.006725f
C3332 vdd.n976 gnd 0.006725f
C3333 vdd.n977 gnd 0.006725f
C3334 vdd.n978 gnd 0.006725f
C3335 vdd.n979 gnd 0.687265f
C3336 vdd.n980 gnd 0.006725f
C3337 vdd.n981 gnd 0.006725f
C3338 vdd.t264 gnd 0.343633f
C3339 vdd.n982 gnd 0.006725f
C3340 vdd.n983 gnd 0.006725f
C3341 vdd.n984 gnd 0.006725f
C3342 vdd.n985 gnd 0.006725f
C3343 vdd.n986 gnd 0.475021f
C3344 vdd.n987 gnd 0.006725f
C3345 vdd.n988 gnd 0.006725f
C3346 vdd.n989 gnd 0.006725f
C3347 vdd.n990 gnd 0.006725f
C3348 vdd.n991 gnd 0.006725f
C3349 vdd.t269 gnd 0.343633f
C3350 vdd.n992 gnd 0.006725f
C3351 vdd.n993 gnd 0.006725f
C3352 vdd.t235 gnd 0.343633f
C3353 vdd.n994 gnd 0.006725f
C3354 vdd.n995 gnd 0.006725f
C3355 vdd.n996 gnd 0.006725f
C3356 vdd.t8 gnd 0.343633f
C3357 vdd.n997 gnd 0.006725f
C3358 vdd.n998 gnd 0.006725f
C3359 vdd.t246 gnd 0.343633f
C3360 vdd.n999 gnd 0.006725f
C3361 vdd.n1000 gnd 0.006725f
C3362 vdd.n1001 gnd 0.006725f
C3363 vdd.t9 gnd 0.308259f
C3364 vdd.n1002 gnd 0.006725f
C3365 vdd.n1003 gnd 0.006725f
C3366 vdd.n1004 gnd 0.530609f
C3367 vdd.n1005 gnd 0.006725f
C3368 vdd.n1006 gnd 0.006725f
C3369 vdd.n1007 gnd 0.006725f
C3370 vdd.t255 gnd 0.343633f
C3371 vdd.n1008 gnd 0.006725f
C3372 vdd.n1009 gnd 0.006725f
C3373 vdd.t257 gnd 0.252671f
C3374 vdd.n1010 gnd 0.379006f
C3375 vdd.n1011 gnd 0.006725f
C3376 vdd.n1012 gnd 0.006725f
C3377 vdd.n1013 gnd 0.006725f
C3378 vdd.n1014 gnd 0.611464f
C3379 vdd.n1015 gnd 0.006725f
C3380 vdd.n1016 gnd 0.006725f
C3381 vdd.t141 gnd 0.343633f
C3382 vdd.n1017 gnd 0.006725f
C3383 vdd.n1018 gnd 0.006725f
C3384 vdd.n1019 gnd 0.006725f
C3385 vdd.n1020 gnd 0.687265f
C3386 vdd.n1021 gnd 0.006725f
C3387 vdd.n1022 gnd 0.006725f
C3388 vdd.t249 gnd 0.343633f
C3389 vdd.n1023 gnd 0.006725f
C3390 vdd.n1024 gnd 0.006725f
C3391 vdd.n1025 gnd 0.006725f
C3392 vdd.t248 gnd 0.121282f
C3393 vdd.n1026 gnd 0.006725f
C3394 vdd.n1027 gnd 0.006725f
C3395 vdd.n1028 gnd 0.006725f
C3396 vdd.t206 gnd 0.278177f
C3397 vdd.t204 gnd 0.177413f
C3398 vdd.t207 gnd 0.278177f
C3399 vdd.n1029 gnd 0.156347f
C3400 vdd.n1030 gnd 0.006725f
C3401 vdd.n1031 gnd 0.006725f
C3402 vdd.t259 gnd 0.343633f
C3403 vdd.n1032 gnd 0.006725f
C3404 vdd.n1033 gnd 0.006725f
C3405 vdd.t205 gnd 0.267831f
C3406 vdd.n1034 gnd 0.565983f
C3407 vdd.n1035 gnd 0.006725f
C3408 vdd.n1036 gnd 0.006725f
C3409 vdd.n1037 gnd 0.006725f
C3410 vdd.n1038 gnd 0.379006f
C3411 vdd.n1039 gnd 0.006725f
C3412 vdd.n1040 gnd 0.006725f
C3413 vdd.n1041 gnd 0.459861f
C3414 vdd.n1042 gnd 0.006725f
C3415 vdd.n1043 gnd 0.006725f
C3416 vdd.n1044 gnd 0.006725f
C3417 vdd.n1045 gnd 0.530609f
C3418 vdd.n1046 gnd 0.006725f
C3419 vdd.n1047 gnd 0.006725f
C3420 vdd.t260 gnd 0.343633f
C3421 vdd.n1048 gnd 0.006725f
C3422 vdd.n1049 gnd 0.006725f
C3423 vdd.n1050 gnd 0.006725f
C3424 vdd.n1051 gnd 0.682212f
C3425 vdd.n1052 gnd 0.006725f
C3426 vdd.n1053 gnd 0.006725f
C3427 vdd.t261 gnd 0.343633f
C3428 vdd.n1054 gnd 0.006725f
C3429 vdd.n1055 gnd 0.006725f
C3430 vdd.n1056 gnd 0.006725f
C3431 vdd.n1057 gnd 0.687265f
C3432 vdd.n1058 gnd 0.006725f
C3433 vdd.n1059 gnd 0.006725f
C3434 vdd.t253 gnd 0.343633f
C3435 vdd.n1060 gnd 0.006725f
C3436 vdd.n1061 gnd 0.006725f
C3437 vdd.n1062 gnd 0.006725f
C3438 vdd.n1063 gnd 0.687265f
C3439 vdd.n1064 gnd 0.006725f
C3440 vdd.n1065 gnd 0.006725f
C3441 vdd.n1066 gnd 0.006725f
C3442 vdd.n1067 gnd 0.006725f
C3443 vdd.n1068 gnd 0.006725f
C3444 vdd.n1069 gnd 0.56093f
C3445 vdd.n1070 gnd 0.006725f
C3446 vdd.n1071 gnd 0.006725f
C3447 vdd.n1072 gnd 0.006725f
C3448 vdd.n1073 gnd 0.006725f
C3449 vdd.n1074 gnd 0.006725f
C3450 vdd.n1075 gnd 0.687265f
C3451 vdd.n1076 gnd 0.006725f
C3452 vdd.n1077 gnd 0.006725f
C3453 vdd.t153 gnd 0.343633f
C3454 vdd.n1078 gnd 0.006725f
C3455 vdd.n1079 gnd 0.0155f
C3456 vdd.n1080 gnd 0.0155f
C3457 vdd.n1081 gnd 10.2787f
C3458 vdd.n1082 gnd 0.014565f
C3459 vdd.n1083 gnd 0.014565f
C3460 vdd.n1084 gnd 0.0155f
C3461 vdd.n1085 gnd 0.006725f
C3462 vdd.n1087 gnd 0.006725f
C3463 vdd.n1088 gnd 0.006725f
C3464 vdd.n1089 gnd 0.006725f
C3465 vdd.n1090 gnd 0.006725f
C3466 vdd.n1091 gnd 0.006725f
C3467 vdd.n1092 gnd 0.006725f
C3468 vdd.n1093 gnd 0.035384f
C3469 vdd.n1094 gnd 0.006725f
C3470 vdd.n1095 gnd 0.006725f
C3471 vdd.n1096 gnd 0.006725f
C3472 vdd.n1097 gnd 0.006725f
C3473 vdd.n1098 gnd 0.006725f
C3474 vdd.n1099 gnd 0.006725f
C3475 vdd.n1100 gnd 0.006725f
C3476 vdd.t218 gnd 0.271757f
C3477 vdd.t219 gnd 0.278177f
C3478 vdd.t217 gnd 0.177413f
C3479 vdd.n1101 gnd 0.095882f
C3480 vdd.n1102 gnd 0.054387f
C3481 vdd.n1103 gnd 0.006725f
C3482 vdd.n1104 gnd 0.006725f
C3483 vdd.n1105 gnd 0.006725f
C3484 vdd.n1106 gnd 0.006725f
C3485 vdd.t154 gnd 0.271757f
C3486 vdd.t155 gnd 0.278177f
C3487 vdd.t152 gnd 0.177413f
C3488 vdd.n1107 gnd 0.095882f
C3489 vdd.n1108 gnd 0.054387f
C3490 vdd.n1109 gnd 0.006725f
C3491 vdd.n1110 gnd 0.006725f
C3492 vdd.n1111 gnd 0.006725f
C3493 vdd.n1112 gnd 0.006725f
C3494 vdd.n1113 gnd 0.006725f
C3495 vdd.n1114 gnd 0.006725f
C3496 vdd.n1115 gnd 0.006329f
C3497 vdd.n1118 gnd 0.022675f
C3498 vdd.n1119 gnd 0.00796f
C3499 vdd.n1120 gnd 0.00989f
C3500 vdd.n1122 gnd 0.00989f
C3501 vdd.n1123 gnd 0.006607f
C3502 vdd.n1124 gnd 0.56093f
C3503 vdd.n1125 gnd 10.501f
C3504 vdd.n1126 gnd 0.00989f
C3505 vdd.n1127 gnd 0.022675f
C3506 vdd.n1128 gnd 0.00796f
C3507 vdd.n1129 gnd 0.00989f
C3508 vdd.n1130 gnd 0.00796f
C3509 vdd.n1131 gnd 0.00989f
C3510 vdd.n1132 gnd 1.01068f
C3511 vdd.n1133 gnd 0.00989f
C3512 vdd.n1134 gnd 0.00796f
C3513 vdd.n1135 gnd 0.00796f
C3514 vdd.n1136 gnd 0.00989f
C3515 vdd.n1137 gnd 0.00796f
C3516 vdd.n1138 gnd 0.00989f
C3517 vdd.t95 gnd 0.505342f
C3518 vdd.n1139 gnd 0.00989f
C3519 vdd.n1140 gnd 0.00796f
C3520 vdd.n1141 gnd 0.00989f
C3521 vdd.n1142 gnd 0.00796f
C3522 vdd.n1143 gnd 0.00989f
C3523 vdd.t25 gnd 0.505342f
C3524 vdd.n1144 gnd 0.00989f
C3525 vdd.n1145 gnd 0.00796f
C3526 vdd.n1146 gnd 0.00989f
C3527 vdd.n1147 gnd 0.00796f
C3528 vdd.n1148 gnd 0.00989f
C3529 vdd.t67 gnd 0.505342f
C3530 vdd.n1149 gnd 0.702425f
C3531 vdd.n1150 gnd 0.00989f
C3532 vdd.n1151 gnd 0.00796f
C3533 vdd.n1152 gnd 0.00989f
C3534 vdd.n1153 gnd 0.00796f
C3535 vdd.n1154 gnd 0.00989f
C3536 vdd.n1155 gnd 0.803494f
C3537 vdd.n1156 gnd 0.00989f
C3538 vdd.n1157 gnd 0.00796f
C3539 vdd.n1158 gnd 0.00989f
C3540 vdd.n1159 gnd 0.00796f
C3541 vdd.n1160 gnd 0.00989f
C3542 vdd.n1161 gnd 0.631677f
C3543 vdd.t50 gnd 0.505342f
C3544 vdd.n1162 gnd 0.00989f
C3545 vdd.n1163 gnd 0.00796f
C3546 vdd.n1164 gnd 0.00989f
C3547 vdd.n1165 gnd 0.00796f
C3548 vdd.n1166 gnd 0.00989f
C3549 vdd.t93 gnd 0.505342f
C3550 vdd.n1167 gnd 0.00989f
C3551 vdd.n1168 gnd 0.00796f
C3552 vdd.n1169 gnd 0.00989f
C3553 vdd.n1170 gnd 0.00796f
C3554 vdd.n1171 gnd 0.00989f
C3555 vdd.t23 gnd 0.505342f
C3556 vdd.n1172 gnd 0.550823f
C3557 vdd.n1173 gnd 0.00989f
C3558 vdd.n1174 gnd 0.00796f
C3559 vdd.n1175 gnd 0.00989f
C3560 vdd.n1176 gnd 0.00796f
C3561 vdd.n1177 gnd 0.00989f
C3562 vdd.t46 gnd 0.505342f
C3563 vdd.n1178 gnd 0.00989f
C3564 vdd.n1179 gnd 0.00796f
C3565 vdd.n1180 gnd 0.00989f
C3566 vdd.n1181 gnd 0.00796f
C3567 vdd.n1182 gnd 0.00989f
C3568 vdd.n1183 gnd 0.78328f
C3569 vdd.n1184 gnd 0.838868f
C3570 vdd.t48 gnd 0.505342f
C3571 vdd.n1185 gnd 0.00989f
C3572 vdd.n1186 gnd 0.00796f
C3573 vdd.n1187 gnd 0.00989f
C3574 vdd.n1188 gnd 0.00796f
C3575 vdd.n1189 gnd 0.00989f
C3576 vdd.n1190 gnd 0.611464f
C3577 vdd.n1191 gnd 0.00989f
C3578 vdd.n1192 gnd 0.00796f
C3579 vdd.n1193 gnd 0.00989f
C3580 vdd.n1194 gnd 0.00796f
C3581 vdd.n1195 gnd 0.00989f
C3582 vdd.t69 gnd 0.505342f
C3583 vdd.t19 gnd 0.505342f
C3584 vdd.n1196 gnd 0.00989f
C3585 vdd.n1197 gnd 0.00796f
C3586 vdd.n1198 gnd 0.00989f
C3587 vdd.n1199 gnd 0.00796f
C3588 vdd.n1200 gnd 0.00989f
C3589 vdd.t89 gnd 0.505342f
C3590 vdd.n1201 gnd 0.00989f
C3591 vdd.n1202 gnd 0.00796f
C3592 vdd.n1203 gnd 0.00989f
C3593 vdd.n1204 gnd 0.00796f
C3594 vdd.n1205 gnd 0.00989f
C3595 vdd.t11 gnd 0.505342f
C3596 vdd.n1206 gnd 0.742853f
C3597 vdd.n1207 gnd 0.00989f
C3598 vdd.n1208 gnd 0.00796f
C3599 vdd.n1209 gnd 0.00989f
C3600 vdd.n1210 gnd 0.00796f
C3601 vdd.n1211 gnd 0.00989f
C3602 vdd.n1212 gnd 1.01068f
C3603 vdd.n1213 gnd 0.00989f
C3604 vdd.n1214 gnd 0.00796f
C3605 vdd.n1215 gnd 0.00989f
C3606 vdd.n1216 gnd 0.00796f
C3607 vdd.n1217 gnd 0.00989f
C3608 vdd.n1218 gnd 0.854028f
C3609 vdd.n1219 gnd 0.00989f
C3610 vdd.n1220 gnd 0.00796f
C3611 vdd.n1221 gnd 0.022521f
C3612 vdd.n1222 gnd 0.006607f
C3613 vdd.n1223 gnd 0.022521f
C3614 vdd.n1224 gnd 1.3341f
C3615 vdd.n1225 gnd 0.022521f
C3616 vdd.n1226 gnd 0.006607f
C3617 vdd.n1227 gnd 0.00989f
C3618 vdd.t179 gnd 0.12167f
C3619 vdd.t180 gnd 0.130031f
C3620 vdd.t177 gnd 0.158899f
C3621 vdd.n1228 gnd 0.203686f
C3622 vdd.n1229 gnd 0.171929f
C3623 vdd.n1230 gnd 0.013055f
C3624 vdd.n1231 gnd 0.00989f
C3625 vdd.n1262 gnd 0.00989f
C3626 vdd.n1263 gnd 0.00989f
C3627 vdd.n1264 gnd 0.022675f
C3628 vdd.n1265 gnd 0.00796f
C3629 vdd.n1266 gnd 0.00989f
C3630 vdd.n1267 gnd 0.00989f
C3631 vdd.n1268 gnd 0.00989f
C3632 vdd.n1269 gnd 0.00989f
C3633 vdd.n1270 gnd 0.00796f
C3634 vdd.n1271 gnd 0.00989f
C3635 vdd.n1272 gnd 0.00989f
C3636 vdd.n1273 gnd 0.00989f
C3637 vdd.n1274 gnd 0.00989f
C3638 vdd.n1275 gnd 0.00989f
C3639 vdd.n1276 gnd 0.00796f
C3640 vdd.n1277 gnd 0.00989f
C3641 vdd.n1278 gnd 0.00989f
C3642 vdd.n1279 gnd 0.00989f
C3643 vdd.n1280 gnd 0.00989f
C3644 vdd.n1281 gnd 0.00989f
C3645 vdd.n1282 gnd 0.00796f
C3646 vdd.n1283 gnd 0.00989f
C3647 vdd.n1284 gnd 0.00989f
C3648 vdd.n1285 gnd 0.00989f
C3649 vdd.n1286 gnd 0.00989f
C3650 vdd.n1287 gnd 0.00989f
C3651 vdd.n1288 gnd 0.006647f
C3652 vdd.n1289 gnd 0.00989f
C3653 vdd.n1290 gnd 0.00989f
C3654 vdd.n1291 gnd 0.00989f
C3655 vdd.n1292 gnd 0.00796f
C3656 vdd.n1293 gnd 0.00989f
C3657 vdd.n1294 gnd 0.00989f
C3658 vdd.n1295 gnd 0.00989f
C3659 vdd.n1296 gnd 0.00989f
C3660 vdd.n1297 gnd 0.00989f
C3661 vdd.n1298 gnd 0.00796f
C3662 vdd.n1299 gnd 0.00989f
C3663 vdd.n1300 gnd 0.00989f
C3664 vdd.n1301 gnd 0.00989f
C3665 vdd.n1302 gnd 0.00989f
C3666 vdd.n1303 gnd 0.00989f
C3667 vdd.n1304 gnd 0.00796f
C3668 vdd.n1305 gnd 0.00989f
C3669 vdd.n1306 gnd 0.00989f
C3670 vdd.n1307 gnd 0.00989f
C3671 vdd.n1308 gnd 0.00989f
C3672 vdd.n1309 gnd 0.00989f
C3673 vdd.n1310 gnd 0.00796f
C3674 vdd.n1311 gnd 0.00989f
C3675 vdd.n1312 gnd 0.00989f
C3676 vdd.n1313 gnd 0.00989f
C3677 vdd.n1314 gnd 0.00989f
C3678 vdd.n1315 gnd 0.00989f
C3679 vdd.n1316 gnd 0.00796f
C3680 vdd.n1317 gnd 0.00989f
C3681 vdd.n1318 gnd 0.00989f
C3682 vdd.n1319 gnd 0.00989f
C3683 vdd.n1320 gnd 0.00989f
C3684 vdd.n1321 gnd 0.00788f
C3685 vdd.n1322 gnd 0.00989f
C3686 vdd.n1323 gnd 0.00989f
C3687 vdd.n1324 gnd 0.00989f
C3688 vdd.n1325 gnd 0.00989f
C3689 vdd.n1326 gnd 0.00989f
C3690 vdd.n1327 gnd 0.00796f
C3691 vdd.n1328 gnd 0.00989f
C3692 vdd.n1329 gnd 0.00989f
C3693 vdd.n1330 gnd 0.00989f
C3694 vdd.n1331 gnd 0.00989f
C3695 vdd.n1332 gnd 0.00989f
C3696 vdd.n1333 gnd 0.00796f
C3697 vdd.n1334 gnd 0.00989f
C3698 vdd.n1335 gnd 0.00989f
C3699 vdd.n1336 gnd 0.00989f
C3700 vdd.n1337 gnd 0.00989f
C3701 vdd.n1338 gnd 0.00989f
C3702 vdd.n1339 gnd 0.00796f
C3703 vdd.n1340 gnd 0.00989f
C3704 vdd.n1341 gnd 0.00989f
C3705 vdd.n1342 gnd 0.00989f
C3706 vdd.n1343 gnd 0.00989f
C3707 vdd.n1344 gnd 0.00989f
C3708 vdd.n1345 gnd 0.00796f
C3709 vdd.n1346 gnd 0.00989f
C3710 vdd.n1347 gnd 0.00989f
C3711 vdd.n1348 gnd 0.00989f
C3712 vdd.n1349 gnd 0.00989f
C3713 vdd.n1350 gnd 0.00989f
C3714 vdd.n1351 gnd 0.004179f
C3715 vdd.n1352 gnd 0.00989f
C3716 vdd.n1353 gnd 0.00796f
C3717 vdd.n1354 gnd 0.00796f
C3718 vdd.n1355 gnd 0.00796f
C3719 vdd.n1356 gnd 0.00989f
C3720 vdd.n1357 gnd 0.00989f
C3721 vdd.n1358 gnd 0.00989f
C3722 vdd.n1359 gnd 0.00796f
C3723 vdd.n1360 gnd 0.00796f
C3724 vdd.n1361 gnd 0.00796f
C3725 vdd.n1362 gnd 0.00989f
C3726 vdd.n1363 gnd 0.00989f
C3727 vdd.n1364 gnd 0.00989f
C3728 vdd.n1365 gnd 0.00796f
C3729 vdd.n1366 gnd 0.00796f
C3730 vdd.n1367 gnd 0.00796f
C3731 vdd.n1368 gnd 0.00989f
C3732 vdd.n1369 gnd 0.00989f
C3733 vdd.n1370 gnd 0.00989f
C3734 vdd.n1371 gnd 0.00796f
C3735 vdd.n1372 gnd 0.00796f
C3736 vdd.n1373 gnd 0.00796f
C3737 vdd.n1374 gnd 0.00989f
C3738 vdd.n1375 gnd 0.00989f
C3739 vdd.n1376 gnd 0.00989f
C3740 vdd.n1377 gnd 0.00796f
C3741 vdd.n1378 gnd 0.00796f
C3742 vdd.n1379 gnd 0.00796f
C3743 vdd.n1380 gnd 0.00989f
C3744 vdd.n1381 gnd 0.00989f
C3745 vdd.n1382 gnd 0.00989f
C3746 vdd.n1383 gnd 0.00989f
C3747 vdd.t202 gnd 0.12167f
C3748 vdd.t203 gnd 0.130031f
C3749 vdd.t201 gnd 0.158899f
C3750 vdd.n1384 gnd 0.203686f
C3751 vdd.n1385 gnd 0.171929f
C3752 vdd.n1386 gnd 0.017035f
C3753 vdd.n1387 gnd 0.005413f
C3754 vdd.n1388 gnd 0.00796f
C3755 vdd.n1389 gnd 0.00989f
C3756 vdd.n1390 gnd 0.00989f
C3757 vdd.n1391 gnd 0.00989f
C3758 vdd.n1392 gnd 0.00796f
C3759 vdd.n1393 gnd 0.00796f
C3760 vdd.n1394 gnd 0.00796f
C3761 vdd.n1395 gnd 0.00989f
C3762 vdd.n1396 gnd 0.00989f
C3763 vdd.n1397 gnd 0.00989f
C3764 vdd.n1398 gnd 0.00796f
C3765 vdd.n1399 gnd 0.00796f
C3766 vdd.n1400 gnd 0.00796f
C3767 vdd.n1401 gnd 0.00989f
C3768 vdd.n1402 gnd 0.00989f
C3769 vdd.n1403 gnd 0.00989f
C3770 vdd.n1404 gnd 0.00796f
C3771 vdd.n1405 gnd 0.00796f
C3772 vdd.n1406 gnd 0.00796f
C3773 vdd.n1407 gnd 0.00989f
C3774 vdd.n1408 gnd 0.00989f
C3775 vdd.n1409 gnd 0.00989f
C3776 vdd.n1410 gnd 0.00796f
C3777 vdd.n1411 gnd 0.00796f
C3778 vdd.n1412 gnd 0.00796f
C3779 vdd.n1413 gnd 0.00989f
C3780 vdd.n1414 gnd 0.00989f
C3781 vdd.n1415 gnd 0.00989f
C3782 vdd.n1416 gnd 0.00796f
C3783 vdd.n1417 gnd 0.006647f
C3784 vdd.n1418 gnd 0.00989f
C3785 vdd.n1419 gnd 0.00989f
C3786 vdd.t212 gnd 0.12167f
C3787 vdd.t213 gnd 0.130031f
C3788 vdd.t211 gnd 0.158899f
C3789 vdd.n1420 gnd 0.203686f
C3790 vdd.n1421 gnd 0.171929f
C3791 vdd.n1422 gnd 0.017035f
C3792 vdd.n1423 gnd 0.00989f
C3793 vdd.n1424 gnd 0.00989f
C3794 vdd.n1425 gnd 0.00989f
C3795 vdd.n1426 gnd 0.00796f
C3796 vdd.n1427 gnd 0.00796f
C3797 vdd.n1428 gnd 0.00796f
C3798 vdd.n1429 gnd 0.00989f
C3799 vdd.n1430 gnd 0.00989f
C3800 vdd.n1431 gnd 0.00989f
C3801 vdd.n1432 gnd 0.00796f
C3802 vdd.n1433 gnd 0.00796f
C3803 vdd.n1434 gnd 0.00796f
C3804 vdd.n1435 gnd 0.00989f
C3805 vdd.n1436 gnd 0.00989f
C3806 vdd.n1437 gnd 0.00989f
C3807 vdd.n1438 gnd 0.00796f
C3808 vdd.n1439 gnd 0.00796f
C3809 vdd.n1440 gnd 0.00796f
C3810 vdd.n1441 gnd 0.00989f
C3811 vdd.n1442 gnd 0.00989f
C3812 vdd.n1443 gnd 0.00989f
C3813 vdd.n1444 gnd 0.00796f
C3814 vdd.n1445 gnd 0.00796f
C3815 vdd.n1446 gnd 0.00796f
C3816 vdd.n1447 gnd 0.00989f
C3817 vdd.n1448 gnd 0.00989f
C3818 vdd.n1449 gnd 0.00989f
C3819 vdd.n1450 gnd 0.00796f
C3820 vdd.n1451 gnd 0.006607f
C3821 vdd.n1452 gnd 0.022675f
C3822 vdd.n1454 gnd 2.23361f
C3823 vdd.n1455 gnd 0.022675f
C3824 vdd.n1456 gnd 0.003781f
C3825 vdd.n1457 gnd 0.022675f
C3826 vdd.n1458 gnd 0.022521f
C3827 vdd.n1459 gnd 0.00989f
C3828 vdd.n1460 gnd 0.00796f
C3829 vdd.n1461 gnd 0.00989f
C3830 vdd.t178 gnd 0.505342f
C3831 vdd.n1462 gnd 0.661998f
C3832 vdd.n1463 gnd 0.00989f
C3833 vdd.n1464 gnd 0.00796f
C3834 vdd.n1465 gnd 0.00989f
C3835 vdd.n1466 gnd 0.00989f
C3836 vdd.n1467 gnd 0.00989f
C3837 vdd.n1468 gnd 0.00796f
C3838 vdd.n1469 gnd 0.00989f
C3839 vdd.n1470 gnd 1.01068f
C3840 vdd.n1471 gnd 0.00989f
C3841 vdd.n1472 gnd 0.00796f
C3842 vdd.n1473 gnd 0.00989f
C3843 vdd.n1474 gnd 0.00989f
C3844 vdd.n1475 gnd 0.00989f
C3845 vdd.n1476 gnd 0.00796f
C3846 vdd.n1477 gnd 0.00989f
C3847 vdd.n1478 gnd 0.838868f
C3848 vdd.t13 gnd 0.505342f
C3849 vdd.n1479 gnd 0.581143f
C3850 vdd.n1480 gnd 0.00989f
C3851 vdd.n1481 gnd 0.00796f
C3852 vdd.n1482 gnd 0.00989f
C3853 vdd.n1483 gnd 0.00989f
C3854 vdd.n1484 gnd 0.00989f
C3855 vdd.n1485 gnd 0.00796f
C3856 vdd.n1486 gnd 0.00989f
C3857 vdd.n1487 gnd 0.601357f
C3858 vdd.n1488 gnd 0.00989f
C3859 vdd.n1489 gnd 0.00796f
C3860 vdd.n1490 gnd 0.00989f
C3861 vdd.n1491 gnd 0.00989f
C3862 vdd.n1492 gnd 0.00989f
C3863 vdd.n1493 gnd 0.00796f
C3864 vdd.n1494 gnd 0.00989f
C3865 vdd.n1495 gnd 0.571036f
C3866 vdd.n1496 gnd 0.773173f
C3867 vdd.n1497 gnd 0.00989f
C3868 vdd.n1498 gnd 0.00796f
C3869 vdd.n1499 gnd 0.00989f
C3870 vdd.n1500 gnd 0.00989f
C3871 vdd.n1501 gnd 0.00989f
C3872 vdd.n1502 gnd 0.00796f
C3873 vdd.n1503 gnd 0.00989f
C3874 vdd.n1504 gnd 0.838868f
C3875 vdd.n1505 gnd 0.00989f
C3876 vdd.n1506 gnd 0.00796f
C3877 vdd.n1507 gnd 0.00989f
C3878 vdd.n1508 gnd 0.00989f
C3879 vdd.n1509 gnd 0.00989f
C3880 vdd.n1510 gnd 0.00796f
C3881 vdd.n1511 gnd 0.00989f
C3882 vdd.t15 gnd 0.505342f
C3883 vdd.n1512 gnd 0.732746f
C3884 vdd.n1513 gnd 0.00989f
C3885 vdd.n1514 gnd 0.00796f
C3886 vdd.n1515 gnd 0.00989f
C3887 vdd.n1516 gnd 0.00989f
C3888 vdd.n1517 gnd 0.00989f
C3889 vdd.n1518 gnd 0.00796f
C3890 vdd.n1519 gnd 0.00989f
C3891 vdd.n1520 gnd 0.56093f
C3892 vdd.n1521 gnd 0.00989f
C3893 vdd.n1522 gnd 0.00796f
C3894 vdd.n1523 gnd 0.00989f
C3895 vdd.n1524 gnd 0.00989f
C3896 vdd.n1525 gnd 0.00989f
C3897 vdd.n1526 gnd 0.00796f
C3898 vdd.n1527 gnd 0.00989f
C3899 vdd.n1528 gnd 0.722639f
C3900 vdd.n1529 gnd 0.621571f
C3901 vdd.n1530 gnd 0.00989f
C3902 vdd.n1531 gnd 0.00796f
C3903 vdd.n1532 gnd 0.007601f
C3904 vdd.n1533 gnd 0.005428f
C3905 vdd.n1534 gnd 0.005037f
C3906 vdd.n1535 gnd 0.002786f
C3907 vdd.n1536 gnd 0.006397f
C3908 vdd.n1537 gnd 0.002706f
C3909 vdd.n1538 gnd 0.002866f
C3910 vdd.n1539 gnd 0.005037f
C3911 vdd.n1540 gnd 0.002706f
C3912 vdd.n1541 gnd 0.006397f
C3913 vdd.n1542 gnd 0.002866f
C3914 vdd.n1543 gnd 0.005037f
C3915 vdd.n1544 gnd 0.002706f
C3916 vdd.n1545 gnd 0.004798f
C3917 vdd.n1546 gnd 0.004812f
C3918 vdd.t96 gnd 0.013743f
C3919 vdd.n1547 gnd 0.030579f
C3920 vdd.n1548 gnd 0.159139f
C3921 vdd.n1549 gnd 0.002706f
C3922 vdd.n1550 gnd 0.002866f
C3923 vdd.n1551 gnd 0.006397f
C3924 vdd.n1552 gnd 0.006397f
C3925 vdd.n1553 gnd 0.002866f
C3926 vdd.n1554 gnd 0.002706f
C3927 vdd.n1555 gnd 0.005037f
C3928 vdd.n1556 gnd 0.005037f
C3929 vdd.n1557 gnd 0.002706f
C3930 vdd.n1558 gnd 0.002866f
C3931 vdd.n1559 gnd 0.006397f
C3932 vdd.n1560 gnd 0.006397f
C3933 vdd.n1561 gnd 0.002866f
C3934 vdd.n1562 gnd 0.002706f
C3935 vdd.n1563 gnd 0.005037f
C3936 vdd.n1564 gnd 0.005037f
C3937 vdd.n1565 gnd 0.002706f
C3938 vdd.n1566 gnd 0.002866f
C3939 vdd.n1567 gnd 0.006397f
C3940 vdd.n1568 gnd 0.006397f
C3941 vdd.n1569 gnd 0.015124f
C3942 vdd.n1570 gnd 0.002786f
C3943 vdd.n1571 gnd 0.002706f
C3944 vdd.n1572 gnd 0.013018f
C3945 vdd.n1573 gnd 0.009088f
C3946 vdd.t68 gnd 0.03184f
C3947 vdd.t26 gnd 0.03184f
C3948 vdd.n1574 gnd 0.218827f
C3949 vdd.n1575 gnd 0.172074f
C3950 vdd.t86 gnd 0.03184f
C3951 vdd.t37 gnd 0.03184f
C3952 vdd.n1576 gnd 0.218827f
C3953 vdd.n1577 gnd 0.138863f
C3954 vdd.t125 gnd 0.03184f
C3955 vdd.t136 gnd 0.03184f
C3956 vdd.n1578 gnd 0.218827f
C3957 vdd.n1579 gnd 0.138863f
C3958 vdd.t106 gnd 0.03184f
C3959 vdd.t40 gnd 0.03184f
C3960 vdd.n1580 gnd 0.218827f
C3961 vdd.n1581 gnd 0.138863f
C3962 vdd.t97 gnd 0.03184f
C3963 vdd.t49 gnd 0.03184f
C3964 vdd.n1582 gnd 0.218827f
C3965 vdd.n1583 gnd 0.138863f
C3966 vdd.t129 gnd 0.03184f
C3967 vdd.t74 gnd 0.03184f
C3968 vdd.n1584 gnd 0.218827f
C3969 vdd.n1585 gnd 0.138863f
C3970 vdd.t112 gnd 0.03184f
C3971 vdd.t90 gnd 0.03184f
C3972 vdd.n1586 gnd 0.218827f
C3973 vdd.n1587 gnd 0.138863f
C3974 vdd.n1588 gnd 0.005428f
C3975 vdd.n1589 gnd 0.005037f
C3976 vdd.n1590 gnd 0.002786f
C3977 vdd.n1591 gnd 0.006397f
C3978 vdd.n1592 gnd 0.002706f
C3979 vdd.n1593 gnd 0.002866f
C3980 vdd.n1594 gnd 0.005037f
C3981 vdd.n1595 gnd 0.002706f
C3982 vdd.n1596 gnd 0.006397f
C3983 vdd.n1597 gnd 0.002866f
C3984 vdd.n1598 gnd 0.005037f
C3985 vdd.n1599 gnd 0.002706f
C3986 vdd.n1600 gnd 0.004798f
C3987 vdd.n1601 gnd 0.004812f
C3988 vdd.t14 gnd 0.013743f
C3989 vdd.n1602 gnd 0.030579f
C3990 vdd.n1603 gnd 0.159139f
C3991 vdd.n1604 gnd 0.002706f
C3992 vdd.n1605 gnd 0.002866f
C3993 vdd.n1606 gnd 0.006397f
C3994 vdd.n1607 gnd 0.006397f
C3995 vdd.n1608 gnd 0.002866f
C3996 vdd.n1609 gnd 0.002706f
C3997 vdd.n1610 gnd 0.005037f
C3998 vdd.n1611 gnd 0.005037f
C3999 vdd.n1612 gnd 0.002706f
C4000 vdd.n1613 gnd 0.002866f
C4001 vdd.n1614 gnd 0.006397f
C4002 vdd.n1615 gnd 0.006397f
C4003 vdd.n1616 gnd 0.002866f
C4004 vdd.n1617 gnd 0.002706f
C4005 vdd.n1618 gnd 0.005037f
C4006 vdd.n1619 gnd 0.005037f
C4007 vdd.n1620 gnd 0.002706f
C4008 vdd.n1621 gnd 0.002866f
C4009 vdd.n1622 gnd 0.006397f
C4010 vdd.n1623 gnd 0.006397f
C4011 vdd.n1624 gnd 0.015124f
C4012 vdd.n1625 gnd 0.002786f
C4013 vdd.n1626 gnd 0.002706f
C4014 vdd.n1627 gnd 0.013018f
C4015 vdd.n1628 gnd 0.008803f
C4016 vdd.n1629 gnd 0.103315f
C4017 vdd.n1630 gnd 0.005428f
C4018 vdd.n1631 gnd 0.005037f
C4019 vdd.n1632 gnd 0.002786f
C4020 vdd.n1633 gnd 0.006397f
C4021 vdd.n1634 gnd 0.002706f
C4022 vdd.n1635 gnd 0.002866f
C4023 vdd.n1636 gnd 0.005037f
C4024 vdd.n1637 gnd 0.002706f
C4025 vdd.n1638 gnd 0.006397f
C4026 vdd.n1639 gnd 0.002866f
C4027 vdd.n1640 gnd 0.005037f
C4028 vdd.n1641 gnd 0.002706f
C4029 vdd.n1642 gnd 0.004798f
C4030 vdd.n1643 gnd 0.004812f
C4031 vdd.t130 gnd 0.013743f
C4032 vdd.n1644 gnd 0.030579f
C4033 vdd.n1645 gnd 0.159139f
C4034 vdd.n1646 gnd 0.002706f
C4035 vdd.n1647 gnd 0.002866f
C4036 vdd.n1648 gnd 0.006397f
C4037 vdd.n1649 gnd 0.006397f
C4038 vdd.n1650 gnd 0.002866f
C4039 vdd.n1651 gnd 0.002706f
C4040 vdd.n1652 gnd 0.005037f
C4041 vdd.n1653 gnd 0.005037f
C4042 vdd.n1654 gnd 0.002706f
C4043 vdd.n1655 gnd 0.002866f
C4044 vdd.n1656 gnd 0.006397f
C4045 vdd.n1657 gnd 0.006397f
C4046 vdd.n1658 gnd 0.002866f
C4047 vdd.n1659 gnd 0.002706f
C4048 vdd.n1660 gnd 0.005037f
C4049 vdd.n1661 gnd 0.005037f
C4050 vdd.n1662 gnd 0.002706f
C4051 vdd.n1663 gnd 0.002866f
C4052 vdd.n1664 gnd 0.006397f
C4053 vdd.n1665 gnd 0.006397f
C4054 vdd.n1666 gnd 0.015124f
C4055 vdd.n1667 gnd 0.002786f
C4056 vdd.n1668 gnd 0.002706f
C4057 vdd.n1669 gnd 0.013018f
C4058 vdd.n1670 gnd 0.009088f
C4059 vdd.t102 gnd 0.03184f
C4060 vdd.t53 gnd 0.03184f
C4061 vdd.n1671 gnd 0.218827f
C4062 vdd.n1672 gnd 0.172074f
C4063 vdd.t51 gnd 0.03184f
C4064 vdd.t103 gnd 0.03184f
C4065 vdd.n1673 gnd 0.218827f
C4066 vdd.n1674 gnd 0.138863f
C4067 vdd.t94 gnd 0.03184f
C4068 vdd.t92 gnd 0.03184f
C4069 vdd.n1675 gnd 0.218827f
C4070 vdd.n1676 gnd 0.138863f
C4071 vdd.t47 gnd 0.03184f
C4072 vdd.t24 gnd 0.03184f
C4073 vdd.n1677 gnd 0.218827f
C4074 vdd.n1678 gnd 0.138863f
C4075 vdd.t16 gnd 0.03184f
C4076 vdd.t87 gnd 0.03184f
C4077 vdd.n1679 gnd 0.218827f
C4078 vdd.n1680 gnd 0.138863f
C4079 vdd.t70 gnd 0.03184f
C4080 vdd.t20 gnd 0.03184f
C4081 vdd.n1681 gnd 0.218827f
C4082 vdd.n1682 gnd 0.138863f
C4083 vdd.t12 gnd 0.03184f
C4084 vdd.t107 gnd 0.03184f
C4085 vdd.n1683 gnd 0.218827f
C4086 vdd.n1684 gnd 0.138863f
C4087 vdd.n1685 gnd 0.005428f
C4088 vdd.n1686 gnd 0.005037f
C4089 vdd.n1687 gnd 0.002786f
C4090 vdd.n1688 gnd 0.006397f
C4091 vdd.n1689 gnd 0.002706f
C4092 vdd.n1690 gnd 0.002866f
C4093 vdd.n1691 gnd 0.005037f
C4094 vdd.n1692 gnd 0.002706f
C4095 vdd.n1693 gnd 0.006397f
C4096 vdd.n1694 gnd 0.002866f
C4097 vdd.n1695 gnd 0.005037f
C4098 vdd.n1696 gnd 0.002706f
C4099 vdd.n1697 gnd 0.004798f
C4100 vdd.n1698 gnd 0.004812f
C4101 vdd.t60 gnd 0.013743f
C4102 vdd.n1699 gnd 0.030579f
C4103 vdd.n1700 gnd 0.159139f
C4104 vdd.n1701 gnd 0.002706f
C4105 vdd.n1702 gnd 0.002866f
C4106 vdd.n1703 gnd 0.006397f
C4107 vdd.n1704 gnd 0.006397f
C4108 vdd.n1705 gnd 0.002866f
C4109 vdd.n1706 gnd 0.002706f
C4110 vdd.n1707 gnd 0.005037f
C4111 vdd.n1708 gnd 0.005037f
C4112 vdd.n1709 gnd 0.002706f
C4113 vdd.n1710 gnd 0.002866f
C4114 vdd.n1711 gnd 0.006397f
C4115 vdd.n1712 gnd 0.006397f
C4116 vdd.n1713 gnd 0.002866f
C4117 vdd.n1714 gnd 0.002706f
C4118 vdd.n1715 gnd 0.005037f
C4119 vdd.n1716 gnd 0.005037f
C4120 vdd.n1717 gnd 0.002706f
C4121 vdd.n1718 gnd 0.002866f
C4122 vdd.n1719 gnd 0.006397f
C4123 vdd.n1720 gnd 0.006397f
C4124 vdd.n1721 gnd 0.015124f
C4125 vdd.n1722 gnd 0.002786f
C4126 vdd.n1723 gnd 0.002706f
C4127 vdd.n1724 gnd 0.013018f
C4128 vdd.n1725 gnd 0.008803f
C4129 vdd.n1726 gnd 0.061462f
C4130 vdd.n1727 gnd 0.221463f
C4131 vdd.n1728 gnd 0.005428f
C4132 vdd.n1729 gnd 0.005037f
C4133 vdd.n1730 gnd 0.002786f
C4134 vdd.n1731 gnd 0.006397f
C4135 vdd.n1732 gnd 0.002706f
C4136 vdd.n1733 gnd 0.002866f
C4137 vdd.n1734 gnd 0.005037f
C4138 vdd.n1735 gnd 0.002706f
C4139 vdd.n1736 gnd 0.006397f
C4140 vdd.n1737 gnd 0.002866f
C4141 vdd.n1738 gnd 0.005037f
C4142 vdd.n1739 gnd 0.002706f
C4143 vdd.n1740 gnd 0.004798f
C4144 vdd.n1741 gnd 0.004812f
C4145 vdd.t138 gnd 0.013743f
C4146 vdd.n1742 gnd 0.030579f
C4147 vdd.n1743 gnd 0.159139f
C4148 vdd.n1744 gnd 0.002706f
C4149 vdd.n1745 gnd 0.002866f
C4150 vdd.n1746 gnd 0.006397f
C4151 vdd.n1747 gnd 0.006397f
C4152 vdd.n1748 gnd 0.002866f
C4153 vdd.n1749 gnd 0.002706f
C4154 vdd.n1750 gnd 0.005037f
C4155 vdd.n1751 gnd 0.005037f
C4156 vdd.n1752 gnd 0.002706f
C4157 vdd.n1753 gnd 0.002866f
C4158 vdd.n1754 gnd 0.006397f
C4159 vdd.n1755 gnd 0.006397f
C4160 vdd.n1756 gnd 0.002866f
C4161 vdd.n1757 gnd 0.002706f
C4162 vdd.n1758 gnd 0.005037f
C4163 vdd.n1759 gnd 0.005037f
C4164 vdd.n1760 gnd 0.002706f
C4165 vdd.n1761 gnd 0.002866f
C4166 vdd.n1762 gnd 0.006397f
C4167 vdd.n1763 gnd 0.006397f
C4168 vdd.n1764 gnd 0.015124f
C4169 vdd.n1765 gnd 0.002786f
C4170 vdd.n1766 gnd 0.002706f
C4171 vdd.n1767 gnd 0.013018f
C4172 vdd.n1768 gnd 0.009088f
C4173 vdd.t115 gnd 0.03184f
C4174 vdd.t75 gnd 0.03184f
C4175 vdd.n1769 gnd 0.218827f
C4176 vdd.n1770 gnd 0.172074f
C4177 vdd.t71 gnd 0.03184f
C4178 vdd.t116 gnd 0.03184f
C4179 vdd.n1771 gnd 0.218827f
C4180 vdd.n1772 gnd 0.138863f
C4181 vdd.t101 gnd 0.03184f
C4182 vdd.t100 gnd 0.03184f
C4183 vdd.n1773 gnd 0.218827f
C4184 vdd.n1774 gnd 0.138863f
C4185 vdd.t66 gnd 0.03184f
C4186 vdd.t43 gnd 0.03184f
C4187 vdd.n1775 gnd 0.218827f
C4188 vdd.n1776 gnd 0.138863f
C4189 vdd.t41 gnd 0.03184f
C4190 vdd.t99 gnd 0.03184f
C4191 vdd.n1777 gnd 0.218827f
C4192 vdd.n1778 gnd 0.138863f
C4193 vdd.t81 gnd 0.03184f
C4194 vdd.t42 gnd 0.03184f
C4195 vdd.n1779 gnd 0.218827f
C4196 vdd.n1780 gnd 0.138863f
C4197 vdd.t35 gnd 0.03184f
C4198 vdd.t117 gnd 0.03184f
C4199 vdd.n1781 gnd 0.218827f
C4200 vdd.n1782 gnd 0.138863f
C4201 vdd.n1783 gnd 0.005428f
C4202 vdd.n1784 gnd 0.005037f
C4203 vdd.n1785 gnd 0.002786f
C4204 vdd.n1786 gnd 0.006397f
C4205 vdd.n1787 gnd 0.002706f
C4206 vdd.n1788 gnd 0.002866f
C4207 vdd.n1789 gnd 0.005037f
C4208 vdd.n1790 gnd 0.002706f
C4209 vdd.n1791 gnd 0.006397f
C4210 vdd.n1792 gnd 0.002866f
C4211 vdd.n1793 gnd 0.005037f
C4212 vdd.n1794 gnd 0.002706f
C4213 vdd.n1795 gnd 0.004798f
C4214 vdd.n1796 gnd 0.004812f
C4215 vdd.t78 gnd 0.013743f
C4216 vdd.n1797 gnd 0.030579f
C4217 vdd.n1798 gnd 0.159139f
C4218 vdd.n1799 gnd 0.002706f
C4219 vdd.n1800 gnd 0.002866f
C4220 vdd.n1801 gnd 0.006397f
C4221 vdd.n1802 gnd 0.006397f
C4222 vdd.n1803 gnd 0.002866f
C4223 vdd.n1804 gnd 0.002706f
C4224 vdd.n1805 gnd 0.005037f
C4225 vdd.n1806 gnd 0.005037f
C4226 vdd.n1807 gnd 0.002706f
C4227 vdd.n1808 gnd 0.002866f
C4228 vdd.n1809 gnd 0.006397f
C4229 vdd.n1810 gnd 0.006397f
C4230 vdd.n1811 gnd 0.002866f
C4231 vdd.n1812 gnd 0.002706f
C4232 vdd.n1813 gnd 0.005037f
C4233 vdd.n1814 gnd 0.005037f
C4234 vdd.n1815 gnd 0.002706f
C4235 vdd.n1816 gnd 0.002866f
C4236 vdd.n1817 gnd 0.006397f
C4237 vdd.n1818 gnd 0.006397f
C4238 vdd.n1819 gnd 0.015124f
C4239 vdd.n1820 gnd 0.002786f
C4240 vdd.n1821 gnd 0.002706f
C4241 vdd.n1822 gnd 0.013018f
C4242 vdd.n1823 gnd 0.008803f
C4243 vdd.n1824 gnd 0.061462f
C4244 vdd.n1825 gnd 0.248009f
C4245 vdd.n1826 gnd 2.60479f
C4246 vdd.n1827 gnd 0.583334f
C4247 vdd.n1828 gnd 0.007601f
C4248 vdd.n1829 gnd 0.00989f
C4249 vdd.n1830 gnd 0.00796f
C4250 vdd.n1831 gnd 0.00989f
C4251 vdd.n1832 gnd 0.793387f
C4252 vdd.n1833 gnd 0.00989f
C4253 vdd.n1834 gnd 0.00796f
C4254 vdd.n1835 gnd 0.00989f
C4255 vdd.n1836 gnd 0.00989f
C4256 vdd.n1837 gnd 0.00989f
C4257 vdd.n1838 gnd 0.00796f
C4258 vdd.n1839 gnd 0.00989f
C4259 vdd.t91 gnd 0.505342f
C4260 vdd.n1840 gnd 0.838868f
C4261 vdd.n1841 gnd 0.00989f
C4262 vdd.n1842 gnd 0.00796f
C4263 vdd.n1843 gnd 0.00989f
C4264 vdd.n1844 gnd 0.00989f
C4265 vdd.n1845 gnd 0.00989f
C4266 vdd.n1846 gnd 0.00796f
C4267 vdd.n1847 gnd 0.00989f
C4268 vdd.n1848 gnd 0.712532f
C4269 vdd.n1849 gnd 0.00989f
C4270 vdd.n1850 gnd 0.00796f
C4271 vdd.n1851 gnd 0.00989f
C4272 vdd.n1852 gnd 0.00989f
C4273 vdd.n1853 gnd 0.00989f
C4274 vdd.n1854 gnd 0.00796f
C4275 vdd.n1855 gnd 0.00989f
C4276 vdd.n1856 gnd 0.838868f
C4277 vdd.t36 gnd 0.505342f
C4278 vdd.n1857 gnd 0.540716f
C4279 vdd.n1858 gnd 0.00989f
C4280 vdd.n1859 gnd 0.00796f
C4281 vdd.n1860 gnd 0.00989f
C4282 vdd.n1861 gnd 0.00989f
C4283 vdd.n1862 gnd 0.00989f
C4284 vdd.n1863 gnd 0.00796f
C4285 vdd.n1864 gnd 0.00989f
C4286 vdd.n1865 gnd 0.641784f
C4287 vdd.n1866 gnd 0.00989f
C4288 vdd.n1867 gnd 0.00796f
C4289 vdd.n1868 gnd 0.00989f
C4290 vdd.n1869 gnd 0.00989f
C4291 vdd.n1870 gnd 0.00989f
C4292 vdd.n1871 gnd 0.00796f
C4293 vdd.n1872 gnd 0.00989f
C4294 vdd.n1873 gnd 0.530609f
C4295 vdd.n1874 gnd 0.813601f
C4296 vdd.n1875 gnd 0.00989f
C4297 vdd.n1876 gnd 0.00796f
C4298 vdd.n1877 gnd 0.00989f
C4299 vdd.n1878 gnd 0.00989f
C4300 vdd.n1879 gnd 0.00989f
C4301 vdd.n1880 gnd 0.00796f
C4302 vdd.n1881 gnd 0.00989f
C4303 vdd.n1882 gnd 0.985417f
C4304 vdd.n1883 gnd 0.00989f
C4305 vdd.n1884 gnd 0.00796f
C4306 vdd.n1885 gnd 0.00989f
C4307 vdd.n1886 gnd 0.00989f
C4308 vdd.n1887 gnd 0.022521f
C4309 vdd.n1888 gnd 0.00989f
C4310 vdd.n1889 gnd 0.00989f
C4311 vdd.n1890 gnd 0.00796f
C4312 vdd.n1891 gnd 0.00989f
C4313 vdd.t171 gnd 0.505342f
C4314 vdd.n1892 gnd 0.955096f
C4315 vdd.n1893 gnd 0.00989f
C4316 vdd.n1894 gnd 0.00796f
C4317 vdd.n1895 gnd 0.00989f
C4318 vdd.n1896 gnd 0.00989f
C4319 vdd.n1897 gnd 0.008505f
C4320 vdd.n1898 gnd 0.00796f
C4321 vdd.n1900 gnd 0.00989f
C4322 vdd.n1902 gnd 0.00796f
C4323 vdd.n1903 gnd 0.00989f
C4324 vdd.n1904 gnd 0.00796f
C4325 vdd.n1906 gnd 0.00989f
C4326 vdd.n1907 gnd 0.00796f
C4327 vdd.n1908 gnd 0.00989f
C4328 vdd.n1909 gnd 0.00989f
C4329 vdd.n1910 gnd 0.00989f
C4330 vdd.n1911 gnd 0.00989f
C4331 vdd.n1912 gnd 0.00989f
C4332 vdd.n1913 gnd 0.00796f
C4333 vdd.n1915 gnd 0.00989f
C4334 vdd.n1916 gnd 0.00989f
C4335 vdd.n1917 gnd 0.00989f
C4336 vdd.n1918 gnd 0.00989f
C4337 vdd.n1919 gnd 0.00989f
C4338 vdd.n1920 gnd 0.00796f
C4339 vdd.n1922 gnd 0.00989f
C4340 vdd.n1923 gnd 0.00989f
C4341 vdd.n1924 gnd 0.00989f
C4342 vdd.n1925 gnd 0.00989f
C4343 vdd.n1926 gnd 0.006647f
C4344 vdd.t200 gnd 0.12167f
C4345 vdd.t199 gnd 0.130031f
C4346 vdd.t198 gnd 0.158899f
C4347 vdd.n1927 gnd 0.203686f
C4348 vdd.n1928 gnd 0.171133f
C4349 vdd.n1930 gnd 0.00989f
C4350 vdd.n1931 gnd 0.00989f
C4351 vdd.n1932 gnd 0.00796f
C4352 vdd.n1933 gnd 0.00989f
C4353 vdd.n1935 gnd 0.00989f
C4354 vdd.n1936 gnd 0.00989f
C4355 vdd.n1937 gnd 0.00989f
C4356 vdd.n1938 gnd 0.00989f
C4357 vdd.n1939 gnd 0.00796f
C4358 vdd.n1941 gnd 0.00989f
C4359 vdd.n1942 gnd 0.00989f
C4360 vdd.n1943 gnd 0.00989f
C4361 vdd.n1944 gnd 0.00989f
C4362 vdd.n1945 gnd 0.00989f
C4363 vdd.n1946 gnd 0.00796f
C4364 vdd.n1948 gnd 0.00989f
C4365 vdd.n1949 gnd 0.00989f
C4366 vdd.n1950 gnd 0.00989f
C4367 vdd.n1951 gnd 0.00989f
C4368 vdd.n1952 gnd 0.00989f
C4369 vdd.n1953 gnd 0.00796f
C4370 vdd.n1955 gnd 0.00989f
C4371 vdd.n1956 gnd 0.00989f
C4372 vdd.n1957 gnd 0.00989f
C4373 vdd.n1958 gnd 0.00989f
C4374 vdd.n1959 gnd 0.00989f
C4375 vdd.n1960 gnd 0.00796f
C4376 vdd.n1962 gnd 0.00989f
C4377 vdd.n1963 gnd 0.00989f
C4378 vdd.n1964 gnd 0.00989f
C4379 vdd.n1965 gnd 0.00989f
C4380 vdd.n1966 gnd 0.00788f
C4381 vdd.t189 gnd 0.12167f
C4382 vdd.t188 gnd 0.130031f
C4383 vdd.t187 gnd 0.158899f
C4384 vdd.n1967 gnd 0.203686f
C4385 vdd.n1968 gnd 0.171133f
C4386 vdd.n1970 gnd 0.00989f
C4387 vdd.n1971 gnd 0.00989f
C4388 vdd.n1972 gnd 0.00796f
C4389 vdd.n1973 gnd 0.00989f
C4390 vdd.n1975 gnd 0.00989f
C4391 vdd.n1976 gnd 0.00989f
C4392 vdd.n1977 gnd 0.00989f
C4393 vdd.n1978 gnd 0.00989f
C4394 vdd.n1979 gnd 0.00796f
C4395 vdd.n1981 gnd 0.00989f
C4396 vdd.n1982 gnd 0.00989f
C4397 vdd.n1983 gnd 0.00989f
C4398 vdd.n1984 gnd 0.00989f
C4399 vdd.n1985 gnd 0.00989f
C4400 vdd.n1986 gnd 0.00796f
C4401 vdd.n1988 gnd 0.00989f
C4402 vdd.n1989 gnd 0.00989f
C4403 vdd.n1990 gnd 0.00989f
C4404 vdd.n1991 gnd 0.00989f
C4405 vdd.n1992 gnd 0.00989f
C4406 vdd.n1993 gnd 0.00989f
C4407 vdd.n1994 gnd 0.00796f
C4408 vdd.n1996 gnd 0.00989f
C4409 vdd.n1998 gnd 0.00989f
C4410 vdd.n1999 gnd 0.00796f
C4411 vdd.n2000 gnd 0.00796f
C4412 vdd.n2001 gnd 0.00989f
C4413 vdd.n2003 gnd 0.00989f
C4414 vdd.n2004 gnd 0.00796f
C4415 vdd.n2005 gnd 0.00796f
C4416 vdd.n2006 gnd 0.00989f
C4417 vdd.n2008 gnd 0.00989f
C4418 vdd.n2009 gnd 0.00989f
C4419 vdd.n2010 gnd 0.00796f
C4420 vdd.n2011 gnd 0.00796f
C4421 vdd.n2012 gnd 0.00796f
C4422 vdd.n2013 gnd 0.00989f
C4423 vdd.n2015 gnd 0.00989f
C4424 vdd.n2016 gnd 0.00989f
C4425 vdd.n2017 gnd 0.00796f
C4426 vdd.n2018 gnd 0.00796f
C4427 vdd.n2019 gnd 0.00796f
C4428 vdd.n2020 gnd 0.00989f
C4429 vdd.n2022 gnd 0.00989f
C4430 vdd.n2023 gnd 0.00989f
C4431 vdd.n2024 gnd 0.00796f
C4432 vdd.n2025 gnd 0.00796f
C4433 vdd.n2026 gnd 0.00796f
C4434 vdd.n2027 gnd 0.00989f
C4435 vdd.n2029 gnd 0.00989f
C4436 vdd.n2030 gnd 0.00989f
C4437 vdd.n2031 gnd 0.00796f
C4438 vdd.n2032 gnd 0.00989f
C4439 vdd.n2033 gnd 0.00989f
C4440 vdd.n2034 gnd 0.00989f
C4441 vdd.n2035 gnd 0.016238f
C4442 vdd.n2036 gnd 0.005413f
C4443 vdd.n2037 gnd 0.00796f
C4444 vdd.n2038 gnd 0.00989f
C4445 vdd.n2040 gnd 0.00989f
C4446 vdd.n2041 gnd 0.00989f
C4447 vdd.n2042 gnd 0.00796f
C4448 vdd.n2043 gnd 0.00796f
C4449 vdd.n2044 gnd 0.00796f
C4450 vdd.n2045 gnd 0.00989f
C4451 vdd.n2047 gnd 0.00989f
C4452 vdd.n2048 gnd 0.00989f
C4453 vdd.n2049 gnd 0.00796f
C4454 vdd.n2050 gnd 0.00796f
C4455 vdd.n2051 gnd 0.00796f
C4456 vdd.n2052 gnd 0.00989f
C4457 vdd.n2054 gnd 0.00989f
C4458 vdd.n2055 gnd 0.00989f
C4459 vdd.n2056 gnd 0.00796f
C4460 vdd.n2057 gnd 0.00796f
C4461 vdd.n2058 gnd 0.00796f
C4462 vdd.n2059 gnd 0.00989f
C4463 vdd.n2061 gnd 0.00989f
C4464 vdd.n2062 gnd 0.00989f
C4465 vdd.n2063 gnd 0.00796f
C4466 vdd.n2064 gnd 0.00796f
C4467 vdd.n2065 gnd 0.00796f
C4468 vdd.n2066 gnd 0.00989f
C4469 vdd.n2068 gnd 0.00989f
C4470 vdd.n2069 gnd 0.00989f
C4471 vdd.n2070 gnd 0.00796f
C4472 vdd.n2071 gnd 0.00989f
C4473 vdd.n2072 gnd 0.00989f
C4474 vdd.n2073 gnd 0.00989f
C4475 vdd.n2074 gnd 0.016238f
C4476 vdd.n2075 gnd 0.006647f
C4477 vdd.n2076 gnd 0.00796f
C4478 vdd.n2077 gnd 0.00989f
C4479 vdd.n2079 gnd 0.00989f
C4480 vdd.n2080 gnd 0.00989f
C4481 vdd.n2081 gnd 0.00796f
C4482 vdd.n2082 gnd 0.00796f
C4483 vdd.n2083 gnd 0.00796f
C4484 vdd.n2084 gnd 0.00989f
C4485 vdd.n2086 gnd 0.00989f
C4486 vdd.n2087 gnd 0.00989f
C4487 vdd.n2088 gnd 0.00796f
C4488 vdd.n2089 gnd 0.00796f
C4489 vdd.n2090 gnd 0.00796f
C4490 vdd.n2091 gnd 0.00989f
C4491 vdd.n2093 gnd 0.00989f
C4492 vdd.n2094 gnd 0.00989f
C4493 vdd.n2096 gnd 0.00989f
C4494 vdd.n2097 gnd 0.00796f
C4495 vdd.n2098 gnd 0.006329f
C4496 vdd.n2099 gnd 0.89965f
C4497 vdd.n2101 gnd 0.00796f
C4498 vdd.n2102 gnd 0.00796f
C4499 vdd.n2103 gnd 0.00989f
C4500 vdd.n2105 gnd 0.00989f
C4501 vdd.n2106 gnd 0.00989f
C4502 vdd.n2107 gnd 0.00796f
C4503 vdd.n2108 gnd 0.006607f
C4504 vdd.n2109 gnd 0.022675f
C4505 vdd.n2110 gnd 0.022521f
C4506 vdd.n2111 gnd 0.006607f
C4507 vdd.n2112 gnd 0.022521f
C4508 vdd.n2113 gnd 1.3341f
C4509 vdd.n2114 gnd 0.022521f
C4510 vdd.n2115 gnd 0.022675f
C4511 vdd.n2116 gnd 0.003781f
C4512 vdd.t173 gnd 0.12167f
C4513 vdd.t172 gnd 0.130031f
C4514 vdd.t170 gnd 0.158899f
C4515 vdd.n2117 gnd 0.203686f
C4516 vdd.n2118 gnd 0.171133f
C4517 vdd.n2119 gnd 0.012258f
C4518 vdd.n2120 gnd 0.004179f
C4519 vdd.n2121 gnd 0.008505f
C4520 vdd.n2122 gnd 0.89965f
C4521 vdd.n2123 gnd 0.035384f
C4522 vdd.n2124 gnd 0.006725f
C4523 vdd.n2125 gnd 0.006725f
C4524 vdd.n2126 gnd 0.006725f
C4525 vdd.n2127 gnd 0.006725f
C4526 vdd.n2128 gnd 0.006725f
C4527 vdd.n2129 gnd 0.006725f
C4528 vdd.n2130 gnd 0.006725f
C4529 vdd.n2131 gnd 0.006725f
C4530 vdd.n2133 gnd 0.006725f
C4531 vdd.n2135 gnd 0.006725f
C4532 vdd.n2136 gnd 0.006725f
C4533 vdd.n2137 gnd 0.006725f
C4534 vdd.n2138 gnd 0.006725f
C4535 vdd.n2139 gnd 0.006725f
C4536 vdd.n2141 gnd 0.006725f
C4537 vdd.n2143 gnd 0.006725f
C4538 vdd.n2144 gnd 0.006725f
C4539 vdd.n2145 gnd 0.006725f
C4540 vdd.n2146 gnd 0.006725f
C4541 vdd.n2147 gnd 0.006725f
C4542 vdd.n2149 gnd 0.006725f
C4543 vdd.n2151 gnd 0.006725f
C4544 vdd.n2152 gnd 0.006725f
C4545 vdd.n2153 gnd 0.006725f
C4546 vdd.n2154 gnd 0.006725f
C4547 vdd.n2155 gnd 0.006725f
C4548 vdd.n2157 gnd 0.006725f
C4549 vdd.n2159 gnd 0.006725f
C4550 vdd.n2160 gnd 0.006725f
C4551 vdd.n2161 gnd 0.006725f
C4552 vdd.n2162 gnd 0.006725f
C4553 vdd.n2163 gnd 0.006725f
C4554 vdd.n2165 gnd 0.006725f
C4555 vdd.n2167 gnd 0.006725f
C4556 vdd.n2168 gnd 0.006725f
C4557 vdd.n2169 gnd 0.006725f
C4558 vdd.n2170 gnd 0.006725f
C4559 vdd.n2171 gnd 0.006725f
C4560 vdd.n2173 gnd 0.006725f
C4561 vdd.n2175 gnd 0.006725f
C4562 vdd.n2176 gnd 0.006725f
C4563 vdd.n2177 gnd 0.006725f
C4564 vdd.n2178 gnd 0.006725f
C4565 vdd.n2179 gnd 0.006725f
C4566 vdd.n2181 gnd 0.006725f
C4567 vdd.n2183 gnd 0.006725f
C4568 vdd.n2184 gnd 0.006725f
C4569 vdd.n2185 gnd 0.006725f
C4570 vdd.n2186 gnd 0.006725f
C4571 vdd.n2187 gnd 0.006725f
C4572 vdd.n2189 gnd 0.006725f
C4573 vdd.n2191 gnd 0.006725f
C4574 vdd.n2192 gnd 0.006725f
C4575 vdd.n2193 gnd 0.004895f
C4576 vdd.n2194 gnd 0.009611f
C4577 vdd.n2195 gnd 0.005192f
C4578 vdd.n2196 gnd 0.006725f
C4579 vdd.n2198 gnd 0.006725f
C4580 vdd.n2199 gnd 0.0155f
C4581 vdd.n2200 gnd 0.0155f
C4582 vdd.n2201 gnd 0.014565f
C4583 vdd.n2202 gnd 0.006725f
C4584 vdd.n2203 gnd 0.006725f
C4585 vdd.n2204 gnd 0.006725f
C4586 vdd.n2205 gnd 0.006725f
C4587 vdd.n2206 gnd 0.006725f
C4588 vdd.n2207 gnd 0.006725f
C4589 vdd.n2208 gnd 0.006725f
C4590 vdd.n2209 gnd 0.006725f
C4591 vdd.n2210 gnd 0.006725f
C4592 vdd.n2211 gnd 0.006725f
C4593 vdd.n2212 gnd 0.006725f
C4594 vdd.n2213 gnd 0.006725f
C4595 vdd.n2214 gnd 0.006725f
C4596 vdd.n2215 gnd 0.006725f
C4597 vdd.n2216 gnd 0.006725f
C4598 vdd.n2217 gnd 0.006725f
C4599 vdd.n2218 gnd 0.006725f
C4600 vdd.n2219 gnd 0.006725f
C4601 vdd.n2220 gnd 0.006725f
C4602 vdd.n2221 gnd 0.006725f
C4603 vdd.n2222 gnd 0.006725f
C4604 vdd.n2223 gnd 0.006725f
C4605 vdd.n2224 gnd 0.006725f
C4606 vdd.n2225 gnd 0.006725f
C4607 vdd.n2226 gnd 0.006725f
C4608 vdd.n2227 gnd 0.006725f
C4609 vdd.n2228 gnd 0.006725f
C4610 vdd.n2229 gnd 0.006725f
C4611 vdd.n2230 gnd 0.006725f
C4612 vdd.n2231 gnd 0.006725f
C4613 vdd.n2232 gnd 0.006725f
C4614 vdd.n2233 gnd 0.006725f
C4615 vdd.n2234 gnd 0.006725f
C4616 vdd.n2235 gnd 0.006725f
C4617 vdd.n2236 gnd 0.006725f
C4618 vdd.n2237 gnd 0.006725f
C4619 vdd.n2238 gnd 0.006725f
C4620 vdd.n2239 gnd 0.006725f
C4621 vdd.n2240 gnd 0.006725f
C4622 vdd.n2241 gnd 0.006725f
C4623 vdd.n2242 gnd 0.006725f
C4624 vdd.n2243 gnd 0.006725f
C4625 vdd.n2244 gnd 0.006725f
C4626 vdd.n2245 gnd 0.006725f
C4627 vdd.n2246 gnd 0.006725f
C4628 vdd.n2247 gnd 0.006725f
C4629 vdd.n2248 gnd 0.006725f
C4630 vdd.n2249 gnd 0.006725f
C4631 vdd.n2250 gnd 0.006725f
C4632 vdd.n2251 gnd 0.409327f
C4633 vdd.n2252 gnd 0.006725f
C4634 vdd.n2253 gnd 0.006725f
C4635 vdd.n2254 gnd 0.006725f
C4636 vdd.n2255 gnd 0.006725f
C4637 vdd.n2256 gnd 0.006725f
C4638 vdd.n2257 gnd 0.006725f
C4639 vdd.n2258 gnd 0.006725f
C4640 vdd.n2259 gnd 0.006725f
C4641 vdd.n2260 gnd 0.006725f
C4642 vdd.n2261 gnd 0.006725f
C4643 vdd.n2262 gnd 0.006725f
C4644 vdd.n2263 gnd 0.621571f
C4645 vdd.n2264 gnd 0.006725f
C4646 vdd.n2265 gnd 0.006725f
C4647 vdd.n2266 gnd 0.006725f
C4648 vdd.n2267 gnd 0.006725f
C4649 vdd.n2268 gnd 0.006725f
C4650 vdd.n2269 gnd 0.006725f
C4651 vdd.n2270 gnd 0.006725f
C4652 vdd.n2271 gnd 0.006725f
C4653 vdd.n2272 gnd 0.006725f
C4654 vdd.n2273 gnd 0.006725f
C4655 vdd.n2274 gnd 0.006725f
C4656 vdd.n2275 gnd 0.217297f
C4657 vdd.n2276 gnd 0.006725f
C4658 vdd.n2277 gnd 0.006725f
C4659 vdd.n2278 gnd 0.006725f
C4660 vdd.n2279 gnd 0.006725f
C4661 vdd.n2280 gnd 0.006725f
C4662 vdd.n2281 gnd 0.006725f
C4663 vdd.n2282 gnd 0.006725f
C4664 vdd.n2283 gnd 0.006725f
C4665 vdd.n2284 gnd 0.006725f
C4666 vdd.n2285 gnd 0.006725f
C4667 vdd.n2286 gnd 0.006725f
C4668 vdd.n2287 gnd 0.006725f
C4669 vdd.n2288 gnd 0.006725f
C4670 vdd.n2289 gnd 0.006725f
C4671 vdd.n2290 gnd 0.006725f
C4672 vdd.n2291 gnd 0.006725f
C4673 vdd.n2292 gnd 0.006725f
C4674 vdd.n2293 gnd 0.006725f
C4675 vdd.n2294 gnd 0.006725f
C4676 vdd.n2295 gnd 0.006725f
C4677 vdd.n2296 gnd 0.006725f
C4678 vdd.n2297 gnd 0.006725f
C4679 vdd.n2298 gnd 0.006725f
C4680 vdd.n2299 gnd 0.006725f
C4681 vdd.n2300 gnd 0.006725f
C4682 vdd.n2301 gnd 0.006725f
C4683 vdd.n2302 gnd 0.006725f
C4684 vdd.n2303 gnd 0.006725f
C4685 vdd.n2304 gnd 0.006725f
C4686 vdd.n2305 gnd 0.006725f
C4687 vdd.n2306 gnd 0.006725f
C4688 vdd.n2307 gnd 0.006725f
C4689 vdd.n2308 gnd 0.006725f
C4690 vdd.n2309 gnd 0.006725f
C4691 vdd.n2310 gnd 0.006725f
C4692 vdd.n2311 gnd 0.014565f
C4693 vdd.n2312 gnd 0.0155f
C4694 vdd.n2313 gnd 0.0155f
C4695 vdd.n2315 gnd 0.006725f
C4696 vdd.n2317 gnd 0.006725f
C4697 vdd.n2318 gnd 0.005192f
C4698 vdd.n2319 gnd 0.009611f
C4699 vdd.n2320 gnd 0.004895f
C4700 vdd.n2321 gnd 0.006725f
C4701 vdd.n2322 gnd 0.006725f
C4702 vdd.n2324 gnd 0.006725f
C4703 vdd.n2326 gnd 0.006725f
C4704 vdd.n2327 gnd 0.006725f
C4705 vdd.n2328 gnd 0.006725f
C4706 vdd.n2329 gnd 0.006725f
C4707 vdd.n2330 gnd 0.006725f
C4708 vdd.n2332 gnd 0.006725f
C4709 vdd.n2334 gnd 0.006725f
C4710 vdd.n2335 gnd 0.006725f
C4711 vdd.n2336 gnd 0.006725f
C4712 vdd.n2337 gnd 0.006725f
C4713 vdd.n2338 gnd 0.006725f
C4714 vdd.n2340 gnd 0.006725f
C4715 vdd.n2342 gnd 0.006725f
C4716 vdd.n2343 gnd 0.006725f
C4717 vdd.n2344 gnd 0.006725f
C4718 vdd.n2345 gnd 0.006725f
C4719 vdd.n2346 gnd 0.006725f
C4720 vdd.n2348 gnd 0.006725f
C4721 vdd.n2350 gnd 0.006725f
C4722 vdd.n2351 gnd 0.006725f
C4723 vdd.n2352 gnd 0.006725f
C4724 vdd.n2353 gnd 0.006725f
C4725 vdd.n2354 gnd 0.006725f
C4726 vdd.n2356 gnd 0.006725f
C4727 vdd.n2358 gnd 0.006725f
C4728 vdd.n2359 gnd 0.006725f
C4729 vdd.n2360 gnd 0.006725f
C4730 vdd.n2361 gnd 0.006725f
C4731 vdd.n2362 gnd 0.006725f
C4732 vdd.n2364 gnd 0.006725f
C4733 vdd.n2366 gnd 0.006725f
C4734 vdd.n2367 gnd 0.006725f
C4735 vdd.n2368 gnd 0.006725f
C4736 vdd.n2369 gnd 0.006725f
C4737 vdd.n2370 gnd 0.006725f
C4738 vdd.n2372 gnd 0.006725f
C4739 vdd.n2373 gnd 0.006725f
C4740 vdd.n2374 gnd 0.006725f
C4741 vdd.n2375 gnd 0.006725f
C4742 vdd.n2376 gnd 0.006725f
C4743 vdd.n2377 gnd 0.006725f
C4744 vdd.n2379 gnd 0.006725f
C4745 vdd.n2380 gnd 0.006725f
C4746 vdd.n2381 gnd 0.0155f
C4747 vdd.n2382 gnd 0.014565f
C4748 vdd.n2383 gnd 0.014565f
C4749 vdd.n2384 gnd 0.950043f
C4750 vdd.n2385 gnd 0.014565f
C4751 vdd.n2386 gnd 0.014565f
C4752 vdd.n2387 gnd 0.006725f
C4753 vdd.n2388 gnd 0.006725f
C4754 vdd.n2389 gnd 0.006725f
C4755 vdd.n2390 gnd 0.469968f
C4756 vdd.n2391 gnd 0.006725f
C4757 vdd.n2392 gnd 0.006725f
C4758 vdd.n2393 gnd 0.006725f
C4759 vdd.n2394 gnd 0.006725f
C4760 vdd.n2395 gnd 0.006725f
C4761 vdd.n2396 gnd 0.687265f
C4762 vdd.n2397 gnd 0.006725f
C4763 vdd.n2398 gnd 0.006725f
C4764 vdd.n2399 gnd 0.006725f
C4765 vdd.n2400 gnd 0.006725f
C4766 vdd.n2401 gnd 0.006725f
C4767 vdd.n2402 gnd 0.687265f
C4768 vdd.n2403 gnd 0.006725f
C4769 vdd.n2404 gnd 0.006725f
C4770 vdd.n2405 gnd 0.006725f
C4771 vdd.n2406 gnd 0.006725f
C4772 vdd.n2407 gnd 0.006725f
C4773 vdd.n2408 gnd 0.348686f
C4774 vdd.n2409 gnd 0.006725f
C4775 vdd.n2410 gnd 0.006725f
C4776 vdd.n2411 gnd 0.006725f
C4777 vdd.n2412 gnd 0.006725f
C4778 vdd.n2413 gnd 0.006725f
C4779 vdd.n2414 gnd 0.500289f
C4780 vdd.n2415 gnd 0.006725f
C4781 vdd.n2416 gnd 0.006725f
C4782 vdd.n2417 gnd 0.006725f
C4783 vdd.n2418 gnd 0.006725f
C4784 vdd.n2419 gnd 0.006725f
C4785 vdd.n2420 gnd 0.651891f
C4786 vdd.n2421 gnd 0.006725f
C4787 vdd.n2422 gnd 0.006725f
C4788 vdd.n2423 gnd 0.006725f
C4789 vdd.n2424 gnd 0.006725f
C4790 vdd.n2425 gnd 0.006725f
C4791 vdd.n2426 gnd 0.687265f
C4792 vdd.n2427 gnd 0.006725f
C4793 vdd.n2428 gnd 0.006725f
C4794 vdd.n2429 gnd 0.006725f
C4795 vdd.n2430 gnd 0.006725f
C4796 vdd.n2431 gnd 0.006725f
C4797 vdd.n2432 gnd 0.571036f
C4798 vdd.n2433 gnd 0.006725f
C4799 vdd.n2434 gnd 0.006725f
C4800 vdd.n2435 gnd 0.005538f
C4801 vdd.n2436 gnd 0.019482f
C4802 vdd.n2437 gnd 0.004549f
C4803 vdd.n2438 gnd 0.006725f
C4804 vdd.n2439 gnd 0.419434f
C4805 vdd.n2440 gnd 0.006725f
C4806 vdd.n2441 gnd 0.006725f
C4807 vdd.n2442 gnd 0.006725f
C4808 vdd.n2443 gnd 0.006725f
C4809 vdd.n2444 gnd 0.006725f
C4810 vdd.n2445 gnd 0.419434f
C4811 vdd.n2446 gnd 0.006725f
C4812 vdd.n2447 gnd 0.006725f
C4813 vdd.n2448 gnd 0.006725f
C4814 vdd.n2449 gnd 0.006725f
C4815 vdd.n2450 gnd 0.006725f
C4816 vdd.n2451 gnd 0.571036f
C4817 vdd.n2452 gnd 0.006725f
C4818 vdd.n2453 gnd 0.006725f
C4819 vdd.n2454 gnd 0.006725f
C4820 vdd.n2455 gnd 0.006725f
C4821 vdd.n2456 gnd 0.006725f
C4822 vdd.n2457 gnd 0.586197f
C4823 vdd.n2458 gnd 0.006725f
C4824 vdd.n2459 gnd 0.006725f
C4825 vdd.n2460 gnd 0.006725f
C4826 vdd.n2461 gnd 0.006725f
C4827 vdd.n2462 gnd 0.006725f
C4828 vdd.n2463 gnd 0.434594f
C4829 vdd.n2464 gnd 0.006725f
C4830 vdd.n2465 gnd 0.006725f
C4831 vdd.n2466 gnd 0.006725f
C4832 vdd.n2467 gnd 0.006725f
C4833 vdd.n2468 gnd 0.006725f
C4834 vdd.n2469 gnd 0.217297f
C4835 vdd.n2470 gnd 0.006725f
C4836 vdd.n2471 gnd 0.006725f
C4837 vdd.n2472 gnd 0.006725f
C4838 vdd.n2473 gnd 0.006725f
C4839 vdd.n2474 gnd 0.006725f
C4840 vdd.n2475 gnd 0.217297f
C4841 vdd.n2476 gnd 0.006725f
C4842 vdd.n2477 gnd 0.006725f
C4843 vdd.n2478 gnd 0.006725f
C4844 vdd.n2479 gnd 0.006725f
C4845 vdd.n2480 gnd 0.006725f
C4846 vdd.n2481 gnd 0.687265f
C4847 vdd.n2482 gnd 0.006725f
C4848 vdd.n2483 gnd 0.006725f
C4849 vdd.n2484 gnd 0.006725f
C4850 vdd.n2485 gnd 0.006725f
C4851 vdd.n2486 gnd 0.006725f
C4852 vdd.n2487 gnd 0.006725f
C4853 vdd.n2488 gnd 0.006725f
C4854 vdd.n2489 gnd 0.495235f
C4855 vdd.n2490 gnd 0.006725f
C4856 vdd.n2491 gnd 0.006725f
C4857 vdd.n2492 gnd 0.006725f
C4858 vdd.n2493 gnd 0.006725f
C4859 vdd.n2494 gnd 0.006725f
C4860 vdd.n2495 gnd 0.006725f
C4861 vdd.n2496 gnd 0.429541f
C4862 vdd.n2497 gnd 0.006725f
C4863 vdd.n2498 gnd 0.006725f
C4864 vdd.n2499 gnd 0.006725f
C4865 vdd.n2500 gnd 0.015417f
C4866 vdd.n2501 gnd 0.014648f
C4867 vdd.n2502 gnd 0.006725f
C4868 vdd.n2503 gnd 0.006725f
C4869 vdd.n2504 gnd 0.005192f
C4870 vdd.n2505 gnd 0.006725f
C4871 vdd.n2506 gnd 0.006725f
C4872 vdd.n2507 gnd 0.004895f
C4873 vdd.n2508 gnd 0.006725f
C4874 vdd.n2509 gnd 0.006725f
C4875 vdd.n2510 gnd 0.006725f
C4876 vdd.n2511 gnd 0.006725f
C4877 vdd.n2512 gnd 0.006725f
C4878 vdd.n2513 gnd 0.006725f
C4879 vdd.n2514 gnd 0.006725f
C4880 vdd.n2515 gnd 0.006725f
C4881 vdd.n2516 gnd 0.006725f
C4882 vdd.n2517 gnd 0.006725f
C4883 vdd.n2518 gnd 0.006725f
C4884 vdd.n2519 gnd 0.006725f
C4885 vdd.n2520 gnd 0.006725f
C4886 vdd.n2521 gnd 0.006725f
C4887 vdd.n2522 gnd 0.006725f
C4888 vdd.n2523 gnd 0.006725f
C4889 vdd.n2524 gnd 0.006725f
C4890 vdd.n2525 gnd 0.006725f
C4891 vdd.n2526 gnd 0.006725f
C4892 vdd.n2527 gnd 0.006725f
C4893 vdd.n2528 gnd 0.006725f
C4894 vdd.n2529 gnd 0.006725f
C4895 vdd.n2530 gnd 0.006725f
C4896 vdd.n2531 gnd 0.006725f
C4897 vdd.n2532 gnd 0.006725f
C4898 vdd.n2533 gnd 0.006725f
C4899 vdd.n2534 gnd 0.006725f
C4900 vdd.n2535 gnd 0.006725f
C4901 vdd.n2536 gnd 0.006725f
C4902 vdd.n2537 gnd 0.006725f
C4903 vdd.n2538 gnd 0.006725f
C4904 vdd.n2539 gnd 0.006725f
C4905 vdd.n2540 gnd 0.006725f
C4906 vdd.n2541 gnd 0.006725f
C4907 vdd.n2542 gnd 0.006725f
C4908 vdd.n2543 gnd 0.006725f
C4909 vdd.n2544 gnd 0.006725f
C4910 vdd.n2545 gnd 0.006725f
C4911 vdd.n2546 gnd 0.006725f
C4912 vdd.n2547 gnd 0.006725f
C4913 vdd.n2548 gnd 0.006725f
C4914 vdd.n2549 gnd 0.006725f
C4915 vdd.n2550 gnd 0.006725f
C4916 vdd.n2551 gnd 0.006725f
C4917 vdd.n2552 gnd 0.006725f
C4918 vdd.n2553 gnd 0.006725f
C4919 vdd.n2554 gnd 0.006725f
C4920 vdd.n2555 gnd 0.006725f
C4921 vdd.n2556 gnd 0.006725f
C4922 vdd.n2557 gnd 0.006725f
C4923 vdd.n2558 gnd 0.006725f
C4924 vdd.n2559 gnd 0.006725f
C4925 vdd.n2560 gnd 0.006725f
C4926 vdd.n2561 gnd 0.006725f
C4927 vdd.n2562 gnd 0.006725f
C4928 vdd.n2563 gnd 0.006725f
C4929 vdd.n2564 gnd 0.006725f
C4930 vdd.n2565 gnd 0.006725f
C4931 vdd.n2566 gnd 0.006725f
C4932 vdd.n2567 gnd 0.006725f
C4933 vdd.n2568 gnd 0.0155f
C4934 vdd.n2569 gnd 0.014565f
C4935 vdd.n2570 gnd 0.014565f
C4936 vdd.n2571 gnd 0.79844f
C4937 vdd.n2572 gnd 0.014565f
C4938 vdd.n2573 gnd 0.0155f
C4939 vdd.n2574 gnd 0.014648f
C4940 vdd.n2575 gnd 0.006725f
C4941 vdd.n2576 gnd 0.006725f
C4942 vdd.n2577 gnd 0.006725f
C4943 vdd.n2578 gnd 0.005192f
C4944 vdd.n2579 gnd 0.009611f
C4945 vdd.n2580 gnd 0.004895f
C4946 vdd.n2581 gnd 0.006725f
C4947 vdd.n2582 gnd 0.006725f
C4948 vdd.n2583 gnd 0.006725f
C4949 vdd.n2584 gnd 0.006725f
C4950 vdd.n2585 gnd 0.006725f
C4951 vdd.n2586 gnd 0.006725f
C4952 vdd.n2587 gnd 0.006725f
C4953 vdd.n2588 gnd 0.006725f
C4954 vdd.n2589 gnd 0.006725f
C4955 vdd.n2590 gnd 0.006725f
C4956 vdd.n2591 gnd 0.006725f
C4957 vdd.n2592 gnd 0.006725f
C4958 vdd.n2593 gnd 0.006725f
C4959 vdd.n2594 gnd 0.006725f
C4960 vdd.n2595 gnd 0.006725f
C4961 vdd.n2596 gnd 0.006725f
C4962 vdd.n2597 gnd 0.006725f
C4963 vdd.n2598 gnd 0.006725f
C4964 vdd.n2599 gnd 0.006725f
C4965 vdd.n2600 gnd 0.006725f
C4966 vdd.n2601 gnd 0.006725f
C4967 vdd.n2602 gnd 0.006725f
C4968 vdd.n2603 gnd 0.006725f
C4969 vdd.n2604 gnd 0.006725f
C4970 vdd.n2605 gnd 0.006725f
C4971 vdd.n2606 gnd 0.006725f
C4972 vdd.n2607 gnd 0.006725f
C4973 vdd.n2608 gnd 0.006725f
C4974 vdd.n2609 gnd 0.006725f
C4975 vdd.n2610 gnd 0.006725f
C4976 vdd.n2611 gnd 0.006725f
C4977 vdd.n2612 gnd 0.006725f
C4978 vdd.n2613 gnd 0.006725f
C4979 vdd.n2614 gnd 0.006725f
C4980 vdd.n2615 gnd 0.006725f
C4981 vdd.n2616 gnd 0.006725f
C4982 vdd.n2617 gnd 0.006725f
C4983 vdd.n2618 gnd 0.006725f
C4984 vdd.n2619 gnd 0.006725f
C4985 vdd.n2620 gnd 0.006725f
C4986 vdd.n2621 gnd 0.006725f
C4987 vdd.n2622 gnd 0.006725f
C4988 vdd.n2623 gnd 0.006725f
C4989 vdd.n2624 gnd 0.006725f
C4990 vdd.n2625 gnd 0.006725f
C4991 vdd.n2626 gnd 0.006725f
C4992 vdd.n2627 gnd 0.006725f
C4993 vdd.n2628 gnd 0.006725f
C4994 vdd.n2629 gnd 0.006725f
C4995 vdd.n2630 gnd 0.006725f
C4996 vdd.n2631 gnd 0.006725f
C4997 vdd.n2632 gnd 0.006725f
C4998 vdd.n2633 gnd 0.006725f
C4999 vdd.n2634 gnd 0.006725f
C5000 vdd.n2635 gnd 0.006725f
C5001 vdd.n2636 gnd 0.006725f
C5002 vdd.n2637 gnd 0.006725f
C5003 vdd.n2638 gnd 0.006725f
C5004 vdd.n2639 gnd 0.006725f
C5005 vdd.n2640 gnd 0.006725f
C5006 vdd.n2641 gnd 0.0155f
C5007 vdd.n2642 gnd 0.0155f
C5008 vdd.n2643 gnd 0.838868f
C5009 vdd.t233 gnd 2.98152f
C5010 vdd.t250 gnd 2.98152f
C5011 vdd.n2677 gnd 0.006725f
C5012 vdd.t209 gnd 0.271757f
C5013 vdd.t210 gnd 0.278177f
C5014 vdd.t208 gnd 0.177413f
C5015 vdd.n2678 gnd 0.095882f
C5016 vdd.n2679 gnd 0.054387f
C5017 vdd.n2680 gnd 0.009611f
C5018 vdd.n2681 gnd 0.006725f
C5019 vdd.n2682 gnd 0.006725f
C5020 vdd.n2683 gnd 0.006725f
C5021 vdd.n2684 gnd 0.006725f
C5022 vdd.n2685 gnd 0.006725f
C5023 vdd.n2686 gnd 0.006725f
C5024 vdd.n2687 gnd 0.006725f
C5025 vdd.n2688 gnd 0.006725f
C5026 vdd.n2689 gnd 0.006725f
C5027 vdd.n2690 gnd 0.006725f
C5028 vdd.n2691 gnd 0.006725f
C5029 vdd.n2692 gnd 0.006725f
C5030 vdd.n2693 gnd 0.006725f
C5031 vdd.n2694 gnd 0.006725f
C5032 vdd.n2695 gnd 0.006725f
C5033 vdd.n2696 gnd 0.006725f
C5034 vdd.n2697 gnd 0.006725f
C5035 vdd.n2698 gnd 0.006725f
C5036 vdd.n2699 gnd 0.006725f
C5037 vdd.n2700 gnd 0.006725f
C5038 vdd.n2701 gnd 0.006725f
C5039 vdd.n2702 gnd 0.006725f
C5040 vdd.n2703 gnd 0.006725f
C5041 vdd.n2704 gnd 0.006725f
C5042 vdd.n2705 gnd 0.006725f
C5043 vdd.n2706 gnd 0.006725f
C5044 vdd.n2707 gnd 0.006725f
C5045 vdd.n2708 gnd 0.006725f
C5046 vdd.n2709 gnd 0.006725f
C5047 vdd.n2710 gnd 0.006725f
C5048 vdd.n2711 gnd 0.006725f
C5049 vdd.n2712 gnd 0.006725f
C5050 vdd.n2713 gnd 0.006725f
C5051 vdd.n2714 gnd 0.006725f
C5052 vdd.n2715 gnd 0.006725f
C5053 vdd.n2716 gnd 0.006725f
C5054 vdd.n2717 gnd 0.006725f
C5055 vdd.n2718 gnd 0.006725f
C5056 vdd.n2719 gnd 0.006725f
C5057 vdd.n2720 gnd 0.006725f
C5058 vdd.n2721 gnd 0.006725f
C5059 vdd.n2722 gnd 0.006725f
C5060 vdd.n2723 gnd 0.006725f
C5061 vdd.n2724 gnd 0.006725f
C5062 vdd.n2725 gnd 0.006725f
C5063 vdd.n2726 gnd 0.006725f
C5064 vdd.n2727 gnd 0.006725f
C5065 vdd.n2728 gnd 0.006725f
C5066 vdd.n2729 gnd 0.006725f
C5067 vdd.n2730 gnd 0.006725f
C5068 vdd.n2731 gnd 0.006725f
C5069 vdd.n2732 gnd 0.006725f
C5070 vdd.n2733 gnd 0.006725f
C5071 vdd.n2734 gnd 0.006725f
C5072 vdd.n2735 gnd 0.006725f
C5073 vdd.n2736 gnd 0.006725f
C5074 vdd.n2737 gnd 0.006725f
C5075 vdd.n2738 gnd 0.006725f
C5076 vdd.n2739 gnd 0.006725f
C5077 vdd.n2740 gnd 0.006725f
C5078 vdd.n2741 gnd 0.004895f
C5079 vdd.n2742 gnd 0.006725f
C5080 vdd.n2743 gnd 0.006725f
C5081 vdd.n2744 gnd 0.005192f
C5082 vdd.n2745 gnd 0.006725f
C5083 vdd.n2746 gnd 0.006725f
C5084 vdd.t196 gnd 0.271757f
C5085 vdd.t197 gnd 0.278177f
C5086 vdd.t194 gnd 0.177413f
C5087 vdd.n2747 gnd 0.095882f
C5088 vdd.n2748 gnd 0.054387f
C5089 vdd.n2749 gnd 0.006725f
C5090 vdd.n2750 gnd 0.006725f
C5091 vdd.n2751 gnd 0.006725f
C5092 vdd.n2752 gnd 0.006725f
C5093 vdd.n2753 gnd 0.006725f
C5094 vdd.n2754 gnd 0.006725f
C5095 vdd.n2755 gnd 0.006725f
C5096 vdd.n2756 gnd 0.006725f
C5097 vdd.n2757 gnd 0.006725f
C5098 vdd.n2758 gnd 0.006725f
C5099 vdd.n2759 gnd 0.006725f
C5100 vdd.n2760 gnd 0.006725f
C5101 vdd.n2761 gnd 0.006725f
C5102 vdd.n2762 gnd 0.006725f
C5103 vdd.n2763 gnd 0.006725f
C5104 vdd.n2764 gnd 0.006725f
C5105 vdd.n2765 gnd 0.006725f
C5106 vdd.n2766 gnd 0.006725f
C5107 vdd.n2767 gnd 0.006725f
C5108 vdd.n2768 gnd 0.006725f
C5109 vdd.n2769 gnd 0.006725f
C5110 vdd.n2770 gnd 0.006725f
C5111 vdd.n2771 gnd 0.006725f
C5112 vdd.n2772 gnd 0.006725f
C5113 vdd.n2773 gnd 0.006725f
C5114 vdd.n2774 gnd 0.006725f
C5115 vdd.n2775 gnd 0.006725f
C5116 vdd.n2776 gnd 0.006725f
C5117 vdd.n2777 gnd 0.006725f
C5118 vdd.n2778 gnd 0.006725f
C5119 vdd.n2779 gnd 0.006725f
C5120 vdd.n2780 gnd 0.006725f
C5121 vdd.n2781 gnd 0.006725f
C5122 vdd.n2782 gnd 0.006725f
C5123 vdd.n2783 gnd 0.006725f
C5124 vdd.n2784 gnd 0.006725f
C5125 vdd.n2785 gnd 0.006725f
C5126 vdd.n2786 gnd 0.006725f
C5127 vdd.n2787 gnd 0.006725f
C5128 vdd.n2788 gnd 0.006725f
C5129 vdd.n2789 gnd 0.006725f
C5130 vdd.n2790 gnd 0.006725f
C5131 vdd.n2791 gnd 0.006725f
C5132 vdd.n2792 gnd 0.006725f
C5133 vdd.n2793 gnd 0.006725f
C5134 vdd.n2794 gnd 0.006725f
C5135 vdd.n2795 gnd 0.006725f
C5136 vdd.n2796 gnd 0.006725f
C5137 vdd.n2797 gnd 0.006725f
C5138 vdd.n2798 gnd 0.006725f
C5139 vdd.n2799 gnd 0.006725f
C5140 vdd.n2800 gnd 0.006725f
C5141 vdd.n2801 gnd 0.006725f
C5142 vdd.n2802 gnd 0.006725f
C5143 vdd.n2803 gnd 0.006725f
C5144 vdd.n2804 gnd 0.006725f
C5145 vdd.n2805 gnd 0.006725f
C5146 vdd.n2806 gnd 0.004895f
C5147 vdd.n2807 gnd 0.009611f
C5148 vdd.n2808 gnd 0.005192f
C5149 vdd.n2809 gnd 0.006725f
C5150 vdd.n2810 gnd 0.006725f
C5151 vdd.n2811 gnd 0.006725f
C5152 vdd.n2812 gnd 0.0155f
C5153 vdd.n2813 gnd 0.0155f
C5154 vdd.n2814 gnd 0.014565f
C5155 vdd.n2815 gnd 0.006725f
C5156 vdd.n2816 gnd 0.006725f
C5157 vdd.n2817 gnd 0.006725f
C5158 vdd.n2818 gnd 0.006725f
C5159 vdd.n2819 gnd 0.006725f
C5160 vdd.n2820 gnd 0.006725f
C5161 vdd.n2821 gnd 0.006725f
C5162 vdd.n2822 gnd 0.006725f
C5163 vdd.n2823 gnd 0.006725f
C5164 vdd.n2824 gnd 0.006725f
C5165 vdd.n2825 gnd 0.006725f
C5166 vdd.n2826 gnd 0.006725f
C5167 vdd.n2827 gnd 0.006725f
C5168 vdd.n2828 gnd 0.006725f
C5169 vdd.n2829 gnd 0.006725f
C5170 vdd.n2830 gnd 0.006725f
C5171 vdd.n2831 gnd 0.006725f
C5172 vdd.n2832 gnd 0.006725f
C5173 vdd.n2833 gnd 0.006725f
C5174 vdd.n2834 gnd 0.006725f
C5175 vdd.n2835 gnd 0.006725f
C5176 vdd.n2836 gnd 0.006725f
C5177 vdd.n2837 gnd 0.006725f
C5178 vdd.n2838 gnd 0.006725f
C5179 vdd.n2839 gnd 0.006725f
C5180 vdd.n2840 gnd 0.006725f
C5181 vdd.n2841 gnd 0.006725f
C5182 vdd.n2842 gnd 0.006725f
C5183 vdd.n2843 gnd 0.006725f
C5184 vdd.n2844 gnd 0.006725f
C5185 vdd.n2845 gnd 0.006725f
C5186 vdd.n2846 gnd 0.006725f
C5187 vdd.n2847 gnd 0.006725f
C5188 vdd.n2848 gnd 0.006725f
C5189 vdd.n2849 gnd 0.006725f
C5190 vdd.n2850 gnd 0.006725f
C5191 vdd.n2851 gnd 0.006725f
C5192 vdd.n2852 gnd 0.006725f
C5193 vdd.n2853 gnd 0.006725f
C5194 vdd.n2854 gnd 0.006725f
C5195 vdd.n2855 gnd 0.006725f
C5196 vdd.n2856 gnd 0.006725f
C5197 vdd.n2857 gnd 0.006725f
C5198 vdd.n2858 gnd 0.006725f
C5199 vdd.n2859 gnd 0.006725f
C5200 vdd.n2860 gnd 0.006725f
C5201 vdd.n2861 gnd 0.006725f
C5202 vdd.n2862 gnd 0.006725f
C5203 vdd.n2863 gnd 0.006725f
C5204 vdd.n2864 gnd 0.006725f
C5205 vdd.n2865 gnd 0.006725f
C5206 vdd.n2866 gnd 0.006725f
C5207 vdd.n2867 gnd 0.006725f
C5208 vdd.n2868 gnd 0.006725f
C5209 vdd.n2869 gnd 0.006725f
C5210 vdd.n2870 gnd 0.006725f
C5211 vdd.n2871 gnd 0.006725f
C5212 vdd.n2872 gnd 0.006725f
C5213 vdd.n2873 gnd 0.006725f
C5214 vdd.n2874 gnd 0.006725f
C5215 vdd.n2875 gnd 0.006725f
C5216 vdd.n2876 gnd 0.006725f
C5217 vdd.n2877 gnd 0.006725f
C5218 vdd.n2878 gnd 0.006725f
C5219 vdd.n2879 gnd 0.006725f
C5220 vdd.n2880 gnd 0.006725f
C5221 vdd.n2881 gnd 0.006725f
C5222 vdd.n2882 gnd 0.006725f
C5223 vdd.n2883 gnd 0.006725f
C5224 vdd.n2884 gnd 0.006725f
C5225 vdd.n2885 gnd 0.006725f
C5226 vdd.n2886 gnd 0.006725f
C5227 vdd.n2887 gnd 0.006725f
C5228 vdd.n2888 gnd 0.006725f
C5229 vdd.n2889 gnd 0.006725f
C5230 vdd.n2890 gnd 0.006725f
C5231 vdd.n2891 gnd 0.006725f
C5232 vdd.n2892 gnd 0.006725f
C5233 vdd.n2893 gnd 0.006725f
C5234 vdd.n2894 gnd 0.217297f
C5235 vdd.n2895 gnd 0.006725f
C5236 vdd.n2896 gnd 0.006725f
C5237 vdd.n2897 gnd 0.006725f
C5238 vdd.n2898 gnd 0.006725f
C5239 vdd.n2899 gnd 0.006725f
C5240 vdd.n2900 gnd 0.006725f
C5241 vdd.n2901 gnd 0.006725f
C5242 vdd.n2902 gnd 0.006725f
C5243 vdd.n2903 gnd 0.006725f
C5244 vdd.n2904 gnd 0.006725f
C5245 vdd.n2905 gnd 0.006725f
C5246 vdd.n2906 gnd 0.621571f
C5247 vdd.n2907 gnd 0.006725f
C5248 vdd.n2908 gnd 0.006725f
C5249 vdd.n2909 gnd 0.006725f
C5250 vdd.n2910 gnd 0.006725f
C5251 vdd.n2911 gnd 0.006725f
C5252 vdd.n2912 gnd 0.006725f
C5253 vdd.n2913 gnd 0.006725f
C5254 vdd.n2914 gnd 0.006725f
C5255 vdd.n2915 gnd 0.006725f
C5256 vdd.n2916 gnd 0.006725f
C5257 vdd.n2917 gnd 0.006725f
C5258 vdd.n2918 gnd 0.409327f
C5259 vdd.n2919 gnd 0.006725f
C5260 vdd.n2920 gnd 0.006725f
C5261 vdd.n2921 gnd 0.006725f
C5262 vdd.n2922 gnd 0.006725f
C5263 vdd.n2923 gnd 0.006725f
C5264 vdd.n2924 gnd 0.014565f
C5265 vdd.n2925 gnd 0.0155f
C5266 vdd.n2926 gnd 0.0155f
C5267 vdd.n2927 gnd 0.838868f
C5268 vdd.n2929 gnd 0.006725f
C5269 vdd.n2930 gnd 0.006725f
C5270 vdd.n2931 gnd 0.0155f
C5271 vdd.n2932 gnd 0.014565f
C5272 vdd.n2933 gnd 0.014565f
C5273 vdd.n2934 gnd 0.79844f
C5274 vdd.n2935 gnd 0.014565f
C5275 vdd.n2936 gnd 0.014565f
C5276 vdd.n2937 gnd 0.006725f
C5277 vdd.n2938 gnd 0.006725f
C5278 vdd.n2939 gnd 0.006725f
C5279 vdd.n2940 gnd 0.429541f
C5280 vdd.n2941 gnd 0.006725f
C5281 vdd.n2942 gnd 0.006725f
C5282 vdd.n2943 gnd 0.006725f
C5283 vdd.n2944 gnd 0.006725f
C5284 vdd.n2945 gnd 0.006725f
C5285 vdd.n2946 gnd 0.495235f
C5286 vdd.n2947 gnd 0.006725f
C5287 vdd.n2948 gnd 0.006725f
C5288 vdd.n2949 gnd 0.006725f
C5289 vdd.n2950 gnd 0.006725f
C5290 vdd.n2951 gnd 0.006725f
C5291 vdd.n2952 gnd 0.687265f
C5292 vdd.n2953 gnd 0.006725f
C5293 vdd.n2954 gnd 0.006725f
C5294 vdd.n2955 gnd 0.006725f
C5295 vdd.n2956 gnd 0.006725f
C5296 vdd.n2957 gnd 0.006725f
C5297 vdd.n2958 gnd 0.217297f
C5298 vdd.n2959 gnd 0.006725f
C5299 vdd.n2960 gnd 0.006725f
C5300 vdd.n2961 gnd 0.006725f
C5301 vdd.n2962 gnd 0.006725f
C5302 vdd.n2963 gnd 0.006725f
C5303 vdd.n2964 gnd 0.217297f
C5304 vdd.n2965 gnd 0.006725f
C5305 vdd.n2966 gnd 0.006725f
C5306 vdd.n2967 gnd 0.006725f
C5307 vdd.n2968 gnd 0.006725f
C5308 vdd.n2969 gnd 0.006725f
C5309 vdd.n2970 gnd 0.434594f
C5310 vdd.n2971 gnd 0.006725f
C5311 vdd.n2972 gnd 0.006725f
C5312 vdd.n2973 gnd 0.006725f
C5313 vdd.n2974 gnd 0.006725f
C5314 vdd.n2975 gnd 0.006725f
C5315 vdd.n2976 gnd 0.586197f
C5316 vdd.n2977 gnd 0.006725f
C5317 vdd.n2978 gnd 0.006725f
C5318 vdd.n2979 gnd 0.006725f
C5319 vdd.n2980 gnd 0.006725f
C5320 vdd.n2981 gnd 0.006725f
C5321 vdd.n2982 gnd 0.571036f
C5322 vdd.n2983 gnd 0.006725f
C5323 vdd.n2984 gnd 0.006725f
C5324 vdd.n2985 gnd 0.006725f
C5325 vdd.n2986 gnd 0.006725f
C5326 vdd.n2987 gnd 0.006725f
C5327 vdd.n2988 gnd 0.419434f
C5328 vdd.n2989 gnd 0.006725f
C5329 vdd.n2990 gnd 0.006725f
C5330 vdd.n2991 gnd 0.006725f
C5331 vdd.n2992 gnd 0.006725f
C5332 vdd.n2993 gnd 0.006725f
C5333 vdd.n2994 gnd 0.419434f
C5334 vdd.n2995 gnd 0.006725f
C5335 vdd.n2996 gnd 0.004549f
C5336 vdd.n2997 gnd 0.019482f
C5337 vdd.n2998 gnd 0.005538f
C5338 vdd.n2999 gnd 0.006725f
C5339 vdd.n3000 gnd 0.006725f
C5340 vdd.n3001 gnd 0.571036f
C5341 vdd.n3002 gnd 0.006725f
C5342 vdd.n3003 gnd 0.006725f
C5343 vdd.n3004 gnd 0.006725f
C5344 vdd.n3005 gnd 0.006725f
C5345 vdd.n3006 gnd 0.006725f
C5346 vdd.n3007 gnd 0.687265f
C5347 vdd.n3008 gnd 0.006725f
C5348 vdd.n3009 gnd 0.006725f
C5349 vdd.n3010 gnd 0.006725f
C5350 vdd.n3011 gnd 0.006725f
C5351 vdd.n3012 gnd 0.006725f
C5352 vdd.n3013 gnd 0.651891f
C5353 vdd.n3014 gnd 0.006725f
C5354 vdd.n3015 gnd 0.006725f
C5355 vdd.n3016 gnd 0.006725f
C5356 vdd.n3017 gnd 0.006725f
C5357 vdd.n3018 gnd 0.006725f
C5358 vdd.n3019 gnd 0.500289f
C5359 vdd.n3020 gnd 0.006725f
C5360 vdd.n3021 gnd 0.006725f
C5361 vdd.n3022 gnd 0.006725f
C5362 vdd.n3023 gnd 0.006725f
C5363 vdd.n3024 gnd 0.006725f
C5364 vdd.n3025 gnd 0.348686f
C5365 vdd.n3026 gnd 0.006725f
C5366 vdd.n3027 gnd 0.006725f
C5367 vdd.n3028 gnd 0.006725f
C5368 vdd.n3029 gnd 0.006725f
C5369 vdd.n3030 gnd 0.006725f
C5370 vdd.n3031 gnd 0.687265f
C5371 vdd.n3032 gnd 0.006725f
C5372 vdd.n3033 gnd 0.006725f
C5373 vdd.n3034 gnd 0.006725f
C5374 vdd.n3035 gnd 0.006725f
C5375 vdd.n3036 gnd 0.006725f
C5376 vdd.n3037 gnd 0.006725f
C5377 vdd.n3039 gnd 0.006725f
C5378 vdd.n3040 gnd 0.006725f
C5379 vdd.n3042 gnd 0.006725f
C5380 vdd.n3043 gnd 0.006725f
C5381 vdd.n3046 gnd 0.006725f
C5382 vdd.n3047 gnd 0.006725f
C5383 vdd.n3048 gnd 0.006725f
C5384 vdd.n3049 gnd 0.006725f
C5385 vdd.n3051 gnd 0.006725f
C5386 vdd.n3052 gnd 0.006725f
C5387 vdd.n3053 gnd 0.006725f
C5388 vdd.n3054 gnd 0.006725f
C5389 vdd.n3055 gnd 0.006725f
C5390 vdd.n3056 gnd 0.006725f
C5391 vdd.n3058 gnd 0.006725f
C5392 vdd.n3059 gnd 0.006725f
C5393 vdd.n3060 gnd 0.006725f
C5394 vdd.n3061 gnd 0.006725f
C5395 vdd.n3062 gnd 0.006725f
C5396 vdd.n3063 gnd 0.006725f
C5397 vdd.n3065 gnd 0.006725f
C5398 vdd.n3066 gnd 0.006725f
C5399 vdd.n3067 gnd 0.006725f
C5400 vdd.n3068 gnd 0.006725f
C5401 vdd.n3069 gnd 0.006725f
C5402 vdd.n3070 gnd 0.006725f
C5403 vdd.n3072 gnd 0.006725f
C5404 vdd.n3073 gnd 0.0155f
C5405 vdd.n3074 gnd 0.0155f
C5406 vdd.n3075 gnd 0.014565f
C5407 vdd.n3076 gnd 0.006725f
C5408 vdd.n3077 gnd 0.006725f
C5409 vdd.n3078 gnd 0.006725f
C5410 vdd.n3079 gnd 0.006725f
C5411 vdd.n3080 gnd 0.006725f
C5412 vdd.n3081 gnd 0.006725f
C5413 vdd.n3082 gnd 0.687265f
C5414 vdd.n3083 gnd 0.006725f
C5415 vdd.n3084 gnd 0.006725f
C5416 vdd.n3085 gnd 0.006725f
C5417 vdd.n3086 gnd 0.006725f
C5418 vdd.n3087 gnd 0.006725f
C5419 vdd.n3088 gnd 0.469968f
C5420 vdd.n3089 gnd 0.006725f
C5421 vdd.n3090 gnd 0.006725f
C5422 vdd.n3091 gnd 0.006725f
C5423 vdd.n3092 gnd 0.015417f
C5424 vdd.n3094 gnd 0.0155f
C5425 vdd.n3095 gnd 0.014648f
C5426 vdd.n3096 gnd 0.006725f
C5427 vdd.n3097 gnd 0.005192f
C5428 vdd.n3098 gnd 0.006725f
C5429 vdd.n3100 gnd 0.006725f
C5430 vdd.n3101 gnd 0.006725f
C5431 vdd.n3102 gnd 0.006725f
C5432 vdd.n3103 gnd 0.006725f
C5433 vdd.n3104 gnd 0.006725f
C5434 vdd.n3105 gnd 0.006725f
C5435 vdd.n3107 gnd 0.006725f
C5436 vdd.n3108 gnd 0.006725f
C5437 vdd.n3109 gnd 0.006725f
C5438 vdd.n3110 gnd 0.006725f
C5439 vdd.n3111 gnd 0.006725f
C5440 vdd.n3112 gnd 0.006725f
C5441 vdd.n3114 gnd 0.006725f
C5442 vdd.n3115 gnd 0.006725f
C5443 vdd.n3116 gnd 0.006725f
C5444 vdd.n3117 gnd 0.006725f
C5445 vdd.n3118 gnd 0.006725f
C5446 vdd.n3119 gnd 0.006725f
C5447 vdd.n3121 gnd 0.006725f
C5448 vdd.n3122 gnd 0.006725f
C5449 vdd.n3123 gnd 0.006725f
C5450 vdd.n3124 gnd 0.903467f
C5451 vdd.n3125 gnd 0.031567f
C5452 vdd.n3126 gnd 0.006725f
C5453 vdd.n3127 gnd 0.006725f
C5454 vdd.n3129 gnd 0.006725f
C5455 vdd.n3130 gnd 0.006725f
C5456 vdd.n3131 gnd 0.006725f
C5457 vdd.n3132 gnd 0.006725f
C5458 vdd.n3133 gnd 0.006725f
C5459 vdd.n3134 gnd 0.006725f
C5460 vdd.n3136 gnd 0.006725f
C5461 vdd.n3137 gnd 0.006725f
C5462 vdd.n3138 gnd 0.006725f
C5463 vdd.n3139 gnd 0.006725f
C5464 vdd.n3140 gnd 0.006725f
C5465 vdd.n3141 gnd 0.006725f
C5466 vdd.n3143 gnd 0.006725f
C5467 vdd.n3144 gnd 0.006725f
C5468 vdd.n3145 gnd 0.006725f
C5469 vdd.n3146 gnd 0.006725f
C5470 vdd.n3147 gnd 0.006725f
C5471 vdd.n3148 gnd 0.006725f
C5472 vdd.n3150 gnd 0.006725f
C5473 vdd.n3151 gnd 0.006725f
C5474 vdd.n3153 gnd 0.006725f
C5475 vdd.n3154 gnd 0.006725f
C5476 vdd.n3155 gnd 0.0155f
C5477 vdd.n3156 gnd 0.014565f
C5478 vdd.n3157 gnd 0.014565f
C5479 vdd.n3158 gnd 0.950043f
C5480 vdd.n3159 gnd 0.014565f
C5481 vdd.n3160 gnd 0.0155f
C5482 vdd.n3161 gnd 0.014648f
C5483 vdd.n3162 gnd 0.006725f
C5484 vdd.n3163 gnd 0.005192f
C5485 vdd.n3164 gnd 0.006725f
C5486 vdd.n3166 gnd 0.006725f
C5487 vdd.n3167 gnd 0.006725f
C5488 vdd.n3168 gnd 0.006725f
C5489 vdd.n3169 gnd 0.006725f
C5490 vdd.n3170 gnd 0.006725f
C5491 vdd.n3171 gnd 0.006725f
C5492 vdd.n3173 gnd 0.006725f
C5493 vdd.n3174 gnd 0.006725f
C5494 vdd.n3175 gnd 0.006725f
C5495 vdd.n3176 gnd 0.006725f
C5496 vdd.n3177 gnd 0.006725f
C5497 vdd.n3178 gnd 0.006725f
C5498 vdd.n3180 gnd 0.006725f
C5499 vdd.n3181 gnd 0.006725f
C5500 vdd.n3182 gnd 0.006725f
C5501 vdd.n3183 gnd 0.006725f
C5502 vdd.n3184 gnd 0.006725f
C5503 vdd.n3185 gnd 0.006725f
C5504 vdd.n3187 gnd 0.006725f
C5505 vdd.n3188 gnd 0.006725f
C5506 vdd.n3190 gnd 0.006725f
C5507 vdd.n3191 gnd 0.031567f
C5508 vdd.n3192 gnd 0.903467f
C5509 vdd.n3193 gnd 0.008505f
C5510 vdd.n3194 gnd 0.003781f
C5511 vdd.t168 gnd 0.12167f
C5512 vdd.t169 gnd 0.130031f
C5513 vdd.t167 gnd 0.158899f
C5514 vdd.n3195 gnd 0.203686f
C5515 vdd.n3196 gnd 0.171133f
C5516 vdd.n3197 gnd 0.012258f
C5517 vdd.n3198 gnd 0.00989f
C5518 vdd.n3199 gnd 0.004179f
C5519 vdd.n3200 gnd 0.00796f
C5520 vdd.n3201 gnd 0.00989f
C5521 vdd.n3202 gnd 0.00989f
C5522 vdd.n3203 gnd 0.00796f
C5523 vdd.n3204 gnd 0.00796f
C5524 vdd.n3205 gnd 0.00989f
C5525 vdd.n3207 gnd 0.00989f
C5526 vdd.n3208 gnd 0.00796f
C5527 vdd.n3209 gnd 0.00796f
C5528 vdd.n3210 gnd 0.00796f
C5529 vdd.n3211 gnd 0.00989f
C5530 vdd.n3213 gnd 0.00989f
C5531 vdd.n3215 gnd 0.00989f
C5532 vdd.n3216 gnd 0.00796f
C5533 vdd.n3217 gnd 0.00796f
C5534 vdd.n3218 gnd 0.00796f
C5535 vdd.n3219 gnd 0.00989f
C5536 vdd.n3221 gnd 0.00989f
C5537 vdd.n3223 gnd 0.00989f
C5538 vdd.n3224 gnd 0.00796f
C5539 vdd.n3225 gnd 0.00796f
C5540 vdd.n3226 gnd 0.00796f
C5541 vdd.n3227 gnd 0.00989f
C5542 vdd.n3229 gnd 0.00989f
C5543 vdd.n3230 gnd 0.00989f
C5544 vdd.n3231 gnd 0.00796f
C5545 vdd.n3232 gnd 0.00796f
C5546 vdd.n3233 gnd 0.00989f
C5547 vdd.n3234 gnd 0.00989f
C5548 vdd.n3236 gnd 0.00989f
C5549 vdd.n3237 gnd 0.00796f
C5550 vdd.n3238 gnd 0.00989f
C5551 vdd.n3239 gnd 0.00989f
C5552 vdd.n3240 gnd 0.00989f
C5553 vdd.n3241 gnd 0.016238f
C5554 vdd.n3242 gnd 0.005413f
C5555 vdd.n3243 gnd 0.00989f
C5556 vdd.n3245 gnd 0.00989f
C5557 vdd.n3247 gnd 0.00989f
C5558 vdd.n3248 gnd 0.00796f
C5559 vdd.n3249 gnd 0.00796f
C5560 vdd.n3250 gnd 0.00796f
C5561 vdd.n3251 gnd 0.00989f
C5562 vdd.n3253 gnd 0.00989f
C5563 vdd.n3255 gnd 0.00989f
C5564 vdd.n3256 gnd 0.00796f
C5565 vdd.n3257 gnd 0.00796f
C5566 vdd.n3258 gnd 0.00796f
C5567 vdd.n3259 gnd 0.00989f
C5568 vdd.n3261 gnd 0.00989f
C5569 vdd.n3263 gnd 0.00989f
C5570 vdd.n3264 gnd 0.00796f
C5571 vdd.n3265 gnd 0.00796f
C5572 vdd.n3266 gnd 0.00796f
C5573 vdd.n3267 gnd 0.00989f
C5574 vdd.n3269 gnd 0.00989f
C5575 vdd.n3271 gnd 0.00989f
C5576 vdd.n3272 gnd 0.00796f
C5577 vdd.n3273 gnd 0.00796f
C5578 vdd.n3274 gnd 0.00796f
C5579 vdd.n3275 gnd 0.00989f
C5580 vdd.n3277 gnd 0.00989f
C5581 vdd.n3279 gnd 0.00989f
C5582 vdd.n3280 gnd 0.00796f
C5583 vdd.n3281 gnd 0.00796f
C5584 vdd.n3282 gnd 0.006647f
C5585 vdd.n3283 gnd 0.00989f
C5586 vdd.n3285 gnd 0.00989f
C5587 vdd.n3287 gnd 0.00989f
C5588 vdd.n3288 gnd 0.006647f
C5589 vdd.n3289 gnd 0.00796f
C5590 vdd.n3290 gnd 0.00796f
C5591 vdd.n3291 gnd 0.00989f
C5592 vdd.n3293 gnd 0.00989f
C5593 vdd.n3295 gnd 0.00989f
C5594 vdd.n3296 gnd 0.00796f
C5595 vdd.n3297 gnd 0.00796f
C5596 vdd.n3298 gnd 0.00796f
C5597 vdd.n3299 gnd 0.00989f
C5598 vdd.n3301 gnd 0.00989f
C5599 vdd.n3303 gnd 0.00989f
C5600 vdd.n3304 gnd 0.00796f
C5601 vdd.n3305 gnd 0.00796f
C5602 vdd.n3306 gnd 0.00796f
C5603 vdd.n3307 gnd 0.00989f
C5604 vdd.n3309 gnd 0.00989f
C5605 vdd.n3310 gnd 0.00989f
C5606 vdd.n3311 gnd 0.00796f
C5607 vdd.n3312 gnd 0.00796f
C5608 vdd.n3313 gnd 0.00989f
C5609 vdd.n3314 gnd 0.00989f
C5610 vdd.n3315 gnd 0.00796f
C5611 vdd.n3316 gnd 0.00796f
C5612 vdd.n3317 gnd 0.00989f
C5613 vdd.n3318 gnd 0.00989f
C5614 vdd.n3320 gnd 0.00989f
C5615 vdd.n3321 gnd 0.00796f
C5616 vdd.n3322 gnd 0.006607f
C5617 vdd.n3323 gnd 0.022675f
C5618 vdd.n3324 gnd 0.022521f
C5619 vdd.n3325 gnd 0.006607f
C5620 vdd.n3326 gnd 0.022521f
C5621 vdd.n3327 gnd 1.3341f
C5622 vdd.n3328 gnd 0.022521f
C5623 vdd.n3329 gnd 0.006607f
C5624 vdd.n3330 gnd 0.022521f
C5625 vdd.n3331 gnd 0.00989f
C5626 vdd.n3332 gnd 0.00989f
C5627 vdd.n3333 gnd 0.00796f
C5628 vdd.n3334 gnd 0.00989f
C5629 vdd.n3335 gnd 0.955096f
C5630 vdd.n3336 gnd 0.00989f
C5631 vdd.n3337 gnd 0.00796f
C5632 vdd.n3338 gnd 0.00989f
C5633 vdd.n3339 gnd 0.00989f
C5634 vdd.n3340 gnd 0.00989f
C5635 vdd.n3341 gnd 0.00796f
C5636 vdd.n3342 gnd 0.00989f
C5637 vdd.n3343 gnd 0.985417f
C5638 vdd.n3344 gnd 0.00989f
C5639 vdd.n3345 gnd 0.00796f
C5640 vdd.n3346 gnd 0.00989f
C5641 vdd.n3347 gnd 0.00989f
C5642 vdd.n3348 gnd 0.00989f
C5643 vdd.n3349 gnd 0.00796f
C5644 vdd.n3350 gnd 0.00989f
C5645 vdd.t21 gnd 0.505342f
C5646 vdd.n3351 gnd 0.813601f
C5647 vdd.n3352 gnd 0.00989f
C5648 vdd.n3353 gnd 0.00796f
C5649 vdd.n3354 gnd 0.00989f
C5650 vdd.n3355 gnd 0.00989f
C5651 vdd.n3356 gnd 0.00989f
C5652 vdd.n3357 gnd 0.00796f
C5653 vdd.n3358 gnd 0.00989f
C5654 vdd.n3359 gnd 0.641784f
C5655 vdd.n3360 gnd 0.00989f
C5656 vdd.n3361 gnd 0.00796f
C5657 vdd.n3362 gnd 0.00989f
C5658 vdd.n3363 gnd 0.00989f
C5659 vdd.n3364 gnd 0.00989f
C5660 vdd.n3365 gnd 0.00796f
C5661 vdd.n3366 gnd 0.00989f
C5662 vdd.n3367 gnd 0.803494f
C5663 vdd.n3368 gnd 0.540716f
C5664 vdd.n3369 gnd 0.00989f
C5665 vdd.n3370 gnd 0.00796f
C5666 vdd.n3371 gnd 0.00989f
C5667 vdd.n3372 gnd 0.00989f
C5668 vdd.n3373 gnd 0.00989f
C5669 vdd.n3374 gnd 0.00796f
C5670 vdd.n3375 gnd 0.00989f
C5671 vdd.n3376 gnd 0.712532f
C5672 vdd.n3377 gnd 0.00989f
C5673 vdd.n3378 gnd 0.00796f
C5674 vdd.n3379 gnd 0.00989f
C5675 vdd.n3380 gnd 0.00989f
C5676 vdd.n3381 gnd 0.00989f
C5677 vdd.n3382 gnd 0.00989f
C5678 vdd.n3383 gnd 0.00989f
C5679 vdd.n3384 gnd 0.00796f
C5680 vdd.n3385 gnd 0.00796f
C5681 vdd.n3386 gnd 0.00989f
C5682 vdd.t31 gnd 0.505342f
C5683 vdd.n3387 gnd 0.838868f
C5684 vdd.n3388 gnd 0.00989f
C5685 vdd.n3389 gnd 0.00796f
C5686 vdd.n3390 gnd 0.00989f
C5687 vdd.n3391 gnd 0.00989f
C5688 vdd.n3392 gnd 0.00989f
C5689 vdd.n3393 gnd 0.00796f
C5690 vdd.n3394 gnd 0.00989f
C5691 vdd.n3395 gnd 0.793387f
C5692 vdd.n3396 gnd 0.00989f
C5693 vdd.n3397 gnd 0.00989f
C5694 vdd.n3398 gnd 0.00796f
C5695 vdd.n3399 gnd 0.00796f
C5696 vdd.n3400 gnd 0.00796f
C5697 vdd.n3401 gnd 0.00989f
C5698 vdd.n3402 gnd 0.00989f
C5699 vdd.n3403 gnd 0.00989f
C5700 vdd.n3404 gnd 0.00989f
C5701 vdd.n3405 gnd 0.00796f
C5702 vdd.n3406 gnd 0.00796f
C5703 vdd.n3407 gnd 0.00796f
C5704 vdd.n3408 gnd 0.00989f
C5705 vdd.n3409 gnd 0.00989f
C5706 vdd.n3410 gnd 0.00989f
C5707 vdd.n3411 gnd 0.00989f
C5708 vdd.n3412 gnd 0.00796f
C5709 vdd.n3413 gnd 0.00796f
C5710 vdd.n3414 gnd 0.00796f
C5711 vdd.n3415 gnd 0.00989f
C5712 vdd.n3416 gnd 0.00989f
C5713 vdd.n3417 gnd 0.00989f
C5714 vdd.n3418 gnd 0.838868f
C5715 vdd.n3419 gnd 0.00989f
C5716 vdd.n3420 gnd 0.00796f
C5717 vdd.n3421 gnd 0.00796f
C5718 vdd.n3422 gnd 0.00796f
C5719 vdd.n3423 gnd 0.00989f
C5720 vdd.n3424 gnd 0.00989f
C5721 vdd.n3425 gnd 0.00989f
C5722 vdd.n3426 gnd 0.00989f
C5723 vdd.n3427 gnd 0.00796f
C5724 vdd.n3428 gnd 0.00796f
C5725 vdd.n3429 gnd 0.006607f
C5726 vdd.n3430 gnd 0.022521f
C5727 vdd.n3431 gnd 0.022675f
C5728 vdd.n3432 gnd 0.003781f
C5729 vdd.n3433 gnd 0.022675f
C5730 vdd.n3435 gnd 2.23361f
C5731 vdd.n3436 gnd 1.3341f
C5732 vdd.n3437 gnd 0.661998f
C5733 vdd.n3438 gnd 0.00989f
C5734 vdd.n3439 gnd 0.00796f
C5735 vdd.n3440 gnd 0.00796f
C5736 vdd.n3441 gnd 0.00796f
C5737 vdd.n3442 gnd 0.00989f
C5738 vdd.n3443 gnd 1.01068f
C5739 vdd.n3444 gnd 1.01068f
C5740 vdd.n3445 gnd 0.581143f
C5741 vdd.n3446 gnd 0.00989f
C5742 vdd.n3447 gnd 0.00796f
C5743 vdd.n3448 gnd 0.00796f
C5744 vdd.n3449 gnd 0.00796f
C5745 vdd.n3450 gnd 0.00989f
C5746 vdd.n3451 gnd 0.601357f
C5747 vdd.n3452 gnd 0.742853f
C5748 vdd.t61 gnd 0.505342f
C5749 vdd.n3453 gnd 0.773173f
C5750 vdd.n3454 gnd 0.00989f
C5751 vdd.n3455 gnd 0.00796f
C5752 vdd.n3456 gnd 0.00796f
C5753 vdd.n3457 gnd 0.00796f
C5754 vdd.n3458 gnd 0.00989f
C5755 vdd.n3459 gnd 0.838868f
C5756 vdd.t72 gnd 0.505342f
C5757 vdd.n3460 gnd 0.611464f
C5758 vdd.n3461 gnd 0.732746f
C5759 vdd.n3462 gnd 0.00989f
C5760 vdd.n3463 gnd 0.00796f
C5761 vdd.n3464 gnd 0.00796f
C5762 vdd.n3465 gnd 0.00796f
C5763 vdd.n3466 gnd 0.00989f
C5764 vdd.n3467 gnd 0.56093f
C5765 vdd.t27 gnd 0.505342f
C5766 vdd.n3468 gnd 0.838868f
C5767 vdd.t104 gnd 0.505342f
C5768 vdd.n3469 gnd 0.621571f
C5769 vdd.n3470 gnd 0.00989f
C5770 vdd.n3471 gnd 0.00796f
C5771 vdd.n3472 gnd 0.007601f
C5772 vdd.n3473 gnd 0.583334f
C5773 vdd.n3474 gnd 2.59397f
C5774 a_n8300_8799.t37 gnd 0.112772f
C5775 a_n8300_8799.t27 gnd 0.112772f
C5776 a_n8300_8799.t26 gnd 0.112772f
C5777 a_n8300_8799.n0 gnd 0.998708f
C5778 a_n8300_8799.t32 gnd 0.112772f
C5779 a_n8300_8799.t31 gnd 0.112772f
C5780 a_n8300_8799.n1 gnd 0.996491f
C5781 a_n8300_8799.n2 gnd 0.793753f
C5782 a_n8300_8799.t0 gnd 0.144992f
C5783 a_n8300_8799.t18 gnd 0.144992f
C5784 a_n8300_8799.n3 gnd 1.14358f
C5785 a_n8300_8799.t1 gnd 0.144992f
C5786 a_n8300_8799.t11 gnd 0.144992f
C5787 a_n8300_8799.n4 gnd 1.14169f
C5788 a_n8300_8799.n5 gnd 1.02624f
C5789 a_n8300_8799.t6 gnd 0.144992f
C5790 a_n8300_8799.t7 gnd 0.144992f
C5791 a_n8300_8799.n6 gnd 1.14169f
C5792 a_n8300_8799.n7 gnd 0.505853f
C5793 a_n8300_8799.t14 gnd 0.144992f
C5794 a_n8300_8799.t19 gnd 0.144992f
C5795 a_n8300_8799.n8 gnd 1.14169f
C5796 a_n8300_8799.n9 gnd 0.505853f
C5797 a_n8300_8799.t9 gnd 0.144992f
C5798 a_n8300_8799.t13 gnd 0.144992f
C5799 a_n8300_8799.n10 gnd 1.14169f
C5800 a_n8300_8799.n11 gnd 3.48625f
C5801 a_n8300_8799.t3 gnd 0.144992f
C5802 a_n8300_8799.t12 gnd 0.144992f
C5803 a_n8300_8799.n12 gnd 1.14358f
C5804 a_n8300_8799.t4 gnd 0.144992f
C5805 a_n8300_8799.t10 gnd 0.144992f
C5806 a_n8300_8799.n13 gnd 1.14169f
C5807 a_n8300_8799.n14 gnd 1.02624f
C5808 a_n8300_8799.t16 gnd 0.144992f
C5809 a_n8300_8799.t15 gnd 0.144992f
C5810 a_n8300_8799.n15 gnd 1.14169f
C5811 a_n8300_8799.n16 gnd 0.505853f
C5812 a_n8300_8799.t2 gnd 0.144992f
C5813 a_n8300_8799.t17 gnd 0.144992f
C5814 a_n8300_8799.n17 gnd 1.14169f
C5815 a_n8300_8799.n18 gnd 0.505853f
C5816 a_n8300_8799.t5 gnd 0.144992f
C5817 a_n8300_8799.t8 gnd 0.144992f
C5818 a_n8300_8799.n19 gnd 1.14169f
C5819 a_n8300_8799.n20 gnd 2.26f
C5820 a_n8300_8799.n21 gnd 7.02726f
C5821 a_n8300_8799.n22 gnd 0.05226f
C5822 a_n8300_8799.t68 gnd 0.601206f
C5823 a_n8300_8799.n23 gnd 0.26851f
C5824 a_n8300_8799.n24 gnd 0.05226f
C5825 a_n8300_8799.n25 gnd 0.011859f
C5826 a_n8300_8799.t102 gnd 0.601206f
C5827 a_n8300_8799.n26 gnd 0.05226f
C5828 a_n8300_8799.t122 gnd 0.601206f
C5829 a_n8300_8799.n27 gnd 0.268349f
C5830 a_n8300_8799.t79 gnd 0.601206f
C5831 a_n8300_8799.n28 gnd 0.05226f
C5832 a_n8300_8799.n29 gnd 0.011859f
C5833 a_n8300_8799.t81 gnd 0.601206f
C5834 a_n8300_8799.n30 gnd 0.05226f
C5835 a_n8300_8799.t93 gnd 0.601206f
C5836 a_n8300_8799.n31 gnd 0.263516f
C5837 a_n8300_8799.t123 gnd 0.601206f
C5838 a_n8300_8799.n32 gnd 0.05226f
C5839 a_n8300_8799.t128 gnd 0.601206f
C5840 a_n8300_8799.n33 gnd 0.267705f
C5841 a_n8300_8799.t96 gnd 0.612585f
C5842 a_n8300_8799.n34 gnd 0.252052f
C5843 a_n8300_8799.n35 gnd 0.170881f
C5844 a_n8300_8799.n36 gnd 0.011859f
C5845 a_n8300_8799.t66 gnd 0.601206f
C5846 a_n8300_8799.n37 gnd 0.26851f
C5847 a_n8300_8799.n38 gnd 0.011859f
C5848 a_n8300_8799.n39 gnd 0.05226f
C5849 a_n8300_8799.n40 gnd 0.05226f
C5850 a_n8300_8799.n41 gnd 0.05226f
C5851 a_n8300_8799.n42 gnd 0.268027f
C5852 a_n8300_8799.n43 gnd 0.011859f
C5853 a_n8300_8799.t124 gnd 0.601206f
C5854 a_n8300_8799.n44 gnd 0.26851f
C5855 a_n8300_8799.n45 gnd 0.05226f
C5856 a_n8300_8799.n46 gnd 0.05226f
C5857 a_n8300_8799.n47 gnd 0.05226f
C5858 a_n8300_8799.n48 gnd 0.263194f
C5859 a_n8300_8799.t105 gnd 0.601206f
C5860 a_n8300_8799.n49 gnd 0.268349f
C5861 a_n8300_8799.n50 gnd 0.011859f
C5862 a_n8300_8799.n51 gnd 0.05226f
C5863 a_n8300_8799.n52 gnd 0.05226f
C5864 a_n8300_8799.n53 gnd 0.05226f
C5865 a_n8300_8799.n54 gnd 0.263194f
C5866 a_n8300_8799.n55 gnd 0.011859f
C5867 a_n8300_8799.t80 gnd 0.601206f
C5868 a_n8300_8799.n56 gnd 0.26851f
C5869 a_n8300_8799.n57 gnd 0.05226f
C5870 a_n8300_8799.n58 gnd 0.05226f
C5871 a_n8300_8799.n59 gnd 0.05226f
C5872 a_n8300_8799.n60 gnd 0.268027f
C5873 a_n8300_8799.t67 gnd 0.601206f
C5874 a_n8300_8799.n61 gnd 0.263516f
C5875 a_n8300_8799.n62 gnd 0.011859f
C5876 a_n8300_8799.n63 gnd 0.05226f
C5877 a_n8300_8799.n64 gnd 0.05226f
C5878 a_n8300_8799.n65 gnd 0.05226f
C5879 a_n8300_8799.n66 gnd 0.011859f
C5880 a_n8300_8799.t99 gnd 0.601206f
C5881 a_n8300_8799.n67 gnd 0.267705f
C5882 a_n8300_8799.t44 gnd 0.601206f
C5883 a_n8300_8799.n68 gnd 0.263033f
C5884 a_n8300_8799.n69 gnd 0.301112f
C5885 a_n8300_8799.n70 gnd 0.05226f
C5886 a_n8300_8799.t78 gnd 0.601206f
C5887 a_n8300_8799.n71 gnd 0.26851f
C5888 a_n8300_8799.n72 gnd 0.05226f
C5889 a_n8300_8799.n73 gnd 0.011859f
C5890 a_n8300_8799.t117 gnd 0.601206f
C5891 a_n8300_8799.n74 gnd 0.05226f
C5892 a_n8300_8799.t134 gnd 0.601206f
C5893 a_n8300_8799.n75 gnd 0.268349f
C5894 a_n8300_8799.t85 gnd 0.601206f
C5895 a_n8300_8799.n76 gnd 0.05226f
C5896 a_n8300_8799.n77 gnd 0.011859f
C5897 a_n8300_8799.t89 gnd 0.601206f
C5898 a_n8300_8799.n78 gnd 0.05226f
C5899 a_n8300_8799.t103 gnd 0.601206f
C5900 a_n8300_8799.n79 gnd 0.263516f
C5901 a_n8300_8799.t136 gnd 0.601206f
C5902 a_n8300_8799.n80 gnd 0.05226f
C5903 a_n8300_8799.t139 gnd 0.601206f
C5904 a_n8300_8799.n81 gnd 0.267705f
C5905 a_n8300_8799.t109 gnd 0.612585f
C5906 a_n8300_8799.n82 gnd 0.252052f
C5907 a_n8300_8799.n83 gnd 0.170881f
C5908 a_n8300_8799.n84 gnd 0.011859f
C5909 a_n8300_8799.t74 gnd 0.601206f
C5910 a_n8300_8799.n85 gnd 0.26851f
C5911 a_n8300_8799.n86 gnd 0.011859f
C5912 a_n8300_8799.n87 gnd 0.05226f
C5913 a_n8300_8799.n88 gnd 0.05226f
C5914 a_n8300_8799.n89 gnd 0.05226f
C5915 a_n8300_8799.n90 gnd 0.268027f
C5916 a_n8300_8799.n91 gnd 0.011859f
C5917 a_n8300_8799.t138 gnd 0.601206f
C5918 a_n8300_8799.n92 gnd 0.26851f
C5919 a_n8300_8799.n93 gnd 0.05226f
C5920 a_n8300_8799.n94 gnd 0.05226f
C5921 a_n8300_8799.n95 gnd 0.05226f
C5922 a_n8300_8799.n96 gnd 0.263194f
C5923 a_n8300_8799.t119 gnd 0.601206f
C5924 a_n8300_8799.n97 gnd 0.268349f
C5925 a_n8300_8799.n98 gnd 0.011859f
C5926 a_n8300_8799.n99 gnd 0.05226f
C5927 a_n8300_8799.n100 gnd 0.05226f
C5928 a_n8300_8799.n101 gnd 0.05226f
C5929 a_n8300_8799.n102 gnd 0.263194f
C5930 a_n8300_8799.n103 gnd 0.011859f
C5931 a_n8300_8799.t86 gnd 0.601206f
C5932 a_n8300_8799.n104 gnd 0.26851f
C5933 a_n8300_8799.n105 gnd 0.05226f
C5934 a_n8300_8799.n106 gnd 0.05226f
C5935 a_n8300_8799.n107 gnd 0.05226f
C5936 a_n8300_8799.n108 gnd 0.268027f
C5937 a_n8300_8799.t77 gnd 0.601206f
C5938 a_n8300_8799.n109 gnd 0.263516f
C5939 a_n8300_8799.n110 gnd 0.011859f
C5940 a_n8300_8799.n111 gnd 0.05226f
C5941 a_n8300_8799.n112 gnd 0.05226f
C5942 a_n8300_8799.n113 gnd 0.05226f
C5943 a_n8300_8799.n114 gnd 0.011859f
C5944 a_n8300_8799.t115 gnd 0.601206f
C5945 a_n8300_8799.n115 gnd 0.267705f
C5946 a_n8300_8799.t52 gnd 0.601206f
C5947 a_n8300_8799.n116 gnd 0.263033f
C5948 a_n8300_8799.n117 gnd 0.135393f
C5949 a_n8300_8799.n118 gnd 0.905483f
C5950 a_n8300_8799.n119 gnd 0.05226f
C5951 a_n8300_8799.t104 gnd 0.601206f
C5952 a_n8300_8799.n120 gnd 0.26851f
C5953 a_n8300_8799.n121 gnd 0.05226f
C5954 a_n8300_8799.n122 gnd 0.011859f
C5955 a_n8300_8799.t90 gnd 0.601206f
C5956 a_n8300_8799.n123 gnd 0.05226f
C5957 a_n8300_8799.t125 gnd 0.601206f
C5958 a_n8300_8799.n124 gnd 0.268349f
C5959 a_n8300_8799.t58 gnd 0.601206f
C5960 a_n8300_8799.n125 gnd 0.05226f
C5961 a_n8300_8799.n126 gnd 0.011859f
C5962 a_n8300_8799.t118 gnd 0.601206f
C5963 a_n8300_8799.n127 gnd 0.05226f
C5964 a_n8300_8799.t53 gnd 0.601206f
C5965 a_n8300_8799.n128 gnd 0.263516f
C5966 a_n8300_8799.t100 gnd 0.601206f
C5967 a_n8300_8799.n129 gnd 0.05226f
C5968 a_n8300_8799.t70 gnd 0.601206f
C5969 a_n8300_8799.n130 gnd 0.267705f
C5970 a_n8300_8799.t111 gnd 0.612585f
C5971 a_n8300_8799.n131 gnd 0.252052f
C5972 a_n8300_8799.n132 gnd 0.170881f
C5973 a_n8300_8799.n133 gnd 0.011859f
C5974 a_n8300_8799.t87 gnd 0.601206f
C5975 a_n8300_8799.n134 gnd 0.26851f
C5976 a_n8300_8799.n135 gnd 0.011859f
C5977 a_n8300_8799.n136 gnd 0.05226f
C5978 a_n8300_8799.n137 gnd 0.05226f
C5979 a_n8300_8799.n138 gnd 0.05226f
C5980 a_n8300_8799.n139 gnd 0.268027f
C5981 a_n8300_8799.n140 gnd 0.011859f
C5982 a_n8300_8799.t83 gnd 0.601206f
C5983 a_n8300_8799.n141 gnd 0.26851f
C5984 a_n8300_8799.n142 gnd 0.05226f
C5985 a_n8300_8799.n143 gnd 0.05226f
C5986 a_n8300_8799.n144 gnd 0.05226f
C5987 a_n8300_8799.n145 gnd 0.263194f
C5988 a_n8300_8799.t75 gnd 0.601206f
C5989 a_n8300_8799.n146 gnd 0.268349f
C5990 a_n8300_8799.n147 gnd 0.011859f
C5991 a_n8300_8799.n148 gnd 0.05226f
C5992 a_n8300_8799.n149 gnd 0.05226f
C5993 a_n8300_8799.n150 gnd 0.05226f
C5994 a_n8300_8799.n151 gnd 0.263194f
C5995 a_n8300_8799.n152 gnd 0.011859f
C5996 a_n8300_8799.t45 gnd 0.601206f
C5997 a_n8300_8799.n153 gnd 0.26851f
C5998 a_n8300_8799.n154 gnd 0.05226f
C5999 a_n8300_8799.n155 gnd 0.05226f
C6000 a_n8300_8799.n156 gnd 0.05226f
C6001 a_n8300_8799.n157 gnd 0.268027f
C6002 a_n8300_8799.t127 gnd 0.601206f
C6003 a_n8300_8799.n158 gnd 0.263516f
C6004 a_n8300_8799.n159 gnd 0.011859f
C6005 a_n8300_8799.n160 gnd 0.05226f
C6006 a_n8300_8799.n161 gnd 0.05226f
C6007 a_n8300_8799.n162 gnd 0.05226f
C6008 a_n8300_8799.n163 gnd 0.011859f
C6009 a_n8300_8799.t133 gnd 0.601206f
C6010 a_n8300_8799.n164 gnd 0.267705f
C6011 a_n8300_8799.t84 gnd 0.601206f
C6012 a_n8300_8799.n165 gnd 0.263033f
C6013 a_n8300_8799.n166 gnd 0.135393f
C6014 a_n8300_8799.n167 gnd 1.76515f
C6015 a_n8300_8799.n168 gnd 0.05226f
C6016 a_n8300_8799.t94 gnd 0.601206f
C6017 a_n8300_8799.t47 gnd 0.601206f
C6018 a_n8300_8799.t98 gnd 0.601206f
C6019 a_n8300_8799.n169 gnd 0.26851f
C6020 a_n8300_8799.n170 gnd 0.05226f
C6021 a_n8300_8799.t97 gnd 0.601206f
C6022 a_n8300_8799.t49 gnd 0.601206f
C6023 a_n8300_8799.n171 gnd 0.05226f
C6024 a_n8300_8799.t48 gnd 0.601206f
C6025 a_n8300_8799.n172 gnd 0.26851f
C6026 a_n8300_8799.n173 gnd 0.05226f
C6027 a_n8300_8799.t116 gnd 0.601206f
C6028 a_n8300_8799.t61 gnd 0.601206f
C6029 a_n8300_8799.n174 gnd 0.05226f
C6030 a_n8300_8799.t51 gnd 0.601206f
C6031 a_n8300_8799.n175 gnd 0.268349f
C6032 a_n8300_8799.n176 gnd 0.05226f
C6033 a_n8300_8799.t120 gnd 0.601206f
C6034 a_n8300_8799.t82 gnd 0.601206f
C6035 a_n8300_8799.n177 gnd 0.05226f
C6036 a_n8300_8799.t62 gnd 0.601206f
C6037 a_n8300_8799.n178 gnd 0.268027f
C6038 a_n8300_8799.n179 gnd 0.05226f
C6039 a_n8300_8799.t137 gnd 0.601206f
C6040 a_n8300_8799.t95 gnd 0.601206f
C6041 a_n8300_8799.n180 gnd 0.05226f
C6042 a_n8300_8799.t64 gnd 0.601206f
C6043 a_n8300_8799.n181 gnd 0.267705f
C6044 a_n8300_8799.t131 gnd 0.612585f
C6045 a_n8300_8799.n182 gnd 0.252052f
C6046 a_n8300_8799.n183 gnd 0.170881f
C6047 a_n8300_8799.n184 gnd 0.011859f
C6048 a_n8300_8799.n185 gnd 0.26851f
C6049 a_n8300_8799.n186 gnd 0.011859f
C6050 a_n8300_8799.n187 gnd 0.263516f
C6051 a_n8300_8799.n188 gnd 0.05226f
C6052 a_n8300_8799.n189 gnd 0.05226f
C6053 a_n8300_8799.n190 gnd 0.05226f
C6054 a_n8300_8799.n191 gnd 0.011859f
C6055 a_n8300_8799.n192 gnd 0.26851f
C6056 a_n8300_8799.n193 gnd 0.011859f
C6057 a_n8300_8799.n194 gnd 0.263194f
C6058 a_n8300_8799.n195 gnd 0.05226f
C6059 a_n8300_8799.n196 gnd 0.05226f
C6060 a_n8300_8799.n197 gnd 0.05226f
C6061 a_n8300_8799.n198 gnd 0.011859f
C6062 a_n8300_8799.n199 gnd 0.268349f
C6063 a_n8300_8799.n200 gnd 0.263194f
C6064 a_n8300_8799.n201 gnd 0.011859f
C6065 a_n8300_8799.n202 gnd 0.05226f
C6066 a_n8300_8799.n203 gnd 0.05226f
C6067 a_n8300_8799.n204 gnd 0.05226f
C6068 a_n8300_8799.n205 gnd 0.011859f
C6069 a_n8300_8799.n206 gnd 0.268027f
C6070 a_n8300_8799.n207 gnd 0.263516f
C6071 a_n8300_8799.n208 gnd 0.011859f
C6072 a_n8300_8799.n209 gnd 0.05226f
C6073 a_n8300_8799.n210 gnd 0.05226f
C6074 a_n8300_8799.n211 gnd 0.05226f
C6075 a_n8300_8799.n212 gnd 0.011859f
C6076 a_n8300_8799.n213 gnd 0.267705f
C6077 a_n8300_8799.n214 gnd 0.263033f
C6078 a_n8300_8799.n215 gnd 0.301112f
C6079 a_n8300_8799.n216 gnd 0.05226f
C6080 a_n8300_8799.t107 gnd 0.601206f
C6081 a_n8300_8799.t55 gnd 0.601206f
C6082 a_n8300_8799.t114 gnd 0.601206f
C6083 a_n8300_8799.n217 gnd 0.26851f
C6084 a_n8300_8799.n218 gnd 0.05226f
C6085 a_n8300_8799.t113 gnd 0.601206f
C6086 a_n8300_8799.t57 gnd 0.601206f
C6087 a_n8300_8799.n219 gnd 0.05226f
C6088 a_n8300_8799.t56 gnd 0.601206f
C6089 a_n8300_8799.n220 gnd 0.26851f
C6090 a_n8300_8799.n221 gnd 0.05226f
C6091 a_n8300_8799.t130 gnd 0.601206f
C6092 a_n8300_8799.t69 gnd 0.601206f
C6093 a_n8300_8799.n222 gnd 0.05226f
C6094 a_n8300_8799.t60 gnd 0.601206f
C6095 a_n8300_8799.n223 gnd 0.268349f
C6096 a_n8300_8799.n224 gnd 0.05226f
C6097 a_n8300_8799.t132 gnd 0.601206f
C6098 a_n8300_8799.t92 gnd 0.601206f
C6099 a_n8300_8799.n225 gnd 0.05226f
C6100 a_n8300_8799.t72 gnd 0.601206f
C6101 a_n8300_8799.n226 gnd 0.268027f
C6102 a_n8300_8799.n227 gnd 0.05226f
C6103 a_n8300_8799.t50 gnd 0.601206f
C6104 a_n8300_8799.t108 gnd 0.601206f
C6105 a_n8300_8799.n228 gnd 0.05226f
C6106 a_n8300_8799.t73 gnd 0.601206f
C6107 a_n8300_8799.n229 gnd 0.267705f
C6108 a_n8300_8799.t46 gnd 0.612585f
C6109 a_n8300_8799.n230 gnd 0.252052f
C6110 a_n8300_8799.n231 gnd 0.170881f
C6111 a_n8300_8799.n232 gnd 0.011859f
C6112 a_n8300_8799.n233 gnd 0.26851f
C6113 a_n8300_8799.n234 gnd 0.011859f
C6114 a_n8300_8799.n235 gnd 0.263516f
C6115 a_n8300_8799.n236 gnd 0.05226f
C6116 a_n8300_8799.n237 gnd 0.05226f
C6117 a_n8300_8799.n238 gnd 0.05226f
C6118 a_n8300_8799.n239 gnd 0.011859f
C6119 a_n8300_8799.n240 gnd 0.26851f
C6120 a_n8300_8799.n241 gnd 0.011859f
C6121 a_n8300_8799.n242 gnd 0.263194f
C6122 a_n8300_8799.n243 gnd 0.05226f
C6123 a_n8300_8799.n244 gnd 0.05226f
C6124 a_n8300_8799.n245 gnd 0.05226f
C6125 a_n8300_8799.n246 gnd 0.011859f
C6126 a_n8300_8799.n247 gnd 0.268349f
C6127 a_n8300_8799.n248 gnd 0.263194f
C6128 a_n8300_8799.n249 gnd 0.011859f
C6129 a_n8300_8799.n250 gnd 0.05226f
C6130 a_n8300_8799.n251 gnd 0.05226f
C6131 a_n8300_8799.n252 gnd 0.05226f
C6132 a_n8300_8799.n253 gnd 0.011859f
C6133 a_n8300_8799.n254 gnd 0.268027f
C6134 a_n8300_8799.n255 gnd 0.263516f
C6135 a_n8300_8799.n256 gnd 0.011859f
C6136 a_n8300_8799.n257 gnd 0.05226f
C6137 a_n8300_8799.n258 gnd 0.05226f
C6138 a_n8300_8799.n259 gnd 0.05226f
C6139 a_n8300_8799.n260 gnd 0.011859f
C6140 a_n8300_8799.n261 gnd 0.267705f
C6141 a_n8300_8799.n262 gnd 0.263033f
C6142 a_n8300_8799.n263 gnd 0.135393f
C6143 a_n8300_8799.n264 gnd 0.905483f
C6144 a_n8300_8799.n265 gnd 0.05226f
C6145 a_n8300_8799.t65 gnd 0.601206f
C6146 a_n8300_8799.t135 gnd 0.601206f
C6147 a_n8300_8799.t106 gnd 0.601206f
C6148 a_n8300_8799.n266 gnd 0.26851f
C6149 a_n8300_8799.n267 gnd 0.05226f
C6150 a_n8300_8799.t129 gnd 0.601206f
C6151 a_n8300_8799.t91 gnd 0.601206f
C6152 a_n8300_8799.n268 gnd 0.05226f
C6153 a_n8300_8799.t112 gnd 0.601206f
C6154 a_n8300_8799.n269 gnd 0.26851f
C6155 a_n8300_8799.n270 gnd 0.05226f
C6156 a_n8300_8799.t59 gnd 0.601206f
C6157 a_n8300_8799.t126 gnd 0.601206f
C6158 a_n8300_8799.n271 gnd 0.05226f
C6159 a_n8300_8799.t76 gnd 0.601206f
C6160 a_n8300_8799.n272 gnd 0.268349f
C6161 a_n8300_8799.n273 gnd 0.05226f
C6162 a_n8300_8799.t121 gnd 0.601206f
C6163 a_n8300_8799.t63 gnd 0.601206f
C6164 a_n8300_8799.n274 gnd 0.05226f
C6165 a_n8300_8799.t101 gnd 0.601206f
C6166 a_n8300_8799.n275 gnd 0.268027f
C6167 a_n8300_8799.n276 gnd 0.05226f
C6168 a_n8300_8799.t54 gnd 0.601206f
C6169 a_n8300_8799.t88 gnd 0.601206f
C6170 a_n8300_8799.n277 gnd 0.05226f
C6171 a_n8300_8799.t71 gnd 0.601206f
C6172 a_n8300_8799.n278 gnd 0.267705f
C6173 a_n8300_8799.t110 gnd 0.612585f
C6174 a_n8300_8799.n279 gnd 0.252052f
C6175 a_n8300_8799.n280 gnd 0.170881f
C6176 a_n8300_8799.n281 gnd 0.011859f
C6177 a_n8300_8799.n282 gnd 0.26851f
C6178 a_n8300_8799.n283 gnd 0.011859f
C6179 a_n8300_8799.n284 gnd 0.263516f
C6180 a_n8300_8799.n285 gnd 0.05226f
C6181 a_n8300_8799.n286 gnd 0.05226f
C6182 a_n8300_8799.n287 gnd 0.05226f
C6183 a_n8300_8799.n288 gnd 0.011859f
C6184 a_n8300_8799.n289 gnd 0.26851f
C6185 a_n8300_8799.n290 gnd 0.011859f
C6186 a_n8300_8799.n291 gnd 0.263194f
C6187 a_n8300_8799.n292 gnd 0.05226f
C6188 a_n8300_8799.n293 gnd 0.05226f
C6189 a_n8300_8799.n294 gnd 0.05226f
C6190 a_n8300_8799.n295 gnd 0.011859f
C6191 a_n8300_8799.n296 gnd 0.268349f
C6192 a_n8300_8799.n297 gnd 0.263194f
C6193 a_n8300_8799.n298 gnd 0.011859f
C6194 a_n8300_8799.n299 gnd 0.05226f
C6195 a_n8300_8799.n300 gnd 0.05226f
C6196 a_n8300_8799.n301 gnd 0.05226f
C6197 a_n8300_8799.n302 gnd 0.011859f
C6198 a_n8300_8799.n303 gnd 0.268027f
C6199 a_n8300_8799.n304 gnd 0.263516f
C6200 a_n8300_8799.n305 gnd 0.011859f
C6201 a_n8300_8799.n306 gnd 0.05226f
C6202 a_n8300_8799.n307 gnd 0.05226f
C6203 a_n8300_8799.n308 gnd 0.05226f
C6204 a_n8300_8799.n309 gnd 0.011859f
C6205 a_n8300_8799.n310 gnd 0.267705f
C6206 a_n8300_8799.n311 gnd 0.263033f
C6207 a_n8300_8799.n312 gnd 0.135393f
C6208 a_n8300_8799.n313 gnd 1.28373f
C6209 a_n8300_8799.n314 gnd 15.762001f
C6210 a_n8300_8799.n315 gnd 4.39996f
C6211 a_n8300_8799.t28 gnd 0.112772f
C6212 a_n8300_8799.t29 gnd 0.112772f
C6213 a_n8300_8799.n316 gnd 0.998708f
C6214 a_n8300_8799.t22 gnd 0.112772f
C6215 a_n8300_8799.t23 gnd 0.112772f
C6216 a_n8300_8799.n317 gnd 0.996492f
C6217 a_n8300_8799.n318 gnd 0.793752f
C6218 a_n8300_8799.t21 gnd 0.112772f
C6219 a_n8300_8799.t39 gnd 0.112772f
C6220 a_n8300_8799.n319 gnd 0.996492f
C6221 a_n8300_8799.n320 gnd 0.331444f
C6222 a_n8300_8799.n321 gnd 0.473195f
C6223 a_n8300_8799.t41 gnd 0.112772f
C6224 a_n8300_8799.t34 gnd 0.112772f
C6225 a_n8300_8799.n322 gnd 0.996492f
C6226 a_n8300_8799.n323 gnd 0.331444f
C6227 a_n8300_8799.t36 gnd 0.112772f
C6228 a_n8300_8799.t20 gnd 0.112772f
C6229 a_n8300_8799.n324 gnd 0.996492f
C6230 a_n8300_8799.n325 gnd 0.389772f
C6231 a_n8300_8799.t38 gnd 0.112772f
C6232 a_n8300_8799.t40 gnd 0.112772f
C6233 a_n8300_8799.n326 gnd 0.996492f
C6234 a_n8300_8799.n327 gnd 2.86956f
C6235 a_n8300_8799.t35 gnd 0.112772f
C6236 a_n8300_8799.t33 gnd 0.112772f
C6237 a_n8300_8799.n328 gnd 0.998708f
C6238 a_n8300_8799.t24 gnd 0.112772f
C6239 a_n8300_8799.t30 gnd 0.112772f
C6240 a_n8300_8799.n329 gnd 0.996491f
C6241 a_n8300_8799.n330 gnd 0.793754f
C6242 a_n8300_8799.t42 gnd 0.112772f
C6243 a_n8300_8799.t25 gnd 0.112772f
C6244 a_n8300_8799.n331 gnd 0.996491f
C6245 a_n8300_8799.n332 gnd 0.331445f
C6246 a_n8300_8799.n333 gnd 2.41514f
C6247 a_n8300_8799.n334 gnd 0.331447f
C6248 a_n8300_8799.n335 gnd 0.996489f
C6249 a_n8300_8799.t43 gnd 0.112772f
C6250 a_n3827_n3924.n0 gnd 1.99733f
C6251 a_n3827_n3924.n1 gnd 2.17486f
C6252 a_n3827_n3924.n2 gnd 1.44807f
C6253 a_n3827_n3924.n3 gnd 1.31657f
C6254 a_n3827_n3924.n4 gnd 1.81285f
C6255 a_n3827_n3924.n5 gnd 3.90473f
C6256 a_n3827_n3924.n6 gnd 1.77302f
C6257 a_n3827_n3924.n7 gnd 0.886511f
C6258 a_n3827_n3924.n8 gnd 2.49022f
C6259 a_n3827_n3924.n9 gnd 0.954549f
C6260 a_n3827_n3924.n10 gnd 1.2733f
C6261 a_n3827_n3924.n11 gnd 0.724031f
C6262 a_n3827_n3924.t12 gnd 0.097472f
C6263 a_n3827_n3924.t14 gnd 0.097472f
C6264 a_n3827_n3924.t5 gnd 0.097472f
C6265 a_n3827_n3924.n12 gnd 0.796069f
C6266 a_n3827_n3924.t57 gnd 1.26084f
C6267 a_n3827_n3924.t7 gnd 1.01304f
C6268 a_n3827_n3924.t15 gnd 1.26048f
C6269 a_n3827_n3924.t21 gnd 1.25868f
C6270 a_n3827_n3924.t20 gnd 1.25868f
C6271 a_n3827_n3924.t11 gnd 1.25868f
C6272 a_n3827_n3924.t1 gnd 1.25868f
C6273 a_n3827_n3924.t16 gnd 1.25868f
C6274 a_n3827_n3924.t53 gnd 1.25868f
C6275 a_n3827_n3924.t2 gnd 1.25868f
C6276 a_n3827_n3924.t3 gnd 1.25868f
C6277 a_n3827_n3924.n13 gnd 0.914318f
C6278 a_n3827_n3924.t24 gnd 1.01304f
C6279 a_n3827_n3924.t22 gnd 0.097472f
C6280 a_n3827_n3924.t34 gnd 0.097472f
C6281 a_n3827_n3924.n14 gnd 0.796068f
C6282 a_n3827_n3924.t38 gnd 0.097472f
C6283 a_n3827_n3924.t40 gnd 0.097472f
C6284 a_n3827_n3924.n15 gnd 0.796068f
C6285 a_n3827_n3924.t28 gnd 0.097472f
C6286 a_n3827_n3924.t27 gnd 0.097472f
C6287 a_n3827_n3924.n16 gnd 0.796068f
C6288 a_n3827_n3924.t25 gnd 0.097472f
C6289 a_n3827_n3924.t37 gnd 0.097472f
C6290 a_n3827_n3924.n17 gnd 0.796068f
C6291 a_n3827_n3924.t45 gnd 0.097472f
C6292 a_n3827_n3924.t35 gnd 0.097472f
C6293 a_n3827_n3924.n18 gnd 0.796068f
C6294 a_n3827_n3924.t36 gnd 1.01304f
C6295 a_n3827_n3924.t10 gnd 1.01304f
C6296 a_n3827_n3924.t4 gnd 0.097472f
C6297 a_n3827_n3924.t49 gnd 0.097472f
C6298 a_n3827_n3924.n19 gnd 0.796068f
C6299 a_n3827_n3924.t52 gnd 0.097472f
C6300 a_n3827_n3924.t13 gnd 0.097472f
C6301 a_n3827_n3924.n20 gnd 0.796068f
C6302 a_n3827_n3924.t48 gnd 0.097472f
C6303 a_n3827_n3924.t17 gnd 0.097472f
C6304 a_n3827_n3924.n21 gnd 0.796068f
C6305 a_n3827_n3924.t47 gnd 0.097472f
C6306 a_n3827_n3924.t50 gnd 0.097472f
C6307 a_n3827_n3924.n22 gnd 0.796068f
C6308 a_n3827_n3924.t8 gnd 0.097472f
C6309 a_n3827_n3924.t51 gnd 0.097472f
C6310 a_n3827_n3924.n23 gnd 0.796068f
C6311 a_n3827_n3924.t55 gnd 1.01304f
C6312 a_n3827_n3924.n24 gnd 0.914318f
C6313 a_n3827_n3924.t43 gnd 1.01304f
C6314 a_n3827_n3924.t30 gnd 0.097472f
C6315 a_n3827_n3924.t41 gnd 0.097472f
C6316 a_n3827_n3924.n25 gnd 0.796069f
C6317 a_n3827_n3924.t39 gnd 0.097472f
C6318 a_n3827_n3924.t44 gnd 0.097472f
C6319 a_n3827_n3924.n26 gnd 0.796069f
C6320 a_n3827_n3924.t42 gnd 0.097472f
C6321 a_n3827_n3924.t26 gnd 0.097472f
C6322 a_n3827_n3924.n27 gnd 0.796069f
C6323 a_n3827_n3924.t33 gnd 0.097472f
C6324 a_n3827_n3924.t29 gnd 0.097472f
C6325 a_n3827_n3924.n28 gnd 0.796069f
C6326 a_n3827_n3924.t31 gnd 0.097472f
C6327 a_n3827_n3924.t32 gnd 0.097472f
C6328 a_n3827_n3924.n29 gnd 0.796069f
C6329 a_n3827_n3924.t23 gnd 1.01304f
C6330 a_n3827_n3924.t46 gnd 1.01304f
C6331 a_n3827_n3924.t56 gnd 0.097472f
C6332 a_n3827_n3924.t19 gnd 0.097472f
C6333 a_n3827_n3924.n30 gnd 0.796069f
C6334 a_n3827_n3924.t9 gnd 0.097472f
C6335 a_n3827_n3924.t6 gnd 0.097472f
C6336 a_n3827_n3924.n31 gnd 0.796069f
C6337 a_n3827_n3924.t18 gnd 0.097472f
C6338 a_n3827_n3924.t54 gnd 0.097472f
C6339 a_n3827_n3924.n32 gnd 0.796069f
C6340 a_n3827_n3924.n33 gnd 0.79607f
C6341 a_n3827_n3924.t0 gnd 0.097472f
C6342 plus.n0 gnd 0.022995f
C6343 plus.t21 gnd 0.325242f
C6344 plus.n1 gnd 0.022995f
C6345 plus.t22 gnd 0.325242f
C6346 plus.t16 gnd 0.325242f
C6347 plus.n2 gnd 0.144483f
C6348 plus.n3 gnd 0.022995f
C6349 plus.t17 gnd 0.325242f
C6350 plus.t11 gnd 0.325242f
C6351 plus.n4 gnd 0.144483f
C6352 plus.n5 gnd 0.022995f
C6353 plus.t5 gnd 0.325242f
C6354 plus.t6 gnd 0.325242f
C6355 plus.n6 gnd 0.144483f
C6356 plus.n7 gnd 0.022995f
C6357 plus.t23 gnd 0.325242f
C6358 plus.t24 gnd 0.325242f
C6359 plus.n8 gnd 0.144483f
C6360 plus.n9 gnd 0.022995f
C6361 plus.t18 gnd 0.325242f
C6362 plus.t13 gnd 0.325242f
C6363 plus.n10 gnd 0.149189f
C6364 plus.t15 gnd 0.337048f
C6365 plus.n11 gnd 0.133901f
C6366 plus.n12 gnd 0.098995f
C6367 plus.n13 gnd 0.005218f
C6368 plus.n14 gnd 0.144483f
C6369 plus.n15 gnd 0.005218f
C6370 plus.n16 gnd 0.022995f
C6371 plus.n17 gnd 0.022995f
C6372 plus.n18 gnd 0.022995f
C6373 plus.n19 gnd 0.005218f
C6374 plus.n20 gnd 0.144483f
C6375 plus.n21 gnd 0.005218f
C6376 plus.n22 gnd 0.022995f
C6377 plus.n23 gnd 0.022995f
C6378 plus.n24 gnd 0.022995f
C6379 plus.n25 gnd 0.005218f
C6380 plus.n26 gnd 0.144483f
C6381 plus.n27 gnd 0.005218f
C6382 plus.n28 gnd 0.022995f
C6383 plus.n29 gnd 0.022995f
C6384 plus.n30 gnd 0.022995f
C6385 plus.n31 gnd 0.005218f
C6386 plus.n32 gnd 0.144483f
C6387 plus.n33 gnd 0.005218f
C6388 plus.n34 gnd 0.022995f
C6389 plus.n35 gnd 0.022995f
C6390 plus.n36 gnd 0.022995f
C6391 plus.n37 gnd 0.005218f
C6392 plus.n38 gnd 0.144483f
C6393 plus.n39 gnd 0.005218f
C6394 plus.n40 gnd 0.144695f
C6395 plus.n41 gnd 0.260382f
C6396 plus.n42 gnd 0.022995f
C6397 plus.n43 gnd 0.005218f
C6398 plus.t10 gnd 0.325242f
C6399 plus.n44 gnd 0.022995f
C6400 plus.n45 gnd 0.005218f
C6401 plus.t12 gnd 0.325242f
C6402 plus.n46 gnd 0.022995f
C6403 plus.n47 gnd 0.005218f
C6404 plus.t7 gnd 0.325242f
C6405 plus.n48 gnd 0.022995f
C6406 plus.n49 gnd 0.005218f
C6407 plus.t27 gnd 0.325242f
C6408 plus.n50 gnd 0.022995f
C6409 plus.n51 gnd 0.005218f
C6410 plus.t26 gnd 0.325242f
C6411 plus.t20 gnd 0.337048f
C6412 plus.t19 gnd 0.325242f
C6413 plus.n52 gnd 0.149189f
C6414 plus.n53 gnd 0.133901f
C6415 plus.n54 gnd 0.098994f
C6416 plus.n55 gnd 0.022995f
C6417 plus.n56 gnd 0.144483f
C6418 plus.n57 gnd 0.005218f
C6419 plus.t25 gnd 0.325242f
C6420 plus.n58 gnd 0.144483f
C6421 plus.n59 gnd 0.022995f
C6422 plus.n60 gnd 0.022995f
C6423 plus.n61 gnd 0.022995f
C6424 plus.n62 gnd 0.144483f
C6425 plus.n63 gnd 0.005218f
C6426 plus.t9 gnd 0.325242f
C6427 plus.n64 gnd 0.144483f
C6428 plus.n65 gnd 0.022995f
C6429 plus.n66 gnd 0.022995f
C6430 plus.n67 gnd 0.022995f
C6431 plus.n68 gnd 0.144483f
C6432 plus.n69 gnd 0.005218f
C6433 plus.t14 gnd 0.325242f
C6434 plus.n70 gnd 0.144483f
C6435 plus.n71 gnd 0.022995f
C6436 plus.n72 gnd 0.022995f
C6437 plus.n73 gnd 0.022995f
C6438 plus.n74 gnd 0.144483f
C6439 plus.n75 gnd 0.005218f
C6440 plus.t28 gnd 0.325242f
C6441 plus.n76 gnd 0.144483f
C6442 plus.n77 gnd 0.022995f
C6443 plus.n78 gnd 0.022995f
C6444 plus.n79 gnd 0.022995f
C6445 plus.n80 gnd 0.144483f
C6446 plus.n81 gnd 0.005218f
C6447 plus.t8 gnd 0.325242f
C6448 plus.n82 gnd 0.144695f
C6449 plus.n83 gnd 0.761135f
C6450 plus.n84 gnd 1.13871f
C6451 plus.t2 gnd 0.039696f
C6452 plus.t3 gnd 0.007089f
C6453 plus.t1 gnd 0.007089f
C6454 plus.n85 gnd 0.02299f
C6455 plus.n86 gnd 0.178472f
C6456 plus.t4 gnd 0.007089f
C6457 plus.t0 gnd 0.007089f
C6458 plus.n87 gnd 0.02299f
C6459 plus.n88 gnd 0.133965f
C6460 plus.n89 gnd 3.14792f
.ends

