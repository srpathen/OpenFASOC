* NGSPICE file created from opamp607.ext - technology: sky130A

.subckt opamp607 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 a_n9628_8799.t34 plus.t5 a_n3827_n3924.t38 gnd.t286 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X1 a_n2804_13878.t31 a_n2982_13878.t20 a_n2982_13878.t21 vdd.t290 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X2 a_n2804_13878.t0 a_n2982_13878.t64 vdd.t303 vdd.t302 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 vdd.t247 a_n9628_8799.t40 CSoutput.t168 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X4 outputibias.t7 outputibias.t6 gnd.t289 gnd.t288 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X5 CSoutput.t167 a_n9628_8799.t41 vdd.t246 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X6 a_n3827_n3924.t41 diffpairibias.t20 gnd.t355 gnd.t354 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X7 gnd.t126 commonsourceibias.t80 CSoutput.t41 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 gnd.t260 gnd.t258 gnd.t259 gnd.t230 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X9 commonsourceibias.t79 commonsourceibias.t78 gnd.t312 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X10 a_n3827_n3924.t36 plus.t6 a_n9628_8799.t33 gnd.t104 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X11 commonsourceibias.t77 commonsourceibias.t76 gnd.t7 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X12 plus.t0 gnd.t255 gnd.t257 gnd.t256 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X13 gnd.t254 gnd.t252 gnd.t253 gnd.t230 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X14 vdd.t245 a_n9628_8799.t42 CSoutput.t166 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X15 a_n2982_8322.t37 a_n2982_13878.t65 a_n9628_8799.t0 vdd.t300 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X16 vdd.t84 CSoutput.t200 output.t19 gnd.t39 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X17 gnd.t251 gnd.t249 gnd.t250 gnd.t169 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X18 CSoutput.t42 commonsourceibias.t81 gnd.t127 gnd.t74 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X19 CSoutput.t165 a_n9628_8799.t43 vdd.t244 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X20 vdd.t243 a_n9628_8799.t44 CSoutput.t164 vdd.t227 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X21 CSoutput.t163 a_n9628_8799.t45 vdd.t242 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X22 gnd.t38 commonsourceibias.t74 commonsourceibias.t75 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X23 CSoutput.t196 commonsourceibias.t82 gnd.t345 gnd.t277 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X24 vdd.t241 a_n9628_8799.t46 CSoutput.t162 vdd.t227 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X25 vdd.t240 a_n9628_8799.t47 CSoutput.t161 vdd.t169 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X26 gnd.t248 gnd.t246 gnd.t247 gnd.t169 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X27 CSoutput.t160 a_n9628_8799.t48 vdd.t239 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X28 commonsourceibias.t73 commonsourceibias.t72 gnd.t278 gnd.t277 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X29 vdd.t2 CSoutput.t201 output.t18 gnd.t10 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X30 a_n9628_8799.t16 a_n2982_13878.t66 a_n2982_8322.t36 vdd.t286 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X31 CSoutput.t197 commonsourceibias.t83 gnd.t346 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 vdd.t238 a_n9628_8799.t49 CSoutput.t159 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X33 a_n2982_13878.t3 minus.t5 a_n3827_n3924.t4 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X34 vdd.t237 a_n9628_8799.t50 CSoutput.t158 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X35 CSoutput.t157 a_n9628_8799.t51 vdd.t236 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X36 a_n9628_8799.t7 a_n2982_13878.t67 a_n2982_8322.t35 vdd.t249 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X37 gnd.t245 gnd.t242 gnd.t244 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X38 commonsourceibias.t71 commonsourceibias.t70 gnd.t23 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X39 a_n3827_n3924.t12 minus.t6 a_n2982_13878.t8 gnd.t106 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X40 gnd.t241 gnd.t239 minus.t4 gnd.t240 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X41 CSoutput.t156 a_n9628_8799.t52 vdd.t235 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X42 a_n3827_n3924.t7 diffpairibias.t21 gnd.t72 gnd.t71 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X43 CSoutput.t4 commonsourceibias.t84 gnd.t28 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X44 CSoutput.t155 a_n9628_8799.t53 vdd.t234 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X45 vdd.t233 a_n9628_8799.t54 CSoutput.t154 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X46 gnd.t30 commonsourceibias.t85 CSoutput.t5 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X47 gnd.t238 gnd.t236 gnd.t237 gnd.t204 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X48 vdd.t232 a_n9628_8799.t55 CSoutput.t153 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X49 gnd.t235 gnd.t233 gnd.t234 gnd.t157 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X50 gnd.t279 commonsourceibias.t68 commonsourceibias.t69 gnd.t119 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X51 vdd.t83 vdd.t81 vdd.t82 vdd.t72 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X52 commonsourceibias.t67 commonsourceibias.t66 gnd.t317 gnd.t124 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X53 a_n3827_n3924.t30 plus.t7 a_n9628_8799.t32 gnd.t283 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X54 vdd.t231 a_n9628_8799.t56 CSoutput.t152 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X55 gnd.t269 commonsourceibias.t86 CSoutput.t171 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X56 a_n2804_13878.t30 a_n2982_13878.t42 a_n2982_13878.t43 vdd.t257 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X57 gnd.t270 commonsourceibias.t87 CSoutput.t172 gnd.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X58 a_n2982_13878.t25 a_n2982_13878.t24 a_n2804_13878.t29 vdd.t272 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X59 vdd.t80 vdd.t78 vdd.t79 vdd.t72 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X60 gnd.t94 commonsourceibias.t88 CSoutput.t24 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X61 a_n9628_8799.t31 plus.t8 a_n3827_n3924.t34 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X62 CSoutput.t151 a_n9628_8799.t57 vdd.t230 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X63 vdd.t77 vdd.t75 vdd.t76 vdd.t54 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X64 output.t17 CSoutput.t202 vdd.t3 gnd.t11 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X65 vdd.t229 a_n9628_8799.t58 CSoutput.t150 vdd.t169 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X66 vdd.t228 a_n9628_8799.t59 CSoutput.t149 vdd.t227 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X67 gnd.t98 commonsourceibias.t64 commonsourceibias.t65 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X68 diffpairibias.t19 diffpairibias.t18 gnd.t310 gnd.t309 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X69 commonsourceibias.t63 commonsourceibias.t62 gnd.t271 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X70 CSoutput.t148 a_n9628_8799.t60 vdd.t226 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X71 a_n2982_13878.t15 minus.t7 a_n3827_n3924.t21 gnd.t311 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X72 a_n2982_13878.t55 a_n2982_13878.t54 a_n2804_13878.t28 vdd.t285 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X73 CSoutput.t147 a_n9628_8799.t61 vdd.t225 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X74 a_n9628_8799.t8 a_n2982_13878.t68 a_n2982_8322.t34 vdd.t282 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X75 vdd.t224 a_n9628_8799.t62 CSoutput.t146 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X76 CSoutput.t145 a_n9628_8799.t63 vdd.t223 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X77 commonsourceibias.t61 commonsourceibias.t60 gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X78 a_n2982_13878.t53 a_n2982_13878.t52 a_n2804_13878.t27 vdd.t301 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X79 vdd.t222 a_n9628_8799.t64 CSoutput.t144 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X80 vdd.t221 a_n9628_8799.t65 CSoutput.t143 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X81 a_n9628_8799.t2 a_n2982_13878.t69 a_n2982_8322.t33 vdd.t280 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X82 CSoutput.t142 a_n9628_8799.t66 vdd.t213 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X83 gnd.t232 gnd.t229 gnd.t231 gnd.t230 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X84 diffpairibias.t17 diffpairibias.t16 gnd.t285 gnd.t284 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X85 gnd.t347 commonsourceibias.t58 commonsourceibias.t59 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X86 CSoutput.t141 a_n9628_8799.t67 vdd.t220 vdd.t113 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X87 a_n9628_8799.t36 a_n2982_13878.t70 a_n2982_8322.t32 vdd.t293 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X88 CSoutput.t25 commonsourceibias.t89 gnd.t95 gnd.t74 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 a_n2982_8322.t31 a_n2982_13878.t71 a_n9628_8799.t9 vdd.t301 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X90 CSoutput.t39 commonsourceibias.t90 gnd.t123 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 CSoutput.t140 a_n9628_8799.t68 vdd.t219 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X92 gnd.t64 commonsourceibias.t56 commonsourceibias.t57 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X93 vdd.t4 CSoutput.t203 output.t16 gnd.t12 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X94 CSoutput.t40 commonsourceibias.t91 gnd.t125 gnd.t124 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X95 CSoutput.t175 commonsourceibias.t92 gnd.t275 gnd.t131 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X96 vdd.t74 vdd.t71 vdd.t73 vdd.t72 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X97 a_n3827_n3924.t33 plus.t9 a_n9628_8799.t30 gnd.t137 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X98 CSoutput.t176 commonsourceibias.t93 gnd.t276 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X99 gnd.t228 gnd.t226 minus.t3 gnd.t227 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X100 CSoutput.t173 commonsourceibias.t94 gnd.t272 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X101 a_n3827_n3924.t19 diffpairibias.t22 gnd.t305 gnd.t304 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X102 CSoutput.t139 a_n9628_8799.t69 vdd.t218 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X103 vdd.t216 a_n9628_8799.t70 CSoutput.t138 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X104 vdd.t215 a_n9628_8799.t71 CSoutput.t137 vdd.t205 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X105 a_n2982_13878.t57 a_n2982_13878.t56 a_n2804_13878.t26 vdd.t300 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X106 vdd.t214 a_n9628_8799.t72 CSoutput.t136 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X107 output.t15 CSoutput.t204 vdd.t5 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X108 a_n9628_8799.t13 a_n2982_13878.t72 a_n2982_8322.t30 vdd.t289 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X109 a_n2982_13878.t49 a_n2982_13878.t48 a_n2804_13878.t25 vdd.t252 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X110 gnd.t15 commonsourceibias.t54 commonsourceibias.t55 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X111 gnd.t41 commonsourceibias.t52 commonsourceibias.t53 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X112 gnd.t338 commonsourceibias.t50 commonsourceibias.t51 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X113 output.t3 outputibias.t8 gnd.t152 gnd.t151 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X114 CSoutput.t205 a_n2982_8322.t5 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X115 vdd.t212 a_n9628_8799.t73 CSoutput.t135 vdd.t175 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X116 CSoutput.t134 a_n9628_8799.t74 vdd.t211 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X117 gnd.t225 gnd.t222 gnd.t224 gnd.t223 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X118 CSoutput.t133 a_n9628_8799.t75 vdd.t210 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X119 diffpairibias.t15 diffpairibias.t14 gnd.t150 gnd.t149 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X120 a_n2982_13878.t1 minus.t8 a_n3827_n3924.t2 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X121 output.t2 outputibias.t9 gnd.t262 gnd.t261 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X122 vdd.t70 vdd.t68 vdd.t69 vdd.t61 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X123 CSoutput.t132 a_n9628_8799.t76 vdd.t209 vdd.t113 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X124 gnd.t274 commonsourceibias.t95 CSoutput.t174 gnd.t273 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X125 vdd.t67 vdd.t64 vdd.t66 vdd.t65 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X126 gnd.t120 commonsourceibias.t96 CSoutput.t37 gnd.t119 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X127 gnd.t122 commonsourceibias.t97 CSoutput.t38 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X128 gnd.t218 gnd.t216 gnd.t217 gnd.t161 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X129 gnd.t116 commonsourceibias.t98 CSoutput.t35 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X130 a_n2804_13878.t24 a_n2982_13878.t36 a_n2982_13878.t37 vdd.t262 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X131 a_n3827_n3924.t3 minus.t9 a_n2982_13878.t2 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X132 CSoutput.t131 a_n9628_8799.t77 vdd.t208 vdd.t88 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X133 gnd.t118 commonsourceibias.t99 CSoutput.t36 gnd.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X134 output.t14 CSoutput.t206 vdd.t0 gnd.t8 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X135 vdd.t207 a_n9628_8799.t78 CSoutput.t130 vdd.t205 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X136 vdd.t1 CSoutput.t207 output.t13 gnd.t9 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X137 vdd.t299 a_n2982_13878.t73 a_n2982_8322.t13 vdd.t298 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X138 a_n2982_13878.t35 a_n2982_13878.t34 a_n2804_13878.t23 vdd.t260 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X139 gnd.t113 commonsourceibias.t100 CSoutput.t33 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X140 gnd.t221 gnd.t219 gnd.t220 gnd.t176 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X141 a_n2982_8322.t12 a_n2982_13878.t74 vdd.t297 vdd.t296 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X142 a_n3827_n3924.t5 diffpairibias.t23 gnd.t69 gnd.t68 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X143 CSoutput.t129 a_n9628_8799.t79 vdd.t203 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X144 CSoutput.t34 commonsourceibias.t101 gnd.t115 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X145 a_n3827_n3924.t20 minus.t10 a_n2982_13878.t14 gnd.t308 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X146 gnd.t301 commonsourceibias.t48 commonsourceibias.t49 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X147 gnd.t215 gnd.t213 plus.t2 gnd.t214 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X148 vdd.t295 a_n2982_13878.t75 a_n2804_13878.t4 vdd.t294 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X149 a_n3827_n3924.t29 plus.t10 a_n9628_8799.t29 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X150 gnd.t111 commonsourceibias.t102 CSoutput.t31 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X151 vdd.t63 vdd.t60 vdd.t62 vdd.t61 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X152 a_n2804_13878.t22 a_n2982_13878.t38 a_n2982_13878.t39 vdd.t293 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X153 vdd.t206 a_n9628_8799.t80 CSoutput.t128 vdd.t205 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X154 vdd.t204 a_n9628_8799.t81 CSoutput.t127 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X155 a_n2982_8322.t29 a_n2982_13878.t76 a_n9628_8799.t12 vdd.t281 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X156 gnd.t280 commonsourceibias.t46 commonsourceibias.t47 gnd.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X157 a_n9628_8799.t28 plus.t11 a_n3827_n3924.t27 gnd.t282 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X158 a_n9628_8799.t27 plus.t12 a_n3827_n3924.t26 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X159 vdd.t59 vdd.t57 vdd.t58 vdd.t34 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X160 vdd.t56 vdd.t53 vdd.t55 vdd.t54 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X161 a_n2982_8322.t11 a_n2982_13878.t77 vdd.t292 vdd.t291 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X162 a_n9628_8799.t17 a_n2982_13878.t78 a_n2982_8322.t28 vdd.t259 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X163 CSoutput.t126 a_n9628_8799.t82 vdd.t202 vdd.t125 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X164 diffpairibias.t13 diffpairibias.t12 gnd.t264 gnd.t263 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X165 CSoutput.t208 a_n2982_8322.t4 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X166 vdd.t201 a_n9628_8799.t83 CSoutput.t125 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X167 CSoutput.t32 commonsourceibias.t103 gnd.t112 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X168 a_n2982_13878.t13 minus.t11 a_n3827_n3924.t18 gnd.t287 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X169 a_n2982_13878.t31 a_n2982_13878.t30 a_n2804_13878.t21 vdd.t275 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X170 a_n9628_8799.t3 a_n2982_13878.t79 a_n2982_8322.t27 vdd.t290 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X171 CSoutput.t124 a_n9628_8799.t84 vdd.t199 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X172 CSoutput.t123 a_n9628_8799.t85 vdd.t197 vdd.t162 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X173 CSoutput.t192 commonsourceibias.t104 gnd.t336 gnd.t124 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X174 a_n2804_13878.t20 a_n2982_13878.t40 a_n2982_13878.t41 vdd.t289 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X175 commonsourceibias.t45 commonsourceibias.t44 gnd.t75 gnd.t74 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X176 CSoutput.t193 commonsourceibias.t105 gnd.t337 gnd.t131 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X177 gnd.t334 commonsourceibias.t106 CSoutput.t190 gnd.t50 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X178 a_n3827_n3924.t0 minus.t12 a_n2982_13878.t0 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X179 CSoutput.t191 commonsourceibias.t107 gnd.t335 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X180 vdd.t6 CSoutput.t209 output.t12 gnd.t20 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X181 minus.t2 gnd.t210 gnd.t212 gnd.t211 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X182 CSoutput.t188 commonsourceibias.t108 gnd.t332 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X183 vdd.t52 vdd.t50 vdd.t51 vdd.t13 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X184 CSoutput.t122 a_n9628_8799.t86 vdd.t196 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X185 gnd.t333 commonsourceibias.t109 CSoutput.t189 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X186 gnd.t302 commonsourceibias.t42 commonsourceibias.t43 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X187 vdd.t288 a_n2982_13878.t80 a_n2982_8322.t10 vdd.t287 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X188 a_n2804_13878.t19 a_n2982_13878.t62 a_n2982_13878.t63 vdd.t286 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X189 vdd.t195 a_n9628_8799.t87 CSoutput.t121 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X190 gnd.t324 commonsourceibias.t110 CSoutput.t180 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X191 vdd.t194 a_n9628_8799.t88 CSoutput.t120 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X192 a_n2982_13878.t33 a_n2982_13878.t32 a_n2804_13878.t18 vdd.t256 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X193 commonsourceibias.t41 commonsourceibias.t40 gnd.t281 gnd.t139 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X194 gnd.t76 commonsourceibias.t38 commonsourceibias.t39 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X195 vdd.t193 a_n9628_8799.t89 CSoutput.t119 vdd.t175 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X196 vdd.t187 a_n9628_8799.t90 CSoutput.t118 vdd.t127 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X197 gnd.t303 commonsourceibias.t36 commonsourceibias.t37 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X198 CSoutput.t117 a_n9628_8799.t91 vdd.t192 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X199 a_n3827_n3924.t13 diffpairibias.t24 gnd.t136 gnd.t135 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X200 commonsourceibias.t35 commonsourceibias.t34 gnd.t78 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X201 vdd.t49 vdd.t47 vdd.t48 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X202 a_n3827_n3924.t23 diffpairibias.t25 gnd.t321 gnd.t320 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X203 gnd.t325 commonsourceibias.t111 CSoutput.t181 gnd.t147 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X204 vdd.t191 a_n9628_8799.t92 CSoutput.t116 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X205 vdd.t190 a_n9628_8799.t93 CSoutput.t115 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X206 gnd.t330 commonsourceibias.t112 CSoutput.t186 gnd.t273 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 CSoutput.t114 a_n9628_8799.t94 vdd.t189 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X208 gnd.t331 commonsourceibias.t113 CSoutput.t187 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X209 gnd.t328 commonsourceibias.t114 CSoutput.t184 gnd.t119 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X210 vdd.t46 vdd.t44 vdd.t45 vdd.t34 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X211 gnd.t329 commonsourceibias.t115 CSoutput.t185 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X212 a_n2804_13878.t17 a_n2982_13878.t44 a_n2982_13878.t45 vdd.t261 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X213 CSoutput.t210 a_n2982_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X214 CSoutput.t45 commonsourceibias.t116 gnd.t144 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X215 a_n2982_8322.t26 a_n2982_13878.t81 a_n9628_8799.t4 vdd.t285 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X216 CSoutput.t113 a_n9628_8799.t95 vdd.t188 vdd.t162 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X217 CSoutput.t112 a_n9628_8799.t96 vdd.t186 vdd.t92 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X218 commonsourceibias.t33 commonsourceibias.t32 gnd.t53 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X219 CSoutput.t46 commonsourceibias.t117 gnd.t145 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X220 CSoutput.t211 a_n2982_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X221 gnd.t326 commonsourceibias.t118 CSoutput.t182 gnd.t89 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X222 CSoutput.t183 commonsourceibias.t119 gnd.t327 gnd.t291 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X223 gnd.t209 gnd.t207 gnd.t208 gnd.t157 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X224 diffpairibias.t11 diffpairibias.t10 gnd.t102 gnd.t101 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X225 a_n2804_13878.t3 a_n2982_13878.t82 vdd.t284 vdd.t283 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X226 gnd.t61 commonsourceibias.t120 CSoutput.t17 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X227 vdd.t271 a_n2982_13878.t83 a_n2804_13878.t1 vdd.t270 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X228 output.t1 outputibias.t10 gnd.t266 gnd.t265 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X229 gnd.t290 commonsourceibias.t30 commonsourceibias.t31 gnd.t147 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X230 CSoutput.t111 a_n9628_8799.t97 vdd.t185 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X231 gnd.t85 commonsourceibias.t28 commonsourceibias.t29 gnd.t50 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X232 vdd.t183 a_n9628_8799.t98 CSoutput.t110 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X233 vdd.t181 a_n9628_8799.t99 CSoutput.t109 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X234 commonsourceibias.t27 commonsourceibias.t26 gnd.t128 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 gnd.t206 gnd.t203 gnd.t205 gnd.t204 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X236 gnd.t202 gnd.t200 plus.t1 gnd.t201 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X237 vdd.t179 a_n9628_8799.t100 CSoutput.t108 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X238 CSoutput.t18 commonsourceibias.t121 gnd.t62 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X239 CSoutput.t107 a_n9628_8799.t101 vdd.t177 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X240 a_n2804_13878.t16 a_n2982_13878.t58 a_n2982_13878.t59 vdd.t282 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X241 diffpairibias.t9 diffpairibias.t8 gnd.t36 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X242 a_n3827_n3924.t16 minus.t13 a_n2982_13878.t11 gnd.t283 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X243 vdd.t176 a_n9628_8799.t102 CSoutput.t106 vdd.t175 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X244 vdd.t174 a_n9628_8799.t103 CSoutput.t105 vdd.t127 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X245 gnd.t87 commonsourceibias.t24 commonsourceibias.t25 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X246 CSoutput.t11 commonsourceibias.t122 gnd.t49 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X247 CSoutput.t104 a_n9628_8799.t104 vdd.t173 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X248 a_n2982_8322.t25 a_n2982_13878.t84 a_n9628_8799.t6 vdd.t248 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X249 a_n2982_13878.t19 a_n2982_13878.t18 a_n2804_13878.t15 vdd.t281 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X250 CSoutput.t103 a_n9628_8799.t105 vdd.t171 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X251 diffpairibias.t7 diffpairibias.t6 gnd.t142 gnd.t141 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X252 vdd.t170 a_n9628_8799.t106 CSoutput.t102 vdd.t169 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X253 a_n2804_13878.t14 a_n2982_13878.t22 a_n2982_13878.t23 vdd.t280 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X254 a_n2982_13878.t5 minus.t14 a_n3827_n3924.t8 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X255 a_n2982_13878.t12 minus.t15 a_n3827_n3924.t17 gnd.t286 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X256 gnd.t51 commonsourceibias.t123 CSoutput.t12 gnd.t50 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X257 vdd.t279 a_n2982_13878.t85 a_n2982_8322.t9 vdd.t278 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X258 vdd.t168 a_n9628_8799.t107 CSoutput.t101 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X259 vdd.t7 CSoutput.t212 output.t11 gnd.t21 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X260 CSoutput.t15 commonsourceibias.t124 gnd.t57 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X261 a_n9628_8799.t26 plus.t13 a_n3827_n3924.t28 gnd.t311 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X262 CSoutput.t16 commonsourceibias.t125 gnd.t59 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X263 gnd.t199 gnd.t196 gnd.t198 gnd.t197 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X264 gnd.t48 commonsourceibias.t126 CSoutput.t10 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X265 a_n3827_n3924.t10 minus.t16 a_n2982_13878.t6 gnd.t104 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X266 CSoutput.t100 a_n9628_8799.t108 vdd.t166 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X267 gnd.t195 gnd.t192 gnd.t194 gnd.t193 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X268 gnd.t56 commonsourceibias.t127 CSoutput.t14 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X269 a_n2804_13878.t5 a_n2982_13878.t86 vdd.t277 vdd.t276 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X270 CSoutput.t9 commonsourceibias.t128 gnd.t46 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X271 commonsourceibias.t23 commonsourceibias.t22 gnd.t130 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X272 vdd.t165 a_n9628_8799.t109 CSoutput.t99 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 CSoutput.t47 commonsourceibias.t129 gnd.t146 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X274 CSoutput.t98 a_n9628_8799.t110 vdd.t163 vdd.t162 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X275 CSoutput.t97 a_n9628_8799.t111 vdd.t161 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X276 gnd.t191 gnd.t189 gnd.t190 gnd.t176 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X277 vdd.t43 vdd.t41 vdd.t42 vdd.t17 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X278 vdd.t160 a_n9628_8799.t112 CSoutput.t96 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X279 a_n3827_n3924.t22 diffpairibias.t26 gnd.t319 gnd.t318 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X280 a_n2982_8322.t24 a_n2982_13878.t87 a_n9628_8799.t35 vdd.t275 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X281 vdd.t274 a_n2982_13878.t88 a_n2982_8322.t8 vdd.t273 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X282 gnd.t148 commonsourceibias.t130 CSoutput.t48 gnd.t147 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X283 vdd.t159 a_n9628_8799.t113 CSoutput.t95 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X284 a_n9628_8799.t25 plus.t14 a_n3827_n3924.t39 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X285 gnd.t138 commonsourceibias.t131 CSoutput.t43 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X286 gnd.t188 gnd.t186 plus.t3 gnd.t187 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X287 CSoutput.t179 commonsourceibias.t132 gnd.t300 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X288 vdd.t40 vdd.t37 vdd.t39 vdd.t38 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X289 CSoutput.t178 commonsourceibias.t133 gnd.t299 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X290 vdd.t158 a_n9628_8799.t114 CSoutput.t94 vdd.t120 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X291 a_n3827_n3924.t37 plus.t15 a_n9628_8799.t24 gnd.t106 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X292 vdd.t157 a_n9628_8799.t115 CSoutput.t93 vdd.t90 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X293 vdd.t156 a_n9628_8799.t116 CSoutput.t92 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X294 CSoutput.t91 a_n9628_8799.t117 vdd.t155 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X295 CSoutput.t90 a_n9628_8799.t118 vdd.t153 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X296 CSoutput.t89 a_n9628_8799.t119 vdd.t151 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X297 gnd.t298 commonsourceibias.t134 CSoutput.t177 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X298 gnd.t344 commonsourceibias.t135 CSoutput.t195 gnd.t89 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X299 a_n2804_13878.t13 a_n2982_13878.t28 a_n2982_13878.t29 vdd.t265 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X300 CSoutput.t88 a_n9628_8799.t120 vdd.t150 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X301 vdd.t85 CSoutput.t213 output.t10 gnd.t96 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X302 CSoutput.t199 commonsourceibias.t136 gnd.t351 gnd.t291 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X303 a_n2982_8322.t23 a_n2982_13878.t89 a_n9628_8799.t14 vdd.t272 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X304 diffpairibias.t5 diffpairibias.t4 gnd.t297 gnd.t296 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X305 commonsourceibias.t21 commonsourceibias.t20 gnd.t292 gnd.t291 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X306 gnd.t185 gnd.t182 gnd.t184 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X307 gnd.t268 commonsourceibias.t137 CSoutput.t170 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X308 CSoutput.t44 commonsourceibias.t138 gnd.t140 gnd.t139 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X309 gnd.t293 commonsourceibias.t18 commonsourceibias.t19 gnd.t273 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X310 CSoutput.t87 a_n9628_8799.t121 vdd.t149 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X311 CSoutput.t86 a_n9628_8799.t122 vdd.t147 vdd.t125 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X312 a_n3827_n3924.t9 diffpairibias.t27 gnd.t93 gnd.t92 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X313 vdd.t36 vdd.t33 vdd.t35 vdd.t34 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X314 CSoutput.t30 commonsourceibias.t139 gnd.t110 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X315 vdd.t146 a_n9628_8799.t123 CSoutput.t85 vdd.t120 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X316 CSoutput.t214 a_n2982_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X317 a_n2982_8322.t7 a_n2982_13878.t90 vdd.t269 vdd.t268 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X318 CSoutput.t84 a_n9628_8799.t124 vdd.t145 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X319 gnd.t163 gnd.t160 gnd.t162 gnd.t161 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X320 CSoutput.t8 commonsourceibias.t140 gnd.t45 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X321 vdd.t143 a_n9628_8799.t125 CSoutput.t83 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X322 CSoutput.t82 a_n9628_8799.t126 vdd.t142 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X323 vdd.t267 a_n2982_13878.t91 a_n2804_13878.t7 vdd.t266 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X324 gnd.t88 commonsourceibias.t16 commonsourceibias.t17 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X325 output.t0 outputibias.t11 gnd.t307 gnd.t306 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X326 vdd.t137 a_n9628_8799.t127 CSoutput.t81 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X327 CSoutput.t80 a_n9628_8799.t128 vdd.t141 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X328 CSoutput.t29 commonsourceibias.t141 gnd.t109 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X329 gnd.t84 commonsourceibias.t142 CSoutput.t23 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X330 vdd.t139 a_n9628_8799.t129 CSoutput.t79 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X331 CSoutput.t2 commonsourceibias.t143 gnd.t19 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X332 commonsourceibias.t15 commonsourceibias.t14 gnd.t54 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X333 a_n2982_8322.t22 a_n2982_13878.t92 a_n9628_8799.t37 vdd.t258 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X334 commonsourceibias.t13 commonsourceibias.t12 gnd.t294 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X335 gnd.t181 gnd.t179 minus.t1 gnd.t180 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X336 a_n9628_8799.t10 a_n2982_13878.t93 a_n2982_8322.t21 vdd.t265 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X337 CSoutput.t7 commonsourceibias.t144 gnd.t43 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X338 gnd.t90 commonsourceibias.t10 commonsourceibias.t11 gnd.t89 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X339 output.t9 CSoutput.t215 vdd.t86 gnd.t97 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X340 a_n2804_13878.t6 a_n2982_13878.t94 vdd.t264 vdd.t263 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X341 gnd.t82 commonsourceibias.t145 CSoutput.t22 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X342 CSoutput.t3 commonsourceibias.t146 gnd.t26 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X343 vdd.t135 a_n9628_8799.t130 CSoutput.t78 vdd.t90 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X344 vdd.t32 vdd.t30 vdd.t31 vdd.t9 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X345 vdd.t29 vdd.t27 vdd.t28 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X346 vdd.t134 a_n9628_8799.t131 CSoutput.t77 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X347 a_n2982_13878.t10 minus.t17 a_n3827_n3924.t15 gnd.t282 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X348 CSoutput.t76 a_n9628_8799.t132 vdd.t133 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X349 CSoutput.t75 a_n9628_8799.t133 vdd.t131 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X350 CSoutput.t74 a_n9628_8799.t134 vdd.t129 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X351 a_n2982_13878.t51 a_n2982_13878.t50 a_n2804_13878.t12 vdd.t253 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X352 gnd.t178 gnd.t175 gnd.t177 gnd.t176 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X353 a_n9628_8799.t11 a_n2982_13878.t95 a_n2982_8322.t20 vdd.t262 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X354 minus.t0 gnd.t172 gnd.t174 gnd.t173 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X355 a_n9628_8799.t1 a_n2982_13878.t96 a_n2982_8322.t19 vdd.t261 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X356 commonsourceibias.t9 commonsourceibias.t8 gnd.t132 gnd.t131 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X357 a_n2982_8322.t18 a_n2982_13878.t97 a_n9628_8799.t18 vdd.t260 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X358 a_n9628_8799.t23 plus.t16 a_n3827_n3924.t25 gnd.t287 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X359 a_n3827_n3924.t14 minus.t18 a_n2982_13878.t9 gnd.t137 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X360 vdd.t128 a_n9628_8799.t135 CSoutput.t73 vdd.t127 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X361 CSoutput.t72 a_n9628_8799.t136 vdd.t126 vdd.t125 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X362 CSoutput.t71 a_n9628_8799.t137 vdd.t124 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X363 CSoutput.t70 a_n9628_8799.t138 vdd.t123 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X364 gnd.t295 commonsourceibias.t6 commonsourceibias.t7 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X365 CSoutput.t69 a_n9628_8799.t139 vdd.t122 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X366 a_n2804_13878.t11 a_n2982_13878.t16 a_n2982_13878.t17 vdd.t259 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X367 vdd.t121 a_n9628_8799.t140 CSoutput.t68 vdd.t120 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X368 vdd.t119 a_n9628_8799.t141 CSoutput.t67 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X369 commonsourceibias.t5 commonsourceibias.t4 gnd.t133 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X370 vdd.t118 a_n9628_8799.t142 CSoutput.t66 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X371 a_n3827_n3924.t35 plus.t17 a_n9628_8799.t22 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X372 gnd.t55 commonsourceibias.t147 CSoutput.t13 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X373 CSoutput.t6 commonsourceibias.t148 gnd.t42 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X374 CSoutput.t216 a_n2982_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X375 output.t8 CSoutput.t217 vdd.t304 gnd.t313 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X376 gnd.t17 commonsourceibias.t149 CSoutput.t1 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X377 a_n3827_n3924.t40 diffpairibias.t28 gnd.t340 gnd.t339 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X378 vdd.t117 a_n9628_8799.t143 CSoutput.t65 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X379 gnd.t67 commonsourceibias.t150 CSoutput.t19 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X380 CSoutput.t64 a_n9628_8799.t144 vdd.t116 vdd.t92 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X381 a_n2982_13878.t47 a_n2982_13878.t46 a_n2804_13878.t10 vdd.t258 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X382 gnd.t171 gnd.t168 gnd.t170 gnd.t169 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X383 a_n9628_8799.t5 a_n2982_13878.t98 a_n2982_8322.t17 vdd.t257 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X384 vdd.t115 a_n9628_8799.t145 CSoutput.t63 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X385 output.t7 CSoutput.t218 vdd.t305 gnd.t314 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X386 gnd.t5 commonsourceibias.t151 CSoutput.t0 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X387 CSoutput.t62 a_n9628_8799.t146 vdd.t114 vdd.t113 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X388 vdd.t26 vdd.t24 vdd.t25 vdd.t17 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X389 a_n9628_8799.t21 plus.t18 a_n3827_n3924.t24 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X390 vdd.t306 CSoutput.t219 output.t6 gnd.t315 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X391 gnd.t167 gnd.t164 gnd.t166 gnd.t165 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X392 CSoutput.t194 commonsourceibias.t152 gnd.t343 gnd.t277 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X393 CSoutput.t198 commonsourceibias.t153 gnd.t350 gnd.t139 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X394 commonsourceibias.t3 commonsourceibias.t2 gnd.t34 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X395 outputibias.t5 outputibias.t4 gnd.t353 gnd.t352 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X396 diffpairibias.t3 diffpairibias.t2 gnd.t323 gnd.t322 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X397 CSoutput.t61 a_n9628_8799.t147 vdd.t112 vdd.t88 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X398 a_n2982_8322.t16 a_n2982_13878.t99 a_n9628_8799.t38 vdd.t256 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X399 a_n3827_n3924.t31 plus.t19 a_n9628_8799.t20 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X400 vdd.t111 a_n9628_8799.t148 CSoutput.t60 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X401 vdd.t23 vdd.t20 vdd.t22 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X402 CSoutput.t59 a_n9628_8799.t149 vdd.t109 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X403 outputibias.t3 outputibias.t2 gnd.t349 gnd.t348 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X404 CSoutput.t58 a_n9628_8799.t150 vdd.t107 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X405 diffpairibias.t1 diffpairibias.t0 gnd.t342 gnd.t341 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X406 a_n3827_n3924.t32 plus.t20 a_n9628_8799.t19 gnd.t308 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X407 CSoutput.t169 commonsourceibias.t154 gnd.t267 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X408 outputibias.t1 outputibias.t0 gnd.t100 gnd.t99 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X409 vdd.t255 a_n2982_13878.t100 a_n2804_13878.t2 vdd.t254 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X410 gnd.t108 commonsourceibias.t155 CSoutput.t28 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X411 CSoutput.t57 a_n9628_8799.t151 vdd.t103 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X412 CSoutput.t56 a_n9628_8799.t152 vdd.t105 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X413 a_n3827_n3924.t6 minus.t19 a_n2982_13878.t4 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X414 vdd.t101 a_n9628_8799.t153 CSoutput.t55 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X415 vdd.t99 a_n9628_8799.t154 CSoutput.t54 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X416 CSoutput.t27 commonsourceibias.t156 gnd.t107 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X417 output.t5 CSoutput.t220 vdd.t307 gnd.t316 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X418 gnd.t80 commonsourceibias.t157 CSoutput.t21 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X419 gnd.t159 gnd.t156 gnd.t158 gnd.t157 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X420 a_n2982_8322.t15 a_n2982_13878.t101 a_n9628_8799.t39 vdd.t253 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X421 a_n2982_13878.t7 minus.t20 a_n3827_n3924.t11 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X422 gnd.t103 commonsourceibias.t158 CSoutput.t26 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X423 a_n2982_8322.t14 a_n2982_13878.t102 a_n9628_8799.t15 vdd.t252 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X424 vdd.t97 a_n9628_8799.t155 CSoutput.t53 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X425 vdd.t95 a_n9628_8799.t156 CSoutput.t52 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X426 CSoutput.t51 a_n9628_8799.t157 vdd.t93 vdd.t92 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X427 output.t4 CSoutput.t221 vdd.t87 gnd.t134 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X428 plus.t4 gnd.t153 gnd.t155 gnd.t154 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X429 gnd.t79 commonsourceibias.t159 CSoutput.t20 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X430 vdd.t19 vdd.t16 vdd.t18 vdd.t17 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X431 a_n2982_8322.t6 a_n2982_13878.t103 vdd.t251 vdd.t250 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X432 a_n2804_13878.t9 a_n2982_13878.t26 a_n2982_13878.t27 vdd.t249 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X433 vdd.t15 vdd.t12 vdd.t14 vdd.t13 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X434 commonsourceibias.t1 commonsourceibias.t0 gnd.t91 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X435 a_n3827_n3924.t1 diffpairibias.t29 gnd.t2 gnd.t1 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X436 vdd.t11 vdd.t8 vdd.t10 vdd.t9 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X437 vdd.t91 a_n9628_8799.t158 CSoutput.t50 vdd.t90 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X438 CSoutput.t49 a_n9628_8799.t159 vdd.t89 vdd.t88 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X439 a_n2982_13878.t61 a_n2982_13878.t60 a_n2804_13878.t8 vdd.t248 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 plus.n33 plus.t15 321.495
R1 plus.n7 plus.t12 321.495
R2 plus.n32 plus.t14 297.12
R3 plus.n36 plus.t19 297.12
R4 plus.n38 plus.t18 297.12
R5 plus.n42 plus.t20 297.12
R6 plus.n44 plus.t8 297.12
R7 plus.n48 plus.t7 297.12
R8 plus.n50 plus.t11 297.12
R9 plus.n24 plus.t9 297.12
R10 plus.n22 plus.t5 297.12
R11 plus.n2 plus.t6 297.12
R12 plus.n16 plus.t16 297.12
R13 plus.n4 plus.t17 297.12
R14 plus.n10 plus.t13 297.12
R15 plus.n6 plus.t10 297.12
R16 plus.n54 plus.t2 243.97
R17 plus.n54 plus.n53 223.454
R18 plus.n56 plus.n55 223.454
R19 plus.n51 plus.n50 161.3
R20 plus.n49 plus.n26 161.3
R21 plus.n48 plus.n47 161.3
R22 plus.n46 plus.n27 161.3
R23 plus.n45 plus.n44 161.3
R24 plus.n43 plus.n28 161.3
R25 plus.n42 plus.n41 161.3
R26 plus.n40 plus.n29 161.3
R27 plus.n39 plus.n38 161.3
R28 plus.n37 plus.n30 161.3
R29 plus.n36 plus.n35 161.3
R30 plus.n34 plus.n31 161.3
R31 plus.n9 plus.n8 161.3
R32 plus.n10 plus.n5 161.3
R33 plus.n12 plus.n11 161.3
R34 plus.n13 plus.n4 161.3
R35 plus.n15 plus.n14 161.3
R36 plus.n16 plus.n3 161.3
R37 plus.n18 plus.n17 161.3
R38 plus.n19 plus.n2 161.3
R39 plus.n21 plus.n20 161.3
R40 plus.n22 plus.n1 161.3
R41 plus.n23 plus.n0 161.3
R42 plus.n25 plus.n24 161.3
R43 plus.n34 plus.n33 44.9377
R44 plus.n8 plus.n7 44.9377
R45 plus.n50 plus.n49 37.246
R46 plus.n24 plus.n23 37.246
R47 plus.n32 plus.n31 32.8641
R48 plus.n48 plus.n27 32.8641
R49 plus.n22 plus.n21 32.8641
R50 plus.n9 plus.n6 32.8641
R51 plus.n52 plus.n51 30.0327
R52 plus.n37 plus.n36 28.4823
R53 plus.n44 plus.n43 28.4823
R54 plus.n17 plus.n2 28.4823
R55 plus.n11 plus.n10 28.4823
R56 plus.n38 plus.n29 24.1005
R57 plus.n42 plus.n29 24.1005
R58 plus.n16 plus.n15 24.1005
R59 plus.n15 plus.n4 24.1005
R60 plus.n53 plus.t1 19.8005
R61 plus.n53 plus.t0 19.8005
R62 plus.n55 plus.t3 19.8005
R63 plus.n55 plus.t4 19.8005
R64 plus.n38 plus.n37 19.7187
R65 plus.n43 plus.n42 19.7187
R66 plus.n17 plus.n16 19.7187
R67 plus.n11 plus.n4 19.7187
R68 plus.n33 plus.n32 17.0522
R69 plus.n7 plus.n6 17.0522
R70 plus.n36 plus.n31 15.3369
R71 plus.n44 plus.n27 15.3369
R72 plus.n21 plus.n2 15.3369
R73 plus.n10 plus.n9 15.3369
R74 plus plus.n57 14.9378
R75 plus.n52 plus.n25 11.8547
R76 plus.n49 plus.n48 10.955
R77 plus.n23 plus.n22 10.955
R78 plus.n57 plus.n56 5.40567
R79 plus.n57 plus.n52 1.188
R80 plus.n56 plus.n54 0.716017
R81 plus.n35 plus.n34 0.189894
R82 plus.n35 plus.n30 0.189894
R83 plus.n39 plus.n30 0.189894
R84 plus.n40 plus.n39 0.189894
R85 plus.n41 plus.n40 0.189894
R86 plus.n41 plus.n28 0.189894
R87 plus.n45 plus.n28 0.189894
R88 plus.n46 plus.n45 0.189894
R89 plus.n47 plus.n46 0.189894
R90 plus.n47 plus.n26 0.189894
R91 plus.n51 plus.n26 0.189894
R92 plus.n25 plus.n0 0.189894
R93 plus.n1 plus.n0 0.189894
R94 plus.n20 plus.n1 0.189894
R95 plus.n20 plus.n19 0.189894
R96 plus.n19 plus.n18 0.189894
R97 plus.n18 plus.n3 0.189894
R98 plus.n14 plus.n3 0.189894
R99 plus.n14 plus.n13 0.189894
R100 plus.n13 plus.n12 0.189894
R101 plus.n12 plus.n5 0.189894
R102 plus.n8 plus.n5 0.189894
R103 a_n3827_n3924.n7 a_n3827_n3924.t9 214.994
R104 a_n3827_n3924.n8 a_n3827_n3924.t41 214.994
R105 a_n3827_n3924.n7 a_n3827_n3924.t5 214.321
R106 a_n3827_n3924.n7 a_n3827_n3924.t40 214.321
R107 a_n3827_n3924.n5 a_n3827_n3924.t23 214.321
R108 a_n3827_n3924.n5 a_n3827_n3924.t1 214.321
R109 a_n3827_n3924.n6 a_n3827_n3924.t13 214.321
R110 a_n3827_n3924.n6 a_n3827_n3924.t7 214.321
R111 a_n3827_n3924.n6 a_n3827_n3924.t19 214.321
R112 a_n3827_n3924.n8 a_n3827_n3924.t22 214.321
R113 a_n3827_n3924.n4 a_n3827_n3924.t37 55.8337
R114 a_n3827_n3924.n4 a_n3827_n3924.t11 55.8337
R115 a_n3827_n3924.n3 a_n3827_n3924.t14 55.8337
R116 a_n3827_n3924.n0 a_n3827_n3924.t27 55.8335
R117 a_n3827_n3924.n1 a_n3827_n3924.t15 55.8335
R118 a_n3827_n3924.n9 a_n3827_n3924.t12 55.8335
R119 a_n3827_n3924.n9 a_n3827_n3924.t26 55.8335
R120 a_n3827_n3924.n2 a_n3827_n3924.t33 55.8335
R121 a_n3827_n3924.n0 a_n3827_n3924.n19 53.0052
R122 a_n3827_n3924.n0 a_n3827_n3924.n20 53.0052
R123 a_n3827_n3924.n0 a_n3827_n3924.n21 53.0052
R124 a_n3827_n3924.n4 a_n3827_n3924.n22 53.0052
R125 a_n3827_n3924.n3 a_n3827_n3924.n10 53.0052
R126 a_n3827_n3924.n1 a_n3827_n3924.n17 53.0051
R127 a_n3827_n3924.n1 a_n3827_n3924.n16 53.0051
R128 a_n3827_n3924.n1 a_n3827_n3924.n15 53.0051
R129 a_n3827_n3924.n9 a_n3827_n3924.n14 53.0051
R130 a_n3827_n3924.n2 a_n3827_n3924.n13 53.0051
R131 a_n3827_n3924.n2 a_n3827_n3924.n12 53.0051
R132 a_n3827_n3924.n23 a_n3827_n3924.n4 53.0051
R133 a_n3827_n3924.n11 a_n3827_n3924.n3 12.1986
R134 a_n3827_n3924.n0 a_n3827_n3924.n18 12.1986
R135 a_n3827_n3924.n2 a_n3827_n3924.n11 5.11903
R136 a_n3827_n3924.n18 a_n3827_n3924.n1 5.11903
R137 a_n3827_n3924.n19 a_n3827_n3924.t34 2.82907
R138 a_n3827_n3924.n19 a_n3827_n3924.t30 2.82907
R139 a_n3827_n3924.n20 a_n3827_n3924.t24 2.82907
R140 a_n3827_n3924.n20 a_n3827_n3924.t32 2.82907
R141 a_n3827_n3924.n21 a_n3827_n3924.t39 2.82907
R142 a_n3827_n3924.n21 a_n3827_n3924.t31 2.82907
R143 a_n3827_n3924.n22 a_n3827_n3924.t21 2.82907
R144 a_n3827_n3924.n22 a_n3827_n3924.t6 2.82907
R145 a_n3827_n3924.n10 a_n3827_n3924.t17 2.82907
R146 a_n3827_n3924.n10 a_n3827_n3924.t10 2.82907
R147 a_n3827_n3924.n17 a_n3827_n3924.t8 2.82907
R148 a_n3827_n3924.n17 a_n3827_n3924.t16 2.82907
R149 a_n3827_n3924.n16 a_n3827_n3924.t2 2.82907
R150 a_n3827_n3924.n16 a_n3827_n3924.t20 2.82907
R151 a_n3827_n3924.n15 a_n3827_n3924.t4 2.82907
R152 a_n3827_n3924.n15 a_n3827_n3924.t3 2.82907
R153 a_n3827_n3924.n14 a_n3827_n3924.t28 2.82907
R154 a_n3827_n3924.n14 a_n3827_n3924.t29 2.82907
R155 a_n3827_n3924.n13 a_n3827_n3924.t25 2.82907
R156 a_n3827_n3924.n13 a_n3827_n3924.t35 2.82907
R157 a_n3827_n3924.n12 a_n3827_n3924.t38 2.82907
R158 a_n3827_n3924.n12 a_n3827_n3924.t36 2.82907
R159 a_n3827_n3924.n23 a_n3827_n3924.t18 2.82907
R160 a_n3827_n3924.t0 a_n3827_n3924.n23 2.82907
R161 a_n3827_n3924.n4 a_n3827_n3924.n0 2.45524
R162 a_n3827_n3924.n6 a_n3827_n3924.n8 2.01503
R163 a_n3827_n3924.n1 a_n3827_n3924.n9 2.01128
R164 a_n3827_n3924.n18 a_n3827_n3924.n7 1.95694
R165 a_n3827_n3924.n11 a_n3827_n3924.n6 1.95694
R166 a_n3827_n3924.n9 a_n3827_n3924.n2 1.77636
R167 a_n3827_n3924.n6 a_n3827_n3924.n5 1.34352
R168 a_n3827_n3924.n5 a_n3827_n3924.n7 1.34352
R169 a_n3827_n3924.n4 a_n3827_n3924.n3 1.3324
R170 a_n9628_8799.n228 a_n9628_8799.t137 485.149
R171 a_n9628_8799.n290 a_n9628_8799.t152 485.149
R172 a_n9628_8799.n353 a_n9628_8799.t75 485.149
R173 a_n9628_8799.n38 a_n9628_8799.t89 485.149
R174 a_n9628_8799.n100 a_n9628_8799.t102 485.149
R175 a_n9628_8799.n163 a_n9628_8799.t73 485.149
R176 a_n9628_8799.n271 a_n9628_8799.t47 464.166
R177 a_n9628_8799.n270 a_n9628_8799.t45 464.166
R178 a_n9628_8799.n212 a_n9628_8799.t131 464.166
R179 a_n9628_8799.n264 a_n9628_8799.t67 464.166
R180 a_n9628_8799.n263 a_n9628_8799.t50 464.166
R181 a_n9628_8799.n215 a_n9628_8799.t138 464.166
R182 a_n9628_8799.n257 a_n9628_8799.t93 464.166
R183 a_n9628_8799.n256 a_n9628_8799.t68 464.166
R184 a_n9628_8799.n218 a_n9628_8799.t156 464.166
R185 a_n9628_8799.n250 a_n9628_8799.t111 464.166
R186 a_n9628_8799.n249 a_n9628_8799.t71 464.166
R187 a_n9628_8799.n221 a_n9628_8799.t150 464.166
R188 a_n9628_8799.n243 a_n9628_8799.t113 464.166
R189 a_n9628_8799.n242 a_n9628_8799.t85 464.166
R190 a_n9628_8799.n224 a_n9628_8799.t46 464.166
R191 a_n9628_8799.n236 a_n9628_8799.t134 464.166
R192 a_n9628_8799.n235 a_n9628_8799.t115 464.166
R193 a_n9628_8799.n227 a_n9628_8799.t51 464.166
R194 a_n9628_8799.n229 a_n9628_8799.t141 464.166
R195 a_n9628_8799.n333 a_n9628_8799.t58 464.166
R196 a_n9628_8799.n332 a_n9628_8799.t57 464.166
R197 a_n9628_8799.n274 a_n9628_8799.t148 464.166
R198 a_n9628_8799.n326 a_n9628_8799.t76 464.166
R199 a_n9628_8799.n325 a_n9628_8799.t65 464.166
R200 a_n9628_8799.n277 a_n9628_8799.t151 464.166
R201 a_n9628_8799.n319 a_n9628_8799.t107 464.166
R202 a_n9628_8799.n318 a_n9628_8799.t79 464.166
R203 a_n9628_8799.n280 a_n9628_8799.t49 464.166
R204 a_n9628_8799.n312 a_n9628_8799.t124 464.166
R205 a_n9628_8799.n311 a_n9628_8799.t80 464.166
R206 a_n9628_8799.n283 a_n9628_8799.t41 464.166
R207 a_n9628_8799.n305 a_n9628_8799.t129 464.166
R208 a_n9628_8799.n304 a_n9628_8799.t95 464.166
R209 a_n9628_8799.n286 a_n9628_8799.t59 464.166
R210 a_n9628_8799.n298 a_n9628_8799.t149 464.166
R211 a_n9628_8799.n297 a_n9628_8799.t130 464.166
R212 a_n9628_8799.n289 a_n9628_8799.t66 464.166
R213 a_n9628_8799.n291 a_n9628_8799.t153 464.166
R214 a_n9628_8799.n396 a_n9628_8799.t106 464.166
R215 a_n9628_8799.n395 a_n9628_8799.t128 464.166
R216 a_n9628_8799.n337 a_n9628_8799.t64 464.166
R217 a_n9628_8799.n389 a_n9628_8799.t146 464.166
R218 a_n9628_8799.n388 a_n9628_8799.t83 464.166
R219 a_n9628_8799.n340 a_n9628_8799.t139 464.166
R220 a_n9628_8799.n382 a_n9628_8799.t70 464.166
R221 a_n9628_8799.n381 a_n9628_8799.t118 464.166
R222 a_n9628_8799.n343 a_n9628_8799.t55 464.166
R223 a_n9628_8799.n375 a_n9628_8799.t101 464.166
R224 a_n9628_8799.n374 a_n9628_8799.t78 464.166
R225 a_n9628_8799.n346 a_n9628_8799.t126 464.166
R226 a_n9628_8799.n368 a_n9628_8799.t62 464.166
R227 a_n9628_8799.n367 a_n9628_8799.t110 464.166
R228 a_n9628_8799.n349 a_n9628_8799.t44 464.166
R229 a_n9628_8799.n361 a_n9628_8799.t94 464.166
R230 a_n9628_8799.n360 a_n9628_8799.t158 464.166
R231 a_n9628_8799.n352 a_n9628_8799.t117 464.166
R232 a_n9628_8799.n354 a_n9628_8799.t54 464.166
R233 a_n9628_8799.n39 a_n9628_8799.t91 464.166
R234 a_n9628_8799.n41 a_n9628_8799.t123 464.166
R235 a_n9628_8799.n45 a_n9628_8799.t48 464.166
R236 a_n9628_8799.n46 a_n9628_8799.t88 464.166
R237 a_n9628_8799.n34 a_n9628_8799.t120 464.166
R238 a_n9628_8799.n52 a_n9628_8799.t42 464.166
R239 a_n9628_8799.n53 a_n9628_8799.t74 464.166
R240 a_n9628_8799.n57 a_n9628_8799.t112 464.166
R241 a_n9628_8799.n59 a_n9628_8799.t147 464.166
R242 a_n9628_8799.n30 a_n9628_8799.t72 464.166
R243 a_n9628_8799.n64 a_n9628_8799.t108 464.166
R244 a_n9628_8799.n28 a_n9628_8799.t143 464.166
R245 a_n9628_8799.n69 a_n9628_8799.t144 464.166
R246 a_n9628_8799.n71 a_n9628_8799.t90 464.166
R247 a_n9628_8799.n75 a_n9628_8799.t122 464.166
R248 a_n9628_8799.n76 a_n9628_8799.t142 464.166
R249 a_n9628_8799.n24 a_n9628_8799.t86 464.166
R250 a_n9628_8799.n82 a_n9628_8799.t87 464.166
R251 a_n9628_8799.n83 a_n9628_8799.t119 464.166
R252 a_n9628_8799.n101 a_n9628_8799.t104 464.166
R253 a_n9628_8799.n103 a_n9628_8799.t140 464.166
R254 a_n9628_8799.n107 a_n9628_8799.t60 464.166
R255 a_n9628_8799.n108 a_n9628_8799.t98 464.166
R256 a_n9628_8799.n96 a_n9628_8799.t132 464.166
R257 a_n9628_8799.n114 a_n9628_8799.t56 464.166
R258 a_n9628_8799.n115 a_n9628_8799.t84 464.166
R259 a_n9628_8799.n119 a_n9628_8799.t125 464.166
R260 a_n9628_8799.n121 a_n9628_8799.t159 464.166
R261 a_n9628_8799.n92 a_n9628_8799.t81 464.166
R262 a_n9628_8799.n126 a_n9628_8799.t121 464.166
R263 a_n9628_8799.n90 a_n9628_8799.t155 464.166
R264 a_n9628_8799.n131 a_n9628_8799.t157 464.166
R265 a_n9628_8799.n133 a_n9628_8799.t103 464.166
R266 a_n9628_8799.n137 a_n9628_8799.t136 464.166
R267 a_n9628_8799.n138 a_n9628_8799.t154 464.166
R268 a_n9628_8799.n86 a_n9628_8799.t97 464.166
R269 a_n9628_8799.n144 a_n9628_8799.t99 464.166
R270 a_n9628_8799.n145 a_n9628_8799.t133 464.166
R271 a_n9628_8799.n164 a_n9628_8799.t52 464.166
R272 a_n9628_8799.n166 a_n9628_8799.t114 464.166
R273 a_n9628_8799.n170 a_n9628_8799.t69 464.166
R274 a_n9628_8799.n171 a_n9628_8799.t92 464.166
R275 a_n9628_8799.n159 a_n9628_8799.t43 464.166
R276 a_n9628_8799.n177 a_n9628_8799.t109 464.166
R277 a_n9628_8799.n178 a_n9628_8799.t61 464.166
R278 a_n9628_8799.n182 a_n9628_8799.t127 464.166
R279 a_n9628_8799.n184 a_n9628_8799.t77 464.166
R280 a_n9628_8799.n155 a_n9628_8799.t100 464.166
R281 a_n9628_8799.n189 a_n9628_8799.t53 464.166
R282 a_n9628_8799.n153 a_n9628_8799.t116 464.166
R283 a_n9628_8799.n194 a_n9628_8799.t96 464.166
R284 a_n9628_8799.n196 a_n9628_8799.t135 464.166
R285 a_n9628_8799.n200 a_n9628_8799.t82 464.166
R286 a_n9628_8799.n201 a_n9628_8799.t145 464.166
R287 a_n9628_8799.n149 a_n9628_8799.t63 464.166
R288 a_n9628_8799.n207 a_n9628_8799.t40 464.166
R289 a_n9628_8799.n208 a_n9628_8799.t105 464.166
R290 a_n9628_8799.n231 a_n9628_8799.n230 161.3
R291 a_n9628_8799.n232 a_n9628_8799.n227 161.3
R292 a_n9628_8799.n234 a_n9628_8799.n233 161.3
R293 a_n9628_8799.n235 a_n9628_8799.n226 161.3
R294 a_n9628_8799.n236 a_n9628_8799.n225 161.3
R295 a_n9628_8799.n238 a_n9628_8799.n237 161.3
R296 a_n9628_8799.n239 a_n9628_8799.n224 161.3
R297 a_n9628_8799.n241 a_n9628_8799.n240 161.3
R298 a_n9628_8799.n242 a_n9628_8799.n223 161.3
R299 a_n9628_8799.n243 a_n9628_8799.n222 161.3
R300 a_n9628_8799.n245 a_n9628_8799.n244 161.3
R301 a_n9628_8799.n246 a_n9628_8799.n221 161.3
R302 a_n9628_8799.n248 a_n9628_8799.n247 161.3
R303 a_n9628_8799.n249 a_n9628_8799.n220 161.3
R304 a_n9628_8799.n250 a_n9628_8799.n219 161.3
R305 a_n9628_8799.n252 a_n9628_8799.n251 161.3
R306 a_n9628_8799.n253 a_n9628_8799.n218 161.3
R307 a_n9628_8799.n255 a_n9628_8799.n254 161.3
R308 a_n9628_8799.n256 a_n9628_8799.n217 161.3
R309 a_n9628_8799.n257 a_n9628_8799.n216 161.3
R310 a_n9628_8799.n259 a_n9628_8799.n258 161.3
R311 a_n9628_8799.n260 a_n9628_8799.n215 161.3
R312 a_n9628_8799.n262 a_n9628_8799.n261 161.3
R313 a_n9628_8799.n263 a_n9628_8799.n214 161.3
R314 a_n9628_8799.n264 a_n9628_8799.n213 161.3
R315 a_n9628_8799.n266 a_n9628_8799.n265 161.3
R316 a_n9628_8799.n267 a_n9628_8799.n212 161.3
R317 a_n9628_8799.n269 a_n9628_8799.n268 161.3
R318 a_n9628_8799.n270 a_n9628_8799.n211 161.3
R319 a_n9628_8799.n272 a_n9628_8799.n271 161.3
R320 a_n9628_8799.n293 a_n9628_8799.n292 161.3
R321 a_n9628_8799.n294 a_n9628_8799.n289 161.3
R322 a_n9628_8799.n296 a_n9628_8799.n295 161.3
R323 a_n9628_8799.n297 a_n9628_8799.n288 161.3
R324 a_n9628_8799.n298 a_n9628_8799.n287 161.3
R325 a_n9628_8799.n300 a_n9628_8799.n299 161.3
R326 a_n9628_8799.n301 a_n9628_8799.n286 161.3
R327 a_n9628_8799.n303 a_n9628_8799.n302 161.3
R328 a_n9628_8799.n304 a_n9628_8799.n285 161.3
R329 a_n9628_8799.n305 a_n9628_8799.n284 161.3
R330 a_n9628_8799.n307 a_n9628_8799.n306 161.3
R331 a_n9628_8799.n308 a_n9628_8799.n283 161.3
R332 a_n9628_8799.n310 a_n9628_8799.n309 161.3
R333 a_n9628_8799.n311 a_n9628_8799.n282 161.3
R334 a_n9628_8799.n312 a_n9628_8799.n281 161.3
R335 a_n9628_8799.n314 a_n9628_8799.n313 161.3
R336 a_n9628_8799.n315 a_n9628_8799.n280 161.3
R337 a_n9628_8799.n317 a_n9628_8799.n316 161.3
R338 a_n9628_8799.n318 a_n9628_8799.n279 161.3
R339 a_n9628_8799.n319 a_n9628_8799.n278 161.3
R340 a_n9628_8799.n321 a_n9628_8799.n320 161.3
R341 a_n9628_8799.n322 a_n9628_8799.n277 161.3
R342 a_n9628_8799.n324 a_n9628_8799.n323 161.3
R343 a_n9628_8799.n325 a_n9628_8799.n276 161.3
R344 a_n9628_8799.n326 a_n9628_8799.n275 161.3
R345 a_n9628_8799.n328 a_n9628_8799.n327 161.3
R346 a_n9628_8799.n329 a_n9628_8799.n274 161.3
R347 a_n9628_8799.n331 a_n9628_8799.n330 161.3
R348 a_n9628_8799.n332 a_n9628_8799.n273 161.3
R349 a_n9628_8799.n334 a_n9628_8799.n333 161.3
R350 a_n9628_8799.n356 a_n9628_8799.n355 161.3
R351 a_n9628_8799.n357 a_n9628_8799.n352 161.3
R352 a_n9628_8799.n359 a_n9628_8799.n358 161.3
R353 a_n9628_8799.n360 a_n9628_8799.n351 161.3
R354 a_n9628_8799.n361 a_n9628_8799.n350 161.3
R355 a_n9628_8799.n363 a_n9628_8799.n362 161.3
R356 a_n9628_8799.n364 a_n9628_8799.n349 161.3
R357 a_n9628_8799.n366 a_n9628_8799.n365 161.3
R358 a_n9628_8799.n367 a_n9628_8799.n348 161.3
R359 a_n9628_8799.n368 a_n9628_8799.n347 161.3
R360 a_n9628_8799.n370 a_n9628_8799.n369 161.3
R361 a_n9628_8799.n371 a_n9628_8799.n346 161.3
R362 a_n9628_8799.n373 a_n9628_8799.n372 161.3
R363 a_n9628_8799.n374 a_n9628_8799.n345 161.3
R364 a_n9628_8799.n375 a_n9628_8799.n344 161.3
R365 a_n9628_8799.n377 a_n9628_8799.n376 161.3
R366 a_n9628_8799.n378 a_n9628_8799.n343 161.3
R367 a_n9628_8799.n380 a_n9628_8799.n379 161.3
R368 a_n9628_8799.n381 a_n9628_8799.n342 161.3
R369 a_n9628_8799.n382 a_n9628_8799.n341 161.3
R370 a_n9628_8799.n384 a_n9628_8799.n383 161.3
R371 a_n9628_8799.n385 a_n9628_8799.n340 161.3
R372 a_n9628_8799.n387 a_n9628_8799.n386 161.3
R373 a_n9628_8799.n388 a_n9628_8799.n339 161.3
R374 a_n9628_8799.n389 a_n9628_8799.n338 161.3
R375 a_n9628_8799.n391 a_n9628_8799.n390 161.3
R376 a_n9628_8799.n392 a_n9628_8799.n337 161.3
R377 a_n9628_8799.n394 a_n9628_8799.n393 161.3
R378 a_n9628_8799.n395 a_n9628_8799.n336 161.3
R379 a_n9628_8799.n397 a_n9628_8799.n396 161.3
R380 a_n9628_8799.n84 a_n9628_8799.n83 161.3
R381 a_n9628_8799.n82 a_n9628_8799.n23 161.3
R382 a_n9628_8799.n81 a_n9628_8799.n80 161.3
R383 a_n9628_8799.n79 a_n9628_8799.n24 161.3
R384 a_n9628_8799.n78 a_n9628_8799.n77 161.3
R385 a_n9628_8799.n76 a_n9628_8799.n25 161.3
R386 a_n9628_8799.n75 a_n9628_8799.n74 161.3
R387 a_n9628_8799.n73 a_n9628_8799.n26 161.3
R388 a_n9628_8799.n72 a_n9628_8799.n71 161.3
R389 a_n9628_8799.n70 a_n9628_8799.n27 161.3
R390 a_n9628_8799.n69 a_n9628_8799.n68 161.3
R391 a_n9628_8799.n67 a_n9628_8799.n28 161.3
R392 a_n9628_8799.n66 a_n9628_8799.n65 161.3
R393 a_n9628_8799.n64 a_n9628_8799.n29 161.3
R394 a_n9628_8799.n63 a_n9628_8799.n62 161.3
R395 a_n9628_8799.n61 a_n9628_8799.n30 161.3
R396 a_n9628_8799.n60 a_n9628_8799.n59 161.3
R397 a_n9628_8799.n58 a_n9628_8799.n31 161.3
R398 a_n9628_8799.n57 a_n9628_8799.n56 161.3
R399 a_n9628_8799.n55 a_n9628_8799.n32 161.3
R400 a_n9628_8799.n54 a_n9628_8799.n53 161.3
R401 a_n9628_8799.n52 a_n9628_8799.n33 161.3
R402 a_n9628_8799.n51 a_n9628_8799.n50 161.3
R403 a_n9628_8799.n49 a_n9628_8799.n34 161.3
R404 a_n9628_8799.n48 a_n9628_8799.n47 161.3
R405 a_n9628_8799.n46 a_n9628_8799.n35 161.3
R406 a_n9628_8799.n45 a_n9628_8799.n44 161.3
R407 a_n9628_8799.n43 a_n9628_8799.n36 161.3
R408 a_n9628_8799.n42 a_n9628_8799.n41 161.3
R409 a_n9628_8799.n40 a_n9628_8799.n37 161.3
R410 a_n9628_8799.n146 a_n9628_8799.n145 161.3
R411 a_n9628_8799.n144 a_n9628_8799.n85 161.3
R412 a_n9628_8799.n143 a_n9628_8799.n142 161.3
R413 a_n9628_8799.n141 a_n9628_8799.n86 161.3
R414 a_n9628_8799.n140 a_n9628_8799.n139 161.3
R415 a_n9628_8799.n138 a_n9628_8799.n87 161.3
R416 a_n9628_8799.n137 a_n9628_8799.n136 161.3
R417 a_n9628_8799.n135 a_n9628_8799.n88 161.3
R418 a_n9628_8799.n134 a_n9628_8799.n133 161.3
R419 a_n9628_8799.n132 a_n9628_8799.n89 161.3
R420 a_n9628_8799.n131 a_n9628_8799.n130 161.3
R421 a_n9628_8799.n129 a_n9628_8799.n90 161.3
R422 a_n9628_8799.n128 a_n9628_8799.n127 161.3
R423 a_n9628_8799.n126 a_n9628_8799.n91 161.3
R424 a_n9628_8799.n125 a_n9628_8799.n124 161.3
R425 a_n9628_8799.n123 a_n9628_8799.n92 161.3
R426 a_n9628_8799.n122 a_n9628_8799.n121 161.3
R427 a_n9628_8799.n120 a_n9628_8799.n93 161.3
R428 a_n9628_8799.n119 a_n9628_8799.n118 161.3
R429 a_n9628_8799.n117 a_n9628_8799.n94 161.3
R430 a_n9628_8799.n116 a_n9628_8799.n115 161.3
R431 a_n9628_8799.n114 a_n9628_8799.n95 161.3
R432 a_n9628_8799.n113 a_n9628_8799.n112 161.3
R433 a_n9628_8799.n111 a_n9628_8799.n96 161.3
R434 a_n9628_8799.n110 a_n9628_8799.n109 161.3
R435 a_n9628_8799.n108 a_n9628_8799.n97 161.3
R436 a_n9628_8799.n107 a_n9628_8799.n106 161.3
R437 a_n9628_8799.n105 a_n9628_8799.n98 161.3
R438 a_n9628_8799.n104 a_n9628_8799.n103 161.3
R439 a_n9628_8799.n102 a_n9628_8799.n99 161.3
R440 a_n9628_8799.n209 a_n9628_8799.n208 161.3
R441 a_n9628_8799.n207 a_n9628_8799.n148 161.3
R442 a_n9628_8799.n206 a_n9628_8799.n205 161.3
R443 a_n9628_8799.n204 a_n9628_8799.n149 161.3
R444 a_n9628_8799.n203 a_n9628_8799.n202 161.3
R445 a_n9628_8799.n201 a_n9628_8799.n150 161.3
R446 a_n9628_8799.n200 a_n9628_8799.n199 161.3
R447 a_n9628_8799.n198 a_n9628_8799.n151 161.3
R448 a_n9628_8799.n197 a_n9628_8799.n196 161.3
R449 a_n9628_8799.n195 a_n9628_8799.n152 161.3
R450 a_n9628_8799.n194 a_n9628_8799.n193 161.3
R451 a_n9628_8799.n192 a_n9628_8799.n153 161.3
R452 a_n9628_8799.n191 a_n9628_8799.n190 161.3
R453 a_n9628_8799.n189 a_n9628_8799.n154 161.3
R454 a_n9628_8799.n188 a_n9628_8799.n187 161.3
R455 a_n9628_8799.n186 a_n9628_8799.n155 161.3
R456 a_n9628_8799.n185 a_n9628_8799.n184 161.3
R457 a_n9628_8799.n183 a_n9628_8799.n156 161.3
R458 a_n9628_8799.n182 a_n9628_8799.n181 161.3
R459 a_n9628_8799.n180 a_n9628_8799.n157 161.3
R460 a_n9628_8799.n179 a_n9628_8799.n178 161.3
R461 a_n9628_8799.n177 a_n9628_8799.n158 161.3
R462 a_n9628_8799.n176 a_n9628_8799.n175 161.3
R463 a_n9628_8799.n174 a_n9628_8799.n159 161.3
R464 a_n9628_8799.n173 a_n9628_8799.n172 161.3
R465 a_n9628_8799.n171 a_n9628_8799.n160 161.3
R466 a_n9628_8799.n170 a_n9628_8799.n169 161.3
R467 a_n9628_8799.n168 a_n9628_8799.n161 161.3
R468 a_n9628_8799.n167 a_n9628_8799.n166 161.3
R469 a_n9628_8799.n165 a_n9628_8799.n162 161.3
R470 a_n9628_8799.n13 a_n9628_8799.n11 98.9633
R471 a_n9628_8799.n2 a_n9628_8799.n0 98.9631
R472 a_n9628_8799.n21 a_n9628_8799.n20 98.6055
R473 a_n9628_8799.n19 a_n9628_8799.n18 98.6055
R474 a_n9628_8799.n17 a_n9628_8799.n16 98.6055
R475 a_n9628_8799.n15 a_n9628_8799.n14 98.6055
R476 a_n9628_8799.n13 a_n9628_8799.n12 98.6055
R477 a_n9628_8799.n2 a_n9628_8799.n1 98.6055
R478 a_n9628_8799.n4 a_n9628_8799.n3 98.6055
R479 a_n9628_8799.n6 a_n9628_8799.n5 98.6055
R480 a_n9628_8799.n8 a_n9628_8799.n7 98.6055
R481 a_n9628_8799.n10 a_n9628_8799.n9 98.6055
R482 a_n9628_8799.n415 a_n9628_8799.n414 81.3766
R483 a_n9628_8799.n403 a_n9628_8799.n401 81.3764
R484 a_n9628_8799.n411 a_n9628_8799.n409 81.3764
R485 a_n9628_8799.n408 a_n9628_8799.n407 80.9324
R486 a_n9628_8799.n406 a_n9628_8799.n405 80.9324
R487 a_n9628_8799.n403 a_n9628_8799.n402 80.9324
R488 a_n9628_8799.n411 a_n9628_8799.n410 80.9324
R489 a_n9628_8799.n414 a_n9628_8799.n413 80.9324
R490 a_n9628_8799.n231 a_n9628_8799.n228 70.4033
R491 a_n9628_8799.n293 a_n9628_8799.n290 70.4033
R492 a_n9628_8799.n356 a_n9628_8799.n353 70.4033
R493 a_n9628_8799.n38 a_n9628_8799.n37 70.4033
R494 a_n9628_8799.n100 a_n9628_8799.n99 70.4033
R495 a_n9628_8799.n163 a_n9628_8799.n162 70.4033
R496 a_n9628_8799.n271 a_n9628_8799.n270 48.2005
R497 a_n9628_8799.n264 a_n9628_8799.n263 48.2005
R498 a_n9628_8799.n257 a_n9628_8799.n256 48.2005
R499 a_n9628_8799.n250 a_n9628_8799.n249 48.2005
R500 a_n9628_8799.n243 a_n9628_8799.n242 48.2005
R501 a_n9628_8799.n236 a_n9628_8799.n235 48.2005
R502 a_n9628_8799.n333 a_n9628_8799.n332 48.2005
R503 a_n9628_8799.n326 a_n9628_8799.n325 48.2005
R504 a_n9628_8799.n319 a_n9628_8799.n318 48.2005
R505 a_n9628_8799.n312 a_n9628_8799.n311 48.2005
R506 a_n9628_8799.n305 a_n9628_8799.n304 48.2005
R507 a_n9628_8799.n298 a_n9628_8799.n297 48.2005
R508 a_n9628_8799.n396 a_n9628_8799.n395 48.2005
R509 a_n9628_8799.n389 a_n9628_8799.n388 48.2005
R510 a_n9628_8799.n382 a_n9628_8799.n381 48.2005
R511 a_n9628_8799.n375 a_n9628_8799.n374 48.2005
R512 a_n9628_8799.n368 a_n9628_8799.n367 48.2005
R513 a_n9628_8799.n361 a_n9628_8799.n360 48.2005
R514 a_n9628_8799.n46 a_n9628_8799.n45 48.2005
R515 a_n9628_8799.n53 a_n9628_8799.n52 48.2005
R516 a_n9628_8799.n59 a_n9628_8799.n30 48.2005
R517 a_n9628_8799.n69 a_n9628_8799.n28 48.2005
R518 a_n9628_8799.n76 a_n9628_8799.n75 48.2005
R519 a_n9628_8799.n83 a_n9628_8799.n82 48.2005
R520 a_n9628_8799.n108 a_n9628_8799.n107 48.2005
R521 a_n9628_8799.n115 a_n9628_8799.n114 48.2005
R522 a_n9628_8799.n121 a_n9628_8799.n92 48.2005
R523 a_n9628_8799.n131 a_n9628_8799.n90 48.2005
R524 a_n9628_8799.n138 a_n9628_8799.n137 48.2005
R525 a_n9628_8799.n145 a_n9628_8799.n144 48.2005
R526 a_n9628_8799.n171 a_n9628_8799.n170 48.2005
R527 a_n9628_8799.n178 a_n9628_8799.n177 48.2005
R528 a_n9628_8799.n184 a_n9628_8799.n155 48.2005
R529 a_n9628_8799.n194 a_n9628_8799.n153 48.2005
R530 a_n9628_8799.n201 a_n9628_8799.n200 48.2005
R531 a_n9628_8799.n208 a_n9628_8799.n207 48.2005
R532 a_n9628_8799.n269 a_n9628_8799.n212 40.1672
R533 a_n9628_8799.n230 a_n9628_8799.n227 40.1672
R534 a_n9628_8799.n331 a_n9628_8799.n274 40.1672
R535 a_n9628_8799.n292 a_n9628_8799.n289 40.1672
R536 a_n9628_8799.n394 a_n9628_8799.n337 40.1672
R537 a_n9628_8799.n355 a_n9628_8799.n352 40.1672
R538 a_n9628_8799.n41 a_n9628_8799.n40 40.1672
R539 a_n9628_8799.n81 a_n9628_8799.n24 40.1672
R540 a_n9628_8799.n103 a_n9628_8799.n102 40.1672
R541 a_n9628_8799.n143 a_n9628_8799.n86 40.1672
R542 a_n9628_8799.n166 a_n9628_8799.n165 40.1672
R543 a_n9628_8799.n206 a_n9628_8799.n149 40.1672
R544 a_n9628_8799.n262 a_n9628_8799.n215 38.7066
R545 a_n9628_8799.n237 a_n9628_8799.n224 38.7066
R546 a_n9628_8799.n324 a_n9628_8799.n277 38.7066
R547 a_n9628_8799.n299 a_n9628_8799.n286 38.7066
R548 a_n9628_8799.n387 a_n9628_8799.n340 38.7066
R549 a_n9628_8799.n362 a_n9628_8799.n349 38.7066
R550 a_n9628_8799.n47 a_n9628_8799.n34 38.7066
R551 a_n9628_8799.n71 a_n9628_8799.n26 38.7066
R552 a_n9628_8799.n109 a_n9628_8799.n96 38.7066
R553 a_n9628_8799.n133 a_n9628_8799.n88 38.7066
R554 a_n9628_8799.n172 a_n9628_8799.n159 38.7066
R555 a_n9628_8799.n196 a_n9628_8799.n151 38.7066
R556 a_n9628_8799.n255 a_n9628_8799.n218 37.246
R557 a_n9628_8799.n244 a_n9628_8799.n221 37.246
R558 a_n9628_8799.n317 a_n9628_8799.n280 37.246
R559 a_n9628_8799.n306 a_n9628_8799.n283 37.246
R560 a_n9628_8799.n380 a_n9628_8799.n343 37.246
R561 a_n9628_8799.n369 a_n9628_8799.n346 37.246
R562 a_n9628_8799.n57 a_n9628_8799.n32 37.246
R563 a_n9628_8799.n65 a_n9628_8799.n64 37.246
R564 a_n9628_8799.n119 a_n9628_8799.n94 37.246
R565 a_n9628_8799.n127 a_n9628_8799.n126 37.246
R566 a_n9628_8799.n182 a_n9628_8799.n157 37.246
R567 a_n9628_8799.n190 a_n9628_8799.n189 37.246
R568 a_n9628_8799.n251 a_n9628_8799.n218 35.7853
R569 a_n9628_8799.n248 a_n9628_8799.n221 35.7853
R570 a_n9628_8799.n313 a_n9628_8799.n280 35.7853
R571 a_n9628_8799.n310 a_n9628_8799.n283 35.7853
R572 a_n9628_8799.n376 a_n9628_8799.n343 35.7853
R573 a_n9628_8799.n373 a_n9628_8799.n346 35.7853
R574 a_n9628_8799.n58 a_n9628_8799.n57 35.7853
R575 a_n9628_8799.n64 a_n9628_8799.n63 35.7853
R576 a_n9628_8799.n120 a_n9628_8799.n119 35.7853
R577 a_n9628_8799.n126 a_n9628_8799.n125 35.7853
R578 a_n9628_8799.n183 a_n9628_8799.n182 35.7853
R579 a_n9628_8799.n189 a_n9628_8799.n188 35.7853
R580 a_n9628_8799.n258 a_n9628_8799.n215 34.3247
R581 a_n9628_8799.n241 a_n9628_8799.n224 34.3247
R582 a_n9628_8799.n320 a_n9628_8799.n277 34.3247
R583 a_n9628_8799.n303 a_n9628_8799.n286 34.3247
R584 a_n9628_8799.n383 a_n9628_8799.n340 34.3247
R585 a_n9628_8799.n366 a_n9628_8799.n349 34.3247
R586 a_n9628_8799.n51 a_n9628_8799.n34 34.3247
R587 a_n9628_8799.n71 a_n9628_8799.n70 34.3247
R588 a_n9628_8799.n113 a_n9628_8799.n96 34.3247
R589 a_n9628_8799.n133 a_n9628_8799.n132 34.3247
R590 a_n9628_8799.n176 a_n9628_8799.n159 34.3247
R591 a_n9628_8799.n196 a_n9628_8799.n195 34.3247
R592 a_n9628_8799.n22 a_n9628_8799.n10 33.7114
R593 a_n9628_8799.n265 a_n9628_8799.n212 32.8641
R594 a_n9628_8799.n234 a_n9628_8799.n227 32.8641
R595 a_n9628_8799.n327 a_n9628_8799.n274 32.8641
R596 a_n9628_8799.n296 a_n9628_8799.n289 32.8641
R597 a_n9628_8799.n390 a_n9628_8799.n337 32.8641
R598 a_n9628_8799.n359 a_n9628_8799.n352 32.8641
R599 a_n9628_8799.n41 a_n9628_8799.n36 32.8641
R600 a_n9628_8799.n77 a_n9628_8799.n24 32.8641
R601 a_n9628_8799.n103 a_n9628_8799.n98 32.8641
R602 a_n9628_8799.n139 a_n9628_8799.n86 32.8641
R603 a_n9628_8799.n166 a_n9628_8799.n161 32.8641
R604 a_n9628_8799.n202 a_n9628_8799.n149 32.8641
R605 a_n9628_8799.n412 a_n9628_8799.n408 32.0866
R606 a_n9628_8799.n22 a_n9628_8799.n21 21.1779
R607 a_n9628_8799.n229 a_n9628_8799.n228 20.9576
R608 a_n9628_8799.n291 a_n9628_8799.n290 20.9576
R609 a_n9628_8799.n354 a_n9628_8799.n353 20.9576
R610 a_n9628_8799.n39 a_n9628_8799.n38 20.9576
R611 a_n9628_8799.n101 a_n9628_8799.n100 20.9576
R612 a_n9628_8799.n164 a_n9628_8799.n163 20.9576
R613 a_n9628_8799.n265 a_n9628_8799.n264 15.3369
R614 a_n9628_8799.n235 a_n9628_8799.n234 15.3369
R615 a_n9628_8799.n327 a_n9628_8799.n326 15.3369
R616 a_n9628_8799.n297 a_n9628_8799.n296 15.3369
R617 a_n9628_8799.n390 a_n9628_8799.n389 15.3369
R618 a_n9628_8799.n360 a_n9628_8799.n359 15.3369
R619 a_n9628_8799.n45 a_n9628_8799.n36 15.3369
R620 a_n9628_8799.n77 a_n9628_8799.n76 15.3369
R621 a_n9628_8799.n107 a_n9628_8799.n98 15.3369
R622 a_n9628_8799.n139 a_n9628_8799.n138 15.3369
R623 a_n9628_8799.n170 a_n9628_8799.n161 15.3369
R624 a_n9628_8799.n202 a_n9628_8799.n201 15.3369
R625 a_n9628_8799.n258 a_n9628_8799.n257 13.8763
R626 a_n9628_8799.n242 a_n9628_8799.n241 13.8763
R627 a_n9628_8799.n320 a_n9628_8799.n319 13.8763
R628 a_n9628_8799.n304 a_n9628_8799.n303 13.8763
R629 a_n9628_8799.n383 a_n9628_8799.n382 13.8763
R630 a_n9628_8799.n367 a_n9628_8799.n366 13.8763
R631 a_n9628_8799.n52 a_n9628_8799.n51 13.8763
R632 a_n9628_8799.n70 a_n9628_8799.n69 13.8763
R633 a_n9628_8799.n114 a_n9628_8799.n113 13.8763
R634 a_n9628_8799.n132 a_n9628_8799.n131 13.8763
R635 a_n9628_8799.n177 a_n9628_8799.n176 13.8763
R636 a_n9628_8799.n195 a_n9628_8799.n194 13.8763
R637 a_n9628_8799.n251 a_n9628_8799.n250 12.4157
R638 a_n9628_8799.n249 a_n9628_8799.n248 12.4157
R639 a_n9628_8799.n313 a_n9628_8799.n312 12.4157
R640 a_n9628_8799.n311 a_n9628_8799.n310 12.4157
R641 a_n9628_8799.n376 a_n9628_8799.n375 12.4157
R642 a_n9628_8799.n374 a_n9628_8799.n373 12.4157
R643 a_n9628_8799.n59 a_n9628_8799.n58 12.4157
R644 a_n9628_8799.n63 a_n9628_8799.n30 12.4157
R645 a_n9628_8799.n121 a_n9628_8799.n120 12.4157
R646 a_n9628_8799.n125 a_n9628_8799.n92 12.4157
R647 a_n9628_8799.n184 a_n9628_8799.n183 12.4157
R648 a_n9628_8799.n188 a_n9628_8799.n155 12.4157
R649 a_n9628_8799.n404 a_n9628_8799.n400 12.3339
R650 a_n9628_8799.n400 a_n9628_8799.n22 11.4887
R651 a_n9628_8799.n256 a_n9628_8799.n255 10.955
R652 a_n9628_8799.n244 a_n9628_8799.n243 10.955
R653 a_n9628_8799.n318 a_n9628_8799.n317 10.955
R654 a_n9628_8799.n306 a_n9628_8799.n305 10.955
R655 a_n9628_8799.n381 a_n9628_8799.n380 10.955
R656 a_n9628_8799.n369 a_n9628_8799.n368 10.955
R657 a_n9628_8799.n53 a_n9628_8799.n32 10.955
R658 a_n9628_8799.n65 a_n9628_8799.n28 10.955
R659 a_n9628_8799.n115 a_n9628_8799.n94 10.955
R660 a_n9628_8799.n127 a_n9628_8799.n90 10.955
R661 a_n9628_8799.n178 a_n9628_8799.n157 10.955
R662 a_n9628_8799.n190 a_n9628_8799.n153 10.955
R663 a_n9628_8799.n263 a_n9628_8799.n262 9.49444
R664 a_n9628_8799.n237 a_n9628_8799.n236 9.49444
R665 a_n9628_8799.n325 a_n9628_8799.n324 9.49444
R666 a_n9628_8799.n299 a_n9628_8799.n298 9.49444
R667 a_n9628_8799.n388 a_n9628_8799.n387 9.49444
R668 a_n9628_8799.n362 a_n9628_8799.n361 9.49444
R669 a_n9628_8799.n47 a_n9628_8799.n46 9.49444
R670 a_n9628_8799.n75 a_n9628_8799.n26 9.49444
R671 a_n9628_8799.n109 a_n9628_8799.n108 9.49444
R672 a_n9628_8799.n137 a_n9628_8799.n88 9.49444
R673 a_n9628_8799.n172 a_n9628_8799.n171 9.49444
R674 a_n9628_8799.n200 a_n9628_8799.n151 9.49444
R675 a_n9628_8799.n335 a_n9628_8799.n272 9.04406
R676 a_n9628_8799.n147 a_n9628_8799.n84 9.04406
R677 a_n9628_8799.n270 a_n9628_8799.n269 8.03383
R678 a_n9628_8799.n230 a_n9628_8799.n229 8.03383
R679 a_n9628_8799.n332 a_n9628_8799.n331 8.03383
R680 a_n9628_8799.n292 a_n9628_8799.n291 8.03383
R681 a_n9628_8799.n395 a_n9628_8799.n394 8.03383
R682 a_n9628_8799.n355 a_n9628_8799.n354 8.03383
R683 a_n9628_8799.n40 a_n9628_8799.n39 8.03383
R684 a_n9628_8799.n82 a_n9628_8799.n81 8.03383
R685 a_n9628_8799.n102 a_n9628_8799.n101 8.03383
R686 a_n9628_8799.n144 a_n9628_8799.n143 8.03383
R687 a_n9628_8799.n165 a_n9628_8799.n164 8.03383
R688 a_n9628_8799.n207 a_n9628_8799.n206 8.03383
R689 a_n9628_8799.n399 a_n9628_8799.n210 7.14965
R690 a_n9628_8799.n399 a_n9628_8799.n398 6.85731
R691 a_n9628_8799.n335 a_n9628_8799.n334 4.93611
R692 a_n9628_8799.n398 a_n9628_8799.n397 4.93611
R693 a_n9628_8799.n147 a_n9628_8799.n146 4.93611
R694 a_n9628_8799.n210 a_n9628_8799.n209 4.93611
R695 a_n9628_8799.n398 a_n9628_8799.n335 4.10845
R696 a_n9628_8799.n210 a_n9628_8799.n147 4.10845
R697 a_n9628_8799.n20 a_n9628_8799.t12 3.61217
R698 a_n9628_8799.n20 a_n9628_8799.t11 3.61217
R699 a_n9628_8799.n18 a_n9628_8799.t4 3.61217
R700 a_n9628_8799.n18 a_n9628_8799.t2 3.61217
R701 a_n9628_8799.n16 a_n9628_8799.t38 3.61217
R702 a_n9628_8799.n16 a_n9628_8799.t16 3.61217
R703 a_n9628_8799.n14 a_n9628_8799.t14 3.61217
R704 a_n9628_8799.n14 a_n9628_8799.t5 3.61217
R705 a_n9628_8799.n12 a_n9628_8799.t6 3.61217
R706 a_n9628_8799.n12 a_n9628_8799.t13 3.61217
R707 a_n9628_8799.n11 a_n9628_8799.t15 3.61217
R708 a_n9628_8799.n11 a_n9628_8799.t3 3.61217
R709 a_n9628_8799.n0 a_n9628_8799.t35 3.61217
R710 a_n9628_8799.n0 a_n9628_8799.t7 3.61217
R711 a_n9628_8799.n1 a_n9628_8799.t0 3.61217
R712 a_n9628_8799.n1 a_n9628_8799.t17 3.61217
R713 a_n9628_8799.n3 a_n9628_8799.t37 3.61217
R714 a_n9628_8799.n3 a_n9628_8799.t10 3.61217
R715 a_n9628_8799.n5 a_n9628_8799.t18 3.61217
R716 a_n9628_8799.n5 a_n9628_8799.t8 3.61217
R717 a_n9628_8799.n7 a_n9628_8799.t9 3.61217
R718 a_n9628_8799.n7 a_n9628_8799.t1 3.61217
R719 a_n9628_8799.n9 a_n9628_8799.t39 3.61217
R720 a_n9628_8799.n9 a_n9628_8799.t36 3.61217
R721 a_n9628_8799.n400 a_n9628_8799.n399 3.4105
R722 a_n9628_8799.n409 a_n9628_8799.t29 2.82907
R723 a_n9628_8799.n409 a_n9628_8799.t27 2.82907
R724 a_n9628_8799.n410 a_n9628_8799.t22 2.82907
R725 a_n9628_8799.n410 a_n9628_8799.t26 2.82907
R726 a_n9628_8799.n413 a_n9628_8799.t33 2.82907
R727 a_n9628_8799.n413 a_n9628_8799.t23 2.82907
R728 a_n9628_8799.n407 a_n9628_8799.t32 2.82907
R729 a_n9628_8799.n407 a_n9628_8799.t28 2.82907
R730 a_n9628_8799.n405 a_n9628_8799.t19 2.82907
R731 a_n9628_8799.n405 a_n9628_8799.t31 2.82907
R732 a_n9628_8799.n402 a_n9628_8799.t20 2.82907
R733 a_n9628_8799.n402 a_n9628_8799.t21 2.82907
R734 a_n9628_8799.n401 a_n9628_8799.t24 2.82907
R735 a_n9628_8799.n401 a_n9628_8799.t25 2.82907
R736 a_n9628_8799.n415 a_n9628_8799.t30 2.82907
R737 a_n9628_8799.t34 a_n9628_8799.n415 2.82907
R738 a_n9628_8799.n408 a_n9628_8799.n406 0.444466
R739 a_n9628_8799.n15 a_n9628_8799.n13 0.358259
R740 a_n9628_8799.n17 a_n9628_8799.n15 0.358259
R741 a_n9628_8799.n19 a_n9628_8799.n17 0.358259
R742 a_n9628_8799.n21 a_n9628_8799.n19 0.358259
R743 a_n9628_8799.n10 a_n9628_8799.n8 0.358259
R744 a_n9628_8799.n8 a_n9628_8799.n6 0.358259
R745 a_n9628_8799.n6 a_n9628_8799.n4 0.358259
R746 a_n9628_8799.n4 a_n9628_8799.n2 0.358259
R747 a_n9628_8799.n404 a_n9628_8799.n403 0.222483
R748 a_n9628_8799.n406 a_n9628_8799.n404 0.222483
R749 a_n9628_8799.n414 a_n9628_8799.n412 0.222483
R750 a_n9628_8799.n412 a_n9628_8799.n411 0.222483
R751 a_n9628_8799.n272 a_n9628_8799.n211 0.189894
R752 a_n9628_8799.n268 a_n9628_8799.n211 0.189894
R753 a_n9628_8799.n268 a_n9628_8799.n267 0.189894
R754 a_n9628_8799.n267 a_n9628_8799.n266 0.189894
R755 a_n9628_8799.n266 a_n9628_8799.n213 0.189894
R756 a_n9628_8799.n214 a_n9628_8799.n213 0.189894
R757 a_n9628_8799.n261 a_n9628_8799.n214 0.189894
R758 a_n9628_8799.n261 a_n9628_8799.n260 0.189894
R759 a_n9628_8799.n260 a_n9628_8799.n259 0.189894
R760 a_n9628_8799.n259 a_n9628_8799.n216 0.189894
R761 a_n9628_8799.n217 a_n9628_8799.n216 0.189894
R762 a_n9628_8799.n254 a_n9628_8799.n217 0.189894
R763 a_n9628_8799.n254 a_n9628_8799.n253 0.189894
R764 a_n9628_8799.n253 a_n9628_8799.n252 0.189894
R765 a_n9628_8799.n252 a_n9628_8799.n219 0.189894
R766 a_n9628_8799.n220 a_n9628_8799.n219 0.189894
R767 a_n9628_8799.n247 a_n9628_8799.n220 0.189894
R768 a_n9628_8799.n247 a_n9628_8799.n246 0.189894
R769 a_n9628_8799.n246 a_n9628_8799.n245 0.189894
R770 a_n9628_8799.n245 a_n9628_8799.n222 0.189894
R771 a_n9628_8799.n223 a_n9628_8799.n222 0.189894
R772 a_n9628_8799.n240 a_n9628_8799.n223 0.189894
R773 a_n9628_8799.n240 a_n9628_8799.n239 0.189894
R774 a_n9628_8799.n239 a_n9628_8799.n238 0.189894
R775 a_n9628_8799.n238 a_n9628_8799.n225 0.189894
R776 a_n9628_8799.n226 a_n9628_8799.n225 0.189894
R777 a_n9628_8799.n233 a_n9628_8799.n226 0.189894
R778 a_n9628_8799.n233 a_n9628_8799.n232 0.189894
R779 a_n9628_8799.n232 a_n9628_8799.n231 0.189894
R780 a_n9628_8799.n334 a_n9628_8799.n273 0.189894
R781 a_n9628_8799.n330 a_n9628_8799.n273 0.189894
R782 a_n9628_8799.n330 a_n9628_8799.n329 0.189894
R783 a_n9628_8799.n329 a_n9628_8799.n328 0.189894
R784 a_n9628_8799.n328 a_n9628_8799.n275 0.189894
R785 a_n9628_8799.n276 a_n9628_8799.n275 0.189894
R786 a_n9628_8799.n323 a_n9628_8799.n276 0.189894
R787 a_n9628_8799.n323 a_n9628_8799.n322 0.189894
R788 a_n9628_8799.n322 a_n9628_8799.n321 0.189894
R789 a_n9628_8799.n321 a_n9628_8799.n278 0.189894
R790 a_n9628_8799.n279 a_n9628_8799.n278 0.189894
R791 a_n9628_8799.n316 a_n9628_8799.n279 0.189894
R792 a_n9628_8799.n316 a_n9628_8799.n315 0.189894
R793 a_n9628_8799.n315 a_n9628_8799.n314 0.189894
R794 a_n9628_8799.n314 a_n9628_8799.n281 0.189894
R795 a_n9628_8799.n282 a_n9628_8799.n281 0.189894
R796 a_n9628_8799.n309 a_n9628_8799.n282 0.189894
R797 a_n9628_8799.n309 a_n9628_8799.n308 0.189894
R798 a_n9628_8799.n308 a_n9628_8799.n307 0.189894
R799 a_n9628_8799.n307 a_n9628_8799.n284 0.189894
R800 a_n9628_8799.n285 a_n9628_8799.n284 0.189894
R801 a_n9628_8799.n302 a_n9628_8799.n285 0.189894
R802 a_n9628_8799.n302 a_n9628_8799.n301 0.189894
R803 a_n9628_8799.n301 a_n9628_8799.n300 0.189894
R804 a_n9628_8799.n300 a_n9628_8799.n287 0.189894
R805 a_n9628_8799.n288 a_n9628_8799.n287 0.189894
R806 a_n9628_8799.n295 a_n9628_8799.n288 0.189894
R807 a_n9628_8799.n295 a_n9628_8799.n294 0.189894
R808 a_n9628_8799.n294 a_n9628_8799.n293 0.189894
R809 a_n9628_8799.n397 a_n9628_8799.n336 0.189894
R810 a_n9628_8799.n393 a_n9628_8799.n336 0.189894
R811 a_n9628_8799.n393 a_n9628_8799.n392 0.189894
R812 a_n9628_8799.n392 a_n9628_8799.n391 0.189894
R813 a_n9628_8799.n391 a_n9628_8799.n338 0.189894
R814 a_n9628_8799.n339 a_n9628_8799.n338 0.189894
R815 a_n9628_8799.n386 a_n9628_8799.n339 0.189894
R816 a_n9628_8799.n386 a_n9628_8799.n385 0.189894
R817 a_n9628_8799.n385 a_n9628_8799.n384 0.189894
R818 a_n9628_8799.n384 a_n9628_8799.n341 0.189894
R819 a_n9628_8799.n342 a_n9628_8799.n341 0.189894
R820 a_n9628_8799.n379 a_n9628_8799.n342 0.189894
R821 a_n9628_8799.n379 a_n9628_8799.n378 0.189894
R822 a_n9628_8799.n378 a_n9628_8799.n377 0.189894
R823 a_n9628_8799.n377 a_n9628_8799.n344 0.189894
R824 a_n9628_8799.n345 a_n9628_8799.n344 0.189894
R825 a_n9628_8799.n372 a_n9628_8799.n345 0.189894
R826 a_n9628_8799.n372 a_n9628_8799.n371 0.189894
R827 a_n9628_8799.n371 a_n9628_8799.n370 0.189894
R828 a_n9628_8799.n370 a_n9628_8799.n347 0.189894
R829 a_n9628_8799.n348 a_n9628_8799.n347 0.189894
R830 a_n9628_8799.n365 a_n9628_8799.n348 0.189894
R831 a_n9628_8799.n365 a_n9628_8799.n364 0.189894
R832 a_n9628_8799.n364 a_n9628_8799.n363 0.189894
R833 a_n9628_8799.n363 a_n9628_8799.n350 0.189894
R834 a_n9628_8799.n351 a_n9628_8799.n350 0.189894
R835 a_n9628_8799.n358 a_n9628_8799.n351 0.189894
R836 a_n9628_8799.n358 a_n9628_8799.n357 0.189894
R837 a_n9628_8799.n357 a_n9628_8799.n356 0.189894
R838 a_n9628_8799.n42 a_n9628_8799.n37 0.189894
R839 a_n9628_8799.n43 a_n9628_8799.n42 0.189894
R840 a_n9628_8799.n44 a_n9628_8799.n43 0.189894
R841 a_n9628_8799.n44 a_n9628_8799.n35 0.189894
R842 a_n9628_8799.n48 a_n9628_8799.n35 0.189894
R843 a_n9628_8799.n49 a_n9628_8799.n48 0.189894
R844 a_n9628_8799.n50 a_n9628_8799.n49 0.189894
R845 a_n9628_8799.n50 a_n9628_8799.n33 0.189894
R846 a_n9628_8799.n54 a_n9628_8799.n33 0.189894
R847 a_n9628_8799.n55 a_n9628_8799.n54 0.189894
R848 a_n9628_8799.n56 a_n9628_8799.n55 0.189894
R849 a_n9628_8799.n56 a_n9628_8799.n31 0.189894
R850 a_n9628_8799.n60 a_n9628_8799.n31 0.189894
R851 a_n9628_8799.n61 a_n9628_8799.n60 0.189894
R852 a_n9628_8799.n62 a_n9628_8799.n61 0.189894
R853 a_n9628_8799.n62 a_n9628_8799.n29 0.189894
R854 a_n9628_8799.n66 a_n9628_8799.n29 0.189894
R855 a_n9628_8799.n67 a_n9628_8799.n66 0.189894
R856 a_n9628_8799.n68 a_n9628_8799.n67 0.189894
R857 a_n9628_8799.n68 a_n9628_8799.n27 0.189894
R858 a_n9628_8799.n72 a_n9628_8799.n27 0.189894
R859 a_n9628_8799.n73 a_n9628_8799.n72 0.189894
R860 a_n9628_8799.n74 a_n9628_8799.n73 0.189894
R861 a_n9628_8799.n74 a_n9628_8799.n25 0.189894
R862 a_n9628_8799.n78 a_n9628_8799.n25 0.189894
R863 a_n9628_8799.n79 a_n9628_8799.n78 0.189894
R864 a_n9628_8799.n80 a_n9628_8799.n79 0.189894
R865 a_n9628_8799.n80 a_n9628_8799.n23 0.189894
R866 a_n9628_8799.n84 a_n9628_8799.n23 0.189894
R867 a_n9628_8799.n104 a_n9628_8799.n99 0.189894
R868 a_n9628_8799.n105 a_n9628_8799.n104 0.189894
R869 a_n9628_8799.n106 a_n9628_8799.n105 0.189894
R870 a_n9628_8799.n106 a_n9628_8799.n97 0.189894
R871 a_n9628_8799.n110 a_n9628_8799.n97 0.189894
R872 a_n9628_8799.n111 a_n9628_8799.n110 0.189894
R873 a_n9628_8799.n112 a_n9628_8799.n111 0.189894
R874 a_n9628_8799.n112 a_n9628_8799.n95 0.189894
R875 a_n9628_8799.n116 a_n9628_8799.n95 0.189894
R876 a_n9628_8799.n117 a_n9628_8799.n116 0.189894
R877 a_n9628_8799.n118 a_n9628_8799.n117 0.189894
R878 a_n9628_8799.n118 a_n9628_8799.n93 0.189894
R879 a_n9628_8799.n122 a_n9628_8799.n93 0.189894
R880 a_n9628_8799.n123 a_n9628_8799.n122 0.189894
R881 a_n9628_8799.n124 a_n9628_8799.n123 0.189894
R882 a_n9628_8799.n124 a_n9628_8799.n91 0.189894
R883 a_n9628_8799.n128 a_n9628_8799.n91 0.189894
R884 a_n9628_8799.n129 a_n9628_8799.n128 0.189894
R885 a_n9628_8799.n130 a_n9628_8799.n129 0.189894
R886 a_n9628_8799.n130 a_n9628_8799.n89 0.189894
R887 a_n9628_8799.n134 a_n9628_8799.n89 0.189894
R888 a_n9628_8799.n135 a_n9628_8799.n134 0.189894
R889 a_n9628_8799.n136 a_n9628_8799.n135 0.189894
R890 a_n9628_8799.n136 a_n9628_8799.n87 0.189894
R891 a_n9628_8799.n140 a_n9628_8799.n87 0.189894
R892 a_n9628_8799.n141 a_n9628_8799.n140 0.189894
R893 a_n9628_8799.n142 a_n9628_8799.n141 0.189894
R894 a_n9628_8799.n142 a_n9628_8799.n85 0.189894
R895 a_n9628_8799.n146 a_n9628_8799.n85 0.189894
R896 a_n9628_8799.n167 a_n9628_8799.n162 0.189894
R897 a_n9628_8799.n168 a_n9628_8799.n167 0.189894
R898 a_n9628_8799.n169 a_n9628_8799.n168 0.189894
R899 a_n9628_8799.n169 a_n9628_8799.n160 0.189894
R900 a_n9628_8799.n173 a_n9628_8799.n160 0.189894
R901 a_n9628_8799.n174 a_n9628_8799.n173 0.189894
R902 a_n9628_8799.n175 a_n9628_8799.n174 0.189894
R903 a_n9628_8799.n175 a_n9628_8799.n158 0.189894
R904 a_n9628_8799.n179 a_n9628_8799.n158 0.189894
R905 a_n9628_8799.n180 a_n9628_8799.n179 0.189894
R906 a_n9628_8799.n181 a_n9628_8799.n180 0.189894
R907 a_n9628_8799.n181 a_n9628_8799.n156 0.189894
R908 a_n9628_8799.n185 a_n9628_8799.n156 0.189894
R909 a_n9628_8799.n186 a_n9628_8799.n185 0.189894
R910 a_n9628_8799.n187 a_n9628_8799.n186 0.189894
R911 a_n9628_8799.n187 a_n9628_8799.n154 0.189894
R912 a_n9628_8799.n191 a_n9628_8799.n154 0.189894
R913 a_n9628_8799.n192 a_n9628_8799.n191 0.189894
R914 a_n9628_8799.n193 a_n9628_8799.n192 0.189894
R915 a_n9628_8799.n193 a_n9628_8799.n152 0.189894
R916 a_n9628_8799.n197 a_n9628_8799.n152 0.189894
R917 a_n9628_8799.n198 a_n9628_8799.n197 0.189894
R918 a_n9628_8799.n199 a_n9628_8799.n198 0.189894
R919 a_n9628_8799.n199 a_n9628_8799.n150 0.189894
R920 a_n9628_8799.n203 a_n9628_8799.n150 0.189894
R921 a_n9628_8799.n204 a_n9628_8799.n203 0.189894
R922 a_n9628_8799.n205 a_n9628_8799.n204 0.189894
R923 a_n9628_8799.n205 a_n9628_8799.n148 0.189894
R924 a_n9628_8799.n209 a_n9628_8799.n148 0.189894
R925 gnd.n7396 gnd.n535 1473.65
R926 gnd.n4148 gnd.n4147 939.716
R927 gnd.n4055 gnd.n2674 766.379
R928 gnd.n4058 gnd.n4057 766.379
R929 gnd.n3297 gnd.n3200 766.379
R930 gnd.n3293 gnd.n3198 766.379
R931 gnd.n4146 gnd.n2696 756.769
R932 gnd.n4049 gnd.n4048 756.769
R933 gnd.n3390 gnd.n3107 756.769
R934 gnd.n3388 gnd.n3110 756.769
R935 gnd.n7775 gnd.n129 751.963
R936 gnd.n7919 gnd.n7918 751.963
R937 gnd.n6053 gnd.n1681 751.963
R938 gnd.n1709 gnd.n1482 751.963
R939 gnd.n1252 gnd.n1240 751.963
R940 gnd.n4925 gnd.n4924 751.963
R941 gnd.n4400 gnd.n4150 751.963
R942 gnd.n4441 gnd.n4326 751.963
R943 gnd.n6877 gnd.n848 737.549
R944 gnd.n7397 gnd.n536 737.549
R945 gnd.n7610 gnd.n409 737.549
R946 gnd.n6709 gnd.n1018 737.549
R947 gnd.n7916 gnd.n131 732.745
R948 gnd.n199 gnd.n127 732.745
R949 gnd.n1942 gnd.n1683 732.745
R950 gnd.n6051 gnd.n1685 732.745
R951 gnd.n6578 gnd.n1245 732.745
R952 gnd.n4823 gnd.n2460 732.745
R953 gnd.n4289 gnd.n4149 732.745
R954 gnd.n4443 gnd.n2672 732.745
R955 gnd.n4971 gnd.n2332 711.122
R956 gnd.n6354 gnd.n1476 711.122
R957 gnd.n4851 gnd.n2308 711.122
R958 gnd.n6356 gnd.n1471 711.122
R959 gnd.n6878 gnd.n6877 585
R960 gnd.n6877 gnd.n6876 585
R961 gnd.n852 gnd.n851 585
R962 gnd.n6875 gnd.n852 585
R963 gnd.n6873 gnd.n6872 585
R964 gnd.n6874 gnd.n6873 585
R965 gnd.n6871 gnd.n854 585
R966 gnd.n854 gnd.n853 585
R967 gnd.n6870 gnd.n6869 585
R968 gnd.n6869 gnd.n6868 585
R969 gnd.n859 gnd.n858 585
R970 gnd.n6867 gnd.n859 585
R971 gnd.n6865 gnd.n6864 585
R972 gnd.n6866 gnd.n6865 585
R973 gnd.n6863 gnd.n861 585
R974 gnd.n861 gnd.n860 585
R975 gnd.n6862 gnd.n6861 585
R976 gnd.n6861 gnd.n6860 585
R977 gnd.n867 gnd.n866 585
R978 gnd.n6859 gnd.n867 585
R979 gnd.n6857 gnd.n6856 585
R980 gnd.n6858 gnd.n6857 585
R981 gnd.n6855 gnd.n869 585
R982 gnd.n869 gnd.n868 585
R983 gnd.n6854 gnd.n6853 585
R984 gnd.n6853 gnd.n6852 585
R985 gnd.n875 gnd.n874 585
R986 gnd.n6851 gnd.n875 585
R987 gnd.n6849 gnd.n6848 585
R988 gnd.n6850 gnd.n6849 585
R989 gnd.n6847 gnd.n877 585
R990 gnd.n877 gnd.n876 585
R991 gnd.n6846 gnd.n6845 585
R992 gnd.n6845 gnd.n6844 585
R993 gnd.n883 gnd.n882 585
R994 gnd.n6843 gnd.n883 585
R995 gnd.n6841 gnd.n6840 585
R996 gnd.n6842 gnd.n6841 585
R997 gnd.n6839 gnd.n885 585
R998 gnd.n885 gnd.n884 585
R999 gnd.n6838 gnd.n6837 585
R1000 gnd.n6837 gnd.n6836 585
R1001 gnd.n891 gnd.n890 585
R1002 gnd.n6835 gnd.n891 585
R1003 gnd.n6833 gnd.n6832 585
R1004 gnd.n6834 gnd.n6833 585
R1005 gnd.n6831 gnd.n893 585
R1006 gnd.n893 gnd.n892 585
R1007 gnd.n6830 gnd.n6829 585
R1008 gnd.n6829 gnd.n6828 585
R1009 gnd.n899 gnd.n898 585
R1010 gnd.n6827 gnd.n899 585
R1011 gnd.n6825 gnd.n6824 585
R1012 gnd.n6826 gnd.n6825 585
R1013 gnd.n6823 gnd.n901 585
R1014 gnd.n901 gnd.n900 585
R1015 gnd.n6822 gnd.n6821 585
R1016 gnd.n6821 gnd.n6820 585
R1017 gnd.n907 gnd.n906 585
R1018 gnd.n6819 gnd.n907 585
R1019 gnd.n6817 gnd.n6816 585
R1020 gnd.n6818 gnd.n6817 585
R1021 gnd.n6815 gnd.n909 585
R1022 gnd.n909 gnd.n908 585
R1023 gnd.n6814 gnd.n6813 585
R1024 gnd.n6813 gnd.n6812 585
R1025 gnd.n915 gnd.n914 585
R1026 gnd.n6811 gnd.n915 585
R1027 gnd.n6809 gnd.n6808 585
R1028 gnd.n6810 gnd.n6809 585
R1029 gnd.n6807 gnd.n917 585
R1030 gnd.n917 gnd.n916 585
R1031 gnd.n6806 gnd.n6805 585
R1032 gnd.n6805 gnd.n6804 585
R1033 gnd.n923 gnd.n922 585
R1034 gnd.n6803 gnd.n923 585
R1035 gnd.n6801 gnd.n6800 585
R1036 gnd.n6802 gnd.n6801 585
R1037 gnd.n6799 gnd.n925 585
R1038 gnd.n925 gnd.n924 585
R1039 gnd.n6798 gnd.n6797 585
R1040 gnd.n6797 gnd.n6796 585
R1041 gnd.n931 gnd.n930 585
R1042 gnd.n6795 gnd.n931 585
R1043 gnd.n6793 gnd.n6792 585
R1044 gnd.n6794 gnd.n6793 585
R1045 gnd.n6791 gnd.n933 585
R1046 gnd.n933 gnd.n932 585
R1047 gnd.n6790 gnd.n6789 585
R1048 gnd.n6789 gnd.n6788 585
R1049 gnd.n939 gnd.n938 585
R1050 gnd.n6787 gnd.n939 585
R1051 gnd.n6785 gnd.n6784 585
R1052 gnd.n6786 gnd.n6785 585
R1053 gnd.n6783 gnd.n941 585
R1054 gnd.n941 gnd.n940 585
R1055 gnd.n6782 gnd.n6781 585
R1056 gnd.n6781 gnd.n6780 585
R1057 gnd.n947 gnd.n946 585
R1058 gnd.n6779 gnd.n947 585
R1059 gnd.n6777 gnd.n6776 585
R1060 gnd.n6778 gnd.n6777 585
R1061 gnd.n6775 gnd.n949 585
R1062 gnd.n949 gnd.n948 585
R1063 gnd.n6774 gnd.n6773 585
R1064 gnd.n6773 gnd.n6772 585
R1065 gnd.n955 gnd.n954 585
R1066 gnd.n6771 gnd.n955 585
R1067 gnd.n6769 gnd.n6768 585
R1068 gnd.n6770 gnd.n6769 585
R1069 gnd.n6767 gnd.n957 585
R1070 gnd.n957 gnd.n956 585
R1071 gnd.n6766 gnd.n6765 585
R1072 gnd.n6765 gnd.n6764 585
R1073 gnd.n963 gnd.n962 585
R1074 gnd.n6763 gnd.n963 585
R1075 gnd.n6761 gnd.n6760 585
R1076 gnd.n6762 gnd.n6761 585
R1077 gnd.n6759 gnd.n965 585
R1078 gnd.n965 gnd.n964 585
R1079 gnd.n6758 gnd.n6757 585
R1080 gnd.n6757 gnd.n6756 585
R1081 gnd.n971 gnd.n970 585
R1082 gnd.n6755 gnd.n971 585
R1083 gnd.n6753 gnd.n6752 585
R1084 gnd.n6754 gnd.n6753 585
R1085 gnd.n6751 gnd.n973 585
R1086 gnd.n973 gnd.n972 585
R1087 gnd.n6750 gnd.n6749 585
R1088 gnd.n6749 gnd.n6748 585
R1089 gnd.n979 gnd.n978 585
R1090 gnd.n6747 gnd.n979 585
R1091 gnd.n6745 gnd.n6744 585
R1092 gnd.n6746 gnd.n6745 585
R1093 gnd.n6743 gnd.n981 585
R1094 gnd.n981 gnd.n980 585
R1095 gnd.n6742 gnd.n6741 585
R1096 gnd.n6741 gnd.n6740 585
R1097 gnd.n987 gnd.n986 585
R1098 gnd.n6739 gnd.n987 585
R1099 gnd.n6737 gnd.n6736 585
R1100 gnd.n6738 gnd.n6737 585
R1101 gnd.n6735 gnd.n989 585
R1102 gnd.n989 gnd.n988 585
R1103 gnd.n6734 gnd.n6733 585
R1104 gnd.n6733 gnd.n6732 585
R1105 gnd.n995 gnd.n994 585
R1106 gnd.n6731 gnd.n995 585
R1107 gnd.n6729 gnd.n6728 585
R1108 gnd.n6730 gnd.n6729 585
R1109 gnd.n6727 gnd.n997 585
R1110 gnd.n997 gnd.n996 585
R1111 gnd.n6726 gnd.n6725 585
R1112 gnd.n6725 gnd.n6724 585
R1113 gnd.n1003 gnd.n1002 585
R1114 gnd.n6723 gnd.n1003 585
R1115 gnd.n6721 gnd.n6720 585
R1116 gnd.n6722 gnd.n6721 585
R1117 gnd.n6719 gnd.n1005 585
R1118 gnd.n1005 gnd.n1004 585
R1119 gnd.n6718 gnd.n6717 585
R1120 gnd.n6717 gnd.n6716 585
R1121 gnd.n1011 gnd.n1010 585
R1122 gnd.n6715 gnd.n1011 585
R1123 gnd.n6713 gnd.n6712 585
R1124 gnd.n6714 gnd.n6713 585
R1125 gnd.n6711 gnd.n1013 585
R1126 gnd.n1013 gnd.n1012 585
R1127 gnd.n849 gnd.n848 585
R1128 gnd.n848 gnd.n847 585
R1129 gnd.n6883 gnd.n6882 585
R1130 gnd.n6884 gnd.n6883 585
R1131 gnd.n846 gnd.n845 585
R1132 gnd.n6885 gnd.n846 585
R1133 gnd.n6888 gnd.n6887 585
R1134 gnd.n6887 gnd.n6886 585
R1135 gnd.n843 gnd.n842 585
R1136 gnd.n842 gnd.n841 585
R1137 gnd.n6893 gnd.n6892 585
R1138 gnd.n6894 gnd.n6893 585
R1139 gnd.n840 gnd.n839 585
R1140 gnd.n6895 gnd.n840 585
R1141 gnd.n6898 gnd.n6897 585
R1142 gnd.n6897 gnd.n6896 585
R1143 gnd.n837 gnd.n836 585
R1144 gnd.n836 gnd.n835 585
R1145 gnd.n6903 gnd.n6902 585
R1146 gnd.n6904 gnd.n6903 585
R1147 gnd.n834 gnd.n833 585
R1148 gnd.n6905 gnd.n834 585
R1149 gnd.n6908 gnd.n6907 585
R1150 gnd.n6907 gnd.n6906 585
R1151 gnd.n831 gnd.n830 585
R1152 gnd.n830 gnd.n829 585
R1153 gnd.n6913 gnd.n6912 585
R1154 gnd.n6914 gnd.n6913 585
R1155 gnd.n828 gnd.n827 585
R1156 gnd.n6915 gnd.n828 585
R1157 gnd.n6918 gnd.n6917 585
R1158 gnd.n6917 gnd.n6916 585
R1159 gnd.n825 gnd.n824 585
R1160 gnd.n824 gnd.n823 585
R1161 gnd.n6923 gnd.n6922 585
R1162 gnd.n6924 gnd.n6923 585
R1163 gnd.n822 gnd.n821 585
R1164 gnd.n6925 gnd.n822 585
R1165 gnd.n6928 gnd.n6927 585
R1166 gnd.n6927 gnd.n6926 585
R1167 gnd.n819 gnd.n818 585
R1168 gnd.n818 gnd.n817 585
R1169 gnd.n6933 gnd.n6932 585
R1170 gnd.n6934 gnd.n6933 585
R1171 gnd.n816 gnd.n815 585
R1172 gnd.n6935 gnd.n816 585
R1173 gnd.n6938 gnd.n6937 585
R1174 gnd.n6937 gnd.n6936 585
R1175 gnd.n813 gnd.n812 585
R1176 gnd.n812 gnd.n811 585
R1177 gnd.n6943 gnd.n6942 585
R1178 gnd.n6944 gnd.n6943 585
R1179 gnd.n810 gnd.n809 585
R1180 gnd.n6945 gnd.n810 585
R1181 gnd.n6948 gnd.n6947 585
R1182 gnd.n6947 gnd.n6946 585
R1183 gnd.n807 gnd.n806 585
R1184 gnd.n806 gnd.n805 585
R1185 gnd.n6953 gnd.n6952 585
R1186 gnd.n6954 gnd.n6953 585
R1187 gnd.n804 gnd.n803 585
R1188 gnd.n6955 gnd.n804 585
R1189 gnd.n6958 gnd.n6957 585
R1190 gnd.n6957 gnd.n6956 585
R1191 gnd.n801 gnd.n800 585
R1192 gnd.n800 gnd.n799 585
R1193 gnd.n6963 gnd.n6962 585
R1194 gnd.n6964 gnd.n6963 585
R1195 gnd.n798 gnd.n797 585
R1196 gnd.n6965 gnd.n798 585
R1197 gnd.n6968 gnd.n6967 585
R1198 gnd.n6967 gnd.n6966 585
R1199 gnd.n795 gnd.n794 585
R1200 gnd.n794 gnd.n793 585
R1201 gnd.n6973 gnd.n6972 585
R1202 gnd.n6974 gnd.n6973 585
R1203 gnd.n792 gnd.n791 585
R1204 gnd.n6975 gnd.n792 585
R1205 gnd.n6978 gnd.n6977 585
R1206 gnd.n6977 gnd.n6976 585
R1207 gnd.n789 gnd.n788 585
R1208 gnd.n788 gnd.n787 585
R1209 gnd.n6983 gnd.n6982 585
R1210 gnd.n6984 gnd.n6983 585
R1211 gnd.n786 gnd.n785 585
R1212 gnd.n6985 gnd.n786 585
R1213 gnd.n6988 gnd.n6987 585
R1214 gnd.n6987 gnd.n6986 585
R1215 gnd.n783 gnd.n782 585
R1216 gnd.n782 gnd.n781 585
R1217 gnd.n6993 gnd.n6992 585
R1218 gnd.n6994 gnd.n6993 585
R1219 gnd.n780 gnd.n779 585
R1220 gnd.n6995 gnd.n780 585
R1221 gnd.n6998 gnd.n6997 585
R1222 gnd.n6997 gnd.n6996 585
R1223 gnd.n777 gnd.n776 585
R1224 gnd.n776 gnd.n775 585
R1225 gnd.n7003 gnd.n7002 585
R1226 gnd.n7004 gnd.n7003 585
R1227 gnd.n774 gnd.n773 585
R1228 gnd.n7005 gnd.n774 585
R1229 gnd.n7008 gnd.n7007 585
R1230 gnd.n7007 gnd.n7006 585
R1231 gnd.n771 gnd.n770 585
R1232 gnd.n770 gnd.n769 585
R1233 gnd.n7013 gnd.n7012 585
R1234 gnd.n7014 gnd.n7013 585
R1235 gnd.n768 gnd.n767 585
R1236 gnd.n7015 gnd.n768 585
R1237 gnd.n7018 gnd.n7017 585
R1238 gnd.n7017 gnd.n7016 585
R1239 gnd.n765 gnd.n764 585
R1240 gnd.n764 gnd.n763 585
R1241 gnd.n7023 gnd.n7022 585
R1242 gnd.n7024 gnd.n7023 585
R1243 gnd.n762 gnd.n761 585
R1244 gnd.n7025 gnd.n762 585
R1245 gnd.n7028 gnd.n7027 585
R1246 gnd.n7027 gnd.n7026 585
R1247 gnd.n759 gnd.n758 585
R1248 gnd.n758 gnd.n757 585
R1249 gnd.n7033 gnd.n7032 585
R1250 gnd.n7034 gnd.n7033 585
R1251 gnd.n756 gnd.n755 585
R1252 gnd.n7035 gnd.n756 585
R1253 gnd.n7038 gnd.n7037 585
R1254 gnd.n7037 gnd.n7036 585
R1255 gnd.n753 gnd.n752 585
R1256 gnd.n752 gnd.n751 585
R1257 gnd.n7043 gnd.n7042 585
R1258 gnd.n7044 gnd.n7043 585
R1259 gnd.n750 gnd.n749 585
R1260 gnd.n7045 gnd.n750 585
R1261 gnd.n7048 gnd.n7047 585
R1262 gnd.n7047 gnd.n7046 585
R1263 gnd.n747 gnd.n746 585
R1264 gnd.n746 gnd.n745 585
R1265 gnd.n7053 gnd.n7052 585
R1266 gnd.n7054 gnd.n7053 585
R1267 gnd.n744 gnd.n743 585
R1268 gnd.n7055 gnd.n744 585
R1269 gnd.n7058 gnd.n7057 585
R1270 gnd.n7057 gnd.n7056 585
R1271 gnd.n741 gnd.n740 585
R1272 gnd.n740 gnd.n739 585
R1273 gnd.n7063 gnd.n7062 585
R1274 gnd.n7064 gnd.n7063 585
R1275 gnd.n738 gnd.n737 585
R1276 gnd.n7065 gnd.n738 585
R1277 gnd.n7068 gnd.n7067 585
R1278 gnd.n7067 gnd.n7066 585
R1279 gnd.n735 gnd.n734 585
R1280 gnd.n734 gnd.n733 585
R1281 gnd.n7073 gnd.n7072 585
R1282 gnd.n7074 gnd.n7073 585
R1283 gnd.n732 gnd.n731 585
R1284 gnd.n7075 gnd.n732 585
R1285 gnd.n7078 gnd.n7077 585
R1286 gnd.n7077 gnd.n7076 585
R1287 gnd.n729 gnd.n728 585
R1288 gnd.n728 gnd.n727 585
R1289 gnd.n7083 gnd.n7082 585
R1290 gnd.n7084 gnd.n7083 585
R1291 gnd.n726 gnd.n725 585
R1292 gnd.n7085 gnd.n726 585
R1293 gnd.n7088 gnd.n7087 585
R1294 gnd.n7087 gnd.n7086 585
R1295 gnd.n723 gnd.n722 585
R1296 gnd.n722 gnd.n721 585
R1297 gnd.n7093 gnd.n7092 585
R1298 gnd.n7094 gnd.n7093 585
R1299 gnd.n720 gnd.n719 585
R1300 gnd.n7095 gnd.n720 585
R1301 gnd.n7098 gnd.n7097 585
R1302 gnd.n7097 gnd.n7096 585
R1303 gnd.n717 gnd.n716 585
R1304 gnd.n716 gnd.n715 585
R1305 gnd.n7103 gnd.n7102 585
R1306 gnd.n7104 gnd.n7103 585
R1307 gnd.n714 gnd.n713 585
R1308 gnd.n7105 gnd.n714 585
R1309 gnd.n7108 gnd.n7107 585
R1310 gnd.n7107 gnd.n7106 585
R1311 gnd.n711 gnd.n710 585
R1312 gnd.n710 gnd.n709 585
R1313 gnd.n7113 gnd.n7112 585
R1314 gnd.n7114 gnd.n7113 585
R1315 gnd.n708 gnd.n707 585
R1316 gnd.n7115 gnd.n708 585
R1317 gnd.n7118 gnd.n7117 585
R1318 gnd.n7117 gnd.n7116 585
R1319 gnd.n705 gnd.n704 585
R1320 gnd.n704 gnd.n703 585
R1321 gnd.n7123 gnd.n7122 585
R1322 gnd.n7124 gnd.n7123 585
R1323 gnd.n702 gnd.n701 585
R1324 gnd.n7125 gnd.n702 585
R1325 gnd.n7128 gnd.n7127 585
R1326 gnd.n7127 gnd.n7126 585
R1327 gnd.n699 gnd.n698 585
R1328 gnd.n698 gnd.n697 585
R1329 gnd.n7133 gnd.n7132 585
R1330 gnd.n7134 gnd.n7133 585
R1331 gnd.n696 gnd.n695 585
R1332 gnd.n7135 gnd.n696 585
R1333 gnd.n7138 gnd.n7137 585
R1334 gnd.n7137 gnd.n7136 585
R1335 gnd.n693 gnd.n692 585
R1336 gnd.n692 gnd.n691 585
R1337 gnd.n7143 gnd.n7142 585
R1338 gnd.n7144 gnd.n7143 585
R1339 gnd.n690 gnd.n689 585
R1340 gnd.n7145 gnd.n690 585
R1341 gnd.n7148 gnd.n7147 585
R1342 gnd.n7147 gnd.n7146 585
R1343 gnd.n687 gnd.n686 585
R1344 gnd.n686 gnd.n685 585
R1345 gnd.n7153 gnd.n7152 585
R1346 gnd.n7154 gnd.n7153 585
R1347 gnd.n684 gnd.n683 585
R1348 gnd.n7155 gnd.n684 585
R1349 gnd.n7158 gnd.n7157 585
R1350 gnd.n7157 gnd.n7156 585
R1351 gnd.n681 gnd.n680 585
R1352 gnd.n680 gnd.n679 585
R1353 gnd.n7163 gnd.n7162 585
R1354 gnd.n7164 gnd.n7163 585
R1355 gnd.n678 gnd.n677 585
R1356 gnd.n7165 gnd.n678 585
R1357 gnd.n7168 gnd.n7167 585
R1358 gnd.n7167 gnd.n7166 585
R1359 gnd.n675 gnd.n674 585
R1360 gnd.n674 gnd.n673 585
R1361 gnd.n7173 gnd.n7172 585
R1362 gnd.n7174 gnd.n7173 585
R1363 gnd.n672 gnd.n671 585
R1364 gnd.n7175 gnd.n672 585
R1365 gnd.n7178 gnd.n7177 585
R1366 gnd.n7177 gnd.n7176 585
R1367 gnd.n669 gnd.n668 585
R1368 gnd.n668 gnd.n667 585
R1369 gnd.n7183 gnd.n7182 585
R1370 gnd.n7184 gnd.n7183 585
R1371 gnd.n666 gnd.n665 585
R1372 gnd.n7185 gnd.n666 585
R1373 gnd.n7188 gnd.n7187 585
R1374 gnd.n7187 gnd.n7186 585
R1375 gnd.n663 gnd.n662 585
R1376 gnd.n662 gnd.n661 585
R1377 gnd.n7193 gnd.n7192 585
R1378 gnd.n7194 gnd.n7193 585
R1379 gnd.n660 gnd.n659 585
R1380 gnd.n7195 gnd.n660 585
R1381 gnd.n7198 gnd.n7197 585
R1382 gnd.n7197 gnd.n7196 585
R1383 gnd.n657 gnd.n656 585
R1384 gnd.n656 gnd.n655 585
R1385 gnd.n7203 gnd.n7202 585
R1386 gnd.n7204 gnd.n7203 585
R1387 gnd.n654 gnd.n653 585
R1388 gnd.n7205 gnd.n654 585
R1389 gnd.n7208 gnd.n7207 585
R1390 gnd.n7207 gnd.n7206 585
R1391 gnd.n651 gnd.n650 585
R1392 gnd.n650 gnd.n649 585
R1393 gnd.n7213 gnd.n7212 585
R1394 gnd.n7214 gnd.n7213 585
R1395 gnd.n648 gnd.n647 585
R1396 gnd.n7215 gnd.n648 585
R1397 gnd.n7218 gnd.n7217 585
R1398 gnd.n7217 gnd.n7216 585
R1399 gnd.n645 gnd.n644 585
R1400 gnd.n644 gnd.n643 585
R1401 gnd.n7223 gnd.n7222 585
R1402 gnd.n7224 gnd.n7223 585
R1403 gnd.n642 gnd.n641 585
R1404 gnd.n7225 gnd.n642 585
R1405 gnd.n7228 gnd.n7227 585
R1406 gnd.n7227 gnd.n7226 585
R1407 gnd.n639 gnd.n638 585
R1408 gnd.n638 gnd.n637 585
R1409 gnd.n7233 gnd.n7232 585
R1410 gnd.n7234 gnd.n7233 585
R1411 gnd.n636 gnd.n635 585
R1412 gnd.n7235 gnd.n636 585
R1413 gnd.n7238 gnd.n7237 585
R1414 gnd.n7237 gnd.n7236 585
R1415 gnd.n633 gnd.n632 585
R1416 gnd.n632 gnd.n631 585
R1417 gnd.n7243 gnd.n7242 585
R1418 gnd.n7244 gnd.n7243 585
R1419 gnd.n630 gnd.n629 585
R1420 gnd.n7245 gnd.n630 585
R1421 gnd.n7248 gnd.n7247 585
R1422 gnd.n7247 gnd.n7246 585
R1423 gnd.n627 gnd.n626 585
R1424 gnd.n626 gnd.n625 585
R1425 gnd.n7253 gnd.n7252 585
R1426 gnd.n7254 gnd.n7253 585
R1427 gnd.n624 gnd.n623 585
R1428 gnd.n7255 gnd.n624 585
R1429 gnd.n7258 gnd.n7257 585
R1430 gnd.n7257 gnd.n7256 585
R1431 gnd.n621 gnd.n620 585
R1432 gnd.n620 gnd.n619 585
R1433 gnd.n7263 gnd.n7262 585
R1434 gnd.n7264 gnd.n7263 585
R1435 gnd.n618 gnd.n617 585
R1436 gnd.n7265 gnd.n618 585
R1437 gnd.n7268 gnd.n7267 585
R1438 gnd.n7267 gnd.n7266 585
R1439 gnd.n615 gnd.n614 585
R1440 gnd.n614 gnd.n613 585
R1441 gnd.n7273 gnd.n7272 585
R1442 gnd.n7274 gnd.n7273 585
R1443 gnd.n612 gnd.n611 585
R1444 gnd.n7275 gnd.n612 585
R1445 gnd.n7278 gnd.n7277 585
R1446 gnd.n7277 gnd.n7276 585
R1447 gnd.n609 gnd.n608 585
R1448 gnd.n608 gnd.n607 585
R1449 gnd.n7283 gnd.n7282 585
R1450 gnd.n7284 gnd.n7283 585
R1451 gnd.n606 gnd.n605 585
R1452 gnd.n7285 gnd.n606 585
R1453 gnd.n7288 gnd.n7287 585
R1454 gnd.n7287 gnd.n7286 585
R1455 gnd.n603 gnd.n602 585
R1456 gnd.n602 gnd.n601 585
R1457 gnd.n7293 gnd.n7292 585
R1458 gnd.n7294 gnd.n7293 585
R1459 gnd.n600 gnd.n599 585
R1460 gnd.n7295 gnd.n600 585
R1461 gnd.n7298 gnd.n7297 585
R1462 gnd.n7297 gnd.n7296 585
R1463 gnd.n597 gnd.n596 585
R1464 gnd.n596 gnd.n595 585
R1465 gnd.n7303 gnd.n7302 585
R1466 gnd.n7304 gnd.n7303 585
R1467 gnd.n594 gnd.n593 585
R1468 gnd.n7305 gnd.n594 585
R1469 gnd.n7308 gnd.n7307 585
R1470 gnd.n7307 gnd.n7306 585
R1471 gnd.n591 gnd.n590 585
R1472 gnd.n590 gnd.n589 585
R1473 gnd.n7313 gnd.n7312 585
R1474 gnd.n7314 gnd.n7313 585
R1475 gnd.n588 gnd.n587 585
R1476 gnd.n7315 gnd.n588 585
R1477 gnd.n7318 gnd.n7317 585
R1478 gnd.n7317 gnd.n7316 585
R1479 gnd.n585 gnd.n584 585
R1480 gnd.n584 gnd.n583 585
R1481 gnd.n7323 gnd.n7322 585
R1482 gnd.n7324 gnd.n7323 585
R1483 gnd.n582 gnd.n581 585
R1484 gnd.n7325 gnd.n582 585
R1485 gnd.n7328 gnd.n7327 585
R1486 gnd.n7327 gnd.n7326 585
R1487 gnd.n579 gnd.n578 585
R1488 gnd.n578 gnd.n577 585
R1489 gnd.n7333 gnd.n7332 585
R1490 gnd.n7334 gnd.n7333 585
R1491 gnd.n576 gnd.n575 585
R1492 gnd.n7335 gnd.n576 585
R1493 gnd.n7338 gnd.n7337 585
R1494 gnd.n7337 gnd.n7336 585
R1495 gnd.n573 gnd.n572 585
R1496 gnd.n572 gnd.n571 585
R1497 gnd.n7343 gnd.n7342 585
R1498 gnd.n7344 gnd.n7343 585
R1499 gnd.n570 gnd.n569 585
R1500 gnd.n7345 gnd.n570 585
R1501 gnd.n7348 gnd.n7347 585
R1502 gnd.n7347 gnd.n7346 585
R1503 gnd.n567 gnd.n566 585
R1504 gnd.n566 gnd.n565 585
R1505 gnd.n7353 gnd.n7352 585
R1506 gnd.n7354 gnd.n7353 585
R1507 gnd.n564 gnd.n563 585
R1508 gnd.n7355 gnd.n564 585
R1509 gnd.n7358 gnd.n7357 585
R1510 gnd.n7357 gnd.n7356 585
R1511 gnd.n561 gnd.n560 585
R1512 gnd.n560 gnd.n559 585
R1513 gnd.n7363 gnd.n7362 585
R1514 gnd.n7364 gnd.n7363 585
R1515 gnd.n558 gnd.n557 585
R1516 gnd.n7365 gnd.n558 585
R1517 gnd.n7368 gnd.n7367 585
R1518 gnd.n7367 gnd.n7366 585
R1519 gnd.n555 gnd.n554 585
R1520 gnd.n554 gnd.n553 585
R1521 gnd.n7373 gnd.n7372 585
R1522 gnd.n7374 gnd.n7373 585
R1523 gnd.n552 gnd.n551 585
R1524 gnd.n7375 gnd.n552 585
R1525 gnd.n7378 gnd.n7377 585
R1526 gnd.n7377 gnd.n7376 585
R1527 gnd.n549 gnd.n548 585
R1528 gnd.n548 gnd.n547 585
R1529 gnd.n7383 gnd.n7382 585
R1530 gnd.n7384 gnd.n7383 585
R1531 gnd.n546 gnd.n545 585
R1532 gnd.n7385 gnd.n546 585
R1533 gnd.n7388 gnd.n7387 585
R1534 gnd.n7387 gnd.n7386 585
R1535 gnd.n543 gnd.n542 585
R1536 gnd.n542 gnd.n541 585
R1537 gnd.n7393 gnd.n7392 585
R1538 gnd.n7394 gnd.n7393 585
R1539 gnd.n540 gnd.n539 585
R1540 gnd.n7395 gnd.n540 585
R1541 gnd.n7398 gnd.n7397 585
R1542 gnd.n7397 gnd.n7396 585
R1543 gnd.n7609 gnd.n413 585
R1544 gnd.n7609 gnd.n7608 585
R1545 gnd.n7603 gnd.n414 585
R1546 gnd.n7607 gnd.n414 585
R1547 gnd.n7605 gnd.n7604 585
R1548 gnd.n7606 gnd.n7605 585
R1549 gnd.n417 gnd.n416 585
R1550 gnd.n416 gnd.n415 585
R1551 gnd.n7598 gnd.n7597 585
R1552 gnd.n7597 gnd.n7596 585
R1553 gnd.n420 gnd.n419 585
R1554 gnd.n7595 gnd.n420 585
R1555 gnd.n7593 gnd.n7592 585
R1556 gnd.n7594 gnd.n7593 585
R1557 gnd.n423 gnd.n422 585
R1558 gnd.n422 gnd.n421 585
R1559 gnd.n7588 gnd.n7587 585
R1560 gnd.n7587 gnd.n7586 585
R1561 gnd.n426 gnd.n425 585
R1562 gnd.n7585 gnd.n426 585
R1563 gnd.n7583 gnd.n7582 585
R1564 gnd.n7584 gnd.n7583 585
R1565 gnd.n429 gnd.n428 585
R1566 gnd.n428 gnd.n427 585
R1567 gnd.n7578 gnd.n7577 585
R1568 gnd.n7577 gnd.n7576 585
R1569 gnd.n432 gnd.n431 585
R1570 gnd.n7575 gnd.n432 585
R1571 gnd.n7573 gnd.n7572 585
R1572 gnd.n7574 gnd.n7573 585
R1573 gnd.n435 gnd.n434 585
R1574 gnd.n434 gnd.n433 585
R1575 gnd.n7568 gnd.n7567 585
R1576 gnd.n7567 gnd.n7566 585
R1577 gnd.n438 gnd.n437 585
R1578 gnd.n7565 gnd.n438 585
R1579 gnd.n7563 gnd.n7562 585
R1580 gnd.n7564 gnd.n7563 585
R1581 gnd.n441 gnd.n440 585
R1582 gnd.n440 gnd.n439 585
R1583 gnd.n7558 gnd.n7557 585
R1584 gnd.n7557 gnd.n7556 585
R1585 gnd.n444 gnd.n443 585
R1586 gnd.n7555 gnd.n444 585
R1587 gnd.n7553 gnd.n7552 585
R1588 gnd.n7554 gnd.n7553 585
R1589 gnd.n447 gnd.n446 585
R1590 gnd.n446 gnd.n445 585
R1591 gnd.n7548 gnd.n7547 585
R1592 gnd.n7547 gnd.n7546 585
R1593 gnd.n450 gnd.n449 585
R1594 gnd.n7545 gnd.n450 585
R1595 gnd.n7543 gnd.n7542 585
R1596 gnd.n7544 gnd.n7543 585
R1597 gnd.n453 gnd.n452 585
R1598 gnd.n452 gnd.n451 585
R1599 gnd.n7538 gnd.n7537 585
R1600 gnd.n7537 gnd.n7536 585
R1601 gnd.n456 gnd.n455 585
R1602 gnd.n7535 gnd.n456 585
R1603 gnd.n7533 gnd.n7532 585
R1604 gnd.n7534 gnd.n7533 585
R1605 gnd.n459 gnd.n458 585
R1606 gnd.n458 gnd.n457 585
R1607 gnd.n7528 gnd.n7527 585
R1608 gnd.n7527 gnd.n7526 585
R1609 gnd.n462 gnd.n461 585
R1610 gnd.n7525 gnd.n462 585
R1611 gnd.n7523 gnd.n7522 585
R1612 gnd.n7524 gnd.n7523 585
R1613 gnd.n465 gnd.n464 585
R1614 gnd.n464 gnd.n463 585
R1615 gnd.n7518 gnd.n7517 585
R1616 gnd.n7517 gnd.n7516 585
R1617 gnd.n468 gnd.n467 585
R1618 gnd.n7515 gnd.n468 585
R1619 gnd.n7513 gnd.n7512 585
R1620 gnd.n7514 gnd.n7513 585
R1621 gnd.n471 gnd.n470 585
R1622 gnd.n470 gnd.n469 585
R1623 gnd.n7508 gnd.n7507 585
R1624 gnd.n7507 gnd.n7506 585
R1625 gnd.n474 gnd.n473 585
R1626 gnd.n7505 gnd.n474 585
R1627 gnd.n7503 gnd.n7502 585
R1628 gnd.n7504 gnd.n7503 585
R1629 gnd.n477 gnd.n476 585
R1630 gnd.n476 gnd.n475 585
R1631 gnd.n7498 gnd.n7497 585
R1632 gnd.n7497 gnd.n7496 585
R1633 gnd.n480 gnd.n479 585
R1634 gnd.n7495 gnd.n480 585
R1635 gnd.n7493 gnd.n7492 585
R1636 gnd.n7494 gnd.n7493 585
R1637 gnd.n483 gnd.n482 585
R1638 gnd.n482 gnd.n481 585
R1639 gnd.n7488 gnd.n7487 585
R1640 gnd.n7487 gnd.n7486 585
R1641 gnd.n486 gnd.n485 585
R1642 gnd.n7485 gnd.n486 585
R1643 gnd.n7483 gnd.n7482 585
R1644 gnd.n7484 gnd.n7483 585
R1645 gnd.n489 gnd.n488 585
R1646 gnd.n488 gnd.n487 585
R1647 gnd.n7478 gnd.n7477 585
R1648 gnd.n7477 gnd.n7476 585
R1649 gnd.n492 gnd.n491 585
R1650 gnd.n7475 gnd.n492 585
R1651 gnd.n7473 gnd.n7472 585
R1652 gnd.n7474 gnd.n7473 585
R1653 gnd.n495 gnd.n494 585
R1654 gnd.n494 gnd.n493 585
R1655 gnd.n7468 gnd.n7467 585
R1656 gnd.n7467 gnd.n7466 585
R1657 gnd.n498 gnd.n497 585
R1658 gnd.n7465 gnd.n498 585
R1659 gnd.n7463 gnd.n7462 585
R1660 gnd.n7464 gnd.n7463 585
R1661 gnd.n501 gnd.n500 585
R1662 gnd.n500 gnd.n499 585
R1663 gnd.n7458 gnd.n7457 585
R1664 gnd.n7457 gnd.n7456 585
R1665 gnd.n504 gnd.n503 585
R1666 gnd.n7455 gnd.n504 585
R1667 gnd.n7453 gnd.n7452 585
R1668 gnd.n7454 gnd.n7453 585
R1669 gnd.n507 gnd.n506 585
R1670 gnd.n506 gnd.n505 585
R1671 gnd.n7448 gnd.n7447 585
R1672 gnd.n7447 gnd.n7446 585
R1673 gnd.n510 gnd.n509 585
R1674 gnd.n7445 gnd.n510 585
R1675 gnd.n7443 gnd.n7442 585
R1676 gnd.n7444 gnd.n7443 585
R1677 gnd.n513 gnd.n512 585
R1678 gnd.n512 gnd.n511 585
R1679 gnd.n7438 gnd.n7437 585
R1680 gnd.n7437 gnd.n7436 585
R1681 gnd.n516 gnd.n515 585
R1682 gnd.n7435 gnd.n516 585
R1683 gnd.n7433 gnd.n7432 585
R1684 gnd.n7434 gnd.n7433 585
R1685 gnd.n519 gnd.n518 585
R1686 gnd.n518 gnd.n517 585
R1687 gnd.n7428 gnd.n7427 585
R1688 gnd.n7427 gnd.n7426 585
R1689 gnd.n522 gnd.n521 585
R1690 gnd.n7425 gnd.n522 585
R1691 gnd.n7423 gnd.n7422 585
R1692 gnd.n7424 gnd.n7423 585
R1693 gnd.n525 gnd.n524 585
R1694 gnd.n524 gnd.n523 585
R1695 gnd.n7418 gnd.n7417 585
R1696 gnd.n7417 gnd.n7416 585
R1697 gnd.n528 gnd.n527 585
R1698 gnd.n7415 gnd.n528 585
R1699 gnd.n7413 gnd.n7412 585
R1700 gnd.n7414 gnd.n7413 585
R1701 gnd.n531 gnd.n530 585
R1702 gnd.n530 gnd.n529 585
R1703 gnd.n7408 gnd.n7407 585
R1704 gnd.n7407 gnd.n7406 585
R1705 gnd.n534 gnd.n533 585
R1706 gnd.n7405 gnd.n534 585
R1707 gnd.n7403 gnd.n7402 585
R1708 gnd.n7404 gnd.n7403 585
R1709 gnd.n537 gnd.n536 585
R1710 gnd.n536 gnd.n535 585
R1711 gnd.n1240 gnd.n1239 585
R1712 gnd.n4923 gnd.n1240 585
R1713 gnd.n6587 gnd.n6586 585
R1714 gnd.n6586 gnd.n6585 585
R1715 gnd.n6588 gnd.n1234 585
R1716 gnd.n4831 gnd.n1234 585
R1717 gnd.n6590 gnd.n6589 585
R1718 gnd.n6591 gnd.n6590 585
R1719 gnd.n1218 gnd.n1217 585
R1720 gnd.n4755 gnd.n1218 585
R1721 gnd.n6599 gnd.n6598 585
R1722 gnd.n6598 gnd.n6597 585
R1723 gnd.n6600 gnd.n1212 585
R1724 gnd.n4751 gnd.n1212 585
R1725 gnd.n6602 gnd.n6601 585
R1726 gnd.n6603 gnd.n6602 585
R1727 gnd.n1197 gnd.n1196 585
R1728 gnd.n4745 gnd.n1197 585
R1729 gnd.n6611 gnd.n6610 585
R1730 gnd.n6610 gnd.n6609 585
R1731 gnd.n6612 gnd.n1191 585
R1732 gnd.n4888 gnd.n1191 585
R1733 gnd.n6614 gnd.n6613 585
R1734 gnd.n6615 gnd.n6614 585
R1735 gnd.n1175 gnd.n1174 585
R1736 gnd.n4737 gnd.n1175 585
R1737 gnd.n6623 gnd.n6622 585
R1738 gnd.n6622 gnd.n6621 585
R1739 gnd.n6624 gnd.n1169 585
R1740 gnd.n4729 gnd.n1169 585
R1741 gnd.n6626 gnd.n6625 585
R1742 gnd.n6627 gnd.n6626 585
R1743 gnd.n1154 gnd.n1153 585
R1744 gnd.n4721 gnd.n1154 585
R1745 gnd.n6635 gnd.n6634 585
R1746 gnd.n6634 gnd.n6633 585
R1747 gnd.n6636 gnd.n1148 585
R1748 gnd.n4713 gnd.n1148 585
R1749 gnd.n6638 gnd.n6637 585
R1750 gnd.n6639 gnd.n6638 585
R1751 gnd.n1132 gnd.n1131 585
R1752 gnd.n4662 gnd.n1132 585
R1753 gnd.n6647 gnd.n6646 585
R1754 gnd.n6646 gnd.n6645 585
R1755 gnd.n6648 gnd.n1126 585
R1756 gnd.n4650 gnd.n1126 585
R1757 gnd.n6650 gnd.n6649 585
R1758 gnd.n6651 gnd.n6650 585
R1759 gnd.n1112 gnd.n1111 585
R1760 gnd.n4646 gnd.n1112 585
R1761 gnd.n6659 gnd.n6658 585
R1762 gnd.n6658 gnd.n6657 585
R1763 gnd.n6660 gnd.n1106 585
R1764 gnd.n4676 gnd.n1106 585
R1765 gnd.n6662 gnd.n6661 585
R1766 gnd.n6663 gnd.n6662 585
R1767 gnd.n1107 gnd.n1105 585
R1768 gnd.n4638 gnd.n1105 585
R1769 gnd.n4624 gnd.n4623 585
R1770 gnd.n4625 gnd.n4624 585
R1771 gnd.n2538 gnd.n2535 585
R1772 gnd.n4630 gnd.n2535 585
R1773 gnd.n4618 gnd.n4617 585
R1774 gnd.n4617 gnd.n4616 585
R1775 gnd.n2541 gnd.n2540 585
R1776 gnd.n4597 gnd.n2541 585
R1777 gnd.n4587 gnd.n4583 585
R1778 gnd.n4583 gnd.n2548 585
R1779 gnd.n4589 gnd.n4588 585
R1780 gnd.n4590 gnd.n4589 585
R1781 gnd.n1085 gnd.n1084 585
R1782 gnd.n4563 gnd.n1085 585
R1783 gnd.n6673 gnd.n6672 585
R1784 gnd.n6672 gnd.n6671 585
R1785 gnd.n6674 gnd.n1079 585
R1786 gnd.n4569 gnd.n1079 585
R1787 gnd.n6676 gnd.n6675 585
R1788 gnd.n6677 gnd.n6676 585
R1789 gnd.n1064 gnd.n1063 585
R1790 gnd.n4551 gnd.n1064 585
R1791 gnd.n6685 gnd.n6684 585
R1792 gnd.n6684 gnd.n6683 585
R1793 gnd.n6686 gnd.n1058 585
R1794 gnd.n4542 gnd.n1058 585
R1795 gnd.n6688 gnd.n6687 585
R1796 gnd.n6689 gnd.n6688 585
R1797 gnd.n1043 gnd.n1042 585
R1798 gnd.n4529 gnd.n1043 585
R1799 gnd.n6697 gnd.n6696 585
R1800 gnd.n6696 gnd.n6695 585
R1801 gnd.n6698 gnd.n1037 585
R1802 gnd.n4521 gnd.n1037 585
R1803 gnd.n6700 gnd.n6699 585
R1804 gnd.n6701 gnd.n6700 585
R1805 gnd.n1038 gnd.n1036 585
R1806 gnd.n1036 gnd.n1022 585
R1807 gnd.n4493 gnd.n1023 585
R1808 gnd.n6707 gnd.n1023 585
R1809 gnd.n4495 gnd.n4494 585
R1810 gnd.n4494 gnd.n1019 585
R1811 gnd.n4496 gnd.n2620 585
R1812 gnd.n4509 gnd.n2620 585
R1813 gnd.n4497 gnd.n2630 585
R1814 gnd.n2630 gnd.n2618 585
R1815 gnd.n4499 gnd.n4498 585
R1816 gnd.n4500 gnd.n4499 585
R1817 gnd.n2631 gnd.n2629 585
R1818 gnd.n2629 gnd.n2626 585
R1819 gnd.n4484 gnd.n4483 585
R1820 gnd.n4483 gnd.n4482 585
R1821 gnd.n2634 gnd.n2633 585
R1822 gnd.n2645 gnd.n2634 585
R1823 gnd.n4473 gnd.n4472 585
R1824 gnd.n4474 gnd.n4473 585
R1825 gnd.n2647 gnd.n2646 585
R1826 gnd.n2646 gnd.n2642 585
R1827 gnd.n4468 gnd.n4467 585
R1828 gnd.n4467 gnd.n4466 585
R1829 gnd.n2650 gnd.n2649 585
R1830 gnd.n2651 gnd.n2650 585
R1831 gnd.n4457 gnd.n4456 585
R1832 gnd.n4458 gnd.n4457 585
R1833 gnd.n2663 gnd.n2662 585
R1834 gnd.n2662 gnd.n2659 585
R1835 gnd.n4452 gnd.n4451 585
R1836 gnd.n4451 gnd.n4450 585
R1837 gnd.n2666 gnd.n2665 585
R1838 gnd.n4325 gnd.n2666 585
R1839 gnd.n4441 gnd.n4440 585
R1840 gnd.n4442 gnd.n4441 585
R1841 gnd.n4437 gnd.n4326 585
R1842 gnd.n4436 gnd.n4435 585
R1843 gnd.n4433 gnd.n4328 585
R1844 gnd.n4431 gnd.n4430 585
R1845 gnd.n4429 gnd.n4329 585
R1846 gnd.n4428 gnd.n4427 585
R1847 gnd.n4425 gnd.n4334 585
R1848 gnd.n4423 gnd.n4422 585
R1849 gnd.n4421 gnd.n4335 585
R1850 gnd.n4420 gnd.n4419 585
R1851 gnd.n4417 gnd.n4340 585
R1852 gnd.n4415 gnd.n4414 585
R1853 gnd.n4413 gnd.n4341 585
R1854 gnd.n4412 gnd.n4411 585
R1855 gnd.n4409 gnd.n4346 585
R1856 gnd.n4407 gnd.n4406 585
R1857 gnd.n4405 gnd.n4347 585
R1858 gnd.n4399 gnd.n4352 585
R1859 gnd.n4401 gnd.n4400 585
R1860 gnd.n4400 gnd.n4148 585
R1861 gnd.n4926 gnd.n4925 585
R1862 gnd.n2451 gnd.n2450 585
R1863 gnd.n4933 gnd.n2447 585
R1864 gnd.n4934 gnd.n2446 585
R1865 gnd.n2445 gnd.n2439 585
R1866 gnd.n4941 gnd.n2438 585
R1867 gnd.n4942 gnd.n2437 585
R1868 gnd.n2429 gnd.n2428 585
R1869 gnd.n4949 gnd.n2427 585
R1870 gnd.n4950 gnd.n2426 585
R1871 gnd.n2425 gnd.n2419 585
R1872 gnd.n4957 gnd.n2418 585
R1873 gnd.n4958 gnd.n2417 585
R1874 gnd.n2410 gnd.n2409 585
R1875 gnd.n4965 gnd.n2408 585
R1876 gnd.n4966 gnd.n2407 585
R1877 gnd.n2406 gnd.n2405 585
R1878 gnd.n2404 gnd.n2338 585
R1879 gnd.n2337 gnd.n1252 585
R1880 gnd.n6577 gnd.n1252 585
R1881 gnd.n4924 gnd.n2459 585
R1882 gnd.n4924 gnd.n4923 585
R1883 gnd.n4833 gnd.n1243 585
R1884 gnd.n6585 gnd.n1243 585
R1885 gnd.n4874 gnd.n4832 585
R1886 gnd.n4832 gnd.n4831 585
R1887 gnd.n4875 gnd.n1232 585
R1888 gnd.n6591 gnd.n1232 585
R1889 gnd.n4876 gnd.n2484 585
R1890 gnd.n4755 gnd.n2484 585
R1891 gnd.n2482 gnd.n1221 585
R1892 gnd.n6597 gnd.n1221 585
R1893 gnd.n4880 gnd.n2481 585
R1894 gnd.n4751 gnd.n2481 585
R1895 gnd.n4881 gnd.n1210 585
R1896 gnd.n6603 gnd.n1210 585
R1897 gnd.n4882 gnd.n2480 585
R1898 gnd.n4745 gnd.n2480 585
R1899 gnd.n2477 gnd.n1199 585
R1900 gnd.n6609 gnd.n1199 585
R1901 gnd.n4887 gnd.n4886 585
R1902 gnd.n4888 gnd.n4887 585
R1903 gnd.n2476 gnd.n1189 585
R1904 gnd.n6615 gnd.n1189 585
R1905 gnd.n4736 gnd.n4735 585
R1906 gnd.n4737 gnd.n4736 585
R1907 gnd.n2492 gnd.n1178 585
R1908 gnd.n6621 gnd.n1178 585
R1909 gnd.n4731 gnd.n4730 585
R1910 gnd.n4730 gnd.n4729 585
R1911 gnd.n2494 gnd.n1167 585
R1912 gnd.n6627 gnd.n1167 585
R1913 gnd.n4720 gnd.n4719 585
R1914 gnd.n4721 gnd.n4720 585
R1915 gnd.n2498 gnd.n1156 585
R1916 gnd.n6633 gnd.n1156 585
R1917 gnd.n4715 gnd.n4714 585
R1918 gnd.n4714 gnd.n4713 585
R1919 gnd.n2500 gnd.n1146 585
R1920 gnd.n6639 gnd.n1146 585
R1921 gnd.n4664 gnd.n4663 585
R1922 gnd.n4663 gnd.n4662 585
R1923 gnd.n2520 gnd.n1135 585
R1924 gnd.n6645 gnd.n1135 585
R1925 gnd.n4668 gnd.n2519 585
R1926 gnd.n4650 gnd.n2519 585
R1927 gnd.n4669 gnd.n1124 585
R1928 gnd.n6651 gnd.n1124 585
R1929 gnd.n4670 gnd.n2518 585
R1930 gnd.n4646 gnd.n2518 585
R1931 gnd.n2515 gnd.n1114 585
R1932 gnd.n6657 gnd.n1114 585
R1933 gnd.n4675 gnd.n4674 585
R1934 gnd.n4676 gnd.n4675 585
R1935 gnd.n2514 gnd.n1103 585
R1936 gnd.n6663 gnd.n1103 585
R1937 gnd.n4637 gnd.n4636 585
R1938 gnd.n4638 gnd.n4637 585
R1939 gnd.n2529 gnd.n2528 585
R1940 gnd.n4625 gnd.n2528 585
R1941 gnd.n4632 gnd.n4631 585
R1942 gnd.n4631 gnd.n4630 585
R1943 gnd.n2532 gnd.n2531 585
R1944 gnd.n4616 gnd.n2532 585
R1945 gnd.n4578 gnd.n2550 585
R1946 gnd.n4597 gnd.n2550 585
R1947 gnd.n4579 gnd.n2554 585
R1948 gnd.n2554 gnd.n2548 585
R1949 gnd.n4581 gnd.n4580 585
R1950 gnd.n4590 gnd.n4581 585
R1951 gnd.n2555 gnd.n2553 585
R1952 gnd.n4563 gnd.n2553 585
R1953 gnd.n4572 gnd.n1088 585
R1954 gnd.n6671 gnd.n1088 585
R1955 gnd.n4571 gnd.n4570 585
R1956 gnd.n4570 gnd.n4569 585
R1957 gnd.n2557 gnd.n1077 585
R1958 gnd.n6677 gnd.n1077 585
R1959 gnd.n4550 gnd.n4549 585
R1960 gnd.n4551 gnd.n4550 585
R1961 gnd.n2580 gnd.n1067 585
R1962 gnd.n6683 gnd.n1067 585
R1963 gnd.n4544 gnd.n4543 585
R1964 gnd.n4543 gnd.n4542 585
R1965 gnd.n2582 gnd.n1056 585
R1966 gnd.n6689 gnd.n1056 585
R1967 gnd.n4528 gnd.n4527 585
R1968 gnd.n4529 gnd.n4528 585
R1969 gnd.n2610 gnd.n1046 585
R1970 gnd.n6695 gnd.n1046 585
R1971 gnd.n4523 gnd.n4522 585
R1972 gnd.n4522 gnd.n4521 585
R1973 gnd.n2612 gnd.n1034 585
R1974 gnd.n6701 gnd.n1034 585
R1975 gnd.n4371 gnd.n4370 585
R1976 gnd.n4370 gnd.n1022 585
R1977 gnd.n4372 gnd.n1021 585
R1978 gnd.n6707 gnd.n1021 585
R1979 gnd.n4374 gnd.n4373 585
R1980 gnd.n4373 gnd.n1019 585
R1981 gnd.n4375 gnd.n2619 585
R1982 gnd.n4509 gnd.n2619 585
R1983 gnd.n4377 gnd.n4376 585
R1984 gnd.n4376 gnd.n2618 585
R1985 gnd.n4378 gnd.n2628 585
R1986 gnd.n4500 gnd.n2628 585
R1987 gnd.n4380 gnd.n4379 585
R1988 gnd.n4379 gnd.n2626 585
R1989 gnd.n4381 gnd.n2636 585
R1990 gnd.n4482 gnd.n2636 585
R1991 gnd.n4383 gnd.n4382 585
R1992 gnd.n4382 gnd.n2645 585
R1993 gnd.n4384 gnd.n2644 585
R1994 gnd.n4474 gnd.n2644 585
R1995 gnd.n4386 gnd.n4385 585
R1996 gnd.n4385 gnd.n2642 585
R1997 gnd.n4387 gnd.n2653 585
R1998 gnd.n4466 gnd.n2653 585
R1999 gnd.n4389 gnd.n4388 585
R2000 gnd.n4388 gnd.n2651 585
R2001 gnd.n4390 gnd.n2661 585
R2002 gnd.n4458 gnd.n2661 585
R2003 gnd.n4392 gnd.n4391 585
R2004 gnd.n4391 gnd.n2659 585
R2005 gnd.n4393 gnd.n2668 585
R2006 gnd.n4450 gnd.n2668 585
R2007 gnd.n4395 gnd.n4394 585
R2008 gnd.n4394 gnd.n4325 585
R2009 gnd.n4396 gnd.n4150 585
R2010 gnd.n4442 gnd.n4150 585
R2011 gnd.n208 gnd.n129 585
R2012 gnd.n7917 gnd.n129 585
R2013 gnd.n7837 gnd.n7836 585
R2014 gnd.n7838 gnd.n7837 585
R2015 gnd.n207 gnd.n206 585
R2016 gnd.n215 gnd.n206 585
R2017 gnd.n7771 gnd.n7770 585
R2018 gnd.n7770 gnd.n7769 585
R2019 gnd.n211 gnd.n210 585
R2020 gnd.n213 gnd.n211 585
R2021 gnd.n7758 gnd.n7757 585
R2022 gnd.n7759 gnd.n7758 585
R2023 gnd.n225 gnd.n224 585
R2024 gnd.n224 gnd.n222 585
R2025 gnd.n7753 gnd.n7752 585
R2026 gnd.n7752 gnd.n7751 585
R2027 gnd.n228 gnd.n227 585
R2028 gnd.n230 gnd.n228 585
R2029 gnd.n7742 gnd.n7741 585
R2030 gnd.n7743 gnd.n7742 585
R2031 gnd.n239 gnd.n238 585
R2032 gnd.n246 gnd.n238 585
R2033 gnd.n7737 gnd.n7736 585
R2034 gnd.n7736 gnd.n7735 585
R2035 gnd.n242 gnd.n241 585
R2036 gnd.n244 gnd.n242 585
R2037 gnd.n7726 gnd.n7725 585
R2038 gnd.n7727 gnd.n7726 585
R2039 gnd.n255 gnd.n254 585
R2040 gnd.n254 gnd.n252 585
R2041 gnd.n7721 gnd.n7720 585
R2042 gnd.n7720 gnd.n7719 585
R2043 gnd.n258 gnd.n257 585
R2044 gnd.n269 gnd.n258 585
R2045 gnd.n7710 gnd.n7709 585
R2046 gnd.n7711 gnd.n7710 585
R2047 gnd.n271 gnd.n270 585
R2048 gnd.n393 gnd.n270 585
R2049 gnd.n7705 gnd.n7704 585
R2050 gnd.n7704 gnd.n7703 585
R2051 gnd.n274 gnd.n273 585
R2052 gnd.n398 gnd.n274 585
R2053 gnd.n7694 gnd.n7693 585
R2054 gnd.n7695 gnd.n7694 585
R2055 gnd.n287 gnd.n286 585
R2056 gnd.n7624 gnd.n286 585
R2057 gnd.n7689 gnd.n7688 585
R2058 gnd.n7688 gnd.n7687 585
R2059 gnd.n290 gnd.n289 585
R2060 gnd.n7629 gnd.n290 585
R2061 gnd.n7678 gnd.n7677 585
R2062 gnd.n7679 gnd.n7678 585
R2063 gnd.n302 gnd.n301 585
R2064 gnd.n7633 gnd.n301 585
R2065 gnd.n7673 gnd.n7672 585
R2066 gnd.n7672 gnd.n7671 585
R2067 gnd.n305 gnd.n304 585
R2068 gnd.n7638 gnd.n305 585
R2069 gnd.n7651 gnd.n7650 585
R2070 gnd.n7650 gnd.n7649 585
R2071 gnd.n334 gnd.n333 585
R2072 gnd.n7644 gnd.n334 585
R2073 gnd.n7655 gnd.n332 585
R2074 gnd.n1537 gnd.n332 585
R2075 gnd.n7656 gnd.n331 585
R2076 gnd.n6285 gnd.n331 585
R2077 gnd.n7657 gnd.n330 585
R2078 gnd.n6290 gnd.n330 585
R2079 gnd.n327 gnd.n325 585
R2080 gnd.n6186 gnd.n325 585
R2081 gnd.n7662 gnd.n7661 585
R2082 gnd.n7663 gnd.n7662 585
R2083 gnd.n326 gnd.n324 585
R2084 gnd.n6190 gnd.n324 585
R2085 gnd.n6307 gnd.n6306 585
R2086 gnd.n6306 gnd.n6305 585
R2087 gnd.n6310 gnd.n1514 585
R2088 gnd.n6302 gnd.n1514 585
R2089 gnd.n6311 gnd.n1513 585
R2090 gnd.n6195 gnd.n1513 585
R2091 gnd.n6312 gnd.n1512 585
R2092 gnd.n6242 gnd.n1512 585
R2093 gnd.n1548 gnd.n1510 585
R2094 gnd.n1549 gnd.n1548 585
R2095 gnd.n6316 gnd.n1509 585
R2096 gnd.n6232 gnd.n1509 585
R2097 gnd.n6317 gnd.n1508 585
R2098 gnd.n6204 gnd.n1508 585
R2099 gnd.n6318 gnd.n1507 585
R2100 gnd.n6220 gnd.n1507 585
R2101 gnd.n1577 gnd.n1505 585
R2102 gnd.n1578 gnd.n1577 585
R2103 gnd.n6322 gnd.n1504 585
R2104 gnd.n6212 gnd.n1504 585
R2105 gnd.n6323 gnd.n1503 585
R2106 gnd.n6163 gnd.n1503 585
R2107 gnd.n6324 gnd.n1502 585
R2108 gnd.n1605 gnd.n1502 585
R2109 gnd.n1603 gnd.n1500 585
R2110 gnd.n6154 gnd.n1603 585
R2111 gnd.n6328 gnd.n1499 585
R2112 gnd.n1614 gnd.n1499 585
R2113 gnd.n6329 gnd.n1498 585
R2114 gnd.n6144 gnd.n1498 585
R2115 gnd.n6330 gnd.n1497 585
R2116 gnd.n6125 gnd.n1497 585
R2117 gnd.n1621 gnd.n1495 585
R2118 gnd.n1622 gnd.n1621 585
R2119 gnd.n6334 gnd.n1494 585
R2120 gnd.n6116 gnd.n1494 585
R2121 gnd.n6335 gnd.n1493 585
R2122 gnd.n1642 gnd.n1493 585
R2123 gnd.n6336 gnd.n1492 585
R2124 gnd.n6106 gnd.n1492 585
R2125 gnd.n6093 gnd.n1490 585
R2126 gnd.n6094 gnd.n6093 585
R2127 gnd.n6340 gnd.n1489 585
R2128 gnd.n1931 gnd.n1489 585
R2129 gnd.n6341 gnd.n1488 585
R2130 gnd.n6084 gnd.n1488 585
R2131 gnd.n6342 gnd.n1487 585
R2132 gnd.n1668 gnd.n1487 585
R2133 gnd.n6073 gnd.n1485 585
R2134 gnd.n6074 gnd.n6073 585
R2135 gnd.n6346 gnd.n1484 585
R2136 gnd.n6061 gnd.n1484 585
R2137 gnd.n6347 gnd.n1483 585
R2138 gnd.n1675 gnd.n1483 585
R2139 gnd.n6348 gnd.n1482 585
R2140 gnd.n6052 gnd.n1482 585
R2141 gnd.n1709 gnd.n1480 585
R2142 gnd.n5932 gnd.n5931 585
R2143 gnd.n5934 gnd.n5933 585
R2144 gnd.n5926 gnd.n5925 585
R2145 gnd.n5943 gnd.n5927 585
R2146 gnd.n5946 gnd.n5945 585
R2147 gnd.n5944 gnd.n5919 585
R2148 gnd.n5956 gnd.n5955 585
R2149 gnd.n5958 gnd.n5957 585
R2150 gnd.n5914 gnd.n5913 585
R2151 gnd.n5967 gnd.n5915 585
R2152 gnd.n5970 gnd.n5969 585
R2153 gnd.n5968 gnd.n5907 585
R2154 gnd.n5980 gnd.n5979 585
R2155 gnd.n5982 gnd.n5981 585
R2156 gnd.n5902 gnd.n5901 585
R2157 gnd.n5996 gnd.n5903 585
R2158 gnd.n5997 gnd.n5898 585
R2159 gnd.n5998 gnd.n1681 585
R2160 gnd.n6041 gnd.n1681 585
R2161 gnd.n7920 gnd.n7919 585
R2162 gnd.n7806 gnd.n124 585
R2163 gnd.n7808 gnd.n7807 585
R2164 gnd.n7804 gnd.n7803 585
R2165 gnd.n7812 gnd.n7802 585
R2166 gnd.n7813 gnd.n7800 585
R2167 gnd.n7814 gnd.n7799 585
R2168 gnd.n7797 gnd.n7795 585
R2169 gnd.n7818 gnd.n7794 585
R2170 gnd.n7819 gnd.n7792 585
R2171 gnd.n7820 gnd.n7791 585
R2172 gnd.n7789 gnd.n7787 585
R2173 gnd.n7824 gnd.n7786 585
R2174 gnd.n7825 gnd.n7784 585
R2175 gnd.n7826 gnd.n7783 585
R2176 gnd.n7781 gnd.n7779 585
R2177 gnd.n7830 gnd.n7778 585
R2178 gnd.n7831 gnd.n7776 585
R2179 gnd.n7832 gnd.n7775 585
R2180 gnd.n7775 gnd.n128 585
R2181 gnd.n7918 gnd.n120 585
R2182 gnd.n7918 gnd.n7917 585
R2183 gnd.n7924 gnd.n119 585
R2184 gnd.n7838 gnd.n119 585
R2185 gnd.n7925 gnd.n118 585
R2186 gnd.n215 gnd.n118 585
R2187 gnd.n7926 gnd.n117 585
R2188 gnd.n7769 gnd.n117 585
R2189 gnd.n212 gnd.n115 585
R2190 gnd.n213 gnd.n212 585
R2191 gnd.n7930 gnd.n114 585
R2192 gnd.n7759 gnd.n114 585
R2193 gnd.n7931 gnd.n113 585
R2194 gnd.n222 gnd.n113 585
R2195 gnd.n7932 gnd.n112 585
R2196 gnd.n7751 gnd.n112 585
R2197 gnd.n229 gnd.n110 585
R2198 gnd.n230 gnd.n229 585
R2199 gnd.n7936 gnd.n109 585
R2200 gnd.n7743 gnd.n109 585
R2201 gnd.n7937 gnd.n108 585
R2202 gnd.n246 gnd.n108 585
R2203 gnd.n7938 gnd.n107 585
R2204 gnd.n7735 gnd.n107 585
R2205 gnd.n243 gnd.n105 585
R2206 gnd.n244 gnd.n243 585
R2207 gnd.n7942 gnd.n104 585
R2208 gnd.n7727 gnd.n104 585
R2209 gnd.n7943 gnd.n103 585
R2210 gnd.n252 gnd.n103 585
R2211 gnd.n7944 gnd.n102 585
R2212 gnd.n7719 gnd.n102 585
R2213 gnd.n268 gnd.n100 585
R2214 gnd.n269 gnd.n268 585
R2215 gnd.n7948 gnd.n99 585
R2216 gnd.n7711 gnd.n99 585
R2217 gnd.n7949 gnd.n98 585
R2218 gnd.n393 gnd.n98 585
R2219 gnd.n7950 gnd.n97 585
R2220 gnd.n7703 gnd.n97 585
R2221 gnd.n397 gnd.n95 585
R2222 gnd.n398 gnd.n397 585
R2223 gnd.n7954 gnd.n94 585
R2224 gnd.n7695 gnd.n94 585
R2225 gnd.n7955 gnd.n93 585
R2226 gnd.n7624 gnd.n93 585
R2227 gnd.n7956 gnd.n92 585
R2228 gnd.n7687 gnd.n92 585
R2229 gnd.n7628 gnd.n90 585
R2230 gnd.n7629 gnd.n7628 585
R2231 gnd.n7960 gnd.n89 585
R2232 gnd.n7679 gnd.n89 585
R2233 gnd.n7961 gnd.n88 585
R2234 gnd.n7633 gnd.n88 585
R2235 gnd.n7962 gnd.n87 585
R2236 gnd.n7671 gnd.n87 585
R2237 gnd.n7637 gnd.n85 585
R2238 gnd.n7638 gnd.n7637 585
R2239 gnd.n7966 gnd.n84 585
R2240 gnd.n7649 gnd.n84 585
R2241 gnd.n7967 gnd.n83 585
R2242 gnd.n7644 gnd.n83 585
R2243 gnd.n7968 gnd.n82 585
R2244 gnd.n1537 gnd.n82 585
R2245 gnd.n1530 gnd.n80 585
R2246 gnd.n6285 gnd.n1530 585
R2247 gnd.n6292 gnd.n6291 585
R2248 gnd.n6291 gnd.n6290 585
R2249 gnd.n6294 gnd.n1529 585
R2250 gnd.n6186 gnd.n1529 585
R2251 gnd.n6295 gnd.n322 585
R2252 gnd.n7663 gnd.n322 585
R2253 gnd.n6296 gnd.n1528 585
R2254 gnd.n6190 gnd.n1528 585
R2255 gnd.n1525 gnd.n1517 585
R2256 gnd.n6305 gnd.n1517 585
R2257 gnd.n6301 gnd.n6300 585
R2258 gnd.n6302 gnd.n6301 585
R2259 gnd.n1524 gnd.n1523 585
R2260 gnd.n6195 gnd.n1523 585
R2261 gnd.n6225 gnd.n1551 585
R2262 gnd.n6242 gnd.n1551 585
R2263 gnd.n1563 gnd.n1561 585
R2264 gnd.n1561 gnd.n1549 585
R2265 gnd.n6230 gnd.n6229 585
R2266 gnd.n6232 gnd.n6230 585
R2267 gnd.n1562 gnd.n1560 585
R2268 gnd.n6204 gnd.n1560 585
R2269 gnd.n6222 gnd.n6221 585
R2270 gnd.n6221 gnd.n6220 585
R2271 gnd.n1566 gnd.n1565 585
R2272 gnd.n1578 gnd.n1566 585
R2273 gnd.n1596 gnd.n1576 585
R2274 gnd.n6212 gnd.n1576 585
R2275 gnd.n6162 gnd.n6161 585
R2276 gnd.n6163 gnd.n6162 585
R2277 gnd.n1595 gnd.n1594 585
R2278 gnd.n1605 gnd.n1594 585
R2279 gnd.n6156 gnd.n6155 585
R2280 gnd.n6155 gnd.n6154 585
R2281 gnd.n1599 gnd.n1598 585
R2282 gnd.n1614 gnd.n1599 585
R2283 gnd.n1626 gnd.n1613 585
R2284 gnd.n6144 gnd.n1613 585
R2285 gnd.n6124 gnd.n6123 585
R2286 gnd.n6125 gnd.n6124 585
R2287 gnd.n1625 gnd.n1624 585
R2288 gnd.n1624 gnd.n1622 585
R2289 gnd.n6118 gnd.n6117 585
R2290 gnd.n6117 gnd.n6116 585
R2291 gnd.n1629 gnd.n1628 585
R2292 gnd.n1642 gnd.n1629 585
R2293 gnd.n1652 gnd.n1641 585
R2294 gnd.n6106 gnd.n1641 585
R2295 gnd.n6092 gnd.n6091 585
R2296 gnd.n6094 gnd.n6092 585
R2297 gnd.n1651 gnd.n1650 585
R2298 gnd.n1931 gnd.n1650 585
R2299 gnd.n6086 gnd.n6085 585
R2300 gnd.n6085 gnd.n6084 585
R2301 gnd.n1655 gnd.n1654 585
R2302 gnd.n1668 gnd.n1655 585
R2303 gnd.n1679 gnd.n1667 585
R2304 gnd.n6074 gnd.n1667 585
R2305 gnd.n6060 gnd.n6059 585
R2306 gnd.n6061 gnd.n6060 585
R2307 gnd.n1678 gnd.n1677 585
R2308 gnd.n1677 gnd.n1675 585
R2309 gnd.n6054 gnd.n6053 585
R2310 gnd.n6053 gnd.n6052 585
R2311 gnd.n4055 gnd.n4054 585
R2312 gnd.n4056 gnd.n4055 585
R2313 gnd.n2749 gnd.n2748 585
R2314 gnd.n2755 gnd.n2748 585
R2315 gnd.n4030 gnd.n2767 585
R2316 gnd.n2767 gnd.n2754 585
R2317 gnd.n4032 gnd.n4031 585
R2318 gnd.n4033 gnd.n4032 585
R2319 gnd.n2768 gnd.n2766 585
R2320 gnd.n2766 gnd.n2762 585
R2321 gnd.n3764 gnd.n3763 585
R2322 gnd.n3763 gnd.n3762 585
R2323 gnd.n2773 gnd.n2772 585
R2324 gnd.n3733 gnd.n2773 585
R2325 gnd.n3753 gnd.n3752 585
R2326 gnd.n3752 gnd.n3751 585
R2327 gnd.n2780 gnd.n2779 585
R2328 gnd.n3739 gnd.n2780 585
R2329 gnd.n3709 gnd.n2801 585
R2330 gnd.n2801 gnd.n2800 585
R2331 gnd.n3711 gnd.n3710 585
R2332 gnd.n3712 gnd.n3711 585
R2333 gnd.n2802 gnd.n2799 585
R2334 gnd.n2810 gnd.n2799 585
R2335 gnd.n3687 gnd.n2822 585
R2336 gnd.n2822 gnd.n2809 585
R2337 gnd.n3689 gnd.n3688 585
R2338 gnd.n3690 gnd.n3689 585
R2339 gnd.n2823 gnd.n2821 585
R2340 gnd.n2821 gnd.n2817 585
R2341 gnd.n3675 gnd.n3674 585
R2342 gnd.n3674 gnd.n3673 585
R2343 gnd.n2828 gnd.n2827 585
R2344 gnd.n2838 gnd.n2828 585
R2345 gnd.n3664 gnd.n3663 585
R2346 gnd.n3663 gnd.n3662 585
R2347 gnd.n2835 gnd.n2834 585
R2348 gnd.n3650 gnd.n2835 585
R2349 gnd.n3624 gnd.n2856 585
R2350 gnd.n2856 gnd.n2845 585
R2351 gnd.n3626 gnd.n3625 585
R2352 gnd.n3627 gnd.n3626 585
R2353 gnd.n2857 gnd.n2855 585
R2354 gnd.n2865 gnd.n2855 585
R2355 gnd.n3602 gnd.n2877 585
R2356 gnd.n2877 gnd.n2864 585
R2357 gnd.n3604 gnd.n3603 585
R2358 gnd.n3605 gnd.n3604 585
R2359 gnd.n2878 gnd.n2876 585
R2360 gnd.n2876 gnd.n2872 585
R2361 gnd.n3590 gnd.n3589 585
R2362 gnd.n3589 gnd.n3588 585
R2363 gnd.n2883 gnd.n2882 585
R2364 gnd.n2892 gnd.n2883 585
R2365 gnd.n3579 gnd.n3578 585
R2366 gnd.n3578 gnd.n3577 585
R2367 gnd.n2890 gnd.n2889 585
R2368 gnd.n3565 gnd.n2890 585
R2369 gnd.n3003 gnd.n3002 585
R2370 gnd.n3003 gnd.n2899 585
R2371 gnd.n3522 gnd.n3521 585
R2372 gnd.n3521 gnd.n3520 585
R2373 gnd.n3523 gnd.n2997 585
R2374 gnd.n3008 gnd.n2997 585
R2375 gnd.n3525 gnd.n3524 585
R2376 gnd.n3526 gnd.n3525 585
R2377 gnd.n2998 gnd.n2996 585
R2378 gnd.n3021 gnd.n2996 585
R2379 gnd.n2981 gnd.n2980 585
R2380 gnd.n2984 gnd.n2981 585
R2381 gnd.n3536 gnd.n3535 585
R2382 gnd.n3535 gnd.n3534 585
R2383 gnd.n3537 gnd.n2975 585
R2384 gnd.n3496 gnd.n2975 585
R2385 gnd.n3539 gnd.n3538 585
R2386 gnd.n3540 gnd.n3539 585
R2387 gnd.n2976 gnd.n2974 585
R2388 gnd.n3035 gnd.n2974 585
R2389 gnd.n3488 gnd.n3487 585
R2390 gnd.n3487 gnd.n3486 585
R2391 gnd.n3032 gnd.n3031 585
R2392 gnd.n3470 gnd.n3032 585
R2393 gnd.n3457 gnd.n3051 585
R2394 gnd.n3051 gnd.n3050 585
R2395 gnd.n3459 gnd.n3458 585
R2396 gnd.n3460 gnd.n3459 585
R2397 gnd.n3052 gnd.n3049 585
R2398 gnd.n3058 gnd.n3049 585
R2399 gnd.n3438 gnd.n3437 585
R2400 gnd.n3439 gnd.n3438 585
R2401 gnd.n3069 gnd.n3068 585
R2402 gnd.n3068 gnd.n3064 585
R2403 gnd.n3428 gnd.n3427 585
R2404 gnd.n3429 gnd.n3428 585
R2405 gnd.n3079 gnd.n3078 585
R2406 gnd.n3084 gnd.n3078 585
R2407 gnd.n3406 gnd.n3097 585
R2408 gnd.n3097 gnd.n3083 585
R2409 gnd.n3408 gnd.n3407 585
R2410 gnd.n3409 gnd.n3408 585
R2411 gnd.n3098 gnd.n3096 585
R2412 gnd.n3096 gnd.n3092 585
R2413 gnd.n3397 gnd.n3396 585
R2414 gnd.n3398 gnd.n3397 585
R2415 gnd.n3105 gnd.n3104 585
R2416 gnd.n3109 gnd.n3104 585
R2417 gnd.n3374 gnd.n3126 585
R2418 gnd.n3126 gnd.n3108 585
R2419 gnd.n3376 gnd.n3375 585
R2420 gnd.n3377 gnd.n3376 585
R2421 gnd.n3127 gnd.n3125 585
R2422 gnd.n3125 gnd.n3116 585
R2423 gnd.n3369 gnd.n3368 585
R2424 gnd.n3368 gnd.n3367 585
R2425 gnd.n3174 gnd.n3173 585
R2426 gnd.n3175 gnd.n3174 585
R2427 gnd.n3328 gnd.n3327 585
R2428 gnd.n3329 gnd.n3328 585
R2429 gnd.n3184 gnd.n3183 585
R2430 gnd.n3183 gnd.n3182 585
R2431 gnd.n3323 gnd.n3322 585
R2432 gnd.n3322 gnd.n3321 585
R2433 gnd.n3187 gnd.n3186 585
R2434 gnd.n3188 gnd.n3187 585
R2435 gnd.n3312 gnd.n3311 585
R2436 gnd.n3313 gnd.n3312 585
R2437 gnd.n3195 gnd.n3194 585
R2438 gnd.n3304 gnd.n3194 585
R2439 gnd.n3307 gnd.n3306 585
R2440 gnd.n3306 gnd.n3305 585
R2441 gnd.n3198 gnd.n3197 585
R2442 gnd.n3199 gnd.n3198 585
R2443 gnd.n3293 gnd.n3292 585
R2444 gnd.n3291 gnd.n3217 585
R2445 gnd.n3290 gnd.n3216 585
R2446 gnd.n3295 gnd.n3216 585
R2447 gnd.n3289 gnd.n3288 585
R2448 gnd.n3287 gnd.n3286 585
R2449 gnd.n3285 gnd.n3284 585
R2450 gnd.n3283 gnd.n3282 585
R2451 gnd.n3281 gnd.n3280 585
R2452 gnd.n3279 gnd.n3278 585
R2453 gnd.n3277 gnd.n3276 585
R2454 gnd.n3275 gnd.n3274 585
R2455 gnd.n3273 gnd.n3272 585
R2456 gnd.n3271 gnd.n3270 585
R2457 gnd.n3269 gnd.n3268 585
R2458 gnd.n3267 gnd.n3266 585
R2459 gnd.n3265 gnd.n3264 585
R2460 gnd.n3263 gnd.n3262 585
R2461 gnd.n3261 gnd.n3260 585
R2462 gnd.n3259 gnd.n3258 585
R2463 gnd.n3257 gnd.n3256 585
R2464 gnd.n3255 gnd.n3254 585
R2465 gnd.n3253 gnd.n3252 585
R2466 gnd.n3251 gnd.n3250 585
R2467 gnd.n3249 gnd.n3248 585
R2468 gnd.n3247 gnd.n3246 585
R2469 gnd.n3204 gnd.n3203 585
R2470 gnd.n3298 gnd.n3297 585
R2471 gnd.n4059 gnd.n4058 585
R2472 gnd.n4061 gnd.n4060 585
R2473 gnd.n4063 gnd.n4062 585
R2474 gnd.n4065 gnd.n4064 585
R2475 gnd.n4067 gnd.n4066 585
R2476 gnd.n4069 gnd.n4068 585
R2477 gnd.n4071 gnd.n4070 585
R2478 gnd.n4073 gnd.n4072 585
R2479 gnd.n4075 gnd.n4074 585
R2480 gnd.n4077 gnd.n4076 585
R2481 gnd.n4079 gnd.n4078 585
R2482 gnd.n4081 gnd.n4080 585
R2483 gnd.n4083 gnd.n4082 585
R2484 gnd.n4085 gnd.n4084 585
R2485 gnd.n4087 gnd.n4086 585
R2486 gnd.n4089 gnd.n4088 585
R2487 gnd.n4091 gnd.n4090 585
R2488 gnd.n4093 gnd.n4092 585
R2489 gnd.n4095 gnd.n4094 585
R2490 gnd.n4097 gnd.n4096 585
R2491 gnd.n4099 gnd.n4098 585
R2492 gnd.n4101 gnd.n4100 585
R2493 gnd.n4103 gnd.n4102 585
R2494 gnd.n4105 gnd.n4104 585
R2495 gnd.n4107 gnd.n4106 585
R2496 gnd.n4108 gnd.n2716 585
R2497 gnd.n4109 gnd.n2674 585
R2498 gnd.n4147 gnd.n2674 585
R2499 gnd.n4057 gnd.n2746 585
R2500 gnd.n4057 gnd.n4056 585
R2501 gnd.n3726 gnd.n2745 585
R2502 gnd.n2755 gnd.n2745 585
R2503 gnd.n3728 gnd.n3727 585
R2504 gnd.n3727 gnd.n2754 585
R2505 gnd.n3729 gnd.n2764 585
R2506 gnd.n4033 gnd.n2764 585
R2507 gnd.n3731 gnd.n3730 585
R2508 gnd.n3730 gnd.n2762 585
R2509 gnd.n3732 gnd.n2775 585
R2510 gnd.n3762 gnd.n2775 585
R2511 gnd.n3735 gnd.n3734 585
R2512 gnd.n3734 gnd.n3733 585
R2513 gnd.n3736 gnd.n2782 585
R2514 gnd.n3751 gnd.n2782 585
R2515 gnd.n3738 gnd.n3737 585
R2516 gnd.n3739 gnd.n3738 585
R2517 gnd.n2793 gnd.n2792 585
R2518 gnd.n2800 gnd.n2792 585
R2519 gnd.n3714 gnd.n3713 585
R2520 gnd.n3713 gnd.n3712 585
R2521 gnd.n2796 gnd.n2795 585
R2522 gnd.n2810 gnd.n2796 585
R2523 gnd.n3640 gnd.n3639 585
R2524 gnd.n3639 gnd.n2809 585
R2525 gnd.n3641 gnd.n2819 585
R2526 gnd.n3690 gnd.n2819 585
R2527 gnd.n3643 gnd.n3642 585
R2528 gnd.n3642 gnd.n2817 585
R2529 gnd.n3644 gnd.n2830 585
R2530 gnd.n3673 gnd.n2830 585
R2531 gnd.n3646 gnd.n3645 585
R2532 gnd.n3645 gnd.n2838 585
R2533 gnd.n3647 gnd.n2837 585
R2534 gnd.n3662 gnd.n2837 585
R2535 gnd.n3649 gnd.n3648 585
R2536 gnd.n3650 gnd.n3649 585
R2537 gnd.n2849 gnd.n2848 585
R2538 gnd.n2848 gnd.n2845 585
R2539 gnd.n3629 gnd.n3628 585
R2540 gnd.n3628 gnd.n3627 585
R2541 gnd.n2852 gnd.n2851 585
R2542 gnd.n2865 gnd.n2852 585
R2543 gnd.n3553 gnd.n3552 585
R2544 gnd.n3552 gnd.n2864 585
R2545 gnd.n3554 gnd.n2874 585
R2546 gnd.n3605 gnd.n2874 585
R2547 gnd.n3556 gnd.n3555 585
R2548 gnd.n3555 gnd.n2872 585
R2549 gnd.n3557 gnd.n2885 585
R2550 gnd.n3588 gnd.n2885 585
R2551 gnd.n3559 gnd.n3558 585
R2552 gnd.n3558 gnd.n2892 585
R2553 gnd.n3560 gnd.n2891 585
R2554 gnd.n3577 gnd.n2891 585
R2555 gnd.n3562 gnd.n3561 585
R2556 gnd.n3565 gnd.n3562 585
R2557 gnd.n2902 gnd.n2901 585
R2558 gnd.n2901 gnd.n2899 585
R2559 gnd.n3005 gnd.n3004 585
R2560 gnd.n3520 gnd.n3004 585
R2561 gnd.n3007 gnd.n3006 585
R2562 gnd.n3008 gnd.n3007 585
R2563 gnd.n3018 gnd.n2994 585
R2564 gnd.n3526 gnd.n2994 585
R2565 gnd.n3020 gnd.n3019 585
R2566 gnd.n3021 gnd.n3020 585
R2567 gnd.n3017 gnd.n3016 585
R2568 gnd.n3017 gnd.n2984 585
R2569 gnd.n3015 gnd.n2982 585
R2570 gnd.n3534 gnd.n2982 585
R2571 gnd.n2971 gnd.n2969 585
R2572 gnd.n3496 gnd.n2971 585
R2573 gnd.n3542 gnd.n3541 585
R2574 gnd.n3541 gnd.n3540 585
R2575 gnd.n2970 gnd.n2968 585
R2576 gnd.n3035 gnd.n2970 585
R2577 gnd.n3467 gnd.n3034 585
R2578 gnd.n3486 gnd.n3034 585
R2579 gnd.n3469 gnd.n3468 585
R2580 gnd.n3470 gnd.n3469 585
R2581 gnd.n3044 gnd.n3043 585
R2582 gnd.n3050 gnd.n3043 585
R2583 gnd.n3462 gnd.n3461 585
R2584 gnd.n3461 gnd.n3460 585
R2585 gnd.n3047 gnd.n3046 585
R2586 gnd.n3058 gnd.n3047 585
R2587 gnd.n3347 gnd.n3066 585
R2588 gnd.n3439 gnd.n3066 585
R2589 gnd.n3349 gnd.n3348 585
R2590 gnd.n3348 gnd.n3064 585
R2591 gnd.n3350 gnd.n3077 585
R2592 gnd.n3429 gnd.n3077 585
R2593 gnd.n3352 gnd.n3351 585
R2594 gnd.n3352 gnd.n3084 585
R2595 gnd.n3354 gnd.n3353 585
R2596 gnd.n3353 gnd.n3083 585
R2597 gnd.n3355 gnd.n3094 585
R2598 gnd.n3409 gnd.n3094 585
R2599 gnd.n3357 gnd.n3356 585
R2600 gnd.n3356 gnd.n3092 585
R2601 gnd.n3358 gnd.n3103 585
R2602 gnd.n3398 gnd.n3103 585
R2603 gnd.n3360 gnd.n3359 585
R2604 gnd.n3360 gnd.n3109 585
R2605 gnd.n3362 gnd.n3361 585
R2606 gnd.n3361 gnd.n3108 585
R2607 gnd.n3363 gnd.n3124 585
R2608 gnd.n3377 gnd.n3124 585
R2609 gnd.n3364 gnd.n3177 585
R2610 gnd.n3177 gnd.n3116 585
R2611 gnd.n3366 gnd.n3365 585
R2612 gnd.n3367 gnd.n3366 585
R2613 gnd.n3178 gnd.n3176 585
R2614 gnd.n3176 gnd.n3175 585
R2615 gnd.n3331 gnd.n3330 585
R2616 gnd.n3330 gnd.n3329 585
R2617 gnd.n3181 gnd.n3180 585
R2618 gnd.n3182 gnd.n3181 585
R2619 gnd.n3320 gnd.n3319 585
R2620 gnd.n3321 gnd.n3320 585
R2621 gnd.n3190 gnd.n3189 585
R2622 gnd.n3189 gnd.n3188 585
R2623 gnd.n3315 gnd.n3314 585
R2624 gnd.n3314 gnd.n3313 585
R2625 gnd.n3193 gnd.n3192 585
R2626 gnd.n3304 gnd.n3193 585
R2627 gnd.n3303 gnd.n3302 585
R2628 gnd.n3305 gnd.n3303 585
R2629 gnd.n3201 gnd.n3200 585
R2630 gnd.n3200 gnd.n3199 585
R2631 gnd.n4042 gnd.n2696 585
R2632 gnd.n2696 gnd.n2673 585
R2633 gnd.n4043 gnd.n2757 585
R2634 gnd.n2757 gnd.n2747 585
R2635 gnd.n4045 gnd.n4044 585
R2636 gnd.n4046 gnd.n4045 585
R2637 gnd.n2758 gnd.n2756 585
R2638 gnd.n2765 gnd.n2756 585
R2639 gnd.n4036 gnd.n4035 585
R2640 gnd.n4035 gnd.n4034 585
R2641 gnd.n2761 gnd.n2760 585
R2642 gnd.n3761 gnd.n2761 585
R2643 gnd.n3747 gnd.n2784 585
R2644 gnd.n2784 gnd.n2774 585
R2645 gnd.n3749 gnd.n3748 585
R2646 gnd.n3750 gnd.n3749 585
R2647 gnd.n2785 gnd.n2783 585
R2648 gnd.n2783 gnd.n2781 585
R2649 gnd.n3742 gnd.n3741 585
R2650 gnd.n3741 gnd.n3740 585
R2651 gnd.n2788 gnd.n2787 585
R2652 gnd.n2798 gnd.n2788 585
R2653 gnd.n3698 gnd.n2812 585
R2654 gnd.n2812 gnd.n2797 585
R2655 gnd.n3700 gnd.n3699 585
R2656 gnd.n3701 gnd.n3700 585
R2657 gnd.n2813 gnd.n2811 585
R2658 gnd.n2820 gnd.n2811 585
R2659 gnd.n3693 gnd.n3692 585
R2660 gnd.n3692 gnd.n3691 585
R2661 gnd.n2816 gnd.n2815 585
R2662 gnd.n3672 gnd.n2816 585
R2663 gnd.n3658 gnd.n2840 585
R2664 gnd.n2840 gnd.n2829 585
R2665 gnd.n3660 gnd.n3659 585
R2666 gnd.n3661 gnd.n3660 585
R2667 gnd.n2841 gnd.n2839 585
R2668 gnd.n2839 gnd.n2836 585
R2669 gnd.n3653 gnd.n3652 585
R2670 gnd.n3652 gnd.n3651 585
R2671 gnd.n2844 gnd.n2843 585
R2672 gnd.n2854 gnd.n2844 585
R2673 gnd.n3613 gnd.n2867 585
R2674 gnd.n2867 gnd.n2853 585
R2675 gnd.n3615 gnd.n3614 585
R2676 gnd.n3616 gnd.n3615 585
R2677 gnd.n2868 gnd.n2866 585
R2678 gnd.n2875 gnd.n2866 585
R2679 gnd.n3608 gnd.n3607 585
R2680 gnd.n3607 gnd.n3606 585
R2681 gnd.n2871 gnd.n2870 585
R2682 gnd.n3587 gnd.n2871 585
R2683 gnd.n3573 gnd.n2894 585
R2684 gnd.n2894 gnd.n2884 585
R2685 gnd.n3575 gnd.n3574 585
R2686 gnd.n3576 gnd.n3575 585
R2687 gnd.n2895 gnd.n2893 585
R2688 gnd.n3564 gnd.n2893 585
R2689 gnd.n3568 gnd.n3567 585
R2690 gnd.n3567 gnd.n3566 585
R2691 gnd.n2898 gnd.n2897 585
R2692 gnd.n3519 gnd.n2898 585
R2693 gnd.n3012 gnd.n3011 585
R2694 gnd.n3013 gnd.n3012 585
R2695 gnd.n2992 gnd.n2991 585
R2696 gnd.n2995 gnd.n2992 585
R2697 gnd.n3529 gnd.n3528 585
R2698 gnd.n3528 gnd.n3527 585
R2699 gnd.n3530 gnd.n2986 585
R2700 gnd.n3022 gnd.n2986 585
R2701 gnd.n3532 gnd.n3531 585
R2702 gnd.n3533 gnd.n3532 585
R2703 gnd.n2987 gnd.n2985 585
R2704 gnd.n3497 gnd.n2985 585
R2705 gnd.n3481 gnd.n3480 585
R2706 gnd.n3480 gnd.n2973 585
R2707 gnd.n3482 gnd.n3037 585
R2708 gnd.n3037 gnd.n2972 585
R2709 gnd.n3484 gnd.n3483 585
R2710 gnd.n3485 gnd.n3484 585
R2711 gnd.n3038 gnd.n3036 585
R2712 gnd.n3036 gnd.n3033 585
R2713 gnd.n3473 gnd.n3472 585
R2714 gnd.n3472 gnd.n3471 585
R2715 gnd.n3041 gnd.n3040 585
R2716 gnd.n3048 gnd.n3041 585
R2717 gnd.n3447 gnd.n3446 585
R2718 gnd.n3448 gnd.n3447 585
R2719 gnd.n3060 gnd.n3059 585
R2720 gnd.n3067 gnd.n3059 585
R2721 gnd.n3442 gnd.n3441 585
R2722 gnd.n3441 gnd.n3440 585
R2723 gnd.n3063 gnd.n3062 585
R2724 gnd.n3430 gnd.n3063 585
R2725 gnd.n3417 gnd.n3087 585
R2726 gnd.n3087 gnd.n3086 585
R2727 gnd.n3419 gnd.n3418 585
R2728 gnd.n3420 gnd.n3419 585
R2729 gnd.n3088 gnd.n3085 585
R2730 gnd.n3095 gnd.n3085 585
R2731 gnd.n3412 gnd.n3411 585
R2732 gnd.n3411 gnd.n3410 585
R2733 gnd.n3091 gnd.n3090 585
R2734 gnd.n3399 gnd.n3091 585
R2735 gnd.n3386 gnd.n3112 585
R2736 gnd.n3112 gnd.n3111 585
R2737 gnd.n3388 gnd.n3387 585
R2738 gnd.n3389 gnd.n3388 585
R2739 gnd.n3382 gnd.n3110 585
R2740 gnd.n3381 gnd.n3380 585
R2741 gnd.n3115 gnd.n3114 585
R2742 gnd.n3378 gnd.n3115 585
R2743 gnd.n3137 gnd.n3136 585
R2744 gnd.n3140 gnd.n3139 585
R2745 gnd.n3138 gnd.n3133 585
R2746 gnd.n3145 gnd.n3144 585
R2747 gnd.n3147 gnd.n3146 585
R2748 gnd.n3150 gnd.n3149 585
R2749 gnd.n3148 gnd.n3131 585
R2750 gnd.n3155 gnd.n3154 585
R2751 gnd.n3157 gnd.n3156 585
R2752 gnd.n3160 gnd.n3159 585
R2753 gnd.n3158 gnd.n3129 585
R2754 gnd.n3165 gnd.n3164 585
R2755 gnd.n3169 gnd.n3166 585
R2756 gnd.n3170 gnd.n3107 585
R2757 gnd.n4048 gnd.n2711 585
R2758 gnd.n4115 gnd.n4114 585
R2759 gnd.n4117 gnd.n4116 585
R2760 gnd.n4119 gnd.n4118 585
R2761 gnd.n4121 gnd.n4120 585
R2762 gnd.n4123 gnd.n4122 585
R2763 gnd.n4125 gnd.n4124 585
R2764 gnd.n4127 gnd.n4126 585
R2765 gnd.n4129 gnd.n4128 585
R2766 gnd.n4131 gnd.n4130 585
R2767 gnd.n4133 gnd.n4132 585
R2768 gnd.n4135 gnd.n4134 585
R2769 gnd.n4137 gnd.n4136 585
R2770 gnd.n4140 gnd.n4139 585
R2771 gnd.n4138 gnd.n2699 585
R2772 gnd.n4144 gnd.n2697 585
R2773 gnd.n4146 gnd.n4145 585
R2774 gnd.n4147 gnd.n4146 585
R2775 gnd.n4049 gnd.n2752 585
R2776 gnd.n4049 gnd.n2673 585
R2777 gnd.n4051 gnd.n4050 585
R2778 gnd.n4050 gnd.n2747 585
R2779 gnd.n4047 gnd.n2751 585
R2780 gnd.n4047 gnd.n4046 585
R2781 gnd.n4026 gnd.n2753 585
R2782 gnd.n2765 gnd.n2753 585
R2783 gnd.n4025 gnd.n2763 585
R2784 gnd.n4034 gnd.n2763 585
R2785 gnd.n3760 gnd.n2770 585
R2786 gnd.n3761 gnd.n3760 585
R2787 gnd.n3759 gnd.n3758 585
R2788 gnd.n3759 gnd.n2774 585
R2789 gnd.n3757 gnd.n2776 585
R2790 gnd.n3750 gnd.n2776 585
R2791 gnd.n2790 gnd.n2777 585
R2792 gnd.n2790 gnd.n2781 585
R2793 gnd.n3706 gnd.n2791 585
R2794 gnd.n3740 gnd.n2791 585
R2795 gnd.n3705 gnd.n3704 585
R2796 gnd.n3704 gnd.n2798 585
R2797 gnd.n3703 gnd.n2806 585
R2798 gnd.n3703 gnd.n2797 585
R2799 gnd.n3702 gnd.n2808 585
R2800 gnd.n3702 gnd.n3701 585
R2801 gnd.n3681 gnd.n2807 585
R2802 gnd.n2820 gnd.n2807 585
R2803 gnd.n3680 gnd.n2818 585
R2804 gnd.n3691 gnd.n2818 585
R2805 gnd.n3671 gnd.n2825 585
R2806 gnd.n3672 gnd.n3671 585
R2807 gnd.n3670 gnd.n3669 585
R2808 gnd.n3670 gnd.n2829 585
R2809 gnd.n3668 gnd.n2831 585
R2810 gnd.n3661 gnd.n2831 585
R2811 gnd.n2846 gnd.n2832 585
R2812 gnd.n2846 gnd.n2836 585
R2813 gnd.n3621 gnd.n2847 585
R2814 gnd.n3651 gnd.n2847 585
R2815 gnd.n3620 gnd.n3619 585
R2816 gnd.n3619 gnd.n2854 585
R2817 gnd.n3618 gnd.n2861 585
R2818 gnd.n3618 gnd.n2853 585
R2819 gnd.n3617 gnd.n2863 585
R2820 gnd.n3617 gnd.n3616 585
R2821 gnd.n3596 gnd.n2862 585
R2822 gnd.n2875 gnd.n2862 585
R2823 gnd.n3595 gnd.n2873 585
R2824 gnd.n3606 gnd.n2873 585
R2825 gnd.n3586 gnd.n2880 585
R2826 gnd.n3587 gnd.n3586 585
R2827 gnd.n3585 gnd.n3584 585
R2828 gnd.n3585 gnd.n2884 585
R2829 gnd.n3583 gnd.n2886 585
R2830 gnd.n3576 gnd.n2886 585
R2831 gnd.n3563 gnd.n2887 585
R2832 gnd.n3564 gnd.n3563 585
R2833 gnd.n3516 gnd.n2900 585
R2834 gnd.n3566 gnd.n2900 585
R2835 gnd.n3518 gnd.n3517 585
R2836 gnd.n3519 gnd.n3518 585
R2837 gnd.n3511 gnd.n3014 585
R2838 gnd.n3014 gnd.n3013 585
R2839 gnd.n3509 gnd.n3508 585
R2840 gnd.n3508 gnd.n2995 585
R2841 gnd.n3506 gnd.n2993 585
R2842 gnd.n3527 gnd.n2993 585
R2843 gnd.n3024 gnd.n3023 585
R2844 gnd.n3023 gnd.n3022 585
R2845 gnd.n3500 gnd.n2983 585
R2846 gnd.n3533 gnd.n2983 585
R2847 gnd.n3499 gnd.n3498 585
R2848 gnd.n3498 gnd.n3497 585
R2849 gnd.n3495 gnd.n3026 585
R2850 gnd.n3495 gnd.n2973 585
R2851 gnd.n3494 gnd.n3493 585
R2852 gnd.n3494 gnd.n2972 585
R2853 gnd.n3029 gnd.n3028 585
R2854 gnd.n3485 gnd.n3028 585
R2855 gnd.n3453 gnd.n3452 585
R2856 gnd.n3452 gnd.n3033 585
R2857 gnd.n3454 gnd.n3042 585
R2858 gnd.n3471 gnd.n3042 585
R2859 gnd.n3451 gnd.n3450 585
R2860 gnd.n3450 gnd.n3048 585
R2861 gnd.n3449 gnd.n3056 585
R2862 gnd.n3449 gnd.n3448 585
R2863 gnd.n3434 gnd.n3057 585
R2864 gnd.n3067 gnd.n3057 585
R2865 gnd.n3433 gnd.n3065 585
R2866 gnd.n3440 gnd.n3065 585
R2867 gnd.n3432 gnd.n3431 585
R2868 gnd.n3431 gnd.n3430 585
R2869 gnd.n3076 gnd.n3073 585
R2870 gnd.n3086 gnd.n3076 585
R2871 gnd.n3422 gnd.n3421 585
R2872 gnd.n3421 gnd.n3420 585
R2873 gnd.n3082 gnd.n3081 585
R2874 gnd.n3095 gnd.n3082 585
R2875 gnd.n3402 gnd.n3093 585
R2876 gnd.n3410 gnd.n3093 585
R2877 gnd.n3401 gnd.n3400 585
R2878 gnd.n3400 gnd.n3399 585
R2879 gnd.n3102 gnd.n3100 585
R2880 gnd.n3111 gnd.n3102 585
R2881 gnd.n3391 gnd.n3390 585
R2882 gnd.n3390 gnd.n3389 585
R2883 gnd.n6582 gnd.n1245 585
R2884 gnd.n4923 gnd.n1245 585
R2885 gnd.n6584 gnd.n6583 585
R2886 gnd.n6585 gnd.n6584 585
R2887 gnd.n1229 gnd.n1228 585
R2888 gnd.n4831 gnd.n1229 585
R2889 gnd.n6593 gnd.n6592 585
R2890 gnd.n6592 gnd.n6591 585
R2891 gnd.n6594 gnd.n1223 585
R2892 gnd.n4755 gnd.n1223 585
R2893 gnd.n6596 gnd.n6595 585
R2894 gnd.n6597 gnd.n6596 585
R2895 gnd.n1207 gnd.n1206 585
R2896 gnd.n4751 gnd.n1207 585
R2897 gnd.n6605 gnd.n6604 585
R2898 gnd.n6604 gnd.n6603 585
R2899 gnd.n6606 gnd.n1201 585
R2900 gnd.n4745 gnd.n1201 585
R2901 gnd.n6608 gnd.n6607 585
R2902 gnd.n6609 gnd.n6608 585
R2903 gnd.n1186 gnd.n1185 585
R2904 gnd.n4888 gnd.n1186 585
R2905 gnd.n6617 gnd.n6616 585
R2906 gnd.n6616 gnd.n6615 585
R2907 gnd.n6618 gnd.n1180 585
R2908 gnd.n4737 gnd.n1180 585
R2909 gnd.n6620 gnd.n6619 585
R2910 gnd.n6621 gnd.n6620 585
R2911 gnd.n1164 gnd.n1163 585
R2912 gnd.n4729 gnd.n1164 585
R2913 gnd.n6629 gnd.n6628 585
R2914 gnd.n6628 gnd.n6627 585
R2915 gnd.n6630 gnd.n1158 585
R2916 gnd.n4721 gnd.n1158 585
R2917 gnd.n6632 gnd.n6631 585
R2918 gnd.n6633 gnd.n6632 585
R2919 gnd.n1143 gnd.n1142 585
R2920 gnd.n4713 gnd.n1143 585
R2921 gnd.n6641 gnd.n6640 585
R2922 gnd.n6640 gnd.n6639 585
R2923 gnd.n6642 gnd.n1137 585
R2924 gnd.n4662 gnd.n1137 585
R2925 gnd.n6644 gnd.n6643 585
R2926 gnd.n6645 gnd.n6644 585
R2927 gnd.n1121 gnd.n1120 585
R2928 gnd.n4650 gnd.n1121 585
R2929 gnd.n6653 gnd.n6652 585
R2930 gnd.n6652 gnd.n6651 585
R2931 gnd.n6654 gnd.n1116 585
R2932 gnd.n4646 gnd.n1116 585
R2933 gnd.n6656 gnd.n6655 585
R2934 gnd.n6657 gnd.n6656 585
R2935 gnd.n1100 gnd.n1098 585
R2936 gnd.n4676 gnd.n1100 585
R2937 gnd.n6665 gnd.n6664 585
R2938 gnd.n6664 gnd.n6663 585
R2939 gnd.n1099 gnd.n1097 585
R2940 gnd.n4638 gnd.n1099 585
R2941 gnd.n4627 gnd.n4626 585
R2942 gnd.n4626 gnd.n4625 585
R2943 gnd.n4629 gnd.n4628 585
R2944 gnd.n4630 gnd.n4629 585
R2945 gnd.n4594 gnd.n2536 585
R2946 gnd.n4616 gnd.n2536 585
R2947 gnd.n4596 gnd.n4595 585
R2948 gnd.n4597 gnd.n4596 585
R2949 gnd.n4593 gnd.n4592 585
R2950 gnd.n4593 gnd.n2548 585
R2951 gnd.n4591 gnd.n1091 585
R2952 gnd.n4591 gnd.n4590 585
R2953 gnd.n6668 gnd.n1089 585
R2954 gnd.n4563 gnd.n1089 585
R2955 gnd.n6670 gnd.n6669 585
R2956 gnd.n6671 gnd.n6670 585
R2957 gnd.n1075 gnd.n1074 585
R2958 gnd.n4569 gnd.n1075 585
R2959 gnd.n6679 gnd.n6678 585
R2960 gnd.n6678 gnd.n6677 585
R2961 gnd.n6680 gnd.n1069 585
R2962 gnd.n4551 gnd.n1069 585
R2963 gnd.n6682 gnd.n6681 585
R2964 gnd.n6683 gnd.n6682 585
R2965 gnd.n1053 gnd.n1052 585
R2966 gnd.n4542 gnd.n1053 585
R2967 gnd.n6691 gnd.n6690 585
R2968 gnd.n6690 gnd.n6689 585
R2969 gnd.n6692 gnd.n1047 585
R2970 gnd.n4529 gnd.n1047 585
R2971 gnd.n6694 gnd.n6693 585
R2972 gnd.n6695 gnd.n6694 585
R2973 gnd.n1031 gnd.n1030 585
R2974 gnd.n4521 gnd.n1031 585
R2975 gnd.n6703 gnd.n6702 585
R2976 gnd.n6702 gnd.n6701 585
R2977 gnd.n6704 gnd.n1025 585
R2978 gnd.n1025 gnd.n1022 585
R2979 gnd.n6706 gnd.n6705 585
R2980 gnd.n6707 gnd.n6706 585
R2981 gnd.n1026 gnd.n1024 585
R2982 gnd.n1024 gnd.n1019 585
R2983 gnd.n4508 gnd.n4507 585
R2984 gnd.n4509 gnd.n4508 585
R2985 gnd.n2622 gnd.n2621 585
R2986 gnd.n2621 gnd.n2618 585
R2987 gnd.n4502 gnd.n4501 585
R2988 gnd.n4501 gnd.n4500 585
R2989 gnd.n2625 gnd.n2624 585
R2990 gnd.n2626 gnd.n2625 585
R2991 gnd.n4481 gnd.n4480 585
R2992 gnd.n4482 gnd.n4481 585
R2993 gnd.n2638 gnd.n2637 585
R2994 gnd.n2645 gnd.n2637 585
R2995 gnd.n4476 gnd.n4475 585
R2996 gnd.n4475 gnd.n4474 585
R2997 gnd.n2641 gnd.n2640 585
R2998 gnd.n2642 gnd.n2641 585
R2999 gnd.n4465 gnd.n4464 585
R3000 gnd.n4466 gnd.n4465 585
R3001 gnd.n2655 gnd.n2654 585
R3002 gnd.n2654 gnd.n2651 585
R3003 gnd.n4460 gnd.n4459 585
R3004 gnd.n4459 gnd.n4458 585
R3005 gnd.n2658 gnd.n2657 585
R3006 gnd.n2659 gnd.n2658 585
R3007 gnd.n4449 gnd.n4448 585
R3008 gnd.n4450 gnd.n4449 585
R3009 gnd.n2670 gnd.n2669 585
R3010 gnd.n4325 gnd.n2669 585
R3011 gnd.n4444 gnd.n4443 585
R3012 gnd.n4443 gnd.n4442 585
R3013 gnd.n4195 gnd.n2672 585
R3014 gnd.n4198 gnd.n4197 585
R3015 gnd.n4194 gnd.n4193 585
R3016 gnd.n4193 gnd.n4148 585
R3017 gnd.n4203 gnd.n4202 585
R3018 gnd.n4205 gnd.n4192 585
R3019 gnd.n4208 gnd.n4207 585
R3020 gnd.n4190 gnd.n4189 585
R3021 gnd.n4213 gnd.n4212 585
R3022 gnd.n4215 gnd.n4188 585
R3023 gnd.n4218 gnd.n4217 585
R3024 gnd.n4186 gnd.n4185 585
R3025 gnd.n4223 gnd.n4222 585
R3026 gnd.n4225 gnd.n4184 585
R3027 gnd.n4228 gnd.n4227 585
R3028 gnd.n4182 gnd.n4181 585
R3029 gnd.n4233 gnd.n4232 585
R3030 gnd.n4235 gnd.n4177 585
R3031 gnd.n4238 gnd.n4237 585
R3032 gnd.n4175 gnd.n4174 585
R3033 gnd.n4243 gnd.n4242 585
R3034 gnd.n4245 gnd.n4173 585
R3035 gnd.n4248 gnd.n4247 585
R3036 gnd.n4171 gnd.n4170 585
R3037 gnd.n4253 gnd.n4252 585
R3038 gnd.n4255 gnd.n4169 585
R3039 gnd.n4258 gnd.n4257 585
R3040 gnd.n4167 gnd.n4166 585
R3041 gnd.n4263 gnd.n4262 585
R3042 gnd.n4265 gnd.n4165 585
R3043 gnd.n4268 gnd.n4267 585
R3044 gnd.n4163 gnd.n4162 585
R3045 gnd.n4273 gnd.n4272 585
R3046 gnd.n4275 gnd.n4161 585
R3047 gnd.n4278 gnd.n4277 585
R3048 gnd.n4159 gnd.n4158 585
R3049 gnd.n4284 gnd.n4283 585
R3050 gnd.n4286 gnd.n4157 585
R3051 gnd.n4287 gnd.n4156 585
R3052 gnd.n4290 gnd.n4289 585
R3053 gnd.n4824 gnd.n4823 585
R3054 gnd.n4822 gnd.n4765 585
R3055 gnd.n4821 gnd.n4820 585
R3056 gnd.n4814 gnd.n4766 585
R3057 gnd.n4816 gnd.n4815 585
R3058 gnd.n4813 gnd.n4812 585
R3059 gnd.n4811 gnd.n4810 585
R3060 gnd.n4804 gnd.n4768 585
R3061 gnd.n4806 gnd.n4805 585
R3062 gnd.n4803 gnd.n4802 585
R3063 gnd.n4801 gnd.n4800 585
R3064 gnd.n4794 gnd.n4770 585
R3065 gnd.n4796 gnd.n4795 585
R3066 gnd.n4793 gnd.n4792 585
R3067 gnd.n4791 gnd.n4790 585
R3068 gnd.n4784 gnd.n4772 585
R3069 gnd.n4786 gnd.n4785 585
R3070 gnd.n4783 gnd.n4782 585
R3071 gnd.n4781 gnd.n4780 585
R3072 gnd.n4776 gnd.n4775 585
R3073 gnd.n4774 gnd.n1296 585
R3074 gnd.n6550 gnd.n6549 585
R3075 gnd.n6552 gnd.n6551 585
R3076 gnd.n6554 gnd.n6553 585
R3077 gnd.n6556 gnd.n6555 585
R3078 gnd.n6558 gnd.n6557 585
R3079 gnd.n6560 gnd.n6559 585
R3080 gnd.n6562 gnd.n6561 585
R3081 gnd.n6564 gnd.n6563 585
R3082 gnd.n6566 gnd.n6565 585
R3083 gnd.n6568 gnd.n6567 585
R3084 gnd.n6570 gnd.n6569 585
R3085 gnd.n6572 gnd.n6571 585
R3086 gnd.n6573 gnd.n1281 585
R3087 gnd.n6575 gnd.n6574 585
R3088 gnd.n1250 gnd.n1249 585
R3089 gnd.n6579 gnd.n6578 585
R3090 gnd.n6578 gnd.n6577 585
R3091 gnd.n4827 gnd.n2460 585
R3092 gnd.n4923 gnd.n2460 585
R3093 gnd.n4828 gnd.n1242 585
R3094 gnd.n6585 gnd.n1242 585
R3095 gnd.n4830 gnd.n4829 585
R3096 gnd.n4831 gnd.n4830 585
R3097 gnd.n2485 gnd.n1231 585
R3098 gnd.n6591 gnd.n1231 585
R3099 gnd.n4757 gnd.n4756 585
R3100 gnd.n4756 gnd.n4755 585
R3101 gnd.n4754 gnd.n1220 585
R3102 gnd.n6597 gnd.n1220 585
R3103 gnd.n4753 gnd.n4752 585
R3104 gnd.n4752 gnd.n4751 585
R3105 gnd.n2487 gnd.n1209 585
R3106 gnd.n6603 gnd.n1209 585
R3107 gnd.n4747 gnd.n4746 585
R3108 gnd.n4746 gnd.n4745 585
R3109 gnd.n4744 gnd.n1198 585
R3110 gnd.n6609 gnd.n1198 585
R3111 gnd.n4743 gnd.n2475 585
R3112 gnd.n4888 gnd.n2475 585
R3113 gnd.n2489 gnd.n1188 585
R3114 gnd.n6615 gnd.n1188 585
R3115 gnd.n4739 gnd.n4738 585
R3116 gnd.n4738 gnd.n4737 585
R3117 gnd.n2491 gnd.n1177 585
R3118 gnd.n6621 gnd.n1177 585
R3119 gnd.n4728 gnd.n4727 585
R3120 gnd.n4729 gnd.n4728 585
R3121 gnd.n2495 gnd.n1166 585
R3122 gnd.n6627 gnd.n1166 585
R3123 gnd.n4723 gnd.n4722 585
R3124 gnd.n4722 gnd.n4721 585
R3125 gnd.n2497 gnd.n1155 585
R3126 gnd.n6633 gnd.n1155 585
R3127 gnd.n4658 gnd.n2501 585
R3128 gnd.n4713 gnd.n2501 585
R3129 gnd.n4659 gnd.n1145 585
R3130 gnd.n6639 gnd.n1145 585
R3131 gnd.n4661 gnd.n4660 585
R3132 gnd.n4662 gnd.n4661 585
R3133 gnd.n2521 gnd.n1134 585
R3134 gnd.n6645 gnd.n1134 585
R3135 gnd.n4652 gnd.n4651 585
R3136 gnd.n4651 gnd.n4650 585
R3137 gnd.n4649 gnd.n1123 585
R3138 gnd.n6651 gnd.n1123 585
R3139 gnd.n4648 gnd.n4647 585
R3140 gnd.n4647 gnd.n4646 585
R3141 gnd.n2523 gnd.n1113 585
R3142 gnd.n6657 gnd.n1113 585
R3143 gnd.n4642 gnd.n2513 585
R3144 gnd.n4676 gnd.n2513 585
R3145 gnd.n4641 gnd.n1102 585
R3146 gnd.n6663 gnd.n1102 585
R3147 gnd.n4640 gnd.n4639 585
R3148 gnd.n4639 gnd.n4638 585
R3149 gnd.n2527 gnd.n2525 585
R3150 gnd.n4625 gnd.n2527 585
R3151 gnd.n2568 gnd.n2533 585
R3152 gnd.n4630 gnd.n2533 585
R3153 gnd.n2569 gnd.n2543 585
R3154 gnd.n4616 gnd.n2543 585
R3155 gnd.n2570 gnd.n2549 585
R3156 gnd.n4597 gnd.n2549 585
R3157 gnd.n2572 gnd.n2571 585
R3158 gnd.n2571 gnd.n2548 585
R3159 gnd.n2573 gnd.n2552 585
R3160 gnd.n4590 gnd.n2552 585
R3161 gnd.n4565 gnd.n4564 585
R3162 gnd.n4564 gnd.n4563 585
R3163 gnd.n4566 gnd.n1087 585
R3164 gnd.n6671 gnd.n1087 585
R3165 gnd.n4568 gnd.n4567 585
R3166 gnd.n4569 gnd.n4568 585
R3167 gnd.n2558 gnd.n1076 585
R3168 gnd.n6677 gnd.n1076 585
R3169 gnd.n4538 gnd.n2579 585
R3170 gnd.n4551 gnd.n2579 585
R3171 gnd.n4539 gnd.n1066 585
R3172 gnd.n6683 gnd.n1066 585
R3173 gnd.n4541 gnd.n4540 585
R3174 gnd.n4542 gnd.n4541 585
R3175 gnd.n2583 gnd.n1055 585
R3176 gnd.n6689 gnd.n1055 585
R3177 gnd.n4531 gnd.n4530 585
R3178 gnd.n4530 gnd.n4529 585
R3179 gnd.n2585 gnd.n1045 585
R3180 gnd.n6695 gnd.n1045 585
R3181 gnd.n4520 gnd.n4519 585
R3182 gnd.n4521 gnd.n4520 585
R3183 gnd.n2613 gnd.n1033 585
R3184 gnd.n6701 gnd.n1033 585
R3185 gnd.n4515 gnd.n4514 585
R3186 gnd.n4514 gnd.n1022 585
R3187 gnd.n4513 gnd.n1020 585
R3188 gnd.n6707 gnd.n1020 585
R3189 gnd.n4512 gnd.n4511 585
R3190 gnd.n4511 gnd.n1019 585
R3191 gnd.n4510 gnd.n2615 585
R3192 gnd.n4510 gnd.n4509 585
R3193 gnd.n4304 gnd.n2617 585
R3194 gnd.n2618 gnd.n2617 585
R3195 gnd.n4305 gnd.n2627 585
R3196 gnd.n4500 gnd.n2627 585
R3197 gnd.n4307 gnd.n4306 585
R3198 gnd.n4306 gnd.n2626 585
R3199 gnd.n4308 gnd.n2635 585
R3200 gnd.n4482 gnd.n2635 585
R3201 gnd.n4310 gnd.n4309 585
R3202 gnd.n4309 gnd.n2645 585
R3203 gnd.n4311 gnd.n2643 585
R3204 gnd.n4474 gnd.n2643 585
R3205 gnd.n4313 gnd.n4312 585
R3206 gnd.n4312 gnd.n2642 585
R3207 gnd.n4314 gnd.n2652 585
R3208 gnd.n4466 gnd.n2652 585
R3209 gnd.n4316 gnd.n4315 585
R3210 gnd.n4315 gnd.n2651 585
R3211 gnd.n4317 gnd.n2660 585
R3212 gnd.n4458 gnd.n2660 585
R3213 gnd.n4319 gnd.n4318 585
R3214 gnd.n4318 gnd.n2659 585
R3215 gnd.n4152 gnd.n2667 585
R3216 gnd.n4450 gnd.n2667 585
R3217 gnd.n4324 gnd.n4323 585
R3218 gnd.n4325 gnd.n4324 585
R3219 gnd.n4151 gnd.n4149 585
R3220 gnd.n4442 gnd.n4149 585
R3221 gnd.n7916 gnd.n7915 585
R3222 gnd.n7917 gnd.n7916 585
R3223 gnd.n132 gnd.n130 585
R3224 gnd.n7838 gnd.n130 585
R3225 gnd.n7766 gnd.n217 585
R3226 gnd.n217 gnd.n215 585
R3227 gnd.n7768 gnd.n7767 585
R3228 gnd.n7769 gnd.n7768 585
R3229 gnd.n218 gnd.n216 585
R3230 gnd.n216 gnd.n213 585
R3231 gnd.n7761 gnd.n7760 585
R3232 gnd.n7760 gnd.n7759 585
R3233 gnd.n221 gnd.n220 585
R3234 gnd.n222 gnd.n221 585
R3235 gnd.n7750 gnd.n7749 585
R3236 gnd.n7751 gnd.n7750 585
R3237 gnd.n233 gnd.n232 585
R3238 gnd.n232 gnd.n230 585
R3239 gnd.n7745 gnd.n7744 585
R3240 gnd.n7744 gnd.n7743 585
R3241 gnd.n236 gnd.n235 585
R3242 gnd.n246 gnd.n236 585
R3243 gnd.n7734 gnd.n7733 585
R3244 gnd.n7735 gnd.n7734 585
R3245 gnd.n248 gnd.n247 585
R3246 gnd.n247 gnd.n244 585
R3247 gnd.n7729 gnd.n7728 585
R3248 gnd.n7728 gnd.n7727 585
R3249 gnd.n251 gnd.n250 585
R3250 gnd.n252 gnd.n251 585
R3251 gnd.n7718 gnd.n7717 585
R3252 gnd.n7719 gnd.n7718 585
R3253 gnd.n262 gnd.n261 585
R3254 gnd.n269 gnd.n261 585
R3255 gnd.n7713 gnd.n7712 585
R3256 gnd.n7712 gnd.n7711 585
R3257 gnd.n265 gnd.n264 585
R3258 gnd.n393 gnd.n265 585
R3259 gnd.n7702 gnd.n7701 585
R3260 gnd.n7703 gnd.n7702 585
R3261 gnd.n279 gnd.n278 585
R3262 gnd.n398 gnd.n278 585
R3263 gnd.n7697 gnd.n7696 585
R3264 gnd.n7696 gnd.n7695 585
R3265 gnd.n282 gnd.n281 585
R3266 gnd.n7624 gnd.n282 585
R3267 gnd.n7686 gnd.n7685 585
R3268 gnd.n7687 gnd.n7686 585
R3269 gnd.n294 gnd.n293 585
R3270 gnd.n7629 gnd.n293 585
R3271 gnd.n7681 gnd.n7680 585
R3272 gnd.n7680 gnd.n7679 585
R3273 gnd.n297 gnd.n296 585
R3274 gnd.n7633 gnd.n297 585
R3275 gnd.n7670 gnd.n7669 585
R3276 gnd.n7671 gnd.n7670 585
R3277 gnd.n310 gnd.n309 585
R3278 gnd.n7638 gnd.n309 585
R3279 gnd.n7648 gnd.n7647 585
R3280 gnd.n7649 gnd.n7648 585
R3281 gnd.n7646 gnd.n7645 585
R3282 gnd.n7645 gnd.n7644 585
R3283 gnd.n1534 gnd.n338 585
R3284 gnd.n1537 gnd.n338 585
R3285 gnd.n6286 gnd.n1535 585
R3286 gnd.n6286 gnd.n6285 585
R3287 gnd.n6289 gnd.n6288 585
R3288 gnd.n6290 gnd.n6289 585
R3289 gnd.n6287 gnd.n319 585
R3290 gnd.n6186 gnd.n319 585
R3291 gnd.n7665 gnd.n7664 585
R3292 gnd.n7664 gnd.n7663 585
R3293 gnd.n7666 gnd.n318 585
R3294 gnd.n6190 gnd.n318 585
R3295 gnd.n6304 gnd.n317 585
R3296 gnd.n6305 gnd.n6304 585
R3297 gnd.n6303 gnd.n1520 585
R3298 gnd.n6303 gnd.n6302 585
R3299 gnd.n6239 gnd.n1519 585
R3300 gnd.n6195 gnd.n1519 585
R3301 gnd.n6241 gnd.n6240 585
R3302 gnd.n6242 gnd.n6241 585
R3303 gnd.n1554 gnd.n1553 585
R3304 gnd.n1553 gnd.n1549 585
R3305 gnd.n6234 gnd.n6233 585
R3306 gnd.n6233 gnd.n6232 585
R3307 gnd.n1557 gnd.n1556 585
R3308 gnd.n6204 gnd.n1557 585
R3309 gnd.n6219 gnd.n6218 585
R3310 gnd.n6220 gnd.n6219 585
R3311 gnd.n1570 gnd.n1569 585
R3312 gnd.n1578 gnd.n1569 585
R3313 gnd.n6214 gnd.n6213 585
R3314 gnd.n6213 gnd.n6212 585
R3315 gnd.n1573 gnd.n1572 585
R3316 gnd.n6163 gnd.n1573 585
R3317 gnd.n6151 gnd.n1606 585
R3318 gnd.n1606 gnd.n1605 585
R3319 gnd.n6153 gnd.n6152 585
R3320 gnd.n6154 gnd.n6153 585
R3321 gnd.n1607 gnd.n1604 585
R3322 gnd.n1614 gnd.n1604 585
R3323 gnd.n6146 gnd.n6145 585
R3324 gnd.n6145 gnd.n6144 585
R3325 gnd.n1610 gnd.n1609 585
R3326 gnd.n6125 gnd.n1610 585
R3327 gnd.n6113 gnd.n1634 585
R3328 gnd.n1634 gnd.n1622 585
R3329 gnd.n6115 gnd.n6114 585
R3330 gnd.n6116 gnd.n6115 585
R3331 gnd.n1635 gnd.n1633 585
R3332 gnd.n1642 gnd.n1633 585
R3333 gnd.n6108 gnd.n6107 585
R3334 gnd.n6107 gnd.n6106 585
R3335 gnd.n1638 gnd.n1637 585
R3336 gnd.n6094 gnd.n1638 585
R3337 gnd.n6081 gnd.n1660 585
R3338 gnd.n1931 gnd.n1660 585
R3339 gnd.n6083 gnd.n6082 585
R3340 gnd.n6084 gnd.n6083 585
R3341 gnd.n1661 gnd.n1659 585
R3342 gnd.n1668 gnd.n1659 585
R3343 gnd.n6076 gnd.n6075 585
R3344 gnd.n6075 gnd.n6074 585
R3345 gnd.n1664 gnd.n1663 585
R3346 gnd.n6061 gnd.n1664 585
R3347 gnd.n6049 gnd.n1686 585
R3348 gnd.n1686 gnd.n1675 585
R3349 gnd.n6051 gnd.n6050 585
R3350 gnd.n6052 gnd.n6051 585
R3351 gnd.n6045 gnd.n1685 585
R3352 gnd.n6044 gnd.n6043 585
R3353 gnd.n1689 gnd.n1688 585
R3354 gnd.n6041 gnd.n1689 585
R3355 gnd.n1843 gnd.n1842 585
R3356 gnd.n1848 gnd.n1847 585
R3357 gnd.n1850 gnd.n1849 585
R3358 gnd.n1853 gnd.n1852 585
R3359 gnd.n1851 gnd.n1840 585
R3360 gnd.n1858 gnd.n1857 585
R3361 gnd.n1860 gnd.n1859 585
R3362 gnd.n1863 gnd.n1862 585
R3363 gnd.n1861 gnd.n1838 585
R3364 gnd.n1868 gnd.n1867 585
R3365 gnd.n1870 gnd.n1869 585
R3366 gnd.n1873 gnd.n1872 585
R3367 gnd.n1871 gnd.n1835 585
R3368 gnd.n1983 gnd.n1982 585
R3369 gnd.n1981 gnd.n1980 585
R3370 gnd.n1979 gnd.n1978 585
R3371 gnd.n1977 gnd.n1976 585
R3372 gnd.n1975 gnd.n1974 585
R3373 gnd.n1973 gnd.n1972 585
R3374 gnd.n1971 gnd.n1970 585
R3375 gnd.n1969 gnd.n1968 585
R3376 gnd.n1967 gnd.n1966 585
R3377 gnd.n1965 gnd.n1964 585
R3378 gnd.n1963 gnd.n1962 585
R3379 gnd.n1961 gnd.n1960 585
R3380 gnd.n1959 gnd.n1958 585
R3381 gnd.n1957 gnd.n1956 585
R3382 gnd.n1955 gnd.n1954 585
R3383 gnd.n1953 gnd.n1952 585
R3384 gnd.n1951 gnd.n1950 585
R3385 gnd.n1949 gnd.n1948 585
R3386 gnd.n1947 gnd.n1897 585
R3387 gnd.n1901 gnd.n1898 585
R3388 gnd.n1943 gnd.n1942 585
R3389 gnd.n200 gnd.n199 585
R3390 gnd.n7845 gnd.n195 585
R3391 gnd.n7847 gnd.n7846 585
R3392 gnd.n7849 gnd.n193 585
R3393 gnd.n7851 gnd.n7850 585
R3394 gnd.n7852 gnd.n188 585
R3395 gnd.n7854 gnd.n7853 585
R3396 gnd.n7856 gnd.n186 585
R3397 gnd.n7858 gnd.n7857 585
R3398 gnd.n7859 gnd.n181 585
R3399 gnd.n7861 gnd.n7860 585
R3400 gnd.n7863 gnd.n179 585
R3401 gnd.n7865 gnd.n7864 585
R3402 gnd.n7866 gnd.n174 585
R3403 gnd.n7868 gnd.n7867 585
R3404 gnd.n7870 gnd.n172 585
R3405 gnd.n7872 gnd.n7871 585
R3406 gnd.n7873 gnd.n167 585
R3407 gnd.n7875 gnd.n7874 585
R3408 gnd.n7877 gnd.n165 585
R3409 gnd.n7879 gnd.n7878 585
R3410 gnd.n7883 gnd.n160 585
R3411 gnd.n7885 gnd.n7884 585
R3412 gnd.n7887 gnd.n158 585
R3413 gnd.n7889 gnd.n7888 585
R3414 gnd.n7890 gnd.n153 585
R3415 gnd.n7892 gnd.n7891 585
R3416 gnd.n7894 gnd.n151 585
R3417 gnd.n7896 gnd.n7895 585
R3418 gnd.n7897 gnd.n146 585
R3419 gnd.n7899 gnd.n7898 585
R3420 gnd.n7901 gnd.n144 585
R3421 gnd.n7903 gnd.n7902 585
R3422 gnd.n7904 gnd.n139 585
R3423 gnd.n7906 gnd.n7905 585
R3424 gnd.n7908 gnd.n137 585
R3425 gnd.n7910 gnd.n7909 585
R3426 gnd.n7911 gnd.n135 585
R3427 gnd.n7912 gnd.n131 585
R3428 gnd.n131 gnd.n128 585
R3429 gnd.n7841 gnd.n127 585
R3430 gnd.n7917 gnd.n127 585
R3431 gnd.n7840 gnd.n7839 585
R3432 gnd.n7839 gnd.n7838 585
R3433 gnd.n205 gnd.n204 585
R3434 gnd.n215 gnd.n205 585
R3435 gnd.n371 gnd.n214 585
R3436 gnd.n7769 gnd.n214 585
R3437 gnd.n373 gnd.n372 585
R3438 gnd.n372 gnd.n213 585
R3439 gnd.n374 gnd.n223 585
R3440 gnd.n7759 gnd.n223 585
R3441 gnd.n376 gnd.n375 585
R3442 gnd.n375 gnd.n222 585
R3443 gnd.n377 gnd.n231 585
R3444 gnd.n7751 gnd.n231 585
R3445 gnd.n379 gnd.n378 585
R3446 gnd.n378 gnd.n230 585
R3447 gnd.n380 gnd.n237 585
R3448 gnd.n7743 gnd.n237 585
R3449 gnd.n382 gnd.n381 585
R3450 gnd.n381 gnd.n246 585
R3451 gnd.n383 gnd.n245 585
R3452 gnd.n7735 gnd.n245 585
R3453 gnd.n385 gnd.n384 585
R3454 gnd.n384 gnd.n244 585
R3455 gnd.n386 gnd.n253 585
R3456 gnd.n7727 gnd.n253 585
R3457 gnd.n388 gnd.n387 585
R3458 gnd.n387 gnd.n252 585
R3459 gnd.n389 gnd.n260 585
R3460 gnd.n7719 gnd.n260 585
R3461 gnd.n391 gnd.n390 585
R3462 gnd.n390 gnd.n269 585
R3463 gnd.n392 gnd.n267 585
R3464 gnd.n7711 gnd.n267 585
R3465 gnd.n395 gnd.n394 585
R3466 gnd.n394 gnd.n393 585
R3467 gnd.n396 gnd.n276 585
R3468 gnd.n7703 gnd.n276 585
R3469 gnd.n400 gnd.n399 585
R3470 gnd.n399 gnd.n398 585
R3471 gnd.n401 gnd.n284 585
R3472 gnd.n7695 gnd.n284 585
R3473 gnd.n7626 gnd.n7625 585
R3474 gnd.n7625 gnd.n7624 585
R3475 gnd.n7627 gnd.n292 585
R3476 gnd.n7687 gnd.n292 585
R3477 gnd.n7631 gnd.n7630 585
R3478 gnd.n7630 gnd.n7629 585
R3479 gnd.n7632 gnd.n299 585
R3480 gnd.n7679 gnd.n299 585
R3481 gnd.n7635 gnd.n7634 585
R3482 gnd.n7634 gnd.n7633 585
R3483 gnd.n7636 gnd.n307 585
R3484 gnd.n7671 gnd.n307 585
R3485 gnd.n7640 gnd.n7639 585
R3486 gnd.n7639 gnd.n7638 585
R3487 gnd.n7641 gnd.n336 585
R3488 gnd.n7649 gnd.n336 585
R3489 gnd.n7643 gnd.n7642 585
R3490 gnd.n7644 gnd.n7643 585
R3491 gnd.n341 gnd.n340 585
R3492 gnd.n1537 gnd.n340 585
R3493 gnd.n6184 gnd.n1536 585
R3494 gnd.n6285 gnd.n1536 585
R3495 gnd.n6185 gnd.n1532 585
R3496 gnd.n6290 gnd.n1532 585
R3497 gnd.n6188 gnd.n6187 585
R3498 gnd.n6187 gnd.n6186 585
R3499 gnd.n6189 gnd.n321 585
R3500 gnd.n7663 gnd.n321 585
R3501 gnd.n6192 gnd.n6191 585
R3502 gnd.n6191 gnd.n6190 585
R3503 gnd.n6193 gnd.n1516 585
R3504 gnd.n6305 gnd.n1516 585
R3505 gnd.n6194 gnd.n1522 585
R3506 gnd.n6302 gnd.n1522 585
R3507 gnd.n6197 gnd.n6196 585
R3508 gnd.n6196 gnd.n6195 585
R3509 gnd.n6198 gnd.n1550 585
R3510 gnd.n6242 gnd.n1550 585
R3511 gnd.n6200 gnd.n6199 585
R3512 gnd.n6199 gnd.n1549 585
R3513 gnd.n6201 gnd.n1559 585
R3514 gnd.n6232 gnd.n1559 585
R3515 gnd.n6203 gnd.n6202 585
R3516 gnd.n6204 gnd.n6203 585
R3517 gnd.n1588 gnd.n1568 585
R3518 gnd.n6220 gnd.n1568 585
R3519 gnd.n6168 gnd.n6167 585
R3520 gnd.n6167 gnd.n1578 585
R3521 gnd.n6166 gnd.n1575 585
R3522 gnd.n6212 gnd.n1575 585
R3523 gnd.n6165 gnd.n6164 585
R3524 gnd.n6164 gnd.n6163 585
R3525 gnd.n1592 gnd.n1590 585
R3526 gnd.n1605 gnd.n1592 585
R3527 gnd.n1919 gnd.n1601 585
R3528 gnd.n6154 gnd.n1601 585
R3529 gnd.n1921 gnd.n1920 585
R3530 gnd.n1920 gnd.n1614 585
R3531 gnd.n1922 gnd.n1612 585
R3532 gnd.n6144 gnd.n1612 585
R3533 gnd.n1923 gnd.n1623 585
R3534 gnd.n6125 gnd.n1623 585
R3535 gnd.n1925 gnd.n1924 585
R3536 gnd.n1924 gnd.n1622 585
R3537 gnd.n1926 gnd.n1631 585
R3538 gnd.n6116 gnd.n1631 585
R3539 gnd.n1928 gnd.n1927 585
R3540 gnd.n1927 gnd.n1642 585
R3541 gnd.n1929 gnd.n1640 585
R3542 gnd.n6106 gnd.n1640 585
R3543 gnd.n1930 gnd.n1649 585
R3544 gnd.n6094 gnd.n1649 585
R3545 gnd.n1933 gnd.n1932 585
R3546 gnd.n1932 gnd.n1931 585
R3547 gnd.n1934 gnd.n1657 585
R3548 gnd.n6084 gnd.n1657 585
R3549 gnd.n1936 gnd.n1935 585
R3550 gnd.n1935 gnd.n1668 585
R3551 gnd.n1937 gnd.n1666 585
R3552 gnd.n6074 gnd.n1666 585
R3553 gnd.n1938 gnd.n1676 585
R3554 gnd.n6061 gnd.n1676 585
R3555 gnd.n1939 gnd.n1903 585
R3556 gnd.n1903 gnd.n1675 585
R3557 gnd.n1940 gnd.n1683 585
R3558 gnd.n6052 gnd.n1683 585
R3559 gnd.n5683 gnd.n1994 585
R3560 gnd.n1994 gnd.n1799 585
R3561 gnd.n5685 gnd.n5684 585
R3562 gnd.n5686 gnd.n5685 585
R3563 gnd.n5594 gnd.n1993 585
R3564 gnd.n1993 gnd.n1991 585
R3565 gnd.n5593 gnd.n5592 585
R3566 gnd.n5592 gnd.n5591 585
R3567 gnd.n1996 gnd.n1995 585
R3568 gnd.n5566 gnd.n1996 585
R3569 gnd.n5579 gnd.n5578 585
R3570 gnd.n5580 gnd.n5579 585
R3571 gnd.n5577 gnd.n2007 585
R3572 gnd.n5572 gnd.n2007 585
R3573 gnd.n5576 gnd.n5575 585
R3574 gnd.n5575 gnd.n5574 585
R3575 gnd.n2009 gnd.n2008 585
R3576 gnd.n5560 gnd.n2009 585
R3577 gnd.n5545 gnd.n5544 585
R3578 gnd.n5544 gnd.n2014 585
R3579 gnd.n5546 gnd.n2025 585
R3580 gnd.n2025 gnd.n2023 585
R3581 gnd.n5548 gnd.n5547 585
R3582 gnd.n5549 gnd.n5548 585
R3583 gnd.n5543 gnd.n2024 585
R3584 gnd.n5538 gnd.n2024 585
R3585 gnd.n5542 gnd.n5541 585
R3586 gnd.n5541 gnd.n5540 585
R3587 gnd.n2027 gnd.n2026 585
R3588 gnd.n2028 gnd.n2027 585
R3589 gnd.n5527 gnd.n5526 585
R3590 gnd.n5528 gnd.n5527 585
R3591 gnd.n5525 gnd.n2034 585
R3592 gnd.n5521 gnd.n2034 585
R3593 gnd.n5524 gnd.n5523 585
R3594 gnd.n5523 gnd.n5522 585
R3595 gnd.n2036 gnd.n2035 585
R3596 gnd.n2043 gnd.n2036 585
R3597 gnd.n5513 gnd.n5512 585
R3598 gnd.n5514 gnd.n5513 585
R3599 gnd.n5511 gnd.n2045 585
R3600 gnd.n2045 gnd.n2042 585
R3601 gnd.n5510 gnd.n5509 585
R3602 gnd.n5509 gnd.n5508 585
R3603 gnd.n2047 gnd.n2046 585
R3604 gnd.n2071 gnd.n2047 585
R3605 gnd.n5446 gnd.n2070 585
R3606 gnd.n5460 gnd.n2070 585
R3607 gnd.n5447 gnd.n2084 585
R3608 gnd.n5435 gnd.n2084 585
R3609 gnd.n5449 gnd.n5448 585
R3610 gnd.n5450 gnd.n5449 585
R3611 gnd.n5445 gnd.n2083 585
R3612 gnd.n2083 gnd.n2079 585
R3613 gnd.n5444 gnd.n5443 585
R3614 gnd.n5443 gnd.n5442 585
R3615 gnd.n2086 gnd.n2085 585
R3616 gnd.n2092 gnd.n2086 585
R3617 gnd.n5426 gnd.n5425 585
R3618 gnd.n5427 gnd.n5426 585
R3619 gnd.n5424 gnd.n2095 585
R3620 gnd.n2101 gnd.n2095 585
R3621 gnd.n5423 gnd.n5422 585
R3622 gnd.n5422 gnd.n5421 585
R3623 gnd.n2097 gnd.n2096 585
R3624 gnd.n5338 gnd.n2097 585
R3625 gnd.n5408 gnd.n5407 585
R3626 gnd.n5409 gnd.n5408 585
R3627 gnd.n5406 gnd.n2111 585
R3628 gnd.n2111 gnd.n2108 585
R3629 gnd.n5405 gnd.n5404 585
R3630 gnd.n5404 gnd.n5403 585
R3631 gnd.n2113 gnd.n2112 585
R3632 gnd.n2114 gnd.n2113 585
R3633 gnd.n5361 gnd.n5360 585
R3634 gnd.n5361 gnd.n2123 585
R3635 gnd.n5363 gnd.n5362 585
R3636 gnd.n5362 gnd.n2122 585
R3637 gnd.n5364 gnd.n2136 585
R3638 gnd.n5349 gnd.n2136 585
R3639 gnd.n5366 gnd.n5365 585
R3640 gnd.n5367 gnd.n5366 585
R3641 gnd.n5359 gnd.n2135 585
R3642 gnd.n2135 gnd.n2131 585
R3643 gnd.n5358 gnd.n5357 585
R3644 gnd.n5357 gnd.n5356 585
R3645 gnd.n2138 gnd.n2137 585
R3646 gnd.n2144 gnd.n2138 585
R3647 gnd.n5330 gnd.n5329 585
R3648 gnd.n5331 gnd.n5330 585
R3649 gnd.n5328 gnd.n2146 585
R3650 gnd.n2153 gnd.n2146 585
R3651 gnd.n5327 gnd.n5326 585
R3652 gnd.n5326 gnd.n5325 585
R3653 gnd.n2148 gnd.n2147 585
R3654 gnd.n2164 gnd.n2148 585
R3655 gnd.n5302 gnd.n2161 585
R3656 gnd.n5314 gnd.n2161 585
R3657 gnd.n5303 gnd.n2170 585
R3658 gnd.n2170 gnd.n2160 585
R3659 gnd.n5305 gnd.n5304 585
R3660 gnd.n5306 gnd.n5305 585
R3661 gnd.n5301 gnd.n2169 585
R3662 gnd.n5297 gnd.n2169 585
R3663 gnd.n5300 gnd.n5299 585
R3664 gnd.n5299 gnd.n5298 585
R3665 gnd.n2172 gnd.n2171 585
R3666 gnd.n5287 gnd.n2172 585
R3667 gnd.n5277 gnd.n2189 585
R3668 gnd.n2189 gnd.n2182 585
R3669 gnd.n5279 gnd.n5278 585
R3670 gnd.n5280 gnd.n5279 585
R3671 gnd.n5276 gnd.n2188 585
R3672 gnd.n2195 gnd.n2188 585
R3673 gnd.n5275 gnd.n5274 585
R3674 gnd.n5274 gnd.n5273 585
R3675 gnd.n2191 gnd.n2190 585
R3676 gnd.n2192 gnd.n2191 585
R3677 gnd.n5262 gnd.n5261 585
R3678 gnd.n5263 gnd.n5262 585
R3679 gnd.n5260 gnd.n2205 585
R3680 gnd.n5256 gnd.n2205 585
R3681 gnd.n5259 gnd.n5258 585
R3682 gnd.n5258 gnd.n5257 585
R3683 gnd.n2207 gnd.n2206 585
R3684 gnd.n5246 gnd.n2207 585
R3685 gnd.n5107 gnd.n5106 585
R3686 gnd.n5107 gnd.n2212 585
R3687 gnd.n5189 gnd.n5105 585
R3688 gnd.n5189 gnd.n5188 585
R3689 gnd.n5191 gnd.n5190 585
R3690 gnd.n5190 gnd.n1378 585
R3691 gnd.n5192 gnd.n5103 585
R3692 gnd.n5103 gnd.n1376 585
R3693 gnd.n5194 gnd.n5193 585
R3694 gnd.n5195 gnd.n5194 585
R3695 gnd.n5104 gnd.n5102 585
R3696 gnd.n5102 gnd.n1366 585
R3697 gnd.n1361 gnd.n1360 585
R3698 gnd.n6473 gnd.n1361 585
R3699 gnd.n6476 gnd.n6475 585
R3700 gnd.n6475 gnd.n6474 585
R3701 gnd.n6477 gnd.n1339 585
R3702 gnd.n5175 gnd.n1339 585
R3703 gnd.n6542 gnd.n6541 585
R3704 gnd.n6540 gnd.n1338 585
R3705 gnd.n6539 gnd.n1337 585
R3706 gnd.n6544 gnd.n1337 585
R3707 gnd.n6538 gnd.n6537 585
R3708 gnd.n6536 gnd.n6535 585
R3709 gnd.n6534 gnd.n6533 585
R3710 gnd.n6532 gnd.n6531 585
R3711 gnd.n6530 gnd.n6529 585
R3712 gnd.n6528 gnd.n6527 585
R3713 gnd.n6526 gnd.n6525 585
R3714 gnd.n6524 gnd.n6523 585
R3715 gnd.n6522 gnd.n6521 585
R3716 gnd.n6520 gnd.n6519 585
R3717 gnd.n6518 gnd.n6517 585
R3718 gnd.n6516 gnd.n6515 585
R3719 gnd.n6514 gnd.n6513 585
R3720 gnd.n6512 gnd.n6511 585
R3721 gnd.n6510 gnd.n6509 585
R3722 gnd.n6508 gnd.n6507 585
R3723 gnd.n6506 gnd.n6505 585
R3724 gnd.n6504 gnd.n6503 585
R3725 gnd.n6502 gnd.n6501 585
R3726 gnd.n6500 gnd.n6499 585
R3727 gnd.n6498 gnd.n6497 585
R3728 gnd.n6496 gnd.n6495 585
R3729 gnd.n6494 gnd.n6493 585
R3730 gnd.n6492 gnd.n6491 585
R3731 gnd.n6490 gnd.n6489 585
R3732 gnd.n6488 gnd.n6487 585
R3733 gnd.n6486 gnd.n6485 585
R3734 gnd.n6484 gnd.n6483 585
R3735 gnd.n6482 gnd.n1302 585
R3736 gnd.n6547 gnd.n6546 585
R3737 gnd.n1304 gnd.n1301 585
R3738 gnd.n5113 gnd.n5112 585
R3739 gnd.n5115 gnd.n5114 585
R3740 gnd.n5118 gnd.n5117 585
R3741 gnd.n5120 gnd.n5119 585
R3742 gnd.n5122 gnd.n5121 585
R3743 gnd.n5124 gnd.n5123 585
R3744 gnd.n5126 gnd.n5125 585
R3745 gnd.n5128 gnd.n5127 585
R3746 gnd.n5130 gnd.n5129 585
R3747 gnd.n5132 gnd.n5131 585
R3748 gnd.n5134 gnd.n5133 585
R3749 gnd.n5136 gnd.n5135 585
R3750 gnd.n5138 gnd.n5137 585
R3751 gnd.n5140 gnd.n5139 585
R3752 gnd.n5142 gnd.n5141 585
R3753 gnd.n5144 gnd.n5143 585
R3754 gnd.n5146 gnd.n5145 585
R3755 gnd.n5148 gnd.n5147 585
R3756 gnd.n5150 gnd.n5149 585
R3757 gnd.n5152 gnd.n5151 585
R3758 gnd.n5154 gnd.n5153 585
R3759 gnd.n5156 gnd.n5155 585
R3760 gnd.n5158 gnd.n5157 585
R3761 gnd.n5160 gnd.n5159 585
R3762 gnd.n5162 gnd.n5161 585
R3763 gnd.n5164 gnd.n5163 585
R3764 gnd.n5166 gnd.n5165 585
R3765 gnd.n5168 gnd.n5167 585
R3766 gnd.n5170 gnd.n5169 585
R3767 gnd.n5172 gnd.n5171 585
R3768 gnd.n5174 gnd.n5173 585
R3769 gnd.n5690 gnd.n5689 585
R3770 gnd.n5692 gnd.n5691 585
R3771 gnd.n5694 gnd.n5693 585
R3772 gnd.n5696 gnd.n5695 585
R3773 gnd.n5698 gnd.n5697 585
R3774 gnd.n5700 gnd.n5699 585
R3775 gnd.n5702 gnd.n5701 585
R3776 gnd.n5704 gnd.n5703 585
R3777 gnd.n5706 gnd.n5705 585
R3778 gnd.n5708 gnd.n5707 585
R3779 gnd.n5710 gnd.n5709 585
R3780 gnd.n5712 gnd.n5711 585
R3781 gnd.n5714 gnd.n5713 585
R3782 gnd.n5716 gnd.n5715 585
R3783 gnd.n5718 gnd.n5717 585
R3784 gnd.n5720 gnd.n5719 585
R3785 gnd.n5722 gnd.n5721 585
R3786 gnd.n5724 gnd.n5723 585
R3787 gnd.n5726 gnd.n5725 585
R3788 gnd.n5728 gnd.n5727 585
R3789 gnd.n5730 gnd.n5729 585
R3790 gnd.n5732 gnd.n5731 585
R3791 gnd.n5734 gnd.n5733 585
R3792 gnd.n5736 gnd.n5735 585
R3793 gnd.n5738 gnd.n5737 585
R3794 gnd.n5740 gnd.n5739 585
R3795 gnd.n5742 gnd.n5741 585
R3796 gnd.n5744 gnd.n5743 585
R3797 gnd.n5746 gnd.n5745 585
R3798 gnd.n5749 gnd.n5748 585
R3799 gnd.n5751 gnd.n5750 585
R3800 gnd.n5753 gnd.n5752 585
R3801 gnd.n5755 gnd.n5754 585
R3802 gnd.n5616 gnd.n1985 585
R3803 gnd.n5618 gnd.n5617 585
R3804 gnd.n5620 gnd.n5619 585
R3805 gnd.n5622 gnd.n5621 585
R3806 gnd.n5625 gnd.n5624 585
R3807 gnd.n5627 gnd.n5626 585
R3808 gnd.n5629 gnd.n5628 585
R3809 gnd.n5631 gnd.n5630 585
R3810 gnd.n5633 gnd.n5632 585
R3811 gnd.n5635 gnd.n5634 585
R3812 gnd.n5637 gnd.n5636 585
R3813 gnd.n5639 gnd.n5638 585
R3814 gnd.n5641 gnd.n5640 585
R3815 gnd.n5643 gnd.n5642 585
R3816 gnd.n5645 gnd.n5644 585
R3817 gnd.n5647 gnd.n5646 585
R3818 gnd.n5649 gnd.n5648 585
R3819 gnd.n5651 gnd.n5650 585
R3820 gnd.n5653 gnd.n5652 585
R3821 gnd.n5655 gnd.n5654 585
R3822 gnd.n5657 gnd.n5656 585
R3823 gnd.n5659 gnd.n5658 585
R3824 gnd.n5661 gnd.n5660 585
R3825 gnd.n5663 gnd.n5662 585
R3826 gnd.n5665 gnd.n5664 585
R3827 gnd.n5667 gnd.n5666 585
R3828 gnd.n5669 gnd.n5668 585
R3829 gnd.n5671 gnd.n5670 585
R3830 gnd.n5673 gnd.n5672 585
R3831 gnd.n5675 gnd.n5674 585
R3832 gnd.n5677 gnd.n5676 585
R3833 gnd.n5679 gnd.n5678 585
R3834 gnd.n5681 gnd.n5680 585
R3835 gnd.n5688 gnd.n1988 585
R3836 gnd.n5688 gnd.n1799 585
R3837 gnd.n5687 gnd.n1990 585
R3838 gnd.n5687 gnd.n5686 585
R3839 gnd.n5564 gnd.n1989 585
R3840 gnd.n1991 gnd.n1989 585
R3841 gnd.n5565 gnd.n1998 585
R3842 gnd.n5591 gnd.n1998 585
R3843 gnd.n5568 gnd.n5567 585
R3844 gnd.n5567 gnd.n5566 585
R3845 gnd.n5569 gnd.n2006 585
R3846 gnd.n5580 gnd.n2006 585
R3847 gnd.n5571 gnd.n5570 585
R3848 gnd.n5572 gnd.n5571 585
R3849 gnd.n5563 gnd.n2010 585
R3850 gnd.n5574 gnd.n2010 585
R3851 gnd.n5562 gnd.n5561 585
R3852 gnd.n5561 gnd.n5560 585
R3853 gnd.n2013 gnd.n2012 585
R3854 gnd.n2014 gnd.n2013 585
R3855 gnd.n5534 gnd.n5533 585
R3856 gnd.n5533 gnd.n2023 585
R3857 gnd.n5535 gnd.n2022 585
R3858 gnd.n5549 gnd.n2022 585
R3859 gnd.n5537 gnd.n5536 585
R3860 gnd.n5538 gnd.n5537 585
R3861 gnd.n5532 gnd.n2029 585
R3862 gnd.n5540 gnd.n2029 585
R3863 gnd.n5531 gnd.n5530 585
R3864 gnd.n5530 gnd.n2028 585
R3865 gnd.n5529 gnd.n2031 585
R3866 gnd.n5529 gnd.n5528 585
R3867 gnd.n5518 gnd.n2032 585
R3868 gnd.n5521 gnd.n2032 585
R3869 gnd.n5520 gnd.n5519 585
R3870 gnd.n5522 gnd.n5520 585
R3871 gnd.n5517 gnd.n2039 585
R3872 gnd.n2043 gnd.n2039 585
R3873 gnd.n5516 gnd.n5515 585
R3874 gnd.n5515 gnd.n5514 585
R3875 gnd.n2041 gnd.n2040 585
R3876 gnd.n2042 gnd.n2041 585
R3877 gnd.n5431 gnd.n2049 585
R3878 gnd.n5508 gnd.n2049 585
R3879 gnd.n5433 gnd.n5432 585
R3880 gnd.n5432 gnd.n2071 585
R3881 gnd.n5434 gnd.n2073 585
R3882 gnd.n5460 gnd.n2073 585
R3883 gnd.n5437 gnd.n5436 585
R3884 gnd.n5436 gnd.n5435 585
R3885 gnd.n5438 gnd.n2081 585
R3886 gnd.n5450 gnd.n2081 585
R3887 gnd.n5439 gnd.n2089 585
R3888 gnd.n2089 gnd.n2079 585
R3889 gnd.n5441 gnd.n5440 585
R3890 gnd.n5442 gnd.n5441 585
R3891 gnd.n5430 gnd.n2088 585
R3892 gnd.n2092 gnd.n2088 585
R3893 gnd.n5429 gnd.n5428 585
R3894 gnd.n5428 gnd.n5427 585
R3895 gnd.n2091 gnd.n2090 585
R3896 gnd.n2101 gnd.n2091 585
R3897 gnd.n5337 gnd.n2099 585
R3898 gnd.n5421 gnd.n2099 585
R3899 gnd.n5340 gnd.n5339 585
R3900 gnd.n5339 gnd.n5338 585
R3901 gnd.n5341 gnd.n2110 585
R3902 gnd.n5409 gnd.n2110 585
R3903 gnd.n5343 gnd.n5342 585
R3904 gnd.n5342 gnd.n2108 585
R3905 gnd.n5344 gnd.n2115 585
R3906 gnd.n5403 gnd.n2115 585
R3907 gnd.n5345 gnd.n5336 585
R3908 gnd.n5336 gnd.n2114 585
R3909 gnd.n5347 gnd.n5346 585
R3910 gnd.n5347 gnd.n2123 585
R3911 gnd.n5348 gnd.n5335 585
R3912 gnd.n5348 gnd.n2122 585
R3913 gnd.n5351 gnd.n5350 585
R3914 gnd.n5350 gnd.n5349 585
R3915 gnd.n5352 gnd.n2133 585
R3916 gnd.n5367 gnd.n2133 585
R3917 gnd.n5353 gnd.n2141 585
R3918 gnd.n2141 gnd.n2131 585
R3919 gnd.n5355 gnd.n5354 585
R3920 gnd.n5356 gnd.n5355 585
R3921 gnd.n5334 gnd.n2140 585
R3922 gnd.n2144 gnd.n2140 585
R3923 gnd.n5333 gnd.n5332 585
R3924 gnd.n5332 gnd.n5331 585
R3925 gnd.n2143 gnd.n2142 585
R3926 gnd.n2153 gnd.n2143 585
R3927 gnd.n5310 gnd.n2151 585
R3928 gnd.n5325 gnd.n2151 585
R3929 gnd.n5311 gnd.n2165 585
R3930 gnd.n2165 gnd.n2164 585
R3931 gnd.n5313 gnd.n5312 585
R3932 gnd.n5314 gnd.n5313 585
R3933 gnd.n5309 gnd.n2163 585
R3934 gnd.n2163 gnd.n2160 585
R3935 gnd.n5308 gnd.n5307 585
R3936 gnd.n5307 gnd.n5306 585
R3937 gnd.n2167 gnd.n2166 585
R3938 gnd.n5297 gnd.n2167 585
R3939 gnd.n5284 gnd.n2175 585
R3940 gnd.n5298 gnd.n2175 585
R3941 gnd.n5286 gnd.n5285 585
R3942 gnd.n5287 gnd.n5286 585
R3943 gnd.n5283 gnd.n2184 585
R3944 gnd.n2184 gnd.n2182 585
R3945 gnd.n5282 gnd.n5281 585
R3946 gnd.n5281 gnd.n5280 585
R3947 gnd.n2186 gnd.n2185 585
R3948 gnd.n2195 gnd.n2186 585
R3949 gnd.n5250 gnd.n2193 585
R3950 gnd.n5273 gnd.n2193 585
R3951 gnd.n5252 gnd.n5251 585
R3952 gnd.n5251 gnd.n2192 585
R3953 gnd.n5253 gnd.n2202 585
R3954 gnd.n5263 gnd.n2202 585
R3955 gnd.n5255 gnd.n5254 585
R3956 gnd.n5256 gnd.n5255 585
R3957 gnd.n5249 gnd.n2209 585
R3958 gnd.n5257 gnd.n2209 585
R3959 gnd.n5248 gnd.n5247 585
R3960 gnd.n5247 gnd.n5246 585
R3961 gnd.n2211 gnd.n2210 585
R3962 gnd.n2212 gnd.n2211 585
R3963 gnd.n5187 gnd.n5186 585
R3964 gnd.n5188 gnd.n5187 585
R3965 gnd.n5185 gnd.n5109 585
R3966 gnd.n5109 gnd.n1378 585
R3967 gnd.n5184 gnd.n5183 585
R3968 gnd.n5183 gnd.n1376 585
R3969 gnd.n5182 gnd.n5101 585
R3970 gnd.n5195 gnd.n5101 585
R3971 gnd.n5181 gnd.n5180 585
R3972 gnd.n5180 gnd.n1366 585
R3973 gnd.n5179 gnd.n1364 585
R3974 gnd.n6473 gnd.n1364 585
R3975 gnd.n5178 gnd.n1363 585
R3976 gnd.n6474 gnd.n1363 585
R3977 gnd.n5177 gnd.n5176 585
R3978 gnd.n5176 gnd.n5175 585
R3979 gnd.n6710 gnd.n6709 585
R3980 gnd.n6709 gnd.n6708 585
R3981 gnd.n7611 gnd.n7610 585
R3982 gnd.n7610 gnd.n259 585
R3983 gnd.n7614 gnd.n409 585
R3984 gnd.n409 gnd.n266 585
R3985 gnd.n7616 gnd.n7615 585
R3986 gnd.n7616 gnd.n277 585
R3987 gnd.n7617 gnd.n408 585
R3988 gnd.n7617 gnd.n275 585
R3989 gnd.n7619 gnd.n7618 585
R3990 gnd.n7618 gnd.n285 585
R3991 gnd.n7620 gnd.n403 585
R3992 gnd.n403 gnd.n283 585
R3993 gnd.n7622 gnd.n7621 585
R3994 gnd.n7623 gnd.n7622 585
R3995 gnd.n404 gnd.n402 585
R3996 gnd.n402 gnd.n291 585
R3997 gnd.n6271 gnd.n6270 585
R3998 gnd.n6271 gnd.n300 585
R3999 gnd.n6273 gnd.n6272 585
R4000 gnd.n6272 gnd.n298 585
R4001 gnd.n6274 gnd.n6264 585
R4002 gnd.n6264 gnd.n308 585
R4003 gnd.n6276 gnd.n6275 585
R4004 gnd.n6276 gnd.n306 585
R4005 gnd.n6277 gnd.n6263 585
R4006 gnd.n6277 gnd.n337 585
R4007 gnd.n6279 gnd.n6278 585
R4008 gnd.n6278 gnd.n335 585
R4009 gnd.n6281 gnd.n1539 585
R4010 gnd.n1539 gnd.n339 585
R4011 gnd.n6283 gnd.n6282 585
R4012 gnd.n6284 gnd.n6283 585
R4013 gnd.n6261 gnd.n1538 585
R4014 gnd.n1538 gnd.n1533 585
R4015 gnd.n6260 gnd.n6259 585
R4016 gnd.n6259 gnd.n1531 585
R4017 gnd.n6258 gnd.n6257 585
R4018 gnd.n6258 gnd.n323 585
R4019 gnd.n6256 gnd.n1541 585
R4020 gnd.n1541 gnd.n320 585
R4021 gnd.n6254 gnd.n6253 585
R4022 gnd.n6253 gnd.n1518 585
R4023 gnd.n6252 gnd.n1542 585
R4024 gnd.n6252 gnd.n1515 585
R4025 gnd.n6251 gnd.n6250 585
R4026 gnd.n6251 gnd.n1521 585
R4027 gnd.n1544 gnd.n1543 585
R4028 gnd.n1552 gnd.n1543 585
R4029 gnd.n6245 gnd.n6244 585
R4030 gnd.n6244 gnd.n6243 585
R4031 gnd.n1547 gnd.n1546 585
R4032 gnd.n6231 gnd.n1547 585
R4033 gnd.n1587 gnd.n1586 585
R4034 gnd.n1587 gnd.n1558 585
R4035 gnd.n6207 gnd.n6206 585
R4036 gnd.n6206 gnd.n6205 585
R4037 gnd.n6208 gnd.n1580 585
R4038 gnd.n1580 gnd.n1567 585
R4039 gnd.n6210 gnd.n6209 585
R4040 gnd.n6211 gnd.n6210 585
R4041 gnd.n1581 gnd.n1579 585
R4042 gnd.n1579 gnd.n1574 585
R4043 gnd.n6137 gnd.n6136 585
R4044 gnd.n6137 gnd.n1593 585
R4045 gnd.n6139 gnd.n6138 585
R4046 gnd.n6138 gnd.n1602 585
R4047 gnd.n6140 gnd.n1616 585
R4048 gnd.n1616 gnd.n1600 585
R4049 gnd.n6142 gnd.n6141 585
R4050 gnd.n6143 gnd.n6142 585
R4051 gnd.n1617 gnd.n1615 585
R4052 gnd.n1615 gnd.n1611 585
R4053 gnd.n6128 gnd.n6127 585
R4054 gnd.n6127 gnd.n6126 585
R4055 gnd.n1620 gnd.n1619 585
R4056 gnd.n1632 gnd.n1620 585
R4057 gnd.n6102 gnd.n1644 585
R4058 gnd.n1644 gnd.n1630 585
R4059 gnd.n6104 gnd.n6103 585
R4060 gnd.n6105 gnd.n6104 585
R4061 gnd.n1645 gnd.n1643 585
R4062 gnd.n1643 gnd.n1639 585
R4063 gnd.n6097 gnd.n6096 585
R4064 gnd.n6096 gnd.n6095 585
R4065 gnd.n1648 gnd.n1647 585
R4066 gnd.n1658 gnd.n1648 585
R4067 gnd.n6069 gnd.n1670 585
R4068 gnd.n1670 gnd.n1656 585
R4069 gnd.n6071 gnd.n6070 585
R4070 gnd.n6072 gnd.n6071 585
R4071 gnd.n1671 gnd.n1669 585
R4072 gnd.n1669 gnd.n1665 585
R4073 gnd.n6064 gnd.n6063 585
R4074 gnd.n6063 gnd.n6062 585
R4075 gnd.n1674 gnd.n1673 585
R4076 gnd.n1684 gnd.n1674 585
R4077 gnd.n6037 gnd.n1720 585
R4078 gnd.n1720 gnd.n1682 585
R4079 gnd.n6039 gnd.n6038 585
R4080 gnd.n6040 gnd.n6039 585
R4081 gnd.n1721 gnd.n1719 585
R4082 gnd.n1719 gnd.n1690 585
R4083 gnd.n6032 gnd.n6031 585
R4084 gnd.n6031 gnd.n6030 585
R4085 gnd.n5871 gnd.n1723 585
R4086 gnd.n6029 gnd.n5871 585
R4087 gnd.n5870 gnd.n5869 585
R4088 gnd.n5870 gnd.n1474 585
R4089 gnd.n1724 gnd.n1473 585
R4090 gnd.n6355 gnd.n1473 585
R4091 gnd.n5865 gnd.n5864 585
R4092 gnd.n5864 gnd.n1472 585
R4093 gnd.n5863 gnd.n1726 585
R4094 gnd.n5863 gnd.n5862 585
R4095 gnd.n5850 gnd.n1727 585
R4096 gnd.n1728 gnd.n1727 585
R4097 gnd.n5852 gnd.n5851 585
R4098 gnd.n5853 gnd.n5852 585
R4099 gnd.n1736 gnd.n1735 585
R4100 gnd.n1735 gnd.n1734 585
R4101 gnd.n5845 gnd.n5844 585
R4102 gnd.n5844 gnd.n5843 585
R4103 gnd.n1739 gnd.n1738 585
R4104 gnd.n1746 gnd.n1739 585
R4105 gnd.n5833 gnd.n5832 585
R4106 gnd.n5834 gnd.n5833 585
R4107 gnd.n1748 gnd.n1747 585
R4108 gnd.n1747 gnd.n1745 585
R4109 gnd.n5828 gnd.n5827 585
R4110 gnd.n5827 gnd.n5826 585
R4111 gnd.n1751 gnd.n1750 585
R4112 gnd.n1752 gnd.n1751 585
R4113 gnd.n5816 gnd.n5815 585
R4114 gnd.n5817 gnd.n5816 585
R4115 gnd.n1760 gnd.n1759 585
R4116 gnd.n1759 gnd.n1758 585
R4117 gnd.n5811 gnd.n5810 585
R4118 gnd.n5810 gnd.n5809 585
R4119 gnd.n1763 gnd.n1762 585
R4120 gnd.n1764 gnd.n1763 585
R4121 gnd.n5799 gnd.n5798 585
R4122 gnd.n5800 gnd.n5799 585
R4123 gnd.n1772 gnd.n1771 585
R4124 gnd.n1771 gnd.n1770 585
R4125 gnd.n5794 gnd.n5793 585
R4126 gnd.n5793 gnd.n5792 585
R4127 gnd.n1775 gnd.n1774 585
R4128 gnd.n1776 gnd.n1775 585
R4129 gnd.n5782 gnd.n5781 585
R4130 gnd.n5783 gnd.n5782 585
R4131 gnd.n1783 gnd.n1782 585
R4132 gnd.n5773 gnd.n1782 585
R4133 gnd.n5777 gnd.n5776 585
R4134 gnd.n5776 gnd.n5775 585
R4135 gnd.n1786 gnd.n1785 585
R4136 gnd.n1787 gnd.n1786 585
R4137 gnd.n5764 gnd.n5763 585
R4138 gnd.n5765 gnd.n5764 585
R4139 gnd.n1795 gnd.n1794 585
R4140 gnd.n1794 gnd.n1793 585
R4141 gnd.n5759 gnd.n5758 585
R4142 gnd.n5758 gnd.n5757 585
R4143 gnd.n1798 gnd.n1797 585
R4144 gnd.n1992 gnd.n1798 585
R4145 gnd.n5589 gnd.n5588 585
R4146 gnd.n5590 gnd.n5589 585
R4147 gnd.n2001 gnd.n2000 585
R4148 gnd.n2000 gnd.n1997 585
R4149 gnd.n5584 gnd.n5583 585
R4150 gnd.n5583 gnd.n5582 585
R4151 gnd.n2004 gnd.n2003 585
R4152 gnd.n5573 gnd.n2004 585
R4153 gnd.n5558 gnd.n5557 585
R4154 gnd.n5559 gnd.n5558 585
R4155 gnd.n2017 gnd.n2016 585
R4156 gnd.n5474 gnd.n2016 585
R4157 gnd.n5553 gnd.n5552 585
R4158 gnd.n5552 gnd.n5551 585
R4159 gnd.n2020 gnd.n2019 585
R4160 gnd.n5539 gnd.n2020 585
R4161 gnd.n5500 gnd.n2060 585
R4162 gnd.n5500 gnd.n5499 585
R4163 gnd.n5501 gnd.n2057 585
R4164 gnd.n5501 gnd.n2033 585
R4165 gnd.n5503 gnd.n5502 585
R4166 gnd.n5502 gnd.n2038 585
R4167 gnd.n5504 gnd.n2052 585
R4168 gnd.n2052 gnd.n2044 585
R4169 gnd.n5506 gnd.n5505 585
R4170 gnd.n5507 gnd.n5506 585
R4171 gnd.n2053 gnd.n2051 585
R4172 gnd.n2051 gnd.n2048 585
R4173 gnd.n5459 gnd.n5458 585
R4174 gnd.n5460 gnd.n5459 585
R4175 gnd.n2075 gnd.n2074 585
R4176 gnd.n2082 gnd.n2074 585
R4177 gnd.n5453 gnd.n5452 585
R4178 gnd.n5452 gnd.n5451 585
R4179 gnd.n2078 gnd.n2077 585
R4180 gnd.n2087 gnd.n2078 585
R4181 gnd.n5417 gnd.n2103 585
R4182 gnd.n2103 gnd.n2094 585
R4183 gnd.n5419 gnd.n5418 585
R4184 gnd.n5420 gnd.n5419 585
R4185 gnd.n2104 gnd.n2102 585
R4186 gnd.n2102 gnd.n2098 585
R4187 gnd.n5412 gnd.n5411 585
R4188 gnd.n5411 gnd.n5410 585
R4189 gnd.n2107 gnd.n2106 585
R4190 gnd.n5402 gnd.n2107 585
R4191 gnd.n5376 gnd.n2126 585
R4192 gnd.n2126 gnd.n2125 585
R4193 gnd.n5378 gnd.n5377 585
R4194 gnd.n5379 gnd.n5378 585
R4195 gnd.n2127 gnd.n2124 585
R4196 gnd.n2134 gnd.n2124 585
R4197 gnd.n5371 gnd.n5370 585
R4198 gnd.n5370 gnd.n5369 585
R4199 gnd.n2130 gnd.n2129 585
R4200 gnd.n2139 gnd.n2130 585
R4201 gnd.n5321 gnd.n2155 585
R4202 gnd.n2155 gnd.n2145 585
R4203 gnd.n5323 gnd.n5322 585
R4204 gnd.n5324 gnd.n5323 585
R4205 gnd.n2156 gnd.n2154 585
R4206 gnd.n2154 gnd.n2150 585
R4207 gnd.n5316 gnd.n5315 585
R4208 gnd.n5315 gnd.n5314 585
R4209 gnd.n2159 gnd.n2158 585
R4210 gnd.n2168 gnd.n2159 585
R4211 gnd.n5295 gnd.n5294 585
R4212 gnd.n5296 gnd.n5295 585
R4213 gnd.n2178 gnd.n2177 585
R4214 gnd.n2177 gnd.n2174 585
R4215 gnd.n5290 gnd.n5289 585
R4216 gnd.n5289 gnd.n5288 585
R4217 gnd.n2181 gnd.n2180 585
R4218 gnd.n2187 gnd.n2181 585
R4219 gnd.n5271 gnd.n5270 585
R4220 gnd.n5272 gnd.n5271 585
R4221 gnd.n2197 gnd.n2196 585
R4222 gnd.n2204 gnd.n2196 585
R4223 gnd.n5266 gnd.n5265 585
R4224 gnd.n5265 gnd.n5264 585
R4225 gnd.n2200 gnd.n2199 585
R4226 gnd.n2208 gnd.n2200 585
R4227 gnd.n5244 gnd.n5243 585
R4228 gnd.n5245 gnd.n5244 585
R4229 gnd.n1375 gnd.n1374 585
R4230 gnd.n5108 gnd.n1375 585
R4231 gnd.n6468 gnd.n6467 585
R4232 gnd.n6467 gnd.n6466 585
R4233 gnd.n6469 gnd.n1369 585
R4234 gnd.n5196 gnd.n1369 585
R4235 gnd.n6471 gnd.n6470 585
R4236 gnd.n6472 gnd.n6471 585
R4237 gnd.n1370 gnd.n1368 585
R4238 gnd.n1368 gnd.n1362 585
R4239 gnd.n5089 gnd.n2225 585
R4240 gnd.n2225 gnd.n1336 585
R4241 gnd.n5091 gnd.n5090 585
R4242 gnd.n5092 gnd.n5091 585
R4243 gnd.n2226 gnd.n2224 585
R4244 gnd.n2224 gnd.n2222 585
R4245 gnd.n5083 gnd.n5082 585
R4246 gnd.n5082 gnd.n5081 585
R4247 gnd.n2229 gnd.n2228 585
R4248 gnd.n2230 gnd.n2229 585
R4249 gnd.n5061 gnd.n5060 585
R4250 gnd.n5062 gnd.n5061 585
R4251 gnd.n2241 gnd.n2240 585
R4252 gnd.n2247 gnd.n2240 585
R4253 gnd.n5056 gnd.n5055 585
R4254 gnd.n5055 gnd.n5054 585
R4255 gnd.n2244 gnd.n2243 585
R4256 gnd.n2245 gnd.n2244 585
R4257 gnd.n5045 gnd.n5044 585
R4258 gnd.n5046 gnd.n5045 585
R4259 gnd.n2256 gnd.n2255 585
R4260 gnd.n2255 gnd.n2253 585
R4261 gnd.n5040 gnd.n5039 585
R4262 gnd.n5039 gnd.n5038 585
R4263 gnd.n2259 gnd.n2258 585
R4264 gnd.n2260 gnd.n2259 585
R4265 gnd.n5029 gnd.n5028 585
R4266 gnd.n5030 gnd.n5029 585
R4267 gnd.n2270 gnd.n2269 585
R4268 gnd.n2269 gnd.n2267 585
R4269 gnd.n5024 gnd.n5023 585
R4270 gnd.n5023 gnd.n5022 585
R4271 gnd.n2273 gnd.n2272 585
R4272 gnd.n2274 gnd.n2273 585
R4273 gnd.n5013 gnd.n5012 585
R4274 gnd.n5014 gnd.n5013 585
R4275 gnd.n2284 gnd.n2283 585
R4276 gnd.n2283 gnd.n2281 585
R4277 gnd.n5008 gnd.n5007 585
R4278 gnd.n5007 gnd.n5006 585
R4279 gnd.n2287 gnd.n2286 585
R4280 gnd.n2296 gnd.n2287 585
R4281 gnd.n4997 gnd.n4996 585
R4282 gnd.n4998 gnd.n4997 585
R4283 gnd.n2298 gnd.n2297 585
R4284 gnd.n2297 gnd.n2294 585
R4285 gnd.n4992 gnd.n4991 585
R4286 gnd.n4991 gnd.n4990 585
R4287 gnd.n2301 gnd.n2300 585
R4288 gnd.n2302 gnd.n2301 585
R4289 gnd.n4981 gnd.n4980 585
R4290 gnd.n4982 gnd.n4981 585
R4291 gnd.n2312 gnd.n2311 585
R4292 gnd.n2311 gnd.n2309 585
R4293 gnd.n4976 gnd.n4975 585
R4294 gnd.n4975 gnd.n4974 585
R4295 gnd.n2315 gnd.n2314 585
R4296 gnd.n2316 gnd.n2315 585
R4297 gnd.n4916 gnd.n4914 585
R4298 gnd.n4916 gnd.n4915 585
R4299 gnd.n4918 gnd.n4917 585
R4300 gnd.n4917 gnd.n1262 585
R4301 gnd.n4919 gnd.n2462 585
R4302 gnd.n2462 gnd.n1251 585
R4303 gnd.n4921 gnd.n4920 585
R4304 gnd.n4922 gnd.n4921 585
R4305 gnd.n2463 gnd.n2461 585
R4306 gnd.n2461 gnd.n1244 585
R4307 gnd.n4907 gnd.n4906 585
R4308 gnd.n4906 gnd.n1241 585
R4309 gnd.n4905 gnd.n2465 585
R4310 gnd.n4905 gnd.n1233 585
R4311 gnd.n4904 gnd.n4903 585
R4312 gnd.n4904 gnd.n1230 585
R4313 gnd.n2467 gnd.n2466 585
R4314 gnd.n2466 gnd.n1222 585
R4315 gnd.n4899 gnd.n4898 585
R4316 gnd.n4898 gnd.n1219 585
R4317 gnd.n4897 gnd.n2469 585
R4318 gnd.n4897 gnd.n1211 585
R4319 gnd.n4896 gnd.n4895 585
R4320 gnd.n4896 gnd.n1208 585
R4321 gnd.n2471 gnd.n2470 585
R4322 gnd.n2470 gnd.n1200 585
R4323 gnd.n4891 gnd.n4890 585
R4324 gnd.n4890 gnd.n4889 585
R4325 gnd.n2474 gnd.n2473 585
R4326 gnd.n2474 gnd.n1190 585
R4327 gnd.n4702 gnd.n4701 585
R4328 gnd.n4701 gnd.n1187 585
R4329 gnd.n4703 gnd.n4696 585
R4330 gnd.n4696 gnd.n1179 585
R4331 gnd.n4705 gnd.n4704 585
R4332 gnd.n4705 gnd.n1176 585
R4333 gnd.n4706 gnd.n4695 585
R4334 gnd.n4706 gnd.n1168 585
R4335 gnd.n4708 gnd.n4707 585
R4336 gnd.n4707 gnd.n1165 585
R4337 gnd.n4709 gnd.n2503 585
R4338 gnd.n2503 gnd.n1157 585
R4339 gnd.n4711 gnd.n4710 585
R4340 gnd.n4712 gnd.n4711 585
R4341 gnd.n2504 gnd.n2502 585
R4342 gnd.n2502 gnd.n1147 585
R4343 gnd.n4689 gnd.n4688 585
R4344 gnd.n4688 gnd.n1144 585
R4345 gnd.n4687 gnd.n2506 585
R4346 gnd.n4687 gnd.n1136 585
R4347 gnd.n4686 gnd.n4685 585
R4348 gnd.n4686 gnd.n1133 585
R4349 gnd.n2508 gnd.n2507 585
R4350 gnd.n2507 gnd.n1125 585
R4351 gnd.n4681 gnd.n4680 585
R4352 gnd.n4680 gnd.n1122 585
R4353 gnd.n4679 gnd.n2510 585
R4354 gnd.n4679 gnd.n1115 585
R4355 gnd.n4678 gnd.n2512 585
R4356 gnd.n4678 gnd.n4677 585
R4357 gnd.n4606 gnd.n2511 585
R4358 gnd.n2511 gnd.n1104 585
R4359 gnd.n4608 gnd.n4607 585
R4360 gnd.n4608 gnd.n1101 585
R4361 gnd.n4610 gnd.n4609 585
R4362 gnd.n4609 gnd.n2537 585
R4363 gnd.n4611 gnd.n2545 585
R4364 gnd.n2545 gnd.n2534 585
R4365 gnd.n4614 gnd.n4613 585
R4366 gnd.n4615 gnd.n4614 585
R4367 gnd.n4602 gnd.n2544 585
R4368 gnd.n2544 gnd.n2542 585
R4369 gnd.n4600 gnd.n4599 585
R4370 gnd.n4599 gnd.n4598 585
R4371 gnd.n2547 gnd.n2546 585
R4372 gnd.n4582 gnd.n2547 585
R4373 gnd.n4559 gnd.n2575 585
R4374 gnd.n2575 gnd.n2551 585
R4375 gnd.n4561 gnd.n4560 585
R4376 gnd.n4562 gnd.n4561 585
R4377 gnd.n4556 gnd.n2574 585
R4378 gnd.n2574 gnd.n1086 585
R4379 gnd.n4555 gnd.n4554 585
R4380 gnd.n4554 gnd.n1078 585
R4381 gnd.n4553 gnd.n2576 585
R4382 gnd.n4553 gnd.n4552 585
R4383 gnd.n2601 gnd.n2578 585
R4384 gnd.n2578 gnd.n1068 585
R4385 gnd.n2603 gnd.n2602 585
R4386 gnd.n2603 gnd.n1065 585
R4387 gnd.n2605 gnd.n2604 585
R4388 gnd.n2604 gnd.n1057 585
R4389 gnd.n2606 gnd.n2587 585
R4390 gnd.n2587 gnd.n1054 585
R4391 gnd.n2608 gnd.n2607 585
R4392 gnd.n2609 gnd.n2608 585
R4393 gnd.n2588 gnd.n2586 585
R4394 gnd.n2586 gnd.n1044 585
R4395 gnd.n2592 gnd.n2591 585
R4396 gnd.n2591 gnd.n1035 585
R4397 gnd.n2590 gnd.n1018 585
R4398 gnd.n1032 gnd.n1018 585
R4399 gnd.n6354 gnd.n6353 585
R4400 gnd.n6355 gnd.n6354 585
R4401 gnd.n1477 gnd.n1475 585
R4402 gnd.n1475 gnd.n1472 585
R4403 gnd.n5860 gnd.n5859 585
R4404 gnd.n5862 gnd.n5860 585
R4405 gnd.n1730 gnd.n1729 585
R4406 gnd.n1729 gnd.n1728 585
R4407 gnd.n5855 gnd.n5854 585
R4408 gnd.n5854 gnd.n5853 585
R4409 gnd.n1733 gnd.n1732 585
R4410 gnd.n1734 gnd.n1733 585
R4411 gnd.n5841 gnd.n5840 585
R4412 gnd.n5843 gnd.n5841 585
R4413 gnd.n1741 gnd.n1740 585
R4414 gnd.n1746 gnd.n1740 585
R4415 gnd.n5836 gnd.n5835 585
R4416 gnd.n5835 gnd.n5834 585
R4417 gnd.n1744 gnd.n1743 585
R4418 gnd.n1745 gnd.n1744 585
R4419 gnd.n5824 gnd.n5823 585
R4420 gnd.n5826 gnd.n5824 585
R4421 gnd.n1754 gnd.n1753 585
R4422 gnd.n1753 gnd.n1752 585
R4423 gnd.n5819 gnd.n5818 585
R4424 gnd.n5818 gnd.n5817 585
R4425 gnd.n1757 gnd.n1756 585
R4426 gnd.n1758 gnd.n1757 585
R4427 gnd.n5807 gnd.n5806 585
R4428 gnd.n5809 gnd.n5807 585
R4429 gnd.n1766 gnd.n1765 585
R4430 gnd.n1765 gnd.n1764 585
R4431 gnd.n5802 gnd.n5801 585
R4432 gnd.n5801 gnd.n5800 585
R4433 gnd.n1769 gnd.n1768 585
R4434 gnd.n1770 gnd.n1769 585
R4435 gnd.n5790 gnd.n5789 585
R4436 gnd.n5792 gnd.n5790 585
R4437 gnd.n1778 gnd.n1777 585
R4438 gnd.n1777 gnd.n1776 585
R4439 gnd.n5785 gnd.n5784 585
R4440 gnd.n5784 gnd.n5783 585
R4441 gnd.n1781 gnd.n1780 585
R4442 gnd.n5773 gnd.n1781 585
R4443 gnd.n5772 gnd.n5771 585
R4444 gnd.n5775 gnd.n5772 585
R4445 gnd.n1789 gnd.n1788 585
R4446 gnd.n1788 gnd.n1787 585
R4447 gnd.n5767 gnd.n5766 585
R4448 gnd.n5766 gnd.n5765 585
R4449 gnd.n1792 gnd.n1791 585
R4450 gnd.n1793 gnd.n1792 585
R4451 gnd.n5481 gnd.n1800 585
R4452 gnd.n5757 gnd.n1800 585
R4453 gnd.n5480 gnd.n5479 585
R4454 gnd.n5479 gnd.n1992 585
R4455 gnd.n5485 gnd.n1999 585
R4456 gnd.n5590 gnd.n1999 585
R4457 gnd.n5486 gnd.n5478 585
R4458 gnd.n5478 gnd.n1997 585
R4459 gnd.n5487 gnd.n2005 585
R4460 gnd.n5582 gnd.n2005 585
R4461 gnd.n5476 gnd.n2011 585
R4462 gnd.n5573 gnd.n2011 585
R4463 gnd.n5491 gnd.n2015 585
R4464 gnd.n5559 gnd.n2015 585
R4465 gnd.n5492 gnd.n5475 585
R4466 gnd.n5475 gnd.n5474 585
R4467 gnd.n5493 gnd.n2021 585
R4468 gnd.n5551 gnd.n2021 585
R4469 gnd.n2063 gnd.n2030 585
R4470 gnd.n5539 gnd.n2030 585
R4471 gnd.n5498 gnd.n5497 585
R4472 gnd.n5499 gnd.n5498 585
R4473 gnd.n2062 gnd.n2061 585
R4474 gnd.n2061 gnd.n2033 585
R4475 gnd.n5470 gnd.n5469 585
R4476 gnd.n5469 gnd.n2038 585
R4477 gnd.n5468 gnd.n5467 585
R4478 gnd.n5468 gnd.n2044 585
R4479 gnd.n5466 gnd.n2050 585
R4480 gnd.n5507 gnd.n2050 585
R4481 gnd.n2069 gnd.n2065 585
R4482 gnd.n2069 gnd.n2048 585
R4483 gnd.n5462 gnd.n5461 585
R4484 gnd.n5461 gnd.n5460 585
R4485 gnd.n2068 gnd.n2067 585
R4486 gnd.n2082 gnd.n2068 585
R4487 gnd.n5389 gnd.n2080 585
R4488 gnd.n5451 gnd.n2080 585
R4489 gnd.n5388 gnd.n5387 585
R4490 gnd.n5387 gnd.n2087 585
R4491 gnd.n5393 gnd.n5386 585
R4492 gnd.n5386 gnd.n2094 585
R4493 gnd.n5394 gnd.n2100 585
R4494 gnd.n5420 gnd.n2100 585
R4495 gnd.n5395 gnd.n5385 585
R4496 gnd.n5385 gnd.n2098 585
R4497 gnd.n2118 gnd.n2109 585
R4498 gnd.n5410 gnd.n2109 585
R4499 gnd.n5400 gnd.n5399 585
R4500 gnd.n5402 gnd.n5400 585
R4501 gnd.n2117 gnd.n2116 585
R4502 gnd.n2125 gnd.n2116 585
R4503 gnd.n5381 gnd.n5380 585
R4504 gnd.n5380 gnd.n5379 585
R4505 gnd.n2121 gnd.n2120 585
R4506 gnd.n2134 gnd.n2121 585
R4507 gnd.n5216 gnd.n2132 585
R4508 gnd.n5369 gnd.n2132 585
R4509 gnd.n5217 gnd.n5215 585
R4510 gnd.n5215 gnd.n2139 585
R4511 gnd.n5214 gnd.n5212 585
R4512 gnd.n5214 gnd.n2145 585
R4513 gnd.n5221 gnd.n2152 585
R4514 gnd.n5324 gnd.n2152 585
R4515 gnd.n5222 gnd.n5211 585
R4516 gnd.n5211 gnd.n2150 585
R4517 gnd.n5223 gnd.n2162 585
R4518 gnd.n5314 gnd.n2162 585
R4519 gnd.n5209 gnd.n5208 585
R4520 gnd.n5208 gnd.n2168 585
R4521 gnd.n5227 gnd.n2176 585
R4522 gnd.n5296 gnd.n2176 585
R4523 gnd.n5228 gnd.n5207 585
R4524 gnd.n5207 gnd.n2174 585
R4525 gnd.n5229 gnd.n2183 585
R4526 gnd.n5288 gnd.n2183 585
R4527 gnd.n5205 gnd.n5204 585
R4528 gnd.n5204 gnd.n2187 585
R4529 gnd.n5233 gnd.n2194 585
R4530 gnd.n5272 gnd.n2194 585
R4531 gnd.n5234 gnd.n5203 585
R4532 gnd.n5203 gnd.n2204 585
R4533 gnd.n5235 gnd.n2201 585
R4534 gnd.n5264 gnd.n2201 585
R4535 gnd.n2216 gnd.n2214 585
R4536 gnd.n2214 gnd.n2208 585
R4537 gnd.n5240 gnd.n5239 585
R4538 gnd.n5245 gnd.n5240 585
R4539 gnd.n2215 gnd.n2213 585
R4540 gnd.n5108 gnd.n2213 585
R4541 gnd.n5199 gnd.n1377 585
R4542 gnd.n6466 gnd.n1377 585
R4543 gnd.n5198 gnd.n5197 585
R4544 gnd.n5197 gnd.n5196 585
R4545 gnd.n5100 gnd.n1365 585
R4546 gnd.n6472 gnd.n1365 585
R4547 gnd.n5094 gnd.n2218 585
R4548 gnd.n5094 gnd.n1362 585
R4549 gnd.n5096 gnd.n5095 585
R4550 gnd.n5095 gnd.n1336 585
R4551 gnd.n5093 gnd.n2220 585
R4552 gnd.n5093 gnd.n5092 585
R4553 gnd.n2364 gnd.n2221 585
R4554 gnd.n2222 gnd.n2221 585
R4555 gnd.n2363 gnd.n2231 585
R4556 gnd.n5081 gnd.n2231 585
R4557 gnd.n2368 gnd.n2362 585
R4558 gnd.n2362 gnd.n2230 585
R4559 gnd.n2369 gnd.n2239 585
R4560 gnd.n5062 gnd.n2239 585
R4561 gnd.n2370 gnd.n2361 585
R4562 gnd.n2361 gnd.n2247 585
R4563 gnd.n2359 gnd.n2246 585
R4564 gnd.n5054 gnd.n2246 585
R4565 gnd.n2374 gnd.n2358 585
R4566 gnd.n2358 gnd.n2245 585
R4567 gnd.n2375 gnd.n2254 585
R4568 gnd.n5046 gnd.n2254 585
R4569 gnd.n2376 gnd.n2357 585
R4570 gnd.n2357 gnd.n2253 585
R4571 gnd.n2355 gnd.n2261 585
R4572 gnd.n5038 gnd.n2261 585
R4573 gnd.n2380 gnd.n2354 585
R4574 gnd.n2354 gnd.n2260 585
R4575 gnd.n2381 gnd.n2268 585
R4576 gnd.n5030 gnd.n2268 585
R4577 gnd.n2382 gnd.n2353 585
R4578 gnd.n2353 gnd.n2267 585
R4579 gnd.n2351 gnd.n2275 585
R4580 gnd.n5022 gnd.n2275 585
R4581 gnd.n2386 gnd.n2350 585
R4582 gnd.n2350 gnd.n2274 585
R4583 gnd.n2387 gnd.n2282 585
R4584 gnd.n5014 gnd.n2282 585
R4585 gnd.n2388 gnd.n2349 585
R4586 gnd.n2349 gnd.n2281 585
R4587 gnd.n2347 gnd.n2288 585
R4588 gnd.n5006 gnd.n2288 585
R4589 gnd.n2392 gnd.n2346 585
R4590 gnd.n2346 gnd.n2296 585
R4591 gnd.n2393 gnd.n2295 585
R4592 gnd.n4998 gnd.n2295 585
R4593 gnd.n2394 gnd.n2345 585
R4594 gnd.n2345 gnd.n2294 585
R4595 gnd.n2343 gnd.n2303 585
R4596 gnd.n4990 gnd.n2303 585
R4597 gnd.n2398 gnd.n2342 585
R4598 gnd.n2342 gnd.n2302 585
R4599 gnd.n2399 gnd.n2310 585
R4600 gnd.n4982 gnd.n2310 585
R4601 gnd.n2400 gnd.n2332 585
R4602 gnd.n2332 gnd.n2309 585
R4603 gnd.n4971 gnd.n4970 585
R4604 gnd.n4969 gnd.n2331 585
R4605 gnd.n2334 gnd.n2330 585
R4606 gnd.n4973 gnd.n2330 585
R4607 gnd.n4962 gnd.n2412 585
R4608 gnd.n4961 gnd.n2413 585
R4609 gnd.n2415 gnd.n2414 585
R4610 gnd.n4954 gnd.n2421 585
R4611 gnd.n4953 gnd.n2422 585
R4612 gnd.n2431 gnd.n2423 585
R4613 gnd.n4946 gnd.n2432 585
R4614 gnd.n4945 gnd.n2433 585
R4615 gnd.n2435 gnd.n2434 585
R4616 gnd.n4938 gnd.n2441 585
R4617 gnd.n4937 gnd.n2442 585
R4618 gnd.n2453 gnd.n2443 585
R4619 gnd.n4930 gnd.n2454 585
R4620 gnd.n4929 gnd.n2455 585
R4621 gnd.n2457 gnd.n2456 585
R4622 gnd.n4868 gnd.n4835 585
R4623 gnd.n4867 gnd.n4836 585
R4624 gnd.n4866 gnd.n4837 585
R4625 gnd.n4839 gnd.n4838 585
R4626 gnd.n4862 gnd.n4841 585
R4627 gnd.n4861 gnd.n4842 585
R4628 gnd.n4860 gnd.n4843 585
R4629 gnd.n4857 gnd.n4848 585
R4630 gnd.n4856 gnd.n4849 585
R4631 gnd.n4855 gnd.n4850 585
R4632 gnd.n4852 gnd.n4851 585
R4633 gnd.n6357 gnd.n6356 585
R4634 gnd.n6356 gnd.n6355 585
R4635 gnd.n6358 gnd.n1470 585
R4636 gnd.n1472 gnd.n1470 585
R4637 gnd.n5861 gnd.n1468 585
R4638 gnd.n5862 gnd.n5861 585
R4639 gnd.n6362 gnd.n1467 585
R4640 gnd.n1728 gnd.n1467 585
R4641 gnd.n6363 gnd.n1466 585
R4642 gnd.n5853 gnd.n1466 585
R4643 gnd.n6364 gnd.n1465 585
R4644 gnd.n1734 gnd.n1465 585
R4645 gnd.n5842 gnd.n1463 585
R4646 gnd.n5843 gnd.n5842 585
R4647 gnd.n6368 gnd.n1462 585
R4648 gnd.n1746 gnd.n1462 585
R4649 gnd.n6369 gnd.n1461 585
R4650 gnd.n5834 gnd.n1461 585
R4651 gnd.n6370 gnd.n1460 585
R4652 gnd.n1745 gnd.n1460 585
R4653 gnd.n5825 gnd.n1458 585
R4654 gnd.n5826 gnd.n5825 585
R4655 gnd.n6374 gnd.n1457 585
R4656 gnd.n1752 gnd.n1457 585
R4657 gnd.n6375 gnd.n1456 585
R4658 gnd.n5817 gnd.n1456 585
R4659 gnd.n6376 gnd.n1455 585
R4660 gnd.n1758 gnd.n1455 585
R4661 gnd.n5808 gnd.n1453 585
R4662 gnd.n5809 gnd.n5808 585
R4663 gnd.n6380 gnd.n1452 585
R4664 gnd.n1764 gnd.n1452 585
R4665 gnd.n6381 gnd.n1451 585
R4666 gnd.n5800 gnd.n1451 585
R4667 gnd.n6382 gnd.n1450 585
R4668 gnd.n1770 gnd.n1450 585
R4669 gnd.n5791 gnd.n1448 585
R4670 gnd.n5792 gnd.n5791 585
R4671 gnd.n6386 gnd.n1447 585
R4672 gnd.n1776 gnd.n1447 585
R4673 gnd.n6387 gnd.n1446 585
R4674 gnd.n5783 gnd.n1446 585
R4675 gnd.n6388 gnd.n1445 585
R4676 gnd.n5773 gnd.n1445 585
R4677 gnd.n5774 gnd.n1443 585
R4678 gnd.n5775 gnd.n5774 585
R4679 gnd.n6392 gnd.n1442 585
R4680 gnd.n1787 gnd.n1442 585
R4681 gnd.n6393 gnd.n1441 585
R4682 gnd.n5765 gnd.n1441 585
R4683 gnd.n6394 gnd.n1440 585
R4684 gnd.n1793 gnd.n1440 585
R4685 gnd.n5756 gnd.n1438 585
R4686 gnd.n5757 gnd.n5756 585
R4687 gnd.n6398 gnd.n1437 585
R4688 gnd.n1992 gnd.n1437 585
R4689 gnd.n6399 gnd.n1436 585
R4690 gnd.n5590 gnd.n1436 585
R4691 gnd.n6400 gnd.n1435 585
R4692 gnd.n1997 gnd.n1435 585
R4693 gnd.n5581 gnd.n1433 585
R4694 gnd.n5582 gnd.n5581 585
R4695 gnd.n6404 gnd.n1432 585
R4696 gnd.n5573 gnd.n1432 585
R4697 gnd.n6405 gnd.n1431 585
R4698 gnd.n5559 gnd.n1431 585
R4699 gnd.n6406 gnd.n1430 585
R4700 gnd.n5474 gnd.n1430 585
R4701 gnd.n5550 gnd.n1428 585
R4702 gnd.n5551 gnd.n5550 585
R4703 gnd.n6410 gnd.n1427 585
R4704 gnd.n5539 gnd.n1427 585
R4705 gnd.n6411 gnd.n1426 585
R4706 gnd.n5499 gnd.n1426 585
R4707 gnd.n6412 gnd.n1425 585
R4708 gnd.n2033 gnd.n1425 585
R4709 gnd.n2037 gnd.n1423 585
R4710 gnd.n2038 gnd.n2037 585
R4711 gnd.n6416 gnd.n1422 585
R4712 gnd.n2044 gnd.n1422 585
R4713 gnd.n6417 gnd.n1421 585
R4714 gnd.n5507 gnd.n1421 585
R4715 gnd.n6418 gnd.n1420 585
R4716 gnd.n2048 gnd.n1420 585
R4717 gnd.n2072 gnd.n1418 585
R4718 gnd.n5460 gnd.n2072 585
R4719 gnd.n6422 gnd.n1417 585
R4720 gnd.n2082 gnd.n1417 585
R4721 gnd.n6423 gnd.n1416 585
R4722 gnd.n5451 gnd.n1416 585
R4723 gnd.n6424 gnd.n1415 585
R4724 gnd.n2087 gnd.n1415 585
R4725 gnd.n2093 gnd.n1413 585
R4726 gnd.n2094 gnd.n2093 585
R4727 gnd.n6428 gnd.n1412 585
R4728 gnd.n5420 gnd.n1412 585
R4729 gnd.n6429 gnd.n1411 585
R4730 gnd.n2098 gnd.n1411 585
R4731 gnd.n6430 gnd.n1410 585
R4732 gnd.n5410 gnd.n1410 585
R4733 gnd.n5401 gnd.n1408 585
R4734 gnd.n5402 gnd.n5401 585
R4735 gnd.n6434 gnd.n1407 585
R4736 gnd.n2125 gnd.n1407 585
R4737 gnd.n6435 gnd.n1406 585
R4738 gnd.n5379 gnd.n1406 585
R4739 gnd.n6436 gnd.n1405 585
R4740 gnd.n2134 gnd.n1405 585
R4741 gnd.n5368 gnd.n1403 585
R4742 gnd.n5369 gnd.n5368 585
R4743 gnd.n6440 gnd.n1402 585
R4744 gnd.n2139 gnd.n1402 585
R4745 gnd.n6441 gnd.n1401 585
R4746 gnd.n2145 gnd.n1401 585
R4747 gnd.n6442 gnd.n1400 585
R4748 gnd.n5324 gnd.n1400 585
R4749 gnd.n2149 gnd.n1398 585
R4750 gnd.n2150 gnd.n2149 585
R4751 gnd.n6446 gnd.n1397 585
R4752 gnd.n5314 gnd.n1397 585
R4753 gnd.n6447 gnd.n1396 585
R4754 gnd.n2168 gnd.n1396 585
R4755 gnd.n6448 gnd.n1395 585
R4756 gnd.n5296 gnd.n1395 585
R4757 gnd.n2173 gnd.n1393 585
R4758 gnd.n2174 gnd.n2173 585
R4759 gnd.n6452 gnd.n1392 585
R4760 gnd.n5288 gnd.n1392 585
R4761 gnd.n6453 gnd.n1391 585
R4762 gnd.n2187 gnd.n1391 585
R4763 gnd.n6454 gnd.n1390 585
R4764 gnd.n5272 gnd.n1390 585
R4765 gnd.n2203 gnd.n1388 585
R4766 gnd.n2204 gnd.n2203 585
R4767 gnd.n6458 gnd.n1387 585
R4768 gnd.n5264 gnd.n1387 585
R4769 gnd.n6459 gnd.n1386 585
R4770 gnd.n2208 gnd.n1386 585
R4771 gnd.n6460 gnd.n1385 585
R4772 gnd.n5245 gnd.n1385 585
R4773 gnd.n1382 gnd.n1380 585
R4774 gnd.n5108 gnd.n1380 585
R4775 gnd.n6465 gnd.n6464 585
R4776 gnd.n6466 gnd.n6465 585
R4777 gnd.n1381 gnd.n1379 585
R4778 gnd.n5196 gnd.n1379 585
R4779 gnd.n5070 gnd.n1367 585
R4780 gnd.n6472 gnd.n1367 585
R4781 gnd.n5073 gnd.n5069 585
R4782 gnd.n5069 gnd.n1362 585
R4783 gnd.n5074 gnd.n5068 585
R4784 gnd.n5068 gnd.n1336 585
R4785 gnd.n5075 gnd.n2223 585
R4786 gnd.n5092 gnd.n2223 585
R4787 gnd.n2235 gnd.n2233 585
R4788 gnd.n2233 gnd.n2222 585
R4789 gnd.n5080 gnd.n5079 585
R4790 gnd.n5081 gnd.n5080 585
R4791 gnd.n2234 gnd.n2232 585
R4792 gnd.n2232 gnd.n2230 585
R4793 gnd.n5064 gnd.n5063 585
R4794 gnd.n5063 gnd.n5062 585
R4795 gnd.n2238 gnd.n2237 585
R4796 gnd.n2247 gnd.n2238 585
R4797 gnd.n5053 gnd.n5052 585
R4798 gnd.n5054 gnd.n5053 585
R4799 gnd.n2249 gnd.n2248 585
R4800 gnd.n2248 gnd.n2245 585
R4801 gnd.n5048 gnd.n5047 585
R4802 gnd.n5047 gnd.n5046 585
R4803 gnd.n2252 gnd.n2251 585
R4804 gnd.n2253 gnd.n2252 585
R4805 gnd.n5037 gnd.n5036 585
R4806 gnd.n5038 gnd.n5037 585
R4807 gnd.n2263 gnd.n2262 585
R4808 gnd.n2262 gnd.n2260 585
R4809 gnd.n5032 gnd.n5031 585
R4810 gnd.n5031 gnd.n5030 585
R4811 gnd.n2266 gnd.n2265 585
R4812 gnd.n2267 gnd.n2266 585
R4813 gnd.n5021 gnd.n5020 585
R4814 gnd.n5022 gnd.n5021 585
R4815 gnd.n2277 gnd.n2276 585
R4816 gnd.n2276 gnd.n2274 585
R4817 gnd.n5016 gnd.n5015 585
R4818 gnd.n5015 gnd.n5014 585
R4819 gnd.n2280 gnd.n2279 585
R4820 gnd.n2281 gnd.n2280 585
R4821 gnd.n5005 gnd.n5004 585
R4822 gnd.n5006 gnd.n5005 585
R4823 gnd.n2290 gnd.n2289 585
R4824 gnd.n2296 gnd.n2289 585
R4825 gnd.n5000 gnd.n4999 585
R4826 gnd.n4999 gnd.n4998 585
R4827 gnd.n2293 gnd.n2292 585
R4828 gnd.n2294 gnd.n2293 585
R4829 gnd.n4989 gnd.n4988 585
R4830 gnd.n4990 gnd.n4989 585
R4831 gnd.n2305 gnd.n2304 585
R4832 gnd.n2304 gnd.n2302 585
R4833 gnd.n4984 gnd.n4983 585
R4834 gnd.n4983 gnd.n4982 585
R4835 gnd.n2308 gnd.n2307 585
R4836 gnd.n2309 gnd.n2308 585
R4837 gnd.n5887 gnd.n1471 585
R4838 gnd.n6028 gnd.n1471 585
R4839 gnd.n6026 gnd.n6025 585
R4840 gnd.n5886 gnd.n5885 585
R4841 gnd.n6020 gnd.n6019 585
R4842 gnd.n6017 gnd.n6016 585
R4843 gnd.n6015 gnd.n6014 585
R4844 gnd.n6008 gnd.n5891 585
R4845 gnd.n6010 gnd.n6009 585
R4846 gnd.n6007 gnd.n6006 585
R4847 gnd.n6005 gnd.n6004 585
R4848 gnd.n6002 gnd.n5895 585
R4849 gnd.n5894 gnd.n5893 585
R4850 gnd.n5992 gnd.n5991 585
R4851 gnd.n5993 gnd.n5990 585
R4852 gnd.n5989 gnd.n5988 585
R4853 gnd.n5987 gnd.n5986 585
R4854 gnd.n5974 gnd.n5905 585
R4855 gnd.n5976 gnd.n5975 585
R4856 gnd.n5973 gnd.n5911 585
R4857 gnd.n5910 gnd.n5909 585
R4858 gnd.n5964 gnd.n5963 585
R4859 gnd.n5962 gnd.n5961 585
R4860 gnd.n5950 gnd.n5917 585
R4861 gnd.n5952 gnd.n5951 585
R4862 gnd.n5949 gnd.n5923 585
R4863 gnd.n5922 gnd.n5921 585
R4864 gnd.n5940 gnd.n5939 585
R4865 gnd.n5938 gnd.n5937 585
R4866 gnd.n5929 gnd.n1476 585
R4867 gnd.n6876 gnd.n847 475.807
R4868 gnd.n5680 gnd.n1994 463.671
R4869 gnd.n5689 gnd.n5688 463.671
R4870 gnd.n5176 gnd.n5174 463.671
R4871 gnd.n6542 gnd.n1339 463.671
R4872 gnd.n5110 gnd.t160 443.966
R4873 gnd.n1986 gnd.t203 443.966
R4874 gnd.n6479 gnd.t216 443.966
R4875 gnd.n5614 gnd.t236 443.966
R4876 gnd.n4844 gnd.t192 371.625
R4877 gnd.n122 gnd.t207 371.625
R4878 gnd.n5899 gnd.t219 371.625
R4879 gnd.n2448 gnd.t246 371.625
R4880 gnd.n1877 gnd.t189 371.625
R4881 gnd.n1899 gnd.t175 371.625
R4882 gnd.n201 gnd.t233 371.625
R4883 gnd.n7880 gnd.t156 371.625
R4884 gnd.n4178 gnd.t258 371.625
R4885 gnd.n4154 gnd.t229 371.625
R4886 gnd.n4350 gnd.t252 371.625
R4887 gnd.n4763 gnd.t249 371.625
R4888 gnd.n1297 gnd.t168 371.625
R4889 gnd.n5889 gnd.t164 371.625
R4890 gnd.n3167 gnd.t242 323.425
R4891 gnd.n2712 gnd.t182 323.425
R4892 gnd.n4015 gnd.n3989 289.615
R4893 gnd.n3983 gnd.n3957 289.615
R4894 gnd.n3951 gnd.n3925 289.615
R4895 gnd.n3920 gnd.n3894 289.615
R4896 gnd.n3888 gnd.n3862 289.615
R4897 gnd.n3856 gnd.n3830 289.615
R4898 gnd.n3824 gnd.n3798 289.615
R4899 gnd.n3793 gnd.n3767 289.615
R4900 gnd.n3241 gnd.t222 279.217
R4901 gnd.n2738 gnd.t196 279.217
R4902 gnd.n1346 gnd.t188 260.649
R4903 gnd.n5606 gnd.t181 260.649
R4904 gnd.n6544 gnd.n6543 256.663
R4905 gnd.n6544 gnd.n1305 256.663
R4906 gnd.n6544 gnd.n1306 256.663
R4907 gnd.n6544 gnd.n1307 256.663
R4908 gnd.n6544 gnd.n1308 256.663
R4909 gnd.n6544 gnd.n1309 256.663
R4910 gnd.n6544 gnd.n1310 256.663
R4911 gnd.n6544 gnd.n1311 256.663
R4912 gnd.n6544 gnd.n1312 256.663
R4913 gnd.n6544 gnd.n1313 256.663
R4914 gnd.n6544 gnd.n1314 256.663
R4915 gnd.n6544 gnd.n1315 256.663
R4916 gnd.n6544 gnd.n1316 256.663
R4917 gnd.n6544 gnd.n1317 256.663
R4918 gnd.n6544 gnd.n1318 256.663
R4919 gnd.n6544 gnd.n1319 256.663
R4920 gnd.n6547 gnd.n1303 256.663
R4921 gnd.n6545 gnd.n6544 256.663
R4922 gnd.n6544 gnd.n1320 256.663
R4923 gnd.n6544 gnd.n1321 256.663
R4924 gnd.n6544 gnd.n1322 256.663
R4925 gnd.n6544 gnd.n1323 256.663
R4926 gnd.n6544 gnd.n1324 256.663
R4927 gnd.n6544 gnd.n1325 256.663
R4928 gnd.n6544 gnd.n1326 256.663
R4929 gnd.n6544 gnd.n1327 256.663
R4930 gnd.n6544 gnd.n1328 256.663
R4931 gnd.n6544 gnd.n1329 256.663
R4932 gnd.n6544 gnd.n1330 256.663
R4933 gnd.n6544 gnd.n1331 256.663
R4934 gnd.n6544 gnd.n1332 256.663
R4935 gnd.n6544 gnd.n1333 256.663
R4936 gnd.n6544 gnd.n1334 256.663
R4937 gnd.n6544 gnd.n1335 256.663
R4938 gnd.n5755 gnd.n1818 256.663
R4939 gnd.n5755 gnd.n1819 256.663
R4940 gnd.n5755 gnd.n1820 256.663
R4941 gnd.n5755 gnd.n1821 256.663
R4942 gnd.n5755 gnd.n1822 256.663
R4943 gnd.n5755 gnd.n1823 256.663
R4944 gnd.n5755 gnd.n1824 256.663
R4945 gnd.n5755 gnd.n1825 256.663
R4946 gnd.n5755 gnd.n1826 256.663
R4947 gnd.n5755 gnd.n1827 256.663
R4948 gnd.n5755 gnd.n1828 256.663
R4949 gnd.n5755 gnd.n1829 256.663
R4950 gnd.n5755 gnd.n1830 256.663
R4951 gnd.n5755 gnd.n1831 256.663
R4952 gnd.n5755 gnd.n1832 256.663
R4953 gnd.n5755 gnd.n1833 256.663
R4954 gnd.n1985 gnd.n1834 256.663
R4955 gnd.n5755 gnd.n1817 256.663
R4956 gnd.n5755 gnd.n1816 256.663
R4957 gnd.n5755 gnd.n1815 256.663
R4958 gnd.n5755 gnd.n1814 256.663
R4959 gnd.n5755 gnd.n1813 256.663
R4960 gnd.n5755 gnd.n1812 256.663
R4961 gnd.n5755 gnd.n1811 256.663
R4962 gnd.n5755 gnd.n1810 256.663
R4963 gnd.n5755 gnd.n1809 256.663
R4964 gnd.n5755 gnd.n1808 256.663
R4965 gnd.n5755 gnd.n1807 256.663
R4966 gnd.n5755 gnd.n1806 256.663
R4967 gnd.n5755 gnd.n1805 256.663
R4968 gnd.n5755 gnd.n1804 256.663
R4969 gnd.n5755 gnd.n1803 256.663
R4970 gnd.n5755 gnd.n1802 256.663
R4971 gnd.n5755 gnd.n1801 256.663
R4972 gnd.n4434 gnd.n4148 242.672
R4973 gnd.n4432 gnd.n4148 242.672
R4974 gnd.n4426 gnd.n4148 242.672
R4975 gnd.n4424 gnd.n4148 242.672
R4976 gnd.n4418 gnd.n4148 242.672
R4977 gnd.n4416 gnd.n4148 242.672
R4978 gnd.n4410 gnd.n4148 242.672
R4979 gnd.n4408 gnd.n4148 242.672
R4980 gnd.n4398 gnd.n4148 242.672
R4981 gnd.n6577 gnd.n1261 242.672
R4982 gnd.n6577 gnd.n1260 242.672
R4983 gnd.n6577 gnd.n1259 242.672
R4984 gnd.n6577 gnd.n1258 242.672
R4985 gnd.n6577 gnd.n1257 242.672
R4986 gnd.n6577 gnd.n1256 242.672
R4987 gnd.n6577 gnd.n1255 242.672
R4988 gnd.n6577 gnd.n1254 242.672
R4989 gnd.n6577 gnd.n1253 242.672
R4990 gnd.n6041 gnd.n1710 242.672
R4991 gnd.n6041 gnd.n1711 242.672
R4992 gnd.n6041 gnd.n1712 242.672
R4993 gnd.n6041 gnd.n1713 242.672
R4994 gnd.n6041 gnd.n1714 242.672
R4995 gnd.n6041 gnd.n1715 242.672
R4996 gnd.n6041 gnd.n1716 242.672
R4997 gnd.n6041 gnd.n1717 242.672
R4998 gnd.n6041 gnd.n1718 242.672
R4999 gnd.n128 gnd.n125 242.672
R5000 gnd.n7805 gnd.n128 242.672
R5001 gnd.n7801 gnd.n128 242.672
R5002 gnd.n7798 gnd.n128 242.672
R5003 gnd.n7793 gnd.n128 242.672
R5004 gnd.n7790 gnd.n128 242.672
R5005 gnd.n7785 gnd.n128 242.672
R5006 gnd.n7782 gnd.n128 242.672
R5007 gnd.n7777 gnd.n128 242.672
R5008 gnd.n3295 gnd.n3294 242.672
R5009 gnd.n3295 gnd.n3205 242.672
R5010 gnd.n3295 gnd.n3206 242.672
R5011 gnd.n3295 gnd.n3207 242.672
R5012 gnd.n3295 gnd.n3208 242.672
R5013 gnd.n3295 gnd.n3209 242.672
R5014 gnd.n3295 gnd.n3210 242.672
R5015 gnd.n3295 gnd.n3211 242.672
R5016 gnd.n3295 gnd.n3212 242.672
R5017 gnd.n3295 gnd.n3213 242.672
R5018 gnd.n3295 gnd.n3214 242.672
R5019 gnd.n3295 gnd.n3215 242.672
R5020 gnd.n3296 gnd.n3295 242.672
R5021 gnd.n4147 gnd.n2687 242.672
R5022 gnd.n4147 gnd.n2686 242.672
R5023 gnd.n4147 gnd.n2685 242.672
R5024 gnd.n4147 gnd.n2684 242.672
R5025 gnd.n4147 gnd.n2683 242.672
R5026 gnd.n4147 gnd.n2682 242.672
R5027 gnd.n4147 gnd.n2681 242.672
R5028 gnd.n4147 gnd.n2680 242.672
R5029 gnd.n4147 gnd.n2679 242.672
R5030 gnd.n4147 gnd.n2678 242.672
R5031 gnd.n4147 gnd.n2677 242.672
R5032 gnd.n4147 gnd.n2676 242.672
R5033 gnd.n4147 gnd.n2675 242.672
R5034 gnd.n3379 gnd.n3378 242.672
R5035 gnd.n3378 gnd.n3117 242.672
R5036 gnd.n3378 gnd.n3118 242.672
R5037 gnd.n3378 gnd.n3119 242.672
R5038 gnd.n3378 gnd.n3120 242.672
R5039 gnd.n3378 gnd.n3121 242.672
R5040 gnd.n3378 gnd.n3122 242.672
R5041 gnd.n3378 gnd.n3123 242.672
R5042 gnd.n4147 gnd.n2688 242.672
R5043 gnd.n4147 gnd.n2689 242.672
R5044 gnd.n4147 gnd.n2690 242.672
R5045 gnd.n4147 gnd.n2691 242.672
R5046 gnd.n4147 gnd.n2692 242.672
R5047 gnd.n4147 gnd.n2693 242.672
R5048 gnd.n4147 gnd.n2694 242.672
R5049 gnd.n4147 gnd.n2695 242.672
R5050 gnd.n4196 gnd.n4148 242.672
R5051 gnd.n4204 gnd.n4148 242.672
R5052 gnd.n4206 gnd.n4148 242.672
R5053 gnd.n4214 gnd.n4148 242.672
R5054 gnd.n4216 gnd.n4148 242.672
R5055 gnd.n4224 gnd.n4148 242.672
R5056 gnd.n4226 gnd.n4148 242.672
R5057 gnd.n4234 gnd.n4148 242.672
R5058 gnd.n4236 gnd.n4148 242.672
R5059 gnd.n4244 gnd.n4148 242.672
R5060 gnd.n4246 gnd.n4148 242.672
R5061 gnd.n4254 gnd.n4148 242.672
R5062 gnd.n4256 gnd.n4148 242.672
R5063 gnd.n4264 gnd.n4148 242.672
R5064 gnd.n4266 gnd.n4148 242.672
R5065 gnd.n4274 gnd.n4148 242.672
R5066 gnd.n4276 gnd.n4148 242.672
R5067 gnd.n4285 gnd.n4148 242.672
R5068 gnd.n4288 gnd.n4148 242.672
R5069 gnd.n6577 gnd.n1263 242.672
R5070 gnd.n6577 gnd.n1264 242.672
R5071 gnd.n6577 gnd.n1265 242.672
R5072 gnd.n6577 gnd.n1266 242.672
R5073 gnd.n6577 gnd.n1267 242.672
R5074 gnd.n6577 gnd.n1268 242.672
R5075 gnd.n6577 gnd.n1269 242.672
R5076 gnd.n6577 gnd.n1270 242.672
R5077 gnd.n6577 gnd.n1271 242.672
R5078 gnd.n6577 gnd.n1272 242.672
R5079 gnd.n6577 gnd.n1273 242.672
R5080 gnd.n6548 gnd.n1299 242.672
R5081 gnd.n6577 gnd.n1274 242.672
R5082 gnd.n6577 gnd.n1275 242.672
R5083 gnd.n6577 gnd.n1276 242.672
R5084 gnd.n6577 gnd.n1277 242.672
R5085 gnd.n6577 gnd.n1278 242.672
R5086 gnd.n6577 gnd.n1279 242.672
R5087 gnd.n6577 gnd.n1280 242.672
R5088 gnd.n6577 gnd.n6576 242.672
R5089 gnd.n6042 gnd.n6041 242.672
R5090 gnd.n6041 gnd.n1691 242.672
R5091 gnd.n6041 gnd.n1692 242.672
R5092 gnd.n6041 gnd.n1693 242.672
R5093 gnd.n6041 gnd.n1694 242.672
R5094 gnd.n6041 gnd.n1695 242.672
R5095 gnd.n6041 gnd.n1696 242.672
R5096 gnd.n6041 gnd.n1697 242.672
R5097 gnd.n1984 gnd.n1836 242.672
R5098 gnd.n6041 gnd.n1698 242.672
R5099 gnd.n6041 gnd.n1699 242.672
R5100 gnd.n6041 gnd.n1700 242.672
R5101 gnd.n6041 gnd.n1701 242.672
R5102 gnd.n6041 gnd.n1702 242.672
R5103 gnd.n6041 gnd.n1703 242.672
R5104 gnd.n6041 gnd.n1704 242.672
R5105 gnd.n6041 gnd.n1705 242.672
R5106 gnd.n6041 gnd.n1706 242.672
R5107 gnd.n6041 gnd.n1707 242.672
R5108 gnd.n6041 gnd.n1708 242.672
R5109 gnd.n198 gnd.n128 242.672
R5110 gnd.n7848 gnd.n128 242.672
R5111 gnd.n194 gnd.n128 242.672
R5112 gnd.n7855 gnd.n128 242.672
R5113 gnd.n187 gnd.n128 242.672
R5114 gnd.n7862 gnd.n128 242.672
R5115 gnd.n180 gnd.n128 242.672
R5116 gnd.n7869 gnd.n128 242.672
R5117 gnd.n173 gnd.n128 242.672
R5118 gnd.n7876 gnd.n128 242.672
R5119 gnd.n166 gnd.n128 242.672
R5120 gnd.n7886 gnd.n128 242.672
R5121 gnd.n159 gnd.n128 242.672
R5122 gnd.n7893 gnd.n128 242.672
R5123 gnd.n152 gnd.n128 242.672
R5124 gnd.n7900 gnd.n128 242.672
R5125 gnd.n145 gnd.n128 242.672
R5126 gnd.n7907 gnd.n128 242.672
R5127 gnd.n138 gnd.n128 242.672
R5128 gnd.n4973 gnd.n4972 242.672
R5129 gnd.n4973 gnd.n2317 242.672
R5130 gnd.n4973 gnd.n2318 242.672
R5131 gnd.n4973 gnd.n2319 242.672
R5132 gnd.n4973 gnd.n2320 242.672
R5133 gnd.n4973 gnd.n2321 242.672
R5134 gnd.n4973 gnd.n2322 242.672
R5135 gnd.n4973 gnd.n2323 242.672
R5136 gnd.n4973 gnd.n2324 242.672
R5137 gnd.n4973 gnd.n2325 242.672
R5138 gnd.n4973 gnd.n2326 242.672
R5139 gnd.n4973 gnd.n2327 242.672
R5140 gnd.n4973 gnd.n2328 242.672
R5141 gnd.n4973 gnd.n2329 242.672
R5142 gnd.n6028 gnd.n6027 242.672
R5143 gnd.n6028 gnd.n5884 242.672
R5144 gnd.n6028 gnd.n5883 242.672
R5145 gnd.n6028 gnd.n5882 242.672
R5146 gnd.n6028 gnd.n5881 242.672
R5147 gnd.n6028 gnd.n5880 242.672
R5148 gnd.n6028 gnd.n5879 242.672
R5149 gnd.n6028 gnd.n5878 242.672
R5150 gnd.n6028 gnd.n5877 242.672
R5151 gnd.n6028 gnd.n5876 242.672
R5152 gnd.n6028 gnd.n5875 242.672
R5153 gnd.n6028 gnd.n5874 242.672
R5154 gnd.n6028 gnd.n5873 242.672
R5155 gnd.n6028 gnd.n5872 242.672
R5156 gnd.n135 gnd.n131 240.244
R5157 gnd.n7909 gnd.n7908 240.244
R5158 gnd.n7906 gnd.n139 240.244
R5159 gnd.n7902 gnd.n7901 240.244
R5160 gnd.n7899 gnd.n146 240.244
R5161 gnd.n7895 gnd.n7894 240.244
R5162 gnd.n7892 gnd.n153 240.244
R5163 gnd.n7888 gnd.n7887 240.244
R5164 gnd.n7885 gnd.n160 240.244
R5165 gnd.n7878 gnd.n7877 240.244
R5166 gnd.n7875 gnd.n167 240.244
R5167 gnd.n7871 gnd.n7870 240.244
R5168 gnd.n7868 gnd.n174 240.244
R5169 gnd.n7864 gnd.n7863 240.244
R5170 gnd.n7861 gnd.n181 240.244
R5171 gnd.n7857 gnd.n7856 240.244
R5172 gnd.n7854 gnd.n188 240.244
R5173 gnd.n7850 gnd.n7849 240.244
R5174 gnd.n7847 gnd.n195 240.244
R5175 gnd.n1903 gnd.n1683 240.244
R5176 gnd.n1903 gnd.n1676 240.244
R5177 gnd.n1676 gnd.n1666 240.244
R5178 gnd.n1935 gnd.n1666 240.244
R5179 gnd.n1935 gnd.n1657 240.244
R5180 gnd.n1932 gnd.n1657 240.244
R5181 gnd.n1932 gnd.n1649 240.244
R5182 gnd.n1649 gnd.n1640 240.244
R5183 gnd.n1927 gnd.n1640 240.244
R5184 gnd.n1927 gnd.n1631 240.244
R5185 gnd.n1924 gnd.n1631 240.244
R5186 gnd.n1924 gnd.n1623 240.244
R5187 gnd.n1623 gnd.n1612 240.244
R5188 gnd.n1920 gnd.n1612 240.244
R5189 gnd.n1920 gnd.n1601 240.244
R5190 gnd.n1601 gnd.n1592 240.244
R5191 gnd.n6164 gnd.n1592 240.244
R5192 gnd.n6164 gnd.n1575 240.244
R5193 gnd.n6167 gnd.n1575 240.244
R5194 gnd.n6167 gnd.n1568 240.244
R5195 gnd.n6203 gnd.n1568 240.244
R5196 gnd.n6203 gnd.n1559 240.244
R5197 gnd.n6199 gnd.n1559 240.244
R5198 gnd.n6199 gnd.n1550 240.244
R5199 gnd.n6196 gnd.n1550 240.244
R5200 gnd.n6196 gnd.n1522 240.244
R5201 gnd.n1522 gnd.n1516 240.244
R5202 gnd.n6191 gnd.n1516 240.244
R5203 gnd.n6191 gnd.n321 240.244
R5204 gnd.n6187 gnd.n321 240.244
R5205 gnd.n6187 gnd.n1532 240.244
R5206 gnd.n1536 gnd.n1532 240.244
R5207 gnd.n1536 gnd.n340 240.244
R5208 gnd.n7643 gnd.n340 240.244
R5209 gnd.n7643 gnd.n336 240.244
R5210 gnd.n7639 gnd.n336 240.244
R5211 gnd.n7639 gnd.n307 240.244
R5212 gnd.n7634 gnd.n307 240.244
R5213 gnd.n7634 gnd.n299 240.244
R5214 gnd.n7630 gnd.n299 240.244
R5215 gnd.n7630 gnd.n292 240.244
R5216 gnd.n7625 gnd.n292 240.244
R5217 gnd.n7625 gnd.n284 240.244
R5218 gnd.n399 gnd.n284 240.244
R5219 gnd.n399 gnd.n276 240.244
R5220 gnd.n394 gnd.n276 240.244
R5221 gnd.n394 gnd.n267 240.244
R5222 gnd.n390 gnd.n267 240.244
R5223 gnd.n390 gnd.n260 240.244
R5224 gnd.n387 gnd.n260 240.244
R5225 gnd.n387 gnd.n253 240.244
R5226 gnd.n384 gnd.n253 240.244
R5227 gnd.n384 gnd.n245 240.244
R5228 gnd.n381 gnd.n245 240.244
R5229 gnd.n381 gnd.n237 240.244
R5230 gnd.n378 gnd.n237 240.244
R5231 gnd.n378 gnd.n231 240.244
R5232 gnd.n375 gnd.n231 240.244
R5233 gnd.n375 gnd.n223 240.244
R5234 gnd.n372 gnd.n223 240.244
R5235 gnd.n372 gnd.n214 240.244
R5236 gnd.n214 gnd.n205 240.244
R5237 gnd.n7839 gnd.n205 240.244
R5238 gnd.n7839 gnd.n127 240.244
R5239 gnd.n6043 gnd.n1689 240.244
R5240 gnd.n1842 gnd.n1689 240.244
R5241 gnd.n1849 gnd.n1848 240.244
R5242 gnd.n1852 gnd.n1851 240.244
R5243 gnd.n1859 gnd.n1858 240.244
R5244 gnd.n1862 gnd.n1861 240.244
R5245 gnd.n1869 gnd.n1868 240.244
R5246 gnd.n1872 gnd.n1871 240.244
R5247 gnd.n1982 gnd.n1981 240.244
R5248 gnd.n1978 gnd.n1977 240.244
R5249 gnd.n1974 gnd.n1973 240.244
R5250 gnd.n1970 gnd.n1969 240.244
R5251 gnd.n1966 gnd.n1965 240.244
R5252 gnd.n1962 gnd.n1961 240.244
R5253 gnd.n1958 gnd.n1957 240.244
R5254 gnd.n1954 gnd.n1953 240.244
R5255 gnd.n1950 gnd.n1949 240.244
R5256 gnd.n1898 gnd.n1897 240.244
R5257 gnd.n6051 gnd.n1686 240.244
R5258 gnd.n1686 gnd.n1664 240.244
R5259 gnd.n6075 gnd.n1664 240.244
R5260 gnd.n6075 gnd.n1659 240.244
R5261 gnd.n6083 gnd.n1659 240.244
R5262 gnd.n6083 gnd.n1660 240.244
R5263 gnd.n1660 gnd.n1638 240.244
R5264 gnd.n6107 gnd.n1638 240.244
R5265 gnd.n6107 gnd.n1633 240.244
R5266 gnd.n6115 gnd.n1633 240.244
R5267 gnd.n6115 gnd.n1634 240.244
R5268 gnd.n1634 gnd.n1610 240.244
R5269 gnd.n6145 gnd.n1610 240.244
R5270 gnd.n6145 gnd.n1604 240.244
R5271 gnd.n6153 gnd.n1604 240.244
R5272 gnd.n6153 gnd.n1606 240.244
R5273 gnd.n1606 gnd.n1573 240.244
R5274 gnd.n6213 gnd.n1573 240.244
R5275 gnd.n6213 gnd.n1569 240.244
R5276 gnd.n6219 gnd.n1569 240.244
R5277 gnd.n6219 gnd.n1557 240.244
R5278 gnd.n6233 gnd.n1557 240.244
R5279 gnd.n6233 gnd.n1553 240.244
R5280 gnd.n6241 gnd.n1553 240.244
R5281 gnd.n6241 gnd.n1519 240.244
R5282 gnd.n6303 gnd.n1519 240.244
R5283 gnd.n6304 gnd.n6303 240.244
R5284 gnd.n6304 gnd.n318 240.244
R5285 gnd.n7664 gnd.n318 240.244
R5286 gnd.n7664 gnd.n319 240.244
R5287 gnd.n6289 gnd.n319 240.244
R5288 gnd.n6289 gnd.n6286 240.244
R5289 gnd.n6286 gnd.n338 240.244
R5290 gnd.n7645 gnd.n338 240.244
R5291 gnd.n7648 gnd.n7645 240.244
R5292 gnd.n7648 gnd.n309 240.244
R5293 gnd.n7670 gnd.n309 240.244
R5294 gnd.n7670 gnd.n297 240.244
R5295 gnd.n7680 gnd.n297 240.244
R5296 gnd.n7680 gnd.n293 240.244
R5297 gnd.n7686 gnd.n293 240.244
R5298 gnd.n7686 gnd.n282 240.244
R5299 gnd.n7696 gnd.n282 240.244
R5300 gnd.n7696 gnd.n278 240.244
R5301 gnd.n7702 gnd.n278 240.244
R5302 gnd.n7702 gnd.n265 240.244
R5303 gnd.n7712 gnd.n265 240.244
R5304 gnd.n7712 gnd.n261 240.244
R5305 gnd.n7718 gnd.n261 240.244
R5306 gnd.n7718 gnd.n251 240.244
R5307 gnd.n7728 gnd.n251 240.244
R5308 gnd.n7728 gnd.n247 240.244
R5309 gnd.n7734 gnd.n247 240.244
R5310 gnd.n7734 gnd.n236 240.244
R5311 gnd.n7744 gnd.n236 240.244
R5312 gnd.n7744 gnd.n232 240.244
R5313 gnd.n7750 gnd.n232 240.244
R5314 gnd.n7750 gnd.n221 240.244
R5315 gnd.n7760 gnd.n221 240.244
R5316 gnd.n7760 gnd.n216 240.244
R5317 gnd.n7768 gnd.n216 240.244
R5318 gnd.n7768 gnd.n217 240.244
R5319 gnd.n217 gnd.n130 240.244
R5320 gnd.n7916 gnd.n130 240.244
R5321 gnd.n6578 gnd.n1250 240.244
R5322 gnd.n6575 gnd.n1281 240.244
R5323 gnd.n6571 gnd.n6570 240.244
R5324 gnd.n6567 gnd.n6566 240.244
R5325 gnd.n6563 gnd.n6562 240.244
R5326 gnd.n6559 gnd.n6558 240.244
R5327 gnd.n6555 gnd.n6554 240.244
R5328 gnd.n6551 gnd.n6550 240.244
R5329 gnd.n4775 gnd.n4774 240.244
R5330 gnd.n4782 gnd.n4781 240.244
R5331 gnd.n4785 gnd.n4784 240.244
R5332 gnd.n4792 gnd.n4791 240.244
R5333 gnd.n4795 gnd.n4794 240.244
R5334 gnd.n4802 gnd.n4801 240.244
R5335 gnd.n4805 gnd.n4804 240.244
R5336 gnd.n4812 gnd.n4811 240.244
R5337 gnd.n4815 gnd.n4814 240.244
R5338 gnd.n4820 gnd.n4765 240.244
R5339 gnd.n4324 gnd.n4149 240.244
R5340 gnd.n4324 gnd.n2667 240.244
R5341 gnd.n4318 gnd.n2667 240.244
R5342 gnd.n4318 gnd.n2660 240.244
R5343 gnd.n4315 gnd.n2660 240.244
R5344 gnd.n4315 gnd.n2652 240.244
R5345 gnd.n4312 gnd.n2652 240.244
R5346 gnd.n4312 gnd.n2643 240.244
R5347 gnd.n4309 gnd.n2643 240.244
R5348 gnd.n4309 gnd.n2635 240.244
R5349 gnd.n4306 gnd.n2635 240.244
R5350 gnd.n4306 gnd.n2627 240.244
R5351 gnd.n2627 gnd.n2617 240.244
R5352 gnd.n4510 gnd.n2617 240.244
R5353 gnd.n4511 gnd.n4510 240.244
R5354 gnd.n4511 gnd.n1020 240.244
R5355 gnd.n4514 gnd.n1020 240.244
R5356 gnd.n4514 gnd.n1033 240.244
R5357 gnd.n4520 gnd.n1033 240.244
R5358 gnd.n4520 gnd.n1045 240.244
R5359 gnd.n4530 gnd.n1045 240.244
R5360 gnd.n4530 gnd.n1055 240.244
R5361 gnd.n4541 gnd.n1055 240.244
R5362 gnd.n4541 gnd.n1066 240.244
R5363 gnd.n2579 gnd.n1066 240.244
R5364 gnd.n2579 gnd.n1076 240.244
R5365 gnd.n4568 gnd.n1076 240.244
R5366 gnd.n4568 gnd.n1087 240.244
R5367 gnd.n4564 gnd.n1087 240.244
R5368 gnd.n4564 gnd.n2552 240.244
R5369 gnd.n2571 gnd.n2552 240.244
R5370 gnd.n2571 gnd.n2549 240.244
R5371 gnd.n2549 gnd.n2543 240.244
R5372 gnd.n2543 gnd.n2533 240.244
R5373 gnd.n2533 gnd.n2527 240.244
R5374 gnd.n4639 gnd.n2527 240.244
R5375 gnd.n4639 gnd.n1102 240.244
R5376 gnd.n2513 gnd.n1102 240.244
R5377 gnd.n2513 gnd.n1113 240.244
R5378 gnd.n4647 gnd.n1113 240.244
R5379 gnd.n4647 gnd.n1123 240.244
R5380 gnd.n4651 gnd.n1123 240.244
R5381 gnd.n4651 gnd.n1134 240.244
R5382 gnd.n4661 gnd.n1134 240.244
R5383 gnd.n4661 gnd.n1145 240.244
R5384 gnd.n2501 gnd.n1145 240.244
R5385 gnd.n2501 gnd.n1155 240.244
R5386 gnd.n4722 gnd.n1155 240.244
R5387 gnd.n4722 gnd.n1166 240.244
R5388 gnd.n4728 gnd.n1166 240.244
R5389 gnd.n4728 gnd.n1177 240.244
R5390 gnd.n4738 gnd.n1177 240.244
R5391 gnd.n4738 gnd.n1188 240.244
R5392 gnd.n2475 gnd.n1188 240.244
R5393 gnd.n2475 gnd.n1198 240.244
R5394 gnd.n4746 gnd.n1198 240.244
R5395 gnd.n4746 gnd.n1209 240.244
R5396 gnd.n4752 gnd.n1209 240.244
R5397 gnd.n4752 gnd.n1220 240.244
R5398 gnd.n4756 gnd.n1220 240.244
R5399 gnd.n4756 gnd.n1231 240.244
R5400 gnd.n4830 gnd.n1231 240.244
R5401 gnd.n4830 gnd.n1242 240.244
R5402 gnd.n2460 gnd.n1242 240.244
R5403 gnd.n4197 gnd.n4193 240.244
R5404 gnd.n4203 gnd.n4193 240.244
R5405 gnd.n4207 gnd.n4205 240.244
R5406 gnd.n4213 gnd.n4189 240.244
R5407 gnd.n4217 gnd.n4215 240.244
R5408 gnd.n4223 gnd.n4185 240.244
R5409 gnd.n4227 gnd.n4225 240.244
R5410 gnd.n4233 gnd.n4181 240.244
R5411 gnd.n4237 gnd.n4235 240.244
R5412 gnd.n4243 gnd.n4174 240.244
R5413 gnd.n4247 gnd.n4245 240.244
R5414 gnd.n4253 gnd.n4170 240.244
R5415 gnd.n4257 gnd.n4255 240.244
R5416 gnd.n4263 gnd.n4166 240.244
R5417 gnd.n4267 gnd.n4265 240.244
R5418 gnd.n4273 gnd.n4162 240.244
R5419 gnd.n4277 gnd.n4275 240.244
R5420 gnd.n4284 gnd.n4158 240.244
R5421 gnd.n4287 gnd.n4286 240.244
R5422 gnd.n4443 gnd.n2669 240.244
R5423 gnd.n4449 gnd.n2669 240.244
R5424 gnd.n4449 gnd.n2658 240.244
R5425 gnd.n4459 gnd.n2658 240.244
R5426 gnd.n4459 gnd.n2654 240.244
R5427 gnd.n4465 gnd.n2654 240.244
R5428 gnd.n4465 gnd.n2641 240.244
R5429 gnd.n4475 gnd.n2641 240.244
R5430 gnd.n4475 gnd.n2637 240.244
R5431 gnd.n4481 gnd.n2637 240.244
R5432 gnd.n4481 gnd.n2625 240.244
R5433 gnd.n4501 gnd.n2625 240.244
R5434 gnd.n4501 gnd.n2621 240.244
R5435 gnd.n4508 gnd.n2621 240.244
R5436 gnd.n4508 gnd.n1024 240.244
R5437 gnd.n6706 gnd.n1024 240.244
R5438 gnd.n6706 gnd.n1025 240.244
R5439 gnd.n6702 gnd.n1025 240.244
R5440 gnd.n6702 gnd.n1031 240.244
R5441 gnd.n6694 gnd.n1031 240.244
R5442 gnd.n6694 gnd.n1047 240.244
R5443 gnd.n6690 gnd.n1047 240.244
R5444 gnd.n6690 gnd.n1053 240.244
R5445 gnd.n6682 gnd.n1053 240.244
R5446 gnd.n6682 gnd.n1069 240.244
R5447 gnd.n6678 gnd.n1069 240.244
R5448 gnd.n6678 gnd.n1075 240.244
R5449 gnd.n6670 gnd.n1075 240.244
R5450 gnd.n6670 gnd.n1089 240.244
R5451 gnd.n4591 gnd.n1089 240.244
R5452 gnd.n4593 gnd.n4591 240.244
R5453 gnd.n4596 gnd.n4593 240.244
R5454 gnd.n4596 gnd.n2536 240.244
R5455 gnd.n4629 gnd.n2536 240.244
R5456 gnd.n4629 gnd.n4626 240.244
R5457 gnd.n4626 gnd.n1099 240.244
R5458 gnd.n6664 gnd.n1099 240.244
R5459 gnd.n6664 gnd.n1100 240.244
R5460 gnd.n6656 gnd.n1100 240.244
R5461 gnd.n6656 gnd.n1116 240.244
R5462 gnd.n6652 gnd.n1116 240.244
R5463 gnd.n6652 gnd.n1121 240.244
R5464 gnd.n6644 gnd.n1121 240.244
R5465 gnd.n6644 gnd.n1137 240.244
R5466 gnd.n6640 gnd.n1137 240.244
R5467 gnd.n6640 gnd.n1143 240.244
R5468 gnd.n6632 gnd.n1143 240.244
R5469 gnd.n6632 gnd.n1158 240.244
R5470 gnd.n6628 gnd.n1158 240.244
R5471 gnd.n6628 gnd.n1164 240.244
R5472 gnd.n6620 gnd.n1164 240.244
R5473 gnd.n6620 gnd.n1180 240.244
R5474 gnd.n6616 gnd.n1180 240.244
R5475 gnd.n6616 gnd.n1186 240.244
R5476 gnd.n6608 gnd.n1186 240.244
R5477 gnd.n6608 gnd.n1201 240.244
R5478 gnd.n6604 gnd.n1201 240.244
R5479 gnd.n6604 gnd.n1207 240.244
R5480 gnd.n6596 gnd.n1207 240.244
R5481 gnd.n6596 gnd.n1223 240.244
R5482 gnd.n6592 gnd.n1223 240.244
R5483 gnd.n6592 gnd.n1229 240.244
R5484 gnd.n6584 gnd.n1229 240.244
R5485 gnd.n6584 gnd.n1245 240.244
R5486 gnd.n4146 gnd.n2697 240.244
R5487 gnd.n4139 gnd.n4138 240.244
R5488 gnd.n4136 gnd.n4135 240.244
R5489 gnd.n4132 gnd.n4131 240.244
R5490 gnd.n4128 gnd.n4127 240.244
R5491 gnd.n4124 gnd.n4123 240.244
R5492 gnd.n4120 gnd.n4119 240.244
R5493 gnd.n4116 gnd.n4115 240.244
R5494 gnd.n3390 gnd.n3102 240.244
R5495 gnd.n3400 gnd.n3102 240.244
R5496 gnd.n3400 gnd.n3093 240.244
R5497 gnd.n3093 gnd.n3082 240.244
R5498 gnd.n3421 gnd.n3082 240.244
R5499 gnd.n3421 gnd.n3076 240.244
R5500 gnd.n3431 gnd.n3076 240.244
R5501 gnd.n3431 gnd.n3065 240.244
R5502 gnd.n3065 gnd.n3057 240.244
R5503 gnd.n3449 gnd.n3057 240.244
R5504 gnd.n3450 gnd.n3449 240.244
R5505 gnd.n3450 gnd.n3042 240.244
R5506 gnd.n3452 gnd.n3042 240.244
R5507 gnd.n3452 gnd.n3028 240.244
R5508 gnd.n3494 gnd.n3028 240.244
R5509 gnd.n3495 gnd.n3494 240.244
R5510 gnd.n3498 gnd.n3495 240.244
R5511 gnd.n3498 gnd.n2983 240.244
R5512 gnd.n3023 gnd.n2983 240.244
R5513 gnd.n3023 gnd.n2993 240.244
R5514 gnd.n3508 gnd.n2993 240.244
R5515 gnd.n3508 gnd.n3014 240.244
R5516 gnd.n3518 gnd.n3014 240.244
R5517 gnd.n3518 gnd.n2900 240.244
R5518 gnd.n3563 gnd.n2900 240.244
R5519 gnd.n3563 gnd.n2886 240.244
R5520 gnd.n3585 gnd.n2886 240.244
R5521 gnd.n3586 gnd.n3585 240.244
R5522 gnd.n3586 gnd.n2873 240.244
R5523 gnd.n2873 gnd.n2862 240.244
R5524 gnd.n3617 gnd.n2862 240.244
R5525 gnd.n3618 gnd.n3617 240.244
R5526 gnd.n3619 gnd.n3618 240.244
R5527 gnd.n3619 gnd.n2847 240.244
R5528 gnd.n2847 gnd.n2846 240.244
R5529 gnd.n2846 gnd.n2831 240.244
R5530 gnd.n3670 gnd.n2831 240.244
R5531 gnd.n3671 gnd.n3670 240.244
R5532 gnd.n3671 gnd.n2818 240.244
R5533 gnd.n2818 gnd.n2807 240.244
R5534 gnd.n3702 gnd.n2807 240.244
R5535 gnd.n3703 gnd.n3702 240.244
R5536 gnd.n3704 gnd.n3703 240.244
R5537 gnd.n3704 gnd.n2791 240.244
R5538 gnd.n2791 gnd.n2790 240.244
R5539 gnd.n2790 gnd.n2776 240.244
R5540 gnd.n3759 gnd.n2776 240.244
R5541 gnd.n3760 gnd.n3759 240.244
R5542 gnd.n3760 gnd.n2763 240.244
R5543 gnd.n2763 gnd.n2753 240.244
R5544 gnd.n4047 gnd.n2753 240.244
R5545 gnd.n4050 gnd.n4047 240.244
R5546 gnd.n4050 gnd.n4049 240.244
R5547 gnd.n3380 gnd.n3115 240.244
R5548 gnd.n3136 gnd.n3115 240.244
R5549 gnd.n3139 gnd.n3138 240.244
R5550 gnd.n3146 gnd.n3145 240.244
R5551 gnd.n3149 gnd.n3148 240.244
R5552 gnd.n3156 gnd.n3155 240.244
R5553 gnd.n3159 gnd.n3158 240.244
R5554 gnd.n3166 gnd.n3165 240.244
R5555 gnd.n3388 gnd.n3112 240.244
R5556 gnd.n3112 gnd.n3091 240.244
R5557 gnd.n3411 gnd.n3091 240.244
R5558 gnd.n3411 gnd.n3085 240.244
R5559 gnd.n3419 gnd.n3085 240.244
R5560 gnd.n3419 gnd.n3087 240.244
R5561 gnd.n3087 gnd.n3063 240.244
R5562 gnd.n3441 gnd.n3063 240.244
R5563 gnd.n3441 gnd.n3059 240.244
R5564 gnd.n3447 gnd.n3059 240.244
R5565 gnd.n3447 gnd.n3041 240.244
R5566 gnd.n3472 gnd.n3041 240.244
R5567 gnd.n3472 gnd.n3036 240.244
R5568 gnd.n3484 gnd.n3036 240.244
R5569 gnd.n3484 gnd.n3037 240.244
R5570 gnd.n3480 gnd.n3037 240.244
R5571 gnd.n3480 gnd.n2985 240.244
R5572 gnd.n3532 gnd.n2985 240.244
R5573 gnd.n3532 gnd.n2986 240.244
R5574 gnd.n3528 gnd.n2986 240.244
R5575 gnd.n3528 gnd.n2992 240.244
R5576 gnd.n3012 gnd.n2992 240.244
R5577 gnd.n3012 gnd.n2898 240.244
R5578 gnd.n3567 gnd.n2898 240.244
R5579 gnd.n3567 gnd.n2893 240.244
R5580 gnd.n3575 gnd.n2893 240.244
R5581 gnd.n3575 gnd.n2894 240.244
R5582 gnd.n2894 gnd.n2871 240.244
R5583 gnd.n3607 gnd.n2871 240.244
R5584 gnd.n3607 gnd.n2866 240.244
R5585 gnd.n3615 gnd.n2866 240.244
R5586 gnd.n3615 gnd.n2867 240.244
R5587 gnd.n2867 gnd.n2844 240.244
R5588 gnd.n3652 gnd.n2844 240.244
R5589 gnd.n3652 gnd.n2839 240.244
R5590 gnd.n3660 gnd.n2839 240.244
R5591 gnd.n3660 gnd.n2840 240.244
R5592 gnd.n2840 gnd.n2816 240.244
R5593 gnd.n3692 gnd.n2816 240.244
R5594 gnd.n3692 gnd.n2811 240.244
R5595 gnd.n3700 gnd.n2811 240.244
R5596 gnd.n3700 gnd.n2812 240.244
R5597 gnd.n2812 gnd.n2788 240.244
R5598 gnd.n3741 gnd.n2788 240.244
R5599 gnd.n3741 gnd.n2783 240.244
R5600 gnd.n3749 gnd.n2783 240.244
R5601 gnd.n3749 gnd.n2784 240.244
R5602 gnd.n2784 gnd.n2761 240.244
R5603 gnd.n4035 gnd.n2761 240.244
R5604 gnd.n4035 gnd.n2756 240.244
R5605 gnd.n4045 gnd.n2756 240.244
R5606 gnd.n4045 gnd.n2757 240.244
R5607 gnd.n2757 gnd.n2696 240.244
R5608 gnd.n2716 gnd.n2674 240.244
R5609 gnd.n4106 gnd.n4105 240.244
R5610 gnd.n4102 gnd.n4101 240.244
R5611 gnd.n4098 gnd.n4097 240.244
R5612 gnd.n4094 gnd.n4093 240.244
R5613 gnd.n4090 gnd.n4089 240.244
R5614 gnd.n4086 gnd.n4085 240.244
R5615 gnd.n4082 gnd.n4081 240.244
R5616 gnd.n4078 gnd.n4077 240.244
R5617 gnd.n4074 gnd.n4073 240.244
R5618 gnd.n4070 gnd.n4069 240.244
R5619 gnd.n4066 gnd.n4065 240.244
R5620 gnd.n4062 gnd.n4061 240.244
R5621 gnd.n3303 gnd.n3200 240.244
R5622 gnd.n3303 gnd.n3193 240.244
R5623 gnd.n3314 gnd.n3193 240.244
R5624 gnd.n3314 gnd.n3189 240.244
R5625 gnd.n3320 gnd.n3189 240.244
R5626 gnd.n3320 gnd.n3181 240.244
R5627 gnd.n3330 gnd.n3181 240.244
R5628 gnd.n3330 gnd.n3176 240.244
R5629 gnd.n3366 gnd.n3176 240.244
R5630 gnd.n3366 gnd.n3177 240.244
R5631 gnd.n3177 gnd.n3124 240.244
R5632 gnd.n3361 gnd.n3124 240.244
R5633 gnd.n3361 gnd.n3360 240.244
R5634 gnd.n3360 gnd.n3103 240.244
R5635 gnd.n3356 gnd.n3103 240.244
R5636 gnd.n3356 gnd.n3094 240.244
R5637 gnd.n3353 gnd.n3094 240.244
R5638 gnd.n3353 gnd.n3352 240.244
R5639 gnd.n3352 gnd.n3077 240.244
R5640 gnd.n3348 gnd.n3077 240.244
R5641 gnd.n3348 gnd.n3066 240.244
R5642 gnd.n3066 gnd.n3047 240.244
R5643 gnd.n3461 gnd.n3047 240.244
R5644 gnd.n3461 gnd.n3043 240.244
R5645 gnd.n3469 gnd.n3043 240.244
R5646 gnd.n3469 gnd.n3034 240.244
R5647 gnd.n3034 gnd.n2970 240.244
R5648 gnd.n3541 gnd.n2970 240.244
R5649 gnd.n3541 gnd.n2971 240.244
R5650 gnd.n2982 gnd.n2971 240.244
R5651 gnd.n3017 gnd.n2982 240.244
R5652 gnd.n3020 gnd.n3017 240.244
R5653 gnd.n3020 gnd.n2994 240.244
R5654 gnd.n3007 gnd.n2994 240.244
R5655 gnd.n3007 gnd.n3004 240.244
R5656 gnd.n3004 gnd.n2901 240.244
R5657 gnd.n3562 gnd.n2901 240.244
R5658 gnd.n3562 gnd.n2891 240.244
R5659 gnd.n3558 gnd.n2891 240.244
R5660 gnd.n3558 gnd.n2885 240.244
R5661 gnd.n3555 gnd.n2885 240.244
R5662 gnd.n3555 gnd.n2874 240.244
R5663 gnd.n3552 gnd.n2874 240.244
R5664 gnd.n3552 gnd.n2852 240.244
R5665 gnd.n3628 gnd.n2852 240.244
R5666 gnd.n3628 gnd.n2848 240.244
R5667 gnd.n3649 gnd.n2848 240.244
R5668 gnd.n3649 gnd.n2837 240.244
R5669 gnd.n3645 gnd.n2837 240.244
R5670 gnd.n3645 gnd.n2830 240.244
R5671 gnd.n3642 gnd.n2830 240.244
R5672 gnd.n3642 gnd.n2819 240.244
R5673 gnd.n3639 gnd.n2819 240.244
R5674 gnd.n3639 gnd.n2796 240.244
R5675 gnd.n3713 gnd.n2796 240.244
R5676 gnd.n3713 gnd.n2792 240.244
R5677 gnd.n3738 gnd.n2792 240.244
R5678 gnd.n3738 gnd.n2782 240.244
R5679 gnd.n3734 gnd.n2782 240.244
R5680 gnd.n3734 gnd.n2775 240.244
R5681 gnd.n3730 gnd.n2775 240.244
R5682 gnd.n3730 gnd.n2764 240.244
R5683 gnd.n3727 gnd.n2764 240.244
R5684 gnd.n3727 gnd.n2745 240.244
R5685 gnd.n4057 gnd.n2745 240.244
R5686 gnd.n3217 gnd.n3216 240.244
R5687 gnd.n3288 gnd.n3216 240.244
R5688 gnd.n3286 gnd.n3285 240.244
R5689 gnd.n3282 gnd.n3281 240.244
R5690 gnd.n3278 gnd.n3277 240.244
R5691 gnd.n3274 gnd.n3273 240.244
R5692 gnd.n3270 gnd.n3269 240.244
R5693 gnd.n3266 gnd.n3265 240.244
R5694 gnd.n3262 gnd.n3261 240.244
R5695 gnd.n3258 gnd.n3257 240.244
R5696 gnd.n3254 gnd.n3253 240.244
R5697 gnd.n3250 gnd.n3249 240.244
R5698 gnd.n3246 gnd.n3204 240.244
R5699 gnd.n3306 gnd.n3198 240.244
R5700 gnd.n3306 gnd.n3194 240.244
R5701 gnd.n3312 gnd.n3194 240.244
R5702 gnd.n3312 gnd.n3187 240.244
R5703 gnd.n3322 gnd.n3187 240.244
R5704 gnd.n3322 gnd.n3183 240.244
R5705 gnd.n3328 gnd.n3183 240.244
R5706 gnd.n3328 gnd.n3174 240.244
R5707 gnd.n3368 gnd.n3174 240.244
R5708 gnd.n3368 gnd.n3125 240.244
R5709 gnd.n3376 gnd.n3125 240.244
R5710 gnd.n3376 gnd.n3126 240.244
R5711 gnd.n3126 gnd.n3104 240.244
R5712 gnd.n3397 gnd.n3104 240.244
R5713 gnd.n3397 gnd.n3096 240.244
R5714 gnd.n3408 gnd.n3096 240.244
R5715 gnd.n3408 gnd.n3097 240.244
R5716 gnd.n3097 gnd.n3078 240.244
R5717 gnd.n3428 gnd.n3078 240.244
R5718 gnd.n3428 gnd.n3068 240.244
R5719 gnd.n3438 gnd.n3068 240.244
R5720 gnd.n3438 gnd.n3049 240.244
R5721 gnd.n3459 gnd.n3049 240.244
R5722 gnd.n3459 gnd.n3051 240.244
R5723 gnd.n3051 gnd.n3032 240.244
R5724 gnd.n3487 gnd.n3032 240.244
R5725 gnd.n3487 gnd.n2974 240.244
R5726 gnd.n3539 gnd.n2974 240.244
R5727 gnd.n3539 gnd.n2975 240.244
R5728 gnd.n3535 gnd.n2975 240.244
R5729 gnd.n3535 gnd.n2981 240.244
R5730 gnd.n2996 gnd.n2981 240.244
R5731 gnd.n3525 gnd.n2996 240.244
R5732 gnd.n3525 gnd.n2997 240.244
R5733 gnd.n3521 gnd.n2997 240.244
R5734 gnd.n3521 gnd.n3003 240.244
R5735 gnd.n3003 gnd.n2890 240.244
R5736 gnd.n3578 gnd.n2890 240.244
R5737 gnd.n3578 gnd.n2883 240.244
R5738 gnd.n3589 gnd.n2883 240.244
R5739 gnd.n3589 gnd.n2876 240.244
R5740 gnd.n3604 gnd.n2876 240.244
R5741 gnd.n3604 gnd.n2877 240.244
R5742 gnd.n2877 gnd.n2855 240.244
R5743 gnd.n3626 gnd.n2855 240.244
R5744 gnd.n3626 gnd.n2856 240.244
R5745 gnd.n2856 gnd.n2835 240.244
R5746 gnd.n3663 gnd.n2835 240.244
R5747 gnd.n3663 gnd.n2828 240.244
R5748 gnd.n3674 gnd.n2828 240.244
R5749 gnd.n3674 gnd.n2821 240.244
R5750 gnd.n3689 gnd.n2821 240.244
R5751 gnd.n3689 gnd.n2822 240.244
R5752 gnd.n2822 gnd.n2799 240.244
R5753 gnd.n3711 gnd.n2799 240.244
R5754 gnd.n3711 gnd.n2801 240.244
R5755 gnd.n2801 gnd.n2780 240.244
R5756 gnd.n3752 gnd.n2780 240.244
R5757 gnd.n3752 gnd.n2773 240.244
R5758 gnd.n3763 gnd.n2773 240.244
R5759 gnd.n3763 gnd.n2766 240.244
R5760 gnd.n4032 gnd.n2766 240.244
R5761 gnd.n4032 gnd.n2767 240.244
R5762 gnd.n2767 gnd.n2748 240.244
R5763 gnd.n4055 gnd.n2748 240.244
R5764 gnd.n7776 gnd.n7775 240.244
R5765 gnd.n7781 gnd.n7778 240.244
R5766 gnd.n7784 gnd.n7783 240.244
R5767 gnd.n7789 gnd.n7786 240.244
R5768 gnd.n7792 gnd.n7791 240.244
R5769 gnd.n7797 gnd.n7794 240.244
R5770 gnd.n7800 gnd.n7799 240.244
R5771 gnd.n7804 gnd.n7802 240.244
R5772 gnd.n7807 gnd.n7806 240.244
R5773 gnd.n6053 gnd.n1677 240.244
R5774 gnd.n6060 gnd.n1677 240.244
R5775 gnd.n6060 gnd.n1667 240.244
R5776 gnd.n1667 gnd.n1655 240.244
R5777 gnd.n6085 gnd.n1655 240.244
R5778 gnd.n6085 gnd.n1650 240.244
R5779 gnd.n6092 gnd.n1650 240.244
R5780 gnd.n6092 gnd.n1641 240.244
R5781 gnd.n1641 gnd.n1629 240.244
R5782 gnd.n6117 gnd.n1629 240.244
R5783 gnd.n6117 gnd.n1624 240.244
R5784 gnd.n6124 gnd.n1624 240.244
R5785 gnd.n6124 gnd.n1613 240.244
R5786 gnd.n1613 gnd.n1599 240.244
R5787 gnd.n6155 gnd.n1599 240.244
R5788 gnd.n6155 gnd.n1594 240.244
R5789 gnd.n6162 gnd.n1594 240.244
R5790 gnd.n6162 gnd.n1576 240.244
R5791 gnd.n1576 gnd.n1566 240.244
R5792 gnd.n6221 gnd.n1566 240.244
R5793 gnd.n6221 gnd.n1560 240.244
R5794 gnd.n6230 gnd.n1560 240.244
R5795 gnd.n6230 gnd.n1561 240.244
R5796 gnd.n1561 gnd.n1551 240.244
R5797 gnd.n1551 gnd.n1523 240.244
R5798 gnd.n6301 gnd.n1523 240.244
R5799 gnd.n6301 gnd.n1517 240.244
R5800 gnd.n1528 gnd.n1517 240.244
R5801 gnd.n1528 gnd.n322 240.244
R5802 gnd.n1529 gnd.n322 240.244
R5803 gnd.n6291 gnd.n1529 240.244
R5804 gnd.n6291 gnd.n1530 240.244
R5805 gnd.n1530 gnd.n82 240.244
R5806 gnd.n83 gnd.n82 240.244
R5807 gnd.n84 gnd.n83 240.244
R5808 gnd.n7637 gnd.n84 240.244
R5809 gnd.n7637 gnd.n87 240.244
R5810 gnd.n88 gnd.n87 240.244
R5811 gnd.n89 gnd.n88 240.244
R5812 gnd.n7628 gnd.n89 240.244
R5813 gnd.n7628 gnd.n92 240.244
R5814 gnd.n93 gnd.n92 240.244
R5815 gnd.n94 gnd.n93 240.244
R5816 gnd.n397 gnd.n94 240.244
R5817 gnd.n397 gnd.n97 240.244
R5818 gnd.n98 gnd.n97 240.244
R5819 gnd.n99 gnd.n98 240.244
R5820 gnd.n268 gnd.n99 240.244
R5821 gnd.n268 gnd.n102 240.244
R5822 gnd.n103 gnd.n102 240.244
R5823 gnd.n104 gnd.n103 240.244
R5824 gnd.n243 gnd.n104 240.244
R5825 gnd.n243 gnd.n107 240.244
R5826 gnd.n108 gnd.n107 240.244
R5827 gnd.n109 gnd.n108 240.244
R5828 gnd.n229 gnd.n109 240.244
R5829 gnd.n229 gnd.n112 240.244
R5830 gnd.n113 gnd.n112 240.244
R5831 gnd.n114 gnd.n113 240.244
R5832 gnd.n212 gnd.n114 240.244
R5833 gnd.n212 gnd.n117 240.244
R5834 gnd.n118 gnd.n117 240.244
R5835 gnd.n119 gnd.n118 240.244
R5836 gnd.n7918 gnd.n119 240.244
R5837 gnd.n5933 gnd.n5932 240.244
R5838 gnd.n5927 gnd.n5926 240.244
R5839 gnd.n5945 gnd.n5944 240.244
R5840 gnd.n5957 gnd.n5956 240.244
R5841 gnd.n5915 gnd.n5914 240.244
R5842 gnd.n5969 gnd.n5968 240.244
R5843 gnd.n5981 gnd.n5980 240.244
R5844 gnd.n5903 gnd.n5902 240.244
R5845 gnd.n5898 gnd.n1681 240.244
R5846 gnd.n1483 gnd.n1482 240.244
R5847 gnd.n1484 gnd.n1483 240.244
R5848 gnd.n6073 gnd.n1484 240.244
R5849 gnd.n6073 gnd.n1487 240.244
R5850 gnd.n1488 gnd.n1487 240.244
R5851 gnd.n1489 gnd.n1488 240.244
R5852 gnd.n6093 gnd.n1489 240.244
R5853 gnd.n6093 gnd.n1492 240.244
R5854 gnd.n1493 gnd.n1492 240.244
R5855 gnd.n1494 gnd.n1493 240.244
R5856 gnd.n1621 gnd.n1494 240.244
R5857 gnd.n1621 gnd.n1497 240.244
R5858 gnd.n1498 gnd.n1497 240.244
R5859 gnd.n1499 gnd.n1498 240.244
R5860 gnd.n1603 gnd.n1499 240.244
R5861 gnd.n1603 gnd.n1502 240.244
R5862 gnd.n1503 gnd.n1502 240.244
R5863 gnd.n1504 gnd.n1503 240.244
R5864 gnd.n1577 gnd.n1504 240.244
R5865 gnd.n1577 gnd.n1507 240.244
R5866 gnd.n1508 gnd.n1507 240.244
R5867 gnd.n1509 gnd.n1508 240.244
R5868 gnd.n1548 gnd.n1509 240.244
R5869 gnd.n1548 gnd.n1512 240.244
R5870 gnd.n1513 gnd.n1512 240.244
R5871 gnd.n1514 gnd.n1513 240.244
R5872 gnd.n6306 gnd.n1514 240.244
R5873 gnd.n6306 gnd.n324 240.244
R5874 gnd.n7662 gnd.n324 240.244
R5875 gnd.n7662 gnd.n325 240.244
R5876 gnd.n330 gnd.n325 240.244
R5877 gnd.n331 gnd.n330 240.244
R5878 gnd.n332 gnd.n331 240.244
R5879 gnd.n334 gnd.n332 240.244
R5880 gnd.n7650 gnd.n334 240.244
R5881 gnd.n7650 gnd.n305 240.244
R5882 gnd.n7672 gnd.n305 240.244
R5883 gnd.n7672 gnd.n301 240.244
R5884 gnd.n7678 gnd.n301 240.244
R5885 gnd.n7678 gnd.n290 240.244
R5886 gnd.n7688 gnd.n290 240.244
R5887 gnd.n7688 gnd.n286 240.244
R5888 gnd.n7694 gnd.n286 240.244
R5889 gnd.n7694 gnd.n274 240.244
R5890 gnd.n7704 gnd.n274 240.244
R5891 gnd.n7704 gnd.n270 240.244
R5892 gnd.n7710 gnd.n270 240.244
R5893 gnd.n7710 gnd.n258 240.244
R5894 gnd.n7720 gnd.n258 240.244
R5895 gnd.n7720 gnd.n254 240.244
R5896 gnd.n7726 gnd.n254 240.244
R5897 gnd.n7726 gnd.n242 240.244
R5898 gnd.n7736 gnd.n242 240.244
R5899 gnd.n7736 gnd.n238 240.244
R5900 gnd.n7742 gnd.n238 240.244
R5901 gnd.n7742 gnd.n228 240.244
R5902 gnd.n7752 gnd.n228 240.244
R5903 gnd.n7752 gnd.n224 240.244
R5904 gnd.n7758 gnd.n224 240.244
R5905 gnd.n7758 gnd.n211 240.244
R5906 gnd.n7770 gnd.n211 240.244
R5907 gnd.n7770 gnd.n206 240.244
R5908 gnd.n7837 gnd.n206 240.244
R5909 gnd.n7837 gnd.n129 240.244
R5910 gnd.n2338 gnd.n1252 240.244
R5911 gnd.n2407 gnd.n2406 240.244
R5912 gnd.n2409 gnd.n2408 240.244
R5913 gnd.n2418 gnd.n2417 240.244
R5914 gnd.n2426 gnd.n2425 240.244
R5915 gnd.n2428 gnd.n2427 240.244
R5916 gnd.n2438 gnd.n2437 240.244
R5917 gnd.n2446 gnd.n2445 240.244
R5918 gnd.n2450 gnd.n2447 240.244
R5919 gnd.n4394 gnd.n4150 240.244
R5920 gnd.n4394 gnd.n2668 240.244
R5921 gnd.n4391 gnd.n2668 240.244
R5922 gnd.n4391 gnd.n2661 240.244
R5923 gnd.n4388 gnd.n2661 240.244
R5924 gnd.n4388 gnd.n2653 240.244
R5925 gnd.n4385 gnd.n2653 240.244
R5926 gnd.n4385 gnd.n2644 240.244
R5927 gnd.n4382 gnd.n2644 240.244
R5928 gnd.n4382 gnd.n2636 240.244
R5929 gnd.n4379 gnd.n2636 240.244
R5930 gnd.n4379 gnd.n2628 240.244
R5931 gnd.n4376 gnd.n2628 240.244
R5932 gnd.n4376 gnd.n2619 240.244
R5933 gnd.n4373 gnd.n2619 240.244
R5934 gnd.n4373 gnd.n1021 240.244
R5935 gnd.n4370 gnd.n1021 240.244
R5936 gnd.n4370 gnd.n1034 240.244
R5937 gnd.n4522 gnd.n1034 240.244
R5938 gnd.n4522 gnd.n1046 240.244
R5939 gnd.n4528 gnd.n1046 240.244
R5940 gnd.n4528 gnd.n1056 240.244
R5941 gnd.n4543 gnd.n1056 240.244
R5942 gnd.n4543 gnd.n1067 240.244
R5943 gnd.n4550 gnd.n1067 240.244
R5944 gnd.n4550 gnd.n1077 240.244
R5945 gnd.n4570 gnd.n1077 240.244
R5946 gnd.n4570 gnd.n1088 240.244
R5947 gnd.n2553 gnd.n1088 240.244
R5948 gnd.n4581 gnd.n2553 240.244
R5949 gnd.n4581 gnd.n2554 240.244
R5950 gnd.n2554 gnd.n2550 240.244
R5951 gnd.n2550 gnd.n2532 240.244
R5952 gnd.n4631 gnd.n2532 240.244
R5953 gnd.n4631 gnd.n2528 240.244
R5954 gnd.n4637 gnd.n2528 240.244
R5955 gnd.n4637 gnd.n1103 240.244
R5956 gnd.n4675 gnd.n1103 240.244
R5957 gnd.n4675 gnd.n1114 240.244
R5958 gnd.n2518 gnd.n1114 240.244
R5959 gnd.n2518 gnd.n1124 240.244
R5960 gnd.n2519 gnd.n1124 240.244
R5961 gnd.n2519 gnd.n1135 240.244
R5962 gnd.n4663 gnd.n1135 240.244
R5963 gnd.n4663 gnd.n1146 240.244
R5964 gnd.n4714 gnd.n1146 240.244
R5965 gnd.n4714 gnd.n1156 240.244
R5966 gnd.n4720 gnd.n1156 240.244
R5967 gnd.n4720 gnd.n1167 240.244
R5968 gnd.n4730 gnd.n1167 240.244
R5969 gnd.n4730 gnd.n1178 240.244
R5970 gnd.n4736 gnd.n1178 240.244
R5971 gnd.n4736 gnd.n1189 240.244
R5972 gnd.n4887 gnd.n1189 240.244
R5973 gnd.n4887 gnd.n1199 240.244
R5974 gnd.n2480 gnd.n1199 240.244
R5975 gnd.n2480 gnd.n1210 240.244
R5976 gnd.n2481 gnd.n1210 240.244
R5977 gnd.n2481 gnd.n1221 240.244
R5978 gnd.n2484 gnd.n1221 240.244
R5979 gnd.n2484 gnd.n1232 240.244
R5980 gnd.n4832 gnd.n1232 240.244
R5981 gnd.n4832 gnd.n1243 240.244
R5982 gnd.n4924 gnd.n1243 240.244
R5983 gnd.n4435 gnd.n4433 240.244
R5984 gnd.n4431 gnd.n4329 240.244
R5985 gnd.n4427 gnd.n4425 240.244
R5986 gnd.n4423 gnd.n4335 240.244
R5987 gnd.n4419 gnd.n4417 240.244
R5988 gnd.n4415 gnd.n4341 240.244
R5989 gnd.n4411 gnd.n4409 240.244
R5990 gnd.n4407 gnd.n4347 240.244
R5991 gnd.n4400 gnd.n4399 240.244
R5992 gnd.n4441 gnd.n2666 240.244
R5993 gnd.n4451 gnd.n2666 240.244
R5994 gnd.n4451 gnd.n2662 240.244
R5995 gnd.n4457 gnd.n2662 240.244
R5996 gnd.n4457 gnd.n2650 240.244
R5997 gnd.n4467 gnd.n2650 240.244
R5998 gnd.n4467 gnd.n2646 240.244
R5999 gnd.n4473 gnd.n2646 240.244
R6000 gnd.n4473 gnd.n2634 240.244
R6001 gnd.n4483 gnd.n2634 240.244
R6002 gnd.n4483 gnd.n2629 240.244
R6003 gnd.n4499 gnd.n2629 240.244
R6004 gnd.n4499 gnd.n2630 240.244
R6005 gnd.n2630 gnd.n2620 240.244
R6006 gnd.n4494 gnd.n2620 240.244
R6007 gnd.n4494 gnd.n1023 240.244
R6008 gnd.n1036 gnd.n1023 240.244
R6009 gnd.n6700 gnd.n1036 240.244
R6010 gnd.n6700 gnd.n1037 240.244
R6011 gnd.n6696 gnd.n1037 240.244
R6012 gnd.n6696 gnd.n1043 240.244
R6013 gnd.n6688 gnd.n1043 240.244
R6014 gnd.n6688 gnd.n1058 240.244
R6015 gnd.n6684 gnd.n1058 240.244
R6016 gnd.n6684 gnd.n1064 240.244
R6017 gnd.n6676 gnd.n1064 240.244
R6018 gnd.n6676 gnd.n1079 240.244
R6019 gnd.n6672 gnd.n1079 240.244
R6020 gnd.n6672 gnd.n1085 240.244
R6021 gnd.n4589 gnd.n1085 240.244
R6022 gnd.n4589 gnd.n4583 240.244
R6023 gnd.n4583 gnd.n2541 240.244
R6024 gnd.n4617 gnd.n2541 240.244
R6025 gnd.n4617 gnd.n2535 240.244
R6026 gnd.n4624 gnd.n2535 240.244
R6027 gnd.n4624 gnd.n1105 240.244
R6028 gnd.n6662 gnd.n1105 240.244
R6029 gnd.n6662 gnd.n1106 240.244
R6030 gnd.n6658 gnd.n1106 240.244
R6031 gnd.n6658 gnd.n1112 240.244
R6032 gnd.n6650 gnd.n1112 240.244
R6033 gnd.n6650 gnd.n1126 240.244
R6034 gnd.n6646 gnd.n1126 240.244
R6035 gnd.n6646 gnd.n1132 240.244
R6036 gnd.n6638 gnd.n1132 240.244
R6037 gnd.n6638 gnd.n1148 240.244
R6038 gnd.n6634 gnd.n1148 240.244
R6039 gnd.n6634 gnd.n1154 240.244
R6040 gnd.n6626 gnd.n1154 240.244
R6041 gnd.n6626 gnd.n1169 240.244
R6042 gnd.n6622 gnd.n1169 240.244
R6043 gnd.n6622 gnd.n1175 240.244
R6044 gnd.n6614 gnd.n1175 240.244
R6045 gnd.n6614 gnd.n1191 240.244
R6046 gnd.n6610 gnd.n1191 240.244
R6047 gnd.n6610 gnd.n1197 240.244
R6048 gnd.n6602 gnd.n1197 240.244
R6049 gnd.n6602 gnd.n1212 240.244
R6050 gnd.n6598 gnd.n1212 240.244
R6051 gnd.n6598 gnd.n1218 240.244
R6052 gnd.n6590 gnd.n1218 240.244
R6053 gnd.n6590 gnd.n1234 240.244
R6054 gnd.n6586 gnd.n1234 240.244
R6055 gnd.n6586 gnd.n1240 240.244
R6056 gnd.n6883 gnd.n848 240.244
R6057 gnd.n6883 gnd.n846 240.244
R6058 gnd.n6887 gnd.n846 240.244
R6059 gnd.n6887 gnd.n842 240.244
R6060 gnd.n6893 gnd.n842 240.244
R6061 gnd.n6893 gnd.n840 240.244
R6062 gnd.n6897 gnd.n840 240.244
R6063 gnd.n6897 gnd.n836 240.244
R6064 gnd.n6903 gnd.n836 240.244
R6065 gnd.n6903 gnd.n834 240.244
R6066 gnd.n6907 gnd.n834 240.244
R6067 gnd.n6907 gnd.n830 240.244
R6068 gnd.n6913 gnd.n830 240.244
R6069 gnd.n6913 gnd.n828 240.244
R6070 gnd.n6917 gnd.n828 240.244
R6071 gnd.n6917 gnd.n824 240.244
R6072 gnd.n6923 gnd.n824 240.244
R6073 gnd.n6923 gnd.n822 240.244
R6074 gnd.n6927 gnd.n822 240.244
R6075 gnd.n6927 gnd.n818 240.244
R6076 gnd.n6933 gnd.n818 240.244
R6077 gnd.n6933 gnd.n816 240.244
R6078 gnd.n6937 gnd.n816 240.244
R6079 gnd.n6937 gnd.n812 240.244
R6080 gnd.n6943 gnd.n812 240.244
R6081 gnd.n6943 gnd.n810 240.244
R6082 gnd.n6947 gnd.n810 240.244
R6083 gnd.n6947 gnd.n806 240.244
R6084 gnd.n6953 gnd.n806 240.244
R6085 gnd.n6953 gnd.n804 240.244
R6086 gnd.n6957 gnd.n804 240.244
R6087 gnd.n6957 gnd.n800 240.244
R6088 gnd.n6963 gnd.n800 240.244
R6089 gnd.n6963 gnd.n798 240.244
R6090 gnd.n6967 gnd.n798 240.244
R6091 gnd.n6967 gnd.n794 240.244
R6092 gnd.n6973 gnd.n794 240.244
R6093 gnd.n6973 gnd.n792 240.244
R6094 gnd.n6977 gnd.n792 240.244
R6095 gnd.n6977 gnd.n788 240.244
R6096 gnd.n6983 gnd.n788 240.244
R6097 gnd.n6983 gnd.n786 240.244
R6098 gnd.n6987 gnd.n786 240.244
R6099 gnd.n6987 gnd.n782 240.244
R6100 gnd.n6993 gnd.n782 240.244
R6101 gnd.n6993 gnd.n780 240.244
R6102 gnd.n6997 gnd.n780 240.244
R6103 gnd.n6997 gnd.n776 240.244
R6104 gnd.n7003 gnd.n776 240.244
R6105 gnd.n7003 gnd.n774 240.244
R6106 gnd.n7007 gnd.n774 240.244
R6107 gnd.n7007 gnd.n770 240.244
R6108 gnd.n7013 gnd.n770 240.244
R6109 gnd.n7013 gnd.n768 240.244
R6110 gnd.n7017 gnd.n768 240.244
R6111 gnd.n7017 gnd.n764 240.244
R6112 gnd.n7023 gnd.n764 240.244
R6113 gnd.n7023 gnd.n762 240.244
R6114 gnd.n7027 gnd.n762 240.244
R6115 gnd.n7027 gnd.n758 240.244
R6116 gnd.n7033 gnd.n758 240.244
R6117 gnd.n7033 gnd.n756 240.244
R6118 gnd.n7037 gnd.n756 240.244
R6119 gnd.n7037 gnd.n752 240.244
R6120 gnd.n7043 gnd.n752 240.244
R6121 gnd.n7043 gnd.n750 240.244
R6122 gnd.n7047 gnd.n750 240.244
R6123 gnd.n7047 gnd.n746 240.244
R6124 gnd.n7053 gnd.n746 240.244
R6125 gnd.n7053 gnd.n744 240.244
R6126 gnd.n7057 gnd.n744 240.244
R6127 gnd.n7057 gnd.n740 240.244
R6128 gnd.n7063 gnd.n740 240.244
R6129 gnd.n7063 gnd.n738 240.244
R6130 gnd.n7067 gnd.n738 240.244
R6131 gnd.n7067 gnd.n734 240.244
R6132 gnd.n7073 gnd.n734 240.244
R6133 gnd.n7073 gnd.n732 240.244
R6134 gnd.n7077 gnd.n732 240.244
R6135 gnd.n7077 gnd.n728 240.244
R6136 gnd.n7083 gnd.n728 240.244
R6137 gnd.n7083 gnd.n726 240.244
R6138 gnd.n7087 gnd.n726 240.244
R6139 gnd.n7087 gnd.n722 240.244
R6140 gnd.n7093 gnd.n722 240.244
R6141 gnd.n7093 gnd.n720 240.244
R6142 gnd.n7097 gnd.n720 240.244
R6143 gnd.n7097 gnd.n716 240.244
R6144 gnd.n7103 gnd.n716 240.244
R6145 gnd.n7103 gnd.n714 240.244
R6146 gnd.n7107 gnd.n714 240.244
R6147 gnd.n7107 gnd.n710 240.244
R6148 gnd.n7113 gnd.n710 240.244
R6149 gnd.n7113 gnd.n708 240.244
R6150 gnd.n7117 gnd.n708 240.244
R6151 gnd.n7117 gnd.n704 240.244
R6152 gnd.n7123 gnd.n704 240.244
R6153 gnd.n7123 gnd.n702 240.244
R6154 gnd.n7127 gnd.n702 240.244
R6155 gnd.n7127 gnd.n698 240.244
R6156 gnd.n7133 gnd.n698 240.244
R6157 gnd.n7133 gnd.n696 240.244
R6158 gnd.n7137 gnd.n696 240.244
R6159 gnd.n7137 gnd.n692 240.244
R6160 gnd.n7143 gnd.n692 240.244
R6161 gnd.n7143 gnd.n690 240.244
R6162 gnd.n7147 gnd.n690 240.244
R6163 gnd.n7147 gnd.n686 240.244
R6164 gnd.n7153 gnd.n686 240.244
R6165 gnd.n7153 gnd.n684 240.244
R6166 gnd.n7157 gnd.n684 240.244
R6167 gnd.n7157 gnd.n680 240.244
R6168 gnd.n7163 gnd.n680 240.244
R6169 gnd.n7163 gnd.n678 240.244
R6170 gnd.n7167 gnd.n678 240.244
R6171 gnd.n7167 gnd.n674 240.244
R6172 gnd.n7173 gnd.n674 240.244
R6173 gnd.n7173 gnd.n672 240.244
R6174 gnd.n7177 gnd.n672 240.244
R6175 gnd.n7177 gnd.n668 240.244
R6176 gnd.n7183 gnd.n668 240.244
R6177 gnd.n7183 gnd.n666 240.244
R6178 gnd.n7187 gnd.n666 240.244
R6179 gnd.n7187 gnd.n662 240.244
R6180 gnd.n7193 gnd.n662 240.244
R6181 gnd.n7193 gnd.n660 240.244
R6182 gnd.n7197 gnd.n660 240.244
R6183 gnd.n7197 gnd.n656 240.244
R6184 gnd.n7203 gnd.n656 240.244
R6185 gnd.n7203 gnd.n654 240.244
R6186 gnd.n7207 gnd.n654 240.244
R6187 gnd.n7207 gnd.n650 240.244
R6188 gnd.n7213 gnd.n650 240.244
R6189 gnd.n7213 gnd.n648 240.244
R6190 gnd.n7217 gnd.n648 240.244
R6191 gnd.n7217 gnd.n644 240.244
R6192 gnd.n7223 gnd.n644 240.244
R6193 gnd.n7223 gnd.n642 240.244
R6194 gnd.n7227 gnd.n642 240.244
R6195 gnd.n7227 gnd.n638 240.244
R6196 gnd.n7233 gnd.n638 240.244
R6197 gnd.n7233 gnd.n636 240.244
R6198 gnd.n7237 gnd.n636 240.244
R6199 gnd.n7237 gnd.n632 240.244
R6200 gnd.n7243 gnd.n632 240.244
R6201 gnd.n7243 gnd.n630 240.244
R6202 gnd.n7247 gnd.n630 240.244
R6203 gnd.n7247 gnd.n626 240.244
R6204 gnd.n7253 gnd.n626 240.244
R6205 gnd.n7253 gnd.n624 240.244
R6206 gnd.n7257 gnd.n624 240.244
R6207 gnd.n7257 gnd.n620 240.244
R6208 gnd.n7263 gnd.n620 240.244
R6209 gnd.n7263 gnd.n618 240.244
R6210 gnd.n7267 gnd.n618 240.244
R6211 gnd.n7267 gnd.n614 240.244
R6212 gnd.n7273 gnd.n614 240.244
R6213 gnd.n7273 gnd.n612 240.244
R6214 gnd.n7277 gnd.n612 240.244
R6215 gnd.n7277 gnd.n608 240.244
R6216 gnd.n7283 gnd.n608 240.244
R6217 gnd.n7283 gnd.n606 240.244
R6218 gnd.n7287 gnd.n606 240.244
R6219 gnd.n7287 gnd.n602 240.244
R6220 gnd.n7293 gnd.n602 240.244
R6221 gnd.n7293 gnd.n600 240.244
R6222 gnd.n7297 gnd.n600 240.244
R6223 gnd.n7297 gnd.n596 240.244
R6224 gnd.n7303 gnd.n596 240.244
R6225 gnd.n7303 gnd.n594 240.244
R6226 gnd.n7307 gnd.n594 240.244
R6227 gnd.n7307 gnd.n590 240.244
R6228 gnd.n7313 gnd.n590 240.244
R6229 gnd.n7313 gnd.n588 240.244
R6230 gnd.n7317 gnd.n588 240.244
R6231 gnd.n7317 gnd.n584 240.244
R6232 gnd.n7323 gnd.n584 240.244
R6233 gnd.n7323 gnd.n582 240.244
R6234 gnd.n7327 gnd.n582 240.244
R6235 gnd.n7327 gnd.n578 240.244
R6236 gnd.n7333 gnd.n578 240.244
R6237 gnd.n7333 gnd.n576 240.244
R6238 gnd.n7337 gnd.n576 240.244
R6239 gnd.n7337 gnd.n572 240.244
R6240 gnd.n7343 gnd.n572 240.244
R6241 gnd.n7343 gnd.n570 240.244
R6242 gnd.n7347 gnd.n570 240.244
R6243 gnd.n7347 gnd.n566 240.244
R6244 gnd.n7353 gnd.n566 240.244
R6245 gnd.n7353 gnd.n564 240.244
R6246 gnd.n7357 gnd.n564 240.244
R6247 gnd.n7357 gnd.n560 240.244
R6248 gnd.n7363 gnd.n560 240.244
R6249 gnd.n7363 gnd.n558 240.244
R6250 gnd.n7367 gnd.n558 240.244
R6251 gnd.n7367 gnd.n554 240.244
R6252 gnd.n7373 gnd.n554 240.244
R6253 gnd.n7373 gnd.n552 240.244
R6254 gnd.n7377 gnd.n552 240.244
R6255 gnd.n7377 gnd.n548 240.244
R6256 gnd.n7383 gnd.n548 240.244
R6257 gnd.n7383 gnd.n546 240.244
R6258 gnd.n7387 gnd.n546 240.244
R6259 gnd.n7387 gnd.n542 240.244
R6260 gnd.n7393 gnd.n542 240.244
R6261 gnd.n7393 gnd.n540 240.244
R6262 gnd.n7397 gnd.n540 240.244
R6263 gnd.n7403 gnd.n536 240.244
R6264 gnd.n7403 gnd.n534 240.244
R6265 gnd.n7407 gnd.n534 240.244
R6266 gnd.n7407 gnd.n530 240.244
R6267 gnd.n7413 gnd.n530 240.244
R6268 gnd.n7413 gnd.n528 240.244
R6269 gnd.n7417 gnd.n528 240.244
R6270 gnd.n7417 gnd.n524 240.244
R6271 gnd.n7423 gnd.n524 240.244
R6272 gnd.n7423 gnd.n522 240.244
R6273 gnd.n7427 gnd.n522 240.244
R6274 gnd.n7427 gnd.n518 240.244
R6275 gnd.n7433 gnd.n518 240.244
R6276 gnd.n7433 gnd.n516 240.244
R6277 gnd.n7437 gnd.n516 240.244
R6278 gnd.n7437 gnd.n512 240.244
R6279 gnd.n7443 gnd.n512 240.244
R6280 gnd.n7443 gnd.n510 240.244
R6281 gnd.n7447 gnd.n510 240.244
R6282 gnd.n7447 gnd.n506 240.244
R6283 gnd.n7453 gnd.n506 240.244
R6284 gnd.n7453 gnd.n504 240.244
R6285 gnd.n7457 gnd.n504 240.244
R6286 gnd.n7457 gnd.n500 240.244
R6287 gnd.n7463 gnd.n500 240.244
R6288 gnd.n7463 gnd.n498 240.244
R6289 gnd.n7467 gnd.n498 240.244
R6290 gnd.n7467 gnd.n494 240.244
R6291 gnd.n7473 gnd.n494 240.244
R6292 gnd.n7473 gnd.n492 240.244
R6293 gnd.n7477 gnd.n492 240.244
R6294 gnd.n7477 gnd.n488 240.244
R6295 gnd.n7483 gnd.n488 240.244
R6296 gnd.n7483 gnd.n486 240.244
R6297 gnd.n7487 gnd.n486 240.244
R6298 gnd.n7487 gnd.n482 240.244
R6299 gnd.n7493 gnd.n482 240.244
R6300 gnd.n7493 gnd.n480 240.244
R6301 gnd.n7497 gnd.n480 240.244
R6302 gnd.n7497 gnd.n476 240.244
R6303 gnd.n7503 gnd.n476 240.244
R6304 gnd.n7503 gnd.n474 240.244
R6305 gnd.n7507 gnd.n474 240.244
R6306 gnd.n7507 gnd.n470 240.244
R6307 gnd.n7513 gnd.n470 240.244
R6308 gnd.n7513 gnd.n468 240.244
R6309 gnd.n7517 gnd.n468 240.244
R6310 gnd.n7517 gnd.n464 240.244
R6311 gnd.n7523 gnd.n464 240.244
R6312 gnd.n7523 gnd.n462 240.244
R6313 gnd.n7527 gnd.n462 240.244
R6314 gnd.n7527 gnd.n458 240.244
R6315 gnd.n7533 gnd.n458 240.244
R6316 gnd.n7533 gnd.n456 240.244
R6317 gnd.n7537 gnd.n456 240.244
R6318 gnd.n7537 gnd.n452 240.244
R6319 gnd.n7543 gnd.n452 240.244
R6320 gnd.n7543 gnd.n450 240.244
R6321 gnd.n7547 gnd.n450 240.244
R6322 gnd.n7547 gnd.n446 240.244
R6323 gnd.n7553 gnd.n446 240.244
R6324 gnd.n7553 gnd.n444 240.244
R6325 gnd.n7557 gnd.n444 240.244
R6326 gnd.n7557 gnd.n440 240.244
R6327 gnd.n7563 gnd.n440 240.244
R6328 gnd.n7563 gnd.n438 240.244
R6329 gnd.n7567 gnd.n438 240.244
R6330 gnd.n7567 gnd.n434 240.244
R6331 gnd.n7573 gnd.n434 240.244
R6332 gnd.n7573 gnd.n432 240.244
R6333 gnd.n7577 gnd.n432 240.244
R6334 gnd.n7577 gnd.n428 240.244
R6335 gnd.n7583 gnd.n428 240.244
R6336 gnd.n7583 gnd.n426 240.244
R6337 gnd.n7587 gnd.n426 240.244
R6338 gnd.n7587 gnd.n422 240.244
R6339 gnd.n7593 gnd.n422 240.244
R6340 gnd.n7593 gnd.n420 240.244
R6341 gnd.n7597 gnd.n420 240.244
R6342 gnd.n7597 gnd.n416 240.244
R6343 gnd.n7605 gnd.n416 240.244
R6344 gnd.n7605 gnd.n414 240.244
R6345 gnd.n7609 gnd.n414 240.244
R6346 gnd.n7610 gnd.n7609 240.244
R6347 gnd.n2591 gnd.n1018 240.244
R6348 gnd.n2591 gnd.n2586 240.244
R6349 gnd.n2608 gnd.n2586 240.244
R6350 gnd.n2608 gnd.n2587 240.244
R6351 gnd.n2604 gnd.n2587 240.244
R6352 gnd.n2604 gnd.n2603 240.244
R6353 gnd.n2603 gnd.n2578 240.244
R6354 gnd.n4553 gnd.n2578 240.244
R6355 gnd.n4554 gnd.n4553 240.244
R6356 gnd.n4554 gnd.n2574 240.244
R6357 gnd.n4561 gnd.n2574 240.244
R6358 gnd.n4561 gnd.n2575 240.244
R6359 gnd.n2575 gnd.n2547 240.244
R6360 gnd.n4599 gnd.n2547 240.244
R6361 gnd.n4599 gnd.n2544 240.244
R6362 gnd.n4614 gnd.n2544 240.244
R6363 gnd.n4614 gnd.n2545 240.244
R6364 gnd.n4609 gnd.n2545 240.244
R6365 gnd.n4609 gnd.n4608 240.244
R6366 gnd.n4608 gnd.n2511 240.244
R6367 gnd.n4678 gnd.n2511 240.244
R6368 gnd.n4679 gnd.n4678 240.244
R6369 gnd.n4680 gnd.n4679 240.244
R6370 gnd.n4680 gnd.n2507 240.244
R6371 gnd.n4686 gnd.n2507 240.244
R6372 gnd.n4687 gnd.n4686 240.244
R6373 gnd.n4688 gnd.n4687 240.244
R6374 gnd.n4688 gnd.n2502 240.244
R6375 gnd.n4711 gnd.n2502 240.244
R6376 gnd.n4711 gnd.n2503 240.244
R6377 gnd.n4707 gnd.n2503 240.244
R6378 gnd.n4707 gnd.n4706 240.244
R6379 gnd.n4706 gnd.n4705 240.244
R6380 gnd.n4705 gnd.n4696 240.244
R6381 gnd.n4701 gnd.n4696 240.244
R6382 gnd.n4701 gnd.n2474 240.244
R6383 gnd.n4890 gnd.n2474 240.244
R6384 gnd.n4890 gnd.n2470 240.244
R6385 gnd.n4896 gnd.n2470 240.244
R6386 gnd.n4897 gnd.n4896 240.244
R6387 gnd.n4898 gnd.n4897 240.244
R6388 gnd.n4898 gnd.n2466 240.244
R6389 gnd.n4904 gnd.n2466 240.244
R6390 gnd.n4905 gnd.n4904 240.244
R6391 gnd.n4906 gnd.n4905 240.244
R6392 gnd.n4906 gnd.n2461 240.244
R6393 gnd.n4921 gnd.n2461 240.244
R6394 gnd.n4921 gnd.n2462 240.244
R6395 gnd.n4917 gnd.n2462 240.244
R6396 gnd.n4917 gnd.n4916 240.244
R6397 gnd.n4916 gnd.n2315 240.244
R6398 gnd.n4975 gnd.n2315 240.244
R6399 gnd.n4975 gnd.n2311 240.244
R6400 gnd.n4981 gnd.n2311 240.244
R6401 gnd.n4981 gnd.n2301 240.244
R6402 gnd.n4991 gnd.n2301 240.244
R6403 gnd.n4991 gnd.n2297 240.244
R6404 gnd.n4997 gnd.n2297 240.244
R6405 gnd.n4997 gnd.n2287 240.244
R6406 gnd.n5007 gnd.n2287 240.244
R6407 gnd.n5007 gnd.n2283 240.244
R6408 gnd.n5013 gnd.n2283 240.244
R6409 gnd.n5013 gnd.n2273 240.244
R6410 gnd.n5023 gnd.n2273 240.244
R6411 gnd.n5023 gnd.n2269 240.244
R6412 gnd.n5029 gnd.n2269 240.244
R6413 gnd.n5029 gnd.n2259 240.244
R6414 gnd.n5039 gnd.n2259 240.244
R6415 gnd.n5039 gnd.n2255 240.244
R6416 gnd.n5045 gnd.n2255 240.244
R6417 gnd.n5045 gnd.n2244 240.244
R6418 gnd.n5055 gnd.n2244 240.244
R6419 gnd.n5055 gnd.n2240 240.244
R6420 gnd.n5061 gnd.n2240 240.244
R6421 gnd.n5061 gnd.n2229 240.244
R6422 gnd.n5082 gnd.n2229 240.244
R6423 gnd.n5082 gnd.n2224 240.244
R6424 gnd.n5091 gnd.n2224 240.244
R6425 gnd.n5091 gnd.n2225 240.244
R6426 gnd.n2225 gnd.n1368 240.244
R6427 gnd.n6471 gnd.n1368 240.244
R6428 gnd.n6471 gnd.n1369 240.244
R6429 gnd.n6467 gnd.n1369 240.244
R6430 gnd.n6467 gnd.n1375 240.244
R6431 gnd.n5244 gnd.n1375 240.244
R6432 gnd.n5244 gnd.n2200 240.244
R6433 gnd.n5265 gnd.n2200 240.244
R6434 gnd.n5265 gnd.n2196 240.244
R6435 gnd.n5271 gnd.n2196 240.244
R6436 gnd.n5271 gnd.n2181 240.244
R6437 gnd.n5289 gnd.n2181 240.244
R6438 gnd.n5289 gnd.n2177 240.244
R6439 gnd.n5295 gnd.n2177 240.244
R6440 gnd.n5295 gnd.n2159 240.244
R6441 gnd.n5315 gnd.n2159 240.244
R6442 gnd.n5315 gnd.n2154 240.244
R6443 gnd.n5323 gnd.n2154 240.244
R6444 gnd.n5323 gnd.n2155 240.244
R6445 gnd.n2155 gnd.n2130 240.244
R6446 gnd.n5370 gnd.n2130 240.244
R6447 gnd.n5370 gnd.n2124 240.244
R6448 gnd.n5378 gnd.n2124 240.244
R6449 gnd.n5378 gnd.n2126 240.244
R6450 gnd.n2126 gnd.n2107 240.244
R6451 gnd.n5411 gnd.n2107 240.244
R6452 gnd.n5411 gnd.n2102 240.244
R6453 gnd.n5419 gnd.n2102 240.244
R6454 gnd.n5419 gnd.n2103 240.244
R6455 gnd.n2103 gnd.n2078 240.244
R6456 gnd.n5452 gnd.n2078 240.244
R6457 gnd.n5452 gnd.n2074 240.244
R6458 gnd.n5459 gnd.n2074 240.244
R6459 gnd.n5459 gnd.n2051 240.244
R6460 gnd.n5506 gnd.n2051 240.244
R6461 gnd.n5506 gnd.n2052 240.244
R6462 gnd.n5502 gnd.n2052 240.244
R6463 gnd.n5502 gnd.n5501 240.244
R6464 gnd.n5501 gnd.n5500 240.244
R6465 gnd.n5500 gnd.n2020 240.244
R6466 gnd.n5552 gnd.n2020 240.244
R6467 gnd.n5552 gnd.n2016 240.244
R6468 gnd.n5558 gnd.n2016 240.244
R6469 gnd.n5558 gnd.n2004 240.244
R6470 gnd.n5583 gnd.n2004 240.244
R6471 gnd.n5583 gnd.n2000 240.244
R6472 gnd.n5589 gnd.n2000 240.244
R6473 gnd.n5589 gnd.n1798 240.244
R6474 gnd.n5758 gnd.n1798 240.244
R6475 gnd.n5758 gnd.n1794 240.244
R6476 gnd.n5764 gnd.n1794 240.244
R6477 gnd.n5764 gnd.n1786 240.244
R6478 gnd.n5776 gnd.n1786 240.244
R6479 gnd.n5776 gnd.n1782 240.244
R6480 gnd.n5782 gnd.n1782 240.244
R6481 gnd.n5782 gnd.n1775 240.244
R6482 gnd.n5793 gnd.n1775 240.244
R6483 gnd.n5793 gnd.n1771 240.244
R6484 gnd.n5799 gnd.n1771 240.244
R6485 gnd.n5799 gnd.n1763 240.244
R6486 gnd.n5810 gnd.n1763 240.244
R6487 gnd.n5810 gnd.n1759 240.244
R6488 gnd.n5816 gnd.n1759 240.244
R6489 gnd.n5816 gnd.n1751 240.244
R6490 gnd.n5827 gnd.n1751 240.244
R6491 gnd.n5827 gnd.n1747 240.244
R6492 gnd.n5833 gnd.n1747 240.244
R6493 gnd.n5833 gnd.n1739 240.244
R6494 gnd.n5844 gnd.n1739 240.244
R6495 gnd.n5844 gnd.n1735 240.244
R6496 gnd.n5852 gnd.n1735 240.244
R6497 gnd.n5852 gnd.n1727 240.244
R6498 gnd.n5863 gnd.n1727 240.244
R6499 gnd.n5864 gnd.n5863 240.244
R6500 gnd.n5864 gnd.n1473 240.244
R6501 gnd.n5870 gnd.n1473 240.244
R6502 gnd.n5871 gnd.n5870 240.244
R6503 gnd.n6031 gnd.n5871 240.244
R6504 gnd.n6031 gnd.n1719 240.244
R6505 gnd.n6039 gnd.n1719 240.244
R6506 gnd.n6039 gnd.n1720 240.244
R6507 gnd.n1720 gnd.n1674 240.244
R6508 gnd.n6063 gnd.n1674 240.244
R6509 gnd.n6063 gnd.n1669 240.244
R6510 gnd.n6071 gnd.n1669 240.244
R6511 gnd.n6071 gnd.n1670 240.244
R6512 gnd.n1670 gnd.n1648 240.244
R6513 gnd.n6096 gnd.n1648 240.244
R6514 gnd.n6096 gnd.n1643 240.244
R6515 gnd.n6104 gnd.n1643 240.244
R6516 gnd.n6104 gnd.n1644 240.244
R6517 gnd.n1644 gnd.n1620 240.244
R6518 gnd.n6127 gnd.n1620 240.244
R6519 gnd.n6127 gnd.n1615 240.244
R6520 gnd.n6142 gnd.n1615 240.244
R6521 gnd.n6142 gnd.n1616 240.244
R6522 gnd.n6138 gnd.n1616 240.244
R6523 gnd.n6138 gnd.n6137 240.244
R6524 gnd.n6137 gnd.n1579 240.244
R6525 gnd.n6210 gnd.n1579 240.244
R6526 gnd.n6210 gnd.n1580 240.244
R6527 gnd.n6206 gnd.n1580 240.244
R6528 gnd.n6206 gnd.n1587 240.244
R6529 gnd.n1587 gnd.n1547 240.244
R6530 gnd.n6244 gnd.n1547 240.244
R6531 gnd.n6244 gnd.n1543 240.244
R6532 gnd.n6251 gnd.n1543 240.244
R6533 gnd.n6252 gnd.n6251 240.244
R6534 gnd.n6253 gnd.n6252 240.244
R6535 gnd.n6253 gnd.n1541 240.244
R6536 gnd.n6258 gnd.n1541 240.244
R6537 gnd.n6259 gnd.n6258 240.244
R6538 gnd.n6259 gnd.n1538 240.244
R6539 gnd.n6283 gnd.n1538 240.244
R6540 gnd.n6283 gnd.n1539 240.244
R6541 gnd.n6278 gnd.n1539 240.244
R6542 gnd.n6278 gnd.n6277 240.244
R6543 gnd.n6277 gnd.n6276 240.244
R6544 gnd.n6276 gnd.n6264 240.244
R6545 gnd.n6272 gnd.n6264 240.244
R6546 gnd.n6272 gnd.n6271 240.244
R6547 gnd.n6271 gnd.n402 240.244
R6548 gnd.n7622 gnd.n402 240.244
R6549 gnd.n7622 gnd.n403 240.244
R6550 gnd.n7618 gnd.n403 240.244
R6551 gnd.n7618 gnd.n7617 240.244
R6552 gnd.n7617 gnd.n7616 240.244
R6553 gnd.n7616 gnd.n409 240.244
R6554 gnd.n6877 gnd.n852 240.244
R6555 gnd.n6873 gnd.n852 240.244
R6556 gnd.n6873 gnd.n854 240.244
R6557 gnd.n6869 gnd.n854 240.244
R6558 gnd.n6869 gnd.n859 240.244
R6559 gnd.n6865 gnd.n859 240.244
R6560 gnd.n6865 gnd.n861 240.244
R6561 gnd.n6861 gnd.n861 240.244
R6562 gnd.n6861 gnd.n867 240.244
R6563 gnd.n6857 gnd.n867 240.244
R6564 gnd.n6857 gnd.n869 240.244
R6565 gnd.n6853 gnd.n869 240.244
R6566 gnd.n6853 gnd.n875 240.244
R6567 gnd.n6849 gnd.n875 240.244
R6568 gnd.n6849 gnd.n877 240.244
R6569 gnd.n6845 gnd.n877 240.244
R6570 gnd.n6845 gnd.n883 240.244
R6571 gnd.n6841 gnd.n883 240.244
R6572 gnd.n6841 gnd.n885 240.244
R6573 gnd.n6837 gnd.n885 240.244
R6574 gnd.n6837 gnd.n891 240.244
R6575 gnd.n6833 gnd.n891 240.244
R6576 gnd.n6833 gnd.n893 240.244
R6577 gnd.n6829 gnd.n893 240.244
R6578 gnd.n6829 gnd.n899 240.244
R6579 gnd.n6825 gnd.n899 240.244
R6580 gnd.n6825 gnd.n901 240.244
R6581 gnd.n6821 gnd.n901 240.244
R6582 gnd.n6821 gnd.n907 240.244
R6583 gnd.n6817 gnd.n907 240.244
R6584 gnd.n6817 gnd.n909 240.244
R6585 gnd.n6813 gnd.n909 240.244
R6586 gnd.n6813 gnd.n915 240.244
R6587 gnd.n6809 gnd.n915 240.244
R6588 gnd.n6809 gnd.n917 240.244
R6589 gnd.n6805 gnd.n917 240.244
R6590 gnd.n6805 gnd.n923 240.244
R6591 gnd.n6801 gnd.n923 240.244
R6592 gnd.n6801 gnd.n925 240.244
R6593 gnd.n6797 gnd.n925 240.244
R6594 gnd.n6797 gnd.n931 240.244
R6595 gnd.n6793 gnd.n931 240.244
R6596 gnd.n6793 gnd.n933 240.244
R6597 gnd.n6789 gnd.n933 240.244
R6598 gnd.n6789 gnd.n939 240.244
R6599 gnd.n6785 gnd.n939 240.244
R6600 gnd.n6785 gnd.n941 240.244
R6601 gnd.n6781 gnd.n941 240.244
R6602 gnd.n6781 gnd.n947 240.244
R6603 gnd.n6777 gnd.n947 240.244
R6604 gnd.n6777 gnd.n949 240.244
R6605 gnd.n6773 gnd.n949 240.244
R6606 gnd.n6773 gnd.n955 240.244
R6607 gnd.n6769 gnd.n955 240.244
R6608 gnd.n6769 gnd.n957 240.244
R6609 gnd.n6765 gnd.n957 240.244
R6610 gnd.n6765 gnd.n963 240.244
R6611 gnd.n6761 gnd.n963 240.244
R6612 gnd.n6761 gnd.n965 240.244
R6613 gnd.n6757 gnd.n965 240.244
R6614 gnd.n6757 gnd.n971 240.244
R6615 gnd.n6753 gnd.n971 240.244
R6616 gnd.n6753 gnd.n973 240.244
R6617 gnd.n6749 gnd.n973 240.244
R6618 gnd.n6749 gnd.n979 240.244
R6619 gnd.n6745 gnd.n979 240.244
R6620 gnd.n6745 gnd.n981 240.244
R6621 gnd.n6741 gnd.n981 240.244
R6622 gnd.n6741 gnd.n987 240.244
R6623 gnd.n6737 gnd.n987 240.244
R6624 gnd.n6737 gnd.n989 240.244
R6625 gnd.n6733 gnd.n989 240.244
R6626 gnd.n6733 gnd.n995 240.244
R6627 gnd.n6729 gnd.n995 240.244
R6628 gnd.n6729 gnd.n997 240.244
R6629 gnd.n6725 gnd.n997 240.244
R6630 gnd.n6725 gnd.n1003 240.244
R6631 gnd.n6721 gnd.n1003 240.244
R6632 gnd.n6721 gnd.n1005 240.244
R6633 gnd.n6717 gnd.n1005 240.244
R6634 gnd.n6717 gnd.n1011 240.244
R6635 gnd.n6713 gnd.n1011 240.244
R6636 gnd.n6713 gnd.n1013 240.244
R6637 gnd.n6709 gnd.n1013 240.244
R6638 gnd.n2332 gnd.n2310 240.244
R6639 gnd.n2342 gnd.n2310 240.244
R6640 gnd.n2342 gnd.n2303 240.244
R6641 gnd.n2345 gnd.n2303 240.244
R6642 gnd.n2345 gnd.n2295 240.244
R6643 gnd.n2346 gnd.n2295 240.244
R6644 gnd.n2346 gnd.n2288 240.244
R6645 gnd.n2349 gnd.n2288 240.244
R6646 gnd.n2349 gnd.n2282 240.244
R6647 gnd.n2350 gnd.n2282 240.244
R6648 gnd.n2350 gnd.n2275 240.244
R6649 gnd.n2353 gnd.n2275 240.244
R6650 gnd.n2353 gnd.n2268 240.244
R6651 gnd.n2354 gnd.n2268 240.244
R6652 gnd.n2354 gnd.n2261 240.244
R6653 gnd.n2357 gnd.n2261 240.244
R6654 gnd.n2357 gnd.n2254 240.244
R6655 gnd.n2358 gnd.n2254 240.244
R6656 gnd.n2358 gnd.n2246 240.244
R6657 gnd.n2361 gnd.n2246 240.244
R6658 gnd.n2361 gnd.n2239 240.244
R6659 gnd.n2362 gnd.n2239 240.244
R6660 gnd.n2362 gnd.n2231 240.244
R6661 gnd.n2231 gnd.n2221 240.244
R6662 gnd.n5093 gnd.n2221 240.244
R6663 gnd.n5095 gnd.n5093 240.244
R6664 gnd.n5095 gnd.n5094 240.244
R6665 gnd.n5094 gnd.n1365 240.244
R6666 gnd.n5197 gnd.n1365 240.244
R6667 gnd.n5197 gnd.n1377 240.244
R6668 gnd.n2213 gnd.n1377 240.244
R6669 gnd.n5240 gnd.n2213 240.244
R6670 gnd.n5240 gnd.n2214 240.244
R6671 gnd.n2214 gnd.n2201 240.244
R6672 gnd.n5203 gnd.n2201 240.244
R6673 gnd.n5203 gnd.n2194 240.244
R6674 gnd.n5204 gnd.n2194 240.244
R6675 gnd.n5204 gnd.n2183 240.244
R6676 gnd.n5207 gnd.n2183 240.244
R6677 gnd.n5207 gnd.n2176 240.244
R6678 gnd.n5208 gnd.n2176 240.244
R6679 gnd.n5208 gnd.n2162 240.244
R6680 gnd.n5211 gnd.n2162 240.244
R6681 gnd.n5211 gnd.n2152 240.244
R6682 gnd.n5214 gnd.n2152 240.244
R6683 gnd.n5215 gnd.n5214 240.244
R6684 gnd.n5215 gnd.n2132 240.244
R6685 gnd.n2132 gnd.n2121 240.244
R6686 gnd.n5380 gnd.n2121 240.244
R6687 gnd.n5380 gnd.n2116 240.244
R6688 gnd.n5400 gnd.n2116 240.244
R6689 gnd.n5400 gnd.n2109 240.244
R6690 gnd.n5385 gnd.n2109 240.244
R6691 gnd.n5385 gnd.n2100 240.244
R6692 gnd.n5386 gnd.n2100 240.244
R6693 gnd.n5387 gnd.n5386 240.244
R6694 gnd.n5387 gnd.n2080 240.244
R6695 gnd.n2080 gnd.n2068 240.244
R6696 gnd.n5461 gnd.n2068 240.244
R6697 gnd.n5461 gnd.n2069 240.244
R6698 gnd.n2069 gnd.n2050 240.244
R6699 gnd.n5468 gnd.n2050 240.244
R6700 gnd.n5469 gnd.n5468 240.244
R6701 gnd.n5469 gnd.n2061 240.244
R6702 gnd.n5498 gnd.n2061 240.244
R6703 gnd.n5498 gnd.n2030 240.244
R6704 gnd.n2030 gnd.n2021 240.244
R6705 gnd.n5475 gnd.n2021 240.244
R6706 gnd.n5475 gnd.n2015 240.244
R6707 gnd.n2015 gnd.n2011 240.244
R6708 gnd.n2011 gnd.n2005 240.244
R6709 gnd.n5478 gnd.n2005 240.244
R6710 gnd.n5478 gnd.n1999 240.244
R6711 gnd.n5479 gnd.n1999 240.244
R6712 gnd.n5479 gnd.n1800 240.244
R6713 gnd.n1800 gnd.n1792 240.244
R6714 gnd.n5766 gnd.n1792 240.244
R6715 gnd.n5766 gnd.n1788 240.244
R6716 gnd.n5772 gnd.n1788 240.244
R6717 gnd.n5772 gnd.n1781 240.244
R6718 gnd.n5784 gnd.n1781 240.244
R6719 gnd.n5784 gnd.n1777 240.244
R6720 gnd.n5790 gnd.n1777 240.244
R6721 gnd.n5790 gnd.n1769 240.244
R6722 gnd.n5801 gnd.n1769 240.244
R6723 gnd.n5801 gnd.n1765 240.244
R6724 gnd.n5807 gnd.n1765 240.244
R6725 gnd.n5807 gnd.n1757 240.244
R6726 gnd.n5818 gnd.n1757 240.244
R6727 gnd.n5818 gnd.n1753 240.244
R6728 gnd.n5824 gnd.n1753 240.244
R6729 gnd.n5824 gnd.n1744 240.244
R6730 gnd.n5835 gnd.n1744 240.244
R6731 gnd.n5835 gnd.n1740 240.244
R6732 gnd.n5841 gnd.n1740 240.244
R6733 gnd.n5841 gnd.n1733 240.244
R6734 gnd.n5854 gnd.n1733 240.244
R6735 gnd.n5854 gnd.n1729 240.244
R6736 gnd.n5860 gnd.n1729 240.244
R6737 gnd.n5860 gnd.n1475 240.244
R6738 gnd.n6354 gnd.n1475 240.244
R6739 gnd.n2331 gnd.n2330 240.244
R6740 gnd.n2412 gnd.n2330 240.244
R6741 gnd.n2414 gnd.n2413 240.244
R6742 gnd.n2422 gnd.n2421 240.244
R6743 gnd.n2432 gnd.n2431 240.244
R6744 gnd.n2434 gnd.n2433 240.244
R6745 gnd.n2442 gnd.n2441 240.244
R6746 gnd.n2454 gnd.n2453 240.244
R6747 gnd.n2456 gnd.n2455 240.244
R6748 gnd.n4836 gnd.n4835 240.244
R6749 gnd.n4838 gnd.n4837 240.244
R6750 gnd.n4842 gnd.n4841 240.244
R6751 gnd.n4848 gnd.n4843 240.244
R6752 gnd.n4850 gnd.n4849 240.244
R6753 gnd.n4983 gnd.n2308 240.244
R6754 gnd.n4983 gnd.n2304 240.244
R6755 gnd.n4989 gnd.n2304 240.244
R6756 gnd.n4989 gnd.n2293 240.244
R6757 gnd.n4999 gnd.n2293 240.244
R6758 gnd.n4999 gnd.n2289 240.244
R6759 gnd.n5005 gnd.n2289 240.244
R6760 gnd.n5005 gnd.n2280 240.244
R6761 gnd.n5015 gnd.n2280 240.244
R6762 gnd.n5015 gnd.n2276 240.244
R6763 gnd.n5021 gnd.n2276 240.244
R6764 gnd.n5021 gnd.n2266 240.244
R6765 gnd.n5031 gnd.n2266 240.244
R6766 gnd.n5031 gnd.n2262 240.244
R6767 gnd.n5037 gnd.n2262 240.244
R6768 gnd.n5037 gnd.n2252 240.244
R6769 gnd.n5047 gnd.n2252 240.244
R6770 gnd.n5047 gnd.n2248 240.244
R6771 gnd.n5053 gnd.n2248 240.244
R6772 gnd.n5053 gnd.n2238 240.244
R6773 gnd.n5063 gnd.n2238 240.244
R6774 gnd.n5063 gnd.n2232 240.244
R6775 gnd.n5080 gnd.n2232 240.244
R6776 gnd.n5080 gnd.n2233 240.244
R6777 gnd.n2233 gnd.n2223 240.244
R6778 gnd.n5068 gnd.n2223 240.244
R6779 gnd.n5069 gnd.n5068 240.244
R6780 gnd.n5069 gnd.n1367 240.244
R6781 gnd.n1379 gnd.n1367 240.244
R6782 gnd.n6465 gnd.n1379 240.244
R6783 gnd.n6465 gnd.n1380 240.244
R6784 gnd.n1385 gnd.n1380 240.244
R6785 gnd.n1386 gnd.n1385 240.244
R6786 gnd.n1387 gnd.n1386 240.244
R6787 gnd.n2203 gnd.n1387 240.244
R6788 gnd.n2203 gnd.n1390 240.244
R6789 gnd.n1391 gnd.n1390 240.244
R6790 gnd.n1392 gnd.n1391 240.244
R6791 gnd.n2173 gnd.n1392 240.244
R6792 gnd.n2173 gnd.n1395 240.244
R6793 gnd.n1396 gnd.n1395 240.244
R6794 gnd.n1397 gnd.n1396 240.244
R6795 gnd.n2149 gnd.n1397 240.244
R6796 gnd.n2149 gnd.n1400 240.244
R6797 gnd.n1401 gnd.n1400 240.244
R6798 gnd.n1402 gnd.n1401 240.244
R6799 gnd.n5368 gnd.n1402 240.244
R6800 gnd.n5368 gnd.n1405 240.244
R6801 gnd.n1406 gnd.n1405 240.244
R6802 gnd.n1407 gnd.n1406 240.244
R6803 gnd.n5401 gnd.n1407 240.244
R6804 gnd.n5401 gnd.n1410 240.244
R6805 gnd.n1411 gnd.n1410 240.244
R6806 gnd.n1412 gnd.n1411 240.244
R6807 gnd.n2093 gnd.n1412 240.244
R6808 gnd.n2093 gnd.n1415 240.244
R6809 gnd.n1416 gnd.n1415 240.244
R6810 gnd.n1417 gnd.n1416 240.244
R6811 gnd.n2072 gnd.n1417 240.244
R6812 gnd.n2072 gnd.n1420 240.244
R6813 gnd.n1421 gnd.n1420 240.244
R6814 gnd.n1422 gnd.n1421 240.244
R6815 gnd.n2037 gnd.n1422 240.244
R6816 gnd.n2037 gnd.n1425 240.244
R6817 gnd.n1426 gnd.n1425 240.244
R6818 gnd.n1427 gnd.n1426 240.244
R6819 gnd.n5550 gnd.n1427 240.244
R6820 gnd.n5550 gnd.n1430 240.244
R6821 gnd.n1431 gnd.n1430 240.244
R6822 gnd.n1432 gnd.n1431 240.244
R6823 gnd.n5581 gnd.n1432 240.244
R6824 gnd.n5581 gnd.n1435 240.244
R6825 gnd.n1436 gnd.n1435 240.244
R6826 gnd.n1437 gnd.n1436 240.244
R6827 gnd.n5756 gnd.n1437 240.244
R6828 gnd.n5756 gnd.n1440 240.244
R6829 gnd.n1441 gnd.n1440 240.244
R6830 gnd.n1442 gnd.n1441 240.244
R6831 gnd.n5774 gnd.n1442 240.244
R6832 gnd.n5774 gnd.n1445 240.244
R6833 gnd.n1446 gnd.n1445 240.244
R6834 gnd.n1447 gnd.n1446 240.244
R6835 gnd.n5791 gnd.n1447 240.244
R6836 gnd.n5791 gnd.n1450 240.244
R6837 gnd.n1451 gnd.n1450 240.244
R6838 gnd.n1452 gnd.n1451 240.244
R6839 gnd.n5808 gnd.n1452 240.244
R6840 gnd.n5808 gnd.n1455 240.244
R6841 gnd.n1456 gnd.n1455 240.244
R6842 gnd.n1457 gnd.n1456 240.244
R6843 gnd.n5825 gnd.n1457 240.244
R6844 gnd.n5825 gnd.n1460 240.244
R6845 gnd.n1461 gnd.n1460 240.244
R6846 gnd.n1462 gnd.n1461 240.244
R6847 gnd.n5842 gnd.n1462 240.244
R6848 gnd.n5842 gnd.n1465 240.244
R6849 gnd.n1466 gnd.n1465 240.244
R6850 gnd.n1467 gnd.n1466 240.244
R6851 gnd.n5861 gnd.n1467 240.244
R6852 gnd.n5861 gnd.n1470 240.244
R6853 gnd.n6356 gnd.n1470 240.244
R6854 gnd.n5939 gnd.n5938 240.244
R6855 gnd.n5923 gnd.n5922 240.244
R6856 gnd.n5951 gnd.n5950 240.244
R6857 gnd.n5963 gnd.n5962 240.244
R6858 gnd.n5911 gnd.n5910 240.244
R6859 gnd.n5975 gnd.n5974 240.244
R6860 gnd.n5988 gnd.n5987 240.244
R6861 gnd.n5991 gnd.n5990 240.244
R6862 gnd.n5895 gnd.n5894 240.244
R6863 gnd.n6006 gnd.n6005 240.244
R6864 gnd.n6009 gnd.n6008 240.244
R6865 gnd.n6016 gnd.n6015 240.244
R6866 gnd.n6019 gnd.n5885 240.244
R6867 gnd.n6026 gnd.n1471 240.244
R6868 gnd.n1346 gnd.n1345 240.132
R6869 gnd.n5606 gnd.n5605 240.132
R6870 gnd.n6884 gnd.n847 225.874
R6871 gnd.n6885 gnd.n6884 225.874
R6872 gnd.n6886 gnd.n6885 225.874
R6873 gnd.n6886 gnd.n841 225.874
R6874 gnd.n6894 gnd.n841 225.874
R6875 gnd.n6895 gnd.n6894 225.874
R6876 gnd.n6896 gnd.n6895 225.874
R6877 gnd.n6896 gnd.n835 225.874
R6878 gnd.n6904 gnd.n835 225.874
R6879 gnd.n6905 gnd.n6904 225.874
R6880 gnd.n6906 gnd.n6905 225.874
R6881 gnd.n6906 gnd.n829 225.874
R6882 gnd.n6914 gnd.n829 225.874
R6883 gnd.n6915 gnd.n6914 225.874
R6884 gnd.n6916 gnd.n6915 225.874
R6885 gnd.n6916 gnd.n823 225.874
R6886 gnd.n6924 gnd.n823 225.874
R6887 gnd.n6925 gnd.n6924 225.874
R6888 gnd.n6926 gnd.n6925 225.874
R6889 gnd.n6926 gnd.n817 225.874
R6890 gnd.n6934 gnd.n817 225.874
R6891 gnd.n6935 gnd.n6934 225.874
R6892 gnd.n6936 gnd.n6935 225.874
R6893 gnd.n6936 gnd.n811 225.874
R6894 gnd.n6944 gnd.n811 225.874
R6895 gnd.n6945 gnd.n6944 225.874
R6896 gnd.n6946 gnd.n6945 225.874
R6897 gnd.n6946 gnd.n805 225.874
R6898 gnd.n6954 gnd.n805 225.874
R6899 gnd.n6955 gnd.n6954 225.874
R6900 gnd.n6956 gnd.n6955 225.874
R6901 gnd.n6956 gnd.n799 225.874
R6902 gnd.n6964 gnd.n799 225.874
R6903 gnd.n6965 gnd.n6964 225.874
R6904 gnd.n6966 gnd.n6965 225.874
R6905 gnd.n6966 gnd.n793 225.874
R6906 gnd.n6974 gnd.n793 225.874
R6907 gnd.n6975 gnd.n6974 225.874
R6908 gnd.n6976 gnd.n6975 225.874
R6909 gnd.n6976 gnd.n787 225.874
R6910 gnd.n6984 gnd.n787 225.874
R6911 gnd.n6985 gnd.n6984 225.874
R6912 gnd.n6986 gnd.n6985 225.874
R6913 gnd.n6986 gnd.n781 225.874
R6914 gnd.n6994 gnd.n781 225.874
R6915 gnd.n6995 gnd.n6994 225.874
R6916 gnd.n6996 gnd.n6995 225.874
R6917 gnd.n6996 gnd.n775 225.874
R6918 gnd.n7004 gnd.n775 225.874
R6919 gnd.n7005 gnd.n7004 225.874
R6920 gnd.n7006 gnd.n7005 225.874
R6921 gnd.n7006 gnd.n769 225.874
R6922 gnd.n7014 gnd.n769 225.874
R6923 gnd.n7015 gnd.n7014 225.874
R6924 gnd.n7016 gnd.n7015 225.874
R6925 gnd.n7016 gnd.n763 225.874
R6926 gnd.n7024 gnd.n763 225.874
R6927 gnd.n7025 gnd.n7024 225.874
R6928 gnd.n7026 gnd.n7025 225.874
R6929 gnd.n7026 gnd.n757 225.874
R6930 gnd.n7034 gnd.n757 225.874
R6931 gnd.n7035 gnd.n7034 225.874
R6932 gnd.n7036 gnd.n7035 225.874
R6933 gnd.n7036 gnd.n751 225.874
R6934 gnd.n7044 gnd.n751 225.874
R6935 gnd.n7045 gnd.n7044 225.874
R6936 gnd.n7046 gnd.n7045 225.874
R6937 gnd.n7046 gnd.n745 225.874
R6938 gnd.n7054 gnd.n745 225.874
R6939 gnd.n7055 gnd.n7054 225.874
R6940 gnd.n7056 gnd.n7055 225.874
R6941 gnd.n7056 gnd.n739 225.874
R6942 gnd.n7064 gnd.n739 225.874
R6943 gnd.n7065 gnd.n7064 225.874
R6944 gnd.n7066 gnd.n7065 225.874
R6945 gnd.n7066 gnd.n733 225.874
R6946 gnd.n7074 gnd.n733 225.874
R6947 gnd.n7075 gnd.n7074 225.874
R6948 gnd.n7076 gnd.n7075 225.874
R6949 gnd.n7076 gnd.n727 225.874
R6950 gnd.n7084 gnd.n727 225.874
R6951 gnd.n7085 gnd.n7084 225.874
R6952 gnd.n7086 gnd.n7085 225.874
R6953 gnd.n7086 gnd.n721 225.874
R6954 gnd.n7094 gnd.n721 225.874
R6955 gnd.n7095 gnd.n7094 225.874
R6956 gnd.n7096 gnd.n7095 225.874
R6957 gnd.n7096 gnd.n715 225.874
R6958 gnd.n7104 gnd.n715 225.874
R6959 gnd.n7105 gnd.n7104 225.874
R6960 gnd.n7106 gnd.n7105 225.874
R6961 gnd.n7106 gnd.n709 225.874
R6962 gnd.n7114 gnd.n709 225.874
R6963 gnd.n7115 gnd.n7114 225.874
R6964 gnd.n7116 gnd.n7115 225.874
R6965 gnd.n7116 gnd.n703 225.874
R6966 gnd.n7124 gnd.n703 225.874
R6967 gnd.n7125 gnd.n7124 225.874
R6968 gnd.n7126 gnd.n7125 225.874
R6969 gnd.n7126 gnd.n697 225.874
R6970 gnd.n7134 gnd.n697 225.874
R6971 gnd.n7135 gnd.n7134 225.874
R6972 gnd.n7136 gnd.n7135 225.874
R6973 gnd.n7136 gnd.n691 225.874
R6974 gnd.n7144 gnd.n691 225.874
R6975 gnd.n7145 gnd.n7144 225.874
R6976 gnd.n7146 gnd.n7145 225.874
R6977 gnd.n7146 gnd.n685 225.874
R6978 gnd.n7154 gnd.n685 225.874
R6979 gnd.n7155 gnd.n7154 225.874
R6980 gnd.n7156 gnd.n7155 225.874
R6981 gnd.n7156 gnd.n679 225.874
R6982 gnd.n7164 gnd.n679 225.874
R6983 gnd.n7165 gnd.n7164 225.874
R6984 gnd.n7166 gnd.n7165 225.874
R6985 gnd.n7166 gnd.n673 225.874
R6986 gnd.n7174 gnd.n673 225.874
R6987 gnd.n7175 gnd.n7174 225.874
R6988 gnd.n7176 gnd.n7175 225.874
R6989 gnd.n7176 gnd.n667 225.874
R6990 gnd.n7184 gnd.n667 225.874
R6991 gnd.n7185 gnd.n7184 225.874
R6992 gnd.n7186 gnd.n7185 225.874
R6993 gnd.n7186 gnd.n661 225.874
R6994 gnd.n7194 gnd.n661 225.874
R6995 gnd.n7195 gnd.n7194 225.874
R6996 gnd.n7196 gnd.n7195 225.874
R6997 gnd.n7196 gnd.n655 225.874
R6998 gnd.n7204 gnd.n655 225.874
R6999 gnd.n7205 gnd.n7204 225.874
R7000 gnd.n7206 gnd.n7205 225.874
R7001 gnd.n7206 gnd.n649 225.874
R7002 gnd.n7214 gnd.n649 225.874
R7003 gnd.n7215 gnd.n7214 225.874
R7004 gnd.n7216 gnd.n7215 225.874
R7005 gnd.n7216 gnd.n643 225.874
R7006 gnd.n7224 gnd.n643 225.874
R7007 gnd.n7225 gnd.n7224 225.874
R7008 gnd.n7226 gnd.n7225 225.874
R7009 gnd.n7226 gnd.n637 225.874
R7010 gnd.n7234 gnd.n637 225.874
R7011 gnd.n7235 gnd.n7234 225.874
R7012 gnd.n7236 gnd.n7235 225.874
R7013 gnd.n7236 gnd.n631 225.874
R7014 gnd.n7244 gnd.n631 225.874
R7015 gnd.n7245 gnd.n7244 225.874
R7016 gnd.n7246 gnd.n7245 225.874
R7017 gnd.n7246 gnd.n625 225.874
R7018 gnd.n7254 gnd.n625 225.874
R7019 gnd.n7255 gnd.n7254 225.874
R7020 gnd.n7256 gnd.n7255 225.874
R7021 gnd.n7256 gnd.n619 225.874
R7022 gnd.n7264 gnd.n619 225.874
R7023 gnd.n7265 gnd.n7264 225.874
R7024 gnd.n7266 gnd.n7265 225.874
R7025 gnd.n7266 gnd.n613 225.874
R7026 gnd.n7274 gnd.n613 225.874
R7027 gnd.n7275 gnd.n7274 225.874
R7028 gnd.n7276 gnd.n7275 225.874
R7029 gnd.n7276 gnd.n607 225.874
R7030 gnd.n7284 gnd.n607 225.874
R7031 gnd.n7285 gnd.n7284 225.874
R7032 gnd.n7286 gnd.n7285 225.874
R7033 gnd.n7286 gnd.n601 225.874
R7034 gnd.n7294 gnd.n601 225.874
R7035 gnd.n7295 gnd.n7294 225.874
R7036 gnd.n7296 gnd.n7295 225.874
R7037 gnd.n7296 gnd.n595 225.874
R7038 gnd.n7304 gnd.n595 225.874
R7039 gnd.n7305 gnd.n7304 225.874
R7040 gnd.n7306 gnd.n7305 225.874
R7041 gnd.n7306 gnd.n589 225.874
R7042 gnd.n7314 gnd.n589 225.874
R7043 gnd.n7315 gnd.n7314 225.874
R7044 gnd.n7316 gnd.n7315 225.874
R7045 gnd.n7316 gnd.n583 225.874
R7046 gnd.n7324 gnd.n583 225.874
R7047 gnd.n7325 gnd.n7324 225.874
R7048 gnd.n7326 gnd.n7325 225.874
R7049 gnd.n7326 gnd.n577 225.874
R7050 gnd.n7334 gnd.n577 225.874
R7051 gnd.n7335 gnd.n7334 225.874
R7052 gnd.n7336 gnd.n7335 225.874
R7053 gnd.n7336 gnd.n571 225.874
R7054 gnd.n7344 gnd.n571 225.874
R7055 gnd.n7345 gnd.n7344 225.874
R7056 gnd.n7346 gnd.n7345 225.874
R7057 gnd.n7346 gnd.n565 225.874
R7058 gnd.n7354 gnd.n565 225.874
R7059 gnd.n7355 gnd.n7354 225.874
R7060 gnd.n7356 gnd.n7355 225.874
R7061 gnd.n7356 gnd.n559 225.874
R7062 gnd.n7364 gnd.n559 225.874
R7063 gnd.n7365 gnd.n7364 225.874
R7064 gnd.n7366 gnd.n7365 225.874
R7065 gnd.n7366 gnd.n553 225.874
R7066 gnd.n7374 gnd.n553 225.874
R7067 gnd.n7375 gnd.n7374 225.874
R7068 gnd.n7376 gnd.n7375 225.874
R7069 gnd.n7376 gnd.n547 225.874
R7070 gnd.n7384 gnd.n547 225.874
R7071 gnd.n7385 gnd.n7384 225.874
R7072 gnd.n7386 gnd.n7385 225.874
R7073 gnd.n7386 gnd.n541 225.874
R7074 gnd.n7394 gnd.n541 225.874
R7075 gnd.n7395 gnd.n7394 225.874
R7076 gnd.n7396 gnd.n7395 225.874
R7077 gnd.n3241 gnd.t225 224.174
R7078 gnd.n2738 gnd.t198 224.174
R7079 gnd.n1836 gnd.n1697 199.319
R7080 gnd.n1836 gnd.n1698 199.319
R7081 gnd.n1299 gnd.n1274 199.319
R7082 gnd.n1299 gnd.n1273 199.319
R7083 gnd.n1985 gnd.n1984 190.912
R7084 gnd.n6548 gnd.n6547 190.912
R7085 gnd.n1347 gnd.n1344 186.49
R7086 gnd.n5607 gnd.n5604 186.49
R7087 gnd.n4016 gnd.n4015 185
R7088 gnd.n4014 gnd.n4013 185
R7089 gnd.n3993 gnd.n3992 185
R7090 gnd.n4008 gnd.n4007 185
R7091 gnd.n4006 gnd.n4005 185
R7092 gnd.n3997 gnd.n3996 185
R7093 gnd.n4000 gnd.n3999 185
R7094 gnd.n3984 gnd.n3983 185
R7095 gnd.n3982 gnd.n3981 185
R7096 gnd.n3961 gnd.n3960 185
R7097 gnd.n3976 gnd.n3975 185
R7098 gnd.n3974 gnd.n3973 185
R7099 gnd.n3965 gnd.n3964 185
R7100 gnd.n3968 gnd.n3967 185
R7101 gnd.n3952 gnd.n3951 185
R7102 gnd.n3950 gnd.n3949 185
R7103 gnd.n3929 gnd.n3928 185
R7104 gnd.n3944 gnd.n3943 185
R7105 gnd.n3942 gnd.n3941 185
R7106 gnd.n3933 gnd.n3932 185
R7107 gnd.n3936 gnd.n3935 185
R7108 gnd.n3921 gnd.n3920 185
R7109 gnd.n3919 gnd.n3918 185
R7110 gnd.n3898 gnd.n3897 185
R7111 gnd.n3913 gnd.n3912 185
R7112 gnd.n3911 gnd.n3910 185
R7113 gnd.n3902 gnd.n3901 185
R7114 gnd.n3905 gnd.n3904 185
R7115 gnd.n3889 gnd.n3888 185
R7116 gnd.n3887 gnd.n3886 185
R7117 gnd.n3866 gnd.n3865 185
R7118 gnd.n3881 gnd.n3880 185
R7119 gnd.n3879 gnd.n3878 185
R7120 gnd.n3870 gnd.n3869 185
R7121 gnd.n3873 gnd.n3872 185
R7122 gnd.n3857 gnd.n3856 185
R7123 gnd.n3855 gnd.n3854 185
R7124 gnd.n3834 gnd.n3833 185
R7125 gnd.n3849 gnd.n3848 185
R7126 gnd.n3847 gnd.n3846 185
R7127 gnd.n3838 gnd.n3837 185
R7128 gnd.n3841 gnd.n3840 185
R7129 gnd.n3825 gnd.n3824 185
R7130 gnd.n3823 gnd.n3822 185
R7131 gnd.n3802 gnd.n3801 185
R7132 gnd.n3817 gnd.n3816 185
R7133 gnd.n3815 gnd.n3814 185
R7134 gnd.n3806 gnd.n3805 185
R7135 gnd.n3809 gnd.n3808 185
R7136 gnd.n3794 gnd.n3793 185
R7137 gnd.n3792 gnd.n3791 185
R7138 gnd.n3771 gnd.n3770 185
R7139 gnd.n3786 gnd.n3785 185
R7140 gnd.n3784 gnd.n3783 185
R7141 gnd.n3775 gnd.n3774 185
R7142 gnd.n3778 gnd.n3777 185
R7143 gnd.n3242 gnd.t224 178.987
R7144 gnd.n2739 gnd.t199 178.987
R7145 gnd.n1 gnd.t355 170.774
R7146 gnd.n9 gnd.t93 170.103
R7147 gnd.n8 gnd.t69 170.103
R7148 gnd.n7 gnd.t340 170.103
R7149 gnd.n6 gnd.t321 170.103
R7150 gnd.n5 gnd.t2 170.103
R7151 gnd.n4 gnd.t136 170.103
R7152 gnd.n3 gnd.t72 170.103
R7153 gnd.n2 gnd.t305 170.103
R7154 gnd.n1 gnd.t319 170.103
R7155 gnd.n5678 gnd.n5677 163.367
R7156 gnd.n5674 gnd.n5673 163.367
R7157 gnd.n5670 gnd.n5669 163.367
R7158 gnd.n5666 gnd.n5665 163.367
R7159 gnd.n5662 gnd.n5661 163.367
R7160 gnd.n5658 gnd.n5657 163.367
R7161 gnd.n5654 gnd.n5653 163.367
R7162 gnd.n5650 gnd.n5649 163.367
R7163 gnd.n5646 gnd.n5645 163.367
R7164 gnd.n5642 gnd.n5641 163.367
R7165 gnd.n5638 gnd.n5637 163.367
R7166 gnd.n5634 gnd.n5633 163.367
R7167 gnd.n5630 gnd.n5629 163.367
R7168 gnd.n5626 gnd.n5625 163.367
R7169 gnd.n5621 gnd.n5620 163.367
R7170 gnd.n5617 gnd.n5616 163.367
R7171 gnd.n5754 gnd.n5753 163.367
R7172 gnd.n5750 gnd.n5749 163.367
R7173 gnd.n5745 gnd.n5744 163.367
R7174 gnd.n5741 gnd.n5740 163.367
R7175 gnd.n5737 gnd.n5736 163.367
R7176 gnd.n5733 gnd.n5732 163.367
R7177 gnd.n5729 gnd.n5728 163.367
R7178 gnd.n5725 gnd.n5724 163.367
R7179 gnd.n5721 gnd.n5720 163.367
R7180 gnd.n5717 gnd.n5716 163.367
R7181 gnd.n5713 gnd.n5712 163.367
R7182 gnd.n5709 gnd.n5708 163.367
R7183 gnd.n5705 gnd.n5704 163.367
R7184 gnd.n5701 gnd.n5700 163.367
R7185 gnd.n5697 gnd.n5696 163.367
R7186 gnd.n5693 gnd.n5692 163.367
R7187 gnd.n5176 gnd.n1363 163.367
R7188 gnd.n1364 gnd.n1363 163.367
R7189 gnd.n5180 gnd.n1364 163.367
R7190 gnd.n5180 gnd.n5101 163.367
R7191 gnd.n5183 gnd.n5101 163.367
R7192 gnd.n5183 gnd.n5109 163.367
R7193 gnd.n5187 gnd.n5109 163.367
R7194 gnd.n5187 gnd.n2211 163.367
R7195 gnd.n5247 gnd.n2211 163.367
R7196 gnd.n5247 gnd.n2209 163.367
R7197 gnd.n5255 gnd.n2209 163.367
R7198 gnd.n5255 gnd.n2202 163.367
R7199 gnd.n5251 gnd.n2202 163.367
R7200 gnd.n5251 gnd.n2193 163.367
R7201 gnd.n2193 gnd.n2186 163.367
R7202 gnd.n5281 gnd.n2186 163.367
R7203 gnd.n5281 gnd.n2184 163.367
R7204 gnd.n5286 gnd.n2184 163.367
R7205 gnd.n5286 gnd.n2175 163.367
R7206 gnd.n2175 gnd.n2167 163.367
R7207 gnd.n5307 gnd.n2167 163.367
R7208 gnd.n5307 gnd.n2163 163.367
R7209 gnd.n5313 gnd.n2163 163.367
R7210 gnd.n5313 gnd.n2165 163.367
R7211 gnd.n2165 gnd.n2151 163.367
R7212 gnd.n2151 gnd.n2143 163.367
R7213 gnd.n5332 gnd.n2143 163.367
R7214 gnd.n5332 gnd.n2140 163.367
R7215 gnd.n5355 gnd.n2140 163.367
R7216 gnd.n5355 gnd.n2141 163.367
R7217 gnd.n2141 gnd.n2133 163.367
R7218 gnd.n5350 gnd.n2133 163.367
R7219 gnd.n5350 gnd.n5348 163.367
R7220 gnd.n5348 gnd.n5347 163.367
R7221 gnd.n5347 gnd.n5336 163.367
R7222 gnd.n5336 gnd.n2115 163.367
R7223 gnd.n5342 gnd.n2115 163.367
R7224 gnd.n5342 gnd.n2110 163.367
R7225 gnd.n5339 gnd.n2110 163.367
R7226 gnd.n5339 gnd.n2099 163.367
R7227 gnd.n2099 gnd.n2091 163.367
R7228 gnd.n5428 gnd.n2091 163.367
R7229 gnd.n5428 gnd.n2088 163.367
R7230 gnd.n5441 gnd.n2088 163.367
R7231 gnd.n5441 gnd.n2089 163.367
R7232 gnd.n2089 gnd.n2081 163.367
R7233 gnd.n5436 gnd.n2081 163.367
R7234 gnd.n5436 gnd.n2073 163.367
R7235 gnd.n5432 gnd.n2073 163.367
R7236 gnd.n5432 gnd.n2049 163.367
R7237 gnd.n2049 gnd.n2041 163.367
R7238 gnd.n5515 gnd.n2041 163.367
R7239 gnd.n5515 gnd.n2039 163.367
R7240 gnd.n5520 gnd.n2039 163.367
R7241 gnd.n5520 gnd.n2032 163.367
R7242 gnd.n5529 gnd.n2032 163.367
R7243 gnd.n5530 gnd.n5529 163.367
R7244 gnd.n5530 gnd.n2029 163.367
R7245 gnd.n5537 gnd.n2029 163.367
R7246 gnd.n5537 gnd.n2022 163.367
R7247 gnd.n5533 gnd.n2022 163.367
R7248 gnd.n5533 gnd.n2013 163.367
R7249 gnd.n5561 gnd.n2013 163.367
R7250 gnd.n5561 gnd.n2010 163.367
R7251 gnd.n5571 gnd.n2010 163.367
R7252 gnd.n5571 gnd.n2006 163.367
R7253 gnd.n5567 gnd.n2006 163.367
R7254 gnd.n5567 gnd.n1998 163.367
R7255 gnd.n1998 gnd.n1989 163.367
R7256 gnd.n5687 gnd.n1989 163.367
R7257 gnd.n5688 gnd.n5687 163.367
R7258 gnd.n1338 gnd.n1337 163.367
R7259 gnd.n6537 gnd.n1337 163.367
R7260 gnd.n6535 gnd.n6534 163.367
R7261 gnd.n6531 gnd.n6530 163.367
R7262 gnd.n6527 gnd.n6526 163.367
R7263 gnd.n6523 gnd.n6522 163.367
R7264 gnd.n6519 gnd.n6518 163.367
R7265 gnd.n6515 gnd.n6514 163.367
R7266 gnd.n6511 gnd.n6510 163.367
R7267 gnd.n6507 gnd.n6506 163.367
R7268 gnd.n6503 gnd.n6502 163.367
R7269 gnd.n6499 gnd.n6498 163.367
R7270 gnd.n6495 gnd.n6494 163.367
R7271 gnd.n6491 gnd.n6490 163.367
R7272 gnd.n6487 gnd.n6486 163.367
R7273 gnd.n6483 gnd.n6482 163.367
R7274 gnd.n6546 gnd.n1304 163.367
R7275 gnd.n5114 gnd.n5113 163.367
R7276 gnd.n5119 gnd.n5118 163.367
R7277 gnd.n5123 gnd.n5122 163.367
R7278 gnd.n5127 gnd.n5126 163.367
R7279 gnd.n5131 gnd.n5130 163.367
R7280 gnd.n5135 gnd.n5134 163.367
R7281 gnd.n5139 gnd.n5138 163.367
R7282 gnd.n5143 gnd.n5142 163.367
R7283 gnd.n5147 gnd.n5146 163.367
R7284 gnd.n5151 gnd.n5150 163.367
R7285 gnd.n5155 gnd.n5154 163.367
R7286 gnd.n5159 gnd.n5158 163.367
R7287 gnd.n5163 gnd.n5162 163.367
R7288 gnd.n5167 gnd.n5166 163.367
R7289 gnd.n5171 gnd.n5170 163.367
R7290 gnd.n6475 gnd.n1339 163.367
R7291 gnd.n6475 gnd.n1361 163.367
R7292 gnd.n5102 gnd.n1361 163.367
R7293 gnd.n5194 gnd.n5102 163.367
R7294 gnd.n5194 gnd.n5103 163.367
R7295 gnd.n5190 gnd.n5103 163.367
R7296 gnd.n5190 gnd.n5189 163.367
R7297 gnd.n5189 gnd.n5107 163.367
R7298 gnd.n5107 gnd.n2207 163.367
R7299 gnd.n5258 gnd.n2207 163.367
R7300 gnd.n5258 gnd.n2205 163.367
R7301 gnd.n5262 gnd.n2205 163.367
R7302 gnd.n5262 gnd.n2191 163.367
R7303 gnd.n5274 gnd.n2191 163.367
R7304 gnd.n5274 gnd.n2188 163.367
R7305 gnd.n5279 gnd.n2188 163.367
R7306 gnd.n5279 gnd.n2189 163.367
R7307 gnd.n2189 gnd.n2172 163.367
R7308 gnd.n5299 gnd.n2172 163.367
R7309 gnd.n5299 gnd.n2169 163.367
R7310 gnd.n5305 gnd.n2169 163.367
R7311 gnd.n5305 gnd.n2170 163.367
R7312 gnd.n2170 gnd.n2161 163.367
R7313 gnd.n2161 gnd.n2148 163.367
R7314 gnd.n5326 gnd.n2148 163.367
R7315 gnd.n5326 gnd.n2146 163.367
R7316 gnd.n5330 gnd.n2146 163.367
R7317 gnd.n5330 gnd.n2138 163.367
R7318 gnd.n5357 gnd.n2138 163.367
R7319 gnd.n5357 gnd.n2135 163.367
R7320 gnd.n5366 gnd.n2135 163.367
R7321 gnd.n5366 gnd.n2136 163.367
R7322 gnd.n5362 gnd.n2136 163.367
R7323 gnd.n5362 gnd.n5361 163.367
R7324 gnd.n5361 gnd.n2113 163.367
R7325 gnd.n5404 gnd.n2113 163.367
R7326 gnd.n5404 gnd.n2111 163.367
R7327 gnd.n5408 gnd.n2111 163.367
R7328 gnd.n5408 gnd.n2097 163.367
R7329 gnd.n5422 gnd.n2097 163.367
R7330 gnd.n5422 gnd.n2095 163.367
R7331 gnd.n5426 gnd.n2095 163.367
R7332 gnd.n5426 gnd.n2086 163.367
R7333 gnd.n5443 gnd.n2086 163.367
R7334 gnd.n5443 gnd.n2083 163.367
R7335 gnd.n5449 gnd.n2083 163.367
R7336 gnd.n5449 gnd.n2084 163.367
R7337 gnd.n2084 gnd.n2070 163.367
R7338 gnd.n2070 gnd.n2047 163.367
R7339 gnd.n5509 gnd.n2047 163.367
R7340 gnd.n5509 gnd.n2045 163.367
R7341 gnd.n5513 gnd.n2045 163.367
R7342 gnd.n5513 gnd.n2036 163.367
R7343 gnd.n5523 gnd.n2036 163.367
R7344 gnd.n5523 gnd.n2034 163.367
R7345 gnd.n5527 gnd.n2034 163.367
R7346 gnd.n5527 gnd.n2027 163.367
R7347 gnd.n5541 gnd.n2027 163.367
R7348 gnd.n5541 gnd.n2024 163.367
R7349 gnd.n5548 gnd.n2024 163.367
R7350 gnd.n5548 gnd.n2025 163.367
R7351 gnd.n5544 gnd.n2025 163.367
R7352 gnd.n5544 gnd.n2009 163.367
R7353 gnd.n5575 gnd.n2009 163.367
R7354 gnd.n5575 gnd.n2007 163.367
R7355 gnd.n5579 gnd.n2007 163.367
R7356 gnd.n5579 gnd.n1996 163.367
R7357 gnd.n5592 gnd.n1996 163.367
R7358 gnd.n5592 gnd.n1993 163.367
R7359 gnd.n5685 gnd.n1993 163.367
R7360 gnd.n5685 gnd.n1994 163.367
R7361 gnd.n5613 gnd.n5612 156.462
R7362 gnd.n3956 gnd.n3924 153.042
R7363 gnd.n4020 gnd.n4019 152.079
R7364 gnd.n3988 gnd.n3987 152.079
R7365 gnd.n3956 gnd.n3955 152.079
R7366 gnd.n1352 gnd.n1351 152
R7367 gnd.n1353 gnd.n1342 152
R7368 gnd.n1355 gnd.n1354 152
R7369 gnd.n1357 gnd.n1340 152
R7370 gnd.n1359 gnd.n1358 152
R7371 gnd.n5611 gnd.n5595 152
R7372 gnd.n5603 gnd.n5596 152
R7373 gnd.n5602 gnd.n5601 152
R7374 gnd.n5600 gnd.n5597 152
R7375 gnd.n5598 gnd.t179 150.546
R7376 gnd.t152 gnd.n3998 147.661
R7377 gnd.t266 gnd.n3966 147.661
R7378 gnd.t262 gnd.n3934 147.661
R7379 gnd.t307 gnd.n3903 147.661
R7380 gnd.t353 gnd.n3871 147.661
R7381 gnd.t349 gnd.n3839 147.661
R7382 gnd.t100 gnd.n3807 147.661
R7383 gnd.t289 gnd.n3776 147.661
R7384 gnd.n1834 gnd.n1817 143.351
R7385 gnd.n1319 gnd.n1303 143.351
R7386 gnd.n6545 gnd.n1303 143.351
R7387 gnd.n7404 gnd.n535 137.802
R7388 gnd.n7405 gnd.n7404 137.802
R7389 gnd.n7406 gnd.n7405 137.802
R7390 gnd.n7406 gnd.n529 137.802
R7391 gnd.n7414 gnd.n529 137.802
R7392 gnd.n7415 gnd.n7414 137.802
R7393 gnd.n7416 gnd.n7415 137.802
R7394 gnd.n7416 gnd.n523 137.802
R7395 gnd.n7424 gnd.n523 137.802
R7396 gnd.n7425 gnd.n7424 137.802
R7397 gnd.n7426 gnd.n7425 137.802
R7398 gnd.n7426 gnd.n517 137.802
R7399 gnd.n7434 gnd.n517 137.802
R7400 gnd.n7435 gnd.n7434 137.802
R7401 gnd.n7436 gnd.n7435 137.802
R7402 gnd.n7436 gnd.n511 137.802
R7403 gnd.n7444 gnd.n511 137.802
R7404 gnd.n7445 gnd.n7444 137.802
R7405 gnd.n7446 gnd.n7445 137.802
R7406 gnd.n7446 gnd.n505 137.802
R7407 gnd.n7454 gnd.n505 137.802
R7408 gnd.n7455 gnd.n7454 137.802
R7409 gnd.n7456 gnd.n7455 137.802
R7410 gnd.n7456 gnd.n499 137.802
R7411 gnd.n7464 gnd.n499 137.802
R7412 gnd.n7465 gnd.n7464 137.802
R7413 gnd.n7466 gnd.n7465 137.802
R7414 gnd.n7466 gnd.n493 137.802
R7415 gnd.n7474 gnd.n493 137.802
R7416 gnd.n7475 gnd.n7474 137.802
R7417 gnd.n7476 gnd.n7475 137.802
R7418 gnd.n7476 gnd.n487 137.802
R7419 gnd.n7484 gnd.n487 137.802
R7420 gnd.n7485 gnd.n7484 137.802
R7421 gnd.n7486 gnd.n7485 137.802
R7422 gnd.n7486 gnd.n481 137.802
R7423 gnd.n7494 gnd.n481 137.802
R7424 gnd.n7495 gnd.n7494 137.802
R7425 gnd.n7496 gnd.n7495 137.802
R7426 gnd.n7496 gnd.n475 137.802
R7427 gnd.n7504 gnd.n475 137.802
R7428 gnd.n7505 gnd.n7504 137.802
R7429 gnd.n7506 gnd.n7505 137.802
R7430 gnd.n7506 gnd.n469 137.802
R7431 gnd.n7514 gnd.n469 137.802
R7432 gnd.n7515 gnd.n7514 137.802
R7433 gnd.n7516 gnd.n7515 137.802
R7434 gnd.n7516 gnd.n463 137.802
R7435 gnd.n7524 gnd.n463 137.802
R7436 gnd.n7525 gnd.n7524 137.802
R7437 gnd.n7526 gnd.n7525 137.802
R7438 gnd.n7526 gnd.n457 137.802
R7439 gnd.n7534 gnd.n457 137.802
R7440 gnd.n7535 gnd.n7534 137.802
R7441 gnd.n7536 gnd.n7535 137.802
R7442 gnd.n7536 gnd.n451 137.802
R7443 gnd.n7544 gnd.n451 137.802
R7444 gnd.n7545 gnd.n7544 137.802
R7445 gnd.n7546 gnd.n7545 137.802
R7446 gnd.n7546 gnd.n445 137.802
R7447 gnd.n7554 gnd.n445 137.802
R7448 gnd.n7555 gnd.n7554 137.802
R7449 gnd.n7556 gnd.n7555 137.802
R7450 gnd.n7556 gnd.n439 137.802
R7451 gnd.n7564 gnd.n439 137.802
R7452 gnd.n7565 gnd.n7564 137.802
R7453 gnd.n7566 gnd.n7565 137.802
R7454 gnd.n7566 gnd.n433 137.802
R7455 gnd.n7574 gnd.n433 137.802
R7456 gnd.n7575 gnd.n7574 137.802
R7457 gnd.n7576 gnd.n7575 137.802
R7458 gnd.n7576 gnd.n427 137.802
R7459 gnd.n7584 gnd.n427 137.802
R7460 gnd.n7585 gnd.n7584 137.802
R7461 gnd.n7586 gnd.n7585 137.802
R7462 gnd.n7586 gnd.n421 137.802
R7463 gnd.n7594 gnd.n421 137.802
R7464 gnd.n7595 gnd.n7594 137.802
R7465 gnd.n7596 gnd.n7595 137.802
R7466 gnd.n7596 gnd.n415 137.802
R7467 gnd.n7606 gnd.n415 137.802
R7468 gnd.n7607 gnd.n7606 137.802
R7469 gnd.n7608 gnd.n7607 137.802
R7470 gnd.n1349 gnd.t213 130.484
R7471 gnd.n1358 gnd.t186 126.766
R7472 gnd.n1356 gnd.t153 126.766
R7473 gnd.n1342 gnd.t200 126.766
R7474 gnd.n1350 gnd.t255 126.766
R7475 gnd.n5599 gnd.t172 126.766
R7476 gnd.n5601 gnd.t226 126.766
R7477 gnd.n5610 gnd.t210 126.766
R7478 gnd.n5612 gnd.t239 126.766
R7479 gnd.n4015 gnd.n4014 104.615
R7480 gnd.n4014 gnd.n3992 104.615
R7481 gnd.n4007 gnd.n3992 104.615
R7482 gnd.n4007 gnd.n4006 104.615
R7483 gnd.n4006 gnd.n3996 104.615
R7484 gnd.n3999 gnd.n3996 104.615
R7485 gnd.n3983 gnd.n3982 104.615
R7486 gnd.n3982 gnd.n3960 104.615
R7487 gnd.n3975 gnd.n3960 104.615
R7488 gnd.n3975 gnd.n3974 104.615
R7489 gnd.n3974 gnd.n3964 104.615
R7490 gnd.n3967 gnd.n3964 104.615
R7491 gnd.n3951 gnd.n3950 104.615
R7492 gnd.n3950 gnd.n3928 104.615
R7493 gnd.n3943 gnd.n3928 104.615
R7494 gnd.n3943 gnd.n3942 104.615
R7495 gnd.n3942 gnd.n3932 104.615
R7496 gnd.n3935 gnd.n3932 104.615
R7497 gnd.n3920 gnd.n3919 104.615
R7498 gnd.n3919 gnd.n3897 104.615
R7499 gnd.n3912 gnd.n3897 104.615
R7500 gnd.n3912 gnd.n3911 104.615
R7501 gnd.n3911 gnd.n3901 104.615
R7502 gnd.n3904 gnd.n3901 104.615
R7503 gnd.n3888 gnd.n3887 104.615
R7504 gnd.n3887 gnd.n3865 104.615
R7505 gnd.n3880 gnd.n3865 104.615
R7506 gnd.n3880 gnd.n3879 104.615
R7507 gnd.n3879 gnd.n3869 104.615
R7508 gnd.n3872 gnd.n3869 104.615
R7509 gnd.n3856 gnd.n3855 104.615
R7510 gnd.n3855 gnd.n3833 104.615
R7511 gnd.n3848 gnd.n3833 104.615
R7512 gnd.n3848 gnd.n3847 104.615
R7513 gnd.n3847 gnd.n3837 104.615
R7514 gnd.n3840 gnd.n3837 104.615
R7515 gnd.n3824 gnd.n3823 104.615
R7516 gnd.n3823 gnd.n3801 104.615
R7517 gnd.n3816 gnd.n3801 104.615
R7518 gnd.n3816 gnd.n3815 104.615
R7519 gnd.n3815 gnd.n3805 104.615
R7520 gnd.n3808 gnd.n3805 104.615
R7521 gnd.n3793 gnd.n3792 104.615
R7522 gnd.n3792 gnd.n3770 104.615
R7523 gnd.n3785 gnd.n3770 104.615
R7524 gnd.n3785 gnd.n3784 104.615
R7525 gnd.n3784 gnd.n3774 104.615
R7526 gnd.n3777 gnd.n3774 104.615
R7527 gnd.n3167 gnd.t245 100.632
R7528 gnd.n2712 gnd.t184 100.632
R7529 gnd.n7909 gnd.n138 99.6594
R7530 gnd.n7907 gnd.n7906 99.6594
R7531 gnd.n7902 gnd.n145 99.6594
R7532 gnd.n7900 gnd.n7899 99.6594
R7533 gnd.n7895 gnd.n152 99.6594
R7534 gnd.n7893 gnd.n7892 99.6594
R7535 gnd.n7888 gnd.n159 99.6594
R7536 gnd.n7886 gnd.n7885 99.6594
R7537 gnd.n7878 gnd.n166 99.6594
R7538 gnd.n7876 gnd.n7875 99.6594
R7539 gnd.n7871 gnd.n173 99.6594
R7540 gnd.n7869 gnd.n7868 99.6594
R7541 gnd.n7864 gnd.n180 99.6594
R7542 gnd.n7862 gnd.n7861 99.6594
R7543 gnd.n7857 gnd.n187 99.6594
R7544 gnd.n7855 gnd.n7854 99.6594
R7545 gnd.n7850 gnd.n194 99.6594
R7546 gnd.n7848 gnd.n7847 99.6594
R7547 gnd.n199 gnd.n198 99.6594
R7548 gnd.n6042 gnd.n1685 99.6594
R7549 gnd.n1842 gnd.n1691 99.6594
R7550 gnd.n1849 gnd.n1692 99.6594
R7551 gnd.n1851 gnd.n1693 99.6594
R7552 gnd.n1859 gnd.n1694 99.6594
R7553 gnd.n1861 gnd.n1695 99.6594
R7554 gnd.n1869 gnd.n1696 99.6594
R7555 gnd.n1871 gnd.n1697 99.6594
R7556 gnd.n1981 gnd.n1699 99.6594
R7557 gnd.n1977 gnd.n1700 99.6594
R7558 gnd.n1973 gnd.n1701 99.6594
R7559 gnd.n1969 gnd.n1702 99.6594
R7560 gnd.n1965 gnd.n1703 99.6594
R7561 gnd.n1961 gnd.n1704 99.6594
R7562 gnd.n1957 gnd.n1705 99.6594
R7563 gnd.n1953 gnd.n1706 99.6594
R7564 gnd.n1949 gnd.n1707 99.6594
R7565 gnd.n1898 gnd.n1708 99.6594
R7566 gnd.n6576 gnd.n6575 99.6594
R7567 gnd.n6571 gnd.n1280 99.6594
R7568 gnd.n6567 gnd.n1279 99.6594
R7569 gnd.n6563 gnd.n1278 99.6594
R7570 gnd.n6559 gnd.n1277 99.6594
R7571 gnd.n6555 gnd.n1276 99.6594
R7572 gnd.n6551 gnd.n1275 99.6594
R7573 gnd.n4774 gnd.n1273 99.6594
R7574 gnd.n4781 gnd.n1272 99.6594
R7575 gnd.n4785 gnd.n1271 99.6594
R7576 gnd.n4791 gnd.n1270 99.6594
R7577 gnd.n4795 gnd.n1269 99.6594
R7578 gnd.n4801 gnd.n1268 99.6594
R7579 gnd.n4805 gnd.n1267 99.6594
R7580 gnd.n4811 gnd.n1266 99.6594
R7581 gnd.n4815 gnd.n1265 99.6594
R7582 gnd.n4820 gnd.n1264 99.6594
R7583 gnd.n4823 gnd.n1263 99.6594
R7584 gnd.n4196 gnd.n2672 99.6594
R7585 gnd.n4204 gnd.n4203 99.6594
R7586 gnd.n4207 gnd.n4206 99.6594
R7587 gnd.n4214 gnd.n4213 99.6594
R7588 gnd.n4217 gnd.n4216 99.6594
R7589 gnd.n4224 gnd.n4223 99.6594
R7590 gnd.n4227 gnd.n4226 99.6594
R7591 gnd.n4234 gnd.n4233 99.6594
R7592 gnd.n4237 gnd.n4236 99.6594
R7593 gnd.n4244 gnd.n4243 99.6594
R7594 gnd.n4247 gnd.n4246 99.6594
R7595 gnd.n4254 gnd.n4253 99.6594
R7596 gnd.n4257 gnd.n4256 99.6594
R7597 gnd.n4264 gnd.n4263 99.6594
R7598 gnd.n4267 gnd.n4266 99.6594
R7599 gnd.n4274 gnd.n4273 99.6594
R7600 gnd.n4277 gnd.n4276 99.6594
R7601 gnd.n4285 gnd.n4284 99.6594
R7602 gnd.n4288 gnd.n4287 99.6594
R7603 gnd.n4138 gnd.n2695 99.6594
R7604 gnd.n4136 gnd.n2694 99.6594
R7605 gnd.n4132 gnd.n2693 99.6594
R7606 gnd.n4128 gnd.n2692 99.6594
R7607 gnd.n4124 gnd.n2691 99.6594
R7608 gnd.n4120 gnd.n2690 99.6594
R7609 gnd.n4116 gnd.n2689 99.6594
R7610 gnd.n4048 gnd.n2688 99.6594
R7611 gnd.n3379 gnd.n3110 99.6594
R7612 gnd.n3136 gnd.n3117 99.6594
R7613 gnd.n3138 gnd.n3118 99.6594
R7614 gnd.n3146 gnd.n3119 99.6594
R7615 gnd.n3148 gnd.n3120 99.6594
R7616 gnd.n3156 gnd.n3121 99.6594
R7617 gnd.n3158 gnd.n3122 99.6594
R7618 gnd.n3166 gnd.n3123 99.6594
R7619 gnd.n4106 gnd.n2675 99.6594
R7620 gnd.n4102 gnd.n2676 99.6594
R7621 gnd.n4098 gnd.n2677 99.6594
R7622 gnd.n4094 gnd.n2678 99.6594
R7623 gnd.n4090 gnd.n2679 99.6594
R7624 gnd.n4086 gnd.n2680 99.6594
R7625 gnd.n4082 gnd.n2681 99.6594
R7626 gnd.n4078 gnd.n2682 99.6594
R7627 gnd.n4074 gnd.n2683 99.6594
R7628 gnd.n4070 gnd.n2684 99.6594
R7629 gnd.n4066 gnd.n2685 99.6594
R7630 gnd.n4062 gnd.n2686 99.6594
R7631 gnd.n4058 gnd.n2687 99.6594
R7632 gnd.n3294 gnd.n3293 99.6594
R7633 gnd.n3288 gnd.n3205 99.6594
R7634 gnd.n3285 gnd.n3206 99.6594
R7635 gnd.n3281 gnd.n3207 99.6594
R7636 gnd.n3277 gnd.n3208 99.6594
R7637 gnd.n3273 gnd.n3209 99.6594
R7638 gnd.n3269 gnd.n3210 99.6594
R7639 gnd.n3265 gnd.n3211 99.6594
R7640 gnd.n3261 gnd.n3212 99.6594
R7641 gnd.n3257 gnd.n3213 99.6594
R7642 gnd.n3253 gnd.n3214 99.6594
R7643 gnd.n3249 gnd.n3215 99.6594
R7644 gnd.n3296 gnd.n3204 99.6594
R7645 gnd.n7778 gnd.n7777 99.6594
R7646 gnd.n7783 gnd.n7782 99.6594
R7647 gnd.n7786 gnd.n7785 99.6594
R7648 gnd.n7791 gnd.n7790 99.6594
R7649 gnd.n7794 gnd.n7793 99.6594
R7650 gnd.n7799 gnd.n7798 99.6594
R7651 gnd.n7802 gnd.n7801 99.6594
R7652 gnd.n7807 gnd.n7805 99.6594
R7653 gnd.n7919 gnd.n125 99.6594
R7654 gnd.n1710 gnd.n1709 99.6594
R7655 gnd.n5933 gnd.n1711 99.6594
R7656 gnd.n5927 gnd.n1712 99.6594
R7657 gnd.n5944 gnd.n1713 99.6594
R7658 gnd.n5957 gnd.n1714 99.6594
R7659 gnd.n5915 gnd.n1715 99.6594
R7660 gnd.n5968 gnd.n1716 99.6594
R7661 gnd.n5981 gnd.n1717 99.6594
R7662 gnd.n5903 gnd.n1718 99.6594
R7663 gnd.n2406 gnd.n1253 99.6594
R7664 gnd.n2408 gnd.n1254 99.6594
R7665 gnd.n2417 gnd.n1255 99.6594
R7666 gnd.n2425 gnd.n1256 99.6594
R7667 gnd.n2427 gnd.n1257 99.6594
R7668 gnd.n2437 gnd.n1258 99.6594
R7669 gnd.n2445 gnd.n1259 99.6594
R7670 gnd.n2447 gnd.n1260 99.6594
R7671 gnd.n4925 gnd.n1261 99.6594
R7672 gnd.n4434 gnd.n4326 99.6594
R7673 gnd.n4433 gnd.n4432 99.6594
R7674 gnd.n4426 gnd.n4329 99.6594
R7675 gnd.n4425 gnd.n4424 99.6594
R7676 gnd.n4418 gnd.n4335 99.6594
R7677 gnd.n4417 gnd.n4416 99.6594
R7678 gnd.n4410 gnd.n4341 99.6594
R7679 gnd.n4409 gnd.n4408 99.6594
R7680 gnd.n4398 gnd.n4347 99.6594
R7681 gnd.n4435 gnd.n4434 99.6594
R7682 gnd.n4432 gnd.n4431 99.6594
R7683 gnd.n4427 gnd.n4426 99.6594
R7684 gnd.n4424 gnd.n4423 99.6594
R7685 gnd.n4419 gnd.n4418 99.6594
R7686 gnd.n4416 gnd.n4415 99.6594
R7687 gnd.n4411 gnd.n4410 99.6594
R7688 gnd.n4408 gnd.n4407 99.6594
R7689 gnd.n4399 gnd.n4398 99.6594
R7690 gnd.n2450 gnd.n1261 99.6594
R7691 gnd.n2446 gnd.n1260 99.6594
R7692 gnd.n2438 gnd.n1259 99.6594
R7693 gnd.n2428 gnd.n1258 99.6594
R7694 gnd.n2426 gnd.n1257 99.6594
R7695 gnd.n2418 gnd.n1256 99.6594
R7696 gnd.n2409 gnd.n1255 99.6594
R7697 gnd.n2407 gnd.n1254 99.6594
R7698 gnd.n2338 gnd.n1253 99.6594
R7699 gnd.n5932 gnd.n1710 99.6594
R7700 gnd.n5926 gnd.n1711 99.6594
R7701 gnd.n5945 gnd.n1712 99.6594
R7702 gnd.n5956 gnd.n1713 99.6594
R7703 gnd.n5914 gnd.n1714 99.6594
R7704 gnd.n5969 gnd.n1715 99.6594
R7705 gnd.n5980 gnd.n1716 99.6594
R7706 gnd.n5902 gnd.n1717 99.6594
R7707 gnd.n5898 gnd.n1718 99.6594
R7708 gnd.n7806 gnd.n125 99.6594
R7709 gnd.n7805 gnd.n7804 99.6594
R7710 gnd.n7801 gnd.n7800 99.6594
R7711 gnd.n7798 gnd.n7797 99.6594
R7712 gnd.n7793 gnd.n7792 99.6594
R7713 gnd.n7790 gnd.n7789 99.6594
R7714 gnd.n7785 gnd.n7784 99.6594
R7715 gnd.n7782 gnd.n7781 99.6594
R7716 gnd.n7777 gnd.n7776 99.6594
R7717 gnd.n3294 gnd.n3217 99.6594
R7718 gnd.n3286 gnd.n3205 99.6594
R7719 gnd.n3282 gnd.n3206 99.6594
R7720 gnd.n3278 gnd.n3207 99.6594
R7721 gnd.n3274 gnd.n3208 99.6594
R7722 gnd.n3270 gnd.n3209 99.6594
R7723 gnd.n3266 gnd.n3210 99.6594
R7724 gnd.n3262 gnd.n3211 99.6594
R7725 gnd.n3258 gnd.n3212 99.6594
R7726 gnd.n3254 gnd.n3213 99.6594
R7727 gnd.n3250 gnd.n3214 99.6594
R7728 gnd.n3246 gnd.n3215 99.6594
R7729 gnd.n3297 gnd.n3296 99.6594
R7730 gnd.n4061 gnd.n2687 99.6594
R7731 gnd.n4065 gnd.n2686 99.6594
R7732 gnd.n4069 gnd.n2685 99.6594
R7733 gnd.n4073 gnd.n2684 99.6594
R7734 gnd.n4077 gnd.n2683 99.6594
R7735 gnd.n4081 gnd.n2682 99.6594
R7736 gnd.n4085 gnd.n2681 99.6594
R7737 gnd.n4089 gnd.n2680 99.6594
R7738 gnd.n4093 gnd.n2679 99.6594
R7739 gnd.n4097 gnd.n2678 99.6594
R7740 gnd.n4101 gnd.n2677 99.6594
R7741 gnd.n4105 gnd.n2676 99.6594
R7742 gnd.n2716 gnd.n2675 99.6594
R7743 gnd.n3380 gnd.n3379 99.6594
R7744 gnd.n3139 gnd.n3117 99.6594
R7745 gnd.n3145 gnd.n3118 99.6594
R7746 gnd.n3149 gnd.n3119 99.6594
R7747 gnd.n3155 gnd.n3120 99.6594
R7748 gnd.n3159 gnd.n3121 99.6594
R7749 gnd.n3165 gnd.n3122 99.6594
R7750 gnd.n3123 gnd.n3107 99.6594
R7751 gnd.n4115 gnd.n2688 99.6594
R7752 gnd.n4119 gnd.n2689 99.6594
R7753 gnd.n4123 gnd.n2690 99.6594
R7754 gnd.n4127 gnd.n2691 99.6594
R7755 gnd.n4131 gnd.n2692 99.6594
R7756 gnd.n4135 gnd.n2693 99.6594
R7757 gnd.n4139 gnd.n2694 99.6594
R7758 gnd.n2697 gnd.n2695 99.6594
R7759 gnd.n4197 gnd.n4196 99.6594
R7760 gnd.n4205 gnd.n4204 99.6594
R7761 gnd.n4206 gnd.n4189 99.6594
R7762 gnd.n4215 gnd.n4214 99.6594
R7763 gnd.n4216 gnd.n4185 99.6594
R7764 gnd.n4225 gnd.n4224 99.6594
R7765 gnd.n4226 gnd.n4181 99.6594
R7766 gnd.n4235 gnd.n4234 99.6594
R7767 gnd.n4236 gnd.n4174 99.6594
R7768 gnd.n4245 gnd.n4244 99.6594
R7769 gnd.n4246 gnd.n4170 99.6594
R7770 gnd.n4255 gnd.n4254 99.6594
R7771 gnd.n4256 gnd.n4166 99.6594
R7772 gnd.n4265 gnd.n4264 99.6594
R7773 gnd.n4266 gnd.n4162 99.6594
R7774 gnd.n4275 gnd.n4274 99.6594
R7775 gnd.n4276 gnd.n4158 99.6594
R7776 gnd.n4286 gnd.n4285 99.6594
R7777 gnd.n4289 gnd.n4288 99.6594
R7778 gnd.n4765 gnd.n1263 99.6594
R7779 gnd.n4814 gnd.n1264 99.6594
R7780 gnd.n4812 gnd.n1265 99.6594
R7781 gnd.n4804 gnd.n1266 99.6594
R7782 gnd.n4802 gnd.n1267 99.6594
R7783 gnd.n4794 gnd.n1268 99.6594
R7784 gnd.n4792 gnd.n1269 99.6594
R7785 gnd.n4784 gnd.n1270 99.6594
R7786 gnd.n4782 gnd.n1271 99.6594
R7787 gnd.n4775 gnd.n1272 99.6594
R7788 gnd.n6550 gnd.n1274 99.6594
R7789 gnd.n6554 gnd.n1275 99.6594
R7790 gnd.n6558 gnd.n1276 99.6594
R7791 gnd.n6562 gnd.n1277 99.6594
R7792 gnd.n6566 gnd.n1278 99.6594
R7793 gnd.n6570 gnd.n1279 99.6594
R7794 gnd.n1281 gnd.n1280 99.6594
R7795 gnd.n6576 gnd.n1250 99.6594
R7796 gnd.n6043 gnd.n6042 99.6594
R7797 gnd.n1848 gnd.n1691 99.6594
R7798 gnd.n1852 gnd.n1692 99.6594
R7799 gnd.n1858 gnd.n1693 99.6594
R7800 gnd.n1862 gnd.n1694 99.6594
R7801 gnd.n1868 gnd.n1695 99.6594
R7802 gnd.n1872 gnd.n1696 99.6594
R7803 gnd.n1982 gnd.n1698 99.6594
R7804 gnd.n1978 gnd.n1699 99.6594
R7805 gnd.n1974 gnd.n1700 99.6594
R7806 gnd.n1970 gnd.n1701 99.6594
R7807 gnd.n1966 gnd.n1702 99.6594
R7808 gnd.n1962 gnd.n1703 99.6594
R7809 gnd.n1958 gnd.n1704 99.6594
R7810 gnd.n1954 gnd.n1705 99.6594
R7811 gnd.n1950 gnd.n1706 99.6594
R7812 gnd.n1897 gnd.n1707 99.6594
R7813 gnd.n1942 gnd.n1708 99.6594
R7814 gnd.n198 gnd.n195 99.6594
R7815 gnd.n7849 gnd.n7848 99.6594
R7816 gnd.n194 gnd.n188 99.6594
R7817 gnd.n7856 gnd.n7855 99.6594
R7818 gnd.n187 gnd.n181 99.6594
R7819 gnd.n7863 gnd.n7862 99.6594
R7820 gnd.n180 gnd.n174 99.6594
R7821 gnd.n7870 gnd.n7869 99.6594
R7822 gnd.n173 gnd.n167 99.6594
R7823 gnd.n7877 gnd.n7876 99.6594
R7824 gnd.n166 gnd.n160 99.6594
R7825 gnd.n7887 gnd.n7886 99.6594
R7826 gnd.n159 gnd.n153 99.6594
R7827 gnd.n7894 gnd.n7893 99.6594
R7828 gnd.n152 gnd.n146 99.6594
R7829 gnd.n7901 gnd.n7900 99.6594
R7830 gnd.n145 gnd.n139 99.6594
R7831 gnd.n7908 gnd.n7907 99.6594
R7832 gnd.n138 gnd.n135 99.6594
R7833 gnd.n4972 gnd.n4971 99.6594
R7834 gnd.n2412 gnd.n2317 99.6594
R7835 gnd.n2414 gnd.n2318 99.6594
R7836 gnd.n2422 gnd.n2319 99.6594
R7837 gnd.n2432 gnd.n2320 99.6594
R7838 gnd.n2434 gnd.n2321 99.6594
R7839 gnd.n2442 gnd.n2322 99.6594
R7840 gnd.n2454 gnd.n2323 99.6594
R7841 gnd.n2456 gnd.n2324 99.6594
R7842 gnd.n4836 gnd.n2325 99.6594
R7843 gnd.n4838 gnd.n2326 99.6594
R7844 gnd.n4842 gnd.n2327 99.6594
R7845 gnd.n4848 gnd.n2328 99.6594
R7846 gnd.n4850 gnd.n2329 99.6594
R7847 gnd.n4972 gnd.n2331 99.6594
R7848 gnd.n2413 gnd.n2317 99.6594
R7849 gnd.n2421 gnd.n2318 99.6594
R7850 gnd.n2431 gnd.n2319 99.6594
R7851 gnd.n2433 gnd.n2320 99.6594
R7852 gnd.n2441 gnd.n2321 99.6594
R7853 gnd.n2453 gnd.n2322 99.6594
R7854 gnd.n2455 gnd.n2323 99.6594
R7855 gnd.n4835 gnd.n2324 99.6594
R7856 gnd.n4837 gnd.n2325 99.6594
R7857 gnd.n4841 gnd.n2326 99.6594
R7858 gnd.n4843 gnd.n2327 99.6594
R7859 gnd.n4849 gnd.n2328 99.6594
R7860 gnd.n4851 gnd.n2329 99.6594
R7861 gnd.n5938 gnd.n5872 99.6594
R7862 gnd.n5922 gnd.n5873 99.6594
R7863 gnd.n5951 gnd.n5874 99.6594
R7864 gnd.n5962 gnd.n5875 99.6594
R7865 gnd.n5910 gnd.n5876 99.6594
R7866 gnd.n5975 gnd.n5877 99.6594
R7867 gnd.n5987 gnd.n5878 99.6594
R7868 gnd.n5990 gnd.n5879 99.6594
R7869 gnd.n5894 gnd.n5880 99.6594
R7870 gnd.n6005 gnd.n5881 99.6594
R7871 gnd.n6009 gnd.n5882 99.6594
R7872 gnd.n6015 gnd.n5883 99.6594
R7873 gnd.n6019 gnd.n5884 99.6594
R7874 gnd.n6027 gnd.n6026 99.6594
R7875 gnd.n6027 gnd.n5885 99.6594
R7876 gnd.n6016 gnd.n5884 99.6594
R7877 gnd.n6008 gnd.n5883 99.6594
R7878 gnd.n6006 gnd.n5882 99.6594
R7879 gnd.n5895 gnd.n5881 99.6594
R7880 gnd.n5991 gnd.n5880 99.6594
R7881 gnd.n5988 gnd.n5879 99.6594
R7882 gnd.n5974 gnd.n5878 99.6594
R7883 gnd.n5911 gnd.n5877 99.6594
R7884 gnd.n5963 gnd.n5876 99.6594
R7885 gnd.n5950 gnd.n5875 99.6594
R7886 gnd.n5923 gnd.n5874 99.6594
R7887 gnd.n5939 gnd.n5873 99.6594
R7888 gnd.n5872 gnd.n1476 99.6594
R7889 gnd.n4844 gnd.t195 98.63
R7890 gnd.n122 gnd.t208 98.63
R7891 gnd.n5899 gnd.t221 98.63
R7892 gnd.n2448 gnd.t247 98.63
R7893 gnd.n1877 gnd.t191 98.63
R7894 gnd.n1899 gnd.t178 98.63
R7895 gnd.n201 gnd.t234 98.63
R7896 gnd.n7880 gnd.t158 98.63
R7897 gnd.n4178 gnd.t260 98.63
R7898 gnd.n4154 gnd.t232 98.63
R7899 gnd.n4350 gnd.t254 98.63
R7900 gnd.n4763 gnd.t250 98.63
R7901 gnd.n1297 gnd.t170 98.63
R7902 gnd.n5889 gnd.t166 98.63
R7903 gnd.n5110 gnd.t163 92.8196
R7904 gnd.n1986 gnd.t205 92.8196
R7905 gnd.n6479 gnd.t218 92.8118
R7906 gnd.n5614 gnd.t237 92.8118
R7907 gnd.n7608 gnd.n126 82.6814
R7908 gnd.n1349 gnd.n1348 81.8399
R7909 gnd.n3168 gnd.t244 74.8376
R7910 gnd.n2713 gnd.t185 74.8376
R7911 gnd.n5111 gnd.t162 72.8438
R7912 gnd.n1987 gnd.t206 72.8438
R7913 gnd.n1350 gnd.n1343 72.8411
R7914 gnd.n1356 gnd.n1341 72.8411
R7915 gnd.n5610 gnd.n5609 72.8411
R7916 gnd.n4845 gnd.t194 72.836
R7917 gnd.n6480 gnd.t217 72.836
R7918 gnd.n5615 gnd.t238 72.836
R7919 gnd.n123 gnd.t209 72.836
R7920 gnd.n5900 gnd.t220 72.836
R7921 gnd.n2449 gnd.t248 72.836
R7922 gnd.n1878 gnd.t190 72.836
R7923 gnd.n1900 gnd.t177 72.836
R7924 gnd.n202 gnd.t235 72.836
R7925 gnd.n7881 gnd.t159 72.836
R7926 gnd.n4179 gnd.t259 72.836
R7927 gnd.n4155 gnd.t231 72.836
R7928 gnd.n4351 gnd.t253 72.836
R7929 gnd.n4764 gnd.t251 72.836
R7930 gnd.n1298 gnd.t171 72.836
R7931 gnd.n5890 gnd.t167 72.836
R7932 gnd.n5678 gnd.n1801 71.676
R7933 gnd.n5674 gnd.n1802 71.676
R7934 gnd.n5670 gnd.n1803 71.676
R7935 gnd.n5666 gnd.n1804 71.676
R7936 gnd.n5662 gnd.n1805 71.676
R7937 gnd.n5658 gnd.n1806 71.676
R7938 gnd.n5654 gnd.n1807 71.676
R7939 gnd.n5650 gnd.n1808 71.676
R7940 gnd.n5646 gnd.n1809 71.676
R7941 gnd.n5642 gnd.n1810 71.676
R7942 gnd.n5638 gnd.n1811 71.676
R7943 gnd.n5634 gnd.n1812 71.676
R7944 gnd.n5630 gnd.n1813 71.676
R7945 gnd.n5626 gnd.n1814 71.676
R7946 gnd.n5621 gnd.n1815 71.676
R7947 gnd.n5617 gnd.n1816 71.676
R7948 gnd.n5754 gnd.n1834 71.676
R7949 gnd.n5750 gnd.n1833 71.676
R7950 gnd.n5745 gnd.n1832 71.676
R7951 gnd.n5741 gnd.n1831 71.676
R7952 gnd.n5737 gnd.n1830 71.676
R7953 gnd.n5733 gnd.n1829 71.676
R7954 gnd.n5729 gnd.n1828 71.676
R7955 gnd.n5725 gnd.n1827 71.676
R7956 gnd.n5721 gnd.n1826 71.676
R7957 gnd.n5717 gnd.n1825 71.676
R7958 gnd.n5713 gnd.n1824 71.676
R7959 gnd.n5709 gnd.n1823 71.676
R7960 gnd.n5705 gnd.n1822 71.676
R7961 gnd.n5701 gnd.n1821 71.676
R7962 gnd.n5697 gnd.n1820 71.676
R7963 gnd.n5693 gnd.n1819 71.676
R7964 gnd.n5689 gnd.n1818 71.676
R7965 gnd.n6543 gnd.n6542 71.676
R7966 gnd.n6537 gnd.n1305 71.676
R7967 gnd.n6534 gnd.n1306 71.676
R7968 gnd.n6530 gnd.n1307 71.676
R7969 gnd.n6526 gnd.n1308 71.676
R7970 gnd.n6522 gnd.n1309 71.676
R7971 gnd.n6518 gnd.n1310 71.676
R7972 gnd.n6514 gnd.n1311 71.676
R7973 gnd.n6510 gnd.n1312 71.676
R7974 gnd.n6506 gnd.n1313 71.676
R7975 gnd.n6502 gnd.n1314 71.676
R7976 gnd.n6498 gnd.n1315 71.676
R7977 gnd.n6494 gnd.n1316 71.676
R7978 gnd.n6490 gnd.n1317 71.676
R7979 gnd.n6486 gnd.n1318 71.676
R7980 gnd.n6482 gnd.n1319 71.676
R7981 gnd.n1320 gnd.n1304 71.676
R7982 gnd.n5114 gnd.n1321 71.676
R7983 gnd.n5119 gnd.n1322 71.676
R7984 gnd.n5123 gnd.n1323 71.676
R7985 gnd.n5127 gnd.n1324 71.676
R7986 gnd.n5131 gnd.n1325 71.676
R7987 gnd.n5135 gnd.n1326 71.676
R7988 gnd.n5139 gnd.n1327 71.676
R7989 gnd.n5143 gnd.n1328 71.676
R7990 gnd.n5147 gnd.n1329 71.676
R7991 gnd.n5151 gnd.n1330 71.676
R7992 gnd.n5155 gnd.n1331 71.676
R7993 gnd.n5159 gnd.n1332 71.676
R7994 gnd.n5163 gnd.n1333 71.676
R7995 gnd.n5167 gnd.n1334 71.676
R7996 gnd.n5171 gnd.n1335 71.676
R7997 gnd.n6543 gnd.n1338 71.676
R7998 gnd.n6535 gnd.n1305 71.676
R7999 gnd.n6531 gnd.n1306 71.676
R8000 gnd.n6527 gnd.n1307 71.676
R8001 gnd.n6523 gnd.n1308 71.676
R8002 gnd.n6519 gnd.n1309 71.676
R8003 gnd.n6515 gnd.n1310 71.676
R8004 gnd.n6511 gnd.n1311 71.676
R8005 gnd.n6507 gnd.n1312 71.676
R8006 gnd.n6503 gnd.n1313 71.676
R8007 gnd.n6499 gnd.n1314 71.676
R8008 gnd.n6495 gnd.n1315 71.676
R8009 gnd.n6491 gnd.n1316 71.676
R8010 gnd.n6487 gnd.n1317 71.676
R8011 gnd.n6483 gnd.n1318 71.676
R8012 gnd.n6546 gnd.n6545 71.676
R8013 gnd.n5113 gnd.n1320 71.676
R8014 gnd.n5118 gnd.n1321 71.676
R8015 gnd.n5122 gnd.n1322 71.676
R8016 gnd.n5126 gnd.n1323 71.676
R8017 gnd.n5130 gnd.n1324 71.676
R8018 gnd.n5134 gnd.n1325 71.676
R8019 gnd.n5138 gnd.n1326 71.676
R8020 gnd.n5142 gnd.n1327 71.676
R8021 gnd.n5146 gnd.n1328 71.676
R8022 gnd.n5150 gnd.n1329 71.676
R8023 gnd.n5154 gnd.n1330 71.676
R8024 gnd.n5158 gnd.n1331 71.676
R8025 gnd.n5162 gnd.n1332 71.676
R8026 gnd.n5166 gnd.n1333 71.676
R8027 gnd.n5170 gnd.n1334 71.676
R8028 gnd.n5174 gnd.n1335 71.676
R8029 gnd.n5692 gnd.n1818 71.676
R8030 gnd.n5696 gnd.n1819 71.676
R8031 gnd.n5700 gnd.n1820 71.676
R8032 gnd.n5704 gnd.n1821 71.676
R8033 gnd.n5708 gnd.n1822 71.676
R8034 gnd.n5712 gnd.n1823 71.676
R8035 gnd.n5716 gnd.n1824 71.676
R8036 gnd.n5720 gnd.n1825 71.676
R8037 gnd.n5724 gnd.n1826 71.676
R8038 gnd.n5728 gnd.n1827 71.676
R8039 gnd.n5732 gnd.n1828 71.676
R8040 gnd.n5736 gnd.n1829 71.676
R8041 gnd.n5740 gnd.n1830 71.676
R8042 gnd.n5744 gnd.n1831 71.676
R8043 gnd.n5749 gnd.n1832 71.676
R8044 gnd.n5753 gnd.n1833 71.676
R8045 gnd.n5616 gnd.n1817 71.676
R8046 gnd.n5620 gnd.n1816 71.676
R8047 gnd.n5625 gnd.n1815 71.676
R8048 gnd.n5629 gnd.n1814 71.676
R8049 gnd.n5633 gnd.n1813 71.676
R8050 gnd.n5637 gnd.n1812 71.676
R8051 gnd.n5641 gnd.n1811 71.676
R8052 gnd.n5645 gnd.n1810 71.676
R8053 gnd.n5649 gnd.n1809 71.676
R8054 gnd.n5653 gnd.n1808 71.676
R8055 gnd.n5657 gnd.n1807 71.676
R8056 gnd.n5661 gnd.n1806 71.676
R8057 gnd.n5665 gnd.n1805 71.676
R8058 gnd.n5669 gnd.n1804 71.676
R8059 gnd.n5673 gnd.n1803 71.676
R8060 gnd.n5677 gnd.n1802 71.676
R8061 gnd.n5680 gnd.n1801 71.676
R8062 gnd.n10 gnd.t36 69.1507
R8063 gnd.n18 gnd.t150 68.4792
R8064 gnd.n17 gnd.t342 68.4792
R8065 gnd.n16 gnd.t102 68.4792
R8066 gnd.n15 gnd.t264 68.4792
R8067 gnd.n14 gnd.t142 68.4792
R8068 gnd.n13 gnd.t323 68.4792
R8069 gnd.n12 gnd.t285 68.4792
R8070 gnd.n11 gnd.t297 68.4792
R8071 gnd.n10 gnd.t310 68.4792
R8072 gnd.n3295 gnd.n3199 64.369
R8073 gnd.n5116 gnd.n5111 59.5399
R8074 gnd.n5747 gnd.n1987 59.5399
R8075 gnd.n6481 gnd.n6480 59.5399
R8076 gnd.n5623 gnd.n5615 59.5399
R8077 gnd.n6478 gnd.n1359 59.1804
R8078 gnd.n4147 gnd.n2673 57.3586
R8079 gnd.n2946 gnd.t54 56.607
R8080 gnd.n60 gnd.t38 56.607
R8081 gnd.n2907 gnd.t49 56.407
R8082 gnd.n2926 gnd.t45 56.407
R8083 gnd.n21 gnd.t113 56.407
R8084 gnd.n40 gnd.t329 56.407
R8085 gnd.n2963 gnd.t85 55.8337
R8086 gnd.n2924 gnd.t334 55.8337
R8087 gnd.n2943 gnd.t51 55.8337
R8088 gnd.n77 gnd.t312 55.8337
R8089 gnd.n38 gnd.t115 55.8337
R8090 gnd.n57 gnd.t145 55.8337
R8091 gnd.n1347 gnd.n1346 54.358
R8092 gnd.n5607 gnd.n5606 54.358
R8093 gnd.n2946 gnd.n2945 53.0052
R8094 gnd.n2948 gnd.n2947 53.0052
R8095 gnd.n2950 gnd.n2949 53.0052
R8096 gnd.n2952 gnd.n2951 53.0052
R8097 gnd.n2954 gnd.n2953 53.0052
R8098 gnd.n2956 gnd.n2955 53.0052
R8099 gnd.n2958 gnd.n2957 53.0052
R8100 gnd.n2960 gnd.n2959 53.0052
R8101 gnd.n2962 gnd.n2961 53.0052
R8102 gnd.n2907 gnd.n2906 53.0052
R8103 gnd.n2909 gnd.n2908 53.0052
R8104 gnd.n2911 gnd.n2910 53.0052
R8105 gnd.n2913 gnd.n2912 53.0052
R8106 gnd.n2915 gnd.n2914 53.0052
R8107 gnd.n2917 gnd.n2916 53.0052
R8108 gnd.n2919 gnd.n2918 53.0052
R8109 gnd.n2921 gnd.n2920 53.0052
R8110 gnd.n2923 gnd.n2922 53.0052
R8111 gnd.n2926 gnd.n2925 53.0052
R8112 gnd.n2928 gnd.n2927 53.0052
R8113 gnd.n2930 gnd.n2929 53.0052
R8114 gnd.n2932 gnd.n2931 53.0052
R8115 gnd.n2934 gnd.n2933 53.0052
R8116 gnd.n2936 gnd.n2935 53.0052
R8117 gnd.n2938 gnd.n2937 53.0052
R8118 gnd.n2940 gnd.n2939 53.0052
R8119 gnd.n2942 gnd.n2941 53.0052
R8120 gnd.n76 gnd.n75 53.0052
R8121 gnd.n74 gnd.n73 53.0052
R8122 gnd.n72 gnd.n71 53.0052
R8123 gnd.n70 gnd.n69 53.0052
R8124 gnd.n68 gnd.n67 53.0052
R8125 gnd.n66 gnd.n65 53.0052
R8126 gnd.n64 gnd.n63 53.0052
R8127 gnd.n62 gnd.n61 53.0052
R8128 gnd.n60 gnd.n59 53.0052
R8129 gnd.n37 gnd.n36 53.0052
R8130 gnd.n35 gnd.n34 53.0052
R8131 gnd.n33 gnd.n32 53.0052
R8132 gnd.n31 gnd.n30 53.0052
R8133 gnd.n29 gnd.n28 53.0052
R8134 gnd.n27 gnd.n26 53.0052
R8135 gnd.n25 gnd.n24 53.0052
R8136 gnd.n23 gnd.n22 53.0052
R8137 gnd.n21 gnd.n20 53.0052
R8138 gnd.n56 gnd.n55 53.0052
R8139 gnd.n54 gnd.n53 53.0052
R8140 gnd.n52 gnd.n51 53.0052
R8141 gnd.n50 gnd.n49 53.0052
R8142 gnd.n48 gnd.n47 53.0052
R8143 gnd.n46 gnd.n45 53.0052
R8144 gnd.n44 gnd.n43 53.0052
R8145 gnd.n42 gnd.n41 53.0052
R8146 gnd.n40 gnd.n39 53.0052
R8147 gnd.n5598 gnd.n5597 52.4801
R8148 gnd.n3999 gnd.t152 52.3082
R8149 gnd.n3967 gnd.t266 52.3082
R8150 gnd.n3935 gnd.t262 52.3082
R8151 gnd.n3904 gnd.t307 52.3082
R8152 gnd.n3872 gnd.t353 52.3082
R8153 gnd.n3840 gnd.t349 52.3082
R8154 gnd.n3808 gnd.t100 52.3082
R8155 gnd.n3777 gnd.t289 52.3082
R8156 gnd.n4442 gnd.n4148 51.6227
R8157 gnd.n7917 gnd.n128 51.6227
R8158 gnd.n3829 gnd.n3797 51.4173
R8159 gnd.n3893 gnd.n3892 50.455
R8160 gnd.n3861 gnd.n3860 50.455
R8161 gnd.n3829 gnd.n3828 50.455
R8162 gnd.n3242 gnd.n3241 45.1884
R8163 gnd.n2739 gnd.n2738 45.1884
R8164 gnd.n5682 gnd.n5613 44.3322
R8165 gnd.n1350 gnd.n1349 44.3189
R8166 gnd.n4846 gnd.n4845 42.4732
R8167 gnd.n6018 gnd.n5890 42.4732
R8168 gnd.n3243 gnd.n3242 42.2793
R8169 gnd.n2740 gnd.n2739 42.2793
R8170 gnd.n3169 gnd.n3168 42.2793
R8171 gnd.n4114 gnd.n2713 42.2793
R8172 gnd.n124 gnd.n123 42.2793
R8173 gnd.n5997 gnd.n5900 42.2793
R8174 gnd.n2451 gnd.n2449 42.2793
R8175 gnd.n1901 gnd.n1900 42.2793
R8176 gnd.n7845 gnd.n202 42.2793
R8177 gnd.n7882 gnd.n7881 42.2793
R8178 gnd.n4180 gnd.n4179 42.2793
R8179 gnd.n4156 gnd.n4155 42.2793
R8180 gnd.n4352 gnd.n4351 42.2793
R8181 gnd.n4822 gnd.n4764 42.2793
R8182 gnd.n1348 gnd.n1347 41.6274
R8183 gnd.n5608 gnd.n5607 41.6274
R8184 gnd.n1357 gnd.n1356 40.8975
R8185 gnd.n5611 gnd.n5610 40.8975
R8186 gnd.n6876 gnd.n6875 37.4155
R8187 gnd.n6875 gnd.n6874 37.4155
R8188 gnd.n6874 gnd.n853 37.4155
R8189 gnd.n6868 gnd.n853 37.4155
R8190 gnd.n6868 gnd.n6867 37.4155
R8191 gnd.n6867 gnd.n6866 37.4155
R8192 gnd.n6866 gnd.n860 37.4155
R8193 gnd.n6860 gnd.n860 37.4155
R8194 gnd.n6860 gnd.n6859 37.4155
R8195 gnd.n6859 gnd.n6858 37.4155
R8196 gnd.n6858 gnd.n868 37.4155
R8197 gnd.n6852 gnd.n868 37.4155
R8198 gnd.n6852 gnd.n6851 37.4155
R8199 gnd.n6851 gnd.n6850 37.4155
R8200 gnd.n6850 gnd.n876 37.4155
R8201 gnd.n6844 gnd.n876 37.4155
R8202 gnd.n6844 gnd.n6843 37.4155
R8203 gnd.n6843 gnd.n6842 37.4155
R8204 gnd.n6842 gnd.n884 37.4155
R8205 gnd.n6836 gnd.n884 37.4155
R8206 gnd.n6836 gnd.n6835 37.4155
R8207 gnd.n6835 gnd.n6834 37.4155
R8208 gnd.n6834 gnd.n892 37.4155
R8209 gnd.n6828 gnd.n892 37.4155
R8210 gnd.n6828 gnd.n6827 37.4155
R8211 gnd.n6827 gnd.n6826 37.4155
R8212 gnd.n6826 gnd.n900 37.4155
R8213 gnd.n6820 gnd.n900 37.4155
R8214 gnd.n6820 gnd.n6819 37.4155
R8215 gnd.n6819 gnd.n6818 37.4155
R8216 gnd.n6818 gnd.n908 37.4155
R8217 gnd.n6812 gnd.n908 37.4155
R8218 gnd.n6812 gnd.n6811 37.4155
R8219 gnd.n6811 gnd.n6810 37.4155
R8220 gnd.n6810 gnd.n916 37.4155
R8221 gnd.n6804 gnd.n916 37.4155
R8222 gnd.n6804 gnd.n6803 37.4155
R8223 gnd.n6803 gnd.n6802 37.4155
R8224 gnd.n6802 gnd.n924 37.4155
R8225 gnd.n6796 gnd.n924 37.4155
R8226 gnd.n6796 gnd.n6795 37.4155
R8227 gnd.n6795 gnd.n6794 37.4155
R8228 gnd.n6794 gnd.n932 37.4155
R8229 gnd.n6788 gnd.n932 37.4155
R8230 gnd.n6788 gnd.n6787 37.4155
R8231 gnd.n6787 gnd.n6786 37.4155
R8232 gnd.n6786 gnd.n940 37.4155
R8233 gnd.n6780 gnd.n940 37.4155
R8234 gnd.n6780 gnd.n6779 37.4155
R8235 gnd.n6779 gnd.n6778 37.4155
R8236 gnd.n6778 gnd.n948 37.4155
R8237 gnd.n6772 gnd.n948 37.4155
R8238 gnd.n6772 gnd.n6771 37.4155
R8239 gnd.n6771 gnd.n6770 37.4155
R8240 gnd.n6770 gnd.n956 37.4155
R8241 gnd.n6764 gnd.n956 37.4155
R8242 gnd.n6764 gnd.n6763 37.4155
R8243 gnd.n6763 gnd.n6762 37.4155
R8244 gnd.n6762 gnd.n964 37.4155
R8245 gnd.n6756 gnd.n964 37.4155
R8246 gnd.n6756 gnd.n6755 37.4155
R8247 gnd.n6755 gnd.n6754 37.4155
R8248 gnd.n6754 gnd.n972 37.4155
R8249 gnd.n6748 gnd.n972 37.4155
R8250 gnd.n6748 gnd.n6747 37.4155
R8251 gnd.n6747 gnd.n6746 37.4155
R8252 gnd.n6746 gnd.n980 37.4155
R8253 gnd.n6740 gnd.n980 37.4155
R8254 gnd.n6740 gnd.n6739 37.4155
R8255 gnd.n6739 gnd.n6738 37.4155
R8256 gnd.n6738 gnd.n988 37.4155
R8257 gnd.n6732 gnd.n988 37.4155
R8258 gnd.n6732 gnd.n6731 37.4155
R8259 gnd.n6731 gnd.n6730 37.4155
R8260 gnd.n6730 gnd.n996 37.4155
R8261 gnd.n6724 gnd.n996 37.4155
R8262 gnd.n6724 gnd.n6723 37.4155
R8263 gnd.n6723 gnd.n6722 37.4155
R8264 gnd.n6722 gnd.n1004 37.4155
R8265 gnd.n6716 gnd.n1004 37.4155
R8266 gnd.n6716 gnd.n6715 37.4155
R8267 gnd.n6715 gnd.n6714 37.4155
R8268 gnd.n6714 gnd.n1012 37.4155
R8269 gnd.n1984 gnd.n1878 36.9518
R8270 gnd.n6548 gnd.n1298 36.9518
R8271 gnd.n1356 gnd.n1355 35.055
R8272 gnd.n1351 gnd.n1350 35.055
R8273 gnd.n5600 gnd.n5599 35.055
R8274 gnd.n5610 gnd.n5596 35.055
R8275 gnd.n3305 gnd.n3199 31.8661
R8276 gnd.n3305 gnd.n3304 31.8661
R8277 gnd.n3313 gnd.n3188 31.8661
R8278 gnd.n3321 gnd.n3188 31.8661
R8279 gnd.n3321 gnd.n3182 31.8661
R8280 gnd.n3329 gnd.n3182 31.8661
R8281 gnd.n3329 gnd.n3175 31.8661
R8282 gnd.n3367 gnd.n3175 31.8661
R8283 gnd.n3377 gnd.n3108 31.8661
R8284 gnd.n4442 gnd.n4325 31.8661
R8285 gnd.n4450 gnd.n2659 31.8661
R8286 gnd.n4458 gnd.n2659 31.8661
R8287 gnd.n4458 gnd.n2651 31.8661
R8288 gnd.n4466 gnd.n2651 31.8661
R8289 gnd.n4474 gnd.n2642 31.8661
R8290 gnd.n4474 gnd.n2645 31.8661
R8291 gnd.n4482 gnd.n2626 31.8661
R8292 gnd.n4500 gnd.n2626 31.8661
R8293 gnd.n4509 gnd.n2618 31.8661
R8294 gnd.n6707 gnd.n1022 31.8661
R8295 gnd.n4922 gnd.n1251 31.8661
R8296 gnd.n4915 gnd.n1262 31.8661
R8297 gnd.n4915 gnd.n2316 31.8661
R8298 gnd.n4974 gnd.n2309 31.8661
R8299 gnd.n4982 gnd.n2309 31.8661
R8300 gnd.n4990 gnd.n2302 31.8661
R8301 gnd.n4990 gnd.n2294 31.8661
R8302 gnd.n4998 gnd.n2294 31.8661
R8303 gnd.n4998 gnd.n2296 31.8661
R8304 gnd.n5006 gnd.n2281 31.8661
R8305 gnd.n5014 gnd.n2281 31.8661
R8306 gnd.n5014 gnd.n2274 31.8661
R8307 gnd.n5022 gnd.n2274 31.8661
R8308 gnd.n5030 gnd.n2267 31.8661
R8309 gnd.n5030 gnd.n2260 31.8661
R8310 gnd.n5038 gnd.n2260 31.8661
R8311 gnd.n5046 gnd.n2253 31.8661
R8312 gnd.n5046 gnd.n2245 31.8661
R8313 gnd.n5054 gnd.n2245 31.8661
R8314 gnd.n5054 gnd.n2247 31.8661
R8315 gnd.n5062 gnd.n2230 31.8661
R8316 gnd.n5081 gnd.n2230 31.8661
R8317 gnd.n5081 gnd.n2222 31.8661
R8318 gnd.n5092 gnd.n2222 31.8661
R8319 gnd.n5765 gnd.n1793 31.8661
R8320 gnd.n5765 gnd.n1787 31.8661
R8321 gnd.n5775 gnd.n1787 31.8661
R8322 gnd.n5775 gnd.n5773 31.8661
R8323 gnd.n5783 gnd.n1776 31.8661
R8324 gnd.n5792 gnd.n1776 31.8661
R8325 gnd.n5792 gnd.n1770 31.8661
R8326 gnd.n5800 gnd.n1770 31.8661
R8327 gnd.n5809 gnd.n1764 31.8661
R8328 gnd.n5809 gnd.n1758 31.8661
R8329 gnd.n5817 gnd.n1758 31.8661
R8330 gnd.n5826 gnd.n1752 31.8661
R8331 gnd.n5826 gnd.n1745 31.8661
R8332 gnd.n5834 gnd.n1745 31.8661
R8333 gnd.n5834 gnd.n1746 31.8661
R8334 gnd.n5843 gnd.n1734 31.8661
R8335 gnd.n5853 gnd.n1734 31.8661
R8336 gnd.n5853 gnd.n1728 31.8661
R8337 gnd.n5862 gnd.n1728 31.8661
R8338 gnd.n6355 gnd.n1472 31.8661
R8339 gnd.n6355 gnd.n1474 31.8661
R8340 gnd.n6030 gnd.n6029 31.8661
R8341 gnd.n6030 gnd.n1690 31.8661
R8342 gnd.n6040 gnd.n1682 31.8661
R8343 gnd.n7711 gnd.n269 31.8661
R8344 gnd.n7727 gnd.n252 31.8661
R8345 gnd.n7735 gnd.n244 31.8661
R8346 gnd.n7735 gnd.n246 31.8661
R8347 gnd.n7743 gnd.n230 31.8661
R8348 gnd.n7751 gnd.n230 31.8661
R8349 gnd.n7759 gnd.n222 31.8661
R8350 gnd.n7759 gnd.n213 31.8661
R8351 gnd.n7769 gnd.n213 31.8661
R8352 gnd.n7769 gnd.n215 31.8661
R8353 gnd.t66 gnd.n2618 30.2728
R8354 gnd.n7727 gnd.t25 30.2728
R8355 gnd.n5690 gnd.n1988 30.1273
R8356 gnd.n5177 gnd.n5173 30.1273
R8357 gnd.n4325 gnd.t230 28.3609
R8358 gnd.n7838 gnd.t157 28.3609
R8359 gnd.n5038 gnd.t318 27.0862
R8360 gnd.t341 gnd.n1764 27.0862
R8361 gnd.n7917 gnd.n126 25.8116
R8362 gnd.n4845 gnd.n4844 25.7944
R8363 gnd.n3168 gnd.n3167 25.7944
R8364 gnd.n2713 gnd.n2712 25.7944
R8365 gnd.n123 gnd.n122 25.7944
R8366 gnd.n5900 gnd.n5899 25.7944
R8367 gnd.n2449 gnd.n2448 25.7944
R8368 gnd.n1878 gnd.n1877 25.7944
R8369 gnd.n1900 gnd.n1899 25.7944
R8370 gnd.n202 gnd.n201 25.7944
R8371 gnd.n7881 gnd.n7880 25.7944
R8372 gnd.n4179 gnd.n4178 25.7944
R8373 gnd.n4155 gnd.n4154 25.7944
R8374 gnd.n4351 gnd.n4350 25.7944
R8375 gnd.n4764 gnd.n4763 25.7944
R8376 gnd.n1298 gnd.n1297 25.7944
R8377 gnd.n5890 gnd.n5889 25.7944
R8378 gnd.n6544 gnd.n1336 25.1743
R8379 gnd.n5757 gnd.n5755 25.1743
R8380 gnd.n3389 gnd.n3109 24.8557
R8381 gnd.n3399 gnd.n3092 24.8557
R8382 gnd.n3095 gnd.n3083 24.8557
R8383 gnd.n3420 gnd.n3084 24.8557
R8384 gnd.n3430 gnd.n3064 24.8557
R8385 gnd.n3440 gnd.n3439 24.8557
R8386 gnd.n3050 gnd.n3048 24.8557
R8387 gnd.n3471 gnd.n3470 24.8557
R8388 gnd.n3486 gnd.n3033 24.8557
R8389 gnd.n3540 gnd.n2972 24.8557
R8390 gnd.n3496 gnd.n2973 24.8557
R8391 gnd.n3533 gnd.n2984 24.8557
R8392 gnd.n3022 gnd.n3021 24.8557
R8393 gnd.n3527 gnd.n3526 24.8557
R8394 gnd.n3008 gnd.n2995 24.8557
R8395 gnd.n3566 gnd.n3565 24.8557
R8396 gnd.n3576 gnd.n2892 24.8557
R8397 gnd.n3588 gnd.n2884 24.8557
R8398 gnd.n3587 gnd.n2872 24.8557
R8399 gnd.n3606 gnd.n3605 24.8557
R8400 gnd.n3616 gnd.n2865 24.8557
R8401 gnd.n3627 gnd.n2853 24.8557
R8402 gnd.n3651 gnd.n3650 24.8557
R8403 gnd.n3662 gnd.n2836 24.8557
R8404 gnd.n3661 gnd.n2838 24.8557
R8405 gnd.n3673 gnd.n2829 24.8557
R8406 gnd.n3691 gnd.n3690 24.8557
R8407 gnd.n2820 gnd.n2809 24.8557
R8408 gnd.n3712 gnd.n2797 24.8557
R8409 gnd.n3740 gnd.n3739 24.8557
R8410 gnd.n3751 gnd.n2781 24.8557
R8411 gnd.n3762 gnd.n2774 24.8557
R8412 gnd.n3761 gnd.n2762 24.8557
R8413 gnd.n4034 gnd.n4033 24.8557
R8414 gnd.n4056 gnd.n2747 24.8557
R8415 gnd.n4982 gnd.t193 24.537
R8416 gnd.t35 gnd.n2267 24.537
R8417 gnd.n5817 gnd.t92 24.537
R8418 gnd.t165 gnd.n1472 24.537
R8419 gnd.n4521 gnd.n1035 24.2183
R8420 gnd.n6695 gnd.n1044 24.2183
R8421 gnd.n4529 gnd.n2609 24.2183
R8422 gnd.n6689 gnd.n1054 24.2183
R8423 gnd.n6683 gnd.n1065 24.2183
R8424 gnd.n4551 gnd.n1068 24.2183
R8425 gnd.n4569 gnd.n1078 24.2183
R8426 gnd.n6671 gnd.n1086 24.2183
R8427 gnd.n4563 gnd.n4562 24.2183
R8428 gnd.n4590 gnd.n2551 24.2183
R8429 gnd.n4598 gnd.n4597 24.2183
R8430 gnd.n4616 gnd.n2542 24.2183
R8431 gnd.n4625 gnd.n2534 24.2183
R8432 gnd.n6663 gnd.n1101 24.2183
R8433 gnd.n4676 gnd.n1104 24.2183
R8434 gnd.n4646 gnd.n1115 24.2183
R8435 gnd.n6651 gnd.n1122 24.2183
R8436 gnd.n6645 gnd.n1133 24.2183
R8437 gnd.n6639 gnd.n1144 24.2183
R8438 gnd.n4713 gnd.n1147 24.2183
R8439 gnd.n4721 gnd.n1157 24.2183
R8440 gnd.n6627 gnd.n1165 24.2183
R8441 gnd.n6621 gnd.n1176 24.2183
R8442 gnd.n6615 gnd.n1187 24.2183
R8443 gnd.n4888 gnd.n1190 24.2183
R8444 gnd.n4745 gnd.n1200 24.2183
R8445 gnd.n6603 gnd.n1208 24.2183
R8446 gnd.n6597 gnd.n1219 24.2183
R8447 gnd.n4755 gnd.n1222 24.2183
R8448 gnd.n6591 gnd.n1230 24.2183
R8449 gnd.n4831 gnd.n1233 24.2183
R8450 gnd.n6585 gnd.n1241 24.2183
R8451 gnd.n4923 gnd.n1244 24.2183
R8452 gnd.n6052 gnd.n1684 24.2183
R8453 gnd.n6062 gnd.n1675 24.2183
R8454 gnd.n6061 gnd.n1665 24.2183
R8455 gnd.n6074 gnd.n6072 24.2183
R8456 gnd.n1668 gnd.n1656 24.2183
R8457 gnd.n6084 gnd.n1658 24.2183
R8458 gnd.n6094 gnd.n1639 24.2183
R8459 gnd.n6106 gnd.n6105 24.2183
R8460 gnd.n6116 gnd.n1632 24.2183
R8461 gnd.n6126 gnd.n1622 24.2183
R8462 gnd.n6144 gnd.n6143 24.2183
R8463 gnd.n6154 gnd.n1602 24.2183
R8464 gnd.n1605 gnd.n1593 24.2183
R8465 gnd.n6212 gnd.n6211 24.2183
R8466 gnd.n1578 gnd.n1567 24.2183
R8467 gnd.n6204 gnd.n1558 24.2183
R8468 gnd.n6243 gnd.n1549 24.2183
R8469 gnd.n6242 gnd.n1552 24.2183
R8470 gnd.n6302 gnd.n1515 24.2183
R8471 gnd.n6305 gnd.n1518 24.2183
R8472 gnd.n7663 gnd.n323 24.2183
R8473 gnd.n6290 gnd.n1533 24.2183
R8474 gnd.n6285 gnd.n6284 24.2183
R8475 gnd.n7644 gnd.n335 24.2183
R8476 gnd.n7649 gnd.n337 24.2183
R8477 gnd.n7638 gnd.n306 24.2183
R8478 gnd.n7671 gnd.n308 24.2183
R8479 gnd.n7679 gnd.n300 24.2183
R8480 gnd.n7629 gnd.n291 24.2183
R8481 gnd.n7624 gnd.n283 24.2183
R8482 gnd.n7695 gnd.n285 24.2183
R8483 gnd.n398 gnd.n275 24.2183
R8484 gnd.n7703 gnd.n277 24.2183
R8485 gnd.n2537 gnd.t52 23.8997
R8486 gnd.n4974 gnd.n4973 23.8997
R8487 gnd.n6028 gnd.n1474 23.8997
R8488 gnd.t89 gnd.n320 23.8997
R8489 gnd.n3410 gnd.t288 23.2624
R8490 gnd.n4466 gnd.t50 23.2624
R8491 gnd.t16 gnd.n1136 23.2624
R8492 gnd.n4751 gnd.t44 23.2624
R8493 gnd.n1931 gnd.t37 23.2624
R8494 gnd.n6205 gnd.t6 23.2624
R8495 gnd.t114 gnd.n222 23.2624
R8496 gnd.n3111 gnd.t243 22.6251
R8497 gnd.n4509 gnd.t143 22.6251
R8498 gnd.n4729 gnd.t147 22.6251
R8499 gnd.t27 gnd.n1179 22.6251
R8500 gnd.t4 gnd.n1611 22.6251
R8501 gnd.n1614 gnd.t131 22.6251
R8502 gnd.t14 gnd.n252 22.6251
R8503 gnd.n2789 gnd.n1012 22.4495
R8504 gnd.n4650 gnd.t74 21.9878
R8505 gnd.n6232 gnd.t86 21.9878
R8506 gnd.n6474 gnd.n6473 21.6691
R8507 gnd.n5257 gnd.n5256 21.6691
R8508 gnd.n5273 gnd.n2192 21.6691
R8509 gnd.n5280 gnd.n2182 21.6691
R8510 gnd.n5298 gnd.n5297 21.6691
R8511 gnd.n5314 gnd.n2160 21.6691
R8512 gnd.n5403 gnd.n2114 21.6691
R8513 gnd.n5460 gnd.n2071 21.6691
R8514 gnd.n5514 gnd.n2042 21.6691
R8515 gnd.n5522 gnd.n5521 21.6691
R8516 gnd.n5540 gnd.n2028 21.6691
R8517 gnd.n5549 gnd.n2023 21.6691
R8518 gnd.n5686 gnd.n1991 21.6691
R8519 gnd.t306 gnd.n3116 21.3504
R8520 gnd.n4630 gnd.t29 21.3504
R8521 gnd.n6186 gnd.t139 21.3504
R8522 gnd.t39 gnd.n2810 20.7131
R8523 gnd.n6677 gnd.t18 20.7131
R8524 gnd.n7633 gnd.t60 20.7131
R8525 gnd.n5175 gnd.n1362 20.3945
R8526 gnd.t316 gnd.n2845 20.0758
R8527 gnd.n6708 gnd.n6707 20.0758
R8528 gnd.n6701 gnd.t119 20.0758
R8529 gnd.n5566 gnd.t339 20.0758
R8530 gnd.n393 gnd.t129 20.0758
R8531 gnd.n269 gnd.n259 20.0758
R8532 gnd.n5111 gnd.n5110 19.9763
R8533 gnd.n1987 gnd.n1986 19.9763
R8534 gnd.n6480 gnd.n6479 19.9763
R8535 gnd.n5615 gnd.n5614 19.9763
R8536 gnd.n1344 gnd.t257 19.8005
R8537 gnd.n1344 gnd.t215 19.8005
R8538 gnd.n1345 gnd.t155 19.8005
R8539 gnd.n1345 gnd.t202 19.8005
R8540 gnd.n5604 gnd.t212 19.8005
R8541 gnd.n5604 gnd.t241 19.8005
R8542 gnd.n5605 gnd.t174 19.8005
R8543 gnd.n5605 gnd.t228 19.8005
R8544 gnd.n6577 gnd.n1262 19.7572
R8545 gnd.t256 gnd.n2212 19.7572
R8546 gnd.n6041 gnd.n1690 19.7572
R8547 gnd.n1341 gnd.n1340 19.5087
R8548 gnd.n1354 gnd.n1341 19.5087
R8549 gnd.n1352 gnd.n1343 19.5087
R8550 gnd.n5609 gnd.n5603 19.5087
R8551 gnd.n3577 gnd.t21 19.4385
R8552 gnd.n4482 gnd.t33 19.4385
R8553 gnd.n2296 gnd.t354 19.4385
R8554 gnd.n5843 gnd.t149 19.4385
R8555 gnd.n246 gnd.t117 19.4385
R8556 gnd.n4984 gnd.n2307 19.3944
R8557 gnd.n4984 gnd.n2305 19.3944
R8558 gnd.n4988 gnd.n2305 19.3944
R8559 gnd.n4988 gnd.n2292 19.3944
R8560 gnd.n5000 gnd.n2292 19.3944
R8561 gnd.n5000 gnd.n2290 19.3944
R8562 gnd.n5004 gnd.n2290 19.3944
R8563 gnd.n5004 gnd.n2279 19.3944
R8564 gnd.n5016 gnd.n2279 19.3944
R8565 gnd.n5016 gnd.n2277 19.3944
R8566 gnd.n5020 gnd.n2277 19.3944
R8567 gnd.n5020 gnd.n2265 19.3944
R8568 gnd.n5032 gnd.n2265 19.3944
R8569 gnd.n5032 gnd.n2263 19.3944
R8570 gnd.n5036 gnd.n2263 19.3944
R8571 gnd.n5036 gnd.n2251 19.3944
R8572 gnd.n5048 gnd.n2251 19.3944
R8573 gnd.n5048 gnd.n2249 19.3944
R8574 gnd.n5052 gnd.n2249 19.3944
R8575 gnd.n5052 gnd.n2237 19.3944
R8576 gnd.n5064 gnd.n2237 19.3944
R8577 gnd.n5064 gnd.n2234 19.3944
R8578 gnd.n5079 gnd.n2234 19.3944
R8579 gnd.n5079 gnd.n2235 19.3944
R8580 gnd.n5075 gnd.n2235 19.3944
R8581 gnd.n5075 gnd.n5074 19.3944
R8582 gnd.n5074 gnd.n5073 19.3944
R8583 gnd.n5073 gnd.n5070 19.3944
R8584 gnd.n5070 gnd.n1381 19.3944
R8585 gnd.n6464 gnd.n1381 19.3944
R8586 gnd.n6464 gnd.n1382 19.3944
R8587 gnd.n6460 gnd.n1382 19.3944
R8588 gnd.n6460 gnd.n6459 19.3944
R8589 gnd.n6459 gnd.n6458 19.3944
R8590 gnd.n6458 gnd.n1388 19.3944
R8591 gnd.n6454 gnd.n1388 19.3944
R8592 gnd.n6454 gnd.n6453 19.3944
R8593 gnd.n6453 gnd.n6452 19.3944
R8594 gnd.n6452 gnd.n1393 19.3944
R8595 gnd.n6448 gnd.n1393 19.3944
R8596 gnd.n6448 gnd.n6447 19.3944
R8597 gnd.n6447 gnd.n6446 19.3944
R8598 gnd.n6446 gnd.n1398 19.3944
R8599 gnd.n6442 gnd.n1398 19.3944
R8600 gnd.n6442 gnd.n6441 19.3944
R8601 gnd.n6441 gnd.n6440 19.3944
R8602 gnd.n6440 gnd.n1403 19.3944
R8603 gnd.n6436 gnd.n1403 19.3944
R8604 gnd.n6436 gnd.n6435 19.3944
R8605 gnd.n6435 gnd.n6434 19.3944
R8606 gnd.n6434 gnd.n1408 19.3944
R8607 gnd.n6430 gnd.n1408 19.3944
R8608 gnd.n6430 gnd.n6429 19.3944
R8609 gnd.n6429 gnd.n6428 19.3944
R8610 gnd.n6428 gnd.n1413 19.3944
R8611 gnd.n6424 gnd.n1413 19.3944
R8612 gnd.n6424 gnd.n6423 19.3944
R8613 gnd.n6423 gnd.n6422 19.3944
R8614 gnd.n6422 gnd.n1418 19.3944
R8615 gnd.n6418 gnd.n1418 19.3944
R8616 gnd.n6418 gnd.n6417 19.3944
R8617 gnd.n6417 gnd.n6416 19.3944
R8618 gnd.n6416 gnd.n1423 19.3944
R8619 gnd.n6412 gnd.n1423 19.3944
R8620 gnd.n6412 gnd.n6411 19.3944
R8621 gnd.n6411 gnd.n6410 19.3944
R8622 gnd.n6410 gnd.n1428 19.3944
R8623 gnd.n6406 gnd.n1428 19.3944
R8624 gnd.n6406 gnd.n6405 19.3944
R8625 gnd.n6405 gnd.n6404 19.3944
R8626 gnd.n6404 gnd.n1433 19.3944
R8627 gnd.n6400 gnd.n1433 19.3944
R8628 gnd.n6400 gnd.n6399 19.3944
R8629 gnd.n6399 gnd.n6398 19.3944
R8630 gnd.n6398 gnd.n1438 19.3944
R8631 gnd.n6394 gnd.n1438 19.3944
R8632 gnd.n6394 gnd.n6393 19.3944
R8633 gnd.n6393 gnd.n6392 19.3944
R8634 gnd.n6392 gnd.n1443 19.3944
R8635 gnd.n6388 gnd.n1443 19.3944
R8636 gnd.n6388 gnd.n6387 19.3944
R8637 gnd.n6387 gnd.n6386 19.3944
R8638 gnd.n6386 gnd.n1448 19.3944
R8639 gnd.n6382 gnd.n1448 19.3944
R8640 gnd.n6382 gnd.n6381 19.3944
R8641 gnd.n6381 gnd.n6380 19.3944
R8642 gnd.n6380 gnd.n1453 19.3944
R8643 gnd.n6376 gnd.n1453 19.3944
R8644 gnd.n6376 gnd.n6375 19.3944
R8645 gnd.n6375 gnd.n6374 19.3944
R8646 gnd.n6374 gnd.n1458 19.3944
R8647 gnd.n6370 gnd.n1458 19.3944
R8648 gnd.n6370 gnd.n6369 19.3944
R8649 gnd.n6369 gnd.n6368 19.3944
R8650 gnd.n6368 gnd.n1463 19.3944
R8651 gnd.n6364 gnd.n1463 19.3944
R8652 gnd.n6364 gnd.n6363 19.3944
R8653 gnd.n6363 gnd.n6362 19.3944
R8654 gnd.n6362 gnd.n1468 19.3944
R8655 gnd.n6358 gnd.n1468 19.3944
R8656 gnd.n6358 gnd.n6357 19.3944
R8657 gnd.n4857 gnd.n4856 19.3944
R8658 gnd.n4856 gnd.n4855 19.3944
R8659 gnd.n4855 gnd.n4852 19.3944
R8660 gnd.n4970 gnd.n4969 19.3944
R8661 gnd.n4969 gnd.n2334 19.3944
R8662 gnd.n4962 gnd.n2334 19.3944
R8663 gnd.n4962 gnd.n4961 19.3944
R8664 gnd.n4961 gnd.n2415 19.3944
R8665 gnd.n4954 gnd.n2415 19.3944
R8666 gnd.n4954 gnd.n4953 19.3944
R8667 gnd.n4953 gnd.n2423 19.3944
R8668 gnd.n4946 gnd.n2423 19.3944
R8669 gnd.n4946 gnd.n4945 19.3944
R8670 gnd.n4945 gnd.n2435 19.3944
R8671 gnd.n4938 gnd.n2435 19.3944
R8672 gnd.n4938 gnd.n4937 19.3944
R8673 gnd.n4937 gnd.n2443 19.3944
R8674 gnd.n4930 gnd.n2443 19.3944
R8675 gnd.n4930 gnd.n4929 19.3944
R8676 gnd.n4929 gnd.n2457 19.3944
R8677 gnd.n4868 gnd.n2457 19.3944
R8678 gnd.n4868 gnd.n4867 19.3944
R8679 gnd.n4867 gnd.n4866 19.3944
R8680 gnd.n4866 gnd.n4839 19.3944
R8681 gnd.n4862 gnd.n4839 19.3944
R8682 gnd.n4862 gnd.n4861 19.3944
R8683 gnd.n4861 gnd.n4860 19.3944
R8684 gnd.n3292 gnd.n3291 19.3944
R8685 gnd.n3291 gnd.n3290 19.3944
R8686 gnd.n3290 gnd.n3289 19.3944
R8687 gnd.n3289 gnd.n3287 19.3944
R8688 gnd.n3287 gnd.n3284 19.3944
R8689 gnd.n3284 gnd.n3283 19.3944
R8690 gnd.n3283 gnd.n3280 19.3944
R8691 gnd.n3280 gnd.n3279 19.3944
R8692 gnd.n3279 gnd.n3276 19.3944
R8693 gnd.n3276 gnd.n3275 19.3944
R8694 gnd.n3275 gnd.n3272 19.3944
R8695 gnd.n3272 gnd.n3271 19.3944
R8696 gnd.n3271 gnd.n3268 19.3944
R8697 gnd.n3268 gnd.n3267 19.3944
R8698 gnd.n3267 gnd.n3264 19.3944
R8699 gnd.n3264 gnd.n3263 19.3944
R8700 gnd.n3263 gnd.n3260 19.3944
R8701 gnd.n3260 gnd.n3259 19.3944
R8702 gnd.n3259 gnd.n3256 19.3944
R8703 gnd.n3256 gnd.n3255 19.3944
R8704 gnd.n3255 gnd.n3252 19.3944
R8705 gnd.n3252 gnd.n3251 19.3944
R8706 gnd.n3248 gnd.n3247 19.3944
R8707 gnd.n3247 gnd.n3203 19.3944
R8708 gnd.n3298 gnd.n3203 19.3944
R8709 gnd.n4064 gnd.n4063 19.3944
R8710 gnd.n4063 gnd.n4060 19.3944
R8711 gnd.n4060 gnd.n4059 19.3944
R8712 gnd.n4109 gnd.n4108 19.3944
R8713 gnd.n4108 gnd.n4107 19.3944
R8714 gnd.n4107 gnd.n4104 19.3944
R8715 gnd.n4104 gnd.n4103 19.3944
R8716 gnd.n4103 gnd.n4100 19.3944
R8717 gnd.n4100 gnd.n4099 19.3944
R8718 gnd.n4099 gnd.n4096 19.3944
R8719 gnd.n4096 gnd.n4095 19.3944
R8720 gnd.n4095 gnd.n4092 19.3944
R8721 gnd.n4092 gnd.n4091 19.3944
R8722 gnd.n4091 gnd.n4088 19.3944
R8723 gnd.n4088 gnd.n4087 19.3944
R8724 gnd.n4087 gnd.n4084 19.3944
R8725 gnd.n4084 gnd.n4083 19.3944
R8726 gnd.n4083 gnd.n4080 19.3944
R8727 gnd.n4080 gnd.n4079 19.3944
R8728 gnd.n4079 gnd.n4076 19.3944
R8729 gnd.n4076 gnd.n4075 19.3944
R8730 gnd.n4075 gnd.n4072 19.3944
R8731 gnd.n4072 gnd.n4071 19.3944
R8732 gnd.n4071 gnd.n4068 19.3944
R8733 gnd.n4068 gnd.n4067 19.3944
R8734 gnd.n3391 gnd.n3100 19.3944
R8735 gnd.n3401 gnd.n3100 19.3944
R8736 gnd.n3402 gnd.n3401 19.3944
R8737 gnd.n3402 gnd.n3081 19.3944
R8738 gnd.n3422 gnd.n3081 19.3944
R8739 gnd.n3422 gnd.n3073 19.3944
R8740 gnd.n3432 gnd.n3073 19.3944
R8741 gnd.n3433 gnd.n3432 19.3944
R8742 gnd.n3434 gnd.n3433 19.3944
R8743 gnd.n3434 gnd.n3056 19.3944
R8744 gnd.n3451 gnd.n3056 19.3944
R8745 gnd.n3454 gnd.n3451 19.3944
R8746 gnd.n3454 gnd.n3453 19.3944
R8747 gnd.n3453 gnd.n3029 19.3944
R8748 gnd.n3493 gnd.n3029 19.3944
R8749 gnd.n3493 gnd.n3026 19.3944
R8750 gnd.n3499 gnd.n3026 19.3944
R8751 gnd.n3500 gnd.n3499 19.3944
R8752 gnd.n3500 gnd.n3024 19.3944
R8753 gnd.n3506 gnd.n3024 19.3944
R8754 gnd.n3509 gnd.n3506 19.3944
R8755 gnd.n3511 gnd.n3509 19.3944
R8756 gnd.n3517 gnd.n3511 19.3944
R8757 gnd.n3517 gnd.n3516 19.3944
R8758 gnd.n3516 gnd.n2887 19.3944
R8759 gnd.n3583 gnd.n2887 19.3944
R8760 gnd.n3584 gnd.n3583 19.3944
R8761 gnd.n3584 gnd.n2880 19.3944
R8762 gnd.n3595 gnd.n2880 19.3944
R8763 gnd.n3596 gnd.n3595 19.3944
R8764 gnd.n3596 gnd.n2863 19.3944
R8765 gnd.n2863 gnd.n2861 19.3944
R8766 gnd.n3620 gnd.n2861 19.3944
R8767 gnd.n3621 gnd.n3620 19.3944
R8768 gnd.n3621 gnd.n2832 19.3944
R8769 gnd.n3668 gnd.n2832 19.3944
R8770 gnd.n3669 gnd.n3668 19.3944
R8771 gnd.n3669 gnd.n2825 19.3944
R8772 gnd.n3680 gnd.n2825 19.3944
R8773 gnd.n3681 gnd.n3680 19.3944
R8774 gnd.n3681 gnd.n2808 19.3944
R8775 gnd.n2808 gnd.n2806 19.3944
R8776 gnd.n3705 gnd.n2806 19.3944
R8777 gnd.n3706 gnd.n3705 19.3944
R8778 gnd.n3706 gnd.n2777 19.3944
R8779 gnd.n3757 gnd.n2777 19.3944
R8780 gnd.n3758 gnd.n3757 19.3944
R8781 gnd.n3758 gnd.n2770 19.3944
R8782 gnd.n4025 gnd.n2770 19.3944
R8783 gnd.n4026 gnd.n4025 19.3944
R8784 gnd.n4026 gnd.n2751 19.3944
R8785 gnd.n4051 gnd.n2751 19.3944
R8786 gnd.n4051 gnd.n2752 19.3944
R8787 gnd.n3382 gnd.n3381 19.3944
R8788 gnd.n3381 gnd.n3114 19.3944
R8789 gnd.n3137 gnd.n3114 19.3944
R8790 gnd.n3140 gnd.n3137 19.3944
R8791 gnd.n3140 gnd.n3133 19.3944
R8792 gnd.n3144 gnd.n3133 19.3944
R8793 gnd.n3147 gnd.n3144 19.3944
R8794 gnd.n3150 gnd.n3147 19.3944
R8795 gnd.n3150 gnd.n3131 19.3944
R8796 gnd.n3154 gnd.n3131 19.3944
R8797 gnd.n3157 gnd.n3154 19.3944
R8798 gnd.n3160 gnd.n3157 19.3944
R8799 gnd.n3160 gnd.n3129 19.3944
R8800 gnd.n3164 gnd.n3129 19.3944
R8801 gnd.n3387 gnd.n3386 19.3944
R8802 gnd.n3386 gnd.n3090 19.3944
R8803 gnd.n3412 gnd.n3090 19.3944
R8804 gnd.n3412 gnd.n3088 19.3944
R8805 gnd.n3418 gnd.n3088 19.3944
R8806 gnd.n3418 gnd.n3417 19.3944
R8807 gnd.n3417 gnd.n3062 19.3944
R8808 gnd.n3442 gnd.n3062 19.3944
R8809 gnd.n3442 gnd.n3060 19.3944
R8810 gnd.n3446 gnd.n3060 19.3944
R8811 gnd.n3446 gnd.n3040 19.3944
R8812 gnd.n3473 gnd.n3040 19.3944
R8813 gnd.n3473 gnd.n3038 19.3944
R8814 gnd.n3483 gnd.n3038 19.3944
R8815 gnd.n3483 gnd.n3482 19.3944
R8816 gnd.n3482 gnd.n3481 19.3944
R8817 gnd.n3481 gnd.n2987 19.3944
R8818 gnd.n3531 gnd.n2987 19.3944
R8819 gnd.n3531 gnd.n3530 19.3944
R8820 gnd.n3530 gnd.n3529 19.3944
R8821 gnd.n3529 gnd.n2991 19.3944
R8822 gnd.n3011 gnd.n2991 19.3944
R8823 gnd.n3011 gnd.n2897 19.3944
R8824 gnd.n3568 gnd.n2897 19.3944
R8825 gnd.n3568 gnd.n2895 19.3944
R8826 gnd.n3574 gnd.n2895 19.3944
R8827 gnd.n3574 gnd.n3573 19.3944
R8828 gnd.n3573 gnd.n2870 19.3944
R8829 gnd.n3608 gnd.n2870 19.3944
R8830 gnd.n3608 gnd.n2868 19.3944
R8831 gnd.n3614 gnd.n2868 19.3944
R8832 gnd.n3614 gnd.n3613 19.3944
R8833 gnd.n3613 gnd.n2843 19.3944
R8834 gnd.n3653 gnd.n2843 19.3944
R8835 gnd.n3653 gnd.n2841 19.3944
R8836 gnd.n3659 gnd.n2841 19.3944
R8837 gnd.n3659 gnd.n3658 19.3944
R8838 gnd.n3658 gnd.n2815 19.3944
R8839 gnd.n3693 gnd.n2815 19.3944
R8840 gnd.n3693 gnd.n2813 19.3944
R8841 gnd.n3699 gnd.n2813 19.3944
R8842 gnd.n3699 gnd.n3698 19.3944
R8843 gnd.n3698 gnd.n2787 19.3944
R8844 gnd.n3742 gnd.n2787 19.3944
R8845 gnd.n3742 gnd.n2785 19.3944
R8846 gnd.n3748 gnd.n2785 19.3944
R8847 gnd.n3748 gnd.n3747 19.3944
R8848 gnd.n3747 gnd.n2760 19.3944
R8849 gnd.n4036 gnd.n2760 19.3944
R8850 gnd.n4036 gnd.n2758 19.3944
R8851 gnd.n4044 gnd.n2758 19.3944
R8852 gnd.n4044 gnd.n4043 19.3944
R8853 gnd.n4043 gnd.n4042 19.3944
R8854 gnd.n4145 gnd.n4144 19.3944
R8855 gnd.n4144 gnd.n2699 19.3944
R8856 gnd.n4140 gnd.n2699 19.3944
R8857 gnd.n4140 gnd.n4137 19.3944
R8858 gnd.n4137 gnd.n4134 19.3944
R8859 gnd.n4134 gnd.n4133 19.3944
R8860 gnd.n4133 gnd.n4130 19.3944
R8861 gnd.n4130 gnd.n4129 19.3944
R8862 gnd.n4129 gnd.n4126 19.3944
R8863 gnd.n4126 gnd.n4125 19.3944
R8864 gnd.n4125 gnd.n4122 19.3944
R8865 gnd.n4122 gnd.n4121 19.3944
R8866 gnd.n4121 gnd.n4118 19.3944
R8867 gnd.n4118 gnd.n4117 19.3944
R8868 gnd.n3302 gnd.n3201 19.3944
R8869 gnd.n3302 gnd.n3192 19.3944
R8870 gnd.n3315 gnd.n3192 19.3944
R8871 gnd.n3315 gnd.n3190 19.3944
R8872 gnd.n3319 gnd.n3190 19.3944
R8873 gnd.n3319 gnd.n3180 19.3944
R8874 gnd.n3331 gnd.n3180 19.3944
R8875 gnd.n3331 gnd.n3178 19.3944
R8876 gnd.n3365 gnd.n3178 19.3944
R8877 gnd.n3365 gnd.n3364 19.3944
R8878 gnd.n3364 gnd.n3363 19.3944
R8879 gnd.n3363 gnd.n3362 19.3944
R8880 gnd.n3362 gnd.n3359 19.3944
R8881 gnd.n3359 gnd.n3358 19.3944
R8882 gnd.n3358 gnd.n3357 19.3944
R8883 gnd.n3357 gnd.n3355 19.3944
R8884 gnd.n3355 gnd.n3354 19.3944
R8885 gnd.n3354 gnd.n3351 19.3944
R8886 gnd.n3351 gnd.n3350 19.3944
R8887 gnd.n3350 gnd.n3349 19.3944
R8888 gnd.n3349 gnd.n3347 19.3944
R8889 gnd.n3347 gnd.n3046 19.3944
R8890 gnd.n3462 gnd.n3046 19.3944
R8891 gnd.n3462 gnd.n3044 19.3944
R8892 gnd.n3468 gnd.n3044 19.3944
R8893 gnd.n3468 gnd.n3467 19.3944
R8894 gnd.n3467 gnd.n2968 19.3944
R8895 gnd.n3542 gnd.n2968 19.3944
R8896 gnd.n3542 gnd.n2969 19.3944
R8897 gnd.n3016 gnd.n3015 19.3944
R8898 gnd.n3019 gnd.n3018 19.3944
R8899 gnd.n3006 gnd.n3005 19.3944
R8900 gnd.n3561 gnd.n2902 19.3944
R8901 gnd.n3561 gnd.n3560 19.3944
R8902 gnd.n3560 gnd.n3559 19.3944
R8903 gnd.n3559 gnd.n3557 19.3944
R8904 gnd.n3557 gnd.n3556 19.3944
R8905 gnd.n3556 gnd.n3554 19.3944
R8906 gnd.n3554 gnd.n3553 19.3944
R8907 gnd.n3553 gnd.n2851 19.3944
R8908 gnd.n3629 gnd.n2851 19.3944
R8909 gnd.n3629 gnd.n2849 19.3944
R8910 gnd.n3648 gnd.n2849 19.3944
R8911 gnd.n3648 gnd.n3647 19.3944
R8912 gnd.n3647 gnd.n3646 19.3944
R8913 gnd.n3646 gnd.n3644 19.3944
R8914 gnd.n3644 gnd.n3643 19.3944
R8915 gnd.n3643 gnd.n3641 19.3944
R8916 gnd.n3641 gnd.n3640 19.3944
R8917 gnd.n3640 gnd.n2795 19.3944
R8918 gnd.n3714 gnd.n2795 19.3944
R8919 gnd.n3714 gnd.n2793 19.3944
R8920 gnd.n3737 gnd.n2793 19.3944
R8921 gnd.n3737 gnd.n3736 19.3944
R8922 gnd.n3736 gnd.n3735 19.3944
R8923 gnd.n3735 gnd.n3732 19.3944
R8924 gnd.n3732 gnd.n3731 19.3944
R8925 gnd.n3731 gnd.n3729 19.3944
R8926 gnd.n3729 gnd.n3728 19.3944
R8927 gnd.n3728 gnd.n3726 19.3944
R8928 gnd.n3726 gnd.n2746 19.3944
R8929 gnd.n3307 gnd.n3197 19.3944
R8930 gnd.n3307 gnd.n3195 19.3944
R8931 gnd.n3311 gnd.n3195 19.3944
R8932 gnd.n3311 gnd.n3186 19.3944
R8933 gnd.n3323 gnd.n3186 19.3944
R8934 gnd.n3323 gnd.n3184 19.3944
R8935 gnd.n3327 gnd.n3184 19.3944
R8936 gnd.n3327 gnd.n3173 19.3944
R8937 gnd.n3369 gnd.n3173 19.3944
R8938 gnd.n3369 gnd.n3127 19.3944
R8939 gnd.n3375 gnd.n3127 19.3944
R8940 gnd.n3375 gnd.n3374 19.3944
R8941 gnd.n3374 gnd.n3105 19.3944
R8942 gnd.n3396 gnd.n3105 19.3944
R8943 gnd.n3396 gnd.n3098 19.3944
R8944 gnd.n3407 gnd.n3098 19.3944
R8945 gnd.n3407 gnd.n3406 19.3944
R8946 gnd.n3406 gnd.n3079 19.3944
R8947 gnd.n3427 gnd.n3079 19.3944
R8948 gnd.n3427 gnd.n3069 19.3944
R8949 gnd.n3437 gnd.n3069 19.3944
R8950 gnd.n3437 gnd.n3052 19.3944
R8951 gnd.n3458 gnd.n3052 19.3944
R8952 gnd.n3458 gnd.n3457 19.3944
R8953 gnd.n3457 gnd.n3031 19.3944
R8954 gnd.n3488 gnd.n3031 19.3944
R8955 gnd.n3488 gnd.n2976 19.3944
R8956 gnd.n3538 gnd.n2976 19.3944
R8957 gnd.n3538 gnd.n3537 19.3944
R8958 gnd.n3537 gnd.n3536 19.3944
R8959 gnd.n3536 gnd.n2980 19.3944
R8960 gnd.n2998 gnd.n2980 19.3944
R8961 gnd.n3524 gnd.n2998 19.3944
R8962 gnd.n3524 gnd.n3523 19.3944
R8963 gnd.n3523 gnd.n3522 19.3944
R8964 gnd.n3522 gnd.n3002 19.3944
R8965 gnd.n3002 gnd.n2889 19.3944
R8966 gnd.n3579 gnd.n2889 19.3944
R8967 gnd.n3579 gnd.n2882 19.3944
R8968 gnd.n3590 gnd.n2882 19.3944
R8969 gnd.n3590 gnd.n2878 19.3944
R8970 gnd.n3603 gnd.n2878 19.3944
R8971 gnd.n3603 gnd.n3602 19.3944
R8972 gnd.n3602 gnd.n2857 19.3944
R8973 gnd.n3625 gnd.n2857 19.3944
R8974 gnd.n3625 gnd.n3624 19.3944
R8975 gnd.n3624 gnd.n2834 19.3944
R8976 gnd.n3664 gnd.n2834 19.3944
R8977 gnd.n3664 gnd.n2827 19.3944
R8978 gnd.n3675 gnd.n2827 19.3944
R8979 gnd.n3675 gnd.n2823 19.3944
R8980 gnd.n3688 gnd.n2823 19.3944
R8981 gnd.n3688 gnd.n3687 19.3944
R8982 gnd.n3687 gnd.n2802 19.3944
R8983 gnd.n3710 gnd.n2802 19.3944
R8984 gnd.n3710 gnd.n3709 19.3944
R8985 gnd.n3709 gnd.n2779 19.3944
R8986 gnd.n3753 gnd.n2779 19.3944
R8987 gnd.n3753 gnd.n2772 19.3944
R8988 gnd.n3764 gnd.n2772 19.3944
R8989 gnd.n3764 gnd.n2768 19.3944
R8990 gnd.n4031 gnd.n2768 19.3944
R8991 gnd.n4031 gnd.n4030 19.3944
R8992 gnd.n4030 gnd.n2749 19.3944
R8993 gnd.n4054 gnd.n2749 19.3944
R8994 gnd.n6054 gnd.n1678 19.3944
R8995 gnd.n6059 gnd.n1678 19.3944
R8996 gnd.n6059 gnd.n1679 19.3944
R8997 gnd.n1679 gnd.n1654 19.3944
R8998 gnd.n6086 gnd.n1654 19.3944
R8999 gnd.n6086 gnd.n1651 19.3944
R9000 gnd.n6091 gnd.n1651 19.3944
R9001 gnd.n6091 gnd.n1652 19.3944
R9002 gnd.n1652 gnd.n1628 19.3944
R9003 gnd.n6118 gnd.n1628 19.3944
R9004 gnd.n6118 gnd.n1625 19.3944
R9005 gnd.n6123 gnd.n1625 19.3944
R9006 gnd.n6123 gnd.n1626 19.3944
R9007 gnd.n1626 gnd.n1598 19.3944
R9008 gnd.n6156 gnd.n1598 19.3944
R9009 gnd.n6156 gnd.n1595 19.3944
R9010 gnd.n6161 gnd.n1595 19.3944
R9011 gnd.n6161 gnd.n1596 19.3944
R9012 gnd.n1596 gnd.n1565 19.3944
R9013 gnd.n6222 gnd.n1565 19.3944
R9014 gnd.n6222 gnd.n1562 19.3944
R9015 gnd.n6229 gnd.n1562 19.3944
R9016 gnd.n6229 gnd.n1563 19.3944
R9017 gnd.n6225 gnd.n1563 19.3944
R9018 gnd.n6225 gnd.n1524 19.3944
R9019 gnd.n6300 gnd.n1524 19.3944
R9020 gnd.n6300 gnd.n1525 19.3944
R9021 gnd.n6296 gnd.n1525 19.3944
R9022 gnd.n6296 gnd.n6295 19.3944
R9023 gnd.n6295 gnd.n6294 19.3944
R9024 gnd.n6294 gnd.n6292 19.3944
R9025 gnd.n6292 gnd.n80 19.3944
R9026 gnd.n7968 gnd.n80 19.3944
R9027 gnd.n7968 gnd.n7967 19.3944
R9028 gnd.n7967 gnd.n7966 19.3944
R9029 gnd.n7966 gnd.n85 19.3944
R9030 gnd.n7962 gnd.n85 19.3944
R9031 gnd.n7962 gnd.n7961 19.3944
R9032 gnd.n7961 gnd.n7960 19.3944
R9033 gnd.n7960 gnd.n90 19.3944
R9034 gnd.n7956 gnd.n90 19.3944
R9035 gnd.n7956 gnd.n7955 19.3944
R9036 gnd.n7955 gnd.n7954 19.3944
R9037 gnd.n7954 gnd.n95 19.3944
R9038 gnd.n7950 gnd.n95 19.3944
R9039 gnd.n7950 gnd.n7949 19.3944
R9040 gnd.n7949 gnd.n7948 19.3944
R9041 gnd.n7948 gnd.n100 19.3944
R9042 gnd.n7944 gnd.n100 19.3944
R9043 gnd.n7944 gnd.n7943 19.3944
R9044 gnd.n7943 gnd.n7942 19.3944
R9045 gnd.n7942 gnd.n105 19.3944
R9046 gnd.n7938 gnd.n105 19.3944
R9047 gnd.n7938 gnd.n7937 19.3944
R9048 gnd.n7937 gnd.n7936 19.3944
R9049 gnd.n7936 gnd.n110 19.3944
R9050 gnd.n7932 gnd.n110 19.3944
R9051 gnd.n7932 gnd.n7931 19.3944
R9052 gnd.n7931 gnd.n7930 19.3944
R9053 gnd.n7930 gnd.n115 19.3944
R9054 gnd.n7926 gnd.n115 19.3944
R9055 gnd.n7926 gnd.n7925 19.3944
R9056 gnd.n7925 gnd.n7924 19.3944
R9057 gnd.n7924 gnd.n120 19.3944
R9058 gnd.n7832 gnd.n7831 19.3944
R9059 gnd.n7831 gnd.n7830 19.3944
R9060 gnd.n7830 gnd.n7779 19.3944
R9061 gnd.n7826 gnd.n7779 19.3944
R9062 gnd.n7826 gnd.n7825 19.3944
R9063 gnd.n7825 gnd.n7824 19.3944
R9064 gnd.n7824 gnd.n7787 19.3944
R9065 gnd.n7820 gnd.n7787 19.3944
R9066 gnd.n7820 gnd.n7819 19.3944
R9067 gnd.n7819 gnd.n7818 19.3944
R9068 gnd.n7818 gnd.n7795 19.3944
R9069 gnd.n7814 gnd.n7795 19.3944
R9070 gnd.n7814 gnd.n7813 19.3944
R9071 gnd.n7813 gnd.n7812 19.3944
R9072 gnd.n7812 gnd.n7803 19.3944
R9073 gnd.n7808 gnd.n7803 19.3944
R9074 gnd.n5931 gnd.n1480 19.3944
R9075 gnd.n5934 gnd.n5931 19.3944
R9076 gnd.n5934 gnd.n5925 19.3944
R9077 gnd.n5943 gnd.n5925 19.3944
R9078 gnd.n5946 gnd.n5943 19.3944
R9079 gnd.n5946 gnd.n5919 19.3944
R9080 gnd.n5955 gnd.n5919 19.3944
R9081 gnd.n5958 gnd.n5955 19.3944
R9082 gnd.n5958 gnd.n5913 19.3944
R9083 gnd.n5967 gnd.n5913 19.3944
R9084 gnd.n5970 gnd.n5967 19.3944
R9085 gnd.n5970 gnd.n5907 19.3944
R9086 gnd.n5979 gnd.n5907 19.3944
R9087 gnd.n5982 gnd.n5979 19.3944
R9088 gnd.n5982 gnd.n5901 19.3944
R9089 gnd.n5996 gnd.n5901 19.3944
R9090 gnd.n6348 gnd.n6347 19.3944
R9091 gnd.n6347 gnd.n6346 19.3944
R9092 gnd.n6346 gnd.n1485 19.3944
R9093 gnd.n6342 gnd.n1485 19.3944
R9094 gnd.n6342 gnd.n6341 19.3944
R9095 gnd.n6341 gnd.n6340 19.3944
R9096 gnd.n6340 gnd.n1490 19.3944
R9097 gnd.n6336 gnd.n1490 19.3944
R9098 gnd.n6336 gnd.n6335 19.3944
R9099 gnd.n6335 gnd.n6334 19.3944
R9100 gnd.n6334 gnd.n1495 19.3944
R9101 gnd.n6330 gnd.n1495 19.3944
R9102 gnd.n6330 gnd.n6329 19.3944
R9103 gnd.n6329 gnd.n6328 19.3944
R9104 gnd.n6328 gnd.n1500 19.3944
R9105 gnd.n6324 gnd.n1500 19.3944
R9106 gnd.n6324 gnd.n6323 19.3944
R9107 gnd.n6323 gnd.n6322 19.3944
R9108 gnd.n6322 gnd.n1505 19.3944
R9109 gnd.n6318 gnd.n1505 19.3944
R9110 gnd.n6318 gnd.n6317 19.3944
R9111 gnd.n6317 gnd.n6316 19.3944
R9112 gnd.n6316 gnd.n1510 19.3944
R9113 gnd.n6312 gnd.n1510 19.3944
R9114 gnd.n6312 gnd.n6311 19.3944
R9115 gnd.n6311 gnd.n6310 19.3944
R9116 gnd.n6310 gnd.n6307 19.3944
R9117 gnd.n6307 gnd.n326 19.3944
R9118 gnd.n7661 gnd.n326 19.3944
R9119 gnd.n7661 gnd.n327 19.3944
R9120 gnd.n7657 gnd.n327 19.3944
R9121 gnd.n7657 gnd.n7656 19.3944
R9122 gnd.n7656 gnd.n7655 19.3944
R9123 gnd.n7655 gnd.n333 19.3944
R9124 gnd.n7651 gnd.n333 19.3944
R9125 gnd.n7651 gnd.n304 19.3944
R9126 gnd.n7673 gnd.n304 19.3944
R9127 gnd.n7673 gnd.n302 19.3944
R9128 gnd.n7677 gnd.n302 19.3944
R9129 gnd.n7677 gnd.n289 19.3944
R9130 gnd.n7689 gnd.n289 19.3944
R9131 gnd.n7689 gnd.n287 19.3944
R9132 gnd.n7693 gnd.n287 19.3944
R9133 gnd.n7693 gnd.n273 19.3944
R9134 gnd.n7705 gnd.n273 19.3944
R9135 gnd.n7705 gnd.n271 19.3944
R9136 gnd.n7709 gnd.n271 19.3944
R9137 gnd.n7709 gnd.n257 19.3944
R9138 gnd.n7721 gnd.n257 19.3944
R9139 gnd.n7721 gnd.n255 19.3944
R9140 gnd.n7725 gnd.n255 19.3944
R9141 gnd.n7725 gnd.n241 19.3944
R9142 gnd.n7737 gnd.n241 19.3944
R9143 gnd.n7737 gnd.n239 19.3944
R9144 gnd.n7741 gnd.n239 19.3944
R9145 gnd.n7741 gnd.n227 19.3944
R9146 gnd.n7753 gnd.n227 19.3944
R9147 gnd.n7753 gnd.n225 19.3944
R9148 gnd.n7757 gnd.n225 19.3944
R9149 gnd.n7757 gnd.n210 19.3944
R9150 gnd.n7771 gnd.n210 19.3944
R9151 gnd.n7771 gnd.n207 19.3944
R9152 gnd.n7836 gnd.n207 19.3944
R9153 gnd.n7836 gnd.n208 19.3944
R9154 gnd.n2404 gnd.n2337 19.3944
R9155 gnd.n2405 gnd.n2404 19.3944
R9156 gnd.n4966 gnd.n2405 19.3944
R9157 gnd.n4966 gnd.n4965 19.3944
R9158 gnd.n4965 gnd.n2410 19.3944
R9159 gnd.n4958 gnd.n2410 19.3944
R9160 gnd.n4958 gnd.n4957 19.3944
R9161 gnd.n4957 gnd.n2419 19.3944
R9162 gnd.n4950 gnd.n2419 19.3944
R9163 gnd.n4950 gnd.n4949 19.3944
R9164 gnd.n4949 gnd.n2429 19.3944
R9165 gnd.n4942 gnd.n2429 19.3944
R9166 gnd.n4942 gnd.n4941 19.3944
R9167 gnd.n4941 gnd.n2439 19.3944
R9168 gnd.n4934 gnd.n2439 19.3944
R9169 gnd.n4934 gnd.n4933 19.3944
R9170 gnd.n7402 gnd.n537 19.3944
R9171 gnd.n7402 gnd.n533 19.3944
R9172 gnd.n7408 gnd.n533 19.3944
R9173 gnd.n7408 gnd.n531 19.3944
R9174 gnd.n7412 gnd.n531 19.3944
R9175 gnd.n7412 gnd.n527 19.3944
R9176 gnd.n7418 gnd.n527 19.3944
R9177 gnd.n7418 gnd.n525 19.3944
R9178 gnd.n7422 gnd.n525 19.3944
R9179 gnd.n7422 gnd.n521 19.3944
R9180 gnd.n7428 gnd.n521 19.3944
R9181 gnd.n7428 gnd.n519 19.3944
R9182 gnd.n7432 gnd.n519 19.3944
R9183 gnd.n7432 gnd.n515 19.3944
R9184 gnd.n7438 gnd.n515 19.3944
R9185 gnd.n7438 gnd.n513 19.3944
R9186 gnd.n7442 gnd.n513 19.3944
R9187 gnd.n7442 gnd.n509 19.3944
R9188 gnd.n7448 gnd.n509 19.3944
R9189 gnd.n7448 gnd.n507 19.3944
R9190 gnd.n7452 gnd.n507 19.3944
R9191 gnd.n7452 gnd.n503 19.3944
R9192 gnd.n7458 gnd.n503 19.3944
R9193 gnd.n7458 gnd.n501 19.3944
R9194 gnd.n7462 gnd.n501 19.3944
R9195 gnd.n7462 gnd.n497 19.3944
R9196 gnd.n7468 gnd.n497 19.3944
R9197 gnd.n7468 gnd.n495 19.3944
R9198 gnd.n7472 gnd.n495 19.3944
R9199 gnd.n7472 gnd.n491 19.3944
R9200 gnd.n7478 gnd.n491 19.3944
R9201 gnd.n7478 gnd.n489 19.3944
R9202 gnd.n7482 gnd.n489 19.3944
R9203 gnd.n7482 gnd.n485 19.3944
R9204 gnd.n7488 gnd.n485 19.3944
R9205 gnd.n7488 gnd.n483 19.3944
R9206 gnd.n7492 gnd.n483 19.3944
R9207 gnd.n7492 gnd.n479 19.3944
R9208 gnd.n7498 gnd.n479 19.3944
R9209 gnd.n7498 gnd.n477 19.3944
R9210 gnd.n7502 gnd.n477 19.3944
R9211 gnd.n7502 gnd.n473 19.3944
R9212 gnd.n7508 gnd.n473 19.3944
R9213 gnd.n7508 gnd.n471 19.3944
R9214 gnd.n7512 gnd.n471 19.3944
R9215 gnd.n7512 gnd.n467 19.3944
R9216 gnd.n7518 gnd.n467 19.3944
R9217 gnd.n7518 gnd.n465 19.3944
R9218 gnd.n7522 gnd.n465 19.3944
R9219 gnd.n7522 gnd.n461 19.3944
R9220 gnd.n7528 gnd.n461 19.3944
R9221 gnd.n7528 gnd.n459 19.3944
R9222 gnd.n7532 gnd.n459 19.3944
R9223 gnd.n7532 gnd.n455 19.3944
R9224 gnd.n7538 gnd.n455 19.3944
R9225 gnd.n7538 gnd.n453 19.3944
R9226 gnd.n7542 gnd.n453 19.3944
R9227 gnd.n7542 gnd.n449 19.3944
R9228 gnd.n7548 gnd.n449 19.3944
R9229 gnd.n7548 gnd.n447 19.3944
R9230 gnd.n7552 gnd.n447 19.3944
R9231 gnd.n7552 gnd.n443 19.3944
R9232 gnd.n7558 gnd.n443 19.3944
R9233 gnd.n7558 gnd.n441 19.3944
R9234 gnd.n7562 gnd.n441 19.3944
R9235 gnd.n7562 gnd.n437 19.3944
R9236 gnd.n7568 gnd.n437 19.3944
R9237 gnd.n7568 gnd.n435 19.3944
R9238 gnd.n7572 gnd.n435 19.3944
R9239 gnd.n7572 gnd.n431 19.3944
R9240 gnd.n7578 gnd.n431 19.3944
R9241 gnd.n7578 gnd.n429 19.3944
R9242 gnd.n7582 gnd.n429 19.3944
R9243 gnd.n7582 gnd.n425 19.3944
R9244 gnd.n7588 gnd.n425 19.3944
R9245 gnd.n7588 gnd.n423 19.3944
R9246 gnd.n7592 gnd.n423 19.3944
R9247 gnd.n7592 gnd.n419 19.3944
R9248 gnd.n7598 gnd.n419 19.3944
R9249 gnd.n7598 gnd.n417 19.3944
R9250 gnd.n7604 gnd.n417 19.3944
R9251 gnd.n7604 gnd.n7603 19.3944
R9252 gnd.n7603 gnd.n413 19.3944
R9253 gnd.n7611 gnd.n413 19.3944
R9254 gnd.n6882 gnd.n849 19.3944
R9255 gnd.n6882 gnd.n845 19.3944
R9256 gnd.n6888 gnd.n845 19.3944
R9257 gnd.n6888 gnd.n843 19.3944
R9258 gnd.n6892 gnd.n843 19.3944
R9259 gnd.n6892 gnd.n839 19.3944
R9260 gnd.n6898 gnd.n839 19.3944
R9261 gnd.n6898 gnd.n837 19.3944
R9262 gnd.n6902 gnd.n837 19.3944
R9263 gnd.n6902 gnd.n833 19.3944
R9264 gnd.n6908 gnd.n833 19.3944
R9265 gnd.n6908 gnd.n831 19.3944
R9266 gnd.n6912 gnd.n831 19.3944
R9267 gnd.n6912 gnd.n827 19.3944
R9268 gnd.n6918 gnd.n827 19.3944
R9269 gnd.n6918 gnd.n825 19.3944
R9270 gnd.n6922 gnd.n825 19.3944
R9271 gnd.n6922 gnd.n821 19.3944
R9272 gnd.n6928 gnd.n821 19.3944
R9273 gnd.n6928 gnd.n819 19.3944
R9274 gnd.n6932 gnd.n819 19.3944
R9275 gnd.n6932 gnd.n815 19.3944
R9276 gnd.n6938 gnd.n815 19.3944
R9277 gnd.n6938 gnd.n813 19.3944
R9278 gnd.n6942 gnd.n813 19.3944
R9279 gnd.n6942 gnd.n809 19.3944
R9280 gnd.n6948 gnd.n809 19.3944
R9281 gnd.n6948 gnd.n807 19.3944
R9282 gnd.n6952 gnd.n807 19.3944
R9283 gnd.n6952 gnd.n803 19.3944
R9284 gnd.n6958 gnd.n803 19.3944
R9285 gnd.n6958 gnd.n801 19.3944
R9286 gnd.n6962 gnd.n801 19.3944
R9287 gnd.n6962 gnd.n797 19.3944
R9288 gnd.n6968 gnd.n797 19.3944
R9289 gnd.n6968 gnd.n795 19.3944
R9290 gnd.n6972 gnd.n795 19.3944
R9291 gnd.n6972 gnd.n791 19.3944
R9292 gnd.n6978 gnd.n791 19.3944
R9293 gnd.n6978 gnd.n789 19.3944
R9294 gnd.n6982 gnd.n789 19.3944
R9295 gnd.n6982 gnd.n785 19.3944
R9296 gnd.n6988 gnd.n785 19.3944
R9297 gnd.n6988 gnd.n783 19.3944
R9298 gnd.n6992 gnd.n783 19.3944
R9299 gnd.n6992 gnd.n779 19.3944
R9300 gnd.n6998 gnd.n779 19.3944
R9301 gnd.n6998 gnd.n777 19.3944
R9302 gnd.n7002 gnd.n777 19.3944
R9303 gnd.n7002 gnd.n773 19.3944
R9304 gnd.n7008 gnd.n773 19.3944
R9305 gnd.n7008 gnd.n771 19.3944
R9306 gnd.n7012 gnd.n771 19.3944
R9307 gnd.n7012 gnd.n767 19.3944
R9308 gnd.n7018 gnd.n767 19.3944
R9309 gnd.n7018 gnd.n765 19.3944
R9310 gnd.n7022 gnd.n765 19.3944
R9311 gnd.n7022 gnd.n761 19.3944
R9312 gnd.n7028 gnd.n761 19.3944
R9313 gnd.n7028 gnd.n759 19.3944
R9314 gnd.n7032 gnd.n759 19.3944
R9315 gnd.n7032 gnd.n755 19.3944
R9316 gnd.n7038 gnd.n755 19.3944
R9317 gnd.n7038 gnd.n753 19.3944
R9318 gnd.n7042 gnd.n753 19.3944
R9319 gnd.n7042 gnd.n749 19.3944
R9320 gnd.n7048 gnd.n749 19.3944
R9321 gnd.n7048 gnd.n747 19.3944
R9322 gnd.n7052 gnd.n747 19.3944
R9323 gnd.n7052 gnd.n743 19.3944
R9324 gnd.n7058 gnd.n743 19.3944
R9325 gnd.n7058 gnd.n741 19.3944
R9326 gnd.n7062 gnd.n741 19.3944
R9327 gnd.n7062 gnd.n737 19.3944
R9328 gnd.n7068 gnd.n737 19.3944
R9329 gnd.n7068 gnd.n735 19.3944
R9330 gnd.n7072 gnd.n735 19.3944
R9331 gnd.n7072 gnd.n731 19.3944
R9332 gnd.n7078 gnd.n731 19.3944
R9333 gnd.n7078 gnd.n729 19.3944
R9334 gnd.n7082 gnd.n729 19.3944
R9335 gnd.n7082 gnd.n725 19.3944
R9336 gnd.n7088 gnd.n725 19.3944
R9337 gnd.n7088 gnd.n723 19.3944
R9338 gnd.n7092 gnd.n723 19.3944
R9339 gnd.n7092 gnd.n719 19.3944
R9340 gnd.n7098 gnd.n719 19.3944
R9341 gnd.n7098 gnd.n717 19.3944
R9342 gnd.n7102 gnd.n717 19.3944
R9343 gnd.n7102 gnd.n713 19.3944
R9344 gnd.n7108 gnd.n713 19.3944
R9345 gnd.n7108 gnd.n711 19.3944
R9346 gnd.n7112 gnd.n711 19.3944
R9347 gnd.n7112 gnd.n707 19.3944
R9348 gnd.n7118 gnd.n707 19.3944
R9349 gnd.n7118 gnd.n705 19.3944
R9350 gnd.n7122 gnd.n705 19.3944
R9351 gnd.n7122 gnd.n701 19.3944
R9352 gnd.n7128 gnd.n701 19.3944
R9353 gnd.n7128 gnd.n699 19.3944
R9354 gnd.n7132 gnd.n699 19.3944
R9355 gnd.n7132 gnd.n695 19.3944
R9356 gnd.n7138 gnd.n695 19.3944
R9357 gnd.n7138 gnd.n693 19.3944
R9358 gnd.n7142 gnd.n693 19.3944
R9359 gnd.n7142 gnd.n689 19.3944
R9360 gnd.n7148 gnd.n689 19.3944
R9361 gnd.n7148 gnd.n687 19.3944
R9362 gnd.n7152 gnd.n687 19.3944
R9363 gnd.n7152 gnd.n683 19.3944
R9364 gnd.n7158 gnd.n683 19.3944
R9365 gnd.n7158 gnd.n681 19.3944
R9366 gnd.n7162 gnd.n681 19.3944
R9367 gnd.n7162 gnd.n677 19.3944
R9368 gnd.n7168 gnd.n677 19.3944
R9369 gnd.n7168 gnd.n675 19.3944
R9370 gnd.n7172 gnd.n675 19.3944
R9371 gnd.n7172 gnd.n671 19.3944
R9372 gnd.n7178 gnd.n671 19.3944
R9373 gnd.n7178 gnd.n669 19.3944
R9374 gnd.n7182 gnd.n669 19.3944
R9375 gnd.n7182 gnd.n665 19.3944
R9376 gnd.n7188 gnd.n665 19.3944
R9377 gnd.n7188 gnd.n663 19.3944
R9378 gnd.n7192 gnd.n663 19.3944
R9379 gnd.n7192 gnd.n659 19.3944
R9380 gnd.n7198 gnd.n659 19.3944
R9381 gnd.n7198 gnd.n657 19.3944
R9382 gnd.n7202 gnd.n657 19.3944
R9383 gnd.n7202 gnd.n653 19.3944
R9384 gnd.n7208 gnd.n653 19.3944
R9385 gnd.n7208 gnd.n651 19.3944
R9386 gnd.n7212 gnd.n651 19.3944
R9387 gnd.n7212 gnd.n647 19.3944
R9388 gnd.n7218 gnd.n647 19.3944
R9389 gnd.n7218 gnd.n645 19.3944
R9390 gnd.n7222 gnd.n645 19.3944
R9391 gnd.n7222 gnd.n641 19.3944
R9392 gnd.n7228 gnd.n641 19.3944
R9393 gnd.n7228 gnd.n639 19.3944
R9394 gnd.n7232 gnd.n639 19.3944
R9395 gnd.n7232 gnd.n635 19.3944
R9396 gnd.n7238 gnd.n635 19.3944
R9397 gnd.n7238 gnd.n633 19.3944
R9398 gnd.n7242 gnd.n633 19.3944
R9399 gnd.n7242 gnd.n629 19.3944
R9400 gnd.n7248 gnd.n629 19.3944
R9401 gnd.n7248 gnd.n627 19.3944
R9402 gnd.n7252 gnd.n627 19.3944
R9403 gnd.n7252 gnd.n623 19.3944
R9404 gnd.n7258 gnd.n623 19.3944
R9405 gnd.n7258 gnd.n621 19.3944
R9406 gnd.n7262 gnd.n621 19.3944
R9407 gnd.n7262 gnd.n617 19.3944
R9408 gnd.n7268 gnd.n617 19.3944
R9409 gnd.n7268 gnd.n615 19.3944
R9410 gnd.n7272 gnd.n615 19.3944
R9411 gnd.n7272 gnd.n611 19.3944
R9412 gnd.n7278 gnd.n611 19.3944
R9413 gnd.n7278 gnd.n609 19.3944
R9414 gnd.n7282 gnd.n609 19.3944
R9415 gnd.n7282 gnd.n605 19.3944
R9416 gnd.n7288 gnd.n605 19.3944
R9417 gnd.n7288 gnd.n603 19.3944
R9418 gnd.n7292 gnd.n603 19.3944
R9419 gnd.n7292 gnd.n599 19.3944
R9420 gnd.n7298 gnd.n599 19.3944
R9421 gnd.n7298 gnd.n597 19.3944
R9422 gnd.n7302 gnd.n597 19.3944
R9423 gnd.n7302 gnd.n593 19.3944
R9424 gnd.n7308 gnd.n593 19.3944
R9425 gnd.n7308 gnd.n591 19.3944
R9426 gnd.n7312 gnd.n591 19.3944
R9427 gnd.n7312 gnd.n587 19.3944
R9428 gnd.n7318 gnd.n587 19.3944
R9429 gnd.n7318 gnd.n585 19.3944
R9430 gnd.n7322 gnd.n585 19.3944
R9431 gnd.n7322 gnd.n581 19.3944
R9432 gnd.n7328 gnd.n581 19.3944
R9433 gnd.n7328 gnd.n579 19.3944
R9434 gnd.n7332 gnd.n579 19.3944
R9435 gnd.n7332 gnd.n575 19.3944
R9436 gnd.n7338 gnd.n575 19.3944
R9437 gnd.n7338 gnd.n573 19.3944
R9438 gnd.n7342 gnd.n573 19.3944
R9439 gnd.n7342 gnd.n569 19.3944
R9440 gnd.n7348 gnd.n569 19.3944
R9441 gnd.n7348 gnd.n567 19.3944
R9442 gnd.n7352 gnd.n567 19.3944
R9443 gnd.n7352 gnd.n563 19.3944
R9444 gnd.n7358 gnd.n563 19.3944
R9445 gnd.n7358 gnd.n561 19.3944
R9446 gnd.n7362 gnd.n561 19.3944
R9447 gnd.n7362 gnd.n557 19.3944
R9448 gnd.n7368 gnd.n557 19.3944
R9449 gnd.n7368 gnd.n555 19.3944
R9450 gnd.n7372 gnd.n555 19.3944
R9451 gnd.n7372 gnd.n551 19.3944
R9452 gnd.n7378 gnd.n551 19.3944
R9453 gnd.n7378 gnd.n549 19.3944
R9454 gnd.n7382 gnd.n549 19.3944
R9455 gnd.n7382 gnd.n545 19.3944
R9456 gnd.n7388 gnd.n545 19.3944
R9457 gnd.n7388 gnd.n543 19.3944
R9458 gnd.n7392 gnd.n543 19.3944
R9459 gnd.n7392 gnd.n539 19.3944
R9460 gnd.n7398 gnd.n539 19.3944
R9461 gnd.n6045 gnd.n6044 19.3944
R9462 gnd.n6044 gnd.n1688 19.3944
R9463 gnd.n1843 gnd.n1688 19.3944
R9464 gnd.n1847 gnd.n1843 19.3944
R9465 gnd.n1850 gnd.n1847 19.3944
R9466 gnd.n1853 gnd.n1850 19.3944
R9467 gnd.n1853 gnd.n1840 19.3944
R9468 gnd.n1857 gnd.n1840 19.3944
R9469 gnd.n1860 gnd.n1857 19.3944
R9470 gnd.n1863 gnd.n1860 19.3944
R9471 gnd.n1863 gnd.n1838 19.3944
R9472 gnd.n1867 gnd.n1838 19.3944
R9473 gnd.n1870 gnd.n1867 19.3944
R9474 gnd.n1873 gnd.n1870 19.3944
R9475 gnd.n1873 gnd.n1835 19.3944
R9476 gnd.n1983 gnd.n1980 19.3944
R9477 gnd.n1980 gnd.n1979 19.3944
R9478 gnd.n1979 gnd.n1976 19.3944
R9479 gnd.n1976 gnd.n1975 19.3944
R9480 gnd.n1975 gnd.n1972 19.3944
R9481 gnd.n1972 gnd.n1971 19.3944
R9482 gnd.n1971 gnd.n1968 19.3944
R9483 gnd.n1968 gnd.n1967 19.3944
R9484 gnd.n1967 gnd.n1964 19.3944
R9485 gnd.n1964 gnd.n1963 19.3944
R9486 gnd.n1963 gnd.n1960 19.3944
R9487 gnd.n1960 gnd.n1959 19.3944
R9488 gnd.n1959 gnd.n1956 19.3944
R9489 gnd.n1956 gnd.n1955 19.3944
R9490 gnd.n1955 gnd.n1952 19.3944
R9491 gnd.n1952 gnd.n1951 19.3944
R9492 gnd.n1951 gnd.n1948 19.3944
R9493 gnd.n1948 gnd.n1947 19.3944
R9494 gnd.n1940 gnd.n1939 19.3944
R9495 gnd.n1939 gnd.n1938 19.3944
R9496 gnd.n1938 gnd.n1937 19.3944
R9497 gnd.n1937 gnd.n1936 19.3944
R9498 gnd.n1936 gnd.n1934 19.3944
R9499 gnd.n1934 gnd.n1933 19.3944
R9500 gnd.n1933 gnd.n1930 19.3944
R9501 gnd.n1930 gnd.n1929 19.3944
R9502 gnd.n1929 gnd.n1928 19.3944
R9503 gnd.n1928 gnd.n1926 19.3944
R9504 gnd.n1926 gnd.n1925 19.3944
R9505 gnd.n1925 gnd.n1923 19.3944
R9506 gnd.n1923 gnd.n1922 19.3944
R9507 gnd.n1922 gnd.n1921 19.3944
R9508 gnd.n1921 gnd.n1919 19.3944
R9509 gnd.n1919 gnd.n1590 19.3944
R9510 gnd.n6165 gnd.n1590 19.3944
R9511 gnd.n6166 gnd.n6165 19.3944
R9512 gnd.n6168 gnd.n6166 19.3944
R9513 gnd.n6168 gnd.n1588 19.3944
R9514 gnd.n6202 gnd.n1588 19.3944
R9515 gnd.n6202 gnd.n6201 19.3944
R9516 gnd.n6201 gnd.n6200 19.3944
R9517 gnd.n6200 gnd.n6198 19.3944
R9518 gnd.n6198 gnd.n6197 19.3944
R9519 gnd.n6197 gnd.n6194 19.3944
R9520 gnd.n6194 gnd.n6193 19.3944
R9521 gnd.n6193 gnd.n6192 19.3944
R9522 gnd.n6192 gnd.n6189 19.3944
R9523 gnd.n6189 gnd.n6188 19.3944
R9524 gnd.n6188 gnd.n6185 19.3944
R9525 gnd.n6185 gnd.n6184 19.3944
R9526 gnd.n6184 gnd.n341 19.3944
R9527 gnd.n7642 gnd.n341 19.3944
R9528 gnd.n7642 gnd.n7641 19.3944
R9529 gnd.n7641 gnd.n7640 19.3944
R9530 gnd.n7640 gnd.n7636 19.3944
R9531 gnd.n7636 gnd.n7635 19.3944
R9532 gnd.n7635 gnd.n7632 19.3944
R9533 gnd.n7632 gnd.n7631 19.3944
R9534 gnd.n7631 gnd.n7627 19.3944
R9535 gnd.n7627 gnd.n7626 19.3944
R9536 gnd.n7626 gnd.n401 19.3944
R9537 gnd.n401 gnd.n400 19.3944
R9538 gnd.n400 gnd.n396 19.3944
R9539 gnd.n396 gnd.n395 19.3944
R9540 gnd.n395 gnd.n392 19.3944
R9541 gnd.n392 gnd.n391 19.3944
R9542 gnd.n391 gnd.n389 19.3944
R9543 gnd.n389 gnd.n388 19.3944
R9544 gnd.n388 gnd.n386 19.3944
R9545 gnd.n386 gnd.n385 19.3944
R9546 gnd.n385 gnd.n383 19.3944
R9547 gnd.n383 gnd.n382 19.3944
R9548 gnd.n382 gnd.n380 19.3944
R9549 gnd.n380 gnd.n379 19.3944
R9550 gnd.n379 gnd.n377 19.3944
R9551 gnd.n377 gnd.n376 19.3944
R9552 gnd.n376 gnd.n374 19.3944
R9553 gnd.n374 gnd.n373 19.3944
R9554 gnd.n373 gnd.n371 19.3944
R9555 gnd.n371 gnd.n204 19.3944
R9556 gnd.n7840 gnd.n204 19.3944
R9557 gnd.n7841 gnd.n7840 19.3944
R9558 gnd.n7879 gnd.n165 19.3944
R9559 gnd.n7874 gnd.n165 19.3944
R9560 gnd.n7874 gnd.n7873 19.3944
R9561 gnd.n7873 gnd.n7872 19.3944
R9562 gnd.n7872 gnd.n172 19.3944
R9563 gnd.n7867 gnd.n172 19.3944
R9564 gnd.n7867 gnd.n7866 19.3944
R9565 gnd.n7866 gnd.n7865 19.3944
R9566 gnd.n7865 gnd.n179 19.3944
R9567 gnd.n7860 gnd.n179 19.3944
R9568 gnd.n7860 gnd.n7859 19.3944
R9569 gnd.n7859 gnd.n7858 19.3944
R9570 gnd.n7858 gnd.n186 19.3944
R9571 gnd.n7853 gnd.n186 19.3944
R9572 gnd.n7853 gnd.n7852 19.3944
R9573 gnd.n7852 gnd.n7851 19.3944
R9574 gnd.n7851 gnd.n193 19.3944
R9575 gnd.n7846 gnd.n193 19.3944
R9576 gnd.n7912 gnd.n7911 19.3944
R9577 gnd.n7911 gnd.n7910 19.3944
R9578 gnd.n7910 gnd.n137 19.3944
R9579 gnd.n7905 gnd.n137 19.3944
R9580 gnd.n7905 gnd.n7904 19.3944
R9581 gnd.n7904 gnd.n7903 19.3944
R9582 gnd.n7903 gnd.n144 19.3944
R9583 gnd.n7898 gnd.n144 19.3944
R9584 gnd.n7898 gnd.n7897 19.3944
R9585 gnd.n7897 gnd.n7896 19.3944
R9586 gnd.n7896 gnd.n151 19.3944
R9587 gnd.n7891 gnd.n151 19.3944
R9588 gnd.n7891 gnd.n7890 19.3944
R9589 gnd.n7890 gnd.n7889 19.3944
R9590 gnd.n7889 gnd.n158 19.3944
R9591 gnd.n7884 gnd.n158 19.3944
R9592 gnd.n7884 gnd.n7883 19.3944
R9593 gnd.n6050 gnd.n6049 19.3944
R9594 gnd.n6049 gnd.n1663 19.3944
R9595 gnd.n6076 gnd.n1663 19.3944
R9596 gnd.n6076 gnd.n1661 19.3944
R9597 gnd.n6082 gnd.n1661 19.3944
R9598 gnd.n6082 gnd.n6081 19.3944
R9599 gnd.n6081 gnd.n1637 19.3944
R9600 gnd.n6108 gnd.n1637 19.3944
R9601 gnd.n6108 gnd.n1635 19.3944
R9602 gnd.n6114 gnd.n1635 19.3944
R9603 gnd.n6114 gnd.n6113 19.3944
R9604 gnd.n6113 gnd.n1609 19.3944
R9605 gnd.n6146 gnd.n1609 19.3944
R9606 gnd.n6146 gnd.n1607 19.3944
R9607 gnd.n6152 gnd.n1607 19.3944
R9608 gnd.n6152 gnd.n6151 19.3944
R9609 gnd.n6151 gnd.n1572 19.3944
R9610 gnd.n6214 gnd.n1572 19.3944
R9611 gnd.n6214 gnd.n1570 19.3944
R9612 gnd.n6218 gnd.n1570 19.3944
R9613 gnd.n6218 gnd.n1556 19.3944
R9614 gnd.n6234 gnd.n1556 19.3944
R9615 gnd.n6234 gnd.n1554 19.3944
R9616 gnd.n6240 gnd.n1554 19.3944
R9617 gnd.n6240 gnd.n6239 19.3944
R9618 gnd.n6239 gnd.n1520 19.3944
R9619 gnd.n1520 gnd.n317 19.3944
R9620 gnd.n7666 gnd.n7665 19.3944
R9621 gnd.n6288 gnd.n6287 19.3944
R9622 gnd.n1535 gnd.n1534 19.3944
R9623 gnd.n7647 gnd.n7646 19.3944
R9624 gnd.n7669 gnd.n310 19.3944
R9625 gnd.n7669 gnd.n296 19.3944
R9626 gnd.n7681 gnd.n296 19.3944
R9627 gnd.n7681 gnd.n294 19.3944
R9628 gnd.n7685 gnd.n294 19.3944
R9629 gnd.n7685 gnd.n281 19.3944
R9630 gnd.n7697 gnd.n281 19.3944
R9631 gnd.n7697 gnd.n279 19.3944
R9632 gnd.n7701 gnd.n279 19.3944
R9633 gnd.n7701 gnd.n264 19.3944
R9634 gnd.n7713 gnd.n264 19.3944
R9635 gnd.n7713 gnd.n262 19.3944
R9636 gnd.n7717 gnd.n262 19.3944
R9637 gnd.n7717 gnd.n250 19.3944
R9638 gnd.n7729 gnd.n250 19.3944
R9639 gnd.n7729 gnd.n248 19.3944
R9640 gnd.n7733 gnd.n248 19.3944
R9641 gnd.n7733 gnd.n235 19.3944
R9642 gnd.n7745 gnd.n235 19.3944
R9643 gnd.n7745 gnd.n233 19.3944
R9644 gnd.n7749 gnd.n233 19.3944
R9645 gnd.n7749 gnd.n220 19.3944
R9646 gnd.n7761 gnd.n220 19.3944
R9647 gnd.n7761 gnd.n218 19.3944
R9648 gnd.n7767 gnd.n218 19.3944
R9649 gnd.n7767 gnd.n7766 19.3944
R9650 gnd.n7766 gnd.n132 19.3944
R9651 gnd.n7915 gnd.n132 19.3944
R9652 gnd.n2592 gnd.n2590 19.3944
R9653 gnd.n2592 gnd.n2588 19.3944
R9654 gnd.n2607 gnd.n2588 19.3944
R9655 gnd.n2607 gnd.n2606 19.3944
R9656 gnd.n2606 gnd.n2605 19.3944
R9657 gnd.n2605 gnd.n2602 19.3944
R9658 gnd.n2602 gnd.n2601 19.3944
R9659 gnd.n2601 gnd.n2576 19.3944
R9660 gnd.n4555 gnd.n2576 19.3944
R9661 gnd.n4556 gnd.n4555 19.3944
R9662 gnd.n4560 gnd.n4559 19.3944
R9663 gnd.n4600 gnd.n2546 19.3944
R9664 gnd.n4613 gnd.n4602 19.3944
R9665 gnd.n4611 gnd.n4610 19.3944
R9666 gnd.n4607 gnd.n4606 19.3944
R9667 gnd.n4606 gnd.n2512 19.3944
R9668 gnd.n2512 gnd.n2510 19.3944
R9669 gnd.n4681 gnd.n2510 19.3944
R9670 gnd.n4681 gnd.n2508 19.3944
R9671 gnd.n4685 gnd.n2508 19.3944
R9672 gnd.n4685 gnd.n2506 19.3944
R9673 gnd.n4689 gnd.n2506 19.3944
R9674 gnd.n4689 gnd.n2504 19.3944
R9675 gnd.n4710 gnd.n2504 19.3944
R9676 gnd.n4710 gnd.n4709 19.3944
R9677 gnd.n4709 gnd.n4708 19.3944
R9678 gnd.n4708 gnd.n4695 19.3944
R9679 gnd.n4704 gnd.n4695 19.3944
R9680 gnd.n4704 gnd.n4703 19.3944
R9681 gnd.n4703 gnd.n4702 19.3944
R9682 gnd.n4702 gnd.n2473 19.3944
R9683 gnd.n4891 gnd.n2473 19.3944
R9684 gnd.n4891 gnd.n2471 19.3944
R9685 gnd.n4895 gnd.n2471 19.3944
R9686 gnd.n4895 gnd.n2469 19.3944
R9687 gnd.n4899 gnd.n2469 19.3944
R9688 gnd.n4899 gnd.n2467 19.3944
R9689 gnd.n4903 gnd.n2467 19.3944
R9690 gnd.n4903 gnd.n2465 19.3944
R9691 gnd.n4907 gnd.n2465 19.3944
R9692 gnd.n4907 gnd.n2463 19.3944
R9693 gnd.n4920 gnd.n2463 19.3944
R9694 gnd.n4920 gnd.n4919 19.3944
R9695 gnd.n4919 gnd.n4918 19.3944
R9696 gnd.n4918 gnd.n4914 19.3944
R9697 gnd.n4914 gnd.n2314 19.3944
R9698 gnd.n4976 gnd.n2314 19.3944
R9699 gnd.n4976 gnd.n2312 19.3944
R9700 gnd.n4980 gnd.n2312 19.3944
R9701 gnd.n4980 gnd.n2300 19.3944
R9702 gnd.n4992 gnd.n2300 19.3944
R9703 gnd.n4992 gnd.n2298 19.3944
R9704 gnd.n4996 gnd.n2298 19.3944
R9705 gnd.n4996 gnd.n2286 19.3944
R9706 gnd.n5008 gnd.n2286 19.3944
R9707 gnd.n5008 gnd.n2284 19.3944
R9708 gnd.n5012 gnd.n2284 19.3944
R9709 gnd.n5012 gnd.n2272 19.3944
R9710 gnd.n5024 gnd.n2272 19.3944
R9711 gnd.n5024 gnd.n2270 19.3944
R9712 gnd.n5028 gnd.n2270 19.3944
R9713 gnd.n5028 gnd.n2258 19.3944
R9714 gnd.n5040 gnd.n2258 19.3944
R9715 gnd.n5040 gnd.n2256 19.3944
R9716 gnd.n5044 gnd.n2256 19.3944
R9717 gnd.n5044 gnd.n2243 19.3944
R9718 gnd.n5056 gnd.n2243 19.3944
R9719 gnd.n5056 gnd.n2241 19.3944
R9720 gnd.n5060 gnd.n2241 19.3944
R9721 gnd.n5060 gnd.n2228 19.3944
R9722 gnd.n5083 gnd.n2228 19.3944
R9723 gnd.n5083 gnd.n2226 19.3944
R9724 gnd.n5090 gnd.n2226 19.3944
R9725 gnd.n5090 gnd.n5089 19.3944
R9726 gnd.n5089 gnd.n1370 19.3944
R9727 gnd.n6470 gnd.n1370 19.3944
R9728 gnd.n6470 gnd.n6469 19.3944
R9729 gnd.n6469 gnd.n6468 19.3944
R9730 gnd.n6468 gnd.n1374 19.3944
R9731 gnd.n5243 gnd.n1374 19.3944
R9732 gnd.n5243 gnd.n2199 19.3944
R9733 gnd.n5266 gnd.n2199 19.3944
R9734 gnd.n5266 gnd.n2197 19.3944
R9735 gnd.n5270 gnd.n2197 19.3944
R9736 gnd.n5270 gnd.n2180 19.3944
R9737 gnd.n5290 gnd.n2180 19.3944
R9738 gnd.n5290 gnd.n2178 19.3944
R9739 gnd.n5294 gnd.n2178 19.3944
R9740 gnd.n5294 gnd.n2158 19.3944
R9741 gnd.n5316 gnd.n2158 19.3944
R9742 gnd.n5316 gnd.n2156 19.3944
R9743 gnd.n5322 gnd.n2156 19.3944
R9744 gnd.n5322 gnd.n5321 19.3944
R9745 gnd.n5321 gnd.n2129 19.3944
R9746 gnd.n5371 gnd.n2129 19.3944
R9747 gnd.n5371 gnd.n2127 19.3944
R9748 gnd.n5377 gnd.n2127 19.3944
R9749 gnd.n5377 gnd.n5376 19.3944
R9750 gnd.n5376 gnd.n2106 19.3944
R9751 gnd.n5412 gnd.n2106 19.3944
R9752 gnd.n5412 gnd.n2104 19.3944
R9753 gnd.n5418 gnd.n2104 19.3944
R9754 gnd.n5418 gnd.n5417 19.3944
R9755 gnd.n5417 gnd.n2077 19.3944
R9756 gnd.n5453 gnd.n2077 19.3944
R9757 gnd.n5453 gnd.n2075 19.3944
R9758 gnd.n5458 gnd.n2075 19.3944
R9759 gnd.n5458 gnd.n2053 19.3944
R9760 gnd.n5505 gnd.n2053 19.3944
R9761 gnd.n5505 gnd.n5504 19.3944
R9762 gnd.n5504 gnd.n5503 19.3944
R9763 gnd.n5503 gnd.n2057 19.3944
R9764 gnd.n2060 gnd.n2057 19.3944
R9765 gnd.n2060 gnd.n2019 19.3944
R9766 gnd.n5553 gnd.n2019 19.3944
R9767 gnd.n5553 gnd.n2017 19.3944
R9768 gnd.n5557 gnd.n2017 19.3944
R9769 gnd.n5557 gnd.n2003 19.3944
R9770 gnd.n5584 gnd.n2003 19.3944
R9771 gnd.n5584 gnd.n2001 19.3944
R9772 gnd.n5588 gnd.n2001 19.3944
R9773 gnd.n5588 gnd.n1797 19.3944
R9774 gnd.n5759 gnd.n1797 19.3944
R9775 gnd.n5759 gnd.n1795 19.3944
R9776 gnd.n5763 gnd.n1795 19.3944
R9777 gnd.n5763 gnd.n1785 19.3944
R9778 gnd.n5777 gnd.n1785 19.3944
R9779 gnd.n5777 gnd.n1783 19.3944
R9780 gnd.n5781 gnd.n1783 19.3944
R9781 gnd.n5781 gnd.n1774 19.3944
R9782 gnd.n5794 gnd.n1774 19.3944
R9783 gnd.n5794 gnd.n1772 19.3944
R9784 gnd.n5798 gnd.n1772 19.3944
R9785 gnd.n5798 gnd.n1762 19.3944
R9786 gnd.n5811 gnd.n1762 19.3944
R9787 gnd.n5811 gnd.n1760 19.3944
R9788 gnd.n5815 gnd.n1760 19.3944
R9789 gnd.n5815 gnd.n1750 19.3944
R9790 gnd.n5828 gnd.n1750 19.3944
R9791 gnd.n5828 gnd.n1748 19.3944
R9792 gnd.n5832 gnd.n1748 19.3944
R9793 gnd.n5832 gnd.n1738 19.3944
R9794 gnd.n5845 gnd.n1738 19.3944
R9795 gnd.n5845 gnd.n1736 19.3944
R9796 gnd.n5851 gnd.n1736 19.3944
R9797 gnd.n5851 gnd.n5850 19.3944
R9798 gnd.n5850 gnd.n1726 19.3944
R9799 gnd.n5865 gnd.n1726 19.3944
R9800 gnd.n5865 gnd.n1724 19.3944
R9801 gnd.n5869 gnd.n1724 19.3944
R9802 gnd.n5869 gnd.n1723 19.3944
R9803 gnd.n6032 gnd.n1723 19.3944
R9804 gnd.n6032 gnd.n1721 19.3944
R9805 gnd.n6038 gnd.n1721 19.3944
R9806 gnd.n6038 gnd.n6037 19.3944
R9807 gnd.n6037 gnd.n1673 19.3944
R9808 gnd.n6064 gnd.n1673 19.3944
R9809 gnd.n6064 gnd.n1671 19.3944
R9810 gnd.n6070 gnd.n1671 19.3944
R9811 gnd.n6070 gnd.n6069 19.3944
R9812 gnd.n6069 gnd.n1647 19.3944
R9813 gnd.n6097 gnd.n1647 19.3944
R9814 gnd.n6097 gnd.n1645 19.3944
R9815 gnd.n6103 gnd.n1645 19.3944
R9816 gnd.n6103 gnd.n6102 19.3944
R9817 gnd.n6102 gnd.n1619 19.3944
R9818 gnd.n6128 gnd.n1619 19.3944
R9819 gnd.n6128 gnd.n1617 19.3944
R9820 gnd.n6141 gnd.n1617 19.3944
R9821 gnd.n6141 gnd.n6140 19.3944
R9822 gnd.n6140 gnd.n6139 19.3944
R9823 gnd.n6139 gnd.n6136 19.3944
R9824 gnd.n6136 gnd.n1581 19.3944
R9825 gnd.n6209 gnd.n1581 19.3944
R9826 gnd.n6209 gnd.n6208 19.3944
R9827 gnd.n6208 gnd.n6207 19.3944
R9828 gnd.n6207 gnd.n1586 19.3944
R9829 gnd.n1586 gnd.n1546 19.3944
R9830 gnd.n6245 gnd.n1546 19.3944
R9831 gnd.n6245 gnd.n1544 19.3944
R9832 gnd.n6250 gnd.n1544 19.3944
R9833 gnd.n6250 gnd.n1542 19.3944
R9834 gnd.n6254 gnd.n1542 19.3944
R9835 gnd.n6257 gnd.n6256 19.3944
R9836 gnd.n6261 gnd.n6260 19.3944
R9837 gnd.n6282 gnd.n6281 19.3944
R9838 gnd.n6279 gnd.n6263 19.3944
R9839 gnd.n6275 gnd.n6274 19.3944
R9840 gnd.n6274 gnd.n6273 19.3944
R9841 gnd.n6273 gnd.n6270 19.3944
R9842 gnd.n6270 gnd.n404 19.3944
R9843 gnd.n7621 gnd.n404 19.3944
R9844 gnd.n7621 gnd.n7620 19.3944
R9845 gnd.n7620 gnd.n7619 19.3944
R9846 gnd.n7619 gnd.n408 19.3944
R9847 gnd.n7615 gnd.n408 19.3944
R9848 gnd.n7615 gnd.n7614 19.3944
R9849 gnd.n4198 gnd.n4195 19.3944
R9850 gnd.n4198 gnd.n4194 19.3944
R9851 gnd.n4202 gnd.n4194 19.3944
R9852 gnd.n4202 gnd.n4192 19.3944
R9853 gnd.n4208 gnd.n4192 19.3944
R9854 gnd.n4208 gnd.n4190 19.3944
R9855 gnd.n4212 gnd.n4190 19.3944
R9856 gnd.n4212 gnd.n4188 19.3944
R9857 gnd.n4218 gnd.n4188 19.3944
R9858 gnd.n4218 gnd.n4186 19.3944
R9859 gnd.n4222 gnd.n4186 19.3944
R9860 gnd.n4222 gnd.n4184 19.3944
R9861 gnd.n4228 gnd.n4184 19.3944
R9862 gnd.n4228 gnd.n4182 19.3944
R9863 gnd.n4232 gnd.n4182 19.3944
R9864 gnd.n4232 gnd.n4177 19.3944
R9865 gnd.n4238 gnd.n4177 19.3944
R9866 gnd.n4242 gnd.n4175 19.3944
R9867 gnd.n4242 gnd.n4173 19.3944
R9868 gnd.n4248 gnd.n4173 19.3944
R9869 gnd.n4248 gnd.n4171 19.3944
R9870 gnd.n4252 gnd.n4171 19.3944
R9871 gnd.n4252 gnd.n4169 19.3944
R9872 gnd.n4258 gnd.n4169 19.3944
R9873 gnd.n4258 gnd.n4167 19.3944
R9874 gnd.n4262 gnd.n4167 19.3944
R9875 gnd.n4262 gnd.n4165 19.3944
R9876 gnd.n4268 gnd.n4165 19.3944
R9877 gnd.n4268 gnd.n4163 19.3944
R9878 gnd.n4272 gnd.n4163 19.3944
R9879 gnd.n4272 gnd.n4161 19.3944
R9880 gnd.n4278 gnd.n4161 19.3944
R9881 gnd.n4278 gnd.n4159 19.3944
R9882 gnd.n4283 gnd.n4159 19.3944
R9883 gnd.n4283 gnd.n4157 19.3944
R9884 gnd.n4440 gnd.n2665 19.3944
R9885 gnd.n4452 gnd.n2665 19.3944
R9886 gnd.n4452 gnd.n2663 19.3944
R9887 gnd.n4456 gnd.n2663 19.3944
R9888 gnd.n4456 gnd.n2649 19.3944
R9889 gnd.n4468 gnd.n2649 19.3944
R9890 gnd.n4468 gnd.n2647 19.3944
R9891 gnd.n4472 gnd.n2647 19.3944
R9892 gnd.n4472 gnd.n2633 19.3944
R9893 gnd.n4484 gnd.n2633 19.3944
R9894 gnd.n4484 gnd.n2631 19.3944
R9895 gnd.n4498 gnd.n2631 19.3944
R9896 gnd.n4498 gnd.n4497 19.3944
R9897 gnd.n4497 gnd.n4496 19.3944
R9898 gnd.n4496 gnd.n4495 19.3944
R9899 gnd.n4495 gnd.n4493 19.3944
R9900 gnd.n4493 gnd.n1038 19.3944
R9901 gnd.n6699 gnd.n1038 19.3944
R9902 gnd.n6699 gnd.n6698 19.3944
R9903 gnd.n6698 gnd.n6697 19.3944
R9904 gnd.n6697 gnd.n1042 19.3944
R9905 gnd.n6687 gnd.n1042 19.3944
R9906 gnd.n6687 gnd.n6686 19.3944
R9907 gnd.n6686 gnd.n6685 19.3944
R9908 gnd.n6685 gnd.n1063 19.3944
R9909 gnd.n6675 gnd.n1063 19.3944
R9910 gnd.n6675 gnd.n6674 19.3944
R9911 gnd.n6674 gnd.n6673 19.3944
R9912 gnd.n6673 gnd.n1084 19.3944
R9913 gnd.n4588 gnd.n1084 19.3944
R9914 gnd.n4588 gnd.n4587 19.3944
R9915 gnd.n4587 gnd.n2540 19.3944
R9916 gnd.n4618 gnd.n2540 19.3944
R9917 gnd.n4618 gnd.n2538 19.3944
R9918 gnd.n4623 gnd.n2538 19.3944
R9919 gnd.n4623 gnd.n1107 19.3944
R9920 gnd.n6661 gnd.n1107 19.3944
R9921 gnd.n6661 gnd.n6660 19.3944
R9922 gnd.n6660 gnd.n6659 19.3944
R9923 gnd.n6659 gnd.n1111 19.3944
R9924 gnd.n6649 gnd.n1111 19.3944
R9925 gnd.n6649 gnd.n6648 19.3944
R9926 gnd.n6648 gnd.n6647 19.3944
R9927 gnd.n6647 gnd.n1131 19.3944
R9928 gnd.n6637 gnd.n1131 19.3944
R9929 gnd.n6637 gnd.n6636 19.3944
R9930 gnd.n6636 gnd.n6635 19.3944
R9931 gnd.n6635 gnd.n1153 19.3944
R9932 gnd.n6625 gnd.n1153 19.3944
R9933 gnd.n6625 gnd.n6624 19.3944
R9934 gnd.n6624 gnd.n6623 19.3944
R9935 gnd.n6623 gnd.n1174 19.3944
R9936 gnd.n6613 gnd.n1174 19.3944
R9937 gnd.n6613 gnd.n6612 19.3944
R9938 gnd.n6612 gnd.n6611 19.3944
R9939 gnd.n6611 gnd.n1196 19.3944
R9940 gnd.n6601 gnd.n1196 19.3944
R9941 gnd.n6601 gnd.n6600 19.3944
R9942 gnd.n6600 gnd.n6599 19.3944
R9943 gnd.n6599 gnd.n1217 19.3944
R9944 gnd.n6589 gnd.n1217 19.3944
R9945 gnd.n6589 gnd.n6588 19.3944
R9946 gnd.n6588 gnd.n6587 19.3944
R9947 gnd.n6587 gnd.n1239 19.3944
R9948 gnd.n4437 gnd.n4436 19.3944
R9949 gnd.n4436 gnd.n4328 19.3944
R9950 gnd.n4430 gnd.n4328 19.3944
R9951 gnd.n4430 gnd.n4429 19.3944
R9952 gnd.n4429 gnd.n4428 19.3944
R9953 gnd.n4428 gnd.n4334 19.3944
R9954 gnd.n4422 gnd.n4334 19.3944
R9955 gnd.n4422 gnd.n4421 19.3944
R9956 gnd.n4421 gnd.n4420 19.3944
R9957 gnd.n4420 gnd.n4340 19.3944
R9958 gnd.n4414 gnd.n4340 19.3944
R9959 gnd.n4414 gnd.n4413 19.3944
R9960 gnd.n4413 gnd.n4412 19.3944
R9961 gnd.n4412 gnd.n4346 19.3944
R9962 gnd.n4406 gnd.n4346 19.3944
R9963 gnd.n4406 gnd.n4405 19.3944
R9964 gnd.n4396 gnd.n4395 19.3944
R9965 gnd.n4395 gnd.n4393 19.3944
R9966 gnd.n4393 gnd.n4392 19.3944
R9967 gnd.n4392 gnd.n4390 19.3944
R9968 gnd.n4390 gnd.n4389 19.3944
R9969 gnd.n4389 gnd.n4387 19.3944
R9970 gnd.n4387 gnd.n4386 19.3944
R9971 gnd.n4386 gnd.n4384 19.3944
R9972 gnd.n4384 gnd.n4383 19.3944
R9973 gnd.n4383 gnd.n4381 19.3944
R9974 gnd.n4381 gnd.n4380 19.3944
R9975 gnd.n4380 gnd.n4378 19.3944
R9976 gnd.n4378 gnd.n4377 19.3944
R9977 gnd.n4377 gnd.n4375 19.3944
R9978 gnd.n4375 gnd.n4374 19.3944
R9979 gnd.n4374 gnd.n4372 19.3944
R9980 gnd.n4372 gnd.n4371 19.3944
R9981 gnd.n4371 gnd.n2612 19.3944
R9982 gnd.n4523 gnd.n2612 19.3944
R9983 gnd.n4523 gnd.n2610 19.3944
R9984 gnd.n4527 gnd.n2610 19.3944
R9985 gnd.n4527 gnd.n2582 19.3944
R9986 gnd.n4544 gnd.n2582 19.3944
R9987 gnd.n4544 gnd.n2580 19.3944
R9988 gnd.n4549 gnd.n2580 19.3944
R9989 gnd.n4549 gnd.n2557 19.3944
R9990 gnd.n4571 gnd.n2557 19.3944
R9991 gnd.n4572 gnd.n4571 19.3944
R9992 gnd.n4572 gnd.n2555 19.3944
R9993 gnd.n4580 gnd.n2555 19.3944
R9994 gnd.n4580 gnd.n4579 19.3944
R9995 gnd.n4579 gnd.n4578 19.3944
R9996 gnd.n4578 gnd.n2531 19.3944
R9997 gnd.n4632 gnd.n2531 19.3944
R9998 gnd.n4632 gnd.n2529 19.3944
R9999 gnd.n4636 gnd.n2529 19.3944
R10000 gnd.n4636 gnd.n2514 19.3944
R10001 gnd.n4674 gnd.n2514 19.3944
R10002 gnd.n4674 gnd.n2515 19.3944
R10003 gnd.n4670 gnd.n2515 19.3944
R10004 gnd.n4670 gnd.n4669 19.3944
R10005 gnd.n4669 gnd.n4668 19.3944
R10006 gnd.n4668 gnd.n2520 19.3944
R10007 gnd.n4664 gnd.n2520 19.3944
R10008 gnd.n4664 gnd.n2500 19.3944
R10009 gnd.n4715 gnd.n2500 19.3944
R10010 gnd.n4715 gnd.n2498 19.3944
R10011 gnd.n4719 gnd.n2498 19.3944
R10012 gnd.n4719 gnd.n2494 19.3944
R10013 gnd.n4731 gnd.n2494 19.3944
R10014 gnd.n4731 gnd.n2492 19.3944
R10015 gnd.n4735 gnd.n2492 19.3944
R10016 gnd.n4735 gnd.n2476 19.3944
R10017 gnd.n4886 gnd.n2476 19.3944
R10018 gnd.n4886 gnd.n2477 19.3944
R10019 gnd.n4882 gnd.n2477 19.3944
R10020 gnd.n4882 gnd.n4881 19.3944
R10021 gnd.n4881 gnd.n4880 19.3944
R10022 gnd.n4880 gnd.n2482 19.3944
R10023 gnd.n4876 gnd.n2482 19.3944
R10024 gnd.n4876 gnd.n4875 19.3944
R10025 gnd.n4875 gnd.n4874 19.3944
R10026 gnd.n4874 gnd.n4833 19.3944
R10027 gnd.n4833 gnd.n2459 19.3944
R10028 gnd.n4323 gnd.n4151 19.3944
R10029 gnd.n4323 gnd.n4152 19.3944
R10030 gnd.n4319 gnd.n4152 19.3944
R10031 gnd.n4319 gnd.n4317 19.3944
R10032 gnd.n4317 gnd.n4316 19.3944
R10033 gnd.n4316 gnd.n4314 19.3944
R10034 gnd.n4314 gnd.n4313 19.3944
R10035 gnd.n4313 gnd.n4311 19.3944
R10036 gnd.n4311 gnd.n4310 19.3944
R10037 gnd.n4310 gnd.n4308 19.3944
R10038 gnd.n4308 gnd.n4307 19.3944
R10039 gnd.n4307 gnd.n4305 19.3944
R10040 gnd.n4305 gnd.n4304 19.3944
R10041 gnd.n4304 gnd.n2615 19.3944
R10042 gnd.n4512 gnd.n2615 19.3944
R10043 gnd.n4513 gnd.n4512 19.3944
R10044 gnd.n4515 gnd.n4513 19.3944
R10045 gnd.n4515 gnd.n2613 19.3944
R10046 gnd.n4519 gnd.n2613 19.3944
R10047 gnd.n4519 gnd.n2585 19.3944
R10048 gnd.n4531 gnd.n2585 19.3944
R10049 gnd.n4531 gnd.n2583 19.3944
R10050 gnd.n4540 gnd.n2583 19.3944
R10051 gnd.n4540 gnd.n4539 19.3944
R10052 gnd.n4539 gnd.n4538 19.3944
R10053 gnd.n4538 gnd.n2558 19.3944
R10054 gnd.n4567 gnd.n2558 19.3944
R10055 gnd.n4567 gnd.n4566 19.3944
R10056 gnd.n4566 gnd.n4565 19.3944
R10057 gnd.n4565 gnd.n2573 19.3944
R10058 gnd.n2573 gnd.n2572 19.3944
R10059 gnd.n2572 gnd.n2570 19.3944
R10060 gnd.n2570 gnd.n2569 19.3944
R10061 gnd.n2569 gnd.n2568 19.3944
R10062 gnd.n2568 gnd.n2525 19.3944
R10063 gnd.n4640 gnd.n2525 19.3944
R10064 gnd.n4641 gnd.n4640 19.3944
R10065 gnd.n4642 gnd.n4641 19.3944
R10066 gnd.n4642 gnd.n2523 19.3944
R10067 gnd.n4648 gnd.n2523 19.3944
R10068 gnd.n4649 gnd.n4648 19.3944
R10069 gnd.n4652 gnd.n4649 19.3944
R10070 gnd.n4652 gnd.n2521 19.3944
R10071 gnd.n4660 gnd.n2521 19.3944
R10072 gnd.n4660 gnd.n4659 19.3944
R10073 gnd.n4659 gnd.n4658 19.3944
R10074 gnd.n4658 gnd.n2497 19.3944
R10075 gnd.n4723 gnd.n2497 19.3944
R10076 gnd.n4723 gnd.n2495 19.3944
R10077 gnd.n4727 gnd.n2495 19.3944
R10078 gnd.n4727 gnd.n2491 19.3944
R10079 gnd.n4739 gnd.n2491 19.3944
R10080 gnd.n4739 gnd.n2489 19.3944
R10081 gnd.n4743 gnd.n2489 19.3944
R10082 gnd.n4744 gnd.n4743 19.3944
R10083 gnd.n4747 gnd.n4744 19.3944
R10084 gnd.n4747 gnd.n2487 19.3944
R10085 gnd.n4753 gnd.n2487 19.3944
R10086 gnd.n4754 gnd.n4753 19.3944
R10087 gnd.n4757 gnd.n4754 19.3944
R10088 gnd.n4757 gnd.n2485 19.3944
R10089 gnd.n4829 gnd.n2485 19.3944
R10090 gnd.n4829 gnd.n4828 19.3944
R10091 gnd.n4828 gnd.n4827 19.3944
R10092 gnd.n4776 gnd.n1296 19.3944
R10093 gnd.n4780 gnd.n4776 19.3944
R10094 gnd.n4783 gnd.n4780 19.3944
R10095 gnd.n4786 gnd.n4783 19.3944
R10096 gnd.n4786 gnd.n4772 19.3944
R10097 gnd.n4790 gnd.n4772 19.3944
R10098 gnd.n4793 gnd.n4790 19.3944
R10099 gnd.n4796 gnd.n4793 19.3944
R10100 gnd.n4796 gnd.n4770 19.3944
R10101 gnd.n4800 gnd.n4770 19.3944
R10102 gnd.n4803 gnd.n4800 19.3944
R10103 gnd.n4806 gnd.n4803 19.3944
R10104 gnd.n4806 gnd.n4768 19.3944
R10105 gnd.n4810 gnd.n4768 19.3944
R10106 gnd.n4813 gnd.n4810 19.3944
R10107 gnd.n4816 gnd.n4813 19.3944
R10108 gnd.n4816 gnd.n4766 19.3944
R10109 gnd.n4821 gnd.n4766 19.3944
R10110 gnd.n6579 gnd.n1249 19.3944
R10111 gnd.n6574 gnd.n1249 19.3944
R10112 gnd.n6574 gnd.n6573 19.3944
R10113 gnd.n6573 gnd.n6572 19.3944
R10114 gnd.n6572 gnd.n6569 19.3944
R10115 gnd.n6569 gnd.n6568 19.3944
R10116 gnd.n6568 gnd.n6565 19.3944
R10117 gnd.n6565 gnd.n6564 19.3944
R10118 gnd.n6564 gnd.n6561 19.3944
R10119 gnd.n6561 gnd.n6560 19.3944
R10120 gnd.n6560 gnd.n6557 19.3944
R10121 gnd.n6557 gnd.n6556 19.3944
R10122 gnd.n6556 gnd.n6553 19.3944
R10123 gnd.n6553 gnd.n6552 19.3944
R10124 gnd.n6552 gnd.n6549 19.3944
R10125 gnd.n4444 gnd.n2670 19.3944
R10126 gnd.n4448 gnd.n2670 19.3944
R10127 gnd.n4448 gnd.n2657 19.3944
R10128 gnd.n4460 gnd.n2657 19.3944
R10129 gnd.n4460 gnd.n2655 19.3944
R10130 gnd.n4464 gnd.n2655 19.3944
R10131 gnd.n4464 gnd.n2640 19.3944
R10132 gnd.n4476 gnd.n2640 19.3944
R10133 gnd.n4476 gnd.n2638 19.3944
R10134 gnd.n4480 gnd.n2638 19.3944
R10135 gnd.n4480 gnd.n2624 19.3944
R10136 gnd.n4502 gnd.n2624 19.3944
R10137 gnd.n4502 gnd.n2622 19.3944
R10138 gnd.n4507 gnd.n2622 19.3944
R10139 gnd.n4507 gnd.n1026 19.3944
R10140 gnd.n6705 gnd.n1026 19.3944
R10141 gnd.n6705 gnd.n6704 19.3944
R10142 gnd.n6704 gnd.n6703 19.3944
R10143 gnd.n6703 gnd.n1030 19.3944
R10144 gnd.n6693 gnd.n1030 19.3944
R10145 gnd.n6693 gnd.n6692 19.3944
R10146 gnd.n6692 gnd.n6691 19.3944
R10147 gnd.n6691 gnd.n1052 19.3944
R10148 gnd.n6681 gnd.n1052 19.3944
R10149 gnd.n6681 gnd.n6680 19.3944
R10150 gnd.n6680 gnd.n6679 19.3944
R10151 gnd.n6679 gnd.n1074 19.3944
R10152 gnd.n6669 gnd.n6668 19.3944
R10153 gnd.n4592 gnd.n1091 19.3944
R10154 gnd.n4595 gnd.n4594 19.3944
R10155 gnd.n4628 gnd.n4627 19.3944
R10156 gnd.n6665 gnd.n1097 19.3944
R10157 gnd.n6665 gnd.n1098 19.3944
R10158 gnd.n6655 gnd.n1098 19.3944
R10159 gnd.n6655 gnd.n6654 19.3944
R10160 gnd.n6654 gnd.n6653 19.3944
R10161 gnd.n6653 gnd.n1120 19.3944
R10162 gnd.n6643 gnd.n1120 19.3944
R10163 gnd.n6643 gnd.n6642 19.3944
R10164 gnd.n6642 gnd.n6641 19.3944
R10165 gnd.n6641 gnd.n1142 19.3944
R10166 gnd.n6631 gnd.n1142 19.3944
R10167 gnd.n6631 gnd.n6630 19.3944
R10168 gnd.n6630 gnd.n6629 19.3944
R10169 gnd.n6629 gnd.n1163 19.3944
R10170 gnd.n6619 gnd.n1163 19.3944
R10171 gnd.n6619 gnd.n6618 19.3944
R10172 gnd.n6618 gnd.n6617 19.3944
R10173 gnd.n6617 gnd.n1185 19.3944
R10174 gnd.n6607 gnd.n1185 19.3944
R10175 gnd.n6607 gnd.n6606 19.3944
R10176 gnd.n6606 gnd.n6605 19.3944
R10177 gnd.n6605 gnd.n1206 19.3944
R10178 gnd.n6595 gnd.n1206 19.3944
R10179 gnd.n6595 gnd.n6594 19.3944
R10180 gnd.n6594 gnd.n6593 19.3944
R10181 gnd.n6593 gnd.n1228 19.3944
R10182 gnd.n6583 gnd.n1228 19.3944
R10183 gnd.n6583 gnd.n6582 19.3944
R10184 gnd.n6878 gnd.n851 19.3944
R10185 gnd.n6872 gnd.n851 19.3944
R10186 gnd.n6872 gnd.n6871 19.3944
R10187 gnd.n6871 gnd.n6870 19.3944
R10188 gnd.n6870 gnd.n858 19.3944
R10189 gnd.n6864 gnd.n858 19.3944
R10190 gnd.n6864 gnd.n6863 19.3944
R10191 gnd.n6863 gnd.n6862 19.3944
R10192 gnd.n6862 gnd.n866 19.3944
R10193 gnd.n6856 gnd.n866 19.3944
R10194 gnd.n6856 gnd.n6855 19.3944
R10195 gnd.n6855 gnd.n6854 19.3944
R10196 gnd.n6854 gnd.n874 19.3944
R10197 gnd.n6848 gnd.n874 19.3944
R10198 gnd.n6848 gnd.n6847 19.3944
R10199 gnd.n6847 gnd.n6846 19.3944
R10200 gnd.n6846 gnd.n882 19.3944
R10201 gnd.n6840 gnd.n882 19.3944
R10202 gnd.n6840 gnd.n6839 19.3944
R10203 gnd.n6839 gnd.n6838 19.3944
R10204 gnd.n6838 gnd.n890 19.3944
R10205 gnd.n6832 gnd.n890 19.3944
R10206 gnd.n6832 gnd.n6831 19.3944
R10207 gnd.n6831 gnd.n6830 19.3944
R10208 gnd.n6830 gnd.n898 19.3944
R10209 gnd.n6824 gnd.n898 19.3944
R10210 gnd.n6824 gnd.n6823 19.3944
R10211 gnd.n6823 gnd.n6822 19.3944
R10212 gnd.n6822 gnd.n906 19.3944
R10213 gnd.n6816 gnd.n906 19.3944
R10214 gnd.n6816 gnd.n6815 19.3944
R10215 gnd.n6815 gnd.n6814 19.3944
R10216 gnd.n6814 gnd.n914 19.3944
R10217 gnd.n6808 gnd.n914 19.3944
R10218 gnd.n6808 gnd.n6807 19.3944
R10219 gnd.n6807 gnd.n6806 19.3944
R10220 gnd.n6806 gnd.n922 19.3944
R10221 gnd.n6800 gnd.n922 19.3944
R10222 gnd.n6800 gnd.n6799 19.3944
R10223 gnd.n6799 gnd.n6798 19.3944
R10224 gnd.n6798 gnd.n930 19.3944
R10225 gnd.n6792 gnd.n930 19.3944
R10226 gnd.n6792 gnd.n6791 19.3944
R10227 gnd.n6791 gnd.n6790 19.3944
R10228 gnd.n6790 gnd.n938 19.3944
R10229 gnd.n6784 gnd.n938 19.3944
R10230 gnd.n6784 gnd.n6783 19.3944
R10231 gnd.n6783 gnd.n6782 19.3944
R10232 gnd.n6782 gnd.n946 19.3944
R10233 gnd.n6776 gnd.n946 19.3944
R10234 gnd.n6776 gnd.n6775 19.3944
R10235 gnd.n6775 gnd.n6774 19.3944
R10236 gnd.n6774 gnd.n954 19.3944
R10237 gnd.n6768 gnd.n954 19.3944
R10238 gnd.n6768 gnd.n6767 19.3944
R10239 gnd.n6767 gnd.n6766 19.3944
R10240 gnd.n6766 gnd.n962 19.3944
R10241 gnd.n6760 gnd.n962 19.3944
R10242 gnd.n6760 gnd.n6759 19.3944
R10243 gnd.n6759 gnd.n6758 19.3944
R10244 gnd.n6758 gnd.n970 19.3944
R10245 gnd.n6752 gnd.n970 19.3944
R10246 gnd.n6752 gnd.n6751 19.3944
R10247 gnd.n6751 gnd.n6750 19.3944
R10248 gnd.n6750 gnd.n978 19.3944
R10249 gnd.n6744 gnd.n978 19.3944
R10250 gnd.n6744 gnd.n6743 19.3944
R10251 gnd.n6743 gnd.n6742 19.3944
R10252 gnd.n6742 gnd.n986 19.3944
R10253 gnd.n6736 gnd.n986 19.3944
R10254 gnd.n6736 gnd.n6735 19.3944
R10255 gnd.n6735 gnd.n6734 19.3944
R10256 gnd.n6734 gnd.n994 19.3944
R10257 gnd.n6728 gnd.n994 19.3944
R10258 gnd.n6728 gnd.n6727 19.3944
R10259 gnd.n6727 gnd.n6726 19.3944
R10260 gnd.n6726 gnd.n1002 19.3944
R10261 gnd.n6720 gnd.n1002 19.3944
R10262 gnd.n6720 gnd.n6719 19.3944
R10263 gnd.n6719 gnd.n6718 19.3944
R10264 gnd.n6718 gnd.n1010 19.3944
R10265 gnd.n6712 gnd.n1010 19.3944
R10266 gnd.n6712 gnd.n6711 19.3944
R10267 gnd.n6711 gnd.n6710 19.3944
R10268 gnd.n2400 gnd.n2399 19.3944
R10269 gnd.n2399 gnd.n2398 19.3944
R10270 gnd.n2398 gnd.n2343 19.3944
R10271 gnd.n2394 gnd.n2343 19.3944
R10272 gnd.n2394 gnd.n2393 19.3944
R10273 gnd.n2393 gnd.n2392 19.3944
R10274 gnd.n2392 gnd.n2347 19.3944
R10275 gnd.n2388 gnd.n2347 19.3944
R10276 gnd.n2388 gnd.n2387 19.3944
R10277 gnd.n2387 gnd.n2386 19.3944
R10278 gnd.n2386 gnd.n2351 19.3944
R10279 gnd.n2382 gnd.n2351 19.3944
R10280 gnd.n2382 gnd.n2381 19.3944
R10281 gnd.n2381 gnd.n2380 19.3944
R10282 gnd.n2380 gnd.n2355 19.3944
R10283 gnd.n2376 gnd.n2355 19.3944
R10284 gnd.n2376 gnd.n2375 19.3944
R10285 gnd.n2375 gnd.n2374 19.3944
R10286 gnd.n2374 gnd.n2359 19.3944
R10287 gnd.n2370 gnd.n2359 19.3944
R10288 gnd.n2370 gnd.n2369 19.3944
R10289 gnd.n2369 gnd.n2368 19.3944
R10290 gnd.n2368 gnd.n2363 19.3944
R10291 gnd.n2364 gnd.n2363 19.3944
R10292 gnd.n2364 gnd.n2220 19.3944
R10293 gnd.n5096 gnd.n2220 19.3944
R10294 gnd.n5096 gnd.n2218 19.3944
R10295 gnd.n5100 gnd.n2218 19.3944
R10296 gnd.n5198 gnd.n5100 19.3944
R10297 gnd.n5199 gnd.n5198 19.3944
R10298 gnd.n5199 gnd.n2215 19.3944
R10299 gnd.n5239 gnd.n2215 19.3944
R10300 gnd.n5239 gnd.n2216 19.3944
R10301 gnd.n5235 gnd.n2216 19.3944
R10302 gnd.n5235 gnd.n5234 19.3944
R10303 gnd.n5234 gnd.n5233 19.3944
R10304 gnd.n5233 gnd.n5205 19.3944
R10305 gnd.n5229 gnd.n5205 19.3944
R10306 gnd.n5229 gnd.n5228 19.3944
R10307 gnd.n5228 gnd.n5227 19.3944
R10308 gnd.n5227 gnd.n5209 19.3944
R10309 gnd.n5223 gnd.n5209 19.3944
R10310 gnd.n5223 gnd.n5222 19.3944
R10311 gnd.n5222 gnd.n5221 19.3944
R10312 gnd.n5221 gnd.n5212 19.3944
R10313 gnd.n5217 gnd.n5212 19.3944
R10314 gnd.n5217 gnd.n5216 19.3944
R10315 gnd.n5216 gnd.n2120 19.3944
R10316 gnd.n5381 gnd.n2120 19.3944
R10317 gnd.n5381 gnd.n2117 19.3944
R10318 gnd.n5399 gnd.n2117 19.3944
R10319 gnd.n5399 gnd.n2118 19.3944
R10320 gnd.n5395 gnd.n2118 19.3944
R10321 gnd.n5395 gnd.n5394 19.3944
R10322 gnd.n5394 gnd.n5393 19.3944
R10323 gnd.n5393 gnd.n5388 19.3944
R10324 gnd.n5389 gnd.n5388 19.3944
R10325 gnd.n5389 gnd.n2067 19.3944
R10326 gnd.n5462 gnd.n2067 19.3944
R10327 gnd.n5462 gnd.n2065 19.3944
R10328 gnd.n5466 gnd.n2065 19.3944
R10329 gnd.n5467 gnd.n5466 19.3944
R10330 gnd.n5470 gnd.n5467 19.3944
R10331 gnd.n5470 gnd.n2062 19.3944
R10332 gnd.n5497 gnd.n2062 19.3944
R10333 gnd.n5497 gnd.n2063 19.3944
R10334 gnd.n5493 gnd.n2063 19.3944
R10335 gnd.n5493 gnd.n5492 19.3944
R10336 gnd.n5492 gnd.n5491 19.3944
R10337 gnd.n5491 gnd.n5476 19.3944
R10338 gnd.n5487 gnd.n5476 19.3944
R10339 gnd.n5487 gnd.n5486 19.3944
R10340 gnd.n5486 gnd.n5485 19.3944
R10341 gnd.n5485 gnd.n5480 19.3944
R10342 gnd.n5481 gnd.n5480 19.3944
R10343 gnd.n5481 gnd.n1791 19.3944
R10344 gnd.n5767 gnd.n1791 19.3944
R10345 gnd.n5767 gnd.n1789 19.3944
R10346 gnd.n5771 gnd.n1789 19.3944
R10347 gnd.n5771 gnd.n1780 19.3944
R10348 gnd.n5785 gnd.n1780 19.3944
R10349 gnd.n5785 gnd.n1778 19.3944
R10350 gnd.n5789 gnd.n1778 19.3944
R10351 gnd.n5789 gnd.n1768 19.3944
R10352 gnd.n5802 gnd.n1768 19.3944
R10353 gnd.n5802 gnd.n1766 19.3944
R10354 gnd.n5806 gnd.n1766 19.3944
R10355 gnd.n5806 gnd.n1756 19.3944
R10356 gnd.n5819 gnd.n1756 19.3944
R10357 gnd.n5819 gnd.n1754 19.3944
R10358 gnd.n5823 gnd.n1754 19.3944
R10359 gnd.n5823 gnd.n1743 19.3944
R10360 gnd.n5836 gnd.n1743 19.3944
R10361 gnd.n5836 gnd.n1741 19.3944
R10362 gnd.n5840 gnd.n1741 19.3944
R10363 gnd.n5840 gnd.n1732 19.3944
R10364 gnd.n5855 gnd.n1732 19.3944
R10365 gnd.n5855 gnd.n1730 19.3944
R10366 gnd.n5859 gnd.n1730 19.3944
R10367 gnd.n5859 gnd.n1477 19.3944
R10368 gnd.n6353 gnd.n1477 19.3944
R10369 gnd.n6020 gnd.n5886 19.3944
R10370 gnd.n6025 gnd.n5886 19.3944
R10371 gnd.n6025 gnd.n5887 19.3944
R10372 gnd.n5937 gnd.n5929 19.3944
R10373 gnd.n5940 gnd.n5937 19.3944
R10374 gnd.n5940 gnd.n5921 19.3944
R10375 gnd.n5949 gnd.n5921 19.3944
R10376 gnd.n5952 gnd.n5949 19.3944
R10377 gnd.n5952 gnd.n5917 19.3944
R10378 gnd.n5961 gnd.n5917 19.3944
R10379 gnd.n5964 gnd.n5961 19.3944
R10380 gnd.n5964 gnd.n5909 19.3944
R10381 gnd.n5973 gnd.n5909 19.3944
R10382 gnd.n5976 gnd.n5973 19.3944
R10383 gnd.n5976 gnd.n5905 19.3944
R10384 gnd.n5986 gnd.n5905 19.3944
R10385 gnd.n5989 gnd.n5986 19.3944
R10386 gnd.n5993 gnd.n5989 19.3944
R10387 gnd.n5993 gnd.n5992 19.3944
R10388 gnd.n5992 gnd.n5893 19.3944
R10389 gnd.n6002 gnd.n5893 19.3944
R10390 gnd.n6004 gnd.n6002 19.3944
R10391 gnd.n6007 gnd.n6004 19.3944
R10392 gnd.n6010 gnd.n6007 19.3944
R10393 gnd.n6010 gnd.n5891 19.3944
R10394 gnd.n6014 gnd.n5891 19.3944
R10395 gnd.n6017 gnd.n6014 19.3944
R10396 gnd.n5196 gnd.n1366 19.1199
R10397 gnd.n2144 gnd.n2139 19.1199
R10398 gnd.n2094 gnd.n2092 19.1199
R10399 gnd.n5591 gnd.n1997 19.1199
R10400 gnd.n3534 gnd.t11 18.8012
R10401 gnd.n3519 gnd.t265 18.8012
R10402 gnd.n3378 gnd.n3377 18.4825
R10403 gnd.n5574 gnd.t180 18.4825
R10404 gnd.n1984 gnd.n1835 18.4247
R10405 gnd.n6549 gnd.n6548 18.4247
R10406 gnd.n7808 gnd.n124 18.2308
R10407 gnd.n5997 gnd.n5996 18.2308
R10408 gnd.n4933 gnd.n2451 18.2308
R10409 gnd.n4405 gnd.n4352 18.2308
R10410 gnd.t10 gnd.n3058 18.1639
R10411 gnd.n6478 gnd.n6477 17.9517
R10412 gnd.n5683 gnd.n5682 17.9517
R10413 gnd.n5108 gnd.n1378 17.8452
R10414 gnd.n5367 gnd.n2134 17.8452
R10415 gnd.n5421 gnd.n2098 17.8452
R10416 gnd.n5573 gnd.n5572 17.8452
R10417 gnd.n3086 gnd.t13 17.5266
R10418 gnd.t286 gnd.n2195 17.2079
R10419 gnd.n5528 gnd.t283 17.2079
R10420 gnd.n3485 gnd.t96 16.8893
R10421 gnd.n5062 gnd.t309 16.8893
R10422 gnd.n5773 gnd.t68 16.8893
R10423 gnd.t104 gnd.n5287 16.5706
R10424 gnd.n2125 gnd.n2123 16.5706
R10425 gnd.n5402 gnd.n2108 16.5706
R10426 gnd.n2043 gnd.t73 16.5706
R10427 gnd.n5474 gnd.n2014 16.5706
R10428 gnd.n3313 gnd.t223 16.2519
R10429 gnd.n3013 gnd.t97 16.2519
R10430 gnd.n5306 gnd.t287 15.9333
R10431 gnd.n5508 gnd.t308 15.9333
R10432 gnd.n4000 gnd.n3998 15.6674
R10433 gnd.n3968 gnd.n3966 15.6674
R10434 gnd.n3936 gnd.n3934 15.6674
R10435 gnd.n3905 gnd.n3903 15.6674
R10436 gnd.n3873 gnd.n3871 15.6674
R10437 gnd.n3841 gnd.n3839 15.6674
R10438 gnd.n3809 gnd.n3807 15.6674
R10439 gnd.n3778 gnd.n3776 15.6674
R10440 gnd.n3304 gnd.t223 15.6146
R10441 gnd.t197 gnd.n2754 15.6146
R10442 gnd.t183 gnd.n2755 15.6146
R10443 gnd.n5246 gnd.n5245 15.296
R10444 gnd.n5263 gnd.n2204 15.296
R10445 gnd.n2164 gnd.t0 15.296
R10446 gnd.n5379 gnd.n2123 15.296
R10447 gnd.n5410 gnd.n2108 15.296
R10448 gnd.n5435 gnd.t3 15.296
R10449 gnd.n5539 gnd.n5538 15.296
R10450 gnd.n5559 gnd.n2014 15.296
R10451 gnd.n5599 gnd.n5598 15.0827
R10452 gnd.n1348 gnd.n1343 15.0481
R10453 gnd.n5609 gnd.n5608 15.0481
R10454 gnd.n3672 gnd.t134 14.9773
R10455 gnd.n2247 gnd.t309 14.9773
R10456 gnd.n5783 gnd.t68 14.9773
R10457 gnd.n5331 gnd.t311 14.6587
R10458 gnd.n5442 gnd.t24 14.6587
R10459 gnd.t352 gnd.n2798 14.34
R10460 gnd.n3750 gnd.t9 14.34
R10461 gnd.t81 gnd.n1057 14.34
R10462 gnd.n7623 gnd.t22 14.34
R10463 gnd.n5195 gnd.t201 14.0214
R10464 gnd.n6466 gnd.n1378 14.0214
R10465 gnd.n2195 gnd.n2187 14.0214
R10466 gnd.t70 gnd.n2131 14.0214
R10467 gnd.n5369 gnd.n5367 14.0214
R10468 gnd.n5421 gnd.n5420 14.0214
R10469 gnd.n2101 gnd.t65 14.0214
R10470 gnd.n5528 gnd.n2033 14.0214
R10471 gnd.n3460 gnd.t261 13.7027
R10472 gnd.n4582 gnd.t277 13.7027
R10473 gnd.t135 gnd.n5324 13.7027
R10474 gnd.n5451 gnd.t141 13.7027
R10475 gnd.t63 gnd.n339 13.7027
R10476 gnd.n3170 gnd.n3169 13.5763
R10477 gnd.n4114 gnd.n2711 13.5763
R10478 gnd.n1947 gnd.n1901 13.5763
R10479 gnd.n7846 gnd.n7845 13.5763
R10480 gnd.n4157 gnd.n4156 13.5763
R10481 gnd.n4822 gnd.n4821 13.5763
R10482 gnd.n3378 gnd.n3116 13.384
R10483 gnd.t105 gnd.n2122 13.384
R10484 gnd.n5409 gnd.t106 13.384
R10485 gnd.n1359 gnd.n1340 13.1884
R10486 gnd.n1354 gnd.n1353 13.1884
R10487 gnd.n1353 gnd.n1352 13.1884
R10488 gnd.n5602 gnd.n5597 13.1884
R10489 gnd.n5603 gnd.n5602 13.1884
R10490 gnd.n1355 gnd.n1342 13.146
R10491 gnd.n1351 gnd.n1342 13.146
R10492 gnd.n5601 gnd.n5600 13.146
R10493 gnd.n5601 gnd.n5596 13.146
R10494 gnd.n4677 gnd.t121 13.0654
R10495 gnd.t77 gnd.n1521 13.0654
R10496 gnd.n4001 gnd.n3997 12.8005
R10497 gnd.n3969 gnd.n3965 12.8005
R10498 gnd.n3937 gnd.n3933 12.8005
R10499 gnd.n3906 gnd.n3902 12.8005
R10500 gnd.n3874 gnd.n3870 12.8005
R10501 gnd.n3842 gnd.n3838 12.8005
R10502 gnd.n3810 gnd.n3806 12.8005
R10503 gnd.n3779 gnd.n3775 12.8005
R10504 gnd.n6472 gnd.n1366 12.7467
R10505 gnd.n2145 gnd.n2144 12.7467
R10506 gnd.n2092 gnd.n2087 12.7467
R10507 gnd.n5572 gnd.t173 12.7467
R10508 gnd.n2645 gnd.t33 12.4281
R10509 gnd.n4712 gnd.t31 12.4281
R10510 gnd.n6609 gnd.t83 12.4281
R10511 gnd.n5006 gnd.t354 12.4281
R10512 gnd.n1746 gnd.t149 12.4281
R10513 gnd.n1642 gnd.t291 12.4281
R10514 gnd.t47 gnd.n1574 12.4281
R10515 gnd.n7743 gnd.t117 12.4281
R10516 gnd.n3169 gnd.n3164 12.4126
R10517 gnd.n4117 gnd.n4114 12.4126
R10518 gnd.n1943 gnd.n1901 12.4126
R10519 gnd.n7845 gnd.n200 12.4126
R10520 gnd.n4290 gnd.n4156 12.4126
R10521 gnd.n4824 gnd.n4822 12.4126
R10522 gnd.n6541 gnd.n6478 12.1761
R10523 gnd.n5682 gnd.n5681 12.1761
R10524 gnd.n6577 gnd.n1251 12.1094
R10525 gnd.t227 gnd.n5590 12.1094
R10526 gnd.n6041 gnd.n6040 12.1094
R10527 gnd.n4005 gnd.n4004 12.0247
R10528 gnd.n3973 gnd.n3972 12.0247
R10529 gnd.n3941 gnd.n3940 12.0247
R10530 gnd.n3910 gnd.n3909 12.0247
R10531 gnd.n3878 gnd.n3877 12.0247
R10532 gnd.n3846 gnd.n3845 12.0247
R10533 gnd.n3814 gnd.n3813 12.0247
R10534 gnd.n3783 gnd.n3782 12.0247
R10535 gnd.n6708 gnd.n1019 11.7908
R10536 gnd.n6633 gnd.t31 11.7908
R10537 gnd.n4889 gnd.t83 11.7908
R10538 gnd.t291 gnd.n1630 11.7908
R10539 gnd.n6163 gnd.t47 11.7908
R10540 gnd.n7719 gnd.n259 11.7908
R10541 gnd.n5246 gnd.t214 11.4721
R10542 gnd.n5306 gnd.n2168 11.4721
R10543 gnd.n5325 gnd.n2150 11.4721
R10544 gnd.n5450 gnd.n2082 11.4721
R10545 gnd.n5508 gnd.n2048 11.4721
R10546 gnd.t211 gnd.n1799 11.4721
R10547 gnd.n5757 gnd.n1799 11.4721
R10548 gnd.n4008 gnd.n3995 11.249
R10549 gnd.n3976 gnd.n3963 11.249
R10550 gnd.n3944 gnd.n3931 11.249
R10551 gnd.n3913 gnd.n3900 11.249
R10552 gnd.n3881 gnd.n3868 11.249
R10553 gnd.n3849 gnd.n3836 11.249
R10554 gnd.n3817 gnd.n3804 11.249
R10555 gnd.n3786 gnd.n3773 11.249
R10556 gnd.n3448 gnd.t261 11.1535
R10557 gnd.n6657 gnd.t121 11.1535
R10558 gnd.n5287 gnd.t284 11.1535
R10559 gnd.t320 gnd.n2043 11.1535
R10560 gnd.n6195 gnd.t77 11.1535
R10561 gnd.n5752 gnd.n5751 10.6151
R10562 gnd.n5751 gnd.n5748 10.6151
R10563 gnd.n5746 gnd.n5743 10.6151
R10564 gnd.n5743 gnd.n5742 10.6151
R10565 gnd.n5742 gnd.n5739 10.6151
R10566 gnd.n5739 gnd.n5738 10.6151
R10567 gnd.n5738 gnd.n5735 10.6151
R10568 gnd.n5735 gnd.n5734 10.6151
R10569 gnd.n5734 gnd.n5731 10.6151
R10570 gnd.n5731 gnd.n5730 10.6151
R10571 gnd.n5730 gnd.n5727 10.6151
R10572 gnd.n5727 gnd.n5726 10.6151
R10573 gnd.n5726 gnd.n5723 10.6151
R10574 gnd.n5723 gnd.n5722 10.6151
R10575 gnd.n5722 gnd.n5719 10.6151
R10576 gnd.n5719 gnd.n5718 10.6151
R10577 gnd.n5718 gnd.n5715 10.6151
R10578 gnd.n5715 gnd.n5714 10.6151
R10579 gnd.n5714 gnd.n5711 10.6151
R10580 gnd.n5711 gnd.n5710 10.6151
R10581 gnd.n5710 gnd.n5707 10.6151
R10582 gnd.n5707 gnd.n5706 10.6151
R10583 gnd.n5706 gnd.n5703 10.6151
R10584 gnd.n5703 gnd.n5702 10.6151
R10585 gnd.n5702 gnd.n5699 10.6151
R10586 gnd.n5699 gnd.n5698 10.6151
R10587 gnd.n5698 gnd.n5695 10.6151
R10588 gnd.n5695 gnd.n5694 10.6151
R10589 gnd.n5694 gnd.n5691 10.6151
R10590 gnd.n5691 gnd.n5690 10.6151
R10591 gnd.n5178 gnd.n5177 10.6151
R10592 gnd.n5179 gnd.n5178 10.6151
R10593 gnd.n5181 gnd.n5179 10.6151
R10594 gnd.n5182 gnd.n5181 10.6151
R10595 gnd.n5184 gnd.n5182 10.6151
R10596 gnd.n5185 gnd.n5184 10.6151
R10597 gnd.n5186 gnd.n5185 10.6151
R10598 gnd.n5186 gnd.n2210 10.6151
R10599 gnd.n5248 gnd.n2210 10.6151
R10600 gnd.n5249 gnd.n5248 10.6151
R10601 gnd.n5254 gnd.n5249 10.6151
R10602 gnd.n5254 gnd.n5253 10.6151
R10603 gnd.n5253 gnd.n5252 10.6151
R10604 gnd.n5252 gnd.n5250 10.6151
R10605 gnd.n5250 gnd.n2185 10.6151
R10606 gnd.n5282 gnd.n2185 10.6151
R10607 gnd.n5283 gnd.n5282 10.6151
R10608 gnd.n5285 gnd.n5283 10.6151
R10609 gnd.n5285 gnd.n5284 10.6151
R10610 gnd.n5284 gnd.n2166 10.6151
R10611 gnd.n5308 gnd.n2166 10.6151
R10612 gnd.n5309 gnd.n5308 10.6151
R10613 gnd.n5312 gnd.n5309 10.6151
R10614 gnd.n5312 gnd.n5311 10.6151
R10615 gnd.n5311 gnd.n5310 10.6151
R10616 gnd.n5310 gnd.n2142 10.6151
R10617 gnd.n5333 gnd.n2142 10.6151
R10618 gnd.n5334 gnd.n5333 10.6151
R10619 gnd.n5354 gnd.n5334 10.6151
R10620 gnd.n5354 gnd.n5353 10.6151
R10621 gnd.n5353 gnd.n5352 10.6151
R10622 gnd.n5352 gnd.n5351 10.6151
R10623 gnd.n5351 gnd.n5335 10.6151
R10624 gnd.n5346 gnd.n5335 10.6151
R10625 gnd.n5346 gnd.n5345 10.6151
R10626 gnd.n5345 gnd.n5344 10.6151
R10627 gnd.n5344 gnd.n5343 10.6151
R10628 gnd.n5343 gnd.n5341 10.6151
R10629 gnd.n5341 gnd.n5340 10.6151
R10630 gnd.n5340 gnd.n5337 10.6151
R10631 gnd.n5337 gnd.n2090 10.6151
R10632 gnd.n5429 gnd.n2090 10.6151
R10633 gnd.n5430 gnd.n5429 10.6151
R10634 gnd.n5440 gnd.n5430 10.6151
R10635 gnd.n5440 gnd.n5439 10.6151
R10636 gnd.n5439 gnd.n5438 10.6151
R10637 gnd.n5438 gnd.n5437 10.6151
R10638 gnd.n5437 gnd.n5434 10.6151
R10639 gnd.n5434 gnd.n5433 10.6151
R10640 gnd.n5433 gnd.n5431 10.6151
R10641 gnd.n5431 gnd.n2040 10.6151
R10642 gnd.n5516 gnd.n2040 10.6151
R10643 gnd.n5517 gnd.n5516 10.6151
R10644 gnd.n5519 gnd.n5517 10.6151
R10645 gnd.n5519 gnd.n5518 10.6151
R10646 gnd.n5518 gnd.n2031 10.6151
R10647 gnd.n5531 gnd.n2031 10.6151
R10648 gnd.n5532 gnd.n5531 10.6151
R10649 gnd.n5536 gnd.n5532 10.6151
R10650 gnd.n5536 gnd.n5535 10.6151
R10651 gnd.n5535 gnd.n5534 10.6151
R10652 gnd.n5534 gnd.n2012 10.6151
R10653 gnd.n5562 gnd.n2012 10.6151
R10654 gnd.n5563 gnd.n5562 10.6151
R10655 gnd.n5570 gnd.n5563 10.6151
R10656 gnd.n5570 gnd.n5569 10.6151
R10657 gnd.n5569 gnd.n5568 10.6151
R10658 gnd.n5568 gnd.n5565 10.6151
R10659 gnd.n5565 gnd.n5564 10.6151
R10660 gnd.n5564 gnd.n1990 10.6151
R10661 gnd.n1990 gnd.n1988 10.6151
R10662 gnd.n5112 gnd.n1301 10.6151
R10663 gnd.n5115 gnd.n5112 10.6151
R10664 gnd.n5120 gnd.n5117 10.6151
R10665 gnd.n5121 gnd.n5120 10.6151
R10666 gnd.n5124 gnd.n5121 10.6151
R10667 gnd.n5125 gnd.n5124 10.6151
R10668 gnd.n5128 gnd.n5125 10.6151
R10669 gnd.n5129 gnd.n5128 10.6151
R10670 gnd.n5132 gnd.n5129 10.6151
R10671 gnd.n5133 gnd.n5132 10.6151
R10672 gnd.n5136 gnd.n5133 10.6151
R10673 gnd.n5137 gnd.n5136 10.6151
R10674 gnd.n5140 gnd.n5137 10.6151
R10675 gnd.n5141 gnd.n5140 10.6151
R10676 gnd.n5144 gnd.n5141 10.6151
R10677 gnd.n5145 gnd.n5144 10.6151
R10678 gnd.n5148 gnd.n5145 10.6151
R10679 gnd.n5149 gnd.n5148 10.6151
R10680 gnd.n5152 gnd.n5149 10.6151
R10681 gnd.n5153 gnd.n5152 10.6151
R10682 gnd.n5156 gnd.n5153 10.6151
R10683 gnd.n5157 gnd.n5156 10.6151
R10684 gnd.n5160 gnd.n5157 10.6151
R10685 gnd.n5161 gnd.n5160 10.6151
R10686 gnd.n5164 gnd.n5161 10.6151
R10687 gnd.n5165 gnd.n5164 10.6151
R10688 gnd.n5168 gnd.n5165 10.6151
R10689 gnd.n5169 gnd.n5168 10.6151
R10690 gnd.n5172 gnd.n5169 10.6151
R10691 gnd.n5173 gnd.n5172 10.6151
R10692 gnd.n6541 gnd.n6540 10.6151
R10693 gnd.n6540 gnd.n6539 10.6151
R10694 gnd.n6539 gnd.n6538 10.6151
R10695 gnd.n6538 gnd.n6536 10.6151
R10696 gnd.n6536 gnd.n6533 10.6151
R10697 gnd.n6533 gnd.n6532 10.6151
R10698 gnd.n6532 gnd.n6529 10.6151
R10699 gnd.n6529 gnd.n6528 10.6151
R10700 gnd.n6528 gnd.n6525 10.6151
R10701 gnd.n6525 gnd.n6524 10.6151
R10702 gnd.n6524 gnd.n6521 10.6151
R10703 gnd.n6521 gnd.n6520 10.6151
R10704 gnd.n6520 gnd.n6517 10.6151
R10705 gnd.n6517 gnd.n6516 10.6151
R10706 gnd.n6516 gnd.n6513 10.6151
R10707 gnd.n6513 gnd.n6512 10.6151
R10708 gnd.n6512 gnd.n6509 10.6151
R10709 gnd.n6509 gnd.n6508 10.6151
R10710 gnd.n6508 gnd.n6505 10.6151
R10711 gnd.n6505 gnd.n6504 10.6151
R10712 gnd.n6504 gnd.n6501 10.6151
R10713 gnd.n6501 gnd.n6500 10.6151
R10714 gnd.n6500 gnd.n6497 10.6151
R10715 gnd.n6497 gnd.n6496 10.6151
R10716 gnd.n6496 gnd.n6493 10.6151
R10717 gnd.n6493 gnd.n6492 10.6151
R10718 gnd.n6492 gnd.n6489 10.6151
R10719 gnd.n6489 gnd.n6488 10.6151
R10720 gnd.n6485 gnd.n6484 10.6151
R10721 gnd.n6484 gnd.n1302 10.6151
R10722 gnd.n5681 gnd.n5679 10.6151
R10723 gnd.n5679 gnd.n5676 10.6151
R10724 gnd.n5676 gnd.n5675 10.6151
R10725 gnd.n5675 gnd.n5672 10.6151
R10726 gnd.n5672 gnd.n5671 10.6151
R10727 gnd.n5671 gnd.n5668 10.6151
R10728 gnd.n5668 gnd.n5667 10.6151
R10729 gnd.n5667 gnd.n5664 10.6151
R10730 gnd.n5664 gnd.n5663 10.6151
R10731 gnd.n5663 gnd.n5660 10.6151
R10732 gnd.n5660 gnd.n5659 10.6151
R10733 gnd.n5659 gnd.n5656 10.6151
R10734 gnd.n5656 gnd.n5655 10.6151
R10735 gnd.n5655 gnd.n5652 10.6151
R10736 gnd.n5652 gnd.n5651 10.6151
R10737 gnd.n5651 gnd.n5648 10.6151
R10738 gnd.n5648 gnd.n5647 10.6151
R10739 gnd.n5647 gnd.n5644 10.6151
R10740 gnd.n5644 gnd.n5643 10.6151
R10741 gnd.n5643 gnd.n5640 10.6151
R10742 gnd.n5640 gnd.n5639 10.6151
R10743 gnd.n5639 gnd.n5636 10.6151
R10744 gnd.n5636 gnd.n5635 10.6151
R10745 gnd.n5635 gnd.n5632 10.6151
R10746 gnd.n5632 gnd.n5631 10.6151
R10747 gnd.n5631 gnd.n5628 10.6151
R10748 gnd.n5628 gnd.n5627 10.6151
R10749 gnd.n5627 gnd.n5624 10.6151
R10750 gnd.n5622 gnd.n5619 10.6151
R10751 gnd.n5619 gnd.n5618 10.6151
R10752 gnd.n6477 gnd.n6476 10.6151
R10753 gnd.n6476 gnd.n1360 10.6151
R10754 gnd.n5104 gnd.n1360 10.6151
R10755 gnd.n5193 gnd.n5104 10.6151
R10756 gnd.n5193 gnd.n5192 10.6151
R10757 gnd.n5192 gnd.n5191 10.6151
R10758 gnd.n5191 gnd.n5105 10.6151
R10759 gnd.n5106 gnd.n5105 10.6151
R10760 gnd.n5106 gnd.n2206 10.6151
R10761 gnd.n5259 gnd.n2206 10.6151
R10762 gnd.n5260 gnd.n5259 10.6151
R10763 gnd.n5261 gnd.n5260 10.6151
R10764 gnd.n5261 gnd.n2190 10.6151
R10765 gnd.n5275 gnd.n2190 10.6151
R10766 gnd.n5276 gnd.n5275 10.6151
R10767 gnd.n5278 gnd.n5276 10.6151
R10768 gnd.n5278 gnd.n5277 10.6151
R10769 gnd.n5277 gnd.n2171 10.6151
R10770 gnd.n5300 gnd.n2171 10.6151
R10771 gnd.n5301 gnd.n5300 10.6151
R10772 gnd.n5304 gnd.n5301 10.6151
R10773 gnd.n5304 gnd.n5303 10.6151
R10774 gnd.n5303 gnd.n5302 10.6151
R10775 gnd.n5302 gnd.n2147 10.6151
R10776 gnd.n5327 gnd.n2147 10.6151
R10777 gnd.n5328 gnd.n5327 10.6151
R10778 gnd.n5329 gnd.n5328 10.6151
R10779 gnd.n5329 gnd.n2137 10.6151
R10780 gnd.n5358 gnd.n2137 10.6151
R10781 gnd.n5359 gnd.n5358 10.6151
R10782 gnd.n5365 gnd.n5359 10.6151
R10783 gnd.n5365 gnd.n5364 10.6151
R10784 gnd.n5364 gnd.n5363 10.6151
R10785 gnd.n5363 gnd.n5360 10.6151
R10786 gnd.n5360 gnd.n2112 10.6151
R10787 gnd.n5405 gnd.n2112 10.6151
R10788 gnd.n5406 gnd.n5405 10.6151
R10789 gnd.n5407 gnd.n5406 10.6151
R10790 gnd.n5407 gnd.n2096 10.6151
R10791 gnd.n5423 gnd.n2096 10.6151
R10792 gnd.n5424 gnd.n5423 10.6151
R10793 gnd.n5425 gnd.n5424 10.6151
R10794 gnd.n5425 gnd.n2085 10.6151
R10795 gnd.n5444 gnd.n2085 10.6151
R10796 gnd.n5445 gnd.n5444 10.6151
R10797 gnd.n5448 gnd.n5445 10.6151
R10798 gnd.n5448 gnd.n5447 10.6151
R10799 gnd.n5447 gnd.n5446 10.6151
R10800 gnd.n5446 gnd.n2046 10.6151
R10801 gnd.n5510 gnd.n2046 10.6151
R10802 gnd.n5511 gnd.n5510 10.6151
R10803 gnd.n5512 gnd.n5511 10.6151
R10804 gnd.n5512 gnd.n2035 10.6151
R10805 gnd.n5524 gnd.n2035 10.6151
R10806 gnd.n5525 gnd.n5524 10.6151
R10807 gnd.n5526 gnd.n5525 10.6151
R10808 gnd.n5526 gnd.n2026 10.6151
R10809 gnd.n5542 gnd.n2026 10.6151
R10810 gnd.n5543 gnd.n5542 10.6151
R10811 gnd.n5547 gnd.n5543 10.6151
R10812 gnd.n5547 gnd.n5546 10.6151
R10813 gnd.n5546 gnd.n5545 10.6151
R10814 gnd.n5545 gnd.n2008 10.6151
R10815 gnd.n5576 gnd.n2008 10.6151
R10816 gnd.n5577 gnd.n5576 10.6151
R10817 gnd.n5578 gnd.n5577 10.6151
R10818 gnd.n5578 gnd.n1995 10.6151
R10819 gnd.n5593 gnd.n1995 10.6151
R10820 gnd.n5594 gnd.n5593 10.6151
R10821 gnd.n5684 gnd.n5594 10.6151
R10822 gnd.n5684 gnd.n5683 10.6151
R10823 gnd.n3367 gnd.t306 10.5161
R10824 gnd.n2800 gnd.t352 10.5161
R10825 gnd.n3733 gnd.t9 10.5161
R10826 gnd.t277 gnd.n2548 10.5161
R10827 gnd.n5264 gnd.t71 10.5161
R10828 gnd.n5551 gnd.t263 10.5161
R10829 gnd.n1537 gnd.t63 10.5161
R10830 gnd.n4009 gnd.n3993 10.4732
R10831 gnd.n3977 gnd.n3961 10.4732
R10832 gnd.n3945 gnd.n3929 10.4732
R10833 gnd.n3914 gnd.n3898 10.4732
R10834 gnd.n3882 gnd.n3866 10.4732
R10835 gnd.n3850 gnd.n3834 10.4732
R10836 gnd.n3818 gnd.n3802 10.4732
R10837 gnd.n3787 gnd.n3771 10.4732
R10838 gnd.n2168 gnd.n2160 10.1975
R10839 gnd.n2164 gnd.n2150 10.1975
R10840 gnd.n5435 gnd.n2082 10.1975
R10841 gnd.n2071 gnd.n2048 10.1975
R10842 gnd.t134 gnd.n2817 9.87883
R10843 gnd.n4542 gnd.t81 9.87883
R10844 gnd.n7687 gnd.t22 9.87883
R10845 gnd.n7971 gnd.n78 9.81789
R10846 gnd.n4013 gnd.n4012 9.69747
R10847 gnd.n3981 gnd.n3980 9.69747
R10848 gnd.n3949 gnd.n3948 9.69747
R10849 gnd.n3918 gnd.n3917 9.69747
R10850 gnd.n3886 gnd.n3885 9.69747
R10851 gnd.n3854 gnd.n3853 9.69747
R10852 gnd.n3822 gnd.n3821 9.69747
R10853 gnd.n3791 gnd.n3790 9.69747
R10854 gnd.n2340 gnd.n2337 9.45751
R10855 gnd.n6350 gnd.n1480 9.45599
R10856 gnd.n4019 gnd.n4018 9.45567
R10857 gnd.n3987 gnd.n3986 9.45567
R10858 gnd.n3955 gnd.n3954 9.45567
R10859 gnd.n3924 gnd.n3923 9.45567
R10860 gnd.n3892 gnd.n3891 9.45567
R10861 gnd.n3860 gnd.n3859 9.45567
R10862 gnd.n3828 gnd.n3827 9.45567
R10863 gnd.n3797 gnd.n3796 9.45567
R10864 gnd.n2965 gnd.n2964 9.39724
R10865 gnd.n4018 gnd.n4017 9.3005
R10866 gnd.n3991 gnd.n3990 9.3005
R10867 gnd.n4012 gnd.n4011 9.3005
R10868 gnd.n4010 gnd.n4009 9.3005
R10869 gnd.n3995 gnd.n3994 9.3005
R10870 gnd.n4004 gnd.n4003 9.3005
R10871 gnd.n4002 gnd.n4001 9.3005
R10872 gnd.n3986 gnd.n3985 9.3005
R10873 gnd.n3959 gnd.n3958 9.3005
R10874 gnd.n3980 gnd.n3979 9.3005
R10875 gnd.n3978 gnd.n3977 9.3005
R10876 gnd.n3963 gnd.n3962 9.3005
R10877 gnd.n3972 gnd.n3971 9.3005
R10878 gnd.n3970 gnd.n3969 9.3005
R10879 gnd.n3954 gnd.n3953 9.3005
R10880 gnd.n3927 gnd.n3926 9.3005
R10881 gnd.n3948 gnd.n3947 9.3005
R10882 gnd.n3946 gnd.n3945 9.3005
R10883 gnd.n3931 gnd.n3930 9.3005
R10884 gnd.n3940 gnd.n3939 9.3005
R10885 gnd.n3938 gnd.n3937 9.3005
R10886 gnd.n3923 gnd.n3922 9.3005
R10887 gnd.n3896 gnd.n3895 9.3005
R10888 gnd.n3917 gnd.n3916 9.3005
R10889 gnd.n3915 gnd.n3914 9.3005
R10890 gnd.n3900 gnd.n3899 9.3005
R10891 gnd.n3909 gnd.n3908 9.3005
R10892 gnd.n3907 gnd.n3906 9.3005
R10893 gnd.n3891 gnd.n3890 9.3005
R10894 gnd.n3864 gnd.n3863 9.3005
R10895 gnd.n3885 gnd.n3884 9.3005
R10896 gnd.n3883 gnd.n3882 9.3005
R10897 gnd.n3868 gnd.n3867 9.3005
R10898 gnd.n3877 gnd.n3876 9.3005
R10899 gnd.n3875 gnd.n3874 9.3005
R10900 gnd.n3859 gnd.n3858 9.3005
R10901 gnd.n3832 gnd.n3831 9.3005
R10902 gnd.n3853 gnd.n3852 9.3005
R10903 gnd.n3851 gnd.n3850 9.3005
R10904 gnd.n3836 gnd.n3835 9.3005
R10905 gnd.n3845 gnd.n3844 9.3005
R10906 gnd.n3843 gnd.n3842 9.3005
R10907 gnd.n3827 gnd.n3826 9.3005
R10908 gnd.n3800 gnd.n3799 9.3005
R10909 gnd.n3821 gnd.n3820 9.3005
R10910 gnd.n3819 gnd.n3818 9.3005
R10911 gnd.n3804 gnd.n3803 9.3005
R10912 gnd.n3813 gnd.n3812 9.3005
R10913 gnd.n3811 gnd.n3810 9.3005
R10914 gnd.n3796 gnd.n3795 9.3005
R10915 gnd.n3769 gnd.n3768 9.3005
R10916 gnd.n3790 gnd.n3789 9.3005
R10917 gnd.n3788 gnd.n3787 9.3005
R10918 gnd.n3773 gnd.n3772 9.3005
R10919 gnd.n3782 gnd.n3781 9.3005
R10920 gnd.n3780 gnd.n3779 9.3005
R10921 gnd.n4144 gnd.n4143 9.3005
R10922 gnd.n4142 gnd.n2699 9.3005
R10923 gnd.n4141 gnd.n4140 9.3005
R10924 gnd.n4137 gnd.n2700 9.3005
R10925 gnd.n4134 gnd.n2701 9.3005
R10926 gnd.n4133 gnd.n2702 9.3005
R10927 gnd.n4130 gnd.n2703 9.3005
R10928 gnd.n4129 gnd.n2704 9.3005
R10929 gnd.n4126 gnd.n2705 9.3005
R10930 gnd.n4125 gnd.n2706 9.3005
R10931 gnd.n4122 gnd.n2707 9.3005
R10932 gnd.n4121 gnd.n2708 9.3005
R10933 gnd.n4118 gnd.n2709 9.3005
R10934 gnd.n4117 gnd.n2710 9.3005
R10935 gnd.n4114 gnd.n4113 9.3005
R10936 gnd.n4112 gnd.n2711 9.3005
R10937 gnd.n4145 gnd.n2698 9.3005
R10938 gnd.n3386 gnd.n3385 9.3005
R10939 gnd.n3090 gnd.n3089 9.3005
R10940 gnd.n3413 gnd.n3412 9.3005
R10941 gnd.n3414 gnd.n3088 9.3005
R10942 gnd.n3418 gnd.n3415 9.3005
R10943 gnd.n3417 gnd.n3416 9.3005
R10944 gnd.n3062 gnd.n3061 9.3005
R10945 gnd.n3443 gnd.n3442 9.3005
R10946 gnd.n3444 gnd.n3060 9.3005
R10947 gnd.n3446 gnd.n3445 9.3005
R10948 gnd.n3040 gnd.n3039 9.3005
R10949 gnd.n3474 gnd.n3473 9.3005
R10950 gnd.n3475 gnd.n3038 9.3005
R10951 gnd.n3483 gnd.n3476 9.3005
R10952 gnd.n3482 gnd.n3477 9.3005
R10953 gnd.n3481 gnd.n3479 9.3005
R10954 gnd.n3478 gnd.n2987 9.3005
R10955 gnd.n3531 gnd.n2988 9.3005
R10956 gnd.n3530 gnd.n2989 9.3005
R10957 gnd.n3529 gnd.n2990 9.3005
R10958 gnd.n3009 gnd.n2991 9.3005
R10959 gnd.n3011 gnd.n3010 9.3005
R10960 gnd.n2897 gnd.n2896 9.3005
R10961 gnd.n3569 gnd.n3568 9.3005
R10962 gnd.n3570 gnd.n2895 9.3005
R10963 gnd.n3574 gnd.n3571 9.3005
R10964 gnd.n3573 gnd.n3572 9.3005
R10965 gnd.n2870 gnd.n2869 9.3005
R10966 gnd.n3609 gnd.n3608 9.3005
R10967 gnd.n3610 gnd.n2868 9.3005
R10968 gnd.n3614 gnd.n3611 9.3005
R10969 gnd.n3613 gnd.n3612 9.3005
R10970 gnd.n2843 gnd.n2842 9.3005
R10971 gnd.n3654 gnd.n3653 9.3005
R10972 gnd.n3655 gnd.n2841 9.3005
R10973 gnd.n3659 gnd.n3656 9.3005
R10974 gnd.n3658 gnd.n3657 9.3005
R10975 gnd.n2815 gnd.n2814 9.3005
R10976 gnd.n3694 gnd.n3693 9.3005
R10977 gnd.n3695 gnd.n2813 9.3005
R10978 gnd.n3699 gnd.n3696 9.3005
R10979 gnd.n3698 gnd.n3697 9.3005
R10980 gnd.n2787 gnd.n2786 9.3005
R10981 gnd.n3743 gnd.n3742 9.3005
R10982 gnd.n3744 gnd.n2785 9.3005
R10983 gnd.n3748 gnd.n3745 9.3005
R10984 gnd.n3747 gnd.n3746 9.3005
R10985 gnd.n2760 gnd.n2759 9.3005
R10986 gnd.n4037 gnd.n4036 9.3005
R10987 gnd.n4038 gnd.n2758 9.3005
R10988 gnd.n4044 gnd.n4039 9.3005
R10989 gnd.n4043 gnd.n4040 9.3005
R10990 gnd.n4042 gnd.n4041 9.3005
R10991 gnd.n3387 gnd.n3384 9.3005
R10992 gnd.n3169 gnd.n3128 9.3005
R10993 gnd.n3164 gnd.n3163 9.3005
R10994 gnd.n3162 gnd.n3129 9.3005
R10995 gnd.n3161 gnd.n3160 9.3005
R10996 gnd.n3157 gnd.n3130 9.3005
R10997 gnd.n3154 gnd.n3153 9.3005
R10998 gnd.n3152 gnd.n3131 9.3005
R10999 gnd.n3151 gnd.n3150 9.3005
R11000 gnd.n3147 gnd.n3132 9.3005
R11001 gnd.n3144 gnd.n3143 9.3005
R11002 gnd.n3142 gnd.n3133 9.3005
R11003 gnd.n3141 gnd.n3140 9.3005
R11004 gnd.n3137 gnd.n3135 9.3005
R11005 gnd.n3134 gnd.n3114 9.3005
R11006 gnd.n3381 gnd.n3113 9.3005
R11007 gnd.n3383 gnd.n3382 9.3005
R11008 gnd.n3171 gnd.n3170 9.3005
R11009 gnd.n3394 gnd.n3100 9.3005
R11010 gnd.n3401 gnd.n3101 9.3005
R11011 gnd.n3403 gnd.n3402 9.3005
R11012 gnd.n3404 gnd.n3081 9.3005
R11013 gnd.n3423 gnd.n3422 9.3005
R11014 gnd.n3425 gnd.n3073 9.3005
R11015 gnd.n3432 gnd.n3075 9.3005
R11016 gnd.n3433 gnd.n3070 9.3005
R11017 gnd.n3435 gnd.n3434 9.3005
R11018 gnd.n3071 gnd.n3056 9.3005
R11019 gnd.n3451 gnd.n3054 9.3005
R11020 gnd.n3455 gnd.n3454 9.3005
R11021 gnd.n3453 gnd.n3030 9.3005
R11022 gnd.n3490 gnd.n3029 9.3005
R11023 gnd.n3493 gnd.n3492 9.3005
R11024 gnd.n3026 gnd.n3025 9.3005
R11025 gnd.n3499 gnd.n3027 9.3005
R11026 gnd.n3501 gnd.n3500 9.3005
R11027 gnd.n3503 gnd.n3024 9.3005
R11028 gnd.n3506 gnd.n3505 9.3005
R11029 gnd.n3509 gnd.n3507 9.3005
R11030 gnd.n3511 gnd.n3510 9.3005
R11031 gnd.n3517 gnd.n3512 9.3005
R11032 gnd.n3516 gnd.n3515 9.3005
R11033 gnd.n2888 gnd.n2887 9.3005
R11034 gnd.n3583 gnd.n3582 9.3005
R11035 gnd.n3584 gnd.n2881 9.3005
R11036 gnd.n3592 gnd.n2880 9.3005
R11037 gnd.n3595 gnd.n3594 9.3005
R11038 gnd.n3597 gnd.n3596 9.3005
R11039 gnd.n3600 gnd.n2863 9.3005
R11040 gnd.n3598 gnd.n2861 9.3005
R11041 gnd.n3620 gnd.n2859 9.3005
R11042 gnd.n3622 gnd.n3621 9.3005
R11043 gnd.n2833 gnd.n2832 9.3005
R11044 gnd.n3668 gnd.n3667 9.3005
R11045 gnd.n3669 gnd.n2826 9.3005
R11046 gnd.n3677 gnd.n2825 9.3005
R11047 gnd.n3680 gnd.n3679 9.3005
R11048 gnd.n3682 gnd.n3681 9.3005
R11049 gnd.n3685 gnd.n2808 9.3005
R11050 gnd.n3683 gnd.n2806 9.3005
R11051 gnd.n3705 gnd.n2804 9.3005
R11052 gnd.n3707 gnd.n3706 9.3005
R11053 gnd.n2778 gnd.n2777 9.3005
R11054 gnd.n3757 gnd.n3756 9.3005
R11055 gnd.n3758 gnd.n2771 9.3005
R11056 gnd.n3766 gnd.n2770 9.3005
R11057 gnd.n4025 gnd.n4024 9.3005
R11058 gnd.n4027 gnd.n4026 9.3005
R11059 gnd.n4028 gnd.n2751 9.3005
R11060 gnd.n4052 gnd.n4051 9.3005
R11061 gnd.n2752 gnd.n2714 9.3005
R11062 gnd.n3392 gnd.n3391 9.3005
R11063 gnd.n4108 gnd.n2715 9.3005
R11064 gnd.n4107 gnd.n2717 9.3005
R11065 gnd.n4104 gnd.n2718 9.3005
R11066 gnd.n4103 gnd.n2719 9.3005
R11067 gnd.n4100 gnd.n2720 9.3005
R11068 gnd.n4099 gnd.n2721 9.3005
R11069 gnd.n4096 gnd.n2722 9.3005
R11070 gnd.n4095 gnd.n2723 9.3005
R11071 gnd.n4092 gnd.n2724 9.3005
R11072 gnd.n4091 gnd.n2725 9.3005
R11073 gnd.n4088 gnd.n2726 9.3005
R11074 gnd.n4087 gnd.n2727 9.3005
R11075 gnd.n4084 gnd.n2728 9.3005
R11076 gnd.n4083 gnd.n2729 9.3005
R11077 gnd.n4080 gnd.n2730 9.3005
R11078 gnd.n4079 gnd.n2731 9.3005
R11079 gnd.n4076 gnd.n2732 9.3005
R11080 gnd.n4075 gnd.n2733 9.3005
R11081 gnd.n4072 gnd.n2734 9.3005
R11082 gnd.n4071 gnd.n2735 9.3005
R11083 gnd.n4068 gnd.n2736 9.3005
R11084 gnd.n4067 gnd.n2737 9.3005
R11085 gnd.n4064 gnd.n2741 9.3005
R11086 gnd.n4063 gnd.n2742 9.3005
R11087 gnd.n4060 gnd.n2743 9.3005
R11088 gnd.n4059 gnd.n2744 9.3005
R11089 gnd.n4110 gnd.n4109 9.3005
R11090 gnd.n3561 gnd.n3545 9.3005
R11091 gnd.n3560 gnd.n3546 9.3005
R11092 gnd.n3559 gnd.n3547 9.3005
R11093 gnd.n3557 gnd.n3548 9.3005
R11094 gnd.n3556 gnd.n3549 9.3005
R11095 gnd.n3554 gnd.n3550 9.3005
R11096 gnd.n3553 gnd.n3551 9.3005
R11097 gnd.n2851 gnd.n2850 9.3005
R11098 gnd.n3630 gnd.n3629 9.3005
R11099 gnd.n3631 gnd.n2849 9.3005
R11100 gnd.n3648 gnd.n3632 9.3005
R11101 gnd.n3647 gnd.n3633 9.3005
R11102 gnd.n3646 gnd.n3634 9.3005
R11103 gnd.n3644 gnd.n3635 9.3005
R11104 gnd.n3643 gnd.n3636 9.3005
R11105 gnd.n3641 gnd.n3637 9.3005
R11106 gnd.n3640 gnd.n3638 9.3005
R11107 gnd.n2795 gnd.n2794 9.3005
R11108 gnd.n3715 gnd.n3714 9.3005
R11109 gnd.n3716 gnd.n2793 9.3005
R11110 gnd.n3737 gnd.n3717 9.3005
R11111 gnd.n3736 gnd.n3718 9.3005
R11112 gnd.n3735 gnd.n3719 9.3005
R11113 gnd.n3732 gnd.n3720 9.3005
R11114 gnd.n3731 gnd.n3721 9.3005
R11115 gnd.n3729 gnd.n3722 9.3005
R11116 gnd.n3728 gnd.n3723 9.3005
R11117 gnd.n3726 gnd.n3725 9.3005
R11118 gnd.n3724 gnd.n2746 9.3005
R11119 gnd.n3302 gnd.n3301 9.3005
R11120 gnd.n3192 gnd.n3191 9.3005
R11121 gnd.n3316 gnd.n3315 9.3005
R11122 gnd.n3317 gnd.n3190 9.3005
R11123 gnd.n3319 gnd.n3318 9.3005
R11124 gnd.n3180 gnd.n3179 9.3005
R11125 gnd.n3332 gnd.n3331 9.3005
R11126 gnd.n3333 gnd.n3178 9.3005
R11127 gnd.n3365 gnd.n3334 9.3005
R11128 gnd.n3364 gnd.n3335 9.3005
R11129 gnd.n3363 gnd.n3336 9.3005
R11130 gnd.n3362 gnd.n3337 9.3005
R11131 gnd.n3359 gnd.n3338 9.3005
R11132 gnd.n3358 gnd.n3339 9.3005
R11133 gnd.n3357 gnd.n3340 9.3005
R11134 gnd.n3355 gnd.n3341 9.3005
R11135 gnd.n3354 gnd.n3342 9.3005
R11136 gnd.n3351 gnd.n3343 9.3005
R11137 gnd.n3350 gnd.n3344 9.3005
R11138 gnd.n3349 gnd.n3345 9.3005
R11139 gnd.n3347 gnd.n3346 9.3005
R11140 gnd.n3046 gnd.n3045 9.3005
R11141 gnd.n3463 gnd.n3462 9.3005
R11142 gnd.n3464 gnd.n3044 9.3005
R11143 gnd.n3468 gnd.n3465 9.3005
R11144 gnd.n3467 gnd.n3466 9.3005
R11145 gnd.n2968 gnd.n2967 9.3005
R11146 gnd.n3543 gnd.n3542 9.3005
R11147 gnd.n3300 gnd.n3201 9.3005
R11148 gnd.n3203 gnd.n3202 9.3005
R11149 gnd.n3247 gnd.n3245 9.3005
R11150 gnd.n3248 gnd.n3244 9.3005
R11151 gnd.n3251 gnd.n3240 9.3005
R11152 gnd.n3252 gnd.n3239 9.3005
R11153 gnd.n3255 gnd.n3238 9.3005
R11154 gnd.n3256 gnd.n3237 9.3005
R11155 gnd.n3259 gnd.n3236 9.3005
R11156 gnd.n3260 gnd.n3235 9.3005
R11157 gnd.n3263 gnd.n3234 9.3005
R11158 gnd.n3264 gnd.n3233 9.3005
R11159 gnd.n3267 gnd.n3232 9.3005
R11160 gnd.n3268 gnd.n3231 9.3005
R11161 gnd.n3271 gnd.n3230 9.3005
R11162 gnd.n3272 gnd.n3229 9.3005
R11163 gnd.n3275 gnd.n3228 9.3005
R11164 gnd.n3276 gnd.n3227 9.3005
R11165 gnd.n3279 gnd.n3226 9.3005
R11166 gnd.n3280 gnd.n3225 9.3005
R11167 gnd.n3283 gnd.n3224 9.3005
R11168 gnd.n3284 gnd.n3223 9.3005
R11169 gnd.n3287 gnd.n3222 9.3005
R11170 gnd.n3289 gnd.n3221 9.3005
R11171 gnd.n3290 gnd.n3220 9.3005
R11172 gnd.n3291 gnd.n3219 9.3005
R11173 gnd.n3292 gnd.n3218 9.3005
R11174 gnd.n3299 gnd.n3298 9.3005
R11175 gnd.n3308 gnd.n3307 9.3005
R11176 gnd.n3309 gnd.n3195 9.3005
R11177 gnd.n3311 gnd.n3310 9.3005
R11178 gnd.n3186 gnd.n3185 9.3005
R11179 gnd.n3324 gnd.n3323 9.3005
R11180 gnd.n3325 gnd.n3184 9.3005
R11181 gnd.n3327 gnd.n3326 9.3005
R11182 gnd.n3173 gnd.n3172 9.3005
R11183 gnd.n3370 gnd.n3369 9.3005
R11184 gnd.n3371 gnd.n3127 9.3005
R11185 gnd.n3375 gnd.n3373 9.3005
R11186 gnd.n3374 gnd.n3106 9.3005
R11187 gnd.n3393 gnd.n3105 9.3005
R11188 gnd.n3396 gnd.n3395 9.3005
R11189 gnd.n3099 gnd.n3098 9.3005
R11190 gnd.n3407 gnd.n3405 9.3005
R11191 gnd.n3406 gnd.n3080 9.3005
R11192 gnd.n3424 gnd.n3079 9.3005
R11193 gnd.n3427 gnd.n3426 9.3005
R11194 gnd.n3074 gnd.n3069 9.3005
R11195 gnd.n3437 gnd.n3436 9.3005
R11196 gnd.n3072 gnd.n3052 9.3005
R11197 gnd.n3458 gnd.n3053 9.3005
R11198 gnd.n3457 gnd.n3456 9.3005
R11199 gnd.n3055 gnd.n3031 9.3005
R11200 gnd.n3489 gnd.n3488 9.3005
R11201 gnd.n3491 gnd.n2976 9.3005
R11202 gnd.n3538 gnd.n2977 9.3005
R11203 gnd.n3537 gnd.n2978 9.3005
R11204 gnd.n3536 gnd.n2979 9.3005
R11205 gnd.n3502 gnd.n2980 9.3005
R11206 gnd.n3504 gnd.n2998 9.3005
R11207 gnd.n3524 gnd.n2999 9.3005
R11208 gnd.n3523 gnd.n3000 9.3005
R11209 gnd.n3522 gnd.n3001 9.3005
R11210 gnd.n3513 gnd.n3002 9.3005
R11211 gnd.n3514 gnd.n2889 9.3005
R11212 gnd.n3580 gnd.n3579 9.3005
R11213 gnd.n3581 gnd.n2882 9.3005
R11214 gnd.n3591 gnd.n3590 9.3005
R11215 gnd.n3593 gnd.n2878 9.3005
R11216 gnd.n3603 gnd.n2879 9.3005
R11217 gnd.n3602 gnd.n3601 9.3005
R11218 gnd.n3599 gnd.n2857 9.3005
R11219 gnd.n3625 gnd.n2858 9.3005
R11220 gnd.n3624 gnd.n3623 9.3005
R11221 gnd.n2860 gnd.n2834 9.3005
R11222 gnd.n3665 gnd.n3664 9.3005
R11223 gnd.n3666 gnd.n2827 9.3005
R11224 gnd.n3676 gnd.n3675 9.3005
R11225 gnd.n3678 gnd.n2823 9.3005
R11226 gnd.n3688 gnd.n2824 9.3005
R11227 gnd.n3687 gnd.n3686 9.3005
R11228 gnd.n3684 gnd.n2802 9.3005
R11229 gnd.n3710 gnd.n2803 9.3005
R11230 gnd.n3709 gnd.n3708 9.3005
R11231 gnd.n2805 gnd.n2779 9.3005
R11232 gnd.n3754 gnd.n3753 9.3005
R11233 gnd.n3755 gnd.n2772 9.3005
R11234 gnd.n3765 gnd.n3764 9.3005
R11235 gnd.n4023 gnd.n2768 9.3005
R11236 gnd.n4031 gnd.n2769 9.3005
R11237 gnd.n4030 gnd.n4029 9.3005
R11238 gnd.n2750 gnd.n2749 9.3005
R11239 gnd.n4054 gnd.n4053 9.3005
R11240 gnd.n3197 gnd.n3196 9.3005
R11241 gnd.n6880 gnd.n849 9.3005
R11242 gnd.n6882 gnd.n6881 9.3005
R11243 gnd.n845 gnd.n844 9.3005
R11244 gnd.n6889 gnd.n6888 9.3005
R11245 gnd.n6890 gnd.n843 9.3005
R11246 gnd.n6892 gnd.n6891 9.3005
R11247 gnd.n839 gnd.n838 9.3005
R11248 gnd.n6899 gnd.n6898 9.3005
R11249 gnd.n6900 gnd.n837 9.3005
R11250 gnd.n6902 gnd.n6901 9.3005
R11251 gnd.n833 gnd.n832 9.3005
R11252 gnd.n6909 gnd.n6908 9.3005
R11253 gnd.n6910 gnd.n831 9.3005
R11254 gnd.n6912 gnd.n6911 9.3005
R11255 gnd.n827 gnd.n826 9.3005
R11256 gnd.n6919 gnd.n6918 9.3005
R11257 gnd.n6920 gnd.n825 9.3005
R11258 gnd.n6922 gnd.n6921 9.3005
R11259 gnd.n821 gnd.n820 9.3005
R11260 gnd.n6929 gnd.n6928 9.3005
R11261 gnd.n6930 gnd.n819 9.3005
R11262 gnd.n6932 gnd.n6931 9.3005
R11263 gnd.n815 gnd.n814 9.3005
R11264 gnd.n6939 gnd.n6938 9.3005
R11265 gnd.n6940 gnd.n813 9.3005
R11266 gnd.n6942 gnd.n6941 9.3005
R11267 gnd.n809 gnd.n808 9.3005
R11268 gnd.n6949 gnd.n6948 9.3005
R11269 gnd.n6950 gnd.n807 9.3005
R11270 gnd.n6952 gnd.n6951 9.3005
R11271 gnd.n803 gnd.n802 9.3005
R11272 gnd.n6959 gnd.n6958 9.3005
R11273 gnd.n6960 gnd.n801 9.3005
R11274 gnd.n6962 gnd.n6961 9.3005
R11275 gnd.n797 gnd.n796 9.3005
R11276 gnd.n6969 gnd.n6968 9.3005
R11277 gnd.n6970 gnd.n795 9.3005
R11278 gnd.n6972 gnd.n6971 9.3005
R11279 gnd.n791 gnd.n790 9.3005
R11280 gnd.n6979 gnd.n6978 9.3005
R11281 gnd.n6980 gnd.n789 9.3005
R11282 gnd.n6982 gnd.n6981 9.3005
R11283 gnd.n785 gnd.n784 9.3005
R11284 gnd.n6989 gnd.n6988 9.3005
R11285 gnd.n6990 gnd.n783 9.3005
R11286 gnd.n6992 gnd.n6991 9.3005
R11287 gnd.n779 gnd.n778 9.3005
R11288 gnd.n6999 gnd.n6998 9.3005
R11289 gnd.n7000 gnd.n777 9.3005
R11290 gnd.n7002 gnd.n7001 9.3005
R11291 gnd.n773 gnd.n772 9.3005
R11292 gnd.n7009 gnd.n7008 9.3005
R11293 gnd.n7010 gnd.n771 9.3005
R11294 gnd.n7012 gnd.n7011 9.3005
R11295 gnd.n767 gnd.n766 9.3005
R11296 gnd.n7019 gnd.n7018 9.3005
R11297 gnd.n7020 gnd.n765 9.3005
R11298 gnd.n7022 gnd.n7021 9.3005
R11299 gnd.n761 gnd.n760 9.3005
R11300 gnd.n7029 gnd.n7028 9.3005
R11301 gnd.n7030 gnd.n759 9.3005
R11302 gnd.n7032 gnd.n7031 9.3005
R11303 gnd.n755 gnd.n754 9.3005
R11304 gnd.n7039 gnd.n7038 9.3005
R11305 gnd.n7040 gnd.n753 9.3005
R11306 gnd.n7042 gnd.n7041 9.3005
R11307 gnd.n749 gnd.n748 9.3005
R11308 gnd.n7049 gnd.n7048 9.3005
R11309 gnd.n7050 gnd.n747 9.3005
R11310 gnd.n7052 gnd.n7051 9.3005
R11311 gnd.n743 gnd.n742 9.3005
R11312 gnd.n7059 gnd.n7058 9.3005
R11313 gnd.n7060 gnd.n741 9.3005
R11314 gnd.n7062 gnd.n7061 9.3005
R11315 gnd.n737 gnd.n736 9.3005
R11316 gnd.n7069 gnd.n7068 9.3005
R11317 gnd.n7070 gnd.n735 9.3005
R11318 gnd.n7072 gnd.n7071 9.3005
R11319 gnd.n731 gnd.n730 9.3005
R11320 gnd.n7079 gnd.n7078 9.3005
R11321 gnd.n7080 gnd.n729 9.3005
R11322 gnd.n7082 gnd.n7081 9.3005
R11323 gnd.n725 gnd.n724 9.3005
R11324 gnd.n7089 gnd.n7088 9.3005
R11325 gnd.n7090 gnd.n723 9.3005
R11326 gnd.n7092 gnd.n7091 9.3005
R11327 gnd.n719 gnd.n718 9.3005
R11328 gnd.n7099 gnd.n7098 9.3005
R11329 gnd.n7100 gnd.n717 9.3005
R11330 gnd.n7102 gnd.n7101 9.3005
R11331 gnd.n713 gnd.n712 9.3005
R11332 gnd.n7109 gnd.n7108 9.3005
R11333 gnd.n7110 gnd.n711 9.3005
R11334 gnd.n7112 gnd.n7111 9.3005
R11335 gnd.n707 gnd.n706 9.3005
R11336 gnd.n7119 gnd.n7118 9.3005
R11337 gnd.n7120 gnd.n705 9.3005
R11338 gnd.n7122 gnd.n7121 9.3005
R11339 gnd.n701 gnd.n700 9.3005
R11340 gnd.n7129 gnd.n7128 9.3005
R11341 gnd.n7130 gnd.n699 9.3005
R11342 gnd.n7132 gnd.n7131 9.3005
R11343 gnd.n695 gnd.n694 9.3005
R11344 gnd.n7139 gnd.n7138 9.3005
R11345 gnd.n7140 gnd.n693 9.3005
R11346 gnd.n7142 gnd.n7141 9.3005
R11347 gnd.n689 gnd.n688 9.3005
R11348 gnd.n7149 gnd.n7148 9.3005
R11349 gnd.n7150 gnd.n687 9.3005
R11350 gnd.n7152 gnd.n7151 9.3005
R11351 gnd.n683 gnd.n682 9.3005
R11352 gnd.n7159 gnd.n7158 9.3005
R11353 gnd.n7160 gnd.n681 9.3005
R11354 gnd.n7162 gnd.n7161 9.3005
R11355 gnd.n677 gnd.n676 9.3005
R11356 gnd.n7169 gnd.n7168 9.3005
R11357 gnd.n7170 gnd.n675 9.3005
R11358 gnd.n7172 gnd.n7171 9.3005
R11359 gnd.n671 gnd.n670 9.3005
R11360 gnd.n7179 gnd.n7178 9.3005
R11361 gnd.n7180 gnd.n669 9.3005
R11362 gnd.n7182 gnd.n7181 9.3005
R11363 gnd.n665 gnd.n664 9.3005
R11364 gnd.n7189 gnd.n7188 9.3005
R11365 gnd.n7190 gnd.n663 9.3005
R11366 gnd.n7192 gnd.n7191 9.3005
R11367 gnd.n659 gnd.n658 9.3005
R11368 gnd.n7199 gnd.n7198 9.3005
R11369 gnd.n7200 gnd.n657 9.3005
R11370 gnd.n7202 gnd.n7201 9.3005
R11371 gnd.n653 gnd.n652 9.3005
R11372 gnd.n7209 gnd.n7208 9.3005
R11373 gnd.n7210 gnd.n651 9.3005
R11374 gnd.n7212 gnd.n7211 9.3005
R11375 gnd.n647 gnd.n646 9.3005
R11376 gnd.n7219 gnd.n7218 9.3005
R11377 gnd.n7220 gnd.n645 9.3005
R11378 gnd.n7222 gnd.n7221 9.3005
R11379 gnd.n641 gnd.n640 9.3005
R11380 gnd.n7229 gnd.n7228 9.3005
R11381 gnd.n7230 gnd.n639 9.3005
R11382 gnd.n7232 gnd.n7231 9.3005
R11383 gnd.n635 gnd.n634 9.3005
R11384 gnd.n7239 gnd.n7238 9.3005
R11385 gnd.n7240 gnd.n633 9.3005
R11386 gnd.n7242 gnd.n7241 9.3005
R11387 gnd.n629 gnd.n628 9.3005
R11388 gnd.n7249 gnd.n7248 9.3005
R11389 gnd.n7250 gnd.n627 9.3005
R11390 gnd.n7252 gnd.n7251 9.3005
R11391 gnd.n623 gnd.n622 9.3005
R11392 gnd.n7259 gnd.n7258 9.3005
R11393 gnd.n7260 gnd.n621 9.3005
R11394 gnd.n7262 gnd.n7261 9.3005
R11395 gnd.n617 gnd.n616 9.3005
R11396 gnd.n7269 gnd.n7268 9.3005
R11397 gnd.n7270 gnd.n615 9.3005
R11398 gnd.n7272 gnd.n7271 9.3005
R11399 gnd.n611 gnd.n610 9.3005
R11400 gnd.n7279 gnd.n7278 9.3005
R11401 gnd.n7280 gnd.n609 9.3005
R11402 gnd.n7282 gnd.n7281 9.3005
R11403 gnd.n605 gnd.n604 9.3005
R11404 gnd.n7289 gnd.n7288 9.3005
R11405 gnd.n7290 gnd.n603 9.3005
R11406 gnd.n7292 gnd.n7291 9.3005
R11407 gnd.n599 gnd.n598 9.3005
R11408 gnd.n7299 gnd.n7298 9.3005
R11409 gnd.n7300 gnd.n597 9.3005
R11410 gnd.n7302 gnd.n7301 9.3005
R11411 gnd.n593 gnd.n592 9.3005
R11412 gnd.n7309 gnd.n7308 9.3005
R11413 gnd.n7310 gnd.n591 9.3005
R11414 gnd.n7312 gnd.n7311 9.3005
R11415 gnd.n587 gnd.n586 9.3005
R11416 gnd.n7319 gnd.n7318 9.3005
R11417 gnd.n7320 gnd.n585 9.3005
R11418 gnd.n7322 gnd.n7321 9.3005
R11419 gnd.n581 gnd.n580 9.3005
R11420 gnd.n7329 gnd.n7328 9.3005
R11421 gnd.n7330 gnd.n579 9.3005
R11422 gnd.n7332 gnd.n7331 9.3005
R11423 gnd.n575 gnd.n574 9.3005
R11424 gnd.n7339 gnd.n7338 9.3005
R11425 gnd.n7340 gnd.n573 9.3005
R11426 gnd.n7342 gnd.n7341 9.3005
R11427 gnd.n569 gnd.n568 9.3005
R11428 gnd.n7349 gnd.n7348 9.3005
R11429 gnd.n7350 gnd.n567 9.3005
R11430 gnd.n7352 gnd.n7351 9.3005
R11431 gnd.n563 gnd.n562 9.3005
R11432 gnd.n7359 gnd.n7358 9.3005
R11433 gnd.n7360 gnd.n561 9.3005
R11434 gnd.n7362 gnd.n7361 9.3005
R11435 gnd.n557 gnd.n556 9.3005
R11436 gnd.n7369 gnd.n7368 9.3005
R11437 gnd.n7370 gnd.n555 9.3005
R11438 gnd.n7372 gnd.n7371 9.3005
R11439 gnd.n551 gnd.n550 9.3005
R11440 gnd.n7379 gnd.n7378 9.3005
R11441 gnd.n7380 gnd.n549 9.3005
R11442 gnd.n7382 gnd.n7381 9.3005
R11443 gnd.n545 gnd.n544 9.3005
R11444 gnd.n7389 gnd.n7388 9.3005
R11445 gnd.n7390 gnd.n543 9.3005
R11446 gnd.n7392 gnd.n7391 9.3005
R11447 gnd.n539 gnd.n538 9.3005
R11448 gnd.n7399 gnd.n7398 9.3005
R11449 gnd.n7402 gnd.n7401 9.3005
R11450 gnd.n533 gnd.n532 9.3005
R11451 gnd.n7409 gnd.n7408 9.3005
R11452 gnd.n7410 gnd.n531 9.3005
R11453 gnd.n7412 gnd.n7411 9.3005
R11454 gnd.n527 gnd.n526 9.3005
R11455 gnd.n7419 gnd.n7418 9.3005
R11456 gnd.n7420 gnd.n525 9.3005
R11457 gnd.n7422 gnd.n7421 9.3005
R11458 gnd.n521 gnd.n520 9.3005
R11459 gnd.n7429 gnd.n7428 9.3005
R11460 gnd.n7430 gnd.n519 9.3005
R11461 gnd.n7432 gnd.n7431 9.3005
R11462 gnd.n515 gnd.n514 9.3005
R11463 gnd.n7439 gnd.n7438 9.3005
R11464 gnd.n7440 gnd.n513 9.3005
R11465 gnd.n7442 gnd.n7441 9.3005
R11466 gnd.n509 gnd.n508 9.3005
R11467 gnd.n7449 gnd.n7448 9.3005
R11468 gnd.n7450 gnd.n507 9.3005
R11469 gnd.n7452 gnd.n7451 9.3005
R11470 gnd.n503 gnd.n502 9.3005
R11471 gnd.n7459 gnd.n7458 9.3005
R11472 gnd.n7460 gnd.n501 9.3005
R11473 gnd.n7462 gnd.n7461 9.3005
R11474 gnd.n497 gnd.n496 9.3005
R11475 gnd.n7469 gnd.n7468 9.3005
R11476 gnd.n7470 gnd.n495 9.3005
R11477 gnd.n7472 gnd.n7471 9.3005
R11478 gnd.n491 gnd.n490 9.3005
R11479 gnd.n7479 gnd.n7478 9.3005
R11480 gnd.n7480 gnd.n489 9.3005
R11481 gnd.n7482 gnd.n7481 9.3005
R11482 gnd.n485 gnd.n484 9.3005
R11483 gnd.n7489 gnd.n7488 9.3005
R11484 gnd.n7490 gnd.n483 9.3005
R11485 gnd.n7492 gnd.n7491 9.3005
R11486 gnd.n479 gnd.n478 9.3005
R11487 gnd.n7499 gnd.n7498 9.3005
R11488 gnd.n7500 gnd.n477 9.3005
R11489 gnd.n7502 gnd.n7501 9.3005
R11490 gnd.n473 gnd.n472 9.3005
R11491 gnd.n7509 gnd.n7508 9.3005
R11492 gnd.n7510 gnd.n471 9.3005
R11493 gnd.n7512 gnd.n7511 9.3005
R11494 gnd.n467 gnd.n466 9.3005
R11495 gnd.n7519 gnd.n7518 9.3005
R11496 gnd.n7520 gnd.n465 9.3005
R11497 gnd.n7522 gnd.n7521 9.3005
R11498 gnd.n461 gnd.n460 9.3005
R11499 gnd.n7529 gnd.n7528 9.3005
R11500 gnd.n7530 gnd.n459 9.3005
R11501 gnd.n7532 gnd.n7531 9.3005
R11502 gnd.n455 gnd.n454 9.3005
R11503 gnd.n7539 gnd.n7538 9.3005
R11504 gnd.n7540 gnd.n453 9.3005
R11505 gnd.n7542 gnd.n7541 9.3005
R11506 gnd.n449 gnd.n448 9.3005
R11507 gnd.n7549 gnd.n7548 9.3005
R11508 gnd.n7550 gnd.n447 9.3005
R11509 gnd.n7552 gnd.n7551 9.3005
R11510 gnd.n443 gnd.n442 9.3005
R11511 gnd.n7559 gnd.n7558 9.3005
R11512 gnd.n7560 gnd.n441 9.3005
R11513 gnd.n7562 gnd.n7561 9.3005
R11514 gnd.n437 gnd.n436 9.3005
R11515 gnd.n7569 gnd.n7568 9.3005
R11516 gnd.n7570 gnd.n435 9.3005
R11517 gnd.n7572 gnd.n7571 9.3005
R11518 gnd.n431 gnd.n430 9.3005
R11519 gnd.n7579 gnd.n7578 9.3005
R11520 gnd.n7580 gnd.n429 9.3005
R11521 gnd.n7582 gnd.n7581 9.3005
R11522 gnd.n425 gnd.n424 9.3005
R11523 gnd.n7589 gnd.n7588 9.3005
R11524 gnd.n7590 gnd.n423 9.3005
R11525 gnd.n7592 gnd.n7591 9.3005
R11526 gnd.n419 gnd.n418 9.3005
R11527 gnd.n7599 gnd.n7598 9.3005
R11528 gnd.n7600 gnd.n417 9.3005
R11529 gnd.n7604 gnd.n7601 9.3005
R11530 gnd.n7603 gnd.n7602 9.3005
R11531 gnd.n413 gnd.n412 9.3005
R11532 gnd.n7612 gnd.n7611 9.3005
R11533 gnd.n7400 gnd.n537 9.3005
R11534 gnd.n7911 gnd.n134 9.3005
R11535 gnd.n7910 gnd.n136 9.3005
R11536 gnd.n140 gnd.n137 9.3005
R11537 gnd.n7905 gnd.n141 9.3005
R11538 gnd.n7904 gnd.n142 9.3005
R11539 gnd.n7903 gnd.n143 9.3005
R11540 gnd.n147 gnd.n144 9.3005
R11541 gnd.n7898 gnd.n148 9.3005
R11542 gnd.n7897 gnd.n149 9.3005
R11543 gnd.n7896 gnd.n150 9.3005
R11544 gnd.n154 gnd.n151 9.3005
R11545 gnd.n7891 gnd.n155 9.3005
R11546 gnd.n7890 gnd.n156 9.3005
R11547 gnd.n7889 gnd.n157 9.3005
R11548 gnd.n161 gnd.n158 9.3005
R11549 gnd.n7884 gnd.n162 9.3005
R11550 gnd.n7883 gnd.n163 9.3005
R11551 gnd.n7879 gnd.n164 9.3005
R11552 gnd.n168 gnd.n165 9.3005
R11553 gnd.n7874 gnd.n169 9.3005
R11554 gnd.n7873 gnd.n170 9.3005
R11555 gnd.n7872 gnd.n171 9.3005
R11556 gnd.n175 gnd.n172 9.3005
R11557 gnd.n7867 gnd.n176 9.3005
R11558 gnd.n7866 gnd.n177 9.3005
R11559 gnd.n7865 gnd.n178 9.3005
R11560 gnd.n182 gnd.n179 9.3005
R11561 gnd.n7860 gnd.n183 9.3005
R11562 gnd.n7859 gnd.n184 9.3005
R11563 gnd.n7858 gnd.n185 9.3005
R11564 gnd.n189 gnd.n186 9.3005
R11565 gnd.n7853 gnd.n190 9.3005
R11566 gnd.n7852 gnd.n191 9.3005
R11567 gnd.n7851 gnd.n192 9.3005
R11568 gnd.n196 gnd.n193 9.3005
R11569 gnd.n7846 gnd.n197 9.3005
R11570 gnd.n7845 gnd.n7844 9.3005
R11571 gnd.n7843 gnd.n200 9.3005
R11572 gnd.n7913 gnd.n7912 9.3005
R11573 gnd.n1939 gnd.n1902 9.3005
R11574 gnd.n1938 gnd.n1904 9.3005
R11575 gnd.n1937 gnd.n1905 9.3005
R11576 gnd.n1936 gnd.n1906 9.3005
R11577 gnd.n1934 gnd.n1907 9.3005
R11578 gnd.n1933 gnd.n1908 9.3005
R11579 gnd.n1930 gnd.n1909 9.3005
R11580 gnd.n1929 gnd.n1910 9.3005
R11581 gnd.n1928 gnd.n1911 9.3005
R11582 gnd.n1926 gnd.n1912 9.3005
R11583 gnd.n1925 gnd.n1913 9.3005
R11584 gnd.n1923 gnd.n1914 9.3005
R11585 gnd.n1922 gnd.n1915 9.3005
R11586 gnd.n1921 gnd.n1916 9.3005
R11587 gnd.n1919 gnd.n1918 9.3005
R11588 gnd.n1917 gnd.n1590 9.3005
R11589 gnd.n6165 gnd.n1591 9.3005
R11590 gnd.n6166 gnd.n1589 9.3005
R11591 gnd.n6169 gnd.n6168 9.3005
R11592 gnd.n6170 gnd.n1588 9.3005
R11593 gnd.n6202 gnd.n6171 9.3005
R11594 gnd.n6201 gnd.n6172 9.3005
R11595 gnd.n6200 gnd.n6173 9.3005
R11596 gnd.n6198 gnd.n6174 9.3005
R11597 gnd.n6197 gnd.n6175 9.3005
R11598 gnd.n6194 gnd.n6176 9.3005
R11599 gnd.n6193 gnd.n6177 9.3005
R11600 gnd.n6192 gnd.n6178 9.3005
R11601 gnd.n6189 gnd.n6179 9.3005
R11602 gnd.n6188 gnd.n6180 9.3005
R11603 gnd.n6185 gnd.n6181 9.3005
R11604 gnd.n6184 gnd.n6183 9.3005
R11605 gnd.n6182 gnd.n341 9.3005
R11606 gnd.n7642 gnd.n342 9.3005
R11607 gnd.n7641 gnd.n343 9.3005
R11608 gnd.n7640 gnd.n344 9.3005
R11609 gnd.n7636 gnd.n345 9.3005
R11610 gnd.n7635 gnd.n346 9.3005
R11611 gnd.n7632 gnd.n347 9.3005
R11612 gnd.n7631 gnd.n348 9.3005
R11613 gnd.n7627 gnd.n349 9.3005
R11614 gnd.n7626 gnd.n350 9.3005
R11615 gnd.n401 gnd.n351 9.3005
R11616 gnd.n400 gnd.n352 9.3005
R11617 gnd.n396 gnd.n353 9.3005
R11618 gnd.n395 gnd.n354 9.3005
R11619 gnd.n392 gnd.n355 9.3005
R11620 gnd.n391 gnd.n356 9.3005
R11621 gnd.n389 gnd.n357 9.3005
R11622 gnd.n388 gnd.n358 9.3005
R11623 gnd.n386 gnd.n359 9.3005
R11624 gnd.n385 gnd.n360 9.3005
R11625 gnd.n383 gnd.n361 9.3005
R11626 gnd.n382 gnd.n362 9.3005
R11627 gnd.n380 gnd.n363 9.3005
R11628 gnd.n379 gnd.n364 9.3005
R11629 gnd.n377 gnd.n365 9.3005
R11630 gnd.n376 gnd.n366 9.3005
R11631 gnd.n374 gnd.n367 9.3005
R11632 gnd.n373 gnd.n368 9.3005
R11633 gnd.n371 gnd.n370 9.3005
R11634 gnd.n369 gnd.n204 9.3005
R11635 gnd.n7840 gnd.n203 9.3005
R11636 gnd.n7842 gnd.n7841 9.3005
R11637 gnd.n1941 gnd.n1940 9.3005
R11638 gnd.n1947 gnd.n1946 9.3005
R11639 gnd.n1948 gnd.n1896 9.3005
R11640 gnd.n1951 gnd.n1895 9.3005
R11641 gnd.n1952 gnd.n1894 9.3005
R11642 gnd.n1955 gnd.n1893 9.3005
R11643 gnd.n1956 gnd.n1892 9.3005
R11644 gnd.n1959 gnd.n1891 9.3005
R11645 gnd.n1960 gnd.n1890 9.3005
R11646 gnd.n1963 gnd.n1889 9.3005
R11647 gnd.n1964 gnd.n1888 9.3005
R11648 gnd.n1967 gnd.n1887 9.3005
R11649 gnd.n1968 gnd.n1886 9.3005
R11650 gnd.n1971 gnd.n1885 9.3005
R11651 gnd.n1972 gnd.n1884 9.3005
R11652 gnd.n1975 gnd.n1883 9.3005
R11653 gnd.n1976 gnd.n1882 9.3005
R11654 gnd.n1979 gnd.n1881 9.3005
R11655 gnd.n1980 gnd.n1880 9.3005
R11656 gnd.n1983 gnd.n1879 9.3005
R11657 gnd.n1875 gnd.n1835 9.3005
R11658 gnd.n1874 gnd.n1873 9.3005
R11659 gnd.n1870 gnd.n1837 9.3005
R11660 gnd.n1867 gnd.n1866 9.3005
R11661 gnd.n1865 gnd.n1838 9.3005
R11662 gnd.n1864 gnd.n1863 9.3005
R11663 gnd.n1860 gnd.n1839 9.3005
R11664 gnd.n1857 gnd.n1856 9.3005
R11665 gnd.n1855 gnd.n1840 9.3005
R11666 gnd.n1854 gnd.n1853 9.3005
R11667 gnd.n1850 gnd.n1841 9.3005
R11668 gnd.n1847 gnd.n1846 9.3005
R11669 gnd.n1845 gnd.n1843 9.3005
R11670 gnd.n1844 gnd.n1688 9.3005
R11671 gnd.n6044 gnd.n1687 9.3005
R11672 gnd.n6046 gnd.n6045 9.3005
R11673 gnd.n1945 gnd.n1901 9.3005
R11674 gnd.n1944 gnd.n1943 9.3005
R11675 gnd.n6049 gnd.n6048 9.3005
R11676 gnd.n1663 gnd.n1662 9.3005
R11677 gnd.n6077 gnd.n6076 9.3005
R11678 gnd.n6078 gnd.n1661 9.3005
R11679 gnd.n6082 gnd.n6079 9.3005
R11680 gnd.n6081 gnd.n6080 9.3005
R11681 gnd.n1637 gnd.n1636 9.3005
R11682 gnd.n6109 gnd.n6108 9.3005
R11683 gnd.n6110 gnd.n1635 9.3005
R11684 gnd.n6114 gnd.n6111 9.3005
R11685 gnd.n6113 gnd.n6112 9.3005
R11686 gnd.n1609 gnd.n1608 9.3005
R11687 gnd.n6147 gnd.n6146 9.3005
R11688 gnd.n6148 gnd.n1607 9.3005
R11689 gnd.n6152 gnd.n6149 9.3005
R11690 gnd.n6151 gnd.n6150 9.3005
R11691 gnd.n1572 gnd.n1571 9.3005
R11692 gnd.n6215 gnd.n6214 9.3005
R11693 gnd.n6216 gnd.n1570 9.3005
R11694 gnd.n6218 gnd.n6217 9.3005
R11695 gnd.n1556 gnd.n1555 9.3005
R11696 gnd.n6235 gnd.n6234 9.3005
R11697 gnd.n6236 gnd.n1554 9.3005
R11698 gnd.n6240 gnd.n6237 9.3005
R11699 gnd.n6239 gnd.n6238 9.3005
R11700 gnd.n1520 gnd.n311 9.3005
R11701 gnd.n296 gnd.n295 9.3005
R11702 gnd.n7682 gnd.n7681 9.3005
R11703 gnd.n7683 gnd.n294 9.3005
R11704 gnd.n7685 gnd.n7684 9.3005
R11705 gnd.n281 gnd.n280 9.3005
R11706 gnd.n7698 gnd.n7697 9.3005
R11707 gnd.n7699 gnd.n279 9.3005
R11708 gnd.n7701 gnd.n7700 9.3005
R11709 gnd.n264 gnd.n263 9.3005
R11710 gnd.n7714 gnd.n7713 9.3005
R11711 gnd.n7715 gnd.n262 9.3005
R11712 gnd.n7717 gnd.n7716 9.3005
R11713 gnd.n250 gnd.n249 9.3005
R11714 gnd.n7730 gnd.n7729 9.3005
R11715 gnd.n7731 gnd.n248 9.3005
R11716 gnd.n7733 gnd.n7732 9.3005
R11717 gnd.n235 gnd.n234 9.3005
R11718 gnd.n7746 gnd.n7745 9.3005
R11719 gnd.n7747 gnd.n233 9.3005
R11720 gnd.n7749 gnd.n7748 9.3005
R11721 gnd.n220 gnd.n219 9.3005
R11722 gnd.n7762 gnd.n7761 9.3005
R11723 gnd.n7763 gnd.n218 9.3005
R11724 gnd.n7767 gnd.n7764 9.3005
R11725 gnd.n7766 gnd.n7765 9.3005
R11726 gnd.n133 gnd.n132 9.3005
R11727 gnd.n7915 gnd.n7914 9.3005
R11728 gnd.n6050 gnd.n6047 9.3005
R11729 gnd.n7669 gnd.n7668 9.3005
R11730 gnd.n4606 gnd.n4605 9.3005
R11731 gnd.n4604 gnd.n2512 9.3005
R11732 gnd.n2510 gnd.n2509 9.3005
R11733 gnd.n4682 gnd.n4681 9.3005
R11734 gnd.n4683 gnd.n2508 9.3005
R11735 gnd.n4685 gnd.n4684 9.3005
R11736 gnd.n2506 gnd.n2505 9.3005
R11737 gnd.n4690 gnd.n4689 9.3005
R11738 gnd.n4691 gnd.n2504 9.3005
R11739 gnd.n4710 gnd.n4692 9.3005
R11740 gnd.n4709 gnd.n4693 9.3005
R11741 gnd.n4708 gnd.n4694 9.3005
R11742 gnd.n4697 gnd.n4695 9.3005
R11743 gnd.n4704 gnd.n4698 9.3005
R11744 gnd.n4703 gnd.n4699 9.3005
R11745 gnd.n4702 gnd.n4700 9.3005
R11746 gnd.n2473 gnd.n2472 9.3005
R11747 gnd.n4892 gnd.n4891 9.3005
R11748 gnd.n4893 gnd.n2471 9.3005
R11749 gnd.n4895 gnd.n4894 9.3005
R11750 gnd.n2469 gnd.n2468 9.3005
R11751 gnd.n4900 gnd.n4899 9.3005
R11752 gnd.n4901 gnd.n2467 9.3005
R11753 gnd.n4903 gnd.n4902 9.3005
R11754 gnd.n2465 gnd.n2464 9.3005
R11755 gnd.n4908 gnd.n4907 9.3005
R11756 gnd.n4909 gnd.n2463 9.3005
R11757 gnd.n4920 gnd.n4910 9.3005
R11758 gnd.n4919 gnd.n4911 9.3005
R11759 gnd.n4918 gnd.n4912 9.3005
R11760 gnd.n4914 gnd.n4913 9.3005
R11761 gnd.n2314 gnd.n2313 9.3005
R11762 gnd.n4977 gnd.n4976 9.3005
R11763 gnd.n4978 gnd.n2312 9.3005
R11764 gnd.n4980 gnd.n4979 9.3005
R11765 gnd.n2300 gnd.n2299 9.3005
R11766 gnd.n4993 gnd.n4992 9.3005
R11767 gnd.n4994 gnd.n2298 9.3005
R11768 gnd.n4996 gnd.n4995 9.3005
R11769 gnd.n2286 gnd.n2285 9.3005
R11770 gnd.n5009 gnd.n5008 9.3005
R11771 gnd.n5010 gnd.n2284 9.3005
R11772 gnd.n5012 gnd.n5011 9.3005
R11773 gnd.n2272 gnd.n2271 9.3005
R11774 gnd.n5025 gnd.n5024 9.3005
R11775 gnd.n5026 gnd.n2270 9.3005
R11776 gnd.n5028 gnd.n5027 9.3005
R11777 gnd.n2258 gnd.n2257 9.3005
R11778 gnd.n5041 gnd.n5040 9.3005
R11779 gnd.n5042 gnd.n2256 9.3005
R11780 gnd.n5044 gnd.n5043 9.3005
R11781 gnd.n2243 gnd.n2242 9.3005
R11782 gnd.n5057 gnd.n5056 9.3005
R11783 gnd.n5058 gnd.n2241 9.3005
R11784 gnd.n5060 gnd.n5059 9.3005
R11785 gnd.n2228 gnd.n2227 9.3005
R11786 gnd.n5084 gnd.n5083 9.3005
R11787 gnd.n5085 gnd.n2226 9.3005
R11788 gnd.n5090 gnd.n5086 9.3005
R11789 gnd.n5089 gnd.n5088 9.3005
R11790 gnd.n5087 gnd.n1370 9.3005
R11791 gnd.n6470 gnd.n1371 9.3005
R11792 gnd.n6469 gnd.n1372 9.3005
R11793 gnd.n6468 gnd.n1373 9.3005
R11794 gnd.n5241 gnd.n1374 9.3005
R11795 gnd.n5243 gnd.n5242 9.3005
R11796 gnd.n2199 gnd.n2198 9.3005
R11797 gnd.n5267 gnd.n5266 9.3005
R11798 gnd.n5268 gnd.n2197 9.3005
R11799 gnd.n5270 gnd.n5269 9.3005
R11800 gnd.n2180 gnd.n2179 9.3005
R11801 gnd.n5291 gnd.n5290 9.3005
R11802 gnd.n5292 gnd.n2178 9.3005
R11803 gnd.n5294 gnd.n5293 9.3005
R11804 gnd.n2158 gnd.n2157 9.3005
R11805 gnd.n5317 gnd.n5316 9.3005
R11806 gnd.n5318 gnd.n2156 9.3005
R11807 gnd.n5322 gnd.n5319 9.3005
R11808 gnd.n5321 gnd.n5320 9.3005
R11809 gnd.n2129 gnd.n2128 9.3005
R11810 gnd.n5372 gnd.n5371 9.3005
R11811 gnd.n5373 gnd.n2127 9.3005
R11812 gnd.n5377 gnd.n5374 9.3005
R11813 gnd.n5376 gnd.n5375 9.3005
R11814 gnd.n2106 gnd.n2105 9.3005
R11815 gnd.n5413 gnd.n5412 9.3005
R11816 gnd.n5414 gnd.n2104 9.3005
R11817 gnd.n5418 gnd.n5415 9.3005
R11818 gnd.n5417 gnd.n5416 9.3005
R11819 gnd.n2077 gnd.n2076 9.3005
R11820 gnd.n5454 gnd.n5453 9.3005
R11821 gnd.n5455 gnd.n2075 9.3005
R11822 gnd.n5458 gnd.n5457 9.3005
R11823 gnd.n5456 gnd.n2053 9.3005
R11824 gnd.n5505 gnd.n2054 9.3005
R11825 gnd.n5504 gnd.n2055 9.3005
R11826 gnd.n5503 gnd.n2056 9.3005
R11827 gnd.n2058 gnd.n2057 9.3005
R11828 gnd.n2060 gnd.n2059 9.3005
R11829 gnd.n2019 gnd.n2018 9.3005
R11830 gnd.n5554 gnd.n5553 9.3005
R11831 gnd.n5555 gnd.n2017 9.3005
R11832 gnd.n5557 gnd.n5556 9.3005
R11833 gnd.n2003 gnd.n2002 9.3005
R11834 gnd.n5585 gnd.n5584 9.3005
R11835 gnd.n5586 gnd.n2001 9.3005
R11836 gnd.n5588 gnd.n5587 9.3005
R11837 gnd.n1797 gnd.n1796 9.3005
R11838 gnd.n5760 gnd.n5759 9.3005
R11839 gnd.n5761 gnd.n1795 9.3005
R11840 gnd.n5763 gnd.n5762 9.3005
R11841 gnd.n1785 gnd.n1784 9.3005
R11842 gnd.n5778 gnd.n5777 9.3005
R11843 gnd.n5779 gnd.n1783 9.3005
R11844 gnd.n5781 gnd.n5780 9.3005
R11845 gnd.n1774 gnd.n1773 9.3005
R11846 gnd.n5795 gnd.n5794 9.3005
R11847 gnd.n5796 gnd.n1772 9.3005
R11848 gnd.n5798 gnd.n5797 9.3005
R11849 gnd.n1762 gnd.n1761 9.3005
R11850 gnd.n5812 gnd.n5811 9.3005
R11851 gnd.n5813 gnd.n1760 9.3005
R11852 gnd.n5815 gnd.n5814 9.3005
R11853 gnd.n1750 gnd.n1749 9.3005
R11854 gnd.n5829 gnd.n5828 9.3005
R11855 gnd.n5830 gnd.n1748 9.3005
R11856 gnd.n5832 gnd.n5831 9.3005
R11857 gnd.n1738 gnd.n1737 9.3005
R11858 gnd.n5846 gnd.n5845 9.3005
R11859 gnd.n5847 gnd.n1736 9.3005
R11860 gnd.n5851 gnd.n5848 9.3005
R11861 gnd.n5850 gnd.n5849 9.3005
R11862 gnd.n1726 gnd.n1725 9.3005
R11863 gnd.n5866 gnd.n5865 9.3005
R11864 gnd.n5867 gnd.n1724 9.3005
R11865 gnd.n5869 gnd.n5868 9.3005
R11866 gnd.n1723 gnd.n1722 9.3005
R11867 gnd.n6033 gnd.n6032 9.3005
R11868 gnd.n6034 gnd.n1721 9.3005
R11869 gnd.n6038 gnd.n6035 9.3005
R11870 gnd.n6037 gnd.n6036 9.3005
R11871 gnd.n1673 gnd.n1672 9.3005
R11872 gnd.n6065 gnd.n6064 9.3005
R11873 gnd.n6066 gnd.n1671 9.3005
R11874 gnd.n6070 gnd.n6067 9.3005
R11875 gnd.n6069 gnd.n6068 9.3005
R11876 gnd.n1647 gnd.n1646 9.3005
R11877 gnd.n6098 gnd.n6097 9.3005
R11878 gnd.n6099 gnd.n1645 9.3005
R11879 gnd.n6103 gnd.n6100 9.3005
R11880 gnd.n6102 gnd.n6101 9.3005
R11881 gnd.n1619 gnd.n1618 9.3005
R11882 gnd.n6129 gnd.n6128 9.3005
R11883 gnd.n6130 gnd.n1617 9.3005
R11884 gnd.n6141 gnd.n6131 9.3005
R11885 gnd.n6140 gnd.n6132 9.3005
R11886 gnd.n6139 gnd.n6133 9.3005
R11887 gnd.n6136 gnd.n6135 9.3005
R11888 gnd.n6134 gnd.n1581 9.3005
R11889 gnd.n6209 gnd.n1582 9.3005
R11890 gnd.n6208 gnd.n1583 9.3005
R11891 gnd.n6207 gnd.n1584 9.3005
R11892 gnd.n1586 gnd.n1585 9.3005
R11893 gnd.n1546 gnd.n1545 9.3005
R11894 gnd.n6246 gnd.n6245 9.3005
R11895 gnd.n6247 gnd.n1544 9.3005
R11896 gnd.n6250 gnd.n6249 9.3005
R11897 gnd.n6248 gnd.n1542 9.3005
R11898 gnd.n6274 gnd.n6266 9.3005
R11899 gnd.n6273 gnd.n6267 9.3005
R11900 gnd.n6270 gnd.n6269 9.3005
R11901 gnd.n6268 gnd.n404 9.3005
R11902 gnd.n7621 gnd.n405 9.3005
R11903 gnd.n7620 gnd.n406 9.3005
R11904 gnd.n7619 gnd.n407 9.3005
R11905 gnd.n410 gnd.n408 9.3005
R11906 gnd.n7615 gnd.n411 9.3005
R11907 gnd.n7614 gnd.n7613 9.3005
R11908 gnd.n4578 gnd.n4577 9.3005
R11909 gnd.n4395 gnd.n4353 9.3005
R11910 gnd.n4393 gnd.n4354 9.3005
R11911 gnd.n4392 gnd.n4355 9.3005
R11912 gnd.n4390 gnd.n4356 9.3005
R11913 gnd.n4389 gnd.n4357 9.3005
R11914 gnd.n4387 gnd.n4358 9.3005
R11915 gnd.n4386 gnd.n4359 9.3005
R11916 gnd.n4384 gnd.n4360 9.3005
R11917 gnd.n4383 gnd.n4361 9.3005
R11918 gnd.n4381 gnd.n4362 9.3005
R11919 gnd.n4380 gnd.n4363 9.3005
R11920 gnd.n4378 gnd.n4364 9.3005
R11921 gnd.n4377 gnd.n4365 9.3005
R11922 gnd.n4375 gnd.n4366 9.3005
R11923 gnd.n4374 gnd.n4367 9.3005
R11924 gnd.n4372 gnd.n4368 9.3005
R11925 gnd.n4371 gnd.n4369 9.3005
R11926 gnd.n2612 gnd.n2611 9.3005
R11927 gnd.n4524 gnd.n4523 9.3005
R11928 gnd.n4525 gnd.n2610 9.3005
R11929 gnd.n4527 gnd.n4526 9.3005
R11930 gnd.n2582 gnd.n2581 9.3005
R11931 gnd.n4545 gnd.n4544 9.3005
R11932 gnd.n4546 gnd.n2580 9.3005
R11933 gnd.n4549 gnd.n4548 9.3005
R11934 gnd.n4547 gnd.n2557 9.3005
R11935 gnd.n4571 gnd.n2556 9.3005
R11936 gnd.n4573 gnd.n4572 9.3005
R11937 gnd.n4574 gnd.n2555 9.3005
R11938 gnd.n4580 gnd.n4575 9.3005
R11939 gnd.n4579 gnd.n4576 9.3005
R11940 gnd.n4397 gnd.n4396 9.3005
R11941 gnd.n4405 gnd.n4404 9.3005
R11942 gnd.n4406 gnd.n4349 9.3005
R11943 gnd.n4348 gnd.n4346 9.3005
R11944 gnd.n4412 gnd.n4345 9.3005
R11945 gnd.n4413 gnd.n4344 9.3005
R11946 gnd.n4414 gnd.n4343 9.3005
R11947 gnd.n4342 gnd.n4340 9.3005
R11948 gnd.n4420 gnd.n4339 9.3005
R11949 gnd.n4421 gnd.n4338 9.3005
R11950 gnd.n4422 gnd.n4337 9.3005
R11951 gnd.n4336 gnd.n4334 9.3005
R11952 gnd.n4428 gnd.n4333 9.3005
R11953 gnd.n4429 gnd.n4332 9.3005
R11954 gnd.n4430 gnd.n4331 9.3005
R11955 gnd.n4330 gnd.n4328 9.3005
R11956 gnd.n4436 gnd.n4327 9.3005
R11957 gnd.n4438 gnd.n4437 9.3005
R11958 gnd.n4403 gnd.n4352 9.3005
R11959 gnd.n4402 gnd.n4401 9.3005
R11960 gnd.n2665 gnd.n2664 9.3005
R11961 gnd.n4453 gnd.n4452 9.3005
R11962 gnd.n4454 gnd.n2663 9.3005
R11963 gnd.n4456 gnd.n4455 9.3005
R11964 gnd.n2649 gnd.n2648 9.3005
R11965 gnd.n4469 gnd.n4468 9.3005
R11966 gnd.n4470 gnd.n2647 9.3005
R11967 gnd.n4472 gnd.n4471 9.3005
R11968 gnd.n2633 gnd.n2632 9.3005
R11969 gnd.n4485 gnd.n4484 9.3005
R11970 gnd.n4486 gnd.n2631 9.3005
R11971 gnd.n4498 gnd.n4487 9.3005
R11972 gnd.n4497 gnd.n4488 9.3005
R11973 gnd.n4496 gnd.n4489 9.3005
R11974 gnd.n4495 gnd.n4490 9.3005
R11975 gnd.n4493 gnd.n4492 9.3005
R11976 gnd.n4491 gnd.n1038 9.3005
R11977 gnd.n6699 gnd.n1039 9.3005
R11978 gnd.n6698 gnd.n1040 9.3005
R11979 gnd.n6697 gnd.n1041 9.3005
R11980 gnd.n1059 gnd.n1042 9.3005
R11981 gnd.n6687 gnd.n1060 9.3005
R11982 gnd.n6686 gnd.n1061 9.3005
R11983 gnd.n6685 gnd.n1062 9.3005
R11984 gnd.n1080 gnd.n1063 9.3005
R11985 gnd.n6675 gnd.n1081 9.3005
R11986 gnd.n6674 gnd.n1082 9.3005
R11987 gnd.n6673 gnd.n1083 9.3005
R11988 gnd.n4584 gnd.n1084 9.3005
R11989 gnd.n4588 gnd.n4585 9.3005
R11990 gnd.n4587 gnd.n4586 9.3005
R11991 gnd.n2540 gnd.n2539 9.3005
R11992 gnd.n4619 gnd.n4618 9.3005
R11993 gnd.n4620 gnd.n2538 9.3005
R11994 gnd.n4623 gnd.n4622 9.3005
R11995 gnd.n4621 gnd.n1107 9.3005
R11996 gnd.n6661 gnd.n1108 9.3005
R11997 gnd.n6660 gnd.n1109 9.3005
R11998 gnd.n6659 gnd.n1110 9.3005
R11999 gnd.n1127 gnd.n1111 9.3005
R12000 gnd.n6649 gnd.n1128 9.3005
R12001 gnd.n6648 gnd.n1129 9.3005
R12002 gnd.n6647 gnd.n1130 9.3005
R12003 gnd.n1149 gnd.n1131 9.3005
R12004 gnd.n6637 gnd.n1150 9.3005
R12005 gnd.n6636 gnd.n1151 9.3005
R12006 gnd.n6635 gnd.n1152 9.3005
R12007 gnd.n1170 gnd.n1153 9.3005
R12008 gnd.n6625 gnd.n1171 9.3005
R12009 gnd.n6624 gnd.n1172 9.3005
R12010 gnd.n6623 gnd.n1173 9.3005
R12011 gnd.n1192 gnd.n1174 9.3005
R12012 gnd.n6613 gnd.n1193 9.3005
R12013 gnd.n6612 gnd.n1194 9.3005
R12014 gnd.n6611 gnd.n1195 9.3005
R12015 gnd.n1213 gnd.n1196 9.3005
R12016 gnd.n6601 gnd.n1214 9.3005
R12017 gnd.n6600 gnd.n1215 9.3005
R12018 gnd.n6599 gnd.n1216 9.3005
R12019 gnd.n1235 gnd.n1217 9.3005
R12020 gnd.n6589 gnd.n1236 9.3005
R12021 gnd.n6588 gnd.n1237 9.3005
R12022 gnd.n6587 gnd.n1238 9.3005
R12023 gnd.n2339 gnd.n1239 9.3005
R12024 gnd.n4440 gnd.n4439 9.3005
R12025 gnd.n6549 gnd.n1295 9.3005
R12026 gnd.n6552 gnd.n1294 9.3005
R12027 gnd.n6553 gnd.n1293 9.3005
R12028 gnd.n6556 gnd.n1292 9.3005
R12029 gnd.n6557 gnd.n1291 9.3005
R12030 gnd.n6560 gnd.n1290 9.3005
R12031 gnd.n6561 gnd.n1289 9.3005
R12032 gnd.n6564 gnd.n1288 9.3005
R12033 gnd.n6565 gnd.n1287 9.3005
R12034 gnd.n6568 gnd.n1286 9.3005
R12035 gnd.n6569 gnd.n1285 9.3005
R12036 gnd.n6572 gnd.n1284 9.3005
R12037 gnd.n6573 gnd.n1283 9.3005
R12038 gnd.n6574 gnd.n1282 9.3005
R12039 gnd.n1249 gnd.n1248 9.3005
R12040 gnd.n6580 gnd.n6579 9.3005
R12041 gnd.n4778 gnd.n4776 9.3005
R12042 gnd.n4780 gnd.n4779 9.3005
R12043 gnd.n4783 gnd.n4773 9.3005
R12044 gnd.n4787 gnd.n4786 9.3005
R12045 gnd.n4788 gnd.n4772 9.3005
R12046 gnd.n4790 gnd.n4789 9.3005
R12047 gnd.n4793 gnd.n4771 9.3005
R12048 gnd.n4797 gnd.n4796 9.3005
R12049 gnd.n4798 gnd.n4770 9.3005
R12050 gnd.n4800 gnd.n4799 9.3005
R12051 gnd.n4803 gnd.n4769 9.3005
R12052 gnd.n4807 gnd.n4806 9.3005
R12053 gnd.n4808 gnd.n4768 9.3005
R12054 gnd.n4810 gnd.n4809 9.3005
R12055 gnd.n4813 gnd.n4767 9.3005
R12056 gnd.n4817 gnd.n4816 9.3005
R12057 gnd.n4818 gnd.n4766 9.3005
R12058 gnd.n4821 gnd.n4819 9.3005
R12059 gnd.n4822 gnd.n4762 9.3005
R12060 gnd.n4825 gnd.n4824 9.3005
R12061 gnd.n4777 gnd.n1296 9.3005
R12062 gnd.n4323 gnd.n4322 9.3005
R12063 gnd.n4321 gnd.n4152 9.3005
R12064 gnd.n4320 gnd.n4319 9.3005
R12065 gnd.n4317 gnd.n4293 9.3005
R12066 gnd.n4316 gnd.n4294 9.3005
R12067 gnd.n4314 gnd.n4295 9.3005
R12068 gnd.n4313 gnd.n4296 9.3005
R12069 gnd.n4311 gnd.n4297 9.3005
R12070 gnd.n4310 gnd.n4298 9.3005
R12071 gnd.n4308 gnd.n4299 9.3005
R12072 gnd.n4307 gnd.n4300 9.3005
R12073 gnd.n4305 gnd.n4301 9.3005
R12074 gnd.n4304 gnd.n4303 9.3005
R12075 gnd.n4302 gnd.n2615 9.3005
R12076 gnd.n4512 gnd.n2616 9.3005
R12077 gnd.n4513 gnd.n2614 9.3005
R12078 gnd.n4516 gnd.n4515 9.3005
R12079 gnd.n4517 gnd.n2613 9.3005
R12080 gnd.n4519 gnd.n4518 9.3005
R12081 gnd.n2585 gnd.n2584 9.3005
R12082 gnd.n4532 gnd.n4531 9.3005
R12083 gnd.n4533 gnd.n2583 9.3005
R12084 gnd.n4540 gnd.n4534 9.3005
R12085 gnd.n4539 gnd.n4535 9.3005
R12086 gnd.n4538 gnd.n4537 9.3005
R12087 gnd.n4536 gnd.n2558 9.3005
R12088 gnd.n4567 gnd.n2559 9.3005
R12089 gnd.n4566 gnd.n2560 9.3005
R12090 gnd.n4565 gnd.n2561 9.3005
R12091 gnd.n2573 gnd.n2562 9.3005
R12092 gnd.n2572 gnd.n2563 9.3005
R12093 gnd.n2570 gnd.n2564 9.3005
R12094 gnd.n2569 gnd.n2565 9.3005
R12095 gnd.n2568 gnd.n2567 9.3005
R12096 gnd.n2566 gnd.n2525 9.3005
R12097 gnd.n4640 gnd.n2526 9.3005
R12098 gnd.n4641 gnd.n2524 9.3005
R12099 gnd.n4643 gnd.n4642 9.3005
R12100 gnd.n4644 gnd.n2523 9.3005
R12101 gnd.n4648 gnd.n4645 9.3005
R12102 gnd.n4649 gnd.n2522 9.3005
R12103 gnd.n4653 gnd.n4652 9.3005
R12104 gnd.n4654 gnd.n2521 9.3005
R12105 gnd.n4660 gnd.n4655 9.3005
R12106 gnd.n4659 gnd.n4656 9.3005
R12107 gnd.n4658 gnd.n4657 9.3005
R12108 gnd.n2497 gnd.n2496 9.3005
R12109 gnd.n4724 gnd.n4723 9.3005
R12110 gnd.n4725 gnd.n2495 9.3005
R12111 gnd.n4727 gnd.n4726 9.3005
R12112 gnd.n2491 gnd.n2490 9.3005
R12113 gnd.n4740 gnd.n4739 9.3005
R12114 gnd.n4741 gnd.n2489 9.3005
R12115 gnd.n4743 gnd.n4742 9.3005
R12116 gnd.n4744 gnd.n2488 9.3005
R12117 gnd.n4748 gnd.n4747 9.3005
R12118 gnd.n4749 gnd.n2487 9.3005
R12119 gnd.n4753 gnd.n4750 9.3005
R12120 gnd.n4754 gnd.n2486 9.3005
R12121 gnd.n4758 gnd.n4757 9.3005
R12122 gnd.n4759 gnd.n2485 9.3005
R12123 gnd.n4829 gnd.n4760 9.3005
R12124 gnd.n4828 gnd.n4761 9.3005
R12125 gnd.n4827 gnd.n4826 9.3005
R12126 gnd.n4292 gnd.n4151 9.3005
R12127 gnd.n4281 gnd.n4157 9.3005
R12128 gnd.n4283 gnd.n4282 9.3005
R12129 gnd.n4280 gnd.n4159 9.3005
R12130 gnd.n4279 gnd.n4278 9.3005
R12131 gnd.n4161 gnd.n4160 9.3005
R12132 gnd.n4272 gnd.n4271 9.3005
R12133 gnd.n4270 gnd.n4163 9.3005
R12134 gnd.n4269 gnd.n4268 9.3005
R12135 gnd.n4165 gnd.n4164 9.3005
R12136 gnd.n4262 gnd.n4261 9.3005
R12137 gnd.n4260 gnd.n4167 9.3005
R12138 gnd.n4259 gnd.n4258 9.3005
R12139 gnd.n4169 gnd.n4168 9.3005
R12140 gnd.n4252 gnd.n4251 9.3005
R12141 gnd.n4250 gnd.n4171 9.3005
R12142 gnd.n4249 gnd.n4248 9.3005
R12143 gnd.n4173 gnd.n4172 9.3005
R12144 gnd.n4242 gnd.n4241 9.3005
R12145 gnd.n4240 gnd.n4175 9.3005
R12146 gnd.n4239 gnd.n4238 9.3005
R12147 gnd.n4177 gnd.n4176 9.3005
R12148 gnd.n4232 gnd.n4231 9.3005
R12149 gnd.n4230 gnd.n4182 9.3005
R12150 gnd.n4229 gnd.n4228 9.3005
R12151 gnd.n4184 gnd.n4183 9.3005
R12152 gnd.n4222 gnd.n4221 9.3005
R12153 gnd.n4220 gnd.n4186 9.3005
R12154 gnd.n4219 gnd.n4218 9.3005
R12155 gnd.n4188 gnd.n4187 9.3005
R12156 gnd.n4212 gnd.n4211 9.3005
R12157 gnd.n4210 gnd.n4190 9.3005
R12158 gnd.n4209 gnd.n4208 9.3005
R12159 gnd.n4192 gnd.n4191 9.3005
R12160 gnd.n4202 gnd.n4201 9.3005
R12161 gnd.n4200 gnd.n4194 9.3005
R12162 gnd.n4199 gnd.n4198 9.3005
R12163 gnd.n4195 gnd.n2671 9.3005
R12164 gnd.n4156 gnd.n4153 9.3005
R12165 gnd.n4291 gnd.n4290 9.3005
R12166 gnd.n4446 gnd.n2670 9.3005
R12167 gnd.n4448 gnd.n4447 9.3005
R12168 gnd.n2657 gnd.n2656 9.3005
R12169 gnd.n4461 gnd.n4460 9.3005
R12170 gnd.n4462 gnd.n2655 9.3005
R12171 gnd.n4464 gnd.n4463 9.3005
R12172 gnd.n2640 gnd.n2639 9.3005
R12173 gnd.n4477 gnd.n4476 9.3005
R12174 gnd.n4478 gnd.n2638 9.3005
R12175 gnd.n4480 gnd.n4479 9.3005
R12176 gnd.n2624 gnd.n2623 9.3005
R12177 gnd.n4503 gnd.n4502 9.3005
R12178 gnd.n4504 gnd.n2622 9.3005
R12179 gnd.n4507 gnd.n4506 9.3005
R12180 gnd.n4505 gnd.n1026 9.3005
R12181 gnd.n6705 gnd.n1027 9.3005
R12182 gnd.n6704 gnd.n1028 9.3005
R12183 gnd.n6703 gnd.n1029 9.3005
R12184 gnd.n1048 gnd.n1030 9.3005
R12185 gnd.n6693 gnd.n1049 9.3005
R12186 gnd.n6692 gnd.n1050 9.3005
R12187 gnd.n6691 gnd.n1051 9.3005
R12188 gnd.n1070 gnd.n1052 9.3005
R12189 gnd.n6681 gnd.n1071 9.3005
R12190 gnd.n6680 gnd.n1072 9.3005
R12191 gnd.n6679 gnd.n1073 9.3005
R12192 gnd.n1098 gnd.n1092 9.3005
R12193 gnd.n6655 gnd.n1117 9.3005
R12194 gnd.n6654 gnd.n1118 9.3005
R12195 gnd.n6653 gnd.n1119 9.3005
R12196 gnd.n1138 gnd.n1120 9.3005
R12197 gnd.n6643 gnd.n1139 9.3005
R12198 gnd.n6642 gnd.n1140 9.3005
R12199 gnd.n6641 gnd.n1141 9.3005
R12200 gnd.n1159 gnd.n1142 9.3005
R12201 gnd.n6631 gnd.n1160 9.3005
R12202 gnd.n6630 gnd.n1161 9.3005
R12203 gnd.n6629 gnd.n1162 9.3005
R12204 gnd.n1181 gnd.n1163 9.3005
R12205 gnd.n6619 gnd.n1182 9.3005
R12206 gnd.n6618 gnd.n1183 9.3005
R12207 gnd.n6617 gnd.n1184 9.3005
R12208 gnd.n1202 gnd.n1185 9.3005
R12209 gnd.n6607 gnd.n1203 9.3005
R12210 gnd.n6606 gnd.n1204 9.3005
R12211 gnd.n6605 gnd.n1205 9.3005
R12212 gnd.n1224 gnd.n1206 9.3005
R12213 gnd.n6595 gnd.n1225 9.3005
R12214 gnd.n6594 gnd.n1226 9.3005
R12215 gnd.n6593 gnd.n1227 9.3005
R12216 gnd.n1246 gnd.n1228 9.3005
R12217 gnd.n6583 gnd.n1247 9.3005
R12218 gnd.n6582 gnd.n6581 9.3005
R12219 gnd.n4445 gnd.n4444 9.3005
R12220 gnd.n6666 gnd.n6665 9.3005
R12221 gnd.n2593 gnd.n2592 9.3005
R12222 gnd.n2594 gnd.n2588 9.3005
R12223 gnd.n2607 gnd.n2595 9.3005
R12224 gnd.n2606 gnd.n2596 9.3005
R12225 gnd.n2605 gnd.n2597 9.3005
R12226 gnd.n2602 gnd.n2598 9.3005
R12227 gnd.n2601 gnd.n2600 9.3005
R12228 gnd.n2599 gnd.n2576 9.3005
R12229 gnd.n4555 gnd.n2577 9.3005
R12230 gnd.n2590 gnd.n2589 9.3005
R12231 gnd.n6711 gnd.n1016 9.3005
R12232 gnd.n6712 gnd.n1015 9.3005
R12233 gnd.n1014 gnd.n1010 9.3005
R12234 gnd.n6718 gnd.n1009 9.3005
R12235 gnd.n6719 gnd.n1008 9.3005
R12236 gnd.n6720 gnd.n1007 9.3005
R12237 gnd.n1006 gnd.n1002 9.3005
R12238 gnd.n6726 gnd.n1001 9.3005
R12239 gnd.n6727 gnd.n1000 9.3005
R12240 gnd.n6728 gnd.n999 9.3005
R12241 gnd.n998 gnd.n994 9.3005
R12242 gnd.n6734 gnd.n993 9.3005
R12243 gnd.n6735 gnd.n992 9.3005
R12244 gnd.n6736 gnd.n991 9.3005
R12245 gnd.n990 gnd.n986 9.3005
R12246 gnd.n6742 gnd.n985 9.3005
R12247 gnd.n6743 gnd.n984 9.3005
R12248 gnd.n6744 gnd.n983 9.3005
R12249 gnd.n982 gnd.n978 9.3005
R12250 gnd.n6750 gnd.n977 9.3005
R12251 gnd.n6751 gnd.n976 9.3005
R12252 gnd.n6752 gnd.n975 9.3005
R12253 gnd.n974 gnd.n970 9.3005
R12254 gnd.n6758 gnd.n969 9.3005
R12255 gnd.n6759 gnd.n968 9.3005
R12256 gnd.n6760 gnd.n967 9.3005
R12257 gnd.n966 gnd.n962 9.3005
R12258 gnd.n6766 gnd.n961 9.3005
R12259 gnd.n6767 gnd.n960 9.3005
R12260 gnd.n6768 gnd.n959 9.3005
R12261 gnd.n958 gnd.n954 9.3005
R12262 gnd.n6774 gnd.n953 9.3005
R12263 gnd.n6775 gnd.n952 9.3005
R12264 gnd.n6776 gnd.n951 9.3005
R12265 gnd.n950 gnd.n946 9.3005
R12266 gnd.n6782 gnd.n945 9.3005
R12267 gnd.n6783 gnd.n944 9.3005
R12268 gnd.n6784 gnd.n943 9.3005
R12269 gnd.n942 gnd.n938 9.3005
R12270 gnd.n6790 gnd.n937 9.3005
R12271 gnd.n6791 gnd.n936 9.3005
R12272 gnd.n6792 gnd.n935 9.3005
R12273 gnd.n934 gnd.n930 9.3005
R12274 gnd.n6798 gnd.n929 9.3005
R12275 gnd.n6799 gnd.n928 9.3005
R12276 gnd.n6800 gnd.n927 9.3005
R12277 gnd.n926 gnd.n922 9.3005
R12278 gnd.n6806 gnd.n921 9.3005
R12279 gnd.n6807 gnd.n920 9.3005
R12280 gnd.n6808 gnd.n919 9.3005
R12281 gnd.n918 gnd.n914 9.3005
R12282 gnd.n6814 gnd.n913 9.3005
R12283 gnd.n6815 gnd.n912 9.3005
R12284 gnd.n6816 gnd.n911 9.3005
R12285 gnd.n910 gnd.n906 9.3005
R12286 gnd.n6822 gnd.n905 9.3005
R12287 gnd.n6823 gnd.n904 9.3005
R12288 gnd.n6824 gnd.n903 9.3005
R12289 gnd.n902 gnd.n898 9.3005
R12290 gnd.n6830 gnd.n897 9.3005
R12291 gnd.n6831 gnd.n896 9.3005
R12292 gnd.n6832 gnd.n895 9.3005
R12293 gnd.n894 gnd.n890 9.3005
R12294 gnd.n6838 gnd.n889 9.3005
R12295 gnd.n6839 gnd.n888 9.3005
R12296 gnd.n6840 gnd.n887 9.3005
R12297 gnd.n886 gnd.n882 9.3005
R12298 gnd.n6846 gnd.n881 9.3005
R12299 gnd.n6847 gnd.n880 9.3005
R12300 gnd.n6848 gnd.n879 9.3005
R12301 gnd.n878 gnd.n874 9.3005
R12302 gnd.n6854 gnd.n873 9.3005
R12303 gnd.n6855 gnd.n872 9.3005
R12304 gnd.n6856 gnd.n871 9.3005
R12305 gnd.n870 gnd.n866 9.3005
R12306 gnd.n6862 gnd.n865 9.3005
R12307 gnd.n6863 gnd.n864 9.3005
R12308 gnd.n6864 gnd.n863 9.3005
R12309 gnd.n862 gnd.n858 9.3005
R12310 gnd.n6870 gnd.n857 9.3005
R12311 gnd.n6871 gnd.n856 9.3005
R12312 gnd.n6872 gnd.n855 9.3005
R12313 gnd.n851 gnd.n850 9.3005
R12314 gnd.n6879 gnd.n6878 9.3005
R12315 gnd.n6710 gnd.n1017 9.3005
R12316 gnd.n5937 gnd.n5936 9.3005
R12317 gnd.n5941 gnd.n5940 9.3005
R12318 gnd.n5924 gnd.n5921 9.3005
R12319 gnd.n5949 gnd.n5948 9.3005
R12320 gnd.n5953 gnd.n5952 9.3005
R12321 gnd.n5918 gnd.n5917 9.3005
R12322 gnd.n5961 gnd.n5960 9.3005
R12323 gnd.n5965 gnd.n5964 9.3005
R12324 gnd.n5912 gnd.n5909 9.3005
R12325 gnd.n5973 gnd.n5972 9.3005
R12326 gnd.n5977 gnd.n5976 9.3005
R12327 gnd.n5906 gnd.n5905 9.3005
R12328 gnd.n5986 gnd.n5985 9.3005
R12329 gnd.n5989 gnd.n5904 9.3005
R12330 gnd.n5994 gnd.n5993 9.3005
R12331 gnd.n5992 gnd.n5896 9.3005
R12332 gnd.n6000 gnd.n5893 9.3005
R12333 gnd.n6002 gnd.n6001 9.3005
R12334 gnd.n5930 gnd.n5929 9.3005
R12335 gnd.n5996 gnd.n5995 9.3005
R12336 gnd.n5984 gnd.n5901 9.3005
R12337 gnd.n5983 gnd.n5982 9.3005
R12338 gnd.n5979 gnd.n5978 9.3005
R12339 gnd.n5908 gnd.n5907 9.3005
R12340 gnd.n5971 gnd.n5970 9.3005
R12341 gnd.n5967 gnd.n5966 9.3005
R12342 gnd.n5916 gnd.n5913 9.3005
R12343 gnd.n5959 gnd.n5958 9.3005
R12344 gnd.n5955 gnd.n5954 9.3005
R12345 gnd.n5920 gnd.n5919 9.3005
R12346 gnd.n5947 gnd.n5946 9.3005
R12347 gnd.n5943 gnd.n5942 9.3005
R12348 gnd.n5928 gnd.n5925 9.3005
R12349 gnd.n5935 gnd.n5934 9.3005
R12350 gnd.n5931 gnd.n1479 9.3005
R12351 gnd.n5997 gnd.n5897 9.3005
R12352 gnd.n5999 gnd.n5998 9.3005
R12353 gnd.n6004 gnd.n6003 9.3005
R12354 gnd.n6007 gnd.n5892 9.3005
R12355 gnd.n6011 gnd.n6010 9.3005
R12356 gnd.n6012 gnd.n5891 9.3005
R12357 gnd.n6014 gnd.n6013 9.3005
R12358 gnd.n6017 gnd.n5888 9.3005
R12359 gnd.n6021 gnd.n6020 9.3005
R12360 gnd.n6022 gnd.n5886 9.3005
R12361 gnd.n6025 gnd.n6024 9.3005
R12362 gnd.n6023 gnd.n5887 9.3005
R12363 gnd.n4985 gnd.n4984 9.3005
R12364 gnd.n4986 gnd.n2305 9.3005
R12365 gnd.n4988 gnd.n4987 9.3005
R12366 gnd.n2292 gnd.n2291 9.3005
R12367 gnd.n5001 gnd.n5000 9.3005
R12368 gnd.n5002 gnd.n2290 9.3005
R12369 gnd.n5004 gnd.n5003 9.3005
R12370 gnd.n2279 gnd.n2278 9.3005
R12371 gnd.n5017 gnd.n5016 9.3005
R12372 gnd.n5018 gnd.n2277 9.3005
R12373 gnd.n5020 gnd.n5019 9.3005
R12374 gnd.n2265 gnd.n2264 9.3005
R12375 gnd.n5033 gnd.n5032 9.3005
R12376 gnd.n5034 gnd.n2263 9.3005
R12377 gnd.n5036 gnd.n5035 9.3005
R12378 gnd.n2251 gnd.n2250 9.3005
R12379 gnd.n5049 gnd.n5048 9.3005
R12380 gnd.n5050 gnd.n2249 9.3005
R12381 gnd.n5052 gnd.n5051 9.3005
R12382 gnd.n2237 gnd.n2236 9.3005
R12383 gnd.n5065 gnd.n5064 9.3005
R12384 gnd.n5066 gnd.n2234 9.3005
R12385 gnd.n5079 gnd.n5078 9.3005
R12386 gnd.n5077 gnd.n2235 9.3005
R12387 gnd.n5076 gnd.n5075 9.3005
R12388 gnd.n5074 gnd.n5067 9.3005
R12389 gnd.n5073 gnd.n5072 9.3005
R12390 gnd.n5071 gnd.n5070 9.3005
R12391 gnd.n1383 gnd.n1381 9.3005
R12392 gnd.n6464 gnd.n6463 9.3005
R12393 gnd.n6462 gnd.n1382 9.3005
R12394 gnd.n6461 gnd.n6460 9.3005
R12395 gnd.n6459 gnd.n1384 9.3005
R12396 gnd.n6458 gnd.n6457 9.3005
R12397 gnd.n6456 gnd.n1388 9.3005
R12398 gnd.n6455 gnd.n6454 9.3005
R12399 gnd.n6453 gnd.n1389 9.3005
R12400 gnd.n6452 gnd.n6451 9.3005
R12401 gnd.n6450 gnd.n1393 9.3005
R12402 gnd.n6449 gnd.n6448 9.3005
R12403 gnd.n6447 gnd.n1394 9.3005
R12404 gnd.n6446 gnd.n6445 9.3005
R12405 gnd.n6444 gnd.n1398 9.3005
R12406 gnd.n6443 gnd.n6442 9.3005
R12407 gnd.n6441 gnd.n1399 9.3005
R12408 gnd.n6440 gnd.n6439 9.3005
R12409 gnd.n6438 gnd.n1403 9.3005
R12410 gnd.n6437 gnd.n6436 9.3005
R12411 gnd.n6435 gnd.n1404 9.3005
R12412 gnd.n6434 gnd.n6433 9.3005
R12413 gnd.n6432 gnd.n1408 9.3005
R12414 gnd.n6431 gnd.n6430 9.3005
R12415 gnd.n6429 gnd.n1409 9.3005
R12416 gnd.n6428 gnd.n6427 9.3005
R12417 gnd.n6426 gnd.n1413 9.3005
R12418 gnd.n6425 gnd.n6424 9.3005
R12419 gnd.n6423 gnd.n1414 9.3005
R12420 gnd.n6422 gnd.n6421 9.3005
R12421 gnd.n6420 gnd.n1418 9.3005
R12422 gnd.n6419 gnd.n6418 9.3005
R12423 gnd.n6417 gnd.n1419 9.3005
R12424 gnd.n6416 gnd.n6415 9.3005
R12425 gnd.n6414 gnd.n1423 9.3005
R12426 gnd.n6413 gnd.n6412 9.3005
R12427 gnd.n6411 gnd.n1424 9.3005
R12428 gnd.n6410 gnd.n6409 9.3005
R12429 gnd.n6408 gnd.n1428 9.3005
R12430 gnd.n6407 gnd.n6406 9.3005
R12431 gnd.n6405 gnd.n1429 9.3005
R12432 gnd.n6404 gnd.n6403 9.3005
R12433 gnd.n6402 gnd.n1433 9.3005
R12434 gnd.n6401 gnd.n6400 9.3005
R12435 gnd.n6399 gnd.n1434 9.3005
R12436 gnd.n6398 gnd.n6397 9.3005
R12437 gnd.n6396 gnd.n1438 9.3005
R12438 gnd.n6395 gnd.n6394 9.3005
R12439 gnd.n6393 gnd.n1439 9.3005
R12440 gnd.n6392 gnd.n6391 9.3005
R12441 gnd.n6390 gnd.n1443 9.3005
R12442 gnd.n6389 gnd.n6388 9.3005
R12443 gnd.n6387 gnd.n1444 9.3005
R12444 gnd.n6386 gnd.n6385 9.3005
R12445 gnd.n6384 gnd.n1448 9.3005
R12446 gnd.n6383 gnd.n6382 9.3005
R12447 gnd.n6381 gnd.n1449 9.3005
R12448 gnd.n6380 gnd.n6379 9.3005
R12449 gnd.n6378 gnd.n1453 9.3005
R12450 gnd.n6377 gnd.n6376 9.3005
R12451 gnd.n6375 gnd.n1454 9.3005
R12452 gnd.n6374 gnd.n6373 9.3005
R12453 gnd.n6372 gnd.n1458 9.3005
R12454 gnd.n6371 gnd.n6370 9.3005
R12455 gnd.n6369 gnd.n1459 9.3005
R12456 gnd.n6368 gnd.n6367 9.3005
R12457 gnd.n6366 gnd.n1463 9.3005
R12458 gnd.n6365 gnd.n6364 9.3005
R12459 gnd.n6363 gnd.n1464 9.3005
R12460 gnd.n6362 gnd.n6361 9.3005
R12461 gnd.n6360 gnd.n1468 9.3005
R12462 gnd.n6359 gnd.n6358 9.3005
R12463 gnd.n6357 gnd.n1469 9.3005
R12464 gnd.n2307 gnd.n2306 9.3005
R12465 gnd.n4855 gnd.n4854 9.3005
R12466 gnd.n4856 gnd.n4847 9.3005
R12467 gnd.n4858 gnd.n4857 9.3005
R12468 gnd.n4860 gnd.n4859 9.3005
R12469 gnd.n4861 gnd.n4840 9.3005
R12470 gnd.n4863 gnd.n4862 9.3005
R12471 gnd.n4864 gnd.n4839 9.3005
R12472 gnd.n4866 gnd.n4865 9.3005
R12473 gnd.n4867 gnd.n4834 9.3005
R12474 gnd.n4853 gnd.n4852 9.3005
R12475 gnd.n2531 gnd.n2530 9.3005
R12476 gnd.n4633 gnd.n4632 9.3005
R12477 gnd.n4634 gnd.n2529 9.3005
R12478 gnd.n4636 gnd.n4635 9.3005
R12479 gnd.n2516 gnd.n2514 9.3005
R12480 gnd.n4674 gnd.n4673 9.3005
R12481 gnd.n4672 gnd.n2515 9.3005
R12482 gnd.n4671 gnd.n4670 9.3005
R12483 gnd.n4669 gnd.n2517 9.3005
R12484 gnd.n4668 gnd.n4667 9.3005
R12485 gnd.n4666 gnd.n2520 9.3005
R12486 gnd.n4665 gnd.n4664 9.3005
R12487 gnd.n2500 gnd.n2499 9.3005
R12488 gnd.n4716 gnd.n4715 9.3005
R12489 gnd.n4717 gnd.n2498 9.3005
R12490 gnd.n4719 gnd.n4718 9.3005
R12491 gnd.n2494 gnd.n2493 9.3005
R12492 gnd.n4732 gnd.n4731 9.3005
R12493 gnd.n4733 gnd.n2492 9.3005
R12494 gnd.n4735 gnd.n4734 9.3005
R12495 gnd.n2478 gnd.n2476 9.3005
R12496 gnd.n4886 gnd.n4885 9.3005
R12497 gnd.n4884 gnd.n2477 9.3005
R12498 gnd.n4883 gnd.n4882 9.3005
R12499 gnd.n4881 gnd.n2479 9.3005
R12500 gnd.n4880 gnd.n4879 9.3005
R12501 gnd.n4878 gnd.n2482 9.3005
R12502 gnd.n4877 gnd.n4876 9.3005
R12503 gnd.n4875 gnd.n2483 9.3005
R12504 gnd.n4874 gnd.n4873 9.3005
R12505 gnd.n4872 gnd.n4833 9.3005
R12506 gnd.n4871 gnd.n2459 9.3005
R12507 gnd.n4869 gnd.n4868 9.3005
R12508 gnd.n2458 gnd.n2457 9.3005
R12509 gnd.n4929 gnd.n4928 9.3005
R12510 gnd.n4931 gnd.n4930 9.3005
R12511 gnd.n2444 gnd.n2443 9.3005
R12512 gnd.n4937 gnd.n4936 9.3005
R12513 gnd.n4939 gnd.n4938 9.3005
R12514 gnd.n2436 gnd.n2435 9.3005
R12515 gnd.n4945 gnd.n4944 9.3005
R12516 gnd.n4947 gnd.n4946 9.3005
R12517 gnd.n2424 gnd.n2423 9.3005
R12518 gnd.n4953 gnd.n4952 9.3005
R12519 gnd.n4955 gnd.n4954 9.3005
R12520 gnd.n2416 gnd.n2415 9.3005
R12521 gnd.n4961 gnd.n4960 9.3005
R12522 gnd.n4963 gnd.n4962 9.3005
R12523 gnd.n2336 gnd.n2334 9.3005
R12524 gnd.n4969 gnd.n4968 9.3005
R12525 gnd.n4970 gnd.n2333 9.3005
R12526 gnd.n2404 gnd.n2403 9.3005
R12527 gnd.n2405 gnd.n2335 9.3005
R12528 gnd.n4967 gnd.n4966 9.3005
R12529 gnd.n4965 gnd.n4964 9.3005
R12530 gnd.n2411 gnd.n2410 9.3005
R12531 gnd.n4959 gnd.n4958 9.3005
R12532 gnd.n4957 gnd.n4956 9.3005
R12533 gnd.n2420 gnd.n2419 9.3005
R12534 gnd.n4951 gnd.n4950 9.3005
R12535 gnd.n4949 gnd.n4948 9.3005
R12536 gnd.n2430 gnd.n2429 9.3005
R12537 gnd.n4943 gnd.n4942 9.3005
R12538 gnd.n4941 gnd.n4940 9.3005
R12539 gnd.n2440 gnd.n2439 9.3005
R12540 gnd.n4935 gnd.n4934 9.3005
R12541 gnd.n4933 gnd.n4932 9.3005
R12542 gnd.n2452 gnd.n2451 9.3005
R12543 gnd.n4927 gnd.n4926 9.3005
R12544 gnd.n2399 gnd.n2341 9.3005
R12545 gnd.n2398 gnd.n2397 9.3005
R12546 gnd.n2396 gnd.n2343 9.3005
R12547 gnd.n2395 gnd.n2394 9.3005
R12548 gnd.n2393 gnd.n2344 9.3005
R12549 gnd.n2392 gnd.n2391 9.3005
R12550 gnd.n2390 gnd.n2347 9.3005
R12551 gnd.n2389 gnd.n2388 9.3005
R12552 gnd.n2387 gnd.n2348 9.3005
R12553 gnd.n2386 gnd.n2385 9.3005
R12554 gnd.n2384 gnd.n2351 9.3005
R12555 gnd.n2383 gnd.n2382 9.3005
R12556 gnd.n2381 gnd.n2352 9.3005
R12557 gnd.n2380 gnd.n2379 9.3005
R12558 gnd.n2378 gnd.n2355 9.3005
R12559 gnd.n2377 gnd.n2376 9.3005
R12560 gnd.n2375 gnd.n2356 9.3005
R12561 gnd.n2374 gnd.n2373 9.3005
R12562 gnd.n2372 gnd.n2359 9.3005
R12563 gnd.n2371 gnd.n2370 9.3005
R12564 gnd.n2369 gnd.n2360 9.3005
R12565 gnd.n2368 gnd.n2367 9.3005
R12566 gnd.n2366 gnd.n2363 9.3005
R12567 gnd.n2365 gnd.n2364 9.3005
R12568 gnd.n2220 gnd.n2219 9.3005
R12569 gnd.n5097 gnd.n5096 9.3005
R12570 gnd.n5098 gnd.n2218 9.3005
R12571 gnd.n5100 gnd.n5099 9.3005
R12572 gnd.n5198 gnd.n2217 9.3005
R12573 gnd.n5200 gnd.n5199 9.3005
R12574 gnd.n5201 gnd.n2215 9.3005
R12575 gnd.n5239 gnd.n5238 9.3005
R12576 gnd.n5237 gnd.n2216 9.3005
R12577 gnd.n5236 gnd.n5235 9.3005
R12578 gnd.n5234 gnd.n5202 9.3005
R12579 gnd.n5233 gnd.n5232 9.3005
R12580 gnd.n5231 gnd.n5205 9.3005
R12581 gnd.n5230 gnd.n5229 9.3005
R12582 gnd.n5228 gnd.n5206 9.3005
R12583 gnd.n5227 gnd.n5226 9.3005
R12584 gnd.n5225 gnd.n5209 9.3005
R12585 gnd.n5224 gnd.n5223 9.3005
R12586 gnd.n5222 gnd.n5210 9.3005
R12587 gnd.n5221 gnd.n5220 9.3005
R12588 gnd.n5219 gnd.n5212 9.3005
R12589 gnd.n5218 gnd.n5217 9.3005
R12590 gnd.n5216 gnd.n5213 9.3005
R12591 gnd.n2120 gnd.n2119 9.3005
R12592 gnd.n5382 gnd.n5381 9.3005
R12593 gnd.n5383 gnd.n2117 9.3005
R12594 gnd.n5399 gnd.n5398 9.3005
R12595 gnd.n5397 gnd.n2118 9.3005
R12596 gnd.n5396 gnd.n5395 9.3005
R12597 gnd.n5394 gnd.n5384 9.3005
R12598 gnd.n5393 gnd.n5392 9.3005
R12599 gnd.n5391 gnd.n5388 9.3005
R12600 gnd.n5390 gnd.n5389 9.3005
R12601 gnd.n2067 gnd.n2066 9.3005
R12602 gnd.n5463 gnd.n5462 9.3005
R12603 gnd.n5464 gnd.n2065 9.3005
R12604 gnd.n5466 gnd.n5465 9.3005
R12605 gnd.n5467 gnd.n2064 9.3005
R12606 gnd.n5471 gnd.n5470 9.3005
R12607 gnd.n5472 gnd.n2062 9.3005
R12608 gnd.n5497 gnd.n5496 9.3005
R12609 gnd.n5495 gnd.n2063 9.3005
R12610 gnd.n5494 gnd.n5493 9.3005
R12611 gnd.n5492 gnd.n5473 9.3005
R12612 gnd.n5491 gnd.n5490 9.3005
R12613 gnd.n5489 gnd.n5476 9.3005
R12614 gnd.n5488 gnd.n5487 9.3005
R12615 gnd.n5486 gnd.n5477 9.3005
R12616 gnd.n5485 gnd.n5484 9.3005
R12617 gnd.n5483 gnd.n5480 9.3005
R12618 gnd.n5482 gnd.n5481 9.3005
R12619 gnd.n1791 gnd.n1790 9.3005
R12620 gnd.n5768 gnd.n5767 9.3005
R12621 gnd.n5769 gnd.n1789 9.3005
R12622 gnd.n5771 gnd.n5770 9.3005
R12623 gnd.n1780 gnd.n1779 9.3005
R12624 gnd.n5786 gnd.n5785 9.3005
R12625 gnd.n5787 gnd.n1778 9.3005
R12626 gnd.n5789 gnd.n5788 9.3005
R12627 gnd.n1768 gnd.n1767 9.3005
R12628 gnd.n5803 gnd.n5802 9.3005
R12629 gnd.n5804 gnd.n1766 9.3005
R12630 gnd.n5806 gnd.n5805 9.3005
R12631 gnd.n1756 gnd.n1755 9.3005
R12632 gnd.n5820 gnd.n5819 9.3005
R12633 gnd.n5821 gnd.n1754 9.3005
R12634 gnd.n5823 gnd.n5822 9.3005
R12635 gnd.n1743 gnd.n1742 9.3005
R12636 gnd.n5837 gnd.n5836 9.3005
R12637 gnd.n5838 gnd.n1741 9.3005
R12638 gnd.n5840 gnd.n5839 9.3005
R12639 gnd.n1732 gnd.n1731 9.3005
R12640 gnd.n5856 gnd.n5855 9.3005
R12641 gnd.n5857 gnd.n1730 9.3005
R12642 gnd.n5859 gnd.n5858 9.3005
R12643 gnd.n1478 gnd.n1477 9.3005
R12644 gnd.n6353 gnd.n6352 9.3005
R12645 gnd.n2401 gnd.n2400 9.3005
R12646 gnd.n6347 gnd.n1481 9.3005
R12647 gnd.n6346 gnd.n6345 9.3005
R12648 gnd.n6344 gnd.n1485 9.3005
R12649 gnd.n6343 gnd.n6342 9.3005
R12650 gnd.n6341 gnd.n1486 9.3005
R12651 gnd.n6340 gnd.n6339 9.3005
R12652 gnd.n6338 gnd.n1490 9.3005
R12653 gnd.n6337 gnd.n6336 9.3005
R12654 gnd.n6335 gnd.n1491 9.3005
R12655 gnd.n6334 gnd.n6333 9.3005
R12656 gnd.n6332 gnd.n1495 9.3005
R12657 gnd.n6331 gnd.n6330 9.3005
R12658 gnd.n6329 gnd.n1496 9.3005
R12659 gnd.n6328 gnd.n6327 9.3005
R12660 gnd.n6326 gnd.n1500 9.3005
R12661 gnd.n6325 gnd.n6324 9.3005
R12662 gnd.n6323 gnd.n1501 9.3005
R12663 gnd.n6322 gnd.n6321 9.3005
R12664 gnd.n6320 gnd.n1505 9.3005
R12665 gnd.n6319 gnd.n6318 9.3005
R12666 gnd.n6317 gnd.n1506 9.3005
R12667 gnd.n6316 gnd.n6315 9.3005
R12668 gnd.n6314 gnd.n1510 9.3005
R12669 gnd.n6313 gnd.n6312 9.3005
R12670 gnd.n6311 gnd.n1511 9.3005
R12671 gnd.n6310 gnd.n6309 9.3005
R12672 gnd.n6308 gnd.n6307 9.3005
R12673 gnd.n328 gnd.n326 9.3005
R12674 gnd.n7661 gnd.n7660 9.3005
R12675 gnd.n7659 gnd.n327 9.3005
R12676 gnd.n7658 gnd.n7657 9.3005
R12677 gnd.n7656 gnd.n329 9.3005
R12678 gnd.n7655 gnd.n7654 9.3005
R12679 gnd.n7653 gnd.n333 9.3005
R12680 gnd.n7652 gnd.n7651 9.3005
R12681 gnd.n304 gnd.n303 9.3005
R12682 gnd.n7674 gnd.n7673 9.3005
R12683 gnd.n7675 gnd.n302 9.3005
R12684 gnd.n7677 gnd.n7676 9.3005
R12685 gnd.n289 gnd.n288 9.3005
R12686 gnd.n7690 gnd.n7689 9.3005
R12687 gnd.n7691 gnd.n287 9.3005
R12688 gnd.n7693 gnd.n7692 9.3005
R12689 gnd.n273 gnd.n272 9.3005
R12690 gnd.n7706 gnd.n7705 9.3005
R12691 gnd.n7707 gnd.n271 9.3005
R12692 gnd.n7709 gnd.n7708 9.3005
R12693 gnd.n257 gnd.n256 9.3005
R12694 gnd.n7722 gnd.n7721 9.3005
R12695 gnd.n7723 gnd.n255 9.3005
R12696 gnd.n7725 gnd.n7724 9.3005
R12697 gnd.n241 gnd.n240 9.3005
R12698 gnd.n7738 gnd.n7737 9.3005
R12699 gnd.n7739 gnd.n239 9.3005
R12700 gnd.n7741 gnd.n7740 9.3005
R12701 gnd.n227 gnd.n226 9.3005
R12702 gnd.n7754 gnd.n7753 9.3005
R12703 gnd.n7755 gnd.n225 9.3005
R12704 gnd.n7757 gnd.n7756 9.3005
R12705 gnd.n210 gnd.n209 9.3005
R12706 gnd.n7772 gnd.n7771 9.3005
R12707 gnd.n7773 gnd.n207 9.3005
R12708 gnd.n7836 gnd.n7835 9.3005
R12709 gnd.n7834 gnd.n208 9.3005
R12710 gnd.n6349 gnd.n6348 9.3005
R12711 gnd.n7831 gnd.n7774 9.3005
R12712 gnd.n7830 gnd.n7829 9.3005
R12713 gnd.n7828 gnd.n7779 9.3005
R12714 gnd.n7827 gnd.n7826 9.3005
R12715 gnd.n7825 gnd.n7780 9.3005
R12716 gnd.n7824 gnd.n7823 9.3005
R12717 gnd.n7822 gnd.n7787 9.3005
R12718 gnd.n7821 gnd.n7820 9.3005
R12719 gnd.n7819 gnd.n7788 9.3005
R12720 gnd.n7818 gnd.n7817 9.3005
R12721 gnd.n7816 gnd.n7795 9.3005
R12722 gnd.n7815 gnd.n7814 9.3005
R12723 gnd.n7813 gnd.n7796 9.3005
R12724 gnd.n7812 gnd.n7811 9.3005
R12725 gnd.n7810 gnd.n7803 9.3005
R12726 gnd.n7809 gnd.n7808 9.3005
R12727 gnd.n124 gnd.n121 9.3005
R12728 gnd.n7921 gnd.n7920 9.3005
R12729 gnd.n7833 gnd.n7832 9.3005
R12730 gnd.n6056 gnd.n1678 9.3005
R12731 gnd.n6059 gnd.n6058 9.3005
R12732 gnd.n6057 gnd.n1679 9.3005
R12733 gnd.n1654 gnd.n1653 9.3005
R12734 gnd.n6087 gnd.n6086 9.3005
R12735 gnd.n6088 gnd.n1651 9.3005
R12736 gnd.n6091 gnd.n6090 9.3005
R12737 gnd.n6089 gnd.n1652 9.3005
R12738 gnd.n1628 gnd.n1627 9.3005
R12739 gnd.n6119 gnd.n6118 9.3005
R12740 gnd.n6120 gnd.n1625 9.3005
R12741 gnd.n6123 gnd.n6122 9.3005
R12742 gnd.n6121 gnd.n1626 9.3005
R12743 gnd.n1598 gnd.n1597 9.3005
R12744 gnd.n6157 gnd.n6156 9.3005
R12745 gnd.n6158 gnd.n1595 9.3005
R12746 gnd.n6161 gnd.n6160 9.3005
R12747 gnd.n6159 gnd.n1596 9.3005
R12748 gnd.n1565 gnd.n1564 9.3005
R12749 gnd.n6223 gnd.n6222 9.3005
R12750 gnd.n6224 gnd.n1562 9.3005
R12751 gnd.n6229 gnd.n6228 9.3005
R12752 gnd.n6227 gnd.n1563 9.3005
R12753 gnd.n6226 gnd.n6225 9.3005
R12754 gnd.n1526 gnd.n1524 9.3005
R12755 gnd.n6300 gnd.n6299 9.3005
R12756 gnd.n6298 gnd.n1525 9.3005
R12757 gnd.n6297 gnd.n6296 9.3005
R12758 gnd.n6295 gnd.n1527 9.3005
R12759 gnd.n6294 gnd.n6293 9.3005
R12760 gnd.n6292 gnd.n79 9.3005
R12761 gnd.n7970 gnd.n80 9.3005
R12762 gnd.n7969 gnd.n7968 9.3005
R12763 gnd.n7967 gnd.n81 9.3005
R12764 gnd.n7966 gnd.n7965 9.3005
R12765 gnd.n7964 gnd.n85 9.3005
R12766 gnd.n7963 gnd.n7962 9.3005
R12767 gnd.n7961 gnd.n86 9.3005
R12768 gnd.n7960 gnd.n7959 9.3005
R12769 gnd.n7958 gnd.n90 9.3005
R12770 gnd.n7957 gnd.n7956 9.3005
R12771 gnd.n7955 gnd.n91 9.3005
R12772 gnd.n7954 gnd.n7953 9.3005
R12773 gnd.n7952 gnd.n95 9.3005
R12774 gnd.n7951 gnd.n7950 9.3005
R12775 gnd.n7949 gnd.n96 9.3005
R12776 gnd.n7948 gnd.n7947 9.3005
R12777 gnd.n7946 gnd.n100 9.3005
R12778 gnd.n7945 gnd.n7944 9.3005
R12779 gnd.n7943 gnd.n101 9.3005
R12780 gnd.n7942 gnd.n7941 9.3005
R12781 gnd.n7940 gnd.n105 9.3005
R12782 gnd.n7939 gnd.n7938 9.3005
R12783 gnd.n7937 gnd.n106 9.3005
R12784 gnd.n7936 gnd.n7935 9.3005
R12785 gnd.n7934 gnd.n110 9.3005
R12786 gnd.n7933 gnd.n7932 9.3005
R12787 gnd.n7931 gnd.n111 9.3005
R12788 gnd.n7930 gnd.n7929 9.3005
R12789 gnd.n7928 gnd.n115 9.3005
R12790 gnd.n7927 gnd.n7926 9.3005
R12791 gnd.n7925 gnd.n116 9.3005
R12792 gnd.n7924 gnd.n7923 9.3005
R12793 gnd.n7922 gnd.n120 9.3005
R12794 gnd.n6055 gnd.n6054 9.3005
R12795 gnd.t315 gnd.n2864 9.24152
R12796 gnd.n2765 gnd.t197 9.24152
R12797 gnd.n4046 gnd.t183 9.24152
R12798 gnd.t143 gnd.n1019 9.24152
R12799 gnd.n7719 gnd.t14 9.24152
R12800 gnd.t348 gnd.t315 8.92286
R12801 gnd.n5298 gnd.n2174 8.92286
R12802 gnd.n5331 gnd.n2145 8.92286
R12803 gnd.n5442 gnd.n2087 8.92286
R12804 gnd.n5514 gnd.n2044 8.92286
R12805 gnd.n5590 gnd.n1991 8.92286
R12806 gnd.n1992 gnd.t211 8.92286
R12807 gnd.n4016 gnd.n3991 8.92171
R12808 gnd.n3984 gnd.n3959 8.92171
R12809 gnd.n3952 gnd.n3927 8.92171
R12810 gnd.n3921 gnd.n3896 8.92171
R12811 gnd.n3889 gnd.n3864 8.92171
R12812 gnd.n3857 gnd.n3832 8.92171
R12813 gnd.n3825 gnd.n3800 8.92171
R12814 gnd.n3794 gnd.n3769 8.92171
R12815 gnd.n5613 gnd.n5595 8.72777
R12816 gnd.n3520 gnd.t97 8.60421
R12817 gnd.t50 gnd.n2642 8.60421
R12818 gnd.n7751 gnd.t114 8.60421
R12819 gnd.n2944 gnd.n2924 8.43467
R12820 gnd.n58 gnd.n38 8.43467
R12821 gnd.n4577 gnd.n0 8.41456
R12822 gnd.n7971 gnd.n7970 8.41456
R12823 gnd.n4017 gnd.n3989 8.14595
R12824 gnd.n3985 gnd.n3957 8.14595
R12825 gnd.n3953 gnd.n3925 8.14595
R12826 gnd.n3922 gnd.n3894 8.14595
R12827 gnd.n3890 gnd.n3862 8.14595
R12828 gnd.n3858 gnd.n3830 8.14595
R12829 gnd.n3826 gnd.n3798 8.14595
R12830 gnd.n3795 gnd.n3767 8.14595
R12831 gnd.n4022 gnd.n4021 7.97301
R12832 gnd.t96 gnd.n3035 7.9669
R12833 gnd.n4973 gnd.n2316 7.9669
R12834 gnd.n6029 gnd.n6028 7.9669
R12835 gnd.n7920 gnd.n124 7.75808
R12836 gnd.n5998 gnd.n5997 7.75808
R12837 gnd.n4926 gnd.n2451 7.75808
R12838 gnd.n4401 gnd.n4352 7.75808
R12839 gnd.n1032 gnd.n1022 7.64824
R12840 gnd.n6701 gnd.n1035 7.64824
R12841 gnd.n4521 gnd.n1044 7.64824
R12842 gnd.n4529 gnd.n1054 7.64824
R12843 gnd.n6689 gnd.n1057 7.64824
R12844 gnd.n4542 gnd.n1065 7.64824
R12845 gnd.n6683 gnd.n1068 7.64824
R12846 gnd.n4552 gnd.n4551 7.64824
R12847 gnd.n6677 gnd.n1078 7.64824
R12848 gnd.n4569 gnd.n1086 7.64824
R12849 gnd.n4563 gnd.n2551 7.64824
R12850 gnd.n4590 gnd.n4582 7.64824
R12851 gnd.n4598 gnd.n2548 7.64824
R12852 gnd.n4597 gnd.n2542 7.64824
R12853 gnd.n4616 gnd.n4615 7.64824
R12854 gnd.n4630 gnd.n2534 7.64824
R12855 gnd.n4625 gnd.n2537 7.64824
R12856 gnd.n4638 gnd.n1101 7.64824
R12857 gnd.n6663 gnd.n1104 7.64824
R12858 gnd.n4677 gnd.n4676 7.64824
R12859 gnd.n6657 gnd.n1115 7.64824
R12860 gnd.n4646 gnd.n1122 7.64824
R12861 gnd.n6651 gnd.n1125 7.64824
R12862 gnd.n4650 gnd.n1133 7.64824
R12863 gnd.n6645 gnd.n1136 7.64824
R12864 gnd.n4662 gnd.n1144 7.64824
R12865 gnd.n6639 gnd.n1147 7.64824
R12866 gnd.n4713 gnd.n4712 7.64824
R12867 gnd.n6633 gnd.n1157 7.64824
R12868 gnd.n4721 gnd.n1165 7.64824
R12869 gnd.n6627 gnd.n1168 7.64824
R12870 gnd.n4729 gnd.n1176 7.64824
R12871 gnd.n6621 gnd.n1179 7.64824
R12872 gnd.n4737 gnd.n1187 7.64824
R12873 gnd.n6615 gnd.n1190 7.64824
R12874 gnd.n4889 gnd.n4888 7.64824
R12875 gnd.n6609 gnd.n1200 7.64824
R12876 gnd.n4745 gnd.n1208 7.64824
R12877 gnd.n6603 gnd.n1211 7.64824
R12878 gnd.n4751 gnd.n1219 7.64824
R12879 gnd.n6597 gnd.n1222 7.64824
R12880 gnd.n4755 gnd.n1230 7.64824
R12881 gnd.n6591 gnd.n1233 7.64824
R12882 gnd.n6585 gnd.n1244 7.64824
R12883 gnd.n4923 gnd.n4922 7.64824
R12884 gnd.n6466 gnd.n1376 7.64824
R12885 gnd.n5280 gnd.n2187 7.64824
R12886 gnd.n5356 gnd.t70 7.64824
R12887 gnd.n5369 gnd.n2131 7.64824
R12888 gnd.n5420 gnd.n2101 7.64824
R12889 gnd.n5427 gnd.t65 7.64824
R12890 gnd.n5521 gnd.n2033 7.64824
R12891 gnd.n5582 gnd.n5580 7.64824
R12892 gnd.n6052 gnd.n1682 7.64824
R12893 gnd.n1684 gnd.n1675 7.64824
R12894 gnd.n6074 gnd.n1665 7.64824
R12895 gnd.n6072 gnd.n1668 7.64824
R12896 gnd.n6084 gnd.n1656 7.64824
R12897 gnd.n1931 gnd.n1658 7.64824
R12898 gnd.n6095 gnd.n6094 7.64824
R12899 gnd.n6106 gnd.n1639 7.64824
R12900 gnd.n6105 gnd.n1642 7.64824
R12901 gnd.n6116 gnd.n1630 7.64824
R12902 gnd.n1632 gnd.n1622 7.64824
R12903 gnd.n6126 gnd.n6125 7.64824
R12904 gnd.n6144 gnd.n1611 7.64824
R12905 gnd.n6143 gnd.n1614 7.64824
R12906 gnd.n6154 gnd.n1600 7.64824
R12907 gnd.n1605 gnd.n1602 7.64824
R12908 gnd.n6163 gnd.n1593 7.64824
R12909 gnd.n6212 gnd.n1574 7.64824
R12910 gnd.n6211 gnd.n1578 7.64824
R12911 gnd.n6220 gnd.n1567 7.64824
R12912 gnd.n6205 gnd.n6204 7.64824
R12913 gnd.n6232 gnd.n1558 7.64824
R12914 gnd.n6231 gnd.n1549 7.64824
R12915 gnd.n6243 gnd.n6242 7.64824
R12916 gnd.n6195 gnd.n1552 7.64824
R12917 gnd.n6302 gnd.n1521 7.64824
R12918 gnd.n6305 gnd.n1515 7.64824
R12919 gnd.n6190 gnd.n1518 7.64824
R12920 gnd.n7663 gnd.n320 7.64824
R12921 gnd.n6186 gnd.n323 7.64824
R12922 gnd.n6290 gnd.n1531 7.64824
R12923 gnd.n6285 gnd.n1533 7.64824
R12924 gnd.n6284 gnd.n1537 7.64824
R12925 gnd.n7644 gnd.n339 7.64824
R12926 gnd.n7649 gnd.n335 7.64824
R12927 gnd.n7671 gnd.n306 7.64824
R12928 gnd.n7633 gnd.n308 7.64824
R12929 gnd.n7679 gnd.n298 7.64824
R12930 gnd.n7629 gnd.n300 7.64824
R12931 gnd.n7687 gnd.n291 7.64824
R12932 gnd.n7624 gnd.n7623 7.64824
R12933 gnd.n7695 gnd.n283 7.64824
R12934 gnd.n7703 gnd.n275 7.64824
R12935 gnd.n393 gnd.n277 7.64824
R12936 gnd.n7711 gnd.n266 7.64824
R12937 gnd.n3429 gnd.t13 7.32958
R12938 gnd.n4562 gnd.t40 7.32958
R12939 gnd.t193 gnd.n2302 7.32958
R12940 gnd.n5022 gnd.t35 7.32958
R12941 gnd.t92 gnd.n1752 7.32958
R12942 gnd.n5862 gnd.t165 7.32958
R12943 gnd.t58 gnd.n337 7.32958
R12944 gnd.n1358 gnd.n1357 7.30353
R12945 gnd.n5612 gnd.n5611 7.30353
R12946 gnd.n3389 gnd.n3108 7.01093
R12947 gnd.n3111 gnd.n3109 7.01093
R12948 gnd.n3399 gnd.n3398 7.01093
R12949 gnd.n3410 gnd.n3092 7.01093
R12950 gnd.n3409 gnd.n3095 7.01093
R12951 gnd.n3420 gnd.n3083 7.01093
R12952 gnd.n3086 gnd.n3084 7.01093
R12953 gnd.n3430 gnd.n3429 7.01093
R12954 gnd.n3440 gnd.n3064 7.01093
R12955 gnd.n3439 gnd.n3067 7.01093
R12956 gnd.n3448 gnd.n3058 7.01093
R12957 gnd.n3460 gnd.n3048 7.01093
R12958 gnd.n3470 gnd.n3033 7.01093
R12959 gnd.n3486 gnd.n3485 7.01093
R12960 gnd.n3035 gnd.n2972 7.01093
R12961 gnd.n3540 gnd.n2973 7.01093
R12962 gnd.n3534 gnd.n3533 7.01093
R12963 gnd.n3022 gnd.n2984 7.01093
R12964 gnd.n3526 gnd.n2995 7.01093
R12965 gnd.n3013 gnd.n3008 7.01093
R12966 gnd.n3520 gnd.n3519 7.01093
R12967 gnd.n3566 gnd.n2899 7.01093
R12968 gnd.n3565 gnd.n3564 7.01093
R12969 gnd.n3577 gnd.n3576 7.01093
R12970 gnd.n2892 gnd.n2884 7.01093
R12971 gnd.n3606 gnd.n2872 7.01093
R12972 gnd.n3605 gnd.n2875 7.01093
R12973 gnd.n3616 gnd.n2864 7.01093
R12974 gnd.n2865 gnd.n2853 7.01093
R12975 gnd.n3627 gnd.n2854 7.01093
R12976 gnd.n3651 gnd.n2845 7.01093
R12977 gnd.n3650 gnd.n2836 7.01093
R12978 gnd.n3673 gnd.n3672 7.01093
R12979 gnd.n3691 gnd.n2817 7.01093
R12980 gnd.n3690 gnd.n2820 7.01093
R12981 gnd.n3701 gnd.n2809 7.01093
R12982 gnd.n2810 gnd.n2797 7.01093
R12983 gnd.n3712 gnd.n2798 7.01093
R12984 gnd.n3739 gnd.n2781 7.01093
R12985 gnd.n3751 gnd.n3750 7.01093
R12986 gnd.n3733 gnd.n2774 7.01093
R12987 gnd.n3762 gnd.n3761 7.01093
R12988 gnd.n4034 gnd.n2762 7.01093
R12989 gnd.n4033 gnd.n2765 7.01093
R12990 gnd.n4046 gnd.n2754 7.01093
R12991 gnd.n2755 gnd.n2747 7.01093
R12992 gnd.n4056 gnd.n2673 7.01093
R12993 gnd.n2153 gnd.t311 7.01093
R12994 gnd.t24 gnd.n2079 7.01093
R12995 gnd.n3067 gnd.t10 6.69227
R12996 gnd.n2875 gnd.t348 6.69227
R12997 gnd.n2609 gnd.t124 6.69227
R12998 gnd.n5325 gnd.t135 6.69227
R12999 gnd.t141 gnd.n5450 6.69227
R13000 gnd.t273 gnd.n285 6.69227
R13001 gnd.n5748 gnd.n5747 6.5566
R13002 gnd.n5116 gnd.n5115 6.5566
R13003 gnd.n6485 gnd.n6481 6.5566
R13004 gnd.n5623 gnd.n5622 6.5566
R13005 gnd.t187 gnd.n1336 6.37362
R13006 gnd.n5245 gnd.n2212 6.37362
R13007 gnd.n2204 gnd.n2192 6.37362
R13008 gnd.n5314 gnd.t0 6.37362
R13009 gnd.n5379 gnd.n2122 6.37362
R13010 gnd.n5410 gnd.n5409 6.37362
R13011 gnd.n5460 gnd.t3 6.37362
R13012 gnd.n5540 gnd.n5539 6.37362
R13013 gnd.n5560 gnd.n5559 6.37362
R13014 gnd.n4857 gnd.n4846 6.20656
R13015 gnd.n7882 gnd.n7879 6.20656
R13016 gnd.n4180 gnd.n4175 6.20656
R13017 gnd.n6020 gnd.n6018 6.20656
R13018 gnd.t99 gnd.n3496 6.05496
R13019 gnd.n3497 gnd.t11 6.05496
R13020 gnd.t265 gnd.n2899 6.05496
R13021 gnd.t20 gnd.n3661 6.05496
R13022 gnd.t201 gnd.t296 6.05496
R13023 gnd.t71 gnd.n5263 6.05496
R13024 gnd.t322 gnd.t105 6.05496
R13025 gnd.t1 gnd.t106 6.05496
R13026 gnd.n5538 gnd.t263 6.05496
R13027 gnd.n7838 gnd.n126 6.05496
R13028 gnd.n4019 gnd.n3989 5.81868
R13029 gnd.n3987 gnd.n3957 5.81868
R13030 gnd.n3955 gnd.n3925 5.81868
R13031 gnd.n3924 gnd.n3894 5.81868
R13032 gnd.n3892 gnd.n3862 5.81868
R13033 gnd.n3860 gnd.n3830 5.81868
R13034 gnd.n3828 gnd.n3798 5.81868
R13035 gnd.n3797 gnd.n3767 5.81868
R13036 gnd.n5752 gnd.n1985 5.62001
R13037 gnd.n6547 gnd.n1301 5.62001
R13038 gnd.n6547 gnd.n1302 5.62001
R13039 gnd.n5618 gnd.n1985 5.62001
R13040 gnd.n3248 gnd.n3243 5.4308
R13041 gnd.n4064 gnd.n2740 5.4308
R13042 gnd.n3564 gnd.t21 5.41765
R13043 gnd.t8 gnd.n3587 5.41765
R13044 gnd.t151 gnd.n2829 5.41765
R13045 gnd.n5175 gnd.t187 5.09899
R13046 gnd.t214 gnd.n2208 5.09899
R13047 gnd.n5257 gnd.n2208 5.09899
R13048 gnd.n2125 gnd.n2114 5.09899
R13049 gnd.n5403 gnd.n5402 5.09899
R13050 gnd.n5474 gnd.n2023 5.09899
R13051 gnd.n4017 gnd.n4016 5.04292
R13052 gnd.n3985 gnd.n3984 5.04292
R13053 gnd.n3953 gnd.n3952 5.04292
R13054 gnd.n3922 gnd.n3921 5.04292
R13055 gnd.n3890 gnd.n3889 5.04292
R13056 gnd.n3858 gnd.n3857 5.04292
R13057 gnd.n3826 gnd.n3825 5.04292
R13058 gnd.n3795 gnd.n3794 5.04292
R13059 gnd.n2964 gnd.n2963 4.82753
R13060 gnd.n78 gnd.n77 4.82753
R13061 gnd.n3527 gnd.t12 4.78034
R13062 gnd.n2854 gnd.t316 4.78034
R13063 gnd.t318 gnd.n2253 4.78034
R13064 gnd.n5800 gnd.t341 4.78034
R13065 gnd.n2969 gnd.n2966 4.74817
R13066 gnd.n3019 gnd.n2905 4.74817
R13067 gnd.n3006 gnd.n2904 4.74817
R13068 gnd.n2903 gnd.n2902 4.74817
R13069 gnd.n3015 gnd.n2966 4.74817
R13070 gnd.n3016 gnd.n2905 4.74817
R13071 gnd.n3018 gnd.n2904 4.74817
R13072 gnd.n3005 gnd.n2903 4.74817
R13073 gnd.n7667 gnd.n7666 4.74817
R13074 gnd.n6287 gnd.n316 4.74817
R13075 gnd.n1535 gnd.n315 4.74817
R13076 gnd.n7646 gnd.n314 4.74817
R13077 gnd.n313 gnd.n310 4.74817
R13078 gnd.n7667 gnd.n317 4.74817
R13079 gnd.n7665 gnd.n316 4.74817
R13080 gnd.n6288 gnd.n315 4.74817
R13081 gnd.n1534 gnd.n314 4.74817
R13082 gnd.n7647 gnd.n313 4.74817
R13083 gnd.n4557 gnd.n4556 4.74817
R13084 gnd.n4558 gnd.n2546 4.74817
R13085 gnd.n4602 gnd.n4601 4.74817
R13086 gnd.n4612 gnd.n4611 4.74817
R13087 gnd.n4607 gnd.n4603 4.74817
R13088 gnd.n6256 gnd.n6255 4.74817
R13089 gnd.n6260 gnd.n1540 4.74817
R13090 gnd.n6282 gnd.n6262 4.74817
R13091 gnd.n6280 gnd.n6279 4.74817
R13092 gnd.n6275 gnd.n6265 4.74817
R13093 gnd.n6255 gnd.n6254 4.74817
R13094 gnd.n6257 gnd.n1540 4.74817
R13095 gnd.n6262 gnd.n6261 4.74817
R13096 gnd.n6281 gnd.n6280 4.74817
R13097 gnd.n6265 gnd.n6263 4.74817
R13098 gnd.n6669 gnd.n1090 4.74817
R13099 gnd.n6667 gnd.n1091 4.74817
R13100 gnd.n4595 gnd.n1096 4.74817
R13101 gnd.n4628 gnd.n1095 4.74817
R13102 gnd.n1097 gnd.n1094 4.74817
R13103 gnd.n1090 gnd.n1074 4.74817
R13104 gnd.n6668 gnd.n6667 4.74817
R13105 gnd.n4592 gnd.n1096 4.74817
R13106 gnd.n4594 gnd.n1095 4.74817
R13107 gnd.n4627 gnd.n1094 4.74817
R13108 gnd.n4560 gnd.n4557 4.74817
R13109 gnd.n4559 gnd.n4558 4.74817
R13110 gnd.n4601 gnd.n4600 4.74817
R13111 gnd.n4613 gnd.n4612 4.74817
R13112 gnd.n4610 gnd.n4603 4.74817
R13113 gnd.n2944 gnd.n2943 4.7074
R13114 gnd.n58 gnd.n57 4.7074
R13115 gnd.n2964 gnd.n2944 4.65959
R13116 gnd.n78 gnd.n58 4.65959
R13117 gnd.n1984 gnd.n1876 4.6132
R13118 gnd.n6548 gnd.n1300 4.6132
R13119 gnd.n6473 gnd.t154 4.46168
R13120 gnd.t154 gnd.n6472 4.46168
R13121 gnd.n5296 gnd.t287 4.46168
R13122 gnd.t308 gnd.n5507 4.46168
R13123 gnd.n5608 gnd.n5595 4.46111
R13124 gnd.n4002 gnd.n3998 4.38594
R13125 gnd.n3970 gnd.n3966 4.38594
R13126 gnd.n3938 gnd.n3934 4.38594
R13127 gnd.n3907 gnd.n3903 4.38594
R13128 gnd.n3875 gnd.n3871 4.38594
R13129 gnd.n3843 gnd.n3839 4.38594
R13130 gnd.n3811 gnd.n3807 4.38594
R13131 gnd.n3780 gnd.n3776 4.38594
R13132 gnd.n4013 gnd.n3991 4.26717
R13133 gnd.n3981 gnd.n3959 4.26717
R13134 gnd.n3949 gnd.n3927 4.26717
R13135 gnd.n3918 gnd.n3896 4.26717
R13136 gnd.n3886 gnd.n3864 4.26717
R13137 gnd.n3854 gnd.n3832 4.26717
R13138 gnd.n3822 gnd.n3800 4.26717
R13139 gnd.n3791 gnd.n3769 4.26717
R13140 gnd.n3471 gnd.t314 4.14303
R13141 gnd.n3701 gnd.t39 4.14303
R13142 gnd.t119 gnd.n1032 4.14303
R13143 gnd.t169 gnd.n1241 4.14303
R13144 gnd.n6062 gnd.t176 4.14303
R13145 gnd.t129 gnd.n266 4.14303
R13146 gnd.n4021 gnd.n4020 4.08274
R13147 gnd.n5747 gnd.n5746 4.05904
R13148 gnd.n5117 gnd.n5116 4.05904
R13149 gnd.n6488 gnd.n6481 4.05904
R13150 gnd.n5624 gnd.n5623 4.05904
R13151 gnd.n19 gnd.n9 3.99943
R13152 gnd.n6544 gnd.t304 3.82437
R13153 gnd.n5188 gnd.n5108 3.82437
R13154 gnd.n5256 gnd.t137 3.82437
R13155 gnd.n5273 gnd.n5272 3.82437
R13156 gnd.n5349 gnd.n2134 3.82437
R13157 gnd.n5338 gnd.n2098 3.82437
R13158 gnd.n5499 gnd.n2028 3.82437
R13159 gnd.t282 gnd.n5549 3.82437
R13160 gnd.n5574 gnd.n5573 3.82437
R13161 gnd.n5755 gnd.t101 3.82437
R13162 gnd.n4021 gnd.n3893 3.70378
R13163 gnd.n3544 gnd.n2965 3.65935
R13164 gnd.n19 gnd.n18 3.60163
R13165 gnd.n3740 gnd.n2789 3.50571
R13166 gnd.n4450 gnd.t230 3.50571
R13167 gnd.n4552 gnd.t18 3.50571
R13168 gnd.n4831 gnd.t169 3.50571
R13169 gnd.t176 gnd.n6061 3.50571
R13170 gnd.t60 gnd.n298 3.50571
R13171 gnd.n215 gnd.t157 3.50571
R13172 gnd.n4012 gnd.n3993 3.49141
R13173 gnd.n3980 gnd.n3961 3.49141
R13174 gnd.n3948 gnd.n3929 3.49141
R13175 gnd.n3917 gnd.n3898 3.49141
R13176 gnd.n3885 gnd.n3866 3.49141
R13177 gnd.n3853 gnd.n3834 3.49141
R13178 gnd.n3821 gnd.n3802 3.49141
R13179 gnd.n3790 gnd.n3771 3.49141
R13180 gnd.t313 gnd.n2789 3.18706
R13181 gnd.n5560 gnd.t180 3.18706
R13182 gnd.n3050 gnd.t314 2.8684
R13183 gnd.n4615 gnd.t29 2.8684
R13184 gnd.n5092 gnd.t304 2.8684
R13185 gnd.t139 gnd.n1531 2.8684
R13186 gnd.n2945 gnd.t91 2.82907
R13187 gnd.n2945 gnd.t302 2.82907
R13188 gnd.n2947 gnd.t32 2.82907
R13189 gnd.n2947 gnd.t290 2.82907
R13190 gnd.n2949 gnd.t75 2.82907
R13191 gnd.n2949 gnd.t88 2.82907
R13192 gnd.n2951 gnd.t53 2.82907
R13193 gnd.n2951 gnd.t347 2.82907
R13194 gnd.n2953 gnd.t278 2.82907
R13195 gnd.n2953 gnd.t98 2.82907
R13196 gnd.n2955 gnd.t271 2.82907
R13197 gnd.n2955 gnd.t41 2.82907
R13198 gnd.n2957 gnd.t317 2.82907
R13199 gnd.n2957 gnd.t295 2.82907
R13200 gnd.n2959 gnd.t294 2.82907
R13201 gnd.n2959 gnd.t279 2.82907
R13202 gnd.n2961 gnd.t34 2.82907
R13203 gnd.n2961 gnd.t301 2.82907
R13204 gnd.n2906 gnd.t107 2.82907
R13205 gnd.n2906 gnd.t84 2.82907
R13206 gnd.n2908 gnd.t300 2.82907
R13207 gnd.n2908 gnd.t325 2.82907
R13208 gnd.n2910 gnd.t127 2.82907
R13209 gnd.n2910 gnd.t17 2.82907
R13210 gnd.n2912 gnd.t109 2.82907
R13211 gnd.n2912 gnd.t122 2.82907
R13212 gnd.n2914 gnd.t343 2.82907
R13213 gnd.n2914 gnd.t80 2.82907
R13214 gnd.n2916 gnd.t57 2.82907
R13215 gnd.n2916 gnd.t138 2.82907
R13216 gnd.n2918 gnd.t125 2.82907
R13217 gnd.n2918 gnd.t82 2.82907
R13218 gnd.n2920 gnd.t144 2.82907
R13219 gnd.n2920 gnd.t120 2.82907
R13220 gnd.n2922 gnd.t123 2.82907
R13221 gnd.n2922 gnd.t298 2.82907
R13222 gnd.n2925 gnd.t28 2.82907
R13223 gnd.n2925 gnd.t108 2.82907
R13224 gnd.n2927 gnd.t42 2.82907
R13225 gnd.n2927 gnd.t148 2.82907
R13226 gnd.n2929 gnd.t95 2.82907
R13227 gnd.n2929 gnd.t126 2.82907
R13228 gnd.n2931 gnd.t267 2.82907
R13229 gnd.n2931 gnd.t331 2.82907
R13230 gnd.n2933 gnd.t345 2.82907
R13231 gnd.n2933 gnd.t30 2.82907
R13232 gnd.n2935 gnd.t19 2.82907
R13233 gnd.n2935 gnd.t55 2.82907
R13234 gnd.n2937 gnd.t336 2.82907
R13235 gnd.n2937 gnd.t103 2.82907
R13236 gnd.n2939 gnd.t299 2.82907
R13237 gnd.n2939 gnd.t328 2.82907
R13238 gnd.n2941 gnd.t112 2.82907
R13239 gnd.n2941 gnd.t67 2.82907
R13240 gnd.n75 gnd.t133 2.82907
R13241 gnd.n75 gnd.t280 2.82907
R13242 gnd.n73 gnd.t130 2.82907
R13243 gnd.n73 gnd.t15 2.82907
R13244 gnd.n71 gnd.t23 2.82907
R13245 gnd.n71 gnd.t293 2.82907
R13246 gnd.n69 gnd.t128 2.82907
R13247 gnd.n69 gnd.t76 2.82907
R13248 gnd.n67 gnd.t281 2.82907
R13249 gnd.n67 gnd.t64 2.82907
R13250 gnd.n65 gnd.t78 2.82907
R13251 gnd.n65 gnd.t90 2.82907
R13252 gnd.n63 gnd.t7 2.82907
R13253 gnd.n63 gnd.t87 2.82907
R13254 gnd.n61 gnd.t132 2.82907
R13255 gnd.n61 gnd.t303 2.82907
R13256 gnd.n59 gnd.t292 2.82907
R13257 gnd.n59 gnd.t338 2.82907
R13258 gnd.n36 gnd.t146 2.82907
R13259 gnd.n36 gnd.t270 2.82907
R13260 gnd.n34 gnd.t276 2.82907
R13261 gnd.n34 gnd.t324 2.82907
R13262 gnd.n32 gnd.t62 2.82907
R13263 gnd.n32 gnd.t274 2.82907
R13264 gnd.n30 gnd.t332 2.82907
R13265 gnd.n30 gnd.t111 2.82907
R13266 gnd.n28 gnd.t140 2.82907
R13267 gnd.n28 gnd.t79 2.82907
R13268 gnd.n26 gnd.t346 2.82907
R13269 gnd.n26 gnd.t326 2.82907
R13270 gnd.n24 gnd.t46 2.82907
R13271 gnd.n24 gnd.t269 2.82907
R13272 gnd.n22 gnd.t275 2.82907
R13273 gnd.n22 gnd.t333 2.82907
R13274 gnd.n20 gnd.t327 2.82907
R13275 gnd.n20 gnd.t268 2.82907
R13276 gnd.n55 gnd.t26 2.82907
R13277 gnd.n55 gnd.t118 2.82907
R13278 gnd.n53 gnd.t335 2.82907
R13279 gnd.n53 gnd.t56 2.82907
R13280 gnd.n51 gnd.t110 2.82907
R13281 gnd.n51 gnd.t330 2.82907
R13282 gnd.n49 gnd.t59 2.82907
R13283 gnd.n49 gnd.t61 2.82907
R13284 gnd.n47 gnd.t350 2.82907
R13285 gnd.n47 gnd.t94 2.82907
R13286 gnd.n45 gnd.t272 2.82907
R13287 gnd.n45 gnd.t344 2.82907
R13288 gnd.n43 gnd.t43 2.82907
R13289 gnd.n43 gnd.t116 2.82907
R13290 gnd.n41 gnd.t337 2.82907
R13291 gnd.n41 gnd.t48 2.82907
R13292 gnd.n39 gnd.t351 2.82907
R13293 gnd.n39 gnd.t5 2.82907
R13294 gnd.n4009 gnd.n4008 2.71565
R13295 gnd.n3977 gnd.n3976 2.71565
R13296 gnd.n3945 gnd.n3944 2.71565
R13297 gnd.n3914 gnd.n3913 2.71565
R13298 gnd.n3882 gnd.n3881 2.71565
R13299 gnd.n3850 gnd.n3849 2.71565
R13300 gnd.n3818 gnd.n3817 2.71565
R13301 gnd.n3787 gnd.n3786 2.71565
R13302 gnd.n5196 gnd.n5195 2.54975
R13303 gnd.n5288 gnd.n2182 2.54975
R13304 gnd.n5288 gnd.t104 2.54975
R13305 gnd.n5356 gnd.n2139 2.54975
R13306 gnd.n5427 gnd.n2094 2.54975
R13307 gnd.t73 gnd.n2038 2.54975
R13308 gnd.n5522 gnd.n2038 2.54975
R13309 gnd.n5566 gnd.n1997 2.54975
R13310 gnd.n3544 gnd.n2966 2.27742
R13311 gnd.n3544 gnd.n2905 2.27742
R13312 gnd.n3544 gnd.n2904 2.27742
R13313 gnd.n3544 gnd.n2903 2.27742
R13314 gnd.n7668 gnd.n7667 2.27742
R13315 gnd.n7668 gnd.n316 2.27742
R13316 gnd.n7668 gnd.n315 2.27742
R13317 gnd.n7668 gnd.n314 2.27742
R13318 gnd.n7668 gnd.n313 2.27742
R13319 gnd.n6255 gnd.n312 2.27742
R13320 gnd.n1540 gnd.n312 2.27742
R13321 gnd.n6262 gnd.n312 2.27742
R13322 gnd.n6280 gnd.n312 2.27742
R13323 gnd.n6265 gnd.n312 2.27742
R13324 gnd.n6666 gnd.n1090 2.27742
R13325 gnd.n6667 gnd.n6666 2.27742
R13326 gnd.n6666 gnd.n1096 2.27742
R13327 gnd.n6666 gnd.n1095 2.27742
R13328 gnd.n6666 gnd.n1094 2.27742
R13329 gnd.n4557 gnd.n1093 2.27742
R13330 gnd.n4558 gnd.n1093 2.27742
R13331 gnd.n4601 gnd.n1093 2.27742
R13332 gnd.n4612 gnd.n1093 2.27742
R13333 gnd.n4603 gnd.n1093 2.27742
R13334 gnd.n3398 gnd.t243 2.23109
R13335 gnd.n3021 gnd.t12 2.23109
R13336 gnd.t74 gnd.n1125 2.23109
R13337 gnd.n5349 gnd.t322 2.23109
R13338 gnd.n5338 gnd.t1 2.23109
R13339 gnd.t86 gnd.n6231 2.23109
R13340 gnd.n4005 gnd.n3995 1.93989
R13341 gnd.n3973 gnd.n3963 1.93989
R13342 gnd.n3941 gnd.n3931 1.93989
R13343 gnd.n3910 gnd.n3900 1.93989
R13344 gnd.n3878 gnd.n3868 1.93989
R13345 gnd.n3846 gnd.n3836 1.93989
R13346 gnd.n3814 gnd.n3804 1.93989
R13347 gnd.n3783 gnd.n3773 1.93989
R13348 gnd.n5188 gnd.t256 1.91244
R13349 gnd.t240 gnd.n1793 1.91244
R13350 gnd.t288 gnd.n3409 1.59378
R13351 gnd.n3588 gnd.t8 1.59378
R13352 gnd.n2838 gnd.t151 1.59378
R13353 gnd.n4500 gnd.t66 1.59378
R13354 gnd.t147 gnd.n1168 1.59378
R13355 gnd.n4737 gnd.t27 1.59378
R13356 gnd.t284 gnd.n2174 1.59378
R13357 gnd.n2044 gnd.t320 1.59378
R13358 gnd.n6125 gnd.t4 1.59378
R13359 gnd.t131 gnd.n1600 1.59378
R13360 gnd.t25 gnd.n244 1.59378
R13361 gnd.n6474 gnd.n1362 1.27512
R13362 gnd.t161 gnd.n1376 1.27512
R13363 gnd.n5264 gnd.t137 1.27512
R13364 gnd.n5297 gnd.n5296 1.27512
R13365 gnd.n5324 gnd.n2153 1.27512
R13366 gnd.n5451 gnd.n2079 1.27512
R13367 gnd.n5507 gnd.n2042 1.27512
R13368 gnd.n5551 gnd.t282 1.27512
R13369 gnd.n5582 gnd.t173 1.27512
R13370 gnd.n5580 gnd.t204 1.27512
R13371 gnd.n5686 gnd.n1992 1.27512
R13372 gnd.n3251 gnd.n3243 1.16414
R13373 gnd.n4067 gnd.n2740 1.16414
R13374 gnd.n4004 gnd.n3997 1.16414
R13375 gnd.n3972 gnd.n3965 1.16414
R13376 gnd.n3940 gnd.n3933 1.16414
R13377 gnd.n3909 gnd.n3902 1.16414
R13378 gnd.n3877 gnd.n3870 1.16414
R13379 gnd.n3845 gnd.n3838 1.16414
R13380 gnd.n3813 gnd.n3806 1.16414
R13381 gnd.n3782 gnd.n3775 1.16414
R13382 gnd.n1984 gnd.n1983 0.970197
R13383 gnd.n6548 gnd.n1296 0.970197
R13384 gnd.n3988 gnd.n3956 0.962709
R13385 gnd.n4020 gnd.n3988 0.962709
R13386 gnd.n3861 gnd.n3829 0.962709
R13387 gnd.n3893 gnd.n3861 0.962709
R13388 gnd.n3497 gnd.t99 0.956468
R13389 gnd.n3662 gnd.t20 0.956468
R13390 gnd.n6695 gnd.t124 0.956468
R13391 gnd.n4662 gnd.t16 0.956468
R13392 gnd.t44 gnd.n1211 0.956468
R13393 gnd.t101 gnd.t240 0.956468
R13394 gnd.n6095 gnd.t37 0.956468
R13395 gnd.n6220 gnd.t6 0.956468
R13396 gnd.n398 gnd.t273 0.956468
R13397 gnd.n2956 gnd.n2954 0.773756
R13398 gnd.n70 gnd.n68 0.773756
R13399 gnd.n2963 gnd.n2962 0.773756
R13400 gnd.n2962 gnd.n2960 0.773756
R13401 gnd.n2960 gnd.n2958 0.773756
R13402 gnd.n2958 gnd.n2956 0.773756
R13403 gnd.n2954 gnd.n2952 0.773756
R13404 gnd.n2952 gnd.n2950 0.773756
R13405 gnd.n2950 gnd.n2948 0.773756
R13406 gnd.n2948 gnd.n2946 0.773756
R13407 gnd.n62 gnd.n60 0.773756
R13408 gnd.n64 gnd.n62 0.773756
R13409 gnd.n66 gnd.n64 0.773756
R13410 gnd.n68 gnd.n66 0.773756
R13411 gnd.n72 gnd.n70 0.773756
R13412 gnd.n74 gnd.n72 0.773756
R13413 gnd.n76 gnd.n74 0.773756
R13414 gnd.n77 gnd.n76 0.773756
R13415 gnd gnd.n0 0.70738
R13416 gnd.n2 gnd.n1 0.672012
R13417 gnd.n3 gnd.n2 0.672012
R13418 gnd.n4 gnd.n3 0.672012
R13419 gnd.n5 gnd.n4 0.672012
R13420 gnd.n6 gnd.n5 0.672012
R13421 gnd.n7 gnd.n6 0.672012
R13422 gnd.n8 gnd.n7 0.672012
R13423 gnd.n9 gnd.n8 0.672012
R13424 gnd.n11 gnd.n10 0.672012
R13425 gnd.n12 gnd.n11 0.672012
R13426 gnd.n13 gnd.n12 0.672012
R13427 gnd.n14 gnd.n13 0.672012
R13428 gnd.n15 gnd.n14 0.672012
R13429 gnd.n16 gnd.n15 0.672012
R13430 gnd.n17 gnd.n16 0.672012
R13431 gnd.n18 gnd.n17 0.672012
R13432 gnd.n5272 gnd.t286 0.637812
R13433 gnd.n5499 gnd.t283 0.637812
R13434 gnd.n5591 gnd.t227 0.637812
R13435 gnd.n7972 gnd.n7971 0.637193
R13436 gnd.n2924 gnd.n2923 0.573776
R13437 gnd.n2923 gnd.n2921 0.573776
R13438 gnd.n2921 gnd.n2919 0.573776
R13439 gnd.n2919 gnd.n2917 0.573776
R13440 gnd.n2917 gnd.n2915 0.573776
R13441 gnd.n2915 gnd.n2913 0.573776
R13442 gnd.n2913 gnd.n2911 0.573776
R13443 gnd.n2911 gnd.n2909 0.573776
R13444 gnd.n2909 gnd.n2907 0.573776
R13445 gnd.n2943 gnd.n2942 0.573776
R13446 gnd.n2942 gnd.n2940 0.573776
R13447 gnd.n2940 gnd.n2938 0.573776
R13448 gnd.n2938 gnd.n2936 0.573776
R13449 gnd.n2936 gnd.n2934 0.573776
R13450 gnd.n2934 gnd.n2932 0.573776
R13451 gnd.n2932 gnd.n2930 0.573776
R13452 gnd.n2930 gnd.n2928 0.573776
R13453 gnd.n2928 gnd.n2926 0.573776
R13454 gnd.n23 gnd.n21 0.573776
R13455 gnd.n25 gnd.n23 0.573776
R13456 gnd.n27 gnd.n25 0.573776
R13457 gnd.n29 gnd.n27 0.573776
R13458 gnd.n31 gnd.n29 0.573776
R13459 gnd.n33 gnd.n31 0.573776
R13460 gnd.n35 gnd.n33 0.573776
R13461 gnd.n37 gnd.n35 0.573776
R13462 gnd.n38 gnd.n37 0.573776
R13463 gnd.n42 gnd.n40 0.573776
R13464 gnd.n44 gnd.n42 0.573776
R13465 gnd.n46 gnd.n44 0.573776
R13466 gnd.n48 gnd.n46 0.573776
R13467 gnd.n50 gnd.n48 0.573776
R13468 gnd.n52 gnd.n50 0.573776
R13469 gnd.n54 gnd.n52 0.573776
R13470 gnd.n56 gnd.n54 0.573776
R13471 gnd.n57 gnd.n56 0.573776
R13472 gnd.n7668 gnd.n312 0.548625
R13473 gnd.n6666 gnd.n1093 0.548625
R13474 gnd.n3724 gnd.n2744 0.486781
R13475 gnd.n6352 gnd.n6351 0.486781
R13476 gnd.n3300 gnd.n3299 0.48678
R13477 gnd.n2402 gnd.n2401 0.485256
R13478 gnd.n4041 gnd.n2698 0.480683
R13479 gnd.n3384 gnd.n3383 0.480683
R13480 gnd.n4402 gnd.n4397 0.477634
R13481 gnd.n4439 gnd.n4438 0.477634
R13482 gnd.n7834 gnd.n7833 0.477634
R13483 gnd.n7922 gnd.n7921 0.477634
R13484 gnd.n6880 gnd.n6879 0.468488
R13485 gnd.n7400 gnd.n7399 0.468488
R13486 gnd.n7613 gnd.n7612 0.468488
R13487 gnd.n2589 gnd.n1017 0.468488
R13488 gnd.n7914 gnd.n7913 0.465439
R13489 gnd.n7843 gnd.n7842 0.465439
R13490 gnd.n1944 gnd.n1941 0.465439
R13491 gnd.n6047 gnd.n6046 0.465439
R13492 gnd.n6581 gnd.n6580 0.465439
R13493 gnd.n4826 gnd.n4825 0.465439
R13494 gnd.n4292 gnd.n4291 0.465439
R13495 gnd.n4445 gnd.n2671 0.465439
R13496 gnd.n6023 gnd.n1469 0.451719
R13497 gnd.n4853 gnd.n2306 0.451719
R13498 gnd.n4860 gnd.n4846 0.388379
R13499 gnd.n4001 gnd.n4000 0.388379
R13500 gnd.n3969 gnd.n3968 0.388379
R13501 gnd.n3937 gnd.n3936 0.388379
R13502 gnd.n3906 gnd.n3905 0.388379
R13503 gnd.n3874 gnd.n3873 0.388379
R13504 gnd.n3842 gnd.n3841 0.388379
R13505 gnd.n3810 gnd.n3809 0.388379
R13506 gnd.n3779 gnd.n3778 0.388379
R13507 gnd.n7883 gnd.n7882 0.388379
R13508 gnd.n4238 gnd.n4180 0.388379
R13509 gnd.n6018 gnd.n6017 0.388379
R13510 gnd.n2340 gnd.n2339 0.378829
R13511 gnd.n6350 gnd.n6349 0.377553
R13512 gnd.n7972 gnd.n19 0.374463
R13513 gnd gnd.n7972 0.367492
R13514 gnd.n2800 gnd.t313 0.319156
R13515 gnd.n6671 gnd.t40 0.319156
R13516 gnd.n4638 gnd.t52 0.319156
R13517 gnd.t296 gnd.t161 0.319156
R13518 gnd.t339 gnd.t204 0.319156
R13519 gnd.n6190 gnd.t89 0.319156
R13520 gnd.n7638 gnd.t58 0.319156
R13521 gnd.n3218 gnd.n3196 0.311721
R13522 gnd.n4112 gnd.n4111 0.268793
R13523 gnd.n4871 gnd.n4870 0.247451
R13524 gnd.n6055 gnd.n1680 0.247451
R13525 gnd.n4111 gnd.n4110 0.241354
R13526 gnd.n1876 gnd.n1875 0.229039
R13527 gnd.n1879 gnd.n1876 0.229039
R13528 gnd.n1300 gnd.n1295 0.229039
R13529 gnd.n4777 gnd.n1300 0.229039
R13530 gnd.n2965 gnd.n0 0.210825
R13531 gnd.n3372 gnd.n3171 0.206293
R13532 gnd.n4018 gnd.n3990 0.155672
R13533 gnd.n4011 gnd.n3990 0.155672
R13534 gnd.n4011 gnd.n4010 0.155672
R13535 gnd.n4010 gnd.n3994 0.155672
R13536 gnd.n4003 gnd.n3994 0.155672
R13537 gnd.n4003 gnd.n4002 0.155672
R13538 gnd.n3986 gnd.n3958 0.155672
R13539 gnd.n3979 gnd.n3958 0.155672
R13540 gnd.n3979 gnd.n3978 0.155672
R13541 gnd.n3978 gnd.n3962 0.155672
R13542 gnd.n3971 gnd.n3962 0.155672
R13543 gnd.n3971 gnd.n3970 0.155672
R13544 gnd.n3954 gnd.n3926 0.155672
R13545 gnd.n3947 gnd.n3926 0.155672
R13546 gnd.n3947 gnd.n3946 0.155672
R13547 gnd.n3946 gnd.n3930 0.155672
R13548 gnd.n3939 gnd.n3930 0.155672
R13549 gnd.n3939 gnd.n3938 0.155672
R13550 gnd.n3923 gnd.n3895 0.155672
R13551 gnd.n3916 gnd.n3895 0.155672
R13552 gnd.n3916 gnd.n3915 0.155672
R13553 gnd.n3915 gnd.n3899 0.155672
R13554 gnd.n3908 gnd.n3899 0.155672
R13555 gnd.n3908 gnd.n3907 0.155672
R13556 gnd.n3891 gnd.n3863 0.155672
R13557 gnd.n3884 gnd.n3863 0.155672
R13558 gnd.n3884 gnd.n3883 0.155672
R13559 gnd.n3883 gnd.n3867 0.155672
R13560 gnd.n3876 gnd.n3867 0.155672
R13561 gnd.n3876 gnd.n3875 0.155672
R13562 gnd.n3859 gnd.n3831 0.155672
R13563 gnd.n3852 gnd.n3831 0.155672
R13564 gnd.n3852 gnd.n3851 0.155672
R13565 gnd.n3851 gnd.n3835 0.155672
R13566 gnd.n3844 gnd.n3835 0.155672
R13567 gnd.n3844 gnd.n3843 0.155672
R13568 gnd.n3827 gnd.n3799 0.155672
R13569 gnd.n3820 gnd.n3799 0.155672
R13570 gnd.n3820 gnd.n3819 0.155672
R13571 gnd.n3819 gnd.n3803 0.155672
R13572 gnd.n3812 gnd.n3803 0.155672
R13573 gnd.n3812 gnd.n3811 0.155672
R13574 gnd.n3796 gnd.n3768 0.155672
R13575 gnd.n3789 gnd.n3768 0.155672
R13576 gnd.n3789 gnd.n3788 0.155672
R13577 gnd.n3788 gnd.n3772 0.155672
R13578 gnd.n3781 gnd.n3772 0.155672
R13579 gnd.n3781 gnd.n3780 0.155672
R13580 gnd.n4143 gnd.n2698 0.152939
R13581 gnd.n4143 gnd.n4142 0.152939
R13582 gnd.n4142 gnd.n4141 0.152939
R13583 gnd.n4141 gnd.n2700 0.152939
R13584 gnd.n2701 gnd.n2700 0.152939
R13585 gnd.n2702 gnd.n2701 0.152939
R13586 gnd.n2703 gnd.n2702 0.152939
R13587 gnd.n2704 gnd.n2703 0.152939
R13588 gnd.n2705 gnd.n2704 0.152939
R13589 gnd.n2706 gnd.n2705 0.152939
R13590 gnd.n2707 gnd.n2706 0.152939
R13591 gnd.n2708 gnd.n2707 0.152939
R13592 gnd.n2709 gnd.n2708 0.152939
R13593 gnd.n2710 gnd.n2709 0.152939
R13594 gnd.n4113 gnd.n2710 0.152939
R13595 gnd.n4113 gnd.n4112 0.152939
R13596 gnd.n3385 gnd.n3384 0.152939
R13597 gnd.n3385 gnd.n3089 0.152939
R13598 gnd.n3413 gnd.n3089 0.152939
R13599 gnd.n3414 gnd.n3413 0.152939
R13600 gnd.n3415 gnd.n3414 0.152939
R13601 gnd.n3416 gnd.n3415 0.152939
R13602 gnd.n3416 gnd.n3061 0.152939
R13603 gnd.n3443 gnd.n3061 0.152939
R13604 gnd.n3444 gnd.n3443 0.152939
R13605 gnd.n3445 gnd.n3444 0.152939
R13606 gnd.n3445 gnd.n3039 0.152939
R13607 gnd.n3474 gnd.n3039 0.152939
R13608 gnd.n3475 gnd.n3474 0.152939
R13609 gnd.n3476 gnd.n3475 0.152939
R13610 gnd.n3477 gnd.n3476 0.152939
R13611 gnd.n3479 gnd.n3477 0.152939
R13612 gnd.n3479 gnd.n3478 0.152939
R13613 gnd.n3478 gnd.n2988 0.152939
R13614 gnd.n2989 gnd.n2988 0.152939
R13615 gnd.n2990 gnd.n2989 0.152939
R13616 gnd.n3009 gnd.n2990 0.152939
R13617 gnd.n3010 gnd.n3009 0.152939
R13618 gnd.n3010 gnd.n2896 0.152939
R13619 gnd.n3569 gnd.n2896 0.152939
R13620 gnd.n3570 gnd.n3569 0.152939
R13621 gnd.n3571 gnd.n3570 0.152939
R13622 gnd.n3572 gnd.n3571 0.152939
R13623 gnd.n3572 gnd.n2869 0.152939
R13624 gnd.n3609 gnd.n2869 0.152939
R13625 gnd.n3610 gnd.n3609 0.152939
R13626 gnd.n3611 gnd.n3610 0.152939
R13627 gnd.n3612 gnd.n3611 0.152939
R13628 gnd.n3612 gnd.n2842 0.152939
R13629 gnd.n3654 gnd.n2842 0.152939
R13630 gnd.n3655 gnd.n3654 0.152939
R13631 gnd.n3656 gnd.n3655 0.152939
R13632 gnd.n3657 gnd.n3656 0.152939
R13633 gnd.n3657 gnd.n2814 0.152939
R13634 gnd.n3694 gnd.n2814 0.152939
R13635 gnd.n3695 gnd.n3694 0.152939
R13636 gnd.n3696 gnd.n3695 0.152939
R13637 gnd.n3697 gnd.n3696 0.152939
R13638 gnd.n3697 gnd.n2786 0.152939
R13639 gnd.n3743 gnd.n2786 0.152939
R13640 gnd.n3744 gnd.n3743 0.152939
R13641 gnd.n3745 gnd.n3744 0.152939
R13642 gnd.n3746 gnd.n3745 0.152939
R13643 gnd.n3746 gnd.n2759 0.152939
R13644 gnd.n4037 gnd.n2759 0.152939
R13645 gnd.n4038 gnd.n4037 0.152939
R13646 gnd.n4039 gnd.n4038 0.152939
R13647 gnd.n4040 gnd.n4039 0.152939
R13648 gnd.n4041 gnd.n4040 0.152939
R13649 gnd.n3383 gnd.n3113 0.152939
R13650 gnd.n3134 gnd.n3113 0.152939
R13651 gnd.n3135 gnd.n3134 0.152939
R13652 gnd.n3141 gnd.n3135 0.152939
R13653 gnd.n3142 gnd.n3141 0.152939
R13654 gnd.n3143 gnd.n3142 0.152939
R13655 gnd.n3143 gnd.n3132 0.152939
R13656 gnd.n3151 gnd.n3132 0.152939
R13657 gnd.n3152 gnd.n3151 0.152939
R13658 gnd.n3153 gnd.n3152 0.152939
R13659 gnd.n3153 gnd.n3130 0.152939
R13660 gnd.n3161 gnd.n3130 0.152939
R13661 gnd.n3162 gnd.n3161 0.152939
R13662 gnd.n3163 gnd.n3162 0.152939
R13663 gnd.n3163 gnd.n3128 0.152939
R13664 gnd.n3171 gnd.n3128 0.152939
R13665 gnd.n4110 gnd.n2715 0.152939
R13666 gnd.n2717 gnd.n2715 0.152939
R13667 gnd.n2718 gnd.n2717 0.152939
R13668 gnd.n2719 gnd.n2718 0.152939
R13669 gnd.n2720 gnd.n2719 0.152939
R13670 gnd.n2721 gnd.n2720 0.152939
R13671 gnd.n2722 gnd.n2721 0.152939
R13672 gnd.n2723 gnd.n2722 0.152939
R13673 gnd.n2724 gnd.n2723 0.152939
R13674 gnd.n2725 gnd.n2724 0.152939
R13675 gnd.n2726 gnd.n2725 0.152939
R13676 gnd.n2727 gnd.n2726 0.152939
R13677 gnd.n2728 gnd.n2727 0.152939
R13678 gnd.n2729 gnd.n2728 0.152939
R13679 gnd.n2730 gnd.n2729 0.152939
R13680 gnd.n2731 gnd.n2730 0.152939
R13681 gnd.n2732 gnd.n2731 0.152939
R13682 gnd.n2733 gnd.n2732 0.152939
R13683 gnd.n2734 gnd.n2733 0.152939
R13684 gnd.n2735 gnd.n2734 0.152939
R13685 gnd.n2736 gnd.n2735 0.152939
R13686 gnd.n2737 gnd.n2736 0.152939
R13687 gnd.n2741 gnd.n2737 0.152939
R13688 gnd.n2742 gnd.n2741 0.152939
R13689 gnd.n2743 gnd.n2742 0.152939
R13690 gnd.n2744 gnd.n2743 0.152939
R13691 gnd.n3546 gnd.n3545 0.152939
R13692 gnd.n3547 gnd.n3546 0.152939
R13693 gnd.n3548 gnd.n3547 0.152939
R13694 gnd.n3549 gnd.n3548 0.152939
R13695 gnd.n3550 gnd.n3549 0.152939
R13696 gnd.n3551 gnd.n3550 0.152939
R13697 gnd.n3551 gnd.n2850 0.152939
R13698 gnd.n3630 gnd.n2850 0.152939
R13699 gnd.n3631 gnd.n3630 0.152939
R13700 gnd.n3632 gnd.n3631 0.152939
R13701 gnd.n3633 gnd.n3632 0.152939
R13702 gnd.n3634 gnd.n3633 0.152939
R13703 gnd.n3635 gnd.n3634 0.152939
R13704 gnd.n3636 gnd.n3635 0.152939
R13705 gnd.n3637 gnd.n3636 0.152939
R13706 gnd.n3638 gnd.n3637 0.152939
R13707 gnd.n3638 gnd.n2794 0.152939
R13708 gnd.n3715 gnd.n2794 0.152939
R13709 gnd.n3716 gnd.n3715 0.152939
R13710 gnd.n3717 gnd.n3716 0.152939
R13711 gnd.n3718 gnd.n3717 0.152939
R13712 gnd.n3719 gnd.n3718 0.152939
R13713 gnd.n3720 gnd.n3719 0.152939
R13714 gnd.n3721 gnd.n3720 0.152939
R13715 gnd.n3722 gnd.n3721 0.152939
R13716 gnd.n3723 gnd.n3722 0.152939
R13717 gnd.n3725 gnd.n3723 0.152939
R13718 gnd.n3725 gnd.n3724 0.152939
R13719 gnd.n3301 gnd.n3300 0.152939
R13720 gnd.n3301 gnd.n3191 0.152939
R13721 gnd.n3316 gnd.n3191 0.152939
R13722 gnd.n3317 gnd.n3316 0.152939
R13723 gnd.n3318 gnd.n3317 0.152939
R13724 gnd.n3318 gnd.n3179 0.152939
R13725 gnd.n3332 gnd.n3179 0.152939
R13726 gnd.n3333 gnd.n3332 0.152939
R13727 gnd.n3334 gnd.n3333 0.152939
R13728 gnd.n3335 gnd.n3334 0.152939
R13729 gnd.n3336 gnd.n3335 0.152939
R13730 gnd.n3337 gnd.n3336 0.152939
R13731 gnd.n3338 gnd.n3337 0.152939
R13732 gnd.n3339 gnd.n3338 0.152939
R13733 gnd.n3340 gnd.n3339 0.152939
R13734 gnd.n3341 gnd.n3340 0.152939
R13735 gnd.n3342 gnd.n3341 0.152939
R13736 gnd.n3343 gnd.n3342 0.152939
R13737 gnd.n3344 gnd.n3343 0.152939
R13738 gnd.n3345 gnd.n3344 0.152939
R13739 gnd.n3346 gnd.n3345 0.152939
R13740 gnd.n3346 gnd.n3045 0.152939
R13741 gnd.n3463 gnd.n3045 0.152939
R13742 gnd.n3464 gnd.n3463 0.152939
R13743 gnd.n3465 gnd.n3464 0.152939
R13744 gnd.n3466 gnd.n3465 0.152939
R13745 gnd.n3466 gnd.n2967 0.152939
R13746 gnd.n3543 gnd.n2967 0.152939
R13747 gnd.n3219 gnd.n3218 0.152939
R13748 gnd.n3220 gnd.n3219 0.152939
R13749 gnd.n3221 gnd.n3220 0.152939
R13750 gnd.n3222 gnd.n3221 0.152939
R13751 gnd.n3223 gnd.n3222 0.152939
R13752 gnd.n3224 gnd.n3223 0.152939
R13753 gnd.n3225 gnd.n3224 0.152939
R13754 gnd.n3226 gnd.n3225 0.152939
R13755 gnd.n3227 gnd.n3226 0.152939
R13756 gnd.n3228 gnd.n3227 0.152939
R13757 gnd.n3229 gnd.n3228 0.152939
R13758 gnd.n3230 gnd.n3229 0.152939
R13759 gnd.n3231 gnd.n3230 0.152939
R13760 gnd.n3232 gnd.n3231 0.152939
R13761 gnd.n3233 gnd.n3232 0.152939
R13762 gnd.n3234 gnd.n3233 0.152939
R13763 gnd.n3235 gnd.n3234 0.152939
R13764 gnd.n3236 gnd.n3235 0.152939
R13765 gnd.n3237 gnd.n3236 0.152939
R13766 gnd.n3238 gnd.n3237 0.152939
R13767 gnd.n3239 gnd.n3238 0.152939
R13768 gnd.n3240 gnd.n3239 0.152939
R13769 gnd.n3244 gnd.n3240 0.152939
R13770 gnd.n3245 gnd.n3244 0.152939
R13771 gnd.n3245 gnd.n3202 0.152939
R13772 gnd.n3299 gnd.n3202 0.152939
R13773 gnd.n6881 gnd.n6880 0.152939
R13774 gnd.n6881 gnd.n844 0.152939
R13775 gnd.n6889 gnd.n844 0.152939
R13776 gnd.n6890 gnd.n6889 0.152939
R13777 gnd.n6891 gnd.n6890 0.152939
R13778 gnd.n6891 gnd.n838 0.152939
R13779 gnd.n6899 gnd.n838 0.152939
R13780 gnd.n6900 gnd.n6899 0.152939
R13781 gnd.n6901 gnd.n6900 0.152939
R13782 gnd.n6901 gnd.n832 0.152939
R13783 gnd.n6909 gnd.n832 0.152939
R13784 gnd.n6910 gnd.n6909 0.152939
R13785 gnd.n6911 gnd.n6910 0.152939
R13786 gnd.n6911 gnd.n826 0.152939
R13787 gnd.n6919 gnd.n826 0.152939
R13788 gnd.n6920 gnd.n6919 0.152939
R13789 gnd.n6921 gnd.n6920 0.152939
R13790 gnd.n6921 gnd.n820 0.152939
R13791 gnd.n6929 gnd.n820 0.152939
R13792 gnd.n6930 gnd.n6929 0.152939
R13793 gnd.n6931 gnd.n6930 0.152939
R13794 gnd.n6931 gnd.n814 0.152939
R13795 gnd.n6939 gnd.n814 0.152939
R13796 gnd.n6940 gnd.n6939 0.152939
R13797 gnd.n6941 gnd.n6940 0.152939
R13798 gnd.n6941 gnd.n808 0.152939
R13799 gnd.n6949 gnd.n808 0.152939
R13800 gnd.n6950 gnd.n6949 0.152939
R13801 gnd.n6951 gnd.n6950 0.152939
R13802 gnd.n6951 gnd.n802 0.152939
R13803 gnd.n6959 gnd.n802 0.152939
R13804 gnd.n6960 gnd.n6959 0.152939
R13805 gnd.n6961 gnd.n6960 0.152939
R13806 gnd.n6961 gnd.n796 0.152939
R13807 gnd.n6969 gnd.n796 0.152939
R13808 gnd.n6970 gnd.n6969 0.152939
R13809 gnd.n6971 gnd.n6970 0.152939
R13810 gnd.n6971 gnd.n790 0.152939
R13811 gnd.n6979 gnd.n790 0.152939
R13812 gnd.n6980 gnd.n6979 0.152939
R13813 gnd.n6981 gnd.n6980 0.152939
R13814 gnd.n6981 gnd.n784 0.152939
R13815 gnd.n6989 gnd.n784 0.152939
R13816 gnd.n6990 gnd.n6989 0.152939
R13817 gnd.n6991 gnd.n6990 0.152939
R13818 gnd.n6991 gnd.n778 0.152939
R13819 gnd.n6999 gnd.n778 0.152939
R13820 gnd.n7000 gnd.n6999 0.152939
R13821 gnd.n7001 gnd.n7000 0.152939
R13822 gnd.n7001 gnd.n772 0.152939
R13823 gnd.n7009 gnd.n772 0.152939
R13824 gnd.n7010 gnd.n7009 0.152939
R13825 gnd.n7011 gnd.n7010 0.152939
R13826 gnd.n7011 gnd.n766 0.152939
R13827 gnd.n7019 gnd.n766 0.152939
R13828 gnd.n7020 gnd.n7019 0.152939
R13829 gnd.n7021 gnd.n7020 0.152939
R13830 gnd.n7021 gnd.n760 0.152939
R13831 gnd.n7029 gnd.n760 0.152939
R13832 gnd.n7030 gnd.n7029 0.152939
R13833 gnd.n7031 gnd.n7030 0.152939
R13834 gnd.n7031 gnd.n754 0.152939
R13835 gnd.n7039 gnd.n754 0.152939
R13836 gnd.n7040 gnd.n7039 0.152939
R13837 gnd.n7041 gnd.n7040 0.152939
R13838 gnd.n7041 gnd.n748 0.152939
R13839 gnd.n7049 gnd.n748 0.152939
R13840 gnd.n7050 gnd.n7049 0.152939
R13841 gnd.n7051 gnd.n7050 0.152939
R13842 gnd.n7051 gnd.n742 0.152939
R13843 gnd.n7059 gnd.n742 0.152939
R13844 gnd.n7060 gnd.n7059 0.152939
R13845 gnd.n7061 gnd.n7060 0.152939
R13846 gnd.n7061 gnd.n736 0.152939
R13847 gnd.n7069 gnd.n736 0.152939
R13848 gnd.n7070 gnd.n7069 0.152939
R13849 gnd.n7071 gnd.n7070 0.152939
R13850 gnd.n7071 gnd.n730 0.152939
R13851 gnd.n7079 gnd.n730 0.152939
R13852 gnd.n7080 gnd.n7079 0.152939
R13853 gnd.n7081 gnd.n7080 0.152939
R13854 gnd.n7081 gnd.n724 0.152939
R13855 gnd.n7089 gnd.n724 0.152939
R13856 gnd.n7090 gnd.n7089 0.152939
R13857 gnd.n7091 gnd.n7090 0.152939
R13858 gnd.n7091 gnd.n718 0.152939
R13859 gnd.n7099 gnd.n718 0.152939
R13860 gnd.n7100 gnd.n7099 0.152939
R13861 gnd.n7101 gnd.n7100 0.152939
R13862 gnd.n7101 gnd.n712 0.152939
R13863 gnd.n7109 gnd.n712 0.152939
R13864 gnd.n7110 gnd.n7109 0.152939
R13865 gnd.n7111 gnd.n7110 0.152939
R13866 gnd.n7111 gnd.n706 0.152939
R13867 gnd.n7119 gnd.n706 0.152939
R13868 gnd.n7120 gnd.n7119 0.152939
R13869 gnd.n7121 gnd.n7120 0.152939
R13870 gnd.n7121 gnd.n700 0.152939
R13871 gnd.n7129 gnd.n700 0.152939
R13872 gnd.n7130 gnd.n7129 0.152939
R13873 gnd.n7131 gnd.n7130 0.152939
R13874 gnd.n7131 gnd.n694 0.152939
R13875 gnd.n7139 gnd.n694 0.152939
R13876 gnd.n7140 gnd.n7139 0.152939
R13877 gnd.n7141 gnd.n7140 0.152939
R13878 gnd.n7141 gnd.n688 0.152939
R13879 gnd.n7149 gnd.n688 0.152939
R13880 gnd.n7150 gnd.n7149 0.152939
R13881 gnd.n7151 gnd.n7150 0.152939
R13882 gnd.n7151 gnd.n682 0.152939
R13883 gnd.n7159 gnd.n682 0.152939
R13884 gnd.n7160 gnd.n7159 0.152939
R13885 gnd.n7161 gnd.n7160 0.152939
R13886 gnd.n7161 gnd.n676 0.152939
R13887 gnd.n7169 gnd.n676 0.152939
R13888 gnd.n7170 gnd.n7169 0.152939
R13889 gnd.n7171 gnd.n7170 0.152939
R13890 gnd.n7171 gnd.n670 0.152939
R13891 gnd.n7179 gnd.n670 0.152939
R13892 gnd.n7180 gnd.n7179 0.152939
R13893 gnd.n7181 gnd.n7180 0.152939
R13894 gnd.n7181 gnd.n664 0.152939
R13895 gnd.n7189 gnd.n664 0.152939
R13896 gnd.n7190 gnd.n7189 0.152939
R13897 gnd.n7191 gnd.n7190 0.152939
R13898 gnd.n7191 gnd.n658 0.152939
R13899 gnd.n7199 gnd.n658 0.152939
R13900 gnd.n7200 gnd.n7199 0.152939
R13901 gnd.n7201 gnd.n7200 0.152939
R13902 gnd.n7201 gnd.n652 0.152939
R13903 gnd.n7209 gnd.n652 0.152939
R13904 gnd.n7210 gnd.n7209 0.152939
R13905 gnd.n7211 gnd.n7210 0.152939
R13906 gnd.n7211 gnd.n646 0.152939
R13907 gnd.n7219 gnd.n646 0.152939
R13908 gnd.n7220 gnd.n7219 0.152939
R13909 gnd.n7221 gnd.n7220 0.152939
R13910 gnd.n7221 gnd.n640 0.152939
R13911 gnd.n7229 gnd.n640 0.152939
R13912 gnd.n7230 gnd.n7229 0.152939
R13913 gnd.n7231 gnd.n7230 0.152939
R13914 gnd.n7231 gnd.n634 0.152939
R13915 gnd.n7239 gnd.n634 0.152939
R13916 gnd.n7240 gnd.n7239 0.152939
R13917 gnd.n7241 gnd.n7240 0.152939
R13918 gnd.n7241 gnd.n628 0.152939
R13919 gnd.n7249 gnd.n628 0.152939
R13920 gnd.n7250 gnd.n7249 0.152939
R13921 gnd.n7251 gnd.n7250 0.152939
R13922 gnd.n7251 gnd.n622 0.152939
R13923 gnd.n7259 gnd.n622 0.152939
R13924 gnd.n7260 gnd.n7259 0.152939
R13925 gnd.n7261 gnd.n7260 0.152939
R13926 gnd.n7261 gnd.n616 0.152939
R13927 gnd.n7269 gnd.n616 0.152939
R13928 gnd.n7270 gnd.n7269 0.152939
R13929 gnd.n7271 gnd.n7270 0.152939
R13930 gnd.n7271 gnd.n610 0.152939
R13931 gnd.n7279 gnd.n610 0.152939
R13932 gnd.n7280 gnd.n7279 0.152939
R13933 gnd.n7281 gnd.n7280 0.152939
R13934 gnd.n7281 gnd.n604 0.152939
R13935 gnd.n7289 gnd.n604 0.152939
R13936 gnd.n7290 gnd.n7289 0.152939
R13937 gnd.n7291 gnd.n7290 0.152939
R13938 gnd.n7291 gnd.n598 0.152939
R13939 gnd.n7299 gnd.n598 0.152939
R13940 gnd.n7300 gnd.n7299 0.152939
R13941 gnd.n7301 gnd.n7300 0.152939
R13942 gnd.n7301 gnd.n592 0.152939
R13943 gnd.n7309 gnd.n592 0.152939
R13944 gnd.n7310 gnd.n7309 0.152939
R13945 gnd.n7311 gnd.n7310 0.152939
R13946 gnd.n7311 gnd.n586 0.152939
R13947 gnd.n7319 gnd.n586 0.152939
R13948 gnd.n7320 gnd.n7319 0.152939
R13949 gnd.n7321 gnd.n7320 0.152939
R13950 gnd.n7321 gnd.n580 0.152939
R13951 gnd.n7329 gnd.n580 0.152939
R13952 gnd.n7330 gnd.n7329 0.152939
R13953 gnd.n7331 gnd.n7330 0.152939
R13954 gnd.n7331 gnd.n574 0.152939
R13955 gnd.n7339 gnd.n574 0.152939
R13956 gnd.n7340 gnd.n7339 0.152939
R13957 gnd.n7341 gnd.n7340 0.152939
R13958 gnd.n7341 gnd.n568 0.152939
R13959 gnd.n7349 gnd.n568 0.152939
R13960 gnd.n7350 gnd.n7349 0.152939
R13961 gnd.n7351 gnd.n7350 0.152939
R13962 gnd.n7351 gnd.n562 0.152939
R13963 gnd.n7359 gnd.n562 0.152939
R13964 gnd.n7360 gnd.n7359 0.152939
R13965 gnd.n7361 gnd.n7360 0.152939
R13966 gnd.n7361 gnd.n556 0.152939
R13967 gnd.n7369 gnd.n556 0.152939
R13968 gnd.n7370 gnd.n7369 0.152939
R13969 gnd.n7371 gnd.n7370 0.152939
R13970 gnd.n7371 gnd.n550 0.152939
R13971 gnd.n7379 gnd.n550 0.152939
R13972 gnd.n7380 gnd.n7379 0.152939
R13973 gnd.n7381 gnd.n7380 0.152939
R13974 gnd.n7381 gnd.n544 0.152939
R13975 gnd.n7389 gnd.n544 0.152939
R13976 gnd.n7390 gnd.n7389 0.152939
R13977 gnd.n7391 gnd.n7390 0.152939
R13978 gnd.n7391 gnd.n538 0.152939
R13979 gnd.n7399 gnd.n538 0.152939
R13980 gnd.n7401 gnd.n7400 0.152939
R13981 gnd.n7401 gnd.n532 0.152939
R13982 gnd.n7409 gnd.n532 0.152939
R13983 gnd.n7410 gnd.n7409 0.152939
R13984 gnd.n7411 gnd.n7410 0.152939
R13985 gnd.n7411 gnd.n526 0.152939
R13986 gnd.n7419 gnd.n526 0.152939
R13987 gnd.n7420 gnd.n7419 0.152939
R13988 gnd.n7421 gnd.n7420 0.152939
R13989 gnd.n7421 gnd.n520 0.152939
R13990 gnd.n7429 gnd.n520 0.152939
R13991 gnd.n7430 gnd.n7429 0.152939
R13992 gnd.n7431 gnd.n7430 0.152939
R13993 gnd.n7431 gnd.n514 0.152939
R13994 gnd.n7439 gnd.n514 0.152939
R13995 gnd.n7440 gnd.n7439 0.152939
R13996 gnd.n7441 gnd.n7440 0.152939
R13997 gnd.n7441 gnd.n508 0.152939
R13998 gnd.n7449 gnd.n508 0.152939
R13999 gnd.n7450 gnd.n7449 0.152939
R14000 gnd.n7451 gnd.n7450 0.152939
R14001 gnd.n7451 gnd.n502 0.152939
R14002 gnd.n7459 gnd.n502 0.152939
R14003 gnd.n7460 gnd.n7459 0.152939
R14004 gnd.n7461 gnd.n7460 0.152939
R14005 gnd.n7461 gnd.n496 0.152939
R14006 gnd.n7469 gnd.n496 0.152939
R14007 gnd.n7470 gnd.n7469 0.152939
R14008 gnd.n7471 gnd.n7470 0.152939
R14009 gnd.n7471 gnd.n490 0.152939
R14010 gnd.n7479 gnd.n490 0.152939
R14011 gnd.n7480 gnd.n7479 0.152939
R14012 gnd.n7481 gnd.n7480 0.152939
R14013 gnd.n7481 gnd.n484 0.152939
R14014 gnd.n7489 gnd.n484 0.152939
R14015 gnd.n7490 gnd.n7489 0.152939
R14016 gnd.n7491 gnd.n7490 0.152939
R14017 gnd.n7491 gnd.n478 0.152939
R14018 gnd.n7499 gnd.n478 0.152939
R14019 gnd.n7500 gnd.n7499 0.152939
R14020 gnd.n7501 gnd.n7500 0.152939
R14021 gnd.n7501 gnd.n472 0.152939
R14022 gnd.n7509 gnd.n472 0.152939
R14023 gnd.n7510 gnd.n7509 0.152939
R14024 gnd.n7511 gnd.n7510 0.152939
R14025 gnd.n7511 gnd.n466 0.152939
R14026 gnd.n7519 gnd.n466 0.152939
R14027 gnd.n7520 gnd.n7519 0.152939
R14028 gnd.n7521 gnd.n7520 0.152939
R14029 gnd.n7521 gnd.n460 0.152939
R14030 gnd.n7529 gnd.n460 0.152939
R14031 gnd.n7530 gnd.n7529 0.152939
R14032 gnd.n7531 gnd.n7530 0.152939
R14033 gnd.n7531 gnd.n454 0.152939
R14034 gnd.n7539 gnd.n454 0.152939
R14035 gnd.n7540 gnd.n7539 0.152939
R14036 gnd.n7541 gnd.n7540 0.152939
R14037 gnd.n7541 gnd.n448 0.152939
R14038 gnd.n7549 gnd.n448 0.152939
R14039 gnd.n7550 gnd.n7549 0.152939
R14040 gnd.n7551 gnd.n7550 0.152939
R14041 gnd.n7551 gnd.n442 0.152939
R14042 gnd.n7559 gnd.n442 0.152939
R14043 gnd.n7560 gnd.n7559 0.152939
R14044 gnd.n7561 gnd.n7560 0.152939
R14045 gnd.n7561 gnd.n436 0.152939
R14046 gnd.n7569 gnd.n436 0.152939
R14047 gnd.n7570 gnd.n7569 0.152939
R14048 gnd.n7571 gnd.n7570 0.152939
R14049 gnd.n7571 gnd.n430 0.152939
R14050 gnd.n7579 gnd.n430 0.152939
R14051 gnd.n7580 gnd.n7579 0.152939
R14052 gnd.n7581 gnd.n7580 0.152939
R14053 gnd.n7581 gnd.n424 0.152939
R14054 gnd.n7589 gnd.n424 0.152939
R14055 gnd.n7590 gnd.n7589 0.152939
R14056 gnd.n7591 gnd.n7590 0.152939
R14057 gnd.n7591 gnd.n418 0.152939
R14058 gnd.n7599 gnd.n418 0.152939
R14059 gnd.n7600 gnd.n7599 0.152939
R14060 gnd.n7601 gnd.n7600 0.152939
R14061 gnd.n7602 gnd.n7601 0.152939
R14062 gnd.n7602 gnd.n412 0.152939
R14063 gnd.n7612 gnd.n412 0.152939
R14064 gnd.n6267 gnd.n6266 0.152939
R14065 gnd.n6269 gnd.n6267 0.152939
R14066 gnd.n6269 gnd.n6268 0.152939
R14067 gnd.n6268 gnd.n405 0.152939
R14068 gnd.n406 gnd.n405 0.152939
R14069 gnd.n407 gnd.n406 0.152939
R14070 gnd.n410 gnd.n407 0.152939
R14071 gnd.n411 gnd.n410 0.152939
R14072 gnd.n7613 gnd.n411 0.152939
R14073 gnd.n7668 gnd.n295 0.152939
R14074 gnd.n7682 gnd.n295 0.152939
R14075 gnd.n7683 gnd.n7682 0.152939
R14076 gnd.n7684 gnd.n7683 0.152939
R14077 gnd.n7684 gnd.n280 0.152939
R14078 gnd.n7698 gnd.n280 0.152939
R14079 gnd.n7699 gnd.n7698 0.152939
R14080 gnd.n7700 gnd.n7699 0.152939
R14081 gnd.n7700 gnd.n263 0.152939
R14082 gnd.n7714 gnd.n263 0.152939
R14083 gnd.n7715 gnd.n7714 0.152939
R14084 gnd.n7716 gnd.n7715 0.152939
R14085 gnd.n7716 gnd.n249 0.152939
R14086 gnd.n7730 gnd.n249 0.152939
R14087 gnd.n7731 gnd.n7730 0.152939
R14088 gnd.n7732 gnd.n7731 0.152939
R14089 gnd.n7732 gnd.n234 0.152939
R14090 gnd.n7746 gnd.n234 0.152939
R14091 gnd.n7747 gnd.n7746 0.152939
R14092 gnd.n7748 gnd.n7747 0.152939
R14093 gnd.n7748 gnd.n219 0.152939
R14094 gnd.n7762 gnd.n219 0.152939
R14095 gnd.n7763 gnd.n7762 0.152939
R14096 gnd.n7764 gnd.n7763 0.152939
R14097 gnd.n7765 gnd.n7764 0.152939
R14098 gnd.n7765 gnd.n133 0.152939
R14099 gnd.n7914 gnd.n133 0.152939
R14100 gnd.n7913 gnd.n134 0.152939
R14101 gnd.n136 gnd.n134 0.152939
R14102 gnd.n140 gnd.n136 0.152939
R14103 gnd.n141 gnd.n140 0.152939
R14104 gnd.n142 gnd.n141 0.152939
R14105 gnd.n143 gnd.n142 0.152939
R14106 gnd.n147 gnd.n143 0.152939
R14107 gnd.n148 gnd.n147 0.152939
R14108 gnd.n149 gnd.n148 0.152939
R14109 gnd.n150 gnd.n149 0.152939
R14110 gnd.n154 gnd.n150 0.152939
R14111 gnd.n155 gnd.n154 0.152939
R14112 gnd.n156 gnd.n155 0.152939
R14113 gnd.n157 gnd.n156 0.152939
R14114 gnd.n161 gnd.n157 0.152939
R14115 gnd.n162 gnd.n161 0.152939
R14116 gnd.n163 gnd.n162 0.152939
R14117 gnd.n164 gnd.n163 0.152939
R14118 gnd.n168 gnd.n164 0.152939
R14119 gnd.n169 gnd.n168 0.152939
R14120 gnd.n170 gnd.n169 0.152939
R14121 gnd.n171 gnd.n170 0.152939
R14122 gnd.n175 gnd.n171 0.152939
R14123 gnd.n176 gnd.n175 0.152939
R14124 gnd.n177 gnd.n176 0.152939
R14125 gnd.n178 gnd.n177 0.152939
R14126 gnd.n182 gnd.n178 0.152939
R14127 gnd.n183 gnd.n182 0.152939
R14128 gnd.n184 gnd.n183 0.152939
R14129 gnd.n185 gnd.n184 0.152939
R14130 gnd.n189 gnd.n185 0.152939
R14131 gnd.n190 gnd.n189 0.152939
R14132 gnd.n191 gnd.n190 0.152939
R14133 gnd.n192 gnd.n191 0.152939
R14134 gnd.n196 gnd.n192 0.152939
R14135 gnd.n197 gnd.n196 0.152939
R14136 gnd.n7844 gnd.n197 0.152939
R14137 gnd.n7844 gnd.n7843 0.152939
R14138 gnd.n1941 gnd.n1902 0.152939
R14139 gnd.n1904 gnd.n1902 0.152939
R14140 gnd.n1905 gnd.n1904 0.152939
R14141 gnd.n1906 gnd.n1905 0.152939
R14142 gnd.n1907 gnd.n1906 0.152939
R14143 gnd.n1908 gnd.n1907 0.152939
R14144 gnd.n1909 gnd.n1908 0.152939
R14145 gnd.n1910 gnd.n1909 0.152939
R14146 gnd.n1911 gnd.n1910 0.152939
R14147 gnd.n1912 gnd.n1911 0.152939
R14148 gnd.n1913 gnd.n1912 0.152939
R14149 gnd.n1914 gnd.n1913 0.152939
R14150 gnd.n1915 gnd.n1914 0.152939
R14151 gnd.n1916 gnd.n1915 0.152939
R14152 gnd.n1918 gnd.n1916 0.152939
R14153 gnd.n1918 gnd.n1917 0.152939
R14154 gnd.n1917 gnd.n1591 0.152939
R14155 gnd.n1591 gnd.n1589 0.152939
R14156 gnd.n6169 gnd.n1589 0.152939
R14157 gnd.n6170 gnd.n6169 0.152939
R14158 gnd.n6171 gnd.n6170 0.152939
R14159 gnd.n6172 gnd.n6171 0.152939
R14160 gnd.n6173 gnd.n6172 0.152939
R14161 gnd.n6174 gnd.n6173 0.152939
R14162 gnd.n6175 gnd.n6174 0.152939
R14163 gnd.n6176 gnd.n6175 0.152939
R14164 gnd.n6177 gnd.n6176 0.152939
R14165 gnd.n6178 gnd.n6177 0.152939
R14166 gnd.n6179 gnd.n6178 0.152939
R14167 gnd.n6180 gnd.n6179 0.152939
R14168 gnd.n6181 gnd.n6180 0.152939
R14169 gnd.n6183 gnd.n6181 0.152939
R14170 gnd.n6183 gnd.n6182 0.152939
R14171 gnd.n6182 gnd.n342 0.152939
R14172 gnd.n343 gnd.n342 0.152939
R14173 gnd.n344 gnd.n343 0.152939
R14174 gnd.n345 gnd.n344 0.152939
R14175 gnd.n346 gnd.n345 0.152939
R14176 gnd.n347 gnd.n346 0.152939
R14177 gnd.n348 gnd.n347 0.152939
R14178 gnd.n349 gnd.n348 0.152939
R14179 gnd.n350 gnd.n349 0.152939
R14180 gnd.n351 gnd.n350 0.152939
R14181 gnd.n352 gnd.n351 0.152939
R14182 gnd.n353 gnd.n352 0.152939
R14183 gnd.n354 gnd.n353 0.152939
R14184 gnd.n355 gnd.n354 0.152939
R14185 gnd.n356 gnd.n355 0.152939
R14186 gnd.n357 gnd.n356 0.152939
R14187 gnd.n358 gnd.n357 0.152939
R14188 gnd.n359 gnd.n358 0.152939
R14189 gnd.n360 gnd.n359 0.152939
R14190 gnd.n361 gnd.n360 0.152939
R14191 gnd.n362 gnd.n361 0.152939
R14192 gnd.n363 gnd.n362 0.152939
R14193 gnd.n364 gnd.n363 0.152939
R14194 gnd.n365 gnd.n364 0.152939
R14195 gnd.n366 gnd.n365 0.152939
R14196 gnd.n367 gnd.n366 0.152939
R14197 gnd.n368 gnd.n367 0.152939
R14198 gnd.n370 gnd.n368 0.152939
R14199 gnd.n370 gnd.n369 0.152939
R14200 gnd.n369 gnd.n203 0.152939
R14201 gnd.n7842 gnd.n203 0.152939
R14202 gnd.n6046 gnd.n1687 0.152939
R14203 gnd.n1844 gnd.n1687 0.152939
R14204 gnd.n1845 gnd.n1844 0.152939
R14205 gnd.n1846 gnd.n1845 0.152939
R14206 gnd.n1846 gnd.n1841 0.152939
R14207 gnd.n1854 gnd.n1841 0.152939
R14208 gnd.n1855 gnd.n1854 0.152939
R14209 gnd.n1856 gnd.n1855 0.152939
R14210 gnd.n1856 gnd.n1839 0.152939
R14211 gnd.n1864 gnd.n1839 0.152939
R14212 gnd.n1865 gnd.n1864 0.152939
R14213 gnd.n1866 gnd.n1865 0.152939
R14214 gnd.n1866 gnd.n1837 0.152939
R14215 gnd.n1874 gnd.n1837 0.152939
R14216 gnd.n1875 gnd.n1874 0.152939
R14217 gnd.n1880 gnd.n1879 0.152939
R14218 gnd.n1881 gnd.n1880 0.152939
R14219 gnd.n1882 gnd.n1881 0.152939
R14220 gnd.n1883 gnd.n1882 0.152939
R14221 gnd.n1884 gnd.n1883 0.152939
R14222 gnd.n1885 gnd.n1884 0.152939
R14223 gnd.n1886 gnd.n1885 0.152939
R14224 gnd.n1887 gnd.n1886 0.152939
R14225 gnd.n1888 gnd.n1887 0.152939
R14226 gnd.n1889 gnd.n1888 0.152939
R14227 gnd.n1890 gnd.n1889 0.152939
R14228 gnd.n1891 gnd.n1890 0.152939
R14229 gnd.n1892 gnd.n1891 0.152939
R14230 gnd.n1893 gnd.n1892 0.152939
R14231 gnd.n1894 gnd.n1893 0.152939
R14232 gnd.n1895 gnd.n1894 0.152939
R14233 gnd.n1896 gnd.n1895 0.152939
R14234 gnd.n1946 gnd.n1896 0.152939
R14235 gnd.n1946 gnd.n1945 0.152939
R14236 gnd.n1945 gnd.n1944 0.152939
R14237 gnd.n6048 gnd.n6047 0.152939
R14238 gnd.n6048 gnd.n1662 0.152939
R14239 gnd.n6077 gnd.n1662 0.152939
R14240 gnd.n6078 gnd.n6077 0.152939
R14241 gnd.n6079 gnd.n6078 0.152939
R14242 gnd.n6080 gnd.n6079 0.152939
R14243 gnd.n6080 gnd.n1636 0.152939
R14244 gnd.n6109 gnd.n1636 0.152939
R14245 gnd.n6110 gnd.n6109 0.152939
R14246 gnd.n6111 gnd.n6110 0.152939
R14247 gnd.n6112 gnd.n6111 0.152939
R14248 gnd.n6112 gnd.n1608 0.152939
R14249 gnd.n6147 gnd.n1608 0.152939
R14250 gnd.n6148 gnd.n6147 0.152939
R14251 gnd.n6149 gnd.n6148 0.152939
R14252 gnd.n6150 gnd.n6149 0.152939
R14253 gnd.n6150 gnd.n1571 0.152939
R14254 gnd.n6215 gnd.n1571 0.152939
R14255 gnd.n6216 gnd.n6215 0.152939
R14256 gnd.n6217 gnd.n6216 0.152939
R14257 gnd.n6217 gnd.n1555 0.152939
R14258 gnd.n6235 gnd.n1555 0.152939
R14259 gnd.n6236 gnd.n6235 0.152939
R14260 gnd.n6237 gnd.n6236 0.152939
R14261 gnd.n6238 gnd.n6237 0.152939
R14262 gnd.n6238 gnd.n311 0.152939
R14263 gnd.n7668 gnd.n311 0.152939
R14264 gnd.n4605 gnd.n4604 0.152939
R14265 gnd.n4604 gnd.n2509 0.152939
R14266 gnd.n4682 gnd.n2509 0.152939
R14267 gnd.n4683 gnd.n4682 0.152939
R14268 gnd.n4684 gnd.n4683 0.152939
R14269 gnd.n4684 gnd.n2505 0.152939
R14270 gnd.n4690 gnd.n2505 0.152939
R14271 gnd.n4691 gnd.n4690 0.152939
R14272 gnd.n4692 gnd.n4691 0.152939
R14273 gnd.n4693 gnd.n4692 0.152939
R14274 gnd.n4694 gnd.n4693 0.152939
R14275 gnd.n4697 gnd.n4694 0.152939
R14276 gnd.n4698 gnd.n4697 0.152939
R14277 gnd.n4699 gnd.n4698 0.152939
R14278 gnd.n4700 gnd.n4699 0.152939
R14279 gnd.n4700 gnd.n2472 0.152939
R14280 gnd.n4892 gnd.n2472 0.152939
R14281 gnd.n4893 gnd.n4892 0.152939
R14282 gnd.n4894 gnd.n4893 0.152939
R14283 gnd.n4894 gnd.n2468 0.152939
R14284 gnd.n4900 gnd.n2468 0.152939
R14285 gnd.n4901 gnd.n4900 0.152939
R14286 gnd.n4902 gnd.n4901 0.152939
R14287 gnd.n4902 gnd.n2464 0.152939
R14288 gnd.n4908 gnd.n2464 0.152939
R14289 gnd.n4909 gnd.n4908 0.152939
R14290 gnd.n4910 gnd.n4909 0.152939
R14291 gnd.n4911 gnd.n4910 0.152939
R14292 gnd.n4912 gnd.n4911 0.152939
R14293 gnd.n4913 gnd.n4912 0.152939
R14294 gnd.n4913 gnd.n2313 0.152939
R14295 gnd.n4977 gnd.n2313 0.152939
R14296 gnd.n4978 gnd.n4977 0.152939
R14297 gnd.n4979 gnd.n4978 0.152939
R14298 gnd.n4979 gnd.n2299 0.152939
R14299 gnd.n4993 gnd.n2299 0.152939
R14300 gnd.n4994 gnd.n4993 0.152939
R14301 gnd.n4995 gnd.n4994 0.152939
R14302 gnd.n4995 gnd.n2285 0.152939
R14303 gnd.n5009 gnd.n2285 0.152939
R14304 gnd.n5010 gnd.n5009 0.152939
R14305 gnd.n5011 gnd.n5010 0.152939
R14306 gnd.n5011 gnd.n2271 0.152939
R14307 gnd.n5025 gnd.n2271 0.152939
R14308 gnd.n5026 gnd.n5025 0.152939
R14309 gnd.n5027 gnd.n5026 0.152939
R14310 gnd.n5027 gnd.n2257 0.152939
R14311 gnd.n5041 gnd.n2257 0.152939
R14312 gnd.n5042 gnd.n5041 0.152939
R14313 gnd.n5043 gnd.n5042 0.152939
R14314 gnd.n5043 gnd.n2242 0.152939
R14315 gnd.n5057 gnd.n2242 0.152939
R14316 gnd.n5058 gnd.n5057 0.152939
R14317 gnd.n5059 gnd.n5058 0.152939
R14318 gnd.n5059 gnd.n2227 0.152939
R14319 gnd.n5084 gnd.n2227 0.152939
R14320 gnd.n5085 gnd.n5084 0.152939
R14321 gnd.n5086 gnd.n5085 0.152939
R14322 gnd.n5088 gnd.n5086 0.152939
R14323 gnd.n5088 gnd.n5087 0.152939
R14324 gnd.n5087 gnd.n1371 0.152939
R14325 gnd.n1372 gnd.n1371 0.152939
R14326 gnd.n1373 gnd.n1372 0.152939
R14327 gnd.n5241 gnd.n1373 0.152939
R14328 gnd.n5242 gnd.n5241 0.152939
R14329 gnd.n5242 gnd.n2198 0.152939
R14330 gnd.n5267 gnd.n2198 0.152939
R14331 gnd.n5268 gnd.n5267 0.152939
R14332 gnd.n5269 gnd.n5268 0.152939
R14333 gnd.n5269 gnd.n2179 0.152939
R14334 gnd.n5291 gnd.n2179 0.152939
R14335 gnd.n5292 gnd.n5291 0.152939
R14336 gnd.n5293 gnd.n5292 0.152939
R14337 gnd.n5293 gnd.n2157 0.152939
R14338 gnd.n5317 gnd.n2157 0.152939
R14339 gnd.n5318 gnd.n5317 0.152939
R14340 gnd.n5319 gnd.n5318 0.152939
R14341 gnd.n5320 gnd.n5319 0.152939
R14342 gnd.n5320 gnd.n2128 0.152939
R14343 gnd.n5372 gnd.n2128 0.152939
R14344 gnd.n5373 gnd.n5372 0.152939
R14345 gnd.n5374 gnd.n5373 0.152939
R14346 gnd.n5375 gnd.n5374 0.152939
R14347 gnd.n5375 gnd.n2105 0.152939
R14348 gnd.n5413 gnd.n2105 0.152939
R14349 gnd.n5414 gnd.n5413 0.152939
R14350 gnd.n5415 gnd.n5414 0.152939
R14351 gnd.n5416 gnd.n5415 0.152939
R14352 gnd.n5416 gnd.n2076 0.152939
R14353 gnd.n5454 gnd.n2076 0.152939
R14354 gnd.n5455 gnd.n5454 0.152939
R14355 gnd.n5457 gnd.n5455 0.152939
R14356 gnd.n5457 gnd.n5456 0.152939
R14357 gnd.n5456 gnd.n2054 0.152939
R14358 gnd.n2055 gnd.n2054 0.152939
R14359 gnd.n2056 gnd.n2055 0.152939
R14360 gnd.n2058 gnd.n2056 0.152939
R14361 gnd.n2059 gnd.n2058 0.152939
R14362 gnd.n2059 gnd.n2018 0.152939
R14363 gnd.n5554 gnd.n2018 0.152939
R14364 gnd.n5555 gnd.n5554 0.152939
R14365 gnd.n5556 gnd.n5555 0.152939
R14366 gnd.n5556 gnd.n2002 0.152939
R14367 gnd.n5585 gnd.n2002 0.152939
R14368 gnd.n5586 gnd.n5585 0.152939
R14369 gnd.n5587 gnd.n5586 0.152939
R14370 gnd.n5587 gnd.n1796 0.152939
R14371 gnd.n5760 gnd.n1796 0.152939
R14372 gnd.n5761 gnd.n5760 0.152939
R14373 gnd.n5762 gnd.n5761 0.152939
R14374 gnd.n5762 gnd.n1784 0.152939
R14375 gnd.n5778 gnd.n1784 0.152939
R14376 gnd.n5779 gnd.n5778 0.152939
R14377 gnd.n5780 gnd.n5779 0.152939
R14378 gnd.n5780 gnd.n1773 0.152939
R14379 gnd.n5795 gnd.n1773 0.152939
R14380 gnd.n5796 gnd.n5795 0.152939
R14381 gnd.n5797 gnd.n5796 0.152939
R14382 gnd.n5797 gnd.n1761 0.152939
R14383 gnd.n5812 gnd.n1761 0.152939
R14384 gnd.n5813 gnd.n5812 0.152939
R14385 gnd.n5814 gnd.n5813 0.152939
R14386 gnd.n5814 gnd.n1749 0.152939
R14387 gnd.n5829 gnd.n1749 0.152939
R14388 gnd.n5830 gnd.n5829 0.152939
R14389 gnd.n5831 gnd.n5830 0.152939
R14390 gnd.n5831 gnd.n1737 0.152939
R14391 gnd.n5846 gnd.n1737 0.152939
R14392 gnd.n5847 gnd.n5846 0.152939
R14393 gnd.n5848 gnd.n5847 0.152939
R14394 gnd.n5849 gnd.n5848 0.152939
R14395 gnd.n5849 gnd.n1725 0.152939
R14396 gnd.n5866 gnd.n1725 0.152939
R14397 gnd.n5867 gnd.n5866 0.152939
R14398 gnd.n5868 gnd.n5867 0.152939
R14399 gnd.n5868 gnd.n1722 0.152939
R14400 gnd.n6033 gnd.n1722 0.152939
R14401 gnd.n6034 gnd.n6033 0.152939
R14402 gnd.n6035 gnd.n6034 0.152939
R14403 gnd.n6036 gnd.n6035 0.152939
R14404 gnd.n6036 gnd.n1672 0.152939
R14405 gnd.n6065 gnd.n1672 0.152939
R14406 gnd.n6066 gnd.n6065 0.152939
R14407 gnd.n6067 gnd.n6066 0.152939
R14408 gnd.n6068 gnd.n6067 0.152939
R14409 gnd.n6068 gnd.n1646 0.152939
R14410 gnd.n6098 gnd.n1646 0.152939
R14411 gnd.n6099 gnd.n6098 0.152939
R14412 gnd.n6100 gnd.n6099 0.152939
R14413 gnd.n6101 gnd.n6100 0.152939
R14414 gnd.n6101 gnd.n1618 0.152939
R14415 gnd.n6129 gnd.n1618 0.152939
R14416 gnd.n6130 gnd.n6129 0.152939
R14417 gnd.n6131 gnd.n6130 0.152939
R14418 gnd.n6132 gnd.n6131 0.152939
R14419 gnd.n6133 gnd.n6132 0.152939
R14420 gnd.n6135 gnd.n6133 0.152939
R14421 gnd.n6135 gnd.n6134 0.152939
R14422 gnd.n6134 gnd.n1582 0.152939
R14423 gnd.n1583 gnd.n1582 0.152939
R14424 gnd.n1584 gnd.n1583 0.152939
R14425 gnd.n1585 gnd.n1584 0.152939
R14426 gnd.n1585 gnd.n1545 0.152939
R14427 gnd.n6246 gnd.n1545 0.152939
R14428 gnd.n6247 gnd.n6246 0.152939
R14429 gnd.n6249 gnd.n6247 0.152939
R14430 gnd.n6249 gnd.n6248 0.152939
R14431 gnd.n4397 gnd.n4353 0.152939
R14432 gnd.n4354 gnd.n4353 0.152939
R14433 gnd.n4355 gnd.n4354 0.152939
R14434 gnd.n4356 gnd.n4355 0.152939
R14435 gnd.n4357 gnd.n4356 0.152939
R14436 gnd.n4358 gnd.n4357 0.152939
R14437 gnd.n4359 gnd.n4358 0.152939
R14438 gnd.n4360 gnd.n4359 0.152939
R14439 gnd.n4361 gnd.n4360 0.152939
R14440 gnd.n4362 gnd.n4361 0.152939
R14441 gnd.n4363 gnd.n4362 0.152939
R14442 gnd.n4364 gnd.n4363 0.152939
R14443 gnd.n4365 gnd.n4364 0.152939
R14444 gnd.n4366 gnd.n4365 0.152939
R14445 gnd.n4367 gnd.n4366 0.152939
R14446 gnd.n4368 gnd.n4367 0.152939
R14447 gnd.n4369 gnd.n4368 0.152939
R14448 gnd.n4369 gnd.n2611 0.152939
R14449 gnd.n4524 gnd.n2611 0.152939
R14450 gnd.n4525 gnd.n4524 0.152939
R14451 gnd.n4526 gnd.n4525 0.152939
R14452 gnd.n4526 gnd.n2581 0.152939
R14453 gnd.n4545 gnd.n2581 0.152939
R14454 gnd.n4546 gnd.n4545 0.152939
R14455 gnd.n4548 gnd.n4546 0.152939
R14456 gnd.n4548 gnd.n4547 0.152939
R14457 gnd.n4547 gnd.n2556 0.152939
R14458 gnd.n4573 gnd.n2556 0.152939
R14459 gnd.n4574 gnd.n4573 0.152939
R14460 gnd.n4575 gnd.n4574 0.152939
R14461 gnd.n4576 gnd.n4575 0.152939
R14462 gnd.n4438 gnd.n4327 0.152939
R14463 gnd.n4330 gnd.n4327 0.152939
R14464 gnd.n4331 gnd.n4330 0.152939
R14465 gnd.n4332 gnd.n4331 0.152939
R14466 gnd.n4333 gnd.n4332 0.152939
R14467 gnd.n4336 gnd.n4333 0.152939
R14468 gnd.n4337 gnd.n4336 0.152939
R14469 gnd.n4338 gnd.n4337 0.152939
R14470 gnd.n4339 gnd.n4338 0.152939
R14471 gnd.n4342 gnd.n4339 0.152939
R14472 gnd.n4343 gnd.n4342 0.152939
R14473 gnd.n4344 gnd.n4343 0.152939
R14474 gnd.n4345 gnd.n4344 0.152939
R14475 gnd.n4348 gnd.n4345 0.152939
R14476 gnd.n4349 gnd.n4348 0.152939
R14477 gnd.n4404 gnd.n4349 0.152939
R14478 gnd.n4404 gnd.n4403 0.152939
R14479 gnd.n4403 gnd.n4402 0.152939
R14480 gnd.n4439 gnd.n2664 0.152939
R14481 gnd.n4453 gnd.n2664 0.152939
R14482 gnd.n4454 gnd.n4453 0.152939
R14483 gnd.n4455 gnd.n4454 0.152939
R14484 gnd.n4455 gnd.n2648 0.152939
R14485 gnd.n4469 gnd.n2648 0.152939
R14486 gnd.n4470 gnd.n4469 0.152939
R14487 gnd.n4471 gnd.n4470 0.152939
R14488 gnd.n4471 gnd.n2632 0.152939
R14489 gnd.n4485 gnd.n2632 0.152939
R14490 gnd.n4486 gnd.n4485 0.152939
R14491 gnd.n4487 gnd.n4486 0.152939
R14492 gnd.n4488 gnd.n4487 0.152939
R14493 gnd.n4489 gnd.n4488 0.152939
R14494 gnd.n4490 gnd.n4489 0.152939
R14495 gnd.n4492 gnd.n4490 0.152939
R14496 gnd.n4492 gnd.n4491 0.152939
R14497 gnd.n4491 gnd.n1039 0.152939
R14498 gnd.n1040 gnd.n1039 0.152939
R14499 gnd.n1041 gnd.n1040 0.152939
R14500 gnd.n1059 gnd.n1041 0.152939
R14501 gnd.n1060 gnd.n1059 0.152939
R14502 gnd.n1061 gnd.n1060 0.152939
R14503 gnd.n1062 gnd.n1061 0.152939
R14504 gnd.n1080 gnd.n1062 0.152939
R14505 gnd.n1081 gnd.n1080 0.152939
R14506 gnd.n1082 gnd.n1081 0.152939
R14507 gnd.n1083 gnd.n1082 0.152939
R14508 gnd.n4584 gnd.n1083 0.152939
R14509 gnd.n4585 gnd.n4584 0.152939
R14510 gnd.n4586 gnd.n4585 0.152939
R14511 gnd.n4586 gnd.n2539 0.152939
R14512 gnd.n4619 gnd.n2539 0.152939
R14513 gnd.n4620 gnd.n4619 0.152939
R14514 gnd.n4622 gnd.n4620 0.152939
R14515 gnd.n4622 gnd.n4621 0.152939
R14516 gnd.n4621 gnd.n1108 0.152939
R14517 gnd.n1109 gnd.n1108 0.152939
R14518 gnd.n1110 gnd.n1109 0.152939
R14519 gnd.n1127 gnd.n1110 0.152939
R14520 gnd.n1128 gnd.n1127 0.152939
R14521 gnd.n1129 gnd.n1128 0.152939
R14522 gnd.n1130 gnd.n1129 0.152939
R14523 gnd.n1149 gnd.n1130 0.152939
R14524 gnd.n1150 gnd.n1149 0.152939
R14525 gnd.n1151 gnd.n1150 0.152939
R14526 gnd.n1152 gnd.n1151 0.152939
R14527 gnd.n1170 gnd.n1152 0.152939
R14528 gnd.n1171 gnd.n1170 0.152939
R14529 gnd.n1172 gnd.n1171 0.152939
R14530 gnd.n1173 gnd.n1172 0.152939
R14531 gnd.n1192 gnd.n1173 0.152939
R14532 gnd.n1193 gnd.n1192 0.152939
R14533 gnd.n1194 gnd.n1193 0.152939
R14534 gnd.n1195 gnd.n1194 0.152939
R14535 gnd.n1213 gnd.n1195 0.152939
R14536 gnd.n1214 gnd.n1213 0.152939
R14537 gnd.n1215 gnd.n1214 0.152939
R14538 gnd.n1216 gnd.n1215 0.152939
R14539 gnd.n1235 gnd.n1216 0.152939
R14540 gnd.n1236 gnd.n1235 0.152939
R14541 gnd.n1237 gnd.n1236 0.152939
R14542 gnd.n1238 gnd.n1237 0.152939
R14543 gnd.n2339 gnd.n1238 0.152939
R14544 gnd.n6666 gnd.n1092 0.152939
R14545 gnd.n1117 gnd.n1092 0.152939
R14546 gnd.n1118 gnd.n1117 0.152939
R14547 gnd.n1119 gnd.n1118 0.152939
R14548 gnd.n1138 gnd.n1119 0.152939
R14549 gnd.n1139 gnd.n1138 0.152939
R14550 gnd.n1140 gnd.n1139 0.152939
R14551 gnd.n1141 gnd.n1140 0.152939
R14552 gnd.n1159 gnd.n1141 0.152939
R14553 gnd.n1160 gnd.n1159 0.152939
R14554 gnd.n1161 gnd.n1160 0.152939
R14555 gnd.n1162 gnd.n1161 0.152939
R14556 gnd.n1181 gnd.n1162 0.152939
R14557 gnd.n1182 gnd.n1181 0.152939
R14558 gnd.n1183 gnd.n1182 0.152939
R14559 gnd.n1184 gnd.n1183 0.152939
R14560 gnd.n1202 gnd.n1184 0.152939
R14561 gnd.n1203 gnd.n1202 0.152939
R14562 gnd.n1204 gnd.n1203 0.152939
R14563 gnd.n1205 gnd.n1204 0.152939
R14564 gnd.n1224 gnd.n1205 0.152939
R14565 gnd.n1225 gnd.n1224 0.152939
R14566 gnd.n1226 gnd.n1225 0.152939
R14567 gnd.n1227 gnd.n1226 0.152939
R14568 gnd.n1246 gnd.n1227 0.152939
R14569 gnd.n1247 gnd.n1246 0.152939
R14570 gnd.n6581 gnd.n1247 0.152939
R14571 gnd.n6580 gnd.n1248 0.152939
R14572 gnd.n1282 gnd.n1248 0.152939
R14573 gnd.n1283 gnd.n1282 0.152939
R14574 gnd.n1284 gnd.n1283 0.152939
R14575 gnd.n1285 gnd.n1284 0.152939
R14576 gnd.n1286 gnd.n1285 0.152939
R14577 gnd.n1287 gnd.n1286 0.152939
R14578 gnd.n1288 gnd.n1287 0.152939
R14579 gnd.n1289 gnd.n1288 0.152939
R14580 gnd.n1290 gnd.n1289 0.152939
R14581 gnd.n1291 gnd.n1290 0.152939
R14582 gnd.n1292 gnd.n1291 0.152939
R14583 gnd.n1293 gnd.n1292 0.152939
R14584 gnd.n1294 gnd.n1293 0.152939
R14585 gnd.n1295 gnd.n1294 0.152939
R14586 gnd.n4778 gnd.n4777 0.152939
R14587 gnd.n4779 gnd.n4778 0.152939
R14588 gnd.n4779 gnd.n4773 0.152939
R14589 gnd.n4787 gnd.n4773 0.152939
R14590 gnd.n4788 gnd.n4787 0.152939
R14591 gnd.n4789 gnd.n4788 0.152939
R14592 gnd.n4789 gnd.n4771 0.152939
R14593 gnd.n4797 gnd.n4771 0.152939
R14594 gnd.n4798 gnd.n4797 0.152939
R14595 gnd.n4799 gnd.n4798 0.152939
R14596 gnd.n4799 gnd.n4769 0.152939
R14597 gnd.n4807 gnd.n4769 0.152939
R14598 gnd.n4808 gnd.n4807 0.152939
R14599 gnd.n4809 gnd.n4808 0.152939
R14600 gnd.n4809 gnd.n4767 0.152939
R14601 gnd.n4817 gnd.n4767 0.152939
R14602 gnd.n4818 gnd.n4817 0.152939
R14603 gnd.n4819 gnd.n4818 0.152939
R14604 gnd.n4819 gnd.n4762 0.152939
R14605 gnd.n4825 gnd.n4762 0.152939
R14606 gnd.n4322 gnd.n4292 0.152939
R14607 gnd.n4322 gnd.n4321 0.152939
R14608 gnd.n4321 gnd.n4320 0.152939
R14609 gnd.n4320 gnd.n4293 0.152939
R14610 gnd.n4294 gnd.n4293 0.152939
R14611 gnd.n4295 gnd.n4294 0.152939
R14612 gnd.n4296 gnd.n4295 0.152939
R14613 gnd.n4297 gnd.n4296 0.152939
R14614 gnd.n4298 gnd.n4297 0.152939
R14615 gnd.n4299 gnd.n4298 0.152939
R14616 gnd.n4300 gnd.n4299 0.152939
R14617 gnd.n4301 gnd.n4300 0.152939
R14618 gnd.n4303 gnd.n4301 0.152939
R14619 gnd.n4303 gnd.n4302 0.152939
R14620 gnd.n4302 gnd.n2616 0.152939
R14621 gnd.n2616 gnd.n2614 0.152939
R14622 gnd.n4516 gnd.n2614 0.152939
R14623 gnd.n4517 gnd.n4516 0.152939
R14624 gnd.n4518 gnd.n4517 0.152939
R14625 gnd.n4518 gnd.n2584 0.152939
R14626 gnd.n4532 gnd.n2584 0.152939
R14627 gnd.n4533 gnd.n4532 0.152939
R14628 gnd.n4534 gnd.n4533 0.152939
R14629 gnd.n4535 gnd.n4534 0.152939
R14630 gnd.n4537 gnd.n4535 0.152939
R14631 gnd.n4537 gnd.n4536 0.152939
R14632 gnd.n4536 gnd.n2559 0.152939
R14633 gnd.n2560 gnd.n2559 0.152939
R14634 gnd.n2561 gnd.n2560 0.152939
R14635 gnd.n2562 gnd.n2561 0.152939
R14636 gnd.n2563 gnd.n2562 0.152939
R14637 gnd.n2564 gnd.n2563 0.152939
R14638 gnd.n2565 gnd.n2564 0.152939
R14639 gnd.n2567 gnd.n2565 0.152939
R14640 gnd.n2567 gnd.n2566 0.152939
R14641 gnd.n2566 gnd.n2526 0.152939
R14642 gnd.n2526 gnd.n2524 0.152939
R14643 gnd.n4643 gnd.n2524 0.152939
R14644 gnd.n4644 gnd.n4643 0.152939
R14645 gnd.n4645 gnd.n4644 0.152939
R14646 gnd.n4645 gnd.n2522 0.152939
R14647 gnd.n4653 gnd.n2522 0.152939
R14648 gnd.n4654 gnd.n4653 0.152939
R14649 gnd.n4655 gnd.n4654 0.152939
R14650 gnd.n4656 gnd.n4655 0.152939
R14651 gnd.n4657 gnd.n4656 0.152939
R14652 gnd.n4657 gnd.n2496 0.152939
R14653 gnd.n4724 gnd.n2496 0.152939
R14654 gnd.n4725 gnd.n4724 0.152939
R14655 gnd.n4726 gnd.n4725 0.152939
R14656 gnd.n4726 gnd.n2490 0.152939
R14657 gnd.n4740 gnd.n2490 0.152939
R14658 gnd.n4741 gnd.n4740 0.152939
R14659 gnd.n4742 gnd.n4741 0.152939
R14660 gnd.n4742 gnd.n2488 0.152939
R14661 gnd.n4748 gnd.n2488 0.152939
R14662 gnd.n4749 gnd.n4748 0.152939
R14663 gnd.n4750 gnd.n4749 0.152939
R14664 gnd.n4750 gnd.n2486 0.152939
R14665 gnd.n4758 gnd.n2486 0.152939
R14666 gnd.n4759 gnd.n4758 0.152939
R14667 gnd.n4760 gnd.n4759 0.152939
R14668 gnd.n4761 gnd.n4760 0.152939
R14669 gnd.n4826 gnd.n4761 0.152939
R14670 gnd.n4199 gnd.n2671 0.152939
R14671 gnd.n4200 gnd.n4199 0.152939
R14672 gnd.n4201 gnd.n4200 0.152939
R14673 gnd.n4201 gnd.n4191 0.152939
R14674 gnd.n4209 gnd.n4191 0.152939
R14675 gnd.n4210 gnd.n4209 0.152939
R14676 gnd.n4211 gnd.n4210 0.152939
R14677 gnd.n4211 gnd.n4187 0.152939
R14678 gnd.n4219 gnd.n4187 0.152939
R14679 gnd.n4220 gnd.n4219 0.152939
R14680 gnd.n4221 gnd.n4220 0.152939
R14681 gnd.n4221 gnd.n4183 0.152939
R14682 gnd.n4229 gnd.n4183 0.152939
R14683 gnd.n4230 gnd.n4229 0.152939
R14684 gnd.n4231 gnd.n4230 0.152939
R14685 gnd.n4231 gnd.n4176 0.152939
R14686 gnd.n4239 gnd.n4176 0.152939
R14687 gnd.n4240 gnd.n4239 0.152939
R14688 gnd.n4241 gnd.n4240 0.152939
R14689 gnd.n4241 gnd.n4172 0.152939
R14690 gnd.n4249 gnd.n4172 0.152939
R14691 gnd.n4250 gnd.n4249 0.152939
R14692 gnd.n4251 gnd.n4250 0.152939
R14693 gnd.n4251 gnd.n4168 0.152939
R14694 gnd.n4259 gnd.n4168 0.152939
R14695 gnd.n4260 gnd.n4259 0.152939
R14696 gnd.n4261 gnd.n4260 0.152939
R14697 gnd.n4261 gnd.n4164 0.152939
R14698 gnd.n4269 gnd.n4164 0.152939
R14699 gnd.n4270 gnd.n4269 0.152939
R14700 gnd.n4271 gnd.n4270 0.152939
R14701 gnd.n4271 gnd.n4160 0.152939
R14702 gnd.n4279 gnd.n4160 0.152939
R14703 gnd.n4280 gnd.n4279 0.152939
R14704 gnd.n4282 gnd.n4280 0.152939
R14705 gnd.n4282 gnd.n4281 0.152939
R14706 gnd.n4281 gnd.n4153 0.152939
R14707 gnd.n4291 gnd.n4153 0.152939
R14708 gnd.n4446 gnd.n4445 0.152939
R14709 gnd.n4447 gnd.n4446 0.152939
R14710 gnd.n4447 gnd.n2656 0.152939
R14711 gnd.n4461 gnd.n2656 0.152939
R14712 gnd.n4462 gnd.n4461 0.152939
R14713 gnd.n4463 gnd.n4462 0.152939
R14714 gnd.n4463 gnd.n2639 0.152939
R14715 gnd.n4477 gnd.n2639 0.152939
R14716 gnd.n4478 gnd.n4477 0.152939
R14717 gnd.n4479 gnd.n4478 0.152939
R14718 gnd.n4479 gnd.n2623 0.152939
R14719 gnd.n4503 gnd.n2623 0.152939
R14720 gnd.n4504 gnd.n4503 0.152939
R14721 gnd.n4506 gnd.n4504 0.152939
R14722 gnd.n4506 gnd.n4505 0.152939
R14723 gnd.n4505 gnd.n1027 0.152939
R14724 gnd.n1028 gnd.n1027 0.152939
R14725 gnd.n1029 gnd.n1028 0.152939
R14726 gnd.n1048 gnd.n1029 0.152939
R14727 gnd.n1049 gnd.n1048 0.152939
R14728 gnd.n1050 gnd.n1049 0.152939
R14729 gnd.n1051 gnd.n1050 0.152939
R14730 gnd.n1070 gnd.n1051 0.152939
R14731 gnd.n1071 gnd.n1070 0.152939
R14732 gnd.n1072 gnd.n1071 0.152939
R14733 gnd.n1073 gnd.n1072 0.152939
R14734 gnd.n6666 gnd.n1073 0.152939
R14735 gnd.n2593 gnd.n2589 0.152939
R14736 gnd.n2594 gnd.n2593 0.152939
R14737 gnd.n2595 gnd.n2594 0.152939
R14738 gnd.n2596 gnd.n2595 0.152939
R14739 gnd.n2597 gnd.n2596 0.152939
R14740 gnd.n2598 gnd.n2597 0.152939
R14741 gnd.n2600 gnd.n2598 0.152939
R14742 gnd.n2600 gnd.n2599 0.152939
R14743 gnd.n2599 gnd.n2577 0.152939
R14744 gnd.n6879 gnd.n850 0.152939
R14745 gnd.n855 gnd.n850 0.152939
R14746 gnd.n856 gnd.n855 0.152939
R14747 gnd.n857 gnd.n856 0.152939
R14748 gnd.n862 gnd.n857 0.152939
R14749 gnd.n863 gnd.n862 0.152939
R14750 gnd.n864 gnd.n863 0.152939
R14751 gnd.n865 gnd.n864 0.152939
R14752 gnd.n870 gnd.n865 0.152939
R14753 gnd.n871 gnd.n870 0.152939
R14754 gnd.n872 gnd.n871 0.152939
R14755 gnd.n873 gnd.n872 0.152939
R14756 gnd.n878 gnd.n873 0.152939
R14757 gnd.n879 gnd.n878 0.152939
R14758 gnd.n880 gnd.n879 0.152939
R14759 gnd.n881 gnd.n880 0.152939
R14760 gnd.n886 gnd.n881 0.152939
R14761 gnd.n887 gnd.n886 0.152939
R14762 gnd.n888 gnd.n887 0.152939
R14763 gnd.n889 gnd.n888 0.152939
R14764 gnd.n894 gnd.n889 0.152939
R14765 gnd.n895 gnd.n894 0.152939
R14766 gnd.n896 gnd.n895 0.152939
R14767 gnd.n897 gnd.n896 0.152939
R14768 gnd.n902 gnd.n897 0.152939
R14769 gnd.n903 gnd.n902 0.152939
R14770 gnd.n904 gnd.n903 0.152939
R14771 gnd.n905 gnd.n904 0.152939
R14772 gnd.n910 gnd.n905 0.152939
R14773 gnd.n911 gnd.n910 0.152939
R14774 gnd.n912 gnd.n911 0.152939
R14775 gnd.n913 gnd.n912 0.152939
R14776 gnd.n918 gnd.n913 0.152939
R14777 gnd.n919 gnd.n918 0.152939
R14778 gnd.n920 gnd.n919 0.152939
R14779 gnd.n921 gnd.n920 0.152939
R14780 gnd.n926 gnd.n921 0.152939
R14781 gnd.n927 gnd.n926 0.152939
R14782 gnd.n928 gnd.n927 0.152939
R14783 gnd.n929 gnd.n928 0.152939
R14784 gnd.n934 gnd.n929 0.152939
R14785 gnd.n935 gnd.n934 0.152939
R14786 gnd.n936 gnd.n935 0.152939
R14787 gnd.n937 gnd.n936 0.152939
R14788 gnd.n942 gnd.n937 0.152939
R14789 gnd.n943 gnd.n942 0.152939
R14790 gnd.n944 gnd.n943 0.152939
R14791 gnd.n945 gnd.n944 0.152939
R14792 gnd.n950 gnd.n945 0.152939
R14793 gnd.n951 gnd.n950 0.152939
R14794 gnd.n952 gnd.n951 0.152939
R14795 gnd.n953 gnd.n952 0.152939
R14796 gnd.n958 gnd.n953 0.152939
R14797 gnd.n959 gnd.n958 0.152939
R14798 gnd.n960 gnd.n959 0.152939
R14799 gnd.n961 gnd.n960 0.152939
R14800 gnd.n966 gnd.n961 0.152939
R14801 gnd.n967 gnd.n966 0.152939
R14802 gnd.n968 gnd.n967 0.152939
R14803 gnd.n969 gnd.n968 0.152939
R14804 gnd.n974 gnd.n969 0.152939
R14805 gnd.n975 gnd.n974 0.152939
R14806 gnd.n976 gnd.n975 0.152939
R14807 gnd.n977 gnd.n976 0.152939
R14808 gnd.n982 gnd.n977 0.152939
R14809 gnd.n983 gnd.n982 0.152939
R14810 gnd.n984 gnd.n983 0.152939
R14811 gnd.n985 gnd.n984 0.152939
R14812 gnd.n990 gnd.n985 0.152939
R14813 gnd.n991 gnd.n990 0.152939
R14814 gnd.n992 gnd.n991 0.152939
R14815 gnd.n993 gnd.n992 0.152939
R14816 gnd.n998 gnd.n993 0.152939
R14817 gnd.n999 gnd.n998 0.152939
R14818 gnd.n1000 gnd.n999 0.152939
R14819 gnd.n1001 gnd.n1000 0.152939
R14820 gnd.n1006 gnd.n1001 0.152939
R14821 gnd.n1007 gnd.n1006 0.152939
R14822 gnd.n1008 gnd.n1007 0.152939
R14823 gnd.n1009 gnd.n1008 0.152939
R14824 gnd.n1014 gnd.n1009 0.152939
R14825 gnd.n1015 gnd.n1014 0.152939
R14826 gnd.n1016 gnd.n1015 0.152939
R14827 gnd.n1017 gnd.n1016 0.152939
R14828 gnd.n6003 gnd.n5892 0.152939
R14829 gnd.n6011 gnd.n5892 0.152939
R14830 gnd.n6012 gnd.n6011 0.152939
R14831 gnd.n6013 gnd.n6012 0.152939
R14832 gnd.n6013 gnd.n5888 0.152939
R14833 gnd.n6021 gnd.n5888 0.152939
R14834 gnd.n6022 gnd.n6021 0.152939
R14835 gnd.n6024 gnd.n6022 0.152939
R14836 gnd.n6024 gnd.n6023 0.152939
R14837 gnd.n4985 gnd.n2306 0.152939
R14838 gnd.n4986 gnd.n4985 0.152939
R14839 gnd.n4987 gnd.n4986 0.152939
R14840 gnd.n4987 gnd.n2291 0.152939
R14841 gnd.n5001 gnd.n2291 0.152939
R14842 gnd.n5002 gnd.n5001 0.152939
R14843 gnd.n5003 gnd.n5002 0.152939
R14844 gnd.n5003 gnd.n2278 0.152939
R14845 gnd.n5017 gnd.n2278 0.152939
R14846 gnd.n5018 gnd.n5017 0.152939
R14847 gnd.n5019 gnd.n5018 0.152939
R14848 gnd.n5019 gnd.n2264 0.152939
R14849 gnd.n5033 gnd.n2264 0.152939
R14850 gnd.n5034 gnd.n5033 0.152939
R14851 gnd.n5035 gnd.n5034 0.152939
R14852 gnd.n5035 gnd.n2250 0.152939
R14853 gnd.n5049 gnd.n2250 0.152939
R14854 gnd.n5050 gnd.n5049 0.152939
R14855 gnd.n5051 gnd.n5050 0.152939
R14856 gnd.n5051 gnd.n2236 0.152939
R14857 gnd.n5065 gnd.n2236 0.152939
R14858 gnd.n5066 gnd.n5065 0.152939
R14859 gnd.n5078 gnd.n5066 0.152939
R14860 gnd.n5078 gnd.n5077 0.152939
R14861 gnd.n5077 gnd.n5076 0.152939
R14862 gnd.n5076 gnd.n5067 0.152939
R14863 gnd.n5072 gnd.n5067 0.152939
R14864 gnd.n5072 gnd.n5071 0.152939
R14865 gnd.n5071 gnd.n1383 0.152939
R14866 gnd.n6463 gnd.n1383 0.152939
R14867 gnd.n6463 gnd.n6462 0.152939
R14868 gnd.n6462 gnd.n6461 0.152939
R14869 gnd.n6461 gnd.n1384 0.152939
R14870 gnd.n6457 gnd.n1384 0.152939
R14871 gnd.n6457 gnd.n6456 0.152939
R14872 gnd.n6456 gnd.n6455 0.152939
R14873 gnd.n6455 gnd.n1389 0.152939
R14874 gnd.n6451 gnd.n1389 0.152939
R14875 gnd.n6451 gnd.n6450 0.152939
R14876 gnd.n6450 gnd.n6449 0.152939
R14877 gnd.n6449 gnd.n1394 0.152939
R14878 gnd.n6445 gnd.n1394 0.152939
R14879 gnd.n6445 gnd.n6444 0.152939
R14880 gnd.n6444 gnd.n6443 0.152939
R14881 gnd.n6443 gnd.n1399 0.152939
R14882 gnd.n6439 gnd.n1399 0.152939
R14883 gnd.n6439 gnd.n6438 0.152939
R14884 gnd.n6438 gnd.n6437 0.152939
R14885 gnd.n6437 gnd.n1404 0.152939
R14886 gnd.n6433 gnd.n1404 0.152939
R14887 gnd.n6433 gnd.n6432 0.152939
R14888 gnd.n6432 gnd.n6431 0.152939
R14889 gnd.n6431 gnd.n1409 0.152939
R14890 gnd.n6427 gnd.n1409 0.152939
R14891 gnd.n6427 gnd.n6426 0.152939
R14892 gnd.n6426 gnd.n6425 0.152939
R14893 gnd.n6425 gnd.n1414 0.152939
R14894 gnd.n6421 gnd.n1414 0.152939
R14895 gnd.n6421 gnd.n6420 0.152939
R14896 gnd.n6420 gnd.n6419 0.152939
R14897 gnd.n6419 gnd.n1419 0.152939
R14898 gnd.n6415 gnd.n1419 0.152939
R14899 gnd.n6415 gnd.n6414 0.152939
R14900 gnd.n6414 gnd.n6413 0.152939
R14901 gnd.n6413 gnd.n1424 0.152939
R14902 gnd.n6409 gnd.n1424 0.152939
R14903 gnd.n6409 gnd.n6408 0.152939
R14904 gnd.n6408 gnd.n6407 0.152939
R14905 gnd.n6407 gnd.n1429 0.152939
R14906 gnd.n6403 gnd.n1429 0.152939
R14907 gnd.n6403 gnd.n6402 0.152939
R14908 gnd.n6402 gnd.n6401 0.152939
R14909 gnd.n6401 gnd.n1434 0.152939
R14910 gnd.n6397 gnd.n1434 0.152939
R14911 gnd.n6397 gnd.n6396 0.152939
R14912 gnd.n6396 gnd.n6395 0.152939
R14913 gnd.n6395 gnd.n1439 0.152939
R14914 gnd.n6391 gnd.n1439 0.152939
R14915 gnd.n6391 gnd.n6390 0.152939
R14916 gnd.n6390 gnd.n6389 0.152939
R14917 gnd.n6389 gnd.n1444 0.152939
R14918 gnd.n6385 gnd.n1444 0.152939
R14919 gnd.n6385 gnd.n6384 0.152939
R14920 gnd.n6384 gnd.n6383 0.152939
R14921 gnd.n6383 gnd.n1449 0.152939
R14922 gnd.n6379 gnd.n1449 0.152939
R14923 gnd.n6379 gnd.n6378 0.152939
R14924 gnd.n6378 gnd.n6377 0.152939
R14925 gnd.n6377 gnd.n1454 0.152939
R14926 gnd.n6373 gnd.n1454 0.152939
R14927 gnd.n6373 gnd.n6372 0.152939
R14928 gnd.n6372 gnd.n6371 0.152939
R14929 gnd.n6371 gnd.n1459 0.152939
R14930 gnd.n6367 gnd.n1459 0.152939
R14931 gnd.n6367 gnd.n6366 0.152939
R14932 gnd.n6366 gnd.n6365 0.152939
R14933 gnd.n6365 gnd.n1464 0.152939
R14934 gnd.n6361 gnd.n1464 0.152939
R14935 gnd.n6361 gnd.n6360 0.152939
R14936 gnd.n6360 gnd.n6359 0.152939
R14937 gnd.n6359 gnd.n1469 0.152939
R14938 gnd.n4865 gnd.n4834 0.152939
R14939 gnd.n4865 gnd.n4864 0.152939
R14940 gnd.n4864 gnd.n4863 0.152939
R14941 gnd.n4863 gnd.n4840 0.152939
R14942 gnd.n4859 gnd.n4840 0.152939
R14943 gnd.n4859 gnd.n4858 0.152939
R14944 gnd.n4858 gnd.n4847 0.152939
R14945 gnd.n4854 gnd.n4847 0.152939
R14946 gnd.n4854 gnd.n4853 0.152939
R14947 gnd.n4633 gnd.n2530 0.152939
R14948 gnd.n4634 gnd.n4633 0.152939
R14949 gnd.n4635 gnd.n4634 0.152939
R14950 gnd.n4635 gnd.n2516 0.152939
R14951 gnd.n4673 gnd.n2516 0.152939
R14952 gnd.n4673 gnd.n4672 0.152939
R14953 gnd.n4672 gnd.n4671 0.152939
R14954 gnd.n4671 gnd.n2517 0.152939
R14955 gnd.n4667 gnd.n2517 0.152939
R14956 gnd.n4667 gnd.n4666 0.152939
R14957 gnd.n4666 gnd.n4665 0.152939
R14958 gnd.n4665 gnd.n2499 0.152939
R14959 gnd.n4716 gnd.n2499 0.152939
R14960 gnd.n4717 gnd.n4716 0.152939
R14961 gnd.n4718 gnd.n4717 0.152939
R14962 gnd.n4718 gnd.n2493 0.152939
R14963 gnd.n4732 gnd.n2493 0.152939
R14964 gnd.n4733 gnd.n4732 0.152939
R14965 gnd.n4734 gnd.n4733 0.152939
R14966 gnd.n4734 gnd.n2478 0.152939
R14967 gnd.n4885 gnd.n2478 0.152939
R14968 gnd.n4885 gnd.n4884 0.152939
R14969 gnd.n4884 gnd.n4883 0.152939
R14970 gnd.n4883 gnd.n2479 0.152939
R14971 gnd.n4879 gnd.n2479 0.152939
R14972 gnd.n4879 gnd.n4878 0.152939
R14973 gnd.n4878 gnd.n4877 0.152939
R14974 gnd.n4877 gnd.n2483 0.152939
R14975 gnd.n4873 gnd.n2483 0.152939
R14976 gnd.n4873 gnd.n4872 0.152939
R14977 gnd.n4872 gnd.n4871 0.152939
R14978 gnd.n2401 gnd.n2341 0.152939
R14979 gnd.n2397 gnd.n2341 0.152939
R14980 gnd.n2397 gnd.n2396 0.152939
R14981 gnd.n2396 gnd.n2395 0.152939
R14982 gnd.n2395 gnd.n2344 0.152939
R14983 gnd.n2391 gnd.n2344 0.152939
R14984 gnd.n2391 gnd.n2390 0.152939
R14985 gnd.n2390 gnd.n2389 0.152939
R14986 gnd.n2389 gnd.n2348 0.152939
R14987 gnd.n2385 gnd.n2348 0.152939
R14988 gnd.n2385 gnd.n2384 0.152939
R14989 gnd.n2384 gnd.n2383 0.152939
R14990 gnd.n2383 gnd.n2352 0.152939
R14991 gnd.n2379 gnd.n2352 0.152939
R14992 gnd.n2379 gnd.n2378 0.152939
R14993 gnd.n2378 gnd.n2377 0.152939
R14994 gnd.n2377 gnd.n2356 0.152939
R14995 gnd.n2373 gnd.n2356 0.152939
R14996 gnd.n2373 gnd.n2372 0.152939
R14997 gnd.n2372 gnd.n2371 0.152939
R14998 gnd.n2371 gnd.n2360 0.152939
R14999 gnd.n2367 gnd.n2360 0.152939
R15000 gnd.n2367 gnd.n2366 0.152939
R15001 gnd.n2366 gnd.n2365 0.152939
R15002 gnd.n2365 gnd.n2219 0.152939
R15003 gnd.n5097 gnd.n2219 0.152939
R15004 gnd.n5098 gnd.n5097 0.152939
R15005 gnd.n5099 gnd.n5098 0.152939
R15006 gnd.n5099 gnd.n2217 0.152939
R15007 gnd.n5200 gnd.n2217 0.152939
R15008 gnd.n5201 gnd.n5200 0.152939
R15009 gnd.n5238 gnd.n5201 0.152939
R15010 gnd.n5238 gnd.n5237 0.152939
R15011 gnd.n5237 gnd.n5236 0.152939
R15012 gnd.n5236 gnd.n5202 0.152939
R15013 gnd.n5232 gnd.n5202 0.152939
R15014 gnd.n5232 gnd.n5231 0.152939
R15015 gnd.n5231 gnd.n5230 0.152939
R15016 gnd.n5230 gnd.n5206 0.152939
R15017 gnd.n5226 gnd.n5206 0.152939
R15018 gnd.n5226 gnd.n5225 0.152939
R15019 gnd.n5225 gnd.n5224 0.152939
R15020 gnd.n5224 gnd.n5210 0.152939
R15021 gnd.n5220 gnd.n5210 0.152939
R15022 gnd.n5220 gnd.n5219 0.152939
R15023 gnd.n5219 gnd.n5218 0.152939
R15024 gnd.n5218 gnd.n5213 0.152939
R15025 gnd.n5213 gnd.n2119 0.152939
R15026 gnd.n5382 gnd.n2119 0.152939
R15027 gnd.n5383 gnd.n5382 0.152939
R15028 gnd.n5398 gnd.n5383 0.152939
R15029 gnd.n5398 gnd.n5397 0.152939
R15030 gnd.n5397 gnd.n5396 0.152939
R15031 gnd.n5396 gnd.n5384 0.152939
R15032 gnd.n5392 gnd.n5384 0.152939
R15033 gnd.n5392 gnd.n5391 0.152939
R15034 gnd.n5391 gnd.n5390 0.152939
R15035 gnd.n5390 gnd.n2066 0.152939
R15036 gnd.n5463 gnd.n2066 0.152939
R15037 gnd.n5464 gnd.n5463 0.152939
R15038 gnd.n5465 gnd.n5464 0.152939
R15039 gnd.n5465 gnd.n2064 0.152939
R15040 gnd.n5471 gnd.n2064 0.152939
R15041 gnd.n5472 gnd.n5471 0.152939
R15042 gnd.n5496 gnd.n5472 0.152939
R15043 gnd.n5496 gnd.n5495 0.152939
R15044 gnd.n5495 gnd.n5494 0.152939
R15045 gnd.n5494 gnd.n5473 0.152939
R15046 gnd.n5490 gnd.n5473 0.152939
R15047 gnd.n5490 gnd.n5489 0.152939
R15048 gnd.n5489 gnd.n5488 0.152939
R15049 gnd.n5488 gnd.n5477 0.152939
R15050 gnd.n5484 gnd.n5477 0.152939
R15051 gnd.n5484 gnd.n5483 0.152939
R15052 gnd.n5483 gnd.n5482 0.152939
R15053 gnd.n5482 gnd.n1790 0.152939
R15054 gnd.n5768 gnd.n1790 0.152939
R15055 gnd.n5769 gnd.n5768 0.152939
R15056 gnd.n5770 gnd.n5769 0.152939
R15057 gnd.n5770 gnd.n1779 0.152939
R15058 gnd.n5786 gnd.n1779 0.152939
R15059 gnd.n5787 gnd.n5786 0.152939
R15060 gnd.n5788 gnd.n5787 0.152939
R15061 gnd.n5788 gnd.n1767 0.152939
R15062 gnd.n5803 gnd.n1767 0.152939
R15063 gnd.n5804 gnd.n5803 0.152939
R15064 gnd.n5805 gnd.n5804 0.152939
R15065 gnd.n5805 gnd.n1755 0.152939
R15066 gnd.n5820 gnd.n1755 0.152939
R15067 gnd.n5821 gnd.n5820 0.152939
R15068 gnd.n5822 gnd.n5821 0.152939
R15069 gnd.n5822 gnd.n1742 0.152939
R15070 gnd.n5837 gnd.n1742 0.152939
R15071 gnd.n5838 gnd.n5837 0.152939
R15072 gnd.n5839 gnd.n5838 0.152939
R15073 gnd.n5839 gnd.n1731 0.152939
R15074 gnd.n5856 gnd.n1731 0.152939
R15075 gnd.n5857 gnd.n5856 0.152939
R15076 gnd.n5858 gnd.n5857 0.152939
R15077 gnd.n5858 gnd.n1478 0.152939
R15078 gnd.n6352 gnd.n1478 0.152939
R15079 gnd.n6349 gnd.n1481 0.152939
R15080 gnd.n6345 gnd.n1481 0.152939
R15081 gnd.n6345 gnd.n6344 0.152939
R15082 gnd.n6344 gnd.n6343 0.152939
R15083 gnd.n6343 gnd.n1486 0.152939
R15084 gnd.n6339 gnd.n1486 0.152939
R15085 gnd.n6339 gnd.n6338 0.152939
R15086 gnd.n6338 gnd.n6337 0.152939
R15087 gnd.n6337 gnd.n1491 0.152939
R15088 gnd.n6333 gnd.n1491 0.152939
R15089 gnd.n6333 gnd.n6332 0.152939
R15090 gnd.n6332 gnd.n6331 0.152939
R15091 gnd.n6331 gnd.n1496 0.152939
R15092 gnd.n6327 gnd.n1496 0.152939
R15093 gnd.n6327 gnd.n6326 0.152939
R15094 gnd.n6326 gnd.n6325 0.152939
R15095 gnd.n6325 gnd.n1501 0.152939
R15096 gnd.n6321 gnd.n1501 0.152939
R15097 gnd.n6321 gnd.n6320 0.152939
R15098 gnd.n6320 gnd.n6319 0.152939
R15099 gnd.n6319 gnd.n1506 0.152939
R15100 gnd.n6315 gnd.n1506 0.152939
R15101 gnd.n6315 gnd.n6314 0.152939
R15102 gnd.n6314 gnd.n6313 0.152939
R15103 gnd.n6313 gnd.n1511 0.152939
R15104 gnd.n6309 gnd.n1511 0.152939
R15105 gnd.n6309 gnd.n6308 0.152939
R15106 gnd.n6308 gnd.n328 0.152939
R15107 gnd.n7660 gnd.n328 0.152939
R15108 gnd.n7660 gnd.n7659 0.152939
R15109 gnd.n7659 gnd.n7658 0.152939
R15110 gnd.n7658 gnd.n329 0.152939
R15111 gnd.n7654 gnd.n329 0.152939
R15112 gnd.n7654 gnd.n7653 0.152939
R15113 gnd.n7653 gnd.n7652 0.152939
R15114 gnd.n7652 gnd.n303 0.152939
R15115 gnd.n7674 gnd.n303 0.152939
R15116 gnd.n7675 gnd.n7674 0.152939
R15117 gnd.n7676 gnd.n7675 0.152939
R15118 gnd.n7676 gnd.n288 0.152939
R15119 gnd.n7690 gnd.n288 0.152939
R15120 gnd.n7691 gnd.n7690 0.152939
R15121 gnd.n7692 gnd.n7691 0.152939
R15122 gnd.n7692 gnd.n272 0.152939
R15123 gnd.n7706 gnd.n272 0.152939
R15124 gnd.n7707 gnd.n7706 0.152939
R15125 gnd.n7708 gnd.n7707 0.152939
R15126 gnd.n7708 gnd.n256 0.152939
R15127 gnd.n7722 gnd.n256 0.152939
R15128 gnd.n7723 gnd.n7722 0.152939
R15129 gnd.n7724 gnd.n7723 0.152939
R15130 gnd.n7724 gnd.n240 0.152939
R15131 gnd.n7738 gnd.n240 0.152939
R15132 gnd.n7739 gnd.n7738 0.152939
R15133 gnd.n7740 gnd.n7739 0.152939
R15134 gnd.n7740 gnd.n226 0.152939
R15135 gnd.n7754 gnd.n226 0.152939
R15136 gnd.n7755 gnd.n7754 0.152939
R15137 gnd.n7756 gnd.n7755 0.152939
R15138 gnd.n7756 gnd.n209 0.152939
R15139 gnd.n7772 gnd.n209 0.152939
R15140 gnd.n7773 gnd.n7772 0.152939
R15141 gnd.n7835 gnd.n7773 0.152939
R15142 gnd.n7835 gnd.n7834 0.152939
R15143 gnd.n7833 gnd.n7774 0.152939
R15144 gnd.n7829 gnd.n7774 0.152939
R15145 gnd.n7829 gnd.n7828 0.152939
R15146 gnd.n7828 gnd.n7827 0.152939
R15147 gnd.n7827 gnd.n7780 0.152939
R15148 gnd.n7823 gnd.n7780 0.152939
R15149 gnd.n7823 gnd.n7822 0.152939
R15150 gnd.n7822 gnd.n7821 0.152939
R15151 gnd.n7821 gnd.n7788 0.152939
R15152 gnd.n7817 gnd.n7788 0.152939
R15153 gnd.n7817 gnd.n7816 0.152939
R15154 gnd.n7816 gnd.n7815 0.152939
R15155 gnd.n7815 gnd.n7796 0.152939
R15156 gnd.n7811 gnd.n7796 0.152939
R15157 gnd.n7811 gnd.n7810 0.152939
R15158 gnd.n7810 gnd.n7809 0.152939
R15159 gnd.n7809 gnd.n121 0.152939
R15160 gnd.n7921 gnd.n121 0.152939
R15161 gnd.n6056 gnd.n6055 0.152939
R15162 gnd.n6058 gnd.n6056 0.152939
R15163 gnd.n6058 gnd.n6057 0.152939
R15164 gnd.n6057 gnd.n1653 0.152939
R15165 gnd.n6087 gnd.n1653 0.152939
R15166 gnd.n6088 gnd.n6087 0.152939
R15167 gnd.n6090 gnd.n6088 0.152939
R15168 gnd.n6090 gnd.n6089 0.152939
R15169 gnd.n6089 gnd.n1627 0.152939
R15170 gnd.n6119 gnd.n1627 0.152939
R15171 gnd.n6120 gnd.n6119 0.152939
R15172 gnd.n6122 gnd.n6120 0.152939
R15173 gnd.n6122 gnd.n6121 0.152939
R15174 gnd.n6121 gnd.n1597 0.152939
R15175 gnd.n6157 gnd.n1597 0.152939
R15176 gnd.n6158 gnd.n6157 0.152939
R15177 gnd.n6160 gnd.n6158 0.152939
R15178 gnd.n6160 gnd.n6159 0.152939
R15179 gnd.n6159 gnd.n1564 0.152939
R15180 gnd.n6223 gnd.n1564 0.152939
R15181 gnd.n6224 gnd.n6223 0.152939
R15182 gnd.n6228 gnd.n6224 0.152939
R15183 gnd.n6228 gnd.n6227 0.152939
R15184 gnd.n6227 gnd.n6226 0.152939
R15185 gnd.n6226 gnd.n1526 0.152939
R15186 gnd.n6299 gnd.n1526 0.152939
R15187 gnd.n6299 gnd.n6298 0.152939
R15188 gnd.n6298 gnd.n6297 0.152939
R15189 gnd.n6297 gnd.n1527 0.152939
R15190 gnd.n6293 gnd.n1527 0.152939
R15191 gnd.n6293 gnd.n79 0.152939
R15192 gnd.n7970 gnd.n79 0.152939
R15193 gnd.n7970 gnd.n7969 0.152939
R15194 gnd.n7969 gnd.n81 0.152939
R15195 gnd.n7965 gnd.n81 0.152939
R15196 gnd.n7965 gnd.n7964 0.152939
R15197 gnd.n7964 gnd.n7963 0.152939
R15198 gnd.n7963 gnd.n86 0.152939
R15199 gnd.n7959 gnd.n86 0.152939
R15200 gnd.n7959 gnd.n7958 0.152939
R15201 gnd.n7958 gnd.n7957 0.152939
R15202 gnd.n7957 gnd.n91 0.152939
R15203 gnd.n7953 gnd.n91 0.152939
R15204 gnd.n7953 gnd.n7952 0.152939
R15205 gnd.n7952 gnd.n7951 0.152939
R15206 gnd.n7951 gnd.n96 0.152939
R15207 gnd.n7947 gnd.n96 0.152939
R15208 gnd.n7947 gnd.n7946 0.152939
R15209 gnd.n7946 gnd.n7945 0.152939
R15210 gnd.n7945 gnd.n101 0.152939
R15211 gnd.n7941 gnd.n101 0.152939
R15212 gnd.n7941 gnd.n7940 0.152939
R15213 gnd.n7940 gnd.n7939 0.152939
R15214 gnd.n7939 gnd.n106 0.152939
R15215 gnd.n7935 gnd.n106 0.152939
R15216 gnd.n7935 gnd.n7934 0.152939
R15217 gnd.n7934 gnd.n7933 0.152939
R15218 gnd.n7933 gnd.n111 0.152939
R15219 gnd.n7929 gnd.n111 0.152939
R15220 gnd.n7929 gnd.n7928 0.152939
R15221 gnd.n7928 gnd.n7927 0.152939
R15222 gnd.n7927 gnd.n116 0.152939
R15223 gnd.n7923 gnd.n116 0.152939
R15224 gnd.n7923 gnd.n7922 0.152939
R15225 gnd.n6003 gnd.n1680 0.151415
R15226 gnd.n4870 gnd.n4834 0.151415
R15227 gnd.n4577 gnd.n4576 0.145814
R15228 gnd.n4577 gnd.n2530 0.145814
R15229 gnd.n6266 gnd.n312 0.116354
R15230 gnd.n2577 gnd.n1093 0.116354
R15231 gnd.n3545 gnd.n3544 0.0767195
R15232 gnd.n3544 gnd.n3543 0.0767195
R15233 gnd.n2402 gnd.n2340 0.063
R15234 gnd.n6351 gnd.n6350 0.063
R15235 gnd.n4111 gnd.n2714 0.0477147
R15236 gnd.n3308 gnd.n3196 0.0442063
R15237 gnd.n3309 gnd.n3308 0.0442063
R15238 gnd.n3310 gnd.n3309 0.0442063
R15239 gnd.n3310 gnd.n3185 0.0442063
R15240 gnd.n3324 gnd.n3185 0.0442063
R15241 gnd.n3325 gnd.n3324 0.0442063
R15242 gnd.n3326 gnd.n3325 0.0442063
R15243 gnd.n3326 gnd.n3172 0.0442063
R15244 gnd.n3370 gnd.n3172 0.0442063
R15245 gnd.n3371 gnd.n3370 0.0442063
R15246 gnd.n4605 gnd.n1093 0.0370854
R15247 gnd.n6248 gnd.n312 0.0370854
R15248 gnd.n3373 gnd.n3106 0.0344674
R15249 gnd.n6001 gnd.n6000 0.0343753
R15250 gnd.n4869 gnd.n2458 0.0343753
R15251 gnd.n3393 gnd.n3392 0.0269946
R15252 gnd.n3395 gnd.n3394 0.0269946
R15253 gnd.n3101 gnd.n3099 0.0269946
R15254 gnd.n3405 gnd.n3403 0.0269946
R15255 gnd.n3404 gnd.n3080 0.0269946
R15256 gnd.n3424 gnd.n3423 0.0269946
R15257 gnd.n3426 gnd.n3425 0.0269946
R15258 gnd.n3075 gnd.n3074 0.0269946
R15259 gnd.n3436 gnd.n3070 0.0269946
R15260 gnd.n3435 gnd.n3072 0.0269946
R15261 gnd.n3071 gnd.n3053 0.0269946
R15262 gnd.n3456 gnd.n3054 0.0269946
R15263 gnd.n3455 gnd.n3055 0.0269946
R15264 gnd.n3489 gnd.n3030 0.0269946
R15265 gnd.n3491 gnd.n3490 0.0269946
R15266 gnd.n3492 gnd.n2977 0.0269946
R15267 gnd.n3025 gnd.n2978 0.0269946
R15268 gnd.n3027 gnd.n2979 0.0269946
R15269 gnd.n3502 gnd.n3501 0.0269946
R15270 gnd.n3504 gnd.n3503 0.0269946
R15271 gnd.n3505 gnd.n2999 0.0269946
R15272 gnd.n3507 gnd.n3000 0.0269946
R15273 gnd.n3510 gnd.n3001 0.0269946
R15274 gnd.n3513 gnd.n3512 0.0269946
R15275 gnd.n3515 gnd.n3514 0.0269946
R15276 gnd.n3580 gnd.n2888 0.0269946
R15277 gnd.n3582 gnd.n3581 0.0269946
R15278 gnd.n3591 gnd.n2881 0.0269946
R15279 gnd.n3593 gnd.n3592 0.0269946
R15280 gnd.n3594 gnd.n2879 0.0269946
R15281 gnd.n3601 gnd.n3597 0.0269946
R15282 gnd.n3600 gnd.n3599 0.0269946
R15283 gnd.n3598 gnd.n2858 0.0269946
R15284 gnd.n3623 gnd.n2859 0.0269946
R15285 gnd.n3622 gnd.n2860 0.0269946
R15286 gnd.n3665 gnd.n2833 0.0269946
R15287 gnd.n3667 gnd.n3666 0.0269946
R15288 gnd.n3676 gnd.n2826 0.0269946
R15289 gnd.n3678 gnd.n3677 0.0269946
R15290 gnd.n3679 gnd.n2824 0.0269946
R15291 gnd.n3686 gnd.n3682 0.0269946
R15292 gnd.n3685 gnd.n3684 0.0269946
R15293 gnd.n3683 gnd.n2803 0.0269946
R15294 gnd.n3708 gnd.n2804 0.0269946
R15295 gnd.n3707 gnd.n2805 0.0269946
R15296 gnd.n3754 gnd.n2778 0.0269946
R15297 gnd.n3756 gnd.n3755 0.0269946
R15298 gnd.n3765 gnd.n2771 0.0269946
R15299 gnd.n4024 gnd.n2769 0.0269946
R15300 gnd.n4029 gnd.n4027 0.0269946
R15301 gnd.n4028 gnd.n2750 0.0269946
R15302 gnd.n4053 gnd.n4052 0.0269946
R15303 gnd.n6351 gnd.n1479 0.0245515
R15304 gnd.n2403 gnd.n2402 0.0245515
R15305 gnd.n3373 gnd.n3372 0.0202011
R15306 gnd.n5930 gnd.n1479 0.0174377
R15307 gnd.n5935 gnd.n5930 0.0174377
R15308 gnd.n5936 gnd.n5935 0.0174377
R15309 gnd.n5936 gnd.n5928 0.0174377
R15310 gnd.n5941 gnd.n5928 0.0174377
R15311 gnd.n5942 gnd.n5941 0.0174377
R15312 gnd.n5942 gnd.n5924 0.0174377
R15313 gnd.n5947 gnd.n5924 0.0174377
R15314 gnd.n5948 gnd.n5947 0.0174377
R15315 gnd.n5948 gnd.n5920 0.0174377
R15316 gnd.n5953 gnd.n5920 0.0174377
R15317 gnd.n5954 gnd.n5953 0.0174377
R15318 gnd.n5954 gnd.n5918 0.0174377
R15319 gnd.n5959 gnd.n5918 0.0174377
R15320 gnd.n5960 gnd.n5959 0.0174377
R15321 gnd.n5960 gnd.n5916 0.0174377
R15322 gnd.n5965 gnd.n5916 0.0174377
R15323 gnd.n5966 gnd.n5965 0.0174377
R15324 gnd.n5966 gnd.n5912 0.0174377
R15325 gnd.n5971 gnd.n5912 0.0174377
R15326 gnd.n5972 gnd.n5971 0.0174377
R15327 gnd.n5972 gnd.n5908 0.0174377
R15328 gnd.n5977 gnd.n5908 0.0174377
R15329 gnd.n5978 gnd.n5977 0.0174377
R15330 gnd.n5978 gnd.n5906 0.0174377
R15331 gnd.n5983 gnd.n5906 0.0174377
R15332 gnd.n5985 gnd.n5983 0.0174377
R15333 gnd.n5985 gnd.n5984 0.0174377
R15334 gnd.n5984 gnd.n5904 0.0174377
R15335 gnd.n5995 gnd.n5904 0.0174377
R15336 gnd.n5995 gnd.n5994 0.0174377
R15337 gnd.n5994 gnd.n5897 0.0174377
R15338 gnd.n5897 gnd.n5896 0.0174377
R15339 gnd.n5999 gnd.n5896 0.0174377
R15340 gnd.n6000 gnd.n5999 0.0174377
R15341 gnd.n2403 gnd.n2333 0.0174377
R15342 gnd.n2335 gnd.n2333 0.0174377
R15343 gnd.n4968 gnd.n2335 0.0174377
R15344 gnd.n4968 gnd.n4967 0.0174377
R15345 gnd.n4967 gnd.n2336 0.0174377
R15346 gnd.n4964 gnd.n2336 0.0174377
R15347 gnd.n4964 gnd.n4963 0.0174377
R15348 gnd.n4963 gnd.n2411 0.0174377
R15349 gnd.n4960 gnd.n2411 0.0174377
R15350 gnd.n4960 gnd.n4959 0.0174377
R15351 gnd.n4959 gnd.n2416 0.0174377
R15352 gnd.n4956 gnd.n2416 0.0174377
R15353 gnd.n4956 gnd.n4955 0.0174377
R15354 gnd.n4955 gnd.n2420 0.0174377
R15355 gnd.n4952 gnd.n2420 0.0174377
R15356 gnd.n4952 gnd.n4951 0.0174377
R15357 gnd.n4951 gnd.n2424 0.0174377
R15358 gnd.n4948 gnd.n2424 0.0174377
R15359 gnd.n4948 gnd.n4947 0.0174377
R15360 gnd.n4947 gnd.n2430 0.0174377
R15361 gnd.n4944 gnd.n2430 0.0174377
R15362 gnd.n4944 gnd.n4943 0.0174377
R15363 gnd.n4943 gnd.n2436 0.0174377
R15364 gnd.n4940 gnd.n2436 0.0174377
R15365 gnd.n4940 gnd.n4939 0.0174377
R15366 gnd.n4939 gnd.n2440 0.0174377
R15367 gnd.n4936 gnd.n2440 0.0174377
R15368 gnd.n4936 gnd.n4935 0.0174377
R15369 gnd.n4935 gnd.n2444 0.0174377
R15370 gnd.n4932 gnd.n2444 0.0174377
R15371 gnd.n4932 gnd.n4931 0.0174377
R15372 gnd.n4931 gnd.n2452 0.0174377
R15373 gnd.n4928 gnd.n2452 0.0174377
R15374 gnd.n4928 gnd.n4927 0.0174377
R15375 gnd.n4927 gnd.n2458 0.0174377
R15376 gnd.n3372 gnd.n3371 0.0148637
R15377 gnd.n4022 gnd.n3766 0.0144266
R15378 gnd.n4023 gnd.n4022 0.0130679
R15379 gnd.n3392 gnd.n3106 0.00797283
R15380 gnd.n3394 gnd.n3393 0.00797283
R15381 gnd.n3395 gnd.n3101 0.00797283
R15382 gnd.n3403 gnd.n3099 0.00797283
R15383 gnd.n3405 gnd.n3404 0.00797283
R15384 gnd.n3423 gnd.n3080 0.00797283
R15385 gnd.n3425 gnd.n3424 0.00797283
R15386 gnd.n3426 gnd.n3075 0.00797283
R15387 gnd.n3074 gnd.n3070 0.00797283
R15388 gnd.n3436 gnd.n3435 0.00797283
R15389 gnd.n3072 gnd.n3071 0.00797283
R15390 gnd.n3054 gnd.n3053 0.00797283
R15391 gnd.n3456 gnd.n3455 0.00797283
R15392 gnd.n3055 gnd.n3030 0.00797283
R15393 gnd.n3490 gnd.n3489 0.00797283
R15394 gnd.n3492 gnd.n3491 0.00797283
R15395 gnd.n3025 gnd.n2977 0.00797283
R15396 gnd.n3027 gnd.n2978 0.00797283
R15397 gnd.n3501 gnd.n2979 0.00797283
R15398 gnd.n3503 gnd.n3502 0.00797283
R15399 gnd.n3505 gnd.n3504 0.00797283
R15400 gnd.n3507 gnd.n2999 0.00797283
R15401 gnd.n3510 gnd.n3000 0.00797283
R15402 gnd.n3512 gnd.n3001 0.00797283
R15403 gnd.n3515 gnd.n3513 0.00797283
R15404 gnd.n3514 gnd.n2888 0.00797283
R15405 gnd.n3582 gnd.n3580 0.00797283
R15406 gnd.n3581 gnd.n2881 0.00797283
R15407 gnd.n3592 gnd.n3591 0.00797283
R15408 gnd.n3594 gnd.n3593 0.00797283
R15409 gnd.n3597 gnd.n2879 0.00797283
R15410 gnd.n3601 gnd.n3600 0.00797283
R15411 gnd.n3599 gnd.n3598 0.00797283
R15412 gnd.n2859 gnd.n2858 0.00797283
R15413 gnd.n3623 gnd.n3622 0.00797283
R15414 gnd.n2860 gnd.n2833 0.00797283
R15415 gnd.n3667 gnd.n3665 0.00797283
R15416 gnd.n3666 gnd.n2826 0.00797283
R15417 gnd.n3677 gnd.n3676 0.00797283
R15418 gnd.n3679 gnd.n3678 0.00797283
R15419 gnd.n3682 gnd.n2824 0.00797283
R15420 gnd.n3686 gnd.n3685 0.00797283
R15421 gnd.n3684 gnd.n3683 0.00797283
R15422 gnd.n2804 gnd.n2803 0.00797283
R15423 gnd.n3708 gnd.n3707 0.00797283
R15424 gnd.n2805 gnd.n2778 0.00797283
R15425 gnd.n3756 gnd.n3754 0.00797283
R15426 gnd.n3755 gnd.n2771 0.00797283
R15427 gnd.n3766 gnd.n3765 0.00797283
R15428 gnd.n4024 gnd.n4023 0.00797283
R15429 gnd.n4027 gnd.n2769 0.00797283
R15430 gnd.n4029 gnd.n4028 0.00797283
R15431 gnd.n4052 gnd.n2750 0.00797283
R15432 gnd.n4053 gnd.n2714 0.00797283
R15433 gnd.n6183 gnd.n329 0.00433921
R15434 gnd.n2564 gnd.n2539 0.00433921
R15435 gnd.n6001 gnd.n1680 0.000838753
R15436 gnd.n4870 gnd.n4869 0.000838753
R15437 a_n2982_13878.n74 a_n2982_13878.t50 532.5
R15438 a_n2982_13878.n149 a_n2982_13878.t38 512.366
R15439 a_n2982_13878.n148 a_n2982_13878.t52 512.366
R15440 a_n2982_13878.n83 a_n2982_13878.t44 512.366
R15441 a_n2982_13878.n147 a_n2982_13878.t34 512.366
R15442 a_n2982_13878.n146 a_n2982_13878.t58 512.366
R15443 a_n2982_13878.n84 a_n2982_13878.t46 512.366
R15444 a_n2982_13878.n145 a_n2982_13878.t28 512.366
R15445 a_n2982_13878.n144 a_n2982_13878.t56 512.366
R15446 a_n2982_13878.n85 a_n2982_13878.t16 512.366
R15447 a_n2982_13878.n143 a_n2982_13878.t30 512.366
R15448 a_n2982_13878.n12 a_n2982_13878.t102 538.698
R15449 a_n2982_13878.n134 a_n2982_13878.t79 512.366
R15450 a_n2982_13878.n133 a_n2982_13878.t84 512.366
R15451 a_n2982_13878.n86 a_n2982_13878.t72 512.366
R15452 a_n2982_13878.n132 a_n2982_13878.t89 512.366
R15453 a_n2982_13878.n131 a_n2982_13878.t98 512.366
R15454 a_n2982_13878.n87 a_n2982_13878.t99 512.366
R15455 a_n2982_13878.n130 a_n2982_13878.t66 512.366
R15456 a_n2982_13878.n129 a_n2982_13878.t81 512.366
R15457 a_n2982_13878.n88 a_n2982_13878.t69 512.366
R15458 a_n2982_13878.n128 a_n2982_13878.t76 512.366
R15459 a_n2982_13878.n27 a_n2982_13878.t48 538.698
R15460 a_n2982_13878.n108 a_n2982_13878.t20 512.366
R15461 a_n2982_13878.n97 a_n2982_13878.t60 512.366
R15462 a_n2982_13878.n109 a_n2982_13878.t40 512.366
R15463 a_n2982_13878.n96 a_n2982_13878.t24 512.366
R15464 a_n2982_13878.n110 a_n2982_13878.t42 512.366
R15465 a_n2982_13878.n111 a_n2982_13878.t32 512.366
R15466 a_n2982_13878.n95 a_n2982_13878.t62 512.366
R15467 a_n2982_13878.n112 a_n2982_13878.t54 512.366
R15468 a_n2982_13878.n94 a_n2982_13878.t22 512.366
R15469 a_n2982_13878.n113 a_n2982_13878.t18 512.366
R15470 a_n2982_13878.n33 a_n2982_13878.t101 538.698
R15471 a_n2982_13878.n102 a_n2982_13878.t70 512.366
R15472 a_n2982_13878.n101 a_n2982_13878.t71 512.366
R15473 a_n2982_13878.n103 a_n2982_13878.t96 512.366
R15474 a_n2982_13878.n100 a_n2982_13878.t97 512.366
R15475 a_n2982_13878.n104 a_n2982_13878.t68 512.366
R15476 a_n2982_13878.n105 a_n2982_13878.t92 512.366
R15477 a_n2982_13878.n99 a_n2982_13878.t93 512.366
R15478 a_n2982_13878.n106 a_n2982_13878.t65 512.366
R15479 a_n2982_13878.n98 a_n2982_13878.t78 512.366
R15480 a_n2982_13878.n107 a_n2982_13878.t87 512.366
R15481 a_n2982_13878.n125 a_n2982_13878.t86 512.366
R15482 a_n2982_13878.n115 a_n2982_13878.t75 512.366
R15483 a_n2982_13878.n126 a_n2982_13878.t64 512.366
R15484 a_n2982_13878.n123 a_n2982_13878.t94 512.366
R15485 a_n2982_13878.n116 a_n2982_13878.t83 512.366
R15486 a_n2982_13878.n124 a_n2982_13878.t82 512.366
R15487 a_n2982_13878.n121 a_n2982_13878.t90 512.366
R15488 a_n2982_13878.n117 a_n2982_13878.t73 512.366
R15489 a_n2982_13878.n122 a_n2982_13878.t74 512.366
R15490 a_n2982_13878.n119 a_n2982_13878.t77 512.366
R15491 a_n2982_13878.n118 a_n2982_13878.t88 512.366
R15492 a_n2982_13878.n120 a_n2982_13878.t103 512.366
R15493 a_n2982_13878.n35 a_n2982_13878.n34 44.7878
R15494 a_n2982_13878.n73 a_n2982_13878.n7 70.5844
R15495 a_n2982_13878.n23 a_n2982_13878.n57 70.5844
R15496 a_n2982_13878.n29 a_n2982_13878.n49 70.5844
R15497 a_n2982_13878.n48 a_n2982_13878.n29 70.1674
R15498 a_n2982_13878.n48 a_n2982_13878.n98 20.9683
R15499 a_n2982_13878.n28 a_n2982_13878.n47 74.73
R15500 a_n2982_13878.n106 a_n2982_13878.n47 11.843
R15501 a_n2982_13878.n46 a_n2982_13878.n28 80.4688
R15502 a_n2982_13878.n46 a_n2982_13878.n99 0.365327
R15503 a_n2982_13878.n30 a_n2982_13878.n45 75.0448
R15504 a_n2982_13878.n44 a_n2982_13878.n30 70.1674
R15505 a_n2982_13878.n44 a_n2982_13878.n100 20.9683
R15506 a_n2982_13878.n31 a_n2982_13878.n43 70.3058
R15507 a_n2982_13878.n103 a_n2982_13878.n43 20.6913
R15508 a_n2982_13878.n42 a_n2982_13878.n31 75.3623
R15509 a_n2982_13878.n42 a_n2982_13878.n101 10.5784
R15510 a_n2982_13878.n33 a_n2982_13878.n32 44.7878
R15511 a_n2982_13878.n56 a_n2982_13878.n23 70.1674
R15512 a_n2982_13878.n56 a_n2982_13878.n94 20.9683
R15513 a_n2982_13878.n22 a_n2982_13878.n55 74.73
R15514 a_n2982_13878.n112 a_n2982_13878.n55 11.843
R15515 a_n2982_13878.n54 a_n2982_13878.n22 80.4688
R15516 a_n2982_13878.n54 a_n2982_13878.n95 0.365327
R15517 a_n2982_13878.n24 a_n2982_13878.n53 75.0448
R15518 a_n2982_13878.n52 a_n2982_13878.n24 70.1674
R15519 a_n2982_13878.n52 a_n2982_13878.n96 20.9683
R15520 a_n2982_13878.n25 a_n2982_13878.n51 70.3058
R15521 a_n2982_13878.n109 a_n2982_13878.n51 20.6913
R15522 a_n2982_13878.n50 a_n2982_13878.n25 75.3623
R15523 a_n2982_13878.n50 a_n2982_13878.n97 10.5784
R15524 a_n2982_13878.n27 a_n2982_13878.n26 44.7878
R15525 a_n2982_13878.n13 a_n2982_13878.n65 70.1674
R15526 a_n2982_13878.n15 a_n2982_13878.n63 70.1674
R15527 a_n2982_13878.n17 a_n2982_13878.n61 70.1674
R15528 a_n2982_13878.n20 a_n2982_13878.n59 70.1674
R15529 a_n2982_13878.n120 a_n2982_13878.n59 20.9683
R15530 a_n2982_13878.n58 a_n2982_13878.n21 75.0448
R15531 a_n2982_13878.n58 a_n2982_13878.n118 11.2134
R15532 a_n2982_13878.n21 a_n2982_13878.n119 161.3
R15533 a_n2982_13878.n122 a_n2982_13878.n61 20.9683
R15534 a_n2982_13878.n60 a_n2982_13878.n18 75.0448
R15535 a_n2982_13878.n60 a_n2982_13878.n117 11.2134
R15536 a_n2982_13878.n18 a_n2982_13878.n121 161.3
R15537 a_n2982_13878.n124 a_n2982_13878.n63 20.9683
R15538 a_n2982_13878.n62 a_n2982_13878.n16 75.0448
R15539 a_n2982_13878.n62 a_n2982_13878.n116 11.2134
R15540 a_n2982_13878.n16 a_n2982_13878.n123 161.3
R15541 a_n2982_13878.n126 a_n2982_13878.n65 20.9683
R15542 a_n2982_13878.n64 a_n2982_13878.n14 75.0448
R15543 a_n2982_13878.n64 a_n2982_13878.n115 11.2134
R15544 a_n2982_13878.n14 a_n2982_13878.n125 161.3
R15545 a_n2982_13878.n7 a_n2982_13878.n72 70.1674
R15546 a_n2982_13878.n72 a_n2982_13878.n88 20.9683
R15547 a_n2982_13878.n71 a_n2982_13878.n8 74.73
R15548 a_n2982_13878.n129 a_n2982_13878.n71 11.843
R15549 a_n2982_13878.n70 a_n2982_13878.n8 80.4688
R15550 a_n2982_13878.n70 a_n2982_13878.n130 0.365327
R15551 a_n2982_13878.n9 a_n2982_13878.n69 75.0448
R15552 a_n2982_13878.n68 a_n2982_13878.n9 70.1674
R15553 a_n2982_13878.n132 a_n2982_13878.n68 20.9683
R15554 a_n2982_13878.n11 a_n2982_13878.n67 70.3058
R15555 a_n2982_13878.n67 a_n2982_13878.n86 20.6913
R15556 a_n2982_13878.n66 a_n2982_13878.n11 75.3623
R15557 a_n2982_13878.n133 a_n2982_13878.n66 10.5784
R15558 a_n2982_13878.n10 a_n2982_13878.n12 44.7878
R15559 a_n2982_13878.n35 a_n2982_13878.n143 14.1668
R15560 a_n2982_13878.n82 a_n2982_13878.n81 75.3623
R15561 a_n2982_13878.n80 a_n2982_13878.n3 70.3058
R15562 a_n2982_13878.n3 a_n2982_13878.n79 70.1674
R15563 a_n2982_13878.n79 a_n2982_13878.n84 20.9683
R15564 a_n2982_13878.n78 a_n2982_13878.n4 75.0448
R15565 a_n2982_13878.n146 a_n2982_13878.n78 11.2134
R15566 a_n2982_13878.n77 a_n2982_13878.n4 80.4688
R15567 a_n2982_13878.n6 a_n2982_13878.n76 74.73
R15568 a_n2982_13878.n75 a_n2982_13878.n6 70.1674
R15569 a_n2982_13878.n149 a_n2982_13878.n75 20.9683
R15570 a_n2982_13878.n5 a_n2982_13878.n74 70.5844
R15571 a_n2982_13878.n1 a_n2982_13878.n141 81.3764
R15572 a_n2982_13878.n2 a_n2982_13878.n137 81.3764
R15573 a_n2982_13878.n2 a_n2982_13878.n135 81.3764
R15574 a_n2982_13878.n1 a_n2982_13878.n142 80.9324
R15575 a_n2982_13878.n1 a_n2982_13878.n140 80.9324
R15576 a_n2982_13878.n0 a_n2982_13878.n139 80.9324
R15577 a_n2982_13878.n2 a_n2982_13878.n138 80.9324
R15578 a_n2982_13878.n2 a_n2982_13878.n136 80.9324
R15579 a_n2982_13878.n41 a_n2982_13878.t27 74.6477
R15580 a_n2982_13878.n36 a_n2982_13878.t49 74.6477
R15581 a_n2982_13878.n39 a_n2982_13878.t51 74.2899
R15582 a_n2982_13878.n38 a_n2982_13878.t37 74.2897
R15583 a_n2982_13878.n41 a_n2982_13878.n154 70.6783
R15584 a_n2982_13878.n40 a_n2982_13878.n153 70.6783
R15585 a_n2982_13878.n40 a_n2982_13878.n152 70.6783
R15586 a_n2982_13878.n39 a_n2982_13878.n151 70.6783
R15587 a_n2982_13878.n38 a_n2982_13878.n93 70.6783
R15588 a_n2982_13878.n37 a_n2982_13878.n92 70.6783
R15589 a_n2982_13878.n37 a_n2982_13878.n91 70.6783
R15590 a_n2982_13878.n36 a_n2982_13878.n90 70.6783
R15591 a_n2982_13878.n36 a_n2982_13878.n89 70.6783
R15592 a_n2982_13878.n155 a_n2982_13878.n41 70.6782
R15593 a_n2982_13878.n75 a_n2982_13878.n148 20.9683
R15594 a_n2982_13878.n147 a_n2982_13878.n146 48.2005
R15595 a_n2982_13878.n145 a_n2982_13878.n79 20.9683
R15596 a_n2982_13878.n143 a_n2982_13878.n85 48.2005
R15597 a_n2982_13878.n134 a_n2982_13878.n133 48.2005
R15598 a_n2982_13878.n68 a_n2982_13878.n131 20.9683
R15599 a_n2982_13878.n130 a_n2982_13878.n87 48.2005
R15600 a_n2982_13878.n128 a_n2982_13878.n72 20.9683
R15601 a_n2982_13878.n108 a_n2982_13878.n97 48.2005
R15602 a_n2982_13878.n110 a_n2982_13878.n52 20.9683
R15603 a_n2982_13878.n111 a_n2982_13878.n95 48.2005
R15604 a_n2982_13878.n113 a_n2982_13878.n56 20.9683
R15605 a_n2982_13878.n102 a_n2982_13878.n101 48.2005
R15606 a_n2982_13878.n104 a_n2982_13878.n44 20.9683
R15607 a_n2982_13878.n105 a_n2982_13878.n99 48.2005
R15608 a_n2982_13878.n107 a_n2982_13878.n48 20.9683
R15609 a_n2982_13878.n125 a_n2982_13878.n115 48.2005
R15610 a_n2982_13878.t91 a_n2982_13878.n65 533.335
R15611 a_n2982_13878.n123 a_n2982_13878.n116 48.2005
R15612 a_n2982_13878.t100 a_n2982_13878.n63 533.335
R15613 a_n2982_13878.n121 a_n2982_13878.n117 48.2005
R15614 a_n2982_13878.t85 a_n2982_13878.n61 533.335
R15615 a_n2982_13878.n119 a_n2982_13878.n118 48.2005
R15616 a_n2982_13878.t80 a_n2982_13878.n59 533.335
R15617 a_n2982_13878.n77 a_n2982_13878.n83 47.835
R15618 a_n2982_13878.n80 a_n2982_13878.n144 20.6913
R15619 a_n2982_13878.n132 a_n2982_13878.n67 21.4216
R15620 a_n2982_13878.n96 a_n2982_13878.n51 21.4216
R15621 a_n2982_13878.n100 a_n2982_13878.n43 21.4216
R15622 a_n2982_13878.n73 a_n2982_13878.t95 532.5
R15623 a_n2982_13878.t36 a_n2982_13878.n57 532.5
R15624 a_n2982_13878.t67 a_n2982_13878.n49 532.5
R15625 a_n2982_13878.n76 a_n2982_13878.n83 11.843
R15626 a_n2982_13878.n144 a_n2982_13878.n81 36.139
R15627 a_n2982_13878.n71 a_n2982_13878.n88 34.4824
R15628 a_n2982_13878.n94 a_n2982_13878.n55 34.4824
R15629 a_n2982_13878.n98 a_n2982_13878.n47 34.4824
R15630 a_n2982_13878.n78 a_n2982_13878.n84 35.3134
R15631 a_n2982_13878.n131 a_n2982_13878.n69 35.3134
R15632 a_n2982_13878.n69 a_n2982_13878.n87 11.2134
R15633 a_n2982_13878.n53 a_n2982_13878.n110 35.3134
R15634 a_n2982_13878.n111 a_n2982_13878.n53 11.2134
R15635 a_n2982_13878.n45 a_n2982_13878.n104 35.3134
R15636 a_n2982_13878.n105 a_n2982_13878.n45 11.2134
R15637 a_n2982_13878.n126 a_n2982_13878.n64 35.3134
R15638 a_n2982_13878.n124 a_n2982_13878.n62 35.3134
R15639 a_n2982_13878.n122 a_n2982_13878.n60 35.3134
R15640 a_n2982_13878.n120 a_n2982_13878.n58 35.3134
R15641 a_n2982_13878.n34 a_n2982_13878.n1 23.891
R15642 a_n2982_13878.n148 a_n2982_13878.n76 34.4824
R15643 a_n2982_13878.n81 a_n2982_13878.n85 10.5784
R15644 a_n2982_13878.n66 a_n2982_13878.n86 36.139
R15645 a_n2982_13878.n109 a_n2982_13878.n50 36.139
R15646 a_n2982_13878.n103 a_n2982_13878.n42 36.139
R15647 a_n2982_13878.n32 a_n2982_13878.n19 13.9285
R15648 a_n2982_13878.n7 a_n2982_13878.n127 13.724
R15649 a_n2982_13878.n150 a_n2982_13878.n5 12.4191
R15650 a_n2982_13878.n21 a_n2982_13878.n19 11.2486
R15651 a_n2982_13878.n127 a_n2982_13878.n13 11.2486
R15652 a_n2982_13878.n114 a_n2982_13878.n38 10.5745
R15653 a_n2982_13878.n114 a_n2982_13878.n23 8.58383
R15654 a_n2982_13878.n39 a_n2982_13878.n150 6.7311
R15655 a_n2982_13878.n127 a_n2982_13878.n114 5.3452
R15656 a_n2982_13878.n26 a_n2982_13878.n29 3.94368
R15657 a_n2982_13878.n34 a_n2982_13878.n10 3.7202
R15658 a_n2982_13878.n154 a_n2982_13878.t29 3.61217
R15659 a_n2982_13878.n154 a_n2982_13878.t57 3.61217
R15660 a_n2982_13878.n153 a_n2982_13878.t59 3.61217
R15661 a_n2982_13878.n153 a_n2982_13878.t47 3.61217
R15662 a_n2982_13878.n152 a_n2982_13878.t45 3.61217
R15663 a_n2982_13878.n152 a_n2982_13878.t35 3.61217
R15664 a_n2982_13878.n151 a_n2982_13878.t39 3.61217
R15665 a_n2982_13878.n151 a_n2982_13878.t53 3.61217
R15666 a_n2982_13878.n93 a_n2982_13878.t23 3.61217
R15667 a_n2982_13878.n93 a_n2982_13878.t19 3.61217
R15668 a_n2982_13878.n92 a_n2982_13878.t63 3.61217
R15669 a_n2982_13878.n92 a_n2982_13878.t55 3.61217
R15670 a_n2982_13878.n91 a_n2982_13878.t43 3.61217
R15671 a_n2982_13878.n91 a_n2982_13878.t33 3.61217
R15672 a_n2982_13878.n90 a_n2982_13878.t41 3.61217
R15673 a_n2982_13878.n90 a_n2982_13878.t25 3.61217
R15674 a_n2982_13878.n89 a_n2982_13878.t21 3.61217
R15675 a_n2982_13878.n89 a_n2982_13878.t61 3.61217
R15676 a_n2982_13878.t17 a_n2982_13878.n155 3.61217
R15677 a_n2982_13878.n155 a_n2982_13878.t31 3.61217
R15678 a_n2982_13878.n141 a_n2982_13878.t4 2.82907
R15679 a_n2982_13878.n141 a_n2982_13878.t7 2.82907
R15680 a_n2982_13878.n142 a_n2982_13878.t0 2.82907
R15681 a_n2982_13878.n142 a_n2982_13878.t15 2.82907
R15682 a_n2982_13878.n140 a_n2982_13878.t6 2.82907
R15683 a_n2982_13878.n140 a_n2982_13878.t13 2.82907
R15684 a_n2982_13878.n139 a_n2982_13878.t9 2.82907
R15685 a_n2982_13878.n139 a_n2982_13878.t12 2.82907
R15686 a_n2982_13878.n137 a_n2982_13878.t11 2.82907
R15687 a_n2982_13878.n137 a_n2982_13878.t10 2.82907
R15688 a_n2982_13878.n138 a_n2982_13878.t14 2.82907
R15689 a_n2982_13878.n138 a_n2982_13878.t5 2.82907
R15690 a_n2982_13878.n136 a_n2982_13878.t2 2.82907
R15691 a_n2982_13878.n136 a_n2982_13878.t1 2.82907
R15692 a_n2982_13878.n135 a_n2982_13878.t8 2.82907
R15693 a_n2982_13878.n135 a_n2982_13878.t3 2.82907
R15694 a_n2982_13878.n74 a_n2982_13878.n149 22.3251
R15695 a_n2982_13878.n35 a_n2982_13878.t26 538.698
R15696 a_n2982_13878.n12 a_n2982_13878.n134 14.1668
R15697 a_n2982_13878.n128 a_n2982_13878.n73 22.3251
R15698 a_n2982_13878.n108 a_n2982_13878.n27 14.1668
R15699 a_n2982_13878.n57 a_n2982_13878.n113 22.3251
R15700 a_n2982_13878.n102 a_n2982_13878.n33 14.1668
R15701 a_n2982_13878.n49 a_n2982_13878.n107 22.3251
R15702 a_n2982_13878.n150 a_n2982_13878.n19 1.30542
R15703 a_n2982_13878.n16 a_n2982_13878.n17 1.04595
R15704 a_n2982_13878.n77 a_n2982_13878.n147 0.365327
R15705 a_n2982_13878.n145 a_n2982_13878.n80 21.4216
R15706 a_n2982_13878.n70 a_n2982_13878.n129 47.835
R15707 a_n2982_13878.n112 a_n2982_13878.n54 47.835
R15708 a_n2982_13878.n106 a_n2982_13878.n46 47.835
R15709 a_n2982_13878.n0 a_n2982_13878.n2 31.7919
R15710 a_n2982_13878.n29 a_n2982_13878.n28 1.13686
R15711 a_n2982_13878.n23 a_n2982_13878.n22 1.13686
R15712 a_n2982_13878.n8 a_n2982_13878.n7 1.13686
R15713 a_n2982_13878.n40 a_n2982_13878.n39 1.07378
R15714 a_n2982_13878.n37 a_n2982_13878.n36 1.07378
R15715 a_n2982_13878.n1 a_n2982_13878.n0 0.888431
R15716 a_n2982_13878.n31 a_n2982_13878.n32 0.758076
R15717 a_n2982_13878.n30 a_n2982_13878.n31 0.758076
R15718 a_n2982_13878.n28 a_n2982_13878.n30 0.758076
R15719 a_n2982_13878.n25 a_n2982_13878.n26 0.758076
R15720 a_n2982_13878.n24 a_n2982_13878.n25 0.758076
R15721 a_n2982_13878.n22 a_n2982_13878.n24 0.758076
R15722 a_n2982_13878.n21 a_n2982_13878.n20 0.758076
R15723 a_n2982_13878.n18 a_n2982_13878.n17 0.758076
R15724 a_n2982_13878.n16 a_n2982_13878.n15 0.758076
R15725 a_n2982_13878.n14 a_n2982_13878.n13 0.758076
R15726 a_n2982_13878.n11 a_n2982_13878.n10 0.758076
R15727 a_n2982_13878.n11 a_n2982_13878.n9 0.758076
R15728 a_n2982_13878.n9 a_n2982_13878.n8 0.758076
R15729 a_n2982_13878.n6 a_n2982_13878.n4 0.758076
R15730 a_n2982_13878.n4 a_n2982_13878.n3 0.758076
R15731 a_n2982_13878.n82 a_n2982_13878.n3 0.758076
R15732 a_n2982_13878.n82 a_n2982_13878.n34 0.754288
R15733 a_n2982_13878.n41 a_n2982_13878.n40 0.716017
R15734 a_n2982_13878.n38 a_n2982_13878.n37 0.716017
R15735 a_n2982_13878.n18 a_n2982_13878.n20 0.67853
R15736 a_n2982_13878.n14 a_n2982_13878.n15 0.67853
R15737 a_n2982_13878.n6 a_n2982_13878.n5 0.568682
R15738 a_n2804_13878.n2 a_n2804_13878.n0 98.9633
R15739 a_n2804_13878.n5 a_n2804_13878.n3 98.7517
R15740 a_n2804_13878.n25 a_n2804_13878.n24 98.6055
R15741 a_n2804_13878.n27 a_n2804_13878.n26 98.6055
R15742 a_n2804_13878.n2 a_n2804_13878.n1 98.6055
R15743 a_n2804_13878.n13 a_n2804_13878.n12 98.6055
R15744 a_n2804_13878.n11 a_n2804_13878.n10 98.6055
R15745 a_n2804_13878.n9 a_n2804_13878.n8 98.6055
R15746 a_n2804_13878.n7 a_n2804_13878.n6 98.6055
R15747 a_n2804_13878.n5 a_n2804_13878.n4 98.6055
R15748 a_n2804_13878.n29 a_n2804_13878.n28 98.6054
R15749 a_n2804_13878.n23 a_n2804_13878.n22 98.6054
R15750 a_n2804_13878.n15 a_n2804_13878.t6 74.6477
R15751 a_n2804_13878.n20 a_n2804_13878.t7 74.2899
R15752 a_n2804_13878.n17 a_n2804_13878.t5 74.2899
R15753 a_n2804_13878.n16 a_n2804_13878.t2 74.2899
R15754 a_n2804_13878.n19 a_n2804_13878.n18 70.6783
R15755 a_n2804_13878.n15 a_n2804_13878.n14 70.6783
R15756 a_n2804_13878.n21 a_n2804_13878.n13 15.7159
R15757 a_n2804_13878.n23 a_n2804_13878.n21 12.6495
R15758 a_n2804_13878.n21 a_n2804_13878.n20 8.38735
R15759 a_n2804_13878.n22 a_n2804_13878.t15 3.61217
R15760 a_n2804_13878.n22 a_n2804_13878.t24 3.61217
R15761 a_n2804_13878.n24 a_n2804_13878.t28 3.61217
R15762 a_n2804_13878.n24 a_n2804_13878.t14 3.61217
R15763 a_n2804_13878.n26 a_n2804_13878.t18 3.61217
R15764 a_n2804_13878.n26 a_n2804_13878.t19 3.61217
R15765 a_n2804_13878.n1 a_n2804_13878.t8 3.61217
R15766 a_n2804_13878.n1 a_n2804_13878.t20 3.61217
R15767 a_n2804_13878.n0 a_n2804_13878.t25 3.61217
R15768 a_n2804_13878.n0 a_n2804_13878.t31 3.61217
R15769 a_n2804_13878.n18 a_n2804_13878.t4 3.61217
R15770 a_n2804_13878.n18 a_n2804_13878.t0 3.61217
R15771 a_n2804_13878.n14 a_n2804_13878.t1 3.61217
R15772 a_n2804_13878.n14 a_n2804_13878.t3 3.61217
R15773 a_n2804_13878.n12 a_n2804_13878.t21 3.61217
R15774 a_n2804_13878.n12 a_n2804_13878.t9 3.61217
R15775 a_n2804_13878.n10 a_n2804_13878.t26 3.61217
R15776 a_n2804_13878.n10 a_n2804_13878.t11 3.61217
R15777 a_n2804_13878.n8 a_n2804_13878.t10 3.61217
R15778 a_n2804_13878.n8 a_n2804_13878.t13 3.61217
R15779 a_n2804_13878.n6 a_n2804_13878.t23 3.61217
R15780 a_n2804_13878.n6 a_n2804_13878.t16 3.61217
R15781 a_n2804_13878.n4 a_n2804_13878.t27 3.61217
R15782 a_n2804_13878.n4 a_n2804_13878.t17 3.61217
R15783 a_n2804_13878.n3 a_n2804_13878.t12 3.61217
R15784 a_n2804_13878.n3 a_n2804_13878.t22 3.61217
R15785 a_n2804_13878.n29 a_n2804_13878.t29 3.61217
R15786 a_n2804_13878.t30 a_n2804_13878.n29 3.61217
R15787 a_n2804_13878.n16 a_n2804_13878.n15 0.358259
R15788 a_n2804_13878.n19 a_n2804_13878.n17 0.358259
R15789 a_n2804_13878.n20 a_n2804_13878.n19 0.358259
R15790 a_n2804_13878.n28 a_n2804_13878.n2 0.358259
R15791 a_n2804_13878.n28 a_n2804_13878.n27 0.358259
R15792 a_n2804_13878.n27 a_n2804_13878.n25 0.358259
R15793 a_n2804_13878.n25 a_n2804_13878.n23 0.358259
R15794 a_n2804_13878.n7 a_n2804_13878.n5 0.146627
R15795 a_n2804_13878.n9 a_n2804_13878.n7 0.146627
R15796 a_n2804_13878.n11 a_n2804_13878.n9 0.146627
R15797 a_n2804_13878.n13 a_n2804_13878.n11 0.146627
R15798 a_n2804_13878.n17 a_n2804_13878.n16 0.101793
R15799 vdd.n327 vdd.n291 756.745
R15800 vdd.n268 vdd.n232 756.745
R15801 vdd.n225 vdd.n189 756.745
R15802 vdd.n166 vdd.n130 756.745
R15803 vdd.n124 vdd.n88 756.745
R15804 vdd.n65 vdd.n29 756.745
R15805 vdd.n2201 vdd.n2165 756.745
R15806 vdd.n2260 vdd.n2224 756.745
R15807 vdd.n2099 vdd.n2063 756.745
R15808 vdd.n2158 vdd.n2122 756.745
R15809 vdd.n1998 vdd.n1962 756.745
R15810 vdd.n2057 vdd.n2021 756.745
R15811 vdd.n1315 vdd.t12 640.208
R15812 vdd.n1010 vdd.t53 640.208
R15813 vdd.n1319 vdd.t50 640.208
R15814 vdd.n1001 vdd.t75 640.208
R15815 vdd.n896 vdd.t37 640.208
R15816 vdd.n2823 vdd.t68 640.208
R15817 vdd.n832 vdd.t30 640.208
R15818 vdd.n2820 vdd.t60 640.208
R15819 vdd.n799 vdd.t8 640.208
R15820 vdd.n1071 vdd.t64 640.208
R15821 vdd.n1772 vdd.t78 592.009
R15822 vdd.n1810 vdd.t71 592.009
R15823 vdd.n1706 vdd.t81 592.009
R15824 vdd.n2362 vdd.t41 592.009
R15825 vdd.n1248 vdd.t16 592.009
R15826 vdd.n1208 vdd.t24 592.009
R15827 vdd.n426 vdd.t47 592.009
R15828 vdd.n440 vdd.t20 592.009
R15829 vdd.n452 vdd.t27 592.009
R15830 vdd.n768 vdd.t44 592.009
R15831 vdd.n3456 vdd.t57 592.009
R15832 vdd.n688 vdd.t33 592.009
R15833 vdd.n328 vdd.n327 585
R15834 vdd.n326 vdd.n293 585
R15835 vdd.n325 vdd.n324 585
R15836 vdd.n296 vdd.n294 585
R15837 vdd.n319 vdd.n318 585
R15838 vdd.n317 vdd.n316 585
R15839 vdd.n300 vdd.n299 585
R15840 vdd.n311 vdd.n310 585
R15841 vdd.n309 vdd.n308 585
R15842 vdd.n304 vdd.n303 585
R15843 vdd.n269 vdd.n268 585
R15844 vdd.n267 vdd.n234 585
R15845 vdd.n266 vdd.n265 585
R15846 vdd.n237 vdd.n235 585
R15847 vdd.n260 vdd.n259 585
R15848 vdd.n258 vdd.n257 585
R15849 vdd.n241 vdd.n240 585
R15850 vdd.n252 vdd.n251 585
R15851 vdd.n250 vdd.n249 585
R15852 vdd.n245 vdd.n244 585
R15853 vdd.n226 vdd.n225 585
R15854 vdd.n224 vdd.n191 585
R15855 vdd.n223 vdd.n222 585
R15856 vdd.n194 vdd.n192 585
R15857 vdd.n217 vdd.n216 585
R15858 vdd.n215 vdd.n214 585
R15859 vdd.n198 vdd.n197 585
R15860 vdd.n209 vdd.n208 585
R15861 vdd.n207 vdd.n206 585
R15862 vdd.n202 vdd.n201 585
R15863 vdd.n167 vdd.n166 585
R15864 vdd.n165 vdd.n132 585
R15865 vdd.n164 vdd.n163 585
R15866 vdd.n135 vdd.n133 585
R15867 vdd.n158 vdd.n157 585
R15868 vdd.n156 vdd.n155 585
R15869 vdd.n139 vdd.n138 585
R15870 vdd.n150 vdd.n149 585
R15871 vdd.n148 vdd.n147 585
R15872 vdd.n143 vdd.n142 585
R15873 vdd.n125 vdd.n124 585
R15874 vdd.n123 vdd.n90 585
R15875 vdd.n122 vdd.n121 585
R15876 vdd.n93 vdd.n91 585
R15877 vdd.n116 vdd.n115 585
R15878 vdd.n114 vdd.n113 585
R15879 vdd.n97 vdd.n96 585
R15880 vdd.n108 vdd.n107 585
R15881 vdd.n106 vdd.n105 585
R15882 vdd.n101 vdd.n100 585
R15883 vdd.n66 vdd.n65 585
R15884 vdd.n64 vdd.n31 585
R15885 vdd.n63 vdd.n62 585
R15886 vdd.n34 vdd.n32 585
R15887 vdd.n57 vdd.n56 585
R15888 vdd.n55 vdd.n54 585
R15889 vdd.n38 vdd.n37 585
R15890 vdd.n49 vdd.n48 585
R15891 vdd.n47 vdd.n46 585
R15892 vdd.n42 vdd.n41 585
R15893 vdd.n2202 vdd.n2201 585
R15894 vdd.n2200 vdd.n2167 585
R15895 vdd.n2199 vdd.n2198 585
R15896 vdd.n2170 vdd.n2168 585
R15897 vdd.n2193 vdd.n2192 585
R15898 vdd.n2191 vdd.n2190 585
R15899 vdd.n2174 vdd.n2173 585
R15900 vdd.n2185 vdd.n2184 585
R15901 vdd.n2183 vdd.n2182 585
R15902 vdd.n2178 vdd.n2177 585
R15903 vdd.n2261 vdd.n2260 585
R15904 vdd.n2259 vdd.n2226 585
R15905 vdd.n2258 vdd.n2257 585
R15906 vdd.n2229 vdd.n2227 585
R15907 vdd.n2252 vdd.n2251 585
R15908 vdd.n2250 vdd.n2249 585
R15909 vdd.n2233 vdd.n2232 585
R15910 vdd.n2244 vdd.n2243 585
R15911 vdd.n2242 vdd.n2241 585
R15912 vdd.n2237 vdd.n2236 585
R15913 vdd.n2100 vdd.n2099 585
R15914 vdd.n2098 vdd.n2065 585
R15915 vdd.n2097 vdd.n2096 585
R15916 vdd.n2068 vdd.n2066 585
R15917 vdd.n2091 vdd.n2090 585
R15918 vdd.n2089 vdd.n2088 585
R15919 vdd.n2072 vdd.n2071 585
R15920 vdd.n2083 vdd.n2082 585
R15921 vdd.n2081 vdd.n2080 585
R15922 vdd.n2076 vdd.n2075 585
R15923 vdd.n2159 vdd.n2158 585
R15924 vdd.n2157 vdd.n2124 585
R15925 vdd.n2156 vdd.n2155 585
R15926 vdd.n2127 vdd.n2125 585
R15927 vdd.n2150 vdd.n2149 585
R15928 vdd.n2148 vdd.n2147 585
R15929 vdd.n2131 vdd.n2130 585
R15930 vdd.n2142 vdd.n2141 585
R15931 vdd.n2140 vdd.n2139 585
R15932 vdd.n2135 vdd.n2134 585
R15933 vdd.n1999 vdd.n1998 585
R15934 vdd.n1997 vdd.n1964 585
R15935 vdd.n1996 vdd.n1995 585
R15936 vdd.n1967 vdd.n1965 585
R15937 vdd.n1990 vdd.n1989 585
R15938 vdd.n1988 vdd.n1987 585
R15939 vdd.n1971 vdd.n1970 585
R15940 vdd.n1982 vdd.n1981 585
R15941 vdd.n1980 vdd.n1979 585
R15942 vdd.n1975 vdd.n1974 585
R15943 vdd.n2058 vdd.n2057 585
R15944 vdd.n2056 vdd.n2023 585
R15945 vdd.n2055 vdd.n2054 585
R15946 vdd.n2026 vdd.n2024 585
R15947 vdd.n2049 vdd.n2048 585
R15948 vdd.n2047 vdd.n2046 585
R15949 vdd.n2030 vdd.n2029 585
R15950 vdd.n2041 vdd.n2040 585
R15951 vdd.n2039 vdd.n2038 585
R15952 vdd.n2034 vdd.n2033 585
R15953 vdd.n3628 vdd.n392 509.269
R15954 vdd.n3624 vdd.n393 509.269
R15955 vdd.n3496 vdd.n685 509.269
R15956 vdd.n3493 vdd.n684 509.269
R15957 vdd.n2357 vdd.n1530 509.269
R15958 vdd.n2360 vdd.n2359 509.269
R15959 vdd.n1679 vdd.n1643 509.269
R15960 vdd.n1875 vdd.n1644 509.269
R15961 vdd.n305 vdd.t124 329.043
R15962 vdd.n246 vdd.t240 329.043
R15963 vdd.n203 vdd.t105 329.043
R15964 vdd.n144 vdd.t229 329.043
R15965 vdd.n102 vdd.t210 329.043
R15966 vdd.n43 vdd.t170 329.043
R15967 vdd.n2179 vdd.t151 329.043
R15968 vdd.n2238 vdd.t193 329.043
R15969 vdd.n2077 vdd.t131 329.043
R15970 vdd.n2136 vdd.t176 329.043
R15971 vdd.n1976 vdd.t171 329.043
R15972 vdd.n2035 vdd.t212 329.043
R15973 vdd.n1772 vdd.t80 319.788
R15974 vdd.n1810 vdd.t74 319.788
R15975 vdd.n1706 vdd.t83 319.788
R15976 vdd.n2362 vdd.t42 319.788
R15977 vdd.n1248 vdd.t18 319.788
R15978 vdd.n1208 vdd.t25 319.788
R15979 vdd.n426 vdd.t48 319.788
R15980 vdd.n440 vdd.t22 319.788
R15981 vdd.n452 vdd.t28 319.788
R15982 vdd.n768 vdd.t46 319.788
R15983 vdd.n3456 vdd.t59 319.788
R15984 vdd.n688 vdd.t36 319.788
R15985 vdd.n1773 vdd.t79 303.69
R15986 vdd.n1811 vdd.t73 303.69
R15987 vdd.n1707 vdd.t82 303.69
R15988 vdd.n2363 vdd.t43 303.69
R15989 vdd.n1249 vdd.t19 303.69
R15990 vdd.n1209 vdd.t26 303.69
R15991 vdd.n427 vdd.t49 303.69
R15992 vdd.n441 vdd.t23 303.69
R15993 vdd.n453 vdd.t29 303.69
R15994 vdd.n769 vdd.t45 303.69
R15995 vdd.n3457 vdd.t58 303.69
R15996 vdd.n689 vdd.t35 303.69
R15997 vdd.n3090 vdd.n960 279.512
R15998 vdd.n3330 vdd.n809 279.512
R15999 vdd.n3267 vdd.n806 279.512
R16000 vdd.n3022 vdd.n3021 279.512
R16001 vdd.n2783 vdd.n998 279.512
R16002 vdd.n2714 vdd.n2713 279.512
R16003 vdd.n1355 vdd.n1354 279.512
R16004 vdd.n2508 vdd.n1138 279.512
R16005 vdd.n3246 vdd.n807 279.512
R16006 vdd.n3333 vdd.n3332 279.512
R16007 vdd.n2895 vdd.n2818 279.512
R16008 vdd.n2826 vdd.n956 279.512
R16009 vdd.n2711 vdd.n1008 279.512
R16010 vdd.n1006 vdd.n980 279.512
R16011 vdd.n1480 vdd.n1175 279.512
R16012 vdd.n1280 vdd.n1133 279.512
R16013 vdd.n2506 vdd.n1141 254.619
R16014 vdd.n3495 vdd.n692 254.619
R16015 vdd.n3248 vdd.n807 185
R16016 vdd.n3331 vdd.n807 185
R16017 vdd.n3250 vdd.n3249 185
R16018 vdd.n3249 vdd.n805 185
R16019 vdd.n3251 vdd.n839 185
R16020 vdd.n3261 vdd.n839 185
R16021 vdd.n3252 vdd.n848 185
R16022 vdd.n848 vdd.n846 185
R16023 vdd.n3254 vdd.n3253 185
R16024 vdd.n3255 vdd.n3254 185
R16025 vdd.n3207 vdd.n847 185
R16026 vdd.n847 vdd.n843 185
R16027 vdd.n3206 vdd.n3205 185
R16028 vdd.n3205 vdd.n3204 185
R16029 vdd.n850 vdd.n849 185
R16030 vdd.n851 vdd.n850 185
R16031 vdd.n3197 vdd.n3196 185
R16032 vdd.n3198 vdd.n3197 185
R16033 vdd.n3195 vdd.n859 185
R16034 vdd.n864 vdd.n859 185
R16035 vdd.n3194 vdd.n3193 185
R16036 vdd.n3193 vdd.n3192 185
R16037 vdd.n861 vdd.n860 185
R16038 vdd.n870 vdd.n861 185
R16039 vdd.n3185 vdd.n3184 185
R16040 vdd.n3186 vdd.n3185 185
R16041 vdd.n3183 vdd.n871 185
R16042 vdd.n877 vdd.n871 185
R16043 vdd.n3182 vdd.n3181 185
R16044 vdd.n3181 vdd.n3180 185
R16045 vdd.n873 vdd.n872 185
R16046 vdd.n874 vdd.n873 185
R16047 vdd.n3173 vdd.n3172 185
R16048 vdd.n3174 vdd.n3173 185
R16049 vdd.n3171 vdd.n884 185
R16050 vdd.n884 vdd.n881 185
R16051 vdd.n3170 vdd.n3169 185
R16052 vdd.n3169 vdd.n3168 185
R16053 vdd.n886 vdd.n885 185
R16054 vdd.n887 vdd.n886 185
R16055 vdd.n3161 vdd.n3160 185
R16056 vdd.n3162 vdd.n3161 185
R16057 vdd.n3159 vdd.n895 185
R16058 vdd.n901 vdd.n895 185
R16059 vdd.n3158 vdd.n3157 185
R16060 vdd.n3157 vdd.n3156 185
R16061 vdd.n3147 vdd.n898 185
R16062 vdd.n908 vdd.n898 185
R16063 vdd.n3149 vdd.n3148 185
R16064 vdd.n3150 vdd.n3149 185
R16065 vdd.n3146 vdd.n909 185
R16066 vdd.n909 vdd.n905 185
R16067 vdd.n3145 vdd.n3144 185
R16068 vdd.n3144 vdd.n3143 185
R16069 vdd.n911 vdd.n910 185
R16070 vdd.n912 vdd.n911 185
R16071 vdd.n3136 vdd.n3135 185
R16072 vdd.n3137 vdd.n3136 185
R16073 vdd.n3134 vdd.n920 185
R16074 vdd.n925 vdd.n920 185
R16075 vdd.n3133 vdd.n3132 185
R16076 vdd.n3132 vdd.n3131 185
R16077 vdd.n922 vdd.n921 185
R16078 vdd.n931 vdd.n922 185
R16079 vdd.n3124 vdd.n3123 185
R16080 vdd.n3125 vdd.n3124 185
R16081 vdd.n3122 vdd.n932 185
R16082 vdd.n2998 vdd.n932 185
R16083 vdd.n3121 vdd.n3120 185
R16084 vdd.n3120 vdd.n3119 185
R16085 vdd.n934 vdd.n933 185
R16086 vdd.n3004 vdd.n934 185
R16087 vdd.n3112 vdd.n3111 185
R16088 vdd.n3113 vdd.n3112 185
R16089 vdd.n3110 vdd.n943 185
R16090 vdd.n943 vdd.n940 185
R16091 vdd.n3109 vdd.n3108 185
R16092 vdd.n3108 vdd.n3107 185
R16093 vdd.n945 vdd.n944 185
R16094 vdd.n946 vdd.n945 185
R16095 vdd.n3100 vdd.n3099 185
R16096 vdd.n3101 vdd.n3100 185
R16097 vdd.n3098 vdd.n954 185
R16098 vdd.n3016 vdd.n954 185
R16099 vdd.n3097 vdd.n3096 185
R16100 vdd.n3096 vdd.n3095 185
R16101 vdd.n956 vdd.n955 185
R16102 vdd.n957 vdd.n956 185
R16103 vdd.n2827 vdd.n2826 185
R16104 vdd.n2829 vdd.n2828 185
R16105 vdd.n2831 vdd.n2830 185
R16106 vdd.n2833 vdd.n2832 185
R16107 vdd.n2835 vdd.n2834 185
R16108 vdd.n2837 vdd.n2836 185
R16109 vdd.n2839 vdd.n2838 185
R16110 vdd.n2841 vdd.n2840 185
R16111 vdd.n2843 vdd.n2842 185
R16112 vdd.n2845 vdd.n2844 185
R16113 vdd.n2847 vdd.n2846 185
R16114 vdd.n2849 vdd.n2848 185
R16115 vdd.n2851 vdd.n2850 185
R16116 vdd.n2853 vdd.n2852 185
R16117 vdd.n2855 vdd.n2854 185
R16118 vdd.n2857 vdd.n2856 185
R16119 vdd.n2859 vdd.n2858 185
R16120 vdd.n2861 vdd.n2860 185
R16121 vdd.n2863 vdd.n2862 185
R16122 vdd.n2865 vdd.n2864 185
R16123 vdd.n2867 vdd.n2866 185
R16124 vdd.n2869 vdd.n2868 185
R16125 vdd.n2871 vdd.n2870 185
R16126 vdd.n2873 vdd.n2872 185
R16127 vdd.n2875 vdd.n2874 185
R16128 vdd.n2877 vdd.n2876 185
R16129 vdd.n2879 vdd.n2878 185
R16130 vdd.n2881 vdd.n2880 185
R16131 vdd.n2883 vdd.n2882 185
R16132 vdd.n2885 vdd.n2884 185
R16133 vdd.n2887 vdd.n2886 185
R16134 vdd.n2889 vdd.n2888 185
R16135 vdd.n2891 vdd.n2890 185
R16136 vdd.n2893 vdd.n2892 185
R16137 vdd.n2894 vdd.n2818 185
R16138 vdd.n3088 vdd.n2818 185
R16139 vdd.n3334 vdd.n3333 185
R16140 vdd.n3335 vdd.n798 185
R16141 vdd.n3337 vdd.n3336 185
R16142 vdd.n3339 vdd.n796 185
R16143 vdd.n3341 vdd.n3340 185
R16144 vdd.n3342 vdd.n795 185
R16145 vdd.n3344 vdd.n3343 185
R16146 vdd.n3346 vdd.n793 185
R16147 vdd.n3348 vdd.n3347 185
R16148 vdd.n3349 vdd.n792 185
R16149 vdd.n3351 vdd.n3350 185
R16150 vdd.n3353 vdd.n790 185
R16151 vdd.n3355 vdd.n3354 185
R16152 vdd.n3356 vdd.n789 185
R16153 vdd.n3358 vdd.n3357 185
R16154 vdd.n3360 vdd.n788 185
R16155 vdd.n3361 vdd.n786 185
R16156 vdd.n3364 vdd.n3363 185
R16157 vdd.n787 vdd.n785 185
R16158 vdd.n3220 vdd.n3219 185
R16159 vdd.n3222 vdd.n3221 185
R16160 vdd.n3224 vdd.n3216 185
R16161 vdd.n3226 vdd.n3225 185
R16162 vdd.n3227 vdd.n3215 185
R16163 vdd.n3229 vdd.n3228 185
R16164 vdd.n3231 vdd.n3213 185
R16165 vdd.n3233 vdd.n3232 185
R16166 vdd.n3234 vdd.n3212 185
R16167 vdd.n3236 vdd.n3235 185
R16168 vdd.n3238 vdd.n3210 185
R16169 vdd.n3240 vdd.n3239 185
R16170 vdd.n3241 vdd.n3209 185
R16171 vdd.n3243 vdd.n3242 185
R16172 vdd.n3245 vdd.n3208 185
R16173 vdd.n3247 vdd.n3246 185
R16174 vdd.n3246 vdd.n692 185
R16175 vdd.n3332 vdd.n802 185
R16176 vdd.n3332 vdd.n3331 185
R16177 vdd.n2949 vdd.n804 185
R16178 vdd.n805 vdd.n804 185
R16179 vdd.n2950 vdd.n838 185
R16180 vdd.n3261 vdd.n838 185
R16181 vdd.n2952 vdd.n2951 185
R16182 vdd.n2951 vdd.n846 185
R16183 vdd.n2953 vdd.n845 185
R16184 vdd.n3255 vdd.n845 185
R16185 vdd.n2955 vdd.n2954 185
R16186 vdd.n2954 vdd.n843 185
R16187 vdd.n2956 vdd.n853 185
R16188 vdd.n3204 vdd.n853 185
R16189 vdd.n2958 vdd.n2957 185
R16190 vdd.n2957 vdd.n851 185
R16191 vdd.n2959 vdd.n858 185
R16192 vdd.n3198 vdd.n858 185
R16193 vdd.n2961 vdd.n2960 185
R16194 vdd.n2960 vdd.n864 185
R16195 vdd.n2962 vdd.n863 185
R16196 vdd.n3192 vdd.n863 185
R16197 vdd.n2964 vdd.n2963 185
R16198 vdd.n2963 vdd.n870 185
R16199 vdd.n2965 vdd.n869 185
R16200 vdd.n3186 vdd.n869 185
R16201 vdd.n2967 vdd.n2966 185
R16202 vdd.n2966 vdd.n877 185
R16203 vdd.n2968 vdd.n876 185
R16204 vdd.n3180 vdd.n876 185
R16205 vdd.n2970 vdd.n2969 185
R16206 vdd.n2969 vdd.n874 185
R16207 vdd.n2971 vdd.n883 185
R16208 vdd.n3174 vdd.n883 185
R16209 vdd.n2973 vdd.n2972 185
R16210 vdd.n2972 vdd.n881 185
R16211 vdd.n2974 vdd.n889 185
R16212 vdd.n3168 vdd.n889 185
R16213 vdd.n2976 vdd.n2975 185
R16214 vdd.n2975 vdd.n887 185
R16215 vdd.n2977 vdd.n894 185
R16216 vdd.n3162 vdd.n894 185
R16217 vdd.n2979 vdd.n2978 185
R16218 vdd.n2978 vdd.n901 185
R16219 vdd.n2980 vdd.n900 185
R16220 vdd.n3156 vdd.n900 185
R16221 vdd.n2982 vdd.n2981 185
R16222 vdd.n2981 vdd.n908 185
R16223 vdd.n2983 vdd.n907 185
R16224 vdd.n3150 vdd.n907 185
R16225 vdd.n2985 vdd.n2984 185
R16226 vdd.n2984 vdd.n905 185
R16227 vdd.n2986 vdd.n914 185
R16228 vdd.n3143 vdd.n914 185
R16229 vdd.n2988 vdd.n2987 185
R16230 vdd.n2987 vdd.n912 185
R16231 vdd.n2989 vdd.n919 185
R16232 vdd.n3137 vdd.n919 185
R16233 vdd.n2991 vdd.n2990 185
R16234 vdd.n2990 vdd.n925 185
R16235 vdd.n2992 vdd.n924 185
R16236 vdd.n3131 vdd.n924 185
R16237 vdd.n2994 vdd.n2993 185
R16238 vdd.n2993 vdd.n931 185
R16239 vdd.n2995 vdd.n930 185
R16240 vdd.n3125 vdd.n930 185
R16241 vdd.n2997 vdd.n2996 185
R16242 vdd.n2998 vdd.n2997 185
R16243 vdd.n2898 vdd.n936 185
R16244 vdd.n3119 vdd.n936 185
R16245 vdd.n3006 vdd.n3005 185
R16246 vdd.n3005 vdd.n3004 185
R16247 vdd.n3007 vdd.n942 185
R16248 vdd.n3113 vdd.n942 185
R16249 vdd.n3009 vdd.n3008 185
R16250 vdd.n3008 vdd.n940 185
R16251 vdd.n3010 vdd.n948 185
R16252 vdd.n3107 vdd.n948 185
R16253 vdd.n3012 vdd.n3011 185
R16254 vdd.n3011 vdd.n946 185
R16255 vdd.n3013 vdd.n953 185
R16256 vdd.n3101 vdd.n953 185
R16257 vdd.n3015 vdd.n3014 185
R16258 vdd.n3016 vdd.n3015 185
R16259 vdd.n2897 vdd.n959 185
R16260 vdd.n3095 vdd.n959 185
R16261 vdd.n2896 vdd.n2895 185
R16262 vdd.n2895 vdd.n957 185
R16263 vdd.n2357 vdd.n2356 185
R16264 vdd.n2358 vdd.n2357 185
R16265 vdd.n1531 vdd.n1529 185
R16266 vdd.n2349 vdd.n1529 185
R16267 vdd.n2352 vdd.n2351 185
R16268 vdd.n2351 vdd.n2350 185
R16269 vdd.n1534 vdd.n1533 185
R16270 vdd.n1535 vdd.n1534 185
R16271 vdd.n2338 vdd.n2337 185
R16272 vdd.n2339 vdd.n2338 185
R16273 vdd.n1543 vdd.n1542 185
R16274 vdd.n2330 vdd.n1542 185
R16275 vdd.n2333 vdd.n2332 185
R16276 vdd.n2332 vdd.n2331 185
R16277 vdd.n1546 vdd.n1545 185
R16278 vdd.n1553 vdd.n1546 185
R16279 vdd.n2321 vdd.n2320 185
R16280 vdd.n2322 vdd.n2321 185
R16281 vdd.n1555 vdd.n1554 185
R16282 vdd.n1554 vdd.n1552 185
R16283 vdd.n2316 vdd.n2315 185
R16284 vdd.n2315 vdd.n2314 185
R16285 vdd.n1558 vdd.n1557 185
R16286 vdd.n1559 vdd.n1558 185
R16287 vdd.n2305 vdd.n2304 185
R16288 vdd.n2306 vdd.n2305 185
R16289 vdd.n1566 vdd.n1565 185
R16290 vdd.n2297 vdd.n1565 185
R16291 vdd.n2300 vdd.n2299 185
R16292 vdd.n2299 vdd.n2298 185
R16293 vdd.n1569 vdd.n1568 185
R16294 vdd.n1575 vdd.n1569 185
R16295 vdd.n2288 vdd.n2287 185
R16296 vdd.n2289 vdd.n2288 185
R16297 vdd.n1577 vdd.n1576 185
R16298 vdd.n2280 vdd.n1576 185
R16299 vdd.n2283 vdd.n2282 185
R16300 vdd.n2282 vdd.n2281 185
R16301 vdd.n1580 vdd.n1579 185
R16302 vdd.n1581 vdd.n1580 185
R16303 vdd.n2271 vdd.n2270 185
R16304 vdd.n2272 vdd.n2271 185
R16305 vdd.n1589 vdd.n1588 185
R16306 vdd.n1588 vdd.n1587 185
R16307 vdd.n1959 vdd.n1958 185
R16308 vdd.n1958 vdd.n1957 185
R16309 vdd.n1592 vdd.n1591 185
R16310 vdd.n1598 vdd.n1592 185
R16311 vdd.n1948 vdd.n1947 185
R16312 vdd.n1949 vdd.n1948 185
R16313 vdd.n1600 vdd.n1599 185
R16314 vdd.n1940 vdd.n1599 185
R16315 vdd.n1943 vdd.n1942 185
R16316 vdd.n1942 vdd.n1941 185
R16317 vdd.n1603 vdd.n1602 185
R16318 vdd.n1610 vdd.n1603 185
R16319 vdd.n1931 vdd.n1930 185
R16320 vdd.n1932 vdd.n1931 185
R16321 vdd.n1612 vdd.n1611 185
R16322 vdd.n1611 vdd.n1609 185
R16323 vdd.n1926 vdd.n1925 185
R16324 vdd.n1925 vdd.n1924 185
R16325 vdd.n1615 vdd.n1614 185
R16326 vdd.n1616 vdd.n1615 185
R16327 vdd.n1915 vdd.n1914 185
R16328 vdd.n1916 vdd.n1915 185
R16329 vdd.n1623 vdd.n1622 185
R16330 vdd.n1907 vdd.n1622 185
R16331 vdd.n1910 vdd.n1909 185
R16332 vdd.n1909 vdd.n1908 185
R16333 vdd.n1626 vdd.n1625 185
R16334 vdd.n1632 vdd.n1626 185
R16335 vdd.n1898 vdd.n1897 185
R16336 vdd.n1899 vdd.n1898 185
R16337 vdd.n1634 vdd.n1633 185
R16338 vdd.n1890 vdd.n1633 185
R16339 vdd.n1893 vdd.n1892 185
R16340 vdd.n1892 vdd.n1891 185
R16341 vdd.n1637 vdd.n1636 185
R16342 vdd.n1638 vdd.n1637 185
R16343 vdd.n1881 vdd.n1880 185
R16344 vdd.n1882 vdd.n1881 185
R16345 vdd.n1645 vdd.n1644 185
R16346 vdd.n1680 vdd.n1644 185
R16347 vdd.n1876 vdd.n1875 185
R16348 vdd.n1648 vdd.n1647 185
R16349 vdd.n1872 vdd.n1871 185
R16350 vdd.n1873 vdd.n1872 185
R16351 vdd.n1682 vdd.n1681 185
R16352 vdd.n1867 vdd.n1684 185
R16353 vdd.n1866 vdd.n1685 185
R16354 vdd.n1865 vdd.n1686 185
R16355 vdd.n1688 vdd.n1687 185
R16356 vdd.n1861 vdd.n1690 185
R16357 vdd.n1860 vdd.n1691 185
R16358 vdd.n1859 vdd.n1692 185
R16359 vdd.n1694 vdd.n1693 185
R16360 vdd.n1855 vdd.n1696 185
R16361 vdd.n1854 vdd.n1697 185
R16362 vdd.n1853 vdd.n1698 185
R16363 vdd.n1700 vdd.n1699 185
R16364 vdd.n1849 vdd.n1702 185
R16365 vdd.n1848 vdd.n1703 185
R16366 vdd.n1847 vdd.n1704 185
R16367 vdd.n1708 vdd.n1705 185
R16368 vdd.n1843 vdd.n1710 185
R16369 vdd.n1842 vdd.n1711 185
R16370 vdd.n1841 vdd.n1712 185
R16371 vdd.n1714 vdd.n1713 185
R16372 vdd.n1837 vdd.n1716 185
R16373 vdd.n1836 vdd.n1717 185
R16374 vdd.n1835 vdd.n1718 185
R16375 vdd.n1720 vdd.n1719 185
R16376 vdd.n1831 vdd.n1722 185
R16377 vdd.n1830 vdd.n1723 185
R16378 vdd.n1829 vdd.n1724 185
R16379 vdd.n1726 vdd.n1725 185
R16380 vdd.n1825 vdd.n1728 185
R16381 vdd.n1824 vdd.n1729 185
R16382 vdd.n1823 vdd.n1730 185
R16383 vdd.n1732 vdd.n1731 185
R16384 vdd.n1819 vdd.n1734 185
R16385 vdd.n1818 vdd.n1735 185
R16386 vdd.n1817 vdd.n1736 185
R16387 vdd.n1738 vdd.n1737 185
R16388 vdd.n1813 vdd.n1740 185
R16389 vdd.n1812 vdd.n1809 185
R16390 vdd.n1808 vdd.n1741 185
R16391 vdd.n1743 vdd.n1742 185
R16392 vdd.n1804 vdd.n1745 185
R16393 vdd.n1803 vdd.n1746 185
R16394 vdd.n1802 vdd.n1747 185
R16395 vdd.n1749 vdd.n1748 185
R16396 vdd.n1798 vdd.n1751 185
R16397 vdd.n1797 vdd.n1752 185
R16398 vdd.n1796 vdd.n1753 185
R16399 vdd.n1755 vdd.n1754 185
R16400 vdd.n1792 vdd.n1757 185
R16401 vdd.n1791 vdd.n1758 185
R16402 vdd.n1790 vdd.n1759 185
R16403 vdd.n1761 vdd.n1760 185
R16404 vdd.n1786 vdd.n1763 185
R16405 vdd.n1785 vdd.n1764 185
R16406 vdd.n1784 vdd.n1765 185
R16407 vdd.n1767 vdd.n1766 185
R16408 vdd.n1780 vdd.n1769 185
R16409 vdd.n1779 vdd.n1770 185
R16410 vdd.n1778 vdd.n1771 185
R16411 vdd.n1775 vdd.n1679 185
R16412 vdd.n1873 vdd.n1679 185
R16413 vdd.n2361 vdd.n2360 185
R16414 vdd.n2365 vdd.n1525 185
R16415 vdd.n1524 vdd.n1518 185
R16416 vdd.n1522 vdd.n1521 185
R16417 vdd.n1520 vdd.n1279 185
R16418 vdd.n2369 vdd.n1276 185
R16419 vdd.n2371 vdd.n2370 185
R16420 vdd.n2373 vdd.n1274 185
R16421 vdd.n2375 vdd.n2374 185
R16422 vdd.n2376 vdd.n1269 185
R16423 vdd.n2378 vdd.n2377 185
R16424 vdd.n2380 vdd.n1267 185
R16425 vdd.n2382 vdd.n2381 185
R16426 vdd.n2383 vdd.n1262 185
R16427 vdd.n2385 vdd.n2384 185
R16428 vdd.n2387 vdd.n1260 185
R16429 vdd.n2389 vdd.n2388 185
R16430 vdd.n2390 vdd.n1256 185
R16431 vdd.n2392 vdd.n2391 185
R16432 vdd.n2394 vdd.n1253 185
R16433 vdd.n2396 vdd.n2395 185
R16434 vdd.n1254 vdd.n1247 185
R16435 vdd.n2400 vdd.n1251 185
R16436 vdd.n2401 vdd.n1243 185
R16437 vdd.n2403 vdd.n2402 185
R16438 vdd.n2405 vdd.n1241 185
R16439 vdd.n2407 vdd.n2406 185
R16440 vdd.n2408 vdd.n1236 185
R16441 vdd.n2410 vdd.n2409 185
R16442 vdd.n2412 vdd.n1234 185
R16443 vdd.n2414 vdd.n2413 185
R16444 vdd.n2415 vdd.n1229 185
R16445 vdd.n2417 vdd.n2416 185
R16446 vdd.n2419 vdd.n1227 185
R16447 vdd.n2421 vdd.n2420 185
R16448 vdd.n2422 vdd.n1222 185
R16449 vdd.n2424 vdd.n2423 185
R16450 vdd.n2426 vdd.n1220 185
R16451 vdd.n2428 vdd.n2427 185
R16452 vdd.n2429 vdd.n1216 185
R16453 vdd.n2431 vdd.n2430 185
R16454 vdd.n2433 vdd.n1213 185
R16455 vdd.n2435 vdd.n2434 185
R16456 vdd.n1214 vdd.n1207 185
R16457 vdd.n2439 vdd.n1211 185
R16458 vdd.n2440 vdd.n1203 185
R16459 vdd.n2442 vdd.n2441 185
R16460 vdd.n2444 vdd.n1201 185
R16461 vdd.n2446 vdd.n2445 185
R16462 vdd.n2447 vdd.n1196 185
R16463 vdd.n2449 vdd.n2448 185
R16464 vdd.n2451 vdd.n1194 185
R16465 vdd.n2453 vdd.n2452 185
R16466 vdd.n2454 vdd.n1189 185
R16467 vdd.n2456 vdd.n2455 185
R16468 vdd.n2458 vdd.n1187 185
R16469 vdd.n2460 vdd.n2459 185
R16470 vdd.n2461 vdd.n1185 185
R16471 vdd.n2463 vdd.n2462 185
R16472 vdd.n2466 vdd.n2465 185
R16473 vdd.n2468 vdd.n2467 185
R16474 vdd.n2470 vdd.n1183 185
R16475 vdd.n2472 vdd.n2471 185
R16476 vdd.n1530 vdd.n1182 185
R16477 vdd.n2359 vdd.n1528 185
R16478 vdd.n2359 vdd.n2358 185
R16479 vdd.n1538 vdd.n1527 185
R16480 vdd.n2349 vdd.n1527 185
R16481 vdd.n2348 vdd.n2347 185
R16482 vdd.n2350 vdd.n2348 185
R16483 vdd.n1537 vdd.n1536 185
R16484 vdd.n1536 vdd.n1535 185
R16485 vdd.n2341 vdd.n2340 185
R16486 vdd.n2340 vdd.n2339 185
R16487 vdd.n1541 vdd.n1540 185
R16488 vdd.n2330 vdd.n1541 185
R16489 vdd.n2329 vdd.n2328 185
R16490 vdd.n2331 vdd.n2329 185
R16491 vdd.n1548 vdd.n1547 185
R16492 vdd.n1553 vdd.n1547 185
R16493 vdd.n2324 vdd.n2323 185
R16494 vdd.n2323 vdd.n2322 185
R16495 vdd.n1551 vdd.n1550 185
R16496 vdd.n1552 vdd.n1551 185
R16497 vdd.n2313 vdd.n2312 185
R16498 vdd.n2314 vdd.n2313 185
R16499 vdd.n1561 vdd.n1560 185
R16500 vdd.n1560 vdd.n1559 185
R16501 vdd.n2308 vdd.n2307 185
R16502 vdd.n2307 vdd.n2306 185
R16503 vdd.n1564 vdd.n1563 185
R16504 vdd.n2297 vdd.n1564 185
R16505 vdd.n2296 vdd.n2295 185
R16506 vdd.n2298 vdd.n2296 185
R16507 vdd.n1571 vdd.n1570 185
R16508 vdd.n1575 vdd.n1570 185
R16509 vdd.n2291 vdd.n2290 185
R16510 vdd.n2290 vdd.n2289 185
R16511 vdd.n1574 vdd.n1573 185
R16512 vdd.n2280 vdd.n1574 185
R16513 vdd.n2279 vdd.n2278 185
R16514 vdd.n2281 vdd.n2279 185
R16515 vdd.n1583 vdd.n1582 185
R16516 vdd.n1582 vdd.n1581 185
R16517 vdd.n2274 vdd.n2273 185
R16518 vdd.n2273 vdd.n2272 185
R16519 vdd.n1586 vdd.n1585 185
R16520 vdd.n1587 vdd.n1586 185
R16521 vdd.n1956 vdd.n1955 185
R16522 vdd.n1957 vdd.n1956 185
R16523 vdd.n1594 vdd.n1593 185
R16524 vdd.n1598 vdd.n1593 185
R16525 vdd.n1951 vdd.n1950 185
R16526 vdd.n1950 vdd.n1949 185
R16527 vdd.n1597 vdd.n1596 185
R16528 vdd.n1940 vdd.n1597 185
R16529 vdd.n1939 vdd.n1938 185
R16530 vdd.n1941 vdd.n1939 185
R16531 vdd.n1605 vdd.n1604 185
R16532 vdd.n1610 vdd.n1604 185
R16533 vdd.n1934 vdd.n1933 185
R16534 vdd.n1933 vdd.n1932 185
R16535 vdd.n1608 vdd.n1607 185
R16536 vdd.n1609 vdd.n1608 185
R16537 vdd.n1923 vdd.n1922 185
R16538 vdd.n1924 vdd.n1923 185
R16539 vdd.n1618 vdd.n1617 185
R16540 vdd.n1617 vdd.n1616 185
R16541 vdd.n1918 vdd.n1917 185
R16542 vdd.n1917 vdd.n1916 185
R16543 vdd.n1621 vdd.n1620 185
R16544 vdd.n1907 vdd.n1621 185
R16545 vdd.n1906 vdd.n1905 185
R16546 vdd.n1908 vdd.n1906 185
R16547 vdd.n1628 vdd.n1627 185
R16548 vdd.n1632 vdd.n1627 185
R16549 vdd.n1901 vdd.n1900 185
R16550 vdd.n1900 vdd.n1899 185
R16551 vdd.n1631 vdd.n1630 185
R16552 vdd.n1890 vdd.n1631 185
R16553 vdd.n1889 vdd.n1888 185
R16554 vdd.n1891 vdd.n1889 185
R16555 vdd.n1640 vdd.n1639 185
R16556 vdd.n1639 vdd.n1638 185
R16557 vdd.n1884 vdd.n1883 185
R16558 vdd.n1883 vdd.n1882 185
R16559 vdd.n1643 vdd.n1642 185
R16560 vdd.n1680 vdd.n1643 185
R16561 vdd.n1000 vdd.n998 185
R16562 vdd.n2712 vdd.n998 185
R16563 vdd.n2634 vdd.n1018 185
R16564 vdd.n1018 vdd.n1005 185
R16565 vdd.n2636 vdd.n2635 185
R16566 vdd.n2637 vdd.n2636 185
R16567 vdd.n2633 vdd.n1017 185
R16568 vdd.n1399 vdd.n1017 185
R16569 vdd.n2632 vdd.n2631 185
R16570 vdd.n2631 vdd.n2630 185
R16571 vdd.n1020 vdd.n1019 185
R16572 vdd.n1021 vdd.n1020 185
R16573 vdd.n2621 vdd.n2620 185
R16574 vdd.n2622 vdd.n2621 185
R16575 vdd.n2619 vdd.n1031 185
R16576 vdd.n1031 vdd.n1028 185
R16577 vdd.n2618 vdd.n2617 185
R16578 vdd.n2617 vdd.n2616 185
R16579 vdd.n1033 vdd.n1032 185
R16580 vdd.n1425 vdd.n1033 185
R16581 vdd.n2609 vdd.n2608 185
R16582 vdd.n2610 vdd.n2609 185
R16583 vdd.n2607 vdd.n1041 185
R16584 vdd.n1046 vdd.n1041 185
R16585 vdd.n2606 vdd.n2605 185
R16586 vdd.n2605 vdd.n2604 185
R16587 vdd.n1043 vdd.n1042 185
R16588 vdd.n1052 vdd.n1043 185
R16589 vdd.n2597 vdd.n2596 185
R16590 vdd.n2598 vdd.n2597 185
R16591 vdd.n2595 vdd.n1053 185
R16592 vdd.n1437 vdd.n1053 185
R16593 vdd.n2594 vdd.n2593 185
R16594 vdd.n2593 vdd.n2592 185
R16595 vdd.n1055 vdd.n1054 185
R16596 vdd.n1056 vdd.n1055 185
R16597 vdd.n2585 vdd.n2584 185
R16598 vdd.n2586 vdd.n2585 185
R16599 vdd.n2583 vdd.n1065 185
R16600 vdd.n1065 vdd.n1062 185
R16601 vdd.n2582 vdd.n2581 185
R16602 vdd.n2581 vdd.n2580 185
R16603 vdd.n1067 vdd.n1066 185
R16604 vdd.n1076 vdd.n1067 185
R16605 vdd.n2572 vdd.n2571 185
R16606 vdd.n2573 vdd.n2572 185
R16607 vdd.n2570 vdd.n1077 185
R16608 vdd.n1083 vdd.n1077 185
R16609 vdd.n2569 vdd.n2568 185
R16610 vdd.n2568 vdd.n2567 185
R16611 vdd.n1079 vdd.n1078 185
R16612 vdd.n1080 vdd.n1079 185
R16613 vdd.n2560 vdd.n2559 185
R16614 vdd.n2561 vdd.n2560 185
R16615 vdd.n2558 vdd.n1090 185
R16616 vdd.n1090 vdd.n1087 185
R16617 vdd.n2557 vdd.n2556 185
R16618 vdd.n2556 vdd.n2555 185
R16619 vdd.n1092 vdd.n1091 185
R16620 vdd.n1093 vdd.n1092 185
R16621 vdd.n2548 vdd.n2547 185
R16622 vdd.n2549 vdd.n2548 185
R16623 vdd.n2546 vdd.n1101 185
R16624 vdd.n1106 vdd.n1101 185
R16625 vdd.n2545 vdd.n2544 185
R16626 vdd.n2544 vdd.n2543 185
R16627 vdd.n1103 vdd.n1102 185
R16628 vdd.n1112 vdd.n1103 185
R16629 vdd.n2536 vdd.n2535 185
R16630 vdd.n2537 vdd.n2536 185
R16631 vdd.n2534 vdd.n1113 185
R16632 vdd.n1119 vdd.n1113 185
R16633 vdd.n2533 vdd.n2532 185
R16634 vdd.n2532 vdd.n2531 185
R16635 vdd.n1115 vdd.n1114 185
R16636 vdd.n1116 vdd.n1115 185
R16637 vdd.n2524 vdd.n2523 185
R16638 vdd.n2525 vdd.n2524 185
R16639 vdd.n2522 vdd.n1126 185
R16640 vdd.n1126 vdd.n1123 185
R16641 vdd.n2521 vdd.n2520 185
R16642 vdd.n2520 vdd.n2519 185
R16643 vdd.n1128 vdd.n1127 185
R16644 vdd.n1137 vdd.n1128 185
R16645 vdd.n2512 vdd.n2511 185
R16646 vdd.n2513 vdd.n2512 185
R16647 vdd.n2510 vdd.n1138 185
R16648 vdd.n1138 vdd.n1134 185
R16649 vdd.n2509 vdd.n2508 185
R16650 vdd.n1140 vdd.n1139 185
R16651 vdd.n2505 vdd.n2504 185
R16652 vdd.n2506 vdd.n2505 185
R16653 vdd.n2503 vdd.n1176 185
R16654 vdd.n2502 vdd.n2501 185
R16655 vdd.n2500 vdd.n2499 185
R16656 vdd.n2498 vdd.n2497 185
R16657 vdd.n2496 vdd.n2495 185
R16658 vdd.n2494 vdd.n2493 185
R16659 vdd.n2492 vdd.n2491 185
R16660 vdd.n2490 vdd.n2489 185
R16661 vdd.n2488 vdd.n2487 185
R16662 vdd.n2486 vdd.n2485 185
R16663 vdd.n2484 vdd.n2483 185
R16664 vdd.n2482 vdd.n2481 185
R16665 vdd.n2480 vdd.n2479 185
R16666 vdd.n2478 vdd.n2477 185
R16667 vdd.n2476 vdd.n2475 185
R16668 vdd.n1321 vdd.n1177 185
R16669 vdd.n1323 vdd.n1322 185
R16670 vdd.n1325 vdd.n1324 185
R16671 vdd.n1327 vdd.n1326 185
R16672 vdd.n1329 vdd.n1328 185
R16673 vdd.n1331 vdd.n1330 185
R16674 vdd.n1333 vdd.n1332 185
R16675 vdd.n1335 vdd.n1334 185
R16676 vdd.n1337 vdd.n1336 185
R16677 vdd.n1339 vdd.n1338 185
R16678 vdd.n1341 vdd.n1340 185
R16679 vdd.n1343 vdd.n1342 185
R16680 vdd.n1345 vdd.n1344 185
R16681 vdd.n1347 vdd.n1346 185
R16682 vdd.n1350 vdd.n1349 185
R16683 vdd.n1352 vdd.n1351 185
R16684 vdd.n1354 vdd.n1353 185
R16685 vdd.n2715 vdd.n2714 185
R16686 vdd.n2717 vdd.n2716 185
R16687 vdd.n2719 vdd.n2718 185
R16688 vdd.n2722 vdd.n2721 185
R16689 vdd.n2724 vdd.n2723 185
R16690 vdd.n2726 vdd.n2725 185
R16691 vdd.n2728 vdd.n2727 185
R16692 vdd.n2730 vdd.n2729 185
R16693 vdd.n2732 vdd.n2731 185
R16694 vdd.n2734 vdd.n2733 185
R16695 vdd.n2736 vdd.n2735 185
R16696 vdd.n2738 vdd.n2737 185
R16697 vdd.n2740 vdd.n2739 185
R16698 vdd.n2742 vdd.n2741 185
R16699 vdd.n2744 vdd.n2743 185
R16700 vdd.n2746 vdd.n2745 185
R16701 vdd.n2748 vdd.n2747 185
R16702 vdd.n2750 vdd.n2749 185
R16703 vdd.n2752 vdd.n2751 185
R16704 vdd.n2754 vdd.n2753 185
R16705 vdd.n2756 vdd.n2755 185
R16706 vdd.n2758 vdd.n2757 185
R16707 vdd.n2760 vdd.n2759 185
R16708 vdd.n2762 vdd.n2761 185
R16709 vdd.n2764 vdd.n2763 185
R16710 vdd.n2766 vdd.n2765 185
R16711 vdd.n2768 vdd.n2767 185
R16712 vdd.n2770 vdd.n2769 185
R16713 vdd.n2772 vdd.n2771 185
R16714 vdd.n2774 vdd.n2773 185
R16715 vdd.n2776 vdd.n2775 185
R16716 vdd.n2778 vdd.n2777 185
R16717 vdd.n2780 vdd.n2779 185
R16718 vdd.n2781 vdd.n999 185
R16719 vdd.n2783 vdd.n2782 185
R16720 vdd.n2784 vdd.n2783 185
R16721 vdd.n2713 vdd.n1003 185
R16722 vdd.n2713 vdd.n2712 185
R16723 vdd.n1397 vdd.n1004 185
R16724 vdd.n1005 vdd.n1004 185
R16725 vdd.n1398 vdd.n1015 185
R16726 vdd.n2637 vdd.n1015 185
R16727 vdd.n1401 vdd.n1400 185
R16728 vdd.n1400 vdd.n1399 185
R16729 vdd.n1402 vdd.n1022 185
R16730 vdd.n2630 vdd.n1022 185
R16731 vdd.n1404 vdd.n1403 185
R16732 vdd.n1403 vdd.n1021 185
R16733 vdd.n1405 vdd.n1029 185
R16734 vdd.n2622 vdd.n1029 185
R16735 vdd.n1407 vdd.n1406 185
R16736 vdd.n1406 vdd.n1028 185
R16737 vdd.n1408 vdd.n1034 185
R16738 vdd.n2616 vdd.n1034 185
R16739 vdd.n1427 vdd.n1426 185
R16740 vdd.n1426 vdd.n1425 185
R16741 vdd.n1428 vdd.n1039 185
R16742 vdd.n2610 vdd.n1039 185
R16743 vdd.n1430 vdd.n1429 185
R16744 vdd.n1429 vdd.n1046 185
R16745 vdd.n1431 vdd.n1044 185
R16746 vdd.n2604 vdd.n1044 185
R16747 vdd.n1433 vdd.n1432 185
R16748 vdd.n1432 vdd.n1052 185
R16749 vdd.n1434 vdd.n1050 185
R16750 vdd.n2598 vdd.n1050 185
R16751 vdd.n1436 vdd.n1435 185
R16752 vdd.n1437 vdd.n1436 185
R16753 vdd.n1396 vdd.n1057 185
R16754 vdd.n2592 vdd.n1057 185
R16755 vdd.n1395 vdd.n1394 185
R16756 vdd.n1394 vdd.n1056 185
R16757 vdd.n1393 vdd.n1063 185
R16758 vdd.n2586 vdd.n1063 185
R16759 vdd.n1392 vdd.n1391 185
R16760 vdd.n1391 vdd.n1062 185
R16761 vdd.n1390 vdd.n1068 185
R16762 vdd.n2580 vdd.n1068 185
R16763 vdd.n1389 vdd.n1388 185
R16764 vdd.n1388 vdd.n1076 185
R16765 vdd.n1387 vdd.n1074 185
R16766 vdd.n2573 vdd.n1074 185
R16767 vdd.n1386 vdd.n1385 185
R16768 vdd.n1385 vdd.n1083 185
R16769 vdd.n1384 vdd.n1081 185
R16770 vdd.n2567 vdd.n1081 185
R16771 vdd.n1383 vdd.n1382 185
R16772 vdd.n1382 vdd.n1080 185
R16773 vdd.n1381 vdd.n1088 185
R16774 vdd.n2561 vdd.n1088 185
R16775 vdd.n1380 vdd.n1379 185
R16776 vdd.n1379 vdd.n1087 185
R16777 vdd.n1378 vdd.n1094 185
R16778 vdd.n2555 vdd.n1094 185
R16779 vdd.n1377 vdd.n1376 185
R16780 vdd.n1376 vdd.n1093 185
R16781 vdd.n1375 vdd.n1099 185
R16782 vdd.n2549 vdd.n1099 185
R16783 vdd.n1374 vdd.n1373 185
R16784 vdd.n1373 vdd.n1106 185
R16785 vdd.n1372 vdd.n1104 185
R16786 vdd.n2543 vdd.n1104 185
R16787 vdd.n1371 vdd.n1370 185
R16788 vdd.n1370 vdd.n1112 185
R16789 vdd.n1369 vdd.n1110 185
R16790 vdd.n2537 vdd.n1110 185
R16791 vdd.n1368 vdd.n1367 185
R16792 vdd.n1367 vdd.n1119 185
R16793 vdd.n1366 vdd.n1117 185
R16794 vdd.n2531 vdd.n1117 185
R16795 vdd.n1365 vdd.n1364 185
R16796 vdd.n1364 vdd.n1116 185
R16797 vdd.n1363 vdd.n1124 185
R16798 vdd.n2525 vdd.n1124 185
R16799 vdd.n1362 vdd.n1361 185
R16800 vdd.n1361 vdd.n1123 185
R16801 vdd.n1360 vdd.n1129 185
R16802 vdd.n2519 vdd.n1129 185
R16803 vdd.n1359 vdd.n1358 185
R16804 vdd.n1358 vdd.n1137 185
R16805 vdd.n1357 vdd.n1135 185
R16806 vdd.n2513 vdd.n1135 185
R16807 vdd.n1356 vdd.n1355 185
R16808 vdd.n1355 vdd.n1134 185
R16809 vdd.n3629 vdd.n3628 185
R16810 vdd.n3628 vdd.n3627 185
R16811 vdd.n3630 vdd.n387 185
R16812 vdd.n387 vdd.n386 185
R16813 vdd.n3632 vdd.n3631 185
R16814 vdd.n3633 vdd.n3632 185
R16815 vdd.n382 vdd.n381 185
R16816 vdd.n3634 vdd.n382 185
R16817 vdd.n3637 vdd.n3636 185
R16818 vdd.n3636 vdd.n3635 185
R16819 vdd.n3638 vdd.n376 185
R16820 vdd.n376 vdd.n375 185
R16821 vdd.n3640 vdd.n3639 185
R16822 vdd.n3641 vdd.n3640 185
R16823 vdd.n371 vdd.n370 185
R16824 vdd.n3642 vdd.n371 185
R16825 vdd.n3645 vdd.n3644 185
R16826 vdd.n3644 vdd.n3643 185
R16827 vdd.n3646 vdd.n365 185
R16828 vdd.n3603 vdd.n365 185
R16829 vdd.n3648 vdd.n3647 185
R16830 vdd.n3649 vdd.n3648 185
R16831 vdd.n360 vdd.n359 185
R16832 vdd.n3650 vdd.n360 185
R16833 vdd.n3653 vdd.n3652 185
R16834 vdd.n3652 vdd.n3651 185
R16835 vdd.n3654 vdd.n354 185
R16836 vdd.n361 vdd.n354 185
R16837 vdd.n3656 vdd.n3655 185
R16838 vdd.n3657 vdd.n3656 185
R16839 vdd.n350 vdd.n349 185
R16840 vdd.n3658 vdd.n350 185
R16841 vdd.n3661 vdd.n3660 185
R16842 vdd.n3660 vdd.n3659 185
R16843 vdd.n3662 vdd.n345 185
R16844 vdd.n345 vdd.n344 185
R16845 vdd.n3664 vdd.n3663 185
R16846 vdd.n3665 vdd.n3664 185
R16847 vdd.n339 vdd.n337 185
R16848 vdd.n3666 vdd.n339 185
R16849 vdd.n3669 vdd.n3668 185
R16850 vdd.n3668 vdd.n3667 185
R16851 vdd.n338 vdd.n336 185
R16852 vdd.n340 vdd.n338 185
R16853 vdd.n3579 vdd.n3578 185
R16854 vdd.n3580 vdd.n3579 185
R16855 vdd.n635 vdd.n634 185
R16856 vdd.n634 vdd.n633 185
R16857 vdd.n3574 vdd.n3573 185
R16858 vdd.n3573 vdd.n3572 185
R16859 vdd.n638 vdd.n637 185
R16860 vdd.n644 vdd.n638 185
R16861 vdd.n3560 vdd.n3559 185
R16862 vdd.n3561 vdd.n3560 185
R16863 vdd.n646 vdd.n645 185
R16864 vdd.n3552 vdd.n645 185
R16865 vdd.n3555 vdd.n3554 185
R16866 vdd.n3554 vdd.n3553 185
R16867 vdd.n649 vdd.n648 185
R16868 vdd.n656 vdd.n649 185
R16869 vdd.n3543 vdd.n3542 185
R16870 vdd.n3544 vdd.n3543 185
R16871 vdd.n658 vdd.n657 185
R16872 vdd.n657 vdd.n655 185
R16873 vdd.n3538 vdd.n3537 185
R16874 vdd.n3537 vdd.n3536 185
R16875 vdd.n661 vdd.n660 185
R16876 vdd.n662 vdd.n661 185
R16877 vdd.n3527 vdd.n3526 185
R16878 vdd.n3528 vdd.n3527 185
R16879 vdd.n669 vdd.n668 185
R16880 vdd.n3519 vdd.n668 185
R16881 vdd.n3522 vdd.n3521 185
R16882 vdd.n3521 vdd.n3520 185
R16883 vdd.n672 vdd.n671 185
R16884 vdd.n679 vdd.n672 185
R16885 vdd.n3510 vdd.n3509 185
R16886 vdd.n3511 vdd.n3510 185
R16887 vdd.n681 vdd.n680 185
R16888 vdd.n680 vdd.n678 185
R16889 vdd.n3505 vdd.n3504 185
R16890 vdd.n3504 vdd.n3503 185
R16891 vdd.n684 vdd.n683 185
R16892 vdd.n723 vdd.n684 185
R16893 vdd.n3493 vdd.n3492 185
R16894 vdd.n3491 vdd.n725 185
R16895 vdd.n3490 vdd.n724 185
R16896 vdd.n3495 vdd.n724 185
R16897 vdd.n729 vdd.n728 185
R16898 vdd.n733 vdd.n732 185
R16899 vdd.n3486 vdd.n734 185
R16900 vdd.n3485 vdd.n3484 185
R16901 vdd.n3483 vdd.n3482 185
R16902 vdd.n3481 vdd.n3480 185
R16903 vdd.n3479 vdd.n3478 185
R16904 vdd.n3477 vdd.n3476 185
R16905 vdd.n3475 vdd.n3474 185
R16906 vdd.n3473 vdd.n3472 185
R16907 vdd.n3471 vdd.n3470 185
R16908 vdd.n3469 vdd.n3468 185
R16909 vdd.n3467 vdd.n3466 185
R16910 vdd.n3465 vdd.n3464 185
R16911 vdd.n3463 vdd.n3462 185
R16912 vdd.n3461 vdd.n3460 185
R16913 vdd.n3459 vdd.n3458 185
R16914 vdd.n3450 vdd.n747 185
R16915 vdd.n3452 vdd.n3451 185
R16916 vdd.n3449 vdd.n3448 185
R16917 vdd.n3447 vdd.n3446 185
R16918 vdd.n3445 vdd.n3444 185
R16919 vdd.n3443 vdd.n3442 185
R16920 vdd.n3441 vdd.n3440 185
R16921 vdd.n3439 vdd.n3438 185
R16922 vdd.n3437 vdd.n3436 185
R16923 vdd.n3435 vdd.n3434 185
R16924 vdd.n3433 vdd.n3432 185
R16925 vdd.n3431 vdd.n3430 185
R16926 vdd.n3429 vdd.n3428 185
R16927 vdd.n3427 vdd.n3426 185
R16928 vdd.n3425 vdd.n3424 185
R16929 vdd.n3423 vdd.n3422 185
R16930 vdd.n3421 vdd.n3420 185
R16931 vdd.n3419 vdd.n3418 185
R16932 vdd.n3417 vdd.n3416 185
R16933 vdd.n3415 vdd.n3414 185
R16934 vdd.n3413 vdd.n3412 185
R16935 vdd.n3411 vdd.n3410 185
R16936 vdd.n3404 vdd.n767 185
R16937 vdd.n3406 vdd.n3405 185
R16938 vdd.n3403 vdd.n3402 185
R16939 vdd.n3401 vdd.n3400 185
R16940 vdd.n3399 vdd.n3398 185
R16941 vdd.n3397 vdd.n3396 185
R16942 vdd.n3395 vdd.n3394 185
R16943 vdd.n3393 vdd.n3392 185
R16944 vdd.n3391 vdd.n3390 185
R16945 vdd.n3389 vdd.n3388 185
R16946 vdd.n3387 vdd.n3386 185
R16947 vdd.n3385 vdd.n3384 185
R16948 vdd.n3383 vdd.n3382 185
R16949 vdd.n3381 vdd.n3380 185
R16950 vdd.n3379 vdd.n3378 185
R16951 vdd.n3377 vdd.n3376 185
R16952 vdd.n3375 vdd.n3374 185
R16953 vdd.n3373 vdd.n3372 185
R16954 vdd.n3371 vdd.n3370 185
R16955 vdd.n3369 vdd.n3368 185
R16956 vdd.n3367 vdd.n691 185
R16957 vdd.n3497 vdd.n3496 185
R16958 vdd.n3496 vdd.n3495 185
R16959 vdd.n3624 vdd.n3623 185
R16960 vdd.n618 vdd.n425 185
R16961 vdd.n617 vdd.n616 185
R16962 vdd.n615 vdd.n614 185
R16963 vdd.n613 vdd.n430 185
R16964 vdd.n609 vdd.n608 185
R16965 vdd.n607 vdd.n606 185
R16966 vdd.n605 vdd.n604 185
R16967 vdd.n603 vdd.n432 185
R16968 vdd.n599 vdd.n598 185
R16969 vdd.n597 vdd.n596 185
R16970 vdd.n595 vdd.n594 185
R16971 vdd.n593 vdd.n434 185
R16972 vdd.n589 vdd.n588 185
R16973 vdd.n587 vdd.n586 185
R16974 vdd.n585 vdd.n584 185
R16975 vdd.n583 vdd.n436 185
R16976 vdd.n579 vdd.n578 185
R16977 vdd.n577 vdd.n576 185
R16978 vdd.n575 vdd.n574 185
R16979 vdd.n573 vdd.n438 185
R16980 vdd.n569 vdd.n568 185
R16981 vdd.n567 vdd.n566 185
R16982 vdd.n565 vdd.n564 185
R16983 vdd.n563 vdd.n442 185
R16984 vdd.n559 vdd.n558 185
R16985 vdd.n557 vdd.n556 185
R16986 vdd.n555 vdd.n554 185
R16987 vdd.n553 vdd.n444 185
R16988 vdd.n549 vdd.n548 185
R16989 vdd.n547 vdd.n546 185
R16990 vdd.n545 vdd.n544 185
R16991 vdd.n543 vdd.n446 185
R16992 vdd.n539 vdd.n538 185
R16993 vdd.n537 vdd.n536 185
R16994 vdd.n535 vdd.n534 185
R16995 vdd.n533 vdd.n448 185
R16996 vdd.n529 vdd.n528 185
R16997 vdd.n527 vdd.n526 185
R16998 vdd.n525 vdd.n524 185
R16999 vdd.n523 vdd.n450 185
R17000 vdd.n519 vdd.n518 185
R17001 vdd.n517 vdd.n516 185
R17002 vdd.n515 vdd.n514 185
R17003 vdd.n513 vdd.n454 185
R17004 vdd.n509 vdd.n508 185
R17005 vdd.n507 vdd.n506 185
R17006 vdd.n505 vdd.n504 185
R17007 vdd.n503 vdd.n456 185
R17008 vdd.n499 vdd.n498 185
R17009 vdd.n497 vdd.n496 185
R17010 vdd.n495 vdd.n494 185
R17011 vdd.n493 vdd.n458 185
R17012 vdd.n489 vdd.n488 185
R17013 vdd.n487 vdd.n486 185
R17014 vdd.n485 vdd.n484 185
R17015 vdd.n483 vdd.n460 185
R17016 vdd.n479 vdd.n478 185
R17017 vdd.n477 vdd.n476 185
R17018 vdd.n475 vdd.n474 185
R17019 vdd.n473 vdd.n462 185
R17020 vdd.n469 vdd.n468 185
R17021 vdd.n467 vdd.n466 185
R17022 vdd.n465 vdd.n392 185
R17023 vdd.n3620 vdd.n393 185
R17024 vdd.n3627 vdd.n393 185
R17025 vdd.n3619 vdd.n3618 185
R17026 vdd.n3618 vdd.n386 185
R17027 vdd.n3617 vdd.n385 185
R17028 vdd.n3633 vdd.n385 185
R17029 vdd.n621 vdd.n384 185
R17030 vdd.n3634 vdd.n384 185
R17031 vdd.n3613 vdd.n383 185
R17032 vdd.n3635 vdd.n383 185
R17033 vdd.n3612 vdd.n3611 185
R17034 vdd.n3611 vdd.n375 185
R17035 vdd.n3610 vdd.n374 185
R17036 vdd.n3641 vdd.n374 185
R17037 vdd.n623 vdd.n373 185
R17038 vdd.n3642 vdd.n373 185
R17039 vdd.n3606 vdd.n372 185
R17040 vdd.n3643 vdd.n372 185
R17041 vdd.n3605 vdd.n3604 185
R17042 vdd.n3604 vdd.n3603 185
R17043 vdd.n3602 vdd.n364 185
R17044 vdd.n3649 vdd.n364 185
R17045 vdd.n625 vdd.n363 185
R17046 vdd.n3650 vdd.n363 185
R17047 vdd.n3598 vdd.n362 185
R17048 vdd.n3651 vdd.n362 185
R17049 vdd.n3597 vdd.n3596 185
R17050 vdd.n3596 vdd.n361 185
R17051 vdd.n3595 vdd.n353 185
R17052 vdd.n3657 vdd.n353 185
R17053 vdd.n627 vdd.n352 185
R17054 vdd.n3658 vdd.n352 185
R17055 vdd.n3591 vdd.n351 185
R17056 vdd.n3659 vdd.n351 185
R17057 vdd.n3590 vdd.n3589 185
R17058 vdd.n3589 vdd.n344 185
R17059 vdd.n3588 vdd.n343 185
R17060 vdd.n3665 vdd.n343 185
R17061 vdd.n629 vdd.n342 185
R17062 vdd.n3666 vdd.n342 185
R17063 vdd.n3584 vdd.n341 185
R17064 vdd.n3667 vdd.n341 185
R17065 vdd.n3583 vdd.n3582 185
R17066 vdd.n3582 vdd.n340 185
R17067 vdd.n3581 vdd.n631 185
R17068 vdd.n3581 vdd.n3580 185
R17069 vdd.n3569 vdd.n632 185
R17070 vdd.n633 vdd.n632 185
R17071 vdd.n3571 vdd.n3570 185
R17072 vdd.n3572 vdd.n3571 185
R17073 vdd.n640 vdd.n639 185
R17074 vdd.n644 vdd.n639 185
R17075 vdd.n3563 vdd.n3562 185
R17076 vdd.n3562 vdd.n3561 185
R17077 vdd.n643 vdd.n642 185
R17078 vdd.n3552 vdd.n643 185
R17079 vdd.n3551 vdd.n3550 185
R17080 vdd.n3553 vdd.n3551 185
R17081 vdd.n651 vdd.n650 185
R17082 vdd.n656 vdd.n650 185
R17083 vdd.n3546 vdd.n3545 185
R17084 vdd.n3545 vdd.n3544 185
R17085 vdd.n654 vdd.n653 185
R17086 vdd.n655 vdd.n654 185
R17087 vdd.n3535 vdd.n3534 185
R17088 vdd.n3536 vdd.n3535 185
R17089 vdd.n664 vdd.n663 185
R17090 vdd.n663 vdd.n662 185
R17091 vdd.n3530 vdd.n3529 185
R17092 vdd.n3529 vdd.n3528 185
R17093 vdd.n667 vdd.n666 185
R17094 vdd.n3519 vdd.n667 185
R17095 vdd.n3518 vdd.n3517 185
R17096 vdd.n3520 vdd.n3518 185
R17097 vdd.n674 vdd.n673 185
R17098 vdd.n679 vdd.n673 185
R17099 vdd.n3513 vdd.n3512 185
R17100 vdd.n3512 vdd.n3511 185
R17101 vdd.n677 vdd.n676 185
R17102 vdd.n678 vdd.n677 185
R17103 vdd.n3502 vdd.n3501 185
R17104 vdd.n3503 vdd.n3502 185
R17105 vdd.n686 vdd.n685 185
R17106 vdd.n723 vdd.n685 185
R17107 vdd.n3091 vdd.n3090 185
R17108 vdd.n962 vdd.n961 185
R17109 vdd.n3087 vdd.n3086 185
R17110 vdd.n3088 vdd.n3087 185
R17111 vdd.n3085 vdd.n2819 185
R17112 vdd.n3084 vdd.n3083 185
R17113 vdd.n3082 vdd.n3081 185
R17114 vdd.n3080 vdd.n3079 185
R17115 vdd.n3078 vdd.n3077 185
R17116 vdd.n3076 vdd.n3075 185
R17117 vdd.n3074 vdd.n3073 185
R17118 vdd.n3072 vdd.n3071 185
R17119 vdd.n3070 vdd.n3069 185
R17120 vdd.n3068 vdd.n3067 185
R17121 vdd.n3066 vdd.n3065 185
R17122 vdd.n3064 vdd.n3063 185
R17123 vdd.n3062 vdd.n3061 185
R17124 vdd.n3060 vdd.n3059 185
R17125 vdd.n3058 vdd.n3057 185
R17126 vdd.n3056 vdd.n3055 185
R17127 vdd.n3054 vdd.n3053 185
R17128 vdd.n3052 vdd.n3051 185
R17129 vdd.n3050 vdd.n3049 185
R17130 vdd.n3048 vdd.n3047 185
R17131 vdd.n3046 vdd.n3045 185
R17132 vdd.n3044 vdd.n3043 185
R17133 vdd.n3042 vdd.n3041 185
R17134 vdd.n3040 vdd.n3039 185
R17135 vdd.n3038 vdd.n3037 185
R17136 vdd.n3036 vdd.n3035 185
R17137 vdd.n3034 vdd.n3033 185
R17138 vdd.n3032 vdd.n3031 185
R17139 vdd.n3030 vdd.n3029 185
R17140 vdd.n3027 vdd.n3026 185
R17141 vdd.n3025 vdd.n3024 185
R17142 vdd.n3023 vdd.n3022 185
R17143 vdd.n3267 vdd.n3266 185
R17144 vdd.n3269 vdd.n834 185
R17145 vdd.n3271 vdd.n3270 185
R17146 vdd.n3273 vdd.n831 185
R17147 vdd.n3275 vdd.n3274 185
R17148 vdd.n3277 vdd.n829 185
R17149 vdd.n3279 vdd.n3278 185
R17150 vdd.n3280 vdd.n828 185
R17151 vdd.n3282 vdd.n3281 185
R17152 vdd.n3284 vdd.n826 185
R17153 vdd.n3286 vdd.n3285 185
R17154 vdd.n3287 vdd.n825 185
R17155 vdd.n3289 vdd.n3288 185
R17156 vdd.n3291 vdd.n823 185
R17157 vdd.n3293 vdd.n3292 185
R17158 vdd.n3294 vdd.n822 185
R17159 vdd.n3296 vdd.n3295 185
R17160 vdd.n3298 vdd.n731 185
R17161 vdd.n3300 vdd.n3299 185
R17162 vdd.n3302 vdd.n820 185
R17163 vdd.n3304 vdd.n3303 185
R17164 vdd.n3305 vdd.n819 185
R17165 vdd.n3307 vdd.n3306 185
R17166 vdd.n3309 vdd.n817 185
R17167 vdd.n3311 vdd.n3310 185
R17168 vdd.n3312 vdd.n816 185
R17169 vdd.n3314 vdd.n3313 185
R17170 vdd.n3316 vdd.n814 185
R17171 vdd.n3318 vdd.n3317 185
R17172 vdd.n3319 vdd.n813 185
R17173 vdd.n3321 vdd.n3320 185
R17174 vdd.n3323 vdd.n812 185
R17175 vdd.n3324 vdd.n811 185
R17176 vdd.n3327 vdd.n3326 185
R17177 vdd.n3328 vdd.n809 185
R17178 vdd.n809 vdd.n692 185
R17179 vdd.n3265 vdd.n806 185
R17180 vdd.n3331 vdd.n806 185
R17181 vdd.n3264 vdd.n3263 185
R17182 vdd.n3263 vdd.n805 185
R17183 vdd.n3262 vdd.n836 185
R17184 vdd.n3262 vdd.n3261 185
R17185 vdd.n2905 vdd.n837 185
R17186 vdd.n846 vdd.n837 185
R17187 vdd.n2906 vdd.n844 185
R17188 vdd.n3255 vdd.n844 185
R17189 vdd.n2908 vdd.n2907 185
R17190 vdd.n2907 vdd.n843 185
R17191 vdd.n2909 vdd.n852 185
R17192 vdd.n3204 vdd.n852 185
R17193 vdd.n2911 vdd.n2910 185
R17194 vdd.n2910 vdd.n851 185
R17195 vdd.n2912 vdd.n857 185
R17196 vdd.n3198 vdd.n857 185
R17197 vdd.n2914 vdd.n2913 185
R17198 vdd.n2913 vdd.n864 185
R17199 vdd.n2915 vdd.n862 185
R17200 vdd.n3192 vdd.n862 185
R17201 vdd.n2917 vdd.n2916 185
R17202 vdd.n2916 vdd.n870 185
R17203 vdd.n2918 vdd.n868 185
R17204 vdd.n3186 vdd.n868 185
R17205 vdd.n2920 vdd.n2919 185
R17206 vdd.n2919 vdd.n877 185
R17207 vdd.n2921 vdd.n875 185
R17208 vdd.n3180 vdd.n875 185
R17209 vdd.n2923 vdd.n2922 185
R17210 vdd.n2922 vdd.n874 185
R17211 vdd.n2924 vdd.n882 185
R17212 vdd.n3174 vdd.n882 185
R17213 vdd.n2926 vdd.n2925 185
R17214 vdd.n2925 vdd.n881 185
R17215 vdd.n2927 vdd.n888 185
R17216 vdd.n3168 vdd.n888 185
R17217 vdd.n2929 vdd.n2928 185
R17218 vdd.n2928 vdd.n887 185
R17219 vdd.n2930 vdd.n893 185
R17220 vdd.n3162 vdd.n893 185
R17221 vdd.n2932 vdd.n2931 185
R17222 vdd.n2931 vdd.n901 185
R17223 vdd.n2933 vdd.n899 185
R17224 vdd.n3156 vdd.n899 185
R17225 vdd.n2935 vdd.n2934 185
R17226 vdd.n2934 vdd.n908 185
R17227 vdd.n2936 vdd.n906 185
R17228 vdd.n3150 vdd.n906 185
R17229 vdd.n2938 vdd.n2937 185
R17230 vdd.n2937 vdd.n905 185
R17231 vdd.n2939 vdd.n913 185
R17232 vdd.n3143 vdd.n913 185
R17233 vdd.n2941 vdd.n2940 185
R17234 vdd.n2940 vdd.n912 185
R17235 vdd.n2942 vdd.n918 185
R17236 vdd.n3137 vdd.n918 185
R17237 vdd.n2944 vdd.n2943 185
R17238 vdd.n2943 vdd.n925 185
R17239 vdd.n2945 vdd.n923 185
R17240 vdd.n3131 vdd.n923 185
R17241 vdd.n2947 vdd.n2946 185
R17242 vdd.n2946 vdd.n931 185
R17243 vdd.n2948 vdd.n929 185
R17244 vdd.n3125 vdd.n929 185
R17245 vdd.n3000 vdd.n2999 185
R17246 vdd.n2999 vdd.n2998 185
R17247 vdd.n3001 vdd.n935 185
R17248 vdd.n3119 vdd.n935 185
R17249 vdd.n3003 vdd.n3002 185
R17250 vdd.n3004 vdd.n3003 185
R17251 vdd.n2904 vdd.n941 185
R17252 vdd.n3113 vdd.n941 185
R17253 vdd.n2903 vdd.n2902 185
R17254 vdd.n2902 vdd.n940 185
R17255 vdd.n2901 vdd.n947 185
R17256 vdd.n3107 vdd.n947 185
R17257 vdd.n2900 vdd.n2899 185
R17258 vdd.n2899 vdd.n946 185
R17259 vdd.n2822 vdd.n952 185
R17260 vdd.n3101 vdd.n952 185
R17261 vdd.n3018 vdd.n3017 185
R17262 vdd.n3017 vdd.n3016 185
R17263 vdd.n3019 vdd.n958 185
R17264 vdd.n3095 vdd.n958 185
R17265 vdd.n3021 vdd.n3020 185
R17266 vdd.n3021 vdd.n957 185
R17267 vdd.n3092 vdd.n960 185
R17268 vdd.n960 vdd.n957 185
R17269 vdd.n3094 vdd.n3093 185
R17270 vdd.n3095 vdd.n3094 185
R17271 vdd.n951 vdd.n950 185
R17272 vdd.n3016 vdd.n951 185
R17273 vdd.n3103 vdd.n3102 185
R17274 vdd.n3102 vdd.n3101 185
R17275 vdd.n3104 vdd.n949 185
R17276 vdd.n949 vdd.n946 185
R17277 vdd.n3106 vdd.n3105 185
R17278 vdd.n3107 vdd.n3106 185
R17279 vdd.n939 vdd.n938 185
R17280 vdd.n940 vdd.n939 185
R17281 vdd.n3115 vdd.n3114 185
R17282 vdd.n3114 vdd.n3113 185
R17283 vdd.n3116 vdd.n937 185
R17284 vdd.n3004 vdd.n937 185
R17285 vdd.n3118 vdd.n3117 185
R17286 vdd.n3119 vdd.n3118 185
R17287 vdd.n928 vdd.n927 185
R17288 vdd.n2998 vdd.n928 185
R17289 vdd.n3127 vdd.n3126 185
R17290 vdd.n3126 vdd.n3125 185
R17291 vdd.n3128 vdd.n926 185
R17292 vdd.n931 vdd.n926 185
R17293 vdd.n3130 vdd.n3129 185
R17294 vdd.n3131 vdd.n3130 185
R17295 vdd.n917 vdd.n916 185
R17296 vdd.n925 vdd.n917 185
R17297 vdd.n3139 vdd.n3138 185
R17298 vdd.n3138 vdd.n3137 185
R17299 vdd.n3140 vdd.n915 185
R17300 vdd.n915 vdd.n912 185
R17301 vdd.n3142 vdd.n3141 185
R17302 vdd.n3143 vdd.n3142 185
R17303 vdd.n904 vdd.n903 185
R17304 vdd.n905 vdd.n904 185
R17305 vdd.n3152 vdd.n3151 185
R17306 vdd.n3151 vdd.n3150 185
R17307 vdd.n3153 vdd.n902 185
R17308 vdd.n908 vdd.n902 185
R17309 vdd.n3155 vdd.n3154 185
R17310 vdd.n3156 vdd.n3155 185
R17311 vdd.n892 vdd.n891 185
R17312 vdd.n901 vdd.n892 185
R17313 vdd.n3164 vdd.n3163 185
R17314 vdd.n3163 vdd.n3162 185
R17315 vdd.n3165 vdd.n890 185
R17316 vdd.n890 vdd.n887 185
R17317 vdd.n3167 vdd.n3166 185
R17318 vdd.n3168 vdd.n3167 185
R17319 vdd.n880 vdd.n879 185
R17320 vdd.n881 vdd.n880 185
R17321 vdd.n3176 vdd.n3175 185
R17322 vdd.n3175 vdd.n3174 185
R17323 vdd.n3177 vdd.n878 185
R17324 vdd.n878 vdd.n874 185
R17325 vdd.n3179 vdd.n3178 185
R17326 vdd.n3180 vdd.n3179 185
R17327 vdd.n867 vdd.n866 185
R17328 vdd.n877 vdd.n867 185
R17329 vdd.n3188 vdd.n3187 185
R17330 vdd.n3187 vdd.n3186 185
R17331 vdd.n3189 vdd.n865 185
R17332 vdd.n870 vdd.n865 185
R17333 vdd.n3191 vdd.n3190 185
R17334 vdd.n3192 vdd.n3191 185
R17335 vdd.n856 vdd.n855 185
R17336 vdd.n864 vdd.n856 185
R17337 vdd.n3200 vdd.n3199 185
R17338 vdd.n3199 vdd.n3198 185
R17339 vdd.n3201 vdd.n854 185
R17340 vdd.n854 vdd.n851 185
R17341 vdd.n3203 vdd.n3202 185
R17342 vdd.n3204 vdd.n3203 185
R17343 vdd.n842 vdd.n841 185
R17344 vdd.n843 vdd.n842 185
R17345 vdd.n3257 vdd.n3256 185
R17346 vdd.n3256 vdd.n3255 185
R17347 vdd.n3258 vdd.n840 185
R17348 vdd.n846 vdd.n840 185
R17349 vdd.n3260 vdd.n3259 185
R17350 vdd.n3261 vdd.n3260 185
R17351 vdd.n810 vdd.n808 185
R17352 vdd.n808 vdd.n805 185
R17353 vdd.n3330 vdd.n3329 185
R17354 vdd.n3331 vdd.n3330 185
R17355 vdd.n2711 vdd.n2710 185
R17356 vdd.n2712 vdd.n2711 185
R17357 vdd.n1009 vdd.n1007 185
R17358 vdd.n1007 vdd.n1005 185
R17359 vdd.n2626 vdd.n1016 185
R17360 vdd.n2637 vdd.n1016 185
R17361 vdd.n2627 vdd.n1025 185
R17362 vdd.n1399 vdd.n1025 185
R17363 vdd.n2629 vdd.n2628 185
R17364 vdd.n2630 vdd.n2629 185
R17365 vdd.n2625 vdd.n1024 185
R17366 vdd.n1024 vdd.n1021 185
R17367 vdd.n2624 vdd.n2623 185
R17368 vdd.n2623 vdd.n2622 185
R17369 vdd.n1027 vdd.n1026 185
R17370 vdd.n1028 vdd.n1027 185
R17371 vdd.n2615 vdd.n2614 185
R17372 vdd.n2616 vdd.n2615 185
R17373 vdd.n2613 vdd.n1036 185
R17374 vdd.n1425 vdd.n1036 185
R17375 vdd.n2612 vdd.n2611 185
R17376 vdd.n2611 vdd.n2610 185
R17377 vdd.n1038 vdd.n1037 185
R17378 vdd.n1046 vdd.n1038 185
R17379 vdd.n2603 vdd.n2602 185
R17380 vdd.n2604 vdd.n2603 185
R17381 vdd.n2601 vdd.n1047 185
R17382 vdd.n1052 vdd.n1047 185
R17383 vdd.n2600 vdd.n2599 185
R17384 vdd.n2599 vdd.n2598 185
R17385 vdd.n1049 vdd.n1048 185
R17386 vdd.n1437 vdd.n1049 185
R17387 vdd.n2591 vdd.n2590 185
R17388 vdd.n2592 vdd.n2591 185
R17389 vdd.n2589 vdd.n1059 185
R17390 vdd.n1059 vdd.n1056 185
R17391 vdd.n2588 vdd.n2587 185
R17392 vdd.n2587 vdd.n2586 185
R17393 vdd.n1061 vdd.n1060 185
R17394 vdd.n1062 vdd.n1061 185
R17395 vdd.n2579 vdd.n2578 185
R17396 vdd.n2580 vdd.n2579 185
R17397 vdd.n2576 vdd.n1070 185
R17398 vdd.n1076 vdd.n1070 185
R17399 vdd.n2575 vdd.n2574 185
R17400 vdd.n2574 vdd.n2573 185
R17401 vdd.n1073 vdd.n1072 185
R17402 vdd.n1083 vdd.n1073 185
R17403 vdd.n2566 vdd.n2565 185
R17404 vdd.n2567 vdd.n2566 185
R17405 vdd.n2564 vdd.n1084 185
R17406 vdd.n1084 vdd.n1080 185
R17407 vdd.n2563 vdd.n2562 185
R17408 vdd.n2562 vdd.n2561 185
R17409 vdd.n1086 vdd.n1085 185
R17410 vdd.n1087 vdd.n1086 185
R17411 vdd.n2554 vdd.n2553 185
R17412 vdd.n2555 vdd.n2554 185
R17413 vdd.n2552 vdd.n1096 185
R17414 vdd.n1096 vdd.n1093 185
R17415 vdd.n2551 vdd.n2550 185
R17416 vdd.n2550 vdd.n2549 185
R17417 vdd.n1098 vdd.n1097 185
R17418 vdd.n1106 vdd.n1098 185
R17419 vdd.n2542 vdd.n2541 185
R17420 vdd.n2543 vdd.n2542 185
R17421 vdd.n2540 vdd.n1107 185
R17422 vdd.n1112 vdd.n1107 185
R17423 vdd.n2539 vdd.n2538 185
R17424 vdd.n2538 vdd.n2537 185
R17425 vdd.n1109 vdd.n1108 185
R17426 vdd.n1119 vdd.n1109 185
R17427 vdd.n2530 vdd.n2529 185
R17428 vdd.n2531 vdd.n2530 185
R17429 vdd.n2528 vdd.n1120 185
R17430 vdd.n1120 vdd.n1116 185
R17431 vdd.n2527 vdd.n2526 185
R17432 vdd.n2526 vdd.n2525 185
R17433 vdd.n1122 vdd.n1121 185
R17434 vdd.n1123 vdd.n1122 185
R17435 vdd.n2518 vdd.n2517 185
R17436 vdd.n2519 vdd.n2518 185
R17437 vdd.n2516 vdd.n1131 185
R17438 vdd.n1137 vdd.n1131 185
R17439 vdd.n2515 vdd.n2514 185
R17440 vdd.n2514 vdd.n2513 185
R17441 vdd.n1133 vdd.n1132 185
R17442 vdd.n1134 vdd.n1133 185
R17443 vdd.n2642 vdd.n980 185
R17444 vdd.n2784 vdd.n980 185
R17445 vdd.n2644 vdd.n2643 185
R17446 vdd.n2646 vdd.n2645 185
R17447 vdd.n2648 vdd.n2647 185
R17448 vdd.n2650 vdd.n2649 185
R17449 vdd.n2652 vdd.n2651 185
R17450 vdd.n2654 vdd.n2653 185
R17451 vdd.n2656 vdd.n2655 185
R17452 vdd.n2658 vdd.n2657 185
R17453 vdd.n2660 vdd.n2659 185
R17454 vdd.n2662 vdd.n2661 185
R17455 vdd.n2664 vdd.n2663 185
R17456 vdd.n2666 vdd.n2665 185
R17457 vdd.n2668 vdd.n2667 185
R17458 vdd.n2670 vdd.n2669 185
R17459 vdd.n2672 vdd.n2671 185
R17460 vdd.n2674 vdd.n2673 185
R17461 vdd.n2676 vdd.n2675 185
R17462 vdd.n2678 vdd.n2677 185
R17463 vdd.n2680 vdd.n2679 185
R17464 vdd.n2682 vdd.n2681 185
R17465 vdd.n2684 vdd.n2683 185
R17466 vdd.n2686 vdd.n2685 185
R17467 vdd.n2688 vdd.n2687 185
R17468 vdd.n2690 vdd.n2689 185
R17469 vdd.n2692 vdd.n2691 185
R17470 vdd.n2694 vdd.n2693 185
R17471 vdd.n2696 vdd.n2695 185
R17472 vdd.n2698 vdd.n2697 185
R17473 vdd.n2700 vdd.n2699 185
R17474 vdd.n2702 vdd.n2701 185
R17475 vdd.n2704 vdd.n2703 185
R17476 vdd.n2706 vdd.n2705 185
R17477 vdd.n2708 vdd.n2707 185
R17478 vdd.n2709 vdd.n1008 185
R17479 vdd.n2641 vdd.n1006 185
R17480 vdd.n2712 vdd.n1006 185
R17481 vdd.n2640 vdd.n2639 185
R17482 vdd.n2639 vdd.n1005 185
R17483 vdd.n2638 vdd.n1013 185
R17484 vdd.n2638 vdd.n2637 185
R17485 vdd.n1415 vdd.n1014 185
R17486 vdd.n1399 vdd.n1014 185
R17487 vdd.n1416 vdd.n1023 185
R17488 vdd.n2630 vdd.n1023 185
R17489 vdd.n1418 vdd.n1417 185
R17490 vdd.n1417 vdd.n1021 185
R17491 vdd.n1419 vdd.n1030 185
R17492 vdd.n2622 vdd.n1030 185
R17493 vdd.n1421 vdd.n1420 185
R17494 vdd.n1420 vdd.n1028 185
R17495 vdd.n1422 vdd.n1035 185
R17496 vdd.n2616 vdd.n1035 185
R17497 vdd.n1424 vdd.n1423 185
R17498 vdd.n1425 vdd.n1424 185
R17499 vdd.n1414 vdd.n1040 185
R17500 vdd.n2610 vdd.n1040 185
R17501 vdd.n1413 vdd.n1412 185
R17502 vdd.n1412 vdd.n1046 185
R17503 vdd.n1411 vdd.n1045 185
R17504 vdd.n2604 vdd.n1045 185
R17505 vdd.n1410 vdd.n1409 185
R17506 vdd.n1409 vdd.n1052 185
R17507 vdd.n1318 vdd.n1051 185
R17508 vdd.n2598 vdd.n1051 185
R17509 vdd.n1439 vdd.n1438 185
R17510 vdd.n1438 vdd.n1437 185
R17511 vdd.n1440 vdd.n1058 185
R17512 vdd.n2592 vdd.n1058 185
R17513 vdd.n1442 vdd.n1441 185
R17514 vdd.n1441 vdd.n1056 185
R17515 vdd.n1443 vdd.n1064 185
R17516 vdd.n2586 vdd.n1064 185
R17517 vdd.n1445 vdd.n1444 185
R17518 vdd.n1444 vdd.n1062 185
R17519 vdd.n1446 vdd.n1069 185
R17520 vdd.n2580 vdd.n1069 185
R17521 vdd.n1448 vdd.n1447 185
R17522 vdd.n1447 vdd.n1076 185
R17523 vdd.n1449 vdd.n1075 185
R17524 vdd.n2573 vdd.n1075 185
R17525 vdd.n1451 vdd.n1450 185
R17526 vdd.n1450 vdd.n1083 185
R17527 vdd.n1452 vdd.n1082 185
R17528 vdd.n2567 vdd.n1082 185
R17529 vdd.n1454 vdd.n1453 185
R17530 vdd.n1453 vdd.n1080 185
R17531 vdd.n1455 vdd.n1089 185
R17532 vdd.n2561 vdd.n1089 185
R17533 vdd.n1457 vdd.n1456 185
R17534 vdd.n1456 vdd.n1087 185
R17535 vdd.n1458 vdd.n1095 185
R17536 vdd.n2555 vdd.n1095 185
R17537 vdd.n1460 vdd.n1459 185
R17538 vdd.n1459 vdd.n1093 185
R17539 vdd.n1461 vdd.n1100 185
R17540 vdd.n2549 vdd.n1100 185
R17541 vdd.n1463 vdd.n1462 185
R17542 vdd.n1462 vdd.n1106 185
R17543 vdd.n1464 vdd.n1105 185
R17544 vdd.n2543 vdd.n1105 185
R17545 vdd.n1466 vdd.n1465 185
R17546 vdd.n1465 vdd.n1112 185
R17547 vdd.n1467 vdd.n1111 185
R17548 vdd.n2537 vdd.n1111 185
R17549 vdd.n1469 vdd.n1468 185
R17550 vdd.n1468 vdd.n1119 185
R17551 vdd.n1470 vdd.n1118 185
R17552 vdd.n2531 vdd.n1118 185
R17553 vdd.n1472 vdd.n1471 185
R17554 vdd.n1471 vdd.n1116 185
R17555 vdd.n1473 vdd.n1125 185
R17556 vdd.n2525 vdd.n1125 185
R17557 vdd.n1475 vdd.n1474 185
R17558 vdd.n1474 vdd.n1123 185
R17559 vdd.n1476 vdd.n1130 185
R17560 vdd.n2519 vdd.n1130 185
R17561 vdd.n1478 vdd.n1477 185
R17562 vdd.n1477 vdd.n1137 185
R17563 vdd.n1479 vdd.n1136 185
R17564 vdd.n2513 vdd.n1136 185
R17565 vdd.n1481 vdd.n1480 185
R17566 vdd.n1480 vdd.n1134 185
R17567 vdd.n1281 vdd.n1280 185
R17568 vdd.n1283 vdd.n1282 185
R17569 vdd.n1285 vdd.n1284 185
R17570 vdd.n1287 vdd.n1286 185
R17571 vdd.n1289 vdd.n1288 185
R17572 vdd.n1291 vdd.n1290 185
R17573 vdd.n1293 vdd.n1292 185
R17574 vdd.n1295 vdd.n1294 185
R17575 vdd.n1297 vdd.n1296 185
R17576 vdd.n1299 vdd.n1298 185
R17577 vdd.n1301 vdd.n1300 185
R17578 vdd.n1303 vdd.n1302 185
R17579 vdd.n1305 vdd.n1304 185
R17580 vdd.n1307 vdd.n1306 185
R17581 vdd.n1309 vdd.n1308 185
R17582 vdd.n1311 vdd.n1310 185
R17583 vdd.n1313 vdd.n1312 185
R17584 vdd.n1515 vdd.n1314 185
R17585 vdd.n1514 vdd.n1513 185
R17586 vdd.n1512 vdd.n1511 185
R17587 vdd.n1510 vdd.n1509 185
R17588 vdd.n1508 vdd.n1507 185
R17589 vdd.n1506 vdd.n1505 185
R17590 vdd.n1504 vdd.n1503 185
R17591 vdd.n1502 vdd.n1501 185
R17592 vdd.n1500 vdd.n1499 185
R17593 vdd.n1498 vdd.n1497 185
R17594 vdd.n1496 vdd.n1495 185
R17595 vdd.n1494 vdd.n1493 185
R17596 vdd.n1492 vdd.n1491 185
R17597 vdd.n1490 vdd.n1489 185
R17598 vdd.n1488 vdd.n1487 185
R17599 vdd.n1486 vdd.n1485 185
R17600 vdd.n1484 vdd.n1483 185
R17601 vdd.n1482 vdd.n1175 185
R17602 vdd.n2506 vdd.n1175 185
R17603 vdd.n327 vdd.n326 171.744
R17604 vdd.n326 vdd.n325 171.744
R17605 vdd.n325 vdd.n294 171.744
R17606 vdd.n318 vdd.n294 171.744
R17607 vdd.n318 vdd.n317 171.744
R17608 vdd.n317 vdd.n299 171.744
R17609 vdd.n310 vdd.n299 171.744
R17610 vdd.n310 vdd.n309 171.744
R17611 vdd.n309 vdd.n303 171.744
R17612 vdd.n268 vdd.n267 171.744
R17613 vdd.n267 vdd.n266 171.744
R17614 vdd.n266 vdd.n235 171.744
R17615 vdd.n259 vdd.n235 171.744
R17616 vdd.n259 vdd.n258 171.744
R17617 vdd.n258 vdd.n240 171.744
R17618 vdd.n251 vdd.n240 171.744
R17619 vdd.n251 vdd.n250 171.744
R17620 vdd.n250 vdd.n244 171.744
R17621 vdd.n225 vdd.n224 171.744
R17622 vdd.n224 vdd.n223 171.744
R17623 vdd.n223 vdd.n192 171.744
R17624 vdd.n216 vdd.n192 171.744
R17625 vdd.n216 vdd.n215 171.744
R17626 vdd.n215 vdd.n197 171.744
R17627 vdd.n208 vdd.n197 171.744
R17628 vdd.n208 vdd.n207 171.744
R17629 vdd.n207 vdd.n201 171.744
R17630 vdd.n166 vdd.n165 171.744
R17631 vdd.n165 vdd.n164 171.744
R17632 vdd.n164 vdd.n133 171.744
R17633 vdd.n157 vdd.n133 171.744
R17634 vdd.n157 vdd.n156 171.744
R17635 vdd.n156 vdd.n138 171.744
R17636 vdd.n149 vdd.n138 171.744
R17637 vdd.n149 vdd.n148 171.744
R17638 vdd.n148 vdd.n142 171.744
R17639 vdd.n124 vdd.n123 171.744
R17640 vdd.n123 vdd.n122 171.744
R17641 vdd.n122 vdd.n91 171.744
R17642 vdd.n115 vdd.n91 171.744
R17643 vdd.n115 vdd.n114 171.744
R17644 vdd.n114 vdd.n96 171.744
R17645 vdd.n107 vdd.n96 171.744
R17646 vdd.n107 vdd.n106 171.744
R17647 vdd.n106 vdd.n100 171.744
R17648 vdd.n65 vdd.n64 171.744
R17649 vdd.n64 vdd.n63 171.744
R17650 vdd.n63 vdd.n32 171.744
R17651 vdd.n56 vdd.n32 171.744
R17652 vdd.n56 vdd.n55 171.744
R17653 vdd.n55 vdd.n37 171.744
R17654 vdd.n48 vdd.n37 171.744
R17655 vdd.n48 vdd.n47 171.744
R17656 vdd.n47 vdd.n41 171.744
R17657 vdd.n2201 vdd.n2200 171.744
R17658 vdd.n2200 vdd.n2199 171.744
R17659 vdd.n2199 vdd.n2168 171.744
R17660 vdd.n2192 vdd.n2168 171.744
R17661 vdd.n2192 vdd.n2191 171.744
R17662 vdd.n2191 vdd.n2173 171.744
R17663 vdd.n2184 vdd.n2173 171.744
R17664 vdd.n2184 vdd.n2183 171.744
R17665 vdd.n2183 vdd.n2177 171.744
R17666 vdd.n2260 vdd.n2259 171.744
R17667 vdd.n2259 vdd.n2258 171.744
R17668 vdd.n2258 vdd.n2227 171.744
R17669 vdd.n2251 vdd.n2227 171.744
R17670 vdd.n2251 vdd.n2250 171.744
R17671 vdd.n2250 vdd.n2232 171.744
R17672 vdd.n2243 vdd.n2232 171.744
R17673 vdd.n2243 vdd.n2242 171.744
R17674 vdd.n2242 vdd.n2236 171.744
R17675 vdd.n2099 vdd.n2098 171.744
R17676 vdd.n2098 vdd.n2097 171.744
R17677 vdd.n2097 vdd.n2066 171.744
R17678 vdd.n2090 vdd.n2066 171.744
R17679 vdd.n2090 vdd.n2089 171.744
R17680 vdd.n2089 vdd.n2071 171.744
R17681 vdd.n2082 vdd.n2071 171.744
R17682 vdd.n2082 vdd.n2081 171.744
R17683 vdd.n2081 vdd.n2075 171.744
R17684 vdd.n2158 vdd.n2157 171.744
R17685 vdd.n2157 vdd.n2156 171.744
R17686 vdd.n2156 vdd.n2125 171.744
R17687 vdd.n2149 vdd.n2125 171.744
R17688 vdd.n2149 vdd.n2148 171.744
R17689 vdd.n2148 vdd.n2130 171.744
R17690 vdd.n2141 vdd.n2130 171.744
R17691 vdd.n2141 vdd.n2140 171.744
R17692 vdd.n2140 vdd.n2134 171.744
R17693 vdd.n1998 vdd.n1997 171.744
R17694 vdd.n1997 vdd.n1996 171.744
R17695 vdd.n1996 vdd.n1965 171.744
R17696 vdd.n1989 vdd.n1965 171.744
R17697 vdd.n1989 vdd.n1988 171.744
R17698 vdd.n1988 vdd.n1970 171.744
R17699 vdd.n1981 vdd.n1970 171.744
R17700 vdd.n1981 vdd.n1980 171.744
R17701 vdd.n1980 vdd.n1974 171.744
R17702 vdd.n2057 vdd.n2056 171.744
R17703 vdd.n2056 vdd.n2055 171.744
R17704 vdd.n2055 vdd.n2024 171.744
R17705 vdd.n2048 vdd.n2024 171.744
R17706 vdd.n2048 vdd.n2047 171.744
R17707 vdd.n2047 vdd.n2029 171.744
R17708 vdd.n2040 vdd.n2029 171.744
R17709 vdd.n2040 vdd.n2039 171.744
R17710 vdd.n2039 vdd.n2033 171.744
R17711 vdd.n468 vdd.n467 146.341
R17712 vdd.n474 vdd.n473 146.341
R17713 vdd.n478 vdd.n477 146.341
R17714 vdd.n484 vdd.n483 146.341
R17715 vdd.n488 vdd.n487 146.341
R17716 vdd.n494 vdd.n493 146.341
R17717 vdd.n498 vdd.n497 146.341
R17718 vdd.n504 vdd.n503 146.341
R17719 vdd.n508 vdd.n507 146.341
R17720 vdd.n514 vdd.n513 146.341
R17721 vdd.n518 vdd.n517 146.341
R17722 vdd.n524 vdd.n523 146.341
R17723 vdd.n528 vdd.n527 146.341
R17724 vdd.n534 vdd.n533 146.341
R17725 vdd.n538 vdd.n537 146.341
R17726 vdd.n544 vdd.n543 146.341
R17727 vdd.n548 vdd.n547 146.341
R17728 vdd.n554 vdd.n553 146.341
R17729 vdd.n558 vdd.n557 146.341
R17730 vdd.n564 vdd.n563 146.341
R17731 vdd.n568 vdd.n567 146.341
R17732 vdd.n574 vdd.n573 146.341
R17733 vdd.n578 vdd.n577 146.341
R17734 vdd.n584 vdd.n583 146.341
R17735 vdd.n588 vdd.n587 146.341
R17736 vdd.n594 vdd.n593 146.341
R17737 vdd.n598 vdd.n597 146.341
R17738 vdd.n604 vdd.n603 146.341
R17739 vdd.n608 vdd.n607 146.341
R17740 vdd.n614 vdd.n613 146.341
R17741 vdd.n616 vdd.n425 146.341
R17742 vdd.n3502 vdd.n685 146.341
R17743 vdd.n3502 vdd.n677 146.341
R17744 vdd.n3512 vdd.n677 146.341
R17745 vdd.n3512 vdd.n673 146.341
R17746 vdd.n3518 vdd.n673 146.341
R17747 vdd.n3518 vdd.n667 146.341
R17748 vdd.n3529 vdd.n667 146.341
R17749 vdd.n3529 vdd.n663 146.341
R17750 vdd.n3535 vdd.n663 146.341
R17751 vdd.n3535 vdd.n654 146.341
R17752 vdd.n3545 vdd.n654 146.341
R17753 vdd.n3545 vdd.n650 146.341
R17754 vdd.n3551 vdd.n650 146.341
R17755 vdd.n3551 vdd.n643 146.341
R17756 vdd.n3562 vdd.n643 146.341
R17757 vdd.n3562 vdd.n639 146.341
R17758 vdd.n3571 vdd.n639 146.341
R17759 vdd.n3571 vdd.n632 146.341
R17760 vdd.n3581 vdd.n632 146.341
R17761 vdd.n3582 vdd.n3581 146.341
R17762 vdd.n3582 vdd.n341 146.341
R17763 vdd.n342 vdd.n341 146.341
R17764 vdd.n343 vdd.n342 146.341
R17765 vdd.n3589 vdd.n343 146.341
R17766 vdd.n3589 vdd.n351 146.341
R17767 vdd.n352 vdd.n351 146.341
R17768 vdd.n353 vdd.n352 146.341
R17769 vdd.n3596 vdd.n353 146.341
R17770 vdd.n3596 vdd.n362 146.341
R17771 vdd.n363 vdd.n362 146.341
R17772 vdd.n364 vdd.n363 146.341
R17773 vdd.n3604 vdd.n364 146.341
R17774 vdd.n3604 vdd.n372 146.341
R17775 vdd.n373 vdd.n372 146.341
R17776 vdd.n374 vdd.n373 146.341
R17777 vdd.n3611 vdd.n374 146.341
R17778 vdd.n3611 vdd.n383 146.341
R17779 vdd.n384 vdd.n383 146.341
R17780 vdd.n385 vdd.n384 146.341
R17781 vdd.n3618 vdd.n385 146.341
R17782 vdd.n3618 vdd.n393 146.341
R17783 vdd.n725 vdd.n724 146.341
R17784 vdd.n728 vdd.n724 146.341
R17785 vdd.n734 vdd.n733 146.341
R17786 vdd.n3484 vdd.n3483 146.341
R17787 vdd.n3480 vdd.n3479 146.341
R17788 vdd.n3476 vdd.n3475 146.341
R17789 vdd.n3472 vdd.n3471 146.341
R17790 vdd.n3468 vdd.n3467 146.341
R17791 vdd.n3464 vdd.n3463 146.341
R17792 vdd.n3460 vdd.n3459 146.341
R17793 vdd.n3451 vdd.n3450 146.341
R17794 vdd.n3448 vdd.n3447 146.341
R17795 vdd.n3444 vdd.n3443 146.341
R17796 vdd.n3440 vdd.n3439 146.341
R17797 vdd.n3436 vdd.n3435 146.341
R17798 vdd.n3432 vdd.n3431 146.341
R17799 vdd.n3428 vdd.n3427 146.341
R17800 vdd.n3424 vdd.n3423 146.341
R17801 vdd.n3420 vdd.n3419 146.341
R17802 vdd.n3416 vdd.n3415 146.341
R17803 vdd.n3412 vdd.n3411 146.341
R17804 vdd.n3405 vdd.n3404 146.341
R17805 vdd.n3402 vdd.n3401 146.341
R17806 vdd.n3398 vdd.n3397 146.341
R17807 vdd.n3394 vdd.n3393 146.341
R17808 vdd.n3390 vdd.n3389 146.341
R17809 vdd.n3386 vdd.n3385 146.341
R17810 vdd.n3382 vdd.n3381 146.341
R17811 vdd.n3378 vdd.n3377 146.341
R17812 vdd.n3374 vdd.n3373 146.341
R17813 vdd.n3370 vdd.n3369 146.341
R17814 vdd.n3496 vdd.n691 146.341
R17815 vdd.n3504 vdd.n684 146.341
R17816 vdd.n3504 vdd.n680 146.341
R17817 vdd.n3510 vdd.n680 146.341
R17818 vdd.n3510 vdd.n672 146.341
R17819 vdd.n3521 vdd.n672 146.341
R17820 vdd.n3521 vdd.n668 146.341
R17821 vdd.n3527 vdd.n668 146.341
R17822 vdd.n3527 vdd.n661 146.341
R17823 vdd.n3537 vdd.n661 146.341
R17824 vdd.n3537 vdd.n657 146.341
R17825 vdd.n3543 vdd.n657 146.341
R17826 vdd.n3543 vdd.n649 146.341
R17827 vdd.n3554 vdd.n649 146.341
R17828 vdd.n3554 vdd.n645 146.341
R17829 vdd.n3560 vdd.n645 146.341
R17830 vdd.n3560 vdd.n638 146.341
R17831 vdd.n3573 vdd.n638 146.341
R17832 vdd.n3573 vdd.n634 146.341
R17833 vdd.n3579 vdd.n634 146.341
R17834 vdd.n3579 vdd.n338 146.341
R17835 vdd.n3668 vdd.n338 146.341
R17836 vdd.n3668 vdd.n339 146.341
R17837 vdd.n3664 vdd.n339 146.341
R17838 vdd.n3664 vdd.n345 146.341
R17839 vdd.n3660 vdd.n345 146.341
R17840 vdd.n3660 vdd.n350 146.341
R17841 vdd.n3656 vdd.n350 146.341
R17842 vdd.n3656 vdd.n354 146.341
R17843 vdd.n3652 vdd.n354 146.341
R17844 vdd.n3652 vdd.n360 146.341
R17845 vdd.n3648 vdd.n360 146.341
R17846 vdd.n3648 vdd.n365 146.341
R17847 vdd.n3644 vdd.n365 146.341
R17848 vdd.n3644 vdd.n371 146.341
R17849 vdd.n3640 vdd.n371 146.341
R17850 vdd.n3640 vdd.n376 146.341
R17851 vdd.n3636 vdd.n376 146.341
R17852 vdd.n3636 vdd.n382 146.341
R17853 vdd.n3632 vdd.n382 146.341
R17854 vdd.n3632 vdd.n387 146.341
R17855 vdd.n3628 vdd.n387 146.341
R17856 vdd.n2471 vdd.n2470 146.341
R17857 vdd.n2468 vdd.n2465 146.341
R17858 vdd.n2463 vdd.n1185 146.341
R17859 vdd.n2459 vdd.n2458 146.341
R17860 vdd.n2456 vdd.n1189 146.341
R17861 vdd.n2452 vdd.n2451 146.341
R17862 vdd.n2449 vdd.n1196 146.341
R17863 vdd.n2445 vdd.n2444 146.341
R17864 vdd.n2442 vdd.n1203 146.341
R17865 vdd.n1214 vdd.n1211 146.341
R17866 vdd.n2434 vdd.n2433 146.341
R17867 vdd.n2431 vdd.n1216 146.341
R17868 vdd.n2427 vdd.n2426 146.341
R17869 vdd.n2424 vdd.n1222 146.341
R17870 vdd.n2420 vdd.n2419 146.341
R17871 vdd.n2417 vdd.n1229 146.341
R17872 vdd.n2413 vdd.n2412 146.341
R17873 vdd.n2410 vdd.n1236 146.341
R17874 vdd.n2406 vdd.n2405 146.341
R17875 vdd.n2403 vdd.n1243 146.341
R17876 vdd.n1254 vdd.n1251 146.341
R17877 vdd.n2395 vdd.n2394 146.341
R17878 vdd.n2392 vdd.n1256 146.341
R17879 vdd.n2388 vdd.n2387 146.341
R17880 vdd.n2385 vdd.n1262 146.341
R17881 vdd.n2381 vdd.n2380 146.341
R17882 vdd.n2378 vdd.n1269 146.341
R17883 vdd.n2374 vdd.n2373 146.341
R17884 vdd.n2371 vdd.n1276 146.341
R17885 vdd.n1522 vdd.n1520 146.341
R17886 vdd.n1525 vdd.n1524 146.341
R17887 vdd.n1883 vdd.n1643 146.341
R17888 vdd.n1883 vdd.n1639 146.341
R17889 vdd.n1889 vdd.n1639 146.341
R17890 vdd.n1889 vdd.n1631 146.341
R17891 vdd.n1900 vdd.n1631 146.341
R17892 vdd.n1900 vdd.n1627 146.341
R17893 vdd.n1906 vdd.n1627 146.341
R17894 vdd.n1906 vdd.n1621 146.341
R17895 vdd.n1917 vdd.n1621 146.341
R17896 vdd.n1917 vdd.n1617 146.341
R17897 vdd.n1923 vdd.n1617 146.341
R17898 vdd.n1923 vdd.n1608 146.341
R17899 vdd.n1933 vdd.n1608 146.341
R17900 vdd.n1933 vdd.n1604 146.341
R17901 vdd.n1939 vdd.n1604 146.341
R17902 vdd.n1939 vdd.n1597 146.341
R17903 vdd.n1950 vdd.n1597 146.341
R17904 vdd.n1950 vdd.n1593 146.341
R17905 vdd.n1956 vdd.n1593 146.341
R17906 vdd.n1956 vdd.n1586 146.341
R17907 vdd.n2273 vdd.n1586 146.341
R17908 vdd.n2273 vdd.n1582 146.341
R17909 vdd.n2279 vdd.n1582 146.341
R17910 vdd.n2279 vdd.n1574 146.341
R17911 vdd.n2290 vdd.n1574 146.341
R17912 vdd.n2290 vdd.n1570 146.341
R17913 vdd.n2296 vdd.n1570 146.341
R17914 vdd.n2296 vdd.n1564 146.341
R17915 vdd.n2307 vdd.n1564 146.341
R17916 vdd.n2307 vdd.n1560 146.341
R17917 vdd.n2313 vdd.n1560 146.341
R17918 vdd.n2313 vdd.n1551 146.341
R17919 vdd.n2323 vdd.n1551 146.341
R17920 vdd.n2323 vdd.n1547 146.341
R17921 vdd.n2329 vdd.n1547 146.341
R17922 vdd.n2329 vdd.n1541 146.341
R17923 vdd.n2340 vdd.n1541 146.341
R17924 vdd.n2340 vdd.n1536 146.341
R17925 vdd.n2348 vdd.n1536 146.341
R17926 vdd.n2348 vdd.n1527 146.341
R17927 vdd.n2359 vdd.n1527 146.341
R17928 vdd.n1872 vdd.n1648 146.341
R17929 vdd.n1872 vdd.n1681 146.341
R17930 vdd.n1685 vdd.n1684 146.341
R17931 vdd.n1687 vdd.n1686 146.341
R17932 vdd.n1691 vdd.n1690 146.341
R17933 vdd.n1693 vdd.n1692 146.341
R17934 vdd.n1697 vdd.n1696 146.341
R17935 vdd.n1699 vdd.n1698 146.341
R17936 vdd.n1703 vdd.n1702 146.341
R17937 vdd.n1705 vdd.n1704 146.341
R17938 vdd.n1711 vdd.n1710 146.341
R17939 vdd.n1713 vdd.n1712 146.341
R17940 vdd.n1717 vdd.n1716 146.341
R17941 vdd.n1719 vdd.n1718 146.341
R17942 vdd.n1723 vdd.n1722 146.341
R17943 vdd.n1725 vdd.n1724 146.341
R17944 vdd.n1729 vdd.n1728 146.341
R17945 vdd.n1731 vdd.n1730 146.341
R17946 vdd.n1735 vdd.n1734 146.341
R17947 vdd.n1737 vdd.n1736 146.341
R17948 vdd.n1809 vdd.n1740 146.341
R17949 vdd.n1742 vdd.n1741 146.341
R17950 vdd.n1746 vdd.n1745 146.341
R17951 vdd.n1748 vdd.n1747 146.341
R17952 vdd.n1752 vdd.n1751 146.341
R17953 vdd.n1754 vdd.n1753 146.341
R17954 vdd.n1758 vdd.n1757 146.341
R17955 vdd.n1760 vdd.n1759 146.341
R17956 vdd.n1764 vdd.n1763 146.341
R17957 vdd.n1766 vdd.n1765 146.341
R17958 vdd.n1770 vdd.n1769 146.341
R17959 vdd.n1771 vdd.n1679 146.341
R17960 vdd.n1881 vdd.n1644 146.341
R17961 vdd.n1881 vdd.n1637 146.341
R17962 vdd.n1892 vdd.n1637 146.341
R17963 vdd.n1892 vdd.n1633 146.341
R17964 vdd.n1898 vdd.n1633 146.341
R17965 vdd.n1898 vdd.n1626 146.341
R17966 vdd.n1909 vdd.n1626 146.341
R17967 vdd.n1909 vdd.n1622 146.341
R17968 vdd.n1915 vdd.n1622 146.341
R17969 vdd.n1915 vdd.n1615 146.341
R17970 vdd.n1925 vdd.n1615 146.341
R17971 vdd.n1925 vdd.n1611 146.341
R17972 vdd.n1931 vdd.n1611 146.341
R17973 vdd.n1931 vdd.n1603 146.341
R17974 vdd.n1942 vdd.n1603 146.341
R17975 vdd.n1942 vdd.n1599 146.341
R17976 vdd.n1948 vdd.n1599 146.341
R17977 vdd.n1948 vdd.n1592 146.341
R17978 vdd.n1958 vdd.n1592 146.341
R17979 vdd.n1958 vdd.n1588 146.341
R17980 vdd.n2271 vdd.n1588 146.341
R17981 vdd.n2271 vdd.n1580 146.341
R17982 vdd.n2282 vdd.n1580 146.341
R17983 vdd.n2282 vdd.n1576 146.341
R17984 vdd.n2288 vdd.n1576 146.341
R17985 vdd.n2288 vdd.n1569 146.341
R17986 vdd.n2299 vdd.n1569 146.341
R17987 vdd.n2299 vdd.n1565 146.341
R17988 vdd.n2305 vdd.n1565 146.341
R17989 vdd.n2305 vdd.n1558 146.341
R17990 vdd.n2315 vdd.n1558 146.341
R17991 vdd.n2315 vdd.n1554 146.341
R17992 vdd.n2321 vdd.n1554 146.341
R17993 vdd.n2321 vdd.n1546 146.341
R17994 vdd.n2332 vdd.n1546 146.341
R17995 vdd.n2332 vdd.n1542 146.341
R17996 vdd.n2338 vdd.n1542 146.341
R17997 vdd.n2338 vdd.n1534 146.341
R17998 vdd.n2351 vdd.n1534 146.341
R17999 vdd.n2351 vdd.n1529 146.341
R18000 vdd.n2357 vdd.n1529 146.341
R18001 vdd.n1315 vdd.t15 127.284
R18002 vdd.n1010 vdd.t55 127.284
R18003 vdd.n1319 vdd.t52 127.284
R18004 vdd.n1001 vdd.t76 127.284
R18005 vdd.n896 vdd.t39 127.284
R18006 vdd.n896 vdd.t40 127.284
R18007 vdd.n2823 vdd.t70 127.284
R18008 vdd.n832 vdd.t31 127.284
R18009 vdd.n2820 vdd.t63 127.284
R18010 vdd.n799 vdd.t10 127.284
R18011 vdd.n1071 vdd.t66 127.284
R18012 vdd.n1071 vdd.t67 127.284
R18013 vdd.n22 vdd.n20 117.314
R18014 vdd.n17 vdd.n15 117.314
R18015 vdd.n27 vdd.n26 116.927
R18016 vdd.n24 vdd.n23 116.927
R18017 vdd.n22 vdd.n21 116.927
R18018 vdd.n17 vdd.n16 116.927
R18019 vdd.n19 vdd.n18 116.927
R18020 vdd.n27 vdd.n25 116.927
R18021 vdd.n1316 vdd.t14 111.188
R18022 vdd.n1011 vdd.t56 111.188
R18023 vdd.n1320 vdd.t51 111.188
R18024 vdd.n1002 vdd.t77 111.188
R18025 vdd.n2824 vdd.t69 111.188
R18026 vdd.n833 vdd.t32 111.188
R18027 vdd.n2821 vdd.t62 111.188
R18028 vdd.n800 vdd.t11 111.188
R18029 vdd.n3094 vdd.n960 99.5127
R18030 vdd.n3094 vdd.n951 99.5127
R18031 vdd.n3102 vdd.n951 99.5127
R18032 vdd.n3102 vdd.n949 99.5127
R18033 vdd.n3106 vdd.n949 99.5127
R18034 vdd.n3106 vdd.n939 99.5127
R18035 vdd.n3114 vdd.n939 99.5127
R18036 vdd.n3114 vdd.n937 99.5127
R18037 vdd.n3118 vdd.n937 99.5127
R18038 vdd.n3118 vdd.n928 99.5127
R18039 vdd.n3126 vdd.n928 99.5127
R18040 vdd.n3126 vdd.n926 99.5127
R18041 vdd.n3130 vdd.n926 99.5127
R18042 vdd.n3130 vdd.n917 99.5127
R18043 vdd.n3138 vdd.n917 99.5127
R18044 vdd.n3138 vdd.n915 99.5127
R18045 vdd.n3142 vdd.n915 99.5127
R18046 vdd.n3142 vdd.n904 99.5127
R18047 vdd.n3151 vdd.n904 99.5127
R18048 vdd.n3151 vdd.n902 99.5127
R18049 vdd.n3155 vdd.n902 99.5127
R18050 vdd.n3155 vdd.n892 99.5127
R18051 vdd.n3163 vdd.n892 99.5127
R18052 vdd.n3163 vdd.n890 99.5127
R18053 vdd.n3167 vdd.n890 99.5127
R18054 vdd.n3167 vdd.n880 99.5127
R18055 vdd.n3175 vdd.n880 99.5127
R18056 vdd.n3175 vdd.n878 99.5127
R18057 vdd.n3179 vdd.n878 99.5127
R18058 vdd.n3179 vdd.n867 99.5127
R18059 vdd.n3187 vdd.n867 99.5127
R18060 vdd.n3187 vdd.n865 99.5127
R18061 vdd.n3191 vdd.n865 99.5127
R18062 vdd.n3191 vdd.n856 99.5127
R18063 vdd.n3199 vdd.n856 99.5127
R18064 vdd.n3199 vdd.n854 99.5127
R18065 vdd.n3203 vdd.n854 99.5127
R18066 vdd.n3203 vdd.n842 99.5127
R18067 vdd.n3256 vdd.n842 99.5127
R18068 vdd.n3256 vdd.n840 99.5127
R18069 vdd.n3260 vdd.n840 99.5127
R18070 vdd.n3260 vdd.n808 99.5127
R18071 vdd.n3330 vdd.n808 99.5127
R18072 vdd.n3326 vdd.n809 99.5127
R18073 vdd.n3324 vdd.n3323 99.5127
R18074 vdd.n3321 vdd.n813 99.5127
R18075 vdd.n3317 vdd.n3316 99.5127
R18076 vdd.n3314 vdd.n816 99.5127
R18077 vdd.n3310 vdd.n3309 99.5127
R18078 vdd.n3307 vdd.n819 99.5127
R18079 vdd.n3303 vdd.n3302 99.5127
R18080 vdd.n3300 vdd.n3298 99.5127
R18081 vdd.n3296 vdd.n822 99.5127
R18082 vdd.n3292 vdd.n3291 99.5127
R18083 vdd.n3289 vdd.n825 99.5127
R18084 vdd.n3285 vdd.n3284 99.5127
R18085 vdd.n3282 vdd.n828 99.5127
R18086 vdd.n3278 vdd.n3277 99.5127
R18087 vdd.n3275 vdd.n831 99.5127
R18088 vdd.n3270 vdd.n3269 99.5127
R18089 vdd.n3021 vdd.n958 99.5127
R18090 vdd.n3017 vdd.n958 99.5127
R18091 vdd.n3017 vdd.n952 99.5127
R18092 vdd.n2899 vdd.n952 99.5127
R18093 vdd.n2899 vdd.n947 99.5127
R18094 vdd.n2902 vdd.n947 99.5127
R18095 vdd.n2902 vdd.n941 99.5127
R18096 vdd.n3003 vdd.n941 99.5127
R18097 vdd.n3003 vdd.n935 99.5127
R18098 vdd.n2999 vdd.n935 99.5127
R18099 vdd.n2999 vdd.n929 99.5127
R18100 vdd.n2946 vdd.n929 99.5127
R18101 vdd.n2946 vdd.n923 99.5127
R18102 vdd.n2943 vdd.n923 99.5127
R18103 vdd.n2943 vdd.n918 99.5127
R18104 vdd.n2940 vdd.n918 99.5127
R18105 vdd.n2940 vdd.n913 99.5127
R18106 vdd.n2937 vdd.n913 99.5127
R18107 vdd.n2937 vdd.n906 99.5127
R18108 vdd.n2934 vdd.n906 99.5127
R18109 vdd.n2934 vdd.n899 99.5127
R18110 vdd.n2931 vdd.n899 99.5127
R18111 vdd.n2931 vdd.n893 99.5127
R18112 vdd.n2928 vdd.n893 99.5127
R18113 vdd.n2928 vdd.n888 99.5127
R18114 vdd.n2925 vdd.n888 99.5127
R18115 vdd.n2925 vdd.n882 99.5127
R18116 vdd.n2922 vdd.n882 99.5127
R18117 vdd.n2922 vdd.n875 99.5127
R18118 vdd.n2919 vdd.n875 99.5127
R18119 vdd.n2919 vdd.n868 99.5127
R18120 vdd.n2916 vdd.n868 99.5127
R18121 vdd.n2916 vdd.n862 99.5127
R18122 vdd.n2913 vdd.n862 99.5127
R18123 vdd.n2913 vdd.n857 99.5127
R18124 vdd.n2910 vdd.n857 99.5127
R18125 vdd.n2910 vdd.n852 99.5127
R18126 vdd.n2907 vdd.n852 99.5127
R18127 vdd.n2907 vdd.n844 99.5127
R18128 vdd.n844 vdd.n837 99.5127
R18129 vdd.n3262 vdd.n837 99.5127
R18130 vdd.n3263 vdd.n3262 99.5127
R18131 vdd.n3263 vdd.n806 99.5127
R18132 vdd.n3087 vdd.n962 99.5127
R18133 vdd.n3087 vdd.n2819 99.5127
R18134 vdd.n3083 vdd.n3082 99.5127
R18135 vdd.n3079 vdd.n3078 99.5127
R18136 vdd.n3075 vdd.n3074 99.5127
R18137 vdd.n3071 vdd.n3070 99.5127
R18138 vdd.n3067 vdd.n3066 99.5127
R18139 vdd.n3063 vdd.n3062 99.5127
R18140 vdd.n3059 vdd.n3058 99.5127
R18141 vdd.n3055 vdd.n3054 99.5127
R18142 vdd.n3051 vdd.n3050 99.5127
R18143 vdd.n3047 vdd.n3046 99.5127
R18144 vdd.n3043 vdd.n3042 99.5127
R18145 vdd.n3039 vdd.n3038 99.5127
R18146 vdd.n3035 vdd.n3034 99.5127
R18147 vdd.n3031 vdd.n3030 99.5127
R18148 vdd.n3026 vdd.n3025 99.5127
R18149 vdd.n2783 vdd.n999 99.5127
R18150 vdd.n2779 vdd.n2778 99.5127
R18151 vdd.n2775 vdd.n2774 99.5127
R18152 vdd.n2771 vdd.n2770 99.5127
R18153 vdd.n2767 vdd.n2766 99.5127
R18154 vdd.n2763 vdd.n2762 99.5127
R18155 vdd.n2759 vdd.n2758 99.5127
R18156 vdd.n2755 vdd.n2754 99.5127
R18157 vdd.n2751 vdd.n2750 99.5127
R18158 vdd.n2747 vdd.n2746 99.5127
R18159 vdd.n2743 vdd.n2742 99.5127
R18160 vdd.n2739 vdd.n2738 99.5127
R18161 vdd.n2735 vdd.n2734 99.5127
R18162 vdd.n2731 vdd.n2730 99.5127
R18163 vdd.n2727 vdd.n2726 99.5127
R18164 vdd.n2723 vdd.n2722 99.5127
R18165 vdd.n2718 vdd.n2717 99.5127
R18166 vdd.n1355 vdd.n1135 99.5127
R18167 vdd.n1358 vdd.n1135 99.5127
R18168 vdd.n1358 vdd.n1129 99.5127
R18169 vdd.n1361 vdd.n1129 99.5127
R18170 vdd.n1361 vdd.n1124 99.5127
R18171 vdd.n1364 vdd.n1124 99.5127
R18172 vdd.n1364 vdd.n1117 99.5127
R18173 vdd.n1367 vdd.n1117 99.5127
R18174 vdd.n1367 vdd.n1110 99.5127
R18175 vdd.n1370 vdd.n1110 99.5127
R18176 vdd.n1370 vdd.n1104 99.5127
R18177 vdd.n1373 vdd.n1104 99.5127
R18178 vdd.n1373 vdd.n1099 99.5127
R18179 vdd.n1376 vdd.n1099 99.5127
R18180 vdd.n1376 vdd.n1094 99.5127
R18181 vdd.n1379 vdd.n1094 99.5127
R18182 vdd.n1379 vdd.n1088 99.5127
R18183 vdd.n1382 vdd.n1088 99.5127
R18184 vdd.n1382 vdd.n1081 99.5127
R18185 vdd.n1385 vdd.n1081 99.5127
R18186 vdd.n1385 vdd.n1074 99.5127
R18187 vdd.n1388 vdd.n1074 99.5127
R18188 vdd.n1388 vdd.n1068 99.5127
R18189 vdd.n1391 vdd.n1068 99.5127
R18190 vdd.n1391 vdd.n1063 99.5127
R18191 vdd.n1394 vdd.n1063 99.5127
R18192 vdd.n1394 vdd.n1057 99.5127
R18193 vdd.n1436 vdd.n1057 99.5127
R18194 vdd.n1436 vdd.n1050 99.5127
R18195 vdd.n1432 vdd.n1050 99.5127
R18196 vdd.n1432 vdd.n1044 99.5127
R18197 vdd.n1429 vdd.n1044 99.5127
R18198 vdd.n1429 vdd.n1039 99.5127
R18199 vdd.n1426 vdd.n1039 99.5127
R18200 vdd.n1426 vdd.n1034 99.5127
R18201 vdd.n1406 vdd.n1034 99.5127
R18202 vdd.n1406 vdd.n1029 99.5127
R18203 vdd.n1403 vdd.n1029 99.5127
R18204 vdd.n1403 vdd.n1022 99.5127
R18205 vdd.n1400 vdd.n1022 99.5127
R18206 vdd.n1400 vdd.n1015 99.5127
R18207 vdd.n1015 vdd.n1004 99.5127
R18208 vdd.n2713 vdd.n1004 99.5127
R18209 vdd.n2505 vdd.n1140 99.5127
R18210 vdd.n2505 vdd.n1176 99.5127
R18211 vdd.n2501 vdd.n2500 99.5127
R18212 vdd.n2497 vdd.n2496 99.5127
R18213 vdd.n2493 vdd.n2492 99.5127
R18214 vdd.n2489 vdd.n2488 99.5127
R18215 vdd.n2485 vdd.n2484 99.5127
R18216 vdd.n2481 vdd.n2480 99.5127
R18217 vdd.n2477 vdd.n2476 99.5127
R18218 vdd.n1322 vdd.n1321 99.5127
R18219 vdd.n1326 vdd.n1325 99.5127
R18220 vdd.n1330 vdd.n1329 99.5127
R18221 vdd.n1334 vdd.n1333 99.5127
R18222 vdd.n1338 vdd.n1337 99.5127
R18223 vdd.n1342 vdd.n1341 99.5127
R18224 vdd.n1346 vdd.n1345 99.5127
R18225 vdd.n1351 vdd.n1350 99.5127
R18226 vdd.n2512 vdd.n1138 99.5127
R18227 vdd.n2512 vdd.n1128 99.5127
R18228 vdd.n2520 vdd.n1128 99.5127
R18229 vdd.n2520 vdd.n1126 99.5127
R18230 vdd.n2524 vdd.n1126 99.5127
R18231 vdd.n2524 vdd.n1115 99.5127
R18232 vdd.n2532 vdd.n1115 99.5127
R18233 vdd.n2532 vdd.n1113 99.5127
R18234 vdd.n2536 vdd.n1113 99.5127
R18235 vdd.n2536 vdd.n1103 99.5127
R18236 vdd.n2544 vdd.n1103 99.5127
R18237 vdd.n2544 vdd.n1101 99.5127
R18238 vdd.n2548 vdd.n1101 99.5127
R18239 vdd.n2548 vdd.n1092 99.5127
R18240 vdd.n2556 vdd.n1092 99.5127
R18241 vdd.n2556 vdd.n1090 99.5127
R18242 vdd.n2560 vdd.n1090 99.5127
R18243 vdd.n2560 vdd.n1079 99.5127
R18244 vdd.n2568 vdd.n1079 99.5127
R18245 vdd.n2568 vdd.n1077 99.5127
R18246 vdd.n2572 vdd.n1077 99.5127
R18247 vdd.n2572 vdd.n1067 99.5127
R18248 vdd.n2581 vdd.n1067 99.5127
R18249 vdd.n2581 vdd.n1065 99.5127
R18250 vdd.n2585 vdd.n1065 99.5127
R18251 vdd.n2585 vdd.n1055 99.5127
R18252 vdd.n2593 vdd.n1055 99.5127
R18253 vdd.n2593 vdd.n1053 99.5127
R18254 vdd.n2597 vdd.n1053 99.5127
R18255 vdd.n2597 vdd.n1043 99.5127
R18256 vdd.n2605 vdd.n1043 99.5127
R18257 vdd.n2605 vdd.n1041 99.5127
R18258 vdd.n2609 vdd.n1041 99.5127
R18259 vdd.n2609 vdd.n1033 99.5127
R18260 vdd.n2617 vdd.n1033 99.5127
R18261 vdd.n2617 vdd.n1031 99.5127
R18262 vdd.n2621 vdd.n1031 99.5127
R18263 vdd.n2621 vdd.n1020 99.5127
R18264 vdd.n2631 vdd.n1020 99.5127
R18265 vdd.n2631 vdd.n1017 99.5127
R18266 vdd.n2636 vdd.n1017 99.5127
R18267 vdd.n2636 vdd.n1018 99.5127
R18268 vdd.n1018 vdd.n998 99.5127
R18269 vdd.n3246 vdd.n3245 99.5127
R18270 vdd.n3243 vdd.n3209 99.5127
R18271 vdd.n3239 vdd.n3238 99.5127
R18272 vdd.n3236 vdd.n3212 99.5127
R18273 vdd.n3232 vdd.n3231 99.5127
R18274 vdd.n3229 vdd.n3215 99.5127
R18275 vdd.n3225 vdd.n3224 99.5127
R18276 vdd.n3222 vdd.n3219 99.5127
R18277 vdd.n3363 vdd.n787 99.5127
R18278 vdd.n3361 vdd.n3360 99.5127
R18279 vdd.n3358 vdd.n789 99.5127
R18280 vdd.n3354 vdd.n3353 99.5127
R18281 vdd.n3351 vdd.n792 99.5127
R18282 vdd.n3347 vdd.n3346 99.5127
R18283 vdd.n3344 vdd.n795 99.5127
R18284 vdd.n3340 vdd.n3339 99.5127
R18285 vdd.n3337 vdd.n798 99.5127
R18286 vdd.n2895 vdd.n959 99.5127
R18287 vdd.n3015 vdd.n959 99.5127
R18288 vdd.n3015 vdd.n953 99.5127
R18289 vdd.n3011 vdd.n953 99.5127
R18290 vdd.n3011 vdd.n948 99.5127
R18291 vdd.n3008 vdd.n948 99.5127
R18292 vdd.n3008 vdd.n942 99.5127
R18293 vdd.n3005 vdd.n942 99.5127
R18294 vdd.n3005 vdd.n936 99.5127
R18295 vdd.n2997 vdd.n936 99.5127
R18296 vdd.n2997 vdd.n930 99.5127
R18297 vdd.n2993 vdd.n930 99.5127
R18298 vdd.n2993 vdd.n924 99.5127
R18299 vdd.n2990 vdd.n924 99.5127
R18300 vdd.n2990 vdd.n919 99.5127
R18301 vdd.n2987 vdd.n919 99.5127
R18302 vdd.n2987 vdd.n914 99.5127
R18303 vdd.n2984 vdd.n914 99.5127
R18304 vdd.n2984 vdd.n907 99.5127
R18305 vdd.n2981 vdd.n907 99.5127
R18306 vdd.n2981 vdd.n900 99.5127
R18307 vdd.n2978 vdd.n900 99.5127
R18308 vdd.n2978 vdd.n894 99.5127
R18309 vdd.n2975 vdd.n894 99.5127
R18310 vdd.n2975 vdd.n889 99.5127
R18311 vdd.n2972 vdd.n889 99.5127
R18312 vdd.n2972 vdd.n883 99.5127
R18313 vdd.n2969 vdd.n883 99.5127
R18314 vdd.n2969 vdd.n876 99.5127
R18315 vdd.n2966 vdd.n876 99.5127
R18316 vdd.n2966 vdd.n869 99.5127
R18317 vdd.n2963 vdd.n869 99.5127
R18318 vdd.n2963 vdd.n863 99.5127
R18319 vdd.n2960 vdd.n863 99.5127
R18320 vdd.n2960 vdd.n858 99.5127
R18321 vdd.n2957 vdd.n858 99.5127
R18322 vdd.n2957 vdd.n853 99.5127
R18323 vdd.n2954 vdd.n853 99.5127
R18324 vdd.n2954 vdd.n845 99.5127
R18325 vdd.n2951 vdd.n845 99.5127
R18326 vdd.n2951 vdd.n838 99.5127
R18327 vdd.n838 vdd.n804 99.5127
R18328 vdd.n3332 vdd.n804 99.5127
R18329 vdd.n2830 vdd.n2829 99.5127
R18330 vdd.n2834 vdd.n2833 99.5127
R18331 vdd.n2838 vdd.n2837 99.5127
R18332 vdd.n2842 vdd.n2841 99.5127
R18333 vdd.n2846 vdd.n2845 99.5127
R18334 vdd.n2850 vdd.n2849 99.5127
R18335 vdd.n2854 vdd.n2853 99.5127
R18336 vdd.n2858 vdd.n2857 99.5127
R18337 vdd.n2862 vdd.n2861 99.5127
R18338 vdd.n2866 vdd.n2865 99.5127
R18339 vdd.n2870 vdd.n2869 99.5127
R18340 vdd.n2874 vdd.n2873 99.5127
R18341 vdd.n2878 vdd.n2877 99.5127
R18342 vdd.n2882 vdd.n2881 99.5127
R18343 vdd.n2886 vdd.n2885 99.5127
R18344 vdd.n2890 vdd.n2889 99.5127
R18345 vdd.n2892 vdd.n2818 99.5127
R18346 vdd.n3096 vdd.n956 99.5127
R18347 vdd.n3096 vdd.n954 99.5127
R18348 vdd.n3100 vdd.n954 99.5127
R18349 vdd.n3100 vdd.n945 99.5127
R18350 vdd.n3108 vdd.n945 99.5127
R18351 vdd.n3108 vdd.n943 99.5127
R18352 vdd.n3112 vdd.n943 99.5127
R18353 vdd.n3112 vdd.n934 99.5127
R18354 vdd.n3120 vdd.n934 99.5127
R18355 vdd.n3120 vdd.n932 99.5127
R18356 vdd.n3124 vdd.n932 99.5127
R18357 vdd.n3124 vdd.n922 99.5127
R18358 vdd.n3132 vdd.n922 99.5127
R18359 vdd.n3132 vdd.n920 99.5127
R18360 vdd.n3136 vdd.n920 99.5127
R18361 vdd.n3136 vdd.n911 99.5127
R18362 vdd.n3144 vdd.n911 99.5127
R18363 vdd.n3144 vdd.n909 99.5127
R18364 vdd.n3149 vdd.n909 99.5127
R18365 vdd.n3149 vdd.n898 99.5127
R18366 vdd.n3157 vdd.n898 99.5127
R18367 vdd.n3157 vdd.n895 99.5127
R18368 vdd.n3161 vdd.n895 99.5127
R18369 vdd.n3161 vdd.n886 99.5127
R18370 vdd.n3169 vdd.n886 99.5127
R18371 vdd.n3169 vdd.n884 99.5127
R18372 vdd.n3173 vdd.n884 99.5127
R18373 vdd.n3173 vdd.n873 99.5127
R18374 vdd.n3181 vdd.n873 99.5127
R18375 vdd.n3181 vdd.n871 99.5127
R18376 vdd.n3185 vdd.n871 99.5127
R18377 vdd.n3185 vdd.n861 99.5127
R18378 vdd.n3193 vdd.n861 99.5127
R18379 vdd.n3193 vdd.n859 99.5127
R18380 vdd.n3197 vdd.n859 99.5127
R18381 vdd.n3197 vdd.n850 99.5127
R18382 vdd.n3205 vdd.n850 99.5127
R18383 vdd.n3205 vdd.n847 99.5127
R18384 vdd.n3254 vdd.n847 99.5127
R18385 vdd.n3254 vdd.n848 99.5127
R18386 vdd.n848 vdd.n839 99.5127
R18387 vdd.n3249 vdd.n839 99.5127
R18388 vdd.n3249 vdd.n807 99.5127
R18389 vdd.n2707 vdd.n2706 99.5127
R18390 vdd.n2703 vdd.n2702 99.5127
R18391 vdd.n2699 vdd.n2698 99.5127
R18392 vdd.n2695 vdd.n2694 99.5127
R18393 vdd.n2691 vdd.n2690 99.5127
R18394 vdd.n2687 vdd.n2686 99.5127
R18395 vdd.n2683 vdd.n2682 99.5127
R18396 vdd.n2679 vdd.n2678 99.5127
R18397 vdd.n2675 vdd.n2674 99.5127
R18398 vdd.n2671 vdd.n2670 99.5127
R18399 vdd.n2667 vdd.n2666 99.5127
R18400 vdd.n2663 vdd.n2662 99.5127
R18401 vdd.n2659 vdd.n2658 99.5127
R18402 vdd.n2655 vdd.n2654 99.5127
R18403 vdd.n2651 vdd.n2650 99.5127
R18404 vdd.n2647 vdd.n2646 99.5127
R18405 vdd.n2643 vdd.n980 99.5127
R18406 vdd.n1480 vdd.n1136 99.5127
R18407 vdd.n1477 vdd.n1136 99.5127
R18408 vdd.n1477 vdd.n1130 99.5127
R18409 vdd.n1474 vdd.n1130 99.5127
R18410 vdd.n1474 vdd.n1125 99.5127
R18411 vdd.n1471 vdd.n1125 99.5127
R18412 vdd.n1471 vdd.n1118 99.5127
R18413 vdd.n1468 vdd.n1118 99.5127
R18414 vdd.n1468 vdd.n1111 99.5127
R18415 vdd.n1465 vdd.n1111 99.5127
R18416 vdd.n1465 vdd.n1105 99.5127
R18417 vdd.n1462 vdd.n1105 99.5127
R18418 vdd.n1462 vdd.n1100 99.5127
R18419 vdd.n1459 vdd.n1100 99.5127
R18420 vdd.n1459 vdd.n1095 99.5127
R18421 vdd.n1456 vdd.n1095 99.5127
R18422 vdd.n1456 vdd.n1089 99.5127
R18423 vdd.n1453 vdd.n1089 99.5127
R18424 vdd.n1453 vdd.n1082 99.5127
R18425 vdd.n1450 vdd.n1082 99.5127
R18426 vdd.n1450 vdd.n1075 99.5127
R18427 vdd.n1447 vdd.n1075 99.5127
R18428 vdd.n1447 vdd.n1069 99.5127
R18429 vdd.n1444 vdd.n1069 99.5127
R18430 vdd.n1444 vdd.n1064 99.5127
R18431 vdd.n1441 vdd.n1064 99.5127
R18432 vdd.n1441 vdd.n1058 99.5127
R18433 vdd.n1438 vdd.n1058 99.5127
R18434 vdd.n1438 vdd.n1051 99.5127
R18435 vdd.n1409 vdd.n1051 99.5127
R18436 vdd.n1409 vdd.n1045 99.5127
R18437 vdd.n1412 vdd.n1045 99.5127
R18438 vdd.n1412 vdd.n1040 99.5127
R18439 vdd.n1424 vdd.n1040 99.5127
R18440 vdd.n1424 vdd.n1035 99.5127
R18441 vdd.n1420 vdd.n1035 99.5127
R18442 vdd.n1420 vdd.n1030 99.5127
R18443 vdd.n1417 vdd.n1030 99.5127
R18444 vdd.n1417 vdd.n1023 99.5127
R18445 vdd.n1023 vdd.n1014 99.5127
R18446 vdd.n2638 vdd.n1014 99.5127
R18447 vdd.n2639 vdd.n2638 99.5127
R18448 vdd.n2639 vdd.n1006 99.5127
R18449 vdd.n1284 vdd.n1283 99.5127
R18450 vdd.n1288 vdd.n1287 99.5127
R18451 vdd.n1292 vdd.n1291 99.5127
R18452 vdd.n1296 vdd.n1295 99.5127
R18453 vdd.n1300 vdd.n1299 99.5127
R18454 vdd.n1304 vdd.n1303 99.5127
R18455 vdd.n1308 vdd.n1307 99.5127
R18456 vdd.n1312 vdd.n1311 99.5127
R18457 vdd.n1513 vdd.n1314 99.5127
R18458 vdd.n1511 vdd.n1510 99.5127
R18459 vdd.n1507 vdd.n1506 99.5127
R18460 vdd.n1503 vdd.n1502 99.5127
R18461 vdd.n1499 vdd.n1498 99.5127
R18462 vdd.n1495 vdd.n1494 99.5127
R18463 vdd.n1491 vdd.n1490 99.5127
R18464 vdd.n1487 vdd.n1486 99.5127
R18465 vdd.n1483 vdd.n1175 99.5127
R18466 vdd.n2514 vdd.n1133 99.5127
R18467 vdd.n2514 vdd.n1131 99.5127
R18468 vdd.n2518 vdd.n1131 99.5127
R18469 vdd.n2518 vdd.n1122 99.5127
R18470 vdd.n2526 vdd.n1122 99.5127
R18471 vdd.n2526 vdd.n1120 99.5127
R18472 vdd.n2530 vdd.n1120 99.5127
R18473 vdd.n2530 vdd.n1109 99.5127
R18474 vdd.n2538 vdd.n1109 99.5127
R18475 vdd.n2538 vdd.n1107 99.5127
R18476 vdd.n2542 vdd.n1107 99.5127
R18477 vdd.n2542 vdd.n1098 99.5127
R18478 vdd.n2550 vdd.n1098 99.5127
R18479 vdd.n2550 vdd.n1096 99.5127
R18480 vdd.n2554 vdd.n1096 99.5127
R18481 vdd.n2554 vdd.n1086 99.5127
R18482 vdd.n2562 vdd.n1086 99.5127
R18483 vdd.n2562 vdd.n1084 99.5127
R18484 vdd.n2566 vdd.n1084 99.5127
R18485 vdd.n2566 vdd.n1073 99.5127
R18486 vdd.n2574 vdd.n1073 99.5127
R18487 vdd.n2574 vdd.n1070 99.5127
R18488 vdd.n2579 vdd.n1070 99.5127
R18489 vdd.n2579 vdd.n1061 99.5127
R18490 vdd.n2587 vdd.n1061 99.5127
R18491 vdd.n2587 vdd.n1059 99.5127
R18492 vdd.n2591 vdd.n1059 99.5127
R18493 vdd.n2591 vdd.n1049 99.5127
R18494 vdd.n2599 vdd.n1049 99.5127
R18495 vdd.n2599 vdd.n1047 99.5127
R18496 vdd.n2603 vdd.n1047 99.5127
R18497 vdd.n2603 vdd.n1038 99.5127
R18498 vdd.n2611 vdd.n1038 99.5127
R18499 vdd.n2611 vdd.n1036 99.5127
R18500 vdd.n2615 vdd.n1036 99.5127
R18501 vdd.n2615 vdd.n1027 99.5127
R18502 vdd.n2623 vdd.n1027 99.5127
R18503 vdd.n2623 vdd.n1024 99.5127
R18504 vdd.n2629 vdd.n1024 99.5127
R18505 vdd.n2629 vdd.n1025 99.5127
R18506 vdd.n1025 vdd.n1016 99.5127
R18507 vdd.n1016 vdd.n1007 99.5127
R18508 vdd.n2711 vdd.n1007 99.5127
R18509 vdd.n9 vdd.n7 98.9633
R18510 vdd.n2 vdd.n0 98.9633
R18511 vdd.n9 vdd.n8 98.6055
R18512 vdd.n11 vdd.n10 98.6055
R18513 vdd.n13 vdd.n12 98.6055
R18514 vdd.n6 vdd.n5 98.6055
R18515 vdd.n4 vdd.n3 98.6055
R18516 vdd.n2 vdd.n1 98.6055
R18517 vdd.t124 vdd.n303 85.8723
R18518 vdd.t240 vdd.n244 85.8723
R18519 vdd.t105 vdd.n201 85.8723
R18520 vdd.t229 vdd.n142 85.8723
R18521 vdd.t210 vdd.n100 85.8723
R18522 vdd.t170 vdd.n41 85.8723
R18523 vdd.t151 vdd.n2177 85.8723
R18524 vdd.t193 vdd.n2236 85.8723
R18525 vdd.t131 vdd.n2075 85.8723
R18526 vdd.t176 vdd.n2134 85.8723
R18527 vdd.t171 vdd.n1974 85.8723
R18528 vdd.t212 vdd.n2033 85.8723
R18529 vdd.n897 vdd.n896 78.546
R18530 vdd.n2577 vdd.n1071 78.546
R18531 vdd.n290 vdd.n289 75.1835
R18532 vdd.n288 vdd.n287 75.1835
R18533 vdd.n286 vdd.n285 75.1835
R18534 vdd.n284 vdd.n283 75.1835
R18535 vdd.n282 vdd.n281 75.1835
R18536 vdd.n280 vdd.n279 75.1835
R18537 vdd.n278 vdd.n277 75.1835
R18538 vdd.n276 vdd.n275 75.1835
R18539 vdd.n274 vdd.n273 75.1835
R18540 vdd.n188 vdd.n187 75.1835
R18541 vdd.n186 vdd.n185 75.1835
R18542 vdd.n184 vdd.n183 75.1835
R18543 vdd.n182 vdd.n181 75.1835
R18544 vdd.n180 vdd.n179 75.1835
R18545 vdd.n178 vdd.n177 75.1835
R18546 vdd.n176 vdd.n175 75.1835
R18547 vdd.n174 vdd.n173 75.1835
R18548 vdd.n172 vdd.n171 75.1835
R18549 vdd.n87 vdd.n86 75.1835
R18550 vdd.n85 vdd.n84 75.1835
R18551 vdd.n83 vdd.n82 75.1835
R18552 vdd.n81 vdd.n80 75.1835
R18553 vdd.n79 vdd.n78 75.1835
R18554 vdd.n77 vdd.n76 75.1835
R18555 vdd.n75 vdd.n74 75.1835
R18556 vdd.n73 vdd.n72 75.1835
R18557 vdd.n71 vdd.n70 75.1835
R18558 vdd.n2207 vdd.n2206 75.1835
R18559 vdd.n2209 vdd.n2208 75.1835
R18560 vdd.n2211 vdd.n2210 75.1835
R18561 vdd.n2213 vdd.n2212 75.1835
R18562 vdd.n2215 vdd.n2214 75.1835
R18563 vdd.n2217 vdd.n2216 75.1835
R18564 vdd.n2219 vdd.n2218 75.1835
R18565 vdd.n2221 vdd.n2220 75.1835
R18566 vdd.n2223 vdd.n2222 75.1835
R18567 vdd.n2105 vdd.n2104 75.1835
R18568 vdd.n2107 vdd.n2106 75.1835
R18569 vdd.n2109 vdd.n2108 75.1835
R18570 vdd.n2111 vdd.n2110 75.1835
R18571 vdd.n2113 vdd.n2112 75.1835
R18572 vdd.n2115 vdd.n2114 75.1835
R18573 vdd.n2117 vdd.n2116 75.1835
R18574 vdd.n2119 vdd.n2118 75.1835
R18575 vdd.n2121 vdd.n2120 75.1835
R18576 vdd.n2004 vdd.n2003 75.1835
R18577 vdd.n2006 vdd.n2005 75.1835
R18578 vdd.n2008 vdd.n2007 75.1835
R18579 vdd.n2010 vdd.n2009 75.1835
R18580 vdd.n2012 vdd.n2011 75.1835
R18581 vdd.n2014 vdd.n2013 75.1835
R18582 vdd.n2016 vdd.n2015 75.1835
R18583 vdd.n2018 vdd.n2017 75.1835
R18584 vdd.n2020 vdd.n2019 75.1835
R18585 vdd.n3088 vdd.n2801 72.8958
R18586 vdd.n3088 vdd.n2802 72.8958
R18587 vdd.n3088 vdd.n2803 72.8958
R18588 vdd.n3088 vdd.n2804 72.8958
R18589 vdd.n3088 vdd.n2805 72.8958
R18590 vdd.n3088 vdd.n2806 72.8958
R18591 vdd.n3088 vdd.n2807 72.8958
R18592 vdd.n3088 vdd.n2808 72.8958
R18593 vdd.n3088 vdd.n2809 72.8958
R18594 vdd.n3088 vdd.n2810 72.8958
R18595 vdd.n3088 vdd.n2811 72.8958
R18596 vdd.n3088 vdd.n2812 72.8958
R18597 vdd.n3088 vdd.n2813 72.8958
R18598 vdd.n3088 vdd.n2814 72.8958
R18599 vdd.n3088 vdd.n2815 72.8958
R18600 vdd.n3088 vdd.n2816 72.8958
R18601 vdd.n3088 vdd.n2817 72.8958
R18602 vdd.n803 vdd.n692 72.8958
R18603 vdd.n3338 vdd.n692 72.8958
R18604 vdd.n797 vdd.n692 72.8958
R18605 vdd.n3345 vdd.n692 72.8958
R18606 vdd.n794 vdd.n692 72.8958
R18607 vdd.n3352 vdd.n692 72.8958
R18608 vdd.n791 vdd.n692 72.8958
R18609 vdd.n3359 vdd.n692 72.8958
R18610 vdd.n3362 vdd.n692 72.8958
R18611 vdd.n3218 vdd.n692 72.8958
R18612 vdd.n3223 vdd.n692 72.8958
R18613 vdd.n3217 vdd.n692 72.8958
R18614 vdd.n3230 vdd.n692 72.8958
R18615 vdd.n3214 vdd.n692 72.8958
R18616 vdd.n3237 vdd.n692 72.8958
R18617 vdd.n3211 vdd.n692 72.8958
R18618 vdd.n3244 vdd.n692 72.8958
R18619 vdd.n2507 vdd.n2506 72.8958
R18620 vdd.n2506 vdd.n1142 72.8958
R18621 vdd.n2506 vdd.n1143 72.8958
R18622 vdd.n2506 vdd.n1144 72.8958
R18623 vdd.n2506 vdd.n1145 72.8958
R18624 vdd.n2506 vdd.n1146 72.8958
R18625 vdd.n2506 vdd.n1147 72.8958
R18626 vdd.n2506 vdd.n1148 72.8958
R18627 vdd.n2506 vdd.n1149 72.8958
R18628 vdd.n2506 vdd.n1150 72.8958
R18629 vdd.n2506 vdd.n1151 72.8958
R18630 vdd.n2506 vdd.n1152 72.8958
R18631 vdd.n2506 vdd.n1153 72.8958
R18632 vdd.n2506 vdd.n1154 72.8958
R18633 vdd.n2506 vdd.n1155 72.8958
R18634 vdd.n2506 vdd.n1156 72.8958
R18635 vdd.n2506 vdd.n1157 72.8958
R18636 vdd.n2784 vdd.n981 72.8958
R18637 vdd.n2784 vdd.n982 72.8958
R18638 vdd.n2784 vdd.n983 72.8958
R18639 vdd.n2784 vdd.n984 72.8958
R18640 vdd.n2784 vdd.n985 72.8958
R18641 vdd.n2784 vdd.n986 72.8958
R18642 vdd.n2784 vdd.n987 72.8958
R18643 vdd.n2784 vdd.n988 72.8958
R18644 vdd.n2784 vdd.n989 72.8958
R18645 vdd.n2784 vdd.n990 72.8958
R18646 vdd.n2784 vdd.n991 72.8958
R18647 vdd.n2784 vdd.n992 72.8958
R18648 vdd.n2784 vdd.n993 72.8958
R18649 vdd.n2784 vdd.n994 72.8958
R18650 vdd.n2784 vdd.n995 72.8958
R18651 vdd.n2784 vdd.n996 72.8958
R18652 vdd.n2784 vdd.n997 72.8958
R18653 vdd.n3089 vdd.n3088 72.8958
R18654 vdd.n3088 vdd.n2785 72.8958
R18655 vdd.n3088 vdd.n2786 72.8958
R18656 vdd.n3088 vdd.n2787 72.8958
R18657 vdd.n3088 vdd.n2788 72.8958
R18658 vdd.n3088 vdd.n2789 72.8958
R18659 vdd.n3088 vdd.n2790 72.8958
R18660 vdd.n3088 vdd.n2791 72.8958
R18661 vdd.n3088 vdd.n2792 72.8958
R18662 vdd.n3088 vdd.n2793 72.8958
R18663 vdd.n3088 vdd.n2794 72.8958
R18664 vdd.n3088 vdd.n2795 72.8958
R18665 vdd.n3088 vdd.n2796 72.8958
R18666 vdd.n3088 vdd.n2797 72.8958
R18667 vdd.n3088 vdd.n2798 72.8958
R18668 vdd.n3088 vdd.n2799 72.8958
R18669 vdd.n3088 vdd.n2800 72.8958
R18670 vdd.n3268 vdd.n692 72.8958
R18671 vdd.n835 vdd.n692 72.8958
R18672 vdd.n3276 vdd.n692 72.8958
R18673 vdd.n830 vdd.n692 72.8958
R18674 vdd.n3283 vdd.n692 72.8958
R18675 vdd.n827 vdd.n692 72.8958
R18676 vdd.n3290 vdd.n692 72.8958
R18677 vdd.n824 vdd.n692 72.8958
R18678 vdd.n3297 vdd.n692 72.8958
R18679 vdd.n3301 vdd.n692 72.8958
R18680 vdd.n821 vdd.n692 72.8958
R18681 vdd.n3308 vdd.n692 72.8958
R18682 vdd.n818 vdd.n692 72.8958
R18683 vdd.n3315 vdd.n692 72.8958
R18684 vdd.n815 vdd.n692 72.8958
R18685 vdd.n3322 vdd.n692 72.8958
R18686 vdd.n3325 vdd.n692 72.8958
R18687 vdd.n2784 vdd.n979 72.8958
R18688 vdd.n2784 vdd.n978 72.8958
R18689 vdd.n2784 vdd.n977 72.8958
R18690 vdd.n2784 vdd.n976 72.8958
R18691 vdd.n2784 vdd.n975 72.8958
R18692 vdd.n2784 vdd.n974 72.8958
R18693 vdd.n2784 vdd.n973 72.8958
R18694 vdd.n2784 vdd.n972 72.8958
R18695 vdd.n2784 vdd.n971 72.8958
R18696 vdd.n2784 vdd.n970 72.8958
R18697 vdd.n2784 vdd.n969 72.8958
R18698 vdd.n2784 vdd.n968 72.8958
R18699 vdd.n2784 vdd.n967 72.8958
R18700 vdd.n2784 vdd.n966 72.8958
R18701 vdd.n2784 vdd.n965 72.8958
R18702 vdd.n2784 vdd.n964 72.8958
R18703 vdd.n2784 vdd.n963 72.8958
R18704 vdd.n2506 vdd.n1158 72.8958
R18705 vdd.n2506 vdd.n1159 72.8958
R18706 vdd.n2506 vdd.n1160 72.8958
R18707 vdd.n2506 vdd.n1161 72.8958
R18708 vdd.n2506 vdd.n1162 72.8958
R18709 vdd.n2506 vdd.n1163 72.8958
R18710 vdd.n2506 vdd.n1164 72.8958
R18711 vdd.n2506 vdd.n1165 72.8958
R18712 vdd.n2506 vdd.n1166 72.8958
R18713 vdd.n2506 vdd.n1167 72.8958
R18714 vdd.n2506 vdd.n1168 72.8958
R18715 vdd.n2506 vdd.n1169 72.8958
R18716 vdd.n2506 vdd.n1170 72.8958
R18717 vdd.n2506 vdd.n1171 72.8958
R18718 vdd.n2506 vdd.n1172 72.8958
R18719 vdd.n2506 vdd.n1173 72.8958
R18720 vdd.n2506 vdd.n1174 72.8958
R18721 vdd.n1874 vdd.n1873 66.2847
R18722 vdd.n1873 vdd.n1649 66.2847
R18723 vdd.n1873 vdd.n1650 66.2847
R18724 vdd.n1873 vdd.n1651 66.2847
R18725 vdd.n1873 vdd.n1652 66.2847
R18726 vdd.n1873 vdd.n1653 66.2847
R18727 vdd.n1873 vdd.n1654 66.2847
R18728 vdd.n1873 vdd.n1655 66.2847
R18729 vdd.n1873 vdd.n1656 66.2847
R18730 vdd.n1873 vdd.n1657 66.2847
R18731 vdd.n1873 vdd.n1658 66.2847
R18732 vdd.n1873 vdd.n1659 66.2847
R18733 vdd.n1873 vdd.n1660 66.2847
R18734 vdd.n1873 vdd.n1661 66.2847
R18735 vdd.n1873 vdd.n1662 66.2847
R18736 vdd.n1873 vdd.n1663 66.2847
R18737 vdd.n1873 vdd.n1664 66.2847
R18738 vdd.n1873 vdd.n1665 66.2847
R18739 vdd.n1873 vdd.n1666 66.2847
R18740 vdd.n1873 vdd.n1667 66.2847
R18741 vdd.n1873 vdd.n1668 66.2847
R18742 vdd.n1873 vdd.n1669 66.2847
R18743 vdd.n1873 vdd.n1670 66.2847
R18744 vdd.n1873 vdd.n1671 66.2847
R18745 vdd.n1873 vdd.n1672 66.2847
R18746 vdd.n1873 vdd.n1673 66.2847
R18747 vdd.n1873 vdd.n1674 66.2847
R18748 vdd.n1873 vdd.n1675 66.2847
R18749 vdd.n1873 vdd.n1676 66.2847
R18750 vdd.n1873 vdd.n1677 66.2847
R18751 vdd.n1873 vdd.n1678 66.2847
R18752 vdd.n1526 vdd.n1141 66.2847
R18753 vdd.n1523 vdd.n1141 66.2847
R18754 vdd.n1519 vdd.n1141 66.2847
R18755 vdd.n2372 vdd.n1141 66.2847
R18756 vdd.n1275 vdd.n1141 66.2847
R18757 vdd.n2379 vdd.n1141 66.2847
R18758 vdd.n1268 vdd.n1141 66.2847
R18759 vdd.n2386 vdd.n1141 66.2847
R18760 vdd.n1261 vdd.n1141 66.2847
R18761 vdd.n2393 vdd.n1141 66.2847
R18762 vdd.n1255 vdd.n1141 66.2847
R18763 vdd.n1250 vdd.n1141 66.2847
R18764 vdd.n2404 vdd.n1141 66.2847
R18765 vdd.n1242 vdd.n1141 66.2847
R18766 vdd.n2411 vdd.n1141 66.2847
R18767 vdd.n1235 vdd.n1141 66.2847
R18768 vdd.n2418 vdd.n1141 66.2847
R18769 vdd.n1228 vdd.n1141 66.2847
R18770 vdd.n2425 vdd.n1141 66.2847
R18771 vdd.n1221 vdd.n1141 66.2847
R18772 vdd.n2432 vdd.n1141 66.2847
R18773 vdd.n1215 vdd.n1141 66.2847
R18774 vdd.n1210 vdd.n1141 66.2847
R18775 vdd.n2443 vdd.n1141 66.2847
R18776 vdd.n1202 vdd.n1141 66.2847
R18777 vdd.n2450 vdd.n1141 66.2847
R18778 vdd.n1195 vdd.n1141 66.2847
R18779 vdd.n2457 vdd.n1141 66.2847
R18780 vdd.n1188 vdd.n1141 66.2847
R18781 vdd.n2464 vdd.n1141 66.2847
R18782 vdd.n2469 vdd.n1141 66.2847
R18783 vdd.n1184 vdd.n1141 66.2847
R18784 vdd.n3495 vdd.n3494 66.2847
R18785 vdd.n3495 vdd.n693 66.2847
R18786 vdd.n3495 vdd.n694 66.2847
R18787 vdd.n3495 vdd.n695 66.2847
R18788 vdd.n3495 vdd.n696 66.2847
R18789 vdd.n3495 vdd.n697 66.2847
R18790 vdd.n3495 vdd.n698 66.2847
R18791 vdd.n3495 vdd.n699 66.2847
R18792 vdd.n3495 vdd.n700 66.2847
R18793 vdd.n3495 vdd.n701 66.2847
R18794 vdd.n3495 vdd.n702 66.2847
R18795 vdd.n3495 vdd.n703 66.2847
R18796 vdd.n3495 vdd.n704 66.2847
R18797 vdd.n3495 vdd.n705 66.2847
R18798 vdd.n3495 vdd.n706 66.2847
R18799 vdd.n3495 vdd.n707 66.2847
R18800 vdd.n3495 vdd.n708 66.2847
R18801 vdd.n3495 vdd.n709 66.2847
R18802 vdd.n3495 vdd.n710 66.2847
R18803 vdd.n3495 vdd.n711 66.2847
R18804 vdd.n3495 vdd.n712 66.2847
R18805 vdd.n3495 vdd.n713 66.2847
R18806 vdd.n3495 vdd.n714 66.2847
R18807 vdd.n3495 vdd.n715 66.2847
R18808 vdd.n3495 vdd.n716 66.2847
R18809 vdd.n3495 vdd.n717 66.2847
R18810 vdd.n3495 vdd.n718 66.2847
R18811 vdd.n3495 vdd.n719 66.2847
R18812 vdd.n3495 vdd.n720 66.2847
R18813 vdd.n3495 vdd.n721 66.2847
R18814 vdd.n3495 vdd.n722 66.2847
R18815 vdd.n3626 vdd.n3625 66.2847
R18816 vdd.n3626 vdd.n424 66.2847
R18817 vdd.n3626 vdd.n423 66.2847
R18818 vdd.n3626 vdd.n422 66.2847
R18819 vdd.n3626 vdd.n421 66.2847
R18820 vdd.n3626 vdd.n420 66.2847
R18821 vdd.n3626 vdd.n419 66.2847
R18822 vdd.n3626 vdd.n418 66.2847
R18823 vdd.n3626 vdd.n417 66.2847
R18824 vdd.n3626 vdd.n416 66.2847
R18825 vdd.n3626 vdd.n415 66.2847
R18826 vdd.n3626 vdd.n414 66.2847
R18827 vdd.n3626 vdd.n413 66.2847
R18828 vdd.n3626 vdd.n412 66.2847
R18829 vdd.n3626 vdd.n411 66.2847
R18830 vdd.n3626 vdd.n410 66.2847
R18831 vdd.n3626 vdd.n409 66.2847
R18832 vdd.n3626 vdd.n408 66.2847
R18833 vdd.n3626 vdd.n407 66.2847
R18834 vdd.n3626 vdd.n406 66.2847
R18835 vdd.n3626 vdd.n405 66.2847
R18836 vdd.n3626 vdd.n404 66.2847
R18837 vdd.n3626 vdd.n403 66.2847
R18838 vdd.n3626 vdd.n402 66.2847
R18839 vdd.n3626 vdd.n401 66.2847
R18840 vdd.n3626 vdd.n400 66.2847
R18841 vdd.n3626 vdd.n399 66.2847
R18842 vdd.n3626 vdd.n398 66.2847
R18843 vdd.n3626 vdd.n397 66.2847
R18844 vdd.n3626 vdd.n396 66.2847
R18845 vdd.n3626 vdd.n395 66.2847
R18846 vdd.n3626 vdd.n394 66.2847
R18847 vdd.n467 vdd.n394 52.4337
R18848 vdd.n473 vdd.n395 52.4337
R18849 vdd.n477 vdd.n396 52.4337
R18850 vdd.n483 vdd.n397 52.4337
R18851 vdd.n487 vdd.n398 52.4337
R18852 vdd.n493 vdd.n399 52.4337
R18853 vdd.n497 vdd.n400 52.4337
R18854 vdd.n503 vdd.n401 52.4337
R18855 vdd.n507 vdd.n402 52.4337
R18856 vdd.n513 vdd.n403 52.4337
R18857 vdd.n517 vdd.n404 52.4337
R18858 vdd.n523 vdd.n405 52.4337
R18859 vdd.n527 vdd.n406 52.4337
R18860 vdd.n533 vdd.n407 52.4337
R18861 vdd.n537 vdd.n408 52.4337
R18862 vdd.n543 vdd.n409 52.4337
R18863 vdd.n547 vdd.n410 52.4337
R18864 vdd.n553 vdd.n411 52.4337
R18865 vdd.n557 vdd.n412 52.4337
R18866 vdd.n563 vdd.n413 52.4337
R18867 vdd.n567 vdd.n414 52.4337
R18868 vdd.n573 vdd.n415 52.4337
R18869 vdd.n577 vdd.n416 52.4337
R18870 vdd.n583 vdd.n417 52.4337
R18871 vdd.n587 vdd.n418 52.4337
R18872 vdd.n593 vdd.n419 52.4337
R18873 vdd.n597 vdd.n420 52.4337
R18874 vdd.n603 vdd.n421 52.4337
R18875 vdd.n607 vdd.n422 52.4337
R18876 vdd.n613 vdd.n423 52.4337
R18877 vdd.n616 vdd.n424 52.4337
R18878 vdd.n3625 vdd.n3624 52.4337
R18879 vdd.n3494 vdd.n3493 52.4337
R18880 vdd.n728 vdd.n693 52.4337
R18881 vdd.n734 vdd.n694 52.4337
R18882 vdd.n3483 vdd.n695 52.4337
R18883 vdd.n3479 vdd.n696 52.4337
R18884 vdd.n3475 vdd.n697 52.4337
R18885 vdd.n3471 vdd.n698 52.4337
R18886 vdd.n3467 vdd.n699 52.4337
R18887 vdd.n3463 vdd.n700 52.4337
R18888 vdd.n3459 vdd.n701 52.4337
R18889 vdd.n3451 vdd.n702 52.4337
R18890 vdd.n3447 vdd.n703 52.4337
R18891 vdd.n3443 vdd.n704 52.4337
R18892 vdd.n3439 vdd.n705 52.4337
R18893 vdd.n3435 vdd.n706 52.4337
R18894 vdd.n3431 vdd.n707 52.4337
R18895 vdd.n3427 vdd.n708 52.4337
R18896 vdd.n3423 vdd.n709 52.4337
R18897 vdd.n3419 vdd.n710 52.4337
R18898 vdd.n3415 vdd.n711 52.4337
R18899 vdd.n3411 vdd.n712 52.4337
R18900 vdd.n3405 vdd.n713 52.4337
R18901 vdd.n3401 vdd.n714 52.4337
R18902 vdd.n3397 vdd.n715 52.4337
R18903 vdd.n3393 vdd.n716 52.4337
R18904 vdd.n3389 vdd.n717 52.4337
R18905 vdd.n3385 vdd.n718 52.4337
R18906 vdd.n3381 vdd.n719 52.4337
R18907 vdd.n3377 vdd.n720 52.4337
R18908 vdd.n3373 vdd.n721 52.4337
R18909 vdd.n3369 vdd.n722 52.4337
R18910 vdd.n2471 vdd.n1184 52.4337
R18911 vdd.n2469 vdd.n2468 52.4337
R18912 vdd.n2464 vdd.n2463 52.4337
R18913 vdd.n2459 vdd.n1188 52.4337
R18914 vdd.n2457 vdd.n2456 52.4337
R18915 vdd.n2452 vdd.n1195 52.4337
R18916 vdd.n2450 vdd.n2449 52.4337
R18917 vdd.n2445 vdd.n1202 52.4337
R18918 vdd.n2443 vdd.n2442 52.4337
R18919 vdd.n1211 vdd.n1210 52.4337
R18920 vdd.n2434 vdd.n1215 52.4337
R18921 vdd.n2432 vdd.n2431 52.4337
R18922 vdd.n2427 vdd.n1221 52.4337
R18923 vdd.n2425 vdd.n2424 52.4337
R18924 vdd.n2420 vdd.n1228 52.4337
R18925 vdd.n2418 vdd.n2417 52.4337
R18926 vdd.n2413 vdd.n1235 52.4337
R18927 vdd.n2411 vdd.n2410 52.4337
R18928 vdd.n2406 vdd.n1242 52.4337
R18929 vdd.n2404 vdd.n2403 52.4337
R18930 vdd.n1251 vdd.n1250 52.4337
R18931 vdd.n2395 vdd.n1255 52.4337
R18932 vdd.n2393 vdd.n2392 52.4337
R18933 vdd.n2388 vdd.n1261 52.4337
R18934 vdd.n2386 vdd.n2385 52.4337
R18935 vdd.n2381 vdd.n1268 52.4337
R18936 vdd.n2379 vdd.n2378 52.4337
R18937 vdd.n2374 vdd.n1275 52.4337
R18938 vdd.n2372 vdd.n2371 52.4337
R18939 vdd.n1520 vdd.n1519 52.4337
R18940 vdd.n1524 vdd.n1523 52.4337
R18941 vdd.n2360 vdd.n1526 52.4337
R18942 vdd.n1875 vdd.n1874 52.4337
R18943 vdd.n1681 vdd.n1649 52.4337
R18944 vdd.n1685 vdd.n1650 52.4337
R18945 vdd.n1687 vdd.n1651 52.4337
R18946 vdd.n1691 vdd.n1652 52.4337
R18947 vdd.n1693 vdd.n1653 52.4337
R18948 vdd.n1697 vdd.n1654 52.4337
R18949 vdd.n1699 vdd.n1655 52.4337
R18950 vdd.n1703 vdd.n1656 52.4337
R18951 vdd.n1705 vdd.n1657 52.4337
R18952 vdd.n1711 vdd.n1658 52.4337
R18953 vdd.n1713 vdd.n1659 52.4337
R18954 vdd.n1717 vdd.n1660 52.4337
R18955 vdd.n1719 vdd.n1661 52.4337
R18956 vdd.n1723 vdd.n1662 52.4337
R18957 vdd.n1725 vdd.n1663 52.4337
R18958 vdd.n1729 vdd.n1664 52.4337
R18959 vdd.n1731 vdd.n1665 52.4337
R18960 vdd.n1735 vdd.n1666 52.4337
R18961 vdd.n1737 vdd.n1667 52.4337
R18962 vdd.n1809 vdd.n1668 52.4337
R18963 vdd.n1742 vdd.n1669 52.4337
R18964 vdd.n1746 vdd.n1670 52.4337
R18965 vdd.n1748 vdd.n1671 52.4337
R18966 vdd.n1752 vdd.n1672 52.4337
R18967 vdd.n1754 vdd.n1673 52.4337
R18968 vdd.n1758 vdd.n1674 52.4337
R18969 vdd.n1760 vdd.n1675 52.4337
R18970 vdd.n1764 vdd.n1676 52.4337
R18971 vdd.n1766 vdd.n1677 52.4337
R18972 vdd.n1770 vdd.n1678 52.4337
R18973 vdd.n1874 vdd.n1648 52.4337
R18974 vdd.n1684 vdd.n1649 52.4337
R18975 vdd.n1686 vdd.n1650 52.4337
R18976 vdd.n1690 vdd.n1651 52.4337
R18977 vdd.n1692 vdd.n1652 52.4337
R18978 vdd.n1696 vdd.n1653 52.4337
R18979 vdd.n1698 vdd.n1654 52.4337
R18980 vdd.n1702 vdd.n1655 52.4337
R18981 vdd.n1704 vdd.n1656 52.4337
R18982 vdd.n1710 vdd.n1657 52.4337
R18983 vdd.n1712 vdd.n1658 52.4337
R18984 vdd.n1716 vdd.n1659 52.4337
R18985 vdd.n1718 vdd.n1660 52.4337
R18986 vdd.n1722 vdd.n1661 52.4337
R18987 vdd.n1724 vdd.n1662 52.4337
R18988 vdd.n1728 vdd.n1663 52.4337
R18989 vdd.n1730 vdd.n1664 52.4337
R18990 vdd.n1734 vdd.n1665 52.4337
R18991 vdd.n1736 vdd.n1666 52.4337
R18992 vdd.n1740 vdd.n1667 52.4337
R18993 vdd.n1741 vdd.n1668 52.4337
R18994 vdd.n1745 vdd.n1669 52.4337
R18995 vdd.n1747 vdd.n1670 52.4337
R18996 vdd.n1751 vdd.n1671 52.4337
R18997 vdd.n1753 vdd.n1672 52.4337
R18998 vdd.n1757 vdd.n1673 52.4337
R18999 vdd.n1759 vdd.n1674 52.4337
R19000 vdd.n1763 vdd.n1675 52.4337
R19001 vdd.n1765 vdd.n1676 52.4337
R19002 vdd.n1769 vdd.n1677 52.4337
R19003 vdd.n1771 vdd.n1678 52.4337
R19004 vdd.n1526 vdd.n1525 52.4337
R19005 vdd.n1523 vdd.n1522 52.4337
R19006 vdd.n1519 vdd.n1276 52.4337
R19007 vdd.n2373 vdd.n2372 52.4337
R19008 vdd.n1275 vdd.n1269 52.4337
R19009 vdd.n2380 vdd.n2379 52.4337
R19010 vdd.n1268 vdd.n1262 52.4337
R19011 vdd.n2387 vdd.n2386 52.4337
R19012 vdd.n1261 vdd.n1256 52.4337
R19013 vdd.n2394 vdd.n2393 52.4337
R19014 vdd.n1255 vdd.n1254 52.4337
R19015 vdd.n1250 vdd.n1243 52.4337
R19016 vdd.n2405 vdd.n2404 52.4337
R19017 vdd.n1242 vdd.n1236 52.4337
R19018 vdd.n2412 vdd.n2411 52.4337
R19019 vdd.n1235 vdd.n1229 52.4337
R19020 vdd.n2419 vdd.n2418 52.4337
R19021 vdd.n1228 vdd.n1222 52.4337
R19022 vdd.n2426 vdd.n2425 52.4337
R19023 vdd.n1221 vdd.n1216 52.4337
R19024 vdd.n2433 vdd.n2432 52.4337
R19025 vdd.n1215 vdd.n1214 52.4337
R19026 vdd.n1210 vdd.n1203 52.4337
R19027 vdd.n2444 vdd.n2443 52.4337
R19028 vdd.n1202 vdd.n1196 52.4337
R19029 vdd.n2451 vdd.n2450 52.4337
R19030 vdd.n1195 vdd.n1189 52.4337
R19031 vdd.n2458 vdd.n2457 52.4337
R19032 vdd.n1188 vdd.n1185 52.4337
R19033 vdd.n2465 vdd.n2464 52.4337
R19034 vdd.n2470 vdd.n2469 52.4337
R19035 vdd.n1530 vdd.n1184 52.4337
R19036 vdd.n3494 vdd.n725 52.4337
R19037 vdd.n733 vdd.n693 52.4337
R19038 vdd.n3484 vdd.n694 52.4337
R19039 vdd.n3480 vdd.n695 52.4337
R19040 vdd.n3476 vdd.n696 52.4337
R19041 vdd.n3472 vdd.n697 52.4337
R19042 vdd.n3468 vdd.n698 52.4337
R19043 vdd.n3464 vdd.n699 52.4337
R19044 vdd.n3460 vdd.n700 52.4337
R19045 vdd.n3450 vdd.n701 52.4337
R19046 vdd.n3448 vdd.n702 52.4337
R19047 vdd.n3444 vdd.n703 52.4337
R19048 vdd.n3440 vdd.n704 52.4337
R19049 vdd.n3436 vdd.n705 52.4337
R19050 vdd.n3432 vdd.n706 52.4337
R19051 vdd.n3428 vdd.n707 52.4337
R19052 vdd.n3424 vdd.n708 52.4337
R19053 vdd.n3420 vdd.n709 52.4337
R19054 vdd.n3416 vdd.n710 52.4337
R19055 vdd.n3412 vdd.n711 52.4337
R19056 vdd.n3404 vdd.n712 52.4337
R19057 vdd.n3402 vdd.n713 52.4337
R19058 vdd.n3398 vdd.n714 52.4337
R19059 vdd.n3394 vdd.n715 52.4337
R19060 vdd.n3390 vdd.n716 52.4337
R19061 vdd.n3386 vdd.n717 52.4337
R19062 vdd.n3382 vdd.n718 52.4337
R19063 vdd.n3378 vdd.n719 52.4337
R19064 vdd.n3374 vdd.n720 52.4337
R19065 vdd.n3370 vdd.n721 52.4337
R19066 vdd.n722 vdd.n691 52.4337
R19067 vdd.n3625 vdd.n425 52.4337
R19068 vdd.n614 vdd.n424 52.4337
R19069 vdd.n608 vdd.n423 52.4337
R19070 vdd.n604 vdd.n422 52.4337
R19071 vdd.n598 vdd.n421 52.4337
R19072 vdd.n594 vdd.n420 52.4337
R19073 vdd.n588 vdd.n419 52.4337
R19074 vdd.n584 vdd.n418 52.4337
R19075 vdd.n578 vdd.n417 52.4337
R19076 vdd.n574 vdd.n416 52.4337
R19077 vdd.n568 vdd.n415 52.4337
R19078 vdd.n564 vdd.n414 52.4337
R19079 vdd.n558 vdd.n413 52.4337
R19080 vdd.n554 vdd.n412 52.4337
R19081 vdd.n548 vdd.n411 52.4337
R19082 vdd.n544 vdd.n410 52.4337
R19083 vdd.n538 vdd.n409 52.4337
R19084 vdd.n534 vdd.n408 52.4337
R19085 vdd.n528 vdd.n407 52.4337
R19086 vdd.n524 vdd.n406 52.4337
R19087 vdd.n518 vdd.n405 52.4337
R19088 vdd.n514 vdd.n404 52.4337
R19089 vdd.n508 vdd.n403 52.4337
R19090 vdd.n504 vdd.n402 52.4337
R19091 vdd.n498 vdd.n401 52.4337
R19092 vdd.n494 vdd.n400 52.4337
R19093 vdd.n488 vdd.n399 52.4337
R19094 vdd.n484 vdd.n398 52.4337
R19095 vdd.n478 vdd.n397 52.4337
R19096 vdd.n474 vdd.n396 52.4337
R19097 vdd.n468 vdd.n395 52.4337
R19098 vdd.n394 vdd.n392 52.4337
R19099 vdd.t263 vdd.t278 51.4683
R19100 vdd.n274 vdd.n272 42.0461
R19101 vdd.n172 vdd.n170 42.0461
R19102 vdd.n71 vdd.n69 42.0461
R19103 vdd.n2207 vdd.n2205 42.0461
R19104 vdd.n2105 vdd.n2103 42.0461
R19105 vdd.n2004 vdd.n2002 42.0461
R19106 vdd.n332 vdd.n331 41.6884
R19107 vdd.n230 vdd.n229 41.6884
R19108 vdd.n129 vdd.n128 41.6884
R19109 vdd.n2265 vdd.n2264 41.6884
R19110 vdd.n2163 vdd.n2162 41.6884
R19111 vdd.n2062 vdd.n2061 41.6884
R19112 vdd.n1774 vdd.n1773 41.1157
R19113 vdd.n1812 vdd.n1811 41.1157
R19114 vdd.n1708 vdd.n1707 41.1157
R19115 vdd.n428 vdd.n427 41.1157
R19116 vdd.n566 vdd.n441 41.1157
R19117 vdd.n454 vdd.n453 41.1157
R19118 vdd.n3325 vdd.n3324 39.2114
R19119 vdd.n3322 vdd.n3321 39.2114
R19120 vdd.n3317 vdd.n815 39.2114
R19121 vdd.n3315 vdd.n3314 39.2114
R19122 vdd.n3310 vdd.n818 39.2114
R19123 vdd.n3308 vdd.n3307 39.2114
R19124 vdd.n3303 vdd.n821 39.2114
R19125 vdd.n3301 vdd.n3300 39.2114
R19126 vdd.n3297 vdd.n3296 39.2114
R19127 vdd.n3292 vdd.n824 39.2114
R19128 vdd.n3290 vdd.n3289 39.2114
R19129 vdd.n3285 vdd.n827 39.2114
R19130 vdd.n3283 vdd.n3282 39.2114
R19131 vdd.n3278 vdd.n830 39.2114
R19132 vdd.n3276 vdd.n3275 39.2114
R19133 vdd.n3270 vdd.n835 39.2114
R19134 vdd.n3268 vdd.n3267 39.2114
R19135 vdd.n3090 vdd.n3089 39.2114
R19136 vdd.n2819 vdd.n2785 39.2114
R19137 vdd.n3082 vdd.n2786 39.2114
R19138 vdd.n3078 vdd.n2787 39.2114
R19139 vdd.n3074 vdd.n2788 39.2114
R19140 vdd.n3070 vdd.n2789 39.2114
R19141 vdd.n3066 vdd.n2790 39.2114
R19142 vdd.n3062 vdd.n2791 39.2114
R19143 vdd.n3058 vdd.n2792 39.2114
R19144 vdd.n3054 vdd.n2793 39.2114
R19145 vdd.n3050 vdd.n2794 39.2114
R19146 vdd.n3046 vdd.n2795 39.2114
R19147 vdd.n3042 vdd.n2796 39.2114
R19148 vdd.n3038 vdd.n2797 39.2114
R19149 vdd.n3034 vdd.n2798 39.2114
R19150 vdd.n3030 vdd.n2799 39.2114
R19151 vdd.n3025 vdd.n2800 39.2114
R19152 vdd.n2779 vdd.n997 39.2114
R19153 vdd.n2775 vdd.n996 39.2114
R19154 vdd.n2771 vdd.n995 39.2114
R19155 vdd.n2767 vdd.n994 39.2114
R19156 vdd.n2763 vdd.n993 39.2114
R19157 vdd.n2759 vdd.n992 39.2114
R19158 vdd.n2755 vdd.n991 39.2114
R19159 vdd.n2751 vdd.n990 39.2114
R19160 vdd.n2747 vdd.n989 39.2114
R19161 vdd.n2743 vdd.n988 39.2114
R19162 vdd.n2739 vdd.n987 39.2114
R19163 vdd.n2735 vdd.n986 39.2114
R19164 vdd.n2731 vdd.n985 39.2114
R19165 vdd.n2727 vdd.n984 39.2114
R19166 vdd.n2723 vdd.n983 39.2114
R19167 vdd.n2718 vdd.n982 39.2114
R19168 vdd.n2714 vdd.n981 39.2114
R19169 vdd.n2508 vdd.n2507 39.2114
R19170 vdd.n1176 vdd.n1142 39.2114
R19171 vdd.n2500 vdd.n1143 39.2114
R19172 vdd.n2496 vdd.n1144 39.2114
R19173 vdd.n2492 vdd.n1145 39.2114
R19174 vdd.n2488 vdd.n1146 39.2114
R19175 vdd.n2484 vdd.n1147 39.2114
R19176 vdd.n2480 vdd.n1148 39.2114
R19177 vdd.n2476 vdd.n1149 39.2114
R19178 vdd.n1322 vdd.n1150 39.2114
R19179 vdd.n1326 vdd.n1151 39.2114
R19180 vdd.n1330 vdd.n1152 39.2114
R19181 vdd.n1334 vdd.n1153 39.2114
R19182 vdd.n1338 vdd.n1154 39.2114
R19183 vdd.n1342 vdd.n1155 39.2114
R19184 vdd.n1346 vdd.n1156 39.2114
R19185 vdd.n1351 vdd.n1157 39.2114
R19186 vdd.n3244 vdd.n3243 39.2114
R19187 vdd.n3239 vdd.n3211 39.2114
R19188 vdd.n3237 vdd.n3236 39.2114
R19189 vdd.n3232 vdd.n3214 39.2114
R19190 vdd.n3230 vdd.n3229 39.2114
R19191 vdd.n3225 vdd.n3217 39.2114
R19192 vdd.n3223 vdd.n3222 39.2114
R19193 vdd.n3218 vdd.n787 39.2114
R19194 vdd.n3362 vdd.n3361 39.2114
R19195 vdd.n3359 vdd.n3358 39.2114
R19196 vdd.n3354 vdd.n791 39.2114
R19197 vdd.n3352 vdd.n3351 39.2114
R19198 vdd.n3347 vdd.n794 39.2114
R19199 vdd.n3345 vdd.n3344 39.2114
R19200 vdd.n3340 vdd.n797 39.2114
R19201 vdd.n3338 vdd.n3337 39.2114
R19202 vdd.n3333 vdd.n803 39.2114
R19203 vdd.n2826 vdd.n2801 39.2114
R19204 vdd.n2830 vdd.n2802 39.2114
R19205 vdd.n2834 vdd.n2803 39.2114
R19206 vdd.n2838 vdd.n2804 39.2114
R19207 vdd.n2842 vdd.n2805 39.2114
R19208 vdd.n2846 vdd.n2806 39.2114
R19209 vdd.n2850 vdd.n2807 39.2114
R19210 vdd.n2854 vdd.n2808 39.2114
R19211 vdd.n2858 vdd.n2809 39.2114
R19212 vdd.n2862 vdd.n2810 39.2114
R19213 vdd.n2866 vdd.n2811 39.2114
R19214 vdd.n2870 vdd.n2812 39.2114
R19215 vdd.n2874 vdd.n2813 39.2114
R19216 vdd.n2878 vdd.n2814 39.2114
R19217 vdd.n2882 vdd.n2815 39.2114
R19218 vdd.n2886 vdd.n2816 39.2114
R19219 vdd.n2890 vdd.n2817 39.2114
R19220 vdd.n2829 vdd.n2801 39.2114
R19221 vdd.n2833 vdd.n2802 39.2114
R19222 vdd.n2837 vdd.n2803 39.2114
R19223 vdd.n2841 vdd.n2804 39.2114
R19224 vdd.n2845 vdd.n2805 39.2114
R19225 vdd.n2849 vdd.n2806 39.2114
R19226 vdd.n2853 vdd.n2807 39.2114
R19227 vdd.n2857 vdd.n2808 39.2114
R19228 vdd.n2861 vdd.n2809 39.2114
R19229 vdd.n2865 vdd.n2810 39.2114
R19230 vdd.n2869 vdd.n2811 39.2114
R19231 vdd.n2873 vdd.n2812 39.2114
R19232 vdd.n2877 vdd.n2813 39.2114
R19233 vdd.n2881 vdd.n2814 39.2114
R19234 vdd.n2885 vdd.n2815 39.2114
R19235 vdd.n2889 vdd.n2816 39.2114
R19236 vdd.n2892 vdd.n2817 39.2114
R19237 vdd.n803 vdd.n798 39.2114
R19238 vdd.n3339 vdd.n3338 39.2114
R19239 vdd.n797 vdd.n795 39.2114
R19240 vdd.n3346 vdd.n3345 39.2114
R19241 vdd.n794 vdd.n792 39.2114
R19242 vdd.n3353 vdd.n3352 39.2114
R19243 vdd.n791 vdd.n789 39.2114
R19244 vdd.n3360 vdd.n3359 39.2114
R19245 vdd.n3363 vdd.n3362 39.2114
R19246 vdd.n3219 vdd.n3218 39.2114
R19247 vdd.n3224 vdd.n3223 39.2114
R19248 vdd.n3217 vdd.n3215 39.2114
R19249 vdd.n3231 vdd.n3230 39.2114
R19250 vdd.n3214 vdd.n3212 39.2114
R19251 vdd.n3238 vdd.n3237 39.2114
R19252 vdd.n3211 vdd.n3209 39.2114
R19253 vdd.n3245 vdd.n3244 39.2114
R19254 vdd.n2507 vdd.n1140 39.2114
R19255 vdd.n2501 vdd.n1142 39.2114
R19256 vdd.n2497 vdd.n1143 39.2114
R19257 vdd.n2493 vdd.n1144 39.2114
R19258 vdd.n2489 vdd.n1145 39.2114
R19259 vdd.n2485 vdd.n1146 39.2114
R19260 vdd.n2481 vdd.n1147 39.2114
R19261 vdd.n2477 vdd.n1148 39.2114
R19262 vdd.n1321 vdd.n1149 39.2114
R19263 vdd.n1325 vdd.n1150 39.2114
R19264 vdd.n1329 vdd.n1151 39.2114
R19265 vdd.n1333 vdd.n1152 39.2114
R19266 vdd.n1337 vdd.n1153 39.2114
R19267 vdd.n1341 vdd.n1154 39.2114
R19268 vdd.n1345 vdd.n1155 39.2114
R19269 vdd.n1350 vdd.n1156 39.2114
R19270 vdd.n1354 vdd.n1157 39.2114
R19271 vdd.n2717 vdd.n981 39.2114
R19272 vdd.n2722 vdd.n982 39.2114
R19273 vdd.n2726 vdd.n983 39.2114
R19274 vdd.n2730 vdd.n984 39.2114
R19275 vdd.n2734 vdd.n985 39.2114
R19276 vdd.n2738 vdd.n986 39.2114
R19277 vdd.n2742 vdd.n987 39.2114
R19278 vdd.n2746 vdd.n988 39.2114
R19279 vdd.n2750 vdd.n989 39.2114
R19280 vdd.n2754 vdd.n990 39.2114
R19281 vdd.n2758 vdd.n991 39.2114
R19282 vdd.n2762 vdd.n992 39.2114
R19283 vdd.n2766 vdd.n993 39.2114
R19284 vdd.n2770 vdd.n994 39.2114
R19285 vdd.n2774 vdd.n995 39.2114
R19286 vdd.n2778 vdd.n996 39.2114
R19287 vdd.n999 vdd.n997 39.2114
R19288 vdd.n3089 vdd.n962 39.2114
R19289 vdd.n3083 vdd.n2785 39.2114
R19290 vdd.n3079 vdd.n2786 39.2114
R19291 vdd.n3075 vdd.n2787 39.2114
R19292 vdd.n3071 vdd.n2788 39.2114
R19293 vdd.n3067 vdd.n2789 39.2114
R19294 vdd.n3063 vdd.n2790 39.2114
R19295 vdd.n3059 vdd.n2791 39.2114
R19296 vdd.n3055 vdd.n2792 39.2114
R19297 vdd.n3051 vdd.n2793 39.2114
R19298 vdd.n3047 vdd.n2794 39.2114
R19299 vdd.n3043 vdd.n2795 39.2114
R19300 vdd.n3039 vdd.n2796 39.2114
R19301 vdd.n3035 vdd.n2797 39.2114
R19302 vdd.n3031 vdd.n2798 39.2114
R19303 vdd.n3026 vdd.n2799 39.2114
R19304 vdd.n3022 vdd.n2800 39.2114
R19305 vdd.n3269 vdd.n3268 39.2114
R19306 vdd.n835 vdd.n831 39.2114
R19307 vdd.n3277 vdd.n3276 39.2114
R19308 vdd.n830 vdd.n828 39.2114
R19309 vdd.n3284 vdd.n3283 39.2114
R19310 vdd.n827 vdd.n825 39.2114
R19311 vdd.n3291 vdd.n3290 39.2114
R19312 vdd.n824 vdd.n822 39.2114
R19313 vdd.n3298 vdd.n3297 39.2114
R19314 vdd.n3302 vdd.n3301 39.2114
R19315 vdd.n821 vdd.n819 39.2114
R19316 vdd.n3309 vdd.n3308 39.2114
R19317 vdd.n818 vdd.n816 39.2114
R19318 vdd.n3316 vdd.n3315 39.2114
R19319 vdd.n815 vdd.n813 39.2114
R19320 vdd.n3323 vdd.n3322 39.2114
R19321 vdd.n3326 vdd.n3325 39.2114
R19322 vdd.n1008 vdd.n963 39.2114
R19323 vdd.n2706 vdd.n964 39.2114
R19324 vdd.n2702 vdd.n965 39.2114
R19325 vdd.n2698 vdd.n966 39.2114
R19326 vdd.n2694 vdd.n967 39.2114
R19327 vdd.n2690 vdd.n968 39.2114
R19328 vdd.n2686 vdd.n969 39.2114
R19329 vdd.n2682 vdd.n970 39.2114
R19330 vdd.n2678 vdd.n971 39.2114
R19331 vdd.n2674 vdd.n972 39.2114
R19332 vdd.n2670 vdd.n973 39.2114
R19333 vdd.n2666 vdd.n974 39.2114
R19334 vdd.n2662 vdd.n975 39.2114
R19335 vdd.n2658 vdd.n976 39.2114
R19336 vdd.n2654 vdd.n977 39.2114
R19337 vdd.n2650 vdd.n978 39.2114
R19338 vdd.n2646 vdd.n979 39.2114
R19339 vdd.n1280 vdd.n1158 39.2114
R19340 vdd.n1284 vdd.n1159 39.2114
R19341 vdd.n1288 vdd.n1160 39.2114
R19342 vdd.n1292 vdd.n1161 39.2114
R19343 vdd.n1296 vdd.n1162 39.2114
R19344 vdd.n1300 vdd.n1163 39.2114
R19345 vdd.n1304 vdd.n1164 39.2114
R19346 vdd.n1308 vdd.n1165 39.2114
R19347 vdd.n1312 vdd.n1166 39.2114
R19348 vdd.n1513 vdd.n1167 39.2114
R19349 vdd.n1510 vdd.n1168 39.2114
R19350 vdd.n1506 vdd.n1169 39.2114
R19351 vdd.n1502 vdd.n1170 39.2114
R19352 vdd.n1498 vdd.n1171 39.2114
R19353 vdd.n1494 vdd.n1172 39.2114
R19354 vdd.n1490 vdd.n1173 39.2114
R19355 vdd.n1486 vdd.n1174 39.2114
R19356 vdd.n2643 vdd.n979 39.2114
R19357 vdd.n2647 vdd.n978 39.2114
R19358 vdd.n2651 vdd.n977 39.2114
R19359 vdd.n2655 vdd.n976 39.2114
R19360 vdd.n2659 vdd.n975 39.2114
R19361 vdd.n2663 vdd.n974 39.2114
R19362 vdd.n2667 vdd.n973 39.2114
R19363 vdd.n2671 vdd.n972 39.2114
R19364 vdd.n2675 vdd.n971 39.2114
R19365 vdd.n2679 vdd.n970 39.2114
R19366 vdd.n2683 vdd.n969 39.2114
R19367 vdd.n2687 vdd.n968 39.2114
R19368 vdd.n2691 vdd.n967 39.2114
R19369 vdd.n2695 vdd.n966 39.2114
R19370 vdd.n2699 vdd.n965 39.2114
R19371 vdd.n2703 vdd.n964 39.2114
R19372 vdd.n2707 vdd.n963 39.2114
R19373 vdd.n1283 vdd.n1158 39.2114
R19374 vdd.n1287 vdd.n1159 39.2114
R19375 vdd.n1291 vdd.n1160 39.2114
R19376 vdd.n1295 vdd.n1161 39.2114
R19377 vdd.n1299 vdd.n1162 39.2114
R19378 vdd.n1303 vdd.n1163 39.2114
R19379 vdd.n1307 vdd.n1164 39.2114
R19380 vdd.n1311 vdd.n1165 39.2114
R19381 vdd.n1314 vdd.n1166 39.2114
R19382 vdd.n1511 vdd.n1167 39.2114
R19383 vdd.n1507 vdd.n1168 39.2114
R19384 vdd.n1503 vdd.n1169 39.2114
R19385 vdd.n1499 vdd.n1170 39.2114
R19386 vdd.n1495 vdd.n1171 39.2114
R19387 vdd.n1491 vdd.n1172 39.2114
R19388 vdd.n1487 vdd.n1173 39.2114
R19389 vdd.n1483 vdd.n1174 39.2114
R19390 vdd.n2364 vdd.n2363 37.2369
R19391 vdd.n2400 vdd.n1249 37.2369
R19392 vdd.n2439 vdd.n1209 37.2369
R19393 vdd.n3410 vdd.n769 37.2369
R19394 vdd.n3458 vdd.n3457 37.2369
R19395 vdd.n690 vdd.n689 37.2369
R19396 vdd.n1317 vdd.n1316 30.449
R19397 vdd.n1012 vdd.n1011 30.449
R19398 vdd.n1348 vdd.n1320 30.449
R19399 vdd.n2720 vdd.n1002 30.449
R19400 vdd.n2825 vdd.n2824 30.449
R19401 vdd.n3272 vdd.n833 30.449
R19402 vdd.n3028 vdd.n2821 30.449
R19403 vdd.n801 vdd.n800 30.449
R19404 vdd.n2510 vdd.n2509 29.8151
R19405 vdd.n2782 vdd.n1000 29.8151
R19406 vdd.n2715 vdd.n1003 29.8151
R19407 vdd.n1356 vdd.n1353 29.8151
R19408 vdd.n3023 vdd.n3020 29.8151
R19409 vdd.n3266 vdd.n3265 29.8151
R19410 vdd.n3092 vdd.n3091 29.8151
R19411 vdd.n3329 vdd.n3328 29.8151
R19412 vdd.n3248 vdd.n3247 29.8151
R19413 vdd.n3334 vdd.n802 29.8151
R19414 vdd.n2896 vdd.n2894 29.8151
R19415 vdd.n2827 vdd.n955 29.8151
R19416 vdd.n1281 vdd.n1132 29.8151
R19417 vdd.n2710 vdd.n2709 29.8151
R19418 vdd.n2642 vdd.n2641 29.8151
R19419 vdd.n1482 vdd.n1481 29.8151
R19420 vdd.n1873 vdd.n1680 22.2201
R19421 vdd.n2358 vdd.n1141 22.2201
R19422 vdd.n3495 vdd.n723 22.2201
R19423 vdd.n3627 vdd.n3626 22.2201
R19424 vdd.n1884 vdd.n1642 19.3944
R19425 vdd.n1884 vdd.n1640 19.3944
R19426 vdd.n1888 vdd.n1640 19.3944
R19427 vdd.n1888 vdd.n1630 19.3944
R19428 vdd.n1901 vdd.n1630 19.3944
R19429 vdd.n1901 vdd.n1628 19.3944
R19430 vdd.n1905 vdd.n1628 19.3944
R19431 vdd.n1905 vdd.n1620 19.3944
R19432 vdd.n1918 vdd.n1620 19.3944
R19433 vdd.n1918 vdd.n1618 19.3944
R19434 vdd.n1922 vdd.n1618 19.3944
R19435 vdd.n1922 vdd.n1607 19.3944
R19436 vdd.n1934 vdd.n1607 19.3944
R19437 vdd.n1934 vdd.n1605 19.3944
R19438 vdd.n1938 vdd.n1605 19.3944
R19439 vdd.n1938 vdd.n1596 19.3944
R19440 vdd.n1951 vdd.n1596 19.3944
R19441 vdd.n1951 vdd.n1594 19.3944
R19442 vdd.n1955 vdd.n1594 19.3944
R19443 vdd.n1955 vdd.n1585 19.3944
R19444 vdd.n2274 vdd.n1585 19.3944
R19445 vdd.n2274 vdd.n1583 19.3944
R19446 vdd.n2278 vdd.n1583 19.3944
R19447 vdd.n2278 vdd.n1573 19.3944
R19448 vdd.n2291 vdd.n1573 19.3944
R19449 vdd.n2291 vdd.n1571 19.3944
R19450 vdd.n2295 vdd.n1571 19.3944
R19451 vdd.n2295 vdd.n1563 19.3944
R19452 vdd.n2308 vdd.n1563 19.3944
R19453 vdd.n2308 vdd.n1561 19.3944
R19454 vdd.n2312 vdd.n1561 19.3944
R19455 vdd.n2312 vdd.n1550 19.3944
R19456 vdd.n2324 vdd.n1550 19.3944
R19457 vdd.n2324 vdd.n1548 19.3944
R19458 vdd.n2328 vdd.n1548 19.3944
R19459 vdd.n2328 vdd.n1540 19.3944
R19460 vdd.n2341 vdd.n1540 19.3944
R19461 vdd.n2341 vdd.n1537 19.3944
R19462 vdd.n2347 vdd.n1537 19.3944
R19463 vdd.n2347 vdd.n1538 19.3944
R19464 vdd.n1538 vdd.n1528 19.3944
R19465 vdd.n1808 vdd.n1743 19.3944
R19466 vdd.n1804 vdd.n1743 19.3944
R19467 vdd.n1804 vdd.n1803 19.3944
R19468 vdd.n1803 vdd.n1802 19.3944
R19469 vdd.n1802 vdd.n1749 19.3944
R19470 vdd.n1798 vdd.n1749 19.3944
R19471 vdd.n1798 vdd.n1797 19.3944
R19472 vdd.n1797 vdd.n1796 19.3944
R19473 vdd.n1796 vdd.n1755 19.3944
R19474 vdd.n1792 vdd.n1755 19.3944
R19475 vdd.n1792 vdd.n1791 19.3944
R19476 vdd.n1791 vdd.n1790 19.3944
R19477 vdd.n1790 vdd.n1761 19.3944
R19478 vdd.n1786 vdd.n1761 19.3944
R19479 vdd.n1786 vdd.n1785 19.3944
R19480 vdd.n1785 vdd.n1784 19.3944
R19481 vdd.n1784 vdd.n1767 19.3944
R19482 vdd.n1780 vdd.n1767 19.3944
R19483 vdd.n1780 vdd.n1779 19.3944
R19484 vdd.n1779 vdd.n1778 19.3944
R19485 vdd.n1843 vdd.n1842 19.3944
R19486 vdd.n1842 vdd.n1841 19.3944
R19487 vdd.n1841 vdd.n1714 19.3944
R19488 vdd.n1837 vdd.n1714 19.3944
R19489 vdd.n1837 vdd.n1836 19.3944
R19490 vdd.n1836 vdd.n1835 19.3944
R19491 vdd.n1835 vdd.n1720 19.3944
R19492 vdd.n1831 vdd.n1720 19.3944
R19493 vdd.n1831 vdd.n1830 19.3944
R19494 vdd.n1830 vdd.n1829 19.3944
R19495 vdd.n1829 vdd.n1726 19.3944
R19496 vdd.n1825 vdd.n1726 19.3944
R19497 vdd.n1825 vdd.n1824 19.3944
R19498 vdd.n1824 vdd.n1823 19.3944
R19499 vdd.n1823 vdd.n1732 19.3944
R19500 vdd.n1819 vdd.n1732 19.3944
R19501 vdd.n1819 vdd.n1818 19.3944
R19502 vdd.n1818 vdd.n1817 19.3944
R19503 vdd.n1817 vdd.n1738 19.3944
R19504 vdd.n1813 vdd.n1738 19.3944
R19505 vdd.n1876 vdd.n1647 19.3944
R19506 vdd.n1871 vdd.n1647 19.3944
R19507 vdd.n1871 vdd.n1682 19.3944
R19508 vdd.n1867 vdd.n1682 19.3944
R19509 vdd.n1867 vdd.n1866 19.3944
R19510 vdd.n1866 vdd.n1865 19.3944
R19511 vdd.n1865 vdd.n1688 19.3944
R19512 vdd.n1861 vdd.n1688 19.3944
R19513 vdd.n1861 vdd.n1860 19.3944
R19514 vdd.n1860 vdd.n1859 19.3944
R19515 vdd.n1859 vdd.n1694 19.3944
R19516 vdd.n1855 vdd.n1694 19.3944
R19517 vdd.n1855 vdd.n1854 19.3944
R19518 vdd.n1854 vdd.n1853 19.3944
R19519 vdd.n1853 vdd.n1700 19.3944
R19520 vdd.n1849 vdd.n1700 19.3944
R19521 vdd.n1849 vdd.n1848 19.3944
R19522 vdd.n1848 vdd.n1847 19.3944
R19523 vdd.n2396 vdd.n1247 19.3944
R19524 vdd.n2396 vdd.n1253 19.3944
R19525 vdd.n2391 vdd.n1253 19.3944
R19526 vdd.n2391 vdd.n2390 19.3944
R19527 vdd.n2390 vdd.n2389 19.3944
R19528 vdd.n2389 vdd.n1260 19.3944
R19529 vdd.n2384 vdd.n1260 19.3944
R19530 vdd.n2384 vdd.n2383 19.3944
R19531 vdd.n2383 vdd.n2382 19.3944
R19532 vdd.n2382 vdd.n1267 19.3944
R19533 vdd.n2377 vdd.n1267 19.3944
R19534 vdd.n2377 vdd.n2376 19.3944
R19535 vdd.n2376 vdd.n2375 19.3944
R19536 vdd.n2375 vdd.n1274 19.3944
R19537 vdd.n2370 vdd.n1274 19.3944
R19538 vdd.n2370 vdd.n2369 19.3944
R19539 vdd.n1521 vdd.n1279 19.3944
R19540 vdd.n2365 vdd.n1518 19.3944
R19541 vdd.n2435 vdd.n1207 19.3944
R19542 vdd.n2435 vdd.n1213 19.3944
R19543 vdd.n2430 vdd.n1213 19.3944
R19544 vdd.n2430 vdd.n2429 19.3944
R19545 vdd.n2429 vdd.n2428 19.3944
R19546 vdd.n2428 vdd.n1220 19.3944
R19547 vdd.n2423 vdd.n1220 19.3944
R19548 vdd.n2423 vdd.n2422 19.3944
R19549 vdd.n2422 vdd.n2421 19.3944
R19550 vdd.n2421 vdd.n1227 19.3944
R19551 vdd.n2416 vdd.n1227 19.3944
R19552 vdd.n2416 vdd.n2415 19.3944
R19553 vdd.n2415 vdd.n2414 19.3944
R19554 vdd.n2414 vdd.n1234 19.3944
R19555 vdd.n2409 vdd.n1234 19.3944
R19556 vdd.n2409 vdd.n2408 19.3944
R19557 vdd.n2408 vdd.n2407 19.3944
R19558 vdd.n2407 vdd.n1241 19.3944
R19559 vdd.n2402 vdd.n1241 19.3944
R19560 vdd.n2402 vdd.n2401 19.3944
R19561 vdd.n2472 vdd.n1182 19.3944
R19562 vdd.n2472 vdd.n1183 19.3944
R19563 vdd.n2467 vdd.n2466 19.3944
R19564 vdd.n2462 vdd.n2461 19.3944
R19565 vdd.n2461 vdd.n2460 19.3944
R19566 vdd.n2460 vdd.n1187 19.3944
R19567 vdd.n2455 vdd.n1187 19.3944
R19568 vdd.n2455 vdd.n2454 19.3944
R19569 vdd.n2454 vdd.n2453 19.3944
R19570 vdd.n2453 vdd.n1194 19.3944
R19571 vdd.n2448 vdd.n1194 19.3944
R19572 vdd.n2448 vdd.n2447 19.3944
R19573 vdd.n2447 vdd.n2446 19.3944
R19574 vdd.n2446 vdd.n1201 19.3944
R19575 vdd.n2441 vdd.n1201 19.3944
R19576 vdd.n2441 vdd.n2440 19.3944
R19577 vdd.n1880 vdd.n1645 19.3944
R19578 vdd.n1880 vdd.n1636 19.3944
R19579 vdd.n1893 vdd.n1636 19.3944
R19580 vdd.n1893 vdd.n1634 19.3944
R19581 vdd.n1897 vdd.n1634 19.3944
R19582 vdd.n1897 vdd.n1625 19.3944
R19583 vdd.n1910 vdd.n1625 19.3944
R19584 vdd.n1910 vdd.n1623 19.3944
R19585 vdd.n1914 vdd.n1623 19.3944
R19586 vdd.n1914 vdd.n1614 19.3944
R19587 vdd.n1926 vdd.n1614 19.3944
R19588 vdd.n1926 vdd.n1612 19.3944
R19589 vdd.n1930 vdd.n1612 19.3944
R19590 vdd.n1930 vdd.n1602 19.3944
R19591 vdd.n1943 vdd.n1602 19.3944
R19592 vdd.n1943 vdd.n1600 19.3944
R19593 vdd.n1947 vdd.n1600 19.3944
R19594 vdd.n1947 vdd.n1591 19.3944
R19595 vdd.n1959 vdd.n1591 19.3944
R19596 vdd.n1959 vdd.n1589 19.3944
R19597 vdd.n2270 vdd.n1589 19.3944
R19598 vdd.n2270 vdd.n1579 19.3944
R19599 vdd.n2283 vdd.n1579 19.3944
R19600 vdd.n2283 vdd.n1577 19.3944
R19601 vdd.n2287 vdd.n1577 19.3944
R19602 vdd.n2287 vdd.n1568 19.3944
R19603 vdd.n2300 vdd.n1568 19.3944
R19604 vdd.n2300 vdd.n1566 19.3944
R19605 vdd.n2304 vdd.n1566 19.3944
R19606 vdd.n2304 vdd.n1557 19.3944
R19607 vdd.n2316 vdd.n1557 19.3944
R19608 vdd.n2316 vdd.n1555 19.3944
R19609 vdd.n2320 vdd.n1555 19.3944
R19610 vdd.n2320 vdd.n1545 19.3944
R19611 vdd.n2333 vdd.n1545 19.3944
R19612 vdd.n2333 vdd.n1543 19.3944
R19613 vdd.n2337 vdd.n1543 19.3944
R19614 vdd.n2337 vdd.n1533 19.3944
R19615 vdd.n2352 vdd.n1533 19.3944
R19616 vdd.n2352 vdd.n1531 19.3944
R19617 vdd.n2356 vdd.n1531 19.3944
R19618 vdd.n3501 vdd.n686 19.3944
R19619 vdd.n3501 vdd.n676 19.3944
R19620 vdd.n3513 vdd.n676 19.3944
R19621 vdd.n3513 vdd.n674 19.3944
R19622 vdd.n3517 vdd.n674 19.3944
R19623 vdd.n3517 vdd.n666 19.3944
R19624 vdd.n3530 vdd.n666 19.3944
R19625 vdd.n3530 vdd.n664 19.3944
R19626 vdd.n3534 vdd.n664 19.3944
R19627 vdd.n3534 vdd.n653 19.3944
R19628 vdd.n3546 vdd.n653 19.3944
R19629 vdd.n3546 vdd.n651 19.3944
R19630 vdd.n3550 vdd.n651 19.3944
R19631 vdd.n3550 vdd.n642 19.3944
R19632 vdd.n3563 vdd.n642 19.3944
R19633 vdd.n3563 vdd.n640 19.3944
R19634 vdd.n3570 vdd.n640 19.3944
R19635 vdd.n3570 vdd.n3569 19.3944
R19636 vdd.n3569 vdd.n631 19.3944
R19637 vdd.n3583 vdd.n631 19.3944
R19638 vdd.n3584 vdd.n3583 19.3944
R19639 vdd.n3584 vdd.n629 19.3944
R19640 vdd.n3588 vdd.n629 19.3944
R19641 vdd.n3590 vdd.n3588 19.3944
R19642 vdd.n3591 vdd.n3590 19.3944
R19643 vdd.n3591 vdd.n627 19.3944
R19644 vdd.n3595 vdd.n627 19.3944
R19645 vdd.n3597 vdd.n3595 19.3944
R19646 vdd.n3598 vdd.n3597 19.3944
R19647 vdd.n3598 vdd.n625 19.3944
R19648 vdd.n3602 vdd.n625 19.3944
R19649 vdd.n3605 vdd.n3602 19.3944
R19650 vdd.n3606 vdd.n3605 19.3944
R19651 vdd.n3606 vdd.n623 19.3944
R19652 vdd.n3610 vdd.n623 19.3944
R19653 vdd.n3612 vdd.n3610 19.3944
R19654 vdd.n3613 vdd.n3612 19.3944
R19655 vdd.n3613 vdd.n621 19.3944
R19656 vdd.n3617 vdd.n621 19.3944
R19657 vdd.n3619 vdd.n3617 19.3944
R19658 vdd.n3620 vdd.n3619 19.3944
R19659 vdd.n569 vdd.n438 19.3944
R19660 vdd.n575 vdd.n438 19.3944
R19661 vdd.n576 vdd.n575 19.3944
R19662 vdd.n579 vdd.n576 19.3944
R19663 vdd.n579 vdd.n436 19.3944
R19664 vdd.n585 vdd.n436 19.3944
R19665 vdd.n586 vdd.n585 19.3944
R19666 vdd.n589 vdd.n586 19.3944
R19667 vdd.n589 vdd.n434 19.3944
R19668 vdd.n595 vdd.n434 19.3944
R19669 vdd.n596 vdd.n595 19.3944
R19670 vdd.n599 vdd.n596 19.3944
R19671 vdd.n599 vdd.n432 19.3944
R19672 vdd.n605 vdd.n432 19.3944
R19673 vdd.n606 vdd.n605 19.3944
R19674 vdd.n609 vdd.n606 19.3944
R19675 vdd.n609 vdd.n430 19.3944
R19676 vdd.n615 vdd.n430 19.3944
R19677 vdd.n617 vdd.n615 19.3944
R19678 vdd.n618 vdd.n617 19.3944
R19679 vdd.n516 vdd.n515 19.3944
R19680 vdd.n519 vdd.n516 19.3944
R19681 vdd.n519 vdd.n450 19.3944
R19682 vdd.n525 vdd.n450 19.3944
R19683 vdd.n526 vdd.n525 19.3944
R19684 vdd.n529 vdd.n526 19.3944
R19685 vdd.n529 vdd.n448 19.3944
R19686 vdd.n535 vdd.n448 19.3944
R19687 vdd.n536 vdd.n535 19.3944
R19688 vdd.n539 vdd.n536 19.3944
R19689 vdd.n539 vdd.n446 19.3944
R19690 vdd.n545 vdd.n446 19.3944
R19691 vdd.n546 vdd.n545 19.3944
R19692 vdd.n549 vdd.n546 19.3944
R19693 vdd.n549 vdd.n444 19.3944
R19694 vdd.n555 vdd.n444 19.3944
R19695 vdd.n556 vdd.n555 19.3944
R19696 vdd.n559 vdd.n556 19.3944
R19697 vdd.n559 vdd.n442 19.3944
R19698 vdd.n565 vdd.n442 19.3944
R19699 vdd.n466 vdd.n465 19.3944
R19700 vdd.n469 vdd.n466 19.3944
R19701 vdd.n469 vdd.n462 19.3944
R19702 vdd.n475 vdd.n462 19.3944
R19703 vdd.n476 vdd.n475 19.3944
R19704 vdd.n479 vdd.n476 19.3944
R19705 vdd.n479 vdd.n460 19.3944
R19706 vdd.n485 vdd.n460 19.3944
R19707 vdd.n486 vdd.n485 19.3944
R19708 vdd.n489 vdd.n486 19.3944
R19709 vdd.n489 vdd.n458 19.3944
R19710 vdd.n495 vdd.n458 19.3944
R19711 vdd.n496 vdd.n495 19.3944
R19712 vdd.n499 vdd.n496 19.3944
R19713 vdd.n499 vdd.n456 19.3944
R19714 vdd.n505 vdd.n456 19.3944
R19715 vdd.n506 vdd.n505 19.3944
R19716 vdd.n509 vdd.n506 19.3944
R19717 vdd.n3505 vdd.n683 19.3944
R19718 vdd.n3505 vdd.n681 19.3944
R19719 vdd.n3509 vdd.n681 19.3944
R19720 vdd.n3509 vdd.n671 19.3944
R19721 vdd.n3522 vdd.n671 19.3944
R19722 vdd.n3522 vdd.n669 19.3944
R19723 vdd.n3526 vdd.n669 19.3944
R19724 vdd.n3526 vdd.n660 19.3944
R19725 vdd.n3538 vdd.n660 19.3944
R19726 vdd.n3538 vdd.n658 19.3944
R19727 vdd.n3542 vdd.n658 19.3944
R19728 vdd.n3542 vdd.n648 19.3944
R19729 vdd.n3555 vdd.n648 19.3944
R19730 vdd.n3555 vdd.n646 19.3944
R19731 vdd.n3559 vdd.n646 19.3944
R19732 vdd.n3559 vdd.n637 19.3944
R19733 vdd.n3574 vdd.n637 19.3944
R19734 vdd.n3574 vdd.n635 19.3944
R19735 vdd.n3578 vdd.n635 19.3944
R19736 vdd.n3578 vdd.n336 19.3944
R19737 vdd.n3669 vdd.n336 19.3944
R19738 vdd.n3669 vdd.n337 19.3944
R19739 vdd.n3663 vdd.n337 19.3944
R19740 vdd.n3663 vdd.n3662 19.3944
R19741 vdd.n3662 vdd.n3661 19.3944
R19742 vdd.n3661 vdd.n349 19.3944
R19743 vdd.n3655 vdd.n349 19.3944
R19744 vdd.n3655 vdd.n3654 19.3944
R19745 vdd.n3654 vdd.n3653 19.3944
R19746 vdd.n3653 vdd.n359 19.3944
R19747 vdd.n3647 vdd.n359 19.3944
R19748 vdd.n3647 vdd.n3646 19.3944
R19749 vdd.n3646 vdd.n3645 19.3944
R19750 vdd.n3645 vdd.n370 19.3944
R19751 vdd.n3639 vdd.n370 19.3944
R19752 vdd.n3639 vdd.n3638 19.3944
R19753 vdd.n3638 vdd.n3637 19.3944
R19754 vdd.n3637 vdd.n381 19.3944
R19755 vdd.n3631 vdd.n381 19.3944
R19756 vdd.n3631 vdd.n3630 19.3944
R19757 vdd.n3630 vdd.n3629 19.3944
R19758 vdd.n3452 vdd.n747 19.3944
R19759 vdd.n3452 vdd.n3449 19.3944
R19760 vdd.n3449 vdd.n3446 19.3944
R19761 vdd.n3446 vdd.n3445 19.3944
R19762 vdd.n3445 vdd.n3442 19.3944
R19763 vdd.n3442 vdd.n3441 19.3944
R19764 vdd.n3441 vdd.n3438 19.3944
R19765 vdd.n3438 vdd.n3437 19.3944
R19766 vdd.n3437 vdd.n3434 19.3944
R19767 vdd.n3434 vdd.n3433 19.3944
R19768 vdd.n3433 vdd.n3430 19.3944
R19769 vdd.n3430 vdd.n3429 19.3944
R19770 vdd.n3429 vdd.n3426 19.3944
R19771 vdd.n3426 vdd.n3425 19.3944
R19772 vdd.n3425 vdd.n3422 19.3944
R19773 vdd.n3422 vdd.n3421 19.3944
R19774 vdd.n3421 vdd.n3418 19.3944
R19775 vdd.n3418 vdd.n3417 19.3944
R19776 vdd.n3417 vdd.n3414 19.3944
R19777 vdd.n3414 vdd.n3413 19.3944
R19778 vdd.n3492 vdd.n3491 19.3944
R19779 vdd.n3491 vdd.n3490 19.3944
R19780 vdd.n732 vdd.n729 19.3944
R19781 vdd.n3486 vdd.n3485 19.3944
R19782 vdd.n3485 vdd.n3482 19.3944
R19783 vdd.n3482 vdd.n3481 19.3944
R19784 vdd.n3481 vdd.n3478 19.3944
R19785 vdd.n3478 vdd.n3477 19.3944
R19786 vdd.n3477 vdd.n3474 19.3944
R19787 vdd.n3474 vdd.n3473 19.3944
R19788 vdd.n3473 vdd.n3470 19.3944
R19789 vdd.n3470 vdd.n3469 19.3944
R19790 vdd.n3469 vdd.n3466 19.3944
R19791 vdd.n3466 vdd.n3465 19.3944
R19792 vdd.n3465 vdd.n3462 19.3944
R19793 vdd.n3462 vdd.n3461 19.3944
R19794 vdd.n3406 vdd.n767 19.3944
R19795 vdd.n3406 vdd.n3403 19.3944
R19796 vdd.n3403 vdd.n3400 19.3944
R19797 vdd.n3400 vdd.n3399 19.3944
R19798 vdd.n3399 vdd.n3396 19.3944
R19799 vdd.n3396 vdd.n3395 19.3944
R19800 vdd.n3395 vdd.n3392 19.3944
R19801 vdd.n3392 vdd.n3391 19.3944
R19802 vdd.n3391 vdd.n3388 19.3944
R19803 vdd.n3388 vdd.n3387 19.3944
R19804 vdd.n3387 vdd.n3384 19.3944
R19805 vdd.n3384 vdd.n3383 19.3944
R19806 vdd.n3383 vdd.n3380 19.3944
R19807 vdd.n3380 vdd.n3379 19.3944
R19808 vdd.n3379 vdd.n3376 19.3944
R19809 vdd.n3376 vdd.n3375 19.3944
R19810 vdd.n3372 vdd.n3371 19.3944
R19811 vdd.n3368 vdd.n3367 19.3944
R19812 vdd.n1812 vdd.n1808 19.0066
R19813 vdd.n2400 vdd.n1247 19.0066
R19814 vdd.n569 vdd.n566 19.0066
R19815 vdd.n3410 vdd.n767 19.0066
R19816 vdd.n1316 vdd.n1315 16.0975
R19817 vdd.n1011 vdd.n1010 16.0975
R19818 vdd.n1773 vdd.n1772 16.0975
R19819 vdd.n1811 vdd.n1810 16.0975
R19820 vdd.n1707 vdd.n1706 16.0975
R19821 vdd.n2363 vdd.n2362 16.0975
R19822 vdd.n1249 vdd.n1248 16.0975
R19823 vdd.n1209 vdd.n1208 16.0975
R19824 vdd.n1320 vdd.n1319 16.0975
R19825 vdd.n1002 vdd.n1001 16.0975
R19826 vdd.n2824 vdd.n2823 16.0975
R19827 vdd.n427 vdd.n426 16.0975
R19828 vdd.n441 vdd.n440 16.0975
R19829 vdd.n453 vdd.n452 16.0975
R19830 vdd.n769 vdd.n768 16.0975
R19831 vdd.n3457 vdd.n3456 16.0975
R19832 vdd.n833 vdd.n832 16.0975
R19833 vdd.n2821 vdd.n2820 16.0975
R19834 vdd.n689 vdd.n688 16.0975
R19835 vdd.n800 vdd.n799 16.0975
R19836 vdd.t278 vdd.n2784 15.4182
R19837 vdd.n3088 vdd.t263 15.4182
R19838 vdd.n28 vdd.n27 15.0023
R19839 vdd.n328 vdd.n293 13.1884
R19840 vdd.n269 vdd.n234 13.1884
R19841 vdd.n226 vdd.n191 13.1884
R19842 vdd.n167 vdd.n132 13.1884
R19843 vdd.n125 vdd.n90 13.1884
R19844 vdd.n66 vdd.n31 13.1884
R19845 vdd.n2202 vdd.n2167 13.1884
R19846 vdd.n2261 vdd.n2226 13.1884
R19847 vdd.n2100 vdd.n2065 13.1884
R19848 vdd.n2159 vdd.n2124 13.1884
R19849 vdd.n1999 vdd.n1964 13.1884
R19850 vdd.n2058 vdd.n2023 13.1884
R19851 vdd.n2506 vdd.n1134 13.1509
R19852 vdd.n3331 vdd.n692 13.1509
R19853 vdd.n1843 vdd.n1708 12.9944
R19854 vdd.n1847 vdd.n1708 12.9944
R19855 vdd.n2439 vdd.n1207 12.9944
R19856 vdd.n2440 vdd.n2439 12.9944
R19857 vdd.n515 vdd.n454 12.9944
R19858 vdd.n509 vdd.n454 12.9944
R19859 vdd.n3458 vdd.n747 12.9944
R19860 vdd.n3461 vdd.n3458 12.9944
R19861 vdd.n329 vdd.n291 12.8005
R19862 vdd.n324 vdd.n295 12.8005
R19863 vdd.n270 vdd.n232 12.8005
R19864 vdd.n265 vdd.n236 12.8005
R19865 vdd.n227 vdd.n189 12.8005
R19866 vdd.n222 vdd.n193 12.8005
R19867 vdd.n168 vdd.n130 12.8005
R19868 vdd.n163 vdd.n134 12.8005
R19869 vdd.n126 vdd.n88 12.8005
R19870 vdd.n121 vdd.n92 12.8005
R19871 vdd.n67 vdd.n29 12.8005
R19872 vdd.n62 vdd.n33 12.8005
R19873 vdd.n2203 vdd.n2165 12.8005
R19874 vdd.n2198 vdd.n2169 12.8005
R19875 vdd.n2262 vdd.n2224 12.8005
R19876 vdd.n2257 vdd.n2228 12.8005
R19877 vdd.n2101 vdd.n2063 12.8005
R19878 vdd.n2096 vdd.n2067 12.8005
R19879 vdd.n2160 vdd.n2122 12.8005
R19880 vdd.n2155 vdd.n2126 12.8005
R19881 vdd.n2000 vdd.n1962 12.8005
R19882 vdd.n1995 vdd.n1966 12.8005
R19883 vdd.n2059 vdd.n2021 12.8005
R19884 vdd.n2054 vdd.n2025 12.8005
R19885 vdd.n323 vdd.n296 12.0247
R19886 vdd.n264 vdd.n237 12.0247
R19887 vdd.n221 vdd.n194 12.0247
R19888 vdd.n162 vdd.n135 12.0247
R19889 vdd.n120 vdd.n93 12.0247
R19890 vdd.n61 vdd.n34 12.0247
R19891 vdd.n2197 vdd.n2170 12.0247
R19892 vdd.n2256 vdd.n2229 12.0247
R19893 vdd.n2095 vdd.n2068 12.0247
R19894 vdd.n2154 vdd.n2127 12.0247
R19895 vdd.n1994 vdd.n1967 12.0247
R19896 vdd.n2053 vdd.n2026 12.0247
R19897 vdd.n1882 vdd.n1638 11.337
R19898 vdd.n1891 vdd.n1638 11.337
R19899 vdd.n1891 vdd.n1890 11.337
R19900 vdd.n1899 vdd.n1632 11.337
R19901 vdd.n1908 vdd.n1907 11.337
R19902 vdd.n1924 vdd.n1616 11.337
R19903 vdd.n1932 vdd.n1609 11.337
R19904 vdd.n1941 vdd.n1940 11.337
R19905 vdd.n1949 vdd.n1598 11.337
R19906 vdd.n2272 vdd.n1587 11.337
R19907 vdd.n2281 vdd.n1581 11.337
R19908 vdd.n2289 vdd.n1575 11.337
R19909 vdd.n2298 vdd.n2297 11.337
R19910 vdd.n2314 vdd.n1559 11.337
R19911 vdd.n2322 vdd.n1552 11.337
R19912 vdd.n2331 vdd.n2330 11.337
R19913 vdd.n2339 vdd.n1535 11.337
R19914 vdd.n2350 vdd.n1535 11.337
R19915 vdd.n2350 vdd.n2349 11.337
R19916 vdd.n3503 vdd.n678 11.337
R19917 vdd.n3511 vdd.n678 11.337
R19918 vdd.n3511 vdd.n679 11.337
R19919 vdd.n3520 vdd.n3519 11.337
R19920 vdd.n3536 vdd.n662 11.337
R19921 vdd.n3544 vdd.n655 11.337
R19922 vdd.n3553 vdd.n3552 11.337
R19923 vdd.n3561 vdd.n644 11.337
R19924 vdd.n3580 vdd.n633 11.337
R19925 vdd.n3667 vdd.n340 11.337
R19926 vdd.n3665 vdd.n344 11.337
R19927 vdd.n3659 vdd.n3658 11.337
R19928 vdd.n3651 vdd.n361 11.337
R19929 vdd.n3650 vdd.n3649 11.337
R19930 vdd.n3643 vdd.n3642 11.337
R19931 vdd.n3641 vdd.n375 11.337
R19932 vdd.n3635 vdd.n3634 11.337
R19933 vdd.n3634 vdd.n3633 11.337
R19934 vdd.n3633 vdd.n386 11.337
R19935 vdd.n320 vdd.n319 11.249
R19936 vdd.n261 vdd.n260 11.249
R19937 vdd.n218 vdd.n217 11.249
R19938 vdd.n159 vdd.n158 11.249
R19939 vdd.n117 vdd.n116 11.249
R19940 vdd.n58 vdd.n57 11.249
R19941 vdd.n2194 vdd.n2193 11.249
R19942 vdd.n2253 vdd.n2252 11.249
R19943 vdd.n2092 vdd.n2091 11.249
R19944 vdd.n2151 vdd.n2150 11.249
R19945 vdd.n1991 vdd.n1990 11.249
R19946 vdd.n2050 vdd.n2049 11.249
R19947 vdd.n1680 vdd.t72 11.2237
R19948 vdd.n3627 vdd.t21 11.2237
R19949 vdd.t184 vdd.n1553 10.7702
R19950 vdd.n3528 vdd.t110 10.7702
R19951 vdd.n305 vdd.n304 10.7238
R19952 vdd.n246 vdd.n245 10.7238
R19953 vdd.n203 vdd.n202 10.7238
R19954 vdd.n144 vdd.n143 10.7238
R19955 vdd.n102 vdd.n101 10.7238
R19956 vdd.n43 vdd.n42 10.7238
R19957 vdd.n2179 vdd.n2178 10.7238
R19958 vdd.n2238 vdd.n2237 10.7238
R19959 vdd.n2077 vdd.n2076 10.7238
R19960 vdd.n2136 vdd.n2135 10.7238
R19961 vdd.n1976 vdd.n1975 10.7238
R19962 vdd.n2035 vdd.n2034 10.7238
R19963 vdd.n2511 vdd.n2510 10.6151
R19964 vdd.n2511 vdd.n1127 10.6151
R19965 vdd.n2521 vdd.n1127 10.6151
R19966 vdd.n2522 vdd.n2521 10.6151
R19967 vdd.n2523 vdd.n2522 10.6151
R19968 vdd.n2523 vdd.n1114 10.6151
R19969 vdd.n2533 vdd.n1114 10.6151
R19970 vdd.n2534 vdd.n2533 10.6151
R19971 vdd.n2535 vdd.n2534 10.6151
R19972 vdd.n2535 vdd.n1102 10.6151
R19973 vdd.n2545 vdd.n1102 10.6151
R19974 vdd.n2546 vdd.n2545 10.6151
R19975 vdd.n2547 vdd.n2546 10.6151
R19976 vdd.n2547 vdd.n1091 10.6151
R19977 vdd.n2557 vdd.n1091 10.6151
R19978 vdd.n2558 vdd.n2557 10.6151
R19979 vdd.n2559 vdd.n2558 10.6151
R19980 vdd.n2559 vdd.n1078 10.6151
R19981 vdd.n2569 vdd.n1078 10.6151
R19982 vdd.n2570 vdd.n2569 10.6151
R19983 vdd.n2571 vdd.n2570 10.6151
R19984 vdd.n2571 vdd.n1066 10.6151
R19985 vdd.n2582 vdd.n1066 10.6151
R19986 vdd.n2583 vdd.n2582 10.6151
R19987 vdd.n2584 vdd.n2583 10.6151
R19988 vdd.n2584 vdd.n1054 10.6151
R19989 vdd.n2594 vdd.n1054 10.6151
R19990 vdd.n2595 vdd.n2594 10.6151
R19991 vdd.n2596 vdd.n2595 10.6151
R19992 vdd.n2596 vdd.n1042 10.6151
R19993 vdd.n2606 vdd.n1042 10.6151
R19994 vdd.n2607 vdd.n2606 10.6151
R19995 vdd.n2608 vdd.n2607 10.6151
R19996 vdd.n2608 vdd.n1032 10.6151
R19997 vdd.n2618 vdd.n1032 10.6151
R19998 vdd.n2619 vdd.n2618 10.6151
R19999 vdd.n2620 vdd.n2619 10.6151
R20000 vdd.n2620 vdd.n1019 10.6151
R20001 vdd.n2632 vdd.n1019 10.6151
R20002 vdd.n2633 vdd.n2632 10.6151
R20003 vdd.n2635 vdd.n2633 10.6151
R20004 vdd.n2635 vdd.n2634 10.6151
R20005 vdd.n2634 vdd.n1000 10.6151
R20006 vdd.n2782 vdd.n2781 10.6151
R20007 vdd.n2781 vdd.n2780 10.6151
R20008 vdd.n2780 vdd.n2777 10.6151
R20009 vdd.n2777 vdd.n2776 10.6151
R20010 vdd.n2776 vdd.n2773 10.6151
R20011 vdd.n2773 vdd.n2772 10.6151
R20012 vdd.n2772 vdd.n2769 10.6151
R20013 vdd.n2769 vdd.n2768 10.6151
R20014 vdd.n2768 vdd.n2765 10.6151
R20015 vdd.n2765 vdd.n2764 10.6151
R20016 vdd.n2764 vdd.n2761 10.6151
R20017 vdd.n2761 vdd.n2760 10.6151
R20018 vdd.n2760 vdd.n2757 10.6151
R20019 vdd.n2757 vdd.n2756 10.6151
R20020 vdd.n2756 vdd.n2753 10.6151
R20021 vdd.n2753 vdd.n2752 10.6151
R20022 vdd.n2752 vdd.n2749 10.6151
R20023 vdd.n2749 vdd.n2748 10.6151
R20024 vdd.n2748 vdd.n2745 10.6151
R20025 vdd.n2745 vdd.n2744 10.6151
R20026 vdd.n2744 vdd.n2741 10.6151
R20027 vdd.n2741 vdd.n2740 10.6151
R20028 vdd.n2740 vdd.n2737 10.6151
R20029 vdd.n2737 vdd.n2736 10.6151
R20030 vdd.n2736 vdd.n2733 10.6151
R20031 vdd.n2733 vdd.n2732 10.6151
R20032 vdd.n2732 vdd.n2729 10.6151
R20033 vdd.n2729 vdd.n2728 10.6151
R20034 vdd.n2728 vdd.n2725 10.6151
R20035 vdd.n2725 vdd.n2724 10.6151
R20036 vdd.n2724 vdd.n2721 10.6151
R20037 vdd.n2719 vdd.n2716 10.6151
R20038 vdd.n2716 vdd.n2715 10.6151
R20039 vdd.n1357 vdd.n1356 10.6151
R20040 vdd.n1359 vdd.n1357 10.6151
R20041 vdd.n1360 vdd.n1359 10.6151
R20042 vdd.n1362 vdd.n1360 10.6151
R20043 vdd.n1363 vdd.n1362 10.6151
R20044 vdd.n1365 vdd.n1363 10.6151
R20045 vdd.n1366 vdd.n1365 10.6151
R20046 vdd.n1368 vdd.n1366 10.6151
R20047 vdd.n1369 vdd.n1368 10.6151
R20048 vdd.n1371 vdd.n1369 10.6151
R20049 vdd.n1372 vdd.n1371 10.6151
R20050 vdd.n1374 vdd.n1372 10.6151
R20051 vdd.n1375 vdd.n1374 10.6151
R20052 vdd.n1377 vdd.n1375 10.6151
R20053 vdd.n1378 vdd.n1377 10.6151
R20054 vdd.n1380 vdd.n1378 10.6151
R20055 vdd.n1381 vdd.n1380 10.6151
R20056 vdd.n1383 vdd.n1381 10.6151
R20057 vdd.n1384 vdd.n1383 10.6151
R20058 vdd.n1386 vdd.n1384 10.6151
R20059 vdd.n1387 vdd.n1386 10.6151
R20060 vdd.n1389 vdd.n1387 10.6151
R20061 vdd.n1390 vdd.n1389 10.6151
R20062 vdd.n1392 vdd.n1390 10.6151
R20063 vdd.n1393 vdd.n1392 10.6151
R20064 vdd.n1395 vdd.n1393 10.6151
R20065 vdd.n1396 vdd.n1395 10.6151
R20066 vdd.n1435 vdd.n1396 10.6151
R20067 vdd.n1435 vdd.n1434 10.6151
R20068 vdd.n1434 vdd.n1433 10.6151
R20069 vdd.n1433 vdd.n1431 10.6151
R20070 vdd.n1431 vdd.n1430 10.6151
R20071 vdd.n1430 vdd.n1428 10.6151
R20072 vdd.n1428 vdd.n1427 10.6151
R20073 vdd.n1427 vdd.n1408 10.6151
R20074 vdd.n1408 vdd.n1407 10.6151
R20075 vdd.n1407 vdd.n1405 10.6151
R20076 vdd.n1405 vdd.n1404 10.6151
R20077 vdd.n1404 vdd.n1402 10.6151
R20078 vdd.n1402 vdd.n1401 10.6151
R20079 vdd.n1401 vdd.n1398 10.6151
R20080 vdd.n1398 vdd.n1397 10.6151
R20081 vdd.n1397 vdd.n1003 10.6151
R20082 vdd.n2509 vdd.n1139 10.6151
R20083 vdd.n2504 vdd.n1139 10.6151
R20084 vdd.n2504 vdd.n2503 10.6151
R20085 vdd.n2503 vdd.n2502 10.6151
R20086 vdd.n2502 vdd.n2499 10.6151
R20087 vdd.n2499 vdd.n2498 10.6151
R20088 vdd.n2498 vdd.n2495 10.6151
R20089 vdd.n2495 vdd.n2494 10.6151
R20090 vdd.n2494 vdd.n2491 10.6151
R20091 vdd.n2491 vdd.n2490 10.6151
R20092 vdd.n2490 vdd.n2487 10.6151
R20093 vdd.n2487 vdd.n2486 10.6151
R20094 vdd.n2486 vdd.n2483 10.6151
R20095 vdd.n2483 vdd.n2482 10.6151
R20096 vdd.n2482 vdd.n2479 10.6151
R20097 vdd.n2479 vdd.n2478 10.6151
R20098 vdd.n2478 vdd.n2475 10.6151
R20099 vdd.n2475 vdd.n1177 10.6151
R20100 vdd.n1323 vdd.n1177 10.6151
R20101 vdd.n1324 vdd.n1323 10.6151
R20102 vdd.n1327 vdd.n1324 10.6151
R20103 vdd.n1328 vdd.n1327 10.6151
R20104 vdd.n1331 vdd.n1328 10.6151
R20105 vdd.n1332 vdd.n1331 10.6151
R20106 vdd.n1335 vdd.n1332 10.6151
R20107 vdd.n1336 vdd.n1335 10.6151
R20108 vdd.n1339 vdd.n1336 10.6151
R20109 vdd.n1340 vdd.n1339 10.6151
R20110 vdd.n1343 vdd.n1340 10.6151
R20111 vdd.n1344 vdd.n1343 10.6151
R20112 vdd.n1347 vdd.n1344 10.6151
R20113 vdd.n1352 vdd.n1349 10.6151
R20114 vdd.n1353 vdd.n1352 10.6151
R20115 vdd.n3020 vdd.n3019 10.6151
R20116 vdd.n3019 vdd.n3018 10.6151
R20117 vdd.n3018 vdd.n2822 10.6151
R20118 vdd.n2900 vdd.n2822 10.6151
R20119 vdd.n2901 vdd.n2900 10.6151
R20120 vdd.n2903 vdd.n2901 10.6151
R20121 vdd.n2904 vdd.n2903 10.6151
R20122 vdd.n3002 vdd.n2904 10.6151
R20123 vdd.n3002 vdd.n3001 10.6151
R20124 vdd.n3001 vdd.n3000 10.6151
R20125 vdd.n3000 vdd.n2948 10.6151
R20126 vdd.n2948 vdd.n2947 10.6151
R20127 vdd.n2947 vdd.n2945 10.6151
R20128 vdd.n2945 vdd.n2944 10.6151
R20129 vdd.n2944 vdd.n2942 10.6151
R20130 vdd.n2942 vdd.n2941 10.6151
R20131 vdd.n2941 vdd.n2939 10.6151
R20132 vdd.n2939 vdd.n2938 10.6151
R20133 vdd.n2938 vdd.n2936 10.6151
R20134 vdd.n2936 vdd.n2935 10.6151
R20135 vdd.n2935 vdd.n2933 10.6151
R20136 vdd.n2933 vdd.n2932 10.6151
R20137 vdd.n2932 vdd.n2930 10.6151
R20138 vdd.n2930 vdd.n2929 10.6151
R20139 vdd.n2929 vdd.n2927 10.6151
R20140 vdd.n2927 vdd.n2926 10.6151
R20141 vdd.n2926 vdd.n2924 10.6151
R20142 vdd.n2924 vdd.n2923 10.6151
R20143 vdd.n2923 vdd.n2921 10.6151
R20144 vdd.n2921 vdd.n2920 10.6151
R20145 vdd.n2920 vdd.n2918 10.6151
R20146 vdd.n2918 vdd.n2917 10.6151
R20147 vdd.n2917 vdd.n2915 10.6151
R20148 vdd.n2915 vdd.n2914 10.6151
R20149 vdd.n2914 vdd.n2912 10.6151
R20150 vdd.n2912 vdd.n2911 10.6151
R20151 vdd.n2911 vdd.n2909 10.6151
R20152 vdd.n2909 vdd.n2908 10.6151
R20153 vdd.n2908 vdd.n2906 10.6151
R20154 vdd.n2906 vdd.n2905 10.6151
R20155 vdd.n2905 vdd.n836 10.6151
R20156 vdd.n3264 vdd.n836 10.6151
R20157 vdd.n3265 vdd.n3264 10.6151
R20158 vdd.n3091 vdd.n961 10.6151
R20159 vdd.n3086 vdd.n961 10.6151
R20160 vdd.n3086 vdd.n3085 10.6151
R20161 vdd.n3085 vdd.n3084 10.6151
R20162 vdd.n3084 vdd.n3081 10.6151
R20163 vdd.n3081 vdd.n3080 10.6151
R20164 vdd.n3080 vdd.n3077 10.6151
R20165 vdd.n3077 vdd.n3076 10.6151
R20166 vdd.n3076 vdd.n3073 10.6151
R20167 vdd.n3073 vdd.n3072 10.6151
R20168 vdd.n3072 vdd.n3069 10.6151
R20169 vdd.n3069 vdd.n3068 10.6151
R20170 vdd.n3068 vdd.n3065 10.6151
R20171 vdd.n3065 vdd.n3064 10.6151
R20172 vdd.n3064 vdd.n3061 10.6151
R20173 vdd.n3061 vdd.n3060 10.6151
R20174 vdd.n3060 vdd.n3057 10.6151
R20175 vdd.n3057 vdd.n3056 10.6151
R20176 vdd.n3056 vdd.n3053 10.6151
R20177 vdd.n3053 vdd.n3052 10.6151
R20178 vdd.n3052 vdd.n3049 10.6151
R20179 vdd.n3049 vdd.n3048 10.6151
R20180 vdd.n3048 vdd.n3045 10.6151
R20181 vdd.n3045 vdd.n3044 10.6151
R20182 vdd.n3044 vdd.n3041 10.6151
R20183 vdd.n3041 vdd.n3040 10.6151
R20184 vdd.n3040 vdd.n3037 10.6151
R20185 vdd.n3037 vdd.n3036 10.6151
R20186 vdd.n3036 vdd.n3033 10.6151
R20187 vdd.n3033 vdd.n3032 10.6151
R20188 vdd.n3032 vdd.n3029 10.6151
R20189 vdd.n3027 vdd.n3024 10.6151
R20190 vdd.n3024 vdd.n3023 10.6151
R20191 vdd.n3093 vdd.n3092 10.6151
R20192 vdd.n3093 vdd.n950 10.6151
R20193 vdd.n3103 vdd.n950 10.6151
R20194 vdd.n3104 vdd.n3103 10.6151
R20195 vdd.n3105 vdd.n3104 10.6151
R20196 vdd.n3105 vdd.n938 10.6151
R20197 vdd.n3115 vdd.n938 10.6151
R20198 vdd.n3116 vdd.n3115 10.6151
R20199 vdd.n3117 vdd.n3116 10.6151
R20200 vdd.n3117 vdd.n927 10.6151
R20201 vdd.n3127 vdd.n927 10.6151
R20202 vdd.n3128 vdd.n3127 10.6151
R20203 vdd.n3129 vdd.n3128 10.6151
R20204 vdd.n3129 vdd.n916 10.6151
R20205 vdd.n3139 vdd.n916 10.6151
R20206 vdd.n3140 vdd.n3139 10.6151
R20207 vdd.n3141 vdd.n3140 10.6151
R20208 vdd.n3141 vdd.n903 10.6151
R20209 vdd.n3152 vdd.n903 10.6151
R20210 vdd.n3153 vdd.n3152 10.6151
R20211 vdd.n3154 vdd.n3153 10.6151
R20212 vdd.n3154 vdd.n891 10.6151
R20213 vdd.n3164 vdd.n891 10.6151
R20214 vdd.n3165 vdd.n3164 10.6151
R20215 vdd.n3166 vdd.n3165 10.6151
R20216 vdd.n3166 vdd.n879 10.6151
R20217 vdd.n3176 vdd.n879 10.6151
R20218 vdd.n3177 vdd.n3176 10.6151
R20219 vdd.n3178 vdd.n3177 10.6151
R20220 vdd.n3178 vdd.n866 10.6151
R20221 vdd.n3188 vdd.n866 10.6151
R20222 vdd.n3189 vdd.n3188 10.6151
R20223 vdd.n3190 vdd.n3189 10.6151
R20224 vdd.n3190 vdd.n855 10.6151
R20225 vdd.n3200 vdd.n855 10.6151
R20226 vdd.n3201 vdd.n3200 10.6151
R20227 vdd.n3202 vdd.n3201 10.6151
R20228 vdd.n3202 vdd.n841 10.6151
R20229 vdd.n3257 vdd.n841 10.6151
R20230 vdd.n3258 vdd.n3257 10.6151
R20231 vdd.n3259 vdd.n3258 10.6151
R20232 vdd.n3259 vdd.n810 10.6151
R20233 vdd.n3329 vdd.n810 10.6151
R20234 vdd.n3328 vdd.n3327 10.6151
R20235 vdd.n3327 vdd.n811 10.6151
R20236 vdd.n812 vdd.n811 10.6151
R20237 vdd.n3320 vdd.n812 10.6151
R20238 vdd.n3320 vdd.n3319 10.6151
R20239 vdd.n3319 vdd.n3318 10.6151
R20240 vdd.n3318 vdd.n814 10.6151
R20241 vdd.n3313 vdd.n814 10.6151
R20242 vdd.n3313 vdd.n3312 10.6151
R20243 vdd.n3312 vdd.n3311 10.6151
R20244 vdd.n3311 vdd.n817 10.6151
R20245 vdd.n3306 vdd.n817 10.6151
R20246 vdd.n3306 vdd.n3305 10.6151
R20247 vdd.n3305 vdd.n3304 10.6151
R20248 vdd.n3304 vdd.n820 10.6151
R20249 vdd.n3299 vdd.n820 10.6151
R20250 vdd.n3299 vdd.n731 10.6151
R20251 vdd.n3295 vdd.n731 10.6151
R20252 vdd.n3295 vdd.n3294 10.6151
R20253 vdd.n3294 vdd.n3293 10.6151
R20254 vdd.n3293 vdd.n823 10.6151
R20255 vdd.n3288 vdd.n823 10.6151
R20256 vdd.n3288 vdd.n3287 10.6151
R20257 vdd.n3287 vdd.n3286 10.6151
R20258 vdd.n3286 vdd.n826 10.6151
R20259 vdd.n3281 vdd.n826 10.6151
R20260 vdd.n3281 vdd.n3280 10.6151
R20261 vdd.n3280 vdd.n3279 10.6151
R20262 vdd.n3279 vdd.n829 10.6151
R20263 vdd.n3274 vdd.n829 10.6151
R20264 vdd.n3274 vdd.n3273 10.6151
R20265 vdd.n3271 vdd.n834 10.6151
R20266 vdd.n3266 vdd.n834 10.6151
R20267 vdd.n3247 vdd.n3208 10.6151
R20268 vdd.n3242 vdd.n3208 10.6151
R20269 vdd.n3242 vdd.n3241 10.6151
R20270 vdd.n3241 vdd.n3240 10.6151
R20271 vdd.n3240 vdd.n3210 10.6151
R20272 vdd.n3235 vdd.n3210 10.6151
R20273 vdd.n3235 vdd.n3234 10.6151
R20274 vdd.n3234 vdd.n3233 10.6151
R20275 vdd.n3233 vdd.n3213 10.6151
R20276 vdd.n3228 vdd.n3213 10.6151
R20277 vdd.n3228 vdd.n3227 10.6151
R20278 vdd.n3227 vdd.n3226 10.6151
R20279 vdd.n3226 vdd.n3216 10.6151
R20280 vdd.n3221 vdd.n3216 10.6151
R20281 vdd.n3221 vdd.n3220 10.6151
R20282 vdd.n3220 vdd.n785 10.6151
R20283 vdd.n3364 vdd.n785 10.6151
R20284 vdd.n3364 vdd.n786 10.6151
R20285 vdd.n788 vdd.n786 10.6151
R20286 vdd.n3357 vdd.n788 10.6151
R20287 vdd.n3357 vdd.n3356 10.6151
R20288 vdd.n3356 vdd.n3355 10.6151
R20289 vdd.n3355 vdd.n790 10.6151
R20290 vdd.n3350 vdd.n790 10.6151
R20291 vdd.n3350 vdd.n3349 10.6151
R20292 vdd.n3349 vdd.n3348 10.6151
R20293 vdd.n3348 vdd.n793 10.6151
R20294 vdd.n3343 vdd.n793 10.6151
R20295 vdd.n3343 vdd.n3342 10.6151
R20296 vdd.n3342 vdd.n3341 10.6151
R20297 vdd.n3341 vdd.n796 10.6151
R20298 vdd.n3336 vdd.n3335 10.6151
R20299 vdd.n3335 vdd.n3334 10.6151
R20300 vdd.n2897 vdd.n2896 10.6151
R20301 vdd.n3014 vdd.n2897 10.6151
R20302 vdd.n3014 vdd.n3013 10.6151
R20303 vdd.n3013 vdd.n3012 10.6151
R20304 vdd.n3012 vdd.n3010 10.6151
R20305 vdd.n3010 vdd.n3009 10.6151
R20306 vdd.n3009 vdd.n3007 10.6151
R20307 vdd.n3007 vdd.n3006 10.6151
R20308 vdd.n3006 vdd.n2898 10.6151
R20309 vdd.n2996 vdd.n2898 10.6151
R20310 vdd.n2996 vdd.n2995 10.6151
R20311 vdd.n2995 vdd.n2994 10.6151
R20312 vdd.n2994 vdd.n2992 10.6151
R20313 vdd.n2992 vdd.n2991 10.6151
R20314 vdd.n2991 vdd.n2989 10.6151
R20315 vdd.n2989 vdd.n2988 10.6151
R20316 vdd.n2988 vdd.n2986 10.6151
R20317 vdd.n2986 vdd.n2985 10.6151
R20318 vdd.n2985 vdd.n2983 10.6151
R20319 vdd.n2983 vdd.n2982 10.6151
R20320 vdd.n2982 vdd.n2980 10.6151
R20321 vdd.n2980 vdd.n2979 10.6151
R20322 vdd.n2979 vdd.n2977 10.6151
R20323 vdd.n2977 vdd.n2976 10.6151
R20324 vdd.n2976 vdd.n2974 10.6151
R20325 vdd.n2974 vdd.n2973 10.6151
R20326 vdd.n2973 vdd.n2971 10.6151
R20327 vdd.n2971 vdd.n2970 10.6151
R20328 vdd.n2970 vdd.n2968 10.6151
R20329 vdd.n2968 vdd.n2967 10.6151
R20330 vdd.n2967 vdd.n2965 10.6151
R20331 vdd.n2965 vdd.n2964 10.6151
R20332 vdd.n2964 vdd.n2962 10.6151
R20333 vdd.n2962 vdd.n2961 10.6151
R20334 vdd.n2961 vdd.n2959 10.6151
R20335 vdd.n2959 vdd.n2958 10.6151
R20336 vdd.n2958 vdd.n2956 10.6151
R20337 vdd.n2956 vdd.n2955 10.6151
R20338 vdd.n2955 vdd.n2953 10.6151
R20339 vdd.n2953 vdd.n2952 10.6151
R20340 vdd.n2952 vdd.n2950 10.6151
R20341 vdd.n2950 vdd.n2949 10.6151
R20342 vdd.n2949 vdd.n802 10.6151
R20343 vdd.n2828 vdd.n2827 10.6151
R20344 vdd.n2831 vdd.n2828 10.6151
R20345 vdd.n2832 vdd.n2831 10.6151
R20346 vdd.n2835 vdd.n2832 10.6151
R20347 vdd.n2836 vdd.n2835 10.6151
R20348 vdd.n2839 vdd.n2836 10.6151
R20349 vdd.n2840 vdd.n2839 10.6151
R20350 vdd.n2843 vdd.n2840 10.6151
R20351 vdd.n2844 vdd.n2843 10.6151
R20352 vdd.n2847 vdd.n2844 10.6151
R20353 vdd.n2848 vdd.n2847 10.6151
R20354 vdd.n2851 vdd.n2848 10.6151
R20355 vdd.n2852 vdd.n2851 10.6151
R20356 vdd.n2855 vdd.n2852 10.6151
R20357 vdd.n2856 vdd.n2855 10.6151
R20358 vdd.n2859 vdd.n2856 10.6151
R20359 vdd.n2860 vdd.n2859 10.6151
R20360 vdd.n2863 vdd.n2860 10.6151
R20361 vdd.n2864 vdd.n2863 10.6151
R20362 vdd.n2867 vdd.n2864 10.6151
R20363 vdd.n2868 vdd.n2867 10.6151
R20364 vdd.n2871 vdd.n2868 10.6151
R20365 vdd.n2872 vdd.n2871 10.6151
R20366 vdd.n2875 vdd.n2872 10.6151
R20367 vdd.n2876 vdd.n2875 10.6151
R20368 vdd.n2879 vdd.n2876 10.6151
R20369 vdd.n2880 vdd.n2879 10.6151
R20370 vdd.n2883 vdd.n2880 10.6151
R20371 vdd.n2884 vdd.n2883 10.6151
R20372 vdd.n2887 vdd.n2884 10.6151
R20373 vdd.n2888 vdd.n2887 10.6151
R20374 vdd.n2893 vdd.n2891 10.6151
R20375 vdd.n2894 vdd.n2893 10.6151
R20376 vdd.n3097 vdd.n955 10.6151
R20377 vdd.n3098 vdd.n3097 10.6151
R20378 vdd.n3099 vdd.n3098 10.6151
R20379 vdd.n3099 vdd.n944 10.6151
R20380 vdd.n3109 vdd.n944 10.6151
R20381 vdd.n3110 vdd.n3109 10.6151
R20382 vdd.n3111 vdd.n3110 10.6151
R20383 vdd.n3111 vdd.n933 10.6151
R20384 vdd.n3121 vdd.n933 10.6151
R20385 vdd.n3122 vdd.n3121 10.6151
R20386 vdd.n3123 vdd.n3122 10.6151
R20387 vdd.n3123 vdd.n921 10.6151
R20388 vdd.n3133 vdd.n921 10.6151
R20389 vdd.n3134 vdd.n3133 10.6151
R20390 vdd.n3135 vdd.n3134 10.6151
R20391 vdd.n3135 vdd.n910 10.6151
R20392 vdd.n3145 vdd.n910 10.6151
R20393 vdd.n3146 vdd.n3145 10.6151
R20394 vdd.n3148 vdd.n3146 10.6151
R20395 vdd.n3148 vdd.n3147 10.6151
R20396 vdd.n3159 vdd.n3158 10.6151
R20397 vdd.n3160 vdd.n3159 10.6151
R20398 vdd.n3160 vdd.n885 10.6151
R20399 vdd.n3170 vdd.n885 10.6151
R20400 vdd.n3171 vdd.n3170 10.6151
R20401 vdd.n3172 vdd.n3171 10.6151
R20402 vdd.n3172 vdd.n872 10.6151
R20403 vdd.n3182 vdd.n872 10.6151
R20404 vdd.n3183 vdd.n3182 10.6151
R20405 vdd.n3184 vdd.n3183 10.6151
R20406 vdd.n3184 vdd.n860 10.6151
R20407 vdd.n3194 vdd.n860 10.6151
R20408 vdd.n3195 vdd.n3194 10.6151
R20409 vdd.n3196 vdd.n3195 10.6151
R20410 vdd.n3196 vdd.n849 10.6151
R20411 vdd.n3206 vdd.n849 10.6151
R20412 vdd.n3207 vdd.n3206 10.6151
R20413 vdd.n3253 vdd.n3207 10.6151
R20414 vdd.n3253 vdd.n3252 10.6151
R20415 vdd.n3252 vdd.n3251 10.6151
R20416 vdd.n3251 vdd.n3250 10.6151
R20417 vdd.n3250 vdd.n3248 10.6151
R20418 vdd.n2515 vdd.n1132 10.6151
R20419 vdd.n2516 vdd.n2515 10.6151
R20420 vdd.n2517 vdd.n2516 10.6151
R20421 vdd.n2517 vdd.n1121 10.6151
R20422 vdd.n2527 vdd.n1121 10.6151
R20423 vdd.n2528 vdd.n2527 10.6151
R20424 vdd.n2529 vdd.n2528 10.6151
R20425 vdd.n2529 vdd.n1108 10.6151
R20426 vdd.n2539 vdd.n1108 10.6151
R20427 vdd.n2540 vdd.n2539 10.6151
R20428 vdd.n2541 vdd.n2540 10.6151
R20429 vdd.n2541 vdd.n1097 10.6151
R20430 vdd.n2551 vdd.n1097 10.6151
R20431 vdd.n2552 vdd.n2551 10.6151
R20432 vdd.n2553 vdd.n2552 10.6151
R20433 vdd.n2553 vdd.n1085 10.6151
R20434 vdd.n2563 vdd.n1085 10.6151
R20435 vdd.n2564 vdd.n2563 10.6151
R20436 vdd.n2565 vdd.n2564 10.6151
R20437 vdd.n2565 vdd.n1072 10.6151
R20438 vdd.n2575 vdd.n1072 10.6151
R20439 vdd.n2576 vdd.n2575 10.6151
R20440 vdd.n2578 vdd.n1060 10.6151
R20441 vdd.n2588 vdd.n1060 10.6151
R20442 vdd.n2589 vdd.n2588 10.6151
R20443 vdd.n2590 vdd.n2589 10.6151
R20444 vdd.n2590 vdd.n1048 10.6151
R20445 vdd.n2600 vdd.n1048 10.6151
R20446 vdd.n2601 vdd.n2600 10.6151
R20447 vdd.n2602 vdd.n2601 10.6151
R20448 vdd.n2602 vdd.n1037 10.6151
R20449 vdd.n2612 vdd.n1037 10.6151
R20450 vdd.n2613 vdd.n2612 10.6151
R20451 vdd.n2614 vdd.n2613 10.6151
R20452 vdd.n2614 vdd.n1026 10.6151
R20453 vdd.n2624 vdd.n1026 10.6151
R20454 vdd.n2625 vdd.n2624 10.6151
R20455 vdd.n2628 vdd.n2625 10.6151
R20456 vdd.n2628 vdd.n2627 10.6151
R20457 vdd.n2627 vdd.n2626 10.6151
R20458 vdd.n2626 vdd.n1009 10.6151
R20459 vdd.n2710 vdd.n1009 10.6151
R20460 vdd.n2709 vdd.n2708 10.6151
R20461 vdd.n2708 vdd.n2705 10.6151
R20462 vdd.n2705 vdd.n2704 10.6151
R20463 vdd.n2704 vdd.n2701 10.6151
R20464 vdd.n2701 vdd.n2700 10.6151
R20465 vdd.n2700 vdd.n2697 10.6151
R20466 vdd.n2697 vdd.n2696 10.6151
R20467 vdd.n2696 vdd.n2693 10.6151
R20468 vdd.n2693 vdd.n2692 10.6151
R20469 vdd.n2692 vdd.n2689 10.6151
R20470 vdd.n2689 vdd.n2688 10.6151
R20471 vdd.n2688 vdd.n2685 10.6151
R20472 vdd.n2685 vdd.n2684 10.6151
R20473 vdd.n2684 vdd.n2681 10.6151
R20474 vdd.n2681 vdd.n2680 10.6151
R20475 vdd.n2680 vdd.n2677 10.6151
R20476 vdd.n2677 vdd.n2676 10.6151
R20477 vdd.n2676 vdd.n2673 10.6151
R20478 vdd.n2673 vdd.n2672 10.6151
R20479 vdd.n2672 vdd.n2669 10.6151
R20480 vdd.n2669 vdd.n2668 10.6151
R20481 vdd.n2668 vdd.n2665 10.6151
R20482 vdd.n2665 vdd.n2664 10.6151
R20483 vdd.n2664 vdd.n2661 10.6151
R20484 vdd.n2661 vdd.n2660 10.6151
R20485 vdd.n2660 vdd.n2657 10.6151
R20486 vdd.n2657 vdd.n2656 10.6151
R20487 vdd.n2656 vdd.n2653 10.6151
R20488 vdd.n2653 vdd.n2652 10.6151
R20489 vdd.n2652 vdd.n2649 10.6151
R20490 vdd.n2649 vdd.n2648 10.6151
R20491 vdd.n2645 vdd.n2644 10.6151
R20492 vdd.n2644 vdd.n2642 10.6151
R20493 vdd.n1481 vdd.n1479 10.6151
R20494 vdd.n1479 vdd.n1478 10.6151
R20495 vdd.n1478 vdd.n1476 10.6151
R20496 vdd.n1476 vdd.n1475 10.6151
R20497 vdd.n1475 vdd.n1473 10.6151
R20498 vdd.n1473 vdd.n1472 10.6151
R20499 vdd.n1472 vdd.n1470 10.6151
R20500 vdd.n1470 vdd.n1469 10.6151
R20501 vdd.n1469 vdd.n1467 10.6151
R20502 vdd.n1467 vdd.n1466 10.6151
R20503 vdd.n1466 vdd.n1464 10.6151
R20504 vdd.n1464 vdd.n1463 10.6151
R20505 vdd.n1463 vdd.n1461 10.6151
R20506 vdd.n1461 vdd.n1460 10.6151
R20507 vdd.n1460 vdd.n1458 10.6151
R20508 vdd.n1458 vdd.n1457 10.6151
R20509 vdd.n1457 vdd.n1455 10.6151
R20510 vdd.n1455 vdd.n1454 10.6151
R20511 vdd.n1454 vdd.n1452 10.6151
R20512 vdd.n1452 vdd.n1451 10.6151
R20513 vdd.n1451 vdd.n1449 10.6151
R20514 vdd.n1449 vdd.n1448 10.6151
R20515 vdd.n1448 vdd.n1446 10.6151
R20516 vdd.n1446 vdd.n1445 10.6151
R20517 vdd.n1445 vdd.n1443 10.6151
R20518 vdd.n1443 vdd.n1442 10.6151
R20519 vdd.n1442 vdd.n1440 10.6151
R20520 vdd.n1440 vdd.n1439 10.6151
R20521 vdd.n1439 vdd.n1318 10.6151
R20522 vdd.n1410 vdd.n1318 10.6151
R20523 vdd.n1411 vdd.n1410 10.6151
R20524 vdd.n1413 vdd.n1411 10.6151
R20525 vdd.n1414 vdd.n1413 10.6151
R20526 vdd.n1423 vdd.n1414 10.6151
R20527 vdd.n1423 vdd.n1422 10.6151
R20528 vdd.n1422 vdd.n1421 10.6151
R20529 vdd.n1421 vdd.n1419 10.6151
R20530 vdd.n1419 vdd.n1418 10.6151
R20531 vdd.n1418 vdd.n1416 10.6151
R20532 vdd.n1416 vdd.n1415 10.6151
R20533 vdd.n1415 vdd.n1013 10.6151
R20534 vdd.n2640 vdd.n1013 10.6151
R20535 vdd.n2641 vdd.n2640 10.6151
R20536 vdd.n1282 vdd.n1281 10.6151
R20537 vdd.n1285 vdd.n1282 10.6151
R20538 vdd.n1286 vdd.n1285 10.6151
R20539 vdd.n1289 vdd.n1286 10.6151
R20540 vdd.n1290 vdd.n1289 10.6151
R20541 vdd.n1293 vdd.n1290 10.6151
R20542 vdd.n1294 vdd.n1293 10.6151
R20543 vdd.n1297 vdd.n1294 10.6151
R20544 vdd.n1298 vdd.n1297 10.6151
R20545 vdd.n1301 vdd.n1298 10.6151
R20546 vdd.n1302 vdd.n1301 10.6151
R20547 vdd.n1305 vdd.n1302 10.6151
R20548 vdd.n1306 vdd.n1305 10.6151
R20549 vdd.n1309 vdd.n1306 10.6151
R20550 vdd.n1310 vdd.n1309 10.6151
R20551 vdd.n1313 vdd.n1310 10.6151
R20552 vdd.n1515 vdd.n1313 10.6151
R20553 vdd.n1515 vdd.n1514 10.6151
R20554 vdd.n1514 vdd.n1512 10.6151
R20555 vdd.n1512 vdd.n1509 10.6151
R20556 vdd.n1509 vdd.n1508 10.6151
R20557 vdd.n1508 vdd.n1505 10.6151
R20558 vdd.n1505 vdd.n1504 10.6151
R20559 vdd.n1504 vdd.n1501 10.6151
R20560 vdd.n1501 vdd.n1500 10.6151
R20561 vdd.n1500 vdd.n1497 10.6151
R20562 vdd.n1497 vdd.n1496 10.6151
R20563 vdd.n1496 vdd.n1493 10.6151
R20564 vdd.n1493 vdd.n1492 10.6151
R20565 vdd.n1492 vdd.n1489 10.6151
R20566 vdd.n1489 vdd.n1488 10.6151
R20567 vdd.n1485 vdd.n1484 10.6151
R20568 vdd.n1484 vdd.n1482 10.6151
R20569 vdd.n2306 vdd.t127 10.5435
R20570 vdd.n656 vdd.t102 10.5435
R20571 vdd.n316 vdd.n298 10.4732
R20572 vdd.n257 vdd.n239 10.4732
R20573 vdd.n214 vdd.n196 10.4732
R20574 vdd.n155 vdd.n137 10.4732
R20575 vdd.n113 vdd.n95 10.4732
R20576 vdd.n54 vdd.n36 10.4732
R20577 vdd.n2190 vdd.n2172 10.4732
R20578 vdd.n2249 vdd.n2231 10.4732
R20579 vdd.n2088 vdd.n2070 10.4732
R20580 vdd.n2147 vdd.n2129 10.4732
R20581 vdd.n1987 vdd.n1969 10.4732
R20582 vdd.n2046 vdd.n2028 10.4732
R20583 vdd.t148 vdd.n2280 10.3167
R20584 vdd.n3572 vdd.t94 10.3167
R20585 vdd.n1957 vdd.t136 10.09
R20586 vdd.n3666 vdd.t106 10.09
R20587 vdd.n2475 vdd.n2474 9.98956
R20588 vdd.n3488 vdd.n731 9.98956
R20589 vdd.n3365 vdd.n3364 9.98956
R20590 vdd.n2367 vdd.n1515 9.98956
R20591 vdd.t132 vdd.n1610 9.86327
R20592 vdd.n3657 vdd.t227 9.86327
R20593 vdd.n2712 vdd.t296 9.7499
R20594 vdd.t270 vdd.n957 9.7499
R20595 vdd.n315 vdd.n300 9.69747
R20596 vdd.n256 vdd.n241 9.69747
R20597 vdd.n213 vdd.n198 9.69747
R20598 vdd.n154 vdd.n139 9.69747
R20599 vdd.n112 vdd.n97 9.69747
R20600 vdd.n53 vdd.n38 9.69747
R20601 vdd.n2189 vdd.n2174 9.69747
R20602 vdd.n2248 vdd.n2233 9.69747
R20603 vdd.n2087 vdd.n2072 9.69747
R20604 vdd.n2146 vdd.n2131 9.69747
R20605 vdd.n1986 vdd.n1971 9.69747
R20606 vdd.n2045 vdd.n2030 9.69747
R20607 vdd.n1916 vdd.t120 9.63654
R20608 vdd.n3603 vdd.t154 9.63654
R20609 vdd.n331 vdd.n330 9.45567
R20610 vdd.n272 vdd.n271 9.45567
R20611 vdd.n229 vdd.n228 9.45567
R20612 vdd.n170 vdd.n169 9.45567
R20613 vdd.n128 vdd.n127 9.45567
R20614 vdd.n69 vdd.n68 9.45567
R20615 vdd.n2205 vdd.n2204 9.45567
R20616 vdd.n2264 vdd.n2263 9.45567
R20617 vdd.n2103 vdd.n2102 9.45567
R20618 vdd.n2162 vdd.n2161 9.45567
R20619 vdd.n2002 vdd.n2001 9.45567
R20620 vdd.n2061 vdd.n2060 9.45567
R20621 vdd.n1890 vdd.t175 9.40981
R20622 vdd.n3635 vdd.t104 9.40981
R20623 vdd.n2437 vdd.n1207 9.3005
R20624 vdd.n2436 vdd.n2435 9.3005
R20625 vdd.n1213 vdd.n1212 9.3005
R20626 vdd.n2430 vdd.n1217 9.3005
R20627 vdd.n2429 vdd.n1218 9.3005
R20628 vdd.n2428 vdd.n1219 9.3005
R20629 vdd.n1223 vdd.n1220 9.3005
R20630 vdd.n2423 vdd.n1224 9.3005
R20631 vdd.n2422 vdd.n1225 9.3005
R20632 vdd.n2421 vdd.n1226 9.3005
R20633 vdd.n1230 vdd.n1227 9.3005
R20634 vdd.n2416 vdd.n1231 9.3005
R20635 vdd.n2415 vdd.n1232 9.3005
R20636 vdd.n2414 vdd.n1233 9.3005
R20637 vdd.n1237 vdd.n1234 9.3005
R20638 vdd.n2409 vdd.n1238 9.3005
R20639 vdd.n2408 vdd.n1239 9.3005
R20640 vdd.n2407 vdd.n1240 9.3005
R20641 vdd.n1244 vdd.n1241 9.3005
R20642 vdd.n2402 vdd.n1245 9.3005
R20643 vdd.n2401 vdd.n1246 9.3005
R20644 vdd.n2400 vdd.n2399 9.3005
R20645 vdd.n2398 vdd.n1247 9.3005
R20646 vdd.n2397 vdd.n2396 9.3005
R20647 vdd.n1253 vdd.n1252 9.3005
R20648 vdd.n2391 vdd.n1257 9.3005
R20649 vdd.n2390 vdd.n1258 9.3005
R20650 vdd.n2389 vdd.n1259 9.3005
R20651 vdd.n1263 vdd.n1260 9.3005
R20652 vdd.n2384 vdd.n1264 9.3005
R20653 vdd.n2383 vdd.n1265 9.3005
R20654 vdd.n2382 vdd.n1266 9.3005
R20655 vdd.n1270 vdd.n1267 9.3005
R20656 vdd.n2377 vdd.n1271 9.3005
R20657 vdd.n2376 vdd.n1272 9.3005
R20658 vdd.n2375 vdd.n1273 9.3005
R20659 vdd.n1277 vdd.n1274 9.3005
R20660 vdd.n2370 vdd.n1278 9.3005
R20661 vdd.n2439 vdd.n2438 9.3005
R20662 vdd.n2461 vdd.n1178 9.3005
R20663 vdd.n2460 vdd.n1186 9.3005
R20664 vdd.n1190 vdd.n1187 9.3005
R20665 vdd.n2455 vdd.n1191 9.3005
R20666 vdd.n2454 vdd.n1192 9.3005
R20667 vdd.n2453 vdd.n1193 9.3005
R20668 vdd.n1197 vdd.n1194 9.3005
R20669 vdd.n2448 vdd.n1198 9.3005
R20670 vdd.n2447 vdd.n1199 9.3005
R20671 vdd.n2446 vdd.n1200 9.3005
R20672 vdd.n1204 vdd.n1201 9.3005
R20673 vdd.n2441 vdd.n1205 9.3005
R20674 vdd.n2440 vdd.n1206 9.3005
R20675 vdd.n2473 vdd.n2472 9.3005
R20676 vdd.n1182 vdd.n1181 9.3005
R20677 vdd.n2270 vdd.n2269 9.3005
R20678 vdd.n1579 vdd.n1578 9.3005
R20679 vdd.n2284 vdd.n2283 9.3005
R20680 vdd.n2285 vdd.n1577 9.3005
R20681 vdd.n2287 vdd.n2286 9.3005
R20682 vdd.n1568 vdd.n1567 9.3005
R20683 vdd.n2301 vdd.n2300 9.3005
R20684 vdd.n2302 vdd.n1566 9.3005
R20685 vdd.n2304 vdd.n2303 9.3005
R20686 vdd.n1557 vdd.n1556 9.3005
R20687 vdd.n2317 vdd.n2316 9.3005
R20688 vdd.n2318 vdd.n1555 9.3005
R20689 vdd.n2320 vdd.n2319 9.3005
R20690 vdd.n1545 vdd.n1544 9.3005
R20691 vdd.n2334 vdd.n2333 9.3005
R20692 vdd.n2335 vdd.n1543 9.3005
R20693 vdd.n2337 vdd.n2336 9.3005
R20694 vdd.n1533 vdd.n1532 9.3005
R20695 vdd.n2353 vdd.n2352 9.3005
R20696 vdd.n2354 vdd.n1531 9.3005
R20697 vdd.n2356 vdd.n2355 9.3005
R20698 vdd.n307 vdd.n306 9.3005
R20699 vdd.n302 vdd.n301 9.3005
R20700 vdd.n313 vdd.n312 9.3005
R20701 vdd.n315 vdd.n314 9.3005
R20702 vdd.n298 vdd.n297 9.3005
R20703 vdd.n321 vdd.n320 9.3005
R20704 vdd.n323 vdd.n322 9.3005
R20705 vdd.n295 vdd.n292 9.3005
R20706 vdd.n330 vdd.n329 9.3005
R20707 vdd.n248 vdd.n247 9.3005
R20708 vdd.n243 vdd.n242 9.3005
R20709 vdd.n254 vdd.n253 9.3005
R20710 vdd.n256 vdd.n255 9.3005
R20711 vdd.n239 vdd.n238 9.3005
R20712 vdd.n262 vdd.n261 9.3005
R20713 vdd.n264 vdd.n263 9.3005
R20714 vdd.n236 vdd.n233 9.3005
R20715 vdd.n271 vdd.n270 9.3005
R20716 vdd.n205 vdd.n204 9.3005
R20717 vdd.n200 vdd.n199 9.3005
R20718 vdd.n211 vdd.n210 9.3005
R20719 vdd.n213 vdd.n212 9.3005
R20720 vdd.n196 vdd.n195 9.3005
R20721 vdd.n219 vdd.n218 9.3005
R20722 vdd.n221 vdd.n220 9.3005
R20723 vdd.n193 vdd.n190 9.3005
R20724 vdd.n228 vdd.n227 9.3005
R20725 vdd.n146 vdd.n145 9.3005
R20726 vdd.n141 vdd.n140 9.3005
R20727 vdd.n152 vdd.n151 9.3005
R20728 vdd.n154 vdd.n153 9.3005
R20729 vdd.n137 vdd.n136 9.3005
R20730 vdd.n160 vdd.n159 9.3005
R20731 vdd.n162 vdd.n161 9.3005
R20732 vdd.n134 vdd.n131 9.3005
R20733 vdd.n169 vdd.n168 9.3005
R20734 vdd.n104 vdd.n103 9.3005
R20735 vdd.n99 vdd.n98 9.3005
R20736 vdd.n110 vdd.n109 9.3005
R20737 vdd.n112 vdd.n111 9.3005
R20738 vdd.n95 vdd.n94 9.3005
R20739 vdd.n118 vdd.n117 9.3005
R20740 vdd.n120 vdd.n119 9.3005
R20741 vdd.n92 vdd.n89 9.3005
R20742 vdd.n127 vdd.n126 9.3005
R20743 vdd.n45 vdd.n44 9.3005
R20744 vdd.n40 vdd.n39 9.3005
R20745 vdd.n51 vdd.n50 9.3005
R20746 vdd.n53 vdd.n52 9.3005
R20747 vdd.n36 vdd.n35 9.3005
R20748 vdd.n59 vdd.n58 9.3005
R20749 vdd.n61 vdd.n60 9.3005
R20750 vdd.n33 vdd.n30 9.3005
R20751 vdd.n68 vdd.n67 9.3005
R20752 vdd.n3410 vdd.n3409 9.3005
R20753 vdd.n3413 vdd.n766 9.3005
R20754 vdd.n3414 vdd.n765 9.3005
R20755 vdd.n3417 vdd.n764 9.3005
R20756 vdd.n3418 vdd.n763 9.3005
R20757 vdd.n3421 vdd.n762 9.3005
R20758 vdd.n3422 vdd.n761 9.3005
R20759 vdd.n3425 vdd.n760 9.3005
R20760 vdd.n3426 vdd.n759 9.3005
R20761 vdd.n3429 vdd.n758 9.3005
R20762 vdd.n3430 vdd.n757 9.3005
R20763 vdd.n3433 vdd.n756 9.3005
R20764 vdd.n3434 vdd.n755 9.3005
R20765 vdd.n3437 vdd.n754 9.3005
R20766 vdd.n3438 vdd.n753 9.3005
R20767 vdd.n3441 vdd.n752 9.3005
R20768 vdd.n3442 vdd.n751 9.3005
R20769 vdd.n3445 vdd.n750 9.3005
R20770 vdd.n3446 vdd.n749 9.3005
R20771 vdd.n3449 vdd.n748 9.3005
R20772 vdd.n3453 vdd.n3452 9.3005
R20773 vdd.n3454 vdd.n747 9.3005
R20774 vdd.n3458 vdd.n3455 9.3005
R20775 vdd.n3461 vdd.n746 9.3005
R20776 vdd.n3462 vdd.n745 9.3005
R20777 vdd.n3465 vdd.n744 9.3005
R20778 vdd.n3466 vdd.n743 9.3005
R20779 vdd.n3469 vdd.n742 9.3005
R20780 vdd.n3470 vdd.n741 9.3005
R20781 vdd.n3473 vdd.n740 9.3005
R20782 vdd.n3474 vdd.n739 9.3005
R20783 vdd.n3477 vdd.n738 9.3005
R20784 vdd.n3478 vdd.n737 9.3005
R20785 vdd.n3481 vdd.n736 9.3005
R20786 vdd.n3482 vdd.n735 9.3005
R20787 vdd.n3485 vdd.n730 9.3005
R20788 vdd.n3491 vdd.n727 9.3005
R20789 vdd.n3492 vdd.n726 9.3005
R20790 vdd.n3506 vdd.n3505 9.3005
R20791 vdd.n3507 vdd.n681 9.3005
R20792 vdd.n3509 vdd.n3508 9.3005
R20793 vdd.n671 vdd.n670 9.3005
R20794 vdd.n3523 vdd.n3522 9.3005
R20795 vdd.n3524 vdd.n669 9.3005
R20796 vdd.n3526 vdd.n3525 9.3005
R20797 vdd.n660 vdd.n659 9.3005
R20798 vdd.n3539 vdd.n3538 9.3005
R20799 vdd.n3540 vdd.n658 9.3005
R20800 vdd.n3542 vdd.n3541 9.3005
R20801 vdd.n648 vdd.n647 9.3005
R20802 vdd.n3556 vdd.n3555 9.3005
R20803 vdd.n3557 vdd.n646 9.3005
R20804 vdd.n3559 vdd.n3558 9.3005
R20805 vdd.n637 vdd.n636 9.3005
R20806 vdd.n3575 vdd.n3574 9.3005
R20807 vdd.n3576 vdd.n635 9.3005
R20808 vdd.n3578 vdd.n3577 9.3005
R20809 vdd.n336 vdd.n334 9.3005
R20810 vdd.n683 vdd.n682 9.3005
R20811 vdd.n3670 vdd.n3669 9.3005
R20812 vdd.n337 vdd.n335 9.3005
R20813 vdd.n3663 vdd.n346 9.3005
R20814 vdd.n3662 vdd.n347 9.3005
R20815 vdd.n3661 vdd.n348 9.3005
R20816 vdd.n355 vdd.n349 9.3005
R20817 vdd.n3655 vdd.n356 9.3005
R20818 vdd.n3654 vdd.n357 9.3005
R20819 vdd.n3653 vdd.n358 9.3005
R20820 vdd.n366 vdd.n359 9.3005
R20821 vdd.n3647 vdd.n367 9.3005
R20822 vdd.n3646 vdd.n368 9.3005
R20823 vdd.n3645 vdd.n369 9.3005
R20824 vdd.n377 vdd.n370 9.3005
R20825 vdd.n3639 vdd.n378 9.3005
R20826 vdd.n3638 vdd.n379 9.3005
R20827 vdd.n3637 vdd.n380 9.3005
R20828 vdd.n388 vdd.n381 9.3005
R20829 vdd.n3631 vdd.n389 9.3005
R20830 vdd.n3630 vdd.n390 9.3005
R20831 vdd.n3629 vdd.n391 9.3005
R20832 vdd.n466 vdd.n463 9.3005
R20833 vdd.n470 vdd.n469 9.3005
R20834 vdd.n471 vdd.n462 9.3005
R20835 vdd.n475 vdd.n472 9.3005
R20836 vdd.n476 vdd.n461 9.3005
R20837 vdd.n480 vdd.n479 9.3005
R20838 vdd.n481 vdd.n460 9.3005
R20839 vdd.n485 vdd.n482 9.3005
R20840 vdd.n486 vdd.n459 9.3005
R20841 vdd.n490 vdd.n489 9.3005
R20842 vdd.n491 vdd.n458 9.3005
R20843 vdd.n495 vdd.n492 9.3005
R20844 vdd.n496 vdd.n457 9.3005
R20845 vdd.n500 vdd.n499 9.3005
R20846 vdd.n501 vdd.n456 9.3005
R20847 vdd.n505 vdd.n502 9.3005
R20848 vdd.n506 vdd.n455 9.3005
R20849 vdd.n510 vdd.n509 9.3005
R20850 vdd.n511 vdd.n454 9.3005
R20851 vdd.n515 vdd.n512 9.3005
R20852 vdd.n516 vdd.n451 9.3005
R20853 vdd.n520 vdd.n519 9.3005
R20854 vdd.n521 vdd.n450 9.3005
R20855 vdd.n525 vdd.n522 9.3005
R20856 vdd.n526 vdd.n449 9.3005
R20857 vdd.n530 vdd.n529 9.3005
R20858 vdd.n531 vdd.n448 9.3005
R20859 vdd.n535 vdd.n532 9.3005
R20860 vdd.n536 vdd.n447 9.3005
R20861 vdd.n540 vdd.n539 9.3005
R20862 vdd.n541 vdd.n446 9.3005
R20863 vdd.n545 vdd.n542 9.3005
R20864 vdd.n546 vdd.n445 9.3005
R20865 vdd.n550 vdd.n549 9.3005
R20866 vdd.n551 vdd.n444 9.3005
R20867 vdd.n555 vdd.n552 9.3005
R20868 vdd.n556 vdd.n443 9.3005
R20869 vdd.n560 vdd.n559 9.3005
R20870 vdd.n561 vdd.n442 9.3005
R20871 vdd.n565 vdd.n562 9.3005
R20872 vdd.n566 vdd.n439 9.3005
R20873 vdd.n570 vdd.n569 9.3005
R20874 vdd.n571 vdd.n438 9.3005
R20875 vdd.n575 vdd.n572 9.3005
R20876 vdd.n576 vdd.n437 9.3005
R20877 vdd.n580 vdd.n579 9.3005
R20878 vdd.n581 vdd.n436 9.3005
R20879 vdd.n585 vdd.n582 9.3005
R20880 vdd.n586 vdd.n435 9.3005
R20881 vdd.n590 vdd.n589 9.3005
R20882 vdd.n591 vdd.n434 9.3005
R20883 vdd.n595 vdd.n592 9.3005
R20884 vdd.n596 vdd.n433 9.3005
R20885 vdd.n600 vdd.n599 9.3005
R20886 vdd.n601 vdd.n432 9.3005
R20887 vdd.n605 vdd.n602 9.3005
R20888 vdd.n606 vdd.n431 9.3005
R20889 vdd.n610 vdd.n609 9.3005
R20890 vdd.n611 vdd.n430 9.3005
R20891 vdd.n615 vdd.n612 9.3005
R20892 vdd.n617 vdd.n429 9.3005
R20893 vdd.n619 vdd.n618 9.3005
R20894 vdd.n3623 vdd.n3622 9.3005
R20895 vdd.n465 vdd.n464 9.3005
R20896 vdd.n3501 vdd.n3500 9.3005
R20897 vdd.n676 vdd.n675 9.3005
R20898 vdd.n3514 vdd.n3513 9.3005
R20899 vdd.n3515 vdd.n674 9.3005
R20900 vdd.n3517 vdd.n3516 9.3005
R20901 vdd.n666 vdd.n665 9.3005
R20902 vdd.n3531 vdd.n3530 9.3005
R20903 vdd.n3532 vdd.n664 9.3005
R20904 vdd.n3534 vdd.n3533 9.3005
R20905 vdd.n653 vdd.n652 9.3005
R20906 vdd.n3547 vdd.n3546 9.3005
R20907 vdd.n3548 vdd.n651 9.3005
R20908 vdd.n3550 vdd.n3549 9.3005
R20909 vdd.n642 vdd.n641 9.3005
R20910 vdd.n3564 vdd.n3563 9.3005
R20911 vdd.n3565 vdd.n640 9.3005
R20912 vdd.n3570 vdd.n3566 9.3005
R20913 vdd.n3569 vdd.n3568 9.3005
R20914 vdd.n3567 vdd.n631 9.3005
R20915 vdd.n3583 vdd.n630 9.3005
R20916 vdd.n3585 vdd.n3584 9.3005
R20917 vdd.n3586 vdd.n629 9.3005
R20918 vdd.n3588 vdd.n3587 9.3005
R20919 vdd.n3590 vdd.n628 9.3005
R20920 vdd.n3592 vdd.n3591 9.3005
R20921 vdd.n3593 vdd.n627 9.3005
R20922 vdd.n3595 vdd.n3594 9.3005
R20923 vdd.n3597 vdd.n626 9.3005
R20924 vdd.n3599 vdd.n3598 9.3005
R20925 vdd.n3600 vdd.n625 9.3005
R20926 vdd.n3602 vdd.n3601 9.3005
R20927 vdd.n3605 vdd.n624 9.3005
R20928 vdd.n3607 vdd.n3606 9.3005
R20929 vdd.n3608 vdd.n623 9.3005
R20930 vdd.n3610 vdd.n3609 9.3005
R20931 vdd.n3612 vdd.n622 9.3005
R20932 vdd.n3614 vdd.n3613 9.3005
R20933 vdd.n3615 vdd.n621 9.3005
R20934 vdd.n3617 vdd.n3616 9.3005
R20935 vdd.n3619 vdd.n620 9.3005
R20936 vdd.n3621 vdd.n3620 9.3005
R20937 vdd.n3499 vdd.n686 9.3005
R20938 vdd.n3498 vdd.n3497 9.3005
R20939 vdd.n3367 vdd.n687 9.3005
R20940 vdd.n3376 vdd.n783 9.3005
R20941 vdd.n3379 vdd.n782 9.3005
R20942 vdd.n3380 vdd.n781 9.3005
R20943 vdd.n3383 vdd.n780 9.3005
R20944 vdd.n3384 vdd.n779 9.3005
R20945 vdd.n3387 vdd.n778 9.3005
R20946 vdd.n3388 vdd.n777 9.3005
R20947 vdd.n3391 vdd.n776 9.3005
R20948 vdd.n3392 vdd.n775 9.3005
R20949 vdd.n3395 vdd.n774 9.3005
R20950 vdd.n3396 vdd.n773 9.3005
R20951 vdd.n3399 vdd.n772 9.3005
R20952 vdd.n3400 vdd.n771 9.3005
R20953 vdd.n3403 vdd.n770 9.3005
R20954 vdd.n3407 vdd.n3406 9.3005
R20955 vdd.n3408 vdd.n767 9.3005
R20956 vdd.n2366 vdd.n2365 9.3005
R20957 vdd.n2361 vdd.n1517 9.3005
R20958 vdd.n1885 vdd.n1884 9.3005
R20959 vdd.n1886 vdd.n1640 9.3005
R20960 vdd.n1888 vdd.n1887 9.3005
R20961 vdd.n1630 vdd.n1629 9.3005
R20962 vdd.n1902 vdd.n1901 9.3005
R20963 vdd.n1903 vdd.n1628 9.3005
R20964 vdd.n1905 vdd.n1904 9.3005
R20965 vdd.n1620 vdd.n1619 9.3005
R20966 vdd.n1919 vdd.n1918 9.3005
R20967 vdd.n1920 vdd.n1618 9.3005
R20968 vdd.n1922 vdd.n1921 9.3005
R20969 vdd.n1607 vdd.n1606 9.3005
R20970 vdd.n1935 vdd.n1934 9.3005
R20971 vdd.n1936 vdd.n1605 9.3005
R20972 vdd.n1938 vdd.n1937 9.3005
R20973 vdd.n1596 vdd.n1595 9.3005
R20974 vdd.n1952 vdd.n1951 9.3005
R20975 vdd.n1953 vdd.n1594 9.3005
R20976 vdd.n1955 vdd.n1954 9.3005
R20977 vdd.n1585 vdd.n1584 9.3005
R20978 vdd.n2275 vdd.n2274 9.3005
R20979 vdd.n2276 vdd.n1583 9.3005
R20980 vdd.n2278 vdd.n2277 9.3005
R20981 vdd.n1573 vdd.n1572 9.3005
R20982 vdd.n2292 vdd.n2291 9.3005
R20983 vdd.n2293 vdd.n1571 9.3005
R20984 vdd.n2295 vdd.n2294 9.3005
R20985 vdd.n1563 vdd.n1562 9.3005
R20986 vdd.n2309 vdd.n2308 9.3005
R20987 vdd.n2310 vdd.n1561 9.3005
R20988 vdd.n2312 vdd.n2311 9.3005
R20989 vdd.n1550 vdd.n1549 9.3005
R20990 vdd.n2325 vdd.n2324 9.3005
R20991 vdd.n2326 vdd.n1548 9.3005
R20992 vdd.n2328 vdd.n2327 9.3005
R20993 vdd.n1540 vdd.n1539 9.3005
R20994 vdd.n2342 vdd.n2341 9.3005
R20995 vdd.n2343 vdd.n1537 9.3005
R20996 vdd.n2347 vdd.n2346 9.3005
R20997 vdd.n2345 vdd.n1538 9.3005
R20998 vdd.n2344 vdd.n1528 9.3005
R20999 vdd.n1642 vdd.n1641 9.3005
R21000 vdd.n1778 vdd.n1777 9.3005
R21001 vdd.n1779 vdd.n1768 9.3005
R21002 vdd.n1781 vdd.n1780 9.3005
R21003 vdd.n1782 vdd.n1767 9.3005
R21004 vdd.n1784 vdd.n1783 9.3005
R21005 vdd.n1785 vdd.n1762 9.3005
R21006 vdd.n1787 vdd.n1786 9.3005
R21007 vdd.n1788 vdd.n1761 9.3005
R21008 vdd.n1790 vdd.n1789 9.3005
R21009 vdd.n1791 vdd.n1756 9.3005
R21010 vdd.n1793 vdd.n1792 9.3005
R21011 vdd.n1794 vdd.n1755 9.3005
R21012 vdd.n1796 vdd.n1795 9.3005
R21013 vdd.n1797 vdd.n1750 9.3005
R21014 vdd.n1799 vdd.n1798 9.3005
R21015 vdd.n1800 vdd.n1749 9.3005
R21016 vdd.n1802 vdd.n1801 9.3005
R21017 vdd.n1803 vdd.n1744 9.3005
R21018 vdd.n1805 vdd.n1804 9.3005
R21019 vdd.n1806 vdd.n1743 9.3005
R21020 vdd.n1808 vdd.n1807 9.3005
R21021 vdd.n1812 vdd.n1739 9.3005
R21022 vdd.n1814 vdd.n1813 9.3005
R21023 vdd.n1815 vdd.n1738 9.3005
R21024 vdd.n1817 vdd.n1816 9.3005
R21025 vdd.n1818 vdd.n1733 9.3005
R21026 vdd.n1820 vdd.n1819 9.3005
R21027 vdd.n1821 vdd.n1732 9.3005
R21028 vdd.n1823 vdd.n1822 9.3005
R21029 vdd.n1824 vdd.n1727 9.3005
R21030 vdd.n1826 vdd.n1825 9.3005
R21031 vdd.n1827 vdd.n1726 9.3005
R21032 vdd.n1829 vdd.n1828 9.3005
R21033 vdd.n1830 vdd.n1721 9.3005
R21034 vdd.n1832 vdd.n1831 9.3005
R21035 vdd.n1833 vdd.n1720 9.3005
R21036 vdd.n1835 vdd.n1834 9.3005
R21037 vdd.n1836 vdd.n1715 9.3005
R21038 vdd.n1838 vdd.n1837 9.3005
R21039 vdd.n1839 vdd.n1714 9.3005
R21040 vdd.n1841 vdd.n1840 9.3005
R21041 vdd.n1842 vdd.n1709 9.3005
R21042 vdd.n1844 vdd.n1843 9.3005
R21043 vdd.n1845 vdd.n1708 9.3005
R21044 vdd.n1847 vdd.n1846 9.3005
R21045 vdd.n1848 vdd.n1701 9.3005
R21046 vdd.n1850 vdd.n1849 9.3005
R21047 vdd.n1851 vdd.n1700 9.3005
R21048 vdd.n1853 vdd.n1852 9.3005
R21049 vdd.n1854 vdd.n1695 9.3005
R21050 vdd.n1856 vdd.n1855 9.3005
R21051 vdd.n1857 vdd.n1694 9.3005
R21052 vdd.n1859 vdd.n1858 9.3005
R21053 vdd.n1860 vdd.n1689 9.3005
R21054 vdd.n1862 vdd.n1861 9.3005
R21055 vdd.n1863 vdd.n1688 9.3005
R21056 vdd.n1865 vdd.n1864 9.3005
R21057 vdd.n1866 vdd.n1683 9.3005
R21058 vdd.n1868 vdd.n1867 9.3005
R21059 vdd.n1869 vdd.n1682 9.3005
R21060 vdd.n1871 vdd.n1870 9.3005
R21061 vdd.n1647 vdd.n1646 9.3005
R21062 vdd.n1877 vdd.n1876 9.3005
R21063 vdd.n1776 vdd.n1775 9.3005
R21064 vdd.n1880 vdd.n1879 9.3005
R21065 vdd.n1636 vdd.n1635 9.3005
R21066 vdd.n1894 vdd.n1893 9.3005
R21067 vdd.n1895 vdd.n1634 9.3005
R21068 vdd.n1897 vdd.n1896 9.3005
R21069 vdd.n1625 vdd.n1624 9.3005
R21070 vdd.n1911 vdd.n1910 9.3005
R21071 vdd.n1912 vdd.n1623 9.3005
R21072 vdd.n1914 vdd.n1913 9.3005
R21073 vdd.n1614 vdd.n1613 9.3005
R21074 vdd.n1927 vdd.n1926 9.3005
R21075 vdd.n1928 vdd.n1612 9.3005
R21076 vdd.n1930 vdd.n1929 9.3005
R21077 vdd.n1602 vdd.n1601 9.3005
R21078 vdd.n1944 vdd.n1943 9.3005
R21079 vdd.n1945 vdd.n1600 9.3005
R21080 vdd.n1947 vdd.n1946 9.3005
R21081 vdd.n1591 vdd.n1590 9.3005
R21082 vdd.n1960 vdd.n1959 9.3005
R21083 vdd.n1961 vdd.n1589 9.3005
R21084 vdd.n1878 vdd.n1645 9.3005
R21085 vdd.n2181 vdd.n2180 9.3005
R21086 vdd.n2176 vdd.n2175 9.3005
R21087 vdd.n2187 vdd.n2186 9.3005
R21088 vdd.n2189 vdd.n2188 9.3005
R21089 vdd.n2172 vdd.n2171 9.3005
R21090 vdd.n2195 vdd.n2194 9.3005
R21091 vdd.n2197 vdd.n2196 9.3005
R21092 vdd.n2169 vdd.n2166 9.3005
R21093 vdd.n2204 vdd.n2203 9.3005
R21094 vdd.n2240 vdd.n2239 9.3005
R21095 vdd.n2235 vdd.n2234 9.3005
R21096 vdd.n2246 vdd.n2245 9.3005
R21097 vdd.n2248 vdd.n2247 9.3005
R21098 vdd.n2231 vdd.n2230 9.3005
R21099 vdd.n2254 vdd.n2253 9.3005
R21100 vdd.n2256 vdd.n2255 9.3005
R21101 vdd.n2228 vdd.n2225 9.3005
R21102 vdd.n2263 vdd.n2262 9.3005
R21103 vdd.n2079 vdd.n2078 9.3005
R21104 vdd.n2074 vdd.n2073 9.3005
R21105 vdd.n2085 vdd.n2084 9.3005
R21106 vdd.n2087 vdd.n2086 9.3005
R21107 vdd.n2070 vdd.n2069 9.3005
R21108 vdd.n2093 vdd.n2092 9.3005
R21109 vdd.n2095 vdd.n2094 9.3005
R21110 vdd.n2067 vdd.n2064 9.3005
R21111 vdd.n2102 vdd.n2101 9.3005
R21112 vdd.n2138 vdd.n2137 9.3005
R21113 vdd.n2133 vdd.n2132 9.3005
R21114 vdd.n2144 vdd.n2143 9.3005
R21115 vdd.n2146 vdd.n2145 9.3005
R21116 vdd.n2129 vdd.n2128 9.3005
R21117 vdd.n2152 vdd.n2151 9.3005
R21118 vdd.n2154 vdd.n2153 9.3005
R21119 vdd.n2126 vdd.n2123 9.3005
R21120 vdd.n2161 vdd.n2160 9.3005
R21121 vdd.n1978 vdd.n1977 9.3005
R21122 vdd.n1973 vdd.n1972 9.3005
R21123 vdd.n1984 vdd.n1983 9.3005
R21124 vdd.n1986 vdd.n1985 9.3005
R21125 vdd.n1969 vdd.n1968 9.3005
R21126 vdd.n1992 vdd.n1991 9.3005
R21127 vdd.n1994 vdd.n1993 9.3005
R21128 vdd.n1966 vdd.n1963 9.3005
R21129 vdd.n2001 vdd.n2000 9.3005
R21130 vdd.n2037 vdd.n2036 9.3005
R21131 vdd.n2032 vdd.n2031 9.3005
R21132 vdd.n2043 vdd.n2042 9.3005
R21133 vdd.n2045 vdd.n2044 9.3005
R21134 vdd.n2028 vdd.n2027 9.3005
R21135 vdd.n2051 vdd.n2050 9.3005
R21136 vdd.n2053 vdd.n2052 9.3005
R21137 vdd.n2025 vdd.n2022 9.3005
R21138 vdd.n2060 vdd.n2059 9.3005
R21139 vdd.n1916 vdd.t217 9.18308
R21140 vdd.n3603 vdd.t90 9.18308
R21141 vdd.n1610 vdd.t164 8.95635
R21142 vdd.n2358 vdd.t17 8.95635
R21143 vdd.n723 vdd.t34 8.95635
R21144 vdd.t162 vdd.n3657 8.95635
R21145 vdd.n312 vdd.n311 8.92171
R21146 vdd.n253 vdd.n252 8.92171
R21147 vdd.n210 vdd.n209 8.92171
R21148 vdd.n151 vdd.n150 8.92171
R21149 vdd.n109 vdd.n108 8.92171
R21150 vdd.n50 vdd.n49 8.92171
R21151 vdd.n2186 vdd.n2185 8.92171
R21152 vdd.n2245 vdd.n2244 8.92171
R21153 vdd.n2084 vdd.n2083 8.92171
R21154 vdd.n2143 vdd.n2142 8.92171
R21155 vdd.n1983 vdd.n1982 8.92171
R21156 vdd.n2042 vdd.n2041 8.92171
R21157 vdd.n231 vdd.n129 8.81535
R21158 vdd.n2164 vdd.n2062 8.81535
R21159 vdd.n1957 vdd.t88 8.72962
R21160 vdd.t205 vdd.n3666 8.72962
R21161 vdd.n2280 vdd.t96 8.50289
R21162 vdd.n3572 vdd.t152 8.50289
R21163 vdd.n28 vdd.n14 8.42249
R21164 vdd.n2306 vdd.t125 8.27616
R21165 vdd.t200 vdd.n656 8.27616
R21166 vdd.n3672 vdd.n3671 8.16225
R21167 vdd.n2268 vdd.n2267 8.16225
R21168 vdd.n308 vdd.n302 8.14595
R21169 vdd.n249 vdd.n243 8.14595
R21170 vdd.n206 vdd.n200 8.14595
R21171 vdd.n147 vdd.n141 8.14595
R21172 vdd.n105 vdd.n99 8.14595
R21173 vdd.n46 vdd.n40 8.14595
R21174 vdd.n2182 vdd.n2176 8.14595
R21175 vdd.n2241 vdd.n2235 8.14595
R21176 vdd.n2080 vdd.n2074 8.14595
R21177 vdd.n2139 vdd.n2133 8.14595
R21178 vdd.n1979 vdd.n1973 8.14595
R21179 vdd.n2038 vdd.n2032 8.14595
R21180 vdd.n1553 vdd.t180 8.04943
R21181 vdd.n3528 vdd.t140 8.04943
R21182 vdd.n2513 vdd.n1134 7.70933
R21183 vdd.n2513 vdd.n1137 7.70933
R21184 vdd.n2519 vdd.n1123 7.70933
R21185 vdd.n2525 vdd.n1123 7.70933
R21186 vdd.n2525 vdd.n1116 7.70933
R21187 vdd.n2531 vdd.n1116 7.70933
R21188 vdd.n2531 vdd.n1119 7.70933
R21189 vdd.n2537 vdd.n1112 7.70933
R21190 vdd.n2543 vdd.n1106 7.70933
R21191 vdd.n2549 vdd.n1093 7.70933
R21192 vdd.n2555 vdd.n1093 7.70933
R21193 vdd.n2561 vdd.n1087 7.70933
R21194 vdd.n2567 vdd.n1080 7.70933
R21195 vdd.n2567 vdd.n1083 7.70933
R21196 vdd.n2573 vdd.n1076 7.70933
R21197 vdd.n2580 vdd.n1062 7.70933
R21198 vdd.n2586 vdd.n1062 7.70933
R21199 vdd.n2592 vdd.n1056 7.70933
R21200 vdd.n2598 vdd.n1052 7.70933
R21201 vdd.n2604 vdd.n1046 7.70933
R21202 vdd.n2622 vdd.n1028 7.70933
R21203 vdd.n2622 vdd.n1021 7.70933
R21204 vdd.n2630 vdd.n1021 7.70933
R21205 vdd.n2712 vdd.n1005 7.70933
R21206 vdd.n3095 vdd.n957 7.70933
R21207 vdd.n3107 vdd.n946 7.70933
R21208 vdd.n3107 vdd.n940 7.70933
R21209 vdd.n3113 vdd.n940 7.70933
R21210 vdd.n3125 vdd.n931 7.70933
R21211 vdd.n3131 vdd.n925 7.70933
R21212 vdd.n3143 vdd.n912 7.70933
R21213 vdd.n3150 vdd.n905 7.70933
R21214 vdd.n3150 vdd.n908 7.70933
R21215 vdd.n3156 vdd.n901 7.70933
R21216 vdd.n3162 vdd.n887 7.70933
R21217 vdd.n3168 vdd.n887 7.70933
R21218 vdd.n3174 vdd.n881 7.70933
R21219 vdd.n3180 vdd.n874 7.70933
R21220 vdd.n3180 vdd.n877 7.70933
R21221 vdd.n3186 vdd.n870 7.70933
R21222 vdd.n3192 vdd.n864 7.70933
R21223 vdd.n3198 vdd.n851 7.70933
R21224 vdd.n3204 vdd.n851 7.70933
R21225 vdd.n3204 vdd.n843 7.70933
R21226 vdd.n3255 vdd.n843 7.70933
R21227 vdd.n3255 vdd.n846 7.70933
R21228 vdd.n3261 vdd.n805 7.70933
R21229 vdd.n3331 vdd.n805 7.70933
R21230 vdd.n307 vdd.n304 7.3702
R21231 vdd.n248 vdd.n245 7.3702
R21232 vdd.n205 vdd.n202 7.3702
R21233 vdd.n146 vdd.n143 7.3702
R21234 vdd.n104 vdd.n101 7.3702
R21235 vdd.n45 vdd.n42 7.3702
R21236 vdd.n2181 vdd.n2178 7.3702
R21237 vdd.n2240 vdd.n2237 7.3702
R21238 vdd.n2079 vdd.n2076 7.3702
R21239 vdd.n2138 vdd.n2135 7.3702
R21240 vdd.n1978 vdd.n1975 7.3702
R21241 vdd.n2037 vdd.n2034 7.3702
R21242 vdd.n1106 vdd.t301 7.36923
R21243 vdd.n3186 vdd.t280 7.36923
R21244 vdd.n2339 vdd.t130 7.1425
R21245 vdd.n2537 vdd.t253 7.1425
R21246 vdd.n1425 vdd.t249 7.1425
R21247 vdd.n3119 vdd.t252 7.1425
R21248 vdd.n864 vdd.t262 7.1425
R21249 vdd.n679 vdd.t169 7.1425
R21250 vdd.n1813 vdd.n1812 6.98232
R21251 vdd.n2401 vdd.n2400 6.98232
R21252 vdd.n566 vdd.n565 6.98232
R21253 vdd.n3413 vdd.n3410 6.98232
R21254 vdd.t98 vdd.n1552 6.91577
R21255 vdd.n3536 vdd.t113 6.91577
R21256 vdd.n1425 vdd.t250 6.80241
R21257 vdd.n3119 vdd.t294 6.80241
R21258 vdd.n2298 vdd.t92 6.68904
R21259 vdd.n3552 vdd.t167 6.68904
R21260 vdd.t178 vdd.n1581 6.46231
R21261 vdd.n2561 vdd.t260 6.46231
R21262 vdd.t265 vdd.n1056 6.46231
R21263 vdd.n3143 vdd.t272 6.46231
R21264 vdd.t286 vdd.n881 6.46231
R21265 vdd.n3580 vdd.t144 6.46231
R21266 vdd.n3672 vdd.n333 6.38151
R21267 vdd.n2267 vdd.n2266 6.38151
R21268 vdd.n2637 vdd.t298 6.34895
R21269 vdd.n3016 vdd.t283 6.34895
R21270 vdd.n3158 vdd.n897 6.2444
R21271 vdd.n2577 vdd.n2576 6.2444
R21272 vdd.n1949 vdd.t198 6.23558
R21273 vdd.t138 vdd.n344 6.23558
R21274 vdd.t182 vdd.n1609 6.00885
R21275 vdd.n3651 vdd.t108 6.00885
R21276 vdd.n2598 vdd.t291 5.89549
R21277 vdd.n925 vdd.t266 5.89549
R21278 vdd.n308 vdd.n307 5.81868
R21279 vdd.n249 vdd.n248 5.81868
R21280 vdd.n206 vdd.n205 5.81868
R21281 vdd.n147 vdd.n146 5.81868
R21282 vdd.n105 vdd.n104 5.81868
R21283 vdd.n46 vdd.n45 5.81868
R21284 vdd.n2182 vdd.n2181 5.81868
R21285 vdd.n2241 vdd.n2240 5.81868
R21286 vdd.n2080 vdd.n2079 5.81868
R21287 vdd.n2139 vdd.n2138 5.81868
R21288 vdd.n1979 vdd.n1978 5.81868
R21289 vdd.n2038 vdd.n2037 5.81868
R21290 vdd.n1908 vdd.t172 5.78212
R21291 vdd.n3642 vdd.t100 5.78212
R21292 vdd.n2720 vdd.n2719 5.77611
R21293 vdd.n1349 vdd.n1348 5.77611
R21294 vdd.n3028 vdd.n3027 5.77611
R21295 vdd.n3272 vdd.n3271 5.77611
R21296 vdd.n3336 vdd.n801 5.77611
R21297 vdd.n2891 vdd.n2825 5.77611
R21298 vdd.n2645 vdd.n1012 5.77611
R21299 vdd.n1485 vdd.n1317 5.77611
R21300 vdd.n1775 vdd.n1774 5.62474
R21301 vdd.n2364 vdd.n2361 5.62474
R21302 vdd.n3623 vdd.n428 5.62474
R21303 vdd.n3497 vdd.n690 5.62474
R21304 vdd.n1632 vdd.t172 5.55539
R21305 vdd.n2573 vdd.t282 5.55539
R21306 vdd.n901 vdd.t256 5.55539
R21307 vdd.t100 vdd.n3641 5.55539
R21308 vdd.n1924 vdd.t182 5.32866
R21309 vdd.t108 vdd.n3650 5.32866
R21310 vdd.n1940 vdd.t198 5.10193
R21311 vdd.n3659 vdd.t138 5.10193
R21312 vdd.n311 vdd.n302 5.04292
R21313 vdd.n252 vdd.n243 5.04292
R21314 vdd.n209 vdd.n200 5.04292
R21315 vdd.n150 vdd.n141 5.04292
R21316 vdd.n108 vdd.n99 5.04292
R21317 vdd.n49 vdd.n40 5.04292
R21318 vdd.n2185 vdd.n2176 5.04292
R21319 vdd.n2244 vdd.n2235 5.04292
R21320 vdd.n2083 vdd.n2074 5.04292
R21321 vdd.n2142 vdd.n2133 5.04292
R21322 vdd.n1982 vdd.n1973 5.04292
R21323 vdd.n2041 vdd.n2032 5.04292
R21324 vdd.n2272 vdd.t178 4.8752
R21325 vdd.t259 vdd.t273 4.8752
R21326 vdd.t302 vdd.t248 4.8752
R21327 vdd.t144 vdd.n340 4.8752
R21328 vdd.n2721 vdd.n2720 4.83952
R21329 vdd.n1348 vdd.n1347 4.83952
R21330 vdd.n3029 vdd.n3028 4.83952
R21331 vdd.n3273 vdd.n3272 4.83952
R21332 vdd.n801 vdd.n796 4.83952
R21333 vdd.n2888 vdd.n2825 4.83952
R21334 vdd.n2648 vdd.n1012 4.83952
R21335 vdd.n1488 vdd.n1317 4.83952
R21336 vdd.n1399 vdd.t268 4.76184
R21337 vdd.n3101 vdd.t254 4.76184
R21338 vdd.n2369 vdd.n2368 4.74817
R21339 vdd.n1521 vdd.n1516 4.74817
R21340 vdd.n1183 vdd.n1180 4.74817
R21341 vdd.n2462 vdd.n1179 4.74817
R21342 vdd.n2467 vdd.n1180 4.74817
R21343 vdd.n2466 vdd.n1179 4.74817
R21344 vdd.n3490 vdd.n3489 4.74817
R21345 vdd.n3487 vdd.n3486 4.74817
R21346 vdd.n3487 vdd.n732 4.74817
R21347 vdd.n3489 vdd.n729 4.74817
R21348 vdd.n3372 vdd.n784 4.74817
R21349 vdd.n3368 vdd.n3366 4.74817
R21350 vdd.n3371 vdd.n3366 4.74817
R21351 vdd.n3375 vdd.n784 4.74817
R21352 vdd.n2368 vdd.n1279 4.74817
R21353 vdd.n1518 vdd.n1516 4.74817
R21354 vdd.n333 vdd.n332 4.7074
R21355 vdd.n231 vdd.n230 4.7074
R21356 vdd.n2266 vdd.n2265 4.7074
R21357 vdd.n2164 vdd.n2163 4.7074
R21358 vdd.n1575 vdd.t92 4.64847
R21359 vdd.t261 vdd.n1087 4.64847
R21360 vdd.n2592 vdd.t300 4.64847
R21361 vdd.t289 vdd.n912 4.64847
R21362 vdd.n3174 vdd.t285 4.64847
R21363 vdd.n3561 vdd.t167 4.64847
R21364 vdd.n1076 vdd.t65 4.53511
R21365 vdd.n3156 vdd.t38 4.53511
R21366 vdd.n2314 vdd.t98 4.42174
R21367 vdd.n2519 vdd.t13 4.42174
R21368 vdd.n1399 vdd.t54 4.42174
R21369 vdd.n3101 vdd.t61 4.42174
R21370 vdd.n846 vdd.t9 4.42174
R21371 vdd.t113 vdd.n655 4.42174
R21372 vdd.n3147 vdd.n897 4.37123
R21373 vdd.n2578 vdd.n2577 4.37123
R21374 vdd.n2616 vdd.t287 4.30838
R21375 vdd.n3004 vdd.t276 4.30838
R21376 vdd.n312 vdd.n300 4.26717
R21377 vdd.n253 vdd.n241 4.26717
R21378 vdd.n210 vdd.n198 4.26717
R21379 vdd.n151 vdd.n139 4.26717
R21380 vdd.n109 vdd.n97 4.26717
R21381 vdd.n50 vdd.n38 4.26717
R21382 vdd.n2186 vdd.n2174 4.26717
R21383 vdd.n2245 vdd.n2233 4.26717
R21384 vdd.n2084 vdd.n2072 4.26717
R21385 vdd.n2143 vdd.n2131 4.26717
R21386 vdd.n1983 vdd.n1971 4.26717
R21387 vdd.n2042 vdd.n2030 4.26717
R21388 vdd.n2330 vdd.t130 4.19501
R21389 vdd.n3520 vdd.t169 4.19501
R21390 vdd.n333 vdd.n231 4.10845
R21391 vdd.n2266 vdd.n2164 4.10845
R21392 vdd.n289 vdd.t236 4.06363
R21393 vdd.n289 vdd.t119 4.06363
R21394 vdd.n287 vdd.t129 4.06363
R21395 vdd.n287 vdd.t157 4.06363
R21396 vdd.n285 vdd.t197 4.06363
R21397 vdd.n285 vdd.t241 4.06363
R21398 vdd.n283 vdd.t107 4.06363
R21399 vdd.n283 vdd.t159 4.06363
R21400 vdd.n281 vdd.t161 4.06363
R21401 vdd.n281 vdd.t215 4.06363
R21402 vdd.n279 vdd.t219 4.06363
R21403 vdd.n279 vdd.t95 4.06363
R21404 vdd.n277 vdd.t123 4.06363
R21405 vdd.n277 vdd.t190 4.06363
R21406 vdd.n275 vdd.t220 4.06363
R21407 vdd.n275 vdd.t237 4.06363
R21408 vdd.n273 vdd.t242 4.06363
R21409 vdd.n273 vdd.t134 4.06363
R21410 vdd.n187 vdd.t213 4.06363
R21411 vdd.n187 vdd.t101 4.06363
R21412 vdd.n185 vdd.t109 4.06363
R21413 vdd.n185 vdd.t135 4.06363
R21414 vdd.n183 vdd.t188 4.06363
R21415 vdd.n183 vdd.t228 4.06363
R21416 vdd.n181 vdd.t246 4.06363
R21417 vdd.n181 vdd.t139 4.06363
R21418 vdd.n179 vdd.t145 4.06363
R21419 vdd.n179 vdd.t206 4.06363
R21420 vdd.n177 vdd.t203 4.06363
R21421 vdd.n177 vdd.t238 4.06363
R21422 vdd.n175 vdd.t103 4.06363
R21423 vdd.n175 vdd.t168 4.06363
R21424 vdd.n173 vdd.t209 4.06363
R21425 vdd.n173 vdd.t221 4.06363
R21426 vdd.n171 vdd.t230 4.06363
R21427 vdd.n171 vdd.t111 4.06363
R21428 vdd.n86 vdd.t155 4.06363
R21429 vdd.n86 vdd.t233 4.06363
R21430 vdd.n84 vdd.t189 4.06363
R21431 vdd.n84 vdd.t91 4.06363
R21432 vdd.n82 vdd.t163 4.06363
R21433 vdd.n82 vdd.t243 4.06363
R21434 vdd.n80 vdd.t142 4.06363
R21435 vdd.n80 vdd.t224 4.06363
R21436 vdd.n78 vdd.t177 4.06363
R21437 vdd.n78 vdd.t207 4.06363
R21438 vdd.n76 vdd.t153 4.06363
R21439 vdd.n76 vdd.t232 4.06363
R21440 vdd.n74 vdd.t122 4.06363
R21441 vdd.n74 vdd.t216 4.06363
R21442 vdd.n72 vdd.t114 4.06363
R21443 vdd.n72 vdd.t201 4.06363
R21444 vdd.n70 vdd.t141 4.06363
R21445 vdd.n70 vdd.t222 4.06363
R21446 vdd.n2206 vdd.t196 4.06363
R21447 vdd.n2206 vdd.t195 4.06363
R21448 vdd.n2208 vdd.t147 4.06363
R21449 vdd.n2208 vdd.t118 4.06363
R21450 vdd.n2210 vdd.t116 4.06363
R21451 vdd.n2210 vdd.t187 4.06363
R21452 vdd.n2212 vdd.t166 4.06363
R21453 vdd.n2212 vdd.t117 4.06363
R21454 vdd.n2214 vdd.t112 4.06363
R21455 vdd.n2214 vdd.t214 4.06363
R21456 vdd.n2216 vdd.t211 4.06363
R21457 vdd.n2216 vdd.t160 4.06363
R21458 vdd.n2218 vdd.t150 4.06363
R21459 vdd.n2218 vdd.t245 4.06363
R21460 vdd.n2220 vdd.t239 4.06363
R21461 vdd.n2220 vdd.t194 4.06363
R21462 vdd.n2222 vdd.t192 4.06363
R21463 vdd.n2222 vdd.t146 4.06363
R21464 vdd.n2104 vdd.t185 4.06363
R21465 vdd.n2104 vdd.t181 4.06363
R21466 vdd.n2106 vdd.t126 4.06363
R21467 vdd.n2106 vdd.t99 4.06363
R21468 vdd.n2108 vdd.t93 4.06363
R21469 vdd.n2108 vdd.t174 4.06363
R21470 vdd.n2110 vdd.t149 4.06363
R21471 vdd.n2110 vdd.t97 4.06363
R21472 vdd.n2112 vdd.t89 4.06363
R21473 vdd.n2112 vdd.t204 4.06363
R21474 vdd.n2114 vdd.t199 4.06363
R21475 vdd.n2114 vdd.t143 4.06363
R21476 vdd.n2116 vdd.t133 4.06363
R21477 vdd.n2116 vdd.t231 4.06363
R21478 vdd.n2118 vdd.t226 4.06363
R21479 vdd.n2118 vdd.t183 4.06363
R21480 vdd.n2120 vdd.t173 4.06363
R21481 vdd.n2120 vdd.t121 4.06363
R21482 vdd.n2003 vdd.t223 4.06363
R21483 vdd.n2003 vdd.t247 4.06363
R21484 vdd.n2005 vdd.t202 4.06363
R21485 vdd.n2005 vdd.t115 4.06363
R21486 vdd.n2007 vdd.t186 4.06363
R21487 vdd.n2007 vdd.t128 4.06363
R21488 vdd.n2009 vdd.t234 4.06363
R21489 vdd.n2009 vdd.t156 4.06363
R21490 vdd.n2011 vdd.t208 4.06363
R21491 vdd.n2011 vdd.t179 4.06363
R21492 vdd.n2013 vdd.t225 4.06363
R21493 vdd.n2013 vdd.t137 4.06363
R21494 vdd.n2015 vdd.t244 4.06363
R21495 vdd.n2015 vdd.t165 4.06363
R21496 vdd.n2017 vdd.t218 4.06363
R21497 vdd.n2017 vdd.t191 4.06363
R21498 vdd.n2019 vdd.t235 4.06363
R21499 vdd.n2019 vdd.t158 4.06363
R21500 vdd.n1112 vdd.t293 3.96828
R21501 vdd.n2610 vdd.t275 3.96828
R21502 vdd.n2998 vdd.t290 3.96828
R21503 vdd.n3192 vdd.t281 3.96828
R21504 vdd.n26 vdd.t0 3.9605
R21505 vdd.n26 vdd.t306 3.9605
R21506 vdd.n23 vdd.t3 3.9605
R21507 vdd.n23 vdd.t4 3.9605
R21508 vdd.n21 vdd.t305 3.9605
R21509 vdd.n21 vdd.t85 3.9605
R21510 vdd.n20 vdd.t5 3.9605
R21511 vdd.n20 vdd.t2 3.9605
R21512 vdd.n15 vdd.t304 3.9605
R21513 vdd.n15 vdd.t1 3.9605
R21514 vdd.n16 vdd.t87 3.9605
R21515 vdd.n16 vdd.t84 3.9605
R21516 vdd.n18 vdd.t307 3.9605
R21517 vdd.n18 vdd.t6 3.9605
R21518 vdd.n25 vdd.t86 3.9605
R21519 vdd.n25 vdd.t7 3.9605
R21520 vdd.n2543 vdd.t293 3.74155
R21521 vdd.n1046 vdd.t275 3.74155
R21522 vdd.n3125 vdd.t290 3.74155
R21523 vdd.n870 vdd.t281 3.74155
R21524 vdd.n7 vdd.t303 3.61217
R21525 vdd.n7 vdd.t267 3.61217
R21526 vdd.n8 vdd.t277 3.61217
R21527 vdd.n8 vdd.t295 3.61217
R21528 vdd.n10 vdd.t284 3.61217
R21529 vdd.n10 vdd.t255 3.61217
R21530 vdd.n12 vdd.t264 3.61217
R21531 vdd.n12 vdd.t271 3.61217
R21532 vdd.n5 vdd.t297 3.61217
R21533 vdd.n5 vdd.t279 3.61217
R21534 vdd.n3 vdd.t269 3.61217
R21535 vdd.n3 vdd.t299 3.61217
R21536 vdd.n1 vdd.t251 3.61217
R21537 vdd.n1 vdd.t288 3.61217
R21538 vdd.n0 vdd.t292 3.61217
R21539 vdd.n0 vdd.t274 3.61217
R21540 vdd.n316 vdd.n315 3.49141
R21541 vdd.n257 vdd.n256 3.49141
R21542 vdd.n214 vdd.n213 3.49141
R21543 vdd.n155 vdd.n154 3.49141
R21544 vdd.n113 vdd.n112 3.49141
R21545 vdd.n54 vdd.n53 3.49141
R21546 vdd.n2190 vdd.n2189 3.49141
R21547 vdd.n2249 vdd.n2248 3.49141
R21548 vdd.n2088 vdd.n2087 3.49141
R21549 vdd.n2147 vdd.n2146 3.49141
R21550 vdd.n1987 vdd.n1986 3.49141
R21551 vdd.n2046 vdd.n2045 3.49141
R21552 vdd.t287 vdd.n1028 3.40145
R21553 vdd.n2784 vdd.t296 3.40145
R21554 vdd.n3088 vdd.t270 3.40145
R21555 vdd.n3113 vdd.t276 3.40145
R21556 vdd.n2331 vdd.t180 3.28809
R21557 vdd.n1137 vdd.t13 3.28809
R21558 vdd.n2637 vdd.t54 3.28809
R21559 vdd.n3016 vdd.t61 3.28809
R21560 vdd.n3261 vdd.t9 3.28809
R21561 vdd.n3519 vdd.t140 3.28809
R21562 vdd.t125 vdd.n1559 3.06136
R21563 vdd.n2555 vdd.t261 3.06136
R21564 vdd.n1437 vdd.t300 3.06136
R21565 vdd.n3137 vdd.t289 3.06136
R21566 vdd.t285 vdd.n874 3.06136
R21567 vdd.n3544 vdd.t200 3.06136
R21568 vdd.n2630 vdd.t268 2.94799
R21569 vdd.t254 vdd.n946 2.94799
R21570 vdd.n2289 vdd.t96 2.83463
R21571 vdd.n644 vdd.t152 2.83463
R21572 vdd.n319 vdd.n298 2.71565
R21573 vdd.n260 vdd.n239 2.71565
R21574 vdd.n217 vdd.n196 2.71565
R21575 vdd.n158 vdd.n137 2.71565
R21576 vdd.n116 vdd.n95 2.71565
R21577 vdd.n57 vdd.n36 2.71565
R21578 vdd.n2193 vdd.n2172 2.71565
R21579 vdd.n2252 vdd.n2231 2.71565
R21580 vdd.n2091 vdd.n2070 2.71565
R21581 vdd.n2150 vdd.n2129 2.71565
R21582 vdd.n1990 vdd.n1969 2.71565
R21583 vdd.n2049 vdd.n2028 2.71565
R21584 vdd.t88 vdd.n1587 2.6079
R21585 vdd.n3667 vdd.t205 2.6079
R21586 vdd.n2604 vdd.t273 2.49453
R21587 vdd.n931 vdd.t302 2.49453
R21588 vdd.n306 vdd.n305 2.4129
R21589 vdd.n247 vdd.n246 2.4129
R21590 vdd.n204 vdd.n203 2.4129
R21591 vdd.n145 vdd.n144 2.4129
R21592 vdd.n103 vdd.n102 2.4129
R21593 vdd.n44 vdd.n43 2.4129
R21594 vdd.n2180 vdd.n2179 2.4129
R21595 vdd.n2239 vdd.n2238 2.4129
R21596 vdd.n2078 vdd.n2077 2.4129
R21597 vdd.n2137 vdd.n2136 2.4129
R21598 vdd.n1977 vdd.n1976 2.4129
R21599 vdd.n2036 vdd.n2035 2.4129
R21600 vdd.n1941 vdd.t164 2.38117
R21601 vdd.n2349 vdd.t17 2.38117
R21602 vdd.n3503 vdd.t34 2.38117
R21603 vdd.n3658 vdd.t162 2.38117
R21604 vdd.n2474 vdd.n1180 2.27742
R21605 vdd.n2474 vdd.n1179 2.27742
R21606 vdd.n3488 vdd.n3487 2.27742
R21607 vdd.n3489 vdd.n3488 2.27742
R21608 vdd.n3366 vdd.n3365 2.27742
R21609 vdd.n3365 vdd.n784 2.27742
R21610 vdd.n2368 vdd.n2367 2.27742
R21611 vdd.n2367 vdd.n1516 2.27742
R21612 vdd.t217 vdd.n1616 2.15444
R21613 vdd.n1083 vdd.t282 2.15444
R21614 vdd.n2580 vdd.t258 2.15444
R21615 vdd.n908 vdd.t257 2.15444
R21616 vdd.n3162 vdd.t256 2.15444
R21617 vdd.n3649 vdd.t90 2.15444
R21618 vdd.n320 vdd.n296 1.93989
R21619 vdd.n261 vdd.n237 1.93989
R21620 vdd.n218 vdd.n194 1.93989
R21621 vdd.n159 vdd.n135 1.93989
R21622 vdd.n117 vdd.n93 1.93989
R21623 vdd.n58 vdd.n34 1.93989
R21624 vdd.n2194 vdd.n2170 1.93989
R21625 vdd.n2253 vdd.n2229 1.93989
R21626 vdd.n2092 vdd.n2068 1.93989
R21627 vdd.n2151 vdd.n2127 1.93989
R21628 vdd.n1991 vdd.n1967 1.93989
R21629 vdd.n2050 vdd.n2026 1.93989
R21630 vdd.n1899 vdd.t175 1.92771
R21631 vdd.t104 vdd.n375 1.92771
R21632 vdd.n1437 vdd.t291 1.81434
R21633 vdd.n3137 vdd.t266 1.81434
R21634 vdd.n1907 vdd.t120 1.70098
R21635 vdd.n3643 vdd.t154 1.70098
R21636 vdd.n1932 vdd.t132 1.47425
R21637 vdd.n361 vdd.t227 1.47425
R21638 vdd.t298 vdd.n1005 1.36088
R21639 vdd.n3095 vdd.t283 1.36088
R21640 vdd.n1598 vdd.t136 1.24752
R21641 vdd.t260 vdd.n1080 1.24752
R21642 vdd.n2586 vdd.t265 1.24752
R21643 vdd.t272 vdd.n905 1.24752
R21644 vdd.n3168 vdd.t286 1.24752
R21645 vdd.t106 vdd.n3665 1.24752
R21646 vdd.n2267 vdd.n28 1.21639
R21647 vdd vdd.n3672 1.20856
R21648 vdd.n331 vdd.n291 1.16414
R21649 vdd.n324 vdd.n323 1.16414
R21650 vdd.n272 vdd.n232 1.16414
R21651 vdd.n265 vdd.n264 1.16414
R21652 vdd.n229 vdd.n189 1.16414
R21653 vdd.n222 vdd.n221 1.16414
R21654 vdd.n170 vdd.n130 1.16414
R21655 vdd.n163 vdd.n162 1.16414
R21656 vdd.n128 vdd.n88 1.16414
R21657 vdd.n121 vdd.n120 1.16414
R21658 vdd.n69 vdd.n29 1.16414
R21659 vdd.n62 vdd.n61 1.16414
R21660 vdd.n2205 vdd.n2165 1.16414
R21661 vdd.n2198 vdd.n2197 1.16414
R21662 vdd.n2264 vdd.n2224 1.16414
R21663 vdd.n2257 vdd.n2256 1.16414
R21664 vdd.n2103 vdd.n2063 1.16414
R21665 vdd.n2096 vdd.n2095 1.16414
R21666 vdd.n2162 vdd.n2122 1.16414
R21667 vdd.n2155 vdd.n2154 1.16414
R21668 vdd.n2002 vdd.n1962 1.16414
R21669 vdd.n1995 vdd.n1994 1.16414
R21670 vdd.n2061 vdd.n2021 1.16414
R21671 vdd.n2054 vdd.n2053 1.16414
R21672 vdd.n2281 vdd.t148 1.02079
R21673 vdd.t65 vdd.t258 1.02079
R21674 vdd.t257 vdd.t38 1.02079
R21675 vdd.t94 vdd.n633 1.02079
R21676 vdd.n1778 vdd.n1774 0.970197
R21677 vdd.n2365 vdd.n2364 0.970197
R21678 vdd.n618 vdd.n428 0.970197
R21679 vdd.n3367 vdd.n690 0.970197
R21680 vdd.n2610 vdd.t250 0.907421
R21681 vdd.n2998 vdd.t294 0.907421
R21682 vdd.n2297 vdd.t127 0.794056
R21683 vdd.n3553 vdd.t102 0.794056
R21684 vdd.n2322 vdd.t184 0.567326
R21685 vdd.n1119 vdd.t253 0.567326
R21686 vdd.n2616 vdd.t249 0.567326
R21687 vdd.n3004 vdd.t252 0.567326
R21688 vdd.n3198 vdd.t262 0.567326
R21689 vdd.t110 vdd.n662 0.567326
R21690 vdd.n2355 vdd.n1181 0.530988
R21691 vdd.n726 vdd.n682 0.530988
R21692 vdd.n464 vdd.n391 0.530988
R21693 vdd.n3622 vdd.n3621 0.530988
R21694 vdd.n3499 vdd.n3498 0.530988
R21695 vdd.n2344 vdd.n1517 0.530988
R21696 vdd.n1776 vdd.n1641 0.530988
R21697 vdd.n1878 vdd.n1877 0.530988
R21698 vdd.n4 vdd.n2 0.459552
R21699 vdd.n11 vdd.n9 0.459552
R21700 vdd.n329 vdd.n328 0.388379
R21701 vdd.n295 vdd.n293 0.388379
R21702 vdd.n270 vdd.n269 0.388379
R21703 vdd.n236 vdd.n234 0.388379
R21704 vdd.n227 vdd.n226 0.388379
R21705 vdd.n193 vdd.n191 0.388379
R21706 vdd.n168 vdd.n167 0.388379
R21707 vdd.n134 vdd.n132 0.388379
R21708 vdd.n126 vdd.n125 0.388379
R21709 vdd.n92 vdd.n90 0.388379
R21710 vdd.n67 vdd.n66 0.388379
R21711 vdd.n33 vdd.n31 0.388379
R21712 vdd.n2203 vdd.n2202 0.388379
R21713 vdd.n2169 vdd.n2167 0.388379
R21714 vdd.n2262 vdd.n2261 0.388379
R21715 vdd.n2228 vdd.n2226 0.388379
R21716 vdd.n2101 vdd.n2100 0.388379
R21717 vdd.n2067 vdd.n2065 0.388379
R21718 vdd.n2160 vdd.n2159 0.388379
R21719 vdd.n2126 vdd.n2124 0.388379
R21720 vdd.n2000 vdd.n1999 0.388379
R21721 vdd.n1966 vdd.n1964 0.388379
R21722 vdd.n2059 vdd.n2058 0.388379
R21723 vdd.n2025 vdd.n2023 0.388379
R21724 vdd.n19 vdd.n17 0.387128
R21725 vdd.n24 vdd.n22 0.387128
R21726 vdd.n6 vdd.n4 0.358259
R21727 vdd.n13 vdd.n11 0.358259
R21728 vdd.n276 vdd.n274 0.358259
R21729 vdd.n278 vdd.n276 0.358259
R21730 vdd.n280 vdd.n278 0.358259
R21731 vdd.n282 vdd.n280 0.358259
R21732 vdd.n284 vdd.n282 0.358259
R21733 vdd.n286 vdd.n284 0.358259
R21734 vdd.n288 vdd.n286 0.358259
R21735 vdd.n290 vdd.n288 0.358259
R21736 vdd.n332 vdd.n290 0.358259
R21737 vdd.n174 vdd.n172 0.358259
R21738 vdd.n176 vdd.n174 0.358259
R21739 vdd.n178 vdd.n176 0.358259
R21740 vdd.n180 vdd.n178 0.358259
R21741 vdd.n182 vdd.n180 0.358259
R21742 vdd.n184 vdd.n182 0.358259
R21743 vdd.n186 vdd.n184 0.358259
R21744 vdd.n188 vdd.n186 0.358259
R21745 vdd.n230 vdd.n188 0.358259
R21746 vdd.n73 vdd.n71 0.358259
R21747 vdd.n75 vdd.n73 0.358259
R21748 vdd.n77 vdd.n75 0.358259
R21749 vdd.n79 vdd.n77 0.358259
R21750 vdd.n81 vdd.n79 0.358259
R21751 vdd.n83 vdd.n81 0.358259
R21752 vdd.n85 vdd.n83 0.358259
R21753 vdd.n87 vdd.n85 0.358259
R21754 vdd.n129 vdd.n87 0.358259
R21755 vdd.n2265 vdd.n2223 0.358259
R21756 vdd.n2223 vdd.n2221 0.358259
R21757 vdd.n2221 vdd.n2219 0.358259
R21758 vdd.n2219 vdd.n2217 0.358259
R21759 vdd.n2217 vdd.n2215 0.358259
R21760 vdd.n2215 vdd.n2213 0.358259
R21761 vdd.n2213 vdd.n2211 0.358259
R21762 vdd.n2211 vdd.n2209 0.358259
R21763 vdd.n2209 vdd.n2207 0.358259
R21764 vdd.n2163 vdd.n2121 0.358259
R21765 vdd.n2121 vdd.n2119 0.358259
R21766 vdd.n2119 vdd.n2117 0.358259
R21767 vdd.n2117 vdd.n2115 0.358259
R21768 vdd.n2115 vdd.n2113 0.358259
R21769 vdd.n2113 vdd.n2111 0.358259
R21770 vdd.n2111 vdd.n2109 0.358259
R21771 vdd.n2109 vdd.n2107 0.358259
R21772 vdd.n2107 vdd.n2105 0.358259
R21773 vdd.n2062 vdd.n2020 0.358259
R21774 vdd.n2020 vdd.n2018 0.358259
R21775 vdd.n2018 vdd.n2016 0.358259
R21776 vdd.n2016 vdd.n2014 0.358259
R21777 vdd.n2014 vdd.n2012 0.358259
R21778 vdd.n2012 vdd.n2010 0.358259
R21779 vdd.n2010 vdd.n2008 0.358259
R21780 vdd.n2008 vdd.n2006 0.358259
R21781 vdd.n2006 vdd.n2004 0.358259
R21782 vdd.n2549 vdd.t301 0.340595
R21783 vdd.n1052 vdd.t259 0.340595
R21784 vdd.n3131 vdd.t248 0.340595
R21785 vdd.n877 vdd.t280 0.340595
R21786 vdd.n14 vdd.n6 0.334552
R21787 vdd.n14 vdd.n13 0.334552
R21788 vdd.n27 vdd.n19 0.21707
R21789 vdd.n27 vdd.n24 0.21707
R21790 vdd.n330 vdd.n292 0.155672
R21791 vdd.n322 vdd.n292 0.155672
R21792 vdd.n322 vdd.n321 0.155672
R21793 vdd.n321 vdd.n297 0.155672
R21794 vdd.n314 vdd.n297 0.155672
R21795 vdd.n314 vdd.n313 0.155672
R21796 vdd.n313 vdd.n301 0.155672
R21797 vdd.n306 vdd.n301 0.155672
R21798 vdd.n271 vdd.n233 0.155672
R21799 vdd.n263 vdd.n233 0.155672
R21800 vdd.n263 vdd.n262 0.155672
R21801 vdd.n262 vdd.n238 0.155672
R21802 vdd.n255 vdd.n238 0.155672
R21803 vdd.n255 vdd.n254 0.155672
R21804 vdd.n254 vdd.n242 0.155672
R21805 vdd.n247 vdd.n242 0.155672
R21806 vdd.n228 vdd.n190 0.155672
R21807 vdd.n220 vdd.n190 0.155672
R21808 vdd.n220 vdd.n219 0.155672
R21809 vdd.n219 vdd.n195 0.155672
R21810 vdd.n212 vdd.n195 0.155672
R21811 vdd.n212 vdd.n211 0.155672
R21812 vdd.n211 vdd.n199 0.155672
R21813 vdd.n204 vdd.n199 0.155672
R21814 vdd.n169 vdd.n131 0.155672
R21815 vdd.n161 vdd.n131 0.155672
R21816 vdd.n161 vdd.n160 0.155672
R21817 vdd.n160 vdd.n136 0.155672
R21818 vdd.n153 vdd.n136 0.155672
R21819 vdd.n153 vdd.n152 0.155672
R21820 vdd.n152 vdd.n140 0.155672
R21821 vdd.n145 vdd.n140 0.155672
R21822 vdd.n127 vdd.n89 0.155672
R21823 vdd.n119 vdd.n89 0.155672
R21824 vdd.n119 vdd.n118 0.155672
R21825 vdd.n118 vdd.n94 0.155672
R21826 vdd.n111 vdd.n94 0.155672
R21827 vdd.n111 vdd.n110 0.155672
R21828 vdd.n110 vdd.n98 0.155672
R21829 vdd.n103 vdd.n98 0.155672
R21830 vdd.n68 vdd.n30 0.155672
R21831 vdd.n60 vdd.n30 0.155672
R21832 vdd.n60 vdd.n59 0.155672
R21833 vdd.n59 vdd.n35 0.155672
R21834 vdd.n52 vdd.n35 0.155672
R21835 vdd.n52 vdd.n51 0.155672
R21836 vdd.n51 vdd.n39 0.155672
R21837 vdd.n44 vdd.n39 0.155672
R21838 vdd.n2204 vdd.n2166 0.155672
R21839 vdd.n2196 vdd.n2166 0.155672
R21840 vdd.n2196 vdd.n2195 0.155672
R21841 vdd.n2195 vdd.n2171 0.155672
R21842 vdd.n2188 vdd.n2171 0.155672
R21843 vdd.n2188 vdd.n2187 0.155672
R21844 vdd.n2187 vdd.n2175 0.155672
R21845 vdd.n2180 vdd.n2175 0.155672
R21846 vdd.n2263 vdd.n2225 0.155672
R21847 vdd.n2255 vdd.n2225 0.155672
R21848 vdd.n2255 vdd.n2254 0.155672
R21849 vdd.n2254 vdd.n2230 0.155672
R21850 vdd.n2247 vdd.n2230 0.155672
R21851 vdd.n2247 vdd.n2246 0.155672
R21852 vdd.n2246 vdd.n2234 0.155672
R21853 vdd.n2239 vdd.n2234 0.155672
R21854 vdd.n2102 vdd.n2064 0.155672
R21855 vdd.n2094 vdd.n2064 0.155672
R21856 vdd.n2094 vdd.n2093 0.155672
R21857 vdd.n2093 vdd.n2069 0.155672
R21858 vdd.n2086 vdd.n2069 0.155672
R21859 vdd.n2086 vdd.n2085 0.155672
R21860 vdd.n2085 vdd.n2073 0.155672
R21861 vdd.n2078 vdd.n2073 0.155672
R21862 vdd.n2161 vdd.n2123 0.155672
R21863 vdd.n2153 vdd.n2123 0.155672
R21864 vdd.n2153 vdd.n2152 0.155672
R21865 vdd.n2152 vdd.n2128 0.155672
R21866 vdd.n2145 vdd.n2128 0.155672
R21867 vdd.n2145 vdd.n2144 0.155672
R21868 vdd.n2144 vdd.n2132 0.155672
R21869 vdd.n2137 vdd.n2132 0.155672
R21870 vdd.n2001 vdd.n1963 0.155672
R21871 vdd.n1993 vdd.n1963 0.155672
R21872 vdd.n1993 vdd.n1992 0.155672
R21873 vdd.n1992 vdd.n1968 0.155672
R21874 vdd.n1985 vdd.n1968 0.155672
R21875 vdd.n1985 vdd.n1984 0.155672
R21876 vdd.n1984 vdd.n1972 0.155672
R21877 vdd.n1977 vdd.n1972 0.155672
R21878 vdd.n2060 vdd.n2022 0.155672
R21879 vdd.n2052 vdd.n2022 0.155672
R21880 vdd.n2052 vdd.n2051 0.155672
R21881 vdd.n2051 vdd.n2027 0.155672
R21882 vdd.n2044 vdd.n2027 0.155672
R21883 vdd.n2044 vdd.n2043 0.155672
R21884 vdd.n2043 vdd.n2031 0.155672
R21885 vdd.n2036 vdd.n2031 0.155672
R21886 vdd.n1186 vdd.n1178 0.152939
R21887 vdd.n1190 vdd.n1186 0.152939
R21888 vdd.n1191 vdd.n1190 0.152939
R21889 vdd.n1192 vdd.n1191 0.152939
R21890 vdd.n1193 vdd.n1192 0.152939
R21891 vdd.n1197 vdd.n1193 0.152939
R21892 vdd.n1198 vdd.n1197 0.152939
R21893 vdd.n1199 vdd.n1198 0.152939
R21894 vdd.n1200 vdd.n1199 0.152939
R21895 vdd.n1204 vdd.n1200 0.152939
R21896 vdd.n1205 vdd.n1204 0.152939
R21897 vdd.n1206 vdd.n1205 0.152939
R21898 vdd.n2438 vdd.n1206 0.152939
R21899 vdd.n2438 vdd.n2437 0.152939
R21900 vdd.n2437 vdd.n2436 0.152939
R21901 vdd.n2436 vdd.n1212 0.152939
R21902 vdd.n1217 vdd.n1212 0.152939
R21903 vdd.n1218 vdd.n1217 0.152939
R21904 vdd.n1219 vdd.n1218 0.152939
R21905 vdd.n1223 vdd.n1219 0.152939
R21906 vdd.n1224 vdd.n1223 0.152939
R21907 vdd.n1225 vdd.n1224 0.152939
R21908 vdd.n1226 vdd.n1225 0.152939
R21909 vdd.n1230 vdd.n1226 0.152939
R21910 vdd.n1231 vdd.n1230 0.152939
R21911 vdd.n1232 vdd.n1231 0.152939
R21912 vdd.n1233 vdd.n1232 0.152939
R21913 vdd.n1237 vdd.n1233 0.152939
R21914 vdd.n1238 vdd.n1237 0.152939
R21915 vdd.n1239 vdd.n1238 0.152939
R21916 vdd.n1240 vdd.n1239 0.152939
R21917 vdd.n1244 vdd.n1240 0.152939
R21918 vdd.n1245 vdd.n1244 0.152939
R21919 vdd.n1246 vdd.n1245 0.152939
R21920 vdd.n2399 vdd.n1246 0.152939
R21921 vdd.n2399 vdd.n2398 0.152939
R21922 vdd.n2398 vdd.n2397 0.152939
R21923 vdd.n2397 vdd.n1252 0.152939
R21924 vdd.n1257 vdd.n1252 0.152939
R21925 vdd.n1258 vdd.n1257 0.152939
R21926 vdd.n1259 vdd.n1258 0.152939
R21927 vdd.n1263 vdd.n1259 0.152939
R21928 vdd.n1264 vdd.n1263 0.152939
R21929 vdd.n1265 vdd.n1264 0.152939
R21930 vdd.n1266 vdd.n1265 0.152939
R21931 vdd.n1270 vdd.n1266 0.152939
R21932 vdd.n1271 vdd.n1270 0.152939
R21933 vdd.n1272 vdd.n1271 0.152939
R21934 vdd.n1273 vdd.n1272 0.152939
R21935 vdd.n1277 vdd.n1273 0.152939
R21936 vdd.n1278 vdd.n1277 0.152939
R21937 vdd.n2473 vdd.n1181 0.152939
R21938 vdd.n2269 vdd.n1578 0.152939
R21939 vdd.n2284 vdd.n1578 0.152939
R21940 vdd.n2285 vdd.n2284 0.152939
R21941 vdd.n2286 vdd.n2285 0.152939
R21942 vdd.n2286 vdd.n1567 0.152939
R21943 vdd.n2301 vdd.n1567 0.152939
R21944 vdd.n2302 vdd.n2301 0.152939
R21945 vdd.n2303 vdd.n2302 0.152939
R21946 vdd.n2303 vdd.n1556 0.152939
R21947 vdd.n2317 vdd.n1556 0.152939
R21948 vdd.n2318 vdd.n2317 0.152939
R21949 vdd.n2319 vdd.n2318 0.152939
R21950 vdd.n2319 vdd.n1544 0.152939
R21951 vdd.n2334 vdd.n1544 0.152939
R21952 vdd.n2335 vdd.n2334 0.152939
R21953 vdd.n2336 vdd.n2335 0.152939
R21954 vdd.n2336 vdd.n1532 0.152939
R21955 vdd.n2353 vdd.n1532 0.152939
R21956 vdd.n2354 vdd.n2353 0.152939
R21957 vdd.n2355 vdd.n2354 0.152939
R21958 vdd.n735 vdd.n730 0.152939
R21959 vdd.n736 vdd.n735 0.152939
R21960 vdd.n737 vdd.n736 0.152939
R21961 vdd.n738 vdd.n737 0.152939
R21962 vdd.n739 vdd.n738 0.152939
R21963 vdd.n740 vdd.n739 0.152939
R21964 vdd.n741 vdd.n740 0.152939
R21965 vdd.n742 vdd.n741 0.152939
R21966 vdd.n743 vdd.n742 0.152939
R21967 vdd.n744 vdd.n743 0.152939
R21968 vdd.n745 vdd.n744 0.152939
R21969 vdd.n746 vdd.n745 0.152939
R21970 vdd.n3455 vdd.n746 0.152939
R21971 vdd.n3455 vdd.n3454 0.152939
R21972 vdd.n3454 vdd.n3453 0.152939
R21973 vdd.n3453 vdd.n748 0.152939
R21974 vdd.n749 vdd.n748 0.152939
R21975 vdd.n750 vdd.n749 0.152939
R21976 vdd.n751 vdd.n750 0.152939
R21977 vdd.n752 vdd.n751 0.152939
R21978 vdd.n753 vdd.n752 0.152939
R21979 vdd.n754 vdd.n753 0.152939
R21980 vdd.n755 vdd.n754 0.152939
R21981 vdd.n756 vdd.n755 0.152939
R21982 vdd.n757 vdd.n756 0.152939
R21983 vdd.n758 vdd.n757 0.152939
R21984 vdd.n759 vdd.n758 0.152939
R21985 vdd.n760 vdd.n759 0.152939
R21986 vdd.n761 vdd.n760 0.152939
R21987 vdd.n762 vdd.n761 0.152939
R21988 vdd.n763 vdd.n762 0.152939
R21989 vdd.n764 vdd.n763 0.152939
R21990 vdd.n765 vdd.n764 0.152939
R21991 vdd.n766 vdd.n765 0.152939
R21992 vdd.n3409 vdd.n766 0.152939
R21993 vdd.n3409 vdd.n3408 0.152939
R21994 vdd.n3408 vdd.n3407 0.152939
R21995 vdd.n3407 vdd.n770 0.152939
R21996 vdd.n771 vdd.n770 0.152939
R21997 vdd.n772 vdd.n771 0.152939
R21998 vdd.n773 vdd.n772 0.152939
R21999 vdd.n774 vdd.n773 0.152939
R22000 vdd.n775 vdd.n774 0.152939
R22001 vdd.n776 vdd.n775 0.152939
R22002 vdd.n777 vdd.n776 0.152939
R22003 vdd.n778 vdd.n777 0.152939
R22004 vdd.n779 vdd.n778 0.152939
R22005 vdd.n780 vdd.n779 0.152939
R22006 vdd.n781 vdd.n780 0.152939
R22007 vdd.n782 vdd.n781 0.152939
R22008 vdd.n783 vdd.n782 0.152939
R22009 vdd.n727 vdd.n726 0.152939
R22010 vdd.n3506 vdd.n682 0.152939
R22011 vdd.n3507 vdd.n3506 0.152939
R22012 vdd.n3508 vdd.n3507 0.152939
R22013 vdd.n3508 vdd.n670 0.152939
R22014 vdd.n3523 vdd.n670 0.152939
R22015 vdd.n3524 vdd.n3523 0.152939
R22016 vdd.n3525 vdd.n3524 0.152939
R22017 vdd.n3525 vdd.n659 0.152939
R22018 vdd.n3539 vdd.n659 0.152939
R22019 vdd.n3540 vdd.n3539 0.152939
R22020 vdd.n3541 vdd.n3540 0.152939
R22021 vdd.n3541 vdd.n647 0.152939
R22022 vdd.n3556 vdd.n647 0.152939
R22023 vdd.n3557 vdd.n3556 0.152939
R22024 vdd.n3558 vdd.n3557 0.152939
R22025 vdd.n3558 vdd.n636 0.152939
R22026 vdd.n3575 vdd.n636 0.152939
R22027 vdd.n3576 vdd.n3575 0.152939
R22028 vdd.n3577 vdd.n3576 0.152939
R22029 vdd.n3577 vdd.n334 0.152939
R22030 vdd.n3670 vdd.n335 0.152939
R22031 vdd.n346 vdd.n335 0.152939
R22032 vdd.n347 vdd.n346 0.152939
R22033 vdd.n348 vdd.n347 0.152939
R22034 vdd.n355 vdd.n348 0.152939
R22035 vdd.n356 vdd.n355 0.152939
R22036 vdd.n357 vdd.n356 0.152939
R22037 vdd.n358 vdd.n357 0.152939
R22038 vdd.n366 vdd.n358 0.152939
R22039 vdd.n367 vdd.n366 0.152939
R22040 vdd.n368 vdd.n367 0.152939
R22041 vdd.n369 vdd.n368 0.152939
R22042 vdd.n377 vdd.n369 0.152939
R22043 vdd.n378 vdd.n377 0.152939
R22044 vdd.n379 vdd.n378 0.152939
R22045 vdd.n380 vdd.n379 0.152939
R22046 vdd.n388 vdd.n380 0.152939
R22047 vdd.n389 vdd.n388 0.152939
R22048 vdd.n390 vdd.n389 0.152939
R22049 vdd.n391 vdd.n390 0.152939
R22050 vdd.n464 vdd.n463 0.152939
R22051 vdd.n470 vdd.n463 0.152939
R22052 vdd.n471 vdd.n470 0.152939
R22053 vdd.n472 vdd.n471 0.152939
R22054 vdd.n472 vdd.n461 0.152939
R22055 vdd.n480 vdd.n461 0.152939
R22056 vdd.n481 vdd.n480 0.152939
R22057 vdd.n482 vdd.n481 0.152939
R22058 vdd.n482 vdd.n459 0.152939
R22059 vdd.n490 vdd.n459 0.152939
R22060 vdd.n491 vdd.n490 0.152939
R22061 vdd.n492 vdd.n491 0.152939
R22062 vdd.n492 vdd.n457 0.152939
R22063 vdd.n500 vdd.n457 0.152939
R22064 vdd.n501 vdd.n500 0.152939
R22065 vdd.n502 vdd.n501 0.152939
R22066 vdd.n502 vdd.n455 0.152939
R22067 vdd.n510 vdd.n455 0.152939
R22068 vdd.n511 vdd.n510 0.152939
R22069 vdd.n512 vdd.n511 0.152939
R22070 vdd.n512 vdd.n451 0.152939
R22071 vdd.n520 vdd.n451 0.152939
R22072 vdd.n521 vdd.n520 0.152939
R22073 vdd.n522 vdd.n521 0.152939
R22074 vdd.n522 vdd.n449 0.152939
R22075 vdd.n530 vdd.n449 0.152939
R22076 vdd.n531 vdd.n530 0.152939
R22077 vdd.n532 vdd.n531 0.152939
R22078 vdd.n532 vdd.n447 0.152939
R22079 vdd.n540 vdd.n447 0.152939
R22080 vdd.n541 vdd.n540 0.152939
R22081 vdd.n542 vdd.n541 0.152939
R22082 vdd.n542 vdd.n445 0.152939
R22083 vdd.n550 vdd.n445 0.152939
R22084 vdd.n551 vdd.n550 0.152939
R22085 vdd.n552 vdd.n551 0.152939
R22086 vdd.n552 vdd.n443 0.152939
R22087 vdd.n560 vdd.n443 0.152939
R22088 vdd.n561 vdd.n560 0.152939
R22089 vdd.n562 vdd.n561 0.152939
R22090 vdd.n562 vdd.n439 0.152939
R22091 vdd.n570 vdd.n439 0.152939
R22092 vdd.n571 vdd.n570 0.152939
R22093 vdd.n572 vdd.n571 0.152939
R22094 vdd.n572 vdd.n437 0.152939
R22095 vdd.n580 vdd.n437 0.152939
R22096 vdd.n581 vdd.n580 0.152939
R22097 vdd.n582 vdd.n581 0.152939
R22098 vdd.n582 vdd.n435 0.152939
R22099 vdd.n590 vdd.n435 0.152939
R22100 vdd.n591 vdd.n590 0.152939
R22101 vdd.n592 vdd.n591 0.152939
R22102 vdd.n592 vdd.n433 0.152939
R22103 vdd.n600 vdd.n433 0.152939
R22104 vdd.n601 vdd.n600 0.152939
R22105 vdd.n602 vdd.n601 0.152939
R22106 vdd.n602 vdd.n431 0.152939
R22107 vdd.n610 vdd.n431 0.152939
R22108 vdd.n611 vdd.n610 0.152939
R22109 vdd.n612 vdd.n611 0.152939
R22110 vdd.n612 vdd.n429 0.152939
R22111 vdd.n619 vdd.n429 0.152939
R22112 vdd.n3622 vdd.n619 0.152939
R22113 vdd.n3500 vdd.n3499 0.152939
R22114 vdd.n3500 vdd.n675 0.152939
R22115 vdd.n3514 vdd.n675 0.152939
R22116 vdd.n3515 vdd.n3514 0.152939
R22117 vdd.n3516 vdd.n3515 0.152939
R22118 vdd.n3516 vdd.n665 0.152939
R22119 vdd.n3531 vdd.n665 0.152939
R22120 vdd.n3532 vdd.n3531 0.152939
R22121 vdd.n3533 vdd.n3532 0.152939
R22122 vdd.n3533 vdd.n652 0.152939
R22123 vdd.n3547 vdd.n652 0.152939
R22124 vdd.n3548 vdd.n3547 0.152939
R22125 vdd.n3549 vdd.n3548 0.152939
R22126 vdd.n3549 vdd.n641 0.152939
R22127 vdd.n3564 vdd.n641 0.152939
R22128 vdd.n3565 vdd.n3564 0.152939
R22129 vdd.n3566 vdd.n3565 0.152939
R22130 vdd.n3568 vdd.n3566 0.152939
R22131 vdd.n3568 vdd.n3567 0.152939
R22132 vdd.n3567 vdd.n630 0.152939
R22133 vdd.n3585 vdd.n630 0.152939
R22134 vdd.n3586 vdd.n3585 0.152939
R22135 vdd.n3587 vdd.n3586 0.152939
R22136 vdd.n3587 vdd.n628 0.152939
R22137 vdd.n3592 vdd.n628 0.152939
R22138 vdd.n3593 vdd.n3592 0.152939
R22139 vdd.n3594 vdd.n3593 0.152939
R22140 vdd.n3594 vdd.n626 0.152939
R22141 vdd.n3599 vdd.n626 0.152939
R22142 vdd.n3600 vdd.n3599 0.152939
R22143 vdd.n3601 vdd.n3600 0.152939
R22144 vdd.n3601 vdd.n624 0.152939
R22145 vdd.n3607 vdd.n624 0.152939
R22146 vdd.n3608 vdd.n3607 0.152939
R22147 vdd.n3609 vdd.n3608 0.152939
R22148 vdd.n3609 vdd.n622 0.152939
R22149 vdd.n3614 vdd.n622 0.152939
R22150 vdd.n3615 vdd.n3614 0.152939
R22151 vdd.n3616 vdd.n3615 0.152939
R22152 vdd.n3616 vdd.n620 0.152939
R22153 vdd.n3621 vdd.n620 0.152939
R22154 vdd.n3498 vdd.n687 0.152939
R22155 vdd.n2366 vdd.n1517 0.152939
R22156 vdd.n1885 vdd.n1641 0.152939
R22157 vdd.n1886 vdd.n1885 0.152939
R22158 vdd.n1887 vdd.n1886 0.152939
R22159 vdd.n1887 vdd.n1629 0.152939
R22160 vdd.n1902 vdd.n1629 0.152939
R22161 vdd.n1903 vdd.n1902 0.152939
R22162 vdd.n1904 vdd.n1903 0.152939
R22163 vdd.n1904 vdd.n1619 0.152939
R22164 vdd.n1919 vdd.n1619 0.152939
R22165 vdd.n1920 vdd.n1919 0.152939
R22166 vdd.n1921 vdd.n1920 0.152939
R22167 vdd.n1921 vdd.n1606 0.152939
R22168 vdd.n1935 vdd.n1606 0.152939
R22169 vdd.n1936 vdd.n1935 0.152939
R22170 vdd.n1937 vdd.n1936 0.152939
R22171 vdd.n1937 vdd.n1595 0.152939
R22172 vdd.n1952 vdd.n1595 0.152939
R22173 vdd.n1953 vdd.n1952 0.152939
R22174 vdd.n1954 vdd.n1953 0.152939
R22175 vdd.n1954 vdd.n1584 0.152939
R22176 vdd.n2275 vdd.n1584 0.152939
R22177 vdd.n2276 vdd.n2275 0.152939
R22178 vdd.n2277 vdd.n2276 0.152939
R22179 vdd.n2277 vdd.n1572 0.152939
R22180 vdd.n2292 vdd.n1572 0.152939
R22181 vdd.n2293 vdd.n2292 0.152939
R22182 vdd.n2294 vdd.n2293 0.152939
R22183 vdd.n2294 vdd.n1562 0.152939
R22184 vdd.n2309 vdd.n1562 0.152939
R22185 vdd.n2310 vdd.n2309 0.152939
R22186 vdd.n2311 vdd.n2310 0.152939
R22187 vdd.n2311 vdd.n1549 0.152939
R22188 vdd.n2325 vdd.n1549 0.152939
R22189 vdd.n2326 vdd.n2325 0.152939
R22190 vdd.n2327 vdd.n2326 0.152939
R22191 vdd.n2327 vdd.n1539 0.152939
R22192 vdd.n2342 vdd.n1539 0.152939
R22193 vdd.n2343 vdd.n2342 0.152939
R22194 vdd.n2346 vdd.n2343 0.152939
R22195 vdd.n2346 vdd.n2345 0.152939
R22196 vdd.n2345 vdd.n2344 0.152939
R22197 vdd.n1877 vdd.n1646 0.152939
R22198 vdd.n1870 vdd.n1646 0.152939
R22199 vdd.n1870 vdd.n1869 0.152939
R22200 vdd.n1869 vdd.n1868 0.152939
R22201 vdd.n1868 vdd.n1683 0.152939
R22202 vdd.n1864 vdd.n1683 0.152939
R22203 vdd.n1864 vdd.n1863 0.152939
R22204 vdd.n1863 vdd.n1862 0.152939
R22205 vdd.n1862 vdd.n1689 0.152939
R22206 vdd.n1858 vdd.n1689 0.152939
R22207 vdd.n1858 vdd.n1857 0.152939
R22208 vdd.n1857 vdd.n1856 0.152939
R22209 vdd.n1856 vdd.n1695 0.152939
R22210 vdd.n1852 vdd.n1695 0.152939
R22211 vdd.n1852 vdd.n1851 0.152939
R22212 vdd.n1851 vdd.n1850 0.152939
R22213 vdd.n1850 vdd.n1701 0.152939
R22214 vdd.n1846 vdd.n1701 0.152939
R22215 vdd.n1846 vdd.n1845 0.152939
R22216 vdd.n1845 vdd.n1844 0.152939
R22217 vdd.n1844 vdd.n1709 0.152939
R22218 vdd.n1840 vdd.n1709 0.152939
R22219 vdd.n1840 vdd.n1839 0.152939
R22220 vdd.n1839 vdd.n1838 0.152939
R22221 vdd.n1838 vdd.n1715 0.152939
R22222 vdd.n1834 vdd.n1715 0.152939
R22223 vdd.n1834 vdd.n1833 0.152939
R22224 vdd.n1833 vdd.n1832 0.152939
R22225 vdd.n1832 vdd.n1721 0.152939
R22226 vdd.n1828 vdd.n1721 0.152939
R22227 vdd.n1828 vdd.n1827 0.152939
R22228 vdd.n1827 vdd.n1826 0.152939
R22229 vdd.n1826 vdd.n1727 0.152939
R22230 vdd.n1822 vdd.n1727 0.152939
R22231 vdd.n1822 vdd.n1821 0.152939
R22232 vdd.n1821 vdd.n1820 0.152939
R22233 vdd.n1820 vdd.n1733 0.152939
R22234 vdd.n1816 vdd.n1733 0.152939
R22235 vdd.n1816 vdd.n1815 0.152939
R22236 vdd.n1815 vdd.n1814 0.152939
R22237 vdd.n1814 vdd.n1739 0.152939
R22238 vdd.n1807 vdd.n1739 0.152939
R22239 vdd.n1807 vdd.n1806 0.152939
R22240 vdd.n1806 vdd.n1805 0.152939
R22241 vdd.n1805 vdd.n1744 0.152939
R22242 vdd.n1801 vdd.n1744 0.152939
R22243 vdd.n1801 vdd.n1800 0.152939
R22244 vdd.n1800 vdd.n1799 0.152939
R22245 vdd.n1799 vdd.n1750 0.152939
R22246 vdd.n1795 vdd.n1750 0.152939
R22247 vdd.n1795 vdd.n1794 0.152939
R22248 vdd.n1794 vdd.n1793 0.152939
R22249 vdd.n1793 vdd.n1756 0.152939
R22250 vdd.n1789 vdd.n1756 0.152939
R22251 vdd.n1789 vdd.n1788 0.152939
R22252 vdd.n1788 vdd.n1787 0.152939
R22253 vdd.n1787 vdd.n1762 0.152939
R22254 vdd.n1783 vdd.n1762 0.152939
R22255 vdd.n1783 vdd.n1782 0.152939
R22256 vdd.n1782 vdd.n1781 0.152939
R22257 vdd.n1781 vdd.n1768 0.152939
R22258 vdd.n1777 vdd.n1768 0.152939
R22259 vdd.n1777 vdd.n1776 0.152939
R22260 vdd.n1879 vdd.n1878 0.152939
R22261 vdd.n1879 vdd.n1635 0.152939
R22262 vdd.n1894 vdd.n1635 0.152939
R22263 vdd.n1895 vdd.n1894 0.152939
R22264 vdd.n1896 vdd.n1895 0.152939
R22265 vdd.n1896 vdd.n1624 0.152939
R22266 vdd.n1911 vdd.n1624 0.152939
R22267 vdd.n1912 vdd.n1911 0.152939
R22268 vdd.n1913 vdd.n1912 0.152939
R22269 vdd.n1913 vdd.n1613 0.152939
R22270 vdd.n1927 vdd.n1613 0.152939
R22271 vdd.n1928 vdd.n1927 0.152939
R22272 vdd.n1929 vdd.n1928 0.152939
R22273 vdd.n1929 vdd.n1601 0.152939
R22274 vdd.n1944 vdd.n1601 0.152939
R22275 vdd.n1945 vdd.n1944 0.152939
R22276 vdd.n1946 vdd.n1945 0.152939
R22277 vdd.n1946 vdd.n1590 0.152939
R22278 vdd.n1960 vdd.n1590 0.152939
R22279 vdd.n1961 vdd.n1960 0.152939
R22280 vdd.n1882 vdd.t72 0.113865
R22281 vdd.t21 vdd.n386 0.113865
R22282 vdd.n2474 vdd.n2473 0.110256
R22283 vdd.n3488 vdd.n727 0.110256
R22284 vdd.n3365 vdd.n687 0.110256
R22285 vdd.n2367 vdd.n2366 0.110256
R22286 vdd.n2269 vdd.n2268 0.0695946
R22287 vdd.n3671 vdd.n334 0.0695946
R22288 vdd.n3671 vdd.n3670 0.0695946
R22289 vdd.n2268 vdd.n1961 0.0695946
R22290 vdd.n2474 vdd.n1178 0.0431829
R22291 vdd.n2367 vdd.n1278 0.0431829
R22292 vdd.n3488 vdd.n730 0.0431829
R22293 vdd.n3365 vdd.n783 0.0431829
R22294 vdd vdd.n28 0.00833333
R22295 CSoutput.n19 CSoutput.t204 184.661
R22296 CSoutput.n78 CSoutput.n77 165.8
R22297 CSoutput.n76 CSoutput.n0 165.8
R22298 CSoutput.n75 CSoutput.n74 165.8
R22299 CSoutput.n73 CSoutput.n72 165.8
R22300 CSoutput.n71 CSoutput.n2 165.8
R22301 CSoutput.n69 CSoutput.n68 165.8
R22302 CSoutput.n67 CSoutput.n3 165.8
R22303 CSoutput.n66 CSoutput.n65 165.8
R22304 CSoutput.n63 CSoutput.n4 165.8
R22305 CSoutput.n61 CSoutput.n60 165.8
R22306 CSoutput.n59 CSoutput.n5 165.8
R22307 CSoutput.n58 CSoutput.n57 165.8
R22308 CSoutput.n55 CSoutput.n6 165.8
R22309 CSoutput.n54 CSoutput.n53 165.8
R22310 CSoutput.n52 CSoutput.n51 165.8
R22311 CSoutput.n50 CSoutput.n8 165.8
R22312 CSoutput.n48 CSoutput.n47 165.8
R22313 CSoutput.n46 CSoutput.n9 165.8
R22314 CSoutput.n45 CSoutput.n44 165.8
R22315 CSoutput.n42 CSoutput.n10 165.8
R22316 CSoutput.n41 CSoutput.n40 165.8
R22317 CSoutput.n39 CSoutput.n38 165.8
R22318 CSoutput.n37 CSoutput.n12 165.8
R22319 CSoutput.n35 CSoutput.n34 165.8
R22320 CSoutput.n33 CSoutput.n13 165.8
R22321 CSoutput.n32 CSoutput.n31 165.8
R22322 CSoutput.n29 CSoutput.n14 165.8
R22323 CSoutput.n28 CSoutput.n27 165.8
R22324 CSoutput.n26 CSoutput.n25 165.8
R22325 CSoutput.n24 CSoutput.n16 165.8
R22326 CSoutput.n22 CSoutput.n21 165.8
R22327 CSoutput.n20 CSoutput.n17 165.8
R22328 CSoutput.n77 CSoutput.t207 162.194
R22329 CSoutput.n18 CSoutput.t201 120.501
R22330 CSoutput.n23 CSoutput.t218 120.501
R22331 CSoutput.n15 CSoutput.t213 120.501
R22332 CSoutput.n30 CSoutput.t202 120.501
R22333 CSoutput.n36 CSoutput.t203 120.501
R22334 CSoutput.n11 CSoutput.t215 120.501
R22335 CSoutput.n43 CSoutput.t212 120.501
R22336 CSoutput.n49 CSoutput.t206 120.501
R22337 CSoutput.n7 CSoutput.t219 120.501
R22338 CSoutput.n56 CSoutput.t220 120.501
R22339 CSoutput.n62 CSoutput.t209 120.501
R22340 CSoutput.n64 CSoutput.t221 120.501
R22341 CSoutput.n70 CSoutput.t200 120.501
R22342 CSoutput.n1 CSoutput.t217 120.501
R22343 CSoutput.n330 CSoutput.n328 103.469
R22344 CSoutput.n310 CSoutput.n308 103.469
R22345 CSoutput.n291 CSoutput.n289 103.469
R22346 CSoutput.n120 CSoutput.n118 103.469
R22347 CSoutput.n100 CSoutput.n98 103.469
R22348 CSoutput.n81 CSoutput.n79 103.469
R22349 CSoutput.n344 CSoutput.n343 103.111
R22350 CSoutput.n342 CSoutput.n341 103.111
R22351 CSoutput.n340 CSoutput.n339 103.111
R22352 CSoutput.n338 CSoutput.n337 103.111
R22353 CSoutput.n336 CSoutput.n335 103.111
R22354 CSoutput.n334 CSoutput.n333 103.111
R22355 CSoutput.n332 CSoutput.n331 103.111
R22356 CSoutput.n330 CSoutput.n329 103.111
R22357 CSoutput.n326 CSoutput.n325 103.111
R22358 CSoutput.n324 CSoutput.n323 103.111
R22359 CSoutput.n322 CSoutput.n321 103.111
R22360 CSoutput.n320 CSoutput.n319 103.111
R22361 CSoutput.n318 CSoutput.n317 103.111
R22362 CSoutput.n316 CSoutput.n315 103.111
R22363 CSoutput.n314 CSoutput.n313 103.111
R22364 CSoutput.n312 CSoutput.n311 103.111
R22365 CSoutput.n310 CSoutput.n309 103.111
R22366 CSoutput.n307 CSoutput.n306 103.111
R22367 CSoutput.n305 CSoutput.n304 103.111
R22368 CSoutput.n303 CSoutput.n302 103.111
R22369 CSoutput.n301 CSoutput.n300 103.111
R22370 CSoutput.n299 CSoutput.n298 103.111
R22371 CSoutput.n297 CSoutput.n296 103.111
R22372 CSoutput.n295 CSoutput.n294 103.111
R22373 CSoutput.n293 CSoutput.n292 103.111
R22374 CSoutput.n291 CSoutput.n290 103.111
R22375 CSoutput.n120 CSoutput.n119 103.111
R22376 CSoutput.n122 CSoutput.n121 103.111
R22377 CSoutput.n124 CSoutput.n123 103.111
R22378 CSoutput.n126 CSoutput.n125 103.111
R22379 CSoutput.n128 CSoutput.n127 103.111
R22380 CSoutput.n130 CSoutput.n129 103.111
R22381 CSoutput.n132 CSoutput.n131 103.111
R22382 CSoutput.n134 CSoutput.n133 103.111
R22383 CSoutput.n136 CSoutput.n135 103.111
R22384 CSoutput.n100 CSoutput.n99 103.111
R22385 CSoutput.n102 CSoutput.n101 103.111
R22386 CSoutput.n104 CSoutput.n103 103.111
R22387 CSoutput.n106 CSoutput.n105 103.111
R22388 CSoutput.n108 CSoutput.n107 103.111
R22389 CSoutput.n110 CSoutput.n109 103.111
R22390 CSoutput.n112 CSoutput.n111 103.111
R22391 CSoutput.n114 CSoutput.n113 103.111
R22392 CSoutput.n116 CSoutput.n115 103.111
R22393 CSoutput.n81 CSoutput.n80 103.111
R22394 CSoutput.n83 CSoutput.n82 103.111
R22395 CSoutput.n85 CSoutput.n84 103.111
R22396 CSoutput.n87 CSoutput.n86 103.111
R22397 CSoutput.n89 CSoutput.n88 103.111
R22398 CSoutput.n91 CSoutput.n90 103.111
R22399 CSoutput.n93 CSoutput.n92 103.111
R22400 CSoutput.n95 CSoutput.n94 103.111
R22401 CSoutput.n97 CSoutput.n96 103.111
R22402 CSoutput.n346 CSoutput.n345 103.111
R22403 CSoutput.n370 CSoutput.n368 81.5057
R22404 CSoutput.n351 CSoutput.n349 81.5057
R22405 CSoutput.n410 CSoutput.n408 81.5057
R22406 CSoutput.n391 CSoutput.n389 81.5057
R22407 CSoutput.n386 CSoutput.n385 80.9324
R22408 CSoutput.n384 CSoutput.n383 80.9324
R22409 CSoutput.n382 CSoutput.n381 80.9324
R22410 CSoutput.n380 CSoutput.n379 80.9324
R22411 CSoutput.n378 CSoutput.n377 80.9324
R22412 CSoutput.n376 CSoutput.n375 80.9324
R22413 CSoutput.n374 CSoutput.n373 80.9324
R22414 CSoutput.n372 CSoutput.n371 80.9324
R22415 CSoutput.n370 CSoutput.n369 80.9324
R22416 CSoutput.n367 CSoutput.n366 80.9324
R22417 CSoutput.n365 CSoutput.n364 80.9324
R22418 CSoutput.n363 CSoutput.n362 80.9324
R22419 CSoutput.n361 CSoutput.n360 80.9324
R22420 CSoutput.n359 CSoutput.n358 80.9324
R22421 CSoutput.n357 CSoutput.n356 80.9324
R22422 CSoutput.n355 CSoutput.n354 80.9324
R22423 CSoutput.n353 CSoutput.n352 80.9324
R22424 CSoutput.n351 CSoutput.n350 80.9324
R22425 CSoutput.n410 CSoutput.n409 80.9324
R22426 CSoutput.n412 CSoutput.n411 80.9324
R22427 CSoutput.n414 CSoutput.n413 80.9324
R22428 CSoutput.n416 CSoutput.n415 80.9324
R22429 CSoutput.n418 CSoutput.n417 80.9324
R22430 CSoutput.n420 CSoutput.n419 80.9324
R22431 CSoutput.n422 CSoutput.n421 80.9324
R22432 CSoutput.n424 CSoutput.n423 80.9324
R22433 CSoutput.n426 CSoutput.n425 80.9324
R22434 CSoutput.n391 CSoutput.n390 80.9324
R22435 CSoutput.n393 CSoutput.n392 80.9324
R22436 CSoutput.n395 CSoutput.n394 80.9324
R22437 CSoutput.n397 CSoutput.n396 80.9324
R22438 CSoutput.n399 CSoutput.n398 80.9324
R22439 CSoutput.n401 CSoutput.n400 80.9324
R22440 CSoutput.n403 CSoutput.n402 80.9324
R22441 CSoutput.n405 CSoutput.n404 80.9324
R22442 CSoutput.n407 CSoutput.n406 80.9324
R22443 CSoutput.n25 CSoutput.n24 48.1486
R22444 CSoutput.n69 CSoutput.n3 48.1486
R22445 CSoutput.n38 CSoutput.n37 48.1486
R22446 CSoutput.n42 CSoutput.n41 48.1486
R22447 CSoutput.n51 CSoutput.n50 48.1486
R22448 CSoutput.n55 CSoutput.n54 48.1486
R22449 CSoutput.n22 CSoutput.n17 46.462
R22450 CSoutput.n72 CSoutput.n71 46.462
R22451 CSoutput.n20 CSoutput.n19 44.9055
R22452 CSoutput.n29 CSoutput.n28 43.7635
R22453 CSoutput.n65 CSoutput.n63 43.7635
R22454 CSoutput.n35 CSoutput.n13 41.7396
R22455 CSoutput.n57 CSoutput.n5 41.7396
R22456 CSoutput.n44 CSoutput.n9 37.0171
R22457 CSoutput.n48 CSoutput.n9 37.0171
R22458 CSoutput.n76 CSoutput.n75 34.9932
R22459 CSoutput.n31 CSoutput.n13 32.2947
R22460 CSoutput.n61 CSoutput.n5 32.2947
R22461 CSoutput.n30 CSoutput.n29 29.6014
R22462 CSoutput.n63 CSoutput.n62 29.6014
R22463 CSoutput.n19 CSoutput.n18 28.4085
R22464 CSoutput.n18 CSoutput.n17 25.1176
R22465 CSoutput.n72 CSoutput.n1 25.1176
R22466 CSoutput.n43 CSoutput.n42 22.0922
R22467 CSoutput.n50 CSoutput.n49 22.0922
R22468 CSoutput.n77 CSoutput.n76 21.8586
R22469 CSoutput.n37 CSoutput.n36 18.9681
R22470 CSoutput.n56 CSoutput.n55 18.9681
R22471 CSoutput.n25 CSoutput.n15 17.6292
R22472 CSoutput.n64 CSoutput.n3 17.6292
R22473 CSoutput.n24 CSoutput.n23 15.844
R22474 CSoutput.n70 CSoutput.n69 15.844
R22475 CSoutput.n38 CSoutput.n11 14.5051
R22476 CSoutput.n54 CSoutput.n7 14.5051
R22477 CSoutput.n429 CSoutput.n78 11.6139
R22478 CSoutput.n41 CSoutput.n11 11.3811
R22479 CSoutput.n51 CSoutput.n7 11.3811
R22480 CSoutput.n23 CSoutput.n22 10.0422
R22481 CSoutput.n71 CSoutput.n70 10.0422
R22482 CSoutput.n327 CSoutput.n307 9.25285
R22483 CSoutput.n117 CSoutput.n97 9.25285
R22484 CSoutput.n387 CSoutput.n367 8.97993
R22485 CSoutput.n427 CSoutput.n407 8.97993
R22486 CSoutput.n388 CSoutput.n348 8.78259
R22487 CSoutput.n28 CSoutput.n15 8.25698
R22488 CSoutput.n65 CSoutput.n64 8.25698
R22489 CSoutput.n388 CSoutput.n387 7.89345
R22490 CSoutput.n428 CSoutput.n427 7.89345
R22491 CSoutput.n348 CSoutput.n347 7.12641
R22492 CSoutput.n138 CSoutput.n137 7.12641
R22493 CSoutput.n36 CSoutput.n35 6.91809
R22494 CSoutput.n57 CSoutput.n56 6.91809
R22495 CSoutput.n387 CSoutput.n386 5.25266
R22496 CSoutput.n427 CSoutput.n426 5.25266
R22497 CSoutput.n429 CSoutput.n138 5.19015
R22498 CSoutput.n347 CSoutput.n346 5.1449
R22499 CSoutput.n327 CSoutput.n326 5.1449
R22500 CSoutput.n137 CSoutput.n136 5.1449
R22501 CSoutput.n117 CSoutput.n116 5.1449
R22502 CSoutput.n229 CSoutput.n182 4.5005
R22503 CSoutput.n198 CSoutput.n182 4.5005
R22504 CSoutput.n193 CSoutput.n177 4.5005
R22505 CSoutput.n193 CSoutput.n179 4.5005
R22506 CSoutput.n193 CSoutput.n176 4.5005
R22507 CSoutput.n193 CSoutput.n180 4.5005
R22508 CSoutput.n193 CSoutput.n175 4.5005
R22509 CSoutput.n193 CSoutput.t208 4.5005
R22510 CSoutput.n193 CSoutput.n174 4.5005
R22511 CSoutput.n193 CSoutput.n181 4.5005
R22512 CSoutput.n193 CSoutput.n182 4.5005
R22513 CSoutput.n191 CSoutput.n177 4.5005
R22514 CSoutput.n191 CSoutput.n179 4.5005
R22515 CSoutput.n191 CSoutput.n176 4.5005
R22516 CSoutput.n191 CSoutput.n180 4.5005
R22517 CSoutput.n191 CSoutput.n175 4.5005
R22518 CSoutput.n191 CSoutput.t208 4.5005
R22519 CSoutput.n191 CSoutput.n174 4.5005
R22520 CSoutput.n191 CSoutput.n181 4.5005
R22521 CSoutput.n191 CSoutput.n182 4.5005
R22522 CSoutput.n190 CSoutput.n177 4.5005
R22523 CSoutput.n190 CSoutput.n179 4.5005
R22524 CSoutput.n190 CSoutput.n176 4.5005
R22525 CSoutput.n190 CSoutput.n180 4.5005
R22526 CSoutput.n190 CSoutput.n175 4.5005
R22527 CSoutput.n190 CSoutput.t208 4.5005
R22528 CSoutput.n190 CSoutput.n174 4.5005
R22529 CSoutput.n190 CSoutput.n181 4.5005
R22530 CSoutput.n190 CSoutput.n182 4.5005
R22531 CSoutput.n275 CSoutput.n177 4.5005
R22532 CSoutput.n275 CSoutput.n179 4.5005
R22533 CSoutput.n275 CSoutput.n176 4.5005
R22534 CSoutput.n275 CSoutput.n180 4.5005
R22535 CSoutput.n275 CSoutput.n175 4.5005
R22536 CSoutput.n275 CSoutput.t208 4.5005
R22537 CSoutput.n275 CSoutput.n174 4.5005
R22538 CSoutput.n275 CSoutput.n181 4.5005
R22539 CSoutput.n275 CSoutput.n182 4.5005
R22540 CSoutput.n273 CSoutput.n177 4.5005
R22541 CSoutput.n273 CSoutput.n179 4.5005
R22542 CSoutput.n273 CSoutput.n176 4.5005
R22543 CSoutput.n273 CSoutput.n180 4.5005
R22544 CSoutput.n273 CSoutput.n175 4.5005
R22545 CSoutput.n273 CSoutput.t208 4.5005
R22546 CSoutput.n273 CSoutput.n174 4.5005
R22547 CSoutput.n273 CSoutput.n181 4.5005
R22548 CSoutput.n271 CSoutput.n177 4.5005
R22549 CSoutput.n271 CSoutput.n179 4.5005
R22550 CSoutput.n271 CSoutput.n176 4.5005
R22551 CSoutput.n271 CSoutput.n180 4.5005
R22552 CSoutput.n271 CSoutput.n175 4.5005
R22553 CSoutput.n271 CSoutput.t208 4.5005
R22554 CSoutput.n271 CSoutput.n174 4.5005
R22555 CSoutput.n271 CSoutput.n181 4.5005
R22556 CSoutput.n201 CSoutput.n177 4.5005
R22557 CSoutput.n201 CSoutput.n179 4.5005
R22558 CSoutput.n201 CSoutput.n176 4.5005
R22559 CSoutput.n201 CSoutput.n180 4.5005
R22560 CSoutput.n201 CSoutput.n175 4.5005
R22561 CSoutput.n201 CSoutput.t208 4.5005
R22562 CSoutput.n201 CSoutput.n174 4.5005
R22563 CSoutput.n201 CSoutput.n181 4.5005
R22564 CSoutput.n201 CSoutput.n182 4.5005
R22565 CSoutput.n200 CSoutput.n177 4.5005
R22566 CSoutput.n200 CSoutput.n179 4.5005
R22567 CSoutput.n200 CSoutput.n176 4.5005
R22568 CSoutput.n200 CSoutput.n180 4.5005
R22569 CSoutput.n200 CSoutput.n175 4.5005
R22570 CSoutput.n200 CSoutput.t208 4.5005
R22571 CSoutput.n200 CSoutput.n174 4.5005
R22572 CSoutput.n200 CSoutput.n181 4.5005
R22573 CSoutput.n200 CSoutput.n182 4.5005
R22574 CSoutput.n204 CSoutput.n177 4.5005
R22575 CSoutput.n204 CSoutput.n179 4.5005
R22576 CSoutput.n204 CSoutput.n176 4.5005
R22577 CSoutput.n204 CSoutput.n180 4.5005
R22578 CSoutput.n204 CSoutput.n175 4.5005
R22579 CSoutput.n204 CSoutput.t208 4.5005
R22580 CSoutput.n204 CSoutput.n174 4.5005
R22581 CSoutput.n204 CSoutput.n181 4.5005
R22582 CSoutput.n204 CSoutput.n182 4.5005
R22583 CSoutput.n203 CSoutput.n177 4.5005
R22584 CSoutput.n203 CSoutput.n179 4.5005
R22585 CSoutput.n203 CSoutput.n176 4.5005
R22586 CSoutput.n203 CSoutput.n180 4.5005
R22587 CSoutput.n203 CSoutput.n175 4.5005
R22588 CSoutput.n203 CSoutput.t208 4.5005
R22589 CSoutput.n203 CSoutput.n174 4.5005
R22590 CSoutput.n203 CSoutput.n181 4.5005
R22591 CSoutput.n203 CSoutput.n182 4.5005
R22592 CSoutput.n186 CSoutput.n177 4.5005
R22593 CSoutput.n186 CSoutput.n179 4.5005
R22594 CSoutput.n186 CSoutput.n176 4.5005
R22595 CSoutput.n186 CSoutput.n180 4.5005
R22596 CSoutput.n186 CSoutput.n175 4.5005
R22597 CSoutput.n186 CSoutput.t208 4.5005
R22598 CSoutput.n186 CSoutput.n174 4.5005
R22599 CSoutput.n186 CSoutput.n181 4.5005
R22600 CSoutput.n186 CSoutput.n182 4.5005
R22601 CSoutput.n278 CSoutput.n177 4.5005
R22602 CSoutput.n278 CSoutput.n179 4.5005
R22603 CSoutput.n278 CSoutput.n176 4.5005
R22604 CSoutput.n278 CSoutput.n180 4.5005
R22605 CSoutput.n278 CSoutput.n175 4.5005
R22606 CSoutput.n278 CSoutput.t208 4.5005
R22607 CSoutput.n278 CSoutput.n174 4.5005
R22608 CSoutput.n278 CSoutput.n181 4.5005
R22609 CSoutput.n278 CSoutput.n182 4.5005
R22610 CSoutput.n265 CSoutput.n236 4.5005
R22611 CSoutput.n265 CSoutput.n242 4.5005
R22612 CSoutput.n223 CSoutput.n212 4.5005
R22613 CSoutput.n223 CSoutput.n214 4.5005
R22614 CSoutput.n223 CSoutput.n211 4.5005
R22615 CSoutput.n223 CSoutput.n215 4.5005
R22616 CSoutput.n223 CSoutput.n210 4.5005
R22617 CSoutput.n223 CSoutput.t210 4.5005
R22618 CSoutput.n223 CSoutput.n209 4.5005
R22619 CSoutput.n223 CSoutput.n216 4.5005
R22620 CSoutput.n265 CSoutput.n223 4.5005
R22621 CSoutput.n244 CSoutput.n212 4.5005
R22622 CSoutput.n244 CSoutput.n214 4.5005
R22623 CSoutput.n244 CSoutput.n211 4.5005
R22624 CSoutput.n244 CSoutput.n215 4.5005
R22625 CSoutput.n244 CSoutput.n210 4.5005
R22626 CSoutput.n244 CSoutput.t210 4.5005
R22627 CSoutput.n244 CSoutput.n209 4.5005
R22628 CSoutput.n244 CSoutput.n216 4.5005
R22629 CSoutput.n265 CSoutput.n244 4.5005
R22630 CSoutput.n222 CSoutput.n212 4.5005
R22631 CSoutput.n222 CSoutput.n214 4.5005
R22632 CSoutput.n222 CSoutput.n211 4.5005
R22633 CSoutput.n222 CSoutput.n215 4.5005
R22634 CSoutput.n222 CSoutput.n210 4.5005
R22635 CSoutput.n222 CSoutput.t210 4.5005
R22636 CSoutput.n222 CSoutput.n209 4.5005
R22637 CSoutput.n222 CSoutput.n216 4.5005
R22638 CSoutput.n265 CSoutput.n222 4.5005
R22639 CSoutput.n246 CSoutput.n212 4.5005
R22640 CSoutput.n246 CSoutput.n214 4.5005
R22641 CSoutput.n246 CSoutput.n211 4.5005
R22642 CSoutput.n246 CSoutput.n215 4.5005
R22643 CSoutput.n246 CSoutput.n210 4.5005
R22644 CSoutput.n246 CSoutput.t210 4.5005
R22645 CSoutput.n246 CSoutput.n209 4.5005
R22646 CSoutput.n246 CSoutput.n216 4.5005
R22647 CSoutput.n265 CSoutput.n246 4.5005
R22648 CSoutput.n212 CSoutput.n207 4.5005
R22649 CSoutput.n214 CSoutput.n207 4.5005
R22650 CSoutput.n211 CSoutput.n207 4.5005
R22651 CSoutput.n215 CSoutput.n207 4.5005
R22652 CSoutput.n210 CSoutput.n207 4.5005
R22653 CSoutput.t210 CSoutput.n207 4.5005
R22654 CSoutput.n209 CSoutput.n207 4.5005
R22655 CSoutput.n216 CSoutput.n207 4.5005
R22656 CSoutput.n268 CSoutput.n212 4.5005
R22657 CSoutput.n268 CSoutput.n214 4.5005
R22658 CSoutput.n268 CSoutput.n211 4.5005
R22659 CSoutput.n268 CSoutput.n215 4.5005
R22660 CSoutput.n268 CSoutput.n210 4.5005
R22661 CSoutput.n268 CSoutput.t210 4.5005
R22662 CSoutput.n268 CSoutput.n209 4.5005
R22663 CSoutput.n268 CSoutput.n216 4.5005
R22664 CSoutput.n266 CSoutput.n212 4.5005
R22665 CSoutput.n266 CSoutput.n214 4.5005
R22666 CSoutput.n266 CSoutput.n211 4.5005
R22667 CSoutput.n266 CSoutput.n215 4.5005
R22668 CSoutput.n266 CSoutput.n210 4.5005
R22669 CSoutput.n266 CSoutput.t210 4.5005
R22670 CSoutput.n266 CSoutput.n209 4.5005
R22671 CSoutput.n266 CSoutput.n216 4.5005
R22672 CSoutput.n266 CSoutput.n265 4.5005
R22673 CSoutput.n248 CSoutput.n212 4.5005
R22674 CSoutput.n248 CSoutput.n214 4.5005
R22675 CSoutput.n248 CSoutput.n211 4.5005
R22676 CSoutput.n248 CSoutput.n215 4.5005
R22677 CSoutput.n248 CSoutput.n210 4.5005
R22678 CSoutput.n248 CSoutput.t210 4.5005
R22679 CSoutput.n248 CSoutput.n209 4.5005
R22680 CSoutput.n248 CSoutput.n216 4.5005
R22681 CSoutput.n265 CSoutput.n248 4.5005
R22682 CSoutput.n220 CSoutput.n212 4.5005
R22683 CSoutput.n220 CSoutput.n214 4.5005
R22684 CSoutput.n220 CSoutput.n211 4.5005
R22685 CSoutput.n220 CSoutput.n215 4.5005
R22686 CSoutput.n220 CSoutput.n210 4.5005
R22687 CSoutput.n220 CSoutput.t210 4.5005
R22688 CSoutput.n220 CSoutput.n209 4.5005
R22689 CSoutput.n220 CSoutput.n216 4.5005
R22690 CSoutput.n265 CSoutput.n220 4.5005
R22691 CSoutput.n250 CSoutput.n212 4.5005
R22692 CSoutput.n250 CSoutput.n214 4.5005
R22693 CSoutput.n250 CSoutput.n211 4.5005
R22694 CSoutput.n250 CSoutput.n215 4.5005
R22695 CSoutput.n250 CSoutput.n210 4.5005
R22696 CSoutput.n250 CSoutput.t210 4.5005
R22697 CSoutput.n250 CSoutput.n209 4.5005
R22698 CSoutput.n250 CSoutput.n216 4.5005
R22699 CSoutput.n265 CSoutput.n250 4.5005
R22700 CSoutput.n219 CSoutput.n212 4.5005
R22701 CSoutput.n219 CSoutput.n214 4.5005
R22702 CSoutput.n219 CSoutput.n211 4.5005
R22703 CSoutput.n219 CSoutput.n215 4.5005
R22704 CSoutput.n219 CSoutput.n210 4.5005
R22705 CSoutput.n219 CSoutput.t210 4.5005
R22706 CSoutput.n219 CSoutput.n209 4.5005
R22707 CSoutput.n219 CSoutput.n216 4.5005
R22708 CSoutput.n265 CSoutput.n219 4.5005
R22709 CSoutput.n264 CSoutput.n212 4.5005
R22710 CSoutput.n264 CSoutput.n214 4.5005
R22711 CSoutput.n264 CSoutput.n211 4.5005
R22712 CSoutput.n264 CSoutput.n215 4.5005
R22713 CSoutput.n264 CSoutput.n210 4.5005
R22714 CSoutput.n264 CSoutput.t210 4.5005
R22715 CSoutput.n264 CSoutput.n209 4.5005
R22716 CSoutput.n264 CSoutput.n216 4.5005
R22717 CSoutput.n265 CSoutput.n264 4.5005
R22718 CSoutput.n263 CSoutput.n148 4.5005
R22719 CSoutput.n164 CSoutput.n148 4.5005
R22720 CSoutput.n159 CSoutput.n143 4.5005
R22721 CSoutput.n159 CSoutput.n145 4.5005
R22722 CSoutput.n159 CSoutput.n142 4.5005
R22723 CSoutput.n159 CSoutput.n146 4.5005
R22724 CSoutput.n159 CSoutput.n141 4.5005
R22725 CSoutput.n159 CSoutput.t211 4.5005
R22726 CSoutput.n159 CSoutput.n140 4.5005
R22727 CSoutput.n159 CSoutput.n147 4.5005
R22728 CSoutput.n159 CSoutput.n148 4.5005
R22729 CSoutput.n157 CSoutput.n143 4.5005
R22730 CSoutput.n157 CSoutput.n145 4.5005
R22731 CSoutput.n157 CSoutput.n142 4.5005
R22732 CSoutput.n157 CSoutput.n146 4.5005
R22733 CSoutput.n157 CSoutput.n141 4.5005
R22734 CSoutput.n157 CSoutput.t211 4.5005
R22735 CSoutput.n157 CSoutput.n140 4.5005
R22736 CSoutput.n157 CSoutput.n147 4.5005
R22737 CSoutput.n157 CSoutput.n148 4.5005
R22738 CSoutput.n156 CSoutput.n143 4.5005
R22739 CSoutput.n156 CSoutput.n145 4.5005
R22740 CSoutput.n156 CSoutput.n142 4.5005
R22741 CSoutput.n156 CSoutput.n146 4.5005
R22742 CSoutput.n156 CSoutput.n141 4.5005
R22743 CSoutput.n156 CSoutput.t211 4.5005
R22744 CSoutput.n156 CSoutput.n140 4.5005
R22745 CSoutput.n156 CSoutput.n147 4.5005
R22746 CSoutput.n156 CSoutput.n148 4.5005
R22747 CSoutput.n285 CSoutput.n143 4.5005
R22748 CSoutput.n285 CSoutput.n145 4.5005
R22749 CSoutput.n285 CSoutput.n142 4.5005
R22750 CSoutput.n285 CSoutput.n146 4.5005
R22751 CSoutput.n285 CSoutput.n141 4.5005
R22752 CSoutput.n285 CSoutput.t211 4.5005
R22753 CSoutput.n285 CSoutput.n140 4.5005
R22754 CSoutput.n285 CSoutput.n147 4.5005
R22755 CSoutput.n285 CSoutput.n148 4.5005
R22756 CSoutput.n283 CSoutput.n143 4.5005
R22757 CSoutput.n283 CSoutput.n145 4.5005
R22758 CSoutput.n283 CSoutput.n142 4.5005
R22759 CSoutput.n283 CSoutput.n146 4.5005
R22760 CSoutput.n283 CSoutput.n141 4.5005
R22761 CSoutput.n283 CSoutput.t211 4.5005
R22762 CSoutput.n283 CSoutput.n140 4.5005
R22763 CSoutput.n283 CSoutput.n147 4.5005
R22764 CSoutput.n281 CSoutput.n143 4.5005
R22765 CSoutput.n281 CSoutput.n145 4.5005
R22766 CSoutput.n281 CSoutput.n142 4.5005
R22767 CSoutput.n281 CSoutput.n146 4.5005
R22768 CSoutput.n281 CSoutput.n141 4.5005
R22769 CSoutput.n281 CSoutput.t211 4.5005
R22770 CSoutput.n281 CSoutput.n140 4.5005
R22771 CSoutput.n281 CSoutput.n147 4.5005
R22772 CSoutput.n167 CSoutput.n143 4.5005
R22773 CSoutput.n167 CSoutput.n145 4.5005
R22774 CSoutput.n167 CSoutput.n142 4.5005
R22775 CSoutput.n167 CSoutput.n146 4.5005
R22776 CSoutput.n167 CSoutput.n141 4.5005
R22777 CSoutput.n167 CSoutput.t211 4.5005
R22778 CSoutput.n167 CSoutput.n140 4.5005
R22779 CSoutput.n167 CSoutput.n147 4.5005
R22780 CSoutput.n167 CSoutput.n148 4.5005
R22781 CSoutput.n166 CSoutput.n143 4.5005
R22782 CSoutput.n166 CSoutput.n145 4.5005
R22783 CSoutput.n166 CSoutput.n142 4.5005
R22784 CSoutput.n166 CSoutput.n146 4.5005
R22785 CSoutput.n166 CSoutput.n141 4.5005
R22786 CSoutput.n166 CSoutput.t211 4.5005
R22787 CSoutput.n166 CSoutput.n140 4.5005
R22788 CSoutput.n166 CSoutput.n147 4.5005
R22789 CSoutput.n166 CSoutput.n148 4.5005
R22790 CSoutput.n170 CSoutput.n143 4.5005
R22791 CSoutput.n170 CSoutput.n145 4.5005
R22792 CSoutput.n170 CSoutput.n142 4.5005
R22793 CSoutput.n170 CSoutput.n146 4.5005
R22794 CSoutput.n170 CSoutput.n141 4.5005
R22795 CSoutput.n170 CSoutput.t211 4.5005
R22796 CSoutput.n170 CSoutput.n140 4.5005
R22797 CSoutput.n170 CSoutput.n147 4.5005
R22798 CSoutput.n170 CSoutput.n148 4.5005
R22799 CSoutput.n169 CSoutput.n143 4.5005
R22800 CSoutput.n169 CSoutput.n145 4.5005
R22801 CSoutput.n169 CSoutput.n142 4.5005
R22802 CSoutput.n169 CSoutput.n146 4.5005
R22803 CSoutput.n169 CSoutput.n141 4.5005
R22804 CSoutput.n169 CSoutput.t211 4.5005
R22805 CSoutput.n169 CSoutput.n140 4.5005
R22806 CSoutput.n169 CSoutput.n147 4.5005
R22807 CSoutput.n169 CSoutput.n148 4.5005
R22808 CSoutput.n152 CSoutput.n143 4.5005
R22809 CSoutput.n152 CSoutput.n145 4.5005
R22810 CSoutput.n152 CSoutput.n142 4.5005
R22811 CSoutput.n152 CSoutput.n146 4.5005
R22812 CSoutput.n152 CSoutput.n141 4.5005
R22813 CSoutput.n152 CSoutput.t211 4.5005
R22814 CSoutput.n152 CSoutput.n140 4.5005
R22815 CSoutput.n152 CSoutput.n147 4.5005
R22816 CSoutput.n152 CSoutput.n148 4.5005
R22817 CSoutput.n288 CSoutput.n143 4.5005
R22818 CSoutput.n288 CSoutput.n145 4.5005
R22819 CSoutput.n288 CSoutput.n142 4.5005
R22820 CSoutput.n288 CSoutput.n146 4.5005
R22821 CSoutput.n288 CSoutput.n141 4.5005
R22822 CSoutput.n288 CSoutput.t211 4.5005
R22823 CSoutput.n288 CSoutput.n140 4.5005
R22824 CSoutput.n288 CSoutput.n147 4.5005
R22825 CSoutput.n288 CSoutput.n148 4.5005
R22826 CSoutput.n347 CSoutput.n327 4.10845
R22827 CSoutput.n137 CSoutput.n117 4.10845
R22828 CSoutput.n345 CSoutput.t67 4.06363
R22829 CSoutput.n345 CSoutput.t71 4.06363
R22830 CSoutput.n343 CSoutput.t93 4.06363
R22831 CSoutput.n343 CSoutput.t157 4.06363
R22832 CSoutput.n341 CSoutput.t162 4.06363
R22833 CSoutput.n341 CSoutput.t74 4.06363
R22834 CSoutput.n339 CSoutput.t95 4.06363
R22835 CSoutput.n339 CSoutput.t123 4.06363
R22836 CSoutput.n337 CSoutput.t137 4.06363
R22837 CSoutput.n337 CSoutput.t58 4.06363
R22838 CSoutput.n335 CSoutput.t52 4.06363
R22839 CSoutput.n335 CSoutput.t97 4.06363
R22840 CSoutput.n333 CSoutput.t115 4.06363
R22841 CSoutput.n333 CSoutput.t140 4.06363
R22842 CSoutput.n331 CSoutput.t158 4.06363
R22843 CSoutput.n331 CSoutput.t70 4.06363
R22844 CSoutput.n329 CSoutput.t77 4.06363
R22845 CSoutput.n329 CSoutput.t141 4.06363
R22846 CSoutput.n328 CSoutput.t161 4.06363
R22847 CSoutput.n328 CSoutput.t163 4.06363
R22848 CSoutput.n325 CSoutput.t55 4.06363
R22849 CSoutput.n325 CSoutput.t56 4.06363
R22850 CSoutput.n323 CSoutput.t78 4.06363
R22851 CSoutput.n323 CSoutput.t142 4.06363
R22852 CSoutput.n321 CSoutput.t149 4.06363
R22853 CSoutput.n321 CSoutput.t59 4.06363
R22854 CSoutput.n319 CSoutput.t79 4.06363
R22855 CSoutput.n319 CSoutput.t113 4.06363
R22856 CSoutput.n317 CSoutput.t128 4.06363
R22857 CSoutput.n317 CSoutput.t167 4.06363
R22858 CSoutput.n315 CSoutput.t159 4.06363
R22859 CSoutput.n315 CSoutput.t84 4.06363
R22860 CSoutput.n313 CSoutput.t101 4.06363
R22861 CSoutput.n313 CSoutput.t129 4.06363
R22862 CSoutput.n311 CSoutput.t143 4.06363
R22863 CSoutput.n311 CSoutput.t57 4.06363
R22864 CSoutput.n309 CSoutput.t60 4.06363
R22865 CSoutput.n309 CSoutput.t132 4.06363
R22866 CSoutput.n308 CSoutput.t150 4.06363
R22867 CSoutput.n308 CSoutput.t151 4.06363
R22868 CSoutput.n306 CSoutput.t154 4.06363
R22869 CSoutput.n306 CSoutput.t133 4.06363
R22870 CSoutput.n304 CSoutput.t50 4.06363
R22871 CSoutput.n304 CSoutput.t91 4.06363
R22872 CSoutput.n302 CSoutput.t164 4.06363
R22873 CSoutput.n302 CSoutput.t114 4.06363
R22874 CSoutput.n300 CSoutput.t146 4.06363
R22875 CSoutput.n300 CSoutput.t98 4.06363
R22876 CSoutput.n298 CSoutput.t130 4.06363
R22877 CSoutput.n298 CSoutput.t82 4.06363
R22878 CSoutput.n296 CSoutput.t153 4.06363
R22879 CSoutput.n296 CSoutput.t107 4.06363
R22880 CSoutput.n294 CSoutput.t138 4.06363
R22881 CSoutput.n294 CSoutput.t90 4.06363
R22882 CSoutput.n292 CSoutput.t125 4.06363
R22883 CSoutput.n292 CSoutput.t69 4.06363
R22884 CSoutput.n290 CSoutput.t144 4.06363
R22885 CSoutput.n290 CSoutput.t62 4.06363
R22886 CSoutput.n289 CSoutput.t102 4.06363
R22887 CSoutput.n289 CSoutput.t80 4.06363
R22888 CSoutput.n118 CSoutput.t121 4.06363
R22889 CSoutput.n118 CSoutput.t89 4.06363
R22890 CSoutput.n119 CSoutput.t66 4.06363
R22891 CSoutput.n119 CSoutput.t122 4.06363
R22892 CSoutput.n121 CSoutput.t118 4.06363
R22893 CSoutput.n121 CSoutput.t86 4.06363
R22894 CSoutput.n123 CSoutput.t65 4.06363
R22895 CSoutput.n123 CSoutput.t64 4.06363
R22896 CSoutput.n125 CSoutput.t136 4.06363
R22897 CSoutput.n125 CSoutput.t100 4.06363
R22898 CSoutput.n127 CSoutput.t96 4.06363
R22899 CSoutput.n127 CSoutput.t61 4.06363
R22900 CSoutput.n129 CSoutput.t166 4.06363
R22901 CSoutput.n129 CSoutput.t134 4.06363
R22902 CSoutput.n131 CSoutput.t120 4.06363
R22903 CSoutput.n131 CSoutput.t88 4.06363
R22904 CSoutput.n133 CSoutput.t85 4.06363
R22905 CSoutput.n133 CSoutput.t160 4.06363
R22906 CSoutput.n135 CSoutput.t119 4.06363
R22907 CSoutput.n135 CSoutput.t117 4.06363
R22908 CSoutput.n98 CSoutput.t109 4.06363
R22909 CSoutput.n98 CSoutput.t75 4.06363
R22910 CSoutput.n99 CSoutput.t54 4.06363
R22911 CSoutput.n99 CSoutput.t111 4.06363
R22912 CSoutput.n101 CSoutput.t105 4.06363
R22913 CSoutput.n101 CSoutput.t72 4.06363
R22914 CSoutput.n103 CSoutput.t53 4.06363
R22915 CSoutput.n103 CSoutput.t51 4.06363
R22916 CSoutput.n105 CSoutput.t127 4.06363
R22917 CSoutput.n105 CSoutput.t87 4.06363
R22918 CSoutput.n107 CSoutput.t83 4.06363
R22919 CSoutput.n107 CSoutput.t49 4.06363
R22920 CSoutput.n109 CSoutput.t152 4.06363
R22921 CSoutput.n109 CSoutput.t124 4.06363
R22922 CSoutput.n111 CSoutput.t110 4.06363
R22923 CSoutput.n111 CSoutput.t76 4.06363
R22924 CSoutput.n113 CSoutput.t68 4.06363
R22925 CSoutput.n113 CSoutput.t148 4.06363
R22926 CSoutput.n115 CSoutput.t106 4.06363
R22927 CSoutput.n115 CSoutput.t104 4.06363
R22928 CSoutput.n79 CSoutput.t168 4.06363
R22929 CSoutput.n79 CSoutput.t103 4.06363
R22930 CSoutput.n80 CSoutput.t63 4.06363
R22931 CSoutput.n80 CSoutput.t145 4.06363
R22932 CSoutput.n82 CSoutput.t73 4.06363
R22933 CSoutput.n82 CSoutput.t126 4.06363
R22934 CSoutput.n84 CSoutput.t92 4.06363
R22935 CSoutput.n84 CSoutput.t112 4.06363
R22936 CSoutput.n86 CSoutput.t108 4.06363
R22937 CSoutput.n86 CSoutput.t155 4.06363
R22938 CSoutput.n88 CSoutput.t81 4.06363
R22939 CSoutput.n88 CSoutput.t131 4.06363
R22940 CSoutput.n90 CSoutput.t99 4.06363
R22941 CSoutput.n90 CSoutput.t147 4.06363
R22942 CSoutput.n92 CSoutput.t116 4.06363
R22943 CSoutput.n92 CSoutput.t165 4.06363
R22944 CSoutput.n94 CSoutput.t94 4.06363
R22945 CSoutput.n94 CSoutput.t139 4.06363
R22946 CSoutput.n96 CSoutput.t135 4.06363
R22947 CSoutput.n96 CSoutput.t156 4.06363
R22948 CSoutput.n44 CSoutput.n43 3.79402
R22949 CSoutput.n49 CSoutput.n48 3.79402
R22950 CSoutput.n428 CSoutput.n388 3.71319
R22951 CSoutput.n429 CSoutput.n428 3.57343
R22952 CSoutput.n348 CSoutput.n138 3.19963
R22953 CSoutput.n385 CSoutput.t172 2.82907
R22954 CSoutput.n385 CSoutput.t34 2.82907
R22955 CSoutput.n383 CSoutput.t180 2.82907
R22956 CSoutput.n383 CSoutput.t47 2.82907
R22957 CSoutput.n381 CSoutput.t174 2.82907
R22958 CSoutput.n381 CSoutput.t176 2.82907
R22959 CSoutput.n379 CSoutput.t31 2.82907
R22960 CSoutput.n379 CSoutput.t18 2.82907
R22961 CSoutput.n377 CSoutput.t20 2.82907
R22962 CSoutput.n377 CSoutput.t188 2.82907
R22963 CSoutput.n375 CSoutput.t182 2.82907
R22964 CSoutput.n375 CSoutput.t44 2.82907
R22965 CSoutput.n373 CSoutput.t171 2.82907
R22966 CSoutput.n373 CSoutput.t197 2.82907
R22967 CSoutput.n371 CSoutput.t189 2.82907
R22968 CSoutput.n371 CSoutput.t9 2.82907
R22969 CSoutput.n369 CSoutput.t170 2.82907
R22970 CSoutput.n369 CSoutput.t175 2.82907
R22971 CSoutput.n368 CSoutput.t33 2.82907
R22972 CSoutput.n368 CSoutput.t183 2.82907
R22973 CSoutput.n366 CSoutput.t36 2.82907
R22974 CSoutput.n366 CSoutput.t46 2.82907
R22975 CSoutput.n364 CSoutput.t14 2.82907
R22976 CSoutput.n364 CSoutput.t3 2.82907
R22977 CSoutput.n362 CSoutput.t186 2.82907
R22978 CSoutput.n362 CSoutput.t191 2.82907
R22979 CSoutput.n360 CSoutput.t17 2.82907
R22980 CSoutput.n360 CSoutput.t30 2.82907
R22981 CSoutput.n358 CSoutput.t24 2.82907
R22982 CSoutput.n358 CSoutput.t16 2.82907
R22983 CSoutput.n356 CSoutput.t195 2.82907
R22984 CSoutput.n356 CSoutput.t198 2.82907
R22985 CSoutput.n354 CSoutput.t35 2.82907
R22986 CSoutput.n354 CSoutput.t173 2.82907
R22987 CSoutput.n352 CSoutput.t10 2.82907
R22988 CSoutput.n352 CSoutput.t7 2.82907
R22989 CSoutput.n350 CSoutput.t0 2.82907
R22990 CSoutput.n350 CSoutput.t193 2.82907
R22991 CSoutput.n349 CSoutput.t185 2.82907
R22992 CSoutput.n349 CSoutput.t199 2.82907
R22993 CSoutput.n408 CSoutput.t23 2.82907
R22994 CSoutput.n408 CSoutput.t11 2.82907
R22995 CSoutput.n409 CSoutput.t181 2.82907
R22996 CSoutput.n409 CSoutput.t27 2.82907
R22997 CSoutput.n411 CSoutput.t1 2.82907
R22998 CSoutput.n411 CSoutput.t179 2.82907
R22999 CSoutput.n413 CSoutput.t38 2.82907
R23000 CSoutput.n413 CSoutput.t42 2.82907
R23001 CSoutput.n415 CSoutput.t21 2.82907
R23002 CSoutput.n415 CSoutput.t29 2.82907
R23003 CSoutput.n417 CSoutput.t43 2.82907
R23004 CSoutput.n417 CSoutput.t194 2.82907
R23005 CSoutput.n419 CSoutput.t22 2.82907
R23006 CSoutput.n419 CSoutput.t15 2.82907
R23007 CSoutput.n421 CSoutput.t37 2.82907
R23008 CSoutput.n421 CSoutput.t40 2.82907
R23009 CSoutput.n423 CSoutput.t177 2.82907
R23010 CSoutput.n423 CSoutput.t45 2.82907
R23011 CSoutput.n425 CSoutput.t190 2.82907
R23012 CSoutput.n425 CSoutput.t39 2.82907
R23013 CSoutput.n389 CSoutput.t28 2.82907
R23014 CSoutput.n389 CSoutput.t8 2.82907
R23015 CSoutput.n390 CSoutput.t48 2.82907
R23016 CSoutput.n390 CSoutput.t4 2.82907
R23017 CSoutput.n392 CSoutput.t41 2.82907
R23018 CSoutput.n392 CSoutput.t6 2.82907
R23019 CSoutput.n394 CSoutput.t187 2.82907
R23020 CSoutput.n394 CSoutput.t25 2.82907
R23021 CSoutput.n396 CSoutput.t5 2.82907
R23022 CSoutput.n396 CSoutput.t169 2.82907
R23023 CSoutput.n398 CSoutput.t13 2.82907
R23024 CSoutput.n398 CSoutput.t196 2.82907
R23025 CSoutput.n400 CSoutput.t26 2.82907
R23026 CSoutput.n400 CSoutput.t2 2.82907
R23027 CSoutput.n402 CSoutput.t184 2.82907
R23028 CSoutput.n402 CSoutput.t192 2.82907
R23029 CSoutput.n404 CSoutput.t19 2.82907
R23030 CSoutput.n404 CSoutput.t178 2.82907
R23031 CSoutput.n406 CSoutput.t12 2.82907
R23032 CSoutput.n406 CSoutput.t32 2.82907
R23033 CSoutput.n75 CSoutput.n1 2.45513
R23034 CSoutput.n229 CSoutput.n227 2.251
R23035 CSoutput.n229 CSoutput.n226 2.251
R23036 CSoutput.n229 CSoutput.n225 2.251
R23037 CSoutput.n229 CSoutput.n224 2.251
R23038 CSoutput.n198 CSoutput.n197 2.251
R23039 CSoutput.n198 CSoutput.n196 2.251
R23040 CSoutput.n198 CSoutput.n195 2.251
R23041 CSoutput.n198 CSoutput.n194 2.251
R23042 CSoutput.n271 CSoutput.n270 2.251
R23043 CSoutput.n236 CSoutput.n234 2.251
R23044 CSoutput.n236 CSoutput.n233 2.251
R23045 CSoutput.n236 CSoutput.n232 2.251
R23046 CSoutput.n254 CSoutput.n236 2.251
R23047 CSoutput.n242 CSoutput.n241 2.251
R23048 CSoutput.n242 CSoutput.n240 2.251
R23049 CSoutput.n242 CSoutput.n239 2.251
R23050 CSoutput.n242 CSoutput.n238 2.251
R23051 CSoutput.n268 CSoutput.n208 2.251
R23052 CSoutput.n263 CSoutput.n261 2.251
R23053 CSoutput.n263 CSoutput.n260 2.251
R23054 CSoutput.n263 CSoutput.n259 2.251
R23055 CSoutput.n263 CSoutput.n258 2.251
R23056 CSoutput.n164 CSoutput.n163 2.251
R23057 CSoutput.n164 CSoutput.n162 2.251
R23058 CSoutput.n164 CSoutput.n161 2.251
R23059 CSoutput.n164 CSoutput.n160 2.251
R23060 CSoutput.n281 CSoutput.n280 2.251
R23061 CSoutput.n198 CSoutput.n178 2.2505
R23062 CSoutput.n193 CSoutput.n178 2.2505
R23063 CSoutput.n191 CSoutput.n178 2.2505
R23064 CSoutput.n190 CSoutput.n178 2.2505
R23065 CSoutput.n275 CSoutput.n178 2.2505
R23066 CSoutput.n273 CSoutput.n178 2.2505
R23067 CSoutput.n271 CSoutput.n178 2.2505
R23068 CSoutput.n201 CSoutput.n178 2.2505
R23069 CSoutput.n200 CSoutput.n178 2.2505
R23070 CSoutput.n204 CSoutput.n178 2.2505
R23071 CSoutput.n203 CSoutput.n178 2.2505
R23072 CSoutput.n186 CSoutput.n178 2.2505
R23073 CSoutput.n278 CSoutput.n178 2.2505
R23074 CSoutput.n278 CSoutput.n277 2.2505
R23075 CSoutput.n242 CSoutput.n213 2.2505
R23076 CSoutput.n223 CSoutput.n213 2.2505
R23077 CSoutput.n244 CSoutput.n213 2.2505
R23078 CSoutput.n222 CSoutput.n213 2.2505
R23079 CSoutput.n246 CSoutput.n213 2.2505
R23080 CSoutput.n213 CSoutput.n207 2.2505
R23081 CSoutput.n268 CSoutput.n213 2.2505
R23082 CSoutput.n266 CSoutput.n213 2.2505
R23083 CSoutput.n248 CSoutput.n213 2.2505
R23084 CSoutput.n220 CSoutput.n213 2.2505
R23085 CSoutput.n250 CSoutput.n213 2.2505
R23086 CSoutput.n219 CSoutput.n213 2.2505
R23087 CSoutput.n264 CSoutput.n213 2.2505
R23088 CSoutput.n264 CSoutput.n217 2.2505
R23089 CSoutput.n164 CSoutput.n144 2.2505
R23090 CSoutput.n159 CSoutput.n144 2.2505
R23091 CSoutput.n157 CSoutput.n144 2.2505
R23092 CSoutput.n156 CSoutput.n144 2.2505
R23093 CSoutput.n285 CSoutput.n144 2.2505
R23094 CSoutput.n283 CSoutput.n144 2.2505
R23095 CSoutput.n281 CSoutput.n144 2.2505
R23096 CSoutput.n167 CSoutput.n144 2.2505
R23097 CSoutput.n166 CSoutput.n144 2.2505
R23098 CSoutput.n170 CSoutput.n144 2.2505
R23099 CSoutput.n169 CSoutput.n144 2.2505
R23100 CSoutput.n152 CSoutput.n144 2.2505
R23101 CSoutput.n288 CSoutput.n144 2.2505
R23102 CSoutput.n288 CSoutput.n287 2.2505
R23103 CSoutput.n206 CSoutput.n199 2.25024
R23104 CSoutput.n206 CSoutput.n192 2.25024
R23105 CSoutput.n274 CSoutput.n206 2.25024
R23106 CSoutput.n206 CSoutput.n202 2.25024
R23107 CSoutput.n206 CSoutput.n205 2.25024
R23108 CSoutput.n206 CSoutput.n173 2.25024
R23109 CSoutput.n256 CSoutput.n253 2.25024
R23110 CSoutput.n256 CSoutput.n252 2.25024
R23111 CSoutput.n256 CSoutput.n251 2.25024
R23112 CSoutput.n256 CSoutput.n218 2.25024
R23113 CSoutput.n256 CSoutput.n255 2.25024
R23114 CSoutput.n257 CSoutput.n256 2.25024
R23115 CSoutput.n172 CSoutput.n165 2.25024
R23116 CSoutput.n172 CSoutput.n158 2.25024
R23117 CSoutput.n284 CSoutput.n172 2.25024
R23118 CSoutput.n172 CSoutput.n168 2.25024
R23119 CSoutput.n172 CSoutput.n171 2.25024
R23120 CSoutput.n172 CSoutput.n139 2.25024
R23121 CSoutput.n273 CSoutput.n183 1.50111
R23122 CSoutput.n221 CSoutput.n207 1.50111
R23123 CSoutput.n283 CSoutput.n149 1.50111
R23124 CSoutput.n229 CSoutput.n228 1.501
R23125 CSoutput.n236 CSoutput.n235 1.501
R23126 CSoutput.n263 CSoutput.n262 1.501
R23127 CSoutput.n277 CSoutput.n188 1.12536
R23128 CSoutput.n277 CSoutput.n189 1.12536
R23129 CSoutput.n277 CSoutput.n276 1.12536
R23130 CSoutput.n237 CSoutput.n217 1.12536
R23131 CSoutput.n243 CSoutput.n217 1.12536
R23132 CSoutput.n245 CSoutput.n217 1.12536
R23133 CSoutput.n287 CSoutput.n154 1.12536
R23134 CSoutput.n287 CSoutput.n155 1.12536
R23135 CSoutput.n287 CSoutput.n286 1.12536
R23136 CSoutput.n277 CSoutput.n184 1.12536
R23137 CSoutput.n277 CSoutput.n185 1.12536
R23138 CSoutput.n277 CSoutput.n187 1.12536
R23139 CSoutput.n267 CSoutput.n217 1.12536
R23140 CSoutput.n247 CSoutput.n217 1.12536
R23141 CSoutput.n249 CSoutput.n217 1.12536
R23142 CSoutput.n287 CSoutput.n150 1.12536
R23143 CSoutput.n287 CSoutput.n151 1.12536
R23144 CSoutput.n287 CSoutput.n153 1.12536
R23145 CSoutput.n31 CSoutput.n30 0.669944
R23146 CSoutput.n62 CSoutput.n61 0.669944
R23147 CSoutput.n372 CSoutput.n370 0.573776
R23148 CSoutput.n374 CSoutput.n372 0.573776
R23149 CSoutput.n376 CSoutput.n374 0.573776
R23150 CSoutput.n378 CSoutput.n376 0.573776
R23151 CSoutput.n380 CSoutput.n378 0.573776
R23152 CSoutput.n382 CSoutput.n380 0.573776
R23153 CSoutput.n384 CSoutput.n382 0.573776
R23154 CSoutput.n386 CSoutput.n384 0.573776
R23155 CSoutput.n353 CSoutput.n351 0.573776
R23156 CSoutput.n355 CSoutput.n353 0.573776
R23157 CSoutput.n357 CSoutput.n355 0.573776
R23158 CSoutput.n359 CSoutput.n357 0.573776
R23159 CSoutput.n361 CSoutput.n359 0.573776
R23160 CSoutput.n363 CSoutput.n361 0.573776
R23161 CSoutput.n365 CSoutput.n363 0.573776
R23162 CSoutput.n367 CSoutput.n365 0.573776
R23163 CSoutput.n426 CSoutput.n424 0.573776
R23164 CSoutput.n424 CSoutput.n422 0.573776
R23165 CSoutput.n422 CSoutput.n420 0.573776
R23166 CSoutput.n420 CSoutput.n418 0.573776
R23167 CSoutput.n418 CSoutput.n416 0.573776
R23168 CSoutput.n416 CSoutput.n414 0.573776
R23169 CSoutput.n414 CSoutput.n412 0.573776
R23170 CSoutput.n412 CSoutput.n410 0.573776
R23171 CSoutput.n407 CSoutput.n405 0.573776
R23172 CSoutput.n405 CSoutput.n403 0.573776
R23173 CSoutput.n403 CSoutput.n401 0.573776
R23174 CSoutput.n401 CSoutput.n399 0.573776
R23175 CSoutput.n399 CSoutput.n397 0.573776
R23176 CSoutput.n397 CSoutput.n395 0.573776
R23177 CSoutput.n395 CSoutput.n393 0.573776
R23178 CSoutput.n393 CSoutput.n391 0.573776
R23179 CSoutput.n429 CSoutput.n288 0.53442
R23180 CSoutput.n332 CSoutput.n330 0.358259
R23181 CSoutput.n334 CSoutput.n332 0.358259
R23182 CSoutput.n336 CSoutput.n334 0.358259
R23183 CSoutput.n338 CSoutput.n336 0.358259
R23184 CSoutput.n340 CSoutput.n338 0.358259
R23185 CSoutput.n342 CSoutput.n340 0.358259
R23186 CSoutput.n344 CSoutput.n342 0.358259
R23187 CSoutput.n346 CSoutput.n344 0.358259
R23188 CSoutput.n312 CSoutput.n310 0.358259
R23189 CSoutput.n314 CSoutput.n312 0.358259
R23190 CSoutput.n316 CSoutput.n314 0.358259
R23191 CSoutput.n318 CSoutput.n316 0.358259
R23192 CSoutput.n320 CSoutput.n318 0.358259
R23193 CSoutput.n322 CSoutput.n320 0.358259
R23194 CSoutput.n324 CSoutput.n322 0.358259
R23195 CSoutput.n326 CSoutput.n324 0.358259
R23196 CSoutput.n293 CSoutput.n291 0.358259
R23197 CSoutput.n295 CSoutput.n293 0.358259
R23198 CSoutput.n297 CSoutput.n295 0.358259
R23199 CSoutput.n299 CSoutput.n297 0.358259
R23200 CSoutput.n301 CSoutput.n299 0.358259
R23201 CSoutput.n303 CSoutput.n301 0.358259
R23202 CSoutput.n305 CSoutput.n303 0.358259
R23203 CSoutput.n307 CSoutput.n305 0.358259
R23204 CSoutput.n136 CSoutput.n134 0.358259
R23205 CSoutput.n134 CSoutput.n132 0.358259
R23206 CSoutput.n132 CSoutput.n130 0.358259
R23207 CSoutput.n130 CSoutput.n128 0.358259
R23208 CSoutput.n128 CSoutput.n126 0.358259
R23209 CSoutput.n126 CSoutput.n124 0.358259
R23210 CSoutput.n124 CSoutput.n122 0.358259
R23211 CSoutput.n122 CSoutput.n120 0.358259
R23212 CSoutput.n116 CSoutput.n114 0.358259
R23213 CSoutput.n114 CSoutput.n112 0.358259
R23214 CSoutput.n112 CSoutput.n110 0.358259
R23215 CSoutput.n110 CSoutput.n108 0.358259
R23216 CSoutput.n108 CSoutput.n106 0.358259
R23217 CSoutput.n106 CSoutput.n104 0.358259
R23218 CSoutput.n104 CSoutput.n102 0.358259
R23219 CSoutput.n102 CSoutput.n100 0.358259
R23220 CSoutput.n97 CSoutput.n95 0.358259
R23221 CSoutput.n95 CSoutput.n93 0.358259
R23222 CSoutput.n93 CSoutput.n91 0.358259
R23223 CSoutput.n91 CSoutput.n89 0.358259
R23224 CSoutput.n89 CSoutput.n87 0.358259
R23225 CSoutput.n87 CSoutput.n85 0.358259
R23226 CSoutput.n85 CSoutput.n83 0.358259
R23227 CSoutput.n83 CSoutput.n81 0.358259
R23228 CSoutput.n21 CSoutput.n20 0.169105
R23229 CSoutput.n21 CSoutput.n16 0.169105
R23230 CSoutput.n26 CSoutput.n16 0.169105
R23231 CSoutput.n27 CSoutput.n26 0.169105
R23232 CSoutput.n27 CSoutput.n14 0.169105
R23233 CSoutput.n32 CSoutput.n14 0.169105
R23234 CSoutput.n33 CSoutput.n32 0.169105
R23235 CSoutput.n34 CSoutput.n33 0.169105
R23236 CSoutput.n34 CSoutput.n12 0.169105
R23237 CSoutput.n39 CSoutput.n12 0.169105
R23238 CSoutput.n40 CSoutput.n39 0.169105
R23239 CSoutput.n40 CSoutput.n10 0.169105
R23240 CSoutput.n45 CSoutput.n10 0.169105
R23241 CSoutput.n46 CSoutput.n45 0.169105
R23242 CSoutput.n47 CSoutput.n46 0.169105
R23243 CSoutput.n47 CSoutput.n8 0.169105
R23244 CSoutput.n52 CSoutput.n8 0.169105
R23245 CSoutput.n53 CSoutput.n52 0.169105
R23246 CSoutput.n53 CSoutput.n6 0.169105
R23247 CSoutput.n58 CSoutput.n6 0.169105
R23248 CSoutput.n59 CSoutput.n58 0.169105
R23249 CSoutput.n60 CSoutput.n59 0.169105
R23250 CSoutput.n60 CSoutput.n4 0.169105
R23251 CSoutput.n66 CSoutput.n4 0.169105
R23252 CSoutput.n67 CSoutput.n66 0.169105
R23253 CSoutput.n68 CSoutput.n67 0.169105
R23254 CSoutput.n68 CSoutput.n2 0.169105
R23255 CSoutput.n73 CSoutput.n2 0.169105
R23256 CSoutput.n74 CSoutput.n73 0.169105
R23257 CSoutput.n74 CSoutput.n0 0.169105
R23258 CSoutput.n78 CSoutput.n0 0.169105
R23259 CSoutput.n231 CSoutput.n230 0.0910737
R23260 CSoutput.n282 CSoutput.n279 0.0723685
R23261 CSoutput.n236 CSoutput.n231 0.0522944
R23262 CSoutput.n279 CSoutput.n278 0.0499135
R23263 CSoutput.n230 CSoutput.n229 0.0499135
R23264 CSoutput.n264 CSoutput.n263 0.0464294
R23265 CSoutput.n272 CSoutput.n269 0.0391444
R23266 CSoutput.n231 CSoutput.t216 0.023435
R23267 CSoutput.n279 CSoutput.t205 0.02262
R23268 CSoutput.n230 CSoutput.t214 0.02262
R23269 CSoutput CSoutput.n429 0.0052
R23270 CSoutput.n201 CSoutput.n184 0.00365111
R23271 CSoutput.n204 CSoutput.n185 0.00365111
R23272 CSoutput.n187 CSoutput.n186 0.00365111
R23273 CSoutput.n229 CSoutput.n188 0.00365111
R23274 CSoutput.n193 CSoutput.n189 0.00365111
R23275 CSoutput.n276 CSoutput.n190 0.00365111
R23276 CSoutput.n267 CSoutput.n266 0.00365111
R23277 CSoutput.n247 CSoutput.n220 0.00365111
R23278 CSoutput.n249 CSoutput.n219 0.00365111
R23279 CSoutput.n237 CSoutput.n236 0.00365111
R23280 CSoutput.n243 CSoutput.n223 0.00365111
R23281 CSoutput.n245 CSoutput.n222 0.00365111
R23282 CSoutput.n167 CSoutput.n150 0.00365111
R23283 CSoutput.n170 CSoutput.n151 0.00365111
R23284 CSoutput.n153 CSoutput.n152 0.00365111
R23285 CSoutput.n263 CSoutput.n154 0.00365111
R23286 CSoutput.n159 CSoutput.n155 0.00365111
R23287 CSoutput.n286 CSoutput.n156 0.00365111
R23288 CSoutput.n198 CSoutput.n188 0.00340054
R23289 CSoutput.n191 CSoutput.n189 0.00340054
R23290 CSoutput.n276 CSoutput.n275 0.00340054
R23291 CSoutput.n271 CSoutput.n184 0.00340054
R23292 CSoutput.n200 CSoutput.n185 0.00340054
R23293 CSoutput.n203 CSoutput.n187 0.00340054
R23294 CSoutput.n242 CSoutput.n237 0.00340054
R23295 CSoutput.n244 CSoutput.n243 0.00340054
R23296 CSoutput.n246 CSoutput.n245 0.00340054
R23297 CSoutput.n268 CSoutput.n267 0.00340054
R23298 CSoutput.n248 CSoutput.n247 0.00340054
R23299 CSoutput.n250 CSoutput.n249 0.00340054
R23300 CSoutput.n164 CSoutput.n154 0.00340054
R23301 CSoutput.n157 CSoutput.n155 0.00340054
R23302 CSoutput.n286 CSoutput.n285 0.00340054
R23303 CSoutput.n281 CSoutput.n150 0.00340054
R23304 CSoutput.n166 CSoutput.n151 0.00340054
R23305 CSoutput.n169 CSoutput.n153 0.00340054
R23306 CSoutput.n199 CSoutput.n193 0.00252698
R23307 CSoutput.n192 CSoutput.n190 0.00252698
R23308 CSoutput.n274 CSoutput.n273 0.00252698
R23309 CSoutput.n202 CSoutput.n200 0.00252698
R23310 CSoutput.n205 CSoutput.n203 0.00252698
R23311 CSoutput.n278 CSoutput.n173 0.00252698
R23312 CSoutput.n199 CSoutput.n198 0.00252698
R23313 CSoutput.n192 CSoutput.n191 0.00252698
R23314 CSoutput.n275 CSoutput.n274 0.00252698
R23315 CSoutput.n202 CSoutput.n201 0.00252698
R23316 CSoutput.n205 CSoutput.n204 0.00252698
R23317 CSoutput.n186 CSoutput.n173 0.00252698
R23318 CSoutput.n253 CSoutput.n223 0.00252698
R23319 CSoutput.n252 CSoutput.n222 0.00252698
R23320 CSoutput.n251 CSoutput.n207 0.00252698
R23321 CSoutput.n248 CSoutput.n218 0.00252698
R23322 CSoutput.n255 CSoutput.n250 0.00252698
R23323 CSoutput.n264 CSoutput.n257 0.00252698
R23324 CSoutput.n253 CSoutput.n242 0.00252698
R23325 CSoutput.n252 CSoutput.n244 0.00252698
R23326 CSoutput.n251 CSoutput.n246 0.00252698
R23327 CSoutput.n266 CSoutput.n218 0.00252698
R23328 CSoutput.n255 CSoutput.n220 0.00252698
R23329 CSoutput.n257 CSoutput.n219 0.00252698
R23330 CSoutput.n165 CSoutput.n159 0.00252698
R23331 CSoutput.n158 CSoutput.n156 0.00252698
R23332 CSoutput.n284 CSoutput.n283 0.00252698
R23333 CSoutput.n168 CSoutput.n166 0.00252698
R23334 CSoutput.n171 CSoutput.n169 0.00252698
R23335 CSoutput.n288 CSoutput.n139 0.00252698
R23336 CSoutput.n165 CSoutput.n164 0.00252698
R23337 CSoutput.n158 CSoutput.n157 0.00252698
R23338 CSoutput.n285 CSoutput.n284 0.00252698
R23339 CSoutput.n168 CSoutput.n167 0.00252698
R23340 CSoutput.n171 CSoutput.n170 0.00252698
R23341 CSoutput.n152 CSoutput.n139 0.00252698
R23342 CSoutput.n273 CSoutput.n272 0.0020275
R23343 CSoutput.n272 CSoutput.n271 0.0020275
R23344 CSoutput.n269 CSoutput.n207 0.0020275
R23345 CSoutput.n269 CSoutput.n268 0.0020275
R23346 CSoutput.n283 CSoutput.n282 0.0020275
R23347 CSoutput.n282 CSoutput.n281 0.0020275
R23348 CSoutput.n183 CSoutput.n182 0.00166668
R23349 CSoutput.n265 CSoutput.n221 0.00166668
R23350 CSoutput.n149 CSoutput.n148 0.00166668
R23351 CSoutput.n287 CSoutput.n149 0.00133328
R23352 CSoutput.n221 CSoutput.n217 0.00133328
R23353 CSoutput.n277 CSoutput.n183 0.00133328
R23354 CSoutput.n280 CSoutput.n172 0.001
R23355 CSoutput.n258 CSoutput.n172 0.001
R23356 CSoutput.n160 CSoutput.n140 0.001
R23357 CSoutput.n259 CSoutput.n140 0.001
R23358 CSoutput.n161 CSoutput.n141 0.001
R23359 CSoutput.n260 CSoutput.n141 0.001
R23360 CSoutput.n162 CSoutput.n142 0.001
R23361 CSoutput.n261 CSoutput.n142 0.001
R23362 CSoutput.n163 CSoutput.n143 0.001
R23363 CSoutput.n262 CSoutput.n143 0.001
R23364 CSoutput.n256 CSoutput.n208 0.001
R23365 CSoutput.n256 CSoutput.n254 0.001
R23366 CSoutput.n238 CSoutput.n209 0.001
R23367 CSoutput.n232 CSoutput.n209 0.001
R23368 CSoutput.n239 CSoutput.n210 0.001
R23369 CSoutput.n233 CSoutput.n210 0.001
R23370 CSoutput.n240 CSoutput.n211 0.001
R23371 CSoutput.n234 CSoutput.n211 0.001
R23372 CSoutput.n241 CSoutput.n212 0.001
R23373 CSoutput.n235 CSoutput.n212 0.001
R23374 CSoutput.n270 CSoutput.n206 0.001
R23375 CSoutput.n224 CSoutput.n206 0.001
R23376 CSoutput.n194 CSoutput.n174 0.001
R23377 CSoutput.n225 CSoutput.n174 0.001
R23378 CSoutput.n195 CSoutput.n175 0.001
R23379 CSoutput.n226 CSoutput.n175 0.001
R23380 CSoutput.n196 CSoutput.n176 0.001
R23381 CSoutput.n227 CSoutput.n176 0.001
R23382 CSoutput.n197 CSoutput.n177 0.001
R23383 CSoutput.n228 CSoutput.n177 0.001
R23384 CSoutput.n228 CSoutput.n178 0.001
R23385 CSoutput.n227 CSoutput.n179 0.001
R23386 CSoutput.n226 CSoutput.n180 0.001
R23387 CSoutput.n225 CSoutput.t208 0.001
R23388 CSoutput.n224 CSoutput.n181 0.001
R23389 CSoutput.n197 CSoutput.n179 0.001
R23390 CSoutput.n196 CSoutput.n180 0.001
R23391 CSoutput.n195 CSoutput.t208 0.001
R23392 CSoutput.n194 CSoutput.n181 0.001
R23393 CSoutput.n270 CSoutput.n182 0.001
R23394 CSoutput.n235 CSoutput.n213 0.001
R23395 CSoutput.n234 CSoutput.n214 0.001
R23396 CSoutput.n233 CSoutput.n215 0.001
R23397 CSoutput.n232 CSoutput.t210 0.001
R23398 CSoutput.n254 CSoutput.n216 0.001
R23399 CSoutput.n241 CSoutput.n214 0.001
R23400 CSoutput.n240 CSoutput.n215 0.001
R23401 CSoutput.n239 CSoutput.t210 0.001
R23402 CSoutput.n238 CSoutput.n216 0.001
R23403 CSoutput.n265 CSoutput.n208 0.001
R23404 CSoutput.n262 CSoutput.n144 0.001
R23405 CSoutput.n261 CSoutput.n145 0.001
R23406 CSoutput.n260 CSoutput.n146 0.001
R23407 CSoutput.n259 CSoutput.t211 0.001
R23408 CSoutput.n258 CSoutput.n147 0.001
R23409 CSoutput.n163 CSoutput.n145 0.001
R23410 CSoutput.n162 CSoutput.n146 0.001
R23411 CSoutput.n161 CSoutput.t211 0.001
R23412 CSoutput.n160 CSoutput.n147 0.001
R23413 CSoutput.n280 CSoutput.n148 0.001
R23414 outputibias.n27 outputibias.n1 289.615
R23415 outputibias.n58 outputibias.n32 289.615
R23416 outputibias.n90 outputibias.n64 289.615
R23417 outputibias.n122 outputibias.n96 289.615
R23418 outputibias.n28 outputibias.n27 185
R23419 outputibias.n26 outputibias.n25 185
R23420 outputibias.n5 outputibias.n4 185
R23421 outputibias.n20 outputibias.n19 185
R23422 outputibias.n18 outputibias.n17 185
R23423 outputibias.n9 outputibias.n8 185
R23424 outputibias.n12 outputibias.n11 185
R23425 outputibias.n59 outputibias.n58 185
R23426 outputibias.n57 outputibias.n56 185
R23427 outputibias.n36 outputibias.n35 185
R23428 outputibias.n51 outputibias.n50 185
R23429 outputibias.n49 outputibias.n48 185
R23430 outputibias.n40 outputibias.n39 185
R23431 outputibias.n43 outputibias.n42 185
R23432 outputibias.n91 outputibias.n90 185
R23433 outputibias.n89 outputibias.n88 185
R23434 outputibias.n68 outputibias.n67 185
R23435 outputibias.n83 outputibias.n82 185
R23436 outputibias.n81 outputibias.n80 185
R23437 outputibias.n72 outputibias.n71 185
R23438 outputibias.n75 outputibias.n74 185
R23439 outputibias.n123 outputibias.n122 185
R23440 outputibias.n121 outputibias.n120 185
R23441 outputibias.n100 outputibias.n99 185
R23442 outputibias.n115 outputibias.n114 185
R23443 outputibias.n113 outputibias.n112 185
R23444 outputibias.n104 outputibias.n103 185
R23445 outputibias.n107 outputibias.n106 185
R23446 outputibias.n0 outputibias.t8 178.945
R23447 outputibias.n133 outputibias.t9 177.018
R23448 outputibias.n132 outputibias.t11 177.018
R23449 outputibias.n0 outputibias.t10 177.018
R23450 outputibias.t5 outputibias.n10 147.661
R23451 outputibias.t3 outputibias.n41 147.661
R23452 outputibias.t1 outputibias.n73 147.661
R23453 outputibias.t7 outputibias.n105 147.661
R23454 outputibias.n128 outputibias.t4 132.363
R23455 outputibias.n128 outputibias.t2 130.436
R23456 outputibias.n129 outputibias.t0 130.436
R23457 outputibias.n130 outputibias.t6 130.436
R23458 outputibias.n27 outputibias.n26 104.615
R23459 outputibias.n26 outputibias.n4 104.615
R23460 outputibias.n19 outputibias.n4 104.615
R23461 outputibias.n19 outputibias.n18 104.615
R23462 outputibias.n18 outputibias.n8 104.615
R23463 outputibias.n11 outputibias.n8 104.615
R23464 outputibias.n58 outputibias.n57 104.615
R23465 outputibias.n57 outputibias.n35 104.615
R23466 outputibias.n50 outputibias.n35 104.615
R23467 outputibias.n50 outputibias.n49 104.615
R23468 outputibias.n49 outputibias.n39 104.615
R23469 outputibias.n42 outputibias.n39 104.615
R23470 outputibias.n90 outputibias.n89 104.615
R23471 outputibias.n89 outputibias.n67 104.615
R23472 outputibias.n82 outputibias.n67 104.615
R23473 outputibias.n82 outputibias.n81 104.615
R23474 outputibias.n81 outputibias.n71 104.615
R23475 outputibias.n74 outputibias.n71 104.615
R23476 outputibias.n122 outputibias.n121 104.615
R23477 outputibias.n121 outputibias.n99 104.615
R23478 outputibias.n114 outputibias.n99 104.615
R23479 outputibias.n114 outputibias.n113 104.615
R23480 outputibias.n113 outputibias.n103 104.615
R23481 outputibias.n106 outputibias.n103 104.615
R23482 outputibias.n63 outputibias.n31 95.6354
R23483 outputibias.n63 outputibias.n62 94.6732
R23484 outputibias.n95 outputibias.n94 94.6732
R23485 outputibias.n127 outputibias.n126 94.6732
R23486 outputibias.n11 outputibias.t5 52.3082
R23487 outputibias.n42 outputibias.t3 52.3082
R23488 outputibias.n74 outputibias.t1 52.3082
R23489 outputibias.n106 outputibias.t7 52.3082
R23490 outputibias.n12 outputibias.n10 15.6674
R23491 outputibias.n43 outputibias.n41 15.6674
R23492 outputibias.n75 outputibias.n73 15.6674
R23493 outputibias.n107 outputibias.n105 15.6674
R23494 outputibias.n13 outputibias.n9 12.8005
R23495 outputibias.n44 outputibias.n40 12.8005
R23496 outputibias.n76 outputibias.n72 12.8005
R23497 outputibias.n108 outputibias.n104 12.8005
R23498 outputibias.n17 outputibias.n16 12.0247
R23499 outputibias.n48 outputibias.n47 12.0247
R23500 outputibias.n80 outputibias.n79 12.0247
R23501 outputibias.n112 outputibias.n111 12.0247
R23502 outputibias.n20 outputibias.n7 11.249
R23503 outputibias.n51 outputibias.n38 11.249
R23504 outputibias.n83 outputibias.n70 11.249
R23505 outputibias.n115 outputibias.n102 11.249
R23506 outputibias.n21 outputibias.n5 10.4732
R23507 outputibias.n52 outputibias.n36 10.4732
R23508 outputibias.n84 outputibias.n68 10.4732
R23509 outputibias.n116 outputibias.n100 10.4732
R23510 outputibias.n25 outputibias.n24 9.69747
R23511 outputibias.n56 outputibias.n55 9.69747
R23512 outputibias.n88 outputibias.n87 9.69747
R23513 outputibias.n120 outputibias.n119 9.69747
R23514 outputibias.n31 outputibias.n30 9.45567
R23515 outputibias.n62 outputibias.n61 9.45567
R23516 outputibias.n94 outputibias.n93 9.45567
R23517 outputibias.n126 outputibias.n125 9.45567
R23518 outputibias.n30 outputibias.n29 9.3005
R23519 outputibias.n3 outputibias.n2 9.3005
R23520 outputibias.n24 outputibias.n23 9.3005
R23521 outputibias.n22 outputibias.n21 9.3005
R23522 outputibias.n7 outputibias.n6 9.3005
R23523 outputibias.n16 outputibias.n15 9.3005
R23524 outputibias.n14 outputibias.n13 9.3005
R23525 outputibias.n61 outputibias.n60 9.3005
R23526 outputibias.n34 outputibias.n33 9.3005
R23527 outputibias.n55 outputibias.n54 9.3005
R23528 outputibias.n53 outputibias.n52 9.3005
R23529 outputibias.n38 outputibias.n37 9.3005
R23530 outputibias.n47 outputibias.n46 9.3005
R23531 outputibias.n45 outputibias.n44 9.3005
R23532 outputibias.n93 outputibias.n92 9.3005
R23533 outputibias.n66 outputibias.n65 9.3005
R23534 outputibias.n87 outputibias.n86 9.3005
R23535 outputibias.n85 outputibias.n84 9.3005
R23536 outputibias.n70 outputibias.n69 9.3005
R23537 outputibias.n79 outputibias.n78 9.3005
R23538 outputibias.n77 outputibias.n76 9.3005
R23539 outputibias.n125 outputibias.n124 9.3005
R23540 outputibias.n98 outputibias.n97 9.3005
R23541 outputibias.n119 outputibias.n118 9.3005
R23542 outputibias.n117 outputibias.n116 9.3005
R23543 outputibias.n102 outputibias.n101 9.3005
R23544 outputibias.n111 outputibias.n110 9.3005
R23545 outputibias.n109 outputibias.n108 9.3005
R23546 outputibias.n28 outputibias.n3 8.92171
R23547 outputibias.n59 outputibias.n34 8.92171
R23548 outputibias.n91 outputibias.n66 8.92171
R23549 outputibias.n123 outputibias.n98 8.92171
R23550 outputibias.n29 outputibias.n1 8.14595
R23551 outputibias.n60 outputibias.n32 8.14595
R23552 outputibias.n92 outputibias.n64 8.14595
R23553 outputibias.n124 outputibias.n96 8.14595
R23554 outputibias.n31 outputibias.n1 5.81868
R23555 outputibias.n62 outputibias.n32 5.81868
R23556 outputibias.n94 outputibias.n64 5.81868
R23557 outputibias.n126 outputibias.n96 5.81868
R23558 outputibias.n131 outputibias.n130 5.20947
R23559 outputibias.n29 outputibias.n28 5.04292
R23560 outputibias.n60 outputibias.n59 5.04292
R23561 outputibias.n92 outputibias.n91 5.04292
R23562 outputibias.n124 outputibias.n123 5.04292
R23563 outputibias.n131 outputibias.n127 4.42209
R23564 outputibias.n14 outputibias.n10 4.38594
R23565 outputibias.n45 outputibias.n41 4.38594
R23566 outputibias.n77 outputibias.n73 4.38594
R23567 outputibias.n109 outputibias.n105 4.38594
R23568 outputibias.n132 outputibias.n131 4.28454
R23569 outputibias.n25 outputibias.n3 4.26717
R23570 outputibias.n56 outputibias.n34 4.26717
R23571 outputibias.n88 outputibias.n66 4.26717
R23572 outputibias.n120 outputibias.n98 4.26717
R23573 outputibias.n24 outputibias.n5 3.49141
R23574 outputibias.n55 outputibias.n36 3.49141
R23575 outputibias.n87 outputibias.n68 3.49141
R23576 outputibias.n119 outputibias.n100 3.49141
R23577 outputibias.n21 outputibias.n20 2.71565
R23578 outputibias.n52 outputibias.n51 2.71565
R23579 outputibias.n84 outputibias.n83 2.71565
R23580 outputibias.n116 outputibias.n115 2.71565
R23581 outputibias.n17 outputibias.n7 1.93989
R23582 outputibias.n48 outputibias.n38 1.93989
R23583 outputibias.n80 outputibias.n70 1.93989
R23584 outputibias.n112 outputibias.n102 1.93989
R23585 outputibias.n130 outputibias.n129 1.9266
R23586 outputibias.n129 outputibias.n128 1.9266
R23587 outputibias.n133 outputibias.n132 1.92658
R23588 outputibias.n134 outputibias.n133 1.29913
R23589 outputibias.n16 outputibias.n9 1.16414
R23590 outputibias.n47 outputibias.n40 1.16414
R23591 outputibias.n79 outputibias.n72 1.16414
R23592 outputibias.n111 outputibias.n104 1.16414
R23593 outputibias.n127 outputibias.n95 0.962709
R23594 outputibias.n95 outputibias.n63 0.962709
R23595 outputibias.n13 outputibias.n12 0.388379
R23596 outputibias.n44 outputibias.n43 0.388379
R23597 outputibias.n76 outputibias.n75 0.388379
R23598 outputibias.n108 outputibias.n107 0.388379
R23599 outputibias.n134 outputibias.n0 0.337251
R23600 outputibias outputibias.n134 0.302375
R23601 outputibias.n30 outputibias.n2 0.155672
R23602 outputibias.n23 outputibias.n2 0.155672
R23603 outputibias.n23 outputibias.n22 0.155672
R23604 outputibias.n22 outputibias.n6 0.155672
R23605 outputibias.n15 outputibias.n6 0.155672
R23606 outputibias.n15 outputibias.n14 0.155672
R23607 outputibias.n61 outputibias.n33 0.155672
R23608 outputibias.n54 outputibias.n33 0.155672
R23609 outputibias.n54 outputibias.n53 0.155672
R23610 outputibias.n53 outputibias.n37 0.155672
R23611 outputibias.n46 outputibias.n37 0.155672
R23612 outputibias.n46 outputibias.n45 0.155672
R23613 outputibias.n93 outputibias.n65 0.155672
R23614 outputibias.n86 outputibias.n65 0.155672
R23615 outputibias.n86 outputibias.n85 0.155672
R23616 outputibias.n85 outputibias.n69 0.155672
R23617 outputibias.n78 outputibias.n69 0.155672
R23618 outputibias.n78 outputibias.n77 0.155672
R23619 outputibias.n125 outputibias.n97 0.155672
R23620 outputibias.n118 outputibias.n97 0.155672
R23621 outputibias.n118 outputibias.n117 0.155672
R23622 outputibias.n117 outputibias.n101 0.155672
R23623 outputibias.n110 outputibias.n101 0.155672
R23624 outputibias.n110 outputibias.n109 0.155672
R23625 diffpairibias.n0 diffpairibias.t27 436.822
R23626 diffpairibias.n27 diffpairibias.t24 435.479
R23627 diffpairibias.n26 diffpairibias.t21 435.479
R23628 diffpairibias.n25 diffpairibias.t22 435.479
R23629 diffpairibias.n24 diffpairibias.t26 435.479
R23630 diffpairibias.n23 diffpairibias.t20 435.479
R23631 diffpairibias.n0 diffpairibias.t23 435.479
R23632 diffpairibias.n1 diffpairibias.t28 435.479
R23633 diffpairibias.n2 diffpairibias.t25 435.479
R23634 diffpairibias.n3 diffpairibias.t29 435.479
R23635 diffpairibias.n13 diffpairibias.t14 377.536
R23636 diffpairibias.n13 diffpairibias.t0 376.193
R23637 diffpairibias.n14 diffpairibias.t10 376.193
R23638 diffpairibias.n15 diffpairibias.t12 376.193
R23639 diffpairibias.n16 diffpairibias.t6 376.193
R23640 diffpairibias.n17 diffpairibias.t2 376.193
R23641 diffpairibias.n18 diffpairibias.t16 376.193
R23642 diffpairibias.n19 diffpairibias.t4 376.193
R23643 diffpairibias.n20 diffpairibias.t18 376.193
R23644 diffpairibias.n21 diffpairibias.t8 376.193
R23645 diffpairibias.n4 diffpairibias.t15 113.368
R23646 diffpairibias.n4 diffpairibias.t1 112.698
R23647 diffpairibias.n5 diffpairibias.t11 112.698
R23648 diffpairibias.n6 diffpairibias.t13 112.698
R23649 diffpairibias.n7 diffpairibias.t7 112.698
R23650 diffpairibias.n8 diffpairibias.t3 112.698
R23651 diffpairibias.n9 diffpairibias.t17 112.698
R23652 diffpairibias.n10 diffpairibias.t5 112.698
R23653 diffpairibias.n11 diffpairibias.t19 112.698
R23654 diffpairibias.n12 diffpairibias.t9 112.698
R23655 diffpairibias.n22 diffpairibias.n21 4.77242
R23656 diffpairibias.n22 diffpairibias.n12 4.30807
R23657 diffpairibias.n23 diffpairibias.n22 4.13945
R23658 diffpairibias.n21 diffpairibias.n20 1.34352
R23659 diffpairibias.n20 diffpairibias.n19 1.34352
R23660 diffpairibias.n19 diffpairibias.n18 1.34352
R23661 diffpairibias.n18 diffpairibias.n17 1.34352
R23662 diffpairibias.n17 diffpairibias.n16 1.34352
R23663 diffpairibias.n16 diffpairibias.n15 1.34352
R23664 diffpairibias.n15 diffpairibias.n14 1.34352
R23665 diffpairibias.n14 diffpairibias.n13 1.34352
R23666 diffpairibias.n3 diffpairibias.n2 1.34352
R23667 diffpairibias.n2 diffpairibias.n1 1.34352
R23668 diffpairibias.n1 diffpairibias.n0 1.34352
R23669 diffpairibias.n24 diffpairibias.n23 1.34352
R23670 diffpairibias.n25 diffpairibias.n24 1.34352
R23671 diffpairibias.n26 diffpairibias.n25 1.34352
R23672 diffpairibias.n27 diffpairibias.n26 1.34352
R23673 diffpairibias.n28 diffpairibias.n27 0.862419
R23674 diffpairibias diffpairibias.n28 0.684875
R23675 diffpairibias.n12 diffpairibias.n11 0.672012
R23676 diffpairibias.n11 diffpairibias.n10 0.672012
R23677 diffpairibias.n10 diffpairibias.n9 0.672012
R23678 diffpairibias.n9 diffpairibias.n8 0.672012
R23679 diffpairibias.n8 diffpairibias.n7 0.672012
R23680 diffpairibias.n7 diffpairibias.n6 0.672012
R23681 diffpairibias.n6 diffpairibias.n5 0.672012
R23682 diffpairibias.n5 diffpairibias.n4 0.672012
R23683 diffpairibias.n28 diffpairibias.n3 0.190907
R23684 commonsourceibias.n281 commonsourceibias.t101 222.032
R23685 commonsourceibias.n44 commonsourceibias.t78 222.032
R23686 commonsourceibias.n166 commonsourceibias.t117 222.032
R23687 commonsourceibias.n643 commonsourceibias.t106 222.032
R23688 commonsourceibias.n413 commonsourceibias.t28 222.032
R23689 commonsourceibias.n529 commonsourceibias.t123 222.032
R23690 commonsourceibias.n364 commonsourceibias.t100 207.983
R23691 commonsourceibias.n127 commonsourceibias.t74 207.983
R23692 commonsourceibias.n249 commonsourceibias.t115 207.983
R23693 commonsourceibias.n731 commonsourceibias.t122 207.983
R23694 commonsourceibias.n501 commonsourceibias.t14 207.983
R23695 commonsourceibias.n616 commonsourceibias.t140 207.983
R23696 commonsourceibias.n280 commonsourceibias.t87 168.701
R23697 commonsourceibias.n286 commonsourceibias.t129 168.701
R23698 commonsourceibias.n292 commonsourceibias.t110 168.701
R23699 commonsourceibias.n276 commonsourceibias.t93 168.701
R23700 commonsourceibias.n300 commonsourceibias.t95 168.701
R23701 commonsourceibias.n306 commonsourceibias.t121 168.701
R23702 commonsourceibias.n271 commonsourceibias.t102 168.701
R23703 commonsourceibias.n314 commonsourceibias.t108 168.701
R23704 commonsourceibias.n320 commonsourceibias.t159 168.701
R23705 commonsourceibias.n266 commonsourceibias.t138 168.701
R23706 commonsourceibias.n328 commonsourceibias.t118 168.701
R23707 commonsourceibias.n334 commonsourceibias.t83 168.701
R23708 commonsourceibias.n261 commonsourceibias.t86 168.701
R23709 commonsourceibias.n342 commonsourceibias.t128 168.701
R23710 commonsourceibias.n348 commonsourceibias.t109 168.701
R23711 commonsourceibias.n256 commonsourceibias.t92 168.701
R23712 commonsourceibias.n356 commonsourceibias.t137 168.701
R23713 commonsourceibias.n362 commonsourceibias.t119 168.701
R23714 commonsourceibias.n125 commonsourceibias.t20 168.701
R23715 commonsourceibias.n119 commonsourceibias.t50 168.701
R23716 commonsourceibias.n19 commonsourceibias.t8 168.701
R23717 commonsourceibias.n111 commonsourceibias.t36 168.701
R23718 commonsourceibias.n105 commonsourceibias.t76 168.701
R23719 commonsourceibias.n24 commonsourceibias.t24 168.701
R23720 commonsourceibias.n97 commonsourceibias.t34 168.701
R23721 commonsourceibias.n91 commonsourceibias.t10 168.701
R23722 commonsourceibias.n29 commonsourceibias.t40 168.701
R23723 commonsourceibias.n83 commonsourceibias.t56 168.701
R23724 commonsourceibias.n77 commonsourceibias.t26 168.701
R23725 commonsourceibias.n34 commonsourceibias.t38 168.701
R23726 commonsourceibias.n69 commonsourceibias.t70 168.701
R23727 commonsourceibias.n63 commonsourceibias.t18 168.701
R23728 commonsourceibias.n39 commonsourceibias.t22 168.701
R23729 commonsourceibias.n55 commonsourceibias.t54 168.701
R23730 commonsourceibias.n49 commonsourceibias.t4 168.701
R23731 commonsourceibias.n43 commonsourceibias.t46 168.701
R23732 commonsourceibias.n247 commonsourceibias.t136 168.701
R23733 commonsourceibias.n241 commonsourceibias.t151 168.701
R23734 commonsourceibias.n5 commonsourceibias.t105 168.701
R23735 commonsourceibias.n233 commonsourceibias.t126 168.701
R23736 commonsourceibias.n227 commonsourceibias.t144 168.701
R23737 commonsourceibias.n10 commonsourceibias.t98 168.701
R23738 commonsourceibias.n219 commonsourceibias.t94 168.701
R23739 commonsourceibias.n213 commonsourceibias.t135 168.701
R23740 commonsourceibias.n150 commonsourceibias.t153 168.701
R23741 commonsourceibias.n151 commonsourceibias.t88 168.701
R23742 commonsourceibias.n153 commonsourceibias.t125 168.701
R23743 commonsourceibias.n155 commonsourceibias.t120 168.701
R23744 commonsourceibias.n191 commonsourceibias.t139 168.701
R23745 commonsourceibias.n185 commonsourceibias.t112 168.701
R23746 commonsourceibias.n161 commonsourceibias.t107 168.701
R23747 commonsourceibias.n177 commonsourceibias.t127 168.701
R23748 commonsourceibias.n171 commonsourceibias.t146 168.701
R23749 commonsourceibias.n165 commonsourceibias.t99 168.701
R23750 commonsourceibias.n642 commonsourceibias.t90 168.701
R23751 commonsourceibias.n648 commonsourceibias.t134 168.701
R23752 commonsourceibias.n654 commonsourceibias.t116 168.701
R23753 commonsourceibias.n656 commonsourceibias.t96 168.701
R23754 commonsourceibias.n663 commonsourceibias.t91 168.701
R23755 commonsourceibias.n669 commonsourceibias.t145 168.701
R23756 commonsourceibias.n671 commonsourceibias.t124 168.701
R23757 commonsourceibias.n678 commonsourceibias.t131 168.701
R23758 commonsourceibias.n684 commonsourceibias.t152 168.701
R23759 commonsourceibias.n686 commonsourceibias.t157 168.701
R23760 commonsourceibias.n693 commonsourceibias.t141 168.701
R23761 commonsourceibias.n699 commonsourceibias.t97 168.701
R23762 commonsourceibias.n701 commonsourceibias.t81 168.701
R23763 commonsourceibias.n708 commonsourceibias.t149 168.701
R23764 commonsourceibias.n714 commonsourceibias.t132 168.701
R23765 commonsourceibias.n716 commonsourceibias.t111 168.701
R23766 commonsourceibias.n723 commonsourceibias.t156 168.701
R23767 commonsourceibias.n729 commonsourceibias.t142 168.701
R23768 commonsourceibias.n412 commonsourceibias.t2 168.701
R23769 commonsourceibias.n418 commonsourceibias.t48 168.701
R23770 commonsourceibias.n424 commonsourceibias.t12 168.701
R23771 commonsourceibias.n426 commonsourceibias.t68 168.701
R23772 commonsourceibias.n433 commonsourceibias.t66 168.701
R23773 commonsourceibias.n439 commonsourceibias.t6 168.701
R23774 commonsourceibias.n441 commonsourceibias.t62 168.701
R23775 commonsourceibias.n448 commonsourceibias.t52 168.701
R23776 commonsourceibias.n454 commonsourceibias.t72 168.701
R23777 commonsourceibias.n456 commonsourceibias.t64 168.701
R23778 commonsourceibias.n463 commonsourceibias.t32 168.701
R23779 commonsourceibias.n469 commonsourceibias.t58 168.701
R23780 commonsourceibias.n471 commonsourceibias.t44 168.701
R23781 commonsourceibias.n478 commonsourceibias.t16 168.701
R23782 commonsourceibias.n484 commonsourceibias.t60 168.701
R23783 commonsourceibias.n486 commonsourceibias.t30 168.701
R23784 commonsourceibias.n493 commonsourceibias.t0 168.701
R23785 commonsourceibias.n499 commonsourceibias.t42 168.701
R23786 commonsourceibias.n614 commonsourceibias.t155 168.701
R23787 commonsourceibias.n608 commonsourceibias.t84 168.701
R23788 commonsourceibias.n601 commonsourceibias.t130 168.701
R23789 commonsourceibias.n599 commonsourceibias.t148 168.701
R23790 commonsourceibias.n593 commonsourceibias.t80 168.701
R23791 commonsourceibias.n586 commonsourceibias.t89 168.701
R23792 commonsourceibias.n584 commonsourceibias.t113 168.701
R23793 commonsourceibias.n578 commonsourceibias.t154 168.701
R23794 commonsourceibias.n571 commonsourceibias.t85 168.701
R23795 commonsourceibias.n528 commonsourceibias.t103 168.701
R23796 commonsourceibias.n534 commonsourceibias.t150 168.701
R23797 commonsourceibias.n540 commonsourceibias.t133 168.701
R23798 commonsourceibias.n542 commonsourceibias.t114 168.701
R23799 commonsourceibias.n549 commonsourceibias.t104 168.701
R23800 commonsourceibias.n555 commonsourceibias.t158 168.701
R23801 commonsourceibias.n519 commonsourceibias.t143 168.701
R23802 commonsourceibias.n517 commonsourceibias.t147 168.701
R23803 commonsourceibias.n515 commonsourceibias.t82 168.701
R23804 commonsourceibias.n363 commonsourceibias.n251 161.3
R23805 commonsourceibias.n361 commonsourceibias.n360 161.3
R23806 commonsourceibias.n359 commonsourceibias.n252 161.3
R23807 commonsourceibias.n358 commonsourceibias.n357 161.3
R23808 commonsourceibias.n355 commonsourceibias.n253 161.3
R23809 commonsourceibias.n354 commonsourceibias.n353 161.3
R23810 commonsourceibias.n352 commonsourceibias.n254 161.3
R23811 commonsourceibias.n351 commonsourceibias.n350 161.3
R23812 commonsourceibias.n349 commonsourceibias.n255 161.3
R23813 commonsourceibias.n347 commonsourceibias.n346 161.3
R23814 commonsourceibias.n345 commonsourceibias.n257 161.3
R23815 commonsourceibias.n344 commonsourceibias.n343 161.3
R23816 commonsourceibias.n341 commonsourceibias.n258 161.3
R23817 commonsourceibias.n340 commonsourceibias.n339 161.3
R23818 commonsourceibias.n338 commonsourceibias.n259 161.3
R23819 commonsourceibias.n337 commonsourceibias.n336 161.3
R23820 commonsourceibias.n335 commonsourceibias.n260 161.3
R23821 commonsourceibias.n333 commonsourceibias.n332 161.3
R23822 commonsourceibias.n331 commonsourceibias.n262 161.3
R23823 commonsourceibias.n330 commonsourceibias.n329 161.3
R23824 commonsourceibias.n327 commonsourceibias.n263 161.3
R23825 commonsourceibias.n326 commonsourceibias.n325 161.3
R23826 commonsourceibias.n324 commonsourceibias.n264 161.3
R23827 commonsourceibias.n323 commonsourceibias.n322 161.3
R23828 commonsourceibias.n321 commonsourceibias.n265 161.3
R23829 commonsourceibias.n319 commonsourceibias.n318 161.3
R23830 commonsourceibias.n317 commonsourceibias.n267 161.3
R23831 commonsourceibias.n316 commonsourceibias.n315 161.3
R23832 commonsourceibias.n313 commonsourceibias.n268 161.3
R23833 commonsourceibias.n312 commonsourceibias.n311 161.3
R23834 commonsourceibias.n310 commonsourceibias.n269 161.3
R23835 commonsourceibias.n309 commonsourceibias.n308 161.3
R23836 commonsourceibias.n307 commonsourceibias.n270 161.3
R23837 commonsourceibias.n305 commonsourceibias.n304 161.3
R23838 commonsourceibias.n303 commonsourceibias.n272 161.3
R23839 commonsourceibias.n302 commonsourceibias.n301 161.3
R23840 commonsourceibias.n299 commonsourceibias.n273 161.3
R23841 commonsourceibias.n298 commonsourceibias.n297 161.3
R23842 commonsourceibias.n296 commonsourceibias.n274 161.3
R23843 commonsourceibias.n295 commonsourceibias.n294 161.3
R23844 commonsourceibias.n293 commonsourceibias.n275 161.3
R23845 commonsourceibias.n291 commonsourceibias.n290 161.3
R23846 commonsourceibias.n289 commonsourceibias.n277 161.3
R23847 commonsourceibias.n288 commonsourceibias.n287 161.3
R23848 commonsourceibias.n285 commonsourceibias.n278 161.3
R23849 commonsourceibias.n284 commonsourceibias.n283 161.3
R23850 commonsourceibias.n282 commonsourceibias.n279 161.3
R23851 commonsourceibias.n45 commonsourceibias.n42 161.3
R23852 commonsourceibias.n47 commonsourceibias.n46 161.3
R23853 commonsourceibias.n48 commonsourceibias.n41 161.3
R23854 commonsourceibias.n51 commonsourceibias.n50 161.3
R23855 commonsourceibias.n52 commonsourceibias.n40 161.3
R23856 commonsourceibias.n54 commonsourceibias.n53 161.3
R23857 commonsourceibias.n56 commonsourceibias.n38 161.3
R23858 commonsourceibias.n58 commonsourceibias.n57 161.3
R23859 commonsourceibias.n59 commonsourceibias.n37 161.3
R23860 commonsourceibias.n61 commonsourceibias.n60 161.3
R23861 commonsourceibias.n62 commonsourceibias.n36 161.3
R23862 commonsourceibias.n65 commonsourceibias.n64 161.3
R23863 commonsourceibias.n66 commonsourceibias.n35 161.3
R23864 commonsourceibias.n68 commonsourceibias.n67 161.3
R23865 commonsourceibias.n70 commonsourceibias.n33 161.3
R23866 commonsourceibias.n72 commonsourceibias.n71 161.3
R23867 commonsourceibias.n73 commonsourceibias.n32 161.3
R23868 commonsourceibias.n75 commonsourceibias.n74 161.3
R23869 commonsourceibias.n76 commonsourceibias.n31 161.3
R23870 commonsourceibias.n79 commonsourceibias.n78 161.3
R23871 commonsourceibias.n80 commonsourceibias.n30 161.3
R23872 commonsourceibias.n82 commonsourceibias.n81 161.3
R23873 commonsourceibias.n84 commonsourceibias.n28 161.3
R23874 commonsourceibias.n86 commonsourceibias.n85 161.3
R23875 commonsourceibias.n87 commonsourceibias.n27 161.3
R23876 commonsourceibias.n89 commonsourceibias.n88 161.3
R23877 commonsourceibias.n90 commonsourceibias.n26 161.3
R23878 commonsourceibias.n93 commonsourceibias.n92 161.3
R23879 commonsourceibias.n94 commonsourceibias.n25 161.3
R23880 commonsourceibias.n96 commonsourceibias.n95 161.3
R23881 commonsourceibias.n98 commonsourceibias.n23 161.3
R23882 commonsourceibias.n100 commonsourceibias.n99 161.3
R23883 commonsourceibias.n101 commonsourceibias.n22 161.3
R23884 commonsourceibias.n103 commonsourceibias.n102 161.3
R23885 commonsourceibias.n104 commonsourceibias.n21 161.3
R23886 commonsourceibias.n107 commonsourceibias.n106 161.3
R23887 commonsourceibias.n108 commonsourceibias.n20 161.3
R23888 commonsourceibias.n110 commonsourceibias.n109 161.3
R23889 commonsourceibias.n112 commonsourceibias.n18 161.3
R23890 commonsourceibias.n114 commonsourceibias.n113 161.3
R23891 commonsourceibias.n115 commonsourceibias.n17 161.3
R23892 commonsourceibias.n117 commonsourceibias.n116 161.3
R23893 commonsourceibias.n118 commonsourceibias.n16 161.3
R23894 commonsourceibias.n121 commonsourceibias.n120 161.3
R23895 commonsourceibias.n122 commonsourceibias.n15 161.3
R23896 commonsourceibias.n124 commonsourceibias.n123 161.3
R23897 commonsourceibias.n126 commonsourceibias.n14 161.3
R23898 commonsourceibias.n167 commonsourceibias.n164 161.3
R23899 commonsourceibias.n169 commonsourceibias.n168 161.3
R23900 commonsourceibias.n170 commonsourceibias.n163 161.3
R23901 commonsourceibias.n173 commonsourceibias.n172 161.3
R23902 commonsourceibias.n174 commonsourceibias.n162 161.3
R23903 commonsourceibias.n176 commonsourceibias.n175 161.3
R23904 commonsourceibias.n178 commonsourceibias.n160 161.3
R23905 commonsourceibias.n180 commonsourceibias.n179 161.3
R23906 commonsourceibias.n181 commonsourceibias.n159 161.3
R23907 commonsourceibias.n183 commonsourceibias.n182 161.3
R23908 commonsourceibias.n184 commonsourceibias.n158 161.3
R23909 commonsourceibias.n187 commonsourceibias.n186 161.3
R23910 commonsourceibias.n188 commonsourceibias.n157 161.3
R23911 commonsourceibias.n190 commonsourceibias.n189 161.3
R23912 commonsourceibias.n192 commonsourceibias.n156 161.3
R23913 commonsourceibias.n194 commonsourceibias.n193 161.3
R23914 commonsourceibias.n196 commonsourceibias.n195 161.3
R23915 commonsourceibias.n197 commonsourceibias.n154 161.3
R23916 commonsourceibias.n199 commonsourceibias.n198 161.3
R23917 commonsourceibias.n201 commonsourceibias.n200 161.3
R23918 commonsourceibias.n202 commonsourceibias.n152 161.3
R23919 commonsourceibias.n204 commonsourceibias.n203 161.3
R23920 commonsourceibias.n206 commonsourceibias.n205 161.3
R23921 commonsourceibias.n208 commonsourceibias.n207 161.3
R23922 commonsourceibias.n209 commonsourceibias.n13 161.3
R23923 commonsourceibias.n211 commonsourceibias.n210 161.3
R23924 commonsourceibias.n212 commonsourceibias.n12 161.3
R23925 commonsourceibias.n215 commonsourceibias.n214 161.3
R23926 commonsourceibias.n216 commonsourceibias.n11 161.3
R23927 commonsourceibias.n218 commonsourceibias.n217 161.3
R23928 commonsourceibias.n220 commonsourceibias.n9 161.3
R23929 commonsourceibias.n222 commonsourceibias.n221 161.3
R23930 commonsourceibias.n223 commonsourceibias.n8 161.3
R23931 commonsourceibias.n225 commonsourceibias.n224 161.3
R23932 commonsourceibias.n226 commonsourceibias.n7 161.3
R23933 commonsourceibias.n229 commonsourceibias.n228 161.3
R23934 commonsourceibias.n230 commonsourceibias.n6 161.3
R23935 commonsourceibias.n232 commonsourceibias.n231 161.3
R23936 commonsourceibias.n234 commonsourceibias.n4 161.3
R23937 commonsourceibias.n236 commonsourceibias.n235 161.3
R23938 commonsourceibias.n237 commonsourceibias.n3 161.3
R23939 commonsourceibias.n239 commonsourceibias.n238 161.3
R23940 commonsourceibias.n240 commonsourceibias.n2 161.3
R23941 commonsourceibias.n243 commonsourceibias.n242 161.3
R23942 commonsourceibias.n244 commonsourceibias.n1 161.3
R23943 commonsourceibias.n246 commonsourceibias.n245 161.3
R23944 commonsourceibias.n248 commonsourceibias.n0 161.3
R23945 commonsourceibias.n730 commonsourceibias.n618 161.3
R23946 commonsourceibias.n728 commonsourceibias.n727 161.3
R23947 commonsourceibias.n726 commonsourceibias.n619 161.3
R23948 commonsourceibias.n725 commonsourceibias.n724 161.3
R23949 commonsourceibias.n722 commonsourceibias.n620 161.3
R23950 commonsourceibias.n721 commonsourceibias.n720 161.3
R23951 commonsourceibias.n719 commonsourceibias.n621 161.3
R23952 commonsourceibias.n718 commonsourceibias.n717 161.3
R23953 commonsourceibias.n715 commonsourceibias.n622 161.3
R23954 commonsourceibias.n713 commonsourceibias.n712 161.3
R23955 commonsourceibias.n711 commonsourceibias.n623 161.3
R23956 commonsourceibias.n710 commonsourceibias.n709 161.3
R23957 commonsourceibias.n707 commonsourceibias.n624 161.3
R23958 commonsourceibias.n706 commonsourceibias.n705 161.3
R23959 commonsourceibias.n704 commonsourceibias.n625 161.3
R23960 commonsourceibias.n703 commonsourceibias.n702 161.3
R23961 commonsourceibias.n700 commonsourceibias.n626 161.3
R23962 commonsourceibias.n698 commonsourceibias.n697 161.3
R23963 commonsourceibias.n696 commonsourceibias.n627 161.3
R23964 commonsourceibias.n695 commonsourceibias.n694 161.3
R23965 commonsourceibias.n692 commonsourceibias.n628 161.3
R23966 commonsourceibias.n691 commonsourceibias.n690 161.3
R23967 commonsourceibias.n689 commonsourceibias.n629 161.3
R23968 commonsourceibias.n688 commonsourceibias.n687 161.3
R23969 commonsourceibias.n685 commonsourceibias.n630 161.3
R23970 commonsourceibias.n683 commonsourceibias.n682 161.3
R23971 commonsourceibias.n681 commonsourceibias.n631 161.3
R23972 commonsourceibias.n680 commonsourceibias.n679 161.3
R23973 commonsourceibias.n677 commonsourceibias.n632 161.3
R23974 commonsourceibias.n676 commonsourceibias.n675 161.3
R23975 commonsourceibias.n674 commonsourceibias.n633 161.3
R23976 commonsourceibias.n673 commonsourceibias.n672 161.3
R23977 commonsourceibias.n670 commonsourceibias.n634 161.3
R23978 commonsourceibias.n668 commonsourceibias.n667 161.3
R23979 commonsourceibias.n666 commonsourceibias.n635 161.3
R23980 commonsourceibias.n665 commonsourceibias.n664 161.3
R23981 commonsourceibias.n662 commonsourceibias.n636 161.3
R23982 commonsourceibias.n661 commonsourceibias.n660 161.3
R23983 commonsourceibias.n659 commonsourceibias.n637 161.3
R23984 commonsourceibias.n658 commonsourceibias.n657 161.3
R23985 commonsourceibias.n655 commonsourceibias.n638 161.3
R23986 commonsourceibias.n653 commonsourceibias.n652 161.3
R23987 commonsourceibias.n651 commonsourceibias.n639 161.3
R23988 commonsourceibias.n650 commonsourceibias.n649 161.3
R23989 commonsourceibias.n647 commonsourceibias.n640 161.3
R23990 commonsourceibias.n646 commonsourceibias.n645 161.3
R23991 commonsourceibias.n644 commonsourceibias.n641 161.3
R23992 commonsourceibias.n500 commonsourceibias.n388 161.3
R23993 commonsourceibias.n498 commonsourceibias.n497 161.3
R23994 commonsourceibias.n496 commonsourceibias.n389 161.3
R23995 commonsourceibias.n495 commonsourceibias.n494 161.3
R23996 commonsourceibias.n492 commonsourceibias.n390 161.3
R23997 commonsourceibias.n491 commonsourceibias.n490 161.3
R23998 commonsourceibias.n489 commonsourceibias.n391 161.3
R23999 commonsourceibias.n488 commonsourceibias.n487 161.3
R24000 commonsourceibias.n485 commonsourceibias.n392 161.3
R24001 commonsourceibias.n483 commonsourceibias.n482 161.3
R24002 commonsourceibias.n481 commonsourceibias.n393 161.3
R24003 commonsourceibias.n480 commonsourceibias.n479 161.3
R24004 commonsourceibias.n477 commonsourceibias.n394 161.3
R24005 commonsourceibias.n476 commonsourceibias.n475 161.3
R24006 commonsourceibias.n474 commonsourceibias.n395 161.3
R24007 commonsourceibias.n473 commonsourceibias.n472 161.3
R24008 commonsourceibias.n470 commonsourceibias.n396 161.3
R24009 commonsourceibias.n468 commonsourceibias.n467 161.3
R24010 commonsourceibias.n466 commonsourceibias.n397 161.3
R24011 commonsourceibias.n465 commonsourceibias.n464 161.3
R24012 commonsourceibias.n462 commonsourceibias.n398 161.3
R24013 commonsourceibias.n461 commonsourceibias.n460 161.3
R24014 commonsourceibias.n459 commonsourceibias.n399 161.3
R24015 commonsourceibias.n458 commonsourceibias.n457 161.3
R24016 commonsourceibias.n455 commonsourceibias.n400 161.3
R24017 commonsourceibias.n453 commonsourceibias.n452 161.3
R24018 commonsourceibias.n451 commonsourceibias.n401 161.3
R24019 commonsourceibias.n450 commonsourceibias.n449 161.3
R24020 commonsourceibias.n447 commonsourceibias.n402 161.3
R24021 commonsourceibias.n446 commonsourceibias.n445 161.3
R24022 commonsourceibias.n444 commonsourceibias.n403 161.3
R24023 commonsourceibias.n443 commonsourceibias.n442 161.3
R24024 commonsourceibias.n440 commonsourceibias.n404 161.3
R24025 commonsourceibias.n438 commonsourceibias.n437 161.3
R24026 commonsourceibias.n436 commonsourceibias.n405 161.3
R24027 commonsourceibias.n435 commonsourceibias.n434 161.3
R24028 commonsourceibias.n432 commonsourceibias.n406 161.3
R24029 commonsourceibias.n431 commonsourceibias.n430 161.3
R24030 commonsourceibias.n429 commonsourceibias.n407 161.3
R24031 commonsourceibias.n428 commonsourceibias.n427 161.3
R24032 commonsourceibias.n425 commonsourceibias.n408 161.3
R24033 commonsourceibias.n423 commonsourceibias.n422 161.3
R24034 commonsourceibias.n421 commonsourceibias.n409 161.3
R24035 commonsourceibias.n420 commonsourceibias.n419 161.3
R24036 commonsourceibias.n417 commonsourceibias.n410 161.3
R24037 commonsourceibias.n416 commonsourceibias.n415 161.3
R24038 commonsourceibias.n414 commonsourceibias.n411 161.3
R24039 commonsourceibias.n570 commonsourceibias.n569 161.3
R24040 commonsourceibias.n568 commonsourceibias.n567 161.3
R24041 commonsourceibias.n566 commonsourceibias.n516 161.3
R24042 commonsourceibias.n565 commonsourceibias.n564 161.3
R24043 commonsourceibias.n563 commonsourceibias.n562 161.3
R24044 commonsourceibias.n561 commonsourceibias.n518 161.3
R24045 commonsourceibias.n560 commonsourceibias.n559 161.3
R24046 commonsourceibias.n558 commonsourceibias.n557 161.3
R24047 commonsourceibias.n556 commonsourceibias.n520 161.3
R24048 commonsourceibias.n554 commonsourceibias.n553 161.3
R24049 commonsourceibias.n552 commonsourceibias.n521 161.3
R24050 commonsourceibias.n551 commonsourceibias.n550 161.3
R24051 commonsourceibias.n548 commonsourceibias.n522 161.3
R24052 commonsourceibias.n547 commonsourceibias.n546 161.3
R24053 commonsourceibias.n545 commonsourceibias.n523 161.3
R24054 commonsourceibias.n544 commonsourceibias.n543 161.3
R24055 commonsourceibias.n541 commonsourceibias.n524 161.3
R24056 commonsourceibias.n539 commonsourceibias.n538 161.3
R24057 commonsourceibias.n537 commonsourceibias.n525 161.3
R24058 commonsourceibias.n536 commonsourceibias.n535 161.3
R24059 commonsourceibias.n533 commonsourceibias.n526 161.3
R24060 commonsourceibias.n532 commonsourceibias.n531 161.3
R24061 commonsourceibias.n530 commonsourceibias.n527 161.3
R24062 commonsourceibias.n615 commonsourceibias.n367 161.3
R24063 commonsourceibias.n613 commonsourceibias.n612 161.3
R24064 commonsourceibias.n611 commonsourceibias.n368 161.3
R24065 commonsourceibias.n610 commonsourceibias.n609 161.3
R24066 commonsourceibias.n607 commonsourceibias.n369 161.3
R24067 commonsourceibias.n606 commonsourceibias.n605 161.3
R24068 commonsourceibias.n604 commonsourceibias.n370 161.3
R24069 commonsourceibias.n603 commonsourceibias.n602 161.3
R24070 commonsourceibias.n600 commonsourceibias.n371 161.3
R24071 commonsourceibias.n598 commonsourceibias.n597 161.3
R24072 commonsourceibias.n596 commonsourceibias.n372 161.3
R24073 commonsourceibias.n595 commonsourceibias.n594 161.3
R24074 commonsourceibias.n592 commonsourceibias.n373 161.3
R24075 commonsourceibias.n591 commonsourceibias.n590 161.3
R24076 commonsourceibias.n589 commonsourceibias.n374 161.3
R24077 commonsourceibias.n588 commonsourceibias.n587 161.3
R24078 commonsourceibias.n585 commonsourceibias.n375 161.3
R24079 commonsourceibias.n583 commonsourceibias.n582 161.3
R24080 commonsourceibias.n581 commonsourceibias.n376 161.3
R24081 commonsourceibias.n580 commonsourceibias.n579 161.3
R24082 commonsourceibias.n577 commonsourceibias.n377 161.3
R24083 commonsourceibias.n576 commonsourceibias.n575 161.3
R24084 commonsourceibias.n574 commonsourceibias.n378 161.3
R24085 commonsourceibias.n573 commonsourceibias.n572 161.3
R24086 commonsourceibias.n141 commonsourceibias.n139 81.5057
R24087 commonsourceibias.n381 commonsourceibias.n379 81.5057
R24088 commonsourceibias.n141 commonsourceibias.n140 80.9324
R24089 commonsourceibias.n143 commonsourceibias.n142 80.9324
R24090 commonsourceibias.n145 commonsourceibias.n144 80.9324
R24091 commonsourceibias.n147 commonsourceibias.n146 80.9324
R24092 commonsourceibias.n138 commonsourceibias.n137 80.9324
R24093 commonsourceibias.n136 commonsourceibias.n135 80.9324
R24094 commonsourceibias.n134 commonsourceibias.n133 80.9324
R24095 commonsourceibias.n132 commonsourceibias.n131 80.9324
R24096 commonsourceibias.n130 commonsourceibias.n129 80.9324
R24097 commonsourceibias.n504 commonsourceibias.n503 80.9324
R24098 commonsourceibias.n506 commonsourceibias.n505 80.9324
R24099 commonsourceibias.n508 commonsourceibias.n507 80.9324
R24100 commonsourceibias.n510 commonsourceibias.n509 80.9324
R24101 commonsourceibias.n512 commonsourceibias.n511 80.9324
R24102 commonsourceibias.n387 commonsourceibias.n386 80.9324
R24103 commonsourceibias.n385 commonsourceibias.n384 80.9324
R24104 commonsourceibias.n383 commonsourceibias.n382 80.9324
R24105 commonsourceibias.n381 commonsourceibias.n380 80.9324
R24106 commonsourceibias.n365 commonsourceibias.n364 80.6037
R24107 commonsourceibias.n128 commonsourceibias.n127 80.6037
R24108 commonsourceibias.n250 commonsourceibias.n249 80.6037
R24109 commonsourceibias.n732 commonsourceibias.n731 80.6037
R24110 commonsourceibias.n502 commonsourceibias.n501 80.6037
R24111 commonsourceibias.n617 commonsourceibias.n616 80.6037
R24112 commonsourceibias.n322 commonsourceibias.n321 56.5617
R24113 commonsourceibias.n336 commonsourceibias.n335 56.5617
R24114 commonsourceibias.n85 commonsourceibias.n84 56.5617
R24115 commonsourceibias.n71 commonsourceibias.n70 56.5617
R24116 commonsourceibias.n207 commonsourceibias.n206 56.5617
R24117 commonsourceibias.n193 commonsourceibias.n192 56.5617
R24118 commonsourceibias.n687 commonsourceibias.n685 56.5617
R24119 commonsourceibias.n702 commonsourceibias.n700 56.5617
R24120 commonsourceibias.n457 commonsourceibias.n455 56.5617
R24121 commonsourceibias.n472 commonsourceibias.n470 56.5617
R24122 commonsourceibias.n572 commonsourceibias.n570 56.5617
R24123 commonsourceibias.n294 commonsourceibias.n293 56.5617
R24124 commonsourceibias.n308 commonsourceibias.n307 56.5617
R24125 commonsourceibias.n350 commonsourceibias.n349 56.5617
R24126 commonsourceibias.n113 commonsourceibias.n112 56.5617
R24127 commonsourceibias.n99 commonsourceibias.n98 56.5617
R24128 commonsourceibias.n57 commonsourceibias.n56 56.5617
R24129 commonsourceibias.n235 commonsourceibias.n234 56.5617
R24130 commonsourceibias.n221 commonsourceibias.n220 56.5617
R24131 commonsourceibias.n179 commonsourceibias.n178 56.5617
R24132 commonsourceibias.n657 commonsourceibias.n655 56.5617
R24133 commonsourceibias.n672 commonsourceibias.n670 56.5617
R24134 commonsourceibias.n717 commonsourceibias.n715 56.5617
R24135 commonsourceibias.n427 commonsourceibias.n425 56.5617
R24136 commonsourceibias.n442 commonsourceibias.n440 56.5617
R24137 commonsourceibias.n487 commonsourceibias.n485 56.5617
R24138 commonsourceibias.n602 commonsourceibias.n600 56.5617
R24139 commonsourceibias.n587 commonsourceibias.n585 56.5617
R24140 commonsourceibias.n543 commonsourceibias.n541 56.5617
R24141 commonsourceibias.n557 commonsourceibias.n556 56.5617
R24142 commonsourceibias.n285 commonsourceibias.n284 51.2335
R24143 commonsourceibias.n357 commonsourceibias.n252 51.2335
R24144 commonsourceibias.n120 commonsourceibias.n15 51.2335
R24145 commonsourceibias.n48 commonsourceibias.n47 51.2335
R24146 commonsourceibias.n242 commonsourceibias.n1 51.2335
R24147 commonsourceibias.n170 commonsourceibias.n169 51.2335
R24148 commonsourceibias.n647 commonsourceibias.n646 51.2335
R24149 commonsourceibias.n724 commonsourceibias.n619 51.2335
R24150 commonsourceibias.n417 commonsourceibias.n416 51.2335
R24151 commonsourceibias.n494 commonsourceibias.n389 51.2335
R24152 commonsourceibias.n609 commonsourceibias.n368 51.2335
R24153 commonsourceibias.n533 commonsourceibias.n532 51.2335
R24154 commonsourceibias.n364 commonsourceibias.n363 50.9056
R24155 commonsourceibias.n127 commonsourceibias.n126 50.9056
R24156 commonsourceibias.n249 commonsourceibias.n248 50.9056
R24157 commonsourceibias.n731 commonsourceibias.n730 50.9056
R24158 commonsourceibias.n501 commonsourceibias.n500 50.9056
R24159 commonsourceibias.n616 commonsourceibias.n615 50.9056
R24160 commonsourceibias.n299 commonsourceibias.n298 50.2647
R24161 commonsourceibias.n343 commonsourceibias.n257 50.2647
R24162 commonsourceibias.n106 commonsourceibias.n20 50.2647
R24163 commonsourceibias.n62 commonsourceibias.n61 50.2647
R24164 commonsourceibias.n228 commonsourceibias.n6 50.2647
R24165 commonsourceibias.n184 commonsourceibias.n183 50.2647
R24166 commonsourceibias.n662 commonsourceibias.n661 50.2647
R24167 commonsourceibias.n709 commonsourceibias.n623 50.2647
R24168 commonsourceibias.n432 commonsourceibias.n431 50.2647
R24169 commonsourceibias.n479 commonsourceibias.n393 50.2647
R24170 commonsourceibias.n594 commonsourceibias.n372 50.2647
R24171 commonsourceibias.n548 commonsourceibias.n547 50.2647
R24172 commonsourceibias.n281 commonsourceibias.n280 49.9027
R24173 commonsourceibias.n44 commonsourceibias.n43 49.9027
R24174 commonsourceibias.n166 commonsourceibias.n165 49.9027
R24175 commonsourceibias.n643 commonsourceibias.n642 49.9027
R24176 commonsourceibias.n413 commonsourceibias.n412 49.9027
R24177 commonsourceibias.n529 commonsourceibias.n528 49.9027
R24178 commonsourceibias.n313 commonsourceibias.n312 49.296
R24179 commonsourceibias.n329 commonsourceibias.n262 49.296
R24180 commonsourceibias.n92 commonsourceibias.n25 49.296
R24181 commonsourceibias.n76 commonsourceibias.n75 49.296
R24182 commonsourceibias.n214 commonsourceibias.n11 49.296
R24183 commonsourceibias.n198 commonsourceibias.n197 49.296
R24184 commonsourceibias.n677 commonsourceibias.n676 49.296
R24185 commonsourceibias.n694 commonsourceibias.n627 49.296
R24186 commonsourceibias.n447 commonsourceibias.n446 49.296
R24187 commonsourceibias.n464 commonsourceibias.n397 49.296
R24188 commonsourceibias.n579 commonsourceibias.n376 49.296
R24189 commonsourceibias.n562 commonsourceibias.n561 49.296
R24190 commonsourceibias.n315 commonsourceibias.n267 48.3272
R24191 commonsourceibias.n327 commonsourceibias.n326 48.3272
R24192 commonsourceibias.n90 commonsourceibias.n89 48.3272
R24193 commonsourceibias.n78 commonsourceibias.n30 48.3272
R24194 commonsourceibias.n212 commonsourceibias.n211 48.3272
R24195 commonsourceibias.n202 commonsourceibias.n201 48.3272
R24196 commonsourceibias.n679 commonsourceibias.n631 48.3272
R24197 commonsourceibias.n692 commonsourceibias.n691 48.3272
R24198 commonsourceibias.n449 commonsourceibias.n401 48.3272
R24199 commonsourceibias.n462 commonsourceibias.n461 48.3272
R24200 commonsourceibias.n577 commonsourceibias.n576 48.3272
R24201 commonsourceibias.n566 commonsourceibias.n565 48.3272
R24202 commonsourceibias.n301 commonsourceibias.n272 47.3584
R24203 commonsourceibias.n341 commonsourceibias.n340 47.3584
R24204 commonsourceibias.n104 commonsourceibias.n103 47.3584
R24205 commonsourceibias.n64 commonsourceibias.n35 47.3584
R24206 commonsourceibias.n226 commonsourceibias.n225 47.3584
R24207 commonsourceibias.n186 commonsourceibias.n157 47.3584
R24208 commonsourceibias.n664 commonsourceibias.n635 47.3584
R24209 commonsourceibias.n707 commonsourceibias.n706 47.3584
R24210 commonsourceibias.n434 commonsourceibias.n405 47.3584
R24211 commonsourceibias.n477 commonsourceibias.n476 47.3584
R24212 commonsourceibias.n592 commonsourceibias.n591 47.3584
R24213 commonsourceibias.n550 commonsourceibias.n521 47.3584
R24214 commonsourceibias.n287 commonsourceibias.n277 46.3896
R24215 commonsourceibias.n355 commonsourceibias.n354 46.3896
R24216 commonsourceibias.n118 commonsourceibias.n117 46.3896
R24217 commonsourceibias.n50 commonsourceibias.n40 46.3896
R24218 commonsourceibias.n240 commonsourceibias.n239 46.3896
R24219 commonsourceibias.n172 commonsourceibias.n162 46.3896
R24220 commonsourceibias.n649 commonsourceibias.n639 46.3896
R24221 commonsourceibias.n722 commonsourceibias.n721 46.3896
R24222 commonsourceibias.n419 commonsourceibias.n409 46.3896
R24223 commonsourceibias.n492 commonsourceibias.n491 46.3896
R24224 commonsourceibias.n607 commonsourceibias.n606 46.3896
R24225 commonsourceibias.n535 commonsourceibias.n525 46.3896
R24226 commonsourceibias.n282 commonsourceibias.n281 44.7059
R24227 commonsourceibias.n644 commonsourceibias.n643 44.7059
R24228 commonsourceibias.n414 commonsourceibias.n413 44.7059
R24229 commonsourceibias.n530 commonsourceibias.n529 44.7059
R24230 commonsourceibias.n45 commonsourceibias.n44 44.7059
R24231 commonsourceibias.n167 commonsourceibias.n166 44.7059
R24232 commonsourceibias.n291 commonsourceibias.n277 34.7644
R24233 commonsourceibias.n354 commonsourceibias.n254 34.7644
R24234 commonsourceibias.n117 commonsourceibias.n17 34.7644
R24235 commonsourceibias.n54 commonsourceibias.n40 34.7644
R24236 commonsourceibias.n239 commonsourceibias.n3 34.7644
R24237 commonsourceibias.n176 commonsourceibias.n162 34.7644
R24238 commonsourceibias.n653 commonsourceibias.n639 34.7644
R24239 commonsourceibias.n721 commonsourceibias.n621 34.7644
R24240 commonsourceibias.n423 commonsourceibias.n409 34.7644
R24241 commonsourceibias.n491 commonsourceibias.n391 34.7644
R24242 commonsourceibias.n606 commonsourceibias.n370 34.7644
R24243 commonsourceibias.n539 commonsourceibias.n525 34.7644
R24244 commonsourceibias.n305 commonsourceibias.n272 33.7956
R24245 commonsourceibias.n340 commonsourceibias.n259 33.7956
R24246 commonsourceibias.n103 commonsourceibias.n22 33.7956
R24247 commonsourceibias.n68 commonsourceibias.n35 33.7956
R24248 commonsourceibias.n225 commonsourceibias.n8 33.7956
R24249 commonsourceibias.n190 commonsourceibias.n157 33.7956
R24250 commonsourceibias.n668 commonsourceibias.n635 33.7956
R24251 commonsourceibias.n706 commonsourceibias.n625 33.7956
R24252 commonsourceibias.n438 commonsourceibias.n405 33.7956
R24253 commonsourceibias.n476 commonsourceibias.n395 33.7956
R24254 commonsourceibias.n591 commonsourceibias.n374 33.7956
R24255 commonsourceibias.n554 commonsourceibias.n521 33.7956
R24256 commonsourceibias.n319 commonsourceibias.n267 32.8269
R24257 commonsourceibias.n326 commonsourceibias.n264 32.8269
R24258 commonsourceibias.n89 commonsourceibias.n27 32.8269
R24259 commonsourceibias.n82 commonsourceibias.n30 32.8269
R24260 commonsourceibias.n211 commonsourceibias.n13 32.8269
R24261 commonsourceibias.n203 commonsourceibias.n202 32.8269
R24262 commonsourceibias.n683 commonsourceibias.n631 32.8269
R24263 commonsourceibias.n691 commonsourceibias.n629 32.8269
R24264 commonsourceibias.n453 commonsourceibias.n401 32.8269
R24265 commonsourceibias.n461 commonsourceibias.n399 32.8269
R24266 commonsourceibias.n576 commonsourceibias.n378 32.8269
R24267 commonsourceibias.n567 commonsourceibias.n566 32.8269
R24268 commonsourceibias.n312 commonsourceibias.n269 31.8581
R24269 commonsourceibias.n333 commonsourceibias.n262 31.8581
R24270 commonsourceibias.n96 commonsourceibias.n25 31.8581
R24271 commonsourceibias.n75 commonsourceibias.n32 31.8581
R24272 commonsourceibias.n218 commonsourceibias.n11 31.8581
R24273 commonsourceibias.n197 commonsourceibias.n196 31.8581
R24274 commonsourceibias.n676 commonsourceibias.n633 31.8581
R24275 commonsourceibias.n698 commonsourceibias.n627 31.8581
R24276 commonsourceibias.n446 commonsourceibias.n403 31.8581
R24277 commonsourceibias.n468 commonsourceibias.n397 31.8581
R24278 commonsourceibias.n583 commonsourceibias.n376 31.8581
R24279 commonsourceibias.n561 commonsourceibias.n560 31.8581
R24280 commonsourceibias.n298 commonsourceibias.n274 30.8893
R24281 commonsourceibias.n347 commonsourceibias.n257 30.8893
R24282 commonsourceibias.n110 commonsourceibias.n20 30.8893
R24283 commonsourceibias.n61 commonsourceibias.n37 30.8893
R24284 commonsourceibias.n232 commonsourceibias.n6 30.8893
R24285 commonsourceibias.n183 commonsourceibias.n159 30.8893
R24286 commonsourceibias.n661 commonsourceibias.n637 30.8893
R24287 commonsourceibias.n713 commonsourceibias.n623 30.8893
R24288 commonsourceibias.n431 commonsourceibias.n407 30.8893
R24289 commonsourceibias.n483 commonsourceibias.n393 30.8893
R24290 commonsourceibias.n598 commonsourceibias.n372 30.8893
R24291 commonsourceibias.n547 commonsourceibias.n523 30.8893
R24292 commonsourceibias.n284 commonsourceibias.n279 29.9206
R24293 commonsourceibias.n361 commonsourceibias.n252 29.9206
R24294 commonsourceibias.n124 commonsourceibias.n15 29.9206
R24295 commonsourceibias.n47 commonsourceibias.n42 29.9206
R24296 commonsourceibias.n246 commonsourceibias.n1 29.9206
R24297 commonsourceibias.n169 commonsourceibias.n164 29.9206
R24298 commonsourceibias.n646 commonsourceibias.n641 29.9206
R24299 commonsourceibias.n728 commonsourceibias.n619 29.9206
R24300 commonsourceibias.n416 commonsourceibias.n411 29.9206
R24301 commonsourceibias.n498 commonsourceibias.n389 29.9206
R24302 commonsourceibias.n613 commonsourceibias.n368 29.9206
R24303 commonsourceibias.n532 commonsourceibias.n527 29.9206
R24304 commonsourceibias.n363 commonsourceibias.n362 21.8872
R24305 commonsourceibias.n126 commonsourceibias.n125 21.8872
R24306 commonsourceibias.n248 commonsourceibias.n247 21.8872
R24307 commonsourceibias.n730 commonsourceibias.n729 21.8872
R24308 commonsourceibias.n500 commonsourceibias.n499 21.8872
R24309 commonsourceibias.n615 commonsourceibias.n614 21.8872
R24310 commonsourceibias.n294 commonsourceibias.n276 21.3954
R24311 commonsourceibias.n349 commonsourceibias.n348 21.3954
R24312 commonsourceibias.n112 commonsourceibias.n111 21.3954
R24313 commonsourceibias.n57 commonsourceibias.n39 21.3954
R24314 commonsourceibias.n234 commonsourceibias.n233 21.3954
R24315 commonsourceibias.n179 commonsourceibias.n161 21.3954
R24316 commonsourceibias.n657 commonsourceibias.n656 21.3954
R24317 commonsourceibias.n715 commonsourceibias.n714 21.3954
R24318 commonsourceibias.n427 commonsourceibias.n426 21.3954
R24319 commonsourceibias.n485 commonsourceibias.n484 21.3954
R24320 commonsourceibias.n600 commonsourceibias.n599 21.3954
R24321 commonsourceibias.n543 commonsourceibias.n542 21.3954
R24322 commonsourceibias.n308 commonsourceibias.n271 20.9036
R24323 commonsourceibias.n335 commonsourceibias.n334 20.9036
R24324 commonsourceibias.n98 commonsourceibias.n97 20.9036
R24325 commonsourceibias.n71 commonsourceibias.n34 20.9036
R24326 commonsourceibias.n220 commonsourceibias.n219 20.9036
R24327 commonsourceibias.n193 commonsourceibias.n155 20.9036
R24328 commonsourceibias.n672 commonsourceibias.n671 20.9036
R24329 commonsourceibias.n700 commonsourceibias.n699 20.9036
R24330 commonsourceibias.n442 commonsourceibias.n441 20.9036
R24331 commonsourceibias.n470 commonsourceibias.n469 20.9036
R24332 commonsourceibias.n585 commonsourceibias.n584 20.9036
R24333 commonsourceibias.n557 commonsourceibias.n519 20.9036
R24334 commonsourceibias.n321 commonsourceibias.n320 20.4117
R24335 commonsourceibias.n322 commonsourceibias.n266 20.4117
R24336 commonsourceibias.n85 commonsourceibias.n29 20.4117
R24337 commonsourceibias.n84 commonsourceibias.n83 20.4117
R24338 commonsourceibias.n207 commonsourceibias.n150 20.4117
R24339 commonsourceibias.n206 commonsourceibias.n151 20.4117
R24340 commonsourceibias.n685 commonsourceibias.n684 20.4117
R24341 commonsourceibias.n687 commonsourceibias.n686 20.4117
R24342 commonsourceibias.n455 commonsourceibias.n454 20.4117
R24343 commonsourceibias.n457 commonsourceibias.n456 20.4117
R24344 commonsourceibias.n572 commonsourceibias.n571 20.4117
R24345 commonsourceibias.n570 commonsourceibias.n515 20.4117
R24346 commonsourceibias.n307 commonsourceibias.n306 19.9199
R24347 commonsourceibias.n336 commonsourceibias.n261 19.9199
R24348 commonsourceibias.n99 commonsourceibias.n24 19.9199
R24349 commonsourceibias.n70 commonsourceibias.n69 19.9199
R24350 commonsourceibias.n221 commonsourceibias.n10 19.9199
R24351 commonsourceibias.n192 commonsourceibias.n191 19.9199
R24352 commonsourceibias.n670 commonsourceibias.n669 19.9199
R24353 commonsourceibias.n702 commonsourceibias.n701 19.9199
R24354 commonsourceibias.n440 commonsourceibias.n439 19.9199
R24355 commonsourceibias.n472 commonsourceibias.n471 19.9199
R24356 commonsourceibias.n587 commonsourceibias.n586 19.9199
R24357 commonsourceibias.n556 commonsourceibias.n555 19.9199
R24358 commonsourceibias.n293 commonsourceibias.n292 19.4281
R24359 commonsourceibias.n350 commonsourceibias.n256 19.4281
R24360 commonsourceibias.n113 commonsourceibias.n19 19.4281
R24361 commonsourceibias.n56 commonsourceibias.n55 19.4281
R24362 commonsourceibias.n235 commonsourceibias.n5 19.4281
R24363 commonsourceibias.n178 commonsourceibias.n177 19.4281
R24364 commonsourceibias.n655 commonsourceibias.n654 19.4281
R24365 commonsourceibias.n717 commonsourceibias.n716 19.4281
R24366 commonsourceibias.n425 commonsourceibias.n424 19.4281
R24367 commonsourceibias.n487 commonsourceibias.n486 19.4281
R24368 commonsourceibias.n602 commonsourceibias.n601 19.4281
R24369 commonsourceibias.n541 commonsourceibias.n540 19.4281
R24370 commonsourceibias.n286 commonsourceibias.n285 13.526
R24371 commonsourceibias.n357 commonsourceibias.n356 13.526
R24372 commonsourceibias.n120 commonsourceibias.n119 13.526
R24373 commonsourceibias.n49 commonsourceibias.n48 13.526
R24374 commonsourceibias.n242 commonsourceibias.n241 13.526
R24375 commonsourceibias.n171 commonsourceibias.n170 13.526
R24376 commonsourceibias.n648 commonsourceibias.n647 13.526
R24377 commonsourceibias.n724 commonsourceibias.n723 13.526
R24378 commonsourceibias.n418 commonsourceibias.n417 13.526
R24379 commonsourceibias.n494 commonsourceibias.n493 13.526
R24380 commonsourceibias.n609 commonsourceibias.n608 13.526
R24381 commonsourceibias.n534 commonsourceibias.n533 13.526
R24382 commonsourceibias.n130 commonsourceibias.n128 13.2322
R24383 commonsourceibias.n504 commonsourceibias.n502 13.2322
R24384 commonsourceibias.n300 commonsourceibias.n299 13.0342
R24385 commonsourceibias.n343 commonsourceibias.n342 13.0342
R24386 commonsourceibias.n106 commonsourceibias.n105 13.0342
R24387 commonsourceibias.n63 commonsourceibias.n62 13.0342
R24388 commonsourceibias.n228 commonsourceibias.n227 13.0342
R24389 commonsourceibias.n185 commonsourceibias.n184 13.0342
R24390 commonsourceibias.n663 commonsourceibias.n662 13.0342
R24391 commonsourceibias.n709 commonsourceibias.n708 13.0342
R24392 commonsourceibias.n433 commonsourceibias.n432 13.0342
R24393 commonsourceibias.n479 commonsourceibias.n478 13.0342
R24394 commonsourceibias.n594 commonsourceibias.n593 13.0342
R24395 commonsourceibias.n549 commonsourceibias.n548 13.0342
R24396 commonsourceibias.n314 commonsourceibias.n313 12.5423
R24397 commonsourceibias.n329 commonsourceibias.n328 12.5423
R24398 commonsourceibias.n92 commonsourceibias.n91 12.5423
R24399 commonsourceibias.n77 commonsourceibias.n76 12.5423
R24400 commonsourceibias.n214 commonsourceibias.n213 12.5423
R24401 commonsourceibias.n198 commonsourceibias.n153 12.5423
R24402 commonsourceibias.n678 commonsourceibias.n677 12.5423
R24403 commonsourceibias.n694 commonsourceibias.n693 12.5423
R24404 commonsourceibias.n448 commonsourceibias.n447 12.5423
R24405 commonsourceibias.n464 commonsourceibias.n463 12.5423
R24406 commonsourceibias.n579 commonsourceibias.n578 12.5423
R24407 commonsourceibias.n562 commonsourceibias.n517 12.5423
R24408 commonsourceibias.n734 commonsourceibias.n366 12.2777
R24409 commonsourceibias.n315 commonsourceibias.n314 12.0505
R24410 commonsourceibias.n328 commonsourceibias.n327 12.0505
R24411 commonsourceibias.n91 commonsourceibias.n90 12.0505
R24412 commonsourceibias.n78 commonsourceibias.n77 12.0505
R24413 commonsourceibias.n213 commonsourceibias.n212 12.0505
R24414 commonsourceibias.n201 commonsourceibias.n153 12.0505
R24415 commonsourceibias.n679 commonsourceibias.n678 12.0505
R24416 commonsourceibias.n693 commonsourceibias.n692 12.0505
R24417 commonsourceibias.n449 commonsourceibias.n448 12.0505
R24418 commonsourceibias.n463 commonsourceibias.n462 12.0505
R24419 commonsourceibias.n578 commonsourceibias.n577 12.0505
R24420 commonsourceibias.n565 commonsourceibias.n517 12.0505
R24421 commonsourceibias.n301 commonsourceibias.n300 11.5587
R24422 commonsourceibias.n342 commonsourceibias.n341 11.5587
R24423 commonsourceibias.n105 commonsourceibias.n104 11.5587
R24424 commonsourceibias.n64 commonsourceibias.n63 11.5587
R24425 commonsourceibias.n227 commonsourceibias.n226 11.5587
R24426 commonsourceibias.n186 commonsourceibias.n185 11.5587
R24427 commonsourceibias.n664 commonsourceibias.n663 11.5587
R24428 commonsourceibias.n708 commonsourceibias.n707 11.5587
R24429 commonsourceibias.n434 commonsourceibias.n433 11.5587
R24430 commonsourceibias.n478 commonsourceibias.n477 11.5587
R24431 commonsourceibias.n593 commonsourceibias.n592 11.5587
R24432 commonsourceibias.n550 commonsourceibias.n549 11.5587
R24433 commonsourceibias.n287 commonsourceibias.n286 11.0668
R24434 commonsourceibias.n356 commonsourceibias.n355 11.0668
R24435 commonsourceibias.n119 commonsourceibias.n118 11.0668
R24436 commonsourceibias.n50 commonsourceibias.n49 11.0668
R24437 commonsourceibias.n241 commonsourceibias.n240 11.0668
R24438 commonsourceibias.n172 commonsourceibias.n171 11.0668
R24439 commonsourceibias.n649 commonsourceibias.n648 11.0668
R24440 commonsourceibias.n723 commonsourceibias.n722 11.0668
R24441 commonsourceibias.n419 commonsourceibias.n418 11.0668
R24442 commonsourceibias.n493 commonsourceibias.n492 11.0668
R24443 commonsourceibias.n608 commonsourceibias.n607 11.0668
R24444 commonsourceibias.n535 commonsourceibias.n534 11.0668
R24445 commonsourceibias.n734 commonsourceibias.n733 10.3347
R24446 commonsourceibias.n149 commonsourceibias.n148 9.50363
R24447 commonsourceibias.n514 commonsourceibias.n513 9.50363
R24448 commonsourceibias.n366 commonsourceibias.n250 8.75852
R24449 commonsourceibias.n733 commonsourceibias.n617 8.75852
R24450 commonsourceibias.n292 commonsourceibias.n291 5.16479
R24451 commonsourceibias.n256 commonsourceibias.n254 5.16479
R24452 commonsourceibias.n19 commonsourceibias.n17 5.16479
R24453 commonsourceibias.n55 commonsourceibias.n54 5.16479
R24454 commonsourceibias.n5 commonsourceibias.n3 5.16479
R24455 commonsourceibias.n177 commonsourceibias.n176 5.16479
R24456 commonsourceibias.n654 commonsourceibias.n653 5.16479
R24457 commonsourceibias.n716 commonsourceibias.n621 5.16479
R24458 commonsourceibias.n424 commonsourceibias.n423 5.16479
R24459 commonsourceibias.n486 commonsourceibias.n391 5.16479
R24460 commonsourceibias.n601 commonsourceibias.n370 5.16479
R24461 commonsourceibias.n540 commonsourceibias.n539 5.16479
R24462 commonsourceibias.n366 commonsourceibias.n365 5.03125
R24463 commonsourceibias.n733 commonsourceibias.n732 5.03125
R24464 commonsourceibias.n306 commonsourceibias.n305 4.67295
R24465 commonsourceibias.n261 commonsourceibias.n259 4.67295
R24466 commonsourceibias.n24 commonsourceibias.n22 4.67295
R24467 commonsourceibias.n69 commonsourceibias.n68 4.67295
R24468 commonsourceibias.n10 commonsourceibias.n8 4.67295
R24469 commonsourceibias.n191 commonsourceibias.n190 4.67295
R24470 commonsourceibias.n669 commonsourceibias.n668 4.67295
R24471 commonsourceibias.n701 commonsourceibias.n625 4.67295
R24472 commonsourceibias.n439 commonsourceibias.n438 4.67295
R24473 commonsourceibias.n471 commonsourceibias.n395 4.67295
R24474 commonsourceibias.n586 commonsourceibias.n374 4.67295
R24475 commonsourceibias.n555 commonsourceibias.n554 4.67295
R24476 commonsourceibias commonsourceibias.n734 4.20978
R24477 commonsourceibias.n320 commonsourceibias.n319 4.18111
R24478 commonsourceibias.n266 commonsourceibias.n264 4.18111
R24479 commonsourceibias.n29 commonsourceibias.n27 4.18111
R24480 commonsourceibias.n83 commonsourceibias.n82 4.18111
R24481 commonsourceibias.n150 commonsourceibias.n13 4.18111
R24482 commonsourceibias.n203 commonsourceibias.n151 4.18111
R24483 commonsourceibias.n684 commonsourceibias.n683 4.18111
R24484 commonsourceibias.n686 commonsourceibias.n629 4.18111
R24485 commonsourceibias.n454 commonsourceibias.n453 4.18111
R24486 commonsourceibias.n456 commonsourceibias.n399 4.18111
R24487 commonsourceibias.n571 commonsourceibias.n378 4.18111
R24488 commonsourceibias.n567 commonsourceibias.n515 4.18111
R24489 commonsourceibias.n271 commonsourceibias.n269 3.68928
R24490 commonsourceibias.n334 commonsourceibias.n333 3.68928
R24491 commonsourceibias.n97 commonsourceibias.n96 3.68928
R24492 commonsourceibias.n34 commonsourceibias.n32 3.68928
R24493 commonsourceibias.n219 commonsourceibias.n218 3.68928
R24494 commonsourceibias.n196 commonsourceibias.n155 3.68928
R24495 commonsourceibias.n671 commonsourceibias.n633 3.68928
R24496 commonsourceibias.n699 commonsourceibias.n698 3.68928
R24497 commonsourceibias.n441 commonsourceibias.n403 3.68928
R24498 commonsourceibias.n469 commonsourceibias.n468 3.68928
R24499 commonsourceibias.n584 commonsourceibias.n583 3.68928
R24500 commonsourceibias.n560 commonsourceibias.n519 3.68928
R24501 commonsourceibias.n276 commonsourceibias.n274 3.19744
R24502 commonsourceibias.n348 commonsourceibias.n347 3.19744
R24503 commonsourceibias.n111 commonsourceibias.n110 3.19744
R24504 commonsourceibias.n39 commonsourceibias.n37 3.19744
R24505 commonsourceibias.n233 commonsourceibias.n232 3.19744
R24506 commonsourceibias.n161 commonsourceibias.n159 3.19744
R24507 commonsourceibias.n656 commonsourceibias.n637 3.19744
R24508 commonsourceibias.n714 commonsourceibias.n713 3.19744
R24509 commonsourceibias.n426 commonsourceibias.n407 3.19744
R24510 commonsourceibias.n484 commonsourceibias.n483 3.19744
R24511 commonsourceibias.n599 commonsourceibias.n598 3.19744
R24512 commonsourceibias.n542 commonsourceibias.n523 3.19744
R24513 commonsourceibias.n139 commonsourceibias.t47 2.82907
R24514 commonsourceibias.n139 commonsourceibias.t79 2.82907
R24515 commonsourceibias.n140 commonsourceibias.t55 2.82907
R24516 commonsourceibias.n140 commonsourceibias.t5 2.82907
R24517 commonsourceibias.n142 commonsourceibias.t19 2.82907
R24518 commonsourceibias.n142 commonsourceibias.t23 2.82907
R24519 commonsourceibias.n144 commonsourceibias.t39 2.82907
R24520 commonsourceibias.n144 commonsourceibias.t71 2.82907
R24521 commonsourceibias.n146 commonsourceibias.t57 2.82907
R24522 commonsourceibias.n146 commonsourceibias.t27 2.82907
R24523 commonsourceibias.n137 commonsourceibias.t11 2.82907
R24524 commonsourceibias.n137 commonsourceibias.t41 2.82907
R24525 commonsourceibias.n135 commonsourceibias.t25 2.82907
R24526 commonsourceibias.n135 commonsourceibias.t35 2.82907
R24527 commonsourceibias.n133 commonsourceibias.t37 2.82907
R24528 commonsourceibias.n133 commonsourceibias.t77 2.82907
R24529 commonsourceibias.n131 commonsourceibias.t51 2.82907
R24530 commonsourceibias.n131 commonsourceibias.t9 2.82907
R24531 commonsourceibias.n129 commonsourceibias.t75 2.82907
R24532 commonsourceibias.n129 commonsourceibias.t21 2.82907
R24533 commonsourceibias.n503 commonsourceibias.t43 2.82907
R24534 commonsourceibias.n503 commonsourceibias.t15 2.82907
R24535 commonsourceibias.n505 commonsourceibias.t31 2.82907
R24536 commonsourceibias.n505 commonsourceibias.t1 2.82907
R24537 commonsourceibias.n507 commonsourceibias.t17 2.82907
R24538 commonsourceibias.n507 commonsourceibias.t61 2.82907
R24539 commonsourceibias.n509 commonsourceibias.t59 2.82907
R24540 commonsourceibias.n509 commonsourceibias.t45 2.82907
R24541 commonsourceibias.n511 commonsourceibias.t65 2.82907
R24542 commonsourceibias.n511 commonsourceibias.t33 2.82907
R24543 commonsourceibias.n386 commonsourceibias.t53 2.82907
R24544 commonsourceibias.n386 commonsourceibias.t73 2.82907
R24545 commonsourceibias.n384 commonsourceibias.t7 2.82907
R24546 commonsourceibias.n384 commonsourceibias.t63 2.82907
R24547 commonsourceibias.n382 commonsourceibias.t69 2.82907
R24548 commonsourceibias.n382 commonsourceibias.t67 2.82907
R24549 commonsourceibias.n380 commonsourceibias.t49 2.82907
R24550 commonsourceibias.n380 commonsourceibias.t13 2.82907
R24551 commonsourceibias.n379 commonsourceibias.t29 2.82907
R24552 commonsourceibias.n379 commonsourceibias.t3 2.82907
R24553 commonsourceibias.n280 commonsourceibias.n279 2.7056
R24554 commonsourceibias.n362 commonsourceibias.n361 2.7056
R24555 commonsourceibias.n125 commonsourceibias.n124 2.7056
R24556 commonsourceibias.n43 commonsourceibias.n42 2.7056
R24557 commonsourceibias.n247 commonsourceibias.n246 2.7056
R24558 commonsourceibias.n165 commonsourceibias.n164 2.7056
R24559 commonsourceibias.n642 commonsourceibias.n641 2.7056
R24560 commonsourceibias.n729 commonsourceibias.n728 2.7056
R24561 commonsourceibias.n412 commonsourceibias.n411 2.7056
R24562 commonsourceibias.n499 commonsourceibias.n498 2.7056
R24563 commonsourceibias.n614 commonsourceibias.n613 2.7056
R24564 commonsourceibias.n528 commonsourceibias.n527 2.7056
R24565 commonsourceibias.n132 commonsourceibias.n130 0.573776
R24566 commonsourceibias.n134 commonsourceibias.n132 0.573776
R24567 commonsourceibias.n136 commonsourceibias.n134 0.573776
R24568 commonsourceibias.n138 commonsourceibias.n136 0.573776
R24569 commonsourceibias.n147 commonsourceibias.n145 0.573776
R24570 commonsourceibias.n145 commonsourceibias.n143 0.573776
R24571 commonsourceibias.n143 commonsourceibias.n141 0.573776
R24572 commonsourceibias.n383 commonsourceibias.n381 0.573776
R24573 commonsourceibias.n385 commonsourceibias.n383 0.573776
R24574 commonsourceibias.n387 commonsourceibias.n385 0.573776
R24575 commonsourceibias.n512 commonsourceibias.n510 0.573776
R24576 commonsourceibias.n510 commonsourceibias.n508 0.573776
R24577 commonsourceibias.n508 commonsourceibias.n506 0.573776
R24578 commonsourceibias.n506 commonsourceibias.n504 0.573776
R24579 commonsourceibias.n148 commonsourceibias.n138 0.287138
R24580 commonsourceibias.n148 commonsourceibias.n147 0.287138
R24581 commonsourceibias.n513 commonsourceibias.n387 0.287138
R24582 commonsourceibias.n513 commonsourceibias.n512 0.287138
R24583 commonsourceibias.n365 commonsourceibias.n251 0.285035
R24584 commonsourceibias.n128 commonsourceibias.n14 0.285035
R24585 commonsourceibias.n250 commonsourceibias.n0 0.285035
R24586 commonsourceibias.n732 commonsourceibias.n618 0.285035
R24587 commonsourceibias.n502 commonsourceibias.n388 0.285035
R24588 commonsourceibias.n617 commonsourceibias.n367 0.285035
R24589 commonsourceibias.n360 commonsourceibias.n251 0.189894
R24590 commonsourceibias.n360 commonsourceibias.n359 0.189894
R24591 commonsourceibias.n359 commonsourceibias.n358 0.189894
R24592 commonsourceibias.n358 commonsourceibias.n253 0.189894
R24593 commonsourceibias.n353 commonsourceibias.n253 0.189894
R24594 commonsourceibias.n353 commonsourceibias.n352 0.189894
R24595 commonsourceibias.n352 commonsourceibias.n351 0.189894
R24596 commonsourceibias.n351 commonsourceibias.n255 0.189894
R24597 commonsourceibias.n346 commonsourceibias.n255 0.189894
R24598 commonsourceibias.n346 commonsourceibias.n345 0.189894
R24599 commonsourceibias.n345 commonsourceibias.n344 0.189894
R24600 commonsourceibias.n344 commonsourceibias.n258 0.189894
R24601 commonsourceibias.n339 commonsourceibias.n258 0.189894
R24602 commonsourceibias.n339 commonsourceibias.n338 0.189894
R24603 commonsourceibias.n338 commonsourceibias.n337 0.189894
R24604 commonsourceibias.n337 commonsourceibias.n260 0.189894
R24605 commonsourceibias.n332 commonsourceibias.n260 0.189894
R24606 commonsourceibias.n332 commonsourceibias.n331 0.189894
R24607 commonsourceibias.n331 commonsourceibias.n330 0.189894
R24608 commonsourceibias.n330 commonsourceibias.n263 0.189894
R24609 commonsourceibias.n325 commonsourceibias.n263 0.189894
R24610 commonsourceibias.n325 commonsourceibias.n324 0.189894
R24611 commonsourceibias.n324 commonsourceibias.n323 0.189894
R24612 commonsourceibias.n323 commonsourceibias.n265 0.189894
R24613 commonsourceibias.n318 commonsourceibias.n265 0.189894
R24614 commonsourceibias.n318 commonsourceibias.n317 0.189894
R24615 commonsourceibias.n317 commonsourceibias.n316 0.189894
R24616 commonsourceibias.n316 commonsourceibias.n268 0.189894
R24617 commonsourceibias.n311 commonsourceibias.n268 0.189894
R24618 commonsourceibias.n311 commonsourceibias.n310 0.189894
R24619 commonsourceibias.n310 commonsourceibias.n309 0.189894
R24620 commonsourceibias.n309 commonsourceibias.n270 0.189894
R24621 commonsourceibias.n304 commonsourceibias.n270 0.189894
R24622 commonsourceibias.n304 commonsourceibias.n303 0.189894
R24623 commonsourceibias.n303 commonsourceibias.n302 0.189894
R24624 commonsourceibias.n302 commonsourceibias.n273 0.189894
R24625 commonsourceibias.n297 commonsourceibias.n273 0.189894
R24626 commonsourceibias.n297 commonsourceibias.n296 0.189894
R24627 commonsourceibias.n296 commonsourceibias.n295 0.189894
R24628 commonsourceibias.n295 commonsourceibias.n275 0.189894
R24629 commonsourceibias.n290 commonsourceibias.n275 0.189894
R24630 commonsourceibias.n290 commonsourceibias.n289 0.189894
R24631 commonsourceibias.n289 commonsourceibias.n288 0.189894
R24632 commonsourceibias.n288 commonsourceibias.n278 0.189894
R24633 commonsourceibias.n283 commonsourceibias.n278 0.189894
R24634 commonsourceibias.n283 commonsourceibias.n282 0.189894
R24635 commonsourceibias.n123 commonsourceibias.n14 0.189894
R24636 commonsourceibias.n123 commonsourceibias.n122 0.189894
R24637 commonsourceibias.n122 commonsourceibias.n121 0.189894
R24638 commonsourceibias.n121 commonsourceibias.n16 0.189894
R24639 commonsourceibias.n116 commonsourceibias.n16 0.189894
R24640 commonsourceibias.n116 commonsourceibias.n115 0.189894
R24641 commonsourceibias.n115 commonsourceibias.n114 0.189894
R24642 commonsourceibias.n114 commonsourceibias.n18 0.189894
R24643 commonsourceibias.n109 commonsourceibias.n18 0.189894
R24644 commonsourceibias.n109 commonsourceibias.n108 0.189894
R24645 commonsourceibias.n108 commonsourceibias.n107 0.189894
R24646 commonsourceibias.n107 commonsourceibias.n21 0.189894
R24647 commonsourceibias.n102 commonsourceibias.n21 0.189894
R24648 commonsourceibias.n102 commonsourceibias.n101 0.189894
R24649 commonsourceibias.n101 commonsourceibias.n100 0.189894
R24650 commonsourceibias.n100 commonsourceibias.n23 0.189894
R24651 commonsourceibias.n95 commonsourceibias.n23 0.189894
R24652 commonsourceibias.n95 commonsourceibias.n94 0.189894
R24653 commonsourceibias.n94 commonsourceibias.n93 0.189894
R24654 commonsourceibias.n93 commonsourceibias.n26 0.189894
R24655 commonsourceibias.n88 commonsourceibias.n26 0.189894
R24656 commonsourceibias.n88 commonsourceibias.n87 0.189894
R24657 commonsourceibias.n87 commonsourceibias.n86 0.189894
R24658 commonsourceibias.n86 commonsourceibias.n28 0.189894
R24659 commonsourceibias.n81 commonsourceibias.n28 0.189894
R24660 commonsourceibias.n81 commonsourceibias.n80 0.189894
R24661 commonsourceibias.n80 commonsourceibias.n79 0.189894
R24662 commonsourceibias.n79 commonsourceibias.n31 0.189894
R24663 commonsourceibias.n74 commonsourceibias.n31 0.189894
R24664 commonsourceibias.n74 commonsourceibias.n73 0.189894
R24665 commonsourceibias.n73 commonsourceibias.n72 0.189894
R24666 commonsourceibias.n72 commonsourceibias.n33 0.189894
R24667 commonsourceibias.n67 commonsourceibias.n33 0.189894
R24668 commonsourceibias.n67 commonsourceibias.n66 0.189894
R24669 commonsourceibias.n66 commonsourceibias.n65 0.189894
R24670 commonsourceibias.n65 commonsourceibias.n36 0.189894
R24671 commonsourceibias.n60 commonsourceibias.n36 0.189894
R24672 commonsourceibias.n60 commonsourceibias.n59 0.189894
R24673 commonsourceibias.n59 commonsourceibias.n58 0.189894
R24674 commonsourceibias.n58 commonsourceibias.n38 0.189894
R24675 commonsourceibias.n53 commonsourceibias.n38 0.189894
R24676 commonsourceibias.n53 commonsourceibias.n52 0.189894
R24677 commonsourceibias.n52 commonsourceibias.n51 0.189894
R24678 commonsourceibias.n51 commonsourceibias.n41 0.189894
R24679 commonsourceibias.n46 commonsourceibias.n41 0.189894
R24680 commonsourceibias.n46 commonsourceibias.n45 0.189894
R24681 commonsourceibias.n205 commonsourceibias.n204 0.189894
R24682 commonsourceibias.n204 commonsourceibias.n152 0.189894
R24683 commonsourceibias.n200 commonsourceibias.n152 0.189894
R24684 commonsourceibias.n200 commonsourceibias.n199 0.189894
R24685 commonsourceibias.n199 commonsourceibias.n154 0.189894
R24686 commonsourceibias.n195 commonsourceibias.n154 0.189894
R24687 commonsourceibias.n195 commonsourceibias.n194 0.189894
R24688 commonsourceibias.n194 commonsourceibias.n156 0.189894
R24689 commonsourceibias.n189 commonsourceibias.n156 0.189894
R24690 commonsourceibias.n189 commonsourceibias.n188 0.189894
R24691 commonsourceibias.n188 commonsourceibias.n187 0.189894
R24692 commonsourceibias.n187 commonsourceibias.n158 0.189894
R24693 commonsourceibias.n182 commonsourceibias.n158 0.189894
R24694 commonsourceibias.n182 commonsourceibias.n181 0.189894
R24695 commonsourceibias.n181 commonsourceibias.n180 0.189894
R24696 commonsourceibias.n180 commonsourceibias.n160 0.189894
R24697 commonsourceibias.n175 commonsourceibias.n160 0.189894
R24698 commonsourceibias.n175 commonsourceibias.n174 0.189894
R24699 commonsourceibias.n174 commonsourceibias.n173 0.189894
R24700 commonsourceibias.n173 commonsourceibias.n163 0.189894
R24701 commonsourceibias.n168 commonsourceibias.n163 0.189894
R24702 commonsourceibias.n168 commonsourceibias.n167 0.189894
R24703 commonsourceibias.n245 commonsourceibias.n0 0.189894
R24704 commonsourceibias.n245 commonsourceibias.n244 0.189894
R24705 commonsourceibias.n244 commonsourceibias.n243 0.189894
R24706 commonsourceibias.n243 commonsourceibias.n2 0.189894
R24707 commonsourceibias.n238 commonsourceibias.n2 0.189894
R24708 commonsourceibias.n238 commonsourceibias.n237 0.189894
R24709 commonsourceibias.n237 commonsourceibias.n236 0.189894
R24710 commonsourceibias.n236 commonsourceibias.n4 0.189894
R24711 commonsourceibias.n231 commonsourceibias.n4 0.189894
R24712 commonsourceibias.n231 commonsourceibias.n230 0.189894
R24713 commonsourceibias.n230 commonsourceibias.n229 0.189894
R24714 commonsourceibias.n229 commonsourceibias.n7 0.189894
R24715 commonsourceibias.n224 commonsourceibias.n7 0.189894
R24716 commonsourceibias.n224 commonsourceibias.n223 0.189894
R24717 commonsourceibias.n223 commonsourceibias.n222 0.189894
R24718 commonsourceibias.n222 commonsourceibias.n9 0.189894
R24719 commonsourceibias.n217 commonsourceibias.n9 0.189894
R24720 commonsourceibias.n217 commonsourceibias.n216 0.189894
R24721 commonsourceibias.n216 commonsourceibias.n215 0.189894
R24722 commonsourceibias.n215 commonsourceibias.n12 0.189894
R24723 commonsourceibias.n210 commonsourceibias.n12 0.189894
R24724 commonsourceibias.n210 commonsourceibias.n209 0.189894
R24725 commonsourceibias.n209 commonsourceibias.n208 0.189894
R24726 commonsourceibias.n645 commonsourceibias.n644 0.189894
R24727 commonsourceibias.n645 commonsourceibias.n640 0.189894
R24728 commonsourceibias.n650 commonsourceibias.n640 0.189894
R24729 commonsourceibias.n651 commonsourceibias.n650 0.189894
R24730 commonsourceibias.n652 commonsourceibias.n651 0.189894
R24731 commonsourceibias.n652 commonsourceibias.n638 0.189894
R24732 commonsourceibias.n658 commonsourceibias.n638 0.189894
R24733 commonsourceibias.n659 commonsourceibias.n658 0.189894
R24734 commonsourceibias.n660 commonsourceibias.n659 0.189894
R24735 commonsourceibias.n660 commonsourceibias.n636 0.189894
R24736 commonsourceibias.n665 commonsourceibias.n636 0.189894
R24737 commonsourceibias.n666 commonsourceibias.n665 0.189894
R24738 commonsourceibias.n667 commonsourceibias.n666 0.189894
R24739 commonsourceibias.n667 commonsourceibias.n634 0.189894
R24740 commonsourceibias.n673 commonsourceibias.n634 0.189894
R24741 commonsourceibias.n674 commonsourceibias.n673 0.189894
R24742 commonsourceibias.n675 commonsourceibias.n674 0.189894
R24743 commonsourceibias.n675 commonsourceibias.n632 0.189894
R24744 commonsourceibias.n680 commonsourceibias.n632 0.189894
R24745 commonsourceibias.n681 commonsourceibias.n680 0.189894
R24746 commonsourceibias.n682 commonsourceibias.n681 0.189894
R24747 commonsourceibias.n682 commonsourceibias.n630 0.189894
R24748 commonsourceibias.n688 commonsourceibias.n630 0.189894
R24749 commonsourceibias.n689 commonsourceibias.n688 0.189894
R24750 commonsourceibias.n690 commonsourceibias.n689 0.189894
R24751 commonsourceibias.n690 commonsourceibias.n628 0.189894
R24752 commonsourceibias.n695 commonsourceibias.n628 0.189894
R24753 commonsourceibias.n696 commonsourceibias.n695 0.189894
R24754 commonsourceibias.n697 commonsourceibias.n696 0.189894
R24755 commonsourceibias.n697 commonsourceibias.n626 0.189894
R24756 commonsourceibias.n703 commonsourceibias.n626 0.189894
R24757 commonsourceibias.n704 commonsourceibias.n703 0.189894
R24758 commonsourceibias.n705 commonsourceibias.n704 0.189894
R24759 commonsourceibias.n705 commonsourceibias.n624 0.189894
R24760 commonsourceibias.n710 commonsourceibias.n624 0.189894
R24761 commonsourceibias.n711 commonsourceibias.n710 0.189894
R24762 commonsourceibias.n712 commonsourceibias.n711 0.189894
R24763 commonsourceibias.n712 commonsourceibias.n622 0.189894
R24764 commonsourceibias.n718 commonsourceibias.n622 0.189894
R24765 commonsourceibias.n719 commonsourceibias.n718 0.189894
R24766 commonsourceibias.n720 commonsourceibias.n719 0.189894
R24767 commonsourceibias.n720 commonsourceibias.n620 0.189894
R24768 commonsourceibias.n725 commonsourceibias.n620 0.189894
R24769 commonsourceibias.n726 commonsourceibias.n725 0.189894
R24770 commonsourceibias.n727 commonsourceibias.n726 0.189894
R24771 commonsourceibias.n727 commonsourceibias.n618 0.189894
R24772 commonsourceibias.n415 commonsourceibias.n414 0.189894
R24773 commonsourceibias.n415 commonsourceibias.n410 0.189894
R24774 commonsourceibias.n420 commonsourceibias.n410 0.189894
R24775 commonsourceibias.n421 commonsourceibias.n420 0.189894
R24776 commonsourceibias.n422 commonsourceibias.n421 0.189894
R24777 commonsourceibias.n422 commonsourceibias.n408 0.189894
R24778 commonsourceibias.n428 commonsourceibias.n408 0.189894
R24779 commonsourceibias.n429 commonsourceibias.n428 0.189894
R24780 commonsourceibias.n430 commonsourceibias.n429 0.189894
R24781 commonsourceibias.n430 commonsourceibias.n406 0.189894
R24782 commonsourceibias.n435 commonsourceibias.n406 0.189894
R24783 commonsourceibias.n436 commonsourceibias.n435 0.189894
R24784 commonsourceibias.n437 commonsourceibias.n436 0.189894
R24785 commonsourceibias.n437 commonsourceibias.n404 0.189894
R24786 commonsourceibias.n443 commonsourceibias.n404 0.189894
R24787 commonsourceibias.n444 commonsourceibias.n443 0.189894
R24788 commonsourceibias.n445 commonsourceibias.n444 0.189894
R24789 commonsourceibias.n445 commonsourceibias.n402 0.189894
R24790 commonsourceibias.n450 commonsourceibias.n402 0.189894
R24791 commonsourceibias.n451 commonsourceibias.n450 0.189894
R24792 commonsourceibias.n452 commonsourceibias.n451 0.189894
R24793 commonsourceibias.n452 commonsourceibias.n400 0.189894
R24794 commonsourceibias.n458 commonsourceibias.n400 0.189894
R24795 commonsourceibias.n459 commonsourceibias.n458 0.189894
R24796 commonsourceibias.n460 commonsourceibias.n459 0.189894
R24797 commonsourceibias.n460 commonsourceibias.n398 0.189894
R24798 commonsourceibias.n465 commonsourceibias.n398 0.189894
R24799 commonsourceibias.n466 commonsourceibias.n465 0.189894
R24800 commonsourceibias.n467 commonsourceibias.n466 0.189894
R24801 commonsourceibias.n467 commonsourceibias.n396 0.189894
R24802 commonsourceibias.n473 commonsourceibias.n396 0.189894
R24803 commonsourceibias.n474 commonsourceibias.n473 0.189894
R24804 commonsourceibias.n475 commonsourceibias.n474 0.189894
R24805 commonsourceibias.n475 commonsourceibias.n394 0.189894
R24806 commonsourceibias.n480 commonsourceibias.n394 0.189894
R24807 commonsourceibias.n481 commonsourceibias.n480 0.189894
R24808 commonsourceibias.n482 commonsourceibias.n481 0.189894
R24809 commonsourceibias.n482 commonsourceibias.n392 0.189894
R24810 commonsourceibias.n488 commonsourceibias.n392 0.189894
R24811 commonsourceibias.n489 commonsourceibias.n488 0.189894
R24812 commonsourceibias.n490 commonsourceibias.n489 0.189894
R24813 commonsourceibias.n490 commonsourceibias.n390 0.189894
R24814 commonsourceibias.n495 commonsourceibias.n390 0.189894
R24815 commonsourceibias.n496 commonsourceibias.n495 0.189894
R24816 commonsourceibias.n497 commonsourceibias.n496 0.189894
R24817 commonsourceibias.n497 commonsourceibias.n388 0.189894
R24818 commonsourceibias.n531 commonsourceibias.n530 0.189894
R24819 commonsourceibias.n531 commonsourceibias.n526 0.189894
R24820 commonsourceibias.n536 commonsourceibias.n526 0.189894
R24821 commonsourceibias.n537 commonsourceibias.n536 0.189894
R24822 commonsourceibias.n538 commonsourceibias.n537 0.189894
R24823 commonsourceibias.n538 commonsourceibias.n524 0.189894
R24824 commonsourceibias.n544 commonsourceibias.n524 0.189894
R24825 commonsourceibias.n545 commonsourceibias.n544 0.189894
R24826 commonsourceibias.n546 commonsourceibias.n545 0.189894
R24827 commonsourceibias.n546 commonsourceibias.n522 0.189894
R24828 commonsourceibias.n551 commonsourceibias.n522 0.189894
R24829 commonsourceibias.n552 commonsourceibias.n551 0.189894
R24830 commonsourceibias.n553 commonsourceibias.n552 0.189894
R24831 commonsourceibias.n553 commonsourceibias.n520 0.189894
R24832 commonsourceibias.n558 commonsourceibias.n520 0.189894
R24833 commonsourceibias.n559 commonsourceibias.n558 0.189894
R24834 commonsourceibias.n559 commonsourceibias.n518 0.189894
R24835 commonsourceibias.n563 commonsourceibias.n518 0.189894
R24836 commonsourceibias.n564 commonsourceibias.n563 0.189894
R24837 commonsourceibias.n564 commonsourceibias.n516 0.189894
R24838 commonsourceibias.n568 commonsourceibias.n516 0.189894
R24839 commonsourceibias.n569 commonsourceibias.n568 0.189894
R24840 commonsourceibias.n574 commonsourceibias.n573 0.189894
R24841 commonsourceibias.n575 commonsourceibias.n574 0.189894
R24842 commonsourceibias.n575 commonsourceibias.n377 0.189894
R24843 commonsourceibias.n580 commonsourceibias.n377 0.189894
R24844 commonsourceibias.n581 commonsourceibias.n580 0.189894
R24845 commonsourceibias.n582 commonsourceibias.n581 0.189894
R24846 commonsourceibias.n582 commonsourceibias.n375 0.189894
R24847 commonsourceibias.n588 commonsourceibias.n375 0.189894
R24848 commonsourceibias.n589 commonsourceibias.n588 0.189894
R24849 commonsourceibias.n590 commonsourceibias.n589 0.189894
R24850 commonsourceibias.n590 commonsourceibias.n373 0.189894
R24851 commonsourceibias.n595 commonsourceibias.n373 0.189894
R24852 commonsourceibias.n596 commonsourceibias.n595 0.189894
R24853 commonsourceibias.n597 commonsourceibias.n596 0.189894
R24854 commonsourceibias.n597 commonsourceibias.n371 0.189894
R24855 commonsourceibias.n603 commonsourceibias.n371 0.189894
R24856 commonsourceibias.n604 commonsourceibias.n603 0.189894
R24857 commonsourceibias.n605 commonsourceibias.n604 0.189894
R24858 commonsourceibias.n605 commonsourceibias.n369 0.189894
R24859 commonsourceibias.n610 commonsourceibias.n369 0.189894
R24860 commonsourceibias.n611 commonsourceibias.n610 0.189894
R24861 commonsourceibias.n612 commonsourceibias.n611 0.189894
R24862 commonsourceibias.n612 commonsourceibias.n367 0.189894
R24863 commonsourceibias.n205 commonsourceibias.n149 0.0762576
R24864 commonsourceibias.n208 commonsourceibias.n149 0.0762576
R24865 commonsourceibias.n569 commonsourceibias.n514 0.0762576
R24866 commonsourceibias.n573 commonsourceibias.n514 0.0762576
R24867 a_n2982_8322.n28 a_n2982_8322.t20 74.6477
R24868 a_n2982_8322.n13 a_n2982_8322.t9 74.6477
R24869 a_n2982_8322.n1 a_n2982_8322.t35 74.6474
R24870 a_n2982_8322.n20 a_n2982_8322.t14 74.2899
R24871 a_n2982_8322.n10 a_n2982_8322.t15 74.2899
R24872 a_n2982_8322.n14 a_n2982_8322.t7 74.2899
R24873 a_n2982_8322.n15 a_n2982_8322.t10 74.2899
R24874 a_n2982_8322.n18 a_n2982_8322.t11 74.2899
R24875 a_n2982_8322.n28 a_n2982_8322.n27 70.6783
R24876 a_n2982_8322.n26 a_n2982_8322.n25 70.6783
R24877 a_n2982_8322.n24 a_n2982_8322.n23 70.6783
R24878 a_n2982_8322.n22 a_n2982_8322.n21 70.6783
R24879 a_n2982_8322.n1 a_n2982_8322.n0 70.6783
R24880 a_n2982_8322.n3 a_n2982_8322.n2 70.6783
R24881 a_n2982_8322.n5 a_n2982_8322.n4 70.6783
R24882 a_n2982_8322.n7 a_n2982_8322.n6 70.6783
R24883 a_n2982_8322.n9 a_n2982_8322.n8 70.6783
R24884 a_n2982_8322.n13 a_n2982_8322.n12 70.6783
R24885 a_n2982_8322.n17 a_n2982_8322.n16 70.6783
R24886 a_n2982_8322.n30 a_n2982_8322.n29 70.6782
R24887 a_n2982_8322.n20 a_n2982_8322.n19 24.9022
R24888 a_n2982_8322.n11 a_n2982_8322.t0 9.96358
R24889 a_n2982_8322.n19 a_n2982_8322.n18 8.38735
R24890 a_n2982_8322.n11 a_n2982_8322.n10 6.90998
R24891 a_n2982_8322.n19 a_n2982_8322.n11 5.3452
R24892 a_n2982_8322.n27 a_n2982_8322.t33 3.61217
R24893 a_n2982_8322.n27 a_n2982_8322.t29 3.61217
R24894 a_n2982_8322.n25 a_n2982_8322.t17 3.61217
R24895 a_n2982_8322.n25 a_n2982_8322.t16 3.61217
R24896 a_n2982_8322.n23 a_n2982_8322.t30 3.61217
R24897 a_n2982_8322.n23 a_n2982_8322.t23 3.61217
R24898 a_n2982_8322.n21 a_n2982_8322.t27 3.61217
R24899 a_n2982_8322.n21 a_n2982_8322.t25 3.61217
R24900 a_n2982_8322.n0 a_n2982_8322.t28 3.61217
R24901 a_n2982_8322.n0 a_n2982_8322.t24 3.61217
R24902 a_n2982_8322.n2 a_n2982_8322.t21 3.61217
R24903 a_n2982_8322.n2 a_n2982_8322.t37 3.61217
R24904 a_n2982_8322.n4 a_n2982_8322.t34 3.61217
R24905 a_n2982_8322.n4 a_n2982_8322.t22 3.61217
R24906 a_n2982_8322.n6 a_n2982_8322.t19 3.61217
R24907 a_n2982_8322.n6 a_n2982_8322.t18 3.61217
R24908 a_n2982_8322.n8 a_n2982_8322.t32 3.61217
R24909 a_n2982_8322.n8 a_n2982_8322.t31 3.61217
R24910 a_n2982_8322.n12 a_n2982_8322.t13 3.61217
R24911 a_n2982_8322.n12 a_n2982_8322.t12 3.61217
R24912 a_n2982_8322.n16 a_n2982_8322.t8 3.61217
R24913 a_n2982_8322.n16 a_n2982_8322.t6 3.61217
R24914 a_n2982_8322.t36 a_n2982_8322.n30 3.61217
R24915 a_n2982_8322.n30 a_n2982_8322.t26 3.61217
R24916 a_n2982_8322.n10 a_n2982_8322.n9 0.358259
R24917 a_n2982_8322.n9 a_n2982_8322.n7 0.358259
R24918 a_n2982_8322.n7 a_n2982_8322.n5 0.358259
R24919 a_n2982_8322.n5 a_n2982_8322.n3 0.358259
R24920 a_n2982_8322.n3 a_n2982_8322.n1 0.358259
R24921 a_n2982_8322.n18 a_n2982_8322.n17 0.358259
R24922 a_n2982_8322.n17 a_n2982_8322.n15 0.358259
R24923 a_n2982_8322.n14 a_n2982_8322.n13 0.358259
R24924 a_n2982_8322.n22 a_n2982_8322.n20 0.358259
R24925 a_n2982_8322.n24 a_n2982_8322.n22 0.358259
R24926 a_n2982_8322.n26 a_n2982_8322.n24 0.358259
R24927 a_n2982_8322.n29 a_n2982_8322.n26 0.358259
R24928 a_n2982_8322.n29 a_n2982_8322.n28 0.358259
R24929 a_n2982_8322.n15 a_n2982_8322.n14 0.101793
R24930 a_n2982_8322.t5 a_n2982_8322.t2 0.0788333
R24931 a_n2982_8322.t4 a_n2982_8322.t3 0.0788333
R24932 a_n2982_8322.t0 a_n2982_8322.t1 0.0788333
R24933 a_n2982_8322.t4 a_n2982_8322.t5 0.0318333
R24934 a_n2982_8322.t0 a_n2982_8322.t3 0.0318333
R24935 a_n2982_8322.t2 a_n2982_8322.t3 0.0318333
R24936 a_n2982_8322.t1 a_n2982_8322.t4 0.0318333
R24937 output.n41 output.n15 289.615
R24938 output.n72 output.n46 289.615
R24939 output.n104 output.n78 289.615
R24940 output.n136 output.n110 289.615
R24941 output.n77 output.n45 197.26
R24942 output.n77 output.n76 196.298
R24943 output.n109 output.n108 196.298
R24944 output.n141 output.n140 196.298
R24945 output.n42 output.n41 185
R24946 output.n40 output.n39 185
R24947 output.n19 output.n18 185
R24948 output.n34 output.n33 185
R24949 output.n32 output.n31 185
R24950 output.n23 output.n22 185
R24951 output.n26 output.n25 185
R24952 output.n73 output.n72 185
R24953 output.n71 output.n70 185
R24954 output.n50 output.n49 185
R24955 output.n65 output.n64 185
R24956 output.n63 output.n62 185
R24957 output.n54 output.n53 185
R24958 output.n57 output.n56 185
R24959 output.n105 output.n104 185
R24960 output.n103 output.n102 185
R24961 output.n82 output.n81 185
R24962 output.n97 output.n96 185
R24963 output.n95 output.n94 185
R24964 output.n86 output.n85 185
R24965 output.n89 output.n88 185
R24966 output.n137 output.n136 185
R24967 output.n135 output.n134 185
R24968 output.n114 output.n113 185
R24969 output.n129 output.n128 185
R24970 output.n127 output.n126 185
R24971 output.n118 output.n117 185
R24972 output.n121 output.n120 185
R24973 output.t3 output.n24 147.661
R24974 output.t1 output.n55 147.661
R24975 output.t2 output.n87 147.661
R24976 output.t0 output.n119 147.661
R24977 output.n41 output.n40 104.615
R24978 output.n40 output.n18 104.615
R24979 output.n33 output.n18 104.615
R24980 output.n33 output.n32 104.615
R24981 output.n32 output.n22 104.615
R24982 output.n25 output.n22 104.615
R24983 output.n72 output.n71 104.615
R24984 output.n71 output.n49 104.615
R24985 output.n64 output.n49 104.615
R24986 output.n64 output.n63 104.615
R24987 output.n63 output.n53 104.615
R24988 output.n56 output.n53 104.615
R24989 output.n104 output.n103 104.615
R24990 output.n103 output.n81 104.615
R24991 output.n96 output.n81 104.615
R24992 output.n96 output.n95 104.615
R24993 output.n95 output.n85 104.615
R24994 output.n88 output.n85 104.615
R24995 output.n136 output.n135 104.615
R24996 output.n135 output.n113 104.615
R24997 output.n128 output.n113 104.615
R24998 output.n128 output.n127 104.615
R24999 output.n127 output.n117 104.615
R25000 output.n120 output.n117 104.615
R25001 output.n1 output.t13 77.056
R25002 output.n14 output.t15 76.6694
R25003 output.n1 output.n0 72.7095
R25004 output.n3 output.n2 72.7095
R25005 output.n5 output.n4 72.7095
R25006 output.n7 output.n6 72.7095
R25007 output.n9 output.n8 72.7095
R25008 output.n11 output.n10 72.7095
R25009 output.n13 output.n12 72.7095
R25010 output.n25 output.t3 52.3082
R25011 output.n56 output.t1 52.3082
R25012 output.n88 output.t2 52.3082
R25013 output.n120 output.t0 52.3082
R25014 output.n26 output.n24 15.6674
R25015 output.n57 output.n55 15.6674
R25016 output.n89 output.n87 15.6674
R25017 output.n121 output.n119 15.6674
R25018 output.n27 output.n23 12.8005
R25019 output.n58 output.n54 12.8005
R25020 output.n90 output.n86 12.8005
R25021 output.n122 output.n118 12.8005
R25022 output.n31 output.n30 12.0247
R25023 output.n62 output.n61 12.0247
R25024 output.n94 output.n93 12.0247
R25025 output.n126 output.n125 12.0247
R25026 output.n34 output.n21 11.249
R25027 output.n65 output.n52 11.249
R25028 output.n97 output.n84 11.249
R25029 output.n129 output.n116 11.249
R25030 output.n35 output.n19 10.4732
R25031 output.n66 output.n50 10.4732
R25032 output.n98 output.n82 10.4732
R25033 output.n130 output.n114 10.4732
R25034 output.n39 output.n38 9.69747
R25035 output.n70 output.n69 9.69747
R25036 output.n102 output.n101 9.69747
R25037 output.n134 output.n133 9.69747
R25038 output.n45 output.n44 9.45567
R25039 output.n76 output.n75 9.45567
R25040 output.n108 output.n107 9.45567
R25041 output.n140 output.n139 9.45567
R25042 output.n44 output.n43 9.3005
R25043 output.n17 output.n16 9.3005
R25044 output.n38 output.n37 9.3005
R25045 output.n36 output.n35 9.3005
R25046 output.n21 output.n20 9.3005
R25047 output.n30 output.n29 9.3005
R25048 output.n28 output.n27 9.3005
R25049 output.n75 output.n74 9.3005
R25050 output.n48 output.n47 9.3005
R25051 output.n69 output.n68 9.3005
R25052 output.n67 output.n66 9.3005
R25053 output.n52 output.n51 9.3005
R25054 output.n61 output.n60 9.3005
R25055 output.n59 output.n58 9.3005
R25056 output.n107 output.n106 9.3005
R25057 output.n80 output.n79 9.3005
R25058 output.n101 output.n100 9.3005
R25059 output.n99 output.n98 9.3005
R25060 output.n84 output.n83 9.3005
R25061 output.n93 output.n92 9.3005
R25062 output.n91 output.n90 9.3005
R25063 output.n139 output.n138 9.3005
R25064 output.n112 output.n111 9.3005
R25065 output.n133 output.n132 9.3005
R25066 output.n131 output.n130 9.3005
R25067 output.n116 output.n115 9.3005
R25068 output.n125 output.n124 9.3005
R25069 output.n123 output.n122 9.3005
R25070 output.n42 output.n17 8.92171
R25071 output.n73 output.n48 8.92171
R25072 output.n105 output.n80 8.92171
R25073 output.n137 output.n112 8.92171
R25074 output output.n141 8.15037
R25075 output.n43 output.n15 8.14595
R25076 output.n74 output.n46 8.14595
R25077 output.n106 output.n78 8.14595
R25078 output.n138 output.n110 8.14595
R25079 output.n45 output.n15 5.81868
R25080 output.n76 output.n46 5.81868
R25081 output.n108 output.n78 5.81868
R25082 output.n140 output.n110 5.81868
R25083 output.n43 output.n42 5.04292
R25084 output.n74 output.n73 5.04292
R25085 output.n106 output.n105 5.04292
R25086 output.n138 output.n137 5.04292
R25087 output.n28 output.n24 4.38594
R25088 output.n59 output.n55 4.38594
R25089 output.n91 output.n87 4.38594
R25090 output.n123 output.n119 4.38594
R25091 output.n39 output.n17 4.26717
R25092 output.n70 output.n48 4.26717
R25093 output.n102 output.n80 4.26717
R25094 output.n134 output.n112 4.26717
R25095 output.n0 output.t19 3.9605
R25096 output.n0 output.t8 3.9605
R25097 output.n2 output.t12 3.9605
R25098 output.n2 output.t4 3.9605
R25099 output.n4 output.t6 3.9605
R25100 output.n4 output.t5 3.9605
R25101 output.n6 output.t11 3.9605
R25102 output.n6 output.t14 3.9605
R25103 output.n8 output.t16 3.9605
R25104 output.n8 output.t9 3.9605
R25105 output.n10 output.t10 3.9605
R25106 output.n10 output.t17 3.9605
R25107 output.n12 output.t18 3.9605
R25108 output.n12 output.t7 3.9605
R25109 output.n38 output.n19 3.49141
R25110 output.n69 output.n50 3.49141
R25111 output.n101 output.n82 3.49141
R25112 output.n133 output.n114 3.49141
R25113 output.n35 output.n34 2.71565
R25114 output.n66 output.n65 2.71565
R25115 output.n98 output.n97 2.71565
R25116 output.n130 output.n129 2.71565
R25117 output.n31 output.n21 1.93989
R25118 output.n62 output.n52 1.93989
R25119 output.n94 output.n84 1.93989
R25120 output.n126 output.n116 1.93989
R25121 output.n30 output.n23 1.16414
R25122 output.n61 output.n54 1.16414
R25123 output.n93 output.n86 1.16414
R25124 output.n125 output.n118 1.16414
R25125 output.n141 output.n109 0.962709
R25126 output.n109 output.n77 0.962709
R25127 output.n27 output.n26 0.388379
R25128 output.n58 output.n57 0.388379
R25129 output.n90 output.n89 0.388379
R25130 output.n122 output.n121 0.388379
R25131 output.n14 output.n13 0.387128
R25132 output.n13 output.n11 0.387128
R25133 output.n11 output.n9 0.387128
R25134 output.n9 output.n7 0.387128
R25135 output.n7 output.n5 0.387128
R25136 output.n5 output.n3 0.387128
R25137 output.n3 output.n1 0.387128
R25138 output.n44 output.n16 0.155672
R25139 output.n37 output.n16 0.155672
R25140 output.n37 output.n36 0.155672
R25141 output.n36 output.n20 0.155672
R25142 output.n29 output.n20 0.155672
R25143 output.n29 output.n28 0.155672
R25144 output.n75 output.n47 0.155672
R25145 output.n68 output.n47 0.155672
R25146 output.n68 output.n67 0.155672
R25147 output.n67 output.n51 0.155672
R25148 output.n60 output.n51 0.155672
R25149 output.n60 output.n59 0.155672
R25150 output.n107 output.n79 0.155672
R25151 output.n100 output.n79 0.155672
R25152 output.n100 output.n99 0.155672
R25153 output.n99 output.n83 0.155672
R25154 output.n92 output.n83 0.155672
R25155 output.n92 output.n91 0.155672
R25156 output.n139 output.n111 0.155672
R25157 output.n132 output.n111 0.155672
R25158 output.n132 output.n131 0.155672
R25159 output.n131 output.n115 0.155672
R25160 output.n124 output.n115 0.155672
R25161 output.n124 output.n123 0.155672
R25162 output output.n14 0.126227
R25163 minus.n33 minus.t20 321.495
R25164 minus.n7 minus.t6 321.495
R25165 minus.n50 minus.t18 297.12
R25166 minus.n48 minus.t15 297.12
R25167 minus.n28 minus.t16 297.12
R25168 minus.n42 minus.t11 297.12
R25169 minus.n30 minus.t12 297.12
R25170 minus.n36 minus.t7 297.12
R25171 minus.n32 minus.t19 297.12
R25172 minus.n6 minus.t5 297.12
R25173 minus.n10 minus.t9 297.12
R25174 minus.n12 minus.t8 297.12
R25175 minus.n16 minus.t10 297.12
R25176 minus.n18 minus.t14 297.12
R25177 minus.n22 minus.t13 297.12
R25178 minus.n24 minus.t17 297.12
R25179 minus.n56 minus.t4 243.255
R25180 minus.n55 minus.n53 224.169
R25181 minus.n55 minus.n54 223.454
R25182 minus.n35 minus.n34 161.3
R25183 minus.n36 minus.n31 161.3
R25184 minus.n38 minus.n37 161.3
R25185 minus.n39 minus.n30 161.3
R25186 minus.n41 minus.n40 161.3
R25187 minus.n42 minus.n29 161.3
R25188 minus.n44 minus.n43 161.3
R25189 minus.n45 minus.n28 161.3
R25190 minus.n47 minus.n46 161.3
R25191 minus.n48 minus.n27 161.3
R25192 minus.n49 minus.n26 161.3
R25193 minus.n51 minus.n50 161.3
R25194 minus.n25 minus.n24 161.3
R25195 minus.n23 minus.n0 161.3
R25196 minus.n22 minus.n21 161.3
R25197 minus.n20 minus.n1 161.3
R25198 minus.n19 minus.n18 161.3
R25199 minus.n17 minus.n2 161.3
R25200 minus.n16 minus.n15 161.3
R25201 minus.n14 minus.n3 161.3
R25202 minus.n13 minus.n12 161.3
R25203 minus.n11 minus.n4 161.3
R25204 minus.n10 minus.n9 161.3
R25205 minus.n8 minus.n5 161.3
R25206 minus.n8 minus.n7 44.9377
R25207 minus.n34 minus.n33 44.9377
R25208 minus.n50 minus.n49 37.246
R25209 minus.n24 minus.n23 37.246
R25210 minus.n48 minus.n47 32.8641
R25211 minus.n35 minus.n32 32.8641
R25212 minus.n6 minus.n5 32.8641
R25213 minus.n22 minus.n1 32.8641
R25214 minus.n52 minus.n51 30.2486
R25215 minus.n43 minus.n28 28.4823
R25216 minus.n37 minus.n36 28.4823
R25217 minus.n11 minus.n10 28.4823
R25218 minus.n18 minus.n17 28.4823
R25219 minus.n42 minus.n41 24.1005
R25220 minus.n41 minus.n30 24.1005
R25221 minus.n12 minus.n3 24.1005
R25222 minus.n16 minus.n3 24.1005
R25223 minus.n54 minus.t3 19.8005
R25224 minus.n54 minus.t2 19.8005
R25225 minus.n53 minus.t1 19.8005
R25226 minus.n53 minus.t0 19.8005
R25227 minus.n43 minus.n42 19.7187
R25228 minus.n37 minus.n30 19.7187
R25229 minus.n12 minus.n11 19.7187
R25230 minus.n17 minus.n16 19.7187
R25231 minus.n33 minus.n32 17.0522
R25232 minus.n7 minus.n6 17.0522
R25233 minus.n47 minus.n28 15.3369
R25234 minus.n36 minus.n35 15.3369
R25235 minus.n10 minus.n5 15.3369
R25236 minus.n18 minus.n1 15.3369
R25237 minus minus.n57 12.2906
R25238 minus.n52 minus.n25 12.0706
R25239 minus.n49 minus.n48 10.955
R25240 minus.n23 minus.n22 10.955
R25241 minus.n57 minus.n56 4.80222
R25242 minus.n57 minus.n52 0.972091
R25243 minus.n56 minus.n55 0.716017
R25244 minus.n51 minus.n26 0.189894
R25245 minus.n27 minus.n26 0.189894
R25246 minus.n46 minus.n27 0.189894
R25247 minus.n46 minus.n45 0.189894
R25248 minus.n45 minus.n44 0.189894
R25249 minus.n44 minus.n29 0.189894
R25250 minus.n40 minus.n29 0.189894
R25251 minus.n40 minus.n39 0.189894
R25252 minus.n39 minus.n38 0.189894
R25253 minus.n38 minus.n31 0.189894
R25254 minus.n34 minus.n31 0.189894
R25255 minus.n9 minus.n8 0.189894
R25256 minus.n9 minus.n4 0.189894
R25257 minus.n13 minus.n4 0.189894
R25258 minus.n14 minus.n13 0.189894
R25259 minus.n15 minus.n14 0.189894
R25260 minus.n15 minus.n2 0.189894
R25261 minus.n19 minus.n2 0.189894
R25262 minus.n20 minus.n19 0.189894
R25263 minus.n21 minus.n20 0.189894
R25264 minus.n21 minus.n0 0.189894
R25265 minus.n25 minus.n0 0.189894
C0 output outputibias 2.34152f
C1 vdd output 7.23429f
C2 CSoutput output 6.13571f
C3 CSoutput outputibias 0.032386f
C4 vdd CSoutput 0.14152p
C5 minus diffpairibias 3.1e-19
C6 commonsourceibias output 0.006808f
C7 CSoutput minus 3.37765f
C8 vdd plus 0.098689f
C9 commonsourceibias outputibias 0.003832f
C10 plus diffpairibias 3.12e-19
C11 vdd commonsourceibias 0.004218f
C12 CSoutput plus 0.880209f
C13 commonsourceibias diffpairibias 0.052527f
C14 CSoutput commonsourceibias 45.462303f
C15 minus plus 9.56783f
C16 minus commonsourceibias 0.327654f
C17 plus commonsourceibias 0.273048f
C18 diffpairibias gnd 59.991035f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.182015p
C22 plus gnd 32.471f
C23 minus gnd 28.40805f
C24 CSoutput gnd 0.115023p
C25 vdd gnd 0.543576p
C26 minus.n0 gnd 0.029692f
C27 minus.n1 gnd 0.006738f
C28 minus.n2 gnd 0.029692f
C29 minus.n3 gnd 0.006738f
C30 minus.n4 gnd 0.029692f
C31 minus.n5 gnd 0.006738f
C32 minus.t6 gnd 0.434123f
C33 minus.t5 gnd 0.419969f
C34 minus.n6 gnd 0.190631f
C35 minus.n7 gnd 0.174881f
C36 minus.n8 gnd 0.12565f
C37 minus.n9 gnd 0.029692f
C38 minus.t9 gnd 0.419969f
C39 minus.n10 gnd 0.186564f
C40 minus.n11 gnd 0.006738f
C41 minus.t8 gnd 0.419969f
C42 minus.n12 gnd 0.186564f
C43 minus.n13 gnd 0.029692f
C44 minus.n14 gnd 0.029692f
C45 minus.n15 gnd 0.029692f
C46 minus.t10 gnd 0.419969f
C47 minus.n16 gnd 0.186564f
C48 minus.n17 gnd 0.006738f
C49 minus.t14 gnd 0.419969f
C50 minus.n18 gnd 0.186564f
C51 minus.n19 gnd 0.029692f
C52 minus.n20 gnd 0.029692f
C53 minus.n21 gnd 0.029692f
C54 minus.t13 gnd 0.419969f
C55 minus.n22 gnd 0.186564f
C56 minus.n23 gnd 0.006738f
C57 minus.t17 gnd 0.419969f
C58 minus.n24 gnd 0.18574f
C59 minus.n25 gnd 0.342275f
C60 minus.n26 gnd 0.029692f
C61 minus.t18 gnd 0.419969f
C62 minus.t15 gnd 0.419969f
C63 minus.n27 gnd 0.029692f
C64 minus.t16 gnd 0.419969f
C65 minus.n28 gnd 0.186564f
C66 minus.n29 gnd 0.029692f
C67 minus.t11 gnd 0.419969f
C68 minus.t12 gnd 0.419969f
C69 minus.n30 gnd 0.186564f
C70 minus.n31 gnd 0.029692f
C71 minus.t7 gnd 0.419969f
C72 minus.t19 gnd 0.419969f
C73 minus.n32 gnd 0.190631f
C74 minus.t20 gnd 0.434123f
C75 minus.n33 gnd 0.174881f
C76 minus.n34 gnd 0.12565f
C77 minus.n35 gnd 0.006738f
C78 minus.n36 gnd 0.186564f
C79 minus.n37 gnd 0.006738f
C80 minus.n38 gnd 0.029692f
C81 minus.n39 gnd 0.029692f
C82 minus.n40 gnd 0.029692f
C83 minus.n41 gnd 0.006738f
C84 minus.n42 gnd 0.186564f
C85 minus.n43 gnd 0.006738f
C86 minus.n44 gnd 0.029692f
C87 minus.n45 gnd 0.029692f
C88 minus.n46 gnd 0.029692f
C89 minus.n47 gnd 0.006738f
C90 minus.n48 gnd 0.186564f
C91 minus.n49 gnd 0.006738f
C92 minus.n50 gnd 0.18574f
C93 minus.n51 gnd 0.86182f
C94 minus.n52 gnd 1.31052f
C95 minus.t1 gnd 0.009153f
C96 minus.t0 gnd 0.009153f
C97 minus.n53 gnd 0.030098f
C98 minus.t3 gnd 0.009153f
C99 minus.t2 gnd 0.009153f
C100 minus.n54 gnd 0.029686f
C101 minus.n55 gnd 0.253353f
C102 minus.t4 gnd 0.050946f
C103 minus.n56 gnd 0.138252f
C104 minus.n57 gnd 2.39424f
C105 output.t13 gnd 0.464308f
C106 output.t19 gnd 0.044422f
C107 output.t8 gnd 0.044422f
C108 output.n0 gnd 0.364624f
C109 output.n1 gnd 0.614102f
C110 output.t12 gnd 0.044422f
C111 output.t4 gnd 0.044422f
C112 output.n2 gnd 0.364624f
C113 output.n3 gnd 0.350265f
C114 output.t6 gnd 0.044422f
C115 output.t5 gnd 0.044422f
C116 output.n4 gnd 0.364624f
C117 output.n5 gnd 0.350265f
C118 output.t11 gnd 0.044422f
C119 output.t14 gnd 0.044422f
C120 output.n6 gnd 0.364624f
C121 output.n7 gnd 0.350265f
C122 output.t16 gnd 0.044422f
C123 output.t9 gnd 0.044422f
C124 output.n8 gnd 0.364624f
C125 output.n9 gnd 0.350265f
C126 output.t10 gnd 0.044422f
C127 output.t17 gnd 0.044422f
C128 output.n10 gnd 0.364624f
C129 output.n11 gnd 0.350265f
C130 output.t18 gnd 0.044422f
C131 output.t7 gnd 0.044422f
C132 output.n12 gnd 0.364624f
C133 output.n13 gnd 0.350265f
C134 output.t15 gnd 0.462979f
C135 output.n14 gnd 0.28994f
C136 output.n15 gnd 0.015803f
C137 output.n16 gnd 0.011243f
C138 output.n17 gnd 0.006041f
C139 output.n18 gnd 0.01428f
C140 output.n19 gnd 0.006397f
C141 output.n20 gnd 0.011243f
C142 output.n21 gnd 0.006041f
C143 output.n22 gnd 0.01428f
C144 output.n23 gnd 0.006397f
C145 output.n24 gnd 0.048111f
C146 output.t3 gnd 0.023274f
C147 output.n25 gnd 0.01071f
C148 output.n26 gnd 0.008435f
C149 output.n27 gnd 0.006041f
C150 output.n28 gnd 0.267512f
C151 output.n29 gnd 0.011243f
C152 output.n30 gnd 0.006041f
C153 output.n31 gnd 0.006397f
C154 output.n32 gnd 0.01428f
C155 output.n33 gnd 0.01428f
C156 output.n34 gnd 0.006397f
C157 output.n35 gnd 0.006041f
C158 output.n36 gnd 0.011243f
C159 output.n37 gnd 0.011243f
C160 output.n38 gnd 0.006041f
C161 output.n39 gnd 0.006397f
C162 output.n40 gnd 0.01428f
C163 output.n41 gnd 0.030913f
C164 output.n42 gnd 0.006397f
C165 output.n43 gnd 0.006041f
C166 output.n44 gnd 0.025987f
C167 output.n45 gnd 0.097665f
C168 output.n46 gnd 0.015803f
C169 output.n47 gnd 0.011243f
C170 output.n48 gnd 0.006041f
C171 output.n49 gnd 0.01428f
C172 output.n50 gnd 0.006397f
C173 output.n51 gnd 0.011243f
C174 output.n52 gnd 0.006041f
C175 output.n53 gnd 0.01428f
C176 output.n54 gnd 0.006397f
C177 output.n55 gnd 0.048111f
C178 output.t1 gnd 0.023274f
C179 output.n56 gnd 0.01071f
C180 output.n57 gnd 0.008435f
C181 output.n58 gnd 0.006041f
C182 output.n59 gnd 0.267512f
C183 output.n60 gnd 0.011243f
C184 output.n61 gnd 0.006041f
C185 output.n62 gnd 0.006397f
C186 output.n63 gnd 0.01428f
C187 output.n64 gnd 0.01428f
C188 output.n65 gnd 0.006397f
C189 output.n66 gnd 0.006041f
C190 output.n67 gnd 0.011243f
C191 output.n68 gnd 0.011243f
C192 output.n69 gnd 0.006041f
C193 output.n70 gnd 0.006397f
C194 output.n71 gnd 0.01428f
C195 output.n72 gnd 0.030913f
C196 output.n73 gnd 0.006397f
C197 output.n74 gnd 0.006041f
C198 output.n75 gnd 0.025987f
C199 output.n76 gnd 0.09306f
C200 output.n77 gnd 1.65264f
C201 output.n78 gnd 0.015803f
C202 output.n79 gnd 0.011243f
C203 output.n80 gnd 0.006041f
C204 output.n81 gnd 0.01428f
C205 output.n82 gnd 0.006397f
C206 output.n83 gnd 0.011243f
C207 output.n84 gnd 0.006041f
C208 output.n85 gnd 0.01428f
C209 output.n86 gnd 0.006397f
C210 output.n87 gnd 0.048111f
C211 output.t2 gnd 0.023274f
C212 output.n88 gnd 0.01071f
C213 output.n89 gnd 0.008435f
C214 output.n90 gnd 0.006041f
C215 output.n91 gnd 0.267512f
C216 output.n92 gnd 0.011243f
C217 output.n93 gnd 0.006041f
C218 output.n94 gnd 0.006397f
C219 output.n95 gnd 0.01428f
C220 output.n96 gnd 0.01428f
C221 output.n97 gnd 0.006397f
C222 output.n98 gnd 0.006041f
C223 output.n99 gnd 0.011243f
C224 output.n100 gnd 0.011243f
C225 output.n101 gnd 0.006041f
C226 output.n102 gnd 0.006397f
C227 output.n103 gnd 0.01428f
C228 output.n104 gnd 0.030913f
C229 output.n105 gnd 0.006397f
C230 output.n106 gnd 0.006041f
C231 output.n107 gnd 0.025987f
C232 output.n108 gnd 0.09306f
C233 output.n109 gnd 0.713089f
C234 output.n110 gnd 0.015803f
C235 output.n111 gnd 0.011243f
C236 output.n112 gnd 0.006041f
C237 output.n113 gnd 0.01428f
C238 output.n114 gnd 0.006397f
C239 output.n115 gnd 0.011243f
C240 output.n116 gnd 0.006041f
C241 output.n117 gnd 0.01428f
C242 output.n118 gnd 0.006397f
C243 output.n119 gnd 0.048111f
C244 output.t0 gnd 0.023274f
C245 output.n120 gnd 0.01071f
C246 output.n121 gnd 0.008435f
C247 output.n122 gnd 0.006041f
C248 output.n123 gnd 0.267512f
C249 output.n124 gnd 0.011243f
C250 output.n125 gnd 0.006041f
C251 output.n126 gnd 0.006397f
C252 output.n127 gnd 0.01428f
C253 output.n128 gnd 0.01428f
C254 output.n129 gnd 0.006397f
C255 output.n130 gnd 0.006041f
C256 output.n131 gnd 0.011243f
C257 output.n132 gnd 0.011243f
C258 output.n133 gnd 0.006041f
C259 output.n134 gnd 0.006397f
C260 output.n135 gnd 0.01428f
C261 output.n136 gnd 0.030913f
C262 output.n137 gnd 0.006397f
C263 output.n138 gnd 0.006041f
C264 output.n139 gnd 0.025987f
C265 output.n140 gnd 0.09306f
C266 output.n141 gnd 1.67353f
C267 a_n2982_8322.t26 gnd 0.100069f
C268 a_n2982_8322.t3 gnd 20.7601f
C269 a_n2982_8322.t2 gnd 20.6146f
C270 a_n2982_8322.t5 gnd 20.6146f
C271 a_n2982_8322.t4 gnd 20.7601f
C272 a_n2982_8322.t1 gnd 20.6146f
C273 a_n2982_8322.t0 gnd 30.2036f
C274 a_n2982_8322.t35 gnd 0.936988f
C275 a_n2982_8322.t28 gnd 0.100069f
C276 a_n2982_8322.t24 gnd 0.100069f
C277 a_n2982_8322.n0 gnd 0.704883f
C278 a_n2982_8322.n1 gnd 0.787605f
C279 a_n2982_8322.t21 gnd 0.100069f
C280 a_n2982_8322.t37 gnd 0.100069f
C281 a_n2982_8322.n2 gnd 0.704883f
C282 a_n2982_8322.n3 gnd 0.400171f
C283 a_n2982_8322.t34 gnd 0.100069f
C284 a_n2982_8322.t22 gnd 0.100069f
C285 a_n2982_8322.n4 gnd 0.704883f
C286 a_n2982_8322.n5 gnd 0.400171f
C287 a_n2982_8322.t19 gnd 0.100069f
C288 a_n2982_8322.t18 gnd 0.100069f
C289 a_n2982_8322.n6 gnd 0.704883f
C290 a_n2982_8322.n7 gnd 0.400171f
C291 a_n2982_8322.t32 gnd 0.100069f
C292 a_n2982_8322.t31 gnd 0.100069f
C293 a_n2982_8322.n8 gnd 0.704883f
C294 a_n2982_8322.n9 gnd 0.400171f
C295 a_n2982_8322.t15 gnd 0.935125f
C296 a_n2982_8322.n10 gnd 1.11045f
C297 a_n2982_8322.n11 gnd 3.82915f
C298 a_n2982_8322.t9 gnd 0.936991f
C299 a_n2982_8322.t13 gnd 0.100069f
C300 a_n2982_8322.t12 gnd 0.100069f
C301 a_n2982_8322.n12 gnd 0.704883f
C302 a_n2982_8322.n13 gnd 0.787602f
C303 a_n2982_8322.t7 gnd 0.935125f
C304 a_n2982_8322.n14 gnd 0.396333f
C305 a_n2982_8322.t10 gnd 0.935125f
C306 a_n2982_8322.n15 gnd 0.396333f
C307 a_n2982_8322.t8 gnd 0.100069f
C308 a_n2982_8322.t6 gnd 0.100069f
C309 a_n2982_8322.n16 gnd 0.704883f
C310 a_n2982_8322.n17 gnd 0.400171f
C311 a_n2982_8322.t11 gnd 0.935125f
C312 a_n2982_8322.n18 gnd 1.47007f
C313 a_n2982_8322.n19 gnd 2.34921f
C314 a_n2982_8322.t14 gnd 0.935125f
C315 a_n2982_8322.n20 gnd 1.86969f
C316 a_n2982_8322.t27 gnd 0.100069f
C317 a_n2982_8322.t25 gnd 0.100069f
C318 a_n2982_8322.n21 gnd 0.704883f
C319 a_n2982_8322.n22 gnd 0.400171f
C320 a_n2982_8322.t30 gnd 0.100069f
C321 a_n2982_8322.t23 gnd 0.100069f
C322 a_n2982_8322.n23 gnd 0.704883f
C323 a_n2982_8322.n24 gnd 0.400171f
C324 a_n2982_8322.t17 gnd 0.100069f
C325 a_n2982_8322.t16 gnd 0.100069f
C326 a_n2982_8322.n25 gnd 0.704883f
C327 a_n2982_8322.n26 gnd 0.400171f
C328 a_n2982_8322.t20 gnd 0.936991f
C329 a_n2982_8322.t33 gnd 0.100069f
C330 a_n2982_8322.t29 gnd 0.100069f
C331 a_n2982_8322.n27 gnd 0.704883f
C332 a_n2982_8322.n28 gnd 0.787602f
C333 a_n2982_8322.n29 gnd 0.400169f
C334 a_n2982_8322.n30 gnd 0.704885f
C335 a_n2982_8322.t36 gnd 0.100069f
C336 commonsourceibias.n0 gnd 0.010724f
C337 commonsourceibias.t115 gnd 0.162395f
C338 commonsourceibias.t136 gnd 0.150157f
C339 commonsourceibias.n1 gnd 0.007823f
C340 commonsourceibias.n2 gnd 0.008037f
C341 commonsourceibias.t151 gnd 0.150157f
C342 commonsourceibias.n3 gnd 0.01034f
C343 commonsourceibias.n4 gnd 0.008037f
C344 commonsourceibias.t105 gnd 0.150157f
C345 commonsourceibias.n5 gnd 0.059912f
C346 commonsourceibias.t126 gnd 0.150157f
C347 commonsourceibias.n6 gnd 0.007578f
C348 commonsourceibias.n7 gnd 0.008037f
C349 commonsourceibias.t144 gnd 0.150157f
C350 commonsourceibias.n8 gnd 0.010186f
C351 commonsourceibias.n9 gnd 0.008037f
C352 commonsourceibias.t98 gnd 0.150157f
C353 commonsourceibias.n10 gnd 0.059912f
C354 commonsourceibias.t94 gnd 0.150157f
C355 commonsourceibias.n11 gnd 0.007361f
C356 commonsourceibias.n12 gnd 0.008037f
C357 commonsourceibias.t135 gnd 0.150157f
C358 commonsourceibias.n13 gnd 0.010015f
C359 commonsourceibias.n14 gnd 0.010724f
C360 commonsourceibias.t74 gnd 0.162395f
C361 commonsourceibias.t20 gnd 0.150157f
C362 commonsourceibias.n15 gnd 0.007823f
C363 commonsourceibias.n16 gnd 0.008037f
C364 commonsourceibias.t50 gnd 0.150157f
C365 commonsourceibias.n17 gnd 0.01034f
C366 commonsourceibias.n18 gnd 0.008037f
C367 commonsourceibias.t8 gnd 0.150157f
C368 commonsourceibias.n19 gnd 0.059912f
C369 commonsourceibias.t36 gnd 0.150157f
C370 commonsourceibias.n20 gnd 0.007578f
C371 commonsourceibias.n21 gnd 0.008037f
C372 commonsourceibias.t76 gnd 0.150157f
C373 commonsourceibias.n22 gnd 0.010186f
C374 commonsourceibias.n23 gnd 0.008037f
C375 commonsourceibias.t24 gnd 0.150157f
C376 commonsourceibias.n24 gnd 0.059912f
C377 commonsourceibias.t34 gnd 0.150157f
C378 commonsourceibias.n25 gnd 0.007361f
C379 commonsourceibias.n26 gnd 0.008037f
C380 commonsourceibias.t10 gnd 0.150157f
C381 commonsourceibias.n27 gnd 0.010015f
C382 commonsourceibias.n28 gnd 0.008037f
C383 commonsourceibias.t40 gnd 0.150157f
C384 commonsourceibias.n29 gnd 0.059912f
C385 commonsourceibias.t56 gnd 0.150157f
C386 commonsourceibias.n30 gnd 0.007172f
C387 commonsourceibias.n31 gnd 0.008037f
C388 commonsourceibias.t26 gnd 0.150157f
C389 commonsourceibias.n32 gnd 0.009825f
C390 commonsourceibias.n33 gnd 0.008037f
C391 commonsourceibias.t38 gnd 0.150157f
C392 commonsourceibias.n34 gnd 0.059912f
C393 commonsourceibias.t70 gnd 0.150157f
C394 commonsourceibias.n35 gnd 0.007008f
C395 commonsourceibias.n36 gnd 0.008037f
C396 commonsourceibias.t18 gnd 0.150157f
C397 commonsourceibias.n37 gnd 0.009613f
C398 commonsourceibias.n38 gnd 0.008037f
C399 commonsourceibias.t22 gnd 0.150157f
C400 commonsourceibias.n39 gnd 0.059912f
C401 commonsourceibias.t54 gnd 0.150157f
C402 commonsourceibias.n40 gnd 0.006868f
C403 commonsourceibias.n41 gnd 0.008037f
C404 commonsourceibias.t4 gnd 0.150157f
C405 commonsourceibias.n42 gnd 0.009378f
C406 commonsourceibias.t78 gnd 0.166947f
C407 commonsourceibias.t46 gnd 0.150157f
C408 commonsourceibias.n43 gnd 0.065449f
C409 commonsourceibias.n44 gnd 0.071822f
C410 commonsourceibias.n45 gnd 0.033327f
C411 commonsourceibias.n46 gnd 0.008037f
C412 commonsourceibias.n47 gnd 0.007823f
C413 commonsourceibias.n48 gnd 0.01121f
C414 commonsourceibias.n49 gnd 0.059912f
C415 commonsourceibias.n50 gnd 0.011203f
C416 commonsourceibias.n51 gnd 0.008037f
C417 commonsourceibias.n52 gnd 0.008037f
C418 commonsourceibias.n53 gnd 0.008037f
C419 commonsourceibias.n54 gnd 0.01034f
C420 commonsourceibias.n55 gnd 0.059912f
C421 commonsourceibias.n56 gnd 0.010583f
C422 commonsourceibias.n57 gnd 0.010282f
C423 commonsourceibias.n58 gnd 0.008037f
C424 commonsourceibias.n59 gnd 0.008037f
C425 commonsourceibias.n60 gnd 0.008037f
C426 commonsourceibias.n61 gnd 0.007578f
C427 commonsourceibias.n62 gnd 0.01122f
C428 commonsourceibias.n63 gnd 0.059912f
C429 commonsourceibias.n64 gnd 0.011217f
C430 commonsourceibias.n65 gnd 0.008037f
C431 commonsourceibias.n66 gnd 0.008037f
C432 commonsourceibias.n67 gnd 0.008037f
C433 commonsourceibias.n68 gnd 0.010186f
C434 commonsourceibias.n69 gnd 0.059912f
C435 commonsourceibias.n70 gnd 0.010507f
C436 commonsourceibias.n71 gnd 0.010357f
C437 commonsourceibias.n72 gnd 0.008037f
C438 commonsourceibias.n73 gnd 0.008037f
C439 commonsourceibias.n74 gnd 0.008037f
C440 commonsourceibias.n75 gnd 0.007361f
C441 commonsourceibias.n76 gnd 0.011225f
C442 commonsourceibias.n77 gnd 0.059912f
C443 commonsourceibias.n78 gnd 0.011224f
C444 commonsourceibias.n79 gnd 0.008037f
C445 commonsourceibias.n80 gnd 0.008037f
C446 commonsourceibias.n81 gnd 0.008037f
C447 commonsourceibias.n82 gnd 0.010015f
C448 commonsourceibias.n83 gnd 0.059912f
C449 commonsourceibias.n84 gnd 0.010432f
C450 commonsourceibias.n85 gnd 0.010432f
C451 commonsourceibias.n86 gnd 0.008037f
C452 commonsourceibias.n87 gnd 0.008037f
C453 commonsourceibias.n88 gnd 0.008037f
C454 commonsourceibias.n89 gnd 0.007172f
C455 commonsourceibias.n90 gnd 0.011224f
C456 commonsourceibias.n91 gnd 0.059912f
C457 commonsourceibias.n92 gnd 0.011225f
C458 commonsourceibias.n93 gnd 0.008037f
C459 commonsourceibias.n94 gnd 0.008037f
C460 commonsourceibias.n95 gnd 0.008037f
C461 commonsourceibias.n96 gnd 0.009825f
C462 commonsourceibias.n97 gnd 0.059912f
C463 commonsourceibias.n98 gnd 0.010357f
C464 commonsourceibias.n99 gnd 0.010507f
C465 commonsourceibias.n100 gnd 0.008037f
C466 commonsourceibias.n101 gnd 0.008037f
C467 commonsourceibias.n102 gnd 0.008037f
C468 commonsourceibias.n103 gnd 0.007008f
C469 commonsourceibias.n104 gnd 0.011217f
C470 commonsourceibias.n105 gnd 0.059912f
C471 commonsourceibias.n106 gnd 0.01122f
C472 commonsourceibias.n107 gnd 0.008037f
C473 commonsourceibias.n108 gnd 0.008037f
C474 commonsourceibias.n109 gnd 0.008037f
C475 commonsourceibias.n110 gnd 0.009613f
C476 commonsourceibias.n111 gnd 0.059912f
C477 commonsourceibias.n112 gnd 0.010282f
C478 commonsourceibias.n113 gnd 0.010583f
C479 commonsourceibias.n114 gnd 0.008037f
C480 commonsourceibias.n115 gnd 0.008037f
C481 commonsourceibias.n116 gnd 0.008037f
C482 commonsourceibias.n117 gnd 0.006868f
C483 commonsourceibias.n118 gnd 0.011203f
C484 commonsourceibias.n119 gnd 0.059912f
C485 commonsourceibias.n120 gnd 0.01121f
C486 commonsourceibias.n121 gnd 0.008037f
C487 commonsourceibias.n122 gnd 0.008037f
C488 commonsourceibias.n123 gnd 0.008037f
C489 commonsourceibias.n124 gnd 0.009378f
C490 commonsourceibias.n125 gnd 0.059912f
C491 commonsourceibias.n126 gnd 0.009861f
C492 commonsourceibias.n127 gnd 0.07189f
C493 commonsourceibias.n128 gnd 0.080075f
C494 commonsourceibias.t75 gnd 0.017343f
C495 commonsourceibias.t21 gnd 0.017343f
C496 commonsourceibias.n129 gnd 0.15325f
C497 commonsourceibias.n130 gnd 0.132562f
C498 commonsourceibias.t51 gnd 0.017343f
C499 commonsourceibias.t9 gnd 0.017343f
C500 commonsourceibias.n131 gnd 0.15325f
C501 commonsourceibias.n132 gnd 0.070394f
C502 commonsourceibias.t37 gnd 0.017343f
C503 commonsourceibias.t77 gnd 0.017343f
C504 commonsourceibias.n133 gnd 0.15325f
C505 commonsourceibias.n134 gnd 0.070394f
C506 commonsourceibias.t25 gnd 0.017343f
C507 commonsourceibias.t35 gnd 0.017343f
C508 commonsourceibias.n135 gnd 0.15325f
C509 commonsourceibias.n136 gnd 0.070394f
C510 commonsourceibias.t11 gnd 0.017343f
C511 commonsourceibias.t41 gnd 0.017343f
C512 commonsourceibias.n137 gnd 0.15325f
C513 commonsourceibias.n138 gnd 0.058811f
C514 commonsourceibias.t47 gnd 0.017343f
C515 commonsourceibias.t79 gnd 0.017343f
C516 commonsourceibias.n139 gnd 0.153763f
C517 commonsourceibias.t55 gnd 0.017343f
C518 commonsourceibias.t5 gnd 0.017343f
C519 commonsourceibias.n140 gnd 0.15325f
C520 commonsourceibias.n141 gnd 0.1428f
C521 commonsourceibias.t19 gnd 0.017343f
C522 commonsourceibias.t23 gnd 0.017343f
C523 commonsourceibias.n142 gnd 0.15325f
C524 commonsourceibias.n143 gnd 0.070394f
C525 commonsourceibias.t39 gnd 0.017343f
C526 commonsourceibias.t71 gnd 0.017343f
C527 commonsourceibias.n144 gnd 0.15325f
C528 commonsourceibias.n145 gnd 0.070394f
C529 commonsourceibias.t57 gnd 0.017343f
C530 commonsourceibias.t27 gnd 0.017343f
C531 commonsourceibias.n146 gnd 0.15325f
C532 commonsourceibias.n147 gnd 0.058811f
C533 commonsourceibias.n148 gnd 0.071213f
C534 commonsourceibias.n149 gnd 0.052016f
C535 commonsourceibias.t153 gnd 0.150157f
C536 commonsourceibias.n150 gnd 0.059912f
C537 commonsourceibias.t88 gnd 0.150157f
C538 commonsourceibias.n151 gnd 0.059912f
C539 commonsourceibias.n152 gnd 0.008037f
C540 commonsourceibias.t125 gnd 0.150157f
C541 commonsourceibias.n153 gnd 0.059912f
C542 commonsourceibias.n154 gnd 0.008037f
C543 commonsourceibias.t120 gnd 0.150157f
C544 commonsourceibias.n155 gnd 0.059912f
C545 commonsourceibias.n156 gnd 0.008037f
C546 commonsourceibias.t139 gnd 0.150157f
C547 commonsourceibias.n157 gnd 0.007008f
C548 commonsourceibias.n158 gnd 0.008037f
C549 commonsourceibias.t112 gnd 0.150157f
C550 commonsourceibias.n159 gnd 0.009613f
C551 commonsourceibias.n160 gnd 0.008037f
C552 commonsourceibias.t107 gnd 0.150157f
C553 commonsourceibias.n161 gnd 0.059912f
C554 commonsourceibias.t127 gnd 0.150157f
C555 commonsourceibias.n162 gnd 0.006868f
C556 commonsourceibias.n163 gnd 0.008037f
C557 commonsourceibias.t146 gnd 0.150157f
C558 commonsourceibias.n164 gnd 0.009378f
C559 commonsourceibias.t117 gnd 0.166947f
C560 commonsourceibias.t99 gnd 0.150157f
C561 commonsourceibias.n165 gnd 0.065449f
C562 commonsourceibias.n166 gnd 0.071822f
C563 commonsourceibias.n167 gnd 0.033327f
C564 commonsourceibias.n168 gnd 0.008037f
C565 commonsourceibias.n169 gnd 0.007823f
C566 commonsourceibias.n170 gnd 0.01121f
C567 commonsourceibias.n171 gnd 0.059912f
C568 commonsourceibias.n172 gnd 0.011203f
C569 commonsourceibias.n173 gnd 0.008037f
C570 commonsourceibias.n174 gnd 0.008037f
C571 commonsourceibias.n175 gnd 0.008037f
C572 commonsourceibias.n176 gnd 0.01034f
C573 commonsourceibias.n177 gnd 0.059912f
C574 commonsourceibias.n178 gnd 0.010583f
C575 commonsourceibias.n179 gnd 0.010282f
C576 commonsourceibias.n180 gnd 0.008037f
C577 commonsourceibias.n181 gnd 0.008037f
C578 commonsourceibias.n182 gnd 0.008037f
C579 commonsourceibias.n183 gnd 0.007578f
C580 commonsourceibias.n184 gnd 0.01122f
C581 commonsourceibias.n185 gnd 0.059912f
C582 commonsourceibias.n186 gnd 0.011217f
C583 commonsourceibias.n187 gnd 0.008037f
C584 commonsourceibias.n188 gnd 0.008037f
C585 commonsourceibias.n189 gnd 0.008037f
C586 commonsourceibias.n190 gnd 0.010186f
C587 commonsourceibias.n191 gnd 0.059912f
C588 commonsourceibias.n192 gnd 0.010507f
C589 commonsourceibias.n193 gnd 0.010357f
C590 commonsourceibias.n194 gnd 0.008037f
C591 commonsourceibias.n195 gnd 0.008037f
C592 commonsourceibias.n196 gnd 0.009825f
C593 commonsourceibias.n197 gnd 0.007361f
C594 commonsourceibias.n198 gnd 0.011225f
C595 commonsourceibias.n199 gnd 0.008037f
C596 commonsourceibias.n200 gnd 0.008037f
C597 commonsourceibias.n201 gnd 0.011224f
C598 commonsourceibias.n202 gnd 0.007172f
C599 commonsourceibias.n203 gnd 0.010015f
C600 commonsourceibias.n204 gnd 0.008037f
C601 commonsourceibias.n205 gnd 0.007021f
C602 commonsourceibias.n206 gnd 0.010432f
C603 commonsourceibias.n207 gnd 0.010432f
C604 commonsourceibias.n208 gnd 0.007021f
C605 commonsourceibias.n209 gnd 0.008037f
C606 commonsourceibias.n210 gnd 0.008037f
C607 commonsourceibias.n211 gnd 0.007172f
C608 commonsourceibias.n212 gnd 0.011224f
C609 commonsourceibias.n213 gnd 0.059912f
C610 commonsourceibias.n214 gnd 0.011225f
C611 commonsourceibias.n215 gnd 0.008037f
C612 commonsourceibias.n216 gnd 0.008037f
C613 commonsourceibias.n217 gnd 0.008037f
C614 commonsourceibias.n218 gnd 0.009825f
C615 commonsourceibias.n219 gnd 0.059912f
C616 commonsourceibias.n220 gnd 0.010357f
C617 commonsourceibias.n221 gnd 0.010507f
C618 commonsourceibias.n222 gnd 0.008037f
C619 commonsourceibias.n223 gnd 0.008037f
C620 commonsourceibias.n224 gnd 0.008037f
C621 commonsourceibias.n225 gnd 0.007008f
C622 commonsourceibias.n226 gnd 0.011217f
C623 commonsourceibias.n227 gnd 0.059912f
C624 commonsourceibias.n228 gnd 0.01122f
C625 commonsourceibias.n229 gnd 0.008037f
C626 commonsourceibias.n230 gnd 0.008037f
C627 commonsourceibias.n231 gnd 0.008037f
C628 commonsourceibias.n232 gnd 0.009613f
C629 commonsourceibias.n233 gnd 0.059912f
C630 commonsourceibias.n234 gnd 0.010282f
C631 commonsourceibias.n235 gnd 0.010583f
C632 commonsourceibias.n236 gnd 0.008037f
C633 commonsourceibias.n237 gnd 0.008037f
C634 commonsourceibias.n238 gnd 0.008037f
C635 commonsourceibias.n239 gnd 0.006868f
C636 commonsourceibias.n240 gnd 0.011203f
C637 commonsourceibias.n241 gnd 0.059912f
C638 commonsourceibias.n242 gnd 0.01121f
C639 commonsourceibias.n243 gnd 0.008037f
C640 commonsourceibias.n244 gnd 0.008037f
C641 commonsourceibias.n245 gnd 0.008037f
C642 commonsourceibias.n246 gnd 0.009378f
C643 commonsourceibias.n247 gnd 0.059912f
C644 commonsourceibias.n248 gnd 0.009861f
C645 commonsourceibias.n249 gnd 0.07189f
C646 commonsourceibias.n250 gnd 0.04697f
C647 commonsourceibias.n251 gnd 0.010724f
C648 commonsourceibias.t119 gnd 0.150157f
C649 commonsourceibias.n252 gnd 0.007823f
C650 commonsourceibias.n253 gnd 0.008037f
C651 commonsourceibias.t137 gnd 0.150157f
C652 commonsourceibias.n254 gnd 0.01034f
C653 commonsourceibias.n255 gnd 0.008037f
C654 commonsourceibias.t92 gnd 0.150157f
C655 commonsourceibias.n256 gnd 0.059912f
C656 commonsourceibias.t109 gnd 0.150157f
C657 commonsourceibias.n257 gnd 0.007578f
C658 commonsourceibias.n258 gnd 0.008037f
C659 commonsourceibias.t128 gnd 0.150157f
C660 commonsourceibias.n259 gnd 0.010186f
C661 commonsourceibias.n260 gnd 0.008037f
C662 commonsourceibias.t86 gnd 0.150157f
C663 commonsourceibias.n261 gnd 0.059912f
C664 commonsourceibias.t83 gnd 0.150157f
C665 commonsourceibias.n262 gnd 0.007361f
C666 commonsourceibias.n263 gnd 0.008037f
C667 commonsourceibias.t118 gnd 0.150157f
C668 commonsourceibias.n264 gnd 0.010015f
C669 commonsourceibias.n265 gnd 0.008037f
C670 commonsourceibias.t138 gnd 0.150157f
C671 commonsourceibias.n266 gnd 0.059912f
C672 commonsourceibias.t159 gnd 0.150157f
C673 commonsourceibias.n267 gnd 0.007172f
C674 commonsourceibias.n268 gnd 0.008037f
C675 commonsourceibias.t108 gnd 0.150157f
C676 commonsourceibias.n269 gnd 0.009825f
C677 commonsourceibias.n270 gnd 0.008037f
C678 commonsourceibias.t102 gnd 0.150157f
C679 commonsourceibias.n271 gnd 0.059912f
C680 commonsourceibias.t121 gnd 0.150157f
C681 commonsourceibias.n272 gnd 0.007008f
C682 commonsourceibias.n273 gnd 0.008037f
C683 commonsourceibias.t95 gnd 0.150157f
C684 commonsourceibias.n274 gnd 0.009613f
C685 commonsourceibias.n275 gnd 0.008037f
C686 commonsourceibias.t93 gnd 0.150157f
C687 commonsourceibias.n276 gnd 0.059912f
C688 commonsourceibias.t110 gnd 0.150157f
C689 commonsourceibias.n277 gnd 0.006868f
C690 commonsourceibias.n278 gnd 0.008037f
C691 commonsourceibias.t129 gnd 0.150157f
C692 commonsourceibias.n279 gnd 0.009378f
C693 commonsourceibias.t101 gnd 0.166947f
C694 commonsourceibias.t87 gnd 0.150157f
C695 commonsourceibias.n280 gnd 0.065449f
C696 commonsourceibias.n281 gnd 0.071822f
C697 commonsourceibias.n282 gnd 0.033327f
C698 commonsourceibias.n283 gnd 0.008037f
C699 commonsourceibias.n284 gnd 0.007823f
C700 commonsourceibias.n285 gnd 0.01121f
C701 commonsourceibias.n286 gnd 0.059912f
C702 commonsourceibias.n287 gnd 0.011203f
C703 commonsourceibias.n288 gnd 0.008037f
C704 commonsourceibias.n289 gnd 0.008037f
C705 commonsourceibias.n290 gnd 0.008037f
C706 commonsourceibias.n291 gnd 0.01034f
C707 commonsourceibias.n292 gnd 0.059912f
C708 commonsourceibias.n293 gnd 0.010583f
C709 commonsourceibias.n294 gnd 0.010282f
C710 commonsourceibias.n295 gnd 0.008037f
C711 commonsourceibias.n296 gnd 0.008037f
C712 commonsourceibias.n297 gnd 0.008037f
C713 commonsourceibias.n298 gnd 0.007578f
C714 commonsourceibias.n299 gnd 0.01122f
C715 commonsourceibias.n300 gnd 0.059912f
C716 commonsourceibias.n301 gnd 0.011217f
C717 commonsourceibias.n302 gnd 0.008037f
C718 commonsourceibias.n303 gnd 0.008037f
C719 commonsourceibias.n304 gnd 0.008037f
C720 commonsourceibias.n305 gnd 0.010186f
C721 commonsourceibias.n306 gnd 0.059912f
C722 commonsourceibias.n307 gnd 0.010507f
C723 commonsourceibias.n308 gnd 0.010357f
C724 commonsourceibias.n309 gnd 0.008037f
C725 commonsourceibias.n310 gnd 0.008037f
C726 commonsourceibias.n311 gnd 0.008037f
C727 commonsourceibias.n312 gnd 0.007361f
C728 commonsourceibias.n313 gnd 0.011225f
C729 commonsourceibias.n314 gnd 0.059912f
C730 commonsourceibias.n315 gnd 0.011224f
C731 commonsourceibias.n316 gnd 0.008037f
C732 commonsourceibias.n317 gnd 0.008037f
C733 commonsourceibias.n318 gnd 0.008037f
C734 commonsourceibias.n319 gnd 0.010015f
C735 commonsourceibias.n320 gnd 0.059912f
C736 commonsourceibias.n321 gnd 0.010432f
C737 commonsourceibias.n322 gnd 0.010432f
C738 commonsourceibias.n323 gnd 0.008037f
C739 commonsourceibias.n324 gnd 0.008037f
C740 commonsourceibias.n325 gnd 0.008037f
C741 commonsourceibias.n326 gnd 0.007172f
C742 commonsourceibias.n327 gnd 0.011224f
C743 commonsourceibias.n328 gnd 0.059912f
C744 commonsourceibias.n329 gnd 0.011225f
C745 commonsourceibias.n330 gnd 0.008037f
C746 commonsourceibias.n331 gnd 0.008037f
C747 commonsourceibias.n332 gnd 0.008037f
C748 commonsourceibias.n333 gnd 0.009825f
C749 commonsourceibias.n334 gnd 0.059912f
C750 commonsourceibias.n335 gnd 0.010357f
C751 commonsourceibias.n336 gnd 0.010507f
C752 commonsourceibias.n337 gnd 0.008037f
C753 commonsourceibias.n338 gnd 0.008037f
C754 commonsourceibias.n339 gnd 0.008037f
C755 commonsourceibias.n340 gnd 0.007008f
C756 commonsourceibias.n341 gnd 0.011217f
C757 commonsourceibias.n342 gnd 0.059912f
C758 commonsourceibias.n343 gnd 0.01122f
C759 commonsourceibias.n344 gnd 0.008037f
C760 commonsourceibias.n345 gnd 0.008037f
C761 commonsourceibias.n346 gnd 0.008037f
C762 commonsourceibias.n347 gnd 0.009613f
C763 commonsourceibias.n348 gnd 0.059912f
C764 commonsourceibias.n349 gnd 0.010282f
C765 commonsourceibias.n350 gnd 0.010583f
C766 commonsourceibias.n351 gnd 0.008037f
C767 commonsourceibias.n352 gnd 0.008037f
C768 commonsourceibias.n353 gnd 0.008037f
C769 commonsourceibias.n354 gnd 0.006868f
C770 commonsourceibias.n355 gnd 0.011203f
C771 commonsourceibias.n356 gnd 0.059912f
C772 commonsourceibias.n357 gnd 0.01121f
C773 commonsourceibias.n358 gnd 0.008037f
C774 commonsourceibias.n359 gnd 0.008037f
C775 commonsourceibias.n360 gnd 0.008037f
C776 commonsourceibias.n361 gnd 0.009378f
C777 commonsourceibias.n362 gnd 0.059912f
C778 commonsourceibias.n363 gnd 0.009861f
C779 commonsourceibias.t100 gnd 0.162395f
C780 commonsourceibias.n364 gnd 0.07189f
C781 commonsourceibias.n365 gnd 0.025003f
C782 commonsourceibias.n366 gnd 0.464917f
C783 commonsourceibias.n367 gnd 0.010724f
C784 commonsourceibias.t140 gnd 0.162395f
C785 commonsourceibias.t155 gnd 0.150157f
C786 commonsourceibias.n368 gnd 0.007823f
C787 commonsourceibias.n369 gnd 0.008037f
C788 commonsourceibias.t84 gnd 0.150157f
C789 commonsourceibias.n370 gnd 0.01034f
C790 commonsourceibias.n371 gnd 0.008037f
C791 commonsourceibias.t148 gnd 0.150157f
C792 commonsourceibias.n372 gnd 0.007578f
C793 commonsourceibias.n373 gnd 0.008037f
C794 commonsourceibias.t80 gnd 0.150157f
C795 commonsourceibias.n374 gnd 0.010186f
C796 commonsourceibias.n375 gnd 0.008037f
C797 commonsourceibias.t113 gnd 0.150157f
C798 commonsourceibias.n376 gnd 0.007361f
C799 commonsourceibias.n377 gnd 0.008037f
C800 commonsourceibias.t154 gnd 0.150157f
C801 commonsourceibias.n378 gnd 0.010015f
C802 commonsourceibias.t29 gnd 0.017343f
C803 commonsourceibias.t3 gnd 0.017343f
C804 commonsourceibias.n379 gnd 0.153763f
C805 commonsourceibias.t49 gnd 0.017343f
C806 commonsourceibias.t13 gnd 0.017343f
C807 commonsourceibias.n380 gnd 0.15325f
C808 commonsourceibias.n381 gnd 0.1428f
C809 commonsourceibias.t69 gnd 0.017343f
C810 commonsourceibias.t67 gnd 0.017343f
C811 commonsourceibias.n382 gnd 0.15325f
C812 commonsourceibias.n383 gnd 0.070394f
C813 commonsourceibias.t7 gnd 0.017343f
C814 commonsourceibias.t63 gnd 0.017343f
C815 commonsourceibias.n384 gnd 0.15325f
C816 commonsourceibias.n385 gnd 0.070394f
C817 commonsourceibias.t53 gnd 0.017343f
C818 commonsourceibias.t73 gnd 0.017343f
C819 commonsourceibias.n386 gnd 0.15325f
C820 commonsourceibias.n387 gnd 0.058811f
C821 commonsourceibias.n388 gnd 0.010724f
C822 commonsourceibias.t42 gnd 0.150157f
C823 commonsourceibias.n389 gnd 0.007823f
C824 commonsourceibias.n390 gnd 0.008037f
C825 commonsourceibias.t0 gnd 0.150157f
C826 commonsourceibias.n391 gnd 0.01034f
C827 commonsourceibias.n392 gnd 0.008037f
C828 commonsourceibias.t60 gnd 0.150157f
C829 commonsourceibias.n393 gnd 0.007578f
C830 commonsourceibias.n394 gnd 0.008037f
C831 commonsourceibias.t16 gnd 0.150157f
C832 commonsourceibias.n395 gnd 0.010186f
C833 commonsourceibias.n396 gnd 0.008037f
C834 commonsourceibias.t58 gnd 0.150157f
C835 commonsourceibias.n397 gnd 0.007361f
C836 commonsourceibias.n398 gnd 0.008037f
C837 commonsourceibias.t32 gnd 0.150157f
C838 commonsourceibias.n399 gnd 0.010015f
C839 commonsourceibias.n400 gnd 0.008037f
C840 commonsourceibias.t72 gnd 0.150157f
C841 commonsourceibias.n401 gnd 0.007172f
C842 commonsourceibias.n402 gnd 0.008037f
C843 commonsourceibias.t52 gnd 0.150157f
C844 commonsourceibias.n403 gnd 0.009825f
C845 commonsourceibias.n404 gnd 0.008037f
C846 commonsourceibias.t6 gnd 0.150157f
C847 commonsourceibias.n405 gnd 0.007008f
C848 commonsourceibias.n406 gnd 0.008037f
C849 commonsourceibias.t66 gnd 0.150157f
C850 commonsourceibias.n407 gnd 0.009613f
C851 commonsourceibias.n408 gnd 0.008037f
C852 commonsourceibias.t12 gnd 0.150157f
C853 commonsourceibias.n409 gnd 0.006868f
C854 commonsourceibias.n410 gnd 0.008037f
C855 commonsourceibias.t48 gnd 0.150157f
C856 commonsourceibias.n411 gnd 0.009378f
C857 commonsourceibias.t28 gnd 0.166947f
C858 commonsourceibias.t2 gnd 0.150157f
C859 commonsourceibias.n412 gnd 0.065449f
C860 commonsourceibias.n413 gnd 0.071822f
C861 commonsourceibias.n414 gnd 0.033327f
C862 commonsourceibias.n415 gnd 0.008037f
C863 commonsourceibias.n416 gnd 0.007823f
C864 commonsourceibias.n417 gnd 0.01121f
C865 commonsourceibias.n418 gnd 0.059912f
C866 commonsourceibias.n419 gnd 0.011203f
C867 commonsourceibias.n420 gnd 0.008037f
C868 commonsourceibias.n421 gnd 0.008037f
C869 commonsourceibias.n422 gnd 0.008037f
C870 commonsourceibias.n423 gnd 0.01034f
C871 commonsourceibias.n424 gnd 0.059912f
C872 commonsourceibias.n425 gnd 0.010583f
C873 commonsourceibias.t68 gnd 0.150157f
C874 commonsourceibias.n426 gnd 0.059912f
C875 commonsourceibias.n427 gnd 0.010282f
C876 commonsourceibias.n428 gnd 0.008037f
C877 commonsourceibias.n429 gnd 0.008037f
C878 commonsourceibias.n430 gnd 0.008037f
C879 commonsourceibias.n431 gnd 0.007578f
C880 commonsourceibias.n432 gnd 0.01122f
C881 commonsourceibias.n433 gnd 0.059912f
C882 commonsourceibias.n434 gnd 0.011217f
C883 commonsourceibias.n435 gnd 0.008037f
C884 commonsourceibias.n436 gnd 0.008037f
C885 commonsourceibias.n437 gnd 0.008037f
C886 commonsourceibias.n438 gnd 0.010186f
C887 commonsourceibias.n439 gnd 0.059912f
C888 commonsourceibias.n440 gnd 0.010507f
C889 commonsourceibias.t62 gnd 0.150157f
C890 commonsourceibias.n441 gnd 0.059912f
C891 commonsourceibias.n442 gnd 0.010357f
C892 commonsourceibias.n443 gnd 0.008037f
C893 commonsourceibias.n444 gnd 0.008037f
C894 commonsourceibias.n445 gnd 0.008037f
C895 commonsourceibias.n446 gnd 0.007361f
C896 commonsourceibias.n447 gnd 0.011225f
C897 commonsourceibias.n448 gnd 0.059912f
C898 commonsourceibias.n449 gnd 0.011224f
C899 commonsourceibias.n450 gnd 0.008037f
C900 commonsourceibias.n451 gnd 0.008037f
C901 commonsourceibias.n452 gnd 0.008037f
C902 commonsourceibias.n453 gnd 0.010015f
C903 commonsourceibias.n454 gnd 0.059912f
C904 commonsourceibias.n455 gnd 0.010432f
C905 commonsourceibias.t64 gnd 0.150157f
C906 commonsourceibias.n456 gnd 0.059912f
C907 commonsourceibias.n457 gnd 0.010432f
C908 commonsourceibias.n458 gnd 0.008037f
C909 commonsourceibias.n459 gnd 0.008037f
C910 commonsourceibias.n460 gnd 0.008037f
C911 commonsourceibias.n461 gnd 0.007172f
C912 commonsourceibias.n462 gnd 0.011224f
C913 commonsourceibias.n463 gnd 0.059912f
C914 commonsourceibias.n464 gnd 0.011225f
C915 commonsourceibias.n465 gnd 0.008037f
C916 commonsourceibias.n466 gnd 0.008037f
C917 commonsourceibias.n467 gnd 0.008037f
C918 commonsourceibias.n468 gnd 0.009825f
C919 commonsourceibias.n469 gnd 0.059912f
C920 commonsourceibias.n470 gnd 0.010357f
C921 commonsourceibias.t44 gnd 0.150157f
C922 commonsourceibias.n471 gnd 0.059912f
C923 commonsourceibias.n472 gnd 0.010507f
C924 commonsourceibias.n473 gnd 0.008037f
C925 commonsourceibias.n474 gnd 0.008037f
C926 commonsourceibias.n475 gnd 0.008037f
C927 commonsourceibias.n476 gnd 0.007008f
C928 commonsourceibias.n477 gnd 0.011217f
C929 commonsourceibias.n478 gnd 0.059912f
C930 commonsourceibias.n479 gnd 0.01122f
C931 commonsourceibias.n480 gnd 0.008037f
C932 commonsourceibias.n481 gnd 0.008037f
C933 commonsourceibias.n482 gnd 0.008037f
C934 commonsourceibias.n483 gnd 0.009613f
C935 commonsourceibias.n484 gnd 0.059912f
C936 commonsourceibias.n485 gnd 0.010282f
C937 commonsourceibias.t30 gnd 0.150157f
C938 commonsourceibias.n486 gnd 0.059912f
C939 commonsourceibias.n487 gnd 0.010583f
C940 commonsourceibias.n488 gnd 0.008037f
C941 commonsourceibias.n489 gnd 0.008037f
C942 commonsourceibias.n490 gnd 0.008037f
C943 commonsourceibias.n491 gnd 0.006868f
C944 commonsourceibias.n492 gnd 0.011203f
C945 commonsourceibias.n493 gnd 0.059912f
C946 commonsourceibias.n494 gnd 0.01121f
C947 commonsourceibias.n495 gnd 0.008037f
C948 commonsourceibias.n496 gnd 0.008037f
C949 commonsourceibias.n497 gnd 0.008037f
C950 commonsourceibias.n498 gnd 0.009378f
C951 commonsourceibias.n499 gnd 0.059912f
C952 commonsourceibias.n500 gnd 0.009861f
C953 commonsourceibias.t14 gnd 0.162395f
C954 commonsourceibias.n501 gnd 0.07189f
C955 commonsourceibias.n502 gnd 0.080075f
C956 commonsourceibias.t43 gnd 0.017343f
C957 commonsourceibias.t15 gnd 0.017343f
C958 commonsourceibias.n503 gnd 0.15325f
C959 commonsourceibias.n504 gnd 0.132562f
C960 commonsourceibias.t31 gnd 0.017343f
C961 commonsourceibias.t1 gnd 0.017343f
C962 commonsourceibias.n505 gnd 0.15325f
C963 commonsourceibias.n506 gnd 0.070394f
C964 commonsourceibias.t17 gnd 0.017343f
C965 commonsourceibias.t61 gnd 0.017343f
C966 commonsourceibias.n507 gnd 0.15325f
C967 commonsourceibias.n508 gnd 0.070394f
C968 commonsourceibias.t59 gnd 0.017343f
C969 commonsourceibias.t45 gnd 0.017343f
C970 commonsourceibias.n509 gnd 0.15325f
C971 commonsourceibias.n510 gnd 0.070394f
C972 commonsourceibias.t65 gnd 0.017343f
C973 commonsourceibias.t33 gnd 0.017343f
C974 commonsourceibias.n511 gnd 0.15325f
C975 commonsourceibias.n512 gnd 0.058811f
C976 commonsourceibias.n513 gnd 0.071213f
C977 commonsourceibias.n514 gnd 0.052016f
C978 commonsourceibias.t82 gnd 0.150157f
C979 commonsourceibias.n515 gnd 0.059912f
C980 commonsourceibias.n516 gnd 0.008037f
C981 commonsourceibias.t147 gnd 0.150157f
C982 commonsourceibias.n517 gnd 0.059912f
C983 commonsourceibias.n518 gnd 0.008037f
C984 commonsourceibias.t143 gnd 0.150157f
C985 commonsourceibias.n519 gnd 0.059912f
C986 commonsourceibias.n520 gnd 0.008037f
C987 commonsourceibias.t158 gnd 0.150157f
C988 commonsourceibias.n521 gnd 0.007008f
C989 commonsourceibias.n522 gnd 0.008037f
C990 commonsourceibias.t104 gnd 0.150157f
C991 commonsourceibias.n523 gnd 0.009613f
C992 commonsourceibias.n524 gnd 0.008037f
C993 commonsourceibias.t133 gnd 0.150157f
C994 commonsourceibias.n525 gnd 0.006868f
C995 commonsourceibias.n526 gnd 0.008037f
C996 commonsourceibias.t150 gnd 0.150157f
C997 commonsourceibias.n527 gnd 0.009378f
C998 commonsourceibias.t123 gnd 0.166947f
C999 commonsourceibias.t103 gnd 0.150157f
C1000 commonsourceibias.n528 gnd 0.065449f
C1001 commonsourceibias.n529 gnd 0.071822f
C1002 commonsourceibias.n530 gnd 0.033327f
C1003 commonsourceibias.n531 gnd 0.008037f
C1004 commonsourceibias.n532 gnd 0.007823f
C1005 commonsourceibias.n533 gnd 0.01121f
C1006 commonsourceibias.n534 gnd 0.059912f
C1007 commonsourceibias.n535 gnd 0.011203f
C1008 commonsourceibias.n536 gnd 0.008037f
C1009 commonsourceibias.n537 gnd 0.008037f
C1010 commonsourceibias.n538 gnd 0.008037f
C1011 commonsourceibias.n539 gnd 0.01034f
C1012 commonsourceibias.n540 gnd 0.059912f
C1013 commonsourceibias.n541 gnd 0.010583f
C1014 commonsourceibias.t114 gnd 0.150157f
C1015 commonsourceibias.n542 gnd 0.059912f
C1016 commonsourceibias.n543 gnd 0.010282f
C1017 commonsourceibias.n544 gnd 0.008037f
C1018 commonsourceibias.n545 gnd 0.008037f
C1019 commonsourceibias.n546 gnd 0.008037f
C1020 commonsourceibias.n547 gnd 0.007578f
C1021 commonsourceibias.n548 gnd 0.01122f
C1022 commonsourceibias.n549 gnd 0.059912f
C1023 commonsourceibias.n550 gnd 0.011217f
C1024 commonsourceibias.n551 gnd 0.008037f
C1025 commonsourceibias.n552 gnd 0.008037f
C1026 commonsourceibias.n553 gnd 0.008037f
C1027 commonsourceibias.n554 gnd 0.010186f
C1028 commonsourceibias.n555 gnd 0.059912f
C1029 commonsourceibias.n556 gnd 0.010507f
C1030 commonsourceibias.n557 gnd 0.010357f
C1031 commonsourceibias.n558 gnd 0.008037f
C1032 commonsourceibias.n559 gnd 0.008037f
C1033 commonsourceibias.n560 gnd 0.009825f
C1034 commonsourceibias.n561 gnd 0.007361f
C1035 commonsourceibias.n562 gnd 0.011225f
C1036 commonsourceibias.n563 gnd 0.008037f
C1037 commonsourceibias.n564 gnd 0.008037f
C1038 commonsourceibias.n565 gnd 0.011224f
C1039 commonsourceibias.n566 gnd 0.007172f
C1040 commonsourceibias.n567 gnd 0.010015f
C1041 commonsourceibias.n568 gnd 0.008037f
C1042 commonsourceibias.n569 gnd 0.007021f
C1043 commonsourceibias.n570 gnd 0.010432f
C1044 commonsourceibias.t85 gnd 0.150157f
C1045 commonsourceibias.n571 gnd 0.059912f
C1046 commonsourceibias.n572 gnd 0.010432f
C1047 commonsourceibias.n573 gnd 0.007021f
C1048 commonsourceibias.n574 gnd 0.008037f
C1049 commonsourceibias.n575 gnd 0.008037f
C1050 commonsourceibias.n576 gnd 0.007172f
C1051 commonsourceibias.n577 gnd 0.011224f
C1052 commonsourceibias.n578 gnd 0.059912f
C1053 commonsourceibias.n579 gnd 0.011225f
C1054 commonsourceibias.n580 gnd 0.008037f
C1055 commonsourceibias.n581 gnd 0.008037f
C1056 commonsourceibias.n582 gnd 0.008037f
C1057 commonsourceibias.n583 gnd 0.009825f
C1058 commonsourceibias.n584 gnd 0.059912f
C1059 commonsourceibias.n585 gnd 0.010357f
C1060 commonsourceibias.t89 gnd 0.150157f
C1061 commonsourceibias.n586 gnd 0.059912f
C1062 commonsourceibias.n587 gnd 0.010507f
C1063 commonsourceibias.n588 gnd 0.008037f
C1064 commonsourceibias.n589 gnd 0.008037f
C1065 commonsourceibias.n590 gnd 0.008037f
C1066 commonsourceibias.n591 gnd 0.007008f
C1067 commonsourceibias.n592 gnd 0.011217f
C1068 commonsourceibias.n593 gnd 0.059912f
C1069 commonsourceibias.n594 gnd 0.01122f
C1070 commonsourceibias.n595 gnd 0.008037f
C1071 commonsourceibias.n596 gnd 0.008037f
C1072 commonsourceibias.n597 gnd 0.008037f
C1073 commonsourceibias.n598 gnd 0.009613f
C1074 commonsourceibias.n599 gnd 0.059912f
C1075 commonsourceibias.n600 gnd 0.010282f
C1076 commonsourceibias.t130 gnd 0.150157f
C1077 commonsourceibias.n601 gnd 0.059912f
C1078 commonsourceibias.n602 gnd 0.010583f
C1079 commonsourceibias.n603 gnd 0.008037f
C1080 commonsourceibias.n604 gnd 0.008037f
C1081 commonsourceibias.n605 gnd 0.008037f
C1082 commonsourceibias.n606 gnd 0.006868f
C1083 commonsourceibias.n607 gnd 0.011203f
C1084 commonsourceibias.n608 gnd 0.059912f
C1085 commonsourceibias.n609 gnd 0.01121f
C1086 commonsourceibias.n610 gnd 0.008037f
C1087 commonsourceibias.n611 gnd 0.008037f
C1088 commonsourceibias.n612 gnd 0.008037f
C1089 commonsourceibias.n613 gnd 0.009378f
C1090 commonsourceibias.n614 gnd 0.059912f
C1091 commonsourceibias.n615 gnd 0.009861f
C1092 commonsourceibias.n616 gnd 0.07189f
C1093 commonsourceibias.n617 gnd 0.04697f
C1094 commonsourceibias.n618 gnd 0.010724f
C1095 commonsourceibias.t142 gnd 0.150157f
C1096 commonsourceibias.n619 gnd 0.007823f
C1097 commonsourceibias.n620 gnd 0.008037f
C1098 commonsourceibias.t156 gnd 0.150157f
C1099 commonsourceibias.n621 gnd 0.01034f
C1100 commonsourceibias.n622 gnd 0.008037f
C1101 commonsourceibias.t132 gnd 0.150157f
C1102 commonsourceibias.n623 gnd 0.007578f
C1103 commonsourceibias.n624 gnd 0.008037f
C1104 commonsourceibias.t149 gnd 0.150157f
C1105 commonsourceibias.n625 gnd 0.010186f
C1106 commonsourceibias.n626 gnd 0.008037f
C1107 commonsourceibias.t97 gnd 0.150157f
C1108 commonsourceibias.n627 gnd 0.007361f
C1109 commonsourceibias.n628 gnd 0.008037f
C1110 commonsourceibias.t141 gnd 0.150157f
C1111 commonsourceibias.n629 gnd 0.010015f
C1112 commonsourceibias.n630 gnd 0.008037f
C1113 commonsourceibias.t152 gnd 0.150157f
C1114 commonsourceibias.n631 gnd 0.007172f
C1115 commonsourceibias.n632 gnd 0.008037f
C1116 commonsourceibias.t131 gnd 0.150157f
C1117 commonsourceibias.n633 gnd 0.009825f
C1118 commonsourceibias.n634 gnd 0.008037f
C1119 commonsourceibias.t145 gnd 0.150157f
C1120 commonsourceibias.n635 gnd 0.007008f
C1121 commonsourceibias.n636 gnd 0.008037f
C1122 commonsourceibias.t91 gnd 0.150157f
C1123 commonsourceibias.n637 gnd 0.009613f
C1124 commonsourceibias.n638 gnd 0.008037f
C1125 commonsourceibias.t116 gnd 0.150157f
C1126 commonsourceibias.n639 gnd 0.006868f
C1127 commonsourceibias.n640 gnd 0.008037f
C1128 commonsourceibias.t134 gnd 0.150157f
C1129 commonsourceibias.n641 gnd 0.009378f
C1130 commonsourceibias.t106 gnd 0.166947f
C1131 commonsourceibias.t90 gnd 0.150157f
C1132 commonsourceibias.n642 gnd 0.065449f
C1133 commonsourceibias.n643 gnd 0.071822f
C1134 commonsourceibias.n644 gnd 0.033327f
C1135 commonsourceibias.n645 gnd 0.008037f
C1136 commonsourceibias.n646 gnd 0.007823f
C1137 commonsourceibias.n647 gnd 0.01121f
C1138 commonsourceibias.n648 gnd 0.059912f
C1139 commonsourceibias.n649 gnd 0.011203f
C1140 commonsourceibias.n650 gnd 0.008037f
C1141 commonsourceibias.n651 gnd 0.008037f
C1142 commonsourceibias.n652 gnd 0.008037f
C1143 commonsourceibias.n653 gnd 0.01034f
C1144 commonsourceibias.n654 gnd 0.059912f
C1145 commonsourceibias.n655 gnd 0.010583f
C1146 commonsourceibias.t96 gnd 0.150157f
C1147 commonsourceibias.n656 gnd 0.059912f
C1148 commonsourceibias.n657 gnd 0.010282f
C1149 commonsourceibias.n658 gnd 0.008037f
C1150 commonsourceibias.n659 gnd 0.008037f
C1151 commonsourceibias.n660 gnd 0.008037f
C1152 commonsourceibias.n661 gnd 0.007578f
C1153 commonsourceibias.n662 gnd 0.01122f
C1154 commonsourceibias.n663 gnd 0.059912f
C1155 commonsourceibias.n664 gnd 0.011217f
C1156 commonsourceibias.n665 gnd 0.008037f
C1157 commonsourceibias.n666 gnd 0.008037f
C1158 commonsourceibias.n667 gnd 0.008037f
C1159 commonsourceibias.n668 gnd 0.010186f
C1160 commonsourceibias.n669 gnd 0.059912f
C1161 commonsourceibias.n670 gnd 0.010507f
C1162 commonsourceibias.t124 gnd 0.150157f
C1163 commonsourceibias.n671 gnd 0.059912f
C1164 commonsourceibias.n672 gnd 0.010357f
C1165 commonsourceibias.n673 gnd 0.008037f
C1166 commonsourceibias.n674 gnd 0.008037f
C1167 commonsourceibias.n675 gnd 0.008037f
C1168 commonsourceibias.n676 gnd 0.007361f
C1169 commonsourceibias.n677 gnd 0.011225f
C1170 commonsourceibias.n678 gnd 0.059912f
C1171 commonsourceibias.n679 gnd 0.011224f
C1172 commonsourceibias.n680 gnd 0.008037f
C1173 commonsourceibias.n681 gnd 0.008037f
C1174 commonsourceibias.n682 gnd 0.008037f
C1175 commonsourceibias.n683 gnd 0.010015f
C1176 commonsourceibias.n684 gnd 0.059912f
C1177 commonsourceibias.n685 gnd 0.010432f
C1178 commonsourceibias.t157 gnd 0.150157f
C1179 commonsourceibias.n686 gnd 0.059912f
C1180 commonsourceibias.n687 gnd 0.010432f
C1181 commonsourceibias.n688 gnd 0.008037f
C1182 commonsourceibias.n689 gnd 0.008037f
C1183 commonsourceibias.n690 gnd 0.008037f
C1184 commonsourceibias.n691 gnd 0.007172f
C1185 commonsourceibias.n692 gnd 0.011224f
C1186 commonsourceibias.n693 gnd 0.059912f
C1187 commonsourceibias.n694 gnd 0.011225f
C1188 commonsourceibias.n695 gnd 0.008037f
C1189 commonsourceibias.n696 gnd 0.008037f
C1190 commonsourceibias.n697 gnd 0.008037f
C1191 commonsourceibias.n698 gnd 0.009825f
C1192 commonsourceibias.n699 gnd 0.059912f
C1193 commonsourceibias.n700 gnd 0.010357f
C1194 commonsourceibias.t81 gnd 0.150157f
C1195 commonsourceibias.n701 gnd 0.059912f
C1196 commonsourceibias.n702 gnd 0.010507f
C1197 commonsourceibias.n703 gnd 0.008037f
C1198 commonsourceibias.n704 gnd 0.008037f
C1199 commonsourceibias.n705 gnd 0.008037f
C1200 commonsourceibias.n706 gnd 0.007008f
C1201 commonsourceibias.n707 gnd 0.011217f
C1202 commonsourceibias.n708 gnd 0.059912f
C1203 commonsourceibias.n709 gnd 0.01122f
C1204 commonsourceibias.n710 gnd 0.008037f
C1205 commonsourceibias.n711 gnd 0.008037f
C1206 commonsourceibias.n712 gnd 0.008037f
C1207 commonsourceibias.n713 gnd 0.009613f
C1208 commonsourceibias.n714 gnd 0.059912f
C1209 commonsourceibias.n715 gnd 0.010282f
C1210 commonsourceibias.t111 gnd 0.150157f
C1211 commonsourceibias.n716 gnd 0.059912f
C1212 commonsourceibias.n717 gnd 0.010583f
C1213 commonsourceibias.n718 gnd 0.008037f
C1214 commonsourceibias.n719 gnd 0.008037f
C1215 commonsourceibias.n720 gnd 0.008037f
C1216 commonsourceibias.n721 gnd 0.006868f
C1217 commonsourceibias.n722 gnd 0.011203f
C1218 commonsourceibias.n723 gnd 0.059912f
C1219 commonsourceibias.n724 gnd 0.01121f
C1220 commonsourceibias.n725 gnd 0.008037f
C1221 commonsourceibias.n726 gnd 0.008037f
C1222 commonsourceibias.n727 gnd 0.008037f
C1223 commonsourceibias.n728 gnd 0.009378f
C1224 commonsourceibias.n729 gnd 0.059912f
C1225 commonsourceibias.n730 gnd 0.009861f
C1226 commonsourceibias.t122 gnd 0.162395f
C1227 commonsourceibias.n731 gnd 0.07189f
C1228 commonsourceibias.n732 gnd 0.025003f
C1229 commonsourceibias.n733 gnd 0.221951f
C1230 commonsourceibias.n734 gnd 4.85761f
C1231 diffpairibias.t27 gnd 0.090128f
C1232 diffpairibias.t23 gnd 0.08996f
C1233 diffpairibias.n0 gnd 0.105991f
C1234 diffpairibias.t28 gnd 0.08996f
C1235 diffpairibias.n1 gnd 0.051736f
C1236 diffpairibias.t25 gnd 0.08996f
C1237 diffpairibias.n2 gnd 0.051736f
C1238 diffpairibias.t29 gnd 0.08996f
C1239 diffpairibias.n3 gnd 0.041084f
C1240 diffpairibias.t15 gnd 0.086371f
C1241 diffpairibias.t1 gnd 0.085993f
C1242 diffpairibias.n4 gnd 0.13579f
C1243 diffpairibias.t11 gnd 0.085993f
C1244 diffpairibias.n5 gnd 0.072463f
C1245 diffpairibias.t13 gnd 0.085993f
C1246 diffpairibias.n6 gnd 0.072463f
C1247 diffpairibias.t7 gnd 0.085993f
C1248 diffpairibias.n7 gnd 0.072463f
C1249 diffpairibias.t3 gnd 0.085993f
C1250 diffpairibias.n8 gnd 0.072463f
C1251 diffpairibias.t17 gnd 0.085993f
C1252 diffpairibias.n9 gnd 0.072463f
C1253 diffpairibias.t5 gnd 0.085993f
C1254 diffpairibias.n10 gnd 0.072463f
C1255 diffpairibias.t19 gnd 0.085993f
C1256 diffpairibias.n11 gnd 0.072463f
C1257 diffpairibias.t9 gnd 0.085993f
C1258 diffpairibias.n12 gnd 0.102883f
C1259 diffpairibias.t14 gnd 0.086899f
C1260 diffpairibias.t0 gnd 0.086748f
C1261 diffpairibias.n13 gnd 0.094648f
C1262 diffpairibias.t10 gnd 0.086748f
C1263 diffpairibias.n14 gnd 0.052262f
C1264 diffpairibias.t12 gnd 0.086748f
C1265 diffpairibias.n15 gnd 0.052262f
C1266 diffpairibias.t6 gnd 0.086748f
C1267 diffpairibias.n16 gnd 0.052262f
C1268 diffpairibias.t2 gnd 0.086748f
C1269 diffpairibias.n17 gnd 0.052262f
C1270 diffpairibias.t16 gnd 0.086748f
C1271 diffpairibias.n18 gnd 0.052262f
C1272 diffpairibias.t4 gnd 0.086748f
C1273 diffpairibias.n19 gnd 0.052262f
C1274 diffpairibias.t18 gnd 0.086748f
C1275 diffpairibias.n20 gnd 0.052262f
C1276 diffpairibias.t8 gnd 0.086748f
C1277 diffpairibias.n21 gnd 0.061849f
C1278 diffpairibias.n22 gnd 0.233513f
C1279 diffpairibias.t20 gnd 0.08996f
C1280 diffpairibias.n23 gnd 0.051747f
C1281 diffpairibias.t26 gnd 0.08996f
C1282 diffpairibias.n24 gnd 0.051736f
C1283 diffpairibias.t22 gnd 0.08996f
C1284 diffpairibias.n25 gnd 0.051736f
C1285 diffpairibias.t21 gnd 0.08996f
C1286 diffpairibias.n26 gnd 0.051736f
C1287 diffpairibias.t24 gnd 0.08996f
C1288 diffpairibias.n27 gnd 0.04729f
C1289 diffpairibias.n28 gnd 0.047711f
C1290 outputibias.t10 gnd 0.11477f
C1291 outputibias.t8 gnd 0.115567f
C1292 outputibias.n0 gnd 0.130108f
C1293 outputibias.n1 gnd 0.001372f
C1294 outputibias.n2 gnd 9.76e-19
C1295 outputibias.n3 gnd 5.24e-19
C1296 outputibias.n4 gnd 0.001239f
C1297 outputibias.n5 gnd 5.55e-19
C1298 outputibias.n6 gnd 9.76e-19
C1299 outputibias.n7 gnd 5.24e-19
C1300 outputibias.n8 gnd 0.001239f
C1301 outputibias.n9 gnd 5.55e-19
C1302 outputibias.n10 gnd 0.004176f
C1303 outputibias.t5 gnd 0.00202f
C1304 outputibias.n11 gnd 9.3e-19
C1305 outputibias.n12 gnd 7.32e-19
C1306 outputibias.n13 gnd 5.24e-19
C1307 outputibias.n14 gnd 0.02322f
C1308 outputibias.n15 gnd 9.76e-19
C1309 outputibias.n16 gnd 5.24e-19
C1310 outputibias.n17 gnd 5.55e-19
C1311 outputibias.n18 gnd 0.001239f
C1312 outputibias.n19 gnd 0.001239f
C1313 outputibias.n20 gnd 5.55e-19
C1314 outputibias.n21 gnd 5.24e-19
C1315 outputibias.n22 gnd 9.76e-19
C1316 outputibias.n23 gnd 9.76e-19
C1317 outputibias.n24 gnd 5.24e-19
C1318 outputibias.n25 gnd 5.55e-19
C1319 outputibias.n26 gnd 0.001239f
C1320 outputibias.n27 gnd 0.002683f
C1321 outputibias.n28 gnd 5.55e-19
C1322 outputibias.n29 gnd 5.24e-19
C1323 outputibias.n30 gnd 0.002256f
C1324 outputibias.n31 gnd 0.005781f
C1325 outputibias.n32 gnd 0.001372f
C1326 outputibias.n33 gnd 9.76e-19
C1327 outputibias.n34 gnd 5.24e-19
C1328 outputibias.n35 gnd 0.001239f
C1329 outputibias.n36 gnd 5.55e-19
C1330 outputibias.n37 gnd 9.76e-19
C1331 outputibias.n38 gnd 5.24e-19
C1332 outputibias.n39 gnd 0.001239f
C1333 outputibias.n40 gnd 5.55e-19
C1334 outputibias.n41 gnd 0.004176f
C1335 outputibias.t3 gnd 0.00202f
C1336 outputibias.n42 gnd 9.3e-19
C1337 outputibias.n43 gnd 7.32e-19
C1338 outputibias.n44 gnd 5.24e-19
C1339 outputibias.n45 gnd 0.02322f
C1340 outputibias.n46 gnd 9.76e-19
C1341 outputibias.n47 gnd 5.24e-19
C1342 outputibias.n48 gnd 5.55e-19
C1343 outputibias.n49 gnd 0.001239f
C1344 outputibias.n50 gnd 0.001239f
C1345 outputibias.n51 gnd 5.55e-19
C1346 outputibias.n52 gnd 5.24e-19
C1347 outputibias.n53 gnd 9.76e-19
C1348 outputibias.n54 gnd 9.76e-19
C1349 outputibias.n55 gnd 5.24e-19
C1350 outputibias.n56 gnd 5.55e-19
C1351 outputibias.n57 gnd 0.001239f
C1352 outputibias.n58 gnd 0.002683f
C1353 outputibias.n59 gnd 5.55e-19
C1354 outputibias.n60 gnd 5.24e-19
C1355 outputibias.n61 gnd 0.002256f
C1356 outputibias.n62 gnd 0.005197f
C1357 outputibias.n63 gnd 0.121892f
C1358 outputibias.n64 gnd 0.001372f
C1359 outputibias.n65 gnd 9.76e-19
C1360 outputibias.n66 gnd 5.24e-19
C1361 outputibias.n67 gnd 0.001239f
C1362 outputibias.n68 gnd 5.55e-19
C1363 outputibias.n69 gnd 9.76e-19
C1364 outputibias.n70 gnd 5.24e-19
C1365 outputibias.n71 gnd 0.001239f
C1366 outputibias.n72 gnd 5.55e-19
C1367 outputibias.n73 gnd 0.004176f
C1368 outputibias.t1 gnd 0.00202f
C1369 outputibias.n74 gnd 9.3e-19
C1370 outputibias.n75 gnd 7.32e-19
C1371 outputibias.n76 gnd 5.24e-19
C1372 outputibias.n77 gnd 0.02322f
C1373 outputibias.n78 gnd 9.76e-19
C1374 outputibias.n79 gnd 5.24e-19
C1375 outputibias.n80 gnd 5.55e-19
C1376 outputibias.n81 gnd 0.001239f
C1377 outputibias.n82 gnd 0.001239f
C1378 outputibias.n83 gnd 5.55e-19
C1379 outputibias.n84 gnd 5.24e-19
C1380 outputibias.n85 gnd 9.76e-19
C1381 outputibias.n86 gnd 9.76e-19
C1382 outputibias.n87 gnd 5.24e-19
C1383 outputibias.n88 gnd 5.55e-19
C1384 outputibias.n89 gnd 0.001239f
C1385 outputibias.n90 gnd 0.002683f
C1386 outputibias.n91 gnd 5.55e-19
C1387 outputibias.n92 gnd 5.24e-19
C1388 outputibias.n93 gnd 0.002256f
C1389 outputibias.n94 gnd 0.005197f
C1390 outputibias.n95 gnd 0.064513f
C1391 outputibias.n96 gnd 0.001372f
C1392 outputibias.n97 gnd 9.76e-19
C1393 outputibias.n98 gnd 5.24e-19
C1394 outputibias.n99 gnd 0.001239f
C1395 outputibias.n100 gnd 5.55e-19
C1396 outputibias.n101 gnd 9.76e-19
C1397 outputibias.n102 gnd 5.24e-19
C1398 outputibias.n103 gnd 0.001239f
C1399 outputibias.n104 gnd 5.55e-19
C1400 outputibias.n105 gnd 0.004176f
C1401 outputibias.t7 gnd 0.00202f
C1402 outputibias.n106 gnd 9.3e-19
C1403 outputibias.n107 gnd 7.32e-19
C1404 outputibias.n108 gnd 5.24e-19
C1405 outputibias.n109 gnd 0.02322f
C1406 outputibias.n110 gnd 9.76e-19
C1407 outputibias.n111 gnd 5.24e-19
C1408 outputibias.n112 gnd 5.55e-19
C1409 outputibias.n113 gnd 0.001239f
C1410 outputibias.n114 gnd 0.001239f
C1411 outputibias.n115 gnd 5.55e-19
C1412 outputibias.n116 gnd 5.24e-19
C1413 outputibias.n117 gnd 9.76e-19
C1414 outputibias.n118 gnd 9.76e-19
C1415 outputibias.n119 gnd 5.24e-19
C1416 outputibias.n120 gnd 5.55e-19
C1417 outputibias.n121 gnd 0.001239f
C1418 outputibias.n122 gnd 0.002683f
C1419 outputibias.n123 gnd 5.55e-19
C1420 outputibias.n124 gnd 5.24e-19
C1421 outputibias.n125 gnd 0.002256f
C1422 outputibias.n126 gnd 0.005197f
C1423 outputibias.n127 gnd 0.084814f
C1424 outputibias.t6 gnd 0.108319f
C1425 outputibias.t0 gnd 0.108319f
C1426 outputibias.t2 gnd 0.108319f
C1427 outputibias.t4 gnd 0.109238f
C1428 outputibias.n128 gnd 0.134674f
C1429 outputibias.n129 gnd 0.07244f
C1430 outputibias.n130 gnd 0.079818f
C1431 outputibias.n131 gnd 0.164901f
C1432 outputibias.t11 gnd 0.11477f
C1433 outputibias.n132 gnd 0.067481f
C1434 outputibias.t9 gnd 0.11477f
C1435 outputibias.n133 gnd 0.065115f
C1436 outputibias.n134 gnd 0.029159f
C1437 CSoutput.n0 gnd 0.048248f
C1438 CSoutput.t217 gnd 0.31915f
C1439 CSoutput.n1 gnd 0.144112f
C1440 CSoutput.n2 gnd 0.048248f
C1441 CSoutput.t200 gnd 0.31915f
C1442 CSoutput.n3 gnd 0.03824f
C1443 CSoutput.n4 gnd 0.048248f
C1444 CSoutput.t209 gnd 0.31915f
C1445 CSoutput.n5 gnd 0.032975f
C1446 CSoutput.n6 gnd 0.048248f
C1447 CSoutput.t220 gnd 0.31915f
C1448 CSoutput.t219 gnd 0.31915f
C1449 CSoutput.n7 gnd 0.142542f
C1450 CSoutput.n8 gnd 0.048248f
C1451 CSoutput.t206 gnd 0.31915f
C1452 CSoutput.n9 gnd 0.03144f
C1453 CSoutput.n10 gnd 0.048248f
C1454 CSoutput.t212 gnd 0.31915f
C1455 CSoutput.t215 gnd 0.31915f
C1456 CSoutput.n11 gnd 0.142542f
C1457 CSoutput.n12 gnd 0.048248f
C1458 CSoutput.t203 gnd 0.31915f
C1459 CSoutput.n13 gnd 0.032975f
C1460 CSoutput.n14 gnd 0.048248f
C1461 CSoutput.t202 gnd 0.31915f
C1462 CSoutput.t213 gnd 0.31915f
C1463 CSoutput.n15 gnd 0.142542f
C1464 CSoutput.n16 gnd 0.048248f
C1465 CSoutput.t218 gnd 0.31915f
C1466 CSoutput.n17 gnd 0.035219f
C1467 CSoutput.t204 gnd 0.381393f
C1468 CSoutput.t201 gnd 0.31915f
C1469 CSoutput.n18 gnd 0.18197f
C1470 CSoutput.n19 gnd 0.176574f
C1471 CSoutput.n20 gnd 0.204847f
C1472 CSoutput.n21 gnd 0.048248f
C1473 CSoutput.n22 gnd 0.040268f
C1474 CSoutput.n23 gnd 0.142542f
C1475 CSoutput.n24 gnd 0.038818f
C1476 CSoutput.n25 gnd 0.03824f
C1477 CSoutput.n26 gnd 0.048248f
C1478 CSoutput.n27 gnd 0.048248f
C1479 CSoutput.n28 gnd 0.039959f
C1480 CSoutput.n29 gnd 0.033926f
C1481 CSoutput.n30 gnd 0.145715f
C1482 CSoutput.n31 gnd 0.034393f
C1483 CSoutput.n32 gnd 0.048248f
C1484 CSoutput.n33 gnd 0.048248f
C1485 CSoutput.n34 gnd 0.048248f
C1486 CSoutput.n35 gnd 0.039533f
C1487 CSoutput.n36 gnd 0.142542f
C1488 CSoutput.n37 gnd 0.037808f
C1489 CSoutput.n38 gnd 0.03925f
C1490 CSoutput.n39 gnd 0.048248f
C1491 CSoutput.n40 gnd 0.048248f
C1492 CSoutput.n41 gnd 0.04026f
C1493 CSoutput.n42 gnd 0.036798f
C1494 CSoutput.n43 gnd 0.142542f
C1495 CSoutput.n44 gnd 0.037731f
C1496 CSoutput.n45 gnd 0.048248f
C1497 CSoutput.n46 gnd 0.048248f
C1498 CSoutput.n47 gnd 0.048248f
C1499 CSoutput.n48 gnd 0.037731f
C1500 CSoutput.n49 gnd 0.142542f
C1501 CSoutput.n50 gnd 0.036798f
C1502 CSoutput.n51 gnd 0.04026f
C1503 CSoutput.n52 gnd 0.048248f
C1504 CSoutput.n53 gnd 0.048248f
C1505 CSoutput.n54 gnd 0.03925f
C1506 CSoutput.n55 gnd 0.037808f
C1507 CSoutput.n56 gnd 0.142542f
C1508 CSoutput.n57 gnd 0.039533f
C1509 CSoutput.n58 gnd 0.048248f
C1510 CSoutput.n59 gnd 0.048248f
C1511 CSoutput.n60 gnd 0.048248f
C1512 CSoutput.n61 gnd 0.034393f
C1513 CSoutput.n62 gnd 0.145715f
C1514 CSoutput.n63 gnd 0.033926f
C1515 CSoutput.t221 gnd 0.31915f
C1516 CSoutput.n64 gnd 0.142542f
C1517 CSoutput.n65 gnd 0.039959f
C1518 CSoutput.n66 gnd 0.048248f
C1519 CSoutput.n67 gnd 0.048248f
C1520 CSoutput.n68 gnd 0.048248f
C1521 CSoutput.n69 gnd 0.038818f
C1522 CSoutput.n70 gnd 0.142542f
C1523 CSoutput.n71 gnd 0.040268f
C1524 CSoutput.n72 gnd 0.035219f
C1525 CSoutput.n73 gnd 0.048248f
C1526 CSoutput.n74 gnd 0.048248f
C1527 CSoutput.n75 gnd 0.036525f
C1528 CSoutput.n76 gnd 0.021692f
C1529 CSoutput.t207 gnd 0.358588f
C1530 CSoutput.n77 gnd 0.178132f
C1531 CSoutput.n78 gnd 0.762212f
C1532 CSoutput.t168 gnd 0.060183f
C1533 CSoutput.t103 gnd 0.060183f
C1534 CSoutput.n79 gnd 0.465954f
C1535 CSoutput.t63 gnd 0.060183f
C1536 CSoutput.t145 gnd 0.060183f
C1537 CSoutput.n80 gnd 0.465123f
C1538 CSoutput.n81 gnd 0.472099f
C1539 CSoutput.t73 gnd 0.060183f
C1540 CSoutput.t126 gnd 0.060183f
C1541 CSoutput.n82 gnd 0.465123f
C1542 CSoutput.n83 gnd 0.232631f
C1543 CSoutput.t92 gnd 0.060183f
C1544 CSoutput.t112 gnd 0.060183f
C1545 CSoutput.n84 gnd 0.465123f
C1546 CSoutput.n85 gnd 0.232631f
C1547 CSoutput.t108 gnd 0.060183f
C1548 CSoutput.t155 gnd 0.060183f
C1549 CSoutput.n86 gnd 0.465123f
C1550 CSoutput.n87 gnd 0.232631f
C1551 CSoutput.t81 gnd 0.060183f
C1552 CSoutput.t131 gnd 0.060183f
C1553 CSoutput.n88 gnd 0.465123f
C1554 CSoutput.n89 gnd 0.232631f
C1555 CSoutput.t99 gnd 0.060183f
C1556 CSoutput.t147 gnd 0.060183f
C1557 CSoutput.n90 gnd 0.465123f
C1558 CSoutput.n91 gnd 0.232631f
C1559 CSoutput.t116 gnd 0.060183f
C1560 CSoutput.t165 gnd 0.060183f
C1561 CSoutput.n92 gnd 0.465123f
C1562 CSoutput.n93 gnd 0.232631f
C1563 CSoutput.t94 gnd 0.060183f
C1564 CSoutput.t139 gnd 0.060183f
C1565 CSoutput.n94 gnd 0.465123f
C1566 CSoutput.n95 gnd 0.232631f
C1567 CSoutput.t135 gnd 0.060183f
C1568 CSoutput.t156 gnd 0.060183f
C1569 CSoutput.n96 gnd 0.465123f
C1570 CSoutput.n97 gnd 0.426591f
C1571 CSoutput.t109 gnd 0.060183f
C1572 CSoutput.t75 gnd 0.060183f
C1573 CSoutput.n98 gnd 0.465954f
C1574 CSoutput.t54 gnd 0.060183f
C1575 CSoutput.t111 gnd 0.060183f
C1576 CSoutput.n99 gnd 0.465123f
C1577 CSoutput.n100 gnd 0.472099f
C1578 CSoutput.t105 gnd 0.060183f
C1579 CSoutput.t72 gnd 0.060183f
C1580 CSoutput.n101 gnd 0.465123f
C1581 CSoutput.n102 gnd 0.232631f
C1582 CSoutput.t53 gnd 0.060183f
C1583 CSoutput.t51 gnd 0.060183f
C1584 CSoutput.n103 gnd 0.465123f
C1585 CSoutput.n104 gnd 0.232631f
C1586 CSoutput.t127 gnd 0.060183f
C1587 CSoutput.t87 gnd 0.060183f
C1588 CSoutput.n105 gnd 0.465123f
C1589 CSoutput.n106 gnd 0.232631f
C1590 CSoutput.t83 gnd 0.060183f
C1591 CSoutput.t49 gnd 0.060183f
C1592 CSoutput.n107 gnd 0.465123f
C1593 CSoutput.n108 gnd 0.232631f
C1594 CSoutput.t152 gnd 0.060183f
C1595 CSoutput.t124 gnd 0.060183f
C1596 CSoutput.n109 gnd 0.465123f
C1597 CSoutput.n110 gnd 0.232631f
C1598 CSoutput.t110 gnd 0.060183f
C1599 CSoutput.t76 gnd 0.060183f
C1600 CSoutput.n111 gnd 0.465123f
C1601 CSoutput.n112 gnd 0.232631f
C1602 CSoutput.t68 gnd 0.060183f
C1603 CSoutput.t148 gnd 0.060183f
C1604 CSoutput.n113 gnd 0.465123f
C1605 CSoutput.n114 gnd 0.232631f
C1606 CSoutput.t106 gnd 0.060183f
C1607 CSoutput.t104 gnd 0.060183f
C1608 CSoutput.n115 gnd 0.465123f
C1609 CSoutput.n116 gnd 0.346911f
C1610 CSoutput.n117 gnd 0.437452f
C1611 CSoutput.t121 gnd 0.060183f
C1612 CSoutput.t89 gnd 0.060183f
C1613 CSoutput.n118 gnd 0.465954f
C1614 CSoutput.t66 gnd 0.060183f
C1615 CSoutput.t122 gnd 0.060183f
C1616 CSoutput.n119 gnd 0.465123f
C1617 CSoutput.n120 gnd 0.472099f
C1618 CSoutput.t118 gnd 0.060183f
C1619 CSoutput.t86 gnd 0.060183f
C1620 CSoutput.n121 gnd 0.465123f
C1621 CSoutput.n122 gnd 0.232631f
C1622 CSoutput.t65 gnd 0.060183f
C1623 CSoutput.t64 gnd 0.060183f
C1624 CSoutput.n123 gnd 0.465123f
C1625 CSoutput.n124 gnd 0.232631f
C1626 CSoutput.t136 gnd 0.060183f
C1627 CSoutput.t100 gnd 0.060183f
C1628 CSoutput.n125 gnd 0.465123f
C1629 CSoutput.n126 gnd 0.232631f
C1630 CSoutput.t96 gnd 0.060183f
C1631 CSoutput.t61 gnd 0.060183f
C1632 CSoutput.n127 gnd 0.465123f
C1633 CSoutput.n128 gnd 0.232631f
C1634 CSoutput.t166 gnd 0.060183f
C1635 CSoutput.t134 gnd 0.060183f
C1636 CSoutput.n129 gnd 0.465123f
C1637 CSoutput.n130 gnd 0.232631f
C1638 CSoutput.t120 gnd 0.060183f
C1639 CSoutput.t88 gnd 0.060183f
C1640 CSoutput.n131 gnd 0.465123f
C1641 CSoutput.n132 gnd 0.232631f
C1642 CSoutput.t85 gnd 0.060183f
C1643 CSoutput.t160 gnd 0.060183f
C1644 CSoutput.n133 gnd 0.465123f
C1645 CSoutput.n134 gnd 0.232631f
C1646 CSoutput.t119 gnd 0.060183f
C1647 CSoutput.t117 gnd 0.060183f
C1648 CSoutput.n135 gnd 0.465123f
C1649 CSoutput.n136 gnd 0.346911f
C1650 CSoutput.n137 gnd 0.48896f
C1651 CSoutput.n138 gnd 10.4068f
C1652 CSoutput.n140 gnd 0.853499f
C1653 CSoutput.n141 gnd 0.640125f
C1654 CSoutput.n142 gnd 0.853499f
C1655 CSoutput.n143 gnd 0.853499f
C1656 CSoutput.n144 gnd 2.29788f
C1657 CSoutput.n145 gnd 0.853499f
C1658 CSoutput.n146 gnd 0.853499f
C1659 CSoutput.t211 gnd 1.06687f
C1660 CSoutput.n147 gnd 0.853499f
C1661 CSoutput.n148 gnd 0.853499f
C1662 CSoutput.n152 gnd 0.853499f
C1663 CSoutput.n156 gnd 0.853499f
C1664 CSoutput.n157 gnd 0.853499f
C1665 CSoutput.n159 gnd 0.853499f
C1666 CSoutput.n164 gnd 0.853499f
C1667 CSoutput.n166 gnd 0.853499f
C1668 CSoutput.n167 gnd 0.853499f
C1669 CSoutput.n169 gnd 0.853499f
C1670 CSoutput.n170 gnd 0.853499f
C1671 CSoutput.n172 gnd 0.853499f
C1672 CSoutput.t205 gnd 14.2619f
C1673 CSoutput.n174 gnd 0.853499f
C1674 CSoutput.n175 gnd 0.640125f
C1675 CSoutput.n176 gnd 0.853499f
C1676 CSoutput.n177 gnd 0.853499f
C1677 CSoutput.n178 gnd 2.29788f
C1678 CSoutput.n179 gnd 0.853499f
C1679 CSoutput.n180 gnd 0.853499f
C1680 CSoutput.t208 gnd 1.06687f
C1681 CSoutput.n181 gnd 0.853499f
C1682 CSoutput.n182 gnd 0.853499f
C1683 CSoutput.n186 gnd 0.853499f
C1684 CSoutput.n190 gnd 0.853499f
C1685 CSoutput.n191 gnd 0.853499f
C1686 CSoutput.n193 gnd 0.853499f
C1687 CSoutput.n198 gnd 0.853499f
C1688 CSoutput.n200 gnd 0.853499f
C1689 CSoutput.n201 gnd 0.853499f
C1690 CSoutput.n203 gnd 0.853499f
C1691 CSoutput.n204 gnd 0.853499f
C1692 CSoutput.n206 gnd 0.853499f
C1693 CSoutput.n207 gnd 0.640125f
C1694 CSoutput.n209 gnd 0.853499f
C1695 CSoutput.n210 gnd 0.640125f
C1696 CSoutput.n211 gnd 0.853499f
C1697 CSoutput.n212 gnd 0.853499f
C1698 CSoutput.n213 gnd 2.29788f
C1699 CSoutput.n214 gnd 0.853499f
C1700 CSoutput.n215 gnd 0.853499f
C1701 CSoutput.t210 gnd 1.06687f
C1702 CSoutput.n216 gnd 0.853499f
C1703 CSoutput.n217 gnd 2.29788f
C1704 CSoutput.n219 gnd 0.853499f
C1705 CSoutput.n220 gnd 0.853499f
C1706 CSoutput.n222 gnd 0.853499f
C1707 CSoutput.n223 gnd 0.853499f
C1708 CSoutput.t216 gnd 14.0295f
C1709 CSoutput.t214 gnd 14.2619f
C1710 CSoutput.n229 gnd 2.67755f
C1711 CSoutput.n230 gnd 10.907401f
C1712 CSoutput.n231 gnd 11.3638f
C1713 CSoutput.n236 gnd 2.90051f
C1714 CSoutput.n242 gnd 0.853499f
C1715 CSoutput.n244 gnd 0.853499f
C1716 CSoutput.n246 gnd 0.853499f
C1717 CSoutput.n248 gnd 0.853499f
C1718 CSoutput.n250 gnd 0.853499f
C1719 CSoutput.n256 gnd 0.853499f
C1720 CSoutput.n263 gnd 1.56584f
C1721 CSoutput.n264 gnd 1.56584f
C1722 CSoutput.n265 gnd 0.853499f
C1723 CSoutput.n266 gnd 0.853499f
C1724 CSoutput.n268 gnd 0.640125f
C1725 CSoutput.n269 gnd 0.548209f
C1726 CSoutput.n271 gnd 0.640125f
C1727 CSoutput.n272 gnd 0.548209f
C1728 CSoutput.n273 gnd 0.640125f
C1729 CSoutput.n275 gnd 0.853499f
C1730 CSoutput.n277 gnd 2.29788f
C1731 CSoutput.n278 gnd 2.67755f
C1732 CSoutput.n279 gnd 10.032f
C1733 CSoutput.n281 gnd 0.640125f
C1734 CSoutput.n282 gnd 1.64708f
C1735 CSoutput.n283 gnd 0.640125f
C1736 CSoutput.n285 gnd 0.853499f
C1737 CSoutput.n287 gnd 2.29788f
C1738 CSoutput.n288 gnd 5.00516f
C1739 CSoutput.t102 gnd 0.060183f
C1740 CSoutput.t80 gnd 0.060183f
C1741 CSoutput.n289 gnd 0.465954f
C1742 CSoutput.t144 gnd 0.060183f
C1743 CSoutput.t62 gnd 0.060183f
C1744 CSoutput.n290 gnd 0.465123f
C1745 CSoutput.n291 gnd 0.472099f
C1746 CSoutput.t125 gnd 0.060183f
C1747 CSoutput.t69 gnd 0.060183f
C1748 CSoutput.n292 gnd 0.465123f
C1749 CSoutput.n293 gnd 0.232631f
C1750 CSoutput.t138 gnd 0.060183f
C1751 CSoutput.t90 gnd 0.060183f
C1752 CSoutput.n294 gnd 0.465123f
C1753 CSoutput.n295 gnd 0.232631f
C1754 CSoutput.t153 gnd 0.060183f
C1755 CSoutput.t107 gnd 0.060183f
C1756 CSoutput.n296 gnd 0.465123f
C1757 CSoutput.n297 gnd 0.232631f
C1758 CSoutput.t130 gnd 0.060183f
C1759 CSoutput.t82 gnd 0.060183f
C1760 CSoutput.n298 gnd 0.465123f
C1761 CSoutput.n299 gnd 0.232631f
C1762 CSoutput.t146 gnd 0.060183f
C1763 CSoutput.t98 gnd 0.060183f
C1764 CSoutput.n300 gnd 0.465123f
C1765 CSoutput.n301 gnd 0.232631f
C1766 CSoutput.t164 gnd 0.060183f
C1767 CSoutput.t114 gnd 0.060183f
C1768 CSoutput.n302 gnd 0.465123f
C1769 CSoutput.n303 gnd 0.232631f
C1770 CSoutput.t50 gnd 0.060183f
C1771 CSoutput.t91 gnd 0.060183f
C1772 CSoutput.n304 gnd 0.465123f
C1773 CSoutput.n305 gnd 0.232631f
C1774 CSoutput.t154 gnd 0.060183f
C1775 CSoutput.t133 gnd 0.060183f
C1776 CSoutput.n306 gnd 0.465123f
C1777 CSoutput.n307 gnd 0.426591f
C1778 CSoutput.t150 gnd 0.060183f
C1779 CSoutput.t151 gnd 0.060183f
C1780 CSoutput.n308 gnd 0.465954f
C1781 CSoutput.t60 gnd 0.060183f
C1782 CSoutput.t132 gnd 0.060183f
C1783 CSoutput.n309 gnd 0.465123f
C1784 CSoutput.n310 gnd 0.472099f
C1785 CSoutput.t143 gnd 0.060183f
C1786 CSoutput.t57 gnd 0.060183f
C1787 CSoutput.n311 gnd 0.465123f
C1788 CSoutput.n312 gnd 0.232631f
C1789 CSoutput.t101 gnd 0.060183f
C1790 CSoutput.t129 gnd 0.060183f
C1791 CSoutput.n313 gnd 0.465123f
C1792 CSoutput.n314 gnd 0.232631f
C1793 CSoutput.t159 gnd 0.060183f
C1794 CSoutput.t84 gnd 0.060183f
C1795 CSoutput.n315 gnd 0.465123f
C1796 CSoutput.n316 gnd 0.232631f
C1797 CSoutput.t128 gnd 0.060183f
C1798 CSoutput.t167 gnd 0.060183f
C1799 CSoutput.n317 gnd 0.465123f
C1800 CSoutput.n318 gnd 0.232631f
C1801 CSoutput.t79 gnd 0.060183f
C1802 CSoutput.t113 gnd 0.060183f
C1803 CSoutput.n319 gnd 0.465123f
C1804 CSoutput.n320 gnd 0.232631f
C1805 CSoutput.t149 gnd 0.060183f
C1806 CSoutput.t59 gnd 0.060183f
C1807 CSoutput.n321 gnd 0.465123f
C1808 CSoutput.n322 gnd 0.232631f
C1809 CSoutput.t78 gnd 0.060183f
C1810 CSoutput.t142 gnd 0.060183f
C1811 CSoutput.n323 gnd 0.465123f
C1812 CSoutput.n324 gnd 0.232631f
C1813 CSoutput.t55 gnd 0.060183f
C1814 CSoutput.t56 gnd 0.060183f
C1815 CSoutput.n325 gnd 0.465123f
C1816 CSoutput.n326 gnd 0.346911f
C1817 CSoutput.n327 gnd 0.437452f
C1818 CSoutput.t161 gnd 0.060183f
C1819 CSoutput.t163 gnd 0.060183f
C1820 CSoutput.n328 gnd 0.465954f
C1821 CSoutput.t77 gnd 0.060183f
C1822 CSoutput.t141 gnd 0.060183f
C1823 CSoutput.n329 gnd 0.465123f
C1824 CSoutput.n330 gnd 0.472099f
C1825 CSoutput.t158 gnd 0.060183f
C1826 CSoutput.t70 gnd 0.060183f
C1827 CSoutput.n331 gnd 0.465123f
C1828 CSoutput.n332 gnd 0.232631f
C1829 CSoutput.t115 gnd 0.060183f
C1830 CSoutput.t140 gnd 0.060183f
C1831 CSoutput.n333 gnd 0.465123f
C1832 CSoutput.n334 gnd 0.232631f
C1833 CSoutput.t52 gnd 0.060183f
C1834 CSoutput.t97 gnd 0.060183f
C1835 CSoutput.n335 gnd 0.465123f
C1836 CSoutput.n336 gnd 0.232631f
C1837 CSoutput.t137 gnd 0.060183f
C1838 CSoutput.t58 gnd 0.060183f
C1839 CSoutput.n337 gnd 0.465123f
C1840 CSoutput.n338 gnd 0.232631f
C1841 CSoutput.t95 gnd 0.060183f
C1842 CSoutput.t123 gnd 0.060183f
C1843 CSoutput.n339 gnd 0.465123f
C1844 CSoutput.n340 gnd 0.232631f
C1845 CSoutput.t162 gnd 0.060183f
C1846 CSoutput.t74 gnd 0.060183f
C1847 CSoutput.n341 gnd 0.465123f
C1848 CSoutput.n342 gnd 0.232631f
C1849 CSoutput.t93 gnd 0.060183f
C1850 CSoutput.t157 gnd 0.060183f
C1851 CSoutput.n343 gnd 0.465123f
C1852 CSoutput.n344 gnd 0.232631f
C1853 CSoutput.t67 gnd 0.060183f
C1854 CSoutput.t71 gnd 0.060183f
C1855 CSoutput.n345 gnd 0.465122f
C1856 CSoutput.n346 gnd 0.346913f
C1857 CSoutput.n347 gnd 0.48896f
C1858 CSoutput.n348 gnd 14.284201f
C1859 CSoutput.t185 gnd 0.05266f
C1860 CSoutput.t199 gnd 0.05266f
C1861 CSoutput.n349 gnd 0.466878f
C1862 CSoutput.t0 gnd 0.05266f
C1863 CSoutput.t193 gnd 0.05266f
C1864 CSoutput.n350 gnd 0.465321f
C1865 CSoutput.n351 gnd 0.433592f
C1866 CSoutput.t10 gnd 0.05266f
C1867 CSoutput.t7 gnd 0.05266f
C1868 CSoutput.n352 gnd 0.465321f
C1869 CSoutput.n353 gnd 0.21374f
C1870 CSoutput.t35 gnd 0.05266f
C1871 CSoutput.t173 gnd 0.05266f
C1872 CSoutput.n354 gnd 0.465321f
C1873 CSoutput.n355 gnd 0.21374f
C1874 CSoutput.t195 gnd 0.05266f
C1875 CSoutput.t198 gnd 0.05266f
C1876 CSoutput.n356 gnd 0.465321f
C1877 CSoutput.n357 gnd 0.21374f
C1878 CSoutput.t24 gnd 0.05266f
C1879 CSoutput.t16 gnd 0.05266f
C1880 CSoutput.n358 gnd 0.465321f
C1881 CSoutput.n359 gnd 0.21374f
C1882 CSoutput.t17 gnd 0.05266f
C1883 CSoutput.t30 gnd 0.05266f
C1884 CSoutput.n360 gnd 0.465321f
C1885 CSoutput.n361 gnd 0.21374f
C1886 CSoutput.t186 gnd 0.05266f
C1887 CSoutput.t191 gnd 0.05266f
C1888 CSoutput.n362 gnd 0.465321f
C1889 CSoutput.n363 gnd 0.21374f
C1890 CSoutput.t14 gnd 0.05266f
C1891 CSoutput.t3 gnd 0.05266f
C1892 CSoutput.n364 gnd 0.465321f
C1893 CSoutput.n365 gnd 0.21374f
C1894 CSoutput.t36 gnd 0.05266f
C1895 CSoutput.t46 gnd 0.05266f
C1896 CSoutput.n366 gnd 0.465321f
C1897 CSoutput.n367 gnd 0.39418f
C1898 CSoutput.t33 gnd 0.05266f
C1899 CSoutput.t183 gnd 0.05266f
C1900 CSoutput.n368 gnd 0.466878f
C1901 CSoutput.t170 gnd 0.05266f
C1902 CSoutput.t175 gnd 0.05266f
C1903 CSoutput.n369 gnd 0.465321f
C1904 CSoutput.n370 gnd 0.433592f
C1905 CSoutput.t189 gnd 0.05266f
C1906 CSoutput.t9 gnd 0.05266f
C1907 CSoutput.n371 gnd 0.465321f
C1908 CSoutput.n372 gnd 0.21374f
C1909 CSoutput.t171 gnd 0.05266f
C1910 CSoutput.t197 gnd 0.05266f
C1911 CSoutput.n373 gnd 0.465321f
C1912 CSoutput.n374 gnd 0.21374f
C1913 CSoutput.t182 gnd 0.05266f
C1914 CSoutput.t44 gnd 0.05266f
C1915 CSoutput.n375 gnd 0.465321f
C1916 CSoutput.n376 gnd 0.21374f
C1917 CSoutput.t20 gnd 0.05266f
C1918 CSoutput.t188 gnd 0.05266f
C1919 CSoutput.n377 gnd 0.465321f
C1920 CSoutput.n378 gnd 0.21374f
C1921 CSoutput.t31 gnd 0.05266f
C1922 CSoutput.t18 gnd 0.05266f
C1923 CSoutput.n379 gnd 0.465321f
C1924 CSoutput.n380 gnd 0.21374f
C1925 CSoutput.t174 gnd 0.05266f
C1926 CSoutput.t176 gnd 0.05266f
C1927 CSoutput.n381 gnd 0.465321f
C1928 CSoutput.n382 gnd 0.21374f
C1929 CSoutput.t180 gnd 0.05266f
C1930 CSoutput.t47 gnd 0.05266f
C1931 CSoutput.n383 gnd 0.465321f
C1932 CSoutput.n384 gnd 0.21374f
C1933 CSoutput.t172 gnd 0.05266f
C1934 CSoutput.t34 gnd 0.05266f
C1935 CSoutput.n385 gnd 0.465321f
C1936 CSoutput.n386 gnd 0.324504f
C1937 CSoutput.n387 gnd 0.602953f
C1938 CSoutput.n388 gnd 14.712999f
C1939 CSoutput.t28 gnd 0.05266f
C1940 CSoutput.t8 gnd 0.05266f
C1941 CSoutput.n389 gnd 0.466878f
C1942 CSoutput.t48 gnd 0.05266f
C1943 CSoutput.t4 gnd 0.05266f
C1944 CSoutput.n390 gnd 0.465321f
C1945 CSoutput.n391 gnd 0.433592f
C1946 CSoutput.t41 gnd 0.05266f
C1947 CSoutput.t6 gnd 0.05266f
C1948 CSoutput.n392 gnd 0.465321f
C1949 CSoutput.n393 gnd 0.21374f
C1950 CSoutput.t187 gnd 0.05266f
C1951 CSoutput.t25 gnd 0.05266f
C1952 CSoutput.n394 gnd 0.465321f
C1953 CSoutput.n395 gnd 0.21374f
C1954 CSoutput.t5 gnd 0.05266f
C1955 CSoutput.t169 gnd 0.05266f
C1956 CSoutput.n396 gnd 0.465321f
C1957 CSoutput.n397 gnd 0.21374f
C1958 CSoutput.t13 gnd 0.05266f
C1959 CSoutput.t196 gnd 0.05266f
C1960 CSoutput.n398 gnd 0.465321f
C1961 CSoutput.n399 gnd 0.21374f
C1962 CSoutput.t26 gnd 0.05266f
C1963 CSoutput.t2 gnd 0.05266f
C1964 CSoutput.n400 gnd 0.465321f
C1965 CSoutput.n401 gnd 0.21374f
C1966 CSoutput.t184 gnd 0.05266f
C1967 CSoutput.t192 gnd 0.05266f
C1968 CSoutput.n402 gnd 0.465321f
C1969 CSoutput.n403 gnd 0.21374f
C1970 CSoutput.t19 gnd 0.05266f
C1971 CSoutput.t178 gnd 0.05266f
C1972 CSoutput.n404 gnd 0.465321f
C1973 CSoutput.n405 gnd 0.21374f
C1974 CSoutput.t12 gnd 0.05266f
C1975 CSoutput.t32 gnd 0.05266f
C1976 CSoutput.n406 gnd 0.465321f
C1977 CSoutput.n407 gnd 0.39418f
C1978 CSoutput.t23 gnd 0.05266f
C1979 CSoutput.t11 gnd 0.05266f
C1980 CSoutput.n408 gnd 0.466878f
C1981 CSoutput.t181 gnd 0.05266f
C1982 CSoutput.t27 gnd 0.05266f
C1983 CSoutput.n409 gnd 0.465321f
C1984 CSoutput.n410 gnd 0.433592f
C1985 CSoutput.t1 gnd 0.05266f
C1986 CSoutput.t179 gnd 0.05266f
C1987 CSoutput.n411 gnd 0.465321f
C1988 CSoutput.n412 gnd 0.21374f
C1989 CSoutput.t38 gnd 0.05266f
C1990 CSoutput.t42 gnd 0.05266f
C1991 CSoutput.n413 gnd 0.465321f
C1992 CSoutput.n414 gnd 0.21374f
C1993 CSoutput.t21 gnd 0.05266f
C1994 CSoutput.t29 gnd 0.05266f
C1995 CSoutput.n415 gnd 0.465321f
C1996 CSoutput.n416 gnd 0.21374f
C1997 CSoutput.t43 gnd 0.05266f
C1998 CSoutput.t194 gnd 0.05266f
C1999 CSoutput.n417 gnd 0.465321f
C2000 CSoutput.n418 gnd 0.21374f
C2001 CSoutput.t22 gnd 0.05266f
C2002 CSoutput.t15 gnd 0.05266f
C2003 CSoutput.n419 gnd 0.465321f
C2004 CSoutput.n420 gnd 0.21374f
C2005 CSoutput.t37 gnd 0.05266f
C2006 CSoutput.t40 gnd 0.05266f
C2007 CSoutput.n421 gnd 0.465321f
C2008 CSoutput.n422 gnd 0.21374f
C2009 CSoutput.t177 gnd 0.05266f
C2010 CSoutput.t45 gnd 0.05266f
C2011 CSoutput.n423 gnd 0.465321f
C2012 CSoutput.n424 gnd 0.21374f
C2013 CSoutput.t190 gnd 0.05266f
C2014 CSoutput.t39 gnd 0.05266f
C2015 CSoutput.n425 gnd 0.465321f
C2016 CSoutput.n426 gnd 0.324504f
C2017 CSoutput.n427 gnd 0.602953f
C2018 CSoutput.n428 gnd 9.11085f
C2019 CSoutput.n429 gnd 15.505301f
C2020 vdd.t292 gnd 0.036842f
C2021 vdd.t274 gnd 0.036842f
C2022 vdd.n0 gnd 0.290576f
C2023 vdd.t251 gnd 0.036842f
C2024 vdd.t288 gnd 0.036842f
C2025 vdd.n1 gnd 0.290096f
C2026 vdd.n2 gnd 0.267524f
C2027 vdd.t269 gnd 0.036842f
C2028 vdd.t299 gnd 0.036842f
C2029 vdd.n3 gnd 0.290096f
C2030 vdd.n4 gnd 0.135297f
C2031 vdd.t297 gnd 0.036842f
C2032 vdd.t279 gnd 0.036842f
C2033 vdd.n5 gnd 0.290096f
C2034 vdd.n6 gnd 0.126951f
C2035 vdd.t303 gnd 0.036842f
C2036 vdd.t267 gnd 0.036842f
C2037 vdd.n7 gnd 0.290576f
C2038 vdd.t277 gnd 0.036842f
C2039 vdd.t295 gnd 0.036842f
C2040 vdd.n8 gnd 0.290096f
C2041 vdd.n9 gnd 0.267524f
C2042 vdd.t284 gnd 0.036842f
C2043 vdd.t255 gnd 0.036842f
C2044 vdd.n10 gnd 0.290096f
C2045 vdd.n11 gnd 0.135297f
C2046 vdd.t264 gnd 0.036842f
C2047 vdd.t271 gnd 0.036842f
C2048 vdd.n12 gnd 0.290096f
C2049 vdd.n13 gnd 0.126951f
C2050 vdd.n14 gnd 0.089752f
C2051 vdd.t304 gnd 0.020468f
C2052 vdd.t1 gnd 0.020468f
C2053 vdd.n15 gnd 0.188395f
C2054 vdd.t87 gnd 0.020468f
C2055 vdd.t84 gnd 0.020468f
C2056 vdd.n16 gnd 0.187844f
C2057 vdd.n17 gnd 0.326907f
C2058 vdd.t307 gnd 0.020468f
C2059 vdd.t6 gnd 0.020468f
C2060 vdd.n18 gnd 0.187844f
C2061 vdd.n19 gnd 0.135246f
C2062 vdd.t5 gnd 0.020468f
C2063 vdd.t2 gnd 0.020468f
C2064 vdd.n20 gnd 0.188395f
C2065 vdd.t305 gnd 0.020468f
C2066 vdd.t85 gnd 0.020468f
C2067 vdd.n21 gnd 0.187844f
C2068 vdd.n22 gnd 0.326907f
C2069 vdd.t3 gnd 0.020468f
C2070 vdd.t4 gnd 0.020468f
C2071 vdd.n23 gnd 0.187844f
C2072 vdd.n24 gnd 0.135246f
C2073 vdd.t86 gnd 0.020468f
C2074 vdd.t7 gnd 0.020468f
C2075 vdd.n25 gnd 0.187844f
C2076 vdd.t0 gnd 0.020468f
C2077 vdd.t306 gnd 0.020468f
C2078 vdd.n26 gnd 0.187844f
C2079 vdd.n27 gnd 22.0613f
C2080 vdd.n28 gnd 8.74629f
C2081 vdd.n29 gnd 0.005582f
C2082 vdd.n30 gnd 0.00518f
C2083 vdd.n31 gnd 0.002865f
C2084 vdd.n32 gnd 0.006579f
C2085 vdd.n33 gnd 0.002784f
C2086 vdd.n34 gnd 0.002947f
C2087 vdd.n35 gnd 0.00518f
C2088 vdd.n36 gnd 0.002784f
C2089 vdd.n37 gnd 0.006579f
C2090 vdd.n38 gnd 0.002947f
C2091 vdd.n39 gnd 0.00518f
C2092 vdd.n40 gnd 0.002784f
C2093 vdd.n41 gnd 0.004935f
C2094 vdd.n42 gnd 0.004949f
C2095 vdd.t170 gnd 0.014135f
C2096 vdd.n43 gnd 0.031451f
C2097 vdd.n44 gnd 0.163677f
C2098 vdd.n45 gnd 0.002784f
C2099 vdd.n46 gnd 0.002947f
C2100 vdd.n47 gnd 0.006579f
C2101 vdd.n48 gnd 0.006579f
C2102 vdd.n49 gnd 0.002947f
C2103 vdd.n50 gnd 0.002784f
C2104 vdd.n51 gnd 0.00518f
C2105 vdd.n52 gnd 0.00518f
C2106 vdd.n53 gnd 0.002784f
C2107 vdd.n54 gnd 0.002947f
C2108 vdd.n55 gnd 0.006579f
C2109 vdd.n56 gnd 0.006579f
C2110 vdd.n57 gnd 0.002947f
C2111 vdd.n58 gnd 0.002784f
C2112 vdd.n59 gnd 0.00518f
C2113 vdd.n60 gnd 0.00518f
C2114 vdd.n61 gnd 0.002784f
C2115 vdd.n62 gnd 0.002947f
C2116 vdd.n63 gnd 0.006579f
C2117 vdd.n64 gnd 0.006579f
C2118 vdd.n65 gnd 0.015555f
C2119 vdd.n66 gnd 0.002865f
C2120 vdd.n67 gnd 0.002784f
C2121 vdd.n68 gnd 0.013389f
C2122 vdd.n69 gnd 0.009347f
C2123 vdd.t141 gnd 0.032748f
C2124 vdd.t222 gnd 0.032748f
C2125 vdd.n70 gnd 0.225067f
C2126 vdd.n71 gnd 0.176981f
C2127 vdd.t114 gnd 0.032748f
C2128 vdd.t201 gnd 0.032748f
C2129 vdd.n72 gnd 0.225067f
C2130 vdd.n73 gnd 0.142823f
C2131 vdd.t122 gnd 0.032748f
C2132 vdd.t216 gnd 0.032748f
C2133 vdd.n74 gnd 0.225067f
C2134 vdd.n75 gnd 0.142823f
C2135 vdd.t153 gnd 0.032748f
C2136 vdd.t232 gnd 0.032748f
C2137 vdd.n76 gnd 0.225067f
C2138 vdd.n77 gnd 0.142823f
C2139 vdd.t177 gnd 0.032748f
C2140 vdd.t207 gnd 0.032748f
C2141 vdd.n78 gnd 0.225067f
C2142 vdd.n79 gnd 0.142823f
C2143 vdd.t142 gnd 0.032748f
C2144 vdd.t224 gnd 0.032748f
C2145 vdd.n80 gnd 0.225067f
C2146 vdd.n81 gnd 0.142823f
C2147 vdd.t163 gnd 0.032748f
C2148 vdd.t243 gnd 0.032748f
C2149 vdd.n82 gnd 0.225067f
C2150 vdd.n83 gnd 0.142823f
C2151 vdd.t189 gnd 0.032748f
C2152 vdd.t91 gnd 0.032748f
C2153 vdd.n84 gnd 0.225067f
C2154 vdd.n85 gnd 0.142823f
C2155 vdd.t155 gnd 0.032748f
C2156 vdd.t233 gnd 0.032748f
C2157 vdd.n86 gnd 0.225067f
C2158 vdd.n87 gnd 0.142823f
C2159 vdd.n88 gnd 0.005582f
C2160 vdd.n89 gnd 0.00518f
C2161 vdd.n90 gnd 0.002865f
C2162 vdd.n91 gnd 0.006579f
C2163 vdd.n92 gnd 0.002784f
C2164 vdd.n93 gnd 0.002947f
C2165 vdd.n94 gnd 0.00518f
C2166 vdd.n95 gnd 0.002784f
C2167 vdd.n96 gnd 0.006579f
C2168 vdd.n97 gnd 0.002947f
C2169 vdd.n98 gnd 0.00518f
C2170 vdd.n99 gnd 0.002784f
C2171 vdd.n100 gnd 0.004935f
C2172 vdd.n101 gnd 0.004949f
C2173 vdd.t210 gnd 0.014135f
C2174 vdd.n102 gnd 0.031451f
C2175 vdd.n103 gnd 0.163677f
C2176 vdd.n104 gnd 0.002784f
C2177 vdd.n105 gnd 0.002947f
C2178 vdd.n106 gnd 0.006579f
C2179 vdd.n107 gnd 0.006579f
C2180 vdd.n108 gnd 0.002947f
C2181 vdd.n109 gnd 0.002784f
C2182 vdd.n110 gnd 0.00518f
C2183 vdd.n111 gnd 0.00518f
C2184 vdd.n112 gnd 0.002784f
C2185 vdd.n113 gnd 0.002947f
C2186 vdd.n114 gnd 0.006579f
C2187 vdd.n115 gnd 0.006579f
C2188 vdd.n116 gnd 0.002947f
C2189 vdd.n117 gnd 0.002784f
C2190 vdd.n118 gnd 0.00518f
C2191 vdd.n119 gnd 0.00518f
C2192 vdd.n120 gnd 0.002784f
C2193 vdd.n121 gnd 0.002947f
C2194 vdd.n122 gnd 0.006579f
C2195 vdd.n123 gnd 0.006579f
C2196 vdd.n124 gnd 0.015555f
C2197 vdd.n125 gnd 0.002865f
C2198 vdd.n126 gnd 0.002784f
C2199 vdd.n127 gnd 0.013389f
C2200 vdd.n128 gnd 0.009054f
C2201 vdd.n129 gnd 0.106261f
C2202 vdd.n130 gnd 0.005582f
C2203 vdd.n131 gnd 0.00518f
C2204 vdd.n132 gnd 0.002865f
C2205 vdd.n133 gnd 0.006579f
C2206 vdd.n134 gnd 0.002784f
C2207 vdd.n135 gnd 0.002947f
C2208 vdd.n136 gnd 0.00518f
C2209 vdd.n137 gnd 0.002784f
C2210 vdd.n138 gnd 0.006579f
C2211 vdd.n139 gnd 0.002947f
C2212 vdd.n140 gnd 0.00518f
C2213 vdd.n141 gnd 0.002784f
C2214 vdd.n142 gnd 0.004935f
C2215 vdd.n143 gnd 0.004949f
C2216 vdd.t229 gnd 0.014135f
C2217 vdd.n144 gnd 0.031451f
C2218 vdd.n145 gnd 0.163677f
C2219 vdd.n146 gnd 0.002784f
C2220 vdd.n147 gnd 0.002947f
C2221 vdd.n148 gnd 0.006579f
C2222 vdd.n149 gnd 0.006579f
C2223 vdd.n150 gnd 0.002947f
C2224 vdd.n151 gnd 0.002784f
C2225 vdd.n152 gnd 0.00518f
C2226 vdd.n153 gnd 0.00518f
C2227 vdd.n154 gnd 0.002784f
C2228 vdd.n155 gnd 0.002947f
C2229 vdd.n156 gnd 0.006579f
C2230 vdd.n157 gnd 0.006579f
C2231 vdd.n158 gnd 0.002947f
C2232 vdd.n159 gnd 0.002784f
C2233 vdd.n160 gnd 0.00518f
C2234 vdd.n161 gnd 0.00518f
C2235 vdd.n162 gnd 0.002784f
C2236 vdd.n163 gnd 0.002947f
C2237 vdd.n164 gnd 0.006579f
C2238 vdd.n165 gnd 0.006579f
C2239 vdd.n166 gnd 0.015555f
C2240 vdd.n167 gnd 0.002865f
C2241 vdd.n168 gnd 0.002784f
C2242 vdd.n169 gnd 0.013389f
C2243 vdd.n170 gnd 0.009347f
C2244 vdd.t230 gnd 0.032748f
C2245 vdd.t111 gnd 0.032748f
C2246 vdd.n171 gnd 0.225067f
C2247 vdd.n172 gnd 0.176981f
C2248 vdd.t209 gnd 0.032748f
C2249 vdd.t221 gnd 0.032748f
C2250 vdd.n173 gnd 0.225067f
C2251 vdd.n174 gnd 0.142823f
C2252 vdd.t103 gnd 0.032748f
C2253 vdd.t168 gnd 0.032748f
C2254 vdd.n175 gnd 0.225067f
C2255 vdd.n176 gnd 0.142823f
C2256 vdd.t203 gnd 0.032748f
C2257 vdd.t238 gnd 0.032748f
C2258 vdd.n177 gnd 0.225067f
C2259 vdd.n178 gnd 0.142823f
C2260 vdd.t145 gnd 0.032748f
C2261 vdd.t206 gnd 0.032748f
C2262 vdd.n179 gnd 0.225067f
C2263 vdd.n180 gnd 0.142823f
C2264 vdd.t246 gnd 0.032748f
C2265 vdd.t139 gnd 0.032748f
C2266 vdd.n181 gnd 0.225067f
C2267 vdd.n182 gnd 0.142823f
C2268 vdd.t188 gnd 0.032748f
C2269 vdd.t228 gnd 0.032748f
C2270 vdd.n183 gnd 0.225067f
C2271 vdd.n184 gnd 0.142823f
C2272 vdd.t109 gnd 0.032748f
C2273 vdd.t135 gnd 0.032748f
C2274 vdd.n185 gnd 0.225067f
C2275 vdd.n186 gnd 0.142823f
C2276 vdd.t213 gnd 0.032748f
C2277 vdd.t101 gnd 0.032748f
C2278 vdd.n187 gnd 0.225067f
C2279 vdd.n188 gnd 0.142823f
C2280 vdd.n189 gnd 0.005582f
C2281 vdd.n190 gnd 0.00518f
C2282 vdd.n191 gnd 0.002865f
C2283 vdd.n192 gnd 0.006579f
C2284 vdd.n193 gnd 0.002784f
C2285 vdd.n194 gnd 0.002947f
C2286 vdd.n195 gnd 0.00518f
C2287 vdd.n196 gnd 0.002784f
C2288 vdd.n197 gnd 0.006579f
C2289 vdd.n198 gnd 0.002947f
C2290 vdd.n199 gnd 0.00518f
C2291 vdd.n200 gnd 0.002784f
C2292 vdd.n201 gnd 0.004935f
C2293 vdd.n202 gnd 0.004949f
C2294 vdd.t105 gnd 0.014135f
C2295 vdd.n203 gnd 0.031451f
C2296 vdd.n204 gnd 0.163677f
C2297 vdd.n205 gnd 0.002784f
C2298 vdd.n206 gnd 0.002947f
C2299 vdd.n207 gnd 0.006579f
C2300 vdd.n208 gnd 0.006579f
C2301 vdd.n209 gnd 0.002947f
C2302 vdd.n210 gnd 0.002784f
C2303 vdd.n211 gnd 0.00518f
C2304 vdd.n212 gnd 0.00518f
C2305 vdd.n213 gnd 0.002784f
C2306 vdd.n214 gnd 0.002947f
C2307 vdd.n215 gnd 0.006579f
C2308 vdd.n216 gnd 0.006579f
C2309 vdd.n217 gnd 0.002947f
C2310 vdd.n218 gnd 0.002784f
C2311 vdd.n219 gnd 0.00518f
C2312 vdd.n220 gnd 0.00518f
C2313 vdd.n221 gnd 0.002784f
C2314 vdd.n222 gnd 0.002947f
C2315 vdd.n223 gnd 0.006579f
C2316 vdd.n224 gnd 0.006579f
C2317 vdd.n225 gnd 0.015555f
C2318 vdd.n226 gnd 0.002865f
C2319 vdd.n227 gnd 0.002784f
C2320 vdd.n228 gnd 0.013389f
C2321 vdd.n229 gnd 0.009054f
C2322 vdd.n230 gnd 0.063214f
C2323 vdd.n231 gnd 0.227778f
C2324 vdd.n232 gnd 0.005582f
C2325 vdd.n233 gnd 0.00518f
C2326 vdd.n234 gnd 0.002865f
C2327 vdd.n235 gnd 0.006579f
C2328 vdd.n236 gnd 0.002784f
C2329 vdd.n237 gnd 0.002947f
C2330 vdd.n238 gnd 0.00518f
C2331 vdd.n239 gnd 0.002784f
C2332 vdd.n240 gnd 0.006579f
C2333 vdd.n241 gnd 0.002947f
C2334 vdd.n242 gnd 0.00518f
C2335 vdd.n243 gnd 0.002784f
C2336 vdd.n244 gnd 0.004935f
C2337 vdd.n245 gnd 0.004949f
C2338 vdd.t240 gnd 0.014135f
C2339 vdd.n246 gnd 0.031451f
C2340 vdd.n247 gnd 0.163677f
C2341 vdd.n248 gnd 0.002784f
C2342 vdd.n249 gnd 0.002947f
C2343 vdd.n250 gnd 0.006579f
C2344 vdd.n251 gnd 0.006579f
C2345 vdd.n252 gnd 0.002947f
C2346 vdd.n253 gnd 0.002784f
C2347 vdd.n254 gnd 0.00518f
C2348 vdd.n255 gnd 0.00518f
C2349 vdd.n256 gnd 0.002784f
C2350 vdd.n257 gnd 0.002947f
C2351 vdd.n258 gnd 0.006579f
C2352 vdd.n259 gnd 0.006579f
C2353 vdd.n260 gnd 0.002947f
C2354 vdd.n261 gnd 0.002784f
C2355 vdd.n262 gnd 0.00518f
C2356 vdd.n263 gnd 0.00518f
C2357 vdd.n264 gnd 0.002784f
C2358 vdd.n265 gnd 0.002947f
C2359 vdd.n266 gnd 0.006579f
C2360 vdd.n267 gnd 0.006579f
C2361 vdd.n268 gnd 0.015555f
C2362 vdd.n269 gnd 0.002865f
C2363 vdd.n270 gnd 0.002784f
C2364 vdd.n271 gnd 0.013389f
C2365 vdd.n272 gnd 0.009347f
C2366 vdd.t242 gnd 0.032748f
C2367 vdd.t134 gnd 0.032748f
C2368 vdd.n273 gnd 0.225067f
C2369 vdd.n274 gnd 0.176981f
C2370 vdd.t220 gnd 0.032748f
C2371 vdd.t237 gnd 0.032748f
C2372 vdd.n275 gnd 0.225067f
C2373 vdd.n276 gnd 0.142823f
C2374 vdd.t123 gnd 0.032748f
C2375 vdd.t190 gnd 0.032748f
C2376 vdd.n277 gnd 0.225067f
C2377 vdd.n278 gnd 0.142823f
C2378 vdd.t219 gnd 0.032748f
C2379 vdd.t95 gnd 0.032748f
C2380 vdd.n279 gnd 0.225067f
C2381 vdd.n280 gnd 0.142823f
C2382 vdd.t161 gnd 0.032748f
C2383 vdd.t215 gnd 0.032748f
C2384 vdd.n281 gnd 0.225067f
C2385 vdd.n282 gnd 0.142823f
C2386 vdd.t107 gnd 0.032748f
C2387 vdd.t159 gnd 0.032748f
C2388 vdd.n283 gnd 0.225067f
C2389 vdd.n284 gnd 0.142823f
C2390 vdd.t197 gnd 0.032748f
C2391 vdd.t241 gnd 0.032748f
C2392 vdd.n285 gnd 0.225067f
C2393 vdd.n286 gnd 0.142823f
C2394 vdd.t129 gnd 0.032748f
C2395 vdd.t157 gnd 0.032748f
C2396 vdd.n287 gnd 0.225067f
C2397 vdd.n288 gnd 0.142823f
C2398 vdd.t236 gnd 0.032748f
C2399 vdd.t119 gnd 0.032748f
C2400 vdd.n289 gnd 0.225067f
C2401 vdd.n290 gnd 0.142823f
C2402 vdd.n291 gnd 0.005582f
C2403 vdd.n292 gnd 0.00518f
C2404 vdd.n293 gnd 0.002865f
C2405 vdd.n294 gnd 0.006579f
C2406 vdd.n295 gnd 0.002784f
C2407 vdd.n296 gnd 0.002947f
C2408 vdd.n297 gnd 0.00518f
C2409 vdd.n298 gnd 0.002784f
C2410 vdd.n299 gnd 0.006579f
C2411 vdd.n300 gnd 0.002947f
C2412 vdd.n301 gnd 0.00518f
C2413 vdd.n302 gnd 0.002784f
C2414 vdd.n303 gnd 0.004935f
C2415 vdd.n304 gnd 0.004949f
C2416 vdd.t124 gnd 0.014135f
C2417 vdd.n305 gnd 0.031451f
C2418 vdd.n306 gnd 0.163677f
C2419 vdd.n307 gnd 0.002784f
C2420 vdd.n308 gnd 0.002947f
C2421 vdd.n309 gnd 0.006579f
C2422 vdd.n310 gnd 0.006579f
C2423 vdd.n311 gnd 0.002947f
C2424 vdd.n312 gnd 0.002784f
C2425 vdd.n313 gnd 0.00518f
C2426 vdd.n314 gnd 0.00518f
C2427 vdd.n315 gnd 0.002784f
C2428 vdd.n316 gnd 0.002947f
C2429 vdd.n317 gnd 0.006579f
C2430 vdd.n318 gnd 0.006579f
C2431 vdd.n319 gnd 0.002947f
C2432 vdd.n320 gnd 0.002784f
C2433 vdd.n321 gnd 0.00518f
C2434 vdd.n322 gnd 0.00518f
C2435 vdd.n323 gnd 0.002784f
C2436 vdd.n324 gnd 0.002947f
C2437 vdd.n325 gnd 0.006579f
C2438 vdd.n326 gnd 0.006579f
C2439 vdd.n327 gnd 0.015555f
C2440 vdd.n328 gnd 0.002865f
C2441 vdd.n329 gnd 0.002784f
C2442 vdd.n330 gnd 0.013389f
C2443 vdd.n331 gnd 0.009054f
C2444 vdd.n332 gnd 0.063214f
C2445 vdd.n333 gnd 0.260757f
C2446 vdd.n334 gnd 0.007818f
C2447 vdd.n335 gnd 0.010172f
C2448 vdd.n336 gnd 0.008187f
C2449 vdd.n337 gnd 0.008187f
C2450 vdd.n338 gnd 0.010172f
C2451 vdd.n339 gnd 0.010172f
C2452 vdd.n340 gnd 0.743246f
C2453 vdd.n341 gnd 0.010172f
C2454 vdd.n342 gnd 0.010172f
C2455 vdd.n343 gnd 0.010172f
C2456 vdd.n344 gnd 0.805616f
C2457 vdd.n345 gnd 0.010172f
C2458 vdd.n346 gnd 0.010172f
C2459 vdd.n347 gnd 0.010172f
C2460 vdd.n348 gnd 0.010172f
C2461 vdd.n349 gnd 0.008187f
C2462 vdd.n350 gnd 0.010172f
C2463 vdd.t138 gnd 0.519752f
C2464 vdd.n351 gnd 0.010172f
C2465 vdd.n352 gnd 0.010172f
C2466 vdd.n353 gnd 0.010172f
C2467 vdd.t227 gnd 0.519752f
C2468 vdd.n354 gnd 0.010172f
C2469 vdd.n355 gnd 0.010172f
C2470 vdd.n356 gnd 0.010172f
C2471 vdd.n357 gnd 0.010172f
C2472 vdd.n358 gnd 0.010172f
C2473 vdd.n359 gnd 0.008187f
C2474 vdd.n360 gnd 0.010172f
C2475 vdd.n361 gnd 0.58732f
C2476 vdd.n362 gnd 0.010172f
C2477 vdd.n363 gnd 0.010172f
C2478 vdd.n364 gnd 0.010172f
C2479 vdd.t90 gnd 0.519752f
C2480 vdd.n365 gnd 0.010172f
C2481 vdd.n366 gnd 0.010172f
C2482 vdd.n367 gnd 0.010172f
C2483 vdd.n368 gnd 0.010172f
C2484 vdd.n369 gnd 0.010172f
C2485 vdd.n370 gnd 0.008187f
C2486 vdd.n371 gnd 0.010172f
C2487 vdd.t154 gnd 0.519752f
C2488 vdd.n372 gnd 0.010172f
C2489 vdd.n373 gnd 0.010172f
C2490 vdd.n374 gnd 0.010172f
C2491 vdd.n375 gnd 0.60811f
C2492 vdd.n376 gnd 0.010172f
C2493 vdd.n377 gnd 0.010172f
C2494 vdd.n378 gnd 0.010172f
C2495 vdd.n379 gnd 0.010172f
C2496 vdd.n380 gnd 0.010172f
C2497 vdd.n381 gnd 0.008187f
C2498 vdd.n382 gnd 0.010172f
C2499 vdd.t104 gnd 0.519752f
C2500 vdd.n383 gnd 0.010172f
C2501 vdd.n384 gnd 0.010172f
C2502 vdd.n385 gnd 0.010172f
C2503 vdd.n386 gnd 0.52495f
C2504 vdd.n387 gnd 0.010172f
C2505 vdd.n388 gnd 0.010172f
C2506 vdd.n389 gnd 0.010172f
C2507 vdd.n390 gnd 0.010172f
C2508 vdd.n391 gnd 0.024606f
C2509 vdd.n392 gnd 0.025134f
C2510 vdd.t21 gnd 0.519752f
C2511 vdd.n393 gnd 0.024606f
C2512 vdd.n425 gnd 0.010172f
C2513 vdd.t49 gnd 0.125139f
C2514 vdd.t48 gnd 0.133739f
C2515 vdd.t47 gnd 0.16343f
C2516 vdd.n426 gnd 0.209494f
C2517 vdd.n427 gnd 0.176832f
C2518 vdd.n428 gnd 0.013427f
C2519 vdd.n429 gnd 0.010172f
C2520 vdd.n430 gnd 0.008187f
C2521 vdd.n431 gnd 0.010172f
C2522 vdd.n432 gnd 0.008187f
C2523 vdd.n433 gnd 0.010172f
C2524 vdd.n434 gnd 0.008187f
C2525 vdd.n435 gnd 0.010172f
C2526 vdd.n436 gnd 0.008187f
C2527 vdd.n437 gnd 0.010172f
C2528 vdd.n438 gnd 0.008187f
C2529 vdd.n439 gnd 0.010172f
C2530 vdd.t23 gnd 0.125139f
C2531 vdd.t22 gnd 0.133739f
C2532 vdd.t20 gnd 0.16343f
C2533 vdd.n440 gnd 0.209494f
C2534 vdd.n441 gnd 0.176832f
C2535 vdd.n442 gnd 0.008187f
C2536 vdd.n443 gnd 0.010172f
C2537 vdd.n444 gnd 0.008187f
C2538 vdd.n445 gnd 0.010172f
C2539 vdd.n446 gnd 0.008187f
C2540 vdd.n447 gnd 0.010172f
C2541 vdd.n448 gnd 0.008187f
C2542 vdd.n449 gnd 0.010172f
C2543 vdd.n450 gnd 0.008187f
C2544 vdd.n451 gnd 0.010172f
C2545 vdd.t29 gnd 0.125139f
C2546 vdd.t28 gnd 0.133739f
C2547 vdd.t27 gnd 0.16343f
C2548 vdd.n452 gnd 0.209494f
C2549 vdd.n453 gnd 0.176832f
C2550 vdd.n454 gnd 0.01752f
C2551 vdd.n455 gnd 0.010172f
C2552 vdd.n456 gnd 0.008187f
C2553 vdd.n457 gnd 0.010172f
C2554 vdd.n458 gnd 0.008187f
C2555 vdd.n459 gnd 0.010172f
C2556 vdd.n460 gnd 0.008187f
C2557 vdd.n461 gnd 0.010172f
C2558 vdd.n462 gnd 0.008187f
C2559 vdd.n463 gnd 0.010172f
C2560 vdd.n464 gnd 0.025134f
C2561 vdd.n465 gnd 0.006795f
C2562 vdd.n466 gnd 0.008187f
C2563 vdd.n467 gnd 0.010172f
C2564 vdd.n468 gnd 0.010172f
C2565 vdd.n469 gnd 0.008187f
C2566 vdd.n470 gnd 0.010172f
C2567 vdd.n471 gnd 0.010172f
C2568 vdd.n472 gnd 0.010172f
C2569 vdd.n473 gnd 0.010172f
C2570 vdd.n474 gnd 0.010172f
C2571 vdd.n475 gnd 0.008187f
C2572 vdd.n476 gnd 0.008187f
C2573 vdd.n477 gnd 0.010172f
C2574 vdd.n478 gnd 0.010172f
C2575 vdd.n479 gnd 0.008187f
C2576 vdd.n480 gnd 0.010172f
C2577 vdd.n481 gnd 0.010172f
C2578 vdd.n482 gnd 0.010172f
C2579 vdd.n483 gnd 0.010172f
C2580 vdd.n484 gnd 0.010172f
C2581 vdd.n485 gnd 0.008187f
C2582 vdd.n486 gnd 0.008187f
C2583 vdd.n487 gnd 0.010172f
C2584 vdd.n488 gnd 0.010172f
C2585 vdd.n489 gnd 0.008187f
C2586 vdd.n490 gnd 0.010172f
C2587 vdd.n491 gnd 0.010172f
C2588 vdd.n492 gnd 0.010172f
C2589 vdd.n493 gnd 0.010172f
C2590 vdd.n494 gnd 0.010172f
C2591 vdd.n495 gnd 0.008187f
C2592 vdd.n496 gnd 0.008187f
C2593 vdd.n497 gnd 0.010172f
C2594 vdd.n498 gnd 0.010172f
C2595 vdd.n499 gnd 0.008187f
C2596 vdd.n500 gnd 0.010172f
C2597 vdd.n501 gnd 0.010172f
C2598 vdd.n502 gnd 0.010172f
C2599 vdd.n503 gnd 0.010172f
C2600 vdd.n504 gnd 0.010172f
C2601 vdd.n505 gnd 0.008187f
C2602 vdd.n506 gnd 0.008187f
C2603 vdd.n507 gnd 0.010172f
C2604 vdd.n508 gnd 0.010172f
C2605 vdd.n509 gnd 0.006836f
C2606 vdd.n510 gnd 0.010172f
C2607 vdd.n511 gnd 0.010172f
C2608 vdd.n512 gnd 0.010172f
C2609 vdd.n513 gnd 0.010172f
C2610 vdd.n514 gnd 0.010172f
C2611 vdd.n515 gnd 0.006836f
C2612 vdd.n516 gnd 0.008187f
C2613 vdd.n517 gnd 0.010172f
C2614 vdd.n518 gnd 0.010172f
C2615 vdd.n519 gnd 0.008187f
C2616 vdd.n520 gnd 0.010172f
C2617 vdd.n521 gnd 0.010172f
C2618 vdd.n522 gnd 0.010172f
C2619 vdd.n523 gnd 0.010172f
C2620 vdd.n524 gnd 0.010172f
C2621 vdd.n525 gnd 0.008187f
C2622 vdd.n526 gnd 0.008187f
C2623 vdd.n527 gnd 0.010172f
C2624 vdd.n528 gnd 0.010172f
C2625 vdd.n529 gnd 0.008187f
C2626 vdd.n530 gnd 0.010172f
C2627 vdd.n531 gnd 0.010172f
C2628 vdd.n532 gnd 0.010172f
C2629 vdd.n533 gnd 0.010172f
C2630 vdd.n534 gnd 0.010172f
C2631 vdd.n535 gnd 0.008187f
C2632 vdd.n536 gnd 0.008187f
C2633 vdd.n537 gnd 0.010172f
C2634 vdd.n538 gnd 0.010172f
C2635 vdd.n539 gnd 0.008187f
C2636 vdd.n540 gnd 0.010172f
C2637 vdd.n541 gnd 0.010172f
C2638 vdd.n542 gnd 0.010172f
C2639 vdd.n543 gnd 0.010172f
C2640 vdd.n544 gnd 0.010172f
C2641 vdd.n545 gnd 0.008187f
C2642 vdd.n546 gnd 0.008187f
C2643 vdd.n547 gnd 0.010172f
C2644 vdd.n548 gnd 0.010172f
C2645 vdd.n549 gnd 0.008187f
C2646 vdd.n550 gnd 0.010172f
C2647 vdd.n551 gnd 0.010172f
C2648 vdd.n552 gnd 0.010172f
C2649 vdd.n553 gnd 0.010172f
C2650 vdd.n554 gnd 0.010172f
C2651 vdd.n555 gnd 0.008187f
C2652 vdd.n556 gnd 0.008187f
C2653 vdd.n557 gnd 0.010172f
C2654 vdd.n558 gnd 0.010172f
C2655 vdd.n559 gnd 0.008187f
C2656 vdd.n560 gnd 0.010172f
C2657 vdd.n561 gnd 0.010172f
C2658 vdd.n562 gnd 0.010172f
C2659 vdd.n563 gnd 0.010172f
C2660 vdd.n564 gnd 0.010172f
C2661 vdd.n565 gnd 0.005567f
C2662 vdd.n566 gnd 0.01752f
C2663 vdd.n567 gnd 0.010172f
C2664 vdd.n568 gnd 0.010172f
C2665 vdd.n569 gnd 0.008105f
C2666 vdd.n570 gnd 0.010172f
C2667 vdd.n571 gnd 0.010172f
C2668 vdd.n572 gnd 0.010172f
C2669 vdd.n573 gnd 0.010172f
C2670 vdd.n574 gnd 0.010172f
C2671 vdd.n575 gnd 0.008187f
C2672 vdd.n576 gnd 0.008187f
C2673 vdd.n577 gnd 0.010172f
C2674 vdd.n578 gnd 0.010172f
C2675 vdd.n579 gnd 0.008187f
C2676 vdd.n580 gnd 0.010172f
C2677 vdd.n581 gnd 0.010172f
C2678 vdd.n582 gnd 0.010172f
C2679 vdd.n583 gnd 0.010172f
C2680 vdd.n584 gnd 0.010172f
C2681 vdd.n585 gnd 0.008187f
C2682 vdd.n586 gnd 0.008187f
C2683 vdd.n587 gnd 0.010172f
C2684 vdd.n588 gnd 0.010172f
C2685 vdd.n589 gnd 0.008187f
C2686 vdd.n590 gnd 0.010172f
C2687 vdd.n591 gnd 0.010172f
C2688 vdd.n592 gnd 0.010172f
C2689 vdd.n593 gnd 0.010172f
C2690 vdd.n594 gnd 0.010172f
C2691 vdd.n595 gnd 0.008187f
C2692 vdd.n596 gnd 0.008187f
C2693 vdd.n597 gnd 0.010172f
C2694 vdd.n598 gnd 0.010172f
C2695 vdd.n599 gnd 0.008187f
C2696 vdd.n600 gnd 0.010172f
C2697 vdd.n601 gnd 0.010172f
C2698 vdd.n602 gnd 0.010172f
C2699 vdd.n603 gnd 0.010172f
C2700 vdd.n604 gnd 0.010172f
C2701 vdd.n605 gnd 0.008187f
C2702 vdd.n606 gnd 0.008187f
C2703 vdd.n607 gnd 0.010172f
C2704 vdd.n608 gnd 0.010172f
C2705 vdd.n609 gnd 0.008187f
C2706 vdd.n610 gnd 0.010172f
C2707 vdd.n611 gnd 0.010172f
C2708 vdd.n612 gnd 0.010172f
C2709 vdd.n613 gnd 0.010172f
C2710 vdd.n614 gnd 0.010172f
C2711 vdd.n615 gnd 0.008187f
C2712 vdd.n616 gnd 0.010172f
C2713 vdd.n617 gnd 0.008187f
C2714 vdd.n618 gnd 0.004298f
C2715 vdd.n619 gnd 0.010172f
C2716 vdd.n620 gnd 0.010172f
C2717 vdd.n621 gnd 0.008187f
C2718 vdd.n622 gnd 0.010172f
C2719 vdd.n623 gnd 0.008187f
C2720 vdd.n624 gnd 0.010172f
C2721 vdd.n625 gnd 0.008187f
C2722 vdd.n626 gnd 0.010172f
C2723 vdd.n627 gnd 0.008187f
C2724 vdd.n628 gnd 0.010172f
C2725 vdd.n629 gnd 0.008187f
C2726 vdd.n630 gnd 0.010172f
C2727 vdd.n631 gnd 0.008187f
C2728 vdd.n632 gnd 0.010172f
C2729 vdd.n633 gnd 0.56653f
C2730 vdd.t144 gnd 0.519752f
C2731 vdd.n634 gnd 0.010172f
C2732 vdd.n635 gnd 0.008187f
C2733 vdd.n636 gnd 0.010172f
C2734 vdd.n637 gnd 0.008187f
C2735 vdd.n638 gnd 0.010172f
C2736 vdd.t152 gnd 0.519752f
C2737 vdd.n639 gnd 0.010172f
C2738 vdd.n640 gnd 0.008187f
C2739 vdd.n641 gnd 0.010172f
C2740 vdd.n642 gnd 0.008187f
C2741 vdd.n643 gnd 0.010172f
C2742 vdd.t167 gnd 0.519752f
C2743 vdd.n644 gnd 0.64969f
C2744 vdd.n645 gnd 0.010172f
C2745 vdd.n646 gnd 0.008187f
C2746 vdd.n647 gnd 0.010172f
C2747 vdd.n648 gnd 0.008187f
C2748 vdd.n649 gnd 0.010172f
C2749 vdd.t102 gnd 0.519752f
C2750 vdd.n650 gnd 0.010172f
C2751 vdd.n651 gnd 0.008187f
C2752 vdd.n652 gnd 0.010172f
C2753 vdd.n653 gnd 0.008187f
C2754 vdd.n654 gnd 0.010172f
C2755 vdd.n655 gnd 0.722456f
C2756 vdd.n656 gnd 0.862789f
C2757 vdd.t200 gnd 0.519752f
C2758 vdd.n657 gnd 0.010172f
C2759 vdd.n658 gnd 0.008187f
C2760 vdd.n659 gnd 0.010172f
C2761 vdd.n660 gnd 0.008187f
C2762 vdd.n661 gnd 0.010172f
C2763 vdd.n662 gnd 0.54574f
C2764 vdd.n663 gnd 0.010172f
C2765 vdd.n664 gnd 0.008187f
C2766 vdd.n665 gnd 0.010172f
C2767 vdd.n666 gnd 0.008187f
C2768 vdd.n667 gnd 0.010172f
C2769 vdd.t140 gnd 0.519752f
C2770 vdd.t110 gnd 0.519752f
C2771 vdd.n668 gnd 0.010172f
C2772 vdd.n669 gnd 0.008187f
C2773 vdd.n670 gnd 0.010172f
C2774 vdd.n671 gnd 0.008187f
C2775 vdd.n672 gnd 0.010172f
C2776 vdd.t169 gnd 0.519752f
C2777 vdd.n673 gnd 0.010172f
C2778 vdd.n674 gnd 0.008187f
C2779 vdd.n675 gnd 0.010172f
C2780 vdd.n676 gnd 0.008187f
C2781 vdd.n677 gnd 0.010172f
C2782 vdd.n678 gnd 1.0395f
C2783 vdd.n679 gnd 0.847196f
C2784 vdd.n680 gnd 0.010172f
C2785 vdd.n681 gnd 0.008187f
C2786 vdd.n682 gnd 0.024606f
C2787 vdd.n683 gnd 0.006795f
C2788 vdd.n684 gnd 0.024606f
C2789 vdd.t34 gnd 0.519752f
C2790 vdd.n685 gnd 0.024606f
C2791 vdd.n686 gnd 0.006795f
C2792 vdd.n687 gnd 0.008748f
C2793 vdd.t35 gnd 0.125139f
C2794 vdd.t36 gnd 0.133739f
C2795 vdd.t33 gnd 0.16343f
C2796 vdd.n688 gnd 0.209494f
C2797 vdd.n689 gnd 0.176013f
C2798 vdd.n690 gnd 0.012608f
C2799 vdd.n691 gnd 0.010172f
C2800 vdd.n692 gnd 12.2765f
C2801 vdd.n723 gnd 1.42932f
C2802 vdd.n724 gnd 0.010172f
C2803 vdd.n725 gnd 0.010172f
C2804 vdd.n726 gnd 0.025134f
C2805 vdd.n727 gnd 0.008748f
C2806 vdd.n728 gnd 0.010172f
C2807 vdd.n729 gnd 0.008187f
C2808 vdd.n730 gnd 0.00651f
C2809 vdd.n731 gnd 0.04271f
C2810 vdd.n732 gnd 0.008187f
C2811 vdd.n733 gnd 0.010172f
C2812 vdd.n734 gnd 0.010172f
C2813 vdd.n735 gnd 0.010172f
C2814 vdd.n736 gnd 0.010172f
C2815 vdd.n737 gnd 0.010172f
C2816 vdd.n738 gnd 0.010172f
C2817 vdd.n739 gnd 0.010172f
C2818 vdd.n740 gnd 0.010172f
C2819 vdd.n741 gnd 0.010172f
C2820 vdd.n742 gnd 0.010172f
C2821 vdd.n743 gnd 0.010172f
C2822 vdd.n744 gnd 0.010172f
C2823 vdd.n745 gnd 0.010172f
C2824 vdd.n746 gnd 0.010172f
C2825 vdd.n747 gnd 0.006836f
C2826 vdd.n748 gnd 0.010172f
C2827 vdd.n749 gnd 0.010172f
C2828 vdd.n750 gnd 0.010172f
C2829 vdd.n751 gnd 0.010172f
C2830 vdd.n752 gnd 0.010172f
C2831 vdd.n753 gnd 0.010172f
C2832 vdd.n754 gnd 0.010172f
C2833 vdd.n755 gnd 0.010172f
C2834 vdd.n756 gnd 0.010172f
C2835 vdd.n757 gnd 0.010172f
C2836 vdd.n758 gnd 0.010172f
C2837 vdd.n759 gnd 0.010172f
C2838 vdd.n760 gnd 0.010172f
C2839 vdd.n761 gnd 0.010172f
C2840 vdd.n762 gnd 0.010172f
C2841 vdd.n763 gnd 0.010172f
C2842 vdd.n764 gnd 0.010172f
C2843 vdd.n765 gnd 0.010172f
C2844 vdd.n766 gnd 0.010172f
C2845 vdd.n767 gnd 0.008105f
C2846 vdd.t45 gnd 0.125139f
C2847 vdd.t46 gnd 0.133739f
C2848 vdd.t44 gnd 0.16343f
C2849 vdd.n768 gnd 0.209494f
C2850 vdd.n769 gnd 0.176013f
C2851 vdd.n770 gnd 0.010172f
C2852 vdd.n771 gnd 0.010172f
C2853 vdd.n772 gnd 0.010172f
C2854 vdd.n773 gnd 0.010172f
C2855 vdd.n774 gnd 0.010172f
C2856 vdd.n775 gnd 0.010172f
C2857 vdd.n776 gnd 0.010172f
C2858 vdd.n777 gnd 0.010172f
C2859 vdd.n778 gnd 0.010172f
C2860 vdd.n779 gnd 0.010172f
C2861 vdd.n780 gnd 0.010172f
C2862 vdd.n781 gnd 0.010172f
C2863 vdd.n782 gnd 0.010172f
C2864 vdd.n783 gnd 0.00651f
C2865 vdd.n785 gnd 0.006917f
C2866 vdd.n786 gnd 0.006917f
C2867 vdd.n787 gnd 0.006917f
C2868 vdd.n788 gnd 0.006917f
C2869 vdd.n789 gnd 0.006917f
C2870 vdd.n790 gnd 0.006917f
C2871 vdd.n792 gnd 0.006917f
C2872 vdd.n793 gnd 0.006917f
C2873 vdd.n795 gnd 0.006917f
C2874 vdd.n796 gnd 0.005035f
C2875 vdd.n798 gnd 0.006917f
C2876 vdd.t11 gnd 0.279506f
C2877 vdd.t10 gnd 0.28611f
C2878 vdd.t8 gnd 0.182472f
C2879 vdd.n799 gnd 0.098616f
C2880 vdd.n800 gnd 0.055938f
C2881 vdd.n801 gnd 0.009885f
C2882 vdd.n802 gnd 0.015705f
C2883 vdd.n804 gnd 0.006917f
C2884 vdd.n805 gnd 0.706863f
C2885 vdd.n806 gnd 0.01481f
C2886 vdd.n807 gnd 0.01481f
C2887 vdd.n808 gnd 0.006917f
C2888 vdd.n809 gnd 0.015705f
C2889 vdd.n810 gnd 0.006917f
C2890 vdd.n811 gnd 0.006917f
C2891 vdd.n812 gnd 0.006917f
C2892 vdd.n813 gnd 0.006917f
C2893 vdd.n814 gnd 0.006917f
C2894 vdd.n816 gnd 0.006917f
C2895 vdd.n817 gnd 0.006917f
C2896 vdd.n819 gnd 0.006917f
C2897 vdd.n820 gnd 0.006917f
C2898 vdd.n822 gnd 0.006917f
C2899 vdd.n823 gnd 0.006917f
C2900 vdd.n825 gnd 0.006917f
C2901 vdd.n826 gnd 0.006917f
C2902 vdd.n828 gnd 0.006917f
C2903 vdd.n829 gnd 0.006917f
C2904 vdd.n831 gnd 0.006917f
C2905 vdd.t32 gnd 0.279506f
C2906 vdd.t31 gnd 0.28611f
C2907 vdd.t30 gnd 0.182472f
C2908 vdd.n832 gnd 0.098616f
C2909 vdd.n833 gnd 0.055938f
C2910 vdd.n834 gnd 0.006917f
C2911 vdd.n836 gnd 0.006917f
C2912 vdd.n837 gnd 0.006917f
C2913 vdd.t9 gnd 0.353431f
C2914 vdd.n838 gnd 0.006917f
C2915 vdd.n839 gnd 0.006917f
C2916 vdd.n840 gnd 0.006917f
C2917 vdd.n841 gnd 0.006917f
C2918 vdd.n842 gnd 0.006917f
C2919 vdd.n843 gnd 0.706863f
C2920 vdd.n844 gnd 0.006917f
C2921 vdd.n845 gnd 0.006917f
C2922 vdd.n846 gnd 0.556135f
C2923 vdd.n847 gnd 0.006917f
C2924 vdd.n848 gnd 0.006917f
C2925 vdd.n849 gnd 0.006917f
C2926 vdd.n850 gnd 0.006917f
C2927 vdd.n851 gnd 0.706863f
C2928 vdd.n852 gnd 0.006917f
C2929 vdd.n853 gnd 0.006917f
C2930 vdd.n854 gnd 0.006917f
C2931 vdd.n855 gnd 0.006917f
C2932 vdd.n856 gnd 0.006917f
C2933 vdd.t262 gnd 0.353431f
C2934 vdd.n857 gnd 0.006917f
C2935 vdd.n858 gnd 0.006917f
C2936 vdd.n859 gnd 0.006917f
C2937 vdd.n860 gnd 0.006917f
C2938 vdd.n861 gnd 0.006917f
C2939 vdd.t281 gnd 0.353431f
C2940 vdd.n862 gnd 0.006917f
C2941 vdd.n863 gnd 0.006917f
C2942 vdd.n864 gnd 0.680875f
C2943 vdd.n865 gnd 0.006917f
C2944 vdd.n866 gnd 0.006917f
C2945 vdd.n867 gnd 0.006917f
C2946 vdd.t280 gnd 0.353431f
C2947 vdd.n868 gnd 0.006917f
C2948 vdd.n869 gnd 0.006917f
C2949 vdd.n870 gnd 0.52495f
C2950 vdd.n871 gnd 0.006917f
C2951 vdd.n872 gnd 0.006917f
C2952 vdd.n873 gnd 0.006917f
C2953 vdd.n874 gnd 0.493765f
C2954 vdd.n875 gnd 0.006917f
C2955 vdd.n876 gnd 0.006917f
C2956 vdd.n877 gnd 0.369024f
C2957 vdd.n878 gnd 0.006917f
C2958 vdd.n879 gnd 0.006917f
C2959 vdd.n880 gnd 0.006917f
C2960 vdd.n881 gnd 0.64969f
C2961 vdd.n882 gnd 0.006917f
C2962 vdd.n883 gnd 0.006917f
C2963 vdd.t285 gnd 0.353431f
C2964 vdd.n884 gnd 0.006917f
C2965 vdd.n885 gnd 0.006917f
C2966 vdd.n886 gnd 0.006917f
C2967 vdd.n887 gnd 0.706863f
C2968 vdd.n888 gnd 0.006917f
C2969 vdd.n889 gnd 0.006917f
C2970 vdd.t286 gnd 0.353431f
C2971 vdd.n890 gnd 0.006917f
C2972 vdd.n891 gnd 0.006917f
C2973 vdd.n892 gnd 0.006917f
C2974 vdd.t256 gnd 0.353431f
C2975 vdd.n893 gnd 0.006917f
C2976 vdd.n894 gnd 0.006917f
C2977 vdd.n895 gnd 0.006917f
C2978 vdd.t39 gnd 0.28611f
C2979 vdd.t37 gnd 0.182472f
C2980 vdd.t40 gnd 0.28611f
C2981 vdd.n896 gnd 0.160805f
C2982 vdd.n897 gnd 0.020037f
C2983 vdd.n898 gnd 0.006917f
C2984 vdd.t38 gnd 0.254679f
C2985 vdd.n899 gnd 0.006917f
C2986 vdd.n900 gnd 0.006917f
C2987 vdd.n901 gnd 0.60811f
C2988 vdd.n902 gnd 0.006917f
C2989 vdd.n903 gnd 0.006917f
C2990 vdd.n904 gnd 0.006917f
C2991 vdd.n905 gnd 0.410604f
C2992 vdd.n906 gnd 0.006917f
C2993 vdd.n907 gnd 0.006917f
C2994 vdd.t257 gnd 0.145531f
C2995 vdd.n908 gnd 0.452184f
C2996 vdd.n909 gnd 0.006917f
C2997 vdd.n910 gnd 0.006917f
C2998 vdd.n911 gnd 0.006917f
C2999 vdd.n912 gnd 0.56653f
C3000 vdd.n913 gnd 0.006917f
C3001 vdd.n914 gnd 0.006917f
C3002 vdd.t272 gnd 0.353431f
C3003 vdd.n915 gnd 0.006917f
C3004 vdd.n916 gnd 0.006917f
C3005 vdd.n917 gnd 0.006917f
C3006 vdd.t266 gnd 0.353431f
C3007 vdd.n918 gnd 0.006917f
C3008 vdd.n919 gnd 0.006917f
C3009 vdd.t289 gnd 0.353431f
C3010 vdd.n920 gnd 0.006917f
C3011 vdd.n921 gnd 0.006917f
C3012 vdd.n922 gnd 0.006917f
C3013 vdd.t248 gnd 0.239086f
C3014 vdd.n923 gnd 0.006917f
C3015 vdd.n924 gnd 0.006917f
C3016 vdd.n925 gnd 0.623703f
C3017 vdd.n926 gnd 0.006917f
C3018 vdd.n927 gnd 0.006917f
C3019 vdd.n928 gnd 0.006917f
C3020 vdd.t290 gnd 0.353431f
C3021 vdd.n929 gnd 0.006917f
C3022 vdd.n930 gnd 0.006917f
C3023 vdd.t302 gnd 0.337839f
C3024 vdd.n931 gnd 0.467777f
C3025 vdd.n932 gnd 0.006917f
C3026 vdd.n933 gnd 0.006917f
C3027 vdd.n934 gnd 0.006917f
C3028 vdd.t252 gnd 0.353431f
C3029 vdd.n935 gnd 0.006917f
C3030 vdd.n936 gnd 0.006917f
C3031 vdd.t294 gnd 0.353431f
C3032 vdd.n937 gnd 0.006917f
C3033 vdd.n938 gnd 0.006917f
C3034 vdd.n939 gnd 0.006917f
C3035 vdd.n940 gnd 0.706863f
C3036 vdd.n941 gnd 0.006917f
C3037 vdd.n942 gnd 0.006917f
C3038 vdd.t276 gnd 0.353431f
C3039 vdd.n943 gnd 0.006917f
C3040 vdd.n944 gnd 0.006917f
C3041 vdd.n945 gnd 0.006917f
C3042 vdd.n946 gnd 0.488567f
C3043 vdd.n947 gnd 0.006917f
C3044 vdd.n948 gnd 0.006917f
C3045 vdd.n949 gnd 0.006917f
C3046 vdd.n950 gnd 0.006917f
C3047 vdd.n951 gnd 0.006917f
C3048 vdd.t61 gnd 0.353431f
C3049 vdd.n952 gnd 0.006917f
C3050 vdd.n953 gnd 0.006917f
C3051 vdd.t254 gnd 0.353431f
C3052 vdd.n954 gnd 0.006917f
C3053 vdd.n955 gnd 0.01481f
C3054 vdd.n956 gnd 0.01481f
C3055 vdd.n957 gnd 0.800418f
C3056 vdd.n958 gnd 0.006917f
C3057 vdd.n959 gnd 0.006917f
C3058 vdd.t283 gnd 0.353431f
C3059 vdd.n960 gnd 0.01481f
C3060 vdd.n961 gnd 0.006917f
C3061 vdd.n962 gnd 0.006917f
C3062 vdd.t296 gnd 0.602912f
C3063 vdd.n980 gnd 0.015705f
C3064 vdd.n998 gnd 0.01481f
C3065 vdd.n999 gnd 0.006917f
C3066 vdd.n1000 gnd 0.01481f
C3067 vdd.t77 gnd 0.279506f
C3068 vdd.t76 gnd 0.28611f
C3069 vdd.t75 gnd 0.182472f
C3070 vdd.n1001 gnd 0.098616f
C3071 vdd.n1002 gnd 0.055938f
C3072 vdd.n1003 gnd 0.015705f
C3073 vdd.n1004 gnd 0.006917f
C3074 vdd.n1005 gnd 0.415802f
C3075 vdd.n1006 gnd 0.01481f
C3076 vdd.n1007 gnd 0.006917f
C3077 vdd.n1008 gnd 0.015705f
C3078 vdd.n1009 gnd 0.006917f
C3079 vdd.t56 gnd 0.279506f
C3080 vdd.t55 gnd 0.28611f
C3081 vdd.t53 gnd 0.182472f
C3082 vdd.n1010 gnd 0.098616f
C3083 vdd.n1011 gnd 0.055938f
C3084 vdd.n1012 gnd 0.009885f
C3085 vdd.n1013 gnd 0.006917f
C3086 vdd.n1014 gnd 0.006917f
C3087 vdd.t54 gnd 0.353431f
C3088 vdd.n1015 gnd 0.006917f
C3089 vdd.t298 gnd 0.353431f
C3090 vdd.n1016 gnd 0.006917f
C3091 vdd.n1017 gnd 0.006917f
C3092 vdd.n1018 gnd 0.006917f
C3093 vdd.n1019 gnd 0.006917f
C3094 vdd.n1020 gnd 0.006917f
C3095 vdd.n1021 gnd 0.706863f
C3096 vdd.n1022 gnd 0.006917f
C3097 vdd.n1023 gnd 0.006917f
C3098 vdd.t268 gnd 0.353431f
C3099 vdd.n1024 gnd 0.006917f
C3100 vdd.n1025 gnd 0.006917f
C3101 vdd.n1026 gnd 0.006917f
C3102 vdd.n1027 gnd 0.006917f
C3103 vdd.n1028 gnd 0.509357f
C3104 vdd.n1029 gnd 0.006917f
C3105 vdd.n1030 gnd 0.006917f
C3106 vdd.n1031 gnd 0.006917f
C3107 vdd.n1032 gnd 0.006917f
C3108 vdd.n1033 gnd 0.006917f
C3109 vdd.t249 gnd 0.353431f
C3110 vdd.n1034 gnd 0.006917f
C3111 vdd.n1035 gnd 0.006917f
C3112 vdd.t287 gnd 0.353431f
C3113 vdd.n1036 gnd 0.006917f
C3114 vdd.n1037 gnd 0.006917f
C3115 vdd.n1038 gnd 0.006917f
C3116 vdd.t275 gnd 0.353431f
C3117 vdd.n1039 gnd 0.006917f
C3118 vdd.n1040 gnd 0.006917f
C3119 vdd.t250 gnd 0.353431f
C3120 vdd.n1041 gnd 0.006917f
C3121 vdd.n1042 gnd 0.006917f
C3122 vdd.n1043 gnd 0.006917f
C3123 vdd.t273 gnd 0.337839f
C3124 vdd.n1044 gnd 0.006917f
C3125 vdd.n1045 gnd 0.006917f
C3126 vdd.n1046 gnd 0.52495f
C3127 vdd.n1047 gnd 0.006917f
C3128 vdd.n1048 gnd 0.006917f
C3129 vdd.n1049 gnd 0.006917f
C3130 vdd.t291 gnd 0.353431f
C3131 vdd.n1050 gnd 0.006917f
C3132 vdd.n1051 gnd 0.006917f
C3133 vdd.t259 gnd 0.239086f
C3134 vdd.n1052 gnd 0.369024f
C3135 vdd.n1053 gnd 0.006917f
C3136 vdd.n1054 gnd 0.006917f
C3137 vdd.n1055 gnd 0.006917f
C3138 vdd.n1056 gnd 0.64969f
C3139 vdd.n1057 gnd 0.006917f
C3140 vdd.n1058 gnd 0.006917f
C3141 vdd.t300 gnd 0.353431f
C3142 vdd.n1059 gnd 0.006917f
C3143 vdd.n1060 gnd 0.006917f
C3144 vdd.n1061 gnd 0.006917f
C3145 vdd.n1062 gnd 0.706863f
C3146 vdd.n1063 gnd 0.006917f
C3147 vdd.n1064 gnd 0.006917f
C3148 vdd.t265 gnd 0.353431f
C3149 vdd.n1065 gnd 0.006917f
C3150 vdd.n1066 gnd 0.006917f
C3151 vdd.n1067 gnd 0.006917f
C3152 vdd.t258 gnd 0.145531f
C3153 vdd.n1068 gnd 0.006917f
C3154 vdd.n1069 gnd 0.006917f
C3155 vdd.n1070 gnd 0.006917f
C3156 vdd.t66 gnd 0.28611f
C3157 vdd.t64 gnd 0.182472f
C3158 vdd.t67 gnd 0.28611f
C3159 vdd.n1071 gnd 0.160805f
C3160 vdd.n1072 gnd 0.006917f
C3161 vdd.n1073 gnd 0.006917f
C3162 vdd.t282 gnd 0.353431f
C3163 vdd.n1074 gnd 0.006917f
C3164 vdd.n1075 gnd 0.006917f
C3165 vdd.t65 gnd 0.254679f
C3166 vdd.n1076 gnd 0.561332f
C3167 vdd.n1077 gnd 0.006917f
C3168 vdd.n1078 gnd 0.006917f
C3169 vdd.n1079 gnd 0.006917f
C3170 vdd.n1080 gnd 0.410604f
C3171 vdd.n1081 gnd 0.006917f
C3172 vdd.n1082 gnd 0.006917f
C3173 vdd.n1083 gnd 0.452184f
C3174 vdd.n1084 gnd 0.006917f
C3175 vdd.n1085 gnd 0.006917f
C3176 vdd.n1086 gnd 0.006917f
C3177 vdd.n1087 gnd 0.56653f
C3178 vdd.n1088 gnd 0.006917f
C3179 vdd.n1089 gnd 0.006917f
C3180 vdd.t260 gnd 0.353431f
C3181 vdd.n1090 gnd 0.006917f
C3182 vdd.n1091 gnd 0.006917f
C3183 vdd.n1092 gnd 0.006917f
C3184 vdd.n1093 gnd 0.706863f
C3185 vdd.n1094 gnd 0.006917f
C3186 vdd.n1095 gnd 0.006917f
C3187 vdd.t261 gnd 0.353431f
C3188 vdd.n1096 gnd 0.006917f
C3189 vdd.n1097 gnd 0.006917f
C3190 vdd.n1098 gnd 0.006917f
C3191 vdd.t301 gnd 0.353431f
C3192 vdd.n1099 gnd 0.006917f
C3193 vdd.n1100 gnd 0.006917f
C3194 vdd.n1101 gnd 0.006917f
C3195 vdd.n1102 gnd 0.006917f
C3196 vdd.n1103 gnd 0.006917f
C3197 vdd.t293 gnd 0.353431f
C3198 vdd.n1104 gnd 0.006917f
C3199 vdd.n1105 gnd 0.006917f
C3200 vdd.n1106 gnd 0.69127f
C3201 vdd.n1107 gnd 0.006917f
C3202 vdd.n1108 gnd 0.006917f
C3203 vdd.n1109 gnd 0.006917f
C3204 vdd.t253 gnd 0.353431f
C3205 vdd.n1110 gnd 0.006917f
C3206 vdd.n1111 gnd 0.006917f
C3207 vdd.n1112 gnd 0.535345f
C3208 vdd.n1113 gnd 0.006917f
C3209 vdd.n1114 gnd 0.006917f
C3210 vdd.n1115 gnd 0.006917f
C3211 vdd.n1116 gnd 0.706863f
C3212 vdd.n1117 gnd 0.006917f
C3213 vdd.n1118 gnd 0.006917f
C3214 vdd.n1119 gnd 0.379419f
C3215 vdd.n1120 gnd 0.006917f
C3216 vdd.n1121 gnd 0.006917f
C3217 vdd.n1122 gnd 0.006917f
C3218 vdd.n1123 gnd 0.706863f
C3219 vdd.n1124 gnd 0.006917f
C3220 vdd.n1125 gnd 0.006917f
C3221 vdd.n1126 gnd 0.006917f
C3222 vdd.n1127 gnd 0.006917f
C3223 vdd.n1128 gnd 0.006917f
C3224 vdd.t13 gnd 0.353431f
C3225 vdd.n1129 gnd 0.006917f
C3226 vdd.n1130 gnd 0.006917f
C3227 vdd.n1131 gnd 0.006917f
C3228 vdd.n1132 gnd 0.01481f
C3229 vdd.n1133 gnd 0.01481f
C3230 vdd.n1134 gnd 0.956344f
C3231 vdd.n1135 gnd 0.006917f
C3232 vdd.n1136 gnd 0.006917f
C3233 vdd.n1137 gnd 0.50416f
C3234 vdd.n1138 gnd 0.01481f
C3235 vdd.n1139 gnd 0.006917f
C3236 vdd.n1140 gnd 0.006917f
C3237 vdd.n1141 gnd 12.6923f
C3238 vdd.n1175 gnd 0.015705f
C3239 vdd.n1176 gnd 0.006917f
C3240 vdd.n1177 gnd 0.006917f
C3241 vdd.n1178 gnd 0.00651f
C3242 vdd.n1181 gnd 0.025134f
C3243 vdd.n1182 gnd 0.006795f
C3244 vdd.n1183 gnd 0.008187f
C3245 vdd.n1185 gnd 0.010172f
C3246 vdd.n1186 gnd 0.010172f
C3247 vdd.n1187 gnd 0.008187f
C3248 vdd.n1189 gnd 0.010172f
C3249 vdd.n1190 gnd 0.010172f
C3250 vdd.n1191 gnd 0.010172f
C3251 vdd.n1192 gnd 0.010172f
C3252 vdd.n1193 gnd 0.010172f
C3253 vdd.n1194 gnd 0.008187f
C3254 vdd.n1196 gnd 0.010172f
C3255 vdd.n1197 gnd 0.010172f
C3256 vdd.n1198 gnd 0.010172f
C3257 vdd.n1199 gnd 0.010172f
C3258 vdd.n1200 gnd 0.010172f
C3259 vdd.n1201 gnd 0.008187f
C3260 vdd.n1203 gnd 0.010172f
C3261 vdd.n1204 gnd 0.010172f
C3262 vdd.n1205 gnd 0.010172f
C3263 vdd.n1206 gnd 0.010172f
C3264 vdd.n1207 gnd 0.006836f
C3265 vdd.t26 gnd 0.125139f
C3266 vdd.t25 gnd 0.133739f
C3267 vdd.t24 gnd 0.16343f
C3268 vdd.n1208 gnd 0.209494f
C3269 vdd.n1209 gnd 0.176013f
C3270 vdd.n1211 gnd 0.010172f
C3271 vdd.n1212 gnd 0.010172f
C3272 vdd.n1213 gnd 0.008187f
C3273 vdd.n1214 gnd 0.010172f
C3274 vdd.n1216 gnd 0.010172f
C3275 vdd.n1217 gnd 0.010172f
C3276 vdd.n1218 gnd 0.010172f
C3277 vdd.n1219 gnd 0.010172f
C3278 vdd.n1220 gnd 0.008187f
C3279 vdd.n1222 gnd 0.010172f
C3280 vdd.n1223 gnd 0.010172f
C3281 vdd.n1224 gnd 0.010172f
C3282 vdd.n1225 gnd 0.010172f
C3283 vdd.n1226 gnd 0.010172f
C3284 vdd.n1227 gnd 0.008187f
C3285 vdd.n1229 gnd 0.010172f
C3286 vdd.n1230 gnd 0.010172f
C3287 vdd.n1231 gnd 0.010172f
C3288 vdd.n1232 gnd 0.010172f
C3289 vdd.n1233 gnd 0.010172f
C3290 vdd.n1234 gnd 0.008187f
C3291 vdd.n1236 gnd 0.010172f
C3292 vdd.n1237 gnd 0.010172f
C3293 vdd.n1238 gnd 0.010172f
C3294 vdd.n1239 gnd 0.010172f
C3295 vdd.n1240 gnd 0.010172f
C3296 vdd.n1241 gnd 0.008187f
C3297 vdd.n1243 gnd 0.010172f
C3298 vdd.n1244 gnd 0.010172f
C3299 vdd.n1245 gnd 0.010172f
C3300 vdd.n1246 gnd 0.010172f
C3301 vdd.n1247 gnd 0.008105f
C3302 vdd.t19 gnd 0.125139f
C3303 vdd.t18 gnd 0.133739f
C3304 vdd.t16 gnd 0.16343f
C3305 vdd.n1248 gnd 0.209494f
C3306 vdd.n1249 gnd 0.176013f
C3307 vdd.n1251 gnd 0.010172f
C3308 vdd.n1252 gnd 0.010172f
C3309 vdd.n1253 gnd 0.008187f
C3310 vdd.n1254 gnd 0.010172f
C3311 vdd.n1256 gnd 0.010172f
C3312 vdd.n1257 gnd 0.010172f
C3313 vdd.n1258 gnd 0.010172f
C3314 vdd.n1259 gnd 0.010172f
C3315 vdd.n1260 gnd 0.008187f
C3316 vdd.n1262 gnd 0.010172f
C3317 vdd.n1263 gnd 0.010172f
C3318 vdd.n1264 gnd 0.010172f
C3319 vdd.n1265 gnd 0.010172f
C3320 vdd.n1266 gnd 0.010172f
C3321 vdd.n1267 gnd 0.008187f
C3322 vdd.n1269 gnd 0.010172f
C3323 vdd.n1270 gnd 0.010172f
C3324 vdd.n1271 gnd 0.010172f
C3325 vdd.n1272 gnd 0.010172f
C3326 vdd.n1273 gnd 0.010172f
C3327 vdd.n1274 gnd 0.008187f
C3328 vdd.n1276 gnd 0.010172f
C3329 vdd.n1277 gnd 0.010172f
C3330 vdd.n1278 gnd 0.00651f
C3331 vdd.n1279 gnd 0.008187f
C3332 vdd.n1280 gnd 0.015705f
C3333 vdd.n1281 gnd 0.015705f
C3334 vdd.n1282 gnd 0.006917f
C3335 vdd.n1283 gnd 0.006917f
C3336 vdd.n1284 gnd 0.006917f
C3337 vdd.n1285 gnd 0.006917f
C3338 vdd.n1286 gnd 0.006917f
C3339 vdd.n1287 gnd 0.006917f
C3340 vdd.n1288 gnd 0.006917f
C3341 vdd.n1289 gnd 0.006917f
C3342 vdd.n1290 gnd 0.006917f
C3343 vdd.n1291 gnd 0.006917f
C3344 vdd.n1292 gnd 0.006917f
C3345 vdd.n1293 gnd 0.006917f
C3346 vdd.n1294 gnd 0.006917f
C3347 vdd.n1295 gnd 0.006917f
C3348 vdd.n1296 gnd 0.006917f
C3349 vdd.n1297 gnd 0.006917f
C3350 vdd.n1298 gnd 0.006917f
C3351 vdd.n1299 gnd 0.006917f
C3352 vdd.n1300 gnd 0.006917f
C3353 vdd.n1301 gnd 0.006917f
C3354 vdd.n1302 gnd 0.006917f
C3355 vdd.n1303 gnd 0.006917f
C3356 vdd.n1304 gnd 0.006917f
C3357 vdd.n1305 gnd 0.006917f
C3358 vdd.n1306 gnd 0.006917f
C3359 vdd.n1307 gnd 0.006917f
C3360 vdd.n1308 gnd 0.006917f
C3361 vdd.n1309 gnd 0.006917f
C3362 vdd.n1310 gnd 0.006917f
C3363 vdd.n1311 gnd 0.006917f
C3364 vdd.n1312 gnd 0.006917f
C3365 vdd.n1313 gnd 0.006917f
C3366 vdd.n1314 gnd 0.006917f
C3367 vdd.t14 gnd 0.279506f
C3368 vdd.t15 gnd 0.28611f
C3369 vdd.t12 gnd 0.182472f
C3370 vdd.n1315 gnd 0.098616f
C3371 vdd.n1316 gnd 0.055938f
C3372 vdd.n1317 gnd 0.009885f
C3373 vdd.n1318 gnd 0.006917f
C3374 vdd.t51 gnd 0.279506f
C3375 vdd.t52 gnd 0.28611f
C3376 vdd.t50 gnd 0.182472f
C3377 vdd.n1319 gnd 0.098616f
C3378 vdd.n1320 gnd 0.055938f
C3379 vdd.n1321 gnd 0.006917f
C3380 vdd.n1322 gnd 0.006917f
C3381 vdd.n1323 gnd 0.006917f
C3382 vdd.n1324 gnd 0.006917f
C3383 vdd.n1325 gnd 0.006917f
C3384 vdd.n1326 gnd 0.006917f
C3385 vdd.n1327 gnd 0.006917f
C3386 vdd.n1328 gnd 0.006917f
C3387 vdd.n1329 gnd 0.006917f
C3388 vdd.n1330 gnd 0.006917f
C3389 vdd.n1331 gnd 0.006917f
C3390 vdd.n1332 gnd 0.006917f
C3391 vdd.n1333 gnd 0.006917f
C3392 vdd.n1334 gnd 0.006917f
C3393 vdd.n1335 gnd 0.006917f
C3394 vdd.n1336 gnd 0.006917f
C3395 vdd.n1337 gnd 0.006917f
C3396 vdd.n1338 gnd 0.006917f
C3397 vdd.n1339 gnd 0.006917f
C3398 vdd.n1340 gnd 0.006917f
C3399 vdd.n1341 gnd 0.006917f
C3400 vdd.n1342 gnd 0.006917f
C3401 vdd.n1343 gnd 0.006917f
C3402 vdd.n1344 gnd 0.006917f
C3403 vdd.n1345 gnd 0.006917f
C3404 vdd.n1346 gnd 0.006917f
C3405 vdd.n1347 gnd 0.005035f
C3406 vdd.n1348 gnd 0.009885f
C3407 vdd.n1349 gnd 0.00534f
C3408 vdd.n1350 gnd 0.006917f
C3409 vdd.n1351 gnd 0.006917f
C3410 vdd.n1352 gnd 0.006917f
C3411 vdd.n1353 gnd 0.015705f
C3412 vdd.n1354 gnd 0.015705f
C3413 vdd.n1355 gnd 0.01481f
C3414 vdd.n1356 gnd 0.01481f
C3415 vdd.n1357 gnd 0.006917f
C3416 vdd.n1358 gnd 0.006917f
C3417 vdd.n1359 gnd 0.006917f
C3418 vdd.n1360 gnd 0.006917f
C3419 vdd.n1361 gnd 0.006917f
C3420 vdd.n1362 gnd 0.006917f
C3421 vdd.n1363 gnd 0.006917f
C3422 vdd.n1364 gnd 0.006917f
C3423 vdd.n1365 gnd 0.006917f
C3424 vdd.n1366 gnd 0.006917f
C3425 vdd.n1367 gnd 0.006917f
C3426 vdd.n1368 gnd 0.006917f
C3427 vdd.n1369 gnd 0.006917f
C3428 vdd.n1370 gnd 0.006917f
C3429 vdd.n1371 gnd 0.006917f
C3430 vdd.n1372 gnd 0.006917f
C3431 vdd.n1373 gnd 0.006917f
C3432 vdd.n1374 gnd 0.006917f
C3433 vdd.n1375 gnd 0.006917f
C3434 vdd.n1376 gnd 0.006917f
C3435 vdd.n1377 gnd 0.006917f
C3436 vdd.n1378 gnd 0.006917f
C3437 vdd.n1379 gnd 0.006917f
C3438 vdd.n1380 gnd 0.006917f
C3439 vdd.n1381 gnd 0.006917f
C3440 vdd.n1382 gnd 0.006917f
C3441 vdd.n1383 gnd 0.006917f
C3442 vdd.n1384 gnd 0.006917f
C3443 vdd.n1385 gnd 0.006917f
C3444 vdd.n1386 gnd 0.006917f
C3445 vdd.n1387 gnd 0.006917f
C3446 vdd.n1388 gnd 0.006917f
C3447 vdd.n1389 gnd 0.006917f
C3448 vdd.n1390 gnd 0.006917f
C3449 vdd.n1391 gnd 0.006917f
C3450 vdd.n1392 gnd 0.006917f
C3451 vdd.n1393 gnd 0.006917f
C3452 vdd.n1394 gnd 0.006917f
C3453 vdd.n1395 gnd 0.006917f
C3454 vdd.n1396 gnd 0.006917f
C3455 vdd.n1397 gnd 0.006917f
C3456 vdd.n1398 gnd 0.006917f
C3457 vdd.n1399 gnd 0.420999f
C3458 vdd.n1400 gnd 0.006917f
C3459 vdd.n1401 gnd 0.006917f
C3460 vdd.n1402 gnd 0.006917f
C3461 vdd.n1403 gnd 0.006917f
C3462 vdd.n1404 gnd 0.006917f
C3463 vdd.n1405 gnd 0.006917f
C3464 vdd.n1406 gnd 0.006917f
C3465 vdd.n1407 gnd 0.006917f
C3466 vdd.n1408 gnd 0.006917f
C3467 vdd.n1409 gnd 0.006917f
C3468 vdd.n1410 gnd 0.006917f
C3469 vdd.n1411 gnd 0.006917f
C3470 vdd.n1412 gnd 0.006917f
C3471 vdd.n1413 gnd 0.006917f
C3472 vdd.n1414 gnd 0.006917f
C3473 vdd.n1415 gnd 0.006917f
C3474 vdd.n1416 gnd 0.006917f
C3475 vdd.n1417 gnd 0.006917f
C3476 vdd.n1418 gnd 0.006917f
C3477 vdd.n1419 gnd 0.006917f
C3478 vdd.n1420 gnd 0.006917f
C3479 vdd.n1421 gnd 0.006917f
C3480 vdd.n1422 gnd 0.006917f
C3481 vdd.n1423 gnd 0.006917f
C3482 vdd.n1424 gnd 0.006917f
C3483 vdd.n1425 gnd 0.639295f
C3484 vdd.n1426 gnd 0.006917f
C3485 vdd.n1427 gnd 0.006917f
C3486 vdd.n1428 gnd 0.006917f
C3487 vdd.n1429 gnd 0.006917f
C3488 vdd.n1430 gnd 0.006917f
C3489 vdd.n1431 gnd 0.006917f
C3490 vdd.n1432 gnd 0.006917f
C3491 vdd.n1433 gnd 0.006917f
C3492 vdd.n1434 gnd 0.006917f
C3493 vdd.n1435 gnd 0.006917f
C3494 vdd.n1436 gnd 0.006917f
C3495 vdd.n1437 gnd 0.223493f
C3496 vdd.n1438 gnd 0.006917f
C3497 vdd.n1439 gnd 0.006917f
C3498 vdd.n1440 gnd 0.006917f
C3499 vdd.n1441 gnd 0.006917f
C3500 vdd.n1442 gnd 0.006917f
C3501 vdd.n1443 gnd 0.006917f
C3502 vdd.n1444 gnd 0.006917f
C3503 vdd.n1445 gnd 0.006917f
C3504 vdd.n1446 gnd 0.006917f
C3505 vdd.n1447 gnd 0.006917f
C3506 vdd.n1448 gnd 0.006917f
C3507 vdd.n1449 gnd 0.006917f
C3508 vdd.n1450 gnd 0.006917f
C3509 vdd.n1451 gnd 0.006917f
C3510 vdd.n1452 gnd 0.006917f
C3511 vdd.n1453 gnd 0.006917f
C3512 vdd.n1454 gnd 0.006917f
C3513 vdd.n1455 gnd 0.006917f
C3514 vdd.n1456 gnd 0.006917f
C3515 vdd.n1457 gnd 0.006917f
C3516 vdd.n1458 gnd 0.006917f
C3517 vdd.n1459 gnd 0.006917f
C3518 vdd.n1460 gnd 0.006917f
C3519 vdd.n1461 gnd 0.006917f
C3520 vdd.n1462 gnd 0.006917f
C3521 vdd.n1463 gnd 0.006917f
C3522 vdd.n1464 gnd 0.006917f
C3523 vdd.n1465 gnd 0.006917f
C3524 vdd.n1466 gnd 0.006917f
C3525 vdd.n1467 gnd 0.006917f
C3526 vdd.n1468 gnd 0.006917f
C3527 vdd.n1469 gnd 0.006917f
C3528 vdd.n1470 gnd 0.006917f
C3529 vdd.n1471 gnd 0.006917f
C3530 vdd.n1472 gnd 0.006917f
C3531 vdd.n1473 gnd 0.006917f
C3532 vdd.n1474 gnd 0.006917f
C3533 vdd.n1475 gnd 0.006917f
C3534 vdd.n1476 gnd 0.006917f
C3535 vdd.n1477 gnd 0.006917f
C3536 vdd.n1478 gnd 0.006917f
C3537 vdd.n1479 gnd 0.006917f
C3538 vdd.n1480 gnd 0.01481f
C3539 vdd.n1481 gnd 0.01481f
C3540 vdd.n1482 gnd 0.015705f
C3541 vdd.n1483 gnd 0.006917f
C3542 vdd.n1484 gnd 0.006917f
C3543 vdd.n1485 gnd 0.00534f
C3544 vdd.n1486 gnd 0.006917f
C3545 vdd.n1487 gnd 0.006917f
C3546 vdd.n1488 gnd 0.005035f
C3547 vdd.n1489 gnd 0.006917f
C3548 vdd.n1490 gnd 0.006917f
C3549 vdd.n1491 gnd 0.006917f
C3550 vdd.n1492 gnd 0.006917f
C3551 vdd.n1493 gnd 0.006917f
C3552 vdd.n1494 gnd 0.006917f
C3553 vdd.n1495 gnd 0.006917f
C3554 vdd.n1496 gnd 0.006917f
C3555 vdd.n1497 gnd 0.006917f
C3556 vdd.n1498 gnd 0.006917f
C3557 vdd.n1499 gnd 0.006917f
C3558 vdd.n1500 gnd 0.006917f
C3559 vdd.n1501 gnd 0.006917f
C3560 vdd.n1502 gnd 0.006917f
C3561 vdd.n1503 gnd 0.006917f
C3562 vdd.n1504 gnd 0.006917f
C3563 vdd.n1505 gnd 0.006917f
C3564 vdd.n1506 gnd 0.006917f
C3565 vdd.n1507 gnd 0.006917f
C3566 vdd.n1508 gnd 0.006917f
C3567 vdd.n1509 gnd 0.006917f
C3568 vdd.n1510 gnd 0.006917f
C3569 vdd.n1511 gnd 0.006917f
C3570 vdd.n1512 gnd 0.006917f
C3571 vdd.n1513 gnd 0.006917f
C3572 vdd.n1514 gnd 0.006917f
C3573 vdd.n1515 gnd 0.046595f
C3574 vdd.n1517 gnd 0.025134f
C3575 vdd.n1518 gnd 0.008187f
C3576 vdd.n1520 gnd 0.010172f
C3577 vdd.n1521 gnd 0.008187f
C3578 vdd.n1522 gnd 0.010172f
C3579 vdd.n1524 gnd 0.010172f
C3580 vdd.n1525 gnd 0.010172f
C3581 vdd.n1527 gnd 0.010172f
C3582 vdd.n1528 gnd 0.006795f
C3583 vdd.t17 gnd 0.519752f
C3584 vdd.n1529 gnd 0.010172f
C3585 vdd.n1530 gnd 0.025134f
C3586 vdd.n1531 gnd 0.008187f
C3587 vdd.n1532 gnd 0.010172f
C3588 vdd.n1533 gnd 0.008187f
C3589 vdd.n1534 gnd 0.010172f
C3590 vdd.n1535 gnd 1.0395f
C3591 vdd.n1536 gnd 0.010172f
C3592 vdd.n1537 gnd 0.008187f
C3593 vdd.n1538 gnd 0.008187f
C3594 vdd.n1539 gnd 0.010172f
C3595 vdd.n1540 gnd 0.008187f
C3596 vdd.n1541 gnd 0.010172f
C3597 vdd.t130 gnd 0.519752f
C3598 vdd.n1542 gnd 0.010172f
C3599 vdd.n1543 gnd 0.008187f
C3600 vdd.n1544 gnd 0.010172f
C3601 vdd.n1545 gnd 0.008187f
C3602 vdd.n1546 gnd 0.010172f
C3603 vdd.t180 gnd 0.519752f
C3604 vdd.n1547 gnd 0.010172f
C3605 vdd.n1548 gnd 0.008187f
C3606 vdd.n1549 gnd 0.010172f
C3607 vdd.n1550 gnd 0.008187f
C3608 vdd.n1551 gnd 0.010172f
C3609 vdd.n1552 gnd 0.836801f
C3610 vdd.n1553 gnd 0.862789f
C3611 vdd.t184 gnd 0.519752f
C3612 vdd.n1554 gnd 0.010172f
C3613 vdd.n1555 gnd 0.008187f
C3614 vdd.n1556 gnd 0.010172f
C3615 vdd.n1557 gnd 0.008187f
C3616 vdd.n1558 gnd 0.010172f
C3617 vdd.n1559 gnd 0.660085f
C3618 vdd.n1560 gnd 0.010172f
C3619 vdd.n1561 gnd 0.008187f
C3620 vdd.n1562 gnd 0.010172f
C3621 vdd.n1563 gnd 0.008187f
C3622 vdd.n1564 gnd 0.010172f
C3623 vdd.t127 gnd 0.519752f
C3624 vdd.t125 gnd 0.519752f
C3625 vdd.n1565 gnd 0.010172f
C3626 vdd.n1566 gnd 0.008187f
C3627 vdd.n1567 gnd 0.010172f
C3628 vdd.n1568 gnd 0.008187f
C3629 vdd.n1569 gnd 0.010172f
C3630 vdd.t92 gnd 0.519752f
C3631 vdd.n1570 gnd 0.010172f
C3632 vdd.n1571 gnd 0.008187f
C3633 vdd.n1572 gnd 0.010172f
C3634 vdd.n1573 gnd 0.008187f
C3635 vdd.n1574 gnd 0.010172f
C3636 vdd.t96 gnd 0.519752f
C3637 vdd.n1575 gnd 0.732851f
C3638 vdd.n1576 gnd 0.010172f
C3639 vdd.n1577 gnd 0.008187f
C3640 vdd.n1578 gnd 0.010172f
C3641 vdd.n1579 gnd 0.008187f
C3642 vdd.n1580 gnd 0.010172f
C3643 vdd.n1581 gnd 0.816011f
C3644 vdd.n1582 gnd 0.010172f
C3645 vdd.n1583 gnd 0.008187f
C3646 vdd.n1584 gnd 0.010172f
C3647 vdd.n1585 gnd 0.008187f
C3648 vdd.n1586 gnd 0.010172f
C3649 vdd.n1587 gnd 0.639295f
C3650 vdd.t178 gnd 0.519752f
C3651 vdd.n1588 gnd 0.010172f
C3652 vdd.n1589 gnd 0.008187f
C3653 vdd.n1590 gnd 0.010172f
C3654 vdd.n1591 gnd 0.008187f
C3655 vdd.n1592 gnd 0.010172f
C3656 vdd.t136 gnd 0.519752f
C3657 vdd.n1593 gnd 0.010172f
C3658 vdd.n1594 gnd 0.008187f
C3659 vdd.n1595 gnd 0.010172f
C3660 vdd.n1596 gnd 0.008187f
C3661 vdd.n1597 gnd 0.010172f
C3662 vdd.t198 gnd 0.519752f
C3663 vdd.n1598 gnd 0.576925f
C3664 vdd.n1599 gnd 0.010172f
C3665 vdd.n1600 gnd 0.008187f
C3666 vdd.n1601 gnd 0.010172f
C3667 vdd.n1602 gnd 0.008187f
C3668 vdd.n1603 gnd 0.010172f
C3669 vdd.t164 gnd 0.519752f
C3670 vdd.n1604 gnd 0.010172f
C3671 vdd.n1605 gnd 0.008187f
C3672 vdd.n1606 gnd 0.010172f
C3673 vdd.n1607 gnd 0.008187f
C3674 vdd.n1608 gnd 0.010172f
C3675 vdd.n1609 gnd 0.795221f
C3676 vdd.n1610 gnd 0.862789f
C3677 vdd.t132 gnd 0.519752f
C3678 vdd.n1611 gnd 0.010172f
C3679 vdd.n1612 gnd 0.008187f
C3680 vdd.n1613 gnd 0.010172f
C3681 vdd.n1614 gnd 0.008187f
C3682 vdd.n1615 gnd 0.010172f
C3683 vdd.n1616 gnd 0.618505f
C3684 vdd.n1617 gnd 0.010172f
C3685 vdd.n1618 gnd 0.008187f
C3686 vdd.n1619 gnd 0.010172f
C3687 vdd.n1620 gnd 0.008187f
C3688 vdd.n1621 gnd 0.010172f
C3689 vdd.t120 gnd 0.519752f
C3690 vdd.t217 gnd 0.519752f
C3691 vdd.n1622 gnd 0.010172f
C3692 vdd.n1623 gnd 0.008187f
C3693 vdd.n1624 gnd 0.010172f
C3694 vdd.n1625 gnd 0.008187f
C3695 vdd.n1626 gnd 0.010172f
C3696 vdd.t172 gnd 0.519752f
C3697 vdd.n1627 gnd 0.010172f
C3698 vdd.n1628 gnd 0.008187f
C3699 vdd.n1629 gnd 0.010172f
C3700 vdd.n1630 gnd 0.008187f
C3701 vdd.n1631 gnd 0.010172f
C3702 vdd.t175 gnd 0.519752f
C3703 vdd.n1632 gnd 0.774431f
C3704 vdd.n1633 gnd 0.010172f
C3705 vdd.n1634 gnd 0.008187f
C3706 vdd.n1635 gnd 0.010172f
C3707 vdd.n1636 gnd 0.008187f
C3708 vdd.n1637 gnd 0.010172f
C3709 vdd.n1638 gnd 1.0395f
C3710 vdd.n1639 gnd 0.010172f
C3711 vdd.n1640 gnd 0.008187f
C3712 vdd.n1641 gnd 0.024606f
C3713 vdd.n1642 gnd 0.006795f
C3714 vdd.n1643 gnd 0.024606f
C3715 vdd.t72 gnd 0.519752f
C3716 vdd.n1644 gnd 0.024606f
C3717 vdd.n1645 gnd 0.006795f
C3718 vdd.n1646 gnd 0.010172f
C3719 vdd.n1647 gnd 0.008187f
C3720 vdd.n1648 gnd 0.010172f
C3721 vdd.n1679 gnd 0.025134f
C3722 vdd.n1680 gnd 1.53327f
C3723 vdd.n1681 gnd 0.010172f
C3724 vdd.n1682 gnd 0.008187f
C3725 vdd.n1683 gnd 0.010172f
C3726 vdd.n1684 gnd 0.010172f
C3727 vdd.n1685 gnd 0.010172f
C3728 vdd.n1686 gnd 0.010172f
C3729 vdd.n1687 gnd 0.010172f
C3730 vdd.n1688 gnd 0.008187f
C3731 vdd.n1689 gnd 0.010172f
C3732 vdd.n1690 gnd 0.010172f
C3733 vdd.n1691 gnd 0.010172f
C3734 vdd.n1692 gnd 0.010172f
C3735 vdd.n1693 gnd 0.010172f
C3736 vdd.n1694 gnd 0.008187f
C3737 vdd.n1695 gnd 0.010172f
C3738 vdd.n1696 gnd 0.010172f
C3739 vdd.n1697 gnd 0.010172f
C3740 vdd.n1698 gnd 0.010172f
C3741 vdd.n1699 gnd 0.010172f
C3742 vdd.n1700 gnd 0.008187f
C3743 vdd.n1701 gnd 0.010172f
C3744 vdd.n1702 gnd 0.010172f
C3745 vdd.n1703 gnd 0.010172f
C3746 vdd.n1704 gnd 0.010172f
C3747 vdd.n1705 gnd 0.010172f
C3748 vdd.t82 gnd 0.125139f
C3749 vdd.t83 gnd 0.133739f
C3750 vdd.t81 gnd 0.16343f
C3751 vdd.n1706 gnd 0.209494f
C3752 vdd.n1707 gnd 0.176832f
C3753 vdd.n1708 gnd 0.01752f
C3754 vdd.n1709 gnd 0.010172f
C3755 vdd.n1710 gnd 0.010172f
C3756 vdd.n1711 gnd 0.010172f
C3757 vdd.n1712 gnd 0.010172f
C3758 vdd.n1713 gnd 0.010172f
C3759 vdd.n1714 gnd 0.008187f
C3760 vdd.n1715 gnd 0.010172f
C3761 vdd.n1716 gnd 0.010172f
C3762 vdd.n1717 gnd 0.010172f
C3763 vdd.n1718 gnd 0.010172f
C3764 vdd.n1719 gnd 0.010172f
C3765 vdd.n1720 gnd 0.008187f
C3766 vdd.n1721 gnd 0.010172f
C3767 vdd.n1722 gnd 0.010172f
C3768 vdd.n1723 gnd 0.010172f
C3769 vdd.n1724 gnd 0.010172f
C3770 vdd.n1725 gnd 0.010172f
C3771 vdd.n1726 gnd 0.008187f
C3772 vdd.n1727 gnd 0.010172f
C3773 vdd.n1728 gnd 0.010172f
C3774 vdd.n1729 gnd 0.010172f
C3775 vdd.n1730 gnd 0.010172f
C3776 vdd.n1731 gnd 0.010172f
C3777 vdd.n1732 gnd 0.008187f
C3778 vdd.n1733 gnd 0.010172f
C3779 vdd.n1734 gnd 0.010172f
C3780 vdd.n1735 gnd 0.010172f
C3781 vdd.n1736 gnd 0.010172f
C3782 vdd.n1737 gnd 0.010172f
C3783 vdd.n1738 gnd 0.008187f
C3784 vdd.n1739 gnd 0.010172f
C3785 vdd.n1740 gnd 0.010172f
C3786 vdd.n1741 gnd 0.010172f
C3787 vdd.n1742 gnd 0.010172f
C3788 vdd.n1743 gnd 0.008187f
C3789 vdd.n1744 gnd 0.010172f
C3790 vdd.n1745 gnd 0.010172f
C3791 vdd.n1746 gnd 0.010172f
C3792 vdd.n1747 gnd 0.010172f
C3793 vdd.n1748 gnd 0.010172f
C3794 vdd.n1749 gnd 0.008187f
C3795 vdd.n1750 gnd 0.010172f
C3796 vdd.n1751 gnd 0.010172f
C3797 vdd.n1752 gnd 0.010172f
C3798 vdd.n1753 gnd 0.010172f
C3799 vdd.n1754 gnd 0.010172f
C3800 vdd.n1755 gnd 0.008187f
C3801 vdd.n1756 gnd 0.010172f
C3802 vdd.n1757 gnd 0.010172f
C3803 vdd.n1758 gnd 0.010172f
C3804 vdd.n1759 gnd 0.010172f
C3805 vdd.n1760 gnd 0.010172f
C3806 vdd.n1761 gnd 0.008187f
C3807 vdd.n1762 gnd 0.010172f
C3808 vdd.n1763 gnd 0.010172f
C3809 vdd.n1764 gnd 0.010172f
C3810 vdd.n1765 gnd 0.010172f
C3811 vdd.n1766 gnd 0.010172f
C3812 vdd.n1767 gnd 0.008187f
C3813 vdd.n1768 gnd 0.010172f
C3814 vdd.n1769 gnd 0.010172f
C3815 vdd.n1770 gnd 0.010172f
C3816 vdd.n1771 gnd 0.010172f
C3817 vdd.t79 gnd 0.125139f
C3818 vdd.t80 gnd 0.133739f
C3819 vdd.t78 gnd 0.16343f
C3820 vdd.n1772 gnd 0.209494f
C3821 vdd.n1773 gnd 0.176832f
C3822 vdd.n1774 gnd 0.013427f
C3823 vdd.n1775 gnd 0.003889f
C3824 vdd.n1776 gnd 0.025134f
C3825 vdd.n1777 gnd 0.010172f
C3826 vdd.n1778 gnd 0.004298f
C3827 vdd.n1779 gnd 0.008187f
C3828 vdd.n1780 gnd 0.008187f
C3829 vdd.n1781 gnd 0.010172f
C3830 vdd.n1782 gnd 0.010172f
C3831 vdd.n1783 gnd 0.010172f
C3832 vdd.n1784 gnd 0.008187f
C3833 vdd.n1785 gnd 0.008187f
C3834 vdd.n1786 gnd 0.008187f
C3835 vdd.n1787 gnd 0.010172f
C3836 vdd.n1788 gnd 0.010172f
C3837 vdd.n1789 gnd 0.010172f
C3838 vdd.n1790 gnd 0.008187f
C3839 vdd.n1791 gnd 0.008187f
C3840 vdd.n1792 gnd 0.008187f
C3841 vdd.n1793 gnd 0.010172f
C3842 vdd.n1794 gnd 0.010172f
C3843 vdd.n1795 gnd 0.010172f
C3844 vdd.n1796 gnd 0.008187f
C3845 vdd.n1797 gnd 0.008187f
C3846 vdd.n1798 gnd 0.008187f
C3847 vdd.n1799 gnd 0.010172f
C3848 vdd.n1800 gnd 0.010172f
C3849 vdd.n1801 gnd 0.010172f
C3850 vdd.n1802 gnd 0.008187f
C3851 vdd.n1803 gnd 0.008187f
C3852 vdd.n1804 gnd 0.008187f
C3853 vdd.n1805 gnd 0.010172f
C3854 vdd.n1806 gnd 0.010172f
C3855 vdd.n1807 gnd 0.010172f
C3856 vdd.n1808 gnd 0.008105f
C3857 vdd.n1809 gnd 0.010172f
C3858 vdd.t73 gnd 0.125139f
C3859 vdd.t74 gnd 0.133739f
C3860 vdd.t71 gnd 0.16343f
C3861 vdd.n1810 gnd 0.209494f
C3862 vdd.n1811 gnd 0.176832f
C3863 vdd.n1812 gnd 0.01752f
C3864 vdd.n1813 gnd 0.005567f
C3865 vdd.n1814 gnd 0.010172f
C3866 vdd.n1815 gnd 0.010172f
C3867 vdd.n1816 gnd 0.010172f
C3868 vdd.n1817 gnd 0.008187f
C3869 vdd.n1818 gnd 0.008187f
C3870 vdd.n1819 gnd 0.008187f
C3871 vdd.n1820 gnd 0.010172f
C3872 vdd.n1821 gnd 0.010172f
C3873 vdd.n1822 gnd 0.010172f
C3874 vdd.n1823 gnd 0.008187f
C3875 vdd.n1824 gnd 0.008187f
C3876 vdd.n1825 gnd 0.008187f
C3877 vdd.n1826 gnd 0.010172f
C3878 vdd.n1827 gnd 0.010172f
C3879 vdd.n1828 gnd 0.010172f
C3880 vdd.n1829 gnd 0.008187f
C3881 vdd.n1830 gnd 0.008187f
C3882 vdd.n1831 gnd 0.008187f
C3883 vdd.n1832 gnd 0.010172f
C3884 vdd.n1833 gnd 0.010172f
C3885 vdd.n1834 gnd 0.010172f
C3886 vdd.n1835 gnd 0.008187f
C3887 vdd.n1836 gnd 0.008187f
C3888 vdd.n1837 gnd 0.008187f
C3889 vdd.n1838 gnd 0.010172f
C3890 vdd.n1839 gnd 0.010172f
C3891 vdd.n1840 gnd 0.010172f
C3892 vdd.n1841 gnd 0.008187f
C3893 vdd.n1842 gnd 0.008187f
C3894 vdd.n1843 gnd 0.006836f
C3895 vdd.n1844 gnd 0.010172f
C3896 vdd.n1845 gnd 0.010172f
C3897 vdd.n1846 gnd 0.010172f
C3898 vdd.n1847 gnd 0.006836f
C3899 vdd.n1848 gnd 0.008187f
C3900 vdd.n1849 gnd 0.008187f
C3901 vdd.n1850 gnd 0.010172f
C3902 vdd.n1851 gnd 0.010172f
C3903 vdd.n1852 gnd 0.010172f
C3904 vdd.n1853 gnd 0.008187f
C3905 vdd.n1854 gnd 0.008187f
C3906 vdd.n1855 gnd 0.008187f
C3907 vdd.n1856 gnd 0.010172f
C3908 vdd.n1857 gnd 0.010172f
C3909 vdd.n1858 gnd 0.010172f
C3910 vdd.n1859 gnd 0.008187f
C3911 vdd.n1860 gnd 0.008187f
C3912 vdd.n1861 gnd 0.008187f
C3913 vdd.n1862 gnd 0.010172f
C3914 vdd.n1863 gnd 0.010172f
C3915 vdd.n1864 gnd 0.010172f
C3916 vdd.n1865 gnd 0.008187f
C3917 vdd.n1866 gnd 0.008187f
C3918 vdd.n1867 gnd 0.008187f
C3919 vdd.n1868 gnd 0.010172f
C3920 vdd.n1869 gnd 0.010172f
C3921 vdd.n1870 gnd 0.010172f
C3922 vdd.n1871 gnd 0.008187f
C3923 vdd.n1872 gnd 0.010172f
C3924 vdd.n1873 gnd 2.46363f
C3925 vdd.n1875 gnd 0.025134f
C3926 vdd.n1876 gnd 0.006795f
C3927 vdd.n1877 gnd 0.025134f
C3928 vdd.n1878 gnd 0.024606f
C3929 vdd.n1879 gnd 0.010172f
C3930 vdd.n1880 gnd 0.008187f
C3931 vdd.n1881 gnd 0.010172f
C3932 vdd.n1882 gnd 0.52495f
C3933 vdd.n1883 gnd 0.010172f
C3934 vdd.n1884 gnd 0.008187f
C3935 vdd.n1885 gnd 0.010172f
C3936 vdd.n1886 gnd 0.010172f
C3937 vdd.n1887 gnd 0.010172f
C3938 vdd.n1888 gnd 0.008187f
C3939 vdd.n1889 gnd 0.010172f
C3940 vdd.n1890 gnd 0.951146f
C3941 vdd.n1891 gnd 1.0395f
C3942 vdd.n1892 gnd 0.010172f
C3943 vdd.n1893 gnd 0.008187f
C3944 vdd.n1894 gnd 0.010172f
C3945 vdd.n1895 gnd 0.010172f
C3946 vdd.n1896 gnd 0.010172f
C3947 vdd.n1897 gnd 0.008187f
C3948 vdd.n1898 gnd 0.010172f
C3949 vdd.n1899 gnd 0.60811f
C3950 vdd.n1900 gnd 0.010172f
C3951 vdd.n1901 gnd 0.008187f
C3952 vdd.n1902 gnd 0.010172f
C3953 vdd.n1903 gnd 0.010172f
C3954 vdd.n1904 gnd 0.010172f
C3955 vdd.n1905 gnd 0.008187f
C3956 vdd.n1906 gnd 0.010172f
C3957 vdd.n1907 gnd 0.597715f
C3958 vdd.n1908 gnd 0.784826f
C3959 vdd.n1909 gnd 0.010172f
C3960 vdd.n1910 gnd 0.008187f
C3961 vdd.n1911 gnd 0.010172f
C3962 vdd.n1912 gnd 0.010172f
C3963 vdd.n1913 gnd 0.010172f
C3964 vdd.n1914 gnd 0.008187f
C3965 vdd.n1915 gnd 0.010172f
C3966 vdd.n1916 gnd 0.862789f
C3967 vdd.n1917 gnd 0.010172f
C3968 vdd.n1918 gnd 0.008187f
C3969 vdd.n1919 gnd 0.010172f
C3970 vdd.n1920 gnd 0.010172f
C3971 vdd.n1921 gnd 0.010172f
C3972 vdd.n1922 gnd 0.008187f
C3973 vdd.n1923 gnd 0.010172f
C3974 vdd.t182 gnd 0.519752f
C3975 vdd.n1924 gnd 0.764036f
C3976 vdd.n1925 gnd 0.010172f
C3977 vdd.n1926 gnd 0.008187f
C3978 vdd.n1927 gnd 0.010172f
C3979 vdd.n1928 gnd 0.010172f
C3980 vdd.n1929 gnd 0.010172f
C3981 vdd.n1930 gnd 0.008187f
C3982 vdd.n1931 gnd 0.010172f
C3983 vdd.n1932 gnd 0.58732f
C3984 vdd.n1933 gnd 0.010172f
C3985 vdd.n1934 gnd 0.008187f
C3986 vdd.n1935 gnd 0.010172f
C3987 vdd.n1936 gnd 0.010172f
C3988 vdd.n1937 gnd 0.010172f
C3989 vdd.n1938 gnd 0.008187f
C3990 vdd.n1939 gnd 0.010172f
C3991 vdd.n1940 gnd 0.753641f
C3992 vdd.n1941 gnd 0.6289f
C3993 vdd.n1942 gnd 0.010172f
C3994 vdd.n1943 gnd 0.008187f
C3995 vdd.n1944 gnd 0.010172f
C3996 vdd.n1945 gnd 0.010172f
C3997 vdd.n1946 gnd 0.010172f
C3998 vdd.n1947 gnd 0.008187f
C3999 vdd.n1948 gnd 0.010172f
C4000 vdd.n1949 gnd 0.805616f
C4001 vdd.n1950 gnd 0.010172f
C4002 vdd.n1951 gnd 0.008187f
C4003 vdd.n1952 gnd 0.010172f
C4004 vdd.n1953 gnd 0.010172f
C4005 vdd.n1954 gnd 0.010172f
C4006 vdd.n1955 gnd 0.008187f
C4007 vdd.n1956 gnd 0.010172f
C4008 vdd.t88 gnd 0.519752f
C4009 vdd.n1957 gnd 0.862789f
C4010 vdd.n1958 gnd 0.010172f
C4011 vdd.n1959 gnd 0.008187f
C4012 vdd.n1960 gnd 0.010172f
C4013 vdd.n1961 gnd 0.007818f
C4014 vdd.n1962 gnd 0.005582f
C4015 vdd.n1963 gnd 0.00518f
C4016 vdd.n1964 gnd 0.002865f
C4017 vdd.n1965 gnd 0.006579f
C4018 vdd.n1966 gnd 0.002784f
C4019 vdd.n1967 gnd 0.002947f
C4020 vdd.n1968 gnd 0.00518f
C4021 vdd.n1969 gnd 0.002784f
C4022 vdd.n1970 gnd 0.006579f
C4023 vdd.n1971 gnd 0.002947f
C4024 vdd.n1972 gnd 0.00518f
C4025 vdd.n1973 gnd 0.002784f
C4026 vdd.n1974 gnd 0.004935f
C4027 vdd.n1975 gnd 0.004949f
C4028 vdd.t171 gnd 0.014135f
C4029 vdd.n1976 gnd 0.031451f
C4030 vdd.n1977 gnd 0.163677f
C4031 vdd.n1978 gnd 0.002784f
C4032 vdd.n1979 gnd 0.002947f
C4033 vdd.n1980 gnd 0.006579f
C4034 vdd.n1981 gnd 0.006579f
C4035 vdd.n1982 gnd 0.002947f
C4036 vdd.n1983 gnd 0.002784f
C4037 vdd.n1984 gnd 0.00518f
C4038 vdd.n1985 gnd 0.00518f
C4039 vdd.n1986 gnd 0.002784f
C4040 vdd.n1987 gnd 0.002947f
C4041 vdd.n1988 gnd 0.006579f
C4042 vdd.n1989 gnd 0.006579f
C4043 vdd.n1990 gnd 0.002947f
C4044 vdd.n1991 gnd 0.002784f
C4045 vdd.n1992 gnd 0.00518f
C4046 vdd.n1993 gnd 0.00518f
C4047 vdd.n1994 gnd 0.002784f
C4048 vdd.n1995 gnd 0.002947f
C4049 vdd.n1996 gnd 0.006579f
C4050 vdd.n1997 gnd 0.006579f
C4051 vdd.n1998 gnd 0.015555f
C4052 vdd.n1999 gnd 0.002865f
C4053 vdd.n2000 gnd 0.002784f
C4054 vdd.n2001 gnd 0.013389f
C4055 vdd.n2002 gnd 0.009347f
C4056 vdd.t223 gnd 0.032748f
C4057 vdd.t247 gnd 0.032748f
C4058 vdd.n2003 gnd 0.225067f
C4059 vdd.n2004 gnd 0.176981f
C4060 vdd.t202 gnd 0.032748f
C4061 vdd.t115 gnd 0.032748f
C4062 vdd.n2005 gnd 0.225067f
C4063 vdd.n2006 gnd 0.142823f
C4064 vdd.t186 gnd 0.032748f
C4065 vdd.t128 gnd 0.032748f
C4066 vdd.n2007 gnd 0.225067f
C4067 vdd.n2008 gnd 0.142823f
C4068 vdd.t234 gnd 0.032748f
C4069 vdd.t156 gnd 0.032748f
C4070 vdd.n2009 gnd 0.225067f
C4071 vdd.n2010 gnd 0.142823f
C4072 vdd.t208 gnd 0.032748f
C4073 vdd.t179 gnd 0.032748f
C4074 vdd.n2011 gnd 0.225067f
C4075 vdd.n2012 gnd 0.142823f
C4076 vdd.t225 gnd 0.032748f
C4077 vdd.t137 gnd 0.032748f
C4078 vdd.n2013 gnd 0.225067f
C4079 vdd.n2014 gnd 0.142823f
C4080 vdd.t244 gnd 0.032748f
C4081 vdd.t165 gnd 0.032748f
C4082 vdd.n2015 gnd 0.225067f
C4083 vdd.n2016 gnd 0.142823f
C4084 vdd.t218 gnd 0.032748f
C4085 vdd.t191 gnd 0.032748f
C4086 vdd.n2017 gnd 0.225067f
C4087 vdd.n2018 gnd 0.142823f
C4088 vdd.t235 gnd 0.032748f
C4089 vdd.t158 gnd 0.032748f
C4090 vdd.n2019 gnd 0.225067f
C4091 vdd.n2020 gnd 0.142823f
C4092 vdd.n2021 gnd 0.005582f
C4093 vdd.n2022 gnd 0.00518f
C4094 vdd.n2023 gnd 0.002865f
C4095 vdd.n2024 gnd 0.006579f
C4096 vdd.n2025 gnd 0.002784f
C4097 vdd.n2026 gnd 0.002947f
C4098 vdd.n2027 gnd 0.00518f
C4099 vdd.n2028 gnd 0.002784f
C4100 vdd.n2029 gnd 0.006579f
C4101 vdd.n2030 gnd 0.002947f
C4102 vdd.n2031 gnd 0.00518f
C4103 vdd.n2032 gnd 0.002784f
C4104 vdd.n2033 gnd 0.004935f
C4105 vdd.n2034 gnd 0.004949f
C4106 vdd.t212 gnd 0.014135f
C4107 vdd.n2035 gnd 0.031451f
C4108 vdd.n2036 gnd 0.163677f
C4109 vdd.n2037 gnd 0.002784f
C4110 vdd.n2038 gnd 0.002947f
C4111 vdd.n2039 gnd 0.006579f
C4112 vdd.n2040 gnd 0.006579f
C4113 vdd.n2041 gnd 0.002947f
C4114 vdd.n2042 gnd 0.002784f
C4115 vdd.n2043 gnd 0.00518f
C4116 vdd.n2044 gnd 0.00518f
C4117 vdd.n2045 gnd 0.002784f
C4118 vdd.n2046 gnd 0.002947f
C4119 vdd.n2047 gnd 0.006579f
C4120 vdd.n2048 gnd 0.006579f
C4121 vdd.n2049 gnd 0.002947f
C4122 vdd.n2050 gnd 0.002784f
C4123 vdd.n2051 gnd 0.00518f
C4124 vdd.n2052 gnd 0.00518f
C4125 vdd.n2053 gnd 0.002784f
C4126 vdd.n2054 gnd 0.002947f
C4127 vdd.n2055 gnd 0.006579f
C4128 vdd.n2056 gnd 0.006579f
C4129 vdd.n2057 gnd 0.015555f
C4130 vdd.n2058 gnd 0.002865f
C4131 vdd.n2059 gnd 0.002784f
C4132 vdd.n2060 gnd 0.013389f
C4133 vdd.n2061 gnd 0.009054f
C4134 vdd.n2062 gnd 0.106261f
C4135 vdd.n2063 gnd 0.005582f
C4136 vdd.n2064 gnd 0.00518f
C4137 vdd.n2065 gnd 0.002865f
C4138 vdd.n2066 gnd 0.006579f
C4139 vdd.n2067 gnd 0.002784f
C4140 vdd.n2068 gnd 0.002947f
C4141 vdd.n2069 gnd 0.00518f
C4142 vdd.n2070 gnd 0.002784f
C4143 vdd.n2071 gnd 0.006579f
C4144 vdd.n2072 gnd 0.002947f
C4145 vdd.n2073 gnd 0.00518f
C4146 vdd.n2074 gnd 0.002784f
C4147 vdd.n2075 gnd 0.004935f
C4148 vdd.n2076 gnd 0.004949f
C4149 vdd.t131 gnd 0.014135f
C4150 vdd.n2077 gnd 0.031451f
C4151 vdd.n2078 gnd 0.163677f
C4152 vdd.n2079 gnd 0.002784f
C4153 vdd.n2080 gnd 0.002947f
C4154 vdd.n2081 gnd 0.006579f
C4155 vdd.n2082 gnd 0.006579f
C4156 vdd.n2083 gnd 0.002947f
C4157 vdd.n2084 gnd 0.002784f
C4158 vdd.n2085 gnd 0.00518f
C4159 vdd.n2086 gnd 0.00518f
C4160 vdd.n2087 gnd 0.002784f
C4161 vdd.n2088 gnd 0.002947f
C4162 vdd.n2089 gnd 0.006579f
C4163 vdd.n2090 gnd 0.006579f
C4164 vdd.n2091 gnd 0.002947f
C4165 vdd.n2092 gnd 0.002784f
C4166 vdd.n2093 gnd 0.00518f
C4167 vdd.n2094 gnd 0.00518f
C4168 vdd.n2095 gnd 0.002784f
C4169 vdd.n2096 gnd 0.002947f
C4170 vdd.n2097 gnd 0.006579f
C4171 vdd.n2098 gnd 0.006579f
C4172 vdd.n2099 gnd 0.015555f
C4173 vdd.n2100 gnd 0.002865f
C4174 vdd.n2101 gnd 0.002784f
C4175 vdd.n2102 gnd 0.013389f
C4176 vdd.n2103 gnd 0.009347f
C4177 vdd.t185 gnd 0.032748f
C4178 vdd.t181 gnd 0.032748f
C4179 vdd.n2104 gnd 0.225067f
C4180 vdd.n2105 gnd 0.176981f
C4181 vdd.t126 gnd 0.032748f
C4182 vdd.t99 gnd 0.032748f
C4183 vdd.n2106 gnd 0.225067f
C4184 vdd.n2107 gnd 0.142823f
C4185 vdd.t93 gnd 0.032748f
C4186 vdd.t174 gnd 0.032748f
C4187 vdd.n2108 gnd 0.225067f
C4188 vdd.n2109 gnd 0.142823f
C4189 vdd.t149 gnd 0.032748f
C4190 vdd.t97 gnd 0.032748f
C4191 vdd.n2110 gnd 0.225067f
C4192 vdd.n2111 gnd 0.142823f
C4193 vdd.t89 gnd 0.032748f
C4194 vdd.t204 gnd 0.032748f
C4195 vdd.n2112 gnd 0.225067f
C4196 vdd.n2113 gnd 0.142823f
C4197 vdd.t199 gnd 0.032748f
C4198 vdd.t143 gnd 0.032748f
C4199 vdd.n2114 gnd 0.225067f
C4200 vdd.n2115 gnd 0.142823f
C4201 vdd.t133 gnd 0.032748f
C4202 vdd.t231 gnd 0.032748f
C4203 vdd.n2116 gnd 0.225067f
C4204 vdd.n2117 gnd 0.142823f
C4205 vdd.t226 gnd 0.032748f
C4206 vdd.t183 gnd 0.032748f
C4207 vdd.n2118 gnd 0.225067f
C4208 vdd.n2119 gnd 0.142823f
C4209 vdd.t173 gnd 0.032748f
C4210 vdd.t121 gnd 0.032748f
C4211 vdd.n2120 gnd 0.225067f
C4212 vdd.n2121 gnd 0.142823f
C4213 vdd.n2122 gnd 0.005582f
C4214 vdd.n2123 gnd 0.00518f
C4215 vdd.n2124 gnd 0.002865f
C4216 vdd.n2125 gnd 0.006579f
C4217 vdd.n2126 gnd 0.002784f
C4218 vdd.n2127 gnd 0.002947f
C4219 vdd.n2128 gnd 0.00518f
C4220 vdd.n2129 gnd 0.002784f
C4221 vdd.n2130 gnd 0.006579f
C4222 vdd.n2131 gnd 0.002947f
C4223 vdd.n2132 gnd 0.00518f
C4224 vdd.n2133 gnd 0.002784f
C4225 vdd.n2134 gnd 0.004935f
C4226 vdd.n2135 gnd 0.004949f
C4227 vdd.t176 gnd 0.014135f
C4228 vdd.n2136 gnd 0.031451f
C4229 vdd.n2137 gnd 0.163677f
C4230 vdd.n2138 gnd 0.002784f
C4231 vdd.n2139 gnd 0.002947f
C4232 vdd.n2140 gnd 0.006579f
C4233 vdd.n2141 gnd 0.006579f
C4234 vdd.n2142 gnd 0.002947f
C4235 vdd.n2143 gnd 0.002784f
C4236 vdd.n2144 gnd 0.00518f
C4237 vdd.n2145 gnd 0.00518f
C4238 vdd.n2146 gnd 0.002784f
C4239 vdd.n2147 gnd 0.002947f
C4240 vdd.n2148 gnd 0.006579f
C4241 vdd.n2149 gnd 0.006579f
C4242 vdd.n2150 gnd 0.002947f
C4243 vdd.n2151 gnd 0.002784f
C4244 vdd.n2152 gnd 0.00518f
C4245 vdd.n2153 gnd 0.00518f
C4246 vdd.n2154 gnd 0.002784f
C4247 vdd.n2155 gnd 0.002947f
C4248 vdd.n2156 gnd 0.006579f
C4249 vdd.n2157 gnd 0.006579f
C4250 vdd.n2158 gnd 0.015555f
C4251 vdd.n2159 gnd 0.002865f
C4252 vdd.n2160 gnd 0.002784f
C4253 vdd.n2161 gnd 0.013389f
C4254 vdd.n2162 gnd 0.009054f
C4255 vdd.n2163 gnd 0.063214f
C4256 vdd.n2164 gnd 0.227778f
C4257 vdd.n2165 gnd 0.005582f
C4258 vdd.n2166 gnd 0.00518f
C4259 vdd.n2167 gnd 0.002865f
C4260 vdd.n2168 gnd 0.006579f
C4261 vdd.n2169 gnd 0.002784f
C4262 vdd.n2170 gnd 0.002947f
C4263 vdd.n2171 gnd 0.00518f
C4264 vdd.n2172 gnd 0.002784f
C4265 vdd.n2173 gnd 0.006579f
C4266 vdd.n2174 gnd 0.002947f
C4267 vdd.n2175 gnd 0.00518f
C4268 vdd.n2176 gnd 0.002784f
C4269 vdd.n2177 gnd 0.004935f
C4270 vdd.n2178 gnd 0.004949f
C4271 vdd.t151 gnd 0.014135f
C4272 vdd.n2179 gnd 0.031451f
C4273 vdd.n2180 gnd 0.163677f
C4274 vdd.n2181 gnd 0.002784f
C4275 vdd.n2182 gnd 0.002947f
C4276 vdd.n2183 gnd 0.006579f
C4277 vdd.n2184 gnd 0.006579f
C4278 vdd.n2185 gnd 0.002947f
C4279 vdd.n2186 gnd 0.002784f
C4280 vdd.n2187 gnd 0.00518f
C4281 vdd.n2188 gnd 0.00518f
C4282 vdd.n2189 gnd 0.002784f
C4283 vdd.n2190 gnd 0.002947f
C4284 vdd.n2191 gnd 0.006579f
C4285 vdd.n2192 gnd 0.006579f
C4286 vdd.n2193 gnd 0.002947f
C4287 vdd.n2194 gnd 0.002784f
C4288 vdd.n2195 gnd 0.00518f
C4289 vdd.n2196 gnd 0.00518f
C4290 vdd.n2197 gnd 0.002784f
C4291 vdd.n2198 gnd 0.002947f
C4292 vdd.n2199 gnd 0.006579f
C4293 vdd.n2200 gnd 0.006579f
C4294 vdd.n2201 gnd 0.015555f
C4295 vdd.n2202 gnd 0.002865f
C4296 vdd.n2203 gnd 0.002784f
C4297 vdd.n2204 gnd 0.013389f
C4298 vdd.n2205 gnd 0.009347f
C4299 vdd.t196 gnd 0.032748f
C4300 vdd.t195 gnd 0.032748f
C4301 vdd.n2206 gnd 0.225067f
C4302 vdd.n2207 gnd 0.176981f
C4303 vdd.t147 gnd 0.032748f
C4304 vdd.t118 gnd 0.032748f
C4305 vdd.n2208 gnd 0.225067f
C4306 vdd.n2209 gnd 0.142823f
C4307 vdd.t116 gnd 0.032748f
C4308 vdd.t187 gnd 0.032748f
C4309 vdd.n2210 gnd 0.225067f
C4310 vdd.n2211 gnd 0.142823f
C4311 vdd.t166 gnd 0.032748f
C4312 vdd.t117 gnd 0.032748f
C4313 vdd.n2212 gnd 0.225067f
C4314 vdd.n2213 gnd 0.142823f
C4315 vdd.t112 gnd 0.032748f
C4316 vdd.t214 gnd 0.032748f
C4317 vdd.n2214 gnd 0.225067f
C4318 vdd.n2215 gnd 0.142823f
C4319 vdd.t211 gnd 0.032748f
C4320 vdd.t160 gnd 0.032748f
C4321 vdd.n2216 gnd 0.225067f
C4322 vdd.n2217 gnd 0.142823f
C4323 vdd.t150 gnd 0.032748f
C4324 vdd.t245 gnd 0.032748f
C4325 vdd.n2218 gnd 0.225067f
C4326 vdd.n2219 gnd 0.142823f
C4327 vdd.t239 gnd 0.032748f
C4328 vdd.t194 gnd 0.032748f
C4329 vdd.n2220 gnd 0.225067f
C4330 vdd.n2221 gnd 0.142823f
C4331 vdd.t192 gnd 0.032748f
C4332 vdd.t146 gnd 0.032748f
C4333 vdd.n2222 gnd 0.225067f
C4334 vdd.n2223 gnd 0.142823f
C4335 vdd.n2224 gnd 0.005582f
C4336 vdd.n2225 gnd 0.00518f
C4337 vdd.n2226 gnd 0.002865f
C4338 vdd.n2227 gnd 0.006579f
C4339 vdd.n2228 gnd 0.002784f
C4340 vdd.n2229 gnd 0.002947f
C4341 vdd.n2230 gnd 0.00518f
C4342 vdd.n2231 gnd 0.002784f
C4343 vdd.n2232 gnd 0.006579f
C4344 vdd.n2233 gnd 0.002947f
C4345 vdd.n2234 gnd 0.00518f
C4346 vdd.n2235 gnd 0.002784f
C4347 vdd.n2236 gnd 0.004935f
C4348 vdd.n2237 gnd 0.004949f
C4349 vdd.t193 gnd 0.014135f
C4350 vdd.n2238 gnd 0.031451f
C4351 vdd.n2239 gnd 0.163677f
C4352 vdd.n2240 gnd 0.002784f
C4353 vdd.n2241 gnd 0.002947f
C4354 vdd.n2242 gnd 0.006579f
C4355 vdd.n2243 gnd 0.006579f
C4356 vdd.n2244 gnd 0.002947f
C4357 vdd.n2245 gnd 0.002784f
C4358 vdd.n2246 gnd 0.00518f
C4359 vdd.n2247 gnd 0.00518f
C4360 vdd.n2248 gnd 0.002784f
C4361 vdd.n2249 gnd 0.002947f
C4362 vdd.n2250 gnd 0.006579f
C4363 vdd.n2251 gnd 0.006579f
C4364 vdd.n2252 gnd 0.002947f
C4365 vdd.n2253 gnd 0.002784f
C4366 vdd.n2254 gnd 0.00518f
C4367 vdd.n2255 gnd 0.00518f
C4368 vdd.n2256 gnd 0.002784f
C4369 vdd.n2257 gnd 0.002947f
C4370 vdd.n2258 gnd 0.006579f
C4371 vdd.n2259 gnd 0.006579f
C4372 vdd.n2260 gnd 0.015555f
C4373 vdd.n2261 gnd 0.002865f
C4374 vdd.n2262 gnd 0.002784f
C4375 vdd.n2263 gnd 0.013389f
C4376 vdd.n2264 gnd 0.009054f
C4377 vdd.n2265 gnd 0.063214f
C4378 vdd.n2266 gnd 0.260757f
C4379 vdd.n2267 gnd 2.98161f
C4380 vdd.n2268 gnd 0.599968f
C4381 vdd.n2269 gnd 0.007818f
C4382 vdd.n2270 gnd 0.008187f
C4383 vdd.n2271 gnd 0.010172f
C4384 vdd.n2272 gnd 0.743246f
C4385 vdd.n2273 gnd 0.010172f
C4386 vdd.n2274 gnd 0.008187f
C4387 vdd.n2275 gnd 0.010172f
C4388 vdd.n2276 gnd 0.010172f
C4389 vdd.n2277 gnd 0.010172f
C4390 vdd.n2278 gnd 0.008187f
C4391 vdd.n2279 gnd 0.010172f
C4392 vdd.n2280 gnd 0.862789f
C4393 vdd.t148 gnd 0.519752f
C4394 vdd.n2281 gnd 0.56653f
C4395 vdd.n2282 gnd 0.010172f
C4396 vdd.n2283 gnd 0.008187f
C4397 vdd.n2284 gnd 0.010172f
C4398 vdd.n2285 gnd 0.010172f
C4399 vdd.n2286 gnd 0.010172f
C4400 vdd.n2287 gnd 0.008187f
C4401 vdd.n2288 gnd 0.010172f
C4402 vdd.n2289 gnd 0.64969f
C4403 vdd.n2290 gnd 0.010172f
C4404 vdd.n2291 gnd 0.008187f
C4405 vdd.n2292 gnd 0.010172f
C4406 vdd.n2293 gnd 0.010172f
C4407 vdd.n2294 gnd 0.010172f
C4408 vdd.n2295 gnd 0.008187f
C4409 vdd.n2296 gnd 0.010172f
C4410 vdd.n2297 gnd 0.556135f
C4411 vdd.n2298 gnd 0.826406f
C4412 vdd.n2299 gnd 0.010172f
C4413 vdd.n2300 gnd 0.008187f
C4414 vdd.n2301 gnd 0.010172f
C4415 vdd.n2302 gnd 0.010172f
C4416 vdd.n2303 gnd 0.010172f
C4417 vdd.n2304 gnd 0.008187f
C4418 vdd.n2305 gnd 0.010172f
C4419 vdd.n2306 gnd 0.862789f
C4420 vdd.n2307 gnd 0.010172f
C4421 vdd.n2308 gnd 0.008187f
C4422 vdd.n2309 gnd 0.010172f
C4423 vdd.n2310 gnd 0.010172f
C4424 vdd.n2311 gnd 0.010172f
C4425 vdd.n2312 gnd 0.008187f
C4426 vdd.n2313 gnd 0.010172f
C4427 vdd.t98 gnd 0.519752f
C4428 vdd.n2314 gnd 0.722456f
C4429 vdd.n2315 gnd 0.010172f
C4430 vdd.n2316 gnd 0.008187f
C4431 vdd.n2317 gnd 0.010172f
C4432 vdd.n2318 gnd 0.010172f
C4433 vdd.n2319 gnd 0.010172f
C4434 vdd.n2320 gnd 0.008187f
C4435 vdd.n2321 gnd 0.010172f
C4436 vdd.n2322 gnd 0.54574f
C4437 vdd.n2323 gnd 0.010172f
C4438 vdd.n2324 gnd 0.008187f
C4439 vdd.n2325 gnd 0.010172f
C4440 vdd.n2326 gnd 0.010172f
C4441 vdd.n2327 gnd 0.010172f
C4442 vdd.n2328 gnd 0.008187f
C4443 vdd.n2329 gnd 0.010172f
C4444 vdd.n2330 gnd 0.71206f
C4445 vdd.n2331 gnd 0.67048f
C4446 vdd.n2332 gnd 0.010172f
C4447 vdd.n2333 gnd 0.008187f
C4448 vdd.n2334 gnd 0.010172f
C4449 vdd.n2335 gnd 0.010172f
C4450 vdd.n2336 gnd 0.010172f
C4451 vdd.n2337 gnd 0.008187f
C4452 vdd.n2338 gnd 0.010172f
C4453 vdd.n2339 gnd 0.847196f
C4454 vdd.n2340 gnd 0.010172f
C4455 vdd.n2341 gnd 0.008187f
C4456 vdd.n2342 gnd 0.010172f
C4457 vdd.n2343 gnd 0.010172f
C4458 vdd.n2344 gnd 0.024606f
C4459 vdd.n2345 gnd 0.010172f
C4460 vdd.n2346 gnd 0.010172f
C4461 vdd.n2347 gnd 0.008187f
C4462 vdd.n2348 gnd 0.010172f
C4463 vdd.n2349 gnd 0.6289f
C4464 vdd.n2350 gnd 1.0395f
C4465 vdd.n2351 gnd 0.010172f
C4466 vdd.n2352 gnd 0.008187f
C4467 vdd.n2353 gnd 0.010172f
C4468 vdd.n2354 gnd 0.010172f
C4469 vdd.n2355 gnd 0.024606f
C4470 vdd.n2356 gnd 0.006795f
C4471 vdd.n2357 gnd 0.024606f
C4472 vdd.n2358 gnd 1.42932f
C4473 vdd.n2359 gnd 0.024606f
C4474 vdd.n2360 gnd 0.025134f
C4475 vdd.n2361 gnd 0.003889f
C4476 vdd.t43 gnd 0.125139f
C4477 vdd.t42 gnd 0.133739f
C4478 vdd.t41 gnd 0.16343f
C4479 vdd.n2362 gnd 0.209494f
C4480 vdd.n2363 gnd 0.176013f
C4481 vdd.n2364 gnd 0.012608f
C4482 vdd.n2365 gnd 0.004298f
C4483 vdd.n2366 gnd 0.008748f
C4484 vdd.n2367 gnd 1.07984f
C4485 vdd.n2369 gnd 0.008187f
C4486 vdd.n2370 gnd 0.008187f
C4487 vdd.n2371 gnd 0.010172f
C4488 vdd.n2373 gnd 0.010172f
C4489 vdd.n2374 gnd 0.010172f
C4490 vdd.n2375 gnd 0.008187f
C4491 vdd.n2376 gnd 0.008187f
C4492 vdd.n2377 gnd 0.008187f
C4493 vdd.n2378 gnd 0.010172f
C4494 vdd.n2380 gnd 0.010172f
C4495 vdd.n2381 gnd 0.010172f
C4496 vdd.n2382 gnd 0.008187f
C4497 vdd.n2383 gnd 0.008187f
C4498 vdd.n2384 gnd 0.008187f
C4499 vdd.n2385 gnd 0.010172f
C4500 vdd.n2387 gnd 0.010172f
C4501 vdd.n2388 gnd 0.010172f
C4502 vdd.n2389 gnd 0.008187f
C4503 vdd.n2390 gnd 0.008187f
C4504 vdd.n2391 gnd 0.008187f
C4505 vdd.n2392 gnd 0.010172f
C4506 vdd.n2394 gnd 0.010172f
C4507 vdd.n2395 gnd 0.010172f
C4508 vdd.n2396 gnd 0.008187f
C4509 vdd.n2397 gnd 0.010172f
C4510 vdd.n2398 gnd 0.010172f
C4511 vdd.n2399 gnd 0.010172f
C4512 vdd.n2400 gnd 0.016701f
C4513 vdd.n2401 gnd 0.005567f
C4514 vdd.n2402 gnd 0.008187f
C4515 vdd.n2403 gnd 0.010172f
C4516 vdd.n2405 gnd 0.010172f
C4517 vdd.n2406 gnd 0.010172f
C4518 vdd.n2407 gnd 0.008187f
C4519 vdd.n2408 gnd 0.008187f
C4520 vdd.n2409 gnd 0.008187f
C4521 vdd.n2410 gnd 0.010172f
C4522 vdd.n2412 gnd 0.010172f
C4523 vdd.n2413 gnd 0.010172f
C4524 vdd.n2414 gnd 0.008187f
C4525 vdd.n2415 gnd 0.008187f
C4526 vdd.n2416 gnd 0.008187f
C4527 vdd.n2417 gnd 0.010172f
C4528 vdd.n2419 gnd 0.010172f
C4529 vdd.n2420 gnd 0.010172f
C4530 vdd.n2421 gnd 0.008187f
C4531 vdd.n2422 gnd 0.008187f
C4532 vdd.n2423 gnd 0.008187f
C4533 vdd.n2424 gnd 0.010172f
C4534 vdd.n2426 gnd 0.010172f
C4535 vdd.n2427 gnd 0.010172f
C4536 vdd.n2428 gnd 0.008187f
C4537 vdd.n2429 gnd 0.008187f
C4538 vdd.n2430 gnd 0.008187f
C4539 vdd.n2431 gnd 0.010172f
C4540 vdd.n2433 gnd 0.010172f
C4541 vdd.n2434 gnd 0.010172f
C4542 vdd.n2435 gnd 0.008187f
C4543 vdd.n2436 gnd 0.010172f
C4544 vdd.n2437 gnd 0.010172f
C4545 vdd.n2438 gnd 0.010172f
C4546 vdd.n2439 gnd 0.016701f
C4547 vdd.n2440 gnd 0.006836f
C4548 vdd.n2441 gnd 0.008187f
C4549 vdd.n2442 gnd 0.010172f
C4550 vdd.n2444 gnd 0.010172f
C4551 vdd.n2445 gnd 0.010172f
C4552 vdd.n2446 gnd 0.008187f
C4553 vdd.n2447 gnd 0.008187f
C4554 vdd.n2448 gnd 0.008187f
C4555 vdd.n2449 gnd 0.010172f
C4556 vdd.n2451 gnd 0.010172f
C4557 vdd.n2452 gnd 0.010172f
C4558 vdd.n2453 gnd 0.008187f
C4559 vdd.n2454 gnd 0.008187f
C4560 vdd.n2455 gnd 0.008187f
C4561 vdd.n2456 gnd 0.010172f
C4562 vdd.n2458 gnd 0.010172f
C4563 vdd.n2459 gnd 0.010172f
C4564 vdd.n2460 gnd 0.008187f
C4565 vdd.n2461 gnd 0.008187f
C4566 vdd.n2462 gnd 0.008187f
C4567 vdd.n2463 gnd 0.010172f
C4568 vdd.n2465 gnd 0.010172f
C4569 vdd.n2466 gnd 0.008187f
C4570 vdd.n2467 gnd 0.008187f
C4571 vdd.n2468 gnd 0.010172f
C4572 vdd.n2470 gnd 0.010172f
C4573 vdd.n2471 gnd 0.010172f
C4574 vdd.n2472 gnd 0.008187f
C4575 vdd.n2473 gnd 0.008748f
C4576 vdd.n2474 gnd 1.07984f
C4577 vdd.n2475 gnd 0.046595f
C4578 vdd.n2476 gnd 0.006917f
C4579 vdd.n2477 gnd 0.006917f
C4580 vdd.n2478 gnd 0.006917f
C4581 vdd.n2479 gnd 0.006917f
C4582 vdd.n2480 gnd 0.006917f
C4583 vdd.n2481 gnd 0.006917f
C4584 vdd.n2482 gnd 0.006917f
C4585 vdd.n2483 gnd 0.006917f
C4586 vdd.n2484 gnd 0.006917f
C4587 vdd.n2485 gnd 0.006917f
C4588 vdd.n2486 gnd 0.006917f
C4589 vdd.n2487 gnd 0.006917f
C4590 vdd.n2488 gnd 0.006917f
C4591 vdd.n2489 gnd 0.006917f
C4592 vdd.n2490 gnd 0.006917f
C4593 vdd.n2491 gnd 0.006917f
C4594 vdd.n2492 gnd 0.006917f
C4595 vdd.n2493 gnd 0.006917f
C4596 vdd.n2494 gnd 0.006917f
C4597 vdd.n2495 gnd 0.006917f
C4598 vdd.n2496 gnd 0.006917f
C4599 vdd.n2497 gnd 0.006917f
C4600 vdd.n2498 gnd 0.006917f
C4601 vdd.n2499 gnd 0.006917f
C4602 vdd.n2500 gnd 0.006917f
C4603 vdd.n2501 gnd 0.006917f
C4604 vdd.n2502 gnd 0.006917f
C4605 vdd.n2503 gnd 0.006917f
C4606 vdd.n2504 gnd 0.006917f
C4607 vdd.n2505 gnd 0.006917f
C4608 vdd.n2506 gnd 12.2765f
C4609 vdd.n2508 gnd 0.015705f
C4610 vdd.n2509 gnd 0.015705f
C4611 vdd.n2510 gnd 0.01481f
C4612 vdd.n2511 gnd 0.006917f
C4613 vdd.n2512 gnd 0.006917f
C4614 vdd.n2513 gnd 0.706863f
C4615 vdd.n2514 gnd 0.006917f
C4616 vdd.n2515 gnd 0.006917f
C4617 vdd.n2516 gnd 0.006917f
C4618 vdd.n2517 gnd 0.006917f
C4619 vdd.n2518 gnd 0.006917f
C4620 vdd.n2519 gnd 0.556135f
C4621 vdd.n2520 gnd 0.006917f
C4622 vdd.n2521 gnd 0.006917f
C4623 vdd.n2522 gnd 0.006917f
C4624 vdd.n2523 gnd 0.006917f
C4625 vdd.n2524 gnd 0.006917f
C4626 vdd.n2525 gnd 0.706863f
C4627 vdd.n2526 gnd 0.006917f
C4628 vdd.n2527 gnd 0.006917f
C4629 vdd.n2528 gnd 0.006917f
C4630 vdd.n2529 gnd 0.006917f
C4631 vdd.n2530 gnd 0.006917f
C4632 vdd.n2531 gnd 0.706863f
C4633 vdd.n2532 gnd 0.006917f
C4634 vdd.n2533 gnd 0.006917f
C4635 vdd.n2534 gnd 0.006917f
C4636 vdd.n2535 gnd 0.006917f
C4637 vdd.n2536 gnd 0.006917f
C4638 vdd.n2537 gnd 0.680875f
C4639 vdd.n2538 gnd 0.006917f
C4640 vdd.n2539 gnd 0.006917f
C4641 vdd.n2540 gnd 0.006917f
C4642 vdd.n2541 gnd 0.006917f
C4643 vdd.n2542 gnd 0.006917f
C4644 vdd.n2543 gnd 0.52495f
C4645 vdd.n2544 gnd 0.006917f
C4646 vdd.n2545 gnd 0.006917f
C4647 vdd.n2546 gnd 0.006917f
C4648 vdd.n2547 gnd 0.006917f
C4649 vdd.n2548 gnd 0.006917f
C4650 vdd.n2549 gnd 0.369024f
C4651 vdd.n2550 gnd 0.006917f
C4652 vdd.n2551 gnd 0.006917f
C4653 vdd.n2552 gnd 0.006917f
C4654 vdd.n2553 gnd 0.006917f
C4655 vdd.n2554 gnd 0.006917f
C4656 vdd.n2555 gnd 0.493765f
C4657 vdd.n2556 gnd 0.006917f
C4658 vdd.n2557 gnd 0.006917f
C4659 vdd.n2558 gnd 0.006917f
C4660 vdd.n2559 gnd 0.006917f
C4661 vdd.n2560 gnd 0.006917f
C4662 vdd.n2561 gnd 0.64969f
C4663 vdd.n2562 gnd 0.006917f
C4664 vdd.n2563 gnd 0.006917f
C4665 vdd.n2564 gnd 0.006917f
C4666 vdd.n2565 gnd 0.006917f
C4667 vdd.n2566 gnd 0.006917f
C4668 vdd.n2567 gnd 0.706863f
C4669 vdd.n2568 gnd 0.006917f
C4670 vdd.n2569 gnd 0.006917f
C4671 vdd.n2570 gnd 0.006917f
C4672 vdd.n2571 gnd 0.006917f
C4673 vdd.n2572 gnd 0.006917f
C4674 vdd.n2573 gnd 0.60811f
C4675 vdd.n2574 gnd 0.006917f
C4676 vdd.n2575 gnd 0.006917f
C4677 vdd.n2576 gnd 0.005493f
C4678 vdd.n2577 gnd 0.020037f
C4679 vdd.n2578 gnd 0.004882f
C4680 vdd.n2579 gnd 0.006917f
C4681 vdd.n2580 gnd 0.452184f
C4682 vdd.n2581 gnd 0.006917f
C4683 vdd.n2582 gnd 0.006917f
C4684 vdd.n2583 gnd 0.006917f
C4685 vdd.n2584 gnd 0.006917f
C4686 vdd.n2585 gnd 0.006917f
C4687 vdd.n2586 gnd 0.410604f
C4688 vdd.n2587 gnd 0.006917f
C4689 vdd.n2588 gnd 0.006917f
C4690 vdd.n2589 gnd 0.006917f
C4691 vdd.n2590 gnd 0.006917f
C4692 vdd.n2591 gnd 0.006917f
C4693 vdd.n2592 gnd 0.56653f
C4694 vdd.n2593 gnd 0.006917f
C4695 vdd.n2594 gnd 0.006917f
C4696 vdd.n2595 gnd 0.006917f
C4697 vdd.n2596 gnd 0.006917f
C4698 vdd.n2597 gnd 0.006917f
C4699 vdd.n2598 gnd 0.623703f
C4700 vdd.n2599 gnd 0.006917f
C4701 vdd.n2600 gnd 0.006917f
C4702 vdd.n2601 gnd 0.006917f
C4703 vdd.n2602 gnd 0.006917f
C4704 vdd.n2603 gnd 0.006917f
C4705 vdd.n2604 gnd 0.467777f
C4706 vdd.n2605 gnd 0.006917f
C4707 vdd.n2606 gnd 0.006917f
C4708 vdd.n2607 gnd 0.006917f
C4709 vdd.n2608 gnd 0.006917f
C4710 vdd.n2609 gnd 0.006917f
C4711 vdd.n2610 gnd 0.223493f
C4712 vdd.n2611 gnd 0.006917f
C4713 vdd.n2612 gnd 0.006917f
C4714 vdd.n2613 gnd 0.006917f
C4715 vdd.n2614 gnd 0.006917f
C4716 vdd.n2615 gnd 0.006917f
C4717 vdd.n2616 gnd 0.223493f
C4718 vdd.n2617 gnd 0.006917f
C4719 vdd.n2618 gnd 0.006917f
C4720 vdd.n2619 gnd 0.006917f
C4721 vdd.n2620 gnd 0.006917f
C4722 vdd.n2621 gnd 0.006917f
C4723 vdd.n2622 gnd 0.706863f
C4724 vdd.n2623 gnd 0.006917f
C4725 vdd.n2624 gnd 0.006917f
C4726 vdd.n2625 gnd 0.006917f
C4727 vdd.n2626 gnd 0.006917f
C4728 vdd.n2627 gnd 0.006917f
C4729 vdd.n2628 gnd 0.006917f
C4730 vdd.n2629 gnd 0.006917f
C4731 vdd.n2630 gnd 0.488567f
C4732 vdd.n2631 gnd 0.006917f
C4733 vdd.n2632 gnd 0.006917f
C4734 vdd.n2633 gnd 0.006917f
C4735 vdd.n2634 gnd 0.006917f
C4736 vdd.n2635 gnd 0.006917f
C4737 vdd.n2636 gnd 0.006917f
C4738 vdd.n2637 gnd 0.441789f
C4739 vdd.n2638 gnd 0.006917f
C4740 vdd.n2639 gnd 0.006917f
C4741 vdd.n2640 gnd 0.006917f
C4742 vdd.n2641 gnd 0.015705f
C4743 vdd.n2642 gnd 0.01481f
C4744 vdd.n2643 gnd 0.006917f
C4745 vdd.n2644 gnd 0.006917f
C4746 vdd.n2645 gnd 0.00534f
C4747 vdd.n2646 gnd 0.006917f
C4748 vdd.n2647 gnd 0.006917f
C4749 vdd.n2648 gnd 0.005035f
C4750 vdd.n2649 gnd 0.006917f
C4751 vdd.n2650 gnd 0.006917f
C4752 vdd.n2651 gnd 0.006917f
C4753 vdd.n2652 gnd 0.006917f
C4754 vdd.n2653 gnd 0.006917f
C4755 vdd.n2654 gnd 0.006917f
C4756 vdd.n2655 gnd 0.006917f
C4757 vdd.n2656 gnd 0.006917f
C4758 vdd.n2657 gnd 0.006917f
C4759 vdd.n2658 gnd 0.006917f
C4760 vdd.n2659 gnd 0.006917f
C4761 vdd.n2660 gnd 0.006917f
C4762 vdd.n2661 gnd 0.006917f
C4763 vdd.n2662 gnd 0.006917f
C4764 vdd.n2663 gnd 0.006917f
C4765 vdd.n2664 gnd 0.006917f
C4766 vdd.n2665 gnd 0.006917f
C4767 vdd.n2666 gnd 0.006917f
C4768 vdd.n2667 gnd 0.006917f
C4769 vdd.n2668 gnd 0.006917f
C4770 vdd.n2669 gnd 0.006917f
C4771 vdd.n2670 gnd 0.006917f
C4772 vdd.n2671 gnd 0.006917f
C4773 vdd.n2672 gnd 0.006917f
C4774 vdd.n2673 gnd 0.006917f
C4775 vdd.n2674 gnd 0.006917f
C4776 vdd.n2675 gnd 0.006917f
C4777 vdd.n2676 gnd 0.006917f
C4778 vdd.n2677 gnd 0.006917f
C4779 vdd.n2678 gnd 0.006917f
C4780 vdd.n2679 gnd 0.006917f
C4781 vdd.n2680 gnd 0.006917f
C4782 vdd.n2681 gnd 0.006917f
C4783 vdd.n2682 gnd 0.006917f
C4784 vdd.n2683 gnd 0.006917f
C4785 vdd.n2684 gnd 0.006917f
C4786 vdd.n2685 gnd 0.006917f
C4787 vdd.n2686 gnd 0.006917f
C4788 vdd.n2687 gnd 0.006917f
C4789 vdd.n2688 gnd 0.006917f
C4790 vdd.n2689 gnd 0.006917f
C4791 vdd.n2690 gnd 0.006917f
C4792 vdd.n2691 gnd 0.006917f
C4793 vdd.n2692 gnd 0.006917f
C4794 vdd.n2693 gnd 0.006917f
C4795 vdd.n2694 gnd 0.006917f
C4796 vdd.n2695 gnd 0.006917f
C4797 vdd.n2696 gnd 0.006917f
C4798 vdd.n2697 gnd 0.006917f
C4799 vdd.n2698 gnd 0.006917f
C4800 vdd.n2699 gnd 0.006917f
C4801 vdd.n2700 gnd 0.006917f
C4802 vdd.n2701 gnd 0.006917f
C4803 vdd.n2702 gnd 0.006917f
C4804 vdd.n2703 gnd 0.006917f
C4805 vdd.n2704 gnd 0.006917f
C4806 vdd.n2705 gnd 0.006917f
C4807 vdd.n2706 gnd 0.006917f
C4808 vdd.n2707 gnd 0.006917f
C4809 vdd.n2708 gnd 0.006917f
C4810 vdd.n2709 gnd 0.015705f
C4811 vdd.n2710 gnd 0.01481f
C4812 vdd.n2711 gnd 0.01481f
C4813 vdd.n2712 gnd 0.800418f
C4814 vdd.n2713 gnd 0.01481f
C4815 vdd.n2714 gnd 0.015705f
C4816 vdd.n2715 gnd 0.01481f
C4817 vdd.n2716 gnd 0.006917f
C4818 vdd.n2717 gnd 0.006917f
C4819 vdd.n2718 gnd 0.006917f
C4820 vdd.n2719 gnd 0.00534f
C4821 vdd.n2720 gnd 0.009885f
C4822 vdd.n2721 gnd 0.005035f
C4823 vdd.n2722 gnd 0.006917f
C4824 vdd.n2723 gnd 0.006917f
C4825 vdd.n2724 gnd 0.006917f
C4826 vdd.n2725 gnd 0.006917f
C4827 vdd.n2726 gnd 0.006917f
C4828 vdd.n2727 gnd 0.006917f
C4829 vdd.n2728 gnd 0.006917f
C4830 vdd.n2729 gnd 0.006917f
C4831 vdd.n2730 gnd 0.006917f
C4832 vdd.n2731 gnd 0.006917f
C4833 vdd.n2732 gnd 0.006917f
C4834 vdd.n2733 gnd 0.006917f
C4835 vdd.n2734 gnd 0.006917f
C4836 vdd.n2735 gnd 0.006917f
C4837 vdd.n2736 gnd 0.006917f
C4838 vdd.n2737 gnd 0.006917f
C4839 vdd.n2738 gnd 0.006917f
C4840 vdd.n2739 gnd 0.006917f
C4841 vdd.n2740 gnd 0.006917f
C4842 vdd.n2741 gnd 0.006917f
C4843 vdd.n2742 gnd 0.006917f
C4844 vdd.n2743 gnd 0.006917f
C4845 vdd.n2744 gnd 0.006917f
C4846 vdd.n2745 gnd 0.006917f
C4847 vdd.n2746 gnd 0.006917f
C4848 vdd.n2747 gnd 0.006917f
C4849 vdd.n2748 gnd 0.006917f
C4850 vdd.n2749 gnd 0.006917f
C4851 vdd.n2750 gnd 0.006917f
C4852 vdd.n2751 gnd 0.006917f
C4853 vdd.n2752 gnd 0.006917f
C4854 vdd.n2753 gnd 0.006917f
C4855 vdd.n2754 gnd 0.006917f
C4856 vdd.n2755 gnd 0.006917f
C4857 vdd.n2756 gnd 0.006917f
C4858 vdd.n2757 gnd 0.006917f
C4859 vdd.n2758 gnd 0.006917f
C4860 vdd.n2759 gnd 0.006917f
C4861 vdd.n2760 gnd 0.006917f
C4862 vdd.n2761 gnd 0.006917f
C4863 vdd.n2762 gnd 0.006917f
C4864 vdd.n2763 gnd 0.006917f
C4865 vdd.n2764 gnd 0.006917f
C4866 vdd.n2765 gnd 0.006917f
C4867 vdd.n2766 gnd 0.006917f
C4868 vdd.n2767 gnd 0.006917f
C4869 vdd.n2768 gnd 0.006917f
C4870 vdd.n2769 gnd 0.006917f
C4871 vdd.n2770 gnd 0.006917f
C4872 vdd.n2771 gnd 0.006917f
C4873 vdd.n2772 gnd 0.006917f
C4874 vdd.n2773 gnd 0.006917f
C4875 vdd.n2774 gnd 0.006917f
C4876 vdd.n2775 gnd 0.006917f
C4877 vdd.n2776 gnd 0.006917f
C4878 vdd.n2777 gnd 0.006917f
C4879 vdd.n2778 gnd 0.006917f
C4880 vdd.n2779 gnd 0.006917f
C4881 vdd.n2780 gnd 0.006917f
C4882 vdd.n2781 gnd 0.006917f
C4883 vdd.n2782 gnd 0.015705f
C4884 vdd.n2783 gnd 0.015705f
C4885 vdd.n2784 gnd 0.862789f
C4886 vdd.t278 gnd 3.06654f
C4887 vdd.t263 gnd 3.06654f
C4888 vdd.n2818 gnd 0.015705f
C4889 vdd.t270 gnd 0.602912f
C4890 vdd.n2819 gnd 0.006917f
C4891 vdd.t62 gnd 0.279506f
C4892 vdd.t63 gnd 0.28611f
C4893 vdd.t60 gnd 0.182472f
C4894 vdd.n2820 gnd 0.098616f
C4895 vdd.n2821 gnd 0.055938f
C4896 vdd.n2822 gnd 0.006917f
C4897 vdd.t69 gnd 0.279506f
C4898 vdd.t70 gnd 0.28611f
C4899 vdd.t68 gnd 0.182472f
C4900 vdd.n2823 gnd 0.098616f
C4901 vdd.n2824 gnd 0.055938f
C4902 vdd.n2825 gnd 0.009885f
C4903 vdd.n2826 gnd 0.015705f
C4904 vdd.n2827 gnd 0.015705f
C4905 vdd.n2828 gnd 0.006917f
C4906 vdd.n2829 gnd 0.006917f
C4907 vdd.n2830 gnd 0.006917f
C4908 vdd.n2831 gnd 0.006917f
C4909 vdd.n2832 gnd 0.006917f
C4910 vdd.n2833 gnd 0.006917f
C4911 vdd.n2834 gnd 0.006917f
C4912 vdd.n2835 gnd 0.006917f
C4913 vdd.n2836 gnd 0.006917f
C4914 vdd.n2837 gnd 0.006917f
C4915 vdd.n2838 gnd 0.006917f
C4916 vdd.n2839 gnd 0.006917f
C4917 vdd.n2840 gnd 0.006917f
C4918 vdd.n2841 gnd 0.006917f
C4919 vdd.n2842 gnd 0.006917f
C4920 vdd.n2843 gnd 0.006917f
C4921 vdd.n2844 gnd 0.006917f
C4922 vdd.n2845 gnd 0.006917f
C4923 vdd.n2846 gnd 0.006917f
C4924 vdd.n2847 gnd 0.006917f
C4925 vdd.n2848 gnd 0.006917f
C4926 vdd.n2849 gnd 0.006917f
C4927 vdd.n2850 gnd 0.006917f
C4928 vdd.n2851 gnd 0.006917f
C4929 vdd.n2852 gnd 0.006917f
C4930 vdd.n2853 gnd 0.006917f
C4931 vdd.n2854 gnd 0.006917f
C4932 vdd.n2855 gnd 0.006917f
C4933 vdd.n2856 gnd 0.006917f
C4934 vdd.n2857 gnd 0.006917f
C4935 vdd.n2858 gnd 0.006917f
C4936 vdd.n2859 gnd 0.006917f
C4937 vdd.n2860 gnd 0.006917f
C4938 vdd.n2861 gnd 0.006917f
C4939 vdd.n2862 gnd 0.006917f
C4940 vdd.n2863 gnd 0.006917f
C4941 vdd.n2864 gnd 0.006917f
C4942 vdd.n2865 gnd 0.006917f
C4943 vdd.n2866 gnd 0.006917f
C4944 vdd.n2867 gnd 0.006917f
C4945 vdd.n2868 gnd 0.006917f
C4946 vdd.n2869 gnd 0.006917f
C4947 vdd.n2870 gnd 0.006917f
C4948 vdd.n2871 gnd 0.006917f
C4949 vdd.n2872 gnd 0.006917f
C4950 vdd.n2873 gnd 0.006917f
C4951 vdd.n2874 gnd 0.006917f
C4952 vdd.n2875 gnd 0.006917f
C4953 vdd.n2876 gnd 0.006917f
C4954 vdd.n2877 gnd 0.006917f
C4955 vdd.n2878 gnd 0.006917f
C4956 vdd.n2879 gnd 0.006917f
C4957 vdd.n2880 gnd 0.006917f
C4958 vdd.n2881 gnd 0.006917f
C4959 vdd.n2882 gnd 0.006917f
C4960 vdd.n2883 gnd 0.006917f
C4961 vdd.n2884 gnd 0.006917f
C4962 vdd.n2885 gnd 0.006917f
C4963 vdd.n2886 gnd 0.006917f
C4964 vdd.n2887 gnd 0.006917f
C4965 vdd.n2888 gnd 0.005035f
C4966 vdd.n2889 gnd 0.006917f
C4967 vdd.n2890 gnd 0.006917f
C4968 vdd.n2891 gnd 0.00534f
C4969 vdd.n2892 gnd 0.006917f
C4970 vdd.n2893 gnd 0.006917f
C4971 vdd.n2894 gnd 0.015705f
C4972 vdd.n2895 gnd 0.01481f
C4973 vdd.n2896 gnd 0.01481f
C4974 vdd.n2897 gnd 0.006917f
C4975 vdd.n2898 gnd 0.006917f
C4976 vdd.n2899 gnd 0.006917f
C4977 vdd.n2900 gnd 0.006917f
C4978 vdd.n2901 gnd 0.006917f
C4979 vdd.n2902 gnd 0.006917f
C4980 vdd.n2903 gnd 0.006917f
C4981 vdd.n2904 gnd 0.006917f
C4982 vdd.n2905 gnd 0.006917f
C4983 vdd.n2906 gnd 0.006917f
C4984 vdd.n2907 gnd 0.006917f
C4985 vdd.n2908 gnd 0.006917f
C4986 vdd.n2909 gnd 0.006917f
C4987 vdd.n2910 gnd 0.006917f
C4988 vdd.n2911 gnd 0.006917f
C4989 vdd.n2912 gnd 0.006917f
C4990 vdd.n2913 gnd 0.006917f
C4991 vdd.n2914 gnd 0.006917f
C4992 vdd.n2915 gnd 0.006917f
C4993 vdd.n2916 gnd 0.006917f
C4994 vdd.n2917 gnd 0.006917f
C4995 vdd.n2918 gnd 0.006917f
C4996 vdd.n2919 gnd 0.006917f
C4997 vdd.n2920 gnd 0.006917f
C4998 vdd.n2921 gnd 0.006917f
C4999 vdd.n2922 gnd 0.006917f
C5000 vdd.n2923 gnd 0.006917f
C5001 vdd.n2924 gnd 0.006917f
C5002 vdd.n2925 gnd 0.006917f
C5003 vdd.n2926 gnd 0.006917f
C5004 vdd.n2927 gnd 0.006917f
C5005 vdd.n2928 gnd 0.006917f
C5006 vdd.n2929 gnd 0.006917f
C5007 vdd.n2930 gnd 0.006917f
C5008 vdd.n2931 gnd 0.006917f
C5009 vdd.n2932 gnd 0.006917f
C5010 vdd.n2933 gnd 0.006917f
C5011 vdd.n2934 gnd 0.006917f
C5012 vdd.n2935 gnd 0.006917f
C5013 vdd.n2936 gnd 0.006917f
C5014 vdd.n2937 gnd 0.006917f
C5015 vdd.n2938 gnd 0.006917f
C5016 vdd.n2939 gnd 0.006917f
C5017 vdd.n2940 gnd 0.006917f
C5018 vdd.n2941 gnd 0.006917f
C5019 vdd.n2942 gnd 0.006917f
C5020 vdd.n2943 gnd 0.006917f
C5021 vdd.n2944 gnd 0.006917f
C5022 vdd.n2945 gnd 0.006917f
C5023 vdd.n2946 gnd 0.006917f
C5024 vdd.n2947 gnd 0.006917f
C5025 vdd.n2948 gnd 0.006917f
C5026 vdd.n2949 gnd 0.006917f
C5027 vdd.n2950 gnd 0.006917f
C5028 vdd.n2951 gnd 0.006917f
C5029 vdd.n2952 gnd 0.006917f
C5030 vdd.n2953 gnd 0.006917f
C5031 vdd.n2954 gnd 0.006917f
C5032 vdd.n2955 gnd 0.006917f
C5033 vdd.n2956 gnd 0.006917f
C5034 vdd.n2957 gnd 0.006917f
C5035 vdd.n2958 gnd 0.006917f
C5036 vdd.n2959 gnd 0.006917f
C5037 vdd.n2960 gnd 0.006917f
C5038 vdd.n2961 gnd 0.006917f
C5039 vdd.n2962 gnd 0.006917f
C5040 vdd.n2963 gnd 0.006917f
C5041 vdd.n2964 gnd 0.006917f
C5042 vdd.n2965 gnd 0.006917f
C5043 vdd.n2966 gnd 0.006917f
C5044 vdd.n2967 gnd 0.006917f
C5045 vdd.n2968 gnd 0.006917f
C5046 vdd.n2969 gnd 0.006917f
C5047 vdd.n2970 gnd 0.006917f
C5048 vdd.n2971 gnd 0.006917f
C5049 vdd.n2972 gnd 0.006917f
C5050 vdd.n2973 gnd 0.006917f
C5051 vdd.n2974 gnd 0.006917f
C5052 vdd.n2975 gnd 0.006917f
C5053 vdd.n2976 gnd 0.006917f
C5054 vdd.n2977 gnd 0.006917f
C5055 vdd.n2978 gnd 0.006917f
C5056 vdd.n2979 gnd 0.006917f
C5057 vdd.n2980 gnd 0.006917f
C5058 vdd.n2981 gnd 0.006917f
C5059 vdd.n2982 gnd 0.006917f
C5060 vdd.n2983 gnd 0.006917f
C5061 vdd.n2984 gnd 0.006917f
C5062 vdd.n2985 gnd 0.006917f
C5063 vdd.n2986 gnd 0.006917f
C5064 vdd.n2987 gnd 0.006917f
C5065 vdd.n2988 gnd 0.006917f
C5066 vdd.n2989 gnd 0.006917f
C5067 vdd.n2990 gnd 0.006917f
C5068 vdd.n2991 gnd 0.006917f
C5069 vdd.n2992 gnd 0.006917f
C5070 vdd.n2993 gnd 0.006917f
C5071 vdd.n2994 gnd 0.006917f
C5072 vdd.n2995 gnd 0.006917f
C5073 vdd.n2996 gnd 0.006917f
C5074 vdd.n2997 gnd 0.006917f
C5075 vdd.n2998 gnd 0.223493f
C5076 vdd.n2999 gnd 0.006917f
C5077 vdd.n3000 gnd 0.006917f
C5078 vdd.n3001 gnd 0.006917f
C5079 vdd.n3002 gnd 0.006917f
C5080 vdd.n3003 gnd 0.006917f
C5081 vdd.n3004 gnd 0.223493f
C5082 vdd.n3005 gnd 0.006917f
C5083 vdd.n3006 gnd 0.006917f
C5084 vdd.n3007 gnd 0.006917f
C5085 vdd.n3008 gnd 0.006917f
C5086 vdd.n3009 gnd 0.006917f
C5087 vdd.n3010 gnd 0.006917f
C5088 vdd.n3011 gnd 0.006917f
C5089 vdd.n3012 gnd 0.006917f
C5090 vdd.n3013 gnd 0.006917f
C5091 vdd.n3014 gnd 0.006917f
C5092 vdd.n3015 gnd 0.006917f
C5093 vdd.n3016 gnd 0.441789f
C5094 vdd.n3017 gnd 0.006917f
C5095 vdd.n3018 gnd 0.006917f
C5096 vdd.n3019 gnd 0.006917f
C5097 vdd.n3020 gnd 0.01481f
C5098 vdd.n3021 gnd 0.01481f
C5099 vdd.n3022 gnd 0.015705f
C5100 vdd.n3023 gnd 0.015705f
C5101 vdd.n3024 gnd 0.006917f
C5102 vdd.n3025 gnd 0.006917f
C5103 vdd.n3026 gnd 0.006917f
C5104 vdd.n3027 gnd 0.00534f
C5105 vdd.n3028 gnd 0.009885f
C5106 vdd.n3029 gnd 0.005035f
C5107 vdd.n3030 gnd 0.006917f
C5108 vdd.n3031 gnd 0.006917f
C5109 vdd.n3032 gnd 0.006917f
C5110 vdd.n3033 gnd 0.006917f
C5111 vdd.n3034 gnd 0.006917f
C5112 vdd.n3035 gnd 0.006917f
C5113 vdd.n3036 gnd 0.006917f
C5114 vdd.n3037 gnd 0.006917f
C5115 vdd.n3038 gnd 0.006917f
C5116 vdd.n3039 gnd 0.006917f
C5117 vdd.n3040 gnd 0.006917f
C5118 vdd.n3041 gnd 0.006917f
C5119 vdd.n3042 gnd 0.006917f
C5120 vdd.n3043 gnd 0.006917f
C5121 vdd.n3044 gnd 0.006917f
C5122 vdd.n3045 gnd 0.006917f
C5123 vdd.n3046 gnd 0.006917f
C5124 vdd.n3047 gnd 0.006917f
C5125 vdd.n3048 gnd 0.006917f
C5126 vdd.n3049 gnd 0.006917f
C5127 vdd.n3050 gnd 0.006917f
C5128 vdd.n3051 gnd 0.006917f
C5129 vdd.n3052 gnd 0.006917f
C5130 vdd.n3053 gnd 0.006917f
C5131 vdd.n3054 gnd 0.006917f
C5132 vdd.n3055 gnd 0.006917f
C5133 vdd.n3056 gnd 0.006917f
C5134 vdd.n3057 gnd 0.006917f
C5135 vdd.n3058 gnd 0.006917f
C5136 vdd.n3059 gnd 0.006917f
C5137 vdd.n3060 gnd 0.006917f
C5138 vdd.n3061 gnd 0.006917f
C5139 vdd.n3062 gnd 0.006917f
C5140 vdd.n3063 gnd 0.006917f
C5141 vdd.n3064 gnd 0.006917f
C5142 vdd.n3065 gnd 0.006917f
C5143 vdd.n3066 gnd 0.006917f
C5144 vdd.n3067 gnd 0.006917f
C5145 vdd.n3068 gnd 0.006917f
C5146 vdd.n3069 gnd 0.006917f
C5147 vdd.n3070 gnd 0.006917f
C5148 vdd.n3071 gnd 0.006917f
C5149 vdd.n3072 gnd 0.006917f
C5150 vdd.n3073 gnd 0.006917f
C5151 vdd.n3074 gnd 0.006917f
C5152 vdd.n3075 gnd 0.006917f
C5153 vdd.n3076 gnd 0.006917f
C5154 vdd.n3077 gnd 0.006917f
C5155 vdd.n3078 gnd 0.006917f
C5156 vdd.n3079 gnd 0.006917f
C5157 vdd.n3080 gnd 0.006917f
C5158 vdd.n3081 gnd 0.006917f
C5159 vdd.n3082 gnd 0.006917f
C5160 vdd.n3083 gnd 0.006917f
C5161 vdd.n3084 gnd 0.006917f
C5162 vdd.n3085 gnd 0.006917f
C5163 vdd.n3086 gnd 0.006917f
C5164 vdd.n3087 gnd 0.006917f
C5165 vdd.n3088 gnd 0.862789f
C5166 vdd.n3090 gnd 0.015705f
C5167 vdd.n3091 gnd 0.015705f
C5168 vdd.n3092 gnd 0.01481f
C5169 vdd.n3093 gnd 0.006917f
C5170 vdd.n3094 gnd 0.006917f
C5171 vdd.n3095 gnd 0.415802f
C5172 vdd.n3096 gnd 0.006917f
C5173 vdd.n3097 gnd 0.006917f
C5174 vdd.n3098 gnd 0.006917f
C5175 vdd.n3099 gnd 0.006917f
C5176 vdd.n3100 gnd 0.006917f
C5177 vdd.n3101 gnd 0.420999f
C5178 vdd.n3102 gnd 0.006917f
C5179 vdd.n3103 gnd 0.006917f
C5180 vdd.n3104 gnd 0.006917f
C5181 vdd.n3105 gnd 0.006917f
C5182 vdd.n3106 gnd 0.006917f
C5183 vdd.n3107 gnd 0.706863f
C5184 vdd.n3108 gnd 0.006917f
C5185 vdd.n3109 gnd 0.006917f
C5186 vdd.n3110 gnd 0.006917f
C5187 vdd.n3111 gnd 0.006917f
C5188 vdd.n3112 gnd 0.006917f
C5189 vdd.n3113 gnd 0.509357f
C5190 vdd.n3114 gnd 0.006917f
C5191 vdd.n3115 gnd 0.006917f
C5192 vdd.n3116 gnd 0.006917f
C5193 vdd.n3117 gnd 0.006917f
C5194 vdd.n3118 gnd 0.006917f
C5195 vdd.n3119 gnd 0.639295f
C5196 vdd.n3120 gnd 0.006917f
C5197 vdd.n3121 gnd 0.006917f
C5198 vdd.n3122 gnd 0.006917f
C5199 vdd.n3123 gnd 0.006917f
C5200 vdd.n3124 gnd 0.006917f
C5201 vdd.n3125 gnd 0.52495f
C5202 vdd.n3126 gnd 0.006917f
C5203 vdd.n3127 gnd 0.006917f
C5204 vdd.n3128 gnd 0.006917f
C5205 vdd.n3129 gnd 0.006917f
C5206 vdd.n3130 gnd 0.006917f
C5207 vdd.n3131 gnd 0.369024f
C5208 vdd.n3132 gnd 0.006917f
C5209 vdd.n3133 gnd 0.006917f
C5210 vdd.n3134 gnd 0.006917f
C5211 vdd.n3135 gnd 0.006917f
C5212 vdd.n3136 gnd 0.006917f
C5213 vdd.n3137 gnd 0.223493f
C5214 vdd.n3138 gnd 0.006917f
C5215 vdd.n3139 gnd 0.006917f
C5216 vdd.n3140 gnd 0.006917f
C5217 vdd.n3141 gnd 0.006917f
C5218 vdd.n3142 gnd 0.006917f
C5219 vdd.n3143 gnd 0.64969f
C5220 vdd.n3144 gnd 0.006917f
C5221 vdd.n3145 gnd 0.006917f
C5222 vdd.n3146 gnd 0.006917f
C5223 vdd.n3147 gnd 0.004882f
C5224 vdd.n3148 gnd 0.006917f
C5225 vdd.n3149 gnd 0.006917f
C5226 vdd.n3150 gnd 0.706863f
C5227 vdd.n3151 gnd 0.006917f
C5228 vdd.n3152 gnd 0.006917f
C5229 vdd.n3153 gnd 0.006917f
C5230 vdd.n3154 gnd 0.006917f
C5231 vdd.n3155 gnd 0.006917f
C5232 vdd.n3156 gnd 0.561332f
C5233 vdd.n3157 gnd 0.006917f
C5234 vdd.n3158 gnd 0.005493f
C5235 vdd.n3159 gnd 0.006917f
C5236 vdd.n3160 gnd 0.006917f
C5237 vdd.n3161 gnd 0.006917f
C5238 vdd.n3162 gnd 0.452184f
C5239 vdd.n3163 gnd 0.006917f
C5240 vdd.n3164 gnd 0.006917f
C5241 vdd.n3165 gnd 0.006917f
C5242 vdd.n3166 gnd 0.006917f
C5243 vdd.n3167 gnd 0.006917f
C5244 vdd.n3168 gnd 0.410604f
C5245 vdd.n3169 gnd 0.006917f
C5246 vdd.n3170 gnd 0.006917f
C5247 vdd.n3171 gnd 0.006917f
C5248 vdd.n3172 gnd 0.006917f
C5249 vdd.n3173 gnd 0.006917f
C5250 vdd.n3174 gnd 0.56653f
C5251 vdd.n3175 gnd 0.006917f
C5252 vdd.n3176 gnd 0.006917f
C5253 vdd.n3177 gnd 0.006917f
C5254 vdd.n3178 gnd 0.006917f
C5255 vdd.n3179 gnd 0.006917f
C5256 vdd.n3180 gnd 0.706863f
C5257 vdd.n3181 gnd 0.006917f
C5258 vdd.n3182 gnd 0.006917f
C5259 vdd.n3183 gnd 0.006917f
C5260 vdd.n3184 gnd 0.006917f
C5261 vdd.n3185 gnd 0.006917f
C5262 vdd.n3186 gnd 0.69127f
C5263 vdd.n3187 gnd 0.006917f
C5264 vdd.n3188 gnd 0.006917f
C5265 vdd.n3189 gnd 0.006917f
C5266 vdd.n3190 gnd 0.006917f
C5267 vdd.n3191 gnd 0.006917f
C5268 vdd.n3192 gnd 0.535345f
C5269 vdd.n3193 gnd 0.006917f
C5270 vdd.n3194 gnd 0.006917f
C5271 vdd.n3195 gnd 0.006917f
C5272 vdd.n3196 gnd 0.006917f
C5273 vdd.n3197 gnd 0.006917f
C5274 vdd.n3198 gnd 0.379419f
C5275 vdd.n3199 gnd 0.006917f
C5276 vdd.n3200 gnd 0.006917f
C5277 vdd.n3201 gnd 0.006917f
C5278 vdd.n3202 gnd 0.006917f
C5279 vdd.n3203 gnd 0.006917f
C5280 vdd.n3204 gnd 0.706863f
C5281 vdd.n3205 gnd 0.006917f
C5282 vdd.n3206 gnd 0.006917f
C5283 vdd.n3207 gnd 0.006917f
C5284 vdd.n3208 gnd 0.006917f
C5285 vdd.n3209 gnd 0.006917f
C5286 vdd.n3210 gnd 0.006917f
C5287 vdd.n3212 gnd 0.006917f
C5288 vdd.n3213 gnd 0.006917f
C5289 vdd.n3215 gnd 0.006917f
C5290 vdd.n3216 gnd 0.006917f
C5291 vdd.n3219 gnd 0.006917f
C5292 vdd.n3220 gnd 0.006917f
C5293 vdd.n3221 gnd 0.006917f
C5294 vdd.n3222 gnd 0.006917f
C5295 vdd.n3224 gnd 0.006917f
C5296 vdd.n3225 gnd 0.006917f
C5297 vdd.n3226 gnd 0.006917f
C5298 vdd.n3227 gnd 0.006917f
C5299 vdd.n3228 gnd 0.006917f
C5300 vdd.n3229 gnd 0.006917f
C5301 vdd.n3231 gnd 0.006917f
C5302 vdd.n3232 gnd 0.006917f
C5303 vdd.n3233 gnd 0.006917f
C5304 vdd.n3234 gnd 0.006917f
C5305 vdd.n3235 gnd 0.006917f
C5306 vdd.n3236 gnd 0.006917f
C5307 vdd.n3238 gnd 0.006917f
C5308 vdd.n3239 gnd 0.006917f
C5309 vdd.n3240 gnd 0.006917f
C5310 vdd.n3241 gnd 0.006917f
C5311 vdd.n3242 gnd 0.006917f
C5312 vdd.n3243 gnd 0.006917f
C5313 vdd.n3245 gnd 0.006917f
C5314 vdd.n3246 gnd 0.015705f
C5315 vdd.n3247 gnd 0.015705f
C5316 vdd.n3248 gnd 0.01481f
C5317 vdd.n3249 gnd 0.006917f
C5318 vdd.n3250 gnd 0.006917f
C5319 vdd.n3251 gnd 0.006917f
C5320 vdd.n3252 gnd 0.006917f
C5321 vdd.n3253 gnd 0.006917f
C5322 vdd.n3254 gnd 0.006917f
C5323 vdd.n3255 gnd 0.706863f
C5324 vdd.n3256 gnd 0.006917f
C5325 vdd.n3257 gnd 0.006917f
C5326 vdd.n3258 gnd 0.006917f
C5327 vdd.n3259 gnd 0.006917f
C5328 vdd.n3260 gnd 0.006917f
C5329 vdd.n3261 gnd 0.50416f
C5330 vdd.n3262 gnd 0.006917f
C5331 vdd.n3263 gnd 0.006917f
C5332 vdd.n3264 gnd 0.006917f
C5333 vdd.n3265 gnd 0.015705f
C5334 vdd.n3266 gnd 0.01481f
C5335 vdd.n3267 gnd 0.015705f
C5336 vdd.n3269 gnd 0.006917f
C5337 vdd.n3270 gnd 0.006917f
C5338 vdd.n3271 gnd 0.00534f
C5339 vdd.n3272 gnd 0.009885f
C5340 vdd.n3273 gnd 0.005035f
C5341 vdd.n3274 gnd 0.006917f
C5342 vdd.n3275 gnd 0.006917f
C5343 vdd.n3277 gnd 0.006917f
C5344 vdd.n3278 gnd 0.006917f
C5345 vdd.n3279 gnd 0.006917f
C5346 vdd.n3280 gnd 0.006917f
C5347 vdd.n3281 gnd 0.006917f
C5348 vdd.n3282 gnd 0.006917f
C5349 vdd.n3284 gnd 0.006917f
C5350 vdd.n3285 gnd 0.006917f
C5351 vdd.n3286 gnd 0.006917f
C5352 vdd.n3287 gnd 0.006917f
C5353 vdd.n3288 gnd 0.006917f
C5354 vdd.n3289 gnd 0.006917f
C5355 vdd.n3291 gnd 0.006917f
C5356 vdd.n3292 gnd 0.006917f
C5357 vdd.n3293 gnd 0.006917f
C5358 vdd.n3294 gnd 0.006917f
C5359 vdd.n3295 gnd 0.006917f
C5360 vdd.n3296 gnd 0.006917f
C5361 vdd.n3298 gnd 0.006917f
C5362 vdd.n3299 gnd 0.006917f
C5363 vdd.n3300 gnd 0.006917f
C5364 vdd.n3302 gnd 0.006917f
C5365 vdd.n3303 gnd 0.006917f
C5366 vdd.n3304 gnd 0.006917f
C5367 vdd.n3305 gnd 0.006917f
C5368 vdd.n3306 gnd 0.006917f
C5369 vdd.n3307 gnd 0.006917f
C5370 vdd.n3309 gnd 0.006917f
C5371 vdd.n3310 gnd 0.006917f
C5372 vdd.n3311 gnd 0.006917f
C5373 vdd.n3312 gnd 0.006917f
C5374 vdd.n3313 gnd 0.006917f
C5375 vdd.n3314 gnd 0.006917f
C5376 vdd.n3316 gnd 0.006917f
C5377 vdd.n3317 gnd 0.006917f
C5378 vdd.n3318 gnd 0.006917f
C5379 vdd.n3319 gnd 0.006917f
C5380 vdd.n3320 gnd 0.006917f
C5381 vdd.n3321 gnd 0.006917f
C5382 vdd.n3323 gnd 0.006917f
C5383 vdd.n3324 gnd 0.006917f
C5384 vdd.n3326 gnd 0.006917f
C5385 vdd.n3327 gnd 0.006917f
C5386 vdd.n3328 gnd 0.015705f
C5387 vdd.n3329 gnd 0.01481f
C5388 vdd.n3330 gnd 0.01481f
C5389 vdd.n3331 gnd 0.956344f
C5390 vdd.n3332 gnd 0.01481f
C5391 vdd.n3333 gnd 0.015705f
C5392 vdd.n3334 gnd 0.01481f
C5393 vdd.n3335 gnd 0.006917f
C5394 vdd.n3336 gnd 0.00534f
C5395 vdd.n3337 gnd 0.006917f
C5396 vdd.n3339 gnd 0.006917f
C5397 vdd.n3340 gnd 0.006917f
C5398 vdd.n3341 gnd 0.006917f
C5399 vdd.n3342 gnd 0.006917f
C5400 vdd.n3343 gnd 0.006917f
C5401 vdd.n3344 gnd 0.006917f
C5402 vdd.n3346 gnd 0.006917f
C5403 vdd.n3347 gnd 0.006917f
C5404 vdd.n3348 gnd 0.006917f
C5405 vdd.n3349 gnd 0.006917f
C5406 vdd.n3350 gnd 0.006917f
C5407 vdd.n3351 gnd 0.006917f
C5408 vdd.n3353 gnd 0.006917f
C5409 vdd.n3354 gnd 0.006917f
C5410 vdd.n3355 gnd 0.006917f
C5411 vdd.n3356 gnd 0.006917f
C5412 vdd.n3357 gnd 0.006917f
C5413 vdd.n3358 gnd 0.006917f
C5414 vdd.n3360 gnd 0.006917f
C5415 vdd.n3361 gnd 0.006917f
C5416 vdd.n3363 gnd 0.006917f
C5417 vdd.n3364 gnd 0.04271f
C5418 vdd.n3365 gnd 1.08372f
C5419 vdd.n3367 gnd 0.004298f
C5420 vdd.n3368 gnd 0.008187f
C5421 vdd.n3369 gnd 0.010172f
C5422 vdd.n3370 gnd 0.010172f
C5423 vdd.n3371 gnd 0.008187f
C5424 vdd.n3372 gnd 0.008187f
C5425 vdd.n3373 gnd 0.010172f
C5426 vdd.n3374 gnd 0.010172f
C5427 vdd.n3375 gnd 0.008187f
C5428 vdd.n3376 gnd 0.008187f
C5429 vdd.n3377 gnd 0.010172f
C5430 vdd.n3378 gnd 0.010172f
C5431 vdd.n3379 gnd 0.008187f
C5432 vdd.n3380 gnd 0.008187f
C5433 vdd.n3381 gnd 0.010172f
C5434 vdd.n3382 gnd 0.010172f
C5435 vdd.n3383 gnd 0.008187f
C5436 vdd.n3384 gnd 0.008187f
C5437 vdd.n3385 gnd 0.010172f
C5438 vdd.n3386 gnd 0.010172f
C5439 vdd.n3387 gnd 0.008187f
C5440 vdd.n3388 gnd 0.008187f
C5441 vdd.n3389 gnd 0.010172f
C5442 vdd.n3390 gnd 0.010172f
C5443 vdd.n3391 gnd 0.008187f
C5444 vdd.n3392 gnd 0.008187f
C5445 vdd.n3393 gnd 0.010172f
C5446 vdd.n3394 gnd 0.010172f
C5447 vdd.n3395 gnd 0.008187f
C5448 vdd.n3396 gnd 0.008187f
C5449 vdd.n3397 gnd 0.010172f
C5450 vdd.n3398 gnd 0.010172f
C5451 vdd.n3399 gnd 0.008187f
C5452 vdd.n3400 gnd 0.008187f
C5453 vdd.n3401 gnd 0.010172f
C5454 vdd.n3402 gnd 0.010172f
C5455 vdd.n3403 gnd 0.008187f
C5456 vdd.n3404 gnd 0.010172f
C5457 vdd.n3405 gnd 0.010172f
C5458 vdd.n3406 gnd 0.008187f
C5459 vdd.n3407 gnd 0.010172f
C5460 vdd.n3408 gnd 0.010172f
C5461 vdd.n3409 gnd 0.010172f
C5462 vdd.n3410 gnd 0.016701f
C5463 vdd.n3411 gnd 0.010172f
C5464 vdd.n3412 gnd 0.010172f
C5465 vdd.n3413 gnd 0.005567f
C5466 vdd.n3414 gnd 0.008187f
C5467 vdd.n3415 gnd 0.010172f
C5468 vdd.n3416 gnd 0.010172f
C5469 vdd.n3417 gnd 0.008187f
C5470 vdd.n3418 gnd 0.008187f
C5471 vdd.n3419 gnd 0.010172f
C5472 vdd.n3420 gnd 0.010172f
C5473 vdd.n3421 gnd 0.008187f
C5474 vdd.n3422 gnd 0.008187f
C5475 vdd.n3423 gnd 0.010172f
C5476 vdd.n3424 gnd 0.010172f
C5477 vdd.n3425 gnd 0.008187f
C5478 vdd.n3426 gnd 0.008187f
C5479 vdd.n3427 gnd 0.010172f
C5480 vdd.n3428 gnd 0.010172f
C5481 vdd.n3429 gnd 0.008187f
C5482 vdd.n3430 gnd 0.008187f
C5483 vdd.n3431 gnd 0.010172f
C5484 vdd.n3432 gnd 0.010172f
C5485 vdd.n3433 gnd 0.008187f
C5486 vdd.n3434 gnd 0.008187f
C5487 vdd.n3435 gnd 0.010172f
C5488 vdd.n3436 gnd 0.010172f
C5489 vdd.n3437 gnd 0.008187f
C5490 vdd.n3438 gnd 0.008187f
C5491 vdd.n3439 gnd 0.010172f
C5492 vdd.n3440 gnd 0.010172f
C5493 vdd.n3441 gnd 0.008187f
C5494 vdd.n3442 gnd 0.008187f
C5495 vdd.n3443 gnd 0.010172f
C5496 vdd.n3444 gnd 0.010172f
C5497 vdd.n3445 gnd 0.008187f
C5498 vdd.n3446 gnd 0.008187f
C5499 vdd.n3447 gnd 0.010172f
C5500 vdd.n3448 gnd 0.010172f
C5501 vdd.n3449 gnd 0.008187f
C5502 vdd.n3450 gnd 0.010172f
C5503 vdd.n3451 gnd 0.010172f
C5504 vdd.n3452 gnd 0.008187f
C5505 vdd.n3453 gnd 0.010172f
C5506 vdd.n3454 gnd 0.010172f
C5507 vdd.n3455 gnd 0.010172f
C5508 vdd.t58 gnd 0.125139f
C5509 vdd.t59 gnd 0.133739f
C5510 vdd.t57 gnd 0.16343f
C5511 vdd.n3456 gnd 0.209494f
C5512 vdd.n3457 gnd 0.176013f
C5513 vdd.n3458 gnd 0.016701f
C5514 vdd.n3459 gnd 0.010172f
C5515 vdd.n3460 gnd 0.010172f
C5516 vdd.n3461 gnd 0.006836f
C5517 vdd.n3462 gnd 0.008187f
C5518 vdd.n3463 gnd 0.010172f
C5519 vdd.n3464 gnd 0.010172f
C5520 vdd.n3465 gnd 0.008187f
C5521 vdd.n3466 gnd 0.008187f
C5522 vdd.n3467 gnd 0.010172f
C5523 vdd.n3468 gnd 0.010172f
C5524 vdd.n3469 gnd 0.008187f
C5525 vdd.n3470 gnd 0.008187f
C5526 vdd.n3471 gnd 0.010172f
C5527 vdd.n3472 gnd 0.010172f
C5528 vdd.n3473 gnd 0.008187f
C5529 vdd.n3474 gnd 0.008187f
C5530 vdd.n3475 gnd 0.010172f
C5531 vdd.n3476 gnd 0.010172f
C5532 vdd.n3477 gnd 0.008187f
C5533 vdd.n3478 gnd 0.008187f
C5534 vdd.n3479 gnd 0.010172f
C5535 vdd.n3480 gnd 0.010172f
C5536 vdd.n3481 gnd 0.008187f
C5537 vdd.n3482 gnd 0.008187f
C5538 vdd.n3483 gnd 0.010172f
C5539 vdd.n3484 gnd 0.010172f
C5540 vdd.n3485 gnd 0.008187f
C5541 vdd.n3486 gnd 0.008187f
C5542 vdd.n3488 gnd 1.08372f
C5543 vdd.n3490 gnd 0.008187f
C5544 vdd.n3491 gnd 0.008187f
C5545 vdd.n3492 gnd 0.006795f
C5546 vdd.n3493 gnd 0.025134f
C5547 vdd.n3495 gnd 12.6923f
C5548 vdd.n3496 gnd 0.025134f
C5549 vdd.n3497 gnd 0.003889f
C5550 vdd.n3498 gnd 0.025134f
C5551 vdd.n3499 gnd 0.024606f
C5552 vdd.n3500 gnd 0.010172f
C5553 vdd.n3501 gnd 0.008187f
C5554 vdd.n3502 gnd 0.010172f
C5555 vdd.n3503 gnd 0.6289f
C5556 vdd.n3504 gnd 0.010172f
C5557 vdd.n3505 gnd 0.008187f
C5558 vdd.n3506 gnd 0.010172f
C5559 vdd.n3507 gnd 0.010172f
C5560 vdd.n3508 gnd 0.010172f
C5561 vdd.n3509 gnd 0.008187f
C5562 vdd.n3510 gnd 0.010172f
C5563 vdd.n3511 gnd 1.0395f
C5564 vdd.n3512 gnd 0.010172f
C5565 vdd.n3513 gnd 0.008187f
C5566 vdd.n3514 gnd 0.010172f
C5567 vdd.n3515 gnd 0.010172f
C5568 vdd.n3516 gnd 0.010172f
C5569 vdd.n3517 gnd 0.008187f
C5570 vdd.n3518 gnd 0.010172f
C5571 vdd.n3519 gnd 0.67048f
C5572 vdd.n3520 gnd 0.71206f
C5573 vdd.n3521 gnd 0.010172f
C5574 vdd.n3522 gnd 0.008187f
C5575 vdd.n3523 gnd 0.010172f
C5576 vdd.n3524 gnd 0.010172f
C5577 vdd.n3525 gnd 0.010172f
C5578 vdd.n3526 gnd 0.008187f
C5579 vdd.n3527 gnd 0.010172f
C5580 vdd.n3528 gnd 0.862789f
C5581 vdd.n3529 gnd 0.010172f
C5582 vdd.n3530 gnd 0.008187f
C5583 vdd.n3531 gnd 0.010172f
C5584 vdd.n3532 gnd 0.010172f
C5585 vdd.n3533 gnd 0.010172f
C5586 vdd.n3534 gnd 0.008187f
C5587 vdd.n3535 gnd 0.010172f
C5588 vdd.t113 gnd 0.519752f
C5589 vdd.n3536 gnd 0.836801f
C5590 vdd.n3537 gnd 0.010172f
C5591 vdd.n3538 gnd 0.008187f
C5592 vdd.n3539 gnd 0.010172f
C5593 vdd.n3540 gnd 0.010172f
C5594 vdd.n3541 gnd 0.010172f
C5595 vdd.n3542 gnd 0.008187f
C5596 vdd.n3543 gnd 0.010172f
C5597 vdd.n3544 gnd 0.660085f
C5598 vdd.n3545 gnd 0.010172f
C5599 vdd.n3546 gnd 0.008187f
C5600 vdd.n3547 gnd 0.010172f
C5601 vdd.n3548 gnd 0.010172f
C5602 vdd.n3549 gnd 0.010172f
C5603 vdd.n3550 gnd 0.008187f
C5604 vdd.n3551 gnd 0.010172f
C5605 vdd.n3552 gnd 0.826406f
C5606 vdd.n3553 gnd 0.556135f
C5607 vdd.n3554 gnd 0.010172f
C5608 vdd.n3555 gnd 0.008187f
C5609 vdd.n3556 gnd 0.010172f
C5610 vdd.n3557 gnd 0.010172f
C5611 vdd.n3558 gnd 0.010172f
C5612 vdd.n3559 gnd 0.008187f
C5613 vdd.n3560 gnd 0.010172f
C5614 vdd.n3561 gnd 0.732851f
C5615 vdd.n3562 gnd 0.010172f
C5616 vdd.n3563 gnd 0.008187f
C5617 vdd.n3564 gnd 0.010172f
C5618 vdd.n3565 gnd 0.010172f
C5619 vdd.n3566 gnd 0.010172f
C5620 vdd.n3567 gnd 0.010172f
C5621 vdd.n3568 gnd 0.010172f
C5622 vdd.n3569 gnd 0.008187f
C5623 vdd.n3570 gnd 0.008187f
C5624 vdd.n3571 gnd 0.010172f
C5625 vdd.t94 gnd 0.519752f
C5626 vdd.n3572 gnd 0.862789f
C5627 vdd.n3573 gnd 0.010172f
C5628 vdd.n3574 gnd 0.008187f
C5629 vdd.n3575 gnd 0.010172f
C5630 vdd.n3576 gnd 0.010172f
C5631 vdd.n3577 gnd 0.010172f
C5632 vdd.n3578 gnd 0.008187f
C5633 vdd.n3579 gnd 0.010172f
C5634 vdd.n3580 gnd 0.816011f
C5635 vdd.n3581 gnd 0.010172f
C5636 vdd.n3582 gnd 0.010172f
C5637 vdd.n3583 gnd 0.008187f
C5638 vdd.n3584 gnd 0.008187f
C5639 vdd.n3585 gnd 0.010172f
C5640 vdd.n3586 gnd 0.010172f
C5641 vdd.n3587 gnd 0.010172f
C5642 vdd.n3588 gnd 0.008187f
C5643 vdd.n3589 gnd 0.010172f
C5644 vdd.n3590 gnd 0.008187f
C5645 vdd.n3591 gnd 0.008187f
C5646 vdd.n3592 gnd 0.010172f
C5647 vdd.n3593 gnd 0.010172f
C5648 vdd.n3594 gnd 0.010172f
C5649 vdd.n3595 gnd 0.008187f
C5650 vdd.n3596 gnd 0.010172f
C5651 vdd.n3597 gnd 0.008187f
C5652 vdd.n3598 gnd 0.008187f
C5653 vdd.n3599 gnd 0.010172f
C5654 vdd.n3600 gnd 0.010172f
C5655 vdd.n3601 gnd 0.010172f
C5656 vdd.n3602 gnd 0.008187f
C5657 vdd.n3603 gnd 0.862789f
C5658 vdd.n3604 gnd 0.010172f
C5659 vdd.n3605 gnd 0.008187f
C5660 vdd.n3606 gnd 0.008187f
C5661 vdd.n3607 gnd 0.010172f
C5662 vdd.n3608 gnd 0.010172f
C5663 vdd.n3609 gnd 0.010172f
C5664 vdd.n3610 gnd 0.008187f
C5665 vdd.n3611 gnd 0.010172f
C5666 vdd.n3612 gnd 0.008187f
C5667 vdd.n3613 gnd 0.008187f
C5668 vdd.n3614 gnd 0.010172f
C5669 vdd.n3615 gnd 0.010172f
C5670 vdd.n3616 gnd 0.010172f
C5671 vdd.n3617 gnd 0.008187f
C5672 vdd.n3618 gnd 0.010172f
C5673 vdd.n3619 gnd 0.008187f
C5674 vdd.n3620 gnd 0.006795f
C5675 vdd.n3621 gnd 0.024606f
C5676 vdd.n3622 gnd 0.025134f
C5677 vdd.n3623 gnd 0.003889f
C5678 vdd.n3624 gnd 0.025134f
C5679 vdd.n3626 gnd 2.46363f
C5680 vdd.n3627 gnd 1.53327f
C5681 vdd.n3628 gnd 0.024606f
C5682 vdd.n3629 gnd 0.006795f
C5683 vdd.n3630 gnd 0.008187f
C5684 vdd.n3631 gnd 0.008187f
C5685 vdd.n3632 gnd 0.010172f
C5686 vdd.n3633 gnd 1.0395f
C5687 vdd.n3634 gnd 1.0395f
C5688 vdd.n3635 gnd 0.951146f
C5689 vdd.n3636 gnd 0.010172f
C5690 vdd.n3637 gnd 0.008187f
C5691 vdd.n3638 gnd 0.008187f
C5692 vdd.n3639 gnd 0.008187f
C5693 vdd.n3640 gnd 0.010172f
C5694 vdd.n3641 gnd 0.774431f
C5695 vdd.t100 gnd 0.519752f
C5696 vdd.n3642 gnd 0.784826f
C5697 vdd.n3643 gnd 0.597715f
C5698 vdd.n3644 gnd 0.010172f
C5699 vdd.n3645 gnd 0.008187f
C5700 vdd.n3646 gnd 0.008187f
C5701 vdd.n3647 gnd 0.008187f
C5702 vdd.n3648 gnd 0.010172f
C5703 vdd.n3649 gnd 0.618505f
C5704 vdd.n3650 gnd 0.764036f
C5705 vdd.t108 gnd 0.519752f
C5706 vdd.n3651 gnd 0.795221f
C5707 vdd.n3652 gnd 0.010172f
C5708 vdd.n3653 gnd 0.008187f
C5709 vdd.n3654 gnd 0.008187f
C5710 vdd.n3655 gnd 0.008187f
C5711 vdd.n3656 gnd 0.010172f
C5712 vdd.n3657 gnd 0.862789f
C5713 vdd.t162 gnd 0.519752f
C5714 vdd.n3658 gnd 0.6289f
C5715 vdd.n3659 gnd 0.753641f
C5716 vdd.n3660 gnd 0.010172f
C5717 vdd.n3661 gnd 0.008187f
C5718 vdd.n3662 gnd 0.008187f
C5719 vdd.n3663 gnd 0.008187f
C5720 vdd.n3664 gnd 0.010172f
C5721 vdd.n3665 gnd 0.576925f
C5722 vdd.t106 gnd 0.519752f
C5723 vdd.n3666 gnd 0.862789f
C5724 vdd.t205 gnd 0.519752f
C5725 vdd.n3667 gnd 0.639295f
C5726 vdd.n3668 gnd 0.010172f
C5727 vdd.n3669 gnd 0.008187f
C5728 vdd.n3670 gnd 0.007818f
C5729 vdd.n3671 gnd 0.599968f
C5730 vdd.n3672 gnd 2.9707f
C5731 a_n2804_13878.t29 gnd 0.194556f
C5732 a_n2804_13878.t25 gnd 0.194556f
C5733 a_n2804_13878.t31 gnd 0.194556f
C5734 a_n2804_13878.n0 gnd 1.53449f
C5735 a_n2804_13878.t8 gnd 0.194556f
C5736 a_n2804_13878.t20 gnd 0.194556f
C5737 a_n2804_13878.n1 gnd 1.53196f
C5738 a_n2804_13878.n2 gnd 1.37704f
C5739 a_n2804_13878.t12 gnd 0.194556f
C5740 a_n2804_13878.t22 gnd 0.194556f
C5741 a_n2804_13878.n3 gnd 1.53358f
C5742 a_n2804_13878.t27 gnd 0.194556f
C5743 a_n2804_13878.t17 gnd 0.194556f
C5744 a_n2804_13878.n4 gnd 1.53196f
C5745 a_n2804_13878.n5 gnd 2.14061f
C5746 a_n2804_13878.t23 gnd 0.194556f
C5747 a_n2804_13878.t16 gnd 0.194556f
C5748 a_n2804_13878.n6 gnd 1.53196f
C5749 a_n2804_13878.n7 gnd 1.04414f
C5750 a_n2804_13878.t10 gnd 0.194556f
C5751 a_n2804_13878.t13 gnd 0.194556f
C5752 a_n2804_13878.n8 gnd 1.53196f
C5753 a_n2804_13878.n9 gnd 1.04414f
C5754 a_n2804_13878.t26 gnd 0.194556f
C5755 a_n2804_13878.t11 gnd 0.194556f
C5756 a_n2804_13878.n10 gnd 1.53196f
C5757 a_n2804_13878.n11 gnd 1.04414f
C5758 a_n2804_13878.t21 gnd 0.194556f
C5759 a_n2804_13878.t9 gnd 0.194556f
C5760 a_n2804_13878.n12 gnd 1.53196f
C5761 a_n2804_13878.n13 gnd 4.90178f
C5762 a_n2804_13878.t6 gnd 1.82172f
C5763 a_n2804_13878.t1 gnd 0.194556f
C5764 a_n2804_13878.t3 gnd 0.194556f
C5765 a_n2804_13878.n14 gnd 1.37045f
C5766 a_n2804_13878.n15 gnd 1.53128f
C5767 a_n2804_13878.t2 gnd 1.81809f
C5768 a_n2804_13878.n16 gnd 0.770559f
C5769 a_n2804_13878.t5 gnd 1.81809f
C5770 a_n2804_13878.n17 gnd 0.770559f
C5771 a_n2804_13878.t4 gnd 0.194556f
C5772 a_n2804_13878.t0 gnd 0.194556f
C5773 a_n2804_13878.n18 gnd 1.37045f
C5774 a_n2804_13878.n19 gnd 0.778022f
C5775 a_n2804_13878.t7 gnd 1.81809f
C5776 a_n2804_13878.n20 gnd 2.85814f
C5777 a_n2804_13878.n21 gnd 3.74876f
C5778 a_n2804_13878.t15 gnd 0.194556f
C5779 a_n2804_13878.t24 gnd 0.194556f
C5780 a_n2804_13878.n22 gnd 1.53195f
C5781 a_n2804_13878.n23 gnd 2.50239f
C5782 a_n2804_13878.t28 gnd 0.194556f
C5783 a_n2804_13878.t14 gnd 0.194556f
C5784 a_n2804_13878.n24 gnd 1.53196f
C5785 a_n2804_13878.n25 gnd 0.678771f
C5786 a_n2804_13878.t18 gnd 0.194556f
C5787 a_n2804_13878.t19 gnd 0.194556f
C5788 a_n2804_13878.n26 gnd 1.53196f
C5789 a_n2804_13878.n27 gnd 0.678771f
C5790 a_n2804_13878.n28 gnd 0.678768f
C5791 a_n2804_13878.n29 gnd 1.53196f
C5792 a_n2804_13878.t30 gnd 0.194556f
C5793 a_n2982_13878.n0 gnd 2.53375f
C5794 a_n2982_13878.n1 gnd 3.78544f
C5795 a_n2982_13878.n2 gnd 3.42813f
C5796 a_n2982_13878.n3 gnd 0.20945f
C5797 a_n2982_13878.n4 gnd 0.20945f
C5798 a_n2982_13878.n5 gnd 0.791576f
C5799 a_n2982_13878.n6 gnd 0.20945f
C5800 a_n2982_13878.n7 gnd 0.971817f
C5801 a_n2982_13878.n8 gnd 0.20945f
C5802 a_n2982_13878.n9 gnd 0.20945f
C5803 a_n2982_13878.n10 gnd 0.458033f
C5804 a_n2982_13878.n11 gnd 0.20945f
C5805 a_n2982_13878.n12 gnd 0.27462f
C5806 a_n2982_13878.n13 gnd 0.90404f
C5807 a_n2982_13878.n14 gnd 0.198733f
C5808 a_n2982_13878.n15 gnd 0.146371f
C5809 a_n2982_13878.n16 gnd 0.230048f
C5810 a_n2982_13878.n17 gnd 0.177686f
C5811 a_n2982_13878.n18 gnd 0.198733f
C5812 a_n2982_13878.n19 gnd 1.32386f
C5813 a_n2982_13878.n20 gnd 0.146371f
C5814 a_n2982_13878.n21 gnd 0.956403f
C5815 a_n2982_13878.n22 gnd 0.20945f
C5816 a_n2982_13878.n23 gnd 0.73719f
C5817 a_n2982_13878.n24 gnd 0.20945f
C5818 a_n2982_13878.n25 gnd 0.20945f
C5819 a_n2982_13878.n26 gnd 0.477018f
C5820 a_n2982_13878.n27 gnd 0.27462f
C5821 a_n2982_13878.n28 gnd 0.20945f
C5822 a_n2982_13878.n29 gnd 0.529381f
C5823 a_n2982_13878.n30 gnd 0.20945f
C5824 a_n2982_13878.n31 gnd 0.20945f
C5825 a_n2982_13878.n32 gnd 0.931898f
C5826 a_n2982_13878.n33 gnd 0.27462f
C5827 a_n2982_13878.n34 gnd 3.08362f
C5828 a_n2982_13878.n35 gnd 0.27462f
C5829 a_n2982_13878.n36 gnd 1.72437f
C5830 a_n2982_13878.n37 gnd 1.16191f
C5831 a_n2982_13878.n38 gnd 2.32061f
C5832 a_n2982_13878.n39 gnd 2.12168f
C5833 a_n2982_13878.n40 gnd 1.16191f
C5834 a_n2982_13878.n41 gnd 1.72437f
C5835 a_n2982_13878.n42 gnd 0.008404f
C5836 a_n2982_13878.n43 gnd 4.05e-19
C5837 a_n2982_13878.n45 gnd 0.008109f
C5838 a_n2982_13878.n46 gnd 0.011792f
C5839 a_n2982_13878.n47 gnd 0.007801f
C5840 a_n2982_13878.n49 gnd 0.277816f
C5841 a_n2982_13878.n50 gnd 0.008404f
C5842 a_n2982_13878.n51 gnd 4.05e-19
C5843 a_n2982_13878.n53 gnd 0.008109f
C5844 a_n2982_13878.n54 gnd 0.011792f
C5845 a_n2982_13878.n55 gnd 0.007801f
C5846 a_n2982_13878.n57 gnd 0.277816f
C5847 a_n2982_13878.n58 gnd 0.008109f
C5848 a_n2982_13878.n59 gnd 0.276683f
C5849 a_n2982_13878.n60 gnd 0.008109f
C5850 a_n2982_13878.n61 gnd 0.276683f
C5851 a_n2982_13878.n62 gnd 0.008109f
C5852 a_n2982_13878.n63 gnd 0.276683f
C5853 a_n2982_13878.n64 gnd 0.008109f
C5854 a_n2982_13878.n65 gnd 0.276683f
C5855 a_n2982_13878.n66 gnd 0.008404f
C5856 a_n2982_13878.n67 gnd 4.05e-19
C5857 a_n2982_13878.n69 gnd 0.008109f
C5858 a_n2982_13878.n70 gnd 0.011792f
C5859 a_n2982_13878.n71 gnd 0.007801f
C5860 a_n2982_13878.n73 gnd 0.277816f
C5861 a_n2982_13878.n74 gnd 0.277816f
C5862 a_n2982_13878.n76 gnd 0.007801f
C5863 a_n2982_13878.n77 gnd 0.011792f
C5864 a_n2982_13878.n78 gnd 0.008109f
C5865 a_n2982_13878.n80 gnd 4.05e-19
C5866 a_n2982_13878.n81 gnd 0.008404f
C5867 a_n2982_13878.n82 gnd 0.104725f
C5868 a_n2982_13878.t31 gnd 0.145277f
C5869 a_n2982_13878.t50 gnd 0.686627f
C5870 a_n2982_13878.t38 gnd 0.675756f
C5871 a_n2982_13878.t52 gnd 0.675756f
C5872 a_n2982_13878.t44 gnd 0.675756f
C5873 a_n2982_13878.n83 gnd 0.293584f
C5874 a_n2982_13878.t34 gnd 0.675756f
C5875 a_n2982_13878.t58 gnd 0.675756f
C5876 a_n2982_13878.t46 gnd 0.675756f
C5877 a_n2982_13878.n84 gnd 0.297105f
C5878 a_n2982_13878.t28 gnd 0.675756f
C5879 a_n2982_13878.t56 gnd 0.675756f
C5880 a_n2982_13878.t16 gnd 0.675756f
C5881 a_n2982_13878.n85 gnd 0.293009f
C5882 a_n2982_13878.t30 gnd 0.675756f
C5883 a_n2982_13878.t26 gnd 0.689824f
C5884 a_n2982_13878.t102 gnd 0.689824f
C5885 a_n2982_13878.t79 gnd 0.675756f
C5886 a_n2982_13878.t84 gnd 0.675756f
C5887 a_n2982_13878.t72 gnd 0.675756f
C5888 a_n2982_13878.n86 gnd 0.296971f
C5889 a_n2982_13878.t89 gnd 0.675756f
C5890 a_n2982_13878.t98 gnd 0.675756f
C5891 a_n2982_13878.t99 gnd 0.675756f
C5892 a_n2982_13878.n87 gnd 0.293332f
C5893 a_n2982_13878.t66 gnd 0.675756f
C5894 a_n2982_13878.t81 gnd 0.675756f
C5895 a_n2982_13878.t69 gnd 0.675756f
C5896 a_n2982_13878.n88 gnd 0.29709f
C5897 a_n2982_13878.t76 gnd 0.675756f
C5898 a_n2982_13878.t95 gnd 0.686627f
C5899 a_n2982_13878.t49 gnd 1.3603f
C5900 a_n2982_13878.t21 gnd 0.145277f
C5901 a_n2982_13878.t61 gnd 0.145277f
C5902 a_n2982_13878.n89 gnd 1.02333f
C5903 a_n2982_13878.t41 gnd 0.145277f
C5904 a_n2982_13878.t25 gnd 0.145277f
C5905 a_n2982_13878.n90 gnd 1.02333f
C5906 a_n2982_13878.t43 gnd 0.145277f
C5907 a_n2982_13878.t33 gnd 0.145277f
C5908 a_n2982_13878.n91 gnd 1.02333f
C5909 a_n2982_13878.t63 gnd 0.145277f
C5910 a_n2982_13878.t55 gnd 0.145277f
C5911 a_n2982_13878.n92 gnd 1.02333f
C5912 a_n2982_13878.t23 gnd 0.145277f
C5913 a_n2982_13878.t19 gnd 0.145277f
C5914 a_n2982_13878.n93 gnd 1.02333f
C5915 a_n2982_13878.t37 gnd 1.35758f
C5916 a_n2982_13878.t22 gnd 0.675756f
C5917 a_n2982_13878.n94 gnd 0.29709f
C5918 a_n2982_13878.t18 gnd 0.675756f
C5919 a_n2982_13878.t62 gnd 0.675756f
C5920 a_n2982_13878.n95 gnd 0.288167f
C5921 a_n2982_13878.t24 gnd 0.675756f
C5922 a_n2982_13878.n96 gnd 0.299644f
C5923 a_n2982_13878.t42 gnd 0.675756f
C5924 a_n2982_13878.t60 gnd 0.675756f
C5925 a_n2982_13878.n97 gnd 0.293009f
C5926 a_n2982_13878.t48 gnd 0.689824f
C5927 a_n2982_13878.t78 gnd 0.675756f
C5928 a_n2982_13878.n98 gnd 0.29709f
C5929 a_n2982_13878.t87 gnd 0.675756f
C5930 a_n2982_13878.t93 gnd 0.675756f
C5931 a_n2982_13878.n99 gnd 0.288167f
C5932 a_n2982_13878.t97 gnd 0.675756f
C5933 a_n2982_13878.n100 gnd 0.299644f
C5934 a_n2982_13878.t68 gnd 0.675756f
C5935 a_n2982_13878.t71 gnd 0.675756f
C5936 a_n2982_13878.n101 gnd 0.293009f
C5937 a_n2982_13878.t101 gnd 0.689824f
C5938 a_n2982_13878.t70 gnd 0.675756f
C5939 a_n2982_13878.n102 gnd 0.299205f
C5940 a_n2982_13878.t96 gnd 0.675756f
C5941 a_n2982_13878.n103 gnd 0.296971f
C5942 a_n2982_13878.n104 gnd 0.297105f
C5943 a_n2982_13878.t92 gnd 0.675756f
C5944 a_n2982_13878.n105 gnd 0.293332f
C5945 a_n2982_13878.t65 gnd 0.675756f
C5946 a_n2982_13878.n106 gnd 0.293584f
C5947 a_n2982_13878.n107 gnd 0.299206f
C5948 a_n2982_13878.t67 gnd 0.686627f
C5949 a_n2982_13878.t20 gnd 0.675756f
C5950 a_n2982_13878.n108 gnd 0.299205f
C5951 a_n2982_13878.t40 gnd 0.675756f
C5952 a_n2982_13878.n109 gnd 0.296971f
C5953 a_n2982_13878.n110 gnd 0.297105f
C5954 a_n2982_13878.t32 gnd 0.675756f
C5955 a_n2982_13878.n111 gnd 0.293332f
C5956 a_n2982_13878.t54 gnd 0.675756f
C5957 a_n2982_13878.n112 gnd 0.293584f
C5958 a_n2982_13878.n113 gnd 0.299206f
C5959 a_n2982_13878.t36 gnd 0.686627f
C5960 a_n2982_13878.n114 gnd 1.30834f
C5961 a_n2982_13878.t75 gnd 0.675756f
C5962 a_n2982_13878.n115 gnd 0.293332f
C5963 a_n2982_13878.t83 gnd 0.675756f
C5964 a_n2982_13878.n116 gnd 0.293332f
C5965 a_n2982_13878.t73 gnd 0.675756f
C5966 a_n2982_13878.n117 gnd 0.293332f
C5967 a_n2982_13878.t88 gnd 0.675756f
C5968 a_n2982_13878.n118 gnd 0.293332f
C5969 a_n2982_13878.t77 gnd 0.675756f
C5970 a_n2982_13878.n119 gnd 0.288005f
C5971 a_n2982_13878.t103 gnd 0.675756f
C5972 a_n2982_13878.n120 gnd 0.297105f
C5973 a_n2982_13878.t80 gnd 0.687079f
C5974 a_n2982_13878.t90 gnd 0.675756f
C5975 a_n2982_13878.n121 gnd 0.288005f
C5976 a_n2982_13878.t74 gnd 0.675756f
C5977 a_n2982_13878.n122 gnd 0.297105f
C5978 a_n2982_13878.t85 gnd 0.687079f
C5979 a_n2982_13878.t94 gnd 0.675756f
C5980 a_n2982_13878.n123 gnd 0.288005f
C5981 a_n2982_13878.t82 gnd 0.675756f
C5982 a_n2982_13878.n124 gnd 0.297105f
C5983 a_n2982_13878.t100 gnd 0.687079f
C5984 a_n2982_13878.t86 gnd 0.675756f
C5985 a_n2982_13878.n125 gnd 0.288005f
C5986 a_n2982_13878.t64 gnd 0.675756f
C5987 a_n2982_13878.n126 gnd 0.297105f
C5988 a_n2982_13878.t91 gnd 0.687079f
C5989 a_n2982_13878.n127 gnd 1.64574f
C5990 a_n2982_13878.n128 gnd 0.299206f
C5991 a_n2982_13878.n129 gnd 0.293584f
C5992 a_n2982_13878.n130 gnd 0.288167f
C5993 a_n2982_13878.n131 gnd 0.297105f
C5994 a_n2982_13878.n132 gnd 0.299644f
C5995 a_n2982_13878.n133 gnd 0.293009f
C5996 a_n2982_13878.n134 gnd 0.299205f
C5997 a_n2982_13878.t8 gnd 0.112993f
C5998 a_n2982_13878.t3 gnd 0.112993f
C5999 a_n2982_13878.n135 gnd 1.00066f
C6000 a_n2982_13878.t2 gnd 0.112993f
C6001 a_n2982_13878.t1 gnd 0.112993f
C6002 a_n2982_13878.n136 gnd 0.998444f
C6003 a_n2982_13878.t11 gnd 0.112993f
C6004 a_n2982_13878.t10 gnd 0.112993f
C6005 a_n2982_13878.n137 gnd 1.00066f
C6006 a_n2982_13878.t14 gnd 0.112993f
C6007 a_n2982_13878.t5 gnd 0.112993f
C6008 a_n2982_13878.n138 gnd 0.998444f
C6009 a_n2982_13878.t9 gnd 0.112993f
C6010 a_n2982_13878.t12 gnd 0.112993f
C6011 a_n2982_13878.n139 gnd 0.998444f
C6012 a_n2982_13878.t6 gnd 0.112993f
C6013 a_n2982_13878.t13 gnd 0.112993f
C6014 a_n2982_13878.n140 gnd 0.998444f
C6015 a_n2982_13878.t4 gnd 0.112993f
C6016 a_n2982_13878.t7 gnd 0.112993f
C6017 a_n2982_13878.n141 gnd 1.00066f
C6018 a_n2982_13878.t0 gnd 0.112993f
C6019 a_n2982_13878.t15 gnd 0.112993f
C6020 a_n2982_13878.n142 gnd 0.998444f
C6021 a_n2982_13878.n143 gnd 0.299205f
C6022 a_n2982_13878.n144 gnd 0.296971f
C6023 a_n2982_13878.n145 gnd 0.299644f
C6024 a_n2982_13878.n146 gnd 0.293332f
C6025 a_n2982_13878.n147 gnd 0.288167f
C6026 a_n2982_13878.n148 gnd 0.29709f
C6027 a_n2982_13878.n149 gnd 0.299206f
C6028 a_n2982_13878.n150 gnd 0.994805f
C6029 a_n2982_13878.t51 gnd 1.35759f
C6030 a_n2982_13878.t39 gnd 0.145277f
C6031 a_n2982_13878.t53 gnd 0.145277f
C6032 a_n2982_13878.n151 gnd 1.02333f
C6033 a_n2982_13878.t45 gnd 0.145277f
C6034 a_n2982_13878.t35 gnd 0.145277f
C6035 a_n2982_13878.n152 gnd 1.02333f
C6036 a_n2982_13878.t59 gnd 0.145277f
C6037 a_n2982_13878.t47 gnd 0.145277f
C6038 a_n2982_13878.n153 gnd 1.02333f
C6039 a_n2982_13878.t29 gnd 0.145277f
C6040 a_n2982_13878.t57 gnd 0.145277f
C6041 a_n2982_13878.n154 gnd 1.02333f
C6042 a_n2982_13878.t27 gnd 1.3603f
C6043 a_n2982_13878.n155 gnd 1.02333f
C6044 a_n2982_13878.t17 gnd 0.145277f
C6045 a_n9628_8799.t30 gnd 0.112803f
C6046 a_n9628_8799.t35 gnd 0.145033f
C6047 a_n9628_8799.t7 gnd 0.145033f
C6048 a_n9628_8799.n0 gnd 1.14389f
C6049 a_n9628_8799.t0 gnd 0.145033f
C6050 a_n9628_8799.t17 gnd 0.145033f
C6051 a_n9628_8799.n1 gnd 1.14201f
C6052 a_n9628_8799.n2 gnd 1.02653f
C6053 a_n9628_8799.t37 gnd 0.145033f
C6054 a_n9628_8799.t10 gnd 0.145033f
C6055 a_n9628_8799.n3 gnd 1.14201f
C6056 a_n9628_8799.n4 gnd 0.505994f
C6057 a_n9628_8799.t18 gnd 0.145033f
C6058 a_n9628_8799.t8 gnd 0.145033f
C6059 a_n9628_8799.n5 gnd 1.14201f
C6060 a_n9628_8799.n6 gnd 0.505994f
C6061 a_n9628_8799.t9 gnd 0.145033f
C6062 a_n9628_8799.t1 gnd 0.145033f
C6063 a_n9628_8799.n7 gnd 1.14201f
C6064 a_n9628_8799.n8 gnd 0.505994f
C6065 a_n9628_8799.t39 gnd 0.145033f
C6066 a_n9628_8799.t36 gnd 0.145033f
C6067 a_n9628_8799.n9 gnd 1.14201f
C6068 a_n9628_8799.n10 gnd 3.67671f
C6069 a_n9628_8799.t15 gnd 0.145033f
C6070 a_n9628_8799.t3 gnd 0.145033f
C6071 a_n9628_8799.n11 gnd 1.1439f
C6072 a_n9628_8799.t6 gnd 0.145033f
C6073 a_n9628_8799.t13 gnd 0.145033f
C6074 a_n9628_8799.n12 gnd 1.14201f
C6075 a_n9628_8799.n13 gnd 1.02653f
C6076 a_n9628_8799.t14 gnd 0.145033f
C6077 a_n9628_8799.t5 gnd 0.145033f
C6078 a_n9628_8799.n14 gnd 1.14201f
C6079 a_n9628_8799.n15 gnd 0.505994f
C6080 a_n9628_8799.t38 gnd 0.145033f
C6081 a_n9628_8799.t16 gnd 0.145033f
C6082 a_n9628_8799.n16 gnd 1.14201f
C6083 a_n9628_8799.n17 gnd 0.505994f
C6084 a_n9628_8799.t4 gnd 0.145033f
C6085 a_n9628_8799.t2 gnd 0.145033f
C6086 a_n9628_8799.n18 gnd 1.14201f
C6087 a_n9628_8799.n19 gnd 0.505994f
C6088 a_n9628_8799.t12 gnd 0.145033f
C6089 a_n9628_8799.t11 gnd 0.145033f
C6090 a_n9628_8799.n20 gnd 1.14201f
C6091 a_n9628_8799.n21 gnd 2.55267f
C6092 a_n9628_8799.n22 gnd 7.67608f
C6093 a_n9628_8799.n23 gnd 0.052275f
C6094 a_n9628_8799.t86 gnd 0.601374f
C6095 a_n9628_8799.n24 gnd 0.268585f
C6096 a_n9628_8799.n25 gnd 0.052275f
C6097 a_n9628_8799.n26 gnd 0.011862f
C6098 a_n9628_8799.t122 gnd 0.601374f
C6099 a_n9628_8799.n27 gnd 0.052275f
C6100 a_n9628_8799.t143 gnd 0.601374f
C6101 a_n9628_8799.n28 gnd 0.265523f
C6102 a_n9628_8799.t144 gnd 0.601374f
C6103 a_n9628_8799.n29 gnd 0.052275f
C6104 a_n9628_8799.t72 gnd 0.601374f
C6105 a_n9628_8799.n30 gnd 0.265846f
C6106 a_n9628_8799.n31 gnd 0.052275f
C6107 a_n9628_8799.n32 gnd 0.011862f
C6108 a_n9628_8799.t112 gnd 0.601374f
C6109 a_n9628_8799.n33 gnd 0.052275f
C6110 a_n9628_8799.t120 gnd 0.601374f
C6111 a_n9628_8799.n34 gnd 0.268585f
C6112 a_n9628_8799.n35 gnd 0.052275f
C6113 a_n9628_8799.n36 gnd 0.011862f
C6114 a_n9628_8799.t48 gnd 0.601374f
C6115 a_n9628_8799.n37 gnd 0.16515f
C6116 a_n9628_8799.t91 gnd 0.601374f
C6117 a_n9628_8799.t89 gnd 0.612756f
C6118 a_n9628_8799.n38 gnd 0.2521f
C6119 a_n9628_8799.n39 gnd 0.264879f
C6120 a_n9628_8799.n40 gnd 0.011862f
C6121 a_n9628_8799.t123 gnd 0.601374f
C6122 a_n9628_8799.n41 gnd 0.268585f
C6123 a_n9628_8799.n42 gnd 0.052275f
C6124 a_n9628_8799.n43 gnd 0.052275f
C6125 a_n9628_8799.n44 gnd 0.052275f
C6126 a_n9628_8799.n45 gnd 0.26649f
C6127 a_n9628_8799.t88 gnd 0.601374f
C6128 a_n9628_8799.n46 gnd 0.265201f
C6129 a_n9628_8799.n47 gnd 0.011862f
C6130 a_n9628_8799.n48 gnd 0.052275f
C6131 a_n9628_8799.n49 gnd 0.052275f
C6132 a_n9628_8799.n50 gnd 0.052275f
C6133 a_n9628_8799.n51 gnd 0.011862f
C6134 a_n9628_8799.t42 gnd 0.601374f
C6135 a_n9628_8799.n52 gnd 0.266168f
C6136 a_n9628_8799.t74 gnd 0.601374f
C6137 a_n9628_8799.n53 gnd 0.265523f
C6138 a_n9628_8799.n54 gnd 0.052275f
C6139 a_n9628_8799.n55 gnd 0.052275f
C6140 a_n9628_8799.n56 gnd 0.052275f
C6141 a_n9628_8799.n57 gnd 0.268585f
C6142 a_n9628_8799.n58 gnd 0.011862f
C6143 a_n9628_8799.t147 gnd 0.601374f
C6144 a_n9628_8799.n59 gnd 0.265846f
C6145 a_n9628_8799.n60 gnd 0.052275f
C6146 a_n9628_8799.n61 gnd 0.052275f
C6147 a_n9628_8799.n62 gnd 0.052275f
C6148 a_n9628_8799.n63 gnd 0.011862f
C6149 a_n9628_8799.t108 gnd 0.601374f
C6150 a_n9628_8799.n64 gnd 0.268585f
C6151 a_n9628_8799.n65 gnd 0.011862f
C6152 a_n9628_8799.n66 gnd 0.052275f
C6153 a_n9628_8799.n67 gnd 0.052275f
C6154 a_n9628_8799.n68 gnd 0.052275f
C6155 a_n9628_8799.n69 gnd 0.266168f
C6156 a_n9628_8799.n70 gnd 0.011862f
C6157 a_n9628_8799.t90 gnd 0.601374f
C6158 a_n9628_8799.n71 gnd 0.268585f
C6159 a_n9628_8799.n72 gnd 0.052275f
C6160 a_n9628_8799.n73 gnd 0.052275f
C6161 a_n9628_8799.n74 gnd 0.052275f
C6162 a_n9628_8799.n75 gnd 0.265201f
C6163 a_n9628_8799.t142 gnd 0.601374f
C6164 a_n9628_8799.n76 gnd 0.26649f
C6165 a_n9628_8799.n77 gnd 0.011862f
C6166 a_n9628_8799.n78 gnd 0.052275f
C6167 a_n9628_8799.n79 gnd 0.052275f
C6168 a_n9628_8799.n80 gnd 0.052275f
C6169 a_n9628_8799.n81 gnd 0.011862f
C6170 a_n9628_8799.t87 gnd 0.601374f
C6171 a_n9628_8799.n82 gnd 0.264879f
C6172 a_n9628_8799.t119 gnd 0.601374f
C6173 a_n9628_8799.n83 gnd 0.263106f
C6174 a_n9628_8799.n84 gnd 0.296383f
C6175 a_n9628_8799.n85 gnd 0.052275f
C6176 a_n9628_8799.t97 gnd 0.601374f
C6177 a_n9628_8799.n86 gnd 0.268585f
C6178 a_n9628_8799.n87 gnd 0.052275f
C6179 a_n9628_8799.n88 gnd 0.011862f
C6180 a_n9628_8799.t136 gnd 0.601374f
C6181 a_n9628_8799.n89 gnd 0.052275f
C6182 a_n9628_8799.t155 gnd 0.601374f
C6183 a_n9628_8799.n90 gnd 0.265523f
C6184 a_n9628_8799.t157 gnd 0.601374f
C6185 a_n9628_8799.n91 gnd 0.052275f
C6186 a_n9628_8799.t81 gnd 0.601374f
C6187 a_n9628_8799.n92 gnd 0.265846f
C6188 a_n9628_8799.n93 gnd 0.052275f
C6189 a_n9628_8799.n94 gnd 0.011862f
C6190 a_n9628_8799.t125 gnd 0.601374f
C6191 a_n9628_8799.n95 gnd 0.052275f
C6192 a_n9628_8799.t132 gnd 0.601374f
C6193 a_n9628_8799.n96 gnd 0.268585f
C6194 a_n9628_8799.n97 gnd 0.052275f
C6195 a_n9628_8799.n98 gnd 0.011862f
C6196 a_n9628_8799.t60 gnd 0.601374f
C6197 a_n9628_8799.n99 gnd 0.16515f
C6198 a_n9628_8799.t104 gnd 0.601374f
C6199 a_n9628_8799.t102 gnd 0.612756f
C6200 a_n9628_8799.n100 gnd 0.2521f
C6201 a_n9628_8799.n101 gnd 0.264879f
C6202 a_n9628_8799.n102 gnd 0.011862f
C6203 a_n9628_8799.t140 gnd 0.601374f
C6204 a_n9628_8799.n103 gnd 0.268585f
C6205 a_n9628_8799.n104 gnd 0.052275f
C6206 a_n9628_8799.n105 gnd 0.052275f
C6207 a_n9628_8799.n106 gnd 0.052275f
C6208 a_n9628_8799.n107 gnd 0.26649f
C6209 a_n9628_8799.t98 gnd 0.601374f
C6210 a_n9628_8799.n108 gnd 0.265201f
C6211 a_n9628_8799.n109 gnd 0.011862f
C6212 a_n9628_8799.n110 gnd 0.052275f
C6213 a_n9628_8799.n111 gnd 0.052275f
C6214 a_n9628_8799.n112 gnd 0.052275f
C6215 a_n9628_8799.n113 gnd 0.011862f
C6216 a_n9628_8799.t56 gnd 0.601374f
C6217 a_n9628_8799.n114 gnd 0.266168f
C6218 a_n9628_8799.t84 gnd 0.601374f
C6219 a_n9628_8799.n115 gnd 0.265523f
C6220 a_n9628_8799.n116 gnd 0.052275f
C6221 a_n9628_8799.n117 gnd 0.052275f
C6222 a_n9628_8799.n118 gnd 0.052275f
C6223 a_n9628_8799.n119 gnd 0.268585f
C6224 a_n9628_8799.n120 gnd 0.011862f
C6225 a_n9628_8799.t159 gnd 0.601374f
C6226 a_n9628_8799.n121 gnd 0.265846f
C6227 a_n9628_8799.n122 gnd 0.052275f
C6228 a_n9628_8799.n123 gnd 0.052275f
C6229 a_n9628_8799.n124 gnd 0.052275f
C6230 a_n9628_8799.n125 gnd 0.011862f
C6231 a_n9628_8799.t121 gnd 0.601374f
C6232 a_n9628_8799.n126 gnd 0.268585f
C6233 a_n9628_8799.n127 gnd 0.011862f
C6234 a_n9628_8799.n128 gnd 0.052275f
C6235 a_n9628_8799.n129 gnd 0.052275f
C6236 a_n9628_8799.n130 gnd 0.052275f
C6237 a_n9628_8799.n131 gnd 0.266168f
C6238 a_n9628_8799.n132 gnd 0.011862f
C6239 a_n9628_8799.t103 gnd 0.601374f
C6240 a_n9628_8799.n133 gnd 0.268585f
C6241 a_n9628_8799.n134 gnd 0.052275f
C6242 a_n9628_8799.n135 gnd 0.052275f
C6243 a_n9628_8799.n136 gnd 0.052275f
C6244 a_n9628_8799.n137 gnd 0.265201f
C6245 a_n9628_8799.t154 gnd 0.601374f
C6246 a_n9628_8799.n138 gnd 0.26649f
C6247 a_n9628_8799.n139 gnd 0.011862f
C6248 a_n9628_8799.n140 gnd 0.052275f
C6249 a_n9628_8799.n141 gnd 0.052275f
C6250 a_n9628_8799.n142 gnd 0.052275f
C6251 a_n9628_8799.n143 gnd 0.011862f
C6252 a_n9628_8799.t99 gnd 0.601374f
C6253 a_n9628_8799.n144 gnd 0.264879f
C6254 a_n9628_8799.t133 gnd 0.601374f
C6255 a_n9628_8799.n145 gnd 0.263106f
C6256 a_n9628_8799.n146 gnd 0.130296f
C6257 a_n9628_8799.n147 gnd 0.904082f
C6258 a_n9628_8799.n148 gnd 0.052275f
C6259 a_n9628_8799.t63 gnd 0.601374f
C6260 a_n9628_8799.n149 gnd 0.268585f
C6261 a_n9628_8799.n150 gnd 0.052275f
C6262 a_n9628_8799.n151 gnd 0.011862f
C6263 a_n9628_8799.t82 gnd 0.601374f
C6264 a_n9628_8799.n152 gnd 0.052275f
C6265 a_n9628_8799.t116 gnd 0.601374f
C6266 a_n9628_8799.n153 gnd 0.265523f
C6267 a_n9628_8799.t96 gnd 0.601374f
C6268 a_n9628_8799.n154 gnd 0.052275f
C6269 a_n9628_8799.t100 gnd 0.601374f
C6270 a_n9628_8799.n155 gnd 0.265846f
C6271 a_n9628_8799.n156 gnd 0.052275f
C6272 a_n9628_8799.n157 gnd 0.011862f
C6273 a_n9628_8799.t127 gnd 0.601374f
C6274 a_n9628_8799.n158 gnd 0.052275f
C6275 a_n9628_8799.t43 gnd 0.601374f
C6276 a_n9628_8799.n159 gnd 0.268585f
C6277 a_n9628_8799.n160 gnd 0.052275f
C6278 a_n9628_8799.n161 gnd 0.011862f
C6279 a_n9628_8799.t69 gnd 0.601374f
C6280 a_n9628_8799.n162 gnd 0.16515f
C6281 a_n9628_8799.t52 gnd 0.601374f
C6282 a_n9628_8799.t73 gnd 0.612756f
C6283 a_n9628_8799.n163 gnd 0.2521f
C6284 a_n9628_8799.n164 gnd 0.264879f
C6285 a_n9628_8799.n165 gnd 0.011862f
C6286 a_n9628_8799.t114 gnd 0.601374f
C6287 a_n9628_8799.n166 gnd 0.268585f
C6288 a_n9628_8799.n167 gnd 0.052275f
C6289 a_n9628_8799.n168 gnd 0.052275f
C6290 a_n9628_8799.n169 gnd 0.052275f
C6291 a_n9628_8799.n170 gnd 0.26649f
C6292 a_n9628_8799.t92 gnd 0.601374f
C6293 a_n9628_8799.n171 gnd 0.265201f
C6294 a_n9628_8799.n172 gnd 0.011862f
C6295 a_n9628_8799.n173 gnd 0.052275f
C6296 a_n9628_8799.n174 gnd 0.052275f
C6297 a_n9628_8799.n175 gnd 0.052275f
C6298 a_n9628_8799.n176 gnd 0.011862f
C6299 a_n9628_8799.t109 gnd 0.601374f
C6300 a_n9628_8799.n177 gnd 0.266168f
C6301 a_n9628_8799.t61 gnd 0.601374f
C6302 a_n9628_8799.n178 gnd 0.265523f
C6303 a_n9628_8799.n179 gnd 0.052275f
C6304 a_n9628_8799.n180 gnd 0.052275f
C6305 a_n9628_8799.n181 gnd 0.052275f
C6306 a_n9628_8799.n182 gnd 0.268585f
C6307 a_n9628_8799.n183 gnd 0.011862f
C6308 a_n9628_8799.t77 gnd 0.601374f
C6309 a_n9628_8799.n184 gnd 0.265846f
C6310 a_n9628_8799.n185 gnd 0.052275f
C6311 a_n9628_8799.n186 gnd 0.052275f
C6312 a_n9628_8799.n187 gnd 0.052275f
C6313 a_n9628_8799.n188 gnd 0.011862f
C6314 a_n9628_8799.t53 gnd 0.601374f
C6315 a_n9628_8799.n189 gnd 0.268585f
C6316 a_n9628_8799.n190 gnd 0.011862f
C6317 a_n9628_8799.n191 gnd 0.052275f
C6318 a_n9628_8799.n192 gnd 0.052275f
C6319 a_n9628_8799.n193 gnd 0.052275f
C6320 a_n9628_8799.n194 gnd 0.266168f
C6321 a_n9628_8799.n195 gnd 0.011862f
C6322 a_n9628_8799.t135 gnd 0.601374f
C6323 a_n9628_8799.n196 gnd 0.268585f
C6324 a_n9628_8799.n197 gnd 0.052275f
C6325 a_n9628_8799.n198 gnd 0.052275f
C6326 a_n9628_8799.n199 gnd 0.052275f
C6327 a_n9628_8799.n200 gnd 0.265201f
C6328 a_n9628_8799.t145 gnd 0.601374f
C6329 a_n9628_8799.n201 gnd 0.26649f
C6330 a_n9628_8799.n202 gnd 0.011862f
C6331 a_n9628_8799.n203 gnd 0.052275f
C6332 a_n9628_8799.n204 gnd 0.052275f
C6333 a_n9628_8799.n205 gnd 0.052275f
C6334 a_n9628_8799.n206 gnd 0.011862f
C6335 a_n9628_8799.t40 gnd 0.601374f
C6336 a_n9628_8799.n207 gnd 0.264879f
C6337 a_n9628_8799.t105 gnd 0.601374f
C6338 a_n9628_8799.n208 gnd 0.263106f
C6339 a_n9628_8799.n209 gnd 0.130296f
C6340 a_n9628_8799.n210 gnd 1.81909f
C6341 a_n9628_8799.n211 gnd 0.052275f
C6342 a_n9628_8799.t47 gnd 0.601374f
C6343 a_n9628_8799.t45 gnd 0.601374f
C6344 a_n9628_8799.t131 gnd 0.601374f
C6345 a_n9628_8799.n212 gnd 0.268585f
C6346 a_n9628_8799.n213 gnd 0.052275f
C6347 a_n9628_8799.t67 gnd 0.601374f
C6348 a_n9628_8799.t50 gnd 0.601374f
C6349 a_n9628_8799.n214 gnd 0.052275f
C6350 a_n9628_8799.t138 gnd 0.601374f
C6351 a_n9628_8799.n215 gnd 0.268585f
C6352 a_n9628_8799.n216 gnd 0.052275f
C6353 a_n9628_8799.t93 gnd 0.601374f
C6354 a_n9628_8799.t68 gnd 0.601374f
C6355 a_n9628_8799.n217 gnd 0.052275f
C6356 a_n9628_8799.t156 gnd 0.601374f
C6357 a_n9628_8799.n218 gnd 0.268585f
C6358 a_n9628_8799.n219 gnd 0.052275f
C6359 a_n9628_8799.t111 gnd 0.601374f
C6360 a_n9628_8799.t71 gnd 0.601374f
C6361 a_n9628_8799.n220 gnd 0.052275f
C6362 a_n9628_8799.t150 gnd 0.601374f
C6363 a_n9628_8799.n221 gnd 0.268585f
C6364 a_n9628_8799.n222 gnd 0.052275f
C6365 a_n9628_8799.t113 gnd 0.601374f
C6366 a_n9628_8799.t85 gnd 0.601374f
C6367 a_n9628_8799.n223 gnd 0.052275f
C6368 a_n9628_8799.t46 gnd 0.601374f
C6369 a_n9628_8799.n224 gnd 0.268585f
C6370 a_n9628_8799.n225 gnd 0.052275f
C6371 a_n9628_8799.t134 gnd 0.601374f
C6372 a_n9628_8799.t115 gnd 0.601374f
C6373 a_n9628_8799.n226 gnd 0.052275f
C6374 a_n9628_8799.t51 gnd 0.601374f
C6375 a_n9628_8799.n227 gnd 0.268585f
C6376 a_n9628_8799.t137 gnd 0.612756f
C6377 a_n9628_8799.n228 gnd 0.2521f
C6378 a_n9628_8799.t141 gnd 0.601374f
C6379 a_n9628_8799.n229 gnd 0.264879f
C6380 a_n9628_8799.n230 gnd 0.011862f
C6381 a_n9628_8799.n231 gnd 0.16515f
C6382 a_n9628_8799.n232 gnd 0.052275f
C6383 a_n9628_8799.n233 gnd 0.052275f
C6384 a_n9628_8799.n234 gnd 0.011862f
C6385 a_n9628_8799.n235 gnd 0.26649f
C6386 a_n9628_8799.n236 gnd 0.265201f
C6387 a_n9628_8799.n237 gnd 0.011862f
C6388 a_n9628_8799.n238 gnd 0.052275f
C6389 a_n9628_8799.n239 gnd 0.052275f
C6390 a_n9628_8799.n240 gnd 0.052275f
C6391 a_n9628_8799.n241 gnd 0.011862f
C6392 a_n9628_8799.n242 gnd 0.266168f
C6393 a_n9628_8799.n243 gnd 0.265523f
C6394 a_n9628_8799.n244 gnd 0.011862f
C6395 a_n9628_8799.n245 gnd 0.052275f
C6396 a_n9628_8799.n246 gnd 0.052275f
C6397 a_n9628_8799.n247 gnd 0.052275f
C6398 a_n9628_8799.n248 gnd 0.011862f
C6399 a_n9628_8799.n249 gnd 0.265846f
C6400 a_n9628_8799.n250 gnd 0.265846f
C6401 a_n9628_8799.n251 gnd 0.011862f
C6402 a_n9628_8799.n252 gnd 0.052275f
C6403 a_n9628_8799.n253 gnd 0.052275f
C6404 a_n9628_8799.n254 gnd 0.052275f
C6405 a_n9628_8799.n255 gnd 0.011862f
C6406 a_n9628_8799.n256 gnd 0.265523f
C6407 a_n9628_8799.n257 gnd 0.266168f
C6408 a_n9628_8799.n258 gnd 0.011862f
C6409 a_n9628_8799.n259 gnd 0.052275f
C6410 a_n9628_8799.n260 gnd 0.052275f
C6411 a_n9628_8799.n261 gnd 0.052275f
C6412 a_n9628_8799.n262 gnd 0.011862f
C6413 a_n9628_8799.n263 gnd 0.265201f
C6414 a_n9628_8799.n264 gnd 0.26649f
C6415 a_n9628_8799.n265 gnd 0.011862f
C6416 a_n9628_8799.n266 gnd 0.052275f
C6417 a_n9628_8799.n267 gnd 0.052275f
C6418 a_n9628_8799.n268 gnd 0.052275f
C6419 a_n9628_8799.n269 gnd 0.011862f
C6420 a_n9628_8799.n270 gnd 0.264879f
C6421 a_n9628_8799.n271 gnd 0.263106f
C6422 a_n9628_8799.n272 gnd 0.296383f
C6423 a_n9628_8799.n273 gnd 0.052275f
C6424 a_n9628_8799.t58 gnd 0.601374f
C6425 a_n9628_8799.t57 gnd 0.601374f
C6426 a_n9628_8799.t148 gnd 0.601374f
C6427 a_n9628_8799.n274 gnd 0.268585f
C6428 a_n9628_8799.n275 gnd 0.052275f
C6429 a_n9628_8799.t76 gnd 0.601374f
C6430 a_n9628_8799.t65 gnd 0.601374f
C6431 a_n9628_8799.n276 gnd 0.052275f
C6432 a_n9628_8799.t151 gnd 0.601374f
C6433 a_n9628_8799.n277 gnd 0.268585f
C6434 a_n9628_8799.n278 gnd 0.052275f
C6435 a_n9628_8799.t107 gnd 0.601374f
C6436 a_n9628_8799.t79 gnd 0.601374f
C6437 a_n9628_8799.n279 gnd 0.052275f
C6438 a_n9628_8799.t49 gnd 0.601374f
C6439 a_n9628_8799.n280 gnd 0.268585f
C6440 a_n9628_8799.n281 gnd 0.052275f
C6441 a_n9628_8799.t124 gnd 0.601374f
C6442 a_n9628_8799.t80 gnd 0.601374f
C6443 a_n9628_8799.n282 gnd 0.052275f
C6444 a_n9628_8799.t41 gnd 0.601374f
C6445 a_n9628_8799.n283 gnd 0.268585f
C6446 a_n9628_8799.n284 gnd 0.052275f
C6447 a_n9628_8799.t129 gnd 0.601374f
C6448 a_n9628_8799.t95 gnd 0.601374f
C6449 a_n9628_8799.n285 gnd 0.052275f
C6450 a_n9628_8799.t59 gnd 0.601374f
C6451 a_n9628_8799.n286 gnd 0.268585f
C6452 a_n9628_8799.n287 gnd 0.052275f
C6453 a_n9628_8799.t149 gnd 0.601374f
C6454 a_n9628_8799.t130 gnd 0.601374f
C6455 a_n9628_8799.n288 gnd 0.052275f
C6456 a_n9628_8799.t66 gnd 0.601374f
C6457 a_n9628_8799.n289 gnd 0.268585f
C6458 a_n9628_8799.t152 gnd 0.612756f
C6459 a_n9628_8799.n290 gnd 0.2521f
C6460 a_n9628_8799.t153 gnd 0.601374f
C6461 a_n9628_8799.n291 gnd 0.264879f
C6462 a_n9628_8799.n292 gnd 0.011862f
C6463 a_n9628_8799.n293 gnd 0.16515f
C6464 a_n9628_8799.n294 gnd 0.052275f
C6465 a_n9628_8799.n295 gnd 0.052275f
C6466 a_n9628_8799.n296 gnd 0.011862f
C6467 a_n9628_8799.n297 gnd 0.26649f
C6468 a_n9628_8799.n298 gnd 0.265201f
C6469 a_n9628_8799.n299 gnd 0.011862f
C6470 a_n9628_8799.n300 gnd 0.052275f
C6471 a_n9628_8799.n301 gnd 0.052275f
C6472 a_n9628_8799.n302 gnd 0.052275f
C6473 a_n9628_8799.n303 gnd 0.011862f
C6474 a_n9628_8799.n304 gnd 0.266168f
C6475 a_n9628_8799.n305 gnd 0.265523f
C6476 a_n9628_8799.n306 gnd 0.011862f
C6477 a_n9628_8799.n307 gnd 0.052275f
C6478 a_n9628_8799.n308 gnd 0.052275f
C6479 a_n9628_8799.n309 gnd 0.052275f
C6480 a_n9628_8799.n310 gnd 0.011862f
C6481 a_n9628_8799.n311 gnd 0.265846f
C6482 a_n9628_8799.n312 gnd 0.265846f
C6483 a_n9628_8799.n313 gnd 0.011862f
C6484 a_n9628_8799.n314 gnd 0.052275f
C6485 a_n9628_8799.n315 gnd 0.052275f
C6486 a_n9628_8799.n316 gnd 0.052275f
C6487 a_n9628_8799.n317 gnd 0.011862f
C6488 a_n9628_8799.n318 gnd 0.265523f
C6489 a_n9628_8799.n319 gnd 0.266168f
C6490 a_n9628_8799.n320 gnd 0.011862f
C6491 a_n9628_8799.n321 gnd 0.052275f
C6492 a_n9628_8799.n322 gnd 0.052275f
C6493 a_n9628_8799.n323 gnd 0.052275f
C6494 a_n9628_8799.n324 gnd 0.011862f
C6495 a_n9628_8799.n325 gnd 0.265201f
C6496 a_n9628_8799.n326 gnd 0.26649f
C6497 a_n9628_8799.n327 gnd 0.011862f
C6498 a_n9628_8799.n328 gnd 0.052275f
C6499 a_n9628_8799.n329 gnd 0.052275f
C6500 a_n9628_8799.n330 gnd 0.052275f
C6501 a_n9628_8799.n331 gnd 0.011862f
C6502 a_n9628_8799.n332 gnd 0.264879f
C6503 a_n9628_8799.n333 gnd 0.263106f
C6504 a_n9628_8799.n334 gnd 0.130296f
C6505 a_n9628_8799.n335 gnd 0.904082f
C6506 a_n9628_8799.n336 gnd 0.052275f
C6507 a_n9628_8799.t106 gnd 0.601374f
C6508 a_n9628_8799.t128 gnd 0.601374f
C6509 a_n9628_8799.t64 gnd 0.601374f
C6510 a_n9628_8799.n337 gnd 0.268585f
C6511 a_n9628_8799.n338 gnd 0.052275f
C6512 a_n9628_8799.t146 gnd 0.601374f
C6513 a_n9628_8799.t83 gnd 0.601374f
C6514 a_n9628_8799.n339 gnd 0.052275f
C6515 a_n9628_8799.t139 gnd 0.601374f
C6516 a_n9628_8799.n340 gnd 0.268585f
C6517 a_n9628_8799.n341 gnd 0.052275f
C6518 a_n9628_8799.t70 gnd 0.601374f
C6519 a_n9628_8799.t118 gnd 0.601374f
C6520 a_n9628_8799.n342 gnd 0.052275f
C6521 a_n9628_8799.t55 gnd 0.601374f
C6522 a_n9628_8799.n343 gnd 0.268585f
C6523 a_n9628_8799.n344 gnd 0.052275f
C6524 a_n9628_8799.t101 gnd 0.601374f
C6525 a_n9628_8799.t78 gnd 0.601374f
C6526 a_n9628_8799.n345 gnd 0.052275f
C6527 a_n9628_8799.t126 gnd 0.601374f
C6528 a_n9628_8799.n346 gnd 0.268585f
C6529 a_n9628_8799.n347 gnd 0.052275f
C6530 a_n9628_8799.t62 gnd 0.601374f
C6531 a_n9628_8799.t110 gnd 0.601374f
C6532 a_n9628_8799.n348 gnd 0.052275f
C6533 a_n9628_8799.t44 gnd 0.601374f
C6534 a_n9628_8799.n349 gnd 0.268585f
C6535 a_n9628_8799.n350 gnd 0.052275f
C6536 a_n9628_8799.t94 gnd 0.601374f
C6537 a_n9628_8799.t158 gnd 0.601374f
C6538 a_n9628_8799.n351 gnd 0.052275f
C6539 a_n9628_8799.t117 gnd 0.601374f
C6540 a_n9628_8799.n352 gnd 0.268585f
C6541 a_n9628_8799.t75 gnd 0.612756f
C6542 a_n9628_8799.n353 gnd 0.2521f
C6543 a_n9628_8799.t54 gnd 0.601374f
C6544 a_n9628_8799.n354 gnd 0.264879f
C6545 a_n9628_8799.n355 gnd 0.011862f
C6546 a_n9628_8799.n356 gnd 0.16515f
C6547 a_n9628_8799.n357 gnd 0.052275f
C6548 a_n9628_8799.n358 gnd 0.052275f
C6549 a_n9628_8799.n359 gnd 0.011862f
C6550 a_n9628_8799.n360 gnd 0.26649f
C6551 a_n9628_8799.n361 gnd 0.265201f
C6552 a_n9628_8799.n362 gnd 0.011862f
C6553 a_n9628_8799.n363 gnd 0.052275f
C6554 a_n9628_8799.n364 gnd 0.052275f
C6555 a_n9628_8799.n365 gnd 0.052275f
C6556 a_n9628_8799.n366 gnd 0.011862f
C6557 a_n9628_8799.n367 gnd 0.266168f
C6558 a_n9628_8799.n368 gnd 0.265523f
C6559 a_n9628_8799.n369 gnd 0.011862f
C6560 a_n9628_8799.n370 gnd 0.052275f
C6561 a_n9628_8799.n371 gnd 0.052275f
C6562 a_n9628_8799.n372 gnd 0.052275f
C6563 a_n9628_8799.n373 gnd 0.011862f
C6564 a_n9628_8799.n374 gnd 0.265846f
C6565 a_n9628_8799.n375 gnd 0.265846f
C6566 a_n9628_8799.n376 gnd 0.011862f
C6567 a_n9628_8799.n377 gnd 0.052275f
C6568 a_n9628_8799.n378 gnd 0.052275f
C6569 a_n9628_8799.n379 gnd 0.052275f
C6570 a_n9628_8799.n380 gnd 0.011862f
C6571 a_n9628_8799.n381 gnd 0.265523f
C6572 a_n9628_8799.n382 gnd 0.266168f
C6573 a_n9628_8799.n383 gnd 0.011862f
C6574 a_n9628_8799.n384 gnd 0.052275f
C6575 a_n9628_8799.n385 gnd 0.052275f
C6576 a_n9628_8799.n386 gnd 0.052275f
C6577 a_n9628_8799.n387 gnd 0.011862f
C6578 a_n9628_8799.n388 gnd 0.265201f
C6579 a_n9628_8799.n389 gnd 0.26649f
C6580 a_n9628_8799.n390 gnd 0.011862f
C6581 a_n9628_8799.n391 gnd 0.052275f
C6582 a_n9628_8799.n392 gnd 0.052275f
C6583 a_n9628_8799.n393 gnd 0.052275f
C6584 a_n9628_8799.n394 gnd 0.011862f
C6585 a_n9628_8799.n395 gnd 0.264879f
C6586 a_n9628_8799.n396 gnd 0.263106f
C6587 a_n9628_8799.n397 gnd 0.130296f
C6588 a_n9628_8799.n398 gnd 1.45409f
C6589 a_n9628_8799.n399 gnd 17.4871f
C6590 a_n9628_8799.n400 gnd 4.40119f
C6591 a_n9628_8799.t24 gnd 0.112803f
C6592 a_n9628_8799.t25 gnd 0.112803f
C6593 a_n9628_8799.n401 gnd 0.998987f
C6594 a_n9628_8799.t20 gnd 0.112803f
C6595 a_n9628_8799.t21 gnd 0.112803f
C6596 a_n9628_8799.n402 gnd 0.996771f
C6597 a_n9628_8799.n403 gnd 0.735628f
C6598 a_n9628_8799.n404 gnd 0.473327f
C6599 a_n9628_8799.t19 gnd 0.112803f
C6600 a_n9628_8799.t31 gnd 0.112803f
C6601 a_n9628_8799.n405 gnd 0.996771f
C6602 a_n9628_8799.n406 gnd 0.331536f
C6603 a_n9628_8799.t32 gnd 0.112803f
C6604 a_n9628_8799.t28 gnd 0.112803f
C6605 a_n9628_8799.n407 gnd 0.996771f
C6606 a_n9628_8799.n408 gnd 2.58476f
C6607 a_n9628_8799.t29 gnd 0.112803f
C6608 a_n9628_8799.t27 gnd 0.112803f
C6609 a_n9628_8799.n409 gnd 0.998987f
C6610 a_n9628_8799.t22 gnd 0.112803f
C6611 a_n9628_8799.t26 gnd 0.112803f
C6612 a_n9628_8799.n410 gnd 0.99677f
C6613 a_n9628_8799.n411 gnd 0.73563f
C6614 a_n9628_8799.n412 gnd 2.00128f
C6615 a_n9628_8799.t33 gnd 0.112803f
C6616 a_n9628_8799.t23 gnd 0.112803f
C6617 a_n9628_8799.n413 gnd 0.99677f
C6618 a_n9628_8799.n414 gnd 0.735633f
C6619 a_n9628_8799.n415 gnd 0.998984f
C6620 a_n9628_8799.t34 gnd 0.112803f
C6621 a_n3827_n3924.n0 gnd 1.73844f
C6622 a_n3827_n3924.n1 gnd 1.46101f
C6623 a_n3827_n3924.n2 gnd 1.14592f
C6624 a_n3827_n3924.n3 gnd 1.10826f
C6625 a_n3827_n3924.n4 gnd 1.26277f
C6626 a_n3827_n3924.n5 gnd 1.54321f
C6627 a_n3827_n3924.n6 gnd 2.44001f
C6628 a_n3827_n3924.n7 gnd 2.62589f
C6629 a_n3827_n3924.n8 gnd 1.27065f
C6630 a_n3827_n3924.n9 gnd 0.94769f
C6631 a_n3827_n3924.t18 gnd 0.084838f
C6632 a_n3827_n3924.t17 gnd 0.084838f
C6633 a_n3827_n3924.t10 gnd 0.084838f
C6634 a_n3827_n3924.n10 gnd 0.692885f
C6635 a_n3827_n3924.t9 gnd 1.09854f
C6636 a_n3827_n3924.t5 gnd 1.09554f
C6637 a_n3827_n3924.t14 gnd 0.881736f
C6638 a_n3827_n3924.t41 gnd 1.0971f
C6639 a_n3827_n3924.t22 gnd 1.09554f
C6640 a_n3827_n3924.t19 gnd 1.09554f
C6641 a_n3827_n3924.t40 gnd 1.09554f
C6642 a_n3827_n3924.t23 gnd 1.09554f
C6643 a_n3827_n3924.t1 gnd 1.09554f
C6644 a_n3827_n3924.t13 gnd 1.09554f
C6645 a_n3827_n3924.t7 gnd 1.09554f
C6646 a_n3827_n3924.n11 gnd 0.795808f
C6647 a_n3827_n3924.t33 gnd 0.881733f
C6648 a_n3827_n3924.t38 gnd 0.084838f
C6649 a_n3827_n3924.t36 gnd 0.084838f
C6650 a_n3827_n3924.n12 gnd 0.692884f
C6651 a_n3827_n3924.t25 gnd 0.084838f
C6652 a_n3827_n3924.t35 gnd 0.084838f
C6653 a_n3827_n3924.n13 gnd 0.692884f
C6654 a_n3827_n3924.t28 gnd 0.084838f
C6655 a_n3827_n3924.t29 gnd 0.084838f
C6656 a_n3827_n3924.n14 gnd 0.692884f
C6657 a_n3827_n3924.t26 gnd 0.881733f
C6658 a_n3827_n3924.t12 gnd 0.881733f
C6659 a_n3827_n3924.t4 gnd 0.084838f
C6660 a_n3827_n3924.t3 gnd 0.084838f
C6661 a_n3827_n3924.n15 gnd 0.692884f
C6662 a_n3827_n3924.t2 gnd 0.084838f
C6663 a_n3827_n3924.t20 gnd 0.084838f
C6664 a_n3827_n3924.n16 gnd 0.692884f
C6665 a_n3827_n3924.t8 gnd 0.084838f
C6666 a_n3827_n3924.t16 gnd 0.084838f
C6667 a_n3827_n3924.n17 gnd 0.692884f
C6668 a_n3827_n3924.t15 gnd 0.881733f
C6669 a_n3827_n3924.n18 gnd 0.795808f
C6670 a_n3827_n3924.t27 gnd 0.881733f
C6671 a_n3827_n3924.t34 gnd 0.084838f
C6672 a_n3827_n3924.t30 gnd 0.084838f
C6673 a_n3827_n3924.n19 gnd 0.692885f
C6674 a_n3827_n3924.t24 gnd 0.084838f
C6675 a_n3827_n3924.t32 gnd 0.084838f
C6676 a_n3827_n3924.n20 gnd 0.692885f
C6677 a_n3827_n3924.t39 gnd 0.084838f
C6678 a_n3827_n3924.t31 gnd 0.084838f
C6679 a_n3827_n3924.n21 gnd 0.692885f
C6680 a_n3827_n3924.t37 gnd 0.881736f
C6681 a_n3827_n3924.t11 gnd 0.881736f
C6682 a_n3827_n3924.t21 gnd 0.084838f
C6683 a_n3827_n3924.t6 gnd 0.084838f
C6684 a_n3827_n3924.n22 gnd 0.692885f
C6685 a_n3827_n3924.n23 gnd 0.692886f
C6686 a_n3827_n3924.t0 gnd 0.084838f
C6687 plus.n0 gnd 0.02154f
C6688 plus.t9 gnd 0.304662f
C6689 plus.n1 gnd 0.02154f
C6690 plus.t5 gnd 0.304662f
C6691 plus.t6 gnd 0.304662f
C6692 plus.n2 gnd 0.135341f
C6693 plus.n3 gnd 0.02154f
C6694 plus.t16 gnd 0.304662f
C6695 plus.t17 gnd 0.304662f
C6696 plus.n4 gnd 0.135341f
C6697 plus.n5 gnd 0.02154f
C6698 plus.t13 gnd 0.304662f
C6699 plus.t10 gnd 0.304662f
C6700 plus.n6 gnd 0.138291f
C6701 plus.t12 gnd 0.31493f
C6702 plus.n7 gnd 0.126865f
C6703 plus.n8 gnd 0.091152f
C6704 plus.n9 gnd 0.004888f
C6705 plus.n10 gnd 0.135341f
C6706 plus.n11 gnd 0.004888f
C6707 plus.n12 gnd 0.02154f
C6708 plus.n13 gnd 0.02154f
C6709 plus.n14 gnd 0.02154f
C6710 plus.n15 gnd 0.004888f
C6711 plus.n16 gnd 0.135341f
C6712 plus.n17 gnd 0.004888f
C6713 plus.n18 gnd 0.02154f
C6714 plus.n19 gnd 0.02154f
C6715 plus.n20 gnd 0.02154f
C6716 plus.n21 gnd 0.004888f
C6717 plus.n22 gnd 0.135341f
C6718 plus.n23 gnd 0.004888f
C6719 plus.n24 gnd 0.134743f
C6720 plus.n25 gnd 0.24275f
C6721 plus.n26 gnd 0.02154f
C6722 plus.n27 gnd 0.004888f
C6723 plus.t7 gnd 0.304662f
C6724 plus.n28 gnd 0.02154f
C6725 plus.n29 gnd 0.004888f
C6726 plus.t20 gnd 0.304662f
C6727 plus.n30 gnd 0.02154f
C6728 plus.n31 gnd 0.004888f
C6729 plus.t19 gnd 0.304662f
C6730 plus.t15 gnd 0.31493f
C6731 plus.t14 gnd 0.304662f
C6732 plus.n32 gnd 0.138291f
C6733 plus.n33 gnd 0.126865f
C6734 plus.n34 gnd 0.091152f
C6735 plus.n35 gnd 0.02154f
C6736 plus.n36 gnd 0.135341f
C6737 plus.n37 gnd 0.004888f
C6738 plus.t18 gnd 0.304662f
C6739 plus.n38 gnd 0.135341f
C6740 plus.n39 gnd 0.02154f
C6741 plus.n40 gnd 0.02154f
C6742 plus.n41 gnd 0.02154f
C6743 plus.n42 gnd 0.135341f
C6744 plus.n43 gnd 0.004888f
C6745 plus.t8 gnd 0.304662f
C6746 plus.n44 gnd 0.135341f
C6747 plus.n45 gnd 0.02154f
C6748 plus.n46 gnd 0.02154f
C6749 plus.n47 gnd 0.02154f
C6750 plus.n48 gnd 0.135341f
C6751 plus.n49 gnd 0.004888f
C6752 plus.t11 gnd 0.304662f
C6753 plus.n50 gnd 0.134743f
C6754 plus.n51 gnd 0.616554f
C6755 plus.n52 gnd 0.942186f
C6756 plus.t2 gnd 0.037184f
C6757 plus.t1 gnd 0.00664f
C6758 plus.t0 gnd 0.00664f
C6759 plus.n53 gnd 0.021535f
C6760 plus.n54 gnd 0.167179f
C6761 plus.t3 gnd 0.00664f
C6762 plus.t4 gnd 0.00664f
C6763 plus.n55 gnd 0.021535f
C6764 plus.n56 gnd 0.125488f
C6765 plus.n57 gnd 2.76704f
.ends

