* NGSPICE file created from opamp.ext - technology: sky130A

.subckt opamp output vdd plus minus commonsourceibias outputibias diffpairibias gnd CSoutput
Cload output gnd 0.0p
X0 gnd.t322 gnd.t319 gnd.t321 gnd.t320 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X1 gnd.t194 commonsourceibias.t46 commonsourceibias.t47 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X2 vdd.t180 a_n5644_8799.t36 CSoutput.t72 vdd.t127 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X3 a_n1986_8322.t11 a_n1986_13878.t48 vdd.t26 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 a_n1808_13878.t11 a_n1986_13878.t31 a_n1986_13878.t32 vdd.t30 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X5 commonsourceibias.t45 commonsourceibias.t44 gnd.t328 gnd.t106 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X6 a_n3827_n3924.t20 diffpairibias.t20 gnd.t83 gnd.t82 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X7 a_n1986_13878.t30 a_n1986_13878.t29 a_n1808_13878.t10 vdd.t35 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X8 a_n1808_13878.t9 a_n1986_13878.t15 a_n1986_13878.t16 vdd.t197 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X9 vdd.t116 vdd.t114 vdd.t115 vdd.t89 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X10 a_n1808_13878.t19 a_n1986_13878.t49 vdd.t28 vdd.t27 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X11 CSoutput.t108 a_n5644_8799.t37 vdd.t179 vdd.t123 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X12 gnd.t143 commonsourceibias.t42 commonsourceibias.t43 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X13 gnd.t318 gnd.t316 gnd.t317 gnd.t239 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X14 gnd.t118 commonsourceibias.t48 CSoutput.t71 gnd.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X15 commonsourceibias.t41 commonsourceibias.t40 gnd.t169 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X16 vdd.t113 vdd.t111 vdd.t112 vdd.t64 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X17 minus.t4 gnd.t313 gnd.t315 gnd.t314 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X18 gnd.t312 gnd.t311 plus.t4 gnd.t239 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X19 a_n5644_8799.t26 plus.t5 a_n3827_n3924.t44 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X20 gnd.t310 gnd.t308 gnd.t309 gnd.t235 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X21 output.t19 outputibias.t8 gnd.t138 gnd.t137 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X22 gnd.t307 gnd.t305 gnd.t306 gnd.t231 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X23 a_n1986_8322.t23 a_n1986_13878.t50 a_n5644_8799.t11 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X24 commonsourceibias.t39 commonsourceibias.t38 gnd.t333 gnd.t87 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X25 gnd.t81 commonsourceibias.t49 CSoutput.t70 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X26 CSoutput.t69 commonsourceibias.t50 gnd.t332 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X27 a_n5644_8799.t24 plus.t6 a_n3827_n3924.t42 gnd.t76 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X28 gnd.t304 gnd.t301 gnd.t303 gnd.t302 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X29 CSoutput.t107 a_n5644_8799.t38 vdd.t178 vdd.t136 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X30 vdd.t177 a_n5644_8799.t39 CSoutput.t106 vdd.t154 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X31 gnd.t141 commonsourceibias.t36 commonsourceibias.t37 gnd.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 a_n5644_8799.t12 a_n1986_13878.t51 a_n1986_8322.t22 vdd.t30 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X33 CSoutput.t77 a_n5644_8799.t40 vdd.t176 vdd.t117 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X34 vdd.t175 a_n5644_8799.t41 CSoutput.t76 vdd.t170 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X35 a_n3827_n3924.t37 minus.t5 a_n1986_13878.t40 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X36 a_n3827_n3924.t19 diffpairibias.t21 gnd.t109 gnd.t108 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X37 commonsourceibias.t35 commonsourceibias.t34 gnd.t128 gnd.t99 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X38 a_n1986_13878.t0 minus.t6 a_n3827_n3924.t7 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X39 a_n3827_n3924.t3 plus.t7 a_n5644_8799.t3 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X40 a_n3827_n3924.t0 plus.t8 a_n5644_8799.t0 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X41 a_n3827_n3924.t54 minus.t7 a_n1986_13878.t47 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X42 CSoutput.t75 a_n5644_8799.t42 vdd.t174 vdd.t132 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X43 vdd.t110 vdd.t108 vdd.t109 vdd.t42 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X44 CSoutput.t68 commonsourceibias.t51 gnd.t29 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X45 gnd.t8 commonsourceibias.t32 commonsourceibias.t33 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X46 output.t15 CSoutput.t120 vdd.t5 gnd.t105 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X47 output.t18 outputibias.t9 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X48 a_n3827_n3924.t10 minus.t8 a_n1986_13878.t2 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X49 a_n1808_13878.t8 a_n1986_13878.t35 a_n1986_13878.t36 vdd.t40 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X50 vdd.t173 a_n5644_8799.t43 CSoutput.t85 vdd.t170 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X51 diffpairibias.t19 diffpairibias.t18 gnd.t196 gnd.t195 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X52 a_n1986_13878.t34 a_n1986_13878.t33 a_n1808_13878.t7 vdd.t34 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X53 CSoutput.t84 a_n5644_8799.t44 vdd.t172 vdd.t148 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X54 vdd.t107 vdd.t105 vdd.t106 vdd.t74 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X55 gnd.t300 gnd.t298 plus.t3 gnd.t299 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X56 CSoutput.t67 commonsourceibias.t52 gnd.t101 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X57 gnd.t297 gnd.t295 gnd.t296 gnd.t215 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X58 a_n1986_13878.t41 minus.t9 a_n3827_n3924.t38 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X59 CSoutput.t66 commonsourceibias.t53 gnd.t134 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X60 diffpairibias.t17 diffpairibias.t16 gnd.t123 gnd.t122 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X61 gnd.t294 gnd.t292 gnd.t293 gnd.t215 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X62 vdd.t104 vdd.t102 vdd.t103 vdd.t53 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X63 CSoutput.t121 a_n1986_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X64 vdd.t171 a_n5644_8799.t45 CSoutput.t83 vdd.t170 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X65 CSoutput.t65 commonsourceibias.t54 gnd.t198 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X66 vdd.t169 a_n5644_8799.t46 CSoutput.t93 vdd.t145 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X67 CSoutput.t92 a_n5644_8799.t47 vdd.t168 vdd.t117 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X68 plus.t2 gnd.t289 gnd.t291 gnd.t290 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X69 gnd.t41 commonsourceibias.t55 CSoutput.t64 gnd.t40 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X70 vdd.t167 a_n5644_8799.t48 CSoutput.t113 vdd.t121 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X71 gnd.t116 commonsourceibias.t56 CSoutput.t63 gnd.t50 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X72 a_n5644_8799.t29 plus.t9 a_n3827_n3924.t47 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X73 CSoutput.t62 commonsourceibias.t57 gnd.t132 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X74 CSoutput.t122 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X75 gnd.t288 gnd.t286 gnd.t287 gnd.t231 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X76 CSoutput.t112 a_n5644_8799.t49 vdd.t166 vdd.t132 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X77 CSoutput.t111 a_n5644_8799.t50 vdd.t165 vdd.t158 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X78 output.t14 CSoutput.t123 vdd.t14 gnd.t176 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X79 a_n3827_n3924.t18 diffpairibias.t22 gnd.t203 gnd.t202 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X80 CSoutput.t116 a_n5644_8799.t51 vdd.t164 vdd.t158 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X81 a_n3827_n3924.t51 minus.t10 a_n1986_13878.t44 gnd.t327 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X82 CSoutput.t61 commonsourceibias.t58 gnd.t49 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X83 vdd.t163 a_n5644_8799.t52 CSoutput.t115 vdd.t156 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X84 a_n3827_n3924.t39 plus.t10 a_n5644_8799.t21 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X85 a_n1986_13878.t10 minus.t11 a_n3827_n3924.t29 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X86 outputibias.t7 outputibias.t6 gnd.t39 gnd.t38 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X87 a_n1986_13878.t26 a_n1986_13878.t25 a_n1808_13878.t6 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X88 CSoutput.t60 commonsourceibias.t59 gnd.t323 gnd.t106 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 gnd.t72 commonsourceibias.t60 CSoutput.t59 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 commonsourceibias.t31 commonsourceibias.t30 gnd.t136 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 a_n1986_13878.t14 a_n1986_13878.t13 a_n1808_13878.t5 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X92 vdd.t162 a_n5644_8799.t53 CSoutput.t114 vdd.t154 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X93 a_n5644_8799.t20 a_n1986_13878.t52 a_n1986_8322.t21 vdd.t187 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X94 gnd.t285 gnd.t283 gnd.t284 gnd.t227 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X95 vdd.t161 a_n5644_8799.t54 CSoutput.t80 vdd.t156 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X96 a_n3827_n3924.t36 minus.t12 a_n1986_13878.t39 gnd.t153 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X97 diffpairibias.t15 diffpairibias.t14 gnd.t60 gnd.t59 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X98 outputibias.t5 outputibias.t4 gnd.t140 gnd.t139 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X99 vdd.t101 vdd.t99 vdd.t100 vdd.t53 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X100 vdd.t160 a_n5644_8799.t55 CSoutput.t79 vdd.t145 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X101 vdd.t98 vdd.t96 vdd.t97 vdd.t82 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X102 CSoutput.t58 commonsourceibias.t61 gnd.t88 gnd.t87 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X103 gnd.t199 commonsourceibias.t28 commonsourceibias.t29 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X104 vdd.t95 vdd.t92 vdd.t94 vdd.t93 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X105 a_n1986_13878.t46 minus.t13 a_n3827_n3924.t53 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X106 gnd.t170 commonsourceibias.t62 CSoutput.t57 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X107 output.t13 CSoutput.t124 vdd.t8 gnd.t177 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X108 a_n3827_n3924.t17 diffpairibias.t23 gnd.t62 gnd.t61 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X109 vdd.t91 vdd.t88 vdd.t90 vdd.t89 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X110 vdd.t10 CSoutput.t125 output.t12 gnd.t178 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X111 vdd.t189 a_n1986_13878.t53 a_n1986_8322.t10 vdd.t188 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X112 vdd.t87 vdd.t85 vdd.t86 vdd.t78 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X113 gnd.t282 gnd.t280 minus.t3 gnd.t281 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X114 a_n3827_n3924.t43 plus.t11 a_n5644_8799.t25 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X115 commonsourceibias.t27 commonsourceibias.t26 gnd.t334 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X116 gnd.t174 commonsourceibias.t63 CSoutput.t56 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X117 CSoutput.t78 a_n5644_8799.t56 vdd.t159 vdd.t158 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X118 a_n1986_8322.t9 a_n1986_13878.t54 vdd.t17 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X119 gnd.t279 gnd.t277 gnd.t278 gnd.t205 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X120 gnd.t24 commonsourceibias.t24 commonsourceibias.t25 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X121 gnd.t276 gnd.t274 gnd.t275 gnd.t227 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X122 vdd.t157 a_n5644_8799.t57 CSoutput.t87 vdd.t156 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X123 vdd.t1 CSoutput.t126 output.t11 gnd.t179 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X124 vdd.t19 a_n1986_13878.t55 a_n1808_13878.t18 vdd.t18 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X125 CSoutput.t55 commonsourceibias.t64 gnd.t190 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X126 a_n1986_13878.t9 minus.t14 a_n3827_n3924.t28 gnd.t97 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X127 a_n5644_8799.t23 plus.t12 a_n3827_n3924.t41 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X128 gnd.t160 commonsourceibias.t65 CSoutput.t54 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X129 commonsourceibias.t23 commonsourceibias.t22 gnd.t154 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X130 vdd.t84 vdd.t81 vdd.t83 vdd.t82 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X131 diffpairibias.t13 diffpairibias.t12 gnd.t130 gnd.t129 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X132 vdd.t80 vdd.t77 vdd.t79 vdd.t78 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X133 vdd.t155 a_n5644_8799.t58 CSoutput.t86 vdd.t154 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X134 a_n5644_8799.t7 a_n1986_13878.t56 a_n1986_8322.t20 vdd.t20 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X135 a_n1986_8322.t8 a_n1986_13878.t57 vdd.t22 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X136 vdd.t76 vdd.t73 vdd.t75 vdd.t74 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X137 a_n1986_13878.t18 a_n1986_13878.t17 a_n1808_13878.t4 vdd.t196 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X138 gnd.t90 commonsourceibias.t66 CSoutput.t53 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X139 a_n3827_n3924.t31 minus.t15 a_n1986_13878.t12 gnd.t120 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X140 a_n3827_n3924.t50 minus.t16 a_n1986_13878.t43 gnd.t175 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X141 a_n5644_8799.t22 plus.t13 a_n3827_n3924.t40 gnd.t95 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X142 gnd.t34 commonsourceibias.t67 CSoutput.t52 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X143 a_n5644_8799.t32 a_n1986_13878.t58 a_n1986_8322.t19 vdd.t197 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X144 a_n1986_13878.t1 minus.t17 a_n3827_n3924.t8 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X145 vdd.t11 CSoutput.t127 output.t10 gnd.t180 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X146 a_n1808_13878.t3 a_n1986_13878.t27 a_n1986_13878.t28 vdd.t187 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X147 output.t9 CSoutput.t128 vdd.t4 gnd.t181 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X148 gnd.t273 gnd.t271 gnd.t272 gnd.t231 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X149 CSoutput.t51 commonsourceibias.t68 gnd.t166 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X150 vdd.t199 a_n1986_13878.t59 a_n1986_8322.t7 vdd.t198 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X151 gnd.t167 commonsourceibias.t69 CSoutput.t50 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X152 output.t8 CSoutput.t129 vdd.t13 gnd.t182 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X153 gnd.t184 commonsourceibias.t70 CSoutput.t49 gnd.t40 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X154 vdd.t72 vdd.t70 vdd.t71 vdd.t64 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X155 a_n3827_n3924.t16 diffpairibias.t24 gnd.t15 gnd.t14 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X156 CSoutput.t103 a_n5644_8799.t59 vdd.t153 vdd.t148 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X157 a_n1986_13878.t6 minus.t18 a_n3827_n3924.t25 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X158 a_n3827_n3924.t15 diffpairibias.t25 gnd.t12 gnd.t11 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X159 vdd.t152 a_n5644_8799.t60 CSoutput.t102 vdd.t119 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X160 gnd.t270 gnd.t268 gnd.t269 gnd.t205 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X161 gnd.t267 gnd.t265 minus.t2 gnd.t266 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X162 vdd.t151 a_n5644_8799.t61 CSoutput.t101 vdd.t134 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X163 a_n1986_13878.t4 minus.t19 a_n3827_n3924.t22 gnd.t76 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X164 CSoutput.t48 commonsourceibias.t71 gnd.t43 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 gnd.t264 gnd.t261 gnd.t263 gnd.t262 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X166 gnd.t260 gnd.t258 gnd.t259 gnd.t215 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X167 gnd.t86 commonsourceibias.t72 CSoutput.t47 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X168 diffpairibias.t11 diffpairibias.t10 gnd.t193 gnd.t192 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X169 vdd.t6 CSoutput.t130 output.t7 gnd.t183 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X170 a_n3827_n3924.t4 plus.t14 a_n5644_8799.t4 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X171 gnd.t165 commonsourceibias.t73 CSoutput.t46 gnd.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X172 CSoutput.t45 commonsourceibias.t74 gnd.t110 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X173 CSoutput.t100 a_n5644_8799.t62 vdd.t150 vdd.t138 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X174 vdd.t69 vdd.t67 vdd.t68 vdd.t49 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X175 a_n1808_13878.t17 a_n1986_13878.t60 vdd.t191 vdd.t190 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X176 vdd.t193 a_n1986_13878.t61 a_n1808_13878.t16 vdd.t192 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X177 gnd.t54 commonsourceibias.t75 CSoutput.t44 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X178 a_n3827_n3924.t35 minus.t20 a_n1986_13878.t38 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X179 a_n3827_n3924.t23 plus.t15 a_n5644_8799.t14 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X180 diffpairibias.t9 diffpairibias.t8 gnd.t201 gnd.t200 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X181 a_n5644_8799.t35 plus.t16 a_n3827_n3924.t57 gnd.t147 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X182 a_n3827_n3924.t52 minus.t21 a_n1986_13878.t45 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X183 CSoutput.t131 a_n1986_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X184 vdd.t66 vdd.t63 vdd.t65 vdd.t64 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X185 gnd.t257 gnd.t255 gnd.t256 gnd.t205 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X186 commonsourceibias.t21 commonsourceibias.t20 gnd.t163 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X187 diffpairibias.t7 diffpairibias.t6 gnd.t115 gnd.t114 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X188 CSoutput.t99 a_n5644_8799.t63 vdd.t149 vdd.t148 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X189 vdd.t147 a_n5644_8799.t64 CSoutput.t98 vdd.t119 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X190 CSoutput.t132 a_n1986_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X191 output.t17 outputibias.t10 gnd.t93 gnd.t92 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X192 CSoutput.t43 commonsourceibias.t76 gnd.t329 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X193 a_n1986_8322.t18 a_n1986_13878.t62 a_n5644_8799.t15 vdd.t35 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X194 gnd.t254 gnd.t252 gnd.t253 gnd.t227 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X195 commonsourceibias.t19 commonsourceibias.t18 gnd.t78 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 vdd.t146 a_n5644_8799.t65 CSoutput.t97 vdd.t145 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X197 CSoutput.t95 a_n5644_8799.t66 vdd.t144 vdd.t125 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X198 gnd.t251 gnd.t248 gnd.t250 gnd.t249 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X199 vdd.t143 a_n5644_8799.t67 CSoutput.t94 vdd.t134 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X200 vdd.t37 a_n1986_13878.t63 a_n1986_8322.t6 vdd.t36 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X201 plus.t1 gnd.t245 gnd.t247 gnd.t246 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X202 CSoutput.t42 commonsourceibias.t77 gnd.t98 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X203 output.t16 outputibias.t11 gnd.t158 gnd.t157 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X204 gnd.t71 commonsourceibias.t78 CSoutput.t41 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X205 gnd.t244 gnd.t242 minus.t1 gnd.t243 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X206 CSoutput.t40 commonsourceibias.t79 gnd.t148 gnd.t106 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 gnd.t241 gnd.t238 gnd.t240 gnd.t239 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X208 output.t6 CSoutput.t133 vdd.t3 gnd.t63 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X209 gnd.t162 commonsourceibias.t16 commonsourceibias.t17 gnd.t50 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X210 gnd.t113 commonsourceibias.t80 CSoutput.t39 gnd.t40 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X211 a_n1808_13878.t15 a_n1986_13878.t64 vdd.t195 vdd.t194 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X212 gnd.t237 gnd.t234 gnd.t236 gnd.t235 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X213 gnd.t233 gnd.t230 gnd.t232 gnd.t231 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X214 CSoutput.t38 commonsourceibias.t81 gnd.t331 gnd.t87 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X215 gnd.t325 commonsourceibias.t82 CSoutput.t37 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X216 CSoutput.t36 commonsourceibias.t83 gnd.t104 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X217 commonsourceibias.t15 commonsourceibias.t14 gnd.t161 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X218 a_n3827_n3924.t14 diffpairibias.t26 gnd.t172 gnd.t171 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X219 CSoutput.t119 a_n5644_8799.t68 vdd.t142 vdd.t138 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X220 CSoutput.t35 commonsourceibias.t84 gnd.t68 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X221 gnd.t89 commonsourceibias.t85 CSoutput.t34 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X222 CSoutput.t118 a_n5644_8799.t69 vdd.t141 vdd.t136 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X223 vdd.t62 vdd.t60 vdd.t61 vdd.t49 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X224 gnd.t74 commonsourceibias.t86 CSoutput.t33 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X225 CSoutput.t32 commonsourceibias.t87 gnd.t168 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X226 a_n1986_8322.t17 a_n1986_13878.t65 a_n5644_8799.t30 vdd.t196 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X227 vdd.t186 a_n1986_13878.t66 a_n1986_8322.t5 vdd.t185 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X228 vdd.t140 a_n5644_8799.t70 CSoutput.t117 vdd.t127 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X229 CSoutput.t105 a_n5644_8799.t71 vdd.t139 vdd.t138 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X230 CSoutput.t31 commonsourceibias.t88 gnd.t56 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X231 gnd.t51 commonsourceibias.t89 CSoutput.t30 gnd.t50 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X232 a_n3827_n3924.t56 plus.t17 a_n5644_8799.t34 gnd.t327 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X233 gnd.t229 gnd.t226 gnd.t228 gnd.t227 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X234 a_n3827_n3924.t27 minus.t22 a_n1986_13878.t8 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X235 a_n5644_8799.t1 plus.t18 a_n3827_n3924.t1 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X236 diffpairibias.t5 diffpairibias.t4 gnd.t186 gnd.t185 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X237 CSoutput.t29 commonsourceibias.t90 gnd.t45 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X238 gnd.t135 commonsourceibias.t91 CSoutput.t28 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X239 vdd.t59 vdd.t56 vdd.t58 vdd.t57 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X240 a_n5644_8799.t31 plus.t19 a_n3827_n3924.t48 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X241 a_n3827_n3924.t30 minus.t23 a_n1986_13878.t11 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X242 CSoutput.t27 commonsourceibias.t92 gnd.t111 gnd.t87 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X243 vdd.t55 vdd.t52 vdd.t54 vdd.t53 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X244 a_n1808_13878.t2 a_n1986_13878.t21 a_n1986_13878.t22 vdd.t24 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X245 gnd.t119 commonsourceibias.t93 CSoutput.t26 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X246 vdd.t0 CSoutput.t134 output.t5 gnd.t64 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X247 a_n3827_n3924.t13 diffpairibias.t27 gnd.t125 gnd.t124 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X248 a_n1986_8322.t16 a_n1986_13878.t67 a_n5644_8799.t19 vdd.t34 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X249 gnd.t324 commonsourceibias.t94 CSoutput.t25 gnd.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X250 CSoutput.t24 commonsourceibias.t95 gnd.t100 gnd.t99 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X251 gnd.t47 commonsourceibias.t12 commonsourceibias.t13 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X252 outputibias.t3 outputibias.t2 gnd.t85 gnd.t84 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X253 gnd.t31 commonsourceibias.t96 CSoutput.t23 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X254 a_n3827_n3924.t6 plus.t20 a_n5644_8799.t6 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X255 CSoutput.t104 a_n5644_8799.t72 vdd.t137 vdd.t136 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X256 a_n1986_8322.t4 a_n1986_13878.t68 vdd.t182 vdd.t181 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X257 CSoutput.t22 commonsourceibias.t97 gnd.t326 gnd.t99 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X258 gnd.t94 commonsourceibias.t98 CSoutput.t21 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X259 CSoutput.t20 commonsourceibias.t99 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X260 gnd.t145 commonsourceibias.t100 CSoutput.t19 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X261 gnd.t21 commonsourceibias.t101 CSoutput.t18 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X262 a_n5644_8799.t5 plus.t21 a_n3827_n3924.t5 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X263 commonsourceibias.t11 commonsourceibias.t10 gnd.t144 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X264 a_n3827_n3924.t49 minus.t24 a_n1986_13878.t42 gnd.t159 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X265 gnd.t164 commonsourceibias.t8 commonsourceibias.t9 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X266 vdd.t184 a_n1986_13878.t69 a_n1808_13878.t14 vdd.t183 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X267 output.t4 CSoutput.t135 vdd.t7 gnd.t187 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X268 gnd.t330 commonsourceibias.t102 CSoutput.t17 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X269 CSoutput.t16 commonsourceibias.t103 gnd.t17 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X270 vdd.t51 vdd.t48 vdd.t50 vdd.t49 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X271 a_n1986_8322.t15 a_n1986_13878.t70 a_n5644_8799.t9 vdd.t23 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X272 a_n5644_8799.t17 plus.t22 a_n3827_n3924.t33 gnd.t97 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X273 gnd.t191 commonsourceibias.t6 commonsourceibias.t7 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X274 vdd.t47 vdd.t45 vdd.t46 vdd.t42 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X275 a_n5644_8799.t10 a_n1986_13878.t71 a_n1986_8322.t14 vdd.t24 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X276 a_n1808_13878.t13 a_n1986_13878.t72 vdd.t39 vdd.t38 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X277 vdd.t135 a_n5644_8799.t73 CSoutput.t91 vdd.t134 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X278 CSoutput.t90 a_n5644_8799.t74 vdd.t133 vdd.t132 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X279 CSoutput.t15 commonsourceibias.t104 gnd.t112 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X280 vdd.t15 CSoutput.t136 output.t3 gnd.t188 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X281 output.t2 CSoutput.t137 vdd.t12 gnd.t189 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X282 a_n1986_13878.t5 minus.t25 a_n3827_n3924.t24 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X283 gnd.t53 commonsourceibias.t105 CSoutput.t14 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X284 CSoutput.t13 commonsourceibias.t106 gnd.t197 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X285 a_n3827_n3924.t55 plus.t23 a_n5644_8799.t33 gnd.t120 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X286 gnd.t133 commonsourceibias.t4 commonsourceibias.t5 gnd.t40 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X287 gnd.t22 commonsourceibias.t2 commonsourceibias.t3 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X288 a_n5644_8799.t8 plus.t24 a_n3827_n3924.t9 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X289 CSoutput.t74 a_n5644_8799.t75 vdd.t131 vdd.t125 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X290 a_n1808_13878.t1 a_n1986_13878.t19 a_n1986_13878.t20 vdd.t20 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X291 gnd.t10 commonsourceibias.t107 CSoutput.t12 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X292 CSoutput.t11 commonsourceibias.t108 gnd.t146 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X293 a_n3827_n3924.t12 diffpairibias.t28 gnd.t150 gnd.t149 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X294 a_n3827_n3924.t45 plus.t25 a_n5644_8799.t27 gnd.t153 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X295 vdd.t9 CSoutput.t138 output.t1 gnd.t65 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X296 CSoutput.t73 a_n5644_8799.t76 vdd.t130 vdd.t123 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X297 gnd.t225 gnd.t222 gnd.t224 gnd.t223 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X298 vdd.t129 a_n5644_8799.t77 CSoutput.t110 vdd.t121 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X299 CSoutput.t10 commonsourceibias.t109 gnd.t58 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X300 gnd.t131 commonsourceibias.t110 CSoutput.t9 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X301 diffpairibias.t3 diffpairibias.t2 gnd.t127 gnd.t126 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X302 gnd.t221 gnd.t218 gnd.t220 gnd.t219 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X303 a_n5644_8799.t18 a_n1986_13878.t73 a_n1986_8322.t13 vdd.t40 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X304 a_n1986_13878.t24 a_n1986_13878.t23 a_n1808_13878.t0 vdd.t23 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X305 vdd.t128 a_n5644_8799.t78 CSoutput.t109 vdd.t127 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X306 gnd.t73 commonsourceibias.t111 CSoutput.t8 gnd.t50 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X307 vdd.t2 CSoutput.t139 output.t0 gnd.t66 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X308 CSoutput.t140 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X309 gnd.t217 gnd.t214 gnd.t216 gnd.t215 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X310 vdd.t44 vdd.t41 vdd.t43 vdd.t42 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X311 gnd.t213 gnd.t211 plus.t0 gnd.t212 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X312 CSoutput.t7 commonsourceibias.t112 gnd.t107 gnd.t106 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X313 a_n5644_8799.t16 plus.t26 a_n3827_n3924.t32 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X314 diffpairibias.t1 diffpairibias.t0 gnd.t156 gnd.t155 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X315 minus.t0 gnd.t208 gnd.t210 gnd.t209 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X316 outputibias.t1 outputibias.t0 gnd.t152 gnd.t151 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X317 CSoutput.t141 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X318 gnd.t33 commonsourceibias.t113 CSoutput.t6 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X319 gnd.t207 gnd.t204 gnd.t206 gnd.t205 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X320 vdd.t32 a_n1986_13878.t74 a_n1808_13878.t12 vdd.t31 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X321 CSoutput.t82 a_n5644_8799.t79 vdd.t126 vdd.t125 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X322 a_n1986_13878.t3 minus.t26 a_n3827_n3924.t21 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X323 CSoutput.t5 commonsourceibias.t114 gnd.t91 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X324 gnd.t55 commonsourceibias.t115 CSoutput.t4 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X325 commonsourceibias.t1 commonsourceibias.t0 gnd.t142 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X326 CSoutput.t81 a_n5644_8799.t80 vdd.t124 vdd.t123 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X327 a_n1986_13878.t37 minus.t27 a_n3827_n3924.t34 gnd.t147 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X328 a_n3827_n3924.t2 plus.t27 a_n5644_8799.t2 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X329 CSoutput.t3 commonsourceibias.t116 gnd.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X330 vdd.t122 a_n5644_8799.t81 CSoutput.t89 vdd.t121 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X331 a_n1986_8322.t12 a_n1986_13878.t75 a_n5644_8799.t13 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X332 vdd.t120 a_n5644_8799.t82 CSoutput.t88 vdd.t119 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X333 CSoutput.t96 a_n5644_8799.t83 vdd.t118 vdd.t117 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X334 CSoutput.t2 commonsourceibias.t117 gnd.t173 gnd.t99 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X335 gnd.t69 commonsourceibias.t118 CSoutput.t1 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X336 CSoutput.t0 commonsourceibias.t119 gnd.t37 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X337 a_n3827_n3924.t46 plus.t28 a_n5644_8799.t28 gnd.t175 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X338 a_n1986_13878.t7 minus.t28 a_n3827_n3924.t26 gnd.t95 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X339 a_n3827_n3924.t11 diffpairibias.t29 gnd.t103 gnd.t102 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
R0 gnd.n5604 gnd.n4157 939.716
R1 gnd.n6094 gnd.n643 893.337
R2 gnd.n6724 gnd.n165 838.452
R3 gnd.n6835 gnd.n6734 838.452
R4 gnd.n322 gnd.n273 838.452
R5 gnd.n6328 gnd.n502 838.452
R6 gnd.n1340 gnd.n1329 838.452
R7 gnd.n2600 gnd.n2599 838.452
R8 gnd.n2460 gnd.n1060 838.452
R9 gnd.n4035 gnd.n1133 838.452
R10 gnd.n7041 gnd.n161 783.196
R11 gnd.n7045 gnd.n7044 783.196
R12 gnd.n501 gnd.n500 783.196
R13 gnd.n6532 gnd.n277 783.196
R14 gnd.n3904 gnd.n1333 783.196
R15 gnd.n2296 gnd.n2295 783.196
R16 gnd.n1136 gnd.n1135 783.196
R17 gnd.n4155 gnd.n1064 783.196
R18 gnd.n5512 gnd.n1009 766.379
R19 gnd.n5515 gnd.n5514 766.379
R20 gnd.n4754 gnd.n4657 766.379
R21 gnd.n4750 gnd.n4655 766.379
R22 gnd.n5603 gnd.n4166 756.769
R23 gnd.n5506 gnd.n5505 756.769
R24 gnd.n4847 gnd.n4564 756.769
R25 gnd.n4845 gnd.n4567 756.769
R26 gnd.n2662 gnd.n2104 711.122
R27 gnd.n6354 gnd.n460 711.122
R28 gnd.n2555 gnd.n2101 711.122
R29 gnd.n6356 gnd.n456 711.122
R30 gnd.n5775 gnd.n839 655.866
R31 gnd.n6095 gnd.n644 655.866
R32 gnd.n6309 gnd.n517 655.866
R33 gnd.n2307 gnd.n1007 655.866
R34 gnd.n842 gnd.n839 585
R35 gnd.n5773 gnd.n839 585
R36 gnd.n5771 gnd.n5770 585
R37 gnd.n5772 gnd.n5771 585
R38 gnd.n5769 gnd.n841 585
R39 gnd.n841 gnd.n840 585
R40 gnd.n5768 gnd.n5767 585
R41 gnd.n5767 gnd.n5766 585
R42 gnd.n847 gnd.n846 585
R43 gnd.n5765 gnd.n847 585
R44 gnd.n5763 gnd.n5762 585
R45 gnd.n5764 gnd.n5763 585
R46 gnd.n5761 gnd.n849 585
R47 gnd.n849 gnd.n848 585
R48 gnd.n5760 gnd.n5759 585
R49 gnd.n5759 gnd.n5758 585
R50 gnd.n855 gnd.n854 585
R51 gnd.n5757 gnd.n855 585
R52 gnd.n5755 gnd.n5754 585
R53 gnd.n5756 gnd.n5755 585
R54 gnd.n5753 gnd.n857 585
R55 gnd.n857 gnd.n856 585
R56 gnd.n5752 gnd.n5751 585
R57 gnd.n5751 gnd.n5750 585
R58 gnd.n863 gnd.n862 585
R59 gnd.n5749 gnd.n863 585
R60 gnd.n5747 gnd.n5746 585
R61 gnd.n5748 gnd.n5747 585
R62 gnd.n5745 gnd.n865 585
R63 gnd.n865 gnd.n864 585
R64 gnd.n5744 gnd.n5743 585
R65 gnd.n5743 gnd.n5742 585
R66 gnd.n871 gnd.n870 585
R67 gnd.n5741 gnd.n871 585
R68 gnd.n5739 gnd.n5738 585
R69 gnd.n5740 gnd.n5739 585
R70 gnd.n5737 gnd.n873 585
R71 gnd.n873 gnd.n872 585
R72 gnd.n5736 gnd.n5735 585
R73 gnd.n5735 gnd.n5734 585
R74 gnd.n879 gnd.n878 585
R75 gnd.n5733 gnd.n879 585
R76 gnd.n5731 gnd.n5730 585
R77 gnd.n5732 gnd.n5731 585
R78 gnd.n5729 gnd.n881 585
R79 gnd.n881 gnd.n880 585
R80 gnd.n5728 gnd.n5727 585
R81 gnd.n5727 gnd.n5726 585
R82 gnd.n887 gnd.n886 585
R83 gnd.n5725 gnd.n887 585
R84 gnd.n5723 gnd.n5722 585
R85 gnd.n5724 gnd.n5723 585
R86 gnd.n5721 gnd.n889 585
R87 gnd.n889 gnd.n888 585
R88 gnd.n5720 gnd.n5719 585
R89 gnd.n5719 gnd.n5718 585
R90 gnd.n895 gnd.n894 585
R91 gnd.n5717 gnd.n895 585
R92 gnd.n5715 gnd.n5714 585
R93 gnd.n5716 gnd.n5715 585
R94 gnd.n5713 gnd.n897 585
R95 gnd.n897 gnd.n896 585
R96 gnd.n5712 gnd.n5711 585
R97 gnd.n5711 gnd.n5710 585
R98 gnd.n903 gnd.n902 585
R99 gnd.n5709 gnd.n903 585
R100 gnd.n5707 gnd.n5706 585
R101 gnd.n5708 gnd.n5707 585
R102 gnd.n5705 gnd.n905 585
R103 gnd.n905 gnd.n904 585
R104 gnd.n5704 gnd.n5703 585
R105 gnd.n5703 gnd.n5702 585
R106 gnd.n911 gnd.n910 585
R107 gnd.n5701 gnd.n911 585
R108 gnd.n5699 gnd.n5698 585
R109 gnd.n5700 gnd.n5699 585
R110 gnd.n5697 gnd.n913 585
R111 gnd.n913 gnd.n912 585
R112 gnd.n5696 gnd.n5695 585
R113 gnd.n5695 gnd.n5694 585
R114 gnd.n919 gnd.n918 585
R115 gnd.n5693 gnd.n919 585
R116 gnd.n5691 gnd.n5690 585
R117 gnd.n5692 gnd.n5691 585
R118 gnd.n5689 gnd.n921 585
R119 gnd.n921 gnd.n920 585
R120 gnd.n5688 gnd.n5687 585
R121 gnd.n5687 gnd.n5686 585
R122 gnd.n927 gnd.n926 585
R123 gnd.n5685 gnd.n927 585
R124 gnd.n5683 gnd.n5682 585
R125 gnd.n5684 gnd.n5683 585
R126 gnd.n5681 gnd.n929 585
R127 gnd.n929 gnd.n928 585
R128 gnd.n5680 gnd.n5679 585
R129 gnd.n5679 gnd.n5678 585
R130 gnd.n935 gnd.n934 585
R131 gnd.n5677 gnd.n935 585
R132 gnd.n5675 gnd.n5674 585
R133 gnd.n5676 gnd.n5675 585
R134 gnd.n5673 gnd.n937 585
R135 gnd.n937 gnd.n936 585
R136 gnd.n5672 gnd.n5671 585
R137 gnd.n5671 gnd.n5670 585
R138 gnd.n943 gnd.n942 585
R139 gnd.n5669 gnd.n943 585
R140 gnd.n5667 gnd.n5666 585
R141 gnd.n5668 gnd.n5667 585
R142 gnd.n5665 gnd.n945 585
R143 gnd.n945 gnd.n944 585
R144 gnd.n5664 gnd.n5663 585
R145 gnd.n5663 gnd.n5662 585
R146 gnd.n951 gnd.n950 585
R147 gnd.n5661 gnd.n951 585
R148 gnd.n5659 gnd.n5658 585
R149 gnd.n5660 gnd.n5659 585
R150 gnd.n5657 gnd.n953 585
R151 gnd.n953 gnd.n952 585
R152 gnd.n5656 gnd.n5655 585
R153 gnd.n5655 gnd.n5654 585
R154 gnd.n959 gnd.n958 585
R155 gnd.n5653 gnd.n959 585
R156 gnd.n5651 gnd.n5650 585
R157 gnd.n5652 gnd.n5651 585
R158 gnd.n5649 gnd.n961 585
R159 gnd.n961 gnd.n960 585
R160 gnd.n5648 gnd.n5647 585
R161 gnd.n5647 gnd.n5646 585
R162 gnd.n967 gnd.n966 585
R163 gnd.n5645 gnd.n967 585
R164 gnd.n5643 gnd.n5642 585
R165 gnd.n5644 gnd.n5643 585
R166 gnd.n5641 gnd.n969 585
R167 gnd.n969 gnd.n968 585
R168 gnd.n5640 gnd.n5639 585
R169 gnd.n5639 gnd.n5638 585
R170 gnd.n975 gnd.n974 585
R171 gnd.n5637 gnd.n975 585
R172 gnd.n5635 gnd.n5634 585
R173 gnd.n5636 gnd.n5635 585
R174 gnd.n5633 gnd.n977 585
R175 gnd.n977 gnd.n976 585
R176 gnd.n5632 gnd.n5631 585
R177 gnd.n5631 gnd.n5630 585
R178 gnd.n983 gnd.n982 585
R179 gnd.n5629 gnd.n983 585
R180 gnd.n5627 gnd.n5626 585
R181 gnd.n5628 gnd.n5627 585
R182 gnd.n5625 gnd.n985 585
R183 gnd.n985 gnd.n984 585
R184 gnd.n5624 gnd.n5623 585
R185 gnd.n5623 gnd.n5622 585
R186 gnd.n991 gnd.n990 585
R187 gnd.n5621 gnd.n991 585
R188 gnd.n5619 gnd.n5618 585
R189 gnd.n5620 gnd.n5619 585
R190 gnd.n5617 gnd.n993 585
R191 gnd.n993 gnd.n992 585
R192 gnd.n5616 gnd.n5615 585
R193 gnd.n5615 gnd.n5614 585
R194 gnd.n999 gnd.n998 585
R195 gnd.n5613 gnd.n999 585
R196 gnd.n5611 gnd.n5610 585
R197 gnd.n5612 gnd.n5611 585
R198 gnd.n5609 gnd.n1001 585
R199 gnd.n1001 gnd.n1000 585
R200 gnd.n5608 gnd.n5607 585
R201 gnd.n5607 gnd.n5606 585
R202 gnd.n5776 gnd.n5775 585
R203 gnd.n5775 gnd.n5774 585
R204 gnd.n837 gnd.n836 585
R205 gnd.n836 gnd.n835 585
R206 gnd.n5781 gnd.n5780 585
R207 gnd.n5782 gnd.n5781 585
R208 gnd.n834 gnd.n833 585
R209 gnd.n5783 gnd.n834 585
R210 gnd.n5786 gnd.n5785 585
R211 gnd.n5785 gnd.n5784 585
R212 gnd.n831 gnd.n830 585
R213 gnd.n830 gnd.n829 585
R214 gnd.n5791 gnd.n5790 585
R215 gnd.n5792 gnd.n5791 585
R216 gnd.n828 gnd.n827 585
R217 gnd.n5793 gnd.n828 585
R218 gnd.n5796 gnd.n5795 585
R219 gnd.n5795 gnd.n5794 585
R220 gnd.n825 gnd.n824 585
R221 gnd.n824 gnd.n823 585
R222 gnd.n5801 gnd.n5800 585
R223 gnd.n5802 gnd.n5801 585
R224 gnd.n822 gnd.n821 585
R225 gnd.n5803 gnd.n822 585
R226 gnd.n5806 gnd.n5805 585
R227 gnd.n5805 gnd.n5804 585
R228 gnd.n819 gnd.n818 585
R229 gnd.n818 gnd.n817 585
R230 gnd.n5811 gnd.n5810 585
R231 gnd.n5812 gnd.n5811 585
R232 gnd.n816 gnd.n815 585
R233 gnd.n5813 gnd.n816 585
R234 gnd.n5816 gnd.n5815 585
R235 gnd.n5815 gnd.n5814 585
R236 gnd.n813 gnd.n812 585
R237 gnd.n812 gnd.n811 585
R238 gnd.n5821 gnd.n5820 585
R239 gnd.n5822 gnd.n5821 585
R240 gnd.n810 gnd.n809 585
R241 gnd.n5823 gnd.n810 585
R242 gnd.n5826 gnd.n5825 585
R243 gnd.n5825 gnd.n5824 585
R244 gnd.n807 gnd.n806 585
R245 gnd.n806 gnd.n805 585
R246 gnd.n5831 gnd.n5830 585
R247 gnd.n5832 gnd.n5831 585
R248 gnd.n804 gnd.n803 585
R249 gnd.n5833 gnd.n804 585
R250 gnd.n5836 gnd.n5835 585
R251 gnd.n5835 gnd.n5834 585
R252 gnd.n801 gnd.n800 585
R253 gnd.n800 gnd.n799 585
R254 gnd.n5841 gnd.n5840 585
R255 gnd.n5842 gnd.n5841 585
R256 gnd.n798 gnd.n797 585
R257 gnd.n5843 gnd.n798 585
R258 gnd.n5846 gnd.n5845 585
R259 gnd.n5845 gnd.n5844 585
R260 gnd.n795 gnd.n794 585
R261 gnd.n794 gnd.n793 585
R262 gnd.n5851 gnd.n5850 585
R263 gnd.n5852 gnd.n5851 585
R264 gnd.n792 gnd.n791 585
R265 gnd.n5853 gnd.n792 585
R266 gnd.n5856 gnd.n5855 585
R267 gnd.n5855 gnd.n5854 585
R268 gnd.n789 gnd.n788 585
R269 gnd.n788 gnd.n787 585
R270 gnd.n5861 gnd.n5860 585
R271 gnd.n5862 gnd.n5861 585
R272 gnd.n786 gnd.n785 585
R273 gnd.n5863 gnd.n786 585
R274 gnd.n5866 gnd.n5865 585
R275 gnd.n5865 gnd.n5864 585
R276 gnd.n783 gnd.n782 585
R277 gnd.n782 gnd.n781 585
R278 gnd.n5871 gnd.n5870 585
R279 gnd.n5872 gnd.n5871 585
R280 gnd.n780 gnd.n779 585
R281 gnd.n5873 gnd.n780 585
R282 gnd.n5876 gnd.n5875 585
R283 gnd.n5875 gnd.n5874 585
R284 gnd.n777 gnd.n776 585
R285 gnd.n776 gnd.n775 585
R286 gnd.n5881 gnd.n5880 585
R287 gnd.n5882 gnd.n5881 585
R288 gnd.n774 gnd.n773 585
R289 gnd.n5883 gnd.n774 585
R290 gnd.n5886 gnd.n5885 585
R291 gnd.n5885 gnd.n5884 585
R292 gnd.n771 gnd.n770 585
R293 gnd.n770 gnd.n769 585
R294 gnd.n5891 gnd.n5890 585
R295 gnd.n5892 gnd.n5891 585
R296 gnd.n768 gnd.n767 585
R297 gnd.n5893 gnd.n768 585
R298 gnd.n5896 gnd.n5895 585
R299 gnd.n5895 gnd.n5894 585
R300 gnd.n765 gnd.n764 585
R301 gnd.n764 gnd.n763 585
R302 gnd.n5901 gnd.n5900 585
R303 gnd.n5902 gnd.n5901 585
R304 gnd.n762 gnd.n761 585
R305 gnd.n5903 gnd.n762 585
R306 gnd.n5906 gnd.n5905 585
R307 gnd.n5905 gnd.n5904 585
R308 gnd.n759 gnd.n758 585
R309 gnd.n758 gnd.n757 585
R310 gnd.n5911 gnd.n5910 585
R311 gnd.n5912 gnd.n5911 585
R312 gnd.n756 gnd.n755 585
R313 gnd.n5913 gnd.n756 585
R314 gnd.n5916 gnd.n5915 585
R315 gnd.n5915 gnd.n5914 585
R316 gnd.n753 gnd.n752 585
R317 gnd.n752 gnd.n751 585
R318 gnd.n5921 gnd.n5920 585
R319 gnd.n5922 gnd.n5921 585
R320 gnd.n750 gnd.n749 585
R321 gnd.n5923 gnd.n750 585
R322 gnd.n5926 gnd.n5925 585
R323 gnd.n5925 gnd.n5924 585
R324 gnd.n747 gnd.n746 585
R325 gnd.n746 gnd.n745 585
R326 gnd.n5931 gnd.n5930 585
R327 gnd.n5932 gnd.n5931 585
R328 gnd.n744 gnd.n743 585
R329 gnd.n5933 gnd.n744 585
R330 gnd.n5936 gnd.n5935 585
R331 gnd.n5935 gnd.n5934 585
R332 gnd.n741 gnd.n740 585
R333 gnd.n740 gnd.n739 585
R334 gnd.n5941 gnd.n5940 585
R335 gnd.n5942 gnd.n5941 585
R336 gnd.n738 gnd.n737 585
R337 gnd.n5943 gnd.n738 585
R338 gnd.n5946 gnd.n5945 585
R339 gnd.n5945 gnd.n5944 585
R340 gnd.n735 gnd.n734 585
R341 gnd.n734 gnd.n733 585
R342 gnd.n5951 gnd.n5950 585
R343 gnd.n5952 gnd.n5951 585
R344 gnd.n732 gnd.n731 585
R345 gnd.n5953 gnd.n732 585
R346 gnd.n5956 gnd.n5955 585
R347 gnd.n5955 gnd.n5954 585
R348 gnd.n729 gnd.n728 585
R349 gnd.n728 gnd.n727 585
R350 gnd.n5961 gnd.n5960 585
R351 gnd.n5962 gnd.n5961 585
R352 gnd.n726 gnd.n725 585
R353 gnd.n5963 gnd.n726 585
R354 gnd.n5966 gnd.n5965 585
R355 gnd.n5965 gnd.n5964 585
R356 gnd.n723 gnd.n722 585
R357 gnd.n722 gnd.n721 585
R358 gnd.n5971 gnd.n5970 585
R359 gnd.n5972 gnd.n5971 585
R360 gnd.n720 gnd.n719 585
R361 gnd.n5973 gnd.n720 585
R362 gnd.n5976 gnd.n5975 585
R363 gnd.n5975 gnd.n5974 585
R364 gnd.n717 gnd.n716 585
R365 gnd.n716 gnd.n715 585
R366 gnd.n5981 gnd.n5980 585
R367 gnd.n5982 gnd.n5981 585
R368 gnd.n714 gnd.n713 585
R369 gnd.n5983 gnd.n714 585
R370 gnd.n5986 gnd.n5985 585
R371 gnd.n5985 gnd.n5984 585
R372 gnd.n711 gnd.n710 585
R373 gnd.n710 gnd.n709 585
R374 gnd.n5991 gnd.n5990 585
R375 gnd.n5992 gnd.n5991 585
R376 gnd.n708 gnd.n707 585
R377 gnd.n5993 gnd.n708 585
R378 gnd.n5996 gnd.n5995 585
R379 gnd.n5995 gnd.n5994 585
R380 gnd.n705 gnd.n704 585
R381 gnd.n704 gnd.n703 585
R382 gnd.n6001 gnd.n6000 585
R383 gnd.n6002 gnd.n6001 585
R384 gnd.n702 gnd.n701 585
R385 gnd.n6003 gnd.n702 585
R386 gnd.n6006 gnd.n6005 585
R387 gnd.n6005 gnd.n6004 585
R388 gnd.n699 gnd.n698 585
R389 gnd.n698 gnd.n697 585
R390 gnd.n6011 gnd.n6010 585
R391 gnd.n6012 gnd.n6011 585
R392 gnd.n696 gnd.n695 585
R393 gnd.n6013 gnd.n696 585
R394 gnd.n6016 gnd.n6015 585
R395 gnd.n6015 gnd.n6014 585
R396 gnd.n693 gnd.n692 585
R397 gnd.n692 gnd.n691 585
R398 gnd.n6021 gnd.n6020 585
R399 gnd.n6022 gnd.n6021 585
R400 gnd.n690 gnd.n689 585
R401 gnd.n6023 gnd.n690 585
R402 gnd.n6026 gnd.n6025 585
R403 gnd.n6025 gnd.n6024 585
R404 gnd.n687 gnd.n686 585
R405 gnd.n686 gnd.n685 585
R406 gnd.n6031 gnd.n6030 585
R407 gnd.n6032 gnd.n6031 585
R408 gnd.n684 gnd.n683 585
R409 gnd.n6033 gnd.n684 585
R410 gnd.n6036 gnd.n6035 585
R411 gnd.n6035 gnd.n6034 585
R412 gnd.n681 gnd.n680 585
R413 gnd.n680 gnd.n679 585
R414 gnd.n6041 gnd.n6040 585
R415 gnd.n6042 gnd.n6041 585
R416 gnd.n678 gnd.n677 585
R417 gnd.n6043 gnd.n678 585
R418 gnd.n6046 gnd.n6045 585
R419 gnd.n6045 gnd.n6044 585
R420 gnd.n675 gnd.n674 585
R421 gnd.n674 gnd.n673 585
R422 gnd.n6051 gnd.n6050 585
R423 gnd.n6052 gnd.n6051 585
R424 gnd.n672 gnd.n671 585
R425 gnd.n6053 gnd.n672 585
R426 gnd.n6056 gnd.n6055 585
R427 gnd.n6055 gnd.n6054 585
R428 gnd.n669 gnd.n668 585
R429 gnd.n668 gnd.n667 585
R430 gnd.n6061 gnd.n6060 585
R431 gnd.n6062 gnd.n6061 585
R432 gnd.n666 gnd.n665 585
R433 gnd.n6063 gnd.n666 585
R434 gnd.n6066 gnd.n6065 585
R435 gnd.n6065 gnd.n6064 585
R436 gnd.n663 gnd.n662 585
R437 gnd.n662 gnd.n661 585
R438 gnd.n6071 gnd.n6070 585
R439 gnd.n6072 gnd.n6071 585
R440 gnd.n660 gnd.n659 585
R441 gnd.n6073 gnd.n660 585
R442 gnd.n6076 gnd.n6075 585
R443 gnd.n6075 gnd.n6074 585
R444 gnd.n657 gnd.n656 585
R445 gnd.n656 gnd.n655 585
R446 gnd.n6081 gnd.n6080 585
R447 gnd.n6082 gnd.n6081 585
R448 gnd.n654 gnd.n653 585
R449 gnd.n6083 gnd.n654 585
R450 gnd.n6086 gnd.n6085 585
R451 gnd.n6085 gnd.n6084 585
R452 gnd.n651 gnd.n650 585
R453 gnd.n650 gnd.n649 585
R454 gnd.n6091 gnd.n6090 585
R455 gnd.n6092 gnd.n6091 585
R456 gnd.n648 gnd.n647 585
R457 gnd.n6093 gnd.n648 585
R458 gnd.n6096 gnd.n6095 585
R459 gnd.n6095 gnd.n6094 585
R460 gnd.n6308 gnd.n521 585
R461 gnd.n6308 gnd.n6307 585
R462 gnd.n6301 gnd.n522 585
R463 gnd.n6305 gnd.n522 585
R464 gnd.n6303 gnd.n6302 585
R465 gnd.n6304 gnd.n6303 585
R466 gnd.n525 gnd.n524 585
R467 gnd.n524 gnd.n523 585
R468 gnd.n6296 gnd.n6295 585
R469 gnd.n6295 gnd.n6294 585
R470 gnd.n528 gnd.n527 585
R471 gnd.n6293 gnd.n528 585
R472 gnd.n6291 gnd.n6290 585
R473 gnd.n6292 gnd.n6291 585
R474 gnd.n531 gnd.n530 585
R475 gnd.n530 gnd.n529 585
R476 gnd.n6286 gnd.n6285 585
R477 gnd.n6285 gnd.n6284 585
R478 gnd.n534 gnd.n533 585
R479 gnd.n6283 gnd.n534 585
R480 gnd.n6281 gnd.n6280 585
R481 gnd.n6282 gnd.n6281 585
R482 gnd.n537 gnd.n536 585
R483 gnd.n536 gnd.n535 585
R484 gnd.n6276 gnd.n6275 585
R485 gnd.n6275 gnd.n6274 585
R486 gnd.n540 gnd.n539 585
R487 gnd.n6273 gnd.n540 585
R488 gnd.n6271 gnd.n6270 585
R489 gnd.n6272 gnd.n6271 585
R490 gnd.n543 gnd.n542 585
R491 gnd.n542 gnd.n541 585
R492 gnd.n6266 gnd.n6265 585
R493 gnd.n6265 gnd.n6264 585
R494 gnd.n546 gnd.n545 585
R495 gnd.n6263 gnd.n546 585
R496 gnd.n6261 gnd.n6260 585
R497 gnd.n6262 gnd.n6261 585
R498 gnd.n549 gnd.n548 585
R499 gnd.n548 gnd.n547 585
R500 gnd.n6256 gnd.n6255 585
R501 gnd.n6255 gnd.n6254 585
R502 gnd.n552 gnd.n551 585
R503 gnd.n6253 gnd.n552 585
R504 gnd.n6251 gnd.n6250 585
R505 gnd.n6252 gnd.n6251 585
R506 gnd.n555 gnd.n554 585
R507 gnd.n554 gnd.n553 585
R508 gnd.n6246 gnd.n6245 585
R509 gnd.n6245 gnd.n6244 585
R510 gnd.n558 gnd.n557 585
R511 gnd.n6243 gnd.n558 585
R512 gnd.n6241 gnd.n6240 585
R513 gnd.n6242 gnd.n6241 585
R514 gnd.n561 gnd.n560 585
R515 gnd.n560 gnd.n559 585
R516 gnd.n6236 gnd.n6235 585
R517 gnd.n6235 gnd.n6234 585
R518 gnd.n564 gnd.n563 585
R519 gnd.n6233 gnd.n564 585
R520 gnd.n6231 gnd.n6230 585
R521 gnd.n6232 gnd.n6231 585
R522 gnd.n567 gnd.n566 585
R523 gnd.n566 gnd.n565 585
R524 gnd.n6226 gnd.n6225 585
R525 gnd.n6225 gnd.n6224 585
R526 gnd.n570 gnd.n569 585
R527 gnd.n6223 gnd.n570 585
R528 gnd.n6221 gnd.n6220 585
R529 gnd.n6222 gnd.n6221 585
R530 gnd.n573 gnd.n572 585
R531 gnd.n572 gnd.n571 585
R532 gnd.n6216 gnd.n6215 585
R533 gnd.n6215 gnd.n6214 585
R534 gnd.n576 gnd.n575 585
R535 gnd.n6213 gnd.n576 585
R536 gnd.n6211 gnd.n6210 585
R537 gnd.n6212 gnd.n6211 585
R538 gnd.n579 gnd.n578 585
R539 gnd.n578 gnd.n577 585
R540 gnd.n6206 gnd.n6205 585
R541 gnd.n6205 gnd.n6204 585
R542 gnd.n582 gnd.n581 585
R543 gnd.n6203 gnd.n582 585
R544 gnd.n6201 gnd.n6200 585
R545 gnd.n6202 gnd.n6201 585
R546 gnd.n585 gnd.n584 585
R547 gnd.n584 gnd.n583 585
R548 gnd.n6196 gnd.n6195 585
R549 gnd.n6195 gnd.n6194 585
R550 gnd.n588 gnd.n587 585
R551 gnd.n6193 gnd.n588 585
R552 gnd.n6191 gnd.n6190 585
R553 gnd.n6192 gnd.n6191 585
R554 gnd.n591 gnd.n590 585
R555 gnd.n590 gnd.n589 585
R556 gnd.n6186 gnd.n6185 585
R557 gnd.n6185 gnd.n6184 585
R558 gnd.n594 gnd.n593 585
R559 gnd.n6183 gnd.n594 585
R560 gnd.n6181 gnd.n6180 585
R561 gnd.n6182 gnd.n6181 585
R562 gnd.n597 gnd.n596 585
R563 gnd.n596 gnd.n595 585
R564 gnd.n6176 gnd.n6175 585
R565 gnd.n6175 gnd.n6174 585
R566 gnd.n600 gnd.n599 585
R567 gnd.n6173 gnd.n600 585
R568 gnd.n6171 gnd.n6170 585
R569 gnd.n6172 gnd.n6171 585
R570 gnd.n603 gnd.n602 585
R571 gnd.n602 gnd.n601 585
R572 gnd.n6166 gnd.n6165 585
R573 gnd.n6165 gnd.n6164 585
R574 gnd.n606 gnd.n605 585
R575 gnd.n6163 gnd.n606 585
R576 gnd.n6161 gnd.n6160 585
R577 gnd.n6162 gnd.n6161 585
R578 gnd.n609 gnd.n608 585
R579 gnd.n608 gnd.n607 585
R580 gnd.n6156 gnd.n6155 585
R581 gnd.n6155 gnd.n6154 585
R582 gnd.n612 gnd.n611 585
R583 gnd.n6153 gnd.n612 585
R584 gnd.n6151 gnd.n6150 585
R585 gnd.n6152 gnd.n6151 585
R586 gnd.n615 gnd.n614 585
R587 gnd.n614 gnd.n613 585
R588 gnd.n6146 gnd.n6145 585
R589 gnd.n6145 gnd.n6144 585
R590 gnd.n618 gnd.n617 585
R591 gnd.n6143 gnd.n618 585
R592 gnd.n6141 gnd.n6140 585
R593 gnd.n6142 gnd.n6141 585
R594 gnd.n621 gnd.n620 585
R595 gnd.n620 gnd.n619 585
R596 gnd.n6136 gnd.n6135 585
R597 gnd.n6135 gnd.n6134 585
R598 gnd.n624 gnd.n623 585
R599 gnd.n6133 gnd.n624 585
R600 gnd.n6131 gnd.n6130 585
R601 gnd.n6132 gnd.n6131 585
R602 gnd.n627 gnd.n626 585
R603 gnd.n626 gnd.n625 585
R604 gnd.n6126 gnd.n6125 585
R605 gnd.n6125 gnd.n6124 585
R606 gnd.n630 gnd.n629 585
R607 gnd.n6123 gnd.n630 585
R608 gnd.n6121 gnd.n6120 585
R609 gnd.n6122 gnd.n6121 585
R610 gnd.n633 gnd.n632 585
R611 gnd.n632 gnd.n631 585
R612 gnd.n6116 gnd.n6115 585
R613 gnd.n6115 gnd.n6114 585
R614 gnd.n636 gnd.n635 585
R615 gnd.n6113 gnd.n636 585
R616 gnd.n6111 gnd.n6110 585
R617 gnd.n6112 gnd.n6111 585
R618 gnd.n639 gnd.n638 585
R619 gnd.n638 gnd.n637 585
R620 gnd.n6106 gnd.n6105 585
R621 gnd.n6105 gnd.n6104 585
R622 gnd.n642 gnd.n641 585
R623 gnd.n6103 gnd.n642 585
R624 gnd.n6101 gnd.n6100 585
R625 gnd.n6102 gnd.n6101 585
R626 gnd.n645 gnd.n644 585
R627 gnd.n644 gnd.n643 585
R628 gnd.n1329 gnd.n1328 585
R629 gnd.n2598 gnd.n1329 585
R630 gnd.n3913 gnd.n3912 585
R631 gnd.n3912 gnd.n3911 585
R632 gnd.n3914 gnd.n1324 585
R633 gnd.n2565 gnd.n1324 585
R634 gnd.n3916 gnd.n3915 585
R635 gnd.n3917 gnd.n3916 585
R636 gnd.n1308 gnd.n1307 585
R637 gnd.n2543 gnd.n1308 585
R638 gnd.n3925 gnd.n3924 585
R639 gnd.n3924 gnd.n3923 585
R640 gnd.n3926 gnd.n1303 585
R641 gnd.n2531 gnd.n1303 585
R642 gnd.n3928 gnd.n3927 585
R643 gnd.n3929 gnd.n3928 585
R644 gnd.n1288 gnd.n1287 585
R645 gnd.n1299 gnd.n1288 585
R646 gnd.n3937 gnd.n3936 585
R647 gnd.n3936 gnd.n3935 585
R648 gnd.n3938 gnd.n1283 585
R649 gnd.n1283 gnd.n1282 585
R650 gnd.n3940 gnd.n3939 585
R651 gnd.n3941 gnd.n3940 585
R652 gnd.n1268 gnd.n1267 585
R653 gnd.n1272 gnd.n1268 585
R654 gnd.n3949 gnd.n3948 585
R655 gnd.n3948 gnd.n3947 585
R656 gnd.n3950 gnd.n1263 585
R657 gnd.n1269 gnd.n1263 585
R658 gnd.n3952 gnd.n3951 585
R659 gnd.n3953 gnd.n3952 585
R660 gnd.n1250 gnd.n1249 585
R661 gnd.n1253 gnd.n1250 585
R662 gnd.n3961 gnd.n3960 585
R663 gnd.n3960 gnd.n3959 585
R664 gnd.n3962 gnd.n1245 585
R665 gnd.n1245 gnd.n1244 585
R666 gnd.n3964 gnd.n3963 585
R667 gnd.n3965 gnd.n3964 585
R668 gnd.n1230 gnd.n1229 585
R669 gnd.n1234 gnd.n1230 585
R670 gnd.n3973 gnd.n3972 585
R671 gnd.n3972 gnd.n3971 585
R672 gnd.n3974 gnd.n1225 585
R673 gnd.n1231 gnd.n1225 585
R674 gnd.n3976 gnd.n3975 585
R675 gnd.n3977 gnd.n3976 585
R676 gnd.n1212 gnd.n1211 585
R677 gnd.n1222 gnd.n1212 585
R678 gnd.n3985 gnd.n3984 585
R679 gnd.n3984 gnd.n3983 585
R680 gnd.n3986 gnd.n1207 585
R681 gnd.n1207 gnd.n1206 585
R682 gnd.n3988 gnd.n3987 585
R683 gnd.n3989 gnd.n3988 585
R684 gnd.n1192 gnd.n1191 585
R685 gnd.n1196 gnd.n1192 585
R686 gnd.n3997 gnd.n3996 585
R687 gnd.n3996 gnd.n3995 585
R688 gnd.n3998 gnd.n1187 585
R689 gnd.n1193 gnd.n1187 585
R690 gnd.n4000 gnd.n3999 585
R691 gnd.n4001 gnd.n4000 585
R692 gnd.n1174 gnd.n1173 585
R693 gnd.n1184 gnd.n1174 585
R694 gnd.n4009 gnd.n4008 585
R695 gnd.n4008 gnd.n4007 585
R696 gnd.n4010 gnd.n1169 585
R697 gnd.n1169 gnd.n1168 585
R698 gnd.n4012 gnd.n4011 585
R699 gnd.n4013 gnd.n4012 585
R700 gnd.n1156 gnd.n1155 585
R701 gnd.n1159 gnd.n1156 585
R702 gnd.n4021 gnd.n4020 585
R703 gnd.n4020 gnd.n4019 585
R704 gnd.n4022 gnd.n1150 585
R705 gnd.n1150 gnd.n1149 585
R706 gnd.n4024 gnd.n4023 585
R707 gnd.n4025 gnd.n4024 585
R708 gnd.n1151 gnd.n1134 585
R709 gnd.n1146 gnd.n1134 585
R710 gnd.n4034 gnd.n1132 585
R711 gnd.n4034 gnd.n4033 585
R712 gnd.n4036 gnd.n4035 585
R713 gnd.n4035 gnd.n1061 585
R714 gnd.n2417 gnd.n1133 585
R715 gnd.n2419 gnd.n2418 585
R716 gnd.n2421 gnd.n2420 585
R717 gnd.n2425 gnd.n2415 585
R718 gnd.n2427 gnd.n2426 585
R719 gnd.n2429 gnd.n2428 585
R720 gnd.n2431 gnd.n2430 585
R721 gnd.n2435 gnd.n2413 585
R722 gnd.n2437 gnd.n2436 585
R723 gnd.n2439 gnd.n2438 585
R724 gnd.n2441 gnd.n2440 585
R725 gnd.n2445 gnd.n2411 585
R726 gnd.n2447 gnd.n2446 585
R727 gnd.n2449 gnd.n2448 585
R728 gnd.n2451 gnd.n2450 585
R729 gnd.n2408 gnd.n2407 585
R730 gnd.n2455 gnd.n2409 585
R731 gnd.n2456 gnd.n2404 585
R732 gnd.n2457 gnd.n1060 585
R733 gnd.n4157 gnd.n1060 585
R734 gnd.n2601 gnd.n2600 585
R735 gnd.n2602 gnd.n2197 585
R736 gnd.n2603 gnd.n2193 585
R737 gnd.n2184 gnd.n2183 585
R738 gnd.n2610 gnd.n2182 585
R739 gnd.n2611 gnd.n2181 585
R740 gnd.n2180 gnd.n2174 585
R741 gnd.n2618 gnd.n2173 585
R742 gnd.n2619 gnd.n2172 585
R743 gnd.n2164 gnd.n2163 585
R744 gnd.n2626 gnd.n2162 585
R745 gnd.n2627 gnd.n2161 585
R746 gnd.n2160 gnd.n2154 585
R747 gnd.n2634 gnd.n2153 585
R748 gnd.n2635 gnd.n2152 585
R749 gnd.n2144 gnd.n2143 585
R750 gnd.n2642 gnd.n2142 585
R751 gnd.n2643 gnd.n2141 585
R752 gnd.n2140 gnd.n1340 585
R753 gnd.n3903 gnd.n1340 585
R754 gnd.n2599 gnd.n2199 585
R755 gnd.n2599 gnd.n2598 585
R756 gnd.n2318 gnd.n1331 585
R757 gnd.n3911 gnd.n1331 585
R758 gnd.n2564 gnd.n2563 585
R759 gnd.n2565 gnd.n2564 585
R760 gnd.n2317 gnd.n1322 585
R761 gnd.n3917 gnd.n1322 585
R762 gnd.n2545 gnd.n2544 585
R763 gnd.n2544 gnd.n2543 585
R764 gnd.n2320 gnd.n1311 585
R765 gnd.n3923 gnd.n1311 585
R766 gnd.n2530 gnd.n2529 585
R767 gnd.n2531 gnd.n2530 585
R768 gnd.n2382 gnd.n1301 585
R769 gnd.n3929 gnd.n1301 585
R770 gnd.n2525 gnd.n2524 585
R771 gnd.n2524 gnd.n1299 585
R772 gnd.n2523 gnd.n1290 585
R773 gnd.n3935 gnd.n1290 585
R774 gnd.n2522 gnd.n2385 585
R775 gnd.n2385 gnd.n1282 585
R776 gnd.n2384 gnd.n1281 585
R777 gnd.n3941 gnd.n1281 585
R778 gnd.n2518 gnd.n2517 585
R779 gnd.n2517 gnd.n1272 585
R780 gnd.n2516 gnd.n1271 585
R781 gnd.n3947 gnd.n1271 585
R782 gnd.n2515 gnd.n2388 585
R783 gnd.n2388 gnd.n1269 585
R784 gnd.n2387 gnd.n1262 585
R785 gnd.n3953 gnd.n1262 585
R786 gnd.n2511 gnd.n2510 585
R787 gnd.n2510 gnd.n1253 585
R788 gnd.n2509 gnd.n1252 585
R789 gnd.n3959 gnd.n1252 585
R790 gnd.n2508 gnd.n2391 585
R791 gnd.n2391 gnd.n1244 585
R792 gnd.n2390 gnd.n1243 585
R793 gnd.n3965 gnd.n1243 585
R794 gnd.n2504 gnd.n2503 585
R795 gnd.n2503 gnd.n1234 585
R796 gnd.n2502 gnd.n1233 585
R797 gnd.n3971 gnd.n1233 585
R798 gnd.n2501 gnd.n2500 585
R799 gnd.n2500 gnd.n1231 585
R800 gnd.n2393 gnd.n1224 585
R801 gnd.n3977 gnd.n1224 585
R802 gnd.n2496 gnd.n2495 585
R803 gnd.n2495 gnd.n1222 585
R804 gnd.n2494 gnd.n1214 585
R805 gnd.n3983 gnd.n1214 585
R806 gnd.n2493 gnd.n2492 585
R807 gnd.n2492 gnd.n1206 585
R808 gnd.n2395 gnd.n1205 585
R809 gnd.n3989 gnd.n1205 585
R810 gnd.n2488 gnd.n2487 585
R811 gnd.n2487 gnd.n1196 585
R812 gnd.n2486 gnd.n1195 585
R813 gnd.n3995 gnd.n1195 585
R814 gnd.n2485 gnd.n2484 585
R815 gnd.n2484 gnd.n1193 585
R816 gnd.n2397 gnd.n1186 585
R817 gnd.n4001 gnd.n1186 585
R818 gnd.n2480 gnd.n2479 585
R819 gnd.n2479 gnd.n1184 585
R820 gnd.n2478 gnd.n1176 585
R821 gnd.n4007 gnd.n1176 585
R822 gnd.n2477 gnd.n2476 585
R823 gnd.n2476 gnd.n1168 585
R824 gnd.n2399 gnd.n1167 585
R825 gnd.n4013 gnd.n1167 585
R826 gnd.n2472 gnd.n2471 585
R827 gnd.n2471 gnd.n1159 585
R828 gnd.n2470 gnd.n1158 585
R829 gnd.n4019 gnd.n1158 585
R830 gnd.n2469 gnd.n2468 585
R831 gnd.n2468 gnd.n1149 585
R832 gnd.n2401 gnd.n1148 585
R833 gnd.n4025 gnd.n1148 585
R834 gnd.n2464 gnd.n2463 585
R835 gnd.n2463 gnd.n1146 585
R836 gnd.n2462 gnd.n1138 585
R837 gnd.n4033 gnd.n1138 585
R838 gnd.n2461 gnd.n2460 585
R839 gnd.n2460 gnd.n1061 585
R840 gnd.n5512 gnd.n5511 585
R841 gnd.n5513 gnd.n5512 585
R842 gnd.n4219 gnd.n4218 585
R843 gnd.n4225 gnd.n4218 585
R844 gnd.n5487 gnd.n4237 585
R845 gnd.n4237 gnd.n4224 585
R846 gnd.n5489 gnd.n5488 585
R847 gnd.n5490 gnd.n5489 585
R848 gnd.n4238 gnd.n4236 585
R849 gnd.n4236 gnd.n4232 585
R850 gnd.n5221 gnd.n5220 585
R851 gnd.n5220 gnd.n5219 585
R852 gnd.n4243 gnd.n4242 585
R853 gnd.n5190 gnd.n4243 585
R854 gnd.n5210 gnd.n5209 585
R855 gnd.n5209 gnd.n5208 585
R856 gnd.n4250 gnd.n4249 585
R857 gnd.n5196 gnd.n4250 585
R858 gnd.n5166 gnd.n4270 585
R859 gnd.n4270 gnd.n4269 585
R860 gnd.n5168 gnd.n5167 585
R861 gnd.n5169 gnd.n5168 585
R862 gnd.n4271 gnd.n4268 585
R863 gnd.n4279 gnd.n4268 585
R864 gnd.n5144 gnd.n4291 585
R865 gnd.n4291 gnd.n4278 585
R866 gnd.n5146 gnd.n5145 585
R867 gnd.n5147 gnd.n5146 585
R868 gnd.n4292 gnd.n4290 585
R869 gnd.n4290 gnd.n4286 585
R870 gnd.n5132 gnd.n5131 585
R871 gnd.n5131 gnd.n5130 585
R872 gnd.n4297 gnd.n4296 585
R873 gnd.n4307 gnd.n4297 585
R874 gnd.n5121 gnd.n5120 585
R875 gnd.n5120 gnd.n5119 585
R876 gnd.n4304 gnd.n4303 585
R877 gnd.n5107 gnd.n4304 585
R878 gnd.n5081 gnd.n4325 585
R879 gnd.n4325 gnd.n4314 585
R880 gnd.n5083 gnd.n5082 585
R881 gnd.n5084 gnd.n5083 585
R882 gnd.n4326 gnd.n4324 585
R883 gnd.n4334 gnd.n4324 585
R884 gnd.n5059 gnd.n4346 585
R885 gnd.n4346 gnd.n4333 585
R886 gnd.n5061 gnd.n5060 585
R887 gnd.n5062 gnd.n5061 585
R888 gnd.n4347 gnd.n4345 585
R889 gnd.n4345 gnd.n4341 585
R890 gnd.n5047 gnd.n5046 585
R891 gnd.n5046 gnd.n5045 585
R892 gnd.n4352 gnd.n4351 585
R893 gnd.n4361 gnd.n4352 585
R894 gnd.n5036 gnd.n5035 585
R895 gnd.n5035 gnd.n5034 585
R896 gnd.n4359 gnd.n4358 585
R897 gnd.n5022 gnd.n4359 585
R898 gnd.n4460 gnd.n4459 585
R899 gnd.n4460 gnd.n4368 585
R900 gnd.n4979 gnd.n4978 585
R901 gnd.n4978 gnd.n4977 585
R902 gnd.n4980 gnd.n4454 585
R903 gnd.n4465 gnd.n4454 585
R904 gnd.n4982 gnd.n4981 585
R905 gnd.n4983 gnd.n4982 585
R906 gnd.n4455 gnd.n4453 585
R907 gnd.n4478 gnd.n4453 585
R908 gnd.n4438 gnd.n4437 585
R909 gnd.n4441 gnd.n4438 585
R910 gnd.n4993 gnd.n4992 585
R911 gnd.n4992 gnd.n4991 585
R912 gnd.n4994 gnd.n4432 585
R913 gnd.n4953 gnd.n4432 585
R914 gnd.n4996 gnd.n4995 585
R915 gnd.n4997 gnd.n4996 585
R916 gnd.n4433 gnd.n4431 585
R917 gnd.n4492 gnd.n4431 585
R918 gnd.n4945 gnd.n4944 585
R919 gnd.n4944 gnd.n4943 585
R920 gnd.n4489 gnd.n4488 585
R921 gnd.n4927 gnd.n4489 585
R922 gnd.n4914 gnd.n4508 585
R923 gnd.n4508 gnd.n4507 585
R924 gnd.n4916 gnd.n4915 585
R925 gnd.n4917 gnd.n4916 585
R926 gnd.n4509 gnd.n4506 585
R927 gnd.n4515 gnd.n4506 585
R928 gnd.n4895 gnd.n4894 585
R929 gnd.n4896 gnd.n4895 585
R930 gnd.n4526 gnd.n4525 585
R931 gnd.n4525 gnd.n4521 585
R932 gnd.n4885 gnd.n4884 585
R933 gnd.n4886 gnd.n4885 585
R934 gnd.n4536 gnd.n4535 585
R935 gnd.n4541 gnd.n4535 585
R936 gnd.n4863 gnd.n4554 585
R937 gnd.n4554 gnd.n4540 585
R938 gnd.n4865 gnd.n4864 585
R939 gnd.n4866 gnd.n4865 585
R940 gnd.n4555 gnd.n4553 585
R941 gnd.n4553 gnd.n4549 585
R942 gnd.n4854 gnd.n4853 585
R943 gnd.n4855 gnd.n4854 585
R944 gnd.n4562 gnd.n4561 585
R945 gnd.n4566 gnd.n4561 585
R946 gnd.n4831 gnd.n4583 585
R947 gnd.n4583 gnd.n4565 585
R948 gnd.n4833 gnd.n4832 585
R949 gnd.n4834 gnd.n4833 585
R950 gnd.n4584 gnd.n4582 585
R951 gnd.n4582 gnd.n4573 585
R952 gnd.n4826 gnd.n4825 585
R953 gnd.n4825 gnd.n4824 585
R954 gnd.n4631 gnd.n4630 585
R955 gnd.n4632 gnd.n4631 585
R956 gnd.n4785 gnd.n4784 585
R957 gnd.n4786 gnd.n4785 585
R958 gnd.n4641 gnd.n4640 585
R959 gnd.n4640 gnd.n4639 585
R960 gnd.n4780 gnd.n4779 585
R961 gnd.n4779 gnd.n4778 585
R962 gnd.n4644 gnd.n4643 585
R963 gnd.n4645 gnd.n4644 585
R964 gnd.n4769 gnd.n4768 585
R965 gnd.n4770 gnd.n4769 585
R966 gnd.n4652 gnd.n4651 585
R967 gnd.n4761 gnd.n4651 585
R968 gnd.n4764 gnd.n4763 585
R969 gnd.n4763 gnd.n4762 585
R970 gnd.n4655 gnd.n4654 585
R971 gnd.n4656 gnd.n4655 585
R972 gnd.n4750 gnd.n4749 585
R973 gnd.n4748 gnd.n4674 585
R974 gnd.n4747 gnd.n4673 585
R975 gnd.n4752 gnd.n4673 585
R976 gnd.n4746 gnd.n4745 585
R977 gnd.n4744 gnd.n4743 585
R978 gnd.n4742 gnd.n4741 585
R979 gnd.n4740 gnd.n4739 585
R980 gnd.n4738 gnd.n4737 585
R981 gnd.n4736 gnd.n4735 585
R982 gnd.n4734 gnd.n4733 585
R983 gnd.n4732 gnd.n4731 585
R984 gnd.n4730 gnd.n4729 585
R985 gnd.n4728 gnd.n4727 585
R986 gnd.n4726 gnd.n4725 585
R987 gnd.n4724 gnd.n4723 585
R988 gnd.n4722 gnd.n4721 585
R989 gnd.n4720 gnd.n4719 585
R990 gnd.n4718 gnd.n4717 585
R991 gnd.n4716 gnd.n4715 585
R992 gnd.n4714 gnd.n4713 585
R993 gnd.n4712 gnd.n4711 585
R994 gnd.n4710 gnd.n4709 585
R995 gnd.n4708 gnd.n4707 585
R996 gnd.n4706 gnd.n4705 585
R997 gnd.n4704 gnd.n4703 585
R998 gnd.n4661 gnd.n4660 585
R999 gnd.n4755 gnd.n4754 585
R1000 gnd.n5516 gnd.n5515 585
R1001 gnd.n5518 gnd.n5517 585
R1002 gnd.n5520 gnd.n5519 585
R1003 gnd.n5522 gnd.n5521 585
R1004 gnd.n5524 gnd.n5523 585
R1005 gnd.n5526 gnd.n5525 585
R1006 gnd.n5528 gnd.n5527 585
R1007 gnd.n5530 gnd.n5529 585
R1008 gnd.n5532 gnd.n5531 585
R1009 gnd.n5534 gnd.n5533 585
R1010 gnd.n5536 gnd.n5535 585
R1011 gnd.n5538 gnd.n5537 585
R1012 gnd.n5540 gnd.n5539 585
R1013 gnd.n5542 gnd.n5541 585
R1014 gnd.n5544 gnd.n5543 585
R1015 gnd.n5546 gnd.n5545 585
R1016 gnd.n5548 gnd.n5547 585
R1017 gnd.n5550 gnd.n5549 585
R1018 gnd.n5552 gnd.n5551 585
R1019 gnd.n5554 gnd.n5553 585
R1020 gnd.n5556 gnd.n5555 585
R1021 gnd.n5558 gnd.n5557 585
R1022 gnd.n5560 gnd.n5559 585
R1023 gnd.n5562 gnd.n5561 585
R1024 gnd.n5564 gnd.n5563 585
R1025 gnd.n5565 gnd.n4186 585
R1026 gnd.n5566 gnd.n1009 585
R1027 gnd.n5604 gnd.n1009 585
R1028 gnd.n5514 gnd.n4216 585
R1029 gnd.n5514 gnd.n5513 585
R1030 gnd.n5183 gnd.n4215 585
R1031 gnd.n4225 gnd.n4215 585
R1032 gnd.n5185 gnd.n5184 585
R1033 gnd.n5184 gnd.n4224 585
R1034 gnd.n5186 gnd.n4234 585
R1035 gnd.n5490 gnd.n4234 585
R1036 gnd.n5188 gnd.n5187 585
R1037 gnd.n5187 gnd.n4232 585
R1038 gnd.n5189 gnd.n4245 585
R1039 gnd.n5219 gnd.n4245 585
R1040 gnd.n5192 gnd.n5191 585
R1041 gnd.n5191 gnd.n5190 585
R1042 gnd.n5193 gnd.n4252 585
R1043 gnd.n5208 gnd.n4252 585
R1044 gnd.n5195 gnd.n5194 585
R1045 gnd.n5196 gnd.n5195 585
R1046 gnd.n4262 gnd.n4261 585
R1047 gnd.n4269 gnd.n4261 585
R1048 gnd.n5171 gnd.n5170 585
R1049 gnd.n5170 gnd.n5169 585
R1050 gnd.n4265 gnd.n4264 585
R1051 gnd.n4279 gnd.n4265 585
R1052 gnd.n5097 gnd.n5096 585
R1053 gnd.n5096 gnd.n4278 585
R1054 gnd.n5098 gnd.n4288 585
R1055 gnd.n5147 gnd.n4288 585
R1056 gnd.n5100 gnd.n5099 585
R1057 gnd.n5099 gnd.n4286 585
R1058 gnd.n5101 gnd.n4299 585
R1059 gnd.n5130 gnd.n4299 585
R1060 gnd.n5103 gnd.n5102 585
R1061 gnd.n5102 gnd.n4307 585
R1062 gnd.n5104 gnd.n4306 585
R1063 gnd.n5119 gnd.n4306 585
R1064 gnd.n5106 gnd.n5105 585
R1065 gnd.n5107 gnd.n5106 585
R1066 gnd.n4318 gnd.n4317 585
R1067 gnd.n4317 gnd.n4314 585
R1068 gnd.n5086 gnd.n5085 585
R1069 gnd.n5085 gnd.n5084 585
R1070 gnd.n4321 gnd.n4320 585
R1071 gnd.n4334 gnd.n4321 585
R1072 gnd.n5010 gnd.n5009 585
R1073 gnd.n5009 gnd.n4333 585
R1074 gnd.n5011 gnd.n4343 585
R1075 gnd.n5062 gnd.n4343 585
R1076 gnd.n5013 gnd.n5012 585
R1077 gnd.n5012 gnd.n4341 585
R1078 gnd.n5014 gnd.n4354 585
R1079 gnd.n5045 gnd.n4354 585
R1080 gnd.n5016 gnd.n5015 585
R1081 gnd.n5015 gnd.n4361 585
R1082 gnd.n5017 gnd.n4360 585
R1083 gnd.n5034 gnd.n4360 585
R1084 gnd.n5019 gnd.n5018 585
R1085 gnd.n5022 gnd.n5019 585
R1086 gnd.n4371 gnd.n4370 585
R1087 gnd.n4370 gnd.n4368 585
R1088 gnd.n4462 gnd.n4461 585
R1089 gnd.n4977 gnd.n4461 585
R1090 gnd.n4464 gnd.n4463 585
R1091 gnd.n4465 gnd.n4464 585
R1092 gnd.n4475 gnd.n4451 585
R1093 gnd.n4983 gnd.n4451 585
R1094 gnd.n4477 gnd.n4476 585
R1095 gnd.n4478 gnd.n4477 585
R1096 gnd.n4474 gnd.n4473 585
R1097 gnd.n4474 gnd.n4441 585
R1098 gnd.n4472 gnd.n4439 585
R1099 gnd.n4991 gnd.n4439 585
R1100 gnd.n4428 gnd.n4426 585
R1101 gnd.n4953 gnd.n4428 585
R1102 gnd.n4999 gnd.n4998 585
R1103 gnd.n4998 gnd.n4997 585
R1104 gnd.n4427 gnd.n4425 585
R1105 gnd.n4492 gnd.n4427 585
R1106 gnd.n4924 gnd.n4491 585
R1107 gnd.n4943 gnd.n4491 585
R1108 gnd.n4926 gnd.n4925 585
R1109 gnd.n4927 gnd.n4926 585
R1110 gnd.n4501 gnd.n4500 585
R1111 gnd.n4507 gnd.n4500 585
R1112 gnd.n4919 gnd.n4918 585
R1113 gnd.n4918 gnd.n4917 585
R1114 gnd.n4504 gnd.n4503 585
R1115 gnd.n4515 gnd.n4504 585
R1116 gnd.n4804 gnd.n4523 585
R1117 gnd.n4896 gnd.n4523 585
R1118 gnd.n4806 gnd.n4805 585
R1119 gnd.n4805 gnd.n4521 585
R1120 gnd.n4807 gnd.n4534 585
R1121 gnd.n4886 gnd.n4534 585
R1122 gnd.n4809 gnd.n4808 585
R1123 gnd.n4809 gnd.n4541 585
R1124 gnd.n4811 gnd.n4810 585
R1125 gnd.n4810 gnd.n4540 585
R1126 gnd.n4812 gnd.n4551 585
R1127 gnd.n4866 gnd.n4551 585
R1128 gnd.n4814 gnd.n4813 585
R1129 gnd.n4813 gnd.n4549 585
R1130 gnd.n4815 gnd.n4560 585
R1131 gnd.n4855 gnd.n4560 585
R1132 gnd.n4817 gnd.n4816 585
R1133 gnd.n4817 gnd.n4566 585
R1134 gnd.n4819 gnd.n4818 585
R1135 gnd.n4818 gnd.n4565 585
R1136 gnd.n4820 gnd.n4581 585
R1137 gnd.n4834 gnd.n4581 585
R1138 gnd.n4821 gnd.n4634 585
R1139 gnd.n4634 gnd.n4573 585
R1140 gnd.n4823 gnd.n4822 585
R1141 gnd.n4824 gnd.n4823 585
R1142 gnd.n4635 gnd.n4633 585
R1143 gnd.n4633 gnd.n4632 585
R1144 gnd.n4788 gnd.n4787 585
R1145 gnd.n4787 gnd.n4786 585
R1146 gnd.n4638 gnd.n4637 585
R1147 gnd.n4639 gnd.n4638 585
R1148 gnd.n4777 gnd.n4776 585
R1149 gnd.n4778 gnd.n4777 585
R1150 gnd.n4647 gnd.n4646 585
R1151 gnd.n4646 gnd.n4645 585
R1152 gnd.n4772 gnd.n4771 585
R1153 gnd.n4771 gnd.n4770 585
R1154 gnd.n4650 gnd.n4649 585
R1155 gnd.n4761 gnd.n4650 585
R1156 gnd.n4760 gnd.n4759 585
R1157 gnd.n4762 gnd.n4760 585
R1158 gnd.n4658 gnd.n4657 585
R1159 gnd.n4657 gnd.n4656 585
R1160 gnd.n7050 gnd.n165 585
R1161 gnd.n165 gnd.n164 585
R1162 gnd.n7052 gnd.n7051 585
R1163 gnd.n7053 gnd.n7052 585
R1164 gnd.n151 gnd.n150 585
R1165 gnd.n154 gnd.n151 585
R1166 gnd.n7061 gnd.n7060 585
R1167 gnd.n7060 gnd.n7059 585
R1168 gnd.n7062 gnd.n146 585
R1169 gnd.n146 gnd.n145 585
R1170 gnd.n7064 gnd.n7063 585
R1171 gnd.n7065 gnd.n7064 585
R1172 gnd.n132 gnd.n131 585
R1173 gnd.n142 gnd.n132 585
R1174 gnd.n7073 gnd.n7072 585
R1175 gnd.n7072 gnd.n7071 585
R1176 gnd.n7074 gnd.n127 585
R1177 gnd.n127 gnd.n126 585
R1178 gnd.n7076 gnd.n7075 585
R1179 gnd.n7077 gnd.n7076 585
R1180 gnd.n113 gnd.n112 585
R1181 gnd.n116 gnd.n113 585
R1182 gnd.n7085 gnd.n7084 585
R1183 gnd.n7084 gnd.n7083 585
R1184 gnd.n7086 gnd.n108 585
R1185 gnd.n108 gnd.n107 585
R1186 gnd.n7088 gnd.n7087 585
R1187 gnd.n7089 gnd.n7088 585
R1188 gnd.n94 gnd.n93 585
R1189 gnd.n104 gnd.n94 585
R1190 gnd.n7097 gnd.n7096 585
R1191 gnd.n7096 gnd.n7095 585
R1192 gnd.n7098 gnd.n88 585
R1193 gnd.n88 gnd.n86 585
R1194 gnd.n7100 gnd.n7099 585
R1195 gnd.n7101 gnd.n7100 585
R1196 gnd.n89 gnd.n87 585
R1197 gnd.n87 gnd.n74 585
R1198 gnd.n6683 gnd.n75 585
R1199 gnd.n7107 gnd.n75 585
R1200 gnd.n6682 gnd.n6681 585
R1201 gnd.n6681 gnd.n6680 585
R1202 gnd.n170 gnd.n169 585
R1203 gnd.n171 gnd.n170 585
R1204 gnd.n6674 gnd.n6673 585
R1205 gnd.n6673 gnd.n6672 585
R1206 gnd.n176 gnd.n175 585
R1207 gnd.n188 gnd.n176 585
R1208 gnd.n6660 gnd.n6659 585
R1209 gnd.n6661 gnd.n6660 585
R1210 gnd.n190 gnd.n189 585
R1211 gnd.n6652 gnd.n189 585
R1212 gnd.n6624 gnd.n6623 585
R1213 gnd.n6623 gnd.n194 585
R1214 gnd.n6625 gnd.n202 585
R1215 gnd.n6639 gnd.n202 585
R1216 gnd.n6626 gnd.n214 585
R1217 gnd.n214 gnd.n212 585
R1218 gnd.n6628 gnd.n6627 585
R1219 gnd.n6629 gnd.n6628 585
R1220 gnd.n215 gnd.n213 585
R1221 gnd.n213 gnd.n209 585
R1222 gnd.n6601 gnd.n223 585
R1223 gnd.n6613 gnd.n223 585
R1224 gnd.n6602 gnd.n233 585
R1225 gnd.n233 gnd.n221 585
R1226 gnd.n6604 gnd.n6603 585
R1227 gnd.n6605 gnd.n6604 585
R1228 gnd.n234 gnd.n232 585
R1229 gnd.n6594 gnd.n232 585
R1230 gnd.n6560 gnd.n6559 585
R1231 gnd.n6559 gnd.n239 585
R1232 gnd.n6561 gnd.n248 585
R1233 gnd.n6575 gnd.n248 585
R1234 gnd.n6562 gnd.n260 585
R1235 gnd.n6553 gnd.n260 585
R1236 gnd.n6564 gnd.n6563 585
R1237 gnd.n6565 gnd.n6564 585
R1238 gnd.n261 gnd.n259 585
R1239 gnd.n6549 gnd.n259 585
R1240 gnd.n6325 gnd.n6324 585
R1241 gnd.n6324 gnd.n6323 585
R1242 gnd.n6326 gnd.n276 585
R1243 gnd.n6540 gnd.n276 585
R1244 gnd.n6328 gnd.n6327 585
R1245 gnd.n6329 gnd.n6328 585
R1246 gnd.n502 gnd.n398 585
R1247 gnd.n6410 gnd.n399 585
R1248 gnd.n6409 gnd.n400 585
R1249 gnd.n407 gnd.n401 585
R1250 gnd.n6402 gnd.n408 585
R1251 gnd.n6401 gnd.n409 585
R1252 gnd.n411 gnd.n410 585
R1253 gnd.n6394 gnd.n417 585
R1254 gnd.n6393 gnd.n418 585
R1255 gnd.n425 gnd.n419 585
R1256 gnd.n6386 gnd.n426 585
R1257 gnd.n6385 gnd.n427 585
R1258 gnd.n429 gnd.n428 585
R1259 gnd.n6378 gnd.n435 585
R1260 gnd.n6377 gnd.n436 585
R1261 gnd.n445 gnd.n437 585
R1262 gnd.n6370 gnd.n446 585
R1263 gnd.n6369 gnd.n6366 585
R1264 gnd.n447 gnd.n322 585
R1265 gnd.n6530 gnd.n322 585
R1266 gnd.n6835 gnd.n6834 585
R1267 gnd.n6737 gnd.n6733 585
R1268 gnd.n6785 gnd.n6784 585
R1269 gnd.n6783 gnd.n6782 585
R1270 gnd.n6781 gnd.n6780 585
R1271 gnd.n6774 gnd.n6739 585
R1272 gnd.n6776 gnd.n6775 585
R1273 gnd.n6773 gnd.n6772 585
R1274 gnd.n6771 gnd.n6770 585
R1275 gnd.n6764 gnd.n6741 585
R1276 gnd.n6766 gnd.n6765 585
R1277 gnd.n6763 gnd.n6762 585
R1278 gnd.n6761 gnd.n6760 585
R1279 gnd.n6754 gnd.n6743 585
R1280 gnd.n6756 gnd.n6755 585
R1281 gnd.n6753 gnd.n6752 585
R1282 gnd.n6751 gnd.n6750 585
R1283 gnd.n6747 gnd.n6746 585
R1284 gnd.n6745 gnd.n6724 585
R1285 gnd.n7042 gnd.n6724 585
R1286 gnd.n6831 gnd.n6734 585
R1287 gnd.n6734 gnd.n164 585
R1288 gnd.n6830 gnd.n163 585
R1289 gnd.n7053 gnd.n163 585
R1290 gnd.n6829 gnd.n6828 585
R1291 gnd.n6828 gnd.n154 585
R1292 gnd.n6789 gnd.n153 585
R1293 gnd.n7059 gnd.n153 585
R1294 gnd.n6824 gnd.n6823 585
R1295 gnd.n6823 gnd.n145 585
R1296 gnd.n6822 gnd.n144 585
R1297 gnd.n7065 gnd.n144 585
R1298 gnd.n6821 gnd.n6820 585
R1299 gnd.n6820 gnd.n142 585
R1300 gnd.n6791 gnd.n134 585
R1301 gnd.n7071 gnd.n134 585
R1302 gnd.n6816 gnd.n6815 585
R1303 gnd.n6815 gnd.n126 585
R1304 gnd.n6814 gnd.n125 585
R1305 gnd.n7077 gnd.n125 585
R1306 gnd.n6813 gnd.n6812 585
R1307 gnd.n6812 gnd.n116 585
R1308 gnd.n6793 gnd.n115 585
R1309 gnd.n7083 gnd.n115 585
R1310 gnd.n6808 gnd.n6807 585
R1311 gnd.n6807 gnd.n107 585
R1312 gnd.n6806 gnd.n106 585
R1313 gnd.n7089 gnd.n106 585
R1314 gnd.n6805 gnd.n6804 585
R1315 gnd.n6804 gnd.n104 585
R1316 gnd.n6795 gnd.n96 585
R1317 gnd.n7095 gnd.n96 585
R1318 gnd.n6800 gnd.n6799 585
R1319 gnd.n6799 gnd.n86 585
R1320 gnd.n6798 gnd.n85 585
R1321 gnd.n7101 gnd.n85 585
R1322 gnd.n72 gnd.n71 585
R1323 gnd.n74 gnd.n72 585
R1324 gnd.n7109 gnd.n7108 585
R1325 gnd.n7108 gnd.n7107 585
R1326 gnd.n7110 gnd.n70 585
R1327 gnd.n6680 gnd.n70 585
R1328 gnd.n178 gnd.n68 585
R1329 gnd.n178 gnd.n171 585
R1330 gnd.n6645 gnd.n179 585
R1331 gnd.n6672 gnd.n179 585
R1332 gnd.n6646 gnd.n6644 585
R1333 gnd.n6644 gnd.n188 585
R1334 gnd.n197 gnd.n187 585
R1335 gnd.n6661 gnd.n187 585
R1336 gnd.n6651 gnd.n6650 585
R1337 gnd.n6652 gnd.n6651 585
R1338 gnd.n196 gnd.n195 585
R1339 gnd.n195 gnd.n194 585
R1340 gnd.n6641 gnd.n6640 585
R1341 gnd.n6640 gnd.n6639 585
R1342 gnd.n200 gnd.n199 585
R1343 gnd.n212 gnd.n200 585
R1344 gnd.n6583 gnd.n211 585
R1345 gnd.n6629 gnd.n211 585
R1346 gnd.n6586 gnd.n6582 585
R1347 gnd.n6582 gnd.n209 585
R1348 gnd.n6587 gnd.n222 585
R1349 gnd.n6613 gnd.n222 585
R1350 gnd.n6588 gnd.n6581 585
R1351 gnd.n6581 gnd.n221 585
R1352 gnd.n242 gnd.n231 585
R1353 gnd.n6605 gnd.n231 585
R1354 gnd.n6593 gnd.n6592 585
R1355 gnd.n6594 gnd.n6593 585
R1356 gnd.n241 gnd.n240 585
R1357 gnd.n240 gnd.n239 585
R1358 gnd.n6577 gnd.n6576 585
R1359 gnd.n6576 gnd.n6575 585
R1360 gnd.n245 gnd.n244 585
R1361 gnd.n6553 gnd.n245 585
R1362 gnd.n270 gnd.n257 585
R1363 gnd.n6565 gnd.n257 585
R1364 gnd.n6548 gnd.n6547 585
R1365 gnd.n6549 gnd.n6548 585
R1366 gnd.n269 gnd.n268 585
R1367 gnd.n6323 gnd.n268 585
R1368 gnd.n6542 gnd.n6541 585
R1369 gnd.n6541 gnd.n6540 585
R1370 gnd.n273 gnd.n272 585
R1371 gnd.n6329 gnd.n273 585
R1372 gnd.n5499 gnd.n4166 585
R1373 gnd.n4166 gnd.n1008 585
R1374 gnd.n5500 gnd.n4227 585
R1375 gnd.n4227 gnd.n4217 585
R1376 gnd.n5502 gnd.n5501 585
R1377 gnd.n5503 gnd.n5502 585
R1378 gnd.n4228 gnd.n4226 585
R1379 gnd.n4235 gnd.n4226 585
R1380 gnd.n5493 gnd.n5492 585
R1381 gnd.n5492 gnd.n5491 585
R1382 gnd.n4231 gnd.n4230 585
R1383 gnd.n5218 gnd.n4231 585
R1384 gnd.n5204 gnd.n4254 585
R1385 gnd.n4254 gnd.n4244 585
R1386 gnd.n5206 gnd.n5205 585
R1387 gnd.n5207 gnd.n5206 585
R1388 gnd.n4255 gnd.n4253 585
R1389 gnd.n4253 gnd.n4251 585
R1390 gnd.n5199 gnd.n5198 585
R1391 gnd.n5198 gnd.n5197 585
R1392 gnd.n4258 gnd.n4257 585
R1393 gnd.n4267 gnd.n4258 585
R1394 gnd.n5155 gnd.n4281 585
R1395 gnd.n4281 gnd.n4266 585
R1396 gnd.n5157 gnd.n5156 585
R1397 gnd.n5158 gnd.n5157 585
R1398 gnd.n4282 gnd.n4280 585
R1399 gnd.n4289 gnd.n4280 585
R1400 gnd.n5150 gnd.n5149 585
R1401 gnd.n5149 gnd.n5148 585
R1402 gnd.n4285 gnd.n4284 585
R1403 gnd.n5129 gnd.n4285 585
R1404 gnd.n5115 gnd.n4309 585
R1405 gnd.n4309 gnd.n4298 585
R1406 gnd.n5117 gnd.n5116 585
R1407 gnd.n5118 gnd.n5117 585
R1408 gnd.n4310 gnd.n4308 585
R1409 gnd.n4308 gnd.n4305 585
R1410 gnd.n5110 gnd.n5109 585
R1411 gnd.n5109 gnd.n5108 585
R1412 gnd.n4313 gnd.n4312 585
R1413 gnd.n4323 gnd.n4313 585
R1414 gnd.n5070 gnd.n4336 585
R1415 gnd.n4336 gnd.n4322 585
R1416 gnd.n5072 gnd.n5071 585
R1417 gnd.n5073 gnd.n5072 585
R1418 gnd.n4337 gnd.n4335 585
R1419 gnd.n4344 gnd.n4335 585
R1420 gnd.n5065 gnd.n5064 585
R1421 gnd.n5064 gnd.n5063 585
R1422 gnd.n4340 gnd.n4339 585
R1423 gnd.n5044 gnd.n4340 585
R1424 gnd.n5030 gnd.n4363 585
R1425 gnd.n4363 gnd.n4353 585
R1426 gnd.n5032 gnd.n5031 585
R1427 gnd.n5033 gnd.n5032 585
R1428 gnd.n4364 gnd.n4362 585
R1429 gnd.n5021 gnd.n4362 585
R1430 gnd.n5025 gnd.n5024 585
R1431 gnd.n5024 gnd.n5023 585
R1432 gnd.n4367 gnd.n4366 585
R1433 gnd.n4976 gnd.n4367 585
R1434 gnd.n4469 gnd.n4468 585
R1435 gnd.n4470 gnd.n4469 585
R1436 gnd.n4449 gnd.n4448 585
R1437 gnd.n4452 gnd.n4449 585
R1438 gnd.n4986 gnd.n4985 585
R1439 gnd.n4985 gnd.n4984 585
R1440 gnd.n4987 gnd.n4443 585
R1441 gnd.n4479 gnd.n4443 585
R1442 gnd.n4989 gnd.n4988 585
R1443 gnd.n4990 gnd.n4989 585
R1444 gnd.n4444 gnd.n4442 585
R1445 gnd.n4954 gnd.n4442 585
R1446 gnd.n4938 gnd.n4937 585
R1447 gnd.n4937 gnd.n4430 585
R1448 gnd.n4939 gnd.n4494 585
R1449 gnd.n4494 gnd.n4429 585
R1450 gnd.n4941 gnd.n4940 585
R1451 gnd.n4942 gnd.n4941 585
R1452 gnd.n4495 gnd.n4493 585
R1453 gnd.n4493 gnd.n4490 585
R1454 gnd.n4930 gnd.n4929 585
R1455 gnd.n4929 gnd.n4928 585
R1456 gnd.n4498 gnd.n4497 585
R1457 gnd.n4505 gnd.n4498 585
R1458 gnd.n4904 gnd.n4903 585
R1459 gnd.n4905 gnd.n4904 585
R1460 gnd.n4517 gnd.n4516 585
R1461 gnd.n4524 gnd.n4516 585
R1462 gnd.n4899 gnd.n4898 585
R1463 gnd.n4898 gnd.n4897 585
R1464 gnd.n4520 gnd.n4519 585
R1465 gnd.n4887 gnd.n4520 585
R1466 gnd.n4874 gnd.n4544 585
R1467 gnd.n4544 gnd.n4543 585
R1468 gnd.n4876 gnd.n4875 585
R1469 gnd.n4877 gnd.n4876 585
R1470 gnd.n4545 gnd.n4542 585
R1471 gnd.n4552 gnd.n4542 585
R1472 gnd.n4869 gnd.n4868 585
R1473 gnd.n4868 gnd.n4867 585
R1474 gnd.n4548 gnd.n4547 585
R1475 gnd.n4856 gnd.n4548 585
R1476 gnd.n4843 gnd.n4569 585
R1477 gnd.n4569 gnd.n4568 585
R1478 gnd.n4845 gnd.n4844 585
R1479 gnd.n4846 gnd.n4845 585
R1480 gnd.n4839 gnd.n4567 585
R1481 gnd.n4838 gnd.n4837 585
R1482 gnd.n4572 gnd.n4571 585
R1483 gnd.n4835 gnd.n4572 585
R1484 gnd.n4594 gnd.n4593 585
R1485 gnd.n4597 gnd.n4596 585
R1486 gnd.n4595 gnd.n4590 585
R1487 gnd.n4602 gnd.n4601 585
R1488 gnd.n4604 gnd.n4603 585
R1489 gnd.n4607 gnd.n4606 585
R1490 gnd.n4605 gnd.n4588 585
R1491 gnd.n4612 gnd.n4611 585
R1492 gnd.n4614 gnd.n4613 585
R1493 gnd.n4617 gnd.n4616 585
R1494 gnd.n4615 gnd.n4586 585
R1495 gnd.n4622 gnd.n4621 585
R1496 gnd.n4626 gnd.n4623 585
R1497 gnd.n4627 gnd.n4564 585
R1498 gnd.n5505 gnd.n4181 585
R1499 gnd.n5572 gnd.n5571 585
R1500 gnd.n5574 gnd.n5573 585
R1501 gnd.n5576 gnd.n5575 585
R1502 gnd.n5578 gnd.n5577 585
R1503 gnd.n5580 gnd.n5579 585
R1504 gnd.n5582 gnd.n5581 585
R1505 gnd.n5584 gnd.n5583 585
R1506 gnd.n5586 gnd.n5585 585
R1507 gnd.n5588 gnd.n5587 585
R1508 gnd.n5590 gnd.n5589 585
R1509 gnd.n5592 gnd.n5591 585
R1510 gnd.n5594 gnd.n5593 585
R1511 gnd.n5597 gnd.n5596 585
R1512 gnd.n5595 gnd.n4169 585
R1513 gnd.n5601 gnd.n4167 585
R1514 gnd.n5603 gnd.n5602 585
R1515 gnd.n5604 gnd.n5603 585
R1516 gnd.n5506 gnd.n4222 585
R1517 gnd.n5506 gnd.n1008 585
R1518 gnd.n5508 gnd.n5507 585
R1519 gnd.n5507 gnd.n4217 585
R1520 gnd.n5504 gnd.n4221 585
R1521 gnd.n5504 gnd.n5503 585
R1522 gnd.n5483 gnd.n4223 585
R1523 gnd.n4235 gnd.n4223 585
R1524 gnd.n5482 gnd.n4233 585
R1525 gnd.n5491 gnd.n4233 585
R1526 gnd.n5217 gnd.n4240 585
R1527 gnd.n5218 gnd.n5217 585
R1528 gnd.n5216 gnd.n5215 585
R1529 gnd.n5216 gnd.n4244 585
R1530 gnd.n5214 gnd.n4246 585
R1531 gnd.n5207 gnd.n4246 585
R1532 gnd.n4259 gnd.n4247 585
R1533 gnd.n4259 gnd.n4251 585
R1534 gnd.n5163 gnd.n4260 585
R1535 gnd.n5197 gnd.n4260 585
R1536 gnd.n5162 gnd.n5161 585
R1537 gnd.n5161 gnd.n4267 585
R1538 gnd.n5160 gnd.n4275 585
R1539 gnd.n5160 gnd.n4266 585
R1540 gnd.n5159 gnd.n4277 585
R1541 gnd.n5159 gnd.n5158 585
R1542 gnd.n5138 gnd.n4276 585
R1543 gnd.n4289 gnd.n4276 585
R1544 gnd.n5137 gnd.n4287 585
R1545 gnd.n5148 gnd.n4287 585
R1546 gnd.n5128 gnd.n4294 585
R1547 gnd.n5129 gnd.n5128 585
R1548 gnd.n5127 gnd.n5126 585
R1549 gnd.n5127 gnd.n4298 585
R1550 gnd.n5125 gnd.n4300 585
R1551 gnd.n5118 gnd.n4300 585
R1552 gnd.n4315 gnd.n4301 585
R1553 gnd.n4315 gnd.n4305 585
R1554 gnd.n5078 gnd.n4316 585
R1555 gnd.n5108 gnd.n4316 585
R1556 gnd.n5077 gnd.n5076 585
R1557 gnd.n5076 gnd.n4323 585
R1558 gnd.n5075 gnd.n4330 585
R1559 gnd.n5075 gnd.n4322 585
R1560 gnd.n5074 gnd.n4332 585
R1561 gnd.n5074 gnd.n5073 585
R1562 gnd.n5053 gnd.n4331 585
R1563 gnd.n4344 gnd.n4331 585
R1564 gnd.n5052 gnd.n4342 585
R1565 gnd.n5063 gnd.n4342 585
R1566 gnd.n5043 gnd.n4349 585
R1567 gnd.n5044 gnd.n5043 585
R1568 gnd.n5042 gnd.n5041 585
R1569 gnd.n5042 gnd.n4353 585
R1570 gnd.n5040 gnd.n4355 585
R1571 gnd.n5033 gnd.n4355 585
R1572 gnd.n5020 gnd.n4356 585
R1573 gnd.n5021 gnd.n5020 585
R1574 gnd.n4973 gnd.n4369 585
R1575 gnd.n5023 gnd.n4369 585
R1576 gnd.n4975 gnd.n4974 585
R1577 gnd.n4976 gnd.n4975 585
R1578 gnd.n4968 gnd.n4471 585
R1579 gnd.n4471 gnd.n4470 585
R1580 gnd.n4966 gnd.n4965 585
R1581 gnd.n4965 gnd.n4452 585
R1582 gnd.n4963 gnd.n4450 585
R1583 gnd.n4984 gnd.n4450 585
R1584 gnd.n4481 gnd.n4480 585
R1585 gnd.n4480 gnd.n4479 585
R1586 gnd.n4957 gnd.n4440 585
R1587 gnd.n4990 gnd.n4440 585
R1588 gnd.n4956 gnd.n4955 585
R1589 gnd.n4955 gnd.n4954 585
R1590 gnd.n4952 gnd.n4483 585
R1591 gnd.n4952 gnd.n4430 585
R1592 gnd.n4951 gnd.n4950 585
R1593 gnd.n4951 gnd.n4429 585
R1594 gnd.n4486 gnd.n4485 585
R1595 gnd.n4942 gnd.n4485 585
R1596 gnd.n4910 gnd.n4909 585
R1597 gnd.n4909 gnd.n4490 585
R1598 gnd.n4911 gnd.n4499 585
R1599 gnd.n4928 gnd.n4499 585
R1600 gnd.n4908 gnd.n4907 585
R1601 gnd.n4907 gnd.n4505 585
R1602 gnd.n4906 gnd.n4513 585
R1603 gnd.n4906 gnd.n4905 585
R1604 gnd.n4891 gnd.n4514 585
R1605 gnd.n4524 gnd.n4514 585
R1606 gnd.n4890 gnd.n4522 585
R1607 gnd.n4897 gnd.n4522 585
R1608 gnd.n4889 gnd.n4888 585
R1609 gnd.n4888 gnd.n4887 585
R1610 gnd.n4533 gnd.n4530 585
R1611 gnd.n4543 gnd.n4533 585
R1612 gnd.n4879 gnd.n4878 585
R1613 gnd.n4878 gnd.n4877 585
R1614 gnd.n4539 gnd.n4538 585
R1615 gnd.n4552 gnd.n4539 585
R1616 gnd.n4859 gnd.n4550 585
R1617 gnd.n4867 gnd.n4550 585
R1618 gnd.n4858 gnd.n4857 585
R1619 gnd.n4857 gnd.n4856 585
R1620 gnd.n4559 gnd.n4557 585
R1621 gnd.n4568 gnd.n4559 585
R1622 gnd.n4848 gnd.n4847 585
R1623 gnd.n4847 gnd.n4846 585
R1624 gnd.n3542 gnd.n3541 585
R1625 gnd.n3543 gnd.n3542 585
R1626 gnd.n1649 gnd.n1647 585
R1627 gnd.n3417 gnd.n1647 585
R1628 gnd.n3389 gnd.n3386 585
R1629 gnd.n3389 gnd.n3388 585
R1630 gnd.n3390 gnd.n3385 585
R1631 gnd.n3390 gnd.t266 585
R1632 gnd.n3392 gnd.n3391 585
R1633 gnd.n3391 gnd.n1731 585
R1634 gnd.n3393 gnd.n1741 585
R1635 gnd.n3373 gnd.n1741 585
R1636 gnd.n3395 gnd.n3394 585
R1637 gnd.n3396 gnd.n3395 585
R1638 gnd.n3384 gnd.n1740 585
R1639 gnd.n3379 gnd.n1740 585
R1640 gnd.n3383 gnd.n3382 585
R1641 gnd.n3382 gnd.n3381 585
R1642 gnd.n1743 gnd.n1742 585
R1643 gnd.n3364 gnd.n1743 585
R1644 gnd.n3350 gnd.n3349 585
R1645 gnd.n3349 gnd.n3348 585
R1646 gnd.n3351 gnd.n1756 585
R1647 gnd.n3327 gnd.n1756 585
R1648 gnd.n3353 gnd.n3352 585
R1649 gnd.n3354 gnd.n3353 585
R1650 gnd.n1757 gnd.n1755 585
R1651 gnd.n3333 gnd.n1755 585
R1652 gnd.n3307 gnd.n3306 585
R1653 gnd.n3306 gnd.n3305 585
R1654 gnd.n3308 gnd.n1769 585
R1655 gnd.n3322 gnd.n1769 585
R1656 gnd.n3309 gnd.n1781 585
R1657 gnd.n3290 gnd.n1781 585
R1658 gnd.n3311 gnd.n3310 585
R1659 gnd.n3312 gnd.n3311 585
R1660 gnd.n3304 gnd.n1780 585
R1661 gnd.n1780 gnd.n1776 585
R1662 gnd.n3303 gnd.n3302 585
R1663 gnd.n3302 gnd.n3301 585
R1664 gnd.n1783 gnd.n1782 585
R1665 gnd.n3200 gnd.n1783 585
R1666 gnd.n3283 gnd.n3282 585
R1667 gnd.n3284 gnd.n3283 585
R1668 gnd.n3281 gnd.n1795 585
R1669 gnd.n1795 gnd.n1792 585
R1670 gnd.n3280 gnd.n3279 585
R1671 gnd.n3279 gnd.n3278 585
R1672 gnd.n1797 gnd.n1796 585
R1673 gnd.n3211 gnd.n1797 585
R1674 gnd.n3265 gnd.n3264 585
R1675 gnd.n3266 gnd.n3265 585
R1676 gnd.n3263 gnd.n1807 585
R1677 gnd.n1807 gnd.n1805 585
R1678 gnd.n3262 gnd.n3261 585
R1679 gnd.n3261 gnd.n3260 585
R1680 gnd.n1809 gnd.n1808 585
R1681 gnd.n1820 gnd.n1809 585
R1682 gnd.n3235 gnd.n3234 585
R1683 gnd.n3234 gnd.n1818 585
R1684 gnd.n3236 gnd.n1831 585
R1685 gnd.n3222 gnd.n1831 585
R1686 gnd.n3238 gnd.n3237 585
R1687 gnd.n3239 gnd.n3238 585
R1688 gnd.n3233 gnd.n1830 585
R1689 gnd.n3228 gnd.n1830 585
R1690 gnd.n3232 gnd.n3231 585
R1691 gnd.n3231 gnd.n3230 585
R1692 gnd.n1833 gnd.n1832 585
R1693 gnd.n3190 gnd.n1833 585
R1694 gnd.n3176 gnd.n3175 585
R1695 gnd.n3175 gnd.n3174 585
R1696 gnd.n3177 gnd.n1845 585
R1697 gnd.n3154 gnd.n1845 585
R1698 gnd.n3179 gnd.n3178 585
R1699 gnd.n3180 gnd.n3179 585
R1700 gnd.n1846 gnd.n1844 585
R1701 gnd.n3160 gnd.n1844 585
R1702 gnd.n3132 gnd.n3131 585
R1703 gnd.n3131 gnd.n3130 585
R1704 gnd.n3133 gnd.n1860 585
R1705 gnd.n3148 gnd.n1860 585
R1706 gnd.n3134 gnd.n1873 585
R1707 gnd.n1873 gnd.n1872 585
R1708 gnd.n3136 gnd.n3135 585
R1709 gnd.n3137 gnd.n3136 585
R1710 gnd.n3129 gnd.n1871 585
R1711 gnd.n1871 gnd.n1867 585
R1712 gnd.n3128 gnd.n3127 585
R1713 gnd.n3127 gnd.n3126 585
R1714 gnd.n1875 gnd.n1874 585
R1715 gnd.n3030 gnd.n1875 585
R1716 gnd.n3111 gnd.n3110 585
R1717 gnd.n3112 gnd.n3111 585
R1718 gnd.n3109 gnd.n1887 585
R1719 gnd.n1887 gnd.n1884 585
R1720 gnd.n3108 gnd.n3107 585
R1721 gnd.n3107 gnd.n3106 585
R1722 gnd.n1889 gnd.n1888 585
R1723 gnd.n3038 gnd.n1889 585
R1724 gnd.n3093 gnd.n3092 585
R1725 gnd.n3094 gnd.n3093 585
R1726 gnd.n3091 gnd.n1902 585
R1727 gnd.n1902 gnd.n1899 585
R1728 gnd.n3090 gnd.n3089 585
R1729 gnd.n3089 gnd.n3088 585
R1730 gnd.n1904 gnd.n1903 585
R1731 gnd.n1915 gnd.n1904 585
R1732 gnd.n3062 gnd.n3061 585
R1733 gnd.n3061 gnd.n1914 585
R1734 gnd.n3063 gnd.n1925 585
R1735 gnd.n3049 gnd.n1925 585
R1736 gnd.n3065 gnd.n3064 585
R1737 gnd.n3066 gnd.n3065 585
R1738 gnd.n3060 gnd.n1924 585
R1739 gnd.n3055 gnd.n1924 585
R1740 gnd.n3059 gnd.n3058 585
R1741 gnd.n3058 gnd.n3057 585
R1742 gnd.n1927 gnd.n1926 585
R1743 gnd.n3020 gnd.n1927 585
R1744 gnd.n3006 gnd.n3005 585
R1745 gnd.n3005 gnd.n3004 585
R1746 gnd.n3007 gnd.n1942 585
R1747 gnd.n3002 gnd.n1942 585
R1748 gnd.n3009 gnd.n3008 585
R1749 gnd.n3010 gnd.n3009 585
R1750 gnd.n1943 gnd.n1941 585
R1751 gnd.n2996 gnd.n1941 585
R1752 gnd.n2960 gnd.n2959 585
R1753 gnd.n2959 gnd.n2958 585
R1754 gnd.n2961 gnd.n1955 585
R1755 gnd.n2975 gnd.n1955 585
R1756 gnd.n2962 gnd.n1966 585
R1757 gnd.n1966 gnd.n1954 585
R1758 gnd.n2964 gnd.n2963 585
R1759 gnd.n2965 gnd.n2964 585
R1760 gnd.n2956 gnd.n1965 585
R1761 gnd.n1965 gnd.n1962 585
R1762 gnd.n2955 gnd.n2954 585
R1763 gnd.n2954 gnd.n2953 585
R1764 gnd.n1968 gnd.n1967 585
R1765 gnd.n2901 gnd.n1968 585
R1766 gnd.n2941 gnd.n2940 585
R1767 gnd.n2942 gnd.n2941 585
R1768 gnd.n2939 gnd.n1979 585
R1769 gnd.n1979 gnd.n1976 585
R1770 gnd.n2938 gnd.n2937 585
R1771 gnd.n2937 gnd.n2936 585
R1772 gnd.n1981 gnd.n1980 585
R1773 gnd.n2909 gnd.n1981 585
R1774 gnd.n2923 gnd.n2922 585
R1775 gnd.n2924 gnd.n2923 585
R1776 gnd.n2921 gnd.n1992 585
R1777 gnd.n2915 gnd.n1992 585
R1778 gnd.n2920 gnd.n2919 585
R1779 gnd.n2919 gnd.n2918 585
R1780 gnd.n1470 gnd.n1469 585
R1781 gnd.n2889 gnd.n1470 585
R1782 gnd.n3781 gnd.n3780 585
R1783 gnd.n3780 gnd.n3779 585
R1784 gnd.n3782 gnd.n1448 585
R1785 gnd.n2875 gnd.n1448 585
R1786 gnd.n3847 gnd.n3846 585
R1787 gnd.n3845 gnd.n1447 585
R1788 gnd.n3844 gnd.n1446 585
R1789 gnd.n3849 gnd.n1446 585
R1790 gnd.n3843 gnd.n3842 585
R1791 gnd.n3841 gnd.n3840 585
R1792 gnd.n3839 gnd.n3838 585
R1793 gnd.n3837 gnd.n3836 585
R1794 gnd.n3835 gnd.n3834 585
R1795 gnd.n3833 gnd.n3832 585
R1796 gnd.n3831 gnd.n3830 585
R1797 gnd.n3829 gnd.n3828 585
R1798 gnd.n3827 gnd.n3826 585
R1799 gnd.n3825 gnd.n3824 585
R1800 gnd.n3823 gnd.n3822 585
R1801 gnd.n3821 gnd.n3820 585
R1802 gnd.n3819 gnd.n3818 585
R1803 gnd.n3817 gnd.n3816 585
R1804 gnd.n3815 gnd.n3814 585
R1805 gnd.n3813 gnd.n3812 585
R1806 gnd.n3811 gnd.n3810 585
R1807 gnd.n3809 gnd.n3808 585
R1808 gnd.n3807 gnd.n3806 585
R1809 gnd.n3805 gnd.n3804 585
R1810 gnd.n3803 gnd.n3802 585
R1811 gnd.n3801 gnd.n3800 585
R1812 gnd.n3799 gnd.n3798 585
R1813 gnd.n3797 gnd.n3796 585
R1814 gnd.n3795 gnd.n3794 585
R1815 gnd.n3793 gnd.n3792 585
R1816 gnd.n3791 gnd.n3790 585
R1817 gnd.n3789 gnd.n3788 585
R1818 gnd.n3787 gnd.n1410 585
R1819 gnd.n3852 gnd.n3851 585
R1820 gnd.n1412 gnd.n1409 585
R1821 gnd.n2812 gnd.n2811 585
R1822 gnd.n2814 gnd.n2813 585
R1823 gnd.n2817 gnd.n2816 585
R1824 gnd.n2819 gnd.n2818 585
R1825 gnd.n2821 gnd.n2820 585
R1826 gnd.n2823 gnd.n2822 585
R1827 gnd.n2825 gnd.n2824 585
R1828 gnd.n2827 gnd.n2826 585
R1829 gnd.n2829 gnd.n2828 585
R1830 gnd.n2831 gnd.n2830 585
R1831 gnd.n2833 gnd.n2832 585
R1832 gnd.n2835 gnd.n2834 585
R1833 gnd.n2837 gnd.n2836 585
R1834 gnd.n2839 gnd.n2838 585
R1835 gnd.n2841 gnd.n2840 585
R1836 gnd.n2843 gnd.n2842 585
R1837 gnd.n2845 gnd.n2844 585
R1838 gnd.n2847 gnd.n2846 585
R1839 gnd.n2849 gnd.n2848 585
R1840 gnd.n2851 gnd.n2850 585
R1841 gnd.n2853 gnd.n2852 585
R1842 gnd.n2855 gnd.n2854 585
R1843 gnd.n2857 gnd.n2856 585
R1844 gnd.n2859 gnd.n2858 585
R1845 gnd.n2861 gnd.n2860 585
R1846 gnd.n2863 gnd.n2862 585
R1847 gnd.n2865 gnd.n2864 585
R1848 gnd.n2867 gnd.n2866 585
R1849 gnd.n2869 gnd.n2868 585
R1850 gnd.n2871 gnd.n2870 585
R1851 gnd.n2872 gnd.n2808 585
R1852 gnd.n3423 gnd.n3422 585
R1853 gnd.n3424 gnd.n1720 585
R1854 gnd.n3426 gnd.n3425 585
R1855 gnd.n3428 gnd.n1718 585
R1856 gnd.n3430 gnd.n3429 585
R1857 gnd.n3431 gnd.n1717 585
R1858 gnd.n3433 gnd.n3432 585
R1859 gnd.n3435 gnd.n1715 585
R1860 gnd.n3437 gnd.n3436 585
R1861 gnd.n3438 gnd.n1714 585
R1862 gnd.n3440 gnd.n3439 585
R1863 gnd.n3442 gnd.n1712 585
R1864 gnd.n3444 gnd.n3443 585
R1865 gnd.n3445 gnd.n1711 585
R1866 gnd.n3447 gnd.n3446 585
R1867 gnd.n3449 gnd.n1709 585
R1868 gnd.n3451 gnd.n3450 585
R1869 gnd.n3452 gnd.n1708 585
R1870 gnd.n3454 gnd.n3453 585
R1871 gnd.n3456 gnd.n1706 585
R1872 gnd.n3458 gnd.n3457 585
R1873 gnd.n3459 gnd.n1705 585
R1874 gnd.n3461 gnd.n3460 585
R1875 gnd.n3463 gnd.n1703 585
R1876 gnd.n3465 gnd.n3464 585
R1877 gnd.n3466 gnd.n1702 585
R1878 gnd.n3468 gnd.n3467 585
R1879 gnd.n3470 gnd.n1700 585
R1880 gnd.n3472 gnd.n3471 585
R1881 gnd.n3474 gnd.n1697 585
R1882 gnd.n3476 gnd.n3475 585
R1883 gnd.n3478 gnd.n1696 585
R1884 gnd.n3479 gnd.n1672 585
R1885 gnd.n3482 gnd.n351 585
R1886 gnd.n3484 gnd.n3483 585
R1887 gnd.n3486 gnd.n1694 585
R1888 gnd.n3488 gnd.n3487 585
R1889 gnd.n3490 gnd.n1691 585
R1890 gnd.n3492 gnd.n3491 585
R1891 gnd.n3494 gnd.n1689 585
R1892 gnd.n3496 gnd.n3495 585
R1893 gnd.n3497 gnd.n1688 585
R1894 gnd.n3499 gnd.n3498 585
R1895 gnd.n3501 gnd.n1686 585
R1896 gnd.n3503 gnd.n3502 585
R1897 gnd.n3504 gnd.n1685 585
R1898 gnd.n3506 gnd.n3505 585
R1899 gnd.n3508 gnd.n1683 585
R1900 gnd.n3510 gnd.n3509 585
R1901 gnd.n3511 gnd.n1682 585
R1902 gnd.n3513 gnd.n3512 585
R1903 gnd.n3515 gnd.n1680 585
R1904 gnd.n3517 gnd.n3516 585
R1905 gnd.n3518 gnd.n1679 585
R1906 gnd.n3520 gnd.n3519 585
R1907 gnd.n3522 gnd.n1677 585
R1908 gnd.n3524 gnd.n3523 585
R1909 gnd.n3525 gnd.n1676 585
R1910 gnd.n3527 gnd.n3526 585
R1911 gnd.n3529 gnd.n1674 585
R1912 gnd.n3531 gnd.n3530 585
R1913 gnd.n3532 gnd.n1673 585
R1914 gnd.n3534 gnd.n3533 585
R1915 gnd.n3536 gnd.n1669 585
R1916 gnd.n3538 gnd.n3537 585
R1917 gnd.n3539 gnd.n1648 585
R1918 gnd.n3420 gnd.n1645 585
R1919 gnd.n3543 gnd.n1645 585
R1920 gnd.n3419 gnd.n3418 585
R1921 gnd.n3418 gnd.n3417 585
R1922 gnd.n1722 gnd.n1721 585
R1923 gnd.n3388 gnd.n1722 585
R1924 gnd.n3370 gnd.n3369 585
R1925 gnd.n3370 gnd.t266 585
R1926 gnd.n3371 gnd.n3368 585
R1927 gnd.n3371 gnd.n1731 585
R1928 gnd.n3375 gnd.n3374 585
R1929 gnd.n3374 gnd.n3373 585
R1930 gnd.n3376 gnd.n1739 585
R1931 gnd.n3396 gnd.n1739 585
R1932 gnd.n3378 gnd.n3377 585
R1933 gnd.n3379 gnd.n3378 585
R1934 gnd.n3367 gnd.n1745 585
R1935 gnd.n3381 gnd.n1745 585
R1936 gnd.n3366 gnd.n3365 585
R1937 gnd.n3365 gnd.n3364 585
R1938 gnd.n1747 gnd.n1746 585
R1939 gnd.n3348 gnd.n1747 585
R1940 gnd.n3329 gnd.n3328 585
R1941 gnd.n3328 gnd.n3327 585
R1942 gnd.n3330 gnd.n1753 585
R1943 gnd.n3354 gnd.n1753 585
R1944 gnd.n3332 gnd.n3331 585
R1945 gnd.n3333 gnd.n3332 585
R1946 gnd.n3325 gnd.n1766 585
R1947 gnd.n3305 gnd.n1766 585
R1948 gnd.n3324 gnd.n3323 585
R1949 gnd.n3323 gnd.n3322 585
R1950 gnd.n1768 gnd.n1767 585
R1951 gnd.n3290 gnd.n1768 585
R1952 gnd.n3195 gnd.n1778 585
R1953 gnd.n3312 gnd.n1778 585
R1954 gnd.n3197 gnd.n3196 585
R1955 gnd.n3196 gnd.n1776 585
R1956 gnd.n3198 gnd.n1785 585
R1957 gnd.n3301 gnd.n1785 585
R1958 gnd.n3202 gnd.n3201 585
R1959 gnd.n3201 gnd.n3200 585
R1960 gnd.n3203 gnd.n1793 585
R1961 gnd.n3284 gnd.n1793 585
R1962 gnd.n3205 gnd.n3204 585
R1963 gnd.n3204 gnd.n1792 585
R1964 gnd.n3206 gnd.n1798 585
R1965 gnd.n3278 gnd.n1798 585
R1966 gnd.n3213 gnd.n3212 585
R1967 gnd.n3212 gnd.n3211 585
R1968 gnd.n3214 gnd.n1806 585
R1969 gnd.n3266 gnd.n1806 585
R1970 gnd.n3216 gnd.n3215 585
R1971 gnd.n3215 gnd.n1805 585
R1972 gnd.n3217 gnd.n1810 585
R1973 gnd.n3260 gnd.n1810 585
R1974 gnd.n3219 gnd.n3218 585
R1975 gnd.n3219 gnd.n1820 585
R1976 gnd.n3220 gnd.n3194 585
R1977 gnd.n3220 gnd.n1818 585
R1978 gnd.n3224 gnd.n3223 585
R1979 gnd.n3223 gnd.n3222 585
R1980 gnd.n3225 gnd.n1827 585
R1981 gnd.n3239 gnd.n1827 585
R1982 gnd.n3227 gnd.n3226 585
R1983 gnd.n3228 gnd.n3227 585
R1984 gnd.n3193 gnd.n1835 585
R1985 gnd.n3230 gnd.n1835 585
R1986 gnd.n3192 gnd.n3191 585
R1987 gnd.n3191 gnd.n3190 585
R1988 gnd.n1837 gnd.n1836 585
R1989 gnd.n3174 gnd.n1837 585
R1990 gnd.n3156 gnd.n3155 585
R1991 gnd.n3155 gnd.n3154 585
R1992 gnd.n3157 gnd.n1843 585
R1993 gnd.n3180 gnd.n1843 585
R1994 gnd.n3159 gnd.n3158 585
R1995 gnd.n3160 gnd.n3159 585
R1996 gnd.n3151 gnd.n1856 585
R1997 gnd.n3130 gnd.n1856 585
R1998 gnd.n3150 gnd.n3149 585
R1999 gnd.n3149 gnd.n3148 585
R2000 gnd.n1858 gnd.n1857 585
R2001 gnd.n1872 gnd.n1858 585
R2002 gnd.n3025 gnd.n1869 585
R2003 gnd.n3137 gnd.n1869 585
R2004 gnd.n3027 gnd.n3026 585
R2005 gnd.n3026 gnd.n1867 585
R2006 gnd.n3028 gnd.n1877 585
R2007 gnd.n3126 gnd.n1877 585
R2008 gnd.n3032 gnd.n3031 585
R2009 gnd.n3031 gnd.n3030 585
R2010 gnd.n3033 gnd.n1885 585
R2011 gnd.n3112 gnd.n1885 585
R2012 gnd.n3035 gnd.n3034 585
R2013 gnd.n3034 gnd.n1884 585
R2014 gnd.n3036 gnd.n1892 585
R2015 gnd.n3106 gnd.n1892 585
R2016 gnd.n3040 gnd.n3039 585
R2017 gnd.n3039 gnd.n3038 585
R2018 gnd.n3041 gnd.n1900 585
R2019 gnd.n3094 gnd.n1900 585
R2020 gnd.n3043 gnd.n3042 585
R2021 gnd.n3042 gnd.n1899 585
R2022 gnd.n3044 gnd.n1906 585
R2023 gnd.n3088 gnd.n1906 585
R2024 gnd.n3046 gnd.n3045 585
R2025 gnd.n3046 gnd.n1915 585
R2026 gnd.n3047 gnd.n3024 585
R2027 gnd.n3047 gnd.n1914 585
R2028 gnd.n3051 gnd.n3050 585
R2029 gnd.n3050 gnd.n3049 585
R2030 gnd.n3052 gnd.n1922 585
R2031 gnd.n3066 gnd.n1922 585
R2032 gnd.n3054 gnd.n3053 585
R2033 gnd.n3055 gnd.n3054 585
R2034 gnd.n3023 gnd.n1929 585
R2035 gnd.n3057 gnd.n1929 585
R2036 gnd.n3022 gnd.n3021 585
R2037 gnd.n3021 gnd.n3020 585
R2038 gnd.n1931 gnd.n1930 585
R2039 gnd.n3004 gnd.n1931 585
R2040 gnd.n3001 gnd.n3000 585
R2041 gnd.n3002 gnd.n3001 585
R2042 gnd.n2999 gnd.n1939 585
R2043 gnd.n3010 gnd.n1939 585
R2044 gnd.n2998 gnd.n2997 585
R2045 gnd.n2997 gnd.n2996 585
R2046 gnd.n1945 gnd.n1944 585
R2047 gnd.n2958 gnd.n1945 585
R2048 gnd.n2893 gnd.n1956 585
R2049 gnd.n2975 gnd.n1956 585
R2050 gnd.n2895 gnd.n2894 585
R2051 gnd.n2894 gnd.n1954 585
R2052 gnd.n2896 gnd.n1963 585
R2053 gnd.n2965 gnd.n1963 585
R2054 gnd.n2898 gnd.n2897 585
R2055 gnd.n2897 gnd.n1962 585
R2056 gnd.n2899 gnd.n1970 585
R2057 gnd.n2953 gnd.n1970 585
R2058 gnd.n2903 gnd.n2902 585
R2059 gnd.n2902 gnd.n2901 585
R2060 gnd.n2904 gnd.n1977 585
R2061 gnd.n2942 gnd.n1977 585
R2062 gnd.n2906 gnd.n2905 585
R2063 gnd.n2905 gnd.n1976 585
R2064 gnd.n2907 gnd.n1983 585
R2065 gnd.n2936 gnd.n1983 585
R2066 gnd.n2911 gnd.n2910 585
R2067 gnd.n2910 gnd.n2909 585
R2068 gnd.n2912 gnd.n1990 585
R2069 gnd.n2924 gnd.n1990 585
R2070 gnd.n2914 gnd.n2913 585
R2071 gnd.n2915 gnd.n2914 585
R2072 gnd.n2892 gnd.n1993 585
R2073 gnd.n2918 gnd.n1993 585
R2074 gnd.n2891 gnd.n2890 585
R2075 gnd.n2890 gnd.n2889 585
R2076 gnd.n1995 gnd.n1472 585
R2077 gnd.n3779 gnd.n1472 585
R2078 gnd.n2874 gnd.n2873 585
R2079 gnd.n2875 gnd.n2874 585
R2080 gnd.n3908 gnd.n1333 585
R2081 gnd.n2598 gnd.n1333 585
R2082 gnd.n3910 gnd.n3909 585
R2083 gnd.n3911 gnd.n3910 585
R2084 gnd.n1319 gnd.n1318 585
R2085 gnd.n2565 gnd.n1319 585
R2086 gnd.n3919 gnd.n3918 585
R2087 gnd.n3918 gnd.n3917 585
R2088 gnd.n3920 gnd.n1313 585
R2089 gnd.n2543 gnd.n1313 585
R2090 gnd.n3922 gnd.n3921 585
R2091 gnd.n3923 gnd.n3922 585
R2092 gnd.n1298 gnd.n1297 585
R2093 gnd.n2531 gnd.n1298 585
R2094 gnd.n3931 gnd.n3930 585
R2095 gnd.n3930 gnd.n3929 585
R2096 gnd.n3932 gnd.n1292 585
R2097 gnd.n1299 gnd.n1292 585
R2098 gnd.n3934 gnd.n3933 585
R2099 gnd.n3935 gnd.n3934 585
R2100 gnd.n1279 gnd.n1278 585
R2101 gnd.n1282 gnd.n1279 585
R2102 gnd.n3943 gnd.n3942 585
R2103 gnd.n3942 gnd.n3941 585
R2104 gnd.n3944 gnd.n1273 585
R2105 gnd.n1273 gnd.n1272 585
R2106 gnd.n3946 gnd.n3945 585
R2107 gnd.n3947 gnd.n3946 585
R2108 gnd.n1260 gnd.n1259 585
R2109 gnd.n1269 gnd.n1260 585
R2110 gnd.n3955 gnd.n3954 585
R2111 gnd.n3954 gnd.n3953 585
R2112 gnd.n3956 gnd.n1254 585
R2113 gnd.n1254 gnd.n1253 585
R2114 gnd.n3958 gnd.n3957 585
R2115 gnd.n3959 gnd.n3958 585
R2116 gnd.n1241 gnd.n1240 585
R2117 gnd.n1244 gnd.n1241 585
R2118 gnd.n3967 gnd.n3966 585
R2119 gnd.n3966 gnd.n3965 585
R2120 gnd.n3968 gnd.n1235 585
R2121 gnd.n1235 gnd.n1234 585
R2122 gnd.n3970 gnd.n3969 585
R2123 gnd.n3971 gnd.n3970 585
R2124 gnd.n1221 gnd.n1220 585
R2125 gnd.n1231 gnd.n1221 585
R2126 gnd.n3979 gnd.n3978 585
R2127 gnd.n3978 gnd.n3977 585
R2128 gnd.n3980 gnd.n1215 585
R2129 gnd.n1222 gnd.n1215 585
R2130 gnd.n3982 gnd.n3981 585
R2131 gnd.n3983 gnd.n3982 585
R2132 gnd.n1203 gnd.n1202 585
R2133 gnd.n1206 gnd.n1203 585
R2134 gnd.n3991 gnd.n3990 585
R2135 gnd.n3990 gnd.n3989 585
R2136 gnd.n3992 gnd.n1197 585
R2137 gnd.n1197 gnd.n1196 585
R2138 gnd.n3994 gnd.n3993 585
R2139 gnd.n3995 gnd.n3994 585
R2140 gnd.n1183 gnd.n1182 585
R2141 gnd.n1193 gnd.n1183 585
R2142 gnd.n4003 gnd.n4002 585
R2143 gnd.n4002 gnd.n4001 585
R2144 gnd.n4004 gnd.n1177 585
R2145 gnd.n1184 gnd.n1177 585
R2146 gnd.n4006 gnd.n4005 585
R2147 gnd.n4007 gnd.n4006 585
R2148 gnd.n1165 gnd.n1164 585
R2149 gnd.n1168 gnd.n1165 585
R2150 gnd.n4015 gnd.n4014 585
R2151 gnd.n4014 gnd.n4013 585
R2152 gnd.n4016 gnd.n1160 585
R2153 gnd.n1160 gnd.n1159 585
R2154 gnd.n4018 gnd.n4017 585
R2155 gnd.n4019 gnd.n4018 585
R2156 gnd.n1145 gnd.n1144 585
R2157 gnd.n1149 gnd.n1145 585
R2158 gnd.n4027 gnd.n4026 585
R2159 gnd.n4026 gnd.n4025 585
R2160 gnd.n1141 gnd.n1139 585
R2161 gnd.n1146 gnd.n1139 585
R2162 gnd.n4032 gnd.n4031 585
R2163 gnd.n4033 gnd.n4032 585
R2164 gnd.n1140 gnd.n1064 585
R2165 gnd.n1064 gnd.n1061 585
R2166 gnd.n4155 gnd.n4154 585
R2167 gnd.n4153 gnd.n1063 585
R2168 gnd.n4152 gnd.n1062 585
R2169 gnd.n4157 gnd.n1062 585
R2170 gnd.n4151 gnd.n4150 585
R2171 gnd.n4149 gnd.n4148 585
R2172 gnd.n4147 gnd.n4146 585
R2173 gnd.n4145 gnd.n4144 585
R2174 gnd.n4143 gnd.n4142 585
R2175 gnd.n4141 gnd.n4140 585
R2176 gnd.n4139 gnd.n4138 585
R2177 gnd.n4137 gnd.n4136 585
R2178 gnd.n4135 gnd.n4134 585
R2179 gnd.n4133 gnd.n4132 585
R2180 gnd.n4131 gnd.n4130 585
R2181 gnd.n4129 gnd.n4128 585
R2182 gnd.n4127 gnd.n4126 585
R2183 gnd.n4125 gnd.n4124 585
R2184 gnd.n4123 gnd.n4122 585
R2185 gnd.n4120 gnd.n4119 585
R2186 gnd.n4118 gnd.n4117 585
R2187 gnd.n4116 gnd.n4115 585
R2188 gnd.n4114 gnd.n4113 585
R2189 gnd.n4112 gnd.n4111 585
R2190 gnd.n4110 gnd.n4109 585
R2191 gnd.n4108 gnd.n4107 585
R2192 gnd.n4106 gnd.n4105 585
R2193 gnd.n4104 gnd.n4103 585
R2194 gnd.n4102 gnd.n4101 585
R2195 gnd.n4100 gnd.n4099 585
R2196 gnd.n4098 gnd.n4097 585
R2197 gnd.n4096 gnd.n4095 585
R2198 gnd.n4094 gnd.n4093 585
R2199 gnd.n4092 gnd.n4091 585
R2200 gnd.n4090 gnd.n4089 585
R2201 gnd.n4088 gnd.n4087 585
R2202 gnd.n4086 gnd.n4085 585
R2203 gnd.n4084 gnd.n4083 585
R2204 gnd.n4082 gnd.n4081 585
R2205 gnd.n4080 gnd.n4079 585
R2206 gnd.n4078 gnd.n4077 585
R2207 gnd.n4076 gnd.n4075 585
R2208 gnd.n4074 gnd.n4073 585
R2209 gnd.n4072 gnd.n4071 585
R2210 gnd.n4070 gnd.n4069 585
R2211 gnd.n4068 gnd.n4067 585
R2212 gnd.n4066 gnd.n4065 585
R2213 gnd.n4064 gnd.n4063 585
R2214 gnd.n4062 gnd.n4061 585
R2215 gnd.n4060 gnd.n4059 585
R2216 gnd.n4058 gnd.n4057 585
R2217 gnd.n4056 gnd.n4055 585
R2218 gnd.n4054 gnd.n4053 585
R2219 gnd.n4052 gnd.n4051 585
R2220 gnd.n4050 gnd.n4049 585
R2221 gnd.n4048 gnd.n4047 585
R2222 gnd.n4046 gnd.n4045 585
R2223 gnd.n4044 gnd.n4043 585
R2224 gnd.n4042 gnd.n4041 585
R2225 gnd.n1135 gnd.n1126 585
R2226 gnd.n2295 gnd.n2294 585
R2227 gnd.n2288 gnd.n2202 585
R2228 gnd.n2290 gnd.n2289 585
R2229 gnd.n2287 gnd.n2286 585
R2230 gnd.n2285 gnd.n2284 585
R2231 gnd.n2278 gnd.n2204 585
R2232 gnd.n2280 gnd.n2279 585
R2233 gnd.n2277 gnd.n2276 585
R2234 gnd.n2275 gnd.n2274 585
R2235 gnd.n2268 gnd.n2206 585
R2236 gnd.n2270 gnd.n2269 585
R2237 gnd.n2267 gnd.n2266 585
R2238 gnd.n2265 gnd.n2264 585
R2239 gnd.n2258 gnd.n2208 585
R2240 gnd.n2260 gnd.n2259 585
R2241 gnd.n2257 gnd.n2256 585
R2242 gnd.n2255 gnd.n2254 585
R2243 gnd.n2248 gnd.n2210 585
R2244 gnd.n2250 gnd.n2249 585
R2245 gnd.n2247 gnd.n2246 585
R2246 gnd.n2245 gnd.n2244 585
R2247 gnd.n2238 gnd.n2214 585
R2248 gnd.n2240 gnd.n2239 585
R2249 gnd.n2237 gnd.n2236 585
R2250 gnd.n2235 gnd.n2234 585
R2251 gnd.n2228 gnd.n2216 585
R2252 gnd.n2230 gnd.n2229 585
R2253 gnd.n2227 gnd.n2226 585
R2254 gnd.n2225 gnd.n2224 585
R2255 gnd.n2220 gnd.n2219 585
R2256 gnd.n2218 gnd.n1406 585
R2257 gnd.n3855 gnd.n3854 585
R2258 gnd.n3857 gnd.n3856 585
R2259 gnd.n3859 gnd.n3858 585
R2260 gnd.n3861 gnd.n3860 585
R2261 gnd.n3863 gnd.n3862 585
R2262 gnd.n3865 gnd.n3864 585
R2263 gnd.n3867 gnd.n3866 585
R2264 gnd.n3869 gnd.n3868 585
R2265 gnd.n3872 gnd.n3871 585
R2266 gnd.n3874 gnd.n3873 585
R2267 gnd.n3876 gnd.n3875 585
R2268 gnd.n3878 gnd.n3877 585
R2269 gnd.n3880 gnd.n3879 585
R2270 gnd.n3882 gnd.n3881 585
R2271 gnd.n3884 gnd.n3883 585
R2272 gnd.n3886 gnd.n3885 585
R2273 gnd.n3888 gnd.n3887 585
R2274 gnd.n3890 gnd.n3889 585
R2275 gnd.n3892 gnd.n3891 585
R2276 gnd.n3894 gnd.n3893 585
R2277 gnd.n3896 gnd.n3895 585
R2278 gnd.n3898 gnd.n3897 585
R2279 gnd.n3899 gnd.n1379 585
R2280 gnd.n3901 gnd.n3900 585
R2281 gnd.n1338 gnd.n1337 585
R2282 gnd.n3905 gnd.n3904 585
R2283 gnd.n3904 gnd.n3903 585
R2284 gnd.n2537 gnd.n2296 585
R2285 gnd.n2598 gnd.n2296 585
R2286 gnd.n2538 gnd.n1330 585
R2287 gnd.n3911 gnd.n1330 585
R2288 gnd.n2539 gnd.n2316 585
R2289 gnd.n2565 gnd.n2316 585
R2290 gnd.n2540 gnd.n1321 585
R2291 gnd.n3917 gnd.n1321 585
R2292 gnd.n2542 gnd.n2541 585
R2293 gnd.n2543 gnd.n2542 585
R2294 gnd.n2534 gnd.n1310 585
R2295 gnd.n3923 gnd.n1310 585
R2296 gnd.n2533 gnd.n2532 585
R2297 gnd.n2532 gnd.n2531 585
R2298 gnd.n2381 gnd.n1300 585
R2299 gnd.n3929 gnd.n1300 585
R2300 gnd.n2380 gnd.n2379 585
R2301 gnd.n2379 gnd.n1299 585
R2302 gnd.n2377 gnd.n1289 585
R2303 gnd.n3935 gnd.n1289 585
R2304 gnd.n2376 gnd.n2375 585
R2305 gnd.n2375 gnd.n1282 585
R2306 gnd.n2374 gnd.n1280 585
R2307 gnd.n3941 gnd.n1280 585
R2308 gnd.n2373 gnd.n2372 585
R2309 gnd.n2372 gnd.n1272 585
R2310 gnd.n2370 gnd.n1270 585
R2311 gnd.n3947 gnd.n1270 585
R2312 gnd.n2369 gnd.n2368 585
R2313 gnd.n2368 gnd.n1269 585
R2314 gnd.n2367 gnd.n1261 585
R2315 gnd.n3953 gnd.n1261 585
R2316 gnd.n2366 gnd.n2365 585
R2317 gnd.n2365 gnd.n1253 585
R2318 gnd.n2363 gnd.n1251 585
R2319 gnd.n3959 gnd.n1251 585
R2320 gnd.n2362 gnd.n2361 585
R2321 gnd.n2361 gnd.n1244 585
R2322 gnd.n2360 gnd.n1242 585
R2323 gnd.n3965 gnd.n1242 585
R2324 gnd.n2359 gnd.n2358 585
R2325 gnd.n2358 gnd.n1234 585
R2326 gnd.n2356 gnd.n1232 585
R2327 gnd.n3971 gnd.n1232 585
R2328 gnd.n2355 gnd.n2354 585
R2329 gnd.n2354 gnd.n1231 585
R2330 gnd.n2353 gnd.n1223 585
R2331 gnd.n3977 gnd.n1223 585
R2332 gnd.n2352 gnd.n2351 585
R2333 gnd.n2351 gnd.n1222 585
R2334 gnd.n2349 gnd.n1213 585
R2335 gnd.n3983 gnd.n1213 585
R2336 gnd.n2348 gnd.n2347 585
R2337 gnd.n2347 gnd.n1206 585
R2338 gnd.n2346 gnd.n1204 585
R2339 gnd.n3989 gnd.n1204 585
R2340 gnd.n2345 gnd.n2344 585
R2341 gnd.n2344 gnd.n1196 585
R2342 gnd.n2342 gnd.n1194 585
R2343 gnd.n3995 gnd.n1194 585
R2344 gnd.n2341 gnd.n2340 585
R2345 gnd.n2340 gnd.n1193 585
R2346 gnd.n2339 gnd.n1185 585
R2347 gnd.n4001 gnd.n1185 585
R2348 gnd.n2338 gnd.n2337 585
R2349 gnd.n2337 gnd.n1184 585
R2350 gnd.n2335 gnd.n1175 585
R2351 gnd.n4007 gnd.n1175 585
R2352 gnd.n2334 gnd.n2333 585
R2353 gnd.n2333 gnd.n1168 585
R2354 gnd.n2332 gnd.n1166 585
R2355 gnd.n4013 gnd.n1166 585
R2356 gnd.n2331 gnd.n2330 585
R2357 gnd.n2330 gnd.n1159 585
R2358 gnd.n2328 gnd.n1157 585
R2359 gnd.n4019 gnd.n1157 585
R2360 gnd.n2327 gnd.n2326 585
R2361 gnd.n2326 gnd.n1149 585
R2362 gnd.n2325 gnd.n1147 585
R2363 gnd.n4025 gnd.n1147 585
R2364 gnd.n2324 gnd.n2323 585
R2365 gnd.n2323 gnd.n1146 585
R2366 gnd.n2321 gnd.n1137 585
R2367 gnd.n4033 gnd.n1137 585
R2368 gnd.n1136 gnd.n1130 585
R2369 gnd.n1136 gnd.n1061 585
R2370 gnd.n161 gnd.n160 585
R2371 gnd.n164 gnd.n161 585
R2372 gnd.n7055 gnd.n7054 585
R2373 gnd.n7054 gnd.n7053 585
R2374 gnd.n7056 gnd.n155 585
R2375 gnd.n155 gnd.n154 585
R2376 gnd.n7058 gnd.n7057 585
R2377 gnd.n7059 gnd.n7058 585
R2378 gnd.n141 gnd.n140 585
R2379 gnd.n145 gnd.n141 585
R2380 gnd.n7067 gnd.n7066 585
R2381 gnd.n7066 gnd.n7065 585
R2382 gnd.n7068 gnd.n135 585
R2383 gnd.n142 gnd.n135 585
R2384 gnd.n7070 gnd.n7069 585
R2385 gnd.n7071 gnd.n7070 585
R2386 gnd.n123 gnd.n122 585
R2387 gnd.n126 gnd.n123 585
R2388 gnd.n7079 gnd.n7078 585
R2389 gnd.n7078 gnd.n7077 585
R2390 gnd.n7080 gnd.n117 585
R2391 gnd.n117 gnd.n116 585
R2392 gnd.n7082 gnd.n7081 585
R2393 gnd.n7083 gnd.n7082 585
R2394 gnd.n103 gnd.n102 585
R2395 gnd.n107 gnd.n103 585
R2396 gnd.n7091 gnd.n7090 585
R2397 gnd.n7090 gnd.n7089 585
R2398 gnd.n7092 gnd.n97 585
R2399 gnd.n104 gnd.n97 585
R2400 gnd.n7094 gnd.n7093 585
R2401 gnd.n7095 gnd.n7094 585
R2402 gnd.n83 gnd.n82 585
R2403 gnd.n86 gnd.n83 585
R2404 gnd.n7103 gnd.n7102 585
R2405 gnd.n7102 gnd.n7101 585
R2406 gnd.n7104 gnd.n77 585
R2407 gnd.n77 gnd.n74 585
R2408 gnd.n7106 gnd.n7105 585
R2409 gnd.n7107 gnd.n7106 585
R2410 gnd.n78 gnd.n76 585
R2411 gnd.n6680 gnd.n76 585
R2412 gnd.n6669 gnd.n181 585
R2413 gnd.n181 gnd.n171 585
R2414 gnd.n6671 gnd.n6670 585
R2415 gnd.n6672 gnd.n6671 585
R2416 gnd.n182 gnd.n180 585
R2417 gnd.n188 gnd.n180 585
R2418 gnd.n6663 gnd.n6662 585
R2419 gnd.n6662 gnd.n6661 585
R2420 gnd.n185 gnd.n184 585
R2421 gnd.n6652 gnd.n185 585
R2422 gnd.n6636 gnd.n204 585
R2423 gnd.n204 gnd.n194 585
R2424 gnd.n6638 gnd.n6637 585
R2425 gnd.n6639 gnd.n6638 585
R2426 gnd.n205 gnd.n203 585
R2427 gnd.n212 gnd.n203 585
R2428 gnd.n6631 gnd.n6630 585
R2429 gnd.n6630 gnd.n6629 585
R2430 gnd.n208 gnd.n207 585
R2431 gnd.n209 gnd.n208 585
R2432 gnd.n6612 gnd.n6611 585
R2433 gnd.n6613 gnd.n6612 585
R2434 gnd.n225 gnd.n224 585
R2435 gnd.n224 gnd.n221 585
R2436 gnd.n6607 gnd.n6606 585
R2437 gnd.n6606 gnd.n6605 585
R2438 gnd.n228 gnd.n227 585
R2439 gnd.n6594 gnd.n228 585
R2440 gnd.n6572 gnd.n250 585
R2441 gnd.n250 gnd.n239 585
R2442 gnd.n6574 gnd.n6573 585
R2443 gnd.n6575 gnd.n6574 585
R2444 gnd.n251 gnd.n249 585
R2445 gnd.n6553 gnd.n249 585
R2446 gnd.n6567 gnd.n6566 585
R2447 gnd.n6566 gnd.n6565 585
R2448 gnd.n254 gnd.n253 585
R2449 gnd.n6549 gnd.n254 585
R2450 gnd.n280 gnd.n278 585
R2451 gnd.n6323 gnd.n278 585
R2452 gnd.n6539 gnd.n6538 585
R2453 gnd.n6540 gnd.n6539 585
R2454 gnd.n279 gnd.n277 585
R2455 gnd.n6329 gnd.n277 585
R2456 gnd.n6533 gnd.n6532 585
R2457 gnd.n283 gnd.n282 585
R2458 gnd.n6529 gnd.n6528 585
R2459 gnd.n6530 gnd.n6529 585
R2460 gnd.n6527 gnd.n324 585
R2461 gnd.n6526 gnd.n6525 585
R2462 gnd.n6524 gnd.n6523 585
R2463 gnd.n6522 gnd.n6521 585
R2464 gnd.n6520 gnd.n6519 585
R2465 gnd.n6518 gnd.n6517 585
R2466 gnd.n6516 gnd.n6515 585
R2467 gnd.n6514 gnd.n6513 585
R2468 gnd.n6512 gnd.n6511 585
R2469 gnd.n6510 gnd.n6509 585
R2470 gnd.n6508 gnd.n6507 585
R2471 gnd.n6506 gnd.n6505 585
R2472 gnd.n6504 gnd.n6503 585
R2473 gnd.n6502 gnd.n6501 585
R2474 gnd.n6500 gnd.n6499 585
R2475 gnd.n6497 gnd.n6496 585
R2476 gnd.n6495 gnd.n6494 585
R2477 gnd.n6493 gnd.n6492 585
R2478 gnd.n6491 gnd.n6490 585
R2479 gnd.n6489 gnd.n6488 585
R2480 gnd.n6487 gnd.n6486 585
R2481 gnd.n6485 gnd.n6484 585
R2482 gnd.n6483 gnd.n6482 585
R2483 gnd.n6480 gnd.n6479 585
R2484 gnd.n6478 gnd.n6477 585
R2485 gnd.n6476 gnd.n6475 585
R2486 gnd.n6474 gnd.n6473 585
R2487 gnd.n6472 gnd.n6471 585
R2488 gnd.n6470 gnd.n6469 585
R2489 gnd.n6468 gnd.n6467 585
R2490 gnd.n6466 gnd.n6465 585
R2491 gnd.n6464 gnd.n6463 585
R2492 gnd.n6462 gnd.n6461 585
R2493 gnd.n6460 gnd.n6459 585
R2494 gnd.n6458 gnd.n6457 585
R2495 gnd.n6456 gnd.n6455 585
R2496 gnd.n6454 gnd.n6453 585
R2497 gnd.n6452 gnd.n6451 585
R2498 gnd.n6450 gnd.n6449 585
R2499 gnd.n6448 gnd.n6447 585
R2500 gnd.n6446 gnd.n6445 585
R2501 gnd.n6444 gnd.n6443 585
R2502 gnd.n6442 gnd.n6441 585
R2503 gnd.n6440 gnd.n6439 585
R2504 gnd.n6438 gnd.n6437 585
R2505 gnd.n6436 gnd.n6435 585
R2506 gnd.n6434 gnd.n6433 585
R2507 gnd.n6432 gnd.n6431 585
R2508 gnd.n6430 gnd.n6429 585
R2509 gnd.n6428 gnd.n6427 585
R2510 gnd.n6426 gnd.n6425 585
R2511 gnd.n6424 gnd.n6423 585
R2512 gnd.n6422 gnd.n6421 585
R2513 gnd.n500 gnd.n385 585
R2514 gnd.n7046 gnd.n7045 585
R2515 gnd.n6723 gnd.n6722 585
R2516 gnd.n6923 gnd.n6922 585
R2517 gnd.n6925 gnd.n6924 585
R2518 gnd.n6927 gnd.n6926 585
R2519 gnd.n6929 gnd.n6928 585
R2520 gnd.n6931 gnd.n6930 585
R2521 gnd.n6933 gnd.n6932 585
R2522 gnd.n6935 gnd.n6934 585
R2523 gnd.n6937 gnd.n6936 585
R2524 gnd.n6939 gnd.n6938 585
R2525 gnd.n6941 gnd.n6940 585
R2526 gnd.n6943 gnd.n6942 585
R2527 gnd.n6945 gnd.n6944 585
R2528 gnd.n6947 gnd.n6946 585
R2529 gnd.n6949 gnd.n6948 585
R2530 gnd.n6951 gnd.n6950 585
R2531 gnd.n6953 gnd.n6952 585
R2532 gnd.n6955 gnd.n6954 585
R2533 gnd.n6958 gnd.n6957 585
R2534 gnd.n6956 gnd.n6902 585
R2535 gnd.n6963 gnd.n6962 585
R2536 gnd.n6965 gnd.n6964 585
R2537 gnd.n6967 gnd.n6966 585
R2538 gnd.n6969 gnd.n6968 585
R2539 gnd.n6971 gnd.n6970 585
R2540 gnd.n6973 gnd.n6972 585
R2541 gnd.n6975 gnd.n6974 585
R2542 gnd.n6977 gnd.n6976 585
R2543 gnd.n6979 gnd.n6978 585
R2544 gnd.n6981 gnd.n6980 585
R2545 gnd.n6983 gnd.n6982 585
R2546 gnd.n6985 gnd.n6984 585
R2547 gnd.n6987 gnd.n6986 585
R2548 gnd.n6989 gnd.n6988 585
R2549 gnd.n6991 gnd.n6990 585
R2550 gnd.n6993 gnd.n6992 585
R2551 gnd.n6995 gnd.n6994 585
R2552 gnd.n6997 gnd.n6996 585
R2553 gnd.n6999 gnd.n6998 585
R2554 gnd.n7001 gnd.n7000 585
R2555 gnd.n7006 gnd.n7005 585
R2556 gnd.n7008 gnd.n7007 585
R2557 gnd.n7010 gnd.n7009 585
R2558 gnd.n7012 gnd.n7011 585
R2559 gnd.n7014 gnd.n7013 585
R2560 gnd.n7016 gnd.n7015 585
R2561 gnd.n7018 gnd.n7017 585
R2562 gnd.n7020 gnd.n7019 585
R2563 gnd.n7022 gnd.n7021 585
R2564 gnd.n7024 gnd.n7023 585
R2565 gnd.n7026 gnd.n7025 585
R2566 gnd.n7028 gnd.n7027 585
R2567 gnd.n7030 gnd.n7029 585
R2568 gnd.n7032 gnd.n7031 585
R2569 gnd.n7035 gnd.n7034 585
R2570 gnd.n7033 gnd.n6868 585
R2571 gnd.n7039 gnd.n6865 585
R2572 gnd.n7041 gnd.n7040 585
R2573 gnd.n7042 gnd.n7041 585
R2574 gnd.n7044 gnd.n6717 585
R2575 gnd.n7044 gnd.n164 585
R2576 gnd.n6716 gnd.n162 585
R2577 gnd.n7053 gnd.n162 585
R2578 gnd.n6715 gnd.n6714 585
R2579 gnd.n6714 gnd.n154 585
R2580 gnd.n6712 gnd.n152 585
R2581 gnd.n7059 gnd.n152 585
R2582 gnd.n6711 gnd.n6710 585
R2583 gnd.n6710 gnd.n145 585
R2584 gnd.n6709 gnd.n143 585
R2585 gnd.n7065 gnd.n143 585
R2586 gnd.n6708 gnd.n6707 585
R2587 gnd.n6707 gnd.n142 585
R2588 gnd.n6705 gnd.n133 585
R2589 gnd.n7071 gnd.n133 585
R2590 gnd.n6704 gnd.n6703 585
R2591 gnd.n6703 gnd.n126 585
R2592 gnd.n6702 gnd.n124 585
R2593 gnd.n7077 gnd.n124 585
R2594 gnd.n6701 gnd.n6700 585
R2595 gnd.n6700 gnd.n116 585
R2596 gnd.n6698 gnd.n114 585
R2597 gnd.n7083 gnd.n114 585
R2598 gnd.n6697 gnd.n6696 585
R2599 gnd.n6696 gnd.n107 585
R2600 gnd.n6695 gnd.n105 585
R2601 gnd.n7089 gnd.n105 585
R2602 gnd.n6694 gnd.n6693 585
R2603 gnd.n6693 gnd.n104 585
R2604 gnd.n6691 gnd.n95 585
R2605 gnd.n7095 gnd.n95 585
R2606 gnd.n6690 gnd.n6689 585
R2607 gnd.n6689 gnd.n86 585
R2608 gnd.n6688 gnd.n84 585
R2609 gnd.n7101 gnd.n84 585
R2610 gnd.n6687 gnd.n6686 585
R2611 gnd.n6686 gnd.n74 585
R2612 gnd.n167 gnd.n73 585
R2613 gnd.n7107 gnd.n73 585
R2614 gnd.n6679 gnd.n6678 585
R2615 gnd.n6680 gnd.n6679 585
R2616 gnd.n6677 gnd.n172 585
R2617 gnd.n172 gnd.n171 585
R2618 gnd.n177 gnd.n173 585
R2619 gnd.n6672 gnd.n177 585
R2620 gnd.n6656 gnd.n6655 585
R2621 gnd.n6655 gnd.n188 585
R2622 gnd.n6657 gnd.n186 585
R2623 gnd.n6661 gnd.n186 585
R2624 gnd.n6654 gnd.n6653 585
R2625 gnd.n6653 gnd.n6652 585
R2626 gnd.n193 gnd.n192 585
R2627 gnd.n194 gnd.n193 585
R2628 gnd.n6620 gnd.n201 585
R2629 gnd.n6639 gnd.n201 585
R2630 gnd.n6619 gnd.n6618 585
R2631 gnd.n6618 gnd.n212 585
R2632 gnd.n6617 gnd.n210 585
R2633 gnd.n6629 gnd.n210 585
R2634 gnd.n6616 gnd.n6615 585
R2635 gnd.n6615 gnd.n209 585
R2636 gnd.n6614 gnd.n218 585
R2637 gnd.n6614 gnd.n6613 585
R2638 gnd.n6598 gnd.n220 585
R2639 gnd.n221 gnd.n220 585
R2640 gnd.n6597 gnd.n230 585
R2641 gnd.n6605 gnd.n230 585
R2642 gnd.n6596 gnd.n6595 585
R2643 gnd.n6595 gnd.n6594 585
R2644 gnd.n238 gnd.n236 585
R2645 gnd.n239 gnd.n238 585
R2646 gnd.n6556 gnd.n247 585
R2647 gnd.n6575 gnd.n247 585
R2648 gnd.n6555 gnd.n6554 585
R2649 gnd.n6554 gnd.n6553 585
R2650 gnd.n6552 gnd.n256 585
R2651 gnd.n6565 gnd.n256 585
R2652 gnd.n6551 gnd.n6550 585
R2653 gnd.n6550 gnd.n6549 585
R2654 gnd.n266 gnd.n264 585
R2655 gnd.n6323 gnd.n266 585
R2656 gnd.n504 gnd.n275 585
R2657 gnd.n6540 gnd.n275 585
R2658 gnd.n503 gnd.n501 585
R2659 gnd.n6329 gnd.n501 585
R2660 gnd.n1007 gnd.n1006 585
R2661 gnd.n1291 gnd.n1007 585
R2662 gnd.n6310 gnd.n6309 585
R2663 gnd.n6309 gnd.n229 585
R2664 gnd.n6313 gnd.n517 585
R2665 gnd.n517 gnd.n516 585
R2666 gnd.n6315 gnd.n6314 585
R2667 gnd.n6315 gnd.n246 585
R2668 gnd.n6316 gnd.n515 585
R2669 gnd.n6316 gnd.n258 585
R2670 gnd.n6318 gnd.n6317 585
R2671 gnd.n6317 gnd.n255 585
R2672 gnd.n6319 gnd.n507 585
R2673 gnd.n507 gnd.n267 585
R2674 gnd.n6321 gnd.n6320 585
R2675 gnd.n6322 gnd.n6321 585
R2676 gnd.n508 gnd.n498 585
R2677 gnd.n498 gnd.n274 585
R2678 gnd.n6331 gnd.n499 585
R2679 gnd.n6331 gnd.n6330 585
R2680 gnd.n6332 gnd.n497 585
R2681 gnd.n6332 gnd.n323 585
R2682 gnd.n6334 gnd.n6333 585
R2683 gnd.n6333 gnd.n284 585
R2684 gnd.n6335 gnd.n492 585
R2685 gnd.n492 gnd.n490 585
R2686 gnd.n6337 gnd.n6336 585
R2687 gnd.n6338 gnd.n6337 585
R2688 gnd.n493 gnd.n491 585
R2689 gnd.n491 gnd.n470 585
R2690 gnd.n3656 gnd.n3655 585
R2691 gnd.n3655 gnd.n458 585
R2692 gnd.n3657 gnd.n1576 585
R2693 gnd.n1576 gnd.n457 585
R2694 gnd.n3659 gnd.n3658 585
R2695 gnd.n3660 gnd.n3659 585
R2696 gnd.n1577 gnd.n1575 585
R2697 gnd.n1575 gnd.n1572 585
R2698 gnd.n3648 gnd.n3647 585
R2699 gnd.n3647 gnd.n3646 585
R2700 gnd.n1580 gnd.n1579 585
R2701 gnd.n3635 gnd.n1580 585
R2702 gnd.n3633 gnd.n3632 585
R2703 gnd.n3634 gnd.n3633 585
R2704 gnd.n1591 gnd.n1590 585
R2705 gnd.n3624 gnd.n1590 585
R2706 gnd.n3628 gnd.n3627 585
R2707 gnd.n3627 gnd.n3626 585
R2708 gnd.n1594 gnd.n1593 585
R2709 gnd.n3615 gnd.n1594 585
R2710 gnd.n3613 gnd.n3612 585
R2711 gnd.n3614 gnd.n3613 585
R2712 gnd.n1604 gnd.n1603 585
R2713 gnd.n3604 gnd.n1603 585
R2714 gnd.n3608 gnd.n3607 585
R2715 gnd.n3607 gnd.n3606 585
R2716 gnd.n1607 gnd.n1606 585
R2717 gnd.n3595 gnd.n1607 585
R2718 gnd.n3593 gnd.n3592 585
R2719 gnd.n3594 gnd.n3593 585
R2720 gnd.n1617 gnd.n1616 585
R2721 gnd.n3584 gnd.n1616 585
R2722 gnd.n3588 gnd.n3587 585
R2723 gnd.n3587 gnd.n3586 585
R2724 gnd.n1620 gnd.n1619 585
R2725 gnd.n3575 gnd.n1620 585
R2726 gnd.n3571 gnd.n3570 585
R2727 gnd.n3572 gnd.n3571 585
R2728 gnd.n1628 gnd.n1627 585
R2729 gnd.n3562 gnd.n1627 585
R2730 gnd.n3566 gnd.n3565 585
R2731 gnd.n3565 gnd.n3564 585
R2732 gnd.n1631 gnd.n1630 585
R2733 gnd.n3553 gnd.n1631 585
R2734 gnd.n3551 gnd.n3550 585
R2735 gnd.n3552 gnd.n3551 585
R2736 gnd.n1641 gnd.n1640 585
R2737 gnd.n1671 gnd.n1640 585
R2738 gnd.n3546 gnd.n3545 585
R2739 gnd.n3545 gnd.n3544 585
R2740 gnd.n1644 gnd.n1643 585
R2741 gnd.n1723 gnd.n1644 585
R2742 gnd.n3404 gnd.n3403 585
R2743 gnd.n3405 gnd.n3404 585
R2744 gnd.n1733 gnd.n1732 585
R2745 gnd.n3372 gnd.n1732 585
R2746 gnd.n3399 gnd.n3398 585
R2747 gnd.n3398 gnd.n3397 585
R2748 gnd.n1736 gnd.n1735 585
R2749 gnd.n3380 gnd.n1736 585
R2750 gnd.n3362 gnd.n3361 585
R2751 gnd.n3363 gnd.n3362 585
R2752 gnd.n1749 gnd.n1748 585
R2753 gnd.n3326 gnd.n1748 585
R2754 gnd.n3357 gnd.n3356 585
R2755 gnd.n3356 gnd.n3355 585
R2756 gnd.n1752 gnd.n1751 585
R2757 gnd.n1765 gnd.n1752 585
R2758 gnd.n3321 gnd.n3320 585
R2759 gnd.n3322 gnd.n3321 585
R2760 gnd.n1772 gnd.n1771 585
R2761 gnd.n1779 gnd.n1771 585
R2762 gnd.n3316 gnd.n3315 585
R2763 gnd.n3315 gnd.n3314 585
R2764 gnd.n1775 gnd.n1774 585
R2765 gnd.n1784 gnd.n1775 585
R2766 gnd.n3274 gnd.n1800 585
R2767 gnd.n1800 gnd.n1794 585
R2768 gnd.n3276 gnd.n3275 585
R2769 gnd.n3277 gnd.n3276 585
R2770 gnd.n1801 gnd.n1799 585
R2771 gnd.n3210 gnd.n1799 585
R2772 gnd.n3269 gnd.n3268 585
R2773 gnd.n3268 gnd.n3267 585
R2774 gnd.n1804 gnd.n1803 585
R2775 gnd.n3259 gnd.n1804 585
R2776 gnd.n3247 gnd.n3246 585
R2777 gnd.n3248 gnd.n3247 585
R2778 gnd.n1822 gnd.n1821 585
R2779 gnd.n3221 gnd.n1821 585
R2780 gnd.n3242 gnd.n3241 585
R2781 gnd.n3241 gnd.n3240 585
R2782 gnd.n1825 gnd.n1824 585
R2783 gnd.n3229 gnd.n1825 585
R2784 gnd.n3188 gnd.n3187 585
R2785 gnd.n3189 gnd.n3188 585
R2786 gnd.n1839 gnd.n1838 585
R2787 gnd.n1847 gnd.n1838 585
R2788 gnd.n3183 gnd.n3182 585
R2789 gnd.n3182 gnd.n3181 585
R2790 gnd.n1842 gnd.n1841 585
R2791 gnd.n1855 gnd.n1842 585
R2792 gnd.n3147 gnd.n3146 585
R2793 gnd.n3148 gnd.n3147 585
R2794 gnd.n1863 gnd.n1862 585
R2795 gnd.n1870 gnd.n1862 585
R2796 gnd.n3142 gnd.n3141 585
R2797 gnd.n3141 gnd.n3140 585
R2798 gnd.n1866 gnd.n1865 585
R2799 gnd.n1876 gnd.n1866 585
R2800 gnd.n3102 gnd.n1894 585
R2801 gnd.n1894 gnd.n1886 585
R2802 gnd.n3104 gnd.n3103 585
R2803 gnd.n3105 gnd.n3104 585
R2804 gnd.n1895 gnd.n1893 585
R2805 gnd.n3037 gnd.n1893 585
R2806 gnd.n3097 gnd.n3096 585
R2807 gnd.n3096 gnd.n3095 585
R2808 gnd.n1898 gnd.n1897 585
R2809 gnd.n3087 gnd.n1898 585
R2810 gnd.n3074 gnd.n3073 585
R2811 gnd.n3075 gnd.n3074 585
R2812 gnd.n1917 gnd.n1916 585
R2813 gnd.n3048 gnd.n1916 585
R2814 gnd.n3069 gnd.n3068 585
R2815 gnd.n3068 gnd.n3067 585
R2816 gnd.n1920 gnd.n1919 585
R2817 gnd.n3056 gnd.n1920 585
R2818 gnd.n3018 gnd.n3017 585
R2819 gnd.n3019 gnd.n3018 585
R2820 gnd.n1935 gnd.n1934 585
R2821 gnd.n3003 gnd.n1934 585
R2822 gnd.n3013 gnd.n3012 585
R2823 gnd.n3012 gnd.n3011 585
R2824 gnd.n1938 gnd.n1937 585
R2825 gnd.n1946 gnd.n1938 585
R2826 gnd.n2974 gnd.n2973 585
R2827 gnd.n2975 gnd.n2974 585
R2828 gnd.n1958 gnd.n1957 585
R2829 gnd.n1964 gnd.n1957 585
R2830 gnd.n2969 gnd.n2968 585
R2831 gnd.n2968 gnd.n2967 585
R2832 gnd.n1961 gnd.n1960 585
R2833 gnd.n1969 gnd.n1961 585
R2834 gnd.n2932 gnd.n1985 585
R2835 gnd.n1985 gnd.n1978 585
R2836 gnd.n2934 gnd.n2933 585
R2837 gnd.n2935 gnd.n2934 585
R2838 gnd.n1986 gnd.n1984 585
R2839 gnd.n2908 gnd.n1984 585
R2840 gnd.n2927 gnd.n2926 585
R2841 gnd.n2926 gnd.n2925 585
R2842 gnd.n1989 gnd.n1988 585
R2843 gnd.n2917 gnd.n1989 585
R2844 gnd.n2786 gnd.n2782 585
R2845 gnd.n2782 gnd.n1474 585
R2846 gnd.n2788 gnd.n2787 585
R2847 gnd.n2788 gnd.n1471 585
R2848 gnd.n2789 gnd.n2781 585
R2849 gnd.n2789 gnd.n1445 585
R2850 gnd.n2791 gnd.n2790 585
R2851 gnd.n2790 gnd.n2003 585
R2852 gnd.n2792 gnd.n2015 585
R2853 gnd.n2015 gnd.n2002 585
R2854 gnd.n2794 gnd.n2793 585
R2855 gnd.n2795 gnd.n2794 585
R2856 gnd.n2016 gnd.n2014 585
R2857 gnd.n2014 gnd.n2011 585
R2858 gnd.n2775 gnd.n2774 585
R2859 gnd.n2774 gnd.n2773 585
R2860 gnd.n2019 gnd.n2018 585
R2861 gnd.n2027 gnd.n2019 585
R2862 gnd.n2747 gnd.n2040 585
R2863 gnd.n2040 gnd.n2039 585
R2864 gnd.n2749 gnd.n2748 585
R2865 gnd.n2750 gnd.n2749 585
R2866 gnd.n2041 gnd.n2038 585
R2867 gnd.n2038 gnd.n2035 585
R2868 gnd.n2742 gnd.n2741 585
R2869 gnd.n2741 gnd.n2740 585
R2870 gnd.n2044 gnd.n2043 585
R2871 gnd.n2053 gnd.n2044 585
R2872 gnd.n2717 gnd.n2065 585
R2873 gnd.n2065 gnd.n2052 585
R2874 gnd.n2719 gnd.n2718 585
R2875 gnd.n2720 gnd.n2719 585
R2876 gnd.n2066 gnd.n2064 585
R2877 gnd.n2064 gnd.n2061 585
R2878 gnd.n2712 gnd.n2711 585
R2879 gnd.n2711 gnd.n2710 585
R2880 gnd.n2069 gnd.n2068 585
R2881 gnd.n2078 gnd.n2069 585
R2882 gnd.n2687 gnd.n2090 585
R2883 gnd.n2090 gnd.n2077 585
R2884 gnd.n2689 gnd.n2688 585
R2885 gnd.n2690 gnd.n2689 585
R2886 gnd.n2091 gnd.n2089 585
R2887 gnd.n2089 gnd.n2086 585
R2888 gnd.n2682 gnd.n2681 585
R2889 gnd.n2681 gnd.n2680 585
R2890 gnd.n2094 gnd.n2093 585
R2891 gnd.n2103 gnd.n2094 585
R2892 gnd.n2582 gnd.n2581 585
R2893 gnd.n2582 gnd.n2102 585
R2894 gnd.n2586 gnd.n2585 585
R2895 gnd.n2585 gnd.n2584 585
R2896 gnd.n2587 gnd.n2575 585
R2897 gnd.n2575 gnd.n2125 585
R2898 gnd.n2589 gnd.n2588 585
R2899 gnd.n2589 gnd.n2111 585
R2900 gnd.n2591 gnd.n2574 585
R2901 gnd.n2591 gnd.n2590 585
R2902 gnd.n2593 gnd.n2592 585
R2903 gnd.n2592 gnd.n1350 585
R2904 gnd.n2594 gnd.n2298 585
R2905 gnd.n2298 gnd.n1339 585
R2906 gnd.n2596 gnd.n2595 585
R2907 gnd.n2597 gnd.n2596 585
R2908 gnd.n2299 gnd.n2297 585
R2909 gnd.n2297 gnd.n1332 585
R2910 gnd.n2568 gnd.n2567 585
R2911 gnd.n2567 gnd.n2566 585
R2912 gnd.n2315 gnd.n2301 585
R2913 gnd.n2315 gnd.n1323 585
R2914 gnd.n2314 gnd.n2313 585
R2915 gnd.n2314 gnd.n1320 585
R2916 gnd.n2303 gnd.n2302 585
R2917 gnd.n2302 gnd.n1312 585
R2918 gnd.n2309 gnd.n2308 585
R2919 gnd.n2308 gnd.n1309 585
R2920 gnd.n2307 gnd.n2306 585
R2921 gnd.n2307 gnd.n1302 585
R2922 gnd.n6354 gnd.n6353 585
R2923 gnd.n6355 gnd.n6354 585
R2924 gnd.n461 gnd.n459 585
R2925 gnd.n1574 gnd.n459 585
R2926 gnd.n3663 gnd.n3662 585
R2927 gnd.n3662 gnd.n3661 585
R2928 gnd.n3664 gnd.n1571 585
R2929 gnd.n3645 gnd.n1571 585
R2930 gnd.n1581 gnd.n1569 585
R2931 gnd.n1582 gnd.n1581 585
R2932 gnd.n3668 gnd.n1568 585
R2933 gnd.n3636 gnd.n1568 585
R2934 gnd.n3669 gnd.n1567 585
R2935 gnd.n1589 gnd.n1567 585
R2936 gnd.n3670 gnd.n1566 585
R2937 gnd.n3625 gnd.n1566 585
R2938 gnd.n1595 gnd.n1564 585
R2939 gnd.n1596 gnd.n1595 585
R2940 gnd.n3674 gnd.n1563 585
R2941 gnd.n3616 gnd.n1563 585
R2942 gnd.n3675 gnd.n1562 585
R2943 gnd.n1602 gnd.n1562 585
R2944 gnd.n3676 gnd.n1561 585
R2945 gnd.n3605 gnd.n1561 585
R2946 gnd.n1608 gnd.n1559 585
R2947 gnd.n1609 gnd.n1608 585
R2948 gnd.n3680 gnd.n1558 585
R2949 gnd.n3596 gnd.n1558 585
R2950 gnd.n3681 gnd.n1557 585
R2951 gnd.n1615 gnd.n1557 585
R2952 gnd.n3682 gnd.n1556 585
R2953 gnd.n3585 gnd.n1556 585
R2954 gnd.n3573 gnd.n1554 585
R2955 gnd.n3574 gnd.n3573 585
R2956 gnd.n3686 gnd.n1553 585
R2957 gnd.n3576 gnd.n1553 585
R2958 gnd.n3687 gnd.n1552 585
R2959 gnd.n1626 gnd.n1552 585
R2960 gnd.n3688 gnd.n1551 585
R2961 gnd.n3563 gnd.n1551 585
R2962 gnd.n1632 gnd.n1549 585
R2963 gnd.n1633 gnd.n1632 585
R2964 gnd.n3692 gnd.n1548 585
R2965 gnd.n3554 gnd.n1548 585
R2966 gnd.n3693 gnd.n1547 585
R2967 gnd.n1639 gnd.n1547 585
R2968 gnd.n3694 gnd.n1546 585
R2969 gnd.n1646 gnd.n1546 585
R2970 gnd.n3415 gnd.n1544 585
R2971 gnd.n3416 gnd.n3415 585
R2972 gnd.n3698 gnd.n1543 585
R2973 gnd.n3387 gnd.n1543 585
R2974 gnd.n3699 gnd.n1542 585
R2975 gnd.n3406 gnd.n1542 585
R2976 gnd.n3700 gnd.n1541 585
R2977 gnd.t314 gnd.n1541 585
R2978 gnd.n1737 gnd.n1539 585
R2979 gnd.n1738 gnd.n1737 585
R2980 gnd.n3704 gnd.n1538 585
R2981 gnd.n1744 gnd.n1538 585
R2982 gnd.n3705 gnd.n1537 585
R2983 gnd.n3347 gnd.n1537 585
R2984 gnd.n3706 gnd.n1536 585
R2985 gnd.n1754 gnd.n1536 585
R2986 gnd.n3334 gnd.n1534 585
R2987 gnd.n3335 gnd.n3334 585
R2988 gnd.n3710 gnd.n1533 585
R2989 gnd.n1770 gnd.n1533 585
R2990 gnd.n3711 gnd.n1532 585
R2991 gnd.n3291 gnd.n1532 585
R2992 gnd.n3712 gnd.n1531 585
R2993 gnd.n3313 gnd.n1531 585
R2994 gnd.n3299 gnd.n1529 585
R2995 gnd.n3300 gnd.n3299 585
R2996 gnd.n3716 gnd.n1528 585
R2997 gnd.n3199 gnd.n1528 585
R2998 gnd.n3717 gnd.n1527 585
R2999 gnd.n3285 gnd.n1527 585
R3000 gnd.n3718 gnd.n1526 585
R3001 gnd.n3209 gnd.n1526 585
R3002 gnd.n3207 gnd.n1524 585
R3003 gnd.n3208 gnd.n3207 585
R3004 gnd.n3722 gnd.n1523 585
R3005 gnd.n3258 gnd.n1523 585
R3006 gnd.n3723 gnd.n1522 585
R3007 gnd.n1819 gnd.n1522 585
R3008 gnd.n3724 gnd.n1521 585
R3009 gnd.n3249 gnd.n1521 585
R3010 gnd.n1828 gnd.n1519 585
R3011 gnd.n1829 gnd.n1828 585
R3012 gnd.n3728 gnd.n1518 585
R3013 gnd.n1826 gnd.n1518 585
R3014 gnd.n3729 gnd.n1517 585
R3015 gnd.n1834 gnd.n1517 585
R3016 gnd.n3730 gnd.n1516 585
R3017 gnd.n3173 gnd.n1516 585
R3018 gnd.n3152 gnd.n1514 585
R3019 gnd.n3153 gnd.n3152 585
R3020 gnd.n3734 gnd.n1513 585
R3021 gnd.n3161 gnd.n1513 585
R3022 gnd.n3735 gnd.n1512 585
R3023 gnd.n1861 gnd.n1512 585
R3024 gnd.n3736 gnd.n1511 585
R3025 gnd.n1859 gnd.n1511 585
R3026 gnd.n3138 gnd.n1509 585
R3027 gnd.n3139 gnd.n3138 585
R3028 gnd.n3740 gnd.n1508 585
R3029 gnd.n3125 gnd.n1508 585
R3030 gnd.n3741 gnd.n1507 585
R3031 gnd.n3029 gnd.n1507 585
R3032 gnd.n3742 gnd.n1506 585
R3033 gnd.n3113 gnd.n1506 585
R3034 gnd.n1890 gnd.n1504 585
R3035 gnd.n1891 gnd.n1890 585
R3036 gnd.n3746 gnd.n1503 585
R3037 gnd.n1901 gnd.n1503 585
R3038 gnd.n3747 gnd.n1502 585
R3039 gnd.n3086 gnd.n1502 585
R3040 gnd.n3748 gnd.n1501 585
R3041 gnd.n1905 gnd.n1501 585
R3042 gnd.n3076 gnd.n1499 585
R3043 gnd.n3077 gnd.n3076 585
R3044 gnd.n3752 gnd.n1498 585
R3045 gnd.n1923 gnd.n1498 585
R3046 gnd.n3753 gnd.n1497 585
R3047 gnd.n1921 gnd.n1497 585
R3048 gnd.n3754 gnd.n1496 585
R3049 gnd.n1928 gnd.n1496 585
R3050 gnd.n1932 gnd.n1494 585
R3051 gnd.n1933 gnd.n1932 585
R3052 gnd.n3758 gnd.n1493 585
R3053 gnd.n1940 gnd.n1493 585
R3054 gnd.n3759 gnd.n1492 585
R3055 gnd.n2995 gnd.n1492 585
R3056 gnd.n3760 gnd.n1491 585
R3057 gnd.n2957 gnd.n1491 585
R3058 gnd.n2976 gnd.n1489 585
R3059 gnd.n2977 gnd.n2976 585
R3060 gnd.n3764 gnd.n1488 585
R3061 gnd.n2966 gnd.n1488 585
R3062 gnd.n3765 gnd.n1487 585
R3063 gnd.n2952 gnd.n1487 585
R3064 gnd.n3766 gnd.n1486 585
R3065 gnd.n2900 gnd.n1486 585
R3066 gnd.n2943 gnd.n1484 585
R3067 gnd.n2944 gnd.n2943 585
R3068 gnd.n3770 gnd.n1483 585
R3069 gnd.n1982 gnd.n1483 585
R3070 gnd.n3771 gnd.n1482 585
R3071 gnd.n1991 gnd.n1482 585
R3072 gnd.n3772 gnd.n1481 585
R3073 gnd.n2916 gnd.n1481 585
R3074 gnd.n1478 gnd.n1476 585
R3075 gnd.n2888 gnd.n1476 585
R3076 gnd.n3777 gnd.n3776 585
R3077 gnd.n3778 gnd.n3777 585
R3078 gnd.n1477 gnd.n1475 585
R3079 gnd.n2876 gnd.n1475 585
R3080 gnd.n2007 gnd.n2005 585
R3081 gnd.n2005 gnd.n1413 585
R3082 gnd.n2804 gnd.n2803 585
R3083 gnd.n2805 gnd.n2804 585
R3084 gnd.n2006 gnd.n2004 585
R3085 gnd.n2013 gnd.n2004 585
R3086 gnd.n2798 gnd.n2797 585
R3087 gnd.n2797 gnd.n2796 585
R3088 gnd.n2010 gnd.n2009 585
R3089 gnd.n2772 gnd.n2010 585
R3090 gnd.n2031 gnd.n2029 585
R3091 gnd.n2029 gnd.n2020 585
R3092 gnd.n2759 gnd.n2758 585
R3093 gnd.n2760 gnd.n2759 585
R3094 gnd.n2030 gnd.n2028 585
R3095 gnd.n2037 gnd.n2028 585
R3096 gnd.n2753 gnd.n2752 585
R3097 gnd.n2752 gnd.n2751 585
R3098 gnd.n2034 gnd.n2033 585
R3099 gnd.n2739 gnd.n2034 585
R3100 gnd.n2057 gnd.n2055 585
R3101 gnd.n2055 gnd.n2045 585
R3102 gnd.n2729 gnd.n2728 585
R3103 gnd.n2730 gnd.n2729 585
R3104 gnd.n2056 gnd.n2054 585
R3105 gnd.n2063 gnd.n2054 585
R3106 gnd.n2723 gnd.n2722 585
R3107 gnd.n2722 gnd.n2721 585
R3108 gnd.n2060 gnd.n2059 585
R3109 gnd.n2709 gnd.n2060 585
R3110 gnd.n2082 gnd.n2080 585
R3111 gnd.n2080 gnd.n2070 585
R3112 gnd.n2699 gnd.n2698 585
R3113 gnd.n2700 gnd.n2699 585
R3114 gnd.n2081 gnd.n2079 585
R3115 gnd.n2088 gnd.n2079 585
R3116 gnd.n2693 gnd.n2692 585
R3117 gnd.n2692 gnd.n2691 585
R3118 gnd.n2085 gnd.n2084 585
R3119 gnd.n2679 gnd.n2085 585
R3120 gnd.n2107 gnd.n2105 585
R3121 gnd.n2105 gnd.n2095 585
R3122 gnd.n2669 gnd.n2668 585
R3123 gnd.n2670 gnd.n2669 585
R3124 gnd.n2106 gnd.n2104 585
R3125 gnd.n2583 gnd.n2104 585
R3126 gnd.n2663 gnd.n2662 585
R3127 gnd.n2110 gnd.n2109 585
R3128 gnd.n2659 gnd.n2658 585
R3129 gnd.n2660 gnd.n2659 585
R3130 gnd.n2127 gnd.n2126 585
R3131 gnd.n2654 gnd.n2129 585
R3132 gnd.n2653 gnd.n2130 585
R3133 gnd.n2652 gnd.n2131 585
R3134 gnd.n2133 gnd.n2132 585
R3135 gnd.n2647 gnd.n2136 585
R3136 gnd.n2646 gnd.n2137 585
R3137 gnd.n2146 gnd.n2138 585
R3138 gnd.n2639 gnd.n2147 585
R3139 gnd.n2638 gnd.n2148 585
R3140 gnd.n2150 gnd.n2149 585
R3141 gnd.n2631 gnd.n2156 585
R3142 gnd.n2630 gnd.n2157 585
R3143 gnd.n2166 gnd.n2158 585
R3144 gnd.n2623 gnd.n2167 585
R3145 gnd.n2622 gnd.n2168 585
R3146 gnd.n2170 gnd.n2169 585
R3147 gnd.n2615 gnd.n2176 585
R3148 gnd.n2614 gnd.n2177 585
R3149 gnd.n2186 gnd.n2178 585
R3150 gnd.n2607 gnd.n2187 585
R3151 gnd.n2606 gnd.n2188 585
R3152 gnd.n2550 gnd.n2549 585
R3153 gnd.n2553 gnd.n2552 585
R3154 gnd.n2557 gnd.n2554 585
R3155 gnd.n2556 gnd.n2555 585
R3156 gnd.n6357 gnd.n6356 585
R3157 gnd.n6356 gnd.n6355 585
R3158 gnd.n455 gnd.n454 585
R3159 gnd.n1574 gnd.n455 585
R3160 gnd.n1585 gnd.n1573 585
R3161 gnd.n3661 gnd.n1573 585
R3162 gnd.n3644 gnd.n3643 585
R3163 gnd.n3645 gnd.n3644 585
R3164 gnd.n1584 gnd.n1583 585
R3165 gnd.n1583 gnd.n1582 585
R3166 gnd.n3638 gnd.n3637 585
R3167 gnd.n3637 gnd.n3636 585
R3168 gnd.n1588 gnd.n1587 585
R3169 gnd.n1589 gnd.n1588 585
R3170 gnd.n3623 gnd.n3622 585
R3171 gnd.n3625 gnd.n3623 585
R3172 gnd.n1598 gnd.n1597 585
R3173 gnd.n1597 gnd.n1596 585
R3174 gnd.n3618 gnd.n3617 585
R3175 gnd.n3617 gnd.n3616 585
R3176 gnd.n1601 gnd.n1600 585
R3177 gnd.n1602 gnd.n1601 585
R3178 gnd.n3603 gnd.n3602 585
R3179 gnd.n3605 gnd.n3603 585
R3180 gnd.n1611 gnd.n1610 585
R3181 gnd.n1610 gnd.n1609 585
R3182 gnd.n3598 gnd.n3597 585
R3183 gnd.n3597 gnd.n3596 585
R3184 gnd.n1614 gnd.n1613 585
R3185 gnd.n1615 gnd.n1614 585
R3186 gnd.n3583 gnd.n3582 585
R3187 gnd.n3585 gnd.n3583 585
R3188 gnd.n1622 gnd.n1621 585
R3189 gnd.n3574 gnd.n1621 585
R3190 gnd.n3578 gnd.n3577 585
R3191 gnd.n3577 gnd.n3576 585
R3192 gnd.n1625 gnd.n1624 585
R3193 gnd.n1626 gnd.n1625 585
R3194 gnd.n3561 gnd.n3560 585
R3195 gnd.n3563 gnd.n3561 585
R3196 gnd.n1635 gnd.n1634 585
R3197 gnd.n1634 gnd.n1633 585
R3198 gnd.n3556 gnd.n3555 585
R3199 gnd.n3555 gnd.n3554 585
R3200 gnd.n1638 gnd.n1637 585
R3201 gnd.n1639 gnd.n1638 585
R3202 gnd.n1727 gnd.n1725 585
R3203 gnd.n1725 gnd.n1646 585
R3204 gnd.n3414 gnd.n3413 585
R3205 gnd.n3416 gnd.n3414 585
R3206 gnd.n1726 gnd.n1724 585
R3207 gnd.n3387 gnd.n1724 585
R3208 gnd.n3408 gnd.n3407 585
R3209 gnd.n3407 gnd.n3406 585
R3210 gnd.n1730 gnd.n1729 585
R3211 gnd.t314 gnd.n1730 585
R3212 gnd.n3341 gnd.n3340 585
R3213 gnd.n3340 gnd.n1738 585
R3214 gnd.n1761 gnd.n1759 585
R3215 gnd.n1759 gnd.n1744 585
R3216 gnd.n3346 gnd.n3345 585
R3217 gnd.n3347 gnd.n3346 585
R3218 gnd.n1760 gnd.n1758 585
R3219 gnd.n1758 gnd.n1754 585
R3220 gnd.n3337 gnd.n3336 585
R3221 gnd.n3336 gnd.n3335 585
R3222 gnd.n1764 gnd.n1763 585
R3223 gnd.n1770 gnd.n1764 585
R3224 gnd.n3293 gnd.n3292 585
R3225 gnd.n3292 gnd.n3291 585
R3226 gnd.n1788 gnd.n1777 585
R3227 gnd.n3313 gnd.n1777 585
R3228 gnd.n3298 gnd.n3297 585
R3229 gnd.n3300 gnd.n3298 585
R3230 gnd.n1787 gnd.n1786 585
R3231 gnd.n3199 gnd.n1786 585
R3232 gnd.n3287 gnd.n3286 585
R3233 gnd.n3286 gnd.n3285 585
R3234 gnd.n1791 gnd.n1790 585
R3235 gnd.n3209 gnd.n1791 585
R3236 gnd.n1814 gnd.n1812 585
R3237 gnd.n3208 gnd.n1812 585
R3238 gnd.n3257 gnd.n3256 585
R3239 gnd.n3258 gnd.n3257 585
R3240 gnd.n1813 gnd.n1811 585
R3241 gnd.n1819 gnd.n1811 585
R3242 gnd.n3251 gnd.n3250 585
R3243 gnd.n3250 gnd.n3249 585
R3244 gnd.n1817 gnd.n1816 585
R3245 gnd.n1829 gnd.n1817 585
R3246 gnd.n3167 gnd.n3166 585
R3247 gnd.n3166 gnd.n1826 585
R3248 gnd.n1851 gnd.n1849 585
R3249 gnd.n1849 gnd.n1834 585
R3250 gnd.n3172 gnd.n3171 585
R3251 gnd.n3173 gnd.n3172 585
R3252 gnd.n1850 gnd.n1848 585
R3253 gnd.n3153 gnd.n1848 585
R3254 gnd.n3163 gnd.n3162 585
R3255 gnd.n3162 gnd.n3161 585
R3256 gnd.n1854 gnd.n1853 585
R3257 gnd.n1861 gnd.n1854 585
R3258 gnd.n3119 gnd.n3118 585
R3259 gnd.n3118 gnd.n1859 585
R3260 gnd.n1880 gnd.n1868 585
R3261 gnd.n3139 gnd.n1868 585
R3262 gnd.n3124 gnd.n3123 585
R3263 gnd.n3125 gnd.n3124 585
R3264 gnd.n1879 gnd.n1878 585
R3265 gnd.n3029 gnd.n1878 585
R3266 gnd.n3115 gnd.n3114 585
R3267 gnd.n3114 gnd.n3113 585
R3268 gnd.n1883 gnd.n1882 585
R3269 gnd.n1891 gnd.n1883 585
R3270 gnd.n1910 gnd.n1908 585
R3271 gnd.n1908 gnd.n1901 585
R3272 gnd.n3085 gnd.n3084 585
R3273 gnd.n3086 gnd.n3085 585
R3274 gnd.n1909 gnd.n1907 585
R3275 gnd.n1907 gnd.n1905 585
R3276 gnd.n3079 gnd.n3078 585
R3277 gnd.n3078 gnd.n3077 585
R3278 gnd.n1913 gnd.n1912 585
R3279 gnd.n1923 gnd.n1913 585
R3280 gnd.n2987 gnd.n2985 585
R3281 gnd.n2985 gnd.n1921 585
R3282 gnd.n2988 gnd.n2984 585
R3283 gnd.n2984 gnd.n1928 585
R3284 gnd.n2989 gnd.n2983 585
R3285 gnd.n2983 gnd.n1933 585
R3286 gnd.n1950 gnd.n1948 585
R3287 gnd.n1948 gnd.n1940 585
R3288 gnd.n2994 gnd.n2993 585
R3289 gnd.n2995 gnd.n2994 585
R3290 gnd.n1949 gnd.n1947 585
R3291 gnd.n2957 gnd.n1947 585
R3292 gnd.n2979 gnd.n2978 585
R3293 gnd.n2978 gnd.n2977 585
R3294 gnd.n1953 gnd.n1952 585
R3295 gnd.n2966 gnd.n1953 585
R3296 gnd.n2951 gnd.n2950 585
R3297 gnd.n2952 gnd.n2951 585
R3298 gnd.n1972 gnd.n1971 585
R3299 gnd.n2900 gnd.n1971 585
R3300 gnd.n2946 gnd.n2945 585
R3301 gnd.n2945 gnd.n2944 585
R3302 gnd.n1975 gnd.n1974 585
R3303 gnd.n1982 gnd.n1975 585
R3304 gnd.n2882 gnd.n2881 585
R3305 gnd.n2881 gnd.n1991 585
R3306 gnd.n1997 gnd.n1994 585
R3307 gnd.n2916 gnd.n1994 585
R3308 gnd.n2887 gnd.n2886 585
R3309 gnd.n2888 gnd.n2887 585
R3310 gnd.n1996 gnd.n1473 585
R3311 gnd.n3778 gnd.n1473 585
R3312 gnd.n2878 gnd.n2877 585
R3313 gnd.n2877 gnd.n2876 585
R3314 gnd.n2807 gnd.n1999 585
R3315 gnd.n2807 gnd.n1413 585
R3316 gnd.n2806 gnd.n2001 585
R3317 gnd.n2806 gnd.n2805 585
R3318 gnd.n2766 gnd.n2000 585
R3319 gnd.n2013 gnd.n2000 585
R3320 gnd.n2023 gnd.n2012 585
R3321 gnd.n2796 gnd.n2012 585
R3322 gnd.n2771 gnd.n2770 585
R3323 gnd.n2772 gnd.n2771 585
R3324 gnd.n2022 gnd.n2021 585
R3325 gnd.n2021 gnd.n2020 585
R3326 gnd.n2762 gnd.n2761 585
R3327 gnd.n2761 gnd.n2760 585
R3328 gnd.n2026 gnd.n2025 585
R3329 gnd.n2037 gnd.n2026 585
R3330 gnd.n2048 gnd.n2036 585
R3331 gnd.n2751 gnd.n2036 585
R3332 gnd.n2738 gnd.n2737 585
R3333 gnd.n2739 gnd.n2738 585
R3334 gnd.n2047 gnd.n2046 585
R3335 gnd.n2046 gnd.n2045 585
R3336 gnd.n2732 gnd.n2731 585
R3337 gnd.n2731 gnd.n2730 585
R3338 gnd.n2051 gnd.n2050 585
R3339 gnd.n2063 gnd.n2051 585
R3340 gnd.n2073 gnd.n2062 585
R3341 gnd.n2721 gnd.n2062 585
R3342 gnd.n2708 gnd.n2707 585
R3343 gnd.n2709 gnd.n2708 585
R3344 gnd.n2072 gnd.n2071 585
R3345 gnd.n2071 gnd.n2070 585
R3346 gnd.n2702 gnd.n2701 585
R3347 gnd.n2701 gnd.n2700 585
R3348 gnd.n2076 gnd.n2075 585
R3349 gnd.n2088 gnd.n2076 585
R3350 gnd.n2098 gnd.n2087 585
R3351 gnd.n2691 gnd.n2087 585
R3352 gnd.n2678 gnd.n2677 585
R3353 gnd.n2679 gnd.n2678 585
R3354 gnd.n2097 gnd.n2096 585
R3355 gnd.n2096 gnd.n2095 585
R3356 gnd.n2672 gnd.n2671 585
R3357 gnd.n2671 gnd.n2670 585
R3358 gnd.n2101 gnd.n2100 585
R3359 gnd.n2583 gnd.n2101 585
R3360 gnd.n6373 gnd.n440 585
R3361 gnd.n6339 gnd.n440 585
R3362 gnd.n6374 gnd.n439 585
R3363 gnd.n485 gnd.n433 585
R3364 gnd.n6381 gnd.n432 585
R3365 gnd.n6382 gnd.n431 585
R3366 gnd.n482 gnd.n423 585
R3367 gnd.n6389 gnd.n422 585
R3368 gnd.n6390 gnd.n421 585
R3369 gnd.n480 gnd.n415 585
R3370 gnd.n6397 gnd.n414 585
R3371 gnd.n6398 gnd.n413 585
R3372 gnd.n477 gnd.n405 585
R3373 gnd.n6405 gnd.n404 585
R3374 gnd.n6406 gnd.n403 585
R3375 gnd.n475 gnd.n395 585
R3376 gnd.n6413 gnd.n394 585
R3377 gnd.n6414 gnd.n393 585
R3378 gnd.n6415 gnd.n392 585
R3379 gnd.n6341 gnd.n391 585
R3380 gnd.n6343 gnd.n6342 585
R3381 gnd.n6344 gnd.n468 585
R3382 gnd.n472 gnd.n466 585
R3383 gnd.n6348 gnd.n465 585
R3384 gnd.n6349 gnd.n464 585
R3385 gnd.n6350 gnd.n460 585
R3386 gnd.n456 gnd.n452 585
R3387 gnd.n6362 gnd.n451 585
R3388 gnd.n6363 gnd.n450 585
R3389 gnd.n487 gnd.n449 585
R3390 gnd.n2809 gnd.t316 543.808
R3391 gnd.n1698 gnd.t308 543.808
R3392 gnd.n3784 gnd.t238 543.808
R3393 gnd.n1692 gnd.t234 543.808
R3394 gnd.n3542 gnd.n1648 458.866
R3395 gnd.n3422 gnd.n1645 458.866
R3396 gnd.n2874 gnd.n2808 458.866
R3397 gnd.n3847 gnd.n1448 458.866
R3398 gnd.n2189 gnd.t248 371.625
R3399 gnd.n6367 gnd.t214 371.625
R3400 gnd.n6720 gnd.t255 371.625
R3401 gnd.n6903 gnd.t268 371.625
R3402 gnd.n7002 gnd.t277 371.625
R3403 gnd.n341 gnd.t292 371.625
R3404 gnd.n364 gnd.t295 371.625
R3405 gnd.n386 gnd.t258 371.625
R3406 gnd.n6735 gnd.t204 371.625
R3407 gnd.n2194 gnd.t230 371.625
R3408 gnd.n2405 gnd.t226 371.625
R3409 gnd.n1083 gnd.t252 371.625
R3410 gnd.n1105 gnd.t274 371.625
R3411 gnd.n1127 gnd.t283 371.625
R3412 gnd.n1396 gnd.t271 371.625
R3413 gnd.n2200 gnd.t286 371.625
R3414 gnd.n2212 gnd.t305 371.625
R3415 gnd.n441 gnd.t222 371.625
R3416 gnd.n5774 gnd.n5773 348.315
R3417 gnd.n4624 gnd.t261 323.425
R3418 gnd.n4182 gnd.t319 323.425
R3419 gnd.n5472 gnd.n5446 289.615
R3420 gnd.n5440 gnd.n5414 289.615
R3421 gnd.n5408 gnd.n5382 289.615
R3422 gnd.n5377 gnd.n5351 289.615
R3423 gnd.n5345 gnd.n5319 289.615
R3424 gnd.n5313 gnd.n5287 289.615
R3425 gnd.n5281 gnd.n5255 289.615
R3426 gnd.n5250 gnd.n5224 289.615
R3427 gnd.n4698 gnd.t301 279.217
R3428 gnd.n4208 gnd.t218 279.217
R3429 gnd.n1455 gnd.t213 260.649
R3430 gnd.n1661 gnd.t244 260.649
R3431 gnd.n3849 gnd.n3848 256.663
R3432 gnd.n3849 gnd.n1414 256.663
R3433 gnd.n3849 gnd.n1415 256.663
R3434 gnd.n3849 gnd.n1416 256.663
R3435 gnd.n3849 gnd.n1417 256.663
R3436 gnd.n3849 gnd.n1418 256.663
R3437 gnd.n3849 gnd.n1419 256.663
R3438 gnd.n3849 gnd.n1420 256.663
R3439 gnd.n3849 gnd.n1421 256.663
R3440 gnd.n3849 gnd.n1422 256.663
R3441 gnd.n3849 gnd.n1423 256.663
R3442 gnd.n3849 gnd.n1424 256.663
R3443 gnd.n3849 gnd.n1425 256.663
R3444 gnd.n3849 gnd.n1426 256.663
R3445 gnd.n3849 gnd.n1427 256.663
R3446 gnd.n3849 gnd.n1428 256.663
R3447 gnd.n3852 gnd.n1411 256.663
R3448 gnd.n3850 gnd.n3849 256.663
R3449 gnd.n3849 gnd.n1429 256.663
R3450 gnd.n3849 gnd.n1430 256.663
R3451 gnd.n3849 gnd.n1431 256.663
R3452 gnd.n3849 gnd.n1432 256.663
R3453 gnd.n3849 gnd.n1433 256.663
R3454 gnd.n3849 gnd.n1434 256.663
R3455 gnd.n3849 gnd.n1435 256.663
R3456 gnd.n3849 gnd.n1436 256.663
R3457 gnd.n3849 gnd.n1437 256.663
R3458 gnd.n3849 gnd.n1438 256.663
R3459 gnd.n3849 gnd.n1439 256.663
R3460 gnd.n3849 gnd.n1440 256.663
R3461 gnd.n3849 gnd.n1441 256.663
R3462 gnd.n3849 gnd.n1442 256.663
R3463 gnd.n3849 gnd.n1443 256.663
R3464 gnd.n3849 gnd.n1444 256.663
R3465 gnd.n3421 gnd.n1672 256.663
R3466 gnd.n3427 gnd.n1672 256.663
R3467 gnd.n1719 gnd.n1672 256.663
R3468 gnd.n3434 gnd.n1672 256.663
R3469 gnd.n1716 gnd.n1672 256.663
R3470 gnd.n3441 gnd.n1672 256.663
R3471 gnd.n1713 gnd.n1672 256.663
R3472 gnd.n3448 gnd.n1672 256.663
R3473 gnd.n1710 gnd.n1672 256.663
R3474 gnd.n3455 gnd.n1672 256.663
R3475 gnd.n1707 gnd.n1672 256.663
R3476 gnd.n3462 gnd.n1672 256.663
R3477 gnd.n1704 gnd.n1672 256.663
R3478 gnd.n3469 gnd.n1672 256.663
R3479 gnd.n1701 gnd.n1672 256.663
R3480 gnd.n3477 gnd.n1672 256.663
R3481 gnd.n3480 gnd.n351 256.663
R3482 gnd.n3481 gnd.n1672 256.663
R3483 gnd.n3485 gnd.n1672 256.663
R3484 gnd.n1695 gnd.n1672 256.663
R3485 gnd.n3493 gnd.n1672 256.663
R3486 gnd.n1690 gnd.n1672 256.663
R3487 gnd.n3500 gnd.n1672 256.663
R3488 gnd.n1687 gnd.n1672 256.663
R3489 gnd.n3507 gnd.n1672 256.663
R3490 gnd.n1684 gnd.n1672 256.663
R3491 gnd.n3514 gnd.n1672 256.663
R3492 gnd.n1681 gnd.n1672 256.663
R3493 gnd.n3521 gnd.n1672 256.663
R3494 gnd.n1678 gnd.n1672 256.663
R3495 gnd.n3528 gnd.n1672 256.663
R3496 gnd.n1675 gnd.n1672 256.663
R3497 gnd.n3535 gnd.n1672 256.663
R3498 gnd.n1672 gnd.n1670 256.663
R3499 gnd.n4157 gnd.n1051 242.672
R3500 gnd.n4157 gnd.n1052 242.672
R3501 gnd.n4157 gnd.n1053 242.672
R3502 gnd.n4157 gnd.n1054 242.672
R3503 gnd.n4157 gnd.n1055 242.672
R3504 gnd.n4157 gnd.n1056 242.672
R3505 gnd.n4157 gnd.n1057 242.672
R3506 gnd.n4157 gnd.n1058 242.672
R3507 gnd.n4157 gnd.n1059 242.672
R3508 gnd.n3903 gnd.n1349 242.672
R3509 gnd.n3903 gnd.n1348 242.672
R3510 gnd.n3903 gnd.n1347 242.672
R3511 gnd.n3903 gnd.n1346 242.672
R3512 gnd.n3903 gnd.n1345 242.672
R3513 gnd.n3903 gnd.n1344 242.672
R3514 gnd.n3903 gnd.n1343 242.672
R3515 gnd.n3903 gnd.n1342 242.672
R3516 gnd.n3903 gnd.n1341 242.672
R3517 gnd.n4752 gnd.n4751 242.672
R3518 gnd.n4752 gnd.n4662 242.672
R3519 gnd.n4752 gnd.n4663 242.672
R3520 gnd.n4752 gnd.n4664 242.672
R3521 gnd.n4752 gnd.n4665 242.672
R3522 gnd.n4752 gnd.n4666 242.672
R3523 gnd.n4752 gnd.n4667 242.672
R3524 gnd.n4752 gnd.n4668 242.672
R3525 gnd.n4752 gnd.n4669 242.672
R3526 gnd.n4752 gnd.n4670 242.672
R3527 gnd.n4752 gnd.n4671 242.672
R3528 gnd.n4752 gnd.n4672 242.672
R3529 gnd.n4753 gnd.n4752 242.672
R3530 gnd.n5604 gnd.n1022 242.672
R3531 gnd.n5604 gnd.n1021 242.672
R3532 gnd.n5604 gnd.n1020 242.672
R3533 gnd.n5604 gnd.n1019 242.672
R3534 gnd.n5604 gnd.n1018 242.672
R3535 gnd.n5604 gnd.n1017 242.672
R3536 gnd.n5604 gnd.n1016 242.672
R3537 gnd.n5604 gnd.n1015 242.672
R3538 gnd.n5604 gnd.n1014 242.672
R3539 gnd.n5604 gnd.n1013 242.672
R3540 gnd.n5604 gnd.n1012 242.672
R3541 gnd.n5604 gnd.n1011 242.672
R3542 gnd.n5604 gnd.n1010 242.672
R3543 gnd.n6530 gnd.n313 242.672
R3544 gnd.n6530 gnd.n314 242.672
R3545 gnd.n6530 gnd.n315 242.672
R3546 gnd.n6530 gnd.n316 242.672
R3547 gnd.n6530 gnd.n317 242.672
R3548 gnd.n6530 gnd.n318 242.672
R3549 gnd.n6530 gnd.n319 242.672
R3550 gnd.n6530 gnd.n320 242.672
R3551 gnd.n6530 gnd.n321 242.672
R3552 gnd.n7042 gnd.n6836 242.672
R3553 gnd.n7042 gnd.n6732 242.672
R3554 gnd.n7042 gnd.n6731 242.672
R3555 gnd.n7042 gnd.n6730 242.672
R3556 gnd.n7042 gnd.n6729 242.672
R3557 gnd.n7042 gnd.n6728 242.672
R3558 gnd.n7042 gnd.n6727 242.672
R3559 gnd.n7042 gnd.n6726 242.672
R3560 gnd.n7042 gnd.n6725 242.672
R3561 gnd.n4836 gnd.n4835 242.672
R3562 gnd.n4835 gnd.n4574 242.672
R3563 gnd.n4835 gnd.n4575 242.672
R3564 gnd.n4835 gnd.n4576 242.672
R3565 gnd.n4835 gnd.n4577 242.672
R3566 gnd.n4835 gnd.n4578 242.672
R3567 gnd.n4835 gnd.n4579 242.672
R3568 gnd.n4835 gnd.n4580 242.672
R3569 gnd.n5604 gnd.n4158 242.672
R3570 gnd.n5604 gnd.n4159 242.672
R3571 gnd.n5604 gnd.n4160 242.672
R3572 gnd.n5604 gnd.n4161 242.672
R3573 gnd.n5604 gnd.n4162 242.672
R3574 gnd.n5604 gnd.n4163 242.672
R3575 gnd.n5604 gnd.n4164 242.672
R3576 gnd.n5604 gnd.n4165 242.672
R3577 gnd.n4157 gnd.n4156 242.672
R3578 gnd.n4157 gnd.n1023 242.672
R3579 gnd.n4157 gnd.n1024 242.672
R3580 gnd.n4157 gnd.n1025 242.672
R3581 gnd.n4157 gnd.n1026 242.672
R3582 gnd.n4157 gnd.n1027 242.672
R3583 gnd.n4157 gnd.n1028 242.672
R3584 gnd.n4157 gnd.n1029 242.672
R3585 gnd.n4157 gnd.n1030 242.672
R3586 gnd.n4157 gnd.n1031 242.672
R3587 gnd.n4157 gnd.n1032 242.672
R3588 gnd.n4157 gnd.n1033 242.672
R3589 gnd.n4157 gnd.n1034 242.672
R3590 gnd.n4157 gnd.n1035 242.672
R3591 gnd.n4157 gnd.n1036 242.672
R3592 gnd.n4157 gnd.n1037 242.672
R3593 gnd.n4157 gnd.n1038 242.672
R3594 gnd.n4157 gnd.n1039 242.672
R3595 gnd.n4157 gnd.n1040 242.672
R3596 gnd.n4157 gnd.n1041 242.672
R3597 gnd.n4157 gnd.n1042 242.672
R3598 gnd.n4157 gnd.n1043 242.672
R3599 gnd.n4157 gnd.n1044 242.672
R3600 gnd.n4157 gnd.n1045 242.672
R3601 gnd.n4157 gnd.n1046 242.672
R3602 gnd.n4157 gnd.n1047 242.672
R3603 gnd.n4157 gnd.n1048 242.672
R3604 gnd.n4157 gnd.n1049 242.672
R3605 gnd.n4157 gnd.n1050 242.672
R3606 gnd.n3903 gnd.n1351 242.672
R3607 gnd.n3903 gnd.n1352 242.672
R3608 gnd.n3903 gnd.n1353 242.672
R3609 gnd.n3903 gnd.n1354 242.672
R3610 gnd.n3903 gnd.n1355 242.672
R3611 gnd.n3903 gnd.n1356 242.672
R3612 gnd.n3903 gnd.n1357 242.672
R3613 gnd.n3903 gnd.n1358 242.672
R3614 gnd.n3903 gnd.n1359 242.672
R3615 gnd.n3903 gnd.n1360 242.672
R3616 gnd.n3903 gnd.n1361 242.672
R3617 gnd.n3903 gnd.n1362 242.672
R3618 gnd.n3903 gnd.n1363 242.672
R3619 gnd.n3903 gnd.n1364 242.672
R3620 gnd.n3903 gnd.n1365 242.672
R3621 gnd.n3903 gnd.n1366 242.672
R3622 gnd.n3853 gnd.n1407 242.672
R3623 gnd.n3903 gnd.n1367 242.672
R3624 gnd.n3903 gnd.n1368 242.672
R3625 gnd.n3903 gnd.n1369 242.672
R3626 gnd.n3903 gnd.n1370 242.672
R3627 gnd.n3903 gnd.n1371 242.672
R3628 gnd.n3903 gnd.n1372 242.672
R3629 gnd.n3903 gnd.n1373 242.672
R3630 gnd.n3903 gnd.n1374 242.672
R3631 gnd.n3903 gnd.n1375 242.672
R3632 gnd.n3903 gnd.n1376 242.672
R3633 gnd.n3903 gnd.n1377 242.672
R3634 gnd.n3903 gnd.n1378 242.672
R3635 gnd.n3903 gnd.n3902 242.672
R3636 gnd.n6531 gnd.n6530 242.672
R3637 gnd.n6530 gnd.n285 242.672
R3638 gnd.n6530 gnd.n286 242.672
R3639 gnd.n6530 gnd.n287 242.672
R3640 gnd.n6530 gnd.n288 242.672
R3641 gnd.n6530 gnd.n289 242.672
R3642 gnd.n6530 gnd.n290 242.672
R3643 gnd.n6530 gnd.n291 242.672
R3644 gnd.n6530 gnd.n292 242.672
R3645 gnd.n6530 gnd.n293 242.672
R3646 gnd.n6530 gnd.n294 242.672
R3647 gnd.n6530 gnd.n295 242.672
R3648 gnd.n6530 gnd.n296 242.672
R3649 gnd.n6481 gnd.n352 242.672
R3650 gnd.n6530 gnd.n297 242.672
R3651 gnd.n6530 gnd.n298 242.672
R3652 gnd.n6530 gnd.n299 242.672
R3653 gnd.n6530 gnd.n300 242.672
R3654 gnd.n6530 gnd.n301 242.672
R3655 gnd.n6530 gnd.n302 242.672
R3656 gnd.n6530 gnd.n303 242.672
R3657 gnd.n6530 gnd.n304 242.672
R3658 gnd.n6530 gnd.n305 242.672
R3659 gnd.n6530 gnd.n306 242.672
R3660 gnd.n6530 gnd.n307 242.672
R3661 gnd.n6530 gnd.n308 242.672
R3662 gnd.n6530 gnd.n309 242.672
R3663 gnd.n6530 gnd.n310 242.672
R3664 gnd.n6530 gnd.n311 242.672
R3665 gnd.n6530 gnd.n312 242.672
R3666 gnd.n7043 gnd.n7042 242.672
R3667 gnd.n7042 gnd.n6837 242.672
R3668 gnd.n7042 gnd.n6838 242.672
R3669 gnd.n7042 gnd.n6839 242.672
R3670 gnd.n7042 gnd.n6840 242.672
R3671 gnd.n7042 gnd.n6841 242.672
R3672 gnd.n7042 gnd.n6842 242.672
R3673 gnd.n7042 gnd.n6843 242.672
R3674 gnd.n7042 gnd.n6844 242.672
R3675 gnd.n7042 gnd.n6845 242.672
R3676 gnd.n7042 gnd.n6846 242.672
R3677 gnd.n7042 gnd.n6847 242.672
R3678 gnd.n7042 gnd.n6848 242.672
R3679 gnd.n7042 gnd.n6849 242.672
R3680 gnd.n7042 gnd.n6850 242.672
R3681 gnd.n7042 gnd.n6851 242.672
R3682 gnd.n7042 gnd.n6852 242.672
R3683 gnd.n7042 gnd.n6853 242.672
R3684 gnd.n7042 gnd.n6854 242.672
R3685 gnd.n7042 gnd.n6855 242.672
R3686 gnd.n7042 gnd.n6856 242.672
R3687 gnd.n7042 gnd.n6857 242.672
R3688 gnd.n7042 gnd.n6858 242.672
R3689 gnd.n7042 gnd.n6859 242.672
R3690 gnd.n7042 gnd.n6860 242.672
R3691 gnd.n7042 gnd.n6861 242.672
R3692 gnd.n7042 gnd.n6862 242.672
R3693 gnd.n7042 gnd.n6863 242.672
R3694 gnd.n7042 gnd.n6864 242.672
R3695 gnd.n2661 gnd.n2660 242.672
R3696 gnd.n2660 gnd.n2112 242.672
R3697 gnd.n2660 gnd.n2113 242.672
R3698 gnd.n2660 gnd.n2114 242.672
R3699 gnd.n2660 gnd.n2115 242.672
R3700 gnd.n2660 gnd.n2116 242.672
R3701 gnd.n2660 gnd.n2117 242.672
R3702 gnd.n2660 gnd.n2118 242.672
R3703 gnd.n2660 gnd.n2119 242.672
R3704 gnd.n2660 gnd.n2120 242.672
R3705 gnd.n2660 gnd.n2121 242.672
R3706 gnd.n2660 gnd.n2122 242.672
R3707 gnd.n2660 gnd.n2123 242.672
R3708 gnd.n2660 gnd.n2124 242.672
R3709 gnd.n6339 gnd.n486 242.672
R3710 gnd.n6339 gnd.n484 242.672
R3711 gnd.n6339 gnd.n483 242.672
R3712 gnd.n6339 gnd.n481 242.672
R3713 gnd.n6339 gnd.n479 242.672
R3714 gnd.n6339 gnd.n478 242.672
R3715 gnd.n6339 gnd.n476 242.672
R3716 gnd.n6339 gnd.n474 242.672
R3717 gnd.n6340 gnd.n6339 242.672
R3718 gnd.n6339 gnd.n469 242.672
R3719 gnd.n6339 gnd.n473 242.672
R3720 gnd.n6339 gnd.n471 242.672
R3721 gnd.n6339 gnd.n489 242.672
R3722 gnd.n6339 gnd.n488 242.672
R3723 gnd.n7041 gnd.n6865 240.244
R3724 gnd.n7034 gnd.n7033 240.244
R3725 gnd.n7031 gnd.n7030 240.244
R3726 gnd.n7027 gnd.n7026 240.244
R3727 gnd.n7023 gnd.n7022 240.244
R3728 gnd.n7019 gnd.n7018 240.244
R3729 gnd.n7015 gnd.n7014 240.244
R3730 gnd.n7011 gnd.n7010 240.244
R3731 gnd.n7007 gnd.n7006 240.244
R3732 gnd.n7000 gnd.n6999 240.244
R3733 gnd.n6996 gnd.n6995 240.244
R3734 gnd.n6992 gnd.n6991 240.244
R3735 gnd.n6988 gnd.n6987 240.244
R3736 gnd.n6984 gnd.n6983 240.244
R3737 gnd.n6980 gnd.n6979 240.244
R3738 gnd.n6976 gnd.n6975 240.244
R3739 gnd.n6972 gnd.n6971 240.244
R3740 gnd.n6968 gnd.n6967 240.244
R3741 gnd.n6964 gnd.n6963 240.244
R3742 gnd.n6957 gnd.n6956 240.244
R3743 gnd.n6954 gnd.n6953 240.244
R3744 gnd.n6950 gnd.n6949 240.244
R3745 gnd.n6946 gnd.n6945 240.244
R3746 gnd.n6942 gnd.n6941 240.244
R3747 gnd.n6938 gnd.n6937 240.244
R3748 gnd.n6934 gnd.n6933 240.244
R3749 gnd.n6930 gnd.n6929 240.244
R3750 gnd.n6926 gnd.n6925 240.244
R3751 gnd.n6922 gnd.n6723 240.244
R3752 gnd.n501 gnd.n275 240.244
R3753 gnd.n275 gnd.n266 240.244
R3754 gnd.n6550 gnd.n266 240.244
R3755 gnd.n6550 gnd.n256 240.244
R3756 gnd.n6554 gnd.n256 240.244
R3757 gnd.n6554 gnd.n247 240.244
R3758 gnd.n247 gnd.n238 240.244
R3759 gnd.n6595 gnd.n238 240.244
R3760 gnd.n6595 gnd.n230 240.244
R3761 gnd.n230 gnd.n220 240.244
R3762 gnd.n6614 gnd.n220 240.244
R3763 gnd.n6615 gnd.n6614 240.244
R3764 gnd.n6615 gnd.n210 240.244
R3765 gnd.n6618 gnd.n210 240.244
R3766 gnd.n6618 gnd.n201 240.244
R3767 gnd.n201 gnd.n193 240.244
R3768 gnd.n6653 gnd.n193 240.244
R3769 gnd.n6653 gnd.n186 240.244
R3770 gnd.n6655 gnd.n186 240.244
R3771 gnd.n6655 gnd.n177 240.244
R3772 gnd.n177 gnd.n172 240.244
R3773 gnd.n6679 gnd.n172 240.244
R3774 gnd.n6679 gnd.n73 240.244
R3775 gnd.n6686 gnd.n73 240.244
R3776 gnd.n6686 gnd.n84 240.244
R3777 gnd.n6689 gnd.n84 240.244
R3778 gnd.n6689 gnd.n95 240.244
R3779 gnd.n6693 gnd.n95 240.244
R3780 gnd.n6693 gnd.n105 240.244
R3781 gnd.n6696 gnd.n105 240.244
R3782 gnd.n6696 gnd.n114 240.244
R3783 gnd.n6700 gnd.n114 240.244
R3784 gnd.n6700 gnd.n124 240.244
R3785 gnd.n6703 gnd.n124 240.244
R3786 gnd.n6703 gnd.n133 240.244
R3787 gnd.n6707 gnd.n133 240.244
R3788 gnd.n6707 gnd.n143 240.244
R3789 gnd.n6710 gnd.n143 240.244
R3790 gnd.n6710 gnd.n152 240.244
R3791 gnd.n6714 gnd.n152 240.244
R3792 gnd.n6714 gnd.n162 240.244
R3793 gnd.n7044 gnd.n162 240.244
R3794 gnd.n6529 gnd.n283 240.244
R3795 gnd.n6529 gnd.n324 240.244
R3796 gnd.n6525 gnd.n6524 240.244
R3797 gnd.n6521 gnd.n6520 240.244
R3798 gnd.n6517 gnd.n6516 240.244
R3799 gnd.n6513 gnd.n6512 240.244
R3800 gnd.n6509 gnd.n6508 240.244
R3801 gnd.n6505 gnd.n6504 240.244
R3802 gnd.n6501 gnd.n6500 240.244
R3803 gnd.n6496 gnd.n6495 240.244
R3804 gnd.n6492 gnd.n6491 240.244
R3805 gnd.n6488 gnd.n6487 240.244
R3806 gnd.n6484 gnd.n6483 240.244
R3807 gnd.n6479 gnd.n6478 240.244
R3808 gnd.n6475 gnd.n6474 240.244
R3809 gnd.n6471 gnd.n6470 240.244
R3810 gnd.n6467 gnd.n6466 240.244
R3811 gnd.n6463 gnd.n6462 240.244
R3812 gnd.n6459 gnd.n6458 240.244
R3813 gnd.n6455 gnd.n6454 240.244
R3814 gnd.n6451 gnd.n6450 240.244
R3815 gnd.n6447 gnd.n6446 240.244
R3816 gnd.n6443 gnd.n6442 240.244
R3817 gnd.n6439 gnd.n6438 240.244
R3818 gnd.n6435 gnd.n6434 240.244
R3819 gnd.n6431 gnd.n6430 240.244
R3820 gnd.n6427 gnd.n6426 240.244
R3821 gnd.n6423 gnd.n6422 240.244
R3822 gnd.n6539 gnd.n277 240.244
R3823 gnd.n6539 gnd.n278 240.244
R3824 gnd.n278 gnd.n254 240.244
R3825 gnd.n6566 gnd.n254 240.244
R3826 gnd.n6566 gnd.n249 240.244
R3827 gnd.n6574 gnd.n249 240.244
R3828 gnd.n6574 gnd.n250 240.244
R3829 gnd.n250 gnd.n228 240.244
R3830 gnd.n6606 gnd.n228 240.244
R3831 gnd.n6606 gnd.n224 240.244
R3832 gnd.n6612 gnd.n224 240.244
R3833 gnd.n6612 gnd.n208 240.244
R3834 gnd.n6630 gnd.n208 240.244
R3835 gnd.n6630 gnd.n203 240.244
R3836 gnd.n6638 gnd.n203 240.244
R3837 gnd.n6638 gnd.n204 240.244
R3838 gnd.n204 gnd.n185 240.244
R3839 gnd.n6662 gnd.n185 240.244
R3840 gnd.n6662 gnd.n180 240.244
R3841 gnd.n6671 gnd.n180 240.244
R3842 gnd.n6671 gnd.n181 240.244
R3843 gnd.n181 gnd.n76 240.244
R3844 gnd.n7106 gnd.n76 240.244
R3845 gnd.n7106 gnd.n77 240.244
R3846 gnd.n7102 gnd.n77 240.244
R3847 gnd.n7102 gnd.n83 240.244
R3848 gnd.n7094 gnd.n83 240.244
R3849 gnd.n7094 gnd.n97 240.244
R3850 gnd.n7090 gnd.n97 240.244
R3851 gnd.n7090 gnd.n103 240.244
R3852 gnd.n7082 gnd.n103 240.244
R3853 gnd.n7082 gnd.n117 240.244
R3854 gnd.n7078 gnd.n117 240.244
R3855 gnd.n7078 gnd.n123 240.244
R3856 gnd.n7070 gnd.n123 240.244
R3857 gnd.n7070 gnd.n135 240.244
R3858 gnd.n7066 gnd.n135 240.244
R3859 gnd.n7066 gnd.n141 240.244
R3860 gnd.n7058 gnd.n141 240.244
R3861 gnd.n7058 gnd.n155 240.244
R3862 gnd.n7054 gnd.n155 240.244
R3863 gnd.n7054 gnd.n161 240.244
R3864 gnd.n3904 gnd.n1338 240.244
R3865 gnd.n3901 gnd.n1379 240.244
R3866 gnd.n3897 gnd.n3896 240.244
R3867 gnd.n3893 gnd.n3892 240.244
R3868 gnd.n3889 gnd.n3888 240.244
R3869 gnd.n3885 gnd.n3884 240.244
R3870 gnd.n3881 gnd.n3880 240.244
R3871 gnd.n3877 gnd.n3876 240.244
R3872 gnd.n3873 gnd.n3872 240.244
R3873 gnd.n3868 gnd.n3867 240.244
R3874 gnd.n3864 gnd.n3863 240.244
R3875 gnd.n3860 gnd.n3859 240.244
R3876 gnd.n3856 gnd.n3855 240.244
R3877 gnd.n2219 gnd.n2218 240.244
R3878 gnd.n2226 gnd.n2225 240.244
R3879 gnd.n2229 gnd.n2228 240.244
R3880 gnd.n2236 gnd.n2235 240.244
R3881 gnd.n2239 gnd.n2238 240.244
R3882 gnd.n2246 gnd.n2245 240.244
R3883 gnd.n2249 gnd.n2248 240.244
R3884 gnd.n2256 gnd.n2255 240.244
R3885 gnd.n2259 gnd.n2258 240.244
R3886 gnd.n2266 gnd.n2265 240.244
R3887 gnd.n2269 gnd.n2268 240.244
R3888 gnd.n2276 gnd.n2275 240.244
R3889 gnd.n2279 gnd.n2278 240.244
R3890 gnd.n2286 gnd.n2285 240.244
R3891 gnd.n2289 gnd.n2288 240.244
R3892 gnd.n1137 gnd.n1136 240.244
R3893 gnd.n2323 gnd.n1137 240.244
R3894 gnd.n2323 gnd.n1147 240.244
R3895 gnd.n2326 gnd.n1147 240.244
R3896 gnd.n2326 gnd.n1157 240.244
R3897 gnd.n2330 gnd.n1157 240.244
R3898 gnd.n2330 gnd.n1166 240.244
R3899 gnd.n2333 gnd.n1166 240.244
R3900 gnd.n2333 gnd.n1175 240.244
R3901 gnd.n2337 gnd.n1175 240.244
R3902 gnd.n2337 gnd.n1185 240.244
R3903 gnd.n2340 gnd.n1185 240.244
R3904 gnd.n2340 gnd.n1194 240.244
R3905 gnd.n2344 gnd.n1194 240.244
R3906 gnd.n2344 gnd.n1204 240.244
R3907 gnd.n2347 gnd.n1204 240.244
R3908 gnd.n2347 gnd.n1213 240.244
R3909 gnd.n2351 gnd.n1213 240.244
R3910 gnd.n2351 gnd.n1223 240.244
R3911 gnd.n2354 gnd.n1223 240.244
R3912 gnd.n2354 gnd.n1232 240.244
R3913 gnd.n2358 gnd.n1232 240.244
R3914 gnd.n2358 gnd.n1242 240.244
R3915 gnd.n2361 gnd.n1242 240.244
R3916 gnd.n2361 gnd.n1251 240.244
R3917 gnd.n2365 gnd.n1251 240.244
R3918 gnd.n2365 gnd.n1261 240.244
R3919 gnd.n2368 gnd.n1261 240.244
R3920 gnd.n2368 gnd.n1270 240.244
R3921 gnd.n2372 gnd.n1270 240.244
R3922 gnd.n2372 gnd.n1280 240.244
R3923 gnd.n2375 gnd.n1280 240.244
R3924 gnd.n2375 gnd.n1289 240.244
R3925 gnd.n2379 gnd.n1289 240.244
R3926 gnd.n2379 gnd.n1300 240.244
R3927 gnd.n2532 gnd.n1300 240.244
R3928 gnd.n2532 gnd.n1310 240.244
R3929 gnd.n2542 gnd.n1310 240.244
R3930 gnd.n2542 gnd.n1321 240.244
R3931 gnd.n2316 gnd.n1321 240.244
R3932 gnd.n2316 gnd.n1330 240.244
R3933 gnd.n2296 gnd.n1330 240.244
R3934 gnd.n1063 gnd.n1062 240.244
R3935 gnd.n4150 gnd.n1062 240.244
R3936 gnd.n4148 gnd.n4147 240.244
R3937 gnd.n4144 gnd.n4143 240.244
R3938 gnd.n4140 gnd.n4139 240.244
R3939 gnd.n4136 gnd.n4135 240.244
R3940 gnd.n4132 gnd.n4131 240.244
R3941 gnd.n4128 gnd.n4127 240.244
R3942 gnd.n4124 gnd.n4123 240.244
R3943 gnd.n4119 gnd.n4118 240.244
R3944 gnd.n4115 gnd.n4114 240.244
R3945 gnd.n4111 gnd.n4110 240.244
R3946 gnd.n4107 gnd.n4106 240.244
R3947 gnd.n4103 gnd.n4102 240.244
R3948 gnd.n4099 gnd.n4098 240.244
R3949 gnd.n4095 gnd.n4094 240.244
R3950 gnd.n4091 gnd.n4090 240.244
R3951 gnd.n4087 gnd.n4086 240.244
R3952 gnd.n4083 gnd.n4082 240.244
R3953 gnd.n4079 gnd.n4078 240.244
R3954 gnd.n4075 gnd.n4074 240.244
R3955 gnd.n4071 gnd.n4070 240.244
R3956 gnd.n4067 gnd.n4066 240.244
R3957 gnd.n4063 gnd.n4062 240.244
R3958 gnd.n4059 gnd.n4058 240.244
R3959 gnd.n4055 gnd.n4054 240.244
R3960 gnd.n4051 gnd.n4050 240.244
R3961 gnd.n4047 gnd.n4046 240.244
R3962 gnd.n4043 gnd.n4042 240.244
R3963 gnd.n4032 gnd.n1064 240.244
R3964 gnd.n4032 gnd.n1139 240.244
R3965 gnd.n4026 gnd.n1139 240.244
R3966 gnd.n4026 gnd.n1145 240.244
R3967 gnd.n4018 gnd.n1145 240.244
R3968 gnd.n4018 gnd.n1160 240.244
R3969 gnd.n4014 gnd.n1160 240.244
R3970 gnd.n4014 gnd.n1165 240.244
R3971 gnd.n4006 gnd.n1165 240.244
R3972 gnd.n4006 gnd.n1177 240.244
R3973 gnd.n4002 gnd.n1177 240.244
R3974 gnd.n4002 gnd.n1183 240.244
R3975 gnd.n3994 gnd.n1183 240.244
R3976 gnd.n3994 gnd.n1197 240.244
R3977 gnd.n3990 gnd.n1197 240.244
R3978 gnd.n3990 gnd.n1203 240.244
R3979 gnd.n3982 gnd.n1203 240.244
R3980 gnd.n3982 gnd.n1215 240.244
R3981 gnd.n3978 gnd.n1215 240.244
R3982 gnd.n3978 gnd.n1221 240.244
R3983 gnd.n3970 gnd.n1221 240.244
R3984 gnd.n3970 gnd.n1235 240.244
R3985 gnd.n3966 gnd.n1235 240.244
R3986 gnd.n3966 gnd.n1241 240.244
R3987 gnd.n3958 gnd.n1241 240.244
R3988 gnd.n3958 gnd.n1254 240.244
R3989 gnd.n3954 gnd.n1254 240.244
R3990 gnd.n3954 gnd.n1260 240.244
R3991 gnd.n3946 gnd.n1260 240.244
R3992 gnd.n3946 gnd.n1273 240.244
R3993 gnd.n3942 gnd.n1273 240.244
R3994 gnd.n3942 gnd.n1279 240.244
R3995 gnd.n3934 gnd.n1279 240.244
R3996 gnd.n3934 gnd.n1292 240.244
R3997 gnd.n3930 gnd.n1292 240.244
R3998 gnd.n3930 gnd.n1298 240.244
R3999 gnd.n3922 gnd.n1298 240.244
R4000 gnd.n3922 gnd.n1313 240.244
R4001 gnd.n3918 gnd.n1313 240.244
R4002 gnd.n3918 gnd.n1319 240.244
R4003 gnd.n3910 gnd.n1319 240.244
R4004 gnd.n3910 gnd.n1333 240.244
R4005 gnd.n5603 gnd.n4167 240.244
R4006 gnd.n5596 gnd.n5595 240.244
R4007 gnd.n5593 gnd.n5592 240.244
R4008 gnd.n5589 gnd.n5588 240.244
R4009 gnd.n5585 gnd.n5584 240.244
R4010 gnd.n5581 gnd.n5580 240.244
R4011 gnd.n5577 gnd.n5576 240.244
R4012 gnd.n5573 gnd.n5572 240.244
R4013 gnd.n4847 gnd.n4559 240.244
R4014 gnd.n4857 gnd.n4559 240.244
R4015 gnd.n4857 gnd.n4550 240.244
R4016 gnd.n4550 gnd.n4539 240.244
R4017 gnd.n4878 gnd.n4539 240.244
R4018 gnd.n4878 gnd.n4533 240.244
R4019 gnd.n4888 gnd.n4533 240.244
R4020 gnd.n4888 gnd.n4522 240.244
R4021 gnd.n4522 gnd.n4514 240.244
R4022 gnd.n4906 gnd.n4514 240.244
R4023 gnd.n4907 gnd.n4906 240.244
R4024 gnd.n4907 gnd.n4499 240.244
R4025 gnd.n4909 gnd.n4499 240.244
R4026 gnd.n4909 gnd.n4485 240.244
R4027 gnd.n4951 gnd.n4485 240.244
R4028 gnd.n4952 gnd.n4951 240.244
R4029 gnd.n4955 gnd.n4952 240.244
R4030 gnd.n4955 gnd.n4440 240.244
R4031 gnd.n4480 gnd.n4440 240.244
R4032 gnd.n4480 gnd.n4450 240.244
R4033 gnd.n4965 gnd.n4450 240.244
R4034 gnd.n4965 gnd.n4471 240.244
R4035 gnd.n4975 gnd.n4471 240.244
R4036 gnd.n4975 gnd.n4369 240.244
R4037 gnd.n5020 gnd.n4369 240.244
R4038 gnd.n5020 gnd.n4355 240.244
R4039 gnd.n5042 gnd.n4355 240.244
R4040 gnd.n5043 gnd.n5042 240.244
R4041 gnd.n5043 gnd.n4342 240.244
R4042 gnd.n4342 gnd.n4331 240.244
R4043 gnd.n5074 gnd.n4331 240.244
R4044 gnd.n5075 gnd.n5074 240.244
R4045 gnd.n5076 gnd.n5075 240.244
R4046 gnd.n5076 gnd.n4316 240.244
R4047 gnd.n4316 gnd.n4315 240.244
R4048 gnd.n4315 gnd.n4300 240.244
R4049 gnd.n5127 gnd.n4300 240.244
R4050 gnd.n5128 gnd.n5127 240.244
R4051 gnd.n5128 gnd.n4287 240.244
R4052 gnd.n4287 gnd.n4276 240.244
R4053 gnd.n5159 gnd.n4276 240.244
R4054 gnd.n5160 gnd.n5159 240.244
R4055 gnd.n5161 gnd.n5160 240.244
R4056 gnd.n5161 gnd.n4260 240.244
R4057 gnd.n4260 gnd.n4259 240.244
R4058 gnd.n4259 gnd.n4246 240.244
R4059 gnd.n5216 gnd.n4246 240.244
R4060 gnd.n5217 gnd.n5216 240.244
R4061 gnd.n5217 gnd.n4233 240.244
R4062 gnd.n4233 gnd.n4223 240.244
R4063 gnd.n5504 gnd.n4223 240.244
R4064 gnd.n5507 gnd.n5504 240.244
R4065 gnd.n5507 gnd.n5506 240.244
R4066 gnd.n4837 gnd.n4572 240.244
R4067 gnd.n4593 gnd.n4572 240.244
R4068 gnd.n4596 gnd.n4595 240.244
R4069 gnd.n4603 gnd.n4602 240.244
R4070 gnd.n4606 gnd.n4605 240.244
R4071 gnd.n4613 gnd.n4612 240.244
R4072 gnd.n4616 gnd.n4615 240.244
R4073 gnd.n4623 gnd.n4622 240.244
R4074 gnd.n4845 gnd.n4569 240.244
R4075 gnd.n4569 gnd.n4548 240.244
R4076 gnd.n4868 gnd.n4548 240.244
R4077 gnd.n4868 gnd.n4542 240.244
R4078 gnd.n4876 gnd.n4542 240.244
R4079 gnd.n4876 gnd.n4544 240.244
R4080 gnd.n4544 gnd.n4520 240.244
R4081 gnd.n4898 gnd.n4520 240.244
R4082 gnd.n4898 gnd.n4516 240.244
R4083 gnd.n4904 gnd.n4516 240.244
R4084 gnd.n4904 gnd.n4498 240.244
R4085 gnd.n4929 gnd.n4498 240.244
R4086 gnd.n4929 gnd.n4493 240.244
R4087 gnd.n4941 gnd.n4493 240.244
R4088 gnd.n4941 gnd.n4494 240.244
R4089 gnd.n4937 gnd.n4494 240.244
R4090 gnd.n4937 gnd.n4442 240.244
R4091 gnd.n4989 gnd.n4442 240.244
R4092 gnd.n4989 gnd.n4443 240.244
R4093 gnd.n4985 gnd.n4443 240.244
R4094 gnd.n4985 gnd.n4449 240.244
R4095 gnd.n4469 gnd.n4449 240.244
R4096 gnd.n4469 gnd.n4367 240.244
R4097 gnd.n5024 gnd.n4367 240.244
R4098 gnd.n5024 gnd.n4362 240.244
R4099 gnd.n5032 gnd.n4362 240.244
R4100 gnd.n5032 gnd.n4363 240.244
R4101 gnd.n4363 gnd.n4340 240.244
R4102 gnd.n5064 gnd.n4340 240.244
R4103 gnd.n5064 gnd.n4335 240.244
R4104 gnd.n5072 gnd.n4335 240.244
R4105 gnd.n5072 gnd.n4336 240.244
R4106 gnd.n4336 gnd.n4313 240.244
R4107 gnd.n5109 gnd.n4313 240.244
R4108 gnd.n5109 gnd.n4308 240.244
R4109 gnd.n5117 gnd.n4308 240.244
R4110 gnd.n5117 gnd.n4309 240.244
R4111 gnd.n4309 gnd.n4285 240.244
R4112 gnd.n5149 gnd.n4285 240.244
R4113 gnd.n5149 gnd.n4280 240.244
R4114 gnd.n5157 gnd.n4280 240.244
R4115 gnd.n5157 gnd.n4281 240.244
R4116 gnd.n4281 gnd.n4258 240.244
R4117 gnd.n5198 gnd.n4258 240.244
R4118 gnd.n5198 gnd.n4253 240.244
R4119 gnd.n5206 gnd.n4253 240.244
R4120 gnd.n5206 gnd.n4254 240.244
R4121 gnd.n4254 gnd.n4231 240.244
R4122 gnd.n5492 gnd.n4231 240.244
R4123 gnd.n5492 gnd.n4226 240.244
R4124 gnd.n5502 gnd.n4226 240.244
R4125 gnd.n5502 gnd.n4227 240.244
R4126 gnd.n4227 gnd.n4166 240.244
R4127 gnd.n6746 gnd.n6724 240.244
R4128 gnd.n6752 gnd.n6751 240.244
R4129 gnd.n6755 gnd.n6754 240.244
R4130 gnd.n6762 gnd.n6761 240.244
R4131 gnd.n6765 gnd.n6764 240.244
R4132 gnd.n6772 gnd.n6771 240.244
R4133 gnd.n6775 gnd.n6774 240.244
R4134 gnd.n6782 gnd.n6781 240.244
R4135 gnd.n6784 gnd.n6733 240.244
R4136 gnd.n6541 gnd.n273 240.244
R4137 gnd.n6541 gnd.n268 240.244
R4138 gnd.n6548 gnd.n268 240.244
R4139 gnd.n6548 gnd.n257 240.244
R4140 gnd.n257 gnd.n245 240.244
R4141 gnd.n6576 gnd.n245 240.244
R4142 gnd.n6576 gnd.n240 240.244
R4143 gnd.n6593 gnd.n240 240.244
R4144 gnd.n6593 gnd.n231 240.244
R4145 gnd.n6581 gnd.n231 240.244
R4146 gnd.n6581 gnd.n222 240.244
R4147 gnd.n6582 gnd.n222 240.244
R4148 gnd.n6582 gnd.n211 240.244
R4149 gnd.n211 gnd.n200 240.244
R4150 gnd.n6640 gnd.n200 240.244
R4151 gnd.n6640 gnd.n195 240.244
R4152 gnd.n6651 gnd.n195 240.244
R4153 gnd.n6651 gnd.n187 240.244
R4154 gnd.n6644 gnd.n187 240.244
R4155 gnd.n6644 gnd.n179 240.244
R4156 gnd.n179 gnd.n178 240.244
R4157 gnd.n178 gnd.n70 240.244
R4158 gnd.n7108 gnd.n70 240.244
R4159 gnd.n7108 gnd.n72 240.244
R4160 gnd.n85 gnd.n72 240.244
R4161 gnd.n6799 gnd.n85 240.244
R4162 gnd.n6799 gnd.n96 240.244
R4163 gnd.n6804 gnd.n96 240.244
R4164 gnd.n6804 gnd.n106 240.244
R4165 gnd.n6807 gnd.n106 240.244
R4166 gnd.n6807 gnd.n115 240.244
R4167 gnd.n6812 gnd.n115 240.244
R4168 gnd.n6812 gnd.n125 240.244
R4169 gnd.n6815 gnd.n125 240.244
R4170 gnd.n6815 gnd.n134 240.244
R4171 gnd.n6820 gnd.n134 240.244
R4172 gnd.n6820 gnd.n144 240.244
R4173 gnd.n6823 gnd.n144 240.244
R4174 gnd.n6823 gnd.n153 240.244
R4175 gnd.n6828 gnd.n153 240.244
R4176 gnd.n6828 gnd.n163 240.244
R4177 gnd.n6734 gnd.n163 240.244
R4178 gnd.n400 gnd.n399 240.244
R4179 gnd.n408 gnd.n407 240.244
R4180 gnd.n410 gnd.n409 240.244
R4181 gnd.n418 gnd.n417 240.244
R4182 gnd.n426 gnd.n425 240.244
R4183 gnd.n428 gnd.n427 240.244
R4184 gnd.n436 gnd.n435 240.244
R4185 gnd.n446 gnd.n445 240.244
R4186 gnd.n6366 gnd.n322 240.244
R4187 gnd.n6328 gnd.n276 240.244
R4188 gnd.n6324 gnd.n276 240.244
R4189 gnd.n6324 gnd.n259 240.244
R4190 gnd.n6564 gnd.n259 240.244
R4191 gnd.n6564 gnd.n260 240.244
R4192 gnd.n260 gnd.n248 240.244
R4193 gnd.n6559 gnd.n248 240.244
R4194 gnd.n6559 gnd.n232 240.244
R4195 gnd.n6604 gnd.n232 240.244
R4196 gnd.n6604 gnd.n233 240.244
R4197 gnd.n233 gnd.n223 240.244
R4198 gnd.n223 gnd.n213 240.244
R4199 gnd.n6628 gnd.n213 240.244
R4200 gnd.n6628 gnd.n214 240.244
R4201 gnd.n214 gnd.n202 240.244
R4202 gnd.n6623 gnd.n202 240.244
R4203 gnd.n6623 gnd.n189 240.244
R4204 gnd.n6660 gnd.n189 240.244
R4205 gnd.n6660 gnd.n176 240.244
R4206 gnd.n6673 gnd.n176 240.244
R4207 gnd.n6673 gnd.n170 240.244
R4208 gnd.n6681 gnd.n170 240.244
R4209 gnd.n6681 gnd.n75 240.244
R4210 gnd.n87 gnd.n75 240.244
R4211 gnd.n7100 gnd.n87 240.244
R4212 gnd.n7100 gnd.n88 240.244
R4213 gnd.n7096 gnd.n88 240.244
R4214 gnd.n7096 gnd.n94 240.244
R4215 gnd.n7088 gnd.n94 240.244
R4216 gnd.n7088 gnd.n108 240.244
R4217 gnd.n7084 gnd.n108 240.244
R4218 gnd.n7084 gnd.n113 240.244
R4219 gnd.n7076 gnd.n113 240.244
R4220 gnd.n7076 gnd.n127 240.244
R4221 gnd.n7072 gnd.n127 240.244
R4222 gnd.n7072 gnd.n132 240.244
R4223 gnd.n7064 gnd.n132 240.244
R4224 gnd.n7064 gnd.n146 240.244
R4225 gnd.n7060 gnd.n146 240.244
R4226 gnd.n7060 gnd.n151 240.244
R4227 gnd.n7052 gnd.n151 240.244
R4228 gnd.n7052 gnd.n165 240.244
R4229 gnd.n4186 gnd.n1009 240.244
R4230 gnd.n5563 gnd.n5562 240.244
R4231 gnd.n5559 gnd.n5558 240.244
R4232 gnd.n5555 gnd.n5554 240.244
R4233 gnd.n5551 gnd.n5550 240.244
R4234 gnd.n5547 gnd.n5546 240.244
R4235 gnd.n5543 gnd.n5542 240.244
R4236 gnd.n5539 gnd.n5538 240.244
R4237 gnd.n5535 gnd.n5534 240.244
R4238 gnd.n5531 gnd.n5530 240.244
R4239 gnd.n5527 gnd.n5526 240.244
R4240 gnd.n5523 gnd.n5522 240.244
R4241 gnd.n5519 gnd.n5518 240.244
R4242 gnd.n4760 gnd.n4657 240.244
R4243 gnd.n4760 gnd.n4650 240.244
R4244 gnd.n4771 gnd.n4650 240.244
R4245 gnd.n4771 gnd.n4646 240.244
R4246 gnd.n4777 gnd.n4646 240.244
R4247 gnd.n4777 gnd.n4638 240.244
R4248 gnd.n4787 gnd.n4638 240.244
R4249 gnd.n4787 gnd.n4633 240.244
R4250 gnd.n4823 gnd.n4633 240.244
R4251 gnd.n4823 gnd.n4634 240.244
R4252 gnd.n4634 gnd.n4581 240.244
R4253 gnd.n4818 gnd.n4581 240.244
R4254 gnd.n4818 gnd.n4817 240.244
R4255 gnd.n4817 gnd.n4560 240.244
R4256 gnd.n4813 gnd.n4560 240.244
R4257 gnd.n4813 gnd.n4551 240.244
R4258 gnd.n4810 gnd.n4551 240.244
R4259 gnd.n4810 gnd.n4809 240.244
R4260 gnd.n4809 gnd.n4534 240.244
R4261 gnd.n4805 gnd.n4534 240.244
R4262 gnd.n4805 gnd.n4523 240.244
R4263 gnd.n4523 gnd.n4504 240.244
R4264 gnd.n4918 gnd.n4504 240.244
R4265 gnd.n4918 gnd.n4500 240.244
R4266 gnd.n4926 gnd.n4500 240.244
R4267 gnd.n4926 gnd.n4491 240.244
R4268 gnd.n4491 gnd.n4427 240.244
R4269 gnd.n4998 gnd.n4427 240.244
R4270 gnd.n4998 gnd.n4428 240.244
R4271 gnd.n4439 gnd.n4428 240.244
R4272 gnd.n4474 gnd.n4439 240.244
R4273 gnd.n4477 gnd.n4474 240.244
R4274 gnd.n4477 gnd.n4451 240.244
R4275 gnd.n4464 gnd.n4451 240.244
R4276 gnd.n4464 gnd.n4461 240.244
R4277 gnd.n4461 gnd.n4370 240.244
R4278 gnd.n5019 gnd.n4370 240.244
R4279 gnd.n5019 gnd.n4360 240.244
R4280 gnd.n5015 gnd.n4360 240.244
R4281 gnd.n5015 gnd.n4354 240.244
R4282 gnd.n5012 gnd.n4354 240.244
R4283 gnd.n5012 gnd.n4343 240.244
R4284 gnd.n5009 gnd.n4343 240.244
R4285 gnd.n5009 gnd.n4321 240.244
R4286 gnd.n5085 gnd.n4321 240.244
R4287 gnd.n5085 gnd.n4317 240.244
R4288 gnd.n5106 gnd.n4317 240.244
R4289 gnd.n5106 gnd.n4306 240.244
R4290 gnd.n5102 gnd.n4306 240.244
R4291 gnd.n5102 gnd.n4299 240.244
R4292 gnd.n5099 gnd.n4299 240.244
R4293 gnd.n5099 gnd.n4288 240.244
R4294 gnd.n5096 gnd.n4288 240.244
R4295 gnd.n5096 gnd.n4265 240.244
R4296 gnd.n5170 gnd.n4265 240.244
R4297 gnd.n5170 gnd.n4261 240.244
R4298 gnd.n5195 gnd.n4261 240.244
R4299 gnd.n5195 gnd.n4252 240.244
R4300 gnd.n5191 gnd.n4252 240.244
R4301 gnd.n5191 gnd.n4245 240.244
R4302 gnd.n5187 gnd.n4245 240.244
R4303 gnd.n5187 gnd.n4234 240.244
R4304 gnd.n5184 gnd.n4234 240.244
R4305 gnd.n5184 gnd.n4215 240.244
R4306 gnd.n5514 gnd.n4215 240.244
R4307 gnd.n4674 gnd.n4673 240.244
R4308 gnd.n4745 gnd.n4673 240.244
R4309 gnd.n4743 gnd.n4742 240.244
R4310 gnd.n4739 gnd.n4738 240.244
R4311 gnd.n4735 gnd.n4734 240.244
R4312 gnd.n4731 gnd.n4730 240.244
R4313 gnd.n4727 gnd.n4726 240.244
R4314 gnd.n4723 gnd.n4722 240.244
R4315 gnd.n4719 gnd.n4718 240.244
R4316 gnd.n4715 gnd.n4714 240.244
R4317 gnd.n4711 gnd.n4710 240.244
R4318 gnd.n4707 gnd.n4706 240.244
R4319 gnd.n4703 gnd.n4661 240.244
R4320 gnd.n4763 gnd.n4655 240.244
R4321 gnd.n4763 gnd.n4651 240.244
R4322 gnd.n4769 gnd.n4651 240.244
R4323 gnd.n4769 gnd.n4644 240.244
R4324 gnd.n4779 gnd.n4644 240.244
R4325 gnd.n4779 gnd.n4640 240.244
R4326 gnd.n4785 gnd.n4640 240.244
R4327 gnd.n4785 gnd.n4631 240.244
R4328 gnd.n4825 gnd.n4631 240.244
R4329 gnd.n4825 gnd.n4582 240.244
R4330 gnd.n4833 gnd.n4582 240.244
R4331 gnd.n4833 gnd.n4583 240.244
R4332 gnd.n4583 gnd.n4561 240.244
R4333 gnd.n4854 gnd.n4561 240.244
R4334 gnd.n4854 gnd.n4553 240.244
R4335 gnd.n4865 gnd.n4553 240.244
R4336 gnd.n4865 gnd.n4554 240.244
R4337 gnd.n4554 gnd.n4535 240.244
R4338 gnd.n4885 gnd.n4535 240.244
R4339 gnd.n4885 gnd.n4525 240.244
R4340 gnd.n4895 gnd.n4525 240.244
R4341 gnd.n4895 gnd.n4506 240.244
R4342 gnd.n4916 gnd.n4506 240.244
R4343 gnd.n4916 gnd.n4508 240.244
R4344 gnd.n4508 gnd.n4489 240.244
R4345 gnd.n4944 gnd.n4489 240.244
R4346 gnd.n4944 gnd.n4431 240.244
R4347 gnd.n4996 gnd.n4431 240.244
R4348 gnd.n4996 gnd.n4432 240.244
R4349 gnd.n4992 gnd.n4432 240.244
R4350 gnd.n4992 gnd.n4438 240.244
R4351 gnd.n4453 gnd.n4438 240.244
R4352 gnd.n4982 gnd.n4453 240.244
R4353 gnd.n4982 gnd.n4454 240.244
R4354 gnd.n4978 gnd.n4454 240.244
R4355 gnd.n4978 gnd.n4460 240.244
R4356 gnd.n4460 gnd.n4359 240.244
R4357 gnd.n5035 gnd.n4359 240.244
R4358 gnd.n5035 gnd.n4352 240.244
R4359 gnd.n5046 gnd.n4352 240.244
R4360 gnd.n5046 gnd.n4345 240.244
R4361 gnd.n5061 gnd.n4345 240.244
R4362 gnd.n5061 gnd.n4346 240.244
R4363 gnd.n4346 gnd.n4324 240.244
R4364 gnd.n5083 gnd.n4324 240.244
R4365 gnd.n5083 gnd.n4325 240.244
R4366 gnd.n4325 gnd.n4304 240.244
R4367 gnd.n5120 gnd.n4304 240.244
R4368 gnd.n5120 gnd.n4297 240.244
R4369 gnd.n5131 gnd.n4297 240.244
R4370 gnd.n5131 gnd.n4290 240.244
R4371 gnd.n5146 gnd.n4290 240.244
R4372 gnd.n5146 gnd.n4291 240.244
R4373 gnd.n4291 gnd.n4268 240.244
R4374 gnd.n5168 gnd.n4268 240.244
R4375 gnd.n5168 gnd.n4270 240.244
R4376 gnd.n4270 gnd.n4250 240.244
R4377 gnd.n5209 gnd.n4250 240.244
R4378 gnd.n5209 gnd.n4243 240.244
R4379 gnd.n5220 gnd.n4243 240.244
R4380 gnd.n5220 gnd.n4236 240.244
R4381 gnd.n5489 gnd.n4236 240.244
R4382 gnd.n5489 gnd.n4237 240.244
R4383 gnd.n4237 gnd.n4218 240.244
R4384 gnd.n5512 gnd.n4218 240.244
R4385 gnd.n2141 gnd.n1340 240.244
R4386 gnd.n2143 gnd.n2142 240.244
R4387 gnd.n2153 gnd.n2152 240.244
R4388 gnd.n2161 gnd.n2160 240.244
R4389 gnd.n2163 gnd.n2162 240.244
R4390 gnd.n2173 gnd.n2172 240.244
R4391 gnd.n2181 gnd.n2180 240.244
R4392 gnd.n2183 gnd.n2182 240.244
R4393 gnd.n2197 gnd.n2193 240.244
R4394 gnd.n2460 gnd.n1138 240.244
R4395 gnd.n2463 gnd.n1138 240.244
R4396 gnd.n2463 gnd.n1148 240.244
R4397 gnd.n2468 gnd.n1148 240.244
R4398 gnd.n2468 gnd.n1158 240.244
R4399 gnd.n2471 gnd.n1158 240.244
R4400 gnd.n2471 gnd.n1167 240.244
R4401 gnd.n2476 gnd.n1167 240.244
R4402 gnd.n2476 gnd.n1176 240.244
R4403 gnd.n2479 gnd.n1176 240.244
R4404 gnd.n2479 gnd.n1186 240.244
R4405 gnd.n2484 gnd.n1186 240.244
R4406 gnd.n2484 gnd.n1195 240.244
R4407 gnd.n2487 gnd.n1195 240.244
R4408 gnd.n2487 gnd.n1205 240.244
R4409 gnd.n2492 gnd.n1205 240.244
R4410 gnd.n2492 gnd.n1214 240.244
R4411 gnd.n2495 gnd.n1214 240.244
R4412 gnd.n2495 gnd.n1224 240.244
R4413 gnd.n2500 gnd.n1224 240.244
R4414 gnd.n2500 gnd.n1233 240.244
R4415 gnd.n2503 gnd.n1233 240.244
R4416 gnd.n2503 gnd.n1243 240.244
R4417 gnd.n2391 gnd.n1243 240.244
R4418 gnd.n2391 gnd.n1252 240.244
R4419 gnd.n2510 gnd.n1252 240.244
R4420 gnd.n2510 gnd.n1262 240.244
R4421 gnd.n2388 gnd.n1262 240.244
R4422 gnd.n2388 gnd.n1271 240.244
R4423 gnd.n2517 gnd.n1271 240.244
R4424 gnd.n2517 gnd.n1281 240.244
R4425 gnd.n2385 gnd.n1281 240.244
R4426 gnd.n2385 gnd.n1290 240.244
R4427 gnd.n2524 gnd.n1290 240.244
R4428 gnd.n2524 gnd.n1301 240.244
R4429 gnd.n2530 gnd.n1301 240.244
R4430 gnd.n2530 gnd.n1311 240.244
R4431 gnd.n2544 gnd.n1311 240.244
R4432 gnd.n2544 gnd.n1322 240.244
R4433 gnd.n2564 gnd.n1322 240.244
R4434 gnd.n2564 gnd.n1331 240.244
R4435 gnd.n2599 gnd.n1331 240.244
R4436 gnd.n2420 gnd.n2419 240.244
R4437 gnd.n2426 gnd.n2425 240.244
R4438 gnd.n2430 gnd.n2429 240.244
R4439 gnd.n2436 gnd.n2435 240.244
R4440 gnd.n2440 gnd.n2439 240.244
R4441 gnd.n2446 gnd.n2445 240.244
R4442 gnd.n2450 gnd.n2449 240.244
R4443 gnd.n2409 gnd.n2408 240.244
R4444 gnd.n2404 gnd.n1060 240.244
R4445 gnd.n4035 gnd.n4034 240.244
R4446 gnd.n4034 gnd.n1134 240.244
R4447 gnd.n4024 gnd.n1134 240.244
R4448 gnd.n4024 gnd.n1150 240.244
R4449 gnd.n4020 gnd.n1150 240.244
R4450 gnd.n4020 gnd.n1156 240.244
R4451 gnd.n4012 gnd.n1156 240.244
R4452 gnd.n4012 gnd.n1169 240.244
R4453 gnd.n4008 gnd.n1169 240.244
R4454 gnd.n4008 gnd.n1174 240.244
R4455 gnd.n4000 gnd.n1174 240.244
R4456 gnd.n4000 gnd.n1187 240.244
R4457 gnd.n3996 gnd.n1187 240.244
R4458 gnd.n3996 gnd.n1192 240.244
R4459 gnd.n3988 gnd.n1192 240.244
R4460 gnd.n3988 gnd.n1207 240.244
R4461 gnd.n3984 gnd.n1207 240.244
R4462 gnd.n3984 gnd.n1212 240.244
R4463 gnd.n3976 gnd.n1212 240.244
R4464 gnd.n3976 gnd.n1225 240.244
R4465 gnd.n3972 gnd.n1225 240.244
R4466 gnd.n3972 gnd.n1230 240.244
R4467 gnd.n3964 gnd.n1230 240.244
R4468 gnd.n3964 gnd.n1245 240.244
R4469 gnd.n3960 gnd.n1245 240.244
R4470 gnd.n3960 gnd.n1250 240.244
R4471 gnd.n3952 gnd.n1250 240.244
R4472 gnd.n3952 gnd.n1263 240.244
R4473 gnd.n3948 gnd.n1263 240.244
R4474 gnd.n3948 gnd.n1268 240.244
R4475 gnd.n3940 gnd.n1268 240.244
R4476 gnd.n3940 gnd.n1283 240.244
R4477 gnd.n3936 gnd.n1283 240.244
R4478 gnd.n3936 gnd.n1288 240.244
R4479 gnd.n3928 gnd.n1288 240.244
R4480 gnd.n3928 gnd.n1303 240.244
R4481 gnd.n3924 gnd.n1303 240.244
R4482 gnd.n3924 gnd.n1308 240.244
R4483 gnd.n3916 gnd.n1308 240.244
R4484 gnd.n3916 gnd.n1324 240.244
R4485 gnd.n3912 gnd.n1324 240.244
R4486 gnd.n3912 gnd.n1329 240.244
R4487 gnd.n5775 gnd.n836 240.244
R4488 gnd.n5781 gnd.n836 240.244
R4489 gnd.n5781 gnd.n834 240.244
R4490 gnd.n5785 gnd.n834 240.244
R4491 gnd.n5785 gnd.n830 240.244
R4492 gnd.n5791 gnd.n830 240.244
R4493 gnd.n5791 gnd.n828 240.244
R4494 gnd.n5795 gnd.n828 240.244
R4495 gnd.n5795 gnd.n824 240.244
R4496 gnd.n5801 gnd.n824 240.244
R4497 gnd.n5801 gnd.n822 240.244
R4498 gnd.n5805 gnd.n822 240.244
R4499 gnd.n5805 gnd.n818 240.244
R4500 gnd.n5811 gnd.n818 240.244
R4501 gnd.n5811 gnd.n816 240.244
R4502 gnd.n5815 gnd.n816 240.244
R4503 gnd.n5815 gnd.n812 240.244
R4504 gnd.n5821 gnd.n812 240.244
R4505 gnd.n5821 gnd.n810 240.244
R4506 gnd.n5825 gnd.n810 240.244
R4507 gnd.n5825 gnd.n806 240.244
R4508 gnd.n5831 gnd.n806 240.244
R4509 gnd.n5831 gnd.n804 240.244
R4510 gnd.n5835 gnd.n804 240.244
R4511 gnd.n5835 gnd.n800 240.244
R4512 gnd.n5841 gnd.n800 240.244
R4513 gnd.n5841 gnd.n798 240.244
R4514 gnd.n5845 gnd.n798 240.244
R4515 gnd.n5845 gnd.n794 240.244
R4516 gnd.n5851 gnd.n794 240.244
R4517 gnd.n5851 gnd.n792 240.244
R4518 gnd.n5855 gnd.n792 240.244
R4519 gnd.n5855 gnd.n788 240.244
R4520 gnd.n5861 gnd.n788 240.244
R4521 gnd.n5861 gnd.n786 240.244
R4522 gnd.n5865 gnd.n786 240.244
R4523 gnd.n5865 gnd.n782 240.244
R4524 gnd.n5871 gnd.n782 240.244
R4525 gnd.n5871 gnd.n780 240.244
R4526 gnd.n5875 gnd.n780 240.244
R4527 gnd.n5875 gnd.n776 240.244
R4528 gnd.n5881 gnd.n776 240.244
R4529 gnd.n5881 gnd.n774 240.244
R4530 gnd.n5885 gnd.n774 240.244
R4531 gnd.n5885 gnd.n770 240.244
R4532 gnd.n5891 gnd.n770 240.244
R4533 gnd.n5891 gnd.n768 240.244
R4534 gnd.n5895 gnd.n768 240.244
R4535 gnd.n5895 gnd.n764 240.244
R4536 gnd.n5901 gnd.n764 240.244
R4537 gnd.n5901 gnd.n762 240.244
R4538 gnd.n5905 gnd.n762 240.244
R4539 gnd.n5905 gnd.n758 240.244
R4540 gnd.n5911 gnd.n758 240.244
R4541 gnd.n5911 gnd.n756 240.244
R4542 gnd.n5915 gnd.n756 240.244
R4543 gnd.n5915 gnd.n752 240.244
R4544 gnd.n5921 gnd.n752 240.244
R4545 gnd.n5921 gnd.n750 240.244
R4546 gnd.n5925 gnd.n750 240.244
R4547 gnd.n5925 gnd.n746 240.244
R4548 gnd.n5931 gnd.n746 240.244
R4549 gnd.n5931 gnd.n744 240.244
R4550 gnd.n5935 gnd.n744 240.244
R4551 gnd.n5935 gnd.n740 240.244
R4552 gnd.n5941 gnd.n740 240.244
R4553 gnd.n5941 gnd.n738 240.244
R4554 gnd.n5945 gnd.n738 240.244
R4555 gnd.n5945 gnd.n734 240.244
R4556 gnd.n5951 gnd.n734 240.244
R4557 gnd.n5951 gnd.n732 240.244
R4558 gnd.n5955 gnd.n732 240.244
R4559 gnd.n5955 gnd.n728 240.244
R4560 gnd.n5961 gnd.n728 240.244
R4561 gnd.n5961 gnd.n726 240.244
R4562 gnd.n5965 gnd.n726 240.244
R4563 gnd.n5965 gnd.n722 240.244
R4564 gnd.n5971 gnd.n722 240.244
R4565 gnd.n5971 gnd.n720 240.244
R4566 gnd.n5975 gnd.n720 240.244
R4567 gnd.n5975 gnd.n716 240.244
R4568 gnd.n5981 gnd.n716 240.244
R4569 gnd.n5981 gnd.n714 240.244
R4570 gnd.n5985 gnd.n714 240.244
R4571 gnd.n5985 gnd.n710 240.244
R4572 gnd.n5991 gnd.n710 240.244
R4573 gnd.n5991 gnd.n708 240.244
R4574 gnd.n5995 gnd.n708 240.244
R4575 gnd.n5995 gnd.n704 240.244
R4576 gnd.n6001 gnd.n704 240.244
R4577 gnd.n6001 gnd.n702 240.244
R4578 gnd.n6005 gnd.n702 240.244
R4579 gnd.n6005 gnd.n698 240.244
R4580 gnd.n6011 gnd.n698 240.244
R4581 gnd.n6011 gnd.n696 240.244
R4582 gnd.n6015 gnd.n696 240.244
R4583 gnd.n6015 gnd.n692 240.244
R4584 gnd.n6021 gnd.n692 240.244
R4585 gnd.n6021 gnd.n690 240.244
R4586 gnd.n6025 gnd.n690 240.244
R4587 gnd.n6025 gnd.n686 240.244
R4588 gnd.n6031 gnd.n686 240.244
R4589 gnd.n6031 gnd.n684 240.244
R4590 gnd.n6035 gnd.n684 240.244
R4591 gnd.n6035 gnd.n680 240.244
R4592 gnd.n6041 gnd.n680 240.244
R4593 gnd.n6041 gnd.n678 240.244
R4594 gnd.n6045 gnd.n678 240.244
R4595 gnd.n6045 gnd.n674 240.244
R4596 gnd.n6051 gnd.n674 240.244
R4597 gnd.n6051 gnd.n672 240.244
R4598 gnd.n6055 gnd.n672 240.244
R4599 gnd.n6055 gnd.n668 240.244
R4600 gnd.n6061 gnd.n668 240.244
R4601 gnd.n6061 gnd.n666 240.244
R4602 gnd.n6065 gnd.n666 240.244
R4603 gnd.n6065 gnd.n662 240.244
R4604 gnd.n6071 gnd.n662 240.244
R4605 gnd.n6071 gnd.n660 240.244
R4606 gnd.n6075 gnd.n660 240.244
R4607 gnd.n6075 gnd.n656 240.244
R4608 gnd.n6081 gnd.n656 240.244
R4609 gnd.n6081 gnd.n654 240.244
R4610 gnd.n6085 gnd.n654 240.244
R4611 gnd.n6085 gnd.n650 240.244
R4612 gnd.n6091 gnd.n650 240.244
R4613 gnd.n6091 gnd.n648 240.244
R4614 gnd.n6095 gnd.n648 240.244
R4615 gnd.n6101 gnd.n644 240.244
R4616 gnd.n6101 gnd.n642 240.244
R4617 gnd.n6105 gnd.n642 240.244
R4618 gnd.n6105 gnd.n638 240.244
R4619 gnd.n6111 gnd.n638 240.244
R4620 gnd.n6111 gnd.n636 240.244
R4621 gnd.n6115 gnd.n636 240.244
R4622 gnd.n6115 gnd.n632 240.244
R4623 gnd.n6121 gnd.n632 240.244
R4624 gnd.n6121 gnd.n630 240.244
R4625 gnd.n6125 gnd.n630 240.244
R4626 gnd.n6125 gnd.n626 240.244
R4627 gnd.n6131 gnd.n626 240.244
R4628 gnd.n6131 gnd.n624 240.244
R4629 gnd.n6135 gnd.n624 240.244
R4630 gnd.n6135 gnd.n620 240.244
R4631 gnd.n6141 gnd.n620 240.244
R4632 gnd.n6141 gnd.n618 240.244
R4633 gnd.n6145 gnd.n618 240.244
R4634 gnd.n6145 gnd.n614 240.244
R4635 gnd.n6151 gnd.n614 240.244
R4636 gnd.n6151 gnd.n612 240.244
R4637 gnd.n6155 gnd.n612 240.244
R4638 gnd.n6155 gnd.n608 240.244
R4639 gnd.n6161 gnd.n608 240.244
R4640 gnd.n6161 gnd.n606 240.244
R4641 gnd.n6165 gnd.n606 240.244
R4642 gnd.n6165 gnd.n602 240.244
R4643 gnd.n6171 gnd.n602 240.244
R4644 gnd.n6171 gnd.n600 240.244
R4645 gnd.n6175 gnd.n600 240.244
R4646 gnd.n6175 gnd.n596 240.244
R4647 gnd.n6181 gnd.n596 240.244
R4648 gnd.n6181 gnd.n594 240.244
R4649 gnd.n6185 gnd.n594 240.244
R4650 gnd.n6185 gnd.n590 240.244
R4651 gnd.n6191 gnd.n590 240.244
R4652 gnd.n6191 gnd.n588 240.244
R4653 gnd.n6195 gnd.n588 240.244
R4654 gnd.n6195 gnd.n584 240.244
R4655 gnd.n6201 gnd.n584 240.244
R4656 gnd.n6201 gnd.n582 240.244
R4657 gnd.n6205 gnd.n582 240.244
R4658 gnd.n6205 gnd.n578 240.244
R4659 gnd.n6211 gnd.n578 240.244
R4660 gnd.n6211 gnd.n576 240.244
R4661 gnd.n6215 gnd.n576 240.244
R4662 gnd.n6215 gnd.n572 240.244
R4663 gnd.n6221 gnd.n572 240.244
R4664 gnd.n6221 gnd.n570 240.244
R4665 gnd.n6225 gnd.n570 240.244
R4666 gnd.n6225 gnd.n566 240.244
R4667 gnd.n6231 gnd.n566 240.244
R4668 gnd.n6231 gnd.n564 240.244
R4669 gnd.n6235 gnd.n564 240.244
R4670 gnd.n6235 gnd.n560 240.244
R4671 gnd.n6241 gnd.n560 240.244
R4672 gnd.n6241 gnd.n558 240.244
R4673 gnd.n6245 gnd.n558 240.244
R4674 gnd.n6245 gnd.n554 240.244
R4675 gnd.n6251 gnd.n554 240.244
R4676 gnd.n6251 gnd.n552 240.244
R4677 gnd.n6255 gnd.n552 240.244
R4678 gnd.n6255 gnd.n548 240.244
R4679 gnd.n6261 gnd.n548 240.244
R4680 gnd.n6261 gnd.n546 240.244
R4681 gnd.n6265 gnd.n546 240.244
R4682 gnd.n6265 gnd.n542 240.244
R4683 gnd.n6271 gnd.n542 240.244
R4684 gnd.n6271 gnd.n540 240.244
R4685 gnd.n6275 gnd.n540 240.244
R4686 gnd.n6275 gnd.n536 240.244
R4687 gnd.n6281 gnd.n536 240.244
R4688 gnd.n6281 gnd.n534 240.244
R4689 gnd.n6285 gnd.n534 240.244
R4690 gnd.n6285 gnd.n530 240.244
R4691 gnd.n6291 gnd.n530 240.244
R4692 gnd.n6291 gnd.n528 240.244
R4693 gnd.n6295 gnd.n528 240.244
R4694 gnd.n6295 gnd.n524 240.244
R4695 gnd.n6303 gnd.n524 240.244
R4696 gnd.n6303 gnd.n522 240.244
R4697 gnd.n6308 gnd.n522 240.244
R4698 gnd.n6309 gnd.n6308 240.244
R4699 gnd.n2308 gnd.n2307 240.244
R4700 gnd.n2308 gnd.n2302 240.244
R4701 gnd.n2314 gnd.n2302 240.244
R4702 gnd.n2315 gnd.n2314 240.244
R4703 gnd.n2567 gnd.n2315 240.244
R4704 gnd.n2567 gnd.n2297 240.244
R4705 gnd.n2596 gnd.n2297 240.244
R4706 gnd.n2596 gnd.n2298 240.244
R4707 gnd.n2592 gnd.n2298 240.244
R4708 gnd.n2592 gnd.n2591 240.244
R4709 gnd.n2591 gnd.n2589 240.244
R4710 gnd.n2589 gnd.n2575 240.244
R4711 gnd.n2585 gnd.n2575 240.244
R4712 gnd.n2585 gnd.n2582 240.244
R4713 gnd.n2582 gnd.n2094 240.244
R4714 gnd.n2681 gnd.n2094 240.244
R4715 gnd.n2681 gnd.n2089 240.244
R4716 gnd.n2689 gnd.n2089 240.244
R4717 gnd.n2689 gnd.n2090 240.244
R4718 gnd.n2090 gnd.n2069 240.244
R4719 gnd.n2711 gnd.n2069 240.244
R4720 gnd.n2711 gnd.n2064 240.244
R4721 gnd.n2719 gnd.n2064 240.244
R4722 gnd.n2719 gnd.n2065 240.244
R4723 gnd.n2065 gnd.n2044 240.244
R4724 gnd.n2741 gnd.n2044 240.244
R4725 gnd.n2741 gnd.n2038 240.244
R4726 gnd.n2749 gnd.n2038 240.244
R4727 gnd.n2749 gnd.n2040 240.244
R4728 gnd.n2040 gnd.n2019 240.244
R4729 gnd.n2774 gnd.n2019 240.244
R4730 gnd.n2774 gnd.n2014 240.244
R4731 gnd.n2794 gnd.n2014 240.244
R4732 gnd.n2794 gnd.n2015 240.244
R4733 gnd.n2790 gnd.n2015 240.244
R4734 gnd.n2790 gnd.n2789 240.244
R4735 gnd.n2789 gnd.n2788 240.244
R4736 gnd.n2788 gnd.n2782 240.244
R4737 gnd.n2782 gnd.n1989 240.244
R4738 gnd.n2926 gnd.n1989 240.244
R4739 gnd.n2926 gnd.n1984 240.244
R4740 gnd.n2934 gnd.n1984 240.244
R4741 gnd.n2934 gnd.n1985 240.244
R4742 gnd.n1985 gnd.n1961 240.244
R4743 gnd.n2968 gnd.n1961 240.244
R4744 gnd.n2968 gnd.n1957 240.244
R4745 gnd.n2974 gnd.n1957 240.244
R4746 gnd.n2974 gnd.n1938 240.244
R4747 gnd.n3012 gnd.n1938 240.244
R4748 gnd.n3012 gnd.n1934 240.244
R4749 gnd.n3018 gnd.n1934 240.244
R4750 gnd.n3018 gnd.n1920 240.244
R4751 gnd.n3068 gnd.n1920 240.244
R4752 gnd.n3068 gnd.n1916 240.244
R4753 gnd.n3074 gnd.n1916 240.244
R4754 gnd.n3074 gnd.n1898 240.244
R4755 gnd.n3096 gnd.n1898 240.244
R4756 gnd.n3096 gnd.n1893 240.244
R4757 gnd.n3104 gnd.n1893 240.244
R4758 gnd.n3104 gnd.n1894 240.244
R4759 gnd.n1894 gnd.n1866 240.244
R4760 gnd.n3141 gnd.n1866 240.244
R4761 gnd.n3141 gnd.n1862 240.244
R4762 gnd.n3147 gnd.n1862 240.244
R4763 gnd.n3147 gnd.n1842 240.244
R4764 gnd.n3182 gnd.n1842 240.244
R4765 gnd.n3182 gnd.n1838 240.244
R4766 gnd.n3188 gnd.n1838 240.244
R4767 gnd.n3188 gnd.n1825 240.244
R4768 gnd.n3241 gnd.n1825 240.244
R4769 gnd.n3241 gnd.n1821 240.244
R4770 gnd.n3247 gnd.n1821 240.244
R4771 gnd.n3247 gnd.n1804 240.244
R4772 gnd.n3268 gnd.n1804 240.244
R4773 gnd.n3268 gnd.n1799 240.244
R4774 gnd.n3276 gnd.n1799 240.244
R4775 gnd.n3276 gnd.n1800 240.244
R4776 gnd.n1800 gnd.n1775 240.244
R4777 gnd.n3315 gnd.n1775 240.244
R4778 gnd.n3315 gnd.n1771 240.244
R4779 gnd.n3321 gnd.n1771 240.244
R4780 gnd.n3321 gnd.n1752 240.244
R4781 gnd.n3356 gnd.n1752 240.244
R4782 gnd.n3356 gnd.n1748 240.244
R4783 gnd.n3362 gnd.n1748 240.244
R4784 gnd.n3362 gnd.n1736 240.244
R4785 gnd.n3398 gnd.n1736 240.244
R4786 gnd.n3398 gnd.n1732 240.244
R4787 gnd.n3404 gnd.n1732 240.244
R4788 gnd.n3404 gnd.n1644 240.244
R4789 gnd.n3545 gnd.n1644 240.244
R4790 gnd.n3545 gnd.n1640 240.244
R4791 gnd.n3551 gnd.n1640 240.244
R4792 gnd.n3551 gnd.n1631 240.244
R4793 gnd.n3565 gnd.n1631 240.244
R4794 gnd.n3565 gnd.n1627 240.244
R4795 gnd.n3571 gnd.n1627 240.244
R4796 gnd.n3571 gnd.n1620 240.244
R4797 gnd.n3587 gnd.n1620 240.244
R4798 gnd.n3587 gnd.n1616 240.244
R4799 gnd.n3593 gnd.n1616 240.244
R4800 gnd.n3593 gnd.n1607 240.244
R4801 gnd.n3607 gnd.n1607 240.244
R4802 gnd.n3607 gnd.n1603 240.244
R4803 gnd.n3613 gnd.n1603 240.244
R4804 gnd.n3613 gnd.n1594 240.244
R4805 gnd.n3627 gnd.n1594 240.244
R4806 gnd.n3627 gnd.n1590 240.244
R4807 gnd.n3633 gnd.n1590 240.244
R4808 gnd.n3633 gnd.n1580 240.244
R4809 gnd.n3647 gnd.n1580 240.244
R4810 gnd.n3647 gnd.n1575 240.244
R4811 gnd.n3659 gnd.n1575 240.244
R4812 gnd.n3659 gnd.n1576 240.244
R4813 gnd.n3655 gnd.n1576 240.244
R4814 gnd.n3655 gnd.n491 240.244
R4815 gnd.n6337 gnd.n491 240.244
R4816 gnd.n6337 gnd.n492 240.244
R4817 gnd.n6333 gnd.n492 240.244
R4818 gnd.n6333 gnd.n6332 240.244
R4819 gnd.n6332 gnd.n6331 240.244
R4820 gnd.n6331 gnd.n498 240.244
R4821 gnd.n6321 gnd.n498 240.244
R4822 gnd.n6321 gnd.n507 240.244
R4823 gnd.n6317 gnd.n507 240.244
R4824 gnd.n6317 gnd.n6316 240.244
R4825 gnd.n6316 gnd.n6315 240.244
R4826 gnd.n6315 gnd.n517 240.244
R4827 gnd.n5771 gnd.n839 240.244
R4828 gnd.n5771 gnd.n841 240.244
R4829 gnd.n5767 gnd.n841 240.244
R4830 gnd.n5767 gnd.n847 240.244
R4831 gnd.n5763 gnd.n847 240.244
R4832 gnd.n5763 gnd.n849 240.244
R4833 gnd.n5759 gnd.n849 240.244
R4834 gnd.n5759 gnd.n855 240.244
R4835 gnd.n5755 gnd.n855 240.244
R4836 gnd.n5755 gnd.n857 240.244
R4837 gnd.n5751 gnd.n857 240.244
R4838 gnd.n5751 gnd.n863 240.244
R4839 gnd.n5747 gnd.n863 240.244
R4840 gnd.n5747 gnd.n865 240.244
R4841 gnd.n5743 gnd.n865 240.244
R4842 gnd.n5743 gnd.n871 240.244
R4843 gnd.n5739 gnd.n871 240.244
R4844 gnd.n5739 gnd.n873 240.244
R4845 gnd.n5735 gnd.n873 240.244
R4846 gnd.n5735 gnd.n879 240.244
R4847 gnd.n5731 gnd.n879 240.244
R4848 gnd.n5731 gnd.n881 240.244
R4849 gnd.n5727 gnd.n881 240.244
R4850 gnd.n5727 gnd.n887 240.244
R4851 gnd.n5723 gnd.n887 240.244
R4852 gnd.n5723 gnd.n889 240.244
R4853 gnd.n5719 gnd.n889 240.244
R4854 gnd.n5719 gnd.n895 240.244
R4855 gnd.n5715 gnd.n895 240.244
R4856 gnd.n5715 gnd.n897 240.244
R4857 gnd.n5711 gnd.n897 240.244
R4858 gnd.n5711 gnd.n903 240.244
R4859 gnd.n5707 gnd.n903 240.244
R4860 gnd.n5707 gnd.n905 240.244
R4861 gnd.n5703 gnd.n905 240.244
R4862 gnd.n5703 gnd.n911 240.244
R4863 gnd.n5699 gnd.n911 240.244
R4864 gnd.n5699 gnd.n913 240.244
R4865 gnd.n5695 gnd.n913 240.244
R4866 gnd.n5695 gnd.n919 240.244
R4867 gnd.n5691 gnd.n919 240.244
R4868 gnd.n5691 gnd.n921 240.244
R4869 gnd.n5687 gnd.n921 240.244
R4870 gnd.n5687 gnd.n927 240.244
R4871 gnd.n5683 gnd.n927 240.244
R4872 gnd.n5683 gnd.n929 240.244
R4873 gnd.n5679 gnd.n929 240.244
R4874 gnd.n5679 gnd.n935 240.244
R4875 gnd.n5675 gnd.n935 240.244
R4876 gnd.n5675 gnd.n937 240.244
R4877 gnd.n5671 gnd.n937 240.244
R4878 gnd.n5671 gnd.n943 240.244
R4879 gnd.n5667 gnd.n943 240.244
R4880 gnd.n5667 gnd.n945 240.244
R4881 gnd.n5663 gnd.n945 240.244
R4882 gnd.n5663 gnd.n951 240.244
R4883 gnd.n5659 gnd.n951 240.244
R4884 gnd.n5659 gnd.n953 240.244
R4885 gnd.n5655 gnd.n953 240.244
R4886 gnd.n5655 gnd.n959 240.244
R4887 gnd.n5651 gnd.n959 240.244
R4888 gnd.n5651 gnd.n961 240.244
R4889 gnd.n5647 gnd.n961 240.244
R4890 gnd.n5647 gnd.n967 240.244
R4891 gnd.n5643 gnd.n967 240.244
R4892 gnd.n5643 gnd.n969 240.244
R4893 gnd.n5639 gnd.n969 240.244
R4894 gnd.n5639 gnd.n975 240.244
R4895 gnd.n5635 gnd.n975 240.244
R4896 gnd.n5635 gnd.n977 240.244
R4897 gnd.n5631 gnd.n977 240.244
R4898 gnd.n5631 gnd.n983 240.244
R4899 gnd.n5627 gnd.n983 240.244
R4900 gnd.n5627 gnd.n985 240.244
R4901 gnd.n5623 gnd.n985 240.244
R4902 gnd.n5623 gnd.n991 240.244
R4903 gnd.n5619 gnd.n991 240.244
R4904 gnd.n5619 gnd.n993 240.244
R4905 gnd.n5615 gnd.n993 240.244
R4906 gnd.n5615 gnd.n999 240.244
R4907 gnd.n5611 gnd.n999 240.244
R4908 gnd.n5611 gnd.n1001 240.244
R4909 gnd.n5607 gnd.n1001 240.244
R4910 gnd.n5607 gnd.n1007 240.244
R4911 gnd.n2669 gnd.n2104 240.244
R4912 gnd.n2669 gnd.n2105 240.244
R4913 gnd.n2105 gnd.n2085 240.244
R4914 gnd.n2692 gnd.n2085 240.244
R4915 gnd.n2692 gnd.n2079 240.244
R4916 gnd.n2699 gnd.n2079 240.244
R4917 gnd.n2699 gnd.n2080 240.244
R4918 gnd.n2080 gnd.n2060 240.244
R4919 gnd.n2722 gnd.n2060 240.244
R4920 gnd.n2722 gnd.n2054 240.244
R4921 gnd.n2729 gnd.n2054 240.244
R4922 gnd.n2729 gnd.n2055 240.244
R4923 gnd.n2055 gnd.n2034 240.244
R4924 gnd.n2752 gnd.n2034 240.244
R4925 gnd.n2752 gnd.n2028 240.244
R4926 gnd.n2759 gnd.n2028 240.244
R4927 gnd.n2759 gnd.n2029 240.244
R4928 gnd.n2029 gnd.n2010 240.244
R4929 gnd.n2797 gnd.n2010 240.244
R4930 gnd.n2797 gnd.n2004 240.244
R4931 gnd.n2804 gnd.n2004 240.244
R4932 gnd.n2804 gnd.n2005 240.244
R4933 gnd.n2005 gnd.n1475 240.244
R4934 gnd.n3777 gnd.n1475 240.244
R4935 gnd.n3777 gnd.n1476 240.244
R4936 gnd.n1481 gnd.n1476 240.244
R4937 gnd.n1482 gnd.n1481 240.244
R4938 gnd.n1483 gnd.n1482 240.244
R4939 gnd.n2943 gnd.n1483 240.244
R4940 gnd.n2943 gnd.n1486 240.244
R4941 gnd.n1487 gnd.n1486 240.244
R4942 gnd.n1488 gnd.n1487 240.244
R4943 gnd.n2976 gnd.n1488 240.244
R4944 gnd.n2976 gnd.n1491 240.244
R4945 gnd.n1492 gnd.n1491 240.244
R4946 gnd.n1493 gnd.n1492 240.244
R4947 gnd.n1932 gnd.n1493 240.244
R4948 gnd.n1932 gnd.n1496 240.244
R4949 gnd.n1497 gnd.n1496 240.244
R4950 gnd.n1498 gnd.n1497 240.244
R4951 gnd.n3076 gnd.n1498 240.244
R4952 gnd.n3076 gnd.n1501 240.244
R4953 gnd.n1502 gnd.n1501 240.244
R4954 gnd.n1503 gnd.n1502 240.244
R4955 gnd.n1890 gnd.n1503 240.244
R4956 gnd.n1890 gnd.n1506 240.244
R4957 gnd.n1507 gnd.n1506 240.244
R4958 gnd.n1508 gnd.n1507 240.244
R4959 gnd.n3138 gnd.n1508 240.244
R4960 gnd.n3138 gnd.n1511 240.244
R4961 gnd.n1512 gnd.n1511 240.244
R4962 gnd.n1513 gnd.n1512 240.244
R4963 gnd.n3152 gnd.n1513 240.244
R4964 gnd.n3152 gnd.n1516 240.244
R4965 gnd.n1517 gnd.n1516 240.244
R4966 gnd.n1518 gnd.n1517 240.244
R4967 gnd.n1828 gnd.n1518 240.244
R4968 gnd.n1828 gnd.n1521 240.244
R4969 gnd.n1522 gnd.n1521 240.244
R4970 gnd.n1523 gnd.n1522 240.244
R4971 gnd.n3207 gnd.n1523 240.244
R4972 gnd.n3207 gnd.n1526 240.244
R4973 gnd.n1527 gnd.n1526 240.244
R4974 gnd.n1528 gnd.n1527 240.244
R4975 gnd.n3299 gnd.n1528 240.244
R4976 gnd.n3299 gnd.n1531 240.244
R4977 gnd.n1532 gnd.n1531 240.244
R4978 gnd.n1533 gnd.n1532 240.244
R4979 gnd.n3334 gnd.n1533 240.244
R4980 gnd.n3334 gnd.n1536 240.244
R4981 gnd.n1537 gnd.n1536 240.244
R4982 gnd.n1538 gnd.n1537 240.244
R4983 gnd.n1737 gnd.n1538 240.244
R4984 gnd.n1737 gnd.n1541 240.244
R4985 gnd.n1542 gnd.n1541 240.244
R4986 gnd.n1543 gnd.n1542 240.244
R4987 gnd.n3415 gnd.n1543 240.244
R4988 gnd.n3415 gnd.n1546 240.244
R4989 gnd.n1547 gnd.n1546 240.244
R4990 gnd.n1548 gnd.n1547 240.244
R4991 gnd.n1632 gnd.n1548 240.244
R4992 gnd.n1632 gnd.n1551 240.244
R4993 gnd.n1552 gnd.n1551 240.244
R4994 gnd.n1553 gnd.n1552 240.244
R4995 gnd.n3573 gnd.n1553 240.244
R4996 gnd.n3573 gnd.n1556 240.244
R4997 gnd.n1557 gnd.n1556 240.244
R4998 gnd.n1558 gnd.n1557 240.244
R4999 gnd.n1608 gnd.n1558 240.244
R5000 gnd.n1608 gnd.n1561 240.244
R5001 gnd.n1562 gnd.n1561 240.244
R5002 gnd.n1563 gnd.n1562 240.244
R5003 gnd.n1595 gnd.n1563 240.244
R5004 gnd.n1595 gnd.n1566 240.244
R5005 gnd.n1567 gnd.n1566 240.244
R5006 gnd.n1568 gnd.n1567 240.244
R5007 gnd.n1581 gnd.n1568 240.244
R5008 gnd.n1581 gnd.n1571 240.244
R5009 gnd.n3662 gnd.n1571 240.244
R5010 gnd.n3662 gnd.n459 240.244
R5011 gnd.n6354 gnd.n459 240.244
R5012 gnd.n2659 gnd.n2110 240.244
R5013 gnd.n2659 gnd.n2126 240.244
R5014 gnd.n2130 gnd.n2129 240.244
R5015 gnd.n2132 gnd.n2131 240.244
R5016 gnd.n2137 gnd.n2136 240.244
R5017 gnd.n2147 gnd.n2146 240.244
R5018 gnd.n2149 gnd.n2148 240.244
R5019 gnd.n2157 gnd.n2156 240.244
R5020 gnd.n2167 gnd.n2166 240.244
R5021 gnd.n2169 gnd.n2168 240.244
R5022 gnd.n2177 gnd.n2176 240.244
R5023 gnd.n2187 gnd.n2186 240.244
R5024 gnd.n2549 gnd.n2188 240.244
R5025 gnd.n2554 gnd.n2553 240.244
R5026 gnd.n2671 gnd.n2101 240.244
R5027 gnd.n2671 gnd.n2096 240.244
R5028 gnd.n2678 gnd.n2096 240.244
R5029 gnd.n2678 gnd.n2087 240.244
R5030 gnd.n2087 gnd.n2076 240.244
R5031 gnd.n2701 gnd.n2076 240.244
R5032 gnd.n2701 gnd.n2071 240.244
R5033 gnd.n2708 gnd.n2071 240.244
R5034 gnd.n2708 gnd.n2062 240.244
R5035 gnd.n2062 gnd.n2051 240.244
R5036 gnd.n2731 gnd.n2051 240.244
R5037 gnd.n2731 gnd.n2046 240.244
R5038 gnd.n2738 gnd.n2046 240.244
R5039 gnd.n2738 gnd.n2036 240.244
R5040 gnd.n2036 gnd.n2026 240.244
R5041 gnd.n2761 gnd.n2026 240.244
R5042 gnd.n2761 gnd.n2021 240.244
R5043 gnd.n2771 gnd.n2021 240.244
R5044 gnd.n2771 gnd.n2012 240.244
R5045 gnd.n2012 gnd.n2000 240.244
R5046 gnd.n2806 gnd.n2000 240.244
R5047 gnd.n2807 gnd.n2806 240.244
R5048 gnd.n2877 gnd.n2807 240.244
R5049 gnd.n2877 gnd.n1473 240.244
R5050 gnd.n2887 gnd.n1473 240.244
R5051 gnd.n2887 gnd.n1994 240.244
R5052 gnd.n2881 gnd.n1994 240.244
R5053 gnd.n2881 gnd.n1975 240.244
R5054 gnd.n2945 gnd.n1975 240.244
R5055 gnd.n2945 gnd.n1971 240.244
R5056 gnd.n2951 gnd.n1971 240.244
R5057 gnd.n2951 gnd.n1953 240.244
R5058 gnd.n2978 gnd.n1953 240.244
R5059 gnd.n2978 gnd.n1947 240.244
R5060 gnd.n2994 gnd.n1947 240.244
R5061 gnd.n2994 gnd.n1948 240.244
R5062 gnd.n2983 gnd.n1948 240.244
R5063 gnd.n2984 gnd.n2983 240.244
R5064 gnd.n2985 gnd.n2984 240.244
R5065 gnd.n2985 gnd.n1913 240.244
R5066 gnd.n3078 gnd.n1913 240.244
R5067 gnd.n3078 gnd.n1907 240.244
R5068 gnd.n3085 gnd.n1907 240.244
R5069 gnd.n3085 gnd.n1908 240.244
R5070 gnd.n1908 gnd.n1883 240.244
R5071 gnd.n3114 gnd.n1883 240.244
R5072 gnd.n3114 gnd.n1878 240.244
R5073 gnd.n3124 gnd.n1878 240.244
R5074 gnd.n3124 gnd.n1868 240.244
R5075 gnd.n3118 gnd.n1868 240.244
R5076 gnd.n3118 gnd.n1854 240.244
R5077 gnd.n3162 gnd.n1854 240.244
R5078 gnd.n3162 gnd.n1848 240.244
R5079 gnd.n3172 gnd.n1848 240.244
R5080 gnd.n3172 gnd.n1849 240.244
R5081 gnd.n3166 gnd.n1849 240.244
R5082 gnd.n3166 gnd.n1817 240.244
R5083 gnd.n3250 gnd.n1817 240.244
R5084 gnd.n3250 gnd.n1811 240.244
R5085 gnd.n3257 gnd.n1811 240.244
R5086 gnd.n3257 gnd.n1812 240.244
R5087 gnd.n1812 gnd.n1791 240.244
R5088 gnd.n3286 gnd.n1791 240.244
R5089 gnd.n3286 gnd.n1786 240.244
R5090 gnd.n3298 gnd.n1786 240.244
R5091 gnd.n3298 gnd.n1777 240.244
R5092 gnd.n3292 gnd.n1777 240.244
R5093 gnd.n3292 gnd.n1764 240.244
R5094 gnd.n3336 gnd.n1764 240.244
R5095 gnd.n3336 gnd.n1758 240.244
R5096 gnd.n3346 gnd.n1758 240.244
R5097 gnd.n3346 gnd.n1759 240.244
R5098 gnd.n3340 gnd.n1759 240.244
R5099 gnd.n3340 gnd.n1730 240.244
R5100 gnd.n3407 gnd.n1730 240.244
R5101 gnd.n3407 gnd.n1724 240.244
R5102 gnd.n3414 gnd.n1724 240.244
R5103 gnd.n3414 gnd.n1725 240.244
R5104 gnd.n1725 gnd.n1638 240.244
R5105 gnd.n3555 gnd.n1638 240.244
R5106 gnd.n3555 gnd.n1634 240.244
R5107 gnd.n3561 gnd.n1634 240.244
R5108 gnd.n3561 gnd.n1625 240.244
R5109 gnd.n3577 gnd.n1625 240.244
R5110 gnd.n3577 gnd.n1621 240.244
R5111 gnd.n3583 gnd.n1621 240.244
R5112 gnd.n3583 gnd.n1614 240.244
R5113 gnd.n3597 gnd.n1614 240.244
R5114 gnd.n3597 gnd.n1610 240.244
R5115 gnd.n3603 gnd.n1610 240.244
R5116 gnd.n3603 gnd.n1601 240.244
R5117 gnd.n3617 gnd.n1601 240.244
R5118 gnd.n3617 gnd.n1597 240.244
R5119 gnd.n3623 gnd.n1597 240.244
R5120 gnd.n3623 gnd.n1588 240.244
R5121 gnd.n3637 gnd.n1588 240.244
R5122 gnd.n3637 gnd.n1583 240.244
R5123 gnd.n3644 gnd.n1583 240.244
R5124 gnd.n3644 gnd.n1573 240.244
R5125 gnd.n1573 gnd.n455 240.244
R5126 gnd.n6356 gnd.n455 240.244
R5127 gnd.n465 gnd.n464 240.244
R5128 gnd.n472 gnd.n468 240.244
R5129 gnd.n6342 gnd.n6341 240.244
R5130 gnd.n393 gnd.n392 240.244
R5131 gnd.n475 gnd.n394 240.244
R5132 gnd.n404 gnd.n403 240.244
R5133 gnd.n477 gnd.n413 240.244
R5134 gnd.n480 gnd.n414 240.244
R5135 gnd.n422 gnd.n421 240.244
R5136 gnd.n482 gnd.n431 240.244
R5137 gnd.n485 gnd.n432 240.244
R5138 gnd.n440 gnd.n439 240.244
R5139 gnd.n487 gnd.n440 240.244
R5140 gnd.n451 gnd.n450 240.244
R5141 gnd.n1455 gnd.n1454 240.132
R5142 gnd.n1661 gnd.n1660 240.132
R5143 gnd.n5774 gnd.n835 225.874
R5144 gnd.n5782 gnd.n835 225.874
R5145 gnd.n5783 gnd.n5782 225.874
R5146 gnd.n5784 gnd.n5783 225.874
R5147 gnd.n5784 gnd.n829 225.874
R5148 gnd.n5792 gnd.n829 225.874
R5149 gnd.n5793 gnd.n5792 225.874
R5150 gnd.n5794 gnd.n5793 225.874
R5151 gnd.n5794 gnd.n823 225.874
R5152 gnd.n5802 gnd.n823 225.874
R5153 gnd.n5803 gnd.n5802 225.874
R5154 gnd.n5804 gnd.n5803 225.874
R5155 gnd.n5804 gnd.n817 225.874
R5156 gnd.n5812 gnd.n817 225.874
R5157 gnd.n5813 gnd.n5812 225.874
R5158 gnd.n5814 gnd.n5813 225.874
R5159 gnd.n5814 gnd.n811 225.874
R5160 gnd.n5822 gnd.n811 225.874
R5161 gnd.n5823 gnd.n5822 225.874
R5162 gnd.n5824 gnd.n5823 225.874
R5163 gnd.n5824 gnd.n805 225.874
R5164 gnd.n5832 gnd.n805 225.874
R5165 gnd.n5833 gnd.n5832 225.874
R5166 gnd.n5834 gnd.n5833 225.874
R5167 gnd.n5834 gnd.n799 225.874
R5168 gnd.n5842 gnd.n799 225.874
R5169 gnd.n5843 gnd.n5842 225.874
R5170 gnd.n5844 gnd.n5843 225.874
R5171 gnd.n5844 gnd.n793 225.874
R5172 gnd.n5852 gnd.n793 225.874
R5173 gnd.n5853 gnd.n5852 225.874
R5174 gnd.n5854 gnd.n5853 225.874
R5175 gnd.n5854 gnd.n787 225.874
R5176 gnd.n5862 gnd.n787 225.874
R5177 gnd.n5863 gnd.n5862 225.874
R5178 gnd.n5864 gnd.n5863 225.874
R5179 gnd.n5864 gnd.n781 225.874
R5180 gnd.n5872 gnd.n781 225.874
R5181 gnd.n5873 gnd.n5872 225.874
R5182 gnd.n5874 gnd.n5873 225.874
R5183 gnd.n5874 gnd.n775 225.874
R5184 gnd.n5882 gnd.n775 225.874
R5185 gnd.n5883 gnd.n5882 225.874
R5186 gnd.n5884 gnd.n5883 225.874
R5187 gnd.n5884 gnd.n769 225.874
R5188 gnd.n5892 gnd.n769 225.874
R5189 gnd.n5893 gnd.n5892 225.874
R5190 gnd.n5894 gnd.n5893 225.874
R5191 gnd.n5894 gnd.n763 225.874
R5192 gnd.n5902 gnd.n763 225.874
R5193 gnd.n5903 gnd.n5902 225.874
R5194 gnd.n5904 gnd.n5903 225.874
R5195 gnd.n5904 gnd.n757 225.874
R5196 gnd.n5912 gnd.n757 225.874
R5197 gnd.n5913 gnd.n5912 225.874
R5198 gnd.n5914 gnd.n5913 225.874
R5199 gnd.n5914 gnd.n751 225.874
R5200 gnd.n5922 gnd.n751 225.874
R5201 gnd.n5923 gnd.n5922 225.874
R5202 gnd.n5924 gnd.n5923 225.874
R5203 gnd.n5924 gnd.n745 225.874
R5204 gnd.n5932 gnd.n745 225.874
R5205 gnd.n5933 gnd.n5932 225.874
R5206 gnd.n5934 gnd.n5933 225.874
R5207 gnd.n5934 gnd.n739 225.874
R5208 gnd.n5942 gnd.n739 225.874
R5209 gnd.n5943 gnd.n5942 225.874
R5210 gnd.n5944 gnd.n5943 225.874
R5211 gnd.n5944 gnd.n733 225.874
R5212 gnd.n5952 gnd.n733 225.874
R5213 gnd.n5953 gnd.n5952 225.874
R5214 gnd.n5954 gnd.n5953 225.874
R5215 gnd.n5954 gnd.n727 225.874
R5216 gnd.n5962 gnd.n727 225.874
R5217 gnd.n5963 gnd.n5962 225.874
R5218 gnd.n5964 gnd.n5963 225.874
R5219 gnd.n5964 gnd.n721 225.874
R5220 gnd.n5972 gnd.n721 225.874
R5221 gnd.n5973 gnd.n5972 225.874
R5222 gnd.n5974 gnd.n5973 225.874
R5223 gnd.n5974 gnd.n715 225.874
R5224 gnd.n5982 gnd.n715 225.874
R5225 gnd.n5983 gnd.n5982 225.874
R5226 gnd.n5984 gnd.n5983 225.874
R5227 gnd.n5984 gnd.n709 225.874
R5228 gnd.n5992 gnd.n709 225.874
R5229 gnd.n5993 gnd.n5992 225.874
R5230 gnd.n5994 gnd.n5993 225.874
R5231 gnd.n5994 gnd.n703 225.874
R5232 gnd.n6002 gnd.n703 225.874
R5233 gnd.n6003 gnd.n6002 225.874
R5234 gnd.n6004 gnd.n6003 225.874
R5235 gnd.n6004 gnd.n697 225.874
R5236 gnd.n6012 gnd.n697 225.874
R5237 gnd.n6013 gnd.n6012 225.874
R5238 gnd.n6014 gnd.n6013 225.874
R5239 gnd.n6014 gnd.n691 225.874
R5240 gnd.n6022 gnd.n691 225.874
R5241 gnd.n6023 gnd.n6022 225.874
R5242 gnd.n6024 gnd.n6023 225.874
R5243 gnd.n6024 gnd.n685 225.874
R5244 gnd.n6032 gnd.n685 225.874
R5245 gnd.n6033 gnd.n6032 225.874
R5246 gnd.n6034 gnd.n6033 225.874
R5247 gnd.n6034 gnd.n679 225.874
R5248 gnd.n6042 gnd.n679 225.874
R5249 gnd.n6043 gnd.n6042 225.874
R5250 gnd.n6044 gnd.n6043 225.874
R5251 gnd.n6044 gnd.n673 225.874
R5252 gnd.n6052 gnd.n673 225.874
R5253 gnd.n6053 gnd.n6052 225.874
R5254 gnd.n6054 gnd.n6053 225.874
R5255 gnd.n6054 gnd.n667 225.874
R5256 gnd.n6062 gnd.n667 225.874
R5257 gnd.n6063 gnd.n6062 225.874
R5258 gnd.n6064 gnd.n6063 225.874
R5259 gnd.n6064 gnd.n661 225.874
R5260 gnd.n6072 gnd.n661 225.874
R5261 gnd.n6073 gnd.n6072 225.874
R5262 gnd.n6074 gnd.n6073 225.874
R5263 gnd.n6074 gnd.n655 225.874
R5264 gnd.n6082 gnd.n655 225.874
R5265 gnd.n6083 gnd.n6082 225.874
R5266 gnd.n6084 gnd.n6083 225.874
R5267 gnd.n6084 gnd.n649 225.874
R5268 gnd.n6092 gnd.n649 225.874
R5269 gnd.n6093 gnd.n6092 225.874
R5270 gnd.n6094 gnd.n6093 225.874
R5271 gnd.n4698 gnd.t304 224.174
R5272 gnd.n4208 gnd.t220 224.174
R5273 gnd.n352 gnd.n296 199.319
R5274 gnd.n352 gnd.n297 199.319
R5275 gnd.n1407 gnd.n1367 199.319
R5276 gnd.n1407 gnd.n1366 199.319
R5277 gnd.n1456 gnd.n1453 186.49
R5278 gnd.n1662 gnd.n1659 186.49
R5279 gnd.n5473 gnd.n5472 185
R5280 gnd.n5471 gnd.n5470 185
R5281 gnd.n5450 gnd.n5449 185
R5282 gnd.n5465 gnd.n5464 185
R5283 gnd.n5463 gnd.n5462 185
R5284 gnd.n5454 gnd.n5453 185
R5285 gnd.n5457 gnd.n5456 185
R5286 gnd.n5441 gnd.n5440 185
R5287 gnd.n5439 gnd.n5438 185
R5288 gnd.n5418 gnd.n5417 185
R5289 gnd.n5433 gnd.n5432 185
R5290 gnd.n5431 gnd.n5430 185
R5291 gnd.n5422 gnd.n5421 185
R5292 gnd.n5425 gnd.n5424 185
R5293 gnd.n5409 gnd.n5408 185
R5294 gnd.n5407 gnd.n5406 185
R5295 gnd.n5386 gnd.n5385 185
R5296 gnd.n5401 gnd.n5400 185
R5297 gnd.n5399 gnd.n5398 185
R5298 gnd.n5390 gnd.n5389 185
R5299 gnd.n5393 gnd.n5392 185
R5300 gnd.n5378 gnd.n5377 185
R5301 gnd.n5376 gnd.n5375 185
R5302 gnd.n5355 gnd.n5354 185
R5303 gnd.n5370 gnd.n5369 185
R5304 gnd.n5368 gnd.n5367 185
R5305 gnd.n5359 gnd.n5358 185
R5306 gnd.n5362 gnd.n5361 185
R5307 gnd.n5346 gnd.n5345 185
R5308 gnd.n5344 gnd.n5343 185
R5309 gnd.n5323 gnd.n5322 185
R5310 gnd.n5338 gnd.n5337 185
R5311 gnd.n5336 gnd.n5335 185
R5312 gnd.n5327 gnd.n5326 185
R5313 gnd.n5330 gnd.n5329 185
R5314 gnd.n5314 gnd.n5313 185
R5315 gnd.n5312 gnd.n5311 185
R5316 gnd.n5291 gnd.n5290 185
R5317 gnd.n5306 gnd.n5305 185
R5318 gnd.n5304 gnd.n5303 185
R5319 gnd.n5295 gnd.n5294 185
R5320 gnd.n5298 gnd.n5297 185
R5321 gnd.n5282 gnd.n5281 185
R5322 gnd.n5280 gnd.n5279 185
R5323 gnd.n5259 gnd.n5258 185
R5324 gnd.n5274 gnd.n5273 185
R5325 gnd.n5272 gnd.n5271 185
R5326 gnd.n5263 gnd.n5262 185
R5327 gnd.n5266 gnd.n5265 185
R5328 gnd.n5251 gnd.n5250 185
R5329 gnd.n5249 gnd.n5248 185
R5330 gnd.n5228 gnd.n5227 185
R5331 gnd.n5243 gnd.n5242 185
R5332 gnd.n5241 gnd.n5240 185
R5333 gnd.n5232 gnd.n5231 185
R5334 gnd.n5235 gnd.n5234 185
R5335 gnd.n4699 gnd.t303 178.987
R5336 gnd.n4209 gnd.t221 178.987
R5337 gnd.n6481 gnd.n351 171.457
R5338 gnd.n3853 gnd.n3852 171.457
R5339 gnd.n1 gnd.t83 170.774
R5340 gnd.n9 gnd.t125 170.103
R5341 gnd.n8 gnd.t62 170.103
R5342 gnd.n7 gnd.t150 170.103
R5343 gnd.n6 gnd.t12 170.103
R5344 gnd.n5 gnd.t103 170.103
R5345 gnd.n4 gnd.t15 170.103
R5346 gnd.n3 gnd.t109 170.103
R5347 gnd.n2 gnd.t203 170.103
R5348 gnd.n1 gnd.t172 170.103
R5349 gnd.n3537 gnd.n3536 163.367
R5350 gnd.n3534 gnd.n1673 163.367
R5351 gnd.n3530 gnd.n3529 163.367
R5352 gnd.n3527 gnd.n1676 163.367
R5353 gnd.n3523 gnd.n3522 163.367
R5354 gnd.n3520 gnd.n1679 163.367
R5355 gnd.n3516 gnd.n3515 163.367
R5356 gnd.n3513 gnd.n1682 163.367
R5357 gnd.n3509 gnd.n3508 163.367
R5358 gnd.n3506 gnd.n1685 163.367
R5359 gnd.n3502 gnd.n3501 163.367
R5360 gnd.n3499 gnd.n1688 163.367
R5361 gnd.n3495 gnd.n3494 163.367
R5362 gnd.n3492 gnd.n1691 163.367
R5363 gnd.n3487 gnd.n3486 163.367
R5364 gnd.n3484 gnd.n3482 163.367
R5365 gnd.n3479 gnd.n3478 163.367
R5366 gnd.n3476 gnd.n1697 163.367
R5367 gnd.n3471 gnd.n3470 163.367
R5368 gnd.n3468 gnd.n1702 163.367
R5369 gnd.n3464 gnd.n3463 163.367
R5370 gnd.n3461 gnd.n1705 163.367
R5371 gnd.n3457 gnd.n3456 163.367
R5372 gnd.n3454 gnd.n1708 163.367
R5373 gnd.n3450 gnd.n3449 163.367
R5374 gnd.n3447 gnd.n1711 163.367
R5375 gnd.n3443 gnd.n3442 163.367
R5376 gnd.n3440 gnd.n1714 163.367
R5377 gnd.n3436 gnd.n3435 163.367
R5378 gnd.n3433 gnd.n1717 163.367
R5379 gnd.n3429 gnd.n3428 163.367
R5380 gnd.n3426 gnd.n1720 163.367
R5381 gnd.n2874 gnd.n1472 163.367
R5382 gnd.n2890 gnd.n1472 163.367
R5383 gnd.n2890 gnd.n1993 163.367
R5384 gnd.n2914 gnd.n1993 163.367
R5385 gnd.n2914 gnd.n1990 163.367
R5386 gnd.n2910 gnd.n1990 163.367
R5387 gnd.n2910 gnd.n1983 163.367
R5388 gnd.n2905 gnd.n1983 163.367
R5389 gnd.n2905 gnd.n1977 163.367
R5390 gnd.n2902 gnd.n1977 163.367
R5391 gnd.n2902 gnd.n1970 163.367
R5392 gnd.n2897 gnd.n1970 163.367
R5393 gnd.n2897 gnd.n1963 163.367
R5394 gnd.n2894 gnd.n1963 163.367
R5395 gnd.n2894 gnd.n1956 163.367
R5396 gnd.n1956 gnd.n1945 163.367
R5397 gnd.n2997 gnd.n1945 163.367
R5398 gnd.n2997 gnd.n1939 163.367
R5399 gnd.n3001 gnd.n1939 163.367
R5400 gnd.n3001 gnd.n1931 163.367
R5401 gnd.n3021 gnd.n1931 163.367
R5402 gnd.n3021 gnd.n1929 163.367
R5403 gnd.n3054 gnd.n1929 163.367
R5404 gnd.n3054 gnd.n1922 163.367
R5405 gnd.n3050 gnd.n1922 163.367
R5406 gnd.n3050 gnd.n3047 163.367
R5407 gnd.n3047 gnd.n3046 163.367
R5408 gnd.n3046 gnd.n1906 163.367
R5409 gnd.n3042 gnd.n1906 163.367
R5410 gnd.n3042 gnd.n1900 163.367
R5411 gnd.n3039 gnd.n1900 163.367
R5412 gnd.n3039 gnd.n1892 163.367
R5413 gnd.n3034 gnd.n1892 163.367
R5414 gnd.n3034 gnd.n1885 163.367
R5415 gnd.n3031 gnd.n1885 163.367
R5416 gnd.n3031 gnd.n1877 163.367
R5417 gnd.n3026 gnd.n1877 163.367
R5418 gnd.n3026 gnd.n1869 163.367
R5419 gnd.n1869 gnd.n1858 163.367
R5420 gnd.n3149 gnd.n1858 163.367
R5421 gnd.n3149 gnd.n1856 163.367
R5422 gnd.n3159 gnd.n1856 163.367
R5423 gnd.n3159 gnd.n1843 163.367
R5424 gnd.n3155 gnd.n1843 163.367
R5425 gnd.n3155 gnd.n1837 163.367
R5426 gnd.n3191 gnd.n1837 163.367
R5427 gnd.n3191 gnd.n1835 163.367
R5428 gnd.n3227 gnd.n1835 163.367
R5429 gnd.n3227 gnd.n1827 163.367
R5430 gnd.n3223 gnd.n1827 163.367
R5431 gnd.n3223 gnd.n3220 163.367
R5432 gnd.n3220 gnd.n3219 163.367
R5433 gnd.n3219 gnd.n1810 163.367
R5434 gnd.n3215 gnd.n1810 163.367
R5435 gnd.n3215 gnd.n1806 163.367
R5436 gnd.n3212 gnd.n1806 163.367
R5437 gnd.n3212 gnd.n1798 163.367
R5438 gnd.n3204 gnd.n1798 163.367
R5439 gnd.n3204 gnd.n1793 163.367
R5440 gnd.n3201 gnd.n1793 163.367
R5441 gnd.n3201 gnd.n1785 163.367
R5442 gnd.n3196 gnd.n1785 163.367
R5443 gnd.n3196 gnd.n1778 163.367
R5444 gnd.n1778 gnd.n1768 163.367
R5445 gnd.n3323 gnd.n1768 163.367
R5446 gnd.n3323 gnd.n1766 163.367
R5447 gnd.n3332 gnd.n1766 163.367
R5448 gnd.n3332 gnd.n1753 163.367
R5449 gnd.n3328 gnd.n1753 163.367
R5450 gnd.n3328 gnd.n1747 163.367
R5451 gnd.n3365 gnd.n1747 163.367
R5452 gnd.n3365 gnd.n1745 163.367
R5453 gnd.n3378 gnd.n1745 163.367
R5454 gnd.n3378 gnd.n1739 163.367
R5455 gnd.n3374 gnd.n1739 163.367
R5456 gnd.n3374 gnd.n3371 163.367
R5457 gnd.n3371 gnd.n3370 163.367
R5458 gnd.n3370 gnd.n1722 163.367
R5459 gnd.n3418 gnd.n1722 163.367
R5460 gnd.n3418 gnd.n1645 163.367
R5461 gnd.n1447 gnd.n1446 163.367
R5462 gnd.n3842 gnd.n1446 163.367
R5463 gnd.n3840 gnd.n3839 163.367
R5464 gnd.n3836 gnd.n3835 163.367
R5465 gnd.n3832 gnd.n3831 163.367
R5466 gnd.n3828 gnd.n3827 163.367
R5467 gnd.n3824 gnd.n3823 163.367
R5468 gnd.n3820 gnd.n3819 163.367
R5469 gnd.n3816 gnd.n3815 163.367
R5470 gnd.n3812 gnd.n3811 163.367
R5471 gnd.n3808 gnd.n3807 163.367
R5472 gnd.n3804 gnd.n3803 163.367
R5473 gnd.n3800 gnd.n3799 163.367
R5474 gnd.n3796 gnd.n3795 163.367
R5475 gnd.n3792 gnd.n3791 163.367
R5476 gnd.n3788 gnd.n3787 163.367
R5477 gnd.n3851 gnd.n1412 163.367
R5478 gnd.n2813 gnd.n2812 163.367
R5479 gnd.n2818 gnd.n2817 163.367
R5480 gnd.n2822 gnd.n2821 163.367
R5481 gnd.n2826 gnd.n2825 163.367
R5482 gnd.n2830 gnd.n2829 163.367
R5483 gnd.n2834 gnd.n2833 163.367
R5484 gnd.n2838 gnd.n2837 163.367
R5485 gnd.n2842 gnd.n2841 163.367
R5486 gnd.n2846 gnd.n2845 163.367
R5487 gnd.n2850 gnd.n2849 163.367
R5488 gnd.n2854 gnd.n2853 163.367
R5489 gnd.n2858 gnd.n2857 163.367
R5490 gnd.n2862 gnd.n2861 163.367
R5491 gnd.n2866 gnd.n2865 163.367
R5492 gnd.n2870 gnd.n2869 163.367
R5493 gnd.n3780 gnd.n1448 163.367
R5494 gnd.n3780 gnd.n1470 163.367
R5495 gnd.n2919 gnd.n1470 163.367
R5496 gnd.n2919 gnd.n1992 163.367
R5497 gnd.n2923 gnd.n1992 163.367
R5498 gnd.n2923 gnd.n1981 163.367
R5499 gnd.n2937 gnd.n1981 163.367
R5500 gnd.n2937 gnd.n1979 163.367
R5501 gnd.n2941 gnd.n1979 163.367
R5502 gnd.n2941 gnd.n1968 163.367
R5503 gnd.n2954 gnd.n1968 163.367
R5504 gnd.n2954 gnd.n1965 163.367
R5505 gnd.n2964 gnd.n1965 163.367
R5506 gnd.n2964 gnd.n1966 163.367
R5507 gnd.n1966 gnd.n1955 163.367
R5508 gnd.n2959 gnd.n1955 163.367
R5509 gnd.n2959 gnd.n1941 163.367
R5510 gnd.n3009 gnd.n1941 163.367
R5511 gnd.n3009 gnd.n1942 163.367
R5512 gnd.n3005 gnd.n1942 163.367
R5513 gnd.n3005 gnd.n1927 163.367
R5514 gnd.n3058 gnd.n1927 163.367
R5515 gnd.n3058 gnd.n1924 163.367
R5516 gnd.n3065 gnd.n1924 163.367
R5517 gnd.n3065 gnd.n1925 163.367
R5518 gnd.n3061 gnd.n1925 163.367
R5519 gnd.n3061 gnd.n1904 163.367
R5520 gnd.n3089 gnd.n1904 163.367
R5521 gnd.n3089 gnd.n1902 163.367
R5522 gnd.n3093 gnd.n1902 163.367
R5523 gnd.n3093 gnd.n1889 163.367
R5524 gnd.n3107 gnd.n1889 163.367
R5525 gnd.n3107 gnd.n1887 163.367
R5526 gnd.n3111 gnd.n1887 163.367
R5527 gnd.n3111 gnd.n1875 163.367
R5528 gnd.n3127 gnd.n1875 163.367
R5529 gnd.n3127 gnd.n1871 163.367
R5530 gnd.n3136 gnd.n1871 163.367
R5531 gnd.n3136 gnd.n1873 163.367
R5532 gnd.n1873 gnd.n1860 163.367
R5533 gnd.n3131 gnd.n1860 163.367
R5534 gnd.n3131 gnd.n1844 163.367
R5535 gnd.n3179 gnd.n1844 163.367
R5536 gnd.n3179 gnd.n1845 163.367
R5537 gnd.n3175 gnd.n1845 163.367
R5538 gnd.n3175 gnd.n1833 163.367
R5539 gnd.n3231 gnd.n1833 163.367
R5540 gnd.n3231 gnd.n1830 163.367
R5541 gnd.n3238 gnd.n1830 163.367
R5542 gnd.n3238 gnd.n1831 163.367
R5543 gnd.n3234 gnd.n1831 163.367
R5544 gnd.n3234 gnd.n1809 163.367
R5545 gnd.n3261 gnd.n1809 163.367
R5546 gnd.n3261 gnd.n1807 163.367
R5547 gnd.n3265 gnd.n1807 163.367
R5548 gnd.n3265 gnd.n1797 163.367
R5549 gnd.n3279 gnd.n1797 163.367
R5550 gnd.n3279 gnd.n1795 163.367
R5551 gnd.n3283 gnd.n1795 163.367
R5552 gnd.n3283 gnd.n1783 163.367
R5553 gnd.n3302 gnd.n1783 163.367
R5554 gnd.n3302 gnd.n1780 163.367
R5555 gnd.n3311 gnd.n1780 163.367
R5556 gnd.n3311 gnd.n1781 163.367
R5557 gnd.n1781 gnd.n1769 163.367
R5558 gnd.n3306 gnd.n1769 163.367
R5559 gnd.n3306 gnd.n1755 163.367
R5560 gnd.n3353 gnd.n1755 163.367
R5561 gnd.n3353 gnd.n1756 163.367
R5562 gnd.n3349 gnd.n1756 163.367
R5563 gnd.n3349 gnd.n1743 163.367
R5564 gnd.n3382 gnd.n1743 163.367
R5565 gnd.n3382 gnd.n1740 163.367
R5566 gnd.n3395 gnd.n1740 163.367
R5567 gnd.n3395 gnd.n1741 163.367
R5568 gnd.n3391 gnd.n1741 163.367
R5569 gnd.n3391 gnd.n3390 163.367
R5570 gnd.n3390 gnd.n3389 163.367
R5571 gnd.n3389 gnd.n1647 163.367
R5572 gnd.n3542 gnd.n1647 163.367
R5573 gnd.n1668 gnd.n1667 156.462
R5574 gnd.n5413 gnd.n5381 153.042
R5575 gnd.n5477 gnd.n5476 152.079
R5576 gnd.n5445 gnd.n5444 152.079
R5577 gnd.n5413 gnd.n5412 152.079
R5578 gnd.n1461 gnd.n1460 152
R5579 gnd.n1462 gnd.n1451 152
R5580 gnd.n1464 gnd.n1463 152
R5581 gnd.n1466 gnd.n1449 152
R5582 gnd.n1468 gnd.n1467 152
R5583 gnd.n1666 gnd.n1650 152
R5584 gnd.n1658 gnd.n1651 152
R5585 gnd.n1657 gnd.n1656 152
R5586 gnd.n1655 gnd.n1652 152
R5587 gnd.n1653 gnd.t242 150.546
R5588 gnd.t93 gnd.n5455 147.661
R5589 gnd.t3 gnd.n5423 147.661
R5590 gnd.t138 gnd.n5391 147.661
R5591 gnd.t158 gnd.n5360 147.661
R5592 gnd.t39 gnd.n5328 147.661
R5593 gnd.t152 gnd.n5296 147.661
R5594 gnd.t85 gnd.n5264 147.661
R5595 gnd.t140 gnd.n5233 147.661
R5596 gnd.n3481 gnd.n3480 143.351
R5597 gnd.n1428 gnd.n1411 143.351
R5598 gnd.n3850 gnd.n1411 143.351
R5599 gnd.n1458 gnd.t298 130.484
R5600 gnd.n1467 gnd.t211 126.766
R5601 gnd.n1465 gnd.t289 126.766
R5602 gnd.n1451 gnd.t311 126.766
R5603 gnd.n1459 gnd.t245 126.766
R5604 gnd.n1654 gnd.t313 126.766
R5605 gnd.n1656 gnd.t265 126.766
R5606 gnd.n1665 gnd.t208 126.766
R5607 gnd.n1667 gnd.t280 126.766
R5608 gnd.n5472 gnd.n5471 104.615
R5609 gnd.n5471 gnd.n5449 104.615
R5610 gnd.n5464 gnd.n5449 104.615
R5611 gnd.n5464 gnd.n5463 104.615
R5612 gnd.n5463 gnd.n5453 104.615
R5613 gnd.n5456 gnd.n5453 104.615
R5614 gnd.n5440 gnd.n5439 104.615
R5615 gnd.n5439 gnd.n5417 104.615
R5616 gnd.n5432 gnd.n5417 104.615
R5617 gnd.n5432 gnd.n5431 104.615
R5618 gnd.n5431 gnd.n5421 104.615
R5619 gnd.n5424 gnd.n5421 104.615
R5620 gnd.n5408 gnd.n5407 104.615
R5621 gnd.n5407 gnd.n5385 104.615
R5622 gnd.n5400 gnd.n5385 104.615
R5623 gnd.n5400 gnd.n5399 104.615
R5624 gnd.n5399 gnd.n5389 104.615
R5625 gnd.n5392 gnd.n5389 104.615
R5626 gnd.n5377 gnd.n5376 104.615
R5627 gnd.n5376 gnd.n5354 104.615
R5628 gnd.n5369 gnd.n5354 104.615
R5629 gnd.n5369 gnd.n5368 104.615
R5630 gnd.n5368 gnd.n5358 104.615
R5631 gnd.n5361 gnd.n5358 104.615
R5632 gnd.n5345 gnd.n5344 104.615
R5633 gnd.n5344 gnd.n5322 104.615
R5634 gnd.n5337 gnd.n5322 104.615
R5635 gnd.n5337 gnd.n5336 104.615
R5636 gnd.n5336 gnd.n5326 104.615
R5637 gnd.n5329 gnd.n5326 104.615
R5638 gnd.n5313 gnd.n5312 104.615
R5639 gnd.n5312 gnd.n5290 104.615
R5640 gnd.n5305 gnd.n5290 104.615
R5641 gnd.n5305 gnd.n5304 104.615
R5642 gnd.n5304 gnd.n5294 104.615
R5643 gnd.n5297 gnd.n5294 104.615
R5644 gnd.n5281 gnd.n5280 104.615
R5645 gnd.n5280 gnd.n5258 104.615
R5646 gnd.n5273 gnd.n5258 104.615
R5647 gnd.n5273 gnd.n5272 104.615
R5648 gnd.n5272 gnd.n5262 104.615
R5649 gnd.n5265 gnd.n5262 104.615
R5650 gnd.n5250 gnd.n5249 104.615
R5651 gnd.n5249 gnd.n5227 104.615
R5652 gnd.n5242 gnd.n5227 104.615
R5653 gnd.n5242 gnd.n5241 104.615
R5654 gnd.n5241 gnd.n5231 104.615
R5655 gnd.n5234 gnd.n5231 104.615
R5656 gnd.n4624 gnd.t264 100.632
R5657 gnd.n4182 gnd.t321 100.632
R5658 gnd.n7033 gnd.n6864 99.6594
R5659 gnd.n7031 gnd.n6863 99.6594
R5660 gnd.n7027 gnd.n6862 99.6594
R5661 gnd.n7023 gnd.n6861 99.6594
R5662 gnd.n7019 gnd.n6860 99.6594
R5663 gnd.n7015 gnd.n6859 99.6594
R5664 gnd.n7011 gnd.n6858 99.6594
R5665 gnd.n7007 gnd.n6857 99.6594
R5666 gnd.n7000 gnd.n6856 99.6594
R5667 gnd.n6996 gnd.n6855 99.6594
R5668 gnd.n6992 gnd.n6854 99.6594
R5669 gnd.n6988 gnd.n6853 99.6594
R5670 gnd.n6984 gnd.n6852 99.6594
R5671 gnd.n6980 gnd.n6851 99.6594
R5672 gnd.n6976 gnd.n6850 99.6594
R5673 gnd.n6972 gnd.n6849 99.6594
R5674 gnd.n6968 gnd.n6848 99.6594
R5675 gnd.n6964 gnd.n6847 99.6594
R5676 gnd.n6956 gnd.n6846 99.6594
R5677 gnd.n6954 gnd.n6845 99.6594
R5678 gnd.n6950 gnd.n6844 99.6594
R5679 gnd.n6946 gnd.n6843 99.6594
R5680 gnd.n6942 gnd.n6842 99.6594
R5681 gnd.n6938 gnd.n6841 99.6594
R5682 gnd.n6934 gnd.n6840 99.6594
R5683 gnd.n6930 gnd.n6839 99.6594
R5684 gnd.n6926 gnd.n6838 99.6594
R5685 gnd.n6922 gnd.n6837 99.6594
R5686 gnd.n7045 gnd.n7043 99.6594
R5687 gnd.n6532 gnd.n6531 99.6594
R5688 gnd.n324 gnd.n285 99.6594
R5689 gnd.n6524 gnd.n286 99.6594
R5690 gnd.n6520 gnd.n287 99.6594
R5691 gnd.n6516 gnd.n288 99.6594
R5692 gnd.n6512 gnd.n289 99.6594
R5693 gnd.n6508 gnd.n290 99.6594
R5694 gnd.n6504 gnd.n291 99.6594
R5695 gnd.n6500 gnd.n292 99.6594
R5696 gnd.n6495 gnd.n293 99.6594
R5697 gnd.n6491 gnd.n294 99.6594
R5698 gnd.n6487 gnd.n295 99.6594
R5699 gnd.n6483 gnd.n296 99.6594
R5700 gnd.n6478 gnd.n298 99.6594
R5701 gnd.n6474 gnd.n299 99.6594
R5702 gnd.n6470 gnd.n300 99.6594
R5703 gnd.n6466 gnd.n301 99.6594
R5704 gnd.n6462 gnd.n302 99.6594
R5705 gnd.n6458 gnd.n303 99.6594
R5706 gnd.n6454 gnd.n304 99.6594
R5707 gnd.n6450 gnd.n305 99.6594
R5708 gnd.n6446 gnd.n306 99.6594
R5709 gnd.n6442 gnd.n307 99.6594
R5710 gnd.n6438 gnd.n308 99.6594
R5711 gnd.n6434 gnd.n309 99.6594
R5712 gnd.n6430 gnd.n310 99.6594
R5713 gnd.n6426 gnd.n311 99.6594
R5714 gnd.n6422 gnd.n312 99.6594
R5715 gnd.n3902 gnd.n3901 99.6594
R5716 gnd.n3897 gnd.n1378 99.6594
R5717 gnd.n3893 gnd.n1377 99.6594
R5718 gnd.n3889 gnd.n1376 99.6594
R5719 gnd.n3885 gnd.n1375 99.6594
R5720 gnd.n3881 gnd.n1374 99.6594
R5721 gnd.n3877 gnd.n1373 99.6594
R5722 gnd.n3873 gnd.n1372 99.6594
R5723 gnd.n3868 gnd.n1371 99.6594
R5724 gnd.n3864 gnd.n1370 99.6594
R5725 gnd.n3860 gnd.n1369 99.6594
R5726 gnd.n3856 gnd.n1368 99.6594
R5727 gnd.n2218 gnd.n1366 99.6594
R5728 gnd.n2225 gnd.n1365 99.6594
R5729 gnd.n2229 gnd.n1364 99.6594
R5730 gnd.n2235 gnd.n1363 99.6594
R5731 gnd.n2239 gnd.n1362 99.6594
R5732 gnd.n2245 gnd.n1361 99.6594
R5733 gnd.n2249 gnd.n1360 99.6594
R5734 gnd.n2255 gnd.n1359 99.6594
R5735 gnd.n2259 gnd.n1358 99.6594
R5736 gnd.n2265 gnd.n1357 99.6594
R5737 gnd.n2269 gnd.n1356 99.6594
R5738 gnd.n2275 gnd.n1355 99.6594
R5739 gnd.n2279 gnd.n1354 99.6594
R5740 gnd.n2285 gnd.n1353 99.6594
R5741 gnd.n2289 gnd.n1352 99.6594
R5742 gnd.n2295 gnd.n1351 99.6594
R5743 gnd.n4156 gnd.n4155 99.6594
R5744 gnd.n4150 gnd.n1023 99.6594
R5745 gnd.n4147 gnd.n1024 99.6594
R5746 gnd.n4143 gnd.n1025 99.6594
R5747 gnd.n4139 gnd.n1026 99.6594
R5748 gnd.n4135 gnd.n1027 99.6594
R5749 gnd.n4131 gnd.n1028 99.6594
R5750 gnd.n4127 gnd.n1029 99.6594
R5751 gnd.n4123 gnd.n1030 99.6594
R5752 gnd.n4118 gnd.n1031 99.6594
R5753 gnd.n4114 gnd.n1032 99.6594
R5754 gnd.n4110 gnd.n1033 99.6594
R5755 gnd.n4106 gnd.n1034 99.6594
R5756 gnd.n4102 gnd.n1035 99.6594
R5757 gnd.n4098 gnd.n1036 99.6594
R5758 gnd.n4094 gnd.n1037 99.6594
R5759 gnd.n4090 gnd.n1038 99.6594
R5760 gnd.n4086 gnd.n1039 99.6594
R5761 gnd.n4082 gnd.n1040 99.6594
R5762 gnd.n4078 gnd.n1041 99.6594
R5763 gnd.n4074 gnd.n1042 99.6594
R5764 gnd.n4070 gnd.n1043 99.6594
R5765 gnd.n4066 gnd.n1044 99.6594
R5766 gnd.n4062 gnd.n1045 99.6594
R5767 gnd.n4058 gnd.n1046 99.6594
R5768 gnd.n4054 gnd.n1047 99.6594
R5769 gnd.n4050 gnd.n1048 99.6594
R5770 gnd.n4046 gnd.n1049 99.6594
R5771 gnd.n4042 gnd.n1050 99.6594
R5772 gnd.n5595 gnd.n4165 99.6594
R5773 gnd.n5593 gnd.n4164 99.6594
R5774 gnd.n5589 gnd.n4163 99.6594
R5775 gnd.n5585 gnd.n4162 99.6594
R5776 gnd.n5581 gnd.n4161 99.6594
R5777 gnd.n5577 gnd.n4160 99.6594
R5778 gnd.n5573 gnd.n4159 99.6594
R5779 gnd.n5505 gnd.n4158 99.6594
R5780 gnd.n4836 gnd.n4567 99.6594
R5781 gnd.n4593 gnd.n4574 99.6594
R5782 gnd.n4595 gnd.n4575 99.6594
R5783 gnd.n4603 gnd.n4576 99.6594
R5784 gnd.n4605 gnd.n4577 99.6594
R5785 gnd.n4613 gnd.n4578 99.6594
R5786 gnd.n4615 gnd.n4579 99.6594
R5787 gnd.n4623 gnd.n4580 99.6594
R5788 gnd.n6751 gnd.n6725 99.6594
R5789 gnd.n6755 gnd.n6726 99.6594
R5790 gnd.n6761 gnd.n6727 99.6594
R5791 gnd.n6765 gnd.n6728 99.6594
R5792 gnd.n6771 gnd.n6729 99.6594
R5793 gnd.n6775 gnd.n6730 99.6594
R5794 gnd.n6781 gnd.n6731 99.6594
R5795 gnd.n6784 gnd.n6732 99.6594
R5796 gnd.n6836 gnd.n6835 99.6594
R5797 gnd.n502 gnd.n313 99.6594
R5798 gnd.n400 gnd.n314 99.6594
R5799 gnd.n408 gnd.n315 99.6594
R5800 gnd.n410 gnd.n316 99.6594
R5801 gnd.n418 gnd.n317 99.6594
R5802 gnd.n426 gnd.n318 99.6594
R5803 gnd.n428 gnd.n319 99.6594
R5804 gnd.n436 gnd.n320 99.6594
R5805 gnd.n446 gnd.n321 99.6594
R5806 gnd.n5563 gnd.n1010 99.6594
R5807 gnd.n5559 gnd.n1011 99.6594
R5808 gnd.n5555 gnd.n1012 99.6594
R5809 gnd.n5551 gnd.n1013 99.6594
R5810 gnd.n5547 gnd.n1014 99.6594
R5811 gnd.n5543 gnd.n1015 99.6594
R5812 gnd.n5539 gnd.n1016 99.6594
R5813 gnd.n5535 gnd.n1017 99.6594
R5814 gnd.n5531 gnd.n1018 99.6594
R5815 gnd.n5527 gnd.n1019 99.6594
R5816 gnd.n5523 gnd.n1020 99.6594
R5817 gnd.n5519 gnd.n1021 99.6594
R5818 gnd.n5515 gnd.n1022 99.6594
R5819 gnd.n4751 gnd.n4750 99.6594
R5820 gnd.n4745 gnd.n4662 99.6594
R5821 gnd.n4742 gnd.n4663 99.6594
R5822 gnd.n4738 gnd.n4664 99.6594
R5823 gnd.n4734 gnd.n4665 99.6594
R5824 gnd.n4730 gnd.n4666 99.6594
R5825 gnd.n4726 gnd.n4667 99.6594
R5826 gnd.n4722 gnd.n4668 99.6594
R5827 gnd.n4718 gnd.n4669 99.6594
R5828 gnd.n4714 gnd.n4670 99.6594
R5829 gnd.n4710 gnd.n4671 99.6594
R5830 gnd.n4706 gnd.n4672 99.6594
R5831 gnd.n4753 gnd.n4661 99.6594
R5832 gnd.n2142 gnd.n1341 99.6594
R5833 gnd.n2152 gnd.n1342 99.6594
R5834 gnd.n2160 gnd.n1343 99.6594
R5835 gnd.n2162 gnd.n1344 99.6594
R5836 gnd.n2172 gnd.n1345 99.6594
R5837 gnd.n2180 gnd.n1346 99.6594
R5838 gnd.n2182 gnd.n1347 99.6594
R5839 gnd.n2193 gnd.n1348 99.6594
R5840 gnd.n2600 gnd.n1349 99.6594
R5841 gnd.n1133 gnd.n1051 99.6594
R5842 gnd.n2420 gnd.n1052 99.6594
R5843 gnd.n2426 gnd.n1053 99.6594
R5844 gnd.n2430 gnd.n1054 99.6594
R5845 gnd.n2436 gnd.n1055 99.6594
R5846 gnd.n2440 gnd.n1056 99.6594
R5847 gnd.n2446 gnd.n1057 99.6594
R5848 gnd.n2450 gnd.n1058 99.6594
R5849 gnd.n2409 gnd.n1059 99.6594
R5850 gnd.n2419 gnd.n1051 99.6594
R5851 gnd.n2425 gnd.n1052 99.6594
R5852 gnd.n2429 gnd.n1053 99.6594
R5853 gnd.n2435 gnd.n1054 99.6594
R5854 gnd.n2439 gnd.n1055 99.6594
R5855 gnd.n2445 gnd.n1056 99.6594
R5856 gnd.n2449 gnd.n1057 99.6594
R5857 gnd.n2408 gnd.n1058 99.6594
R5858 gnd.n2404 gnd.n1059 99.6594
R5859 gnd.n2197 gnd.n1349 99.6594
R5860 gnd.n2183 gnd.n1348 99.6594
R5861 gnd.n2181 gnd.n1347 99.6594
R5862 gnd.n2173 gnd.n1346 99.6594
R5863 gnd.n2163 gnd.n1345 99.6594
R5864 gnd.n2161 gnd.n1344 99.6594
R5865 gnd.n2153 gnd.n1343 99.6594
R5866 gnd.n2143 gnd.n1342 99.6594
R5867 gnd.n2141 gnd.n1341 99.6594
R5868 gnd.n4751 gnd.n4674 99.6594
R5869 gnd.n4743 gnd.n4662 99.6594
R5870 gnd.n4739 gnd.n4663 99.6594
R5871 gnd.n4735 gnd.n4664 99.6594
R5872 gnd.n4731 gnd.n4665 99.6594
R5873 gnd.n4727 gnd.n4666 99.6594
R5874 gnd.n4723 gnd.n4667 99.6594
R5875 gnd.n4719 gnd.n4668 99.6594
R5876 gnd.n4715 gnd.n4669 99.6594
R5877 gnd.n4711 gnd.n4670 99.6594
R5878 gnd.n4707 gnd.n4671 99.6594
R5879 gnd.n4703 gnd.n4672 99.6594
R5880 gnd.n4754 gnd.n4753 99.6594
R5881 gnd.n5518 gnd.n1022 99.6594
R5882 gnd.n5522 gnd.n1021 99.6594
R5883 gnd.n5526 gnd.n1020 99.6594
R5884 gnd.n5530 gnd.n1019 99.6594
R5885 gnd.n5534 gnd.n1018 99.6594
R5886 gnd.n5538 gnd.n1017 99.6594
R5887 gnd.n5542 gnd.n1016 99.6594
R5888 gnd.n5546 gnd.n1015 99.6594
R5889 gnd.n5550 gnd.n1014 99.6594
R5890 gnd.n5554 gnd.n1013 99.6594
R5891 gnd.n5558 gnd.n1012 99.6594
R5892 gnd.n5562 gnd.n1011 99.6594
R5893 gnd.n4186 gnd.n1010 99.6594
R5894 gnd.n399 gnd.n313 99.6594
R5895 gnd.n407 gnd.n314 99.6594
R5896 gnd.n409 gnd.n315 99.6594
R5897 gnd.n417 gnd.n316 99.6594
R5898 gnd.n425 gnd.n317 99.6594
R5899 gnd.n427 gnd.n318 99.6594
R5900 gnd.n435 gnd.n319 99.6594
R5901 gnd.n445 gnd.n320 99.6594
R5902 gnd.n6366 gnd.n321 99.6594
R5903 gnd.n6836 gnd.n6733 99.6594
R5904 gnd.n6782 gnd.n6732 99.6594
R5905 gnd.n6774 gnd.n6731 99.6594
R5906 gnd.n6772 gnd.n6730 99.6594
R5907 gnd.n6764 gnd.n6729 99.6594
R5908 gnd.n6762 gnd.n6728 99.6594
R5909 gnd.n6754 gnd.n6727 99.6594
R5910 gnd.n6752 gnd.n6726 99.6594
R5911 gnd.n6746 gnd.n6725 99.6594
R5912 gnd.n4837 gnd.n4836 99.6594
R5913 gnd.n4596 gnd.n4574 99.6594
R5914 gnd.n4602 gnd.n4575 99.6594
R5915 gnd.n4606 gnd.n4576 99.6594
R5916 gnd.n4612 gnd.n4577 99.6594
R5917 gnd.n4616 gnd.n4578 99.6594
R5918 gnd.n4622 gnd.n4579 99.6594
R5919 gnd.n4580 gnd.n4564 99.6594
R5920 gnd.n5572 gnd.n4158 99.6594
R5921 gnd.n5576 gnd.n4159 99.6594
R5922 gnd.n5580 gnd.n4160 99.6594
R5923 gnd.n5584 gnd.n4161 99.6594
R5924 gnd.n5588 gnd.n4162 99.6594
R5925 gnd.n5592 gnd.n4163 99.6594
R5926 gnd.n5596 gnd.n4164 99.6594
R5927 gnd.n4167 gnd.n4165 99.6594
R5928 gnd.n4156 gnd.n1063 99.6594
R5929 gnd.n4148 gnd.n1023 99.6594
R5930 gnd.n4144 gnd.n1024 99.6594
R5931 gnd.n4140 gnd.n1025 99.6594
R5932 gnd.n4136 gnd.n1026 99.6594
R5933 gnd.n4132 gnd.n1027 99.6594
R5934 gnd.n4128 gnd.n1028 99.6594
R5935 gnd.n4124 gnd.n1029 99.6594
R5936 gnd.n4119 gnd.n1030 99.6594
R5937 gnd.n4115 gnd.n1031 99.6594
R5938 gnd.n4111 gnd.n1032 99.6594
R5939 gnd.n4107 gnd.n1033 99.6594
R5940 gnd.n4103 gnd.n1034 99.6594
R5941 gnd.n4099 gnd.n1035 99.6594
R5942 gnd.n4095 gnd.n1036 99.6594
R5943 gnd.n4091 gnd.n1037 99.6594
R5944 gnd.n4087 gnd.n1038 99.6594
R5945 gnd.n4083 gnd.n1039 99.6594
R5946 gnd.n4079 gnd.n1040 99.6594
R5947 gnd.n4075 gnd.n1041 99.6594
R5948 gnd.n4071 gnd.n1042 99.6594
R5949 gnd.n4067 gnd.n1043 99.6594
R5950 gnd.n4063 gnd.n1044 99.6594
R5951 gnd.n4059 gnd.n1045 99.6594
R5952 gnd.n4055 gnd.n1046 99.6594
R5953 gnd.n4051 gnd.n1047 99.6594
R5954 gnd.n4047 gnd.n1048 99.6594
R5955 gnd.n4043 gnd.n1049 99.6594
R5956 gnd.n1135 gnd.n1050 99.6594
R5957 gnd.n2288 gnd.n1351 99.6594
R5958 gnd.n2286 gnd.n1352 99.6594
R5959 gnd.n2278 gnd.n1353 99.6594
R5960 gnd.n2276 gnd.n1354 99.6594
R5961 gnd.n2268 gnd.n1355 99.6594
R5962 gnd.n2266 gnd.n1356 99.6594
R5963 gnd.n2258 gnd.n1357 99.6594
R5964 gnd.n2256 gnd.n1358 99.6594
R5965 gnd.n2248 gnd.n1359 99.6594
R5966 gnd.n2246 gnd.n1360 99.6594
R5967 gnd.n2238 gnd.n1361 99.6594
R5968 gnd.n2236 gnd.n1362 99.6594
R5969 gnd.n2228 gnd.n1363 99.6594
R5970 gnd.n2226 gnd.n1364 99.6594
R5971 gnd.n2219 gnd.n1365 99.6594
R5972 gnd.n3855 gnd.n1367 99.6594
R5973 gnd.n3859 gnd.n1368 99.6594
R5974 gnd.n3863 gnd.n1369 99.6594
R5975 gnd.n3867 gnd.n1370 99.6594
R5976 gnd.n3872 gnd.n1371 99.6594
R5977 gnd.n3876 gnd.n1372 99.6594
R5978 gnd.n3880 gnd.n1373 99.6594
R5979 gnd.n3884 gnd.n1374 99.6594
R5980 gnd.n3888 gnd.n1375 99.6594
R5981 gnd.n3892 gnd.n1376 99.6594
R5982 gnd.n3896 gnd.n1377 99.6594
R5983 gnd.n1379 gnd.n1378 99.6594
R5984 gnd.n3902 gnd.n1338 99.6594
R5985 gnd.n6531 gnd.n283 99.6594
R5986 gnd.n6525 gnd.n285 99.6594
R5987 gnd.n6521 gnd.n286 99.6594
R5988 gnd.n6517 gnd.n287 99.6594
R5989 gnd.n6513 gnd.n288 99.6594
R5990 gnd.n6509 gnd.n289 99.6594
R5991 gnd.n6505 gnd.n290 99.6594
R5992 gnd.n6501 gnd.n291 99.6594
R5993 gnd.n6496 gnd.n292 99.6594
R5994 gnd.n6492 gnd.n293 99.6594
R5995 gnd.n6488 gnd.n294 99.6594
R5996 gnd.n6484 gnd.n295 99.6594
R5997 gnd.n6479 gnd.n297 99.6594
R5998 gnd.n6475 gnd.n298 99.6594
R5999 gnd.n6471 gnd.n299 99.6594
R6000 gnd.n6467 gnd.n300 99.6594
R6001 gnd.n6463 gnd.n301 99.6594
R6002 gnd.n6459 gnd.n302 99.6594
R6003 gnd.n6455 gnd.n303 99.6594
R6004 gnd.n6451 gnd.n304 99.6594
R6005 gnd.n6447 gnd.n305 99.6594
R6006 gnd.n6443 gnd.n306 99.6594
R6007 gnd.n6439 gnd.n307 99.6594
R6008 gnd.n6435 gnd.n308 99.6594
R6009 gnd.n6431 gnd.n309 99.6594
R6010 gnd.n6427 gnd.n310 99.6594
R6011 gnd.n6423 gnd.n311 99.6594
R6012 gnd.n500 gnd.n312 99.6594
R6013 gnd.n7043 gnd.n6723 99.6594
R6014 gnd.n6925 gnd.n6837 99.6594
R6015 gnd.n6929 gnd.n6838 99.6594
R6016 gnd.n6933 gnd.n6839 99.6594
R6017 gnd.n6937 gnd.n6840 99.6594
R6018 gnd.n6941 gnd.n6841 99.6594
R6019 gnd.n6945 gnd.n6842 99.6594
R6020 gnd.n6949 gnd.n6843 99.6594
R6021 gnd.n6953 gnd.n6844 99.6594
R6022 gnd.n6957 gnd.n6845 99.6594
R6023 gnd.n6963 gnd.n6846 99.6594
R6024 gnd.n6967 gnd.n6847 99.6594
R6025 gnd.n6971 gnd.n6848 99.6594
R6026 gnd.n6975 gnd.n6849 99.6594
R6027 gnd.n6979 gnd.n6850 99.6594
R6028 gnd.n6983 gnd.n6851 99.6594
R6029 gnd.n6987 gnd.n6852 99.6594
R6030 gnd.n6991 gnd.n6853 99.6594
R6031 gnd.n6995 gnd.n6854 99.6594
R6032 gnd.n6999 gnd.n6855 99.6594
R6033 gnd.n7006 gnd.n6856 99.6594
R6034 gnd.n7010 gnd.n6857 99.6594
R6035 gnd.n7014 gnd.n6858 99.6594
R6036 gnd.n7018 gnd.n6859 99.6594
R6037 gnd.n7022 gnd.n6860 99.6594
R6038 gnd.n7026 gnd.n6861 99.6594
R6039 gnd.n7030 gnd.n6862 99.6594
R6040 gnd.n7034 gnd.n6863 99.6594
R6041 gnd.n6865 gnd.n6864 99.6594
R6042 gnd.n2662 gnd.n2661 99.6594
R6043 gnd.n2126 gnd.n2112 99.6594
R6044 gnd.n2130 gnd.n2113 99.6594
R6045 gnd.n2132 gnd.n2114 99.6594
R6046 gnd.n2137 gnd.n2115 99.6594
R6047 gnd.n2147 gnd.n2116 99.6594
R6048 gnd.n2149 gnd.n2117 99.6594
R6049 gnd.n2157 gnd.n2118 99.6594
R6050 gnd.n2167 gnd.n2119 99.6594
R6051 gnd.n2169 gnd.n2120 99.6594
R6052 gnd.n2177 gnd.n2121 99.6594
R6053 gnd.n2187 gnd.n2122 99.6594
R6054 gnd.n2549 gnd.n2123 99.6594
R6055 gnd.n2554 gnd.n2124 99.6594
R6056 gnd.n2661 gnd.n2110 99.6594
R6057 gnd.n2129 gnd.n2112 99.6594
R6058 gnd.n2131 gnd.n2113 99.6594
R6059 gnd.n2136 gnd.n2114 99.6594
R6060 gnd.n2146 gnd.n2115 99.6594
R6061 gnd.n2148 gnd.n2116 99.6594
R6062 gnd.n2156 gnd.n2117 99.6594
R6063 gnd.n2166 gnd.n2118 99.6594
R6064 gnd.n2168 gnd.n2119 99.6594
R6065 gnd.n2176 gnd.n2120 99.6594
R6066 gnd.n2186 gnd.n2121 99.6594
R6067 gnd.n2188 gnd.n2122 99.6594
R6068 gnd.n2553 gnd.n2123 99.6594
R6069 gnd.n2555 gnd.n2124 99.6594
R6070 gnd.n471 gnd.n464 99.6594
R6071 gnd.n473 gnd.n472 99.6594
R6072 gnd.n6342 gnd.n469 99.6594
R6073 gnd.n6340 gnd.n392 99.6594
R6074 gnd.n474 gnd.n394 99.6594
R6075 gnd.n476 gnd.n403 99.6594
R6076 gnd.n478 gnd.n477 99.6594
R6077 gnd.n479 gnd.n414 99.6594
R6078 gnd.n481 gnd.n421 99.6594
R6079 gnd.n483 gnd.n482 99.6594
R6080 gnd.n484 gnd.n432 99.6594
R6081 gnd.n486 gnd.n439 99.6594
R6082 gnd.n488 gnd.n487 99.6594
R6083 gnd.n489 gnd.n451 99.6594
R6084 gnd.n486 gnd.n485 99.6594
R6085 gnd.n484 gnd.n431 99.6594
R6086 gnd.n483 gnd.n422 99.6594
R6087 gnd.n481 gnd.n480 99.6594
R6088 gnd.n479 gnd.n413 99.6594
R6089 gnd.n478 gnd.n404 99.6594
R6090 gnd.n476 gnd.n475 99.6594
R6091 gnd.n474 gnd.n393 99.6594
R6092 gnd.n6341 gnd.n6340 99.6594
R6093 gnd.n469 gnd.n468 99.6594
R6094 gnd.n473 gnd.n465 99.6594
R6095 gnd.n471 gnd.n460 99.6594
R6096 gnd.n489 gnd.n456 99.6594
R6097 gnd.n488 gnd.n450 99.6594
R6098 gnd.n2189 gnd.t251 98.63
R6099 gnd.n6367 gnd.t217 98.63
R6100 gnd.n6720 gnd.t256 98.63
R6101 gnd.n6903 gnd.t269 98.63
R6102 gnd.n7002 gnd.t278 98.63
R6103 gnd.n341 gnd.t294 98.63
R6104 gnd.n364 gnd.t297 98.63
R6105 gnd.n386 gnd.t260 98.63
R6106 gnd.n6735 gnd.t206 98.63
R6107 gnd.n2194 gnd.t232 98.63
R6108 gnd.n2405 gnd.t229 98.63
R6109 gnd.n1083 gnd.t254 98.63
R6110 gnd.n1105 gnd.t276 98.63
R6111 gnd.n1127 gnd.t285 98.63
R6112 gnd.n1396 gnd.t272 98.63
R6113 gnd.n2200 gnd.t287 98.63
R6114 gnd.n2212 gnd.t306 98.63
R6115 gnd.n441 gnd.t224 98.63
R6116 gnd.n2809 gnd.t318 88.9408
R6117 gnd.n1698 gnd.t309 88.9408
R6118 gnd.n3784 gnd.t241 88.933
R6119 gnd.n1692 gnd.t236 88.933
R6120 gnd.n6102 gnd.n643 87.1465
R6121 gnd.n6103 gnd.n6102 87.1465
R6122 gnd.n6104 gnd.n6103 87.1465
R6123 gnd.n6104 gnd.n637 87.1465
R6124 gnd.n6112 gnd.n637 87.1465
R6125 gnd.n6113 gnd.n6112 87.1465
R6126 gnd.n6114 gnd.n6113 87.1465
R6127 gnd.n6114 gnd.n631 87.1465
R6128 gnd.n6122 gnd.n631 87.1465
R6129 gnd.n6123 gnd.n6122 87.1465
R6130 gnd.n6124 gnd.n6123 87.1465
R6131 gnd.n6124 gnd.n625 87.1465
R6132 gnd.n6132 gnd.n625 87.1465
R6133 gnd.n6133 gnd.n6132 87.1465
R6134 gnd.n6134 gnd.n6133 87.1465
R6135 gnd.n6134 gnd.n619 87.1465
R6136 gnd.n6142 gnd.n619 87.1465
R6137 gnd.n6143 gnd.n6142 87.1465
R6138 gnd.n6144 gnd.n6143 87.1465
R6139 gnd.n6144 gnd.n613 87.1465
R6140 gnd.n6152 gnd.n613 87.1465
R6141 gnd.n6153 gnd.n6152 87.1465
R6142 gnd.n6154 gnd.n6153 87.1465
R6143 gnd.n6154 gnd.n607 87.1465
R6144 gnd.n6162 gnd.n607 87.1465
R6145 gnd.n6163 gnd.n6162 87.1465
R6146 gnd.n6164 gnd.n6163 87.1465
R6147 gnd.n6164 gnd.n601 87.1465
R6148 gnd.n6172 gnd.n601 87.1465
R6149 gnd.n6173 gnd.n6172 87.1465
R6150 gnd.n6174 gnd.n6173 87.1465
R6151 gnd.n6174 gnd.n595 87.1465
R6152 gnd.n6182 gnd.n595 87.1465
R6153 gnd.n6183 gnd.n6182 87.1465
R6154 gnd.n6184 gnd.n6183 87.1465
R6155 gnd.n6184 gnd.n589 87.1465
R6156 gnd.n6192 gnd.n589 87.1465
R6157 gnd.n6193 gnd.n6192 87.1465
R6158 gnd.n6194 gnd.n6193 87.1465
R6159 gnd.n6194 gnd.n583 87.1465
R6160 gnd.n6202 gnd.n583 87.1465
R6161 gnd.n6203 gnd.n6202 87.1465
R6162 gnd.n6204 gnd.n6203 87.1465
R6163 gnd.n6204 gnd.n577 87.1465
R6164 gnd.n6212 gnd.n577 87.1465
R6165 gnd.n6213 gnd.n6212 87.1465
R6166 gnd.n6214 gnd.n6213 87.1465
R6167 gnd.n6214 gnd.n571 87.1465
R6168 gnd.n6222 gnd.n571 87.1465
R6169 gnd.n6223 gnd.n6222 87.1465
R6170 gnd.n6224 gnd.n6223 87.1465
R6171 gnd.n6224 gnd.n565 87.1465
R6172 gnd.n6232 gnd.n565 87.1465
R6173 gnd.n6233 gnd.n6232 87.1465
R6174 gnd.n6234 gnd.n6233 87.1465
R6175 gnd.n6234 gnd.n559 87.1465
R6176 gnd.n6242 gnd.n559 87.1465
R6177 gnd.n6243 gnd.n6242 87.1465
R6178 gnd.n6244 gnd.n6243 87.1465
R6179 gnd.n6244 gnd.n553 87.1465
R6180 gnd.n6252 gnd.n553 87.1465
R6181 gnd.n6253 gnd.n6252 87.1465
R6182 gnd.n6254 gnd.n6253 87.1465
R6183 gnd.n6254 gnd.n547 87.1465
R6184 gnd.n6262 gnd.n547 87.1465
R6185 gnd.n6263 gnd.n6262 87.1465
R6186 gnd.n6264 gnd.n6263 87.1465
R6187 gnd.n6264 gnd.n541 87.1465
R6188 gnd.n6272 gnd.n541 87.1465
R6189 gnd.n6273 gnd.n6272 87.1465
R6190 gnd.n6274 gnd.n6273 87.1465
R6191 gnd.n6274 gnd.n535 87.1465
R6192 gnd.n6282 gnd.n535 87.1465
R6193 gnd.n6283 gnd.n6282 87.1465
R6194 gnd.n6284 gnd.n6283 87.1465
R6195 gnd.n6284 gnd.n529 87.1465
R6196 gnd.n6292 gnd.n529 87.1465
R6197 gnd.n6293 gnd.n6292 87.1465
R6198 gnd.n6294 gnd.n6293 87.1465
R6199 gnd.n6294 gnd.n523 87.1465
R6200 gnd.n6304 gnd.n523 87.1465
R6201 gnd.n6305 gnd.n6304 87.1465
R6202 gnd.n6307 gnd.n6305 87.1465
R6203 gnd.n1458 gnd.n1457 81.8399
R6204 gnd.n4625 gnd.t263 74.8376
R6205 gnd.n4183 gnd.t322 74.8376
R6206 gnd.n2810 gnd.t317 72.8438
R6207 gnd.n1699 gnd.t310 72.8438
R6208 gnd.n1459 gnd.n1452 72.8411
R6209 gnd.n1465 gnd.n1450 72.8411
R6210 gnd.n1665 gnd.n1664 72.8411
R6211 gnd.n2190 gnd.t250 72.836
R6212 gnd.n3785 gnd.t240 72.836
R6213 gnd.n1693 gnd.t237 72.836
R6214 gnd.n6368 gnd.t216 72.836
R6215 gnd.n6721 gnd.t257 72.836
R6216 gnd.n6904 gnd.t270 72.836
R6217 gnd.n7003 gnd.t279 72.836
R6218 gnd.n342 gnd.t293 72.836
R6219 gnd.n365 gnd.t296 72.836
R6220 gnd.n387 gnd.t259 72.836
R6221 gnd.n6736 gnd.t207 72.836
R6222 gnd.n2195 gnd.t233 72.836
R6223 gnd.n2406 gnd.t228 72.836
R6224 gnd.n1084 gnd.t253 72.836
R6225 gnd.n1106 gnd.t275 72.836
R6226 gnd.n1128 gnd.t284 72.836
R6227 gnd.n1397 gnd.t273 72.836
R6228 gnd.n2201 gnd.t288 72.836
R6229 gnd.n2213 gnd.t307 72.836
R6230 gnd.n442 gnd.t225 72.836
R6231 gnd.n3537 gnd.n1670 71.676
R6232 gnd.n3535 gnd.n3534 71.676
R6233 gnd.n3530 gnd.n1675 71.676
R6234 gnd.n3528 gnd.n3527 71.676
R6235 gnd.n3523 gnd.n1678 71.676
R6236 gnd.n3521 gnd.n3520 71.676
R6237 gnd.n3516 gnd.n1681 71.676
R6238 gnd.n3514 gnd.n3513 71.676
R6239 gnd.n3509 gnd.n1684 71.676
R6240 gnd.n3507 gnd.n3506 71.676
R6241 gnd.n3502 gnd.n1687 71.676
R6242 gnd.n3500 gnd.n3499 71.676
R6243 gnd.n3495 gnd.n1690 71.676
R6244 gnd.n3493 gnd.n3492 71.676
R6245 gnd.n3487 gnd.n1695 71.676
R6246 gnd.n3485 gnd.n3484 71.676
R6247 gnd.n3480 gnd.n3479 71.676
R6248 gnd.n3477 gnd.n3476 71.676
R6249 gnd.n3471 gnd.n1701 71.676
R6250 gnd.n3469 gnd.n3468 71.676
R6251 gnd.n3464 gnd.n1704 71.676
R6252 gnd.n3462 gnd.n3461 71.676
R6253 gnd.n3457 gnd.n1707 71.676
R6254 gnd.n3455 gnd.n3454 71.676
R6255 gnd.n3450 gnd.n1710 71.676
R6256 gnd.n3448 gnd.n3447 71.676
R6257 gnd.n3443 gnd.n1713 71.676
R6258 gnd.n3441 gnd.n3440 71.676
R6259 gnd.n3436 gnd.n1716 71.676
R6260 gnd.n3434 gnd.n3433 71.676
R6261 gnd.n3429 gnd.n1719 71.676
R6262 gnd.n3427 gnd.n3426 71.676
R6263 gnd.n3422 gnd.n3421 71.676
R6264 gnd.n3848 gnd.n3847 71.676
R6265 gnd.n3842 gnd.n1414 71.676
R6266 gnd.n3839 gnd.n1415 71.676
R6267 gnd.n3835 gnd.n1416 71.676
R6268 gnd.n3831 gnd.n1417 71.676
R6269 gnd.n3827 gnd.n1418 71.676
R6270 gnd.n3823 gnd.n1419 71.676
R6271 gnd.n3819 gnd.n1420 71.676
R6272 gnd.n3815 gnd.n1421 71.676
R6273 gnd.n3811 gnd.n1422 71.676
R6274 gnd.n3807 gnd.n1423 71.676
R6275 gnd.n3803 gnd.n1424 71.676
R6276 gnd.n3799 gnd.n1425 71.676
R6277 gnd.n3795 gnd.n1426 71.676
R6278 gnd.n3791 gnd.n1427 71.676
R6279 gnd.n3787 gnd.n1428 71.676
R6280 gnd.n1429 gnd.n1412 71.676
R6281 gnd.n2813 gnd.n1430 71.676
R6282 gnd.n2818 gnd.n1431 71.676
R6283 gnd.n2822 gnd.n1432 71.676
R6284 gnd.n2826 gnd.n1433 71.676
R6285 gnd.n2830 gnd.n1434 71.676
R6286 gnd.n2834 gnd.n1435 71.676
R6287 gnd.n2838 gnd.n1436 71.676
R6288 gnd.n2842 gnd.n1437 71.676
R6289 gnd.n2846 gnd.n1438 71.676
R6290 gnd.n2850 gnd.n1439 71.676
R6291 gnd.n2854 gnd.n1440 71.676
R6292 gnd.n2858 gnd.n1441 71.676
R6293 gnd.n2862 gnd.n1442 71.676
R6294 gnd.n2866 gnd.n1443 71.676
R6295 gnd.n2870 gnd.n1444 71.676
R6296 gnd.n3848 gnd.n1447 71.676
R6297 gnd.n3840 gnd.n1414 71.676
R6298 gnd.n3836 gnd.n1415 71.676
R6299 gnd.n3832 gnd.n1416 71.676
R6300 gnd.n3828 gnd.n1417 71.676
R6301 gnd.n3824 gnd.n1418 71.676
R6302 gnd.n3820 gnd.n1419 71.676
R6303 gnd.n3816 gnd.n1420 71.676
R6304 gnd.n3812 gnd.n1421 71.676
R6305 gnd.n3808 gnd.n1422 71.676
R6306 gnd.n3804 gnd.n1423 71.676
R6307 gnd.n3800 gnd.n1424 71.676
R6308 gnd.n3796 gnd.n1425 71.676
R6309 gnd.n3792 gnd.n1426 71.676
R6310 gnd.n3788 gnd.n1427 71.676
R6311 gnd.n3851 gnd.n3850 71.676
R6312 gnd.n2812 gnd.n1429 71.676
R6313 gnd.n2817 gnd.n1430 71.676
R6314 gnd.n2821 gnd.n1431 71.676
R6315 gnd.n2825 gnd.n1432 71.676
R6316 gnd.n2829 gnd.n1433 71.676
R6317 gnd.n2833 gnd.n1434 71.676
R6318 gnd.n2837 gnd.n1435 71.676
R6319 gnd.n2841 gnd.n1436 71.676
R6320 gnd.n2845 gnd.n1437 71.676
R6321 gnd.n2849 gnd.n1438 71.676
R6322 gnd.n2853 gnd.n1439 71.676
R6323 gnd.n2857 gnd.n1440 71.676
R6324 gnd.n2861 gnd.n1441 71.676
R6325 gnd.n2865 gnd.n1442 71.676
R6326 gnd.n2869 gnd.n1443 71.676
R6327 gnd.n2808 gnd.n1444 71.676
R6328 gnd.n3421 gnd.n1720 71.676
R6329 gnd.n3428 gnd.n3427 71.676
R6330 gnd.n1719 gnd.n1717 71.676
R6331 gnd.n3435 gnd.n3434 71.676
R6332 gnd.n1716 gnd.n1714 71.676
R6333 gnd.n3442 gnd.n3441 71.676
R6334 gnd.n1713 gnd.n1711 71.676
R6335 gnd.n3449 gnd.n3448 71.676
R6336 gnd.n1710 gnd.n1708 71.676
R6337 gnd.n3456 gnd.n3455 71.676
R6338 gnd.n1707 gnd.n1705 71.676
R6339 gnd.n3463 gnd.n3462 71.676
R6340 gnd.n1704 gnd.n1702 71.676
R6341 gnd.n3470 gnd.n3469 71.676
R6342 gnd.n1701 gnd.n1697 71.676
R6343 gnd.n3478 gnd.n3477 71.676
R6344 gnd.n3482 gnd.n3481 71.676
R6345 gnd.n3486 gnd.n3485 71.676
R6346 gnd.n1695 gnd.n1691 71.676
R6347 gnd.n3494 gnd.n3493 71.676
R6348 gnd.n1690 gnd.n1688 71.676
R6349 gnd.n3501 gnd.n3500 71.676
R6350 gnd.n1687 gnd.n1685 71.676
R6351 gnd.n3508 gnd.n3507 71.676
R6352 gnd.n1684 gnd.n1682 71.676
R6353 gnd.n3515 gnd.n3514 71.676
R6354 gnd.n1681 gnd.n1679 71.676
R6355 gnd.n3522 gnd.n3521 71.676
R6356 gnd.n1678 gnd.n1676 71.676
R6357 gnd.n3529 gnd.n3528 71.676
R6358 gnd.n1675 gnd.n1673 71.676
R6359 gnd.n3536 gnd.n3535 71.676
R6360 gnd.n1670 gnd.n1648 71.676
R6361 gnd.n10 gnd.t201 69.1507
R6362 gnd.n18 gnd.t60 68.4792
R6363 gnd.n17 gnd.t156 68.4792
R6364 gnd.n16 gnd.t193 68.4792
R6365 gnd.n15 gnd.t130 68.4792
R6366 gnd.n14 gnd.t115 68.4792
R6367 gnd.n13 gnd.t127 68.4792
R6368 gnd.n12 gnd.t123 68.4792
R6369 gnd.n11 gnd.t186 68.4792
R6370 gnd.n10 gnd.t196 68.4792
R6371 gnd.n4752 gnd.n4656 64.369
R6372 gnd.n4157 gnd.n1061 63.0944
R6373 gnd.n7042 gnd.n164 63.0944
R6374 gnd.n2815 gnd.n2810 59.5399
R6375 gnd.n3473 gnd.n1699 59.5399
R6376 gnd.n3786 gnd.n3785 59.5399
R6377 gnd.n3489 gnd.n1693 59.5399
R6378 gnd.n3783 gnd.n1468 59.1804
R6379 gnd.n4411 gnd.t334 56.407
R6380 gnd.n4376 gnd.t29 56.407
R6381 gnd.n4387 gnd.t110 56.407
R6382 gnd.n4399 gnd.t91 56.407
R6383 gnd.n56 gnd.t162 56.407
R6384 gnd.n21 gnd.t73 56.407
R6385 gnd.n32 gnd.t51 56.407
R6386 gnd.n44 gnd.t116 56.407
R6387 gnd.n4420 gnd.t133 55.8337
R6388 gnd.n4385 gnd.t41 55.8337
R6389 gnd.n4396 gnd.t113 55.8337
R6390 gnd.n4408 gnd.t184 55.8337
R6391 gnd.n65 gnd.t128 55.8337
R6392 gnd.n30 gnd.t173 55.8337
R6393 gnd.n41 gnd.t326 55.8337
R6394 gnd.n53 gnd.t100 55.8337
R6395 gnd.n1456 gnd.n1455 54.358
R6396 gnd.n1662 gnd.n1661 54.358
R6397 gnd.n4411 gnd.n4410 53.0052
R6398 gnd.n4413 gnd.n4412 53.0052
R6399 gnd.n4415 gnd.n4414 53.0052
R6400 gnd.n4417 gnd.n4416 53.0052
R6401 gnd.n4419 gnd.n4418 53.0052
R6402 gnd.n4376 gnd.n4375 53.0052
R6403 gnd.n4378 gnd.n4377 53.0052
R6404 gnd.n4380 gnd.n4379 53.0052
R6405 gnd.n4382 gnd.n4381 53.0052
R6406 gnd.n4384 gnd.n4383 53.0052
R6407 gnd.n4387 gnd.n4386 53.0052
R6408 gnd.n4389 gnd.n4388 53.0052
R6409 gnd.n4391 gnd.n4390 53.0052
R6410 gnd.n4393 gnd.n4392 53.0052
R6411 gnd.n4395 gnd.n4394 53.0052
R6412 gnd.n4399 gnd.n4398 53.0052
R6413 gnd.n4401 gnd.n4400 53.0052
R6414 gnd.n4403 gnd.n4402 53.0052
R6415 gnd.n4405 gnd.n4404 53.0052
R6416 gnd.n4407 gnd.n4406 53.0052
R6417 gnd.n64 gnd.n63 53.0052
R6418 gnd.n62 gnd.n61 53.0052
R6419 gnd.n60 gnd.n59 53.0052
R6420 gnd.n58 gnd.n57 53.0052
R6421 gnd.n56 gnd.n55 53.0052
R6422 gnd.n29 gnd.n28 53.0052
R6423 gnd.n27 gnd.n26 53.0052
R6424 gnd.n25 gnd.n24 53.0052
R6425 gnd.n23 gnd.n22 53.0052
R6426 gnd.n21 gnd.n20 53.0052
R6427 gnd.n40 gnd.n39 53.0052
R6428 gnd.n38 gnd.n37 53.0052
R6429 gnd.n36 gnd.n35 53.0052
R6430 gnd.n34 gnd.n33 53.0052
R6431 gnd.n32 gnd.n31 53.0052
R6432 gnd.n52 gnd.n51 53.0052
R6433 gnd.n50 gnd.n49 53.0052
R6434 gnd.n48 gnd.n47 53.0052
R6435 gnd.n46 gnd.n45 53.0052
R6436 gnd.n44 gnd.n43 53.0052
R6437 gnd.n1653 gnd.n1652 52.4801
R6438 gnd.n5456 gnd.t93 52.3082
R6439 gnd.n5424 gnd.t3 52.3082
R6440 gnd.n5392 gnd.t138 52.3082
R6441 gnd.n5361 gnd.t158 52.3082
R6442 gnd.n5329 gnd.t39 52.3082
R6443 gnd.n5297 gnd.t152 52.3082
R6444 gnd.n5265 gnd.t85 52.3082
R6445 gnd.n5234 gnd.t140 52.3082
R6446 gnd.n6307 gnd.n6306 52.2881
R6447 gnd.n5605 gnd.n5604 51.9414
R6448 gnd.n5286 gnd.n5254 51.4173
R6449 gnd.n5350 gnd.n5349 50.455
R6450 gnd.n5318 gnd.n5317 50.455
R6451 gnd.n5286 gnd.n5285 50.455
R6452 gnd.n4699 gnd.n4698 45.1884
R6453 gnd.n4209 gnd.n4208 45.1884
R6454 gnd.n3540 gnd.n1668 44.3322
R6455 gnd.n1459 gnd.n1458 44.3189
R6456 gnd.n2191 gnd.n2190 42.4732
R6457 gnd.n443 gnd.n442 42.4732
R6458 gnd.n6369 gnd.n6368 42.2793
R6459 gnd.n6722 gnd.n6721 42.2793
R6460 gnd.n6962 gnd.n6904 42.2793
R6461 gnd.n7004 gnd.n7003 42.2793
R6462 gnd.n6498 gnd.n342 42.2793
R6463 gnd.n6461 gnd.n365 42.2793
R6464 gnd.n6421 gnd.n387 42.2793
R6465 gnd.n6737 gnd.n6736 42.2793
R6466 gnd.n4700 gnd.n4699 42.2793
R6467 gnd.n4210 gnd.n4209 42.2793
R6468 gnd.n4626 gnd.n4625 42.2793
R6469 gnd.n5571 gnd.n4183 42.2793
R6470 gnd.n2602 gnd.n2195 42.2793
R6471 gnd.n2456 gnd.n2406 42.2793
R6472 gnd.n4121 gnd.n1084 42.2793
R6473 gnd.n4081 gnd.n1106 42.2793
R6474 gnd.n4041 gnd.n1128 42.2793
R6475 gnd.n3870 gnd.n1397 42.2793
R6476 gnd.n2202 gnd.n2201 42.2793
R6477 gnd.n2214 gnd.n2213 42.2793
R6478 gnd.n1457 gnd.n1456 41.6274
R6479 gnd.n1663 gnd.n1662 41.6274
R6480 gnd.n1466 gnd.n1465 40.8975
R6481 gnd.n1666 gnd.n1665 40.8975
R6482 gnd.n1465 gnd.n1464 35.055
R6483 gnd.n1460 gnd.n1459 35.055
R6484 gnd.n1655 gnd.n1654 35.055
R6485 gnd.n1665 gnd.n1651 35.055
R6486 gnd.n5773 gnd.n5772 32.3154
R6487 gnd.n5772 gnd.n840 32.3154
R6488 gnd.n5766 gnd.n840 32.3154
R6489 gnd.n5766 gnd.n5765 32.3154
R6490 gnd.n5765 gnd.n5764 32.3154
R6491 gnd.n5764 gnd.n848 32.3154
R6492 gnd.n5758 gnd.n848 32.3154
R6493 gnd.n5758 gnd.n5757 32.3154
R6494 gnd.n5757 gnd.n5756 32.3154
R6495 gnd.n5756 gnd.n856 32.3154
R6496 gnd.n5750 gnd.n856 32.3154
R6497 gnd.n5750 gnd.n5749 32.3154
R6498 gnd.n5749 gnd.n5748 32.3154
R6499 gnd.n5748 gnd.n864 32.3154
R6500 gnd.n5742 gnd.n864 32.3154
R6501 gnd.n5742 gnd.n5741 32.3154
R6502 gnd.n5741 gnd.n5740 32.3154
R6503 gnd.n5740 gnd.n872 32.3154
R6504 gnd.n5734 gnd.n872 32.3154
R6505 gnd.n5734 gnd.n5733 32.3154
R6506 gnd.n5733 gnd.n5732 32.3154
R6507 gnd.n5732 gnd.n880 32.3154
R6508 gnd.n5726 gnd.n880 32.3154
R6509 gnd.n5726 gnd.n5725 32.3154
R6510 gnd.n5725 gnd.n5724 32.3154
R6511 gnd.n5724 gnd.n888 32.3154
R6512 gnd.n5718 gnd.n888 32.3154
R6513 gnd.n5718 gnd.n5717 32.3154
R6514 gnd.n5717 gnd.n5716 32.3154
R6515 gnd.n5716 gnd.n896 32.3154
R6516 gnd.n5710 gnd.n896 32.3154
R6517 gnd.n5710 gnd.n5709 32.3154
R6518 gnd.n5709 gnd.n5708 32.3154
R6519 gnd.n5708 gnd.n904 32.3154
R6520 gnd.n5702 gnd.n904 32.3154
R6521 gnd.n5702 gnd.n5701 32.3154
R6522 gnd.n5701 gnd.n5700 32.3154
R6523 gnd.n5700 gnd.n912 32.3154
R6524 gnd.n5694 gnd.n912 32.3154
R6525 gnd.n5694 gnd.n5693 32.3154
R6526 gnd.n5693 gnd.n5692 32.3154
R6527 gnd.n5692 gnd.n920 32.3154
R6528 gnd.n5686 gnd.n920 32.3154
R6529 gnd.n5686 gnd.n5685 32.3154
R6530 gnd.n5685 gnd.n5684 32.3154
R6531 gnd.n5684 gnd.n928 32.3154
R6532 gnd.n5678 gnd.n928 32.3154
R6533 gnd.n5678 gnd.n5677 32.3154
R6534 gnd.n5677 gnd.n5676 32.3154
R6535 gnd.n5676 gnd.n936 32.3154
R6536 gnd.n5670 gnd.n936 32.3154
R6537 gnd.n5670 gnd.n5669 32.3154
R6538 gnd.n5669 gnd.n5668 32.3154
R6539 gnd.n5668 gnd.n944 32.3154
R6540 gnd.n5662 gnd.n944 32.3154
R6541 gnd.n5662 gnd.n5661 32.3154
R6542 gnd.n5661 gnd.n5660 32.3154
R6543 gnd.n5660 gnd.n952 32.3154
R6544 gnd.n5654 gnd.n952 32.3154
R6545 gnd.n5654 gnd.n5653 32.3154
R6546 gnd.n5653 gnd.n5652 32.3154
R6547 gnd.n5652 gnd.n960 32.3154
R6548 gnd.n5646 gnd.n960 32.3154
R6549 gnd.n5646 gnd.n5645 32.3154
R6550 gnd.n5645 gnd.n5644 32.3154
R6551 gnd.n5644 gnd.n968 32.3154
R6552 gnd.n5638 gnd.n968 32.3154
R6553 gnd.n5638 gnd.n5637 32.3154
R6554 gnd.n5637 gnd.n5636 32.3154
R6555 gnd.n5636 gnd.n976 32.3154
R6556 gnd.n5630 gnd.n976 32.3154
R6557 gnd.n5630 gnd.n5629 32.3154
R6558 gnd.n5629 gnd.n5628 32.3154
R6559 gnd.n5628 gnd.n984 32.3154
R6560 gnd.n5622 gnd.n984 32.3154
R6561 gnd.n5622 gnd.n5621 32.3154
R6562 gnd.n5621 gnd.n5620 32.3154
R6563 gnd.n5620 gnd.n992 32.3154
R6564 gnd.n5614 gnd.n992 32.3154
R6565 gnd.n5614 gnd.n5613 32.3154
R6566 gnd.n5613 gnd.n5612 32.3154
R6567 gnd.n5612 gnd.n1000 32.3154
R6568 gnd.n5606 gnd.n1000 32.3154
R6569 gnd.n4762 gnd.n4656 31.8661
R6570 gnd.n4762 gnd.n4761 31.8661
R6571 gnd.n4770 gnd.n4645 31.8661
R6572 gnd.n4778 gnd.n4645 31.8661
R6573 gnd.n4778 gnd.n4639 31.8661
R6574 gnd.n4786 gnd.n4639 31.8661
R6575 gnd.n4786 gnd.n4632 31.8661
R6576 gnd.n4824 gnd.n4632 31.8661
R6577 gnd.n4834 gnd.n4565 31.8661
R6578 gnd.n4033 gnd.n1061 31.8661
R6579 gnd.n4025 gnd.n1146 31.8661
R6580 gnd.n4025 gnd.n1149 31.8661
R6581 gnd.n4019 gnd.n1149 31.8661
R6582 gnd.n4019 gnd.n1159 31.8661
R6583 gnd.n4013 gnd.n1168 31.8661
R6584 gnd.n4007 gnd.n1168 31.8661
R6585 gnd.n4001 gnd.n1184 31.8661
R6586 gnd.n3995 gnd.n1193 31.8661
R6587 gnd.n3995 gnd.n1196 31.8661
R6588 gnd.n3989 gnd.n1206 31.8661
R6589 gnd.n3983 gnd.n1206 31.8661
R6590 gnd.n3977 gnd.n1222 31.8661
R6591 gnd.n3971 gnd.n1231 31.8661
R6592 gnd.n3971 gnd.n1234 31.8661
R6593 gnd.n3965 gnd.n1244 31.8661
R6594 gnd.n3959 gnd.n1253 31.8661
R6595 gnd.n3953 gnd.n1253 31.8661
R6596 gnd.n3947 gnd.n1269 31.8661
R6597 gnd.n3947 gnd.n1272 31.8661
R6598 gnd.n3941 gnd.n1282 31.8661
R6599 gnd.n3929 gnd.n1299 31.8661
R6600 gnd.n2597 gnd.n1339 31.8661
R6601 gnd.n2590 gnd.n1350 31.8661
R6602 gnd.n2590 gnd.n2111 31.8661
R6603 gnd.n2584 gnd.n2125 31.8661
R6604 gnd.n470 gnd.n458 31.8661
R6605 gnd.n6338 gnd.n490 31.8661
R6606 gnd.n490 gnd.n284 31.8661
R6607 gnd.n6330 gnd.n323 31.8661
R6608 gnd.n6594 gnd.n239 31.8661
R6609 gnd.n6613 gnd.n221 31.8661
R6610 gnd.n6629 gnd.n209 31.8661
R6611 gnd.n6629 gnd.n212 31.8661
R6612 gnd.n6639 gnd.n194 31.8661
R6613 gnd.n6652 gnd.n194 31.8661
R6614 gnd.n6661 gnd.n188 31.8661
R6615 gnd.n6672 gnd.n171 31.8661
R6616 gnd.n6680 gnd.n171 31.8661
R6617 gnd.n7107 gnd.n74 31.8661
R6618 gnd.n7101 gnd.n86 31.8661
R6619 gnd.n7095 gnd.n86 31.8661
R6620 gnd.n7089 gnd.n104 31.8661
R6621 gnd.n7089 gnd.n107 31.8661
R6622 gnd.n7083 gnd.n116 31.8661
R6623 gnd.n7077 gnd.n126 31.8661
R6624 gnd.n7071 gnd.n126 31.8661
R6625 gnd.n7065 gnd.n142 31.8661
R6626 gnd.n7065 gnd.n145 31.8661
R6627 gnd.n7059 gnd.n145 31.8661
R6628 gnd.n7059 gnd.n154 31.8661
R6629 gnd.n7053 gnd.n164 31.8661
R6630 gnd.n1222 gnd.t30 31.5474
R6631 gnd.t44 gnd.n1244 31.5474
R6632 gnd.n6661 gnd.t52 31.5474
R6633 gnd.t67 gnd.n74 31.5474
R6634 gnd.n1184 gnd.t4 30.9101
R6635 gnd.t70 gnd.n1282 30.9101
R6636 gnd.t57 gnd.n221 30.9101
R6637 gnd.n3423 gnd.n3420 29.8151
R6638 gnd.n2873 gnd.n2872 29.8151
R6639 gnd.n3923 gnd.n1309 28.6795
R6640 gnd.n2543 gnd.n1312 28.6795
R6641 gnd.n3917 gnd.n1320 28.6795
R6642 gnd.n2565 gnd.n1323 28.6795
R6643 gnd.n2598 gnd.n1332 28.6795
R6644 gnd.n6329 gnd.n274 28.6795
R6645 gnd.n6323 gnd.n267 28.6795
R6646 gnd.n6549 gnd.n255 28.6795
R6647 gnd.n6565 gnd.n258 28.6795
R6648 gnd.n6553 gnd.n246 28.6795
R6649 gnd.n3903 gnd.n1339 28.0422
R6650 gnd.n6530 gnd.n323 28.0422
R6651 gnd.n2190 gnd.n2189 25.7944
R6652 gnd.n6368 gnd.n6367 25.7944
R6653 gnd.n6721 gnd.n6720 25.7944
R6654 gnd.n6904 gnd.n6903 25.7944
R6655 gnd.n7003 gnd.n7002 25.7944
R6656 gnd.n342 gnd.n341 25.7944
R6657 gnd.n365 gnd.n364 25.7944
R6658 gnd.n387 gnd.n386 25.7944
R6659 gnd.n6736 gnd.n6735 25.7944
R6660 gnd.n4625 gnd.n4624 25.7944
R6661 gnd.n4183 gnd.n4182 25.7944
R6662 gnd.n2195 gnd.n2194 25.7944
R6663 gnd.n2406 gnd.n2405 25.7944
R6664 gnd.n1084 gnd.n1083 25.7944
R6665 gnd.n1106 gnd.n1105 25.7944
R6666 gnd.n1128 gnd.n1127 25.7944
R6667 gnd.n1397 gnd.n1396 25.7944
R6668 gnd.n2201 gnd.n2200 25.7944
R6669 gnd.n2213 gnd.n2212 25.7944
R6670 gnd.n442 gnd.n441 25.7944
R6671 gnd.n4846 gnd.n4566 24.8557
R6672 gnd.n4856 gnd.n4549 24.8557
R6673 gnd.n4552 gnd.n4540 24.8557
R6674 gnd.n4877 gnd.n4541 24.8557
R6675 gnd.n4887 gnd.n4521 24.8557
R6676 gnd.n4897 gnd.n4896 24.8557
R6677 gnd.n4507 gnd.n4505 24.8557
R6678 gnd.n4928 gnd.n4927 24.8557
R6679 gnd.n4943 gnd.n4490 24.8557
R6680 gnd.n4997 gnd.n4429 24.8557
R6681 gnd.n4953 gnd.n4430 24.8557
R6682 gnd.n4990 gnd.n4441 24.8557
R6683 gnd.n4479 gnd.n4478 24.8557
R6684 gnd.n4984 gnd.n4983 24.8557
R6685 gnd.n4465 gnd.n4452 24.8557
R6686 gnd.n5023 gnd.n5022 24.8557
R6687 gnd.n5033 gnd.n4361 24.8557
R6688 gnd.n5045 gnd.n4353 24.8557
R6689 gnd.n5044 gnd.n4341 24.8557
R6690 gnd.n5063 gnd.n5062 24.8557
R6691 gnd.n5073 gnd.n4334 24.8557
R6692 gnd.n5084 gnd.n4322 24.8557
R6693 gnd.n5108 gnd.n5107 24.8557
R6694 gnd.n5119 gnd.n4305 24.8557
R6695 gnd.n5118 gnd.n4307 24.8557
R6696 gnd.n5130 gnd.n4298 24.8557
R6697 gnd.n5148 gnd.n5147 24.8557
R6698 gnd.n4289 gnd.n4278 24.8557
R6699 gnd.n5169 gnd.n4266 24.8557
R6700 gnd.n5197 gnd.n5196 24.8557
R6701 gnd.n5208 gnd.n4251 24.8557
R6702 gnd.n5219 gnd.n4244 24.8557
R6703 gnd.n5218 gnd.n4232 24.8557
R6704 gnd.n5491 gnd.n5490 24.8557
R6705 gnd.n5513 gnd.n4217 24.8557
R6706 gnd.n2660 gnd.n2111 23.8997
R6707 gnd.n6339 gnd.n6338 23.8997
R6708 gnd.n4867 gnd.t139 23.2624
R6709 gnd.n4568 gnd.t262 22.6251
R6710 gnd.n6306 gnd.t9 22.3064
R6711 gnd.n4001 gnd.t46 21.9878
R6712 gnd.n3941 gnd.t42 21.9878
R6713 gnd.n6613 gnd.t20 21.9878
R6714 gnd.n7083 gnd.t106 21.9878
R6715 gnd.t157 gnd.n4573 21.3504
R6716 gnd.n3977 gnd.t16 21.3504
R6717 gnd.n3965 gnd.t32 21.3504
R6718 gnd.n188 gnd.t0 21.3504
R6719 gnd.n7107 gnd.t7 21.3504
R6720 gnd.t178 gnd.n4279 20.7131
R6721 gnd.n3989 gnd.t87 20.7131
R6722 gnd.n3953 gnd.t117 20.7131
R6723 gnd.n6639 gnd.t36 20.7131
R6724 gnd.n7095 gnd.t23 20.7131
R6725 gnd.t176 gnd.n4314 20.0758
R6726 gnd.n4013 gnd.t40 20.0758
R6727 gnd.n7071 gnd.t99 20.0758
R6728 gnd.n1454 gnd.t291 19.8005
R6729 gnd.n1454 gnd.t312 19.8005
R6730 gnd.n1453 gnd.t247 19.8005
R6731 gnd.n1453 gnd.t300 19.8005
R6732 gnd.n1660 gnd.t315 19.8005
R6733 gnd.n1660 gnd.t267 19.8005
R6734 gnd.n1659 gnd.t210 19.8005
R6735 gnd.n1659 gnd.t282 19.8005
R6736 gnd.n1450 gnd.n1449 19.5087
R6737 gnd.n1463 gnd.n1450 19.5087
R6738 gnd.n1461 gnd.n1452 19.5087
R6739 gnd.n1664 gnd.n1658 19.5087
R6740 gnd.n5034 gnd.t188 19.4385
R6741 gnd.n2672 gnd.n2100 19.3944
R6742 gnd.n2672 gnd.n2097 19.3944
R6743 gnd.n2677 gnd.n2097 19.3944
R6744 gnd.n2677 gnd.n2098 19.3944
R6745 gnd.n2098 gnd.n2075 19.3944
R6746 gnd.n2702 gnd.n2075 19.3944
R6747 gnd.n2702 gnd.n2072 19.3944
R6748 gnd.n2707 gnd.n2072 19.3944
R6749 gnd.n2707 gnd.n2073 19.3944
R6750 gnd.n2073 gnd.n2050 19.3944
R6751 gnd.n2732 gnd.n2050 19.3944
R6752 gnd.n2732 gnd.n2047 19.3944
R6753 gnd.n2737 gnd.n2047 19.3944
R6754 gnd.n2737 gnd.n2048 19.3944
R6755 gnd.n2048 gnd.n2025 19.3944
R6756 gnd.n2762 gnd.n2025 19.3944
R6757 gnd.n2762 gnd.n2022 19.3944
R6758 gnd.n2770 gnd.n2022 19.3944
R6759 gnd.n2770 gnd.n2023 19.3944
R6760 gnd.n2766 gnd.n2023 19.3944
R6761 gnd.n2766 gnd.n2001 19.3944
R6762 gnd.n2001 gnd.n1999 19.3944
R6763 gnd.n2878 gnd.n1999 19.3944
R6764 gnd.n2878 gnd.n1996 19.3944
R6765 gnd.n2886 gnd.n1996 19.3944
R6766 gnd.n2886 gnd.n1997 19.3944
R6767 gnd.n2882 gnd.n1997 19.3944
R6768 gnd.n2882 gnd.n1974 19.3944
R6769 gnd.n2946 gnd.n1974 19.3944
R6770 gnd.n2946 gnd.n1972 19.3944
R6771 gnd.n2950 gnd.n1972 19.3944
R6772 gnd.n2950 gnd.n1952 19.3944
R6773 gnd.n2979 gnd.n1952 19.3944
R6774 gnd.n2979 gnd.n1949 19.3944
R6775 gnd.n2993 gnd.n1949 19.3944
R6776 gnd.n2993 gnd.n1950 19.3944
R6777 gnd.n2989 gnd.n1950 19.3944
R6778 gnd.n2989 gnd.n2988 19.3944
R6779 gnd.n2988 gnd.n2987 19.3944
R6780 gnd.n2987 gnd.n1912 19.3944
R6781 gnd.n3079 gnd.n1912 19.3944
R6782 gnd.n3079 gnd.n1909 19.3944
R6783 gnd.n3084 gnd.n1909 19.3944
R6784 gnd.n3084 gnd.n1910 19.3944
R6785 gnd.n1910 gnd.n1882 19.3944
R6786 gnd.n3115 gnd.n1882 19.3944
R6787 gnd.n3115 gnd.n1879 19.3944
R6788 gnd.n3123 gnd.n1879 19.3944
R6789 gnd.n3123 gnd.n1880 19.3944
R6790 gnd.n3119 gnd.n1880 19.3944
R6791 gnd.n3119 gnd.n1853 19.3944
R6792 gnd.n3163 gnd.n1853 19.3944
R6793 gnd.n3163 gnd.n1850 19.3944
R6794 gnd.n3171 gnd.n1850 19.3944
R6795 gnd.n3171 gnd.n1851 19.3944
R6796 gnd.n3167 gnd.n1851 19.3944
R6797 gnd.n3167 gnd.n1816 19.3944
R6798 gnd.n3251 gnd.n1816 19.3944
R6799 gnd.n3251 gnd.n1813 19.3944
R6800 gnd.n3256 gnd.n1813 19.3944
R6801 gnd.n3256 gnd.n1814 19.3944
R6802 gnd.n1814 gnd.n1790 19.3944
R6803 gnd.n3287 gnd.n1790 19.3944
R6804 gnd.n3287 gnd.n1787 19.3944
R6805 gnd.n3297 gnd.n1787 19.3944
R6806 gnd.n3297 gnd.n1788 19.3944
R6807 gnd.n3293 gnd.n1788 19.3944
R6808 gnd.n3293 gnd.n1763 19.3944
R6809 gnd.n3337 gnd.n1763 19.3944
R6810 gnd.n3337 gnd.n1760 19.3944
R6811 gnd.n3345 gnd.n1760 19.3944
R6812 gnd.n3345 gnd.n1761 19.3944
R6813 gnd.n3341 gnd.n1761 19.3944
R6814 gnd.n3341 gnd.n1729 19.3944
R6815 gnd.n3408 gnd.n1729 19.3944
R6816 gnd.n3408 gnd.n1726 19.3944
R6817 gnd.n3413 gnd.n1726 19.3944
R6818 gnd.n3413 gnd.n1727 19.3944
R6819 gnd.n1727 gnd.n1637 19.3944
R6820 gnd.n3556 gnd.n1637 19.3944
R6821 gnd.n3556 gnd.n1635 19.3944
R6822 gnd.n3560 gnd.n1635 19.3944
R6823 gnd.n3560 gnd.n1624 19.3944
R6824 gnd.n3578 gnd.n1624 19.3944
R6825 gnd.n3578 gnd.n1622 19.3944
R6826 gnd.n3582 gnd.n1622 19.3944
R6827 gnd.n3582 gnd.n1613 19.3944
R6828 gnd.n3598 gnd.n1613 19.3944
R6829 gnd.n3598 gnd.n1611 19.3944
R6830 gnd.n3602 gnd.n1611 19.3944
R6831 gnd.n3602 gnd.n1600 19.3944
R6832 gnd.n3618 gnd.n1600 19.3944
R6833 gnd.n3618 gnd.n1598 19.3944
R6834 gnd.n3622 gnd.n1598 19.3944
R6835 gnd.n3622 gnd.n1587 19.3944
R6836 gnd.n3638 gnd.n1587 19.3944
R6837 gnd.n3638 gnd.n1584 19.3944
R6838 gnd.n3643 gnd.n1584 19.3944
R6839 gnd.n3643 gnd.n1585 19.3944
R6840 gnd.n1585 gnd.n454 19.3944
R6841 gnd.n6357 gnd.n454 19.3944
R6842 gnd.n2552 gnd.n2550 19.3944
R6843 gnd.n2557 gnd.n2552 19.3944
R6844 gnd.n2557 gnd.n2556 19.3944
R6845 gnd.n2663 gnd.n2109 19.3944
R6846 gnd.n2658 gnd.n2109 19.3944
R6847 gnd.n2658 gnd.n2127 19.3944
R6848 gnd.n2654 gnd.n2127 19.3944
R6849 gnd.n2654 gnd.n2653 19.3944
R6850 gnd.n2653 gnd.n2652 19.3944
R6851 gnd.n2652 gnd.n2133 19.3944
R6852 gnd.n2647 gnd.n2133 19.3944
R6853 gnd.n2647 gnd.n2646 19.3944
R6854 gnd.n2646 gnd.n2138 19.3944
R6855 gnd.n2639 gnd.n2138 19.3944
R6856 gnd.n2639 gnd.n2638 19.3944
R6857 gnd.n2638 gnd.n2150 19.3944
R6858 gnd.n2631 gnd.n2150 19.3944
R6859 gnd.n2631 gnd.n2630 19.3944
R6860 gnd.n2630 gnd.n2158 19.3944
R6861 gnd.n2623 gnd.n2158 19.3944
R6862 gnd.n2623 gnd.n2622 19.3944
R6863 gnd.n2622 gnd.n2170 19.3944
R6864 gnd.n2615 gnd.n2170 19.3944
R6865 gnd.n2615 gnd.n2614 19.3944
R6866 gnd.n2614 gnd.n2178 19.3944
R6867 gnd.n2607 gnd.n2178 19.3944
R6868 gnd.n2607 gnd.n2606 19.3944
R6869 gnd.n6410 gnd.n398 19.3944
R6870 gnd.n6410 gnd.n6409 19.3944
R6871 gnd.n6409 gnd.n401 19.3944
R6872 gnd.n6402 gnd.n401 19.3944
R6873 gnd.n6402 gnd.n6401 19.3944
R6874 gnd.n6401 gnd.n411 19.3944
R6875 gnd.n6394 gnd.n411 19.3944
R6876 gnd.n6394 gnd.n6393 19.3944
R6877 gnd.n6393 gnd.n419 19.3944
R6878 gnd.n6386 gnd.n419 19.3944
R6879 gnd.n6386 gnd.n6385 19.3944
R6880 gnd.n6385 gnd.n429 19.3944
R6881 gnd.n6378 gnd.n429 19.3944
R6882 gnd.n6378 gnd.n6377 19.3944
R6883 gnd.n6377 gnd.n437 19.3944
R6884 gnd.n6370 gnd.n437 19.3944
R6885 gnd.n504 gnd.n503 19.3944
R6886 gnd.n504 gnd.n264 19.3944
R6887 gnd.n6551 gnd.n264 19.3944
R6888 gnd.n6552 gnd.n6551 19.3944
R6889 gnd.n6555 gnd.n6552 19.3944
R6890 gnd.n6556 gnd.n6555 19.3944
R6891 gnd.n6556 gnd.n236 19.3944
R6892 gnd.n6596 gnd.n236 19.3944
R6893 gnd.n6597 gnd.n6596 19.3944
R6894 gnd.n6598 gnd.n6597 19.3944
R6895 gnd.n6598 gnd.n218 19.3944
R6896 gnd.n6616 gnd.n218 19.3944
R6897 gnd.n6617 gnd.n6616 19.3944
R6898 gnd.n6619 gnd.n6617 19.3944
R6899 gnd.n6620 gnd.n6619 19.3944
R6900 gnd.n6620 gnd.n192 19.3944
R6901 gnd.n6654 gnd.n192 19.3944
R6902 gnd.n6657 gnd.n6654 19.3944
R6903 gnd.n6657 gnd.n6656 19.3944
R6904 gnd.n6656 gnd.n173 19.3944
R6905 gnd.n6677 gnd.n173 19.3944
R6906 gnd.n6678 gnd.n6677 19.3944
R6907 gnd.n6678 gnd.n167 19.3944
R6908 gnd.n6687 gnd.n167 19.3944
R6909 gnd.n6688 gnd.n6687 19.3944
R6910 gnd.n6690 gnd.n6688 19.3944
R6911 gnd.n6691 gnd.n6690 19.3944
R6912 gnd.n6694 gnd.n6691 19.3944
R6913 gnd.n6695 gnd.n6694 19.3944
R6914 gnd.n6697 gnd.n6695 19.3944
R6915 gnd.n6698 gnd.n6697 19.3944
R6916 gnd.n6701 gnd.n6698 19.3944
R6917 gnd.n6702 gnd.n6701 19.3944
R6918 gnd.n6704 gnd.n6702 19.3944
R6919 gnd.n6705 gnd.n6704 19.3944
R6920 gnd.n6708 gnd.n6705 19.3944
R6921 gnd.n6709 gnd.n6708 19.3944
R6922 gnd.n6711 gnd.n6709 19.3944
R6923 gnd.n6712 gnd.n6711 19.3944
R6924 gnd.n6715 gnd.n6712 19.3944
R6925 gnd.n6716 gnd.n6715 19.3944
R6926 gnd.n6717 gnd.n6716 19.3944
R6927 gnd.n6958 gnd.n6902 19.3944
R6928 gnd.n6958 gnd.n6955 19.3944
R6929 gnd.n6955 gnd.n6952 19.3944
R6930 gnd.n6952 gnd.n6951 19.3944
R6931 gnd.n6951 gnd.n6948 19.3944
R6932 gnd.n6948 gnd.n6947 19.3944
R6933 gnd.n6947 gnd.n6944 19.3944
R6934 gnd.n6944 gnd.n6943 19.3944
R6935 gnd.n6943 gnd.n6940 19.3944
R6936 gnd.n6940 gnd.n6939 19.3944
R6937 gnd.n6939 gnd.n6936 19.3944
R6938 gnd.n6936 gnd.n6935 19.3944
R6939 gnd.n6935 gnd.n6932 19.3944
R6940 gnd.n6932 gnd.n6931 19.3944
R6941 gnd.n6931 gnd.n6928 19.3944
R6942 gnd.n6928 gnd.n6927 19.3944
R6943 gnd.n6927 gnd.n6924 19.3944
R6944 gnd.n6924 gnd.n6923 19.3944
R6945 gnd.n7001 gnd.n6998 19.3944
R6946 gnd.n6998 gnd.n6997 19.3944
R6947 gnd.n6997 gnd.n6994 19.3944
R6948 gnd.n6994 gnd.n6993 19.3944
R6949 gnd.n6993 gnd.n6990 19.3944
R6950 gnd.n6990 gnd.n6989 19.3944
R6951 gnd.n6989 gnd.n6986 19.3944
R6952 gnd.n6986 gnd.n6985 19.3944
R6953 gnd.n6985 gnd.n6982 19.3944
R6954 gnd.n6982 gnd.n6981 19.3944
R6955 gnd.n6981 gnd.n6978 19.3944
R6956 gnd.n6978 gnd.n6977 19.3944
R6957 gnd.n6977 gnd.n6974 19.3944
R6958 gnd.n6974 gnd.n6973 19.3944
R6959 gnd.n6973 gnd.n6970 19.3944
R6960 gnd.n6970 gnd.n6969 19.3944
R6961 gnd.n6969 gnd.n6966 19.3944
R6962 gnd.n6966 gnd.n6965 19.3944
R6963 gnd.n7040 gnd.n7039 19.3944
R6964 gnd.n7039 gnd.n6868 19.3944
R6965 gnd.n7035 gnd.n6868 19.3944
R6966 gnd.n7035 gnd.n7032 19.3944
R6967 gnd.n7032 gnd.n7029 19.3944
R6968 gnd.n7029 gnd.n7028 19.3944
R6969 gnd.n7028 gnd.n7025 19.3944
R6970 gnd.n7025 gnd.n7024 19.3944
R6971 gnd.n7024 gnd.n7021 19.3944
R6972 gnd.n7021 gnd.n7020 19.3944
R6973 gnd.n7020 gnd.n7017 19.3944
R6974 gnd.n7017 gnd.n7016 19.3944
R6975 gnd.n7016 gnd.n7013 19.3944
R6976 gnd.n7013 gnd.n7012 19.3944
R6977 gnd.n7012 gnd.n7009 19.3944
R6978 gnd.n7009 gnd.n7008 19.3944
R6979 gnd.n7008 gnd.n7005 19.3944
R6980 gnd.n6538 gnd.n279 19.3944
R6981 gnd.n6538 gnd.n280 19.3944
R6982 gnd.n280 gnd.n253 19.3944
R6983 gnd.n6567 gnd.n253 19.3944
R6984 gnd.n6567 gnd.n251 19.3944
R6985 gnd.n6573 gnd.n251 19.3944
R6986 gnd.n6573 gnd.n6572 19.3944
R6987 gnd.n6572 gnd.n227 19.3944
R6988 gnd.n6607 gnd.n227 19.3944
R6989 gnd.n6607 gnd.n225 19.3944
R6990 gnd.n6611 gnd.n225 19.3944
R6991 gnd.n6611 gnd.n207 19.3944
R6992 gnd.n6631 gnd.n207 19.3944
R6993 gnd.n6631 gnd.n205 19.3944
R6994 gnd.n6637 gnd.n205 19.3944
R6995 gnd.n6637 gnd.n6636 19.3944
R6996 gnd.n6636 gnd.n184 19.3944
R6997 gnd.n6663 gnd.n184 19.3944
R6998 gnd.n6663 gnd.n182 19.3944
R6999 gnd.n6670 gnd.n182 19.3944
R7000 gnd.n6670 gnd.n6669 19.3944
R7001 gnd.n6669 gnd.n78 19.3944
R7002 gnd.n7105 gnd.n78 19.3944
R7003 gnd.n7105 gnd.n7104 19.3944
R7004 gnd.n7104 gnd.n7103 19.3944
R7005 gnd.n7103 gnd.n82 19.3944
R7006 gnd.n7093 gnd.n82 19.3944
R7007 gnd.n7093 gnd.n7092 19.3944
R7008 gnd.n7092 gnd.n7091 19.3944
R7009 gnd.n7091 gnd.n102 19.3944
R7010 gnd.n7081 gnd.n102 19.3944
R7011 gnd.n7081 gnd.n7080 19.3944
R7012 gnd.n7080 gnd.n7079 19.3944
R7013 gnd.n7079 gnd.n122 19.3944
R7014 gnd.n7069 gnd.n122 19.3944
R7015 gnd.n7069 gnd.n7068 19.3944
R7016 gnd.n7068 gnd.n7067 19.3944
R7017 gnd.n7067 gnd.n140 19.3944
R7018 gnd.n7057 gnd.n140 19.3944
R7019 gnd.n7057 gnd.n7056 19.3944
R7020 gnd.n7056 gnd.n7055 19.3944
R7021 gnd.n7055 gnd.n160 19.3944
R7022 gnd.n6533 gnd.n282 19.3944
R7023 gnd.n6528 gnd.n282 19.3944
R7024 gnd.n6528 gnd.n6527 19.3944
R7025 gnd.n6527 gnd.n6526 19.3944
R7026 gnd.n6526 gnd.n6523 19.3944
R7027 gnd.n6523 gnd.n6522 19.3944
R7028 gnd.n6522 gnd.n6519 19.3944
R7029 gnd.n6519 gnd.n6518 19.3944
R7030 gnd.n6518 gnd.n6515 19.3944
R7031 gnd.n6515 gnd.n6514 19.3944
R7032 gnd.n6514 gnd.n6511 19.3944
R7033 gnd.n6511 gnd.n6510 19.3944
R7034 gnd.n6510 gnd.n6507 19.3944
R7035 gnd.n6507 gnd.n6506 19.3944
R7036 gnd.n6506 gnd.n6503 19.3944
R7037 gnd.n6503 gnd.n6502 19.3944
R7038 gnd.n6502 gnd.n6499 19.3944
R7039 gnd.n6497 gnd.n6494 19.3944
R7040 gnd.n6494 gnd.n6493 19.3944
R7041 gnd.n6493 gnd.n6490 19.3944
R7042 gnd.n6490 gnd.n6489 19.3944
R7043 gnd.n6489 gnd.n6486 19.3944
R7044 gnd.n6486 gnd.n6485 19.3944
R7045 gnd.n6485 gnd.n6482 19.3944
R7046 gnd.n6480 gnd.n6477 19.3944
R7047 gnd.n6477 gnd.n6476 19.3944
R7048 gnd.n6476 gnd.n6473 19.3944
R7049 gnd.n6473 gnd.n6472 19.3944
R7050 gnd.n6472 gnd.n6469 19.3944
R7051 gnd.n6469 gnd.n6468 19.3944
R7052 gnd.n6468 gnd.n6465 19.3944
R7053 gnd.n6465 gnd.n6464 19.3944
R7054 gnd.n6460 gnd.n6457 19.3944
R7055 gnd.n6457 gnd.n6456 19.3944
R7056 gnd.n6456 gnd.n6453 19.3944
R7057 gnd.n6453 gnd.n6452 19.3944
R7058 gnd.n6452 gnd.n6449 19.3944
R7059 gnd.n6449 gnd.n6448 19.3944
R7060 gnd.n6448 gnd.n6445 19.3944
R7061 gnd.n6445 gnd.n6444 19.3944
R7062 gnd.n6444 gnd.n6441 19.3944
R7063 gnd.n6441 gnd.n6440 19.3944
R7064 gnd.n6440 gnd.n6437 19.3944
R7065 gnd.n6437 gnd.n6436 19.3944
R7066 gnd.n6436 gnd.n6433 19.3944
R7067 gnd.n6433 gnd.n6432 19.3944
R7068 gnd.n6432 gnd.n6429 19.3944
R7069 gnd.n6429 gnd.n6428 19.3944
R7070 gnd.n6428 gnd.n6425 19.3944
R7071 gnd.n6425 gnd.n6424 19.3944
R7072 gnd.n6747 gnd.n6745 19.3944
R7073 gnd.n6750 gnd.n6747 19.3944
R7074 gnd.n6753 gnd.n6750 19.3944
R7075 gnd.n6756 gnd.n6753 19.3944
R7076 gnd.n6756 gnd.n6743 19.3944
R7077 gnd.n6760 gnd.n6743 19.3944
R7078 gnd.n6763 gnd.n6760 19.3944
R7079 gnd.n6766 gnd.n6763 19.3944
R7080 gnd.n6766 gnd.n6741 19.3944
R7081 gnd.n6770 gnd.n6741 19.3944
R7082 gnd.n6773 gnd.n6770 19.3944
R7083 gnd.n6776 gnd.n6773 19.3944
R7084 gnd.n6776 gnd.n6739 19.3944
R7085 gnd.n6780 gnd.n6739 19.3944
R7086 gnd.n6783 gnd.n6780 19.3944
R7087 gnd.n6785 gnd.n6783 19.3944
R7088 gnd.n6542 gnd.n272 19.3944
R7089 gnd.n6542 gnd.n269 19.3944
R7090 gnd.n6547 gnd.n269 19.3944
R7091 gnd.n6547 gnd.n270 19.3944
R7092 gnd.n270 gnd.n244 19.3944
R7093 gnd.n6577 gnd.n244 19.3944
R7094 gnd.n6577 gnd.n241 19.3944
R7095 gnd.n6592 gnd.n241 19.3944
R7096 gnd.n6592 gnd.n242 19.3944
R7097 gnd.n6588 gnd.n242 19.3944
R7098 gnd.n6588 gnd.n6587 19.3944
R7099 gnd.n6587 gnd.n6586 19.3944
R7100 gnd.n6586 gnd.n6583 19.3944
R7101 gnd.n6583 gnd.n199 19.3944
R7102 gnd.n6641 gnd.n199 19.3944
R7103 gnd.n6641 gnd.n196 19.3944
R7104 gnd.n6650 gnd.n196 19.3944
R7105 gnd.n6650 gnd.n197 19.3944
R7106 gnd.n6646 gnd.n197 19.3944
R7107 gnd.n6646 gnd.n6645 19.3944
R7108 gnd.n6645 gnd.n68 19.3944
R7109 gnd.n7110 gnd.n68 19.3944
R7110 gnd.n7110 gnd.n7109 19.3944
R7111 gnd.n7109 gnd.n71 19.3944
R7112 gnd.n6798 gnd.n71 19.3944
R7113 gnd.n6800 gnd.n6798 19.3944
R7114 gnd.n6800 gnd.n6795 19.3944
R7115 gnd.n6805 gnd.n6795 19.3944
R7116 gnd.n6806 gnd.n6805 19.3944
R7117 gnd.n6808 gnd.n6806 19.3944
R7118 gnd.n6808 gnd.n6793 19.3944
R7119 gnd.n6813 gnd.n6793 19.3944
R7120 gnd.n6814 gnd.n6813 19.3944
R7121 gnd.n6816 gnd.n6814 19.3944
R7122 gnd.n6816 gnd.n6791 19.3944
R7123 gnd.n6821 gnd.n6791 19.3944
R7124 gnd.n6822 gnd.n6821 19.3944
R7125 gnd.n6824 gnd.n6822 19.3944
R7126 gnd.n6824 gnd.n6789 19.3944
R7127 gnd.n6829 gnd.n6789 19.3944
R7128 gnd.n6830 gnd.n6829 19.3944
R7129 gnd.n6831 gnd.n6830 19.3944
R7130 gnd.n6327 gnd.n6326 19.3944
R7131 gnd.n6326 gnd.n6325 19.3944
R7132 gnd.n6325 gnd.n261 19.3944
R7133 gnd.n6563 gnd.n261 19.3944
R7134 gnd.n6563 gnd.n6562 19.3944
R7135 gnd.n6562 gnd.n6561 19.3944
R7136 gnd.n6561 gnd.n6560 19.3944
R7137 gnd.n6560 gnd.n234 19.3944
R7138 gnd.n6603 gnd.n234 19.3944
R7139 gnd.n6603 gnd.n6602 19.3944
R7140 gnd.n6602 gnd.n6601 19.3944
R7141 gnd.n6601 gnd.n215 19.3944
R7142 gnd.n6627 gnd.n215 19.3944
R7143 gnd.n6627 gnd.n6626 19.3944
R7144 gnd.n6626 gnd.n6625 19.3944
R7145 gnd.n6625 gnd.n6624 19.3944
R7146 gnd.n6624 gnd.n190 19.3944
R7147 gnd.n6659 gnd.n190 19.3944
R7148 gnd.n6659 gnd.n175 19.3944
R7149 gnd.n6674 gnd.n175 19.3944
R7150 gnd.n6674 gnd.n169 19.3944
R7151 gnd.n6682 gnd.n169 19.3944
R7152 gnd.n6683 gnd.n6682 19.3944
R7153 gnd.n6683 gnd.n89 19.3944
R7154 gnd.n7099 gnd.n89 19.3944
R7155 gnd.n7099 gnd.n7098 19.3944
R7156 gnd.n7098 gnd.n7097 19.3944
R7157 gnd.n7097 gnd.n93 19.3944
R7158 gnd.n7087 gnd.n93 19.3944
R7159 gnd.n7087 gnd.n7086 19.3944
R7160 gnd.n7086 gnd.n7085 19.3944
R7161 gnd.n7085 gnd.n112 19.3944
R7162 gnd.n7075 gnd.n112 19.3944
R7163 gnd.n7075 gnd.n7074 19.3944
R7164 gnd.n7074 gnd.n7073 19.3944
R7165 gnd.n7073 gnd.n131 19.3944
R7166 gnd.n7063 gnd.n131 19.3944
R7167 gnd.n7063 gnd.n7062 19.3944
R7168 gnd.n7062 gnd.n7061 19.3944
R7169 gnd.n7061 gnd.n150 19.3944
R7170 gnd.n7051 gnd.n150 19.3944
R7171 gnd.n7051 gnd.n7050 19.3944
R7172 gnd.n4749 gnd.n4748 19.3944
R7173 gnd.n4748 gnd.n4747 19.3944
R7174 gnd.n4747 gnd.n4746 19.3944
R7175 gnd.n4746 gnd.n4744 19.3944
R7176 gnd.n4744 gnd.n4741 19.3944
R7177 gnd.n4741 gnd.n4740 19.3944
R7178 gnd.n4740 gnd.n4737 19.3944
R7179 gnd.n4737 gnd.n4736 19.3944
R7180 gnd.n4736 gnd.n4733 19.3944
R7181 gnd.n4733 gnd.n4732 19.3944
R7182 gnd.n4732 gnd.n4729 19.3944
R7183 gnd.n4729 gnd.n4728 19.3944
R7184 gnd.n4728 gnd.n4725 19.3944
R7185 gnd.n4725 gnd.n4724 19.3944
R7186 gnd.n4724 gnd.n4721 19.3944
R7187 gnd.n4721 gnd.n4720 19.3944
R7188 gnd.n4720 gnd.n4717 19.3944
R7189 gnd.n4717 gnd.n4716 19.3944
R7190 gnd.n4716 gnd.n4713 19.3944
R7191 gnd.n4713 gnd.n4712 19.3944
R7192 gnd.n4712 gnd.n4709 19.3944
R7193 gnd.n4709 gnd.n4708 19.3944
R7194 gnd.n4705 gnd.n4704 19.3944
R7195 gnd.n4704 gnd.n4660 19.3944
R7196 gnd.n4755 gnd.n4660 19.3944
R7197 gnd.n5521 gnd.n5520 19.3944
R7198 gnd.n5520 gnd.n5517 19.3944
R7199 gnd.n5517 gnd.n5516 19.3944
R7200 gnd.n5566 gnd.n5565 19.3944
R7201 gnd.n5565 gnd.n5564 19.3944
R7202 gnd.n5564 gnd.n5561 19.3944
R7203 gnd.n5561 gnd.n5560 19.3944
R7204 gnd.n5560 gnd.n5557 19.3944
R7205 gnd.n5557 gnd.n5556 19.3944
R7206 gnd.n5556 gnd.n5553 19.3944
R7207 gnd.n5553 gnd.n5552 19.3944
R7208 gnd.n5552 gnd.n5549 19.3944
R7209 gnd.n5549 gnd.n5548 19.3944
R7210 gnd.n5548 gnd.n5545 19.3944
R7211 gnd.n5545 gnd.n5544 19.3944
R7212 gnd.n5544 gnd.n5541 19.3944
R7213 gnd.n5541 gnd.n5540 19.3944
R7214 gnd.n5540 gnd.n5537 19.3944
R7215 gnd.n5537 gnd.n5536 19.3944
R7216 gnd.n5536 gnd.n5533 19.3944
R7217 gnd.n5533 gnd.n5532 19.3944
R7218 gnd.n5532 gnd.n5529 19.3944
R7219 gnd.n5529 gnd.n5528 19.3944
R7220 gnd.n5528 gnd.n5525 19.3944
R7221 gnd.n5525 gnd.n5524 19.3944
R7222 gnd.n4848 gnd.n4557 19.3944
R7223 gnd.n4858 gnd.n4557 19.3944
R7224 gnd.n4859 gnd.n4858 19.3944
R7225 gnd.n4859 gnd.n4538 19.3944
R7226 gnd.n4879 gnd.n4538 19.3944
R7227 gnd.n4879 gnd.n4530 19.3944
R7228 gnd.n4889 gnd.n4530 19.3944
R7229 gnd.n4890 gnd.n4889 19.3944
R7230 gnd.n4891 gnd.n4890 19.3944
R7231 gnd.n4891 gnd.n4513 19.3944
R7232 gnd.n4908 gnd.n4513 19.3944
R7233 gnd.n4911 gnd.n4908 19.3944
R7234 gnd.n4911 gnd.n4910 19.3944
R7235 gnd.n4910 gnd.n4486 19.3944
R7236 gnd.n4950 gnd.n4486 19.3944
R7237 gnd.n4950 gnd.n4483 19.3944
R7238 gnd.n4956 gnd.n4483 19.3944
R7239 gnd.n4957 gnd.n4956 19.3944
R7240 gnd.n4957 gnd.n4481 19.3944
R7241 gnd.n4963 gnd.n4481 19.3944
R7242 gnd.n4966 gnd.n4963 19.3944
R7243 gnd.n4968 gnd.n4966 19.3944
R7244 gnd.n4974 gnd.n4968 19.3944
R7245 gnd.n4974 gnd.n4973 19.3944
R7246 gnd.n4973 gnd.n4356 19.3944
R7247 gnd.n5040 gnd.n4356 19.3944
R7248 gnd.n5041 gnd.n5040 19.3944
R7249 gnd.n5041 gnd.n4349 19.3944
R7250 gnd.n5052 gnd.n4349 19.3944
R7251 gnd.n5053 gnd.n5052 19.3944
R7252 gnd.n5053 gnd.n4332 19.3944
R7253 gnd.n4332 gnd.n4330 19.3944
R7254 gnd.n5077 gnd.n4330 19.3944
R7255 gnd.n5078 gnd.n5077 19.3944
R7256 gnd.n5078 gnd.n4301 19.3944
R7257 gnd.n5125 gnd.n4301 19.3944
R7258 gnd.n5126 gnd.n5125 19.3944
R7259 gnd.n5126 gnd.n4294 19.3944
R7260 gnd.n5137 gnd.n4294 19.3944
R7261 gnd.n5138 gnd.n5137 19.3944
R7262 gnd.n5138 gnd.n4277 19.3944
R7263 gnd.n4277 gnd.n4275 19.3944
R7264 gnd.n5162 gnd.n4275 19.3944
R7265 gnd.n5163 gnd.n5162 19.3944
R7266 gnd.n5163 gnd.n4247 19.3944
R7267 gnd.n5214 gnd.n4247 19.3944
R7268 gnd.n5215 gnd.n5214 19.3944
R7269 gnd.n5215 gnd.n4240 19.3944
R7270 gnd.n5482 gnd.n4240 19.3944
R7271 gnd.n5483 gnd.n5482 19.3944
R7272 gnd.n5483 gnd.n4221 19.3944
R7273 gnd.n5508 gnd.n4221 19.3944
R7274 gnd.n5508 gnd.n4222 19.3944
R7275 gnd.n4839 gnd.n4838 19.3944
R7276 gnd.n4838 gnd.n4571 19.3944
R7277 gnd.n4594 gnd.n4571 19.3944
R7278 gnd.n4597 gnd.n4594 19.3944
R7279 gnd.n4597 gnd.n4590 19.3944
R7280 gnd.n4601 gnd.n4590 19.3944
R7281 gnd.n4604 gnd.n4601 19.3944
R7282 gnd.n4607 gnd.n4604 19.3944
R7283 gnd.n4607 gnd.n4588 19.3944
R7284 gnd.n4611 gnd.n4588 19.3944
R7285 gnd.n4614 gnd.n4611 19.3944
R7286 gnd.n4617 gnd.n4614 19.3944
R7287 gnd.n4617 gnd.n4586 19.3944
R7288 gnd.n4621 gnd.n4586 19.3944
R7289 gnd.n4844 gnd.n4843 19.3944
R7290 gnd.n4843 gnd.n4547 19.3944
R7291 gnd.n4869 gnd.n4547 19.3944
R7292 gnd.n4869 gnd.n4545 19.3944
R7293 gnd.n4875 gnd.n4545 19.3944
R7294 gnd.n4875 gnd.n4874 19.3944
R7295 gnd.n4874 gnd.n4519 19.3944
R7296 gnd.n4899 gnd.n4519 19.3944
R7297 gnd.n4899 gnd.n4517 19.3944
R7298 gnd.n4903 gnd.n4517 19.3944
R7299 gnd.n4903 gnd.n4497 19.3944
R7300 gnd.n4930 gnd.n4497 19.3944
R7301 gnd.n4930 gnd.n4495 19.3944
R7302 gnd.n4940 gnd.n4495 19.3944
R7303 gnd.n4940 gnd.n4939 19.3944
R7304 gnd.n4939 gnd.n4938 19.3944
R7305 gnd.n4938 gnd.n4444 19.3944
R7306 gnd.n4988 gnd.n4444 19.3944
R7307 gnd.n4988 gnd.n4987 19.3944
R7308 gnd.n4987 gnd.n4986 19.3944
R7309 gnd.n4986 gnd.n4448 19.3944
R7310 gnd.n4468 gnd.n4448 19.3944
R7311 gnd.n4468 gnd.n4366 19.3944
R7312 gnd.n5025 gnd.n4366 19.3944
R7313 gnd.n5025 gnd.n4364 19.3944
R7314 gnd.n5031 gnd.n4364 19.3944
R7315 gnd.n5031 gnd.n5030 19.3944
R7316 gnd.n5030 gnd.n4339 19.3944
R7317 gnd.n5065 gnd.n4339 19.3944
R7318 gnd.n5065 gnd.n4337 19.3944
R7319 gnd.n5071 gnd.n4337 19.3944
R7320 gnd.n5071 gnd.n5070 19.3944
R7321 gnd.n5070 gnd.n4312 19.3944
R7322 gnd.n5110 gnd.n4312 19.3944
R7323 gnd.n5110 gnd.n4310 19.3944
R7324 gnd.n5116 gnd.n4310 19.3944
R7325 gnd.n5116 gnd.n5115 19.3944
R7326 gnd.n5115 gnd.n4284 19.3944
R7327 gnd.n5150 gnd.n4284 19.3944
R7328 gnd.n5150 gnd.n4282 19.3944
R7329 gnd.n5156 gnd.n4282 19.3944
R7330 gnd.n5156 gnd.n5155 19.3944
R7331 gnd.n5155 gnd.n4257 19.3944
R7332 gnd.n5199 gnd.n4257 19.3944
R7333 gnd.n5199 gnd.n4255 19.3944
R7334 gnd.n5205 gnd.n4255 19.3944
R7335 gnd.n5205 gnd.n5204 19.3944
R7336 gnd.n5204 gnd.n4230 19.3944
R7337 gnd.n5493 gnd.n4230 19.3944
R7338 gnd.n5493 gnd.n4228 19.3944
R7339 gnd.n5501 gnd.n4228 19.3944
R7340 gnd.n5501 gnd.n5500 19.3944
R7341 gnd.n5500 gnd.n5499 19.3944
R7342 gnd.n5602 gnd.n5601 19.3944
R7343 gnd.n5601 gnd.n4169 19.3944
R7344 gnd.n5597 gnd.n4169 19.3944
R7345 gnd.n5597 gnd.n5594 19.3944
R7346 gnd.n5594 gnd.n5591 19.3944
R7347 gnd.n5591 gnd.n5590 19.3944
R7348 gnd.n5590 gnd.n5587 19.3944
R7349 gnd.n5587 gnd.n5586 19.3944
R7350 gnd.n5586 gnd.n5583 19.3944
R7351 gnd.n5583 gnd.n5582 19.3944
R7352 gnd.n5582 gnd.n5579 19.3944
R7353 gnd.n5579 gnd.n5578 19.3944
R7354 gnd.n5578 gnd.n5575 19.3944
R7355 gnd.n5575 gnd.n5574 19.3944
R7356 gnd.n4759 gnd.n4658 19.3944
R7357 gnd.n4759 gnd.n4649 19.3944
R7358 gnd.n4772 gnd.n4649 19.3944
R7359 gnd.n4772 gnd.n4647 19.3944
R7360 gnd.n4776 gnd.n4647 19.3944
R7361 gnd.n4776 gnd.n4637 19.3944
R7362 gnd.n4788 gnd.n4637 19.3944
R7363 gnd.n4788 gnd.n4635 19.3944
R7364 gnd.n4822 gnd.n4635 19.3944
R7365 gnd.n4822 gnd.n4821 19.3944
R7366 gnd.n4821 gnd.n4820 19.3944
R7367 gnd.n4820 gnd.n4819 19.3944
R7368 gnd.n4819 gnd.n4816 19.3944
R7369 gnd.n4816 gnd.n4815 19.3944
R7370 gnd.n4815 gnd.n4814 19.3944
R7371 gnd.n4814 gnd.n4812 19.3944
R7372 gnd.n4812 gnd.n4811 19.3944
R7373 gnd.n4811 gnd.n4808 19.3944
R7374 gnd.n4808 gnd.n4807 19.3944
R7375 gnd.n4807 gnd.n4806 19.3944
R7376 gnd.n4806 gnd.n4804 19.3944
R7377 gnd.n4804 gnd.n4503 19.3944
R7378 gnd.n4919 gnd.n4503 19.3944
R7379 gnd.n4919 gnd.n4501 19.3944
R7380 gnd.n4925 gnd.n4501 19.3944
R7381 gnd.n4925 gnd.n4924 19.3944
R7382 gnd.n4924 gnd.n4425 19.3944
R7383 gnd.n4999 gnd.n4425 19.3944
R7384 gnd.n4999 gnd.n4426 19.3944
R7385 gnd.n4473 gnd.n4472 19.3944
R7386 gnd.n4476 gnd.n4475 19.3944
R7387 gnd.n4463 gnd.n4462 19.3944
R7388 gnd.n5018 gnd.n4371 19.3944
R7389 gnd.n5018 gnd.n5017 19.3944
R7390 gnd.n5017 gnd.n5016 19.3944
R7391 gnd.n5016 gnd.n5014 19.3944
R7392 gnd.n5014 gnd.n5013 19.3944
R7393 gnd.n5013 gnd.n5011 19.3944
R7394 gnd.n5011 gnd.n5010 19.3944
R7395 gnd.n5010 gnd.n4320 19.3944
R7396 gnd.n5086 gnd.n4320 19.3944
R7397 gnd.n5086 gnd.n4318 19.3944
R7398 gnd.n5105 gnd.n4318 19.3944
R7399 gnd.n5105 gnd.n5104 19.3944
R7400 gnd.n5104 gnd.n5103 19.3944
R7401 gnd.n5103 gnd.n5101 19.3944
R7402 gnd.n5101 gnd.n5100 19.3944
R7403 gnd.n5100 gnd.n5098 19.3944
R7404 gnd.n5098 gnd.n5097 19.3944
R7405 gnd.n5097 gnd.n4264 19.3944
R7406 gnd.n5171 gnd.n4264 19.3944
R7407 gnd.n5171 gnd.n4262 19.3944
R7408 gnd.n5194 gnd.n4262 19.3944
R7409 gnd.n5194 gnd.n5193 19.3944
R7410 gnd.n5193 gnd.n5192 19.3944
R7411 gnd.n5192 gnd.n5189 19.3944
R7412 gnd.n5189 gnd.n5188 19.3944
R7413 gnd.n5188 gnd.n5186 19.3944
R7414 gnd.n5186 gnd.n5185 19.3944
R7415 gnd.n5185 gnd.n5183 19.3944
R7416 gnd.n5183 gnd.n4216 19.3944
R7417 gnd.n4764 gnd.n4654 19.3944
R7418 gnd.n4764 gnd.n4652 19.3944
R7419 gnd.n4768 gnd.n4652 19.3944
R7420 gnd.n4768 gnd.n4643 19.3944
R7421 gnd.n4780 gnd.n4643 19.3944
R7422 gnd.n4780 gnd.n4641 19.3944
R7423 gnd.n4784 gnd.n4641 19.3944
R7424 gnd.n4784 gnd.n4630 19.3944
R7425 gnd.n4826 gnd.n4630 19.3944
R7426 gnd.n4826 gnd.n4584 19.3944
R7427 gnd.n4832 gnd.n4584 19.3944
R7428 gnd.n4832 gnd.n4831 19.3944
R7429 gnd.n4831 gnd.n4562 19.3944
R7430 gnd.n4853 gnd.n4562 19.3944
R7431 gnd.n4853 gnd.n4555 19.3944
R7432 gnd.n4864 gnd.n4555 19.3944
R7433 gnd.n4864 gnd.n4863 19.3944
R7434 gnd.n4863 gnd.n4536 19.3944
R7435 gnd.n4884 gnd.n4536 19.3944
R7436 gnd.n4884 gnd.n4526 19.3944
R7437 gnd.n4894 gnd.n4526 19.3944
R7438 gnd.n4894 gnd.n4509 19.3944
R7439 gnd.n4915 gnd.n4509 19.3944
R7440 gnd.n4915 gnd.n4914 19.3944
R7441 gnd.n4914 gnd.n4488 19.3944
R7442 gnd.n4945 gnd.n4488 19.3944
R7443 gnd.n4945 gnd.n4433 19.3944
R7444 gnd.n4995 gnd.n4433 19.3944
R7445 gnd.n4995 gnd.n4994 19.3944
R7446 gnd.n4994 gnd.n4993 19.3944
R7447 gnd.n4993 gnd.n4437 19.3944
R7448 gnd.n4455 gnd.n4437 19.3944
R7449 gnd.n4981 gnd.n4455 19.3944
R7450 gnd.n4981 gnd.n4980 19.3944
R7451 gnd.n4980 gnd.n4979 19.3944
R7452 gnd.n4979 gnd.n4459 19.3944
R7453 gnd.n4459 gnd.n4358 19.3944
R7454 gnd.n5036 gnd.n4358 19.3944
R7455 gnd.n5036 gnd.n4351 19.3944
R7456 gnd.n5047 gnd.n4351 19.3944
R7457 gnd.n5047 gnd.n4347 19.3944
R7458 gnd.n5060 gnd.n4347 19.3944
R7459 gnd.n5060 gnd.n5059 19.3944
R7460 gnd.n5059 gnd.n4326 19.3944
R7461 gnd.n5082 gnd.n4326 19.3944
R7462 gnd.n5082 gnd.n5081 19.3944
R7463 gnd.n5081 gnd.n4303 19.3944
R7464 gnd.n5121 gnd.n4303 19.3944
R7465 gnd.n5121 gnd.n4296 19.3944
R7466 gnd.n5132 gnd.n4296 19.3944
R7467 gnd.n5132 gnd.n4292 19.3944
R7468 gnd.n5145 gnd.n4292 19.3944
R7469 gnd.n5145 gnd.n5144 19.3944
R7470 gnd.n5144 gnd.n4271 19.3944
R7471 gnd.n5167 gnd.n4271 19.3944
R7472 gnd.n5167 gnd.n5166 19.3944
R7473 gnd.n5166 gnd.n4249 19.3944
R7474 gnd.n5210 gnd.n4249 19.3944
R7475 gnd.n5210 gnd.n4242 19.3944
R7476 gnd.n5221 gnd.n4242 19.3944
R7477 gnd.n5221 gnd.n4238 19.3944
R7478 gnd.n5488 gnd.n4238 19.3944
R7479 gnd.n5488 gnd.n5487 19.3944
R7480 gnd.n5487 gnd.n4219 19.3944
R7481 gnd.n5511 gnd.n4219 19.3944
R7482 gnd.n2643 gnd.n2140 19.3944
R7483 gnd.n2643 gnd.n2642 19.3944
R7484 gnd.n2642 gnd.n2144 19.3944
R7485 gnd.n2635 gnd.n2144 19.3944
R7486 gnd.n2635 gnd.n2634 19.3944
R7487 gnd.n2634 gnd.n2154 19.3944
R7488 gnd.n2627 gnd.n2154 19.3944
R7489 gnd.n2627 gnd.n2626 19.3944
R7490 gnd.n2626 gnd.n2164 19.3944
R7491 gnd.n2619 gnd.n2164 19.3944
R7492 gnd.n2619 gnd.n2618 19.3944
R7493 gnd.n2618 gnd.n2174 19.3944
R7494 gnd.n2611 gnd.n2174 19.3944
R7495 gnd.n2611 gnd.n2610 19.3944
R7496 gnd.n2610 gnd.n2184 19.3944
R7497 gnd.n2603 gnd.n2184 19.3944
R7498 gnd.n2321 gnd.n1130 19.3944
R7499 gnd.n2324 gnd.n2321 19.3944
R7500 gnd.n2325 gnd.n2324 19.3944
R7501 gnd.n2327 gnd.n2325 19.3944
R7502 gnd.n2328 gnd.n2327 19.3944
R7503 gnd.n2331 gnd.n2328 19.3944
R7504 gnd.n2332 gnd.n2331 19.3944
R7505 gnd.n2334 gnd.n2332 19.3944
R7506 gnd.n2335 gnd.n2334 19.3944
R7507 gnd.n2338 gnd.n2335 19.3944
R7508 gnd.n2339 gnd.n2338 19.3944
R7509 gnd.n2341 gnd.n2339 19.3944
R7510 gnd.n2342 gnd.n2341 19.3944
R7511 gnd.n2345 gnd.n2342 19.3944
R7512 gnd.n2346 gnd.n2345 19.3944
R7513 gnd.n2348 gnd.n2346 19.3944
R7514 gnd.n2349 gnd.n2348 19.3944
R7515 gnd.n2352 gnd.n2349 19.3944
R7516 gnd.n2353 gnd.n2352 19.3944
R7517 gnd.n2355 gnd.n2353 19.3944
R7518 gnd.n2356 gnd.n2355 19.3944
R7519 gnd.n2359 gnd.n2356 19.3944
R7520 gnd.n2360 gnd.n2359 19.3944
R7521 gnd.n2362 gnd.n2360 19.3944
R7522 gnd.n2363 gnd.n2362 19.3944
R7523 gnd.n2366 gnd.n2363 19.3944
R7524 gnd.n2367 gnd.n2366 19.3944
R7525 gnd.n2369 gnd.n2367 19.3944
R7526 gnd.n2370 gnd.n2369 19.3944
R7527 gnd.n2373 gnd.n2370 19.3944
R7528 gnd.n2374 gnd.n2373 19.3944
R7529 gnd.n2376 gnd.n2374 19.3944
R7530 gnd.n2377 gnd.n2376 19.3944
R7531 gnd.n2380 gnd.n2377 19.3944
R7532 gnd.n2381 gnd.n2380 19.3944
R7533 gnd.n2533 gnd.n2381 19.3944
R7534 gnd.n2534 gnd.n2533 19.3944
R7535 gnd.n2541 gnd.n2534 19.3944
R7536 gnd.n2541 gnd.n2540 19.3944
R7537 gnd.n2540 gnd.n2539 19.3944
R7538 gnd.n2539 gnd.n2538 19.3944
R7539 gnd.n2538 gnd.n2537 19.3944
R7540 gnd.n2418 gnd.n2417 19.3944
R7541 gnd.n2421 gnd.n2418 19.3944
R7542 gnd.n2421 gnd.n2415 19.3944
R7543 gnd.n2427 gnd.n2415 19.3944
R7544 gnd.n2428 gnd.n2427 19.3944
R7545 gnd.n2431 gnd.n2428 19.3944
R7546 gnd.n2431 gnd.n2413 19.3944
R7547 gnd.n2437 gnd.n2413 19.3944
R7548 gnd.n2438 gnd.n2437 19.3944
R7549 gnd.n2441 gnd.n2438 19.3944
R7550 gnd.n2441 gnd.n2411 19.3944
R7551 gnd.n2447 gnd.n2411 19.3944
R7552 gnd.n2448 gnd.n2447 19.3944
R7553 gnd.n2451 gnd.n2448 19.3944
R7554 gnd.n2451 gnd.n2407 19.3944
R7555 gnd.n2455 gnd.n2407 19.3944
R7556 gnd.n2462 gnd.n2461 19.3944
R7557 gnd.n2464 gnd.n2462 19.3944
R7558 gnd.n2464 gnd.n2401 19.3944
R7559 gnd.n2469 gnd.n2401 19.3944
R7560 gnd.n2470 gnd.n2469 19.3944
R7561 gnd.n2472 gnd.n2470 19.3944
R7562 gnd.n2472 gnd.n2399 19.3944
R7563 gnd.n2477 gnd.n2399 19.3944
R7564 gnd.n2478 gnd.n2477 19.3944
R7565 gnd.n2480 gnd.n2478 19.3944
R7566 gnd.n2480 gnd.n2397 19.3944
R7567 gnd.n2485 gnd.n2397 19.3944
R7568 gnd.n2486 gnd.n2485 19.3944
R7569 gnd.n2488 gnd.n2486 19.3944
R7570 gnd.n2488 gnd.n2395 19.3944
R7571 gnd.n2493 gnd.n2395 19.3944
R7572 gnd.n2494 gnd.n2493 19.3944
R7573 gnd.n2496 gnd.n2494 19.3944
R7574 gnd.n2496 gnd.n2393 19.3944
R7575 gnd.n2501 gnd.n2393 19.3944
R7576 gnd.n2502 gnd.n2501 19.3944
R7577 gnd.n2504 gnd.n2502 19.3944
R7578 gnd.n2504 gnd.n2390 19.3944
R7579 gnd.n2508 gnd.n2390 19.3944
R7580 gnd.n2509 gnd.n2508 19.3944
R7581 gnd.n2511 gnd.n2509 19.3944
R7582 gnd.n2511 gnd.n2387 19.3944
R7583 gnd.n2515 gnd.n2387 19.3944
R7584 gnd.n2516 gnd.n2515 19.3944
R7585 gnd.n2518 gnd.n2516 19.3944
R7586 gnd.n2518 gnd.n2384 19.3944
R7587 gnd.n2522 gnd.n2384 19.3944
R7588 gnd.n2523 gnd.n2522 19.3944
R7589 gnd.n2525 gnd.n2523 19.3944
R7590 gnd.n2525 gnd.n2382 19.3944
R7591 gnd.n2529 gnd.n2382 19.3944
R7592 gnd.n2529 gnd.n2320 19.3944
R7593 gnd.n2545 gnd.n2320 19.3944
R7594 gnd.n2545 gnd.n2317 19.3944
R7595 gnd.n2563 gnd.n2317 19.3944
R7596 gnd.n2563 gnd.n2318 19.3944
R7597 gnd.n2318 gnd.n2199 19.3944
R7598 gnd.n4154 gnd.n4153 19.3944
R7599 gnd.n4153 gnd.n4152 19.3944
R7600 gnd.n4152 gnd.n4151 19.3944
R7601 gnd.n4151 gnd.n4149 19.3944
R7602 gnd.n4149 gnd.n4146 19.3944
R7603 gnd.n4146 gnd.n4145 19.3944
R7604 gnd.n4145 gnd.n4142 19.3944
R7605 gnd.n4142 gnd.n4141 19.3944
R7606 gnd.n4141 gnd.n4138 19.3944
R7607 gnd.n4138 gnd.n4137 19.3944
R7608 gnd.n4137 gnd.n4134 19.3944
R7609 gnd.n4134 gnd.n4133 19.3944
R7610 gnd.n4133 gnd.n4130 19.3944
R7611 gnd.n4130 gnd.n4129 19.3944
R7612 gnd.n4129 gnd.n4126 19.3944
R7613 gnd.n4126 gnd.n4125 19.3944
R7614 gnd.n4125 gnd.n4122 19.3944
R7615 gnd.n4120 gnd.n4117 19.3944
R7616 gnd.n4117 gnd.n4116 19.3944
R7617 gnd.n4116 gnd.n4113 19.3944
R7618 gnd.n4113 gnd.n4112 19.3944
R7619 gnd.n4112 gnd.n4109 19.3944
R7620 gnd.n4109 gnd.n4108 19.3944
R7621 gnd.n4108 gnd.n4105 19.3944
R7622 gnd.n4105 gnd.n4104 19.3944
R7623 gnd.n4104 gnd.n4101 19.3944
R7624 gnd.n4101 gnd.n4100 19.3944
R7625 gnd.n4100 gnd.n4097 19.3944
R7626 gnd.n4097 gnd.n4096 19.3944
R7627 gnd.n4096 gnd.n4093 19.3944
R7628 gnd.n4093 gnd.n4092 19.3944
R7629 gnd.n4092 gnd.n4089 19.3944
R7630 gnd.n4089 gnd.n4088 19.3944
R7631 gnd.n4088 gnd.n4085 19.3944
R7632 gnd.n4085 gnd.n4084 19.3944
R7633 gnd.n4080 gnd.n4077 19.3944
R7634 gnd.n4077 gnd.n4076 19.3944
R7635 gnd.n4076 gnd.n4073 19.3944
R7636 gnd.n4073 gnd.n4072 19.3944
R7637 gnd.n4072 gnd.n4069 19.3944
R7638 gnd.n4069 gnd.n4068 19.3944
R7639 gnd.n4068 gnd.n4065 19.3944
R7640 gnd.n4065 gnd.n4064 19.3944
R7641 gnd.n4064 gnd.n4061 19.3944
R7642 gnd.n4061 gnd.n4060 19.3944
R7643 gnd.n4060 gnd.n4057 19.3944
R7644 gnd.n4057 gnd.n4056 19.3944
R7645 gnd.n4056 gnd.n4053 19.3944
R7646 gnd.n4053 gnd.n4052 19.3944
R7647 gnd.n4052 gnd.n4049 19.3944
R7648 gnd.n4049 gnd.n4048 19.3944
R7649 gnd.n4048 gnd.n4045 19.3944
R7650 gnd.n4045 gnd.n4044 19.3944
R7651 gnd.n3905 gnd.n1337 19.3944
R7652 gnd.n3900 gnd.n1337 19.3944
R7653 gnd.n3900 gnd.n3899 19.3944
R7654 gnd.n3899 gnd.n3898 19.3944
R7655 gnd.n3898 gnd.n3895 19.3944
R7656 gnd.n3895 gnd.n3894 19.3944
R7657 gnd.n3894 gnd.n3891 19.3944
R7658 gnd.n3891 gnd.n3890 19.3944
R7659 gnd.n3890 gnd.n3887 19.3944
R7660 gnd.n3887 gnd.n3886 19.3944
R7661 gnd.n3886 gnd.n3883 19.3944
R7662 gnd.n3883 gnd.n3882 19.3944
R7663 gnd.n3882 gnd.n3879 19.3944
R7664 gnd.n3879 gnd.n3878 19.3944
R7665 gnd.n3878 gnd.n3875 19.3944
R7666 gnd.n3875 gnd.n3874 19.3944
R7667 gnd.n3874 gnd.n3871 19.3944
R7668 gnd.n2247 gnd.n2244 19.3944
R7669 gnd.n2250 gnd.n2247 19.3944
R7670 gnd.n2250 gnd.n2210 19.3944
R7671 gnd.n2254 gnd.n2210 19.3944
R7672 gnd.n2257 gnd.n2254 19.3944
R7673 gnd.n2260 gnd.n2257 19.3944
R7674 gnd.n2260 gnd.n2208 19.3944
R7675 gnd.n2264 gnd.n2208 19.3944
R7676 gnd.n2267 gnd.n2264 19.3944
R7677 gnd.n2270 gnd.n2267 19.3944
R7678 gnd.n2270 gnd.n2206 19.3944
R7679 gnd.n2274 gnd.n2206 19.3944
R7680 gnd.n2277 gnd.n2274 19.3944
R7681 gnd.n2280 gnd.n2277 19.3944
R7682 gnd.n2280 gnd.n2204 19.3944
R7683 gnd.n2284 gnd.n2204 19.3944
R7684 gnd.n2287 gnd.n2284 19.3944
R7685 gnd.n2290 gnd.n2287 19.3944
R7686 gnd.n2220 gnd.n1406 19.3944
R7687 gnd.n2224 gnd.n2220 19.3944
R7688 gnd.n2227 gnd.n2224 19.3944
R7689 gnd.n2230 gnd.n2227 19.3944
R7690 gnd.n2230 gnd.n2216 19.3944
R7691 gnd.n2234 gnd.n2216 19.3944
R7692 gnd.n2237 gnd.n2234 19.3944
R7693 gnd.n2240 gnd.n2237 19.3944
R7694 gnd.n3869 gnd.n3866 19.3944
R7695 gnd.n3866 gnd.n3865 19.3944
R7696 gnd.n3865 gnd.n3862 19.3944
R7697 gnd.n3862 gnd.n3861 19.3944
R7698 gnd.n3861 gnd.n3858 19.3944
R7699 gnd.n3858 gnd.n3857 19.3944
R7700 gnd.n3857 gnd.n3854 19.3944
R7701 gnd.n4031 gnd.n1140 19.3944
R7702 gnd.n4031 gnd.n1141 19.3944
R7703 gnd.n4027 gnd.n1141 19.3944
R7704 gnd.n4027 gnd.n1144 19.3944
R7705 gnd.n4017 gnd.n1144 19.3944
R7706 gnd.n4017 gnd.n4016 19.3944
R7707 gnd.n4016 gnd.n4015 19.3944
R7708 gnd.n4015 gnd.n1164 19.3944
R7709 gnd.n4005 gnd.n1164 19.3944
R7710 gnd.n4005 gnd.n4004 19.3944
R7711 gnd.n4004 gnd.n4003 19.3944
R7712 gnd.n4003 gnd.n1182 19.3944
R7713 gnd.n3993 gnd.n1182 19.3944
R7714 gnd.n3993 gnd.n3992 19.3944
R7715 gnd.n3992 gnd.n3991 19.3944
R7716 gnd.n3991 gnd.n1202 19.3944
R7717 gnd.n3981 gnd.n1202 19.3944
R7718 gnd.n3981 gnd.n3980 19.3944
R7719 gnd.n3980 gnd.n3979 19.3944
R7720 gnd.n3979 gnd.n1220 19.3944
R7721 gnd.n3969 gnd.n1220 19.3944
R7722 gnd.n3969 gnd.n3968 19.3944
R7723 gnd.n3968 gnd.n3967 19.3944
R7724 gnd.n3967 gnd.n1240 19.3944
R7725 gnd.n3957 gnd.n1240 19.3944
R7726 gnd.n3957 gnd.n3956 19.3944
R7727 gnd.n3956 gnd.n3955 19.3944
R7728 gnd.n3955 gnd.n1259 19.3944
R7729 gnd.n3945 gnd.n1259 19.3944
R7730 gnd.n3945 gnd.n3944 19.3944
R7731 gnd.n3944 gnd.n3943 19.3944
R7732 gnd.n3943 gnd.n1278 19.3944
R7733 gnd.n3933 gnd.n1278 19.3944
R7734 gnd.n3933 gnd.n3932 19.3944
R7735 gnd.n3932 gnd.n3931 19.3944
R7736 gnd.n3931 gnd.n1297 19.3944
R7737 gnd.n3921 gnd.n1297 19.3944
R7738 gnd.n3921 gnd.n3920 19.3944
R7739 gnd.n3920 gnd.n3919 19.3944
R7740 gnd.n3919 gnd.n1318 19.3944
R7741 gnd.n3909 gnd.n1318 19.3944
R7742 gnd.n3909 gnd.n3908 19.3944
R7743 gnd.n4036 gnd.n1132 19.3944
R7744 gnd.n1151 gnd.n1132 19.3944
R7745 gnd.n4023 gnd.n1151 19.3944
R7746 gnd.n4023 gnd.n4022 19.3944
R7747 gnd.n4022 gnd.n4021 19.3944
R7748 gnd.n4021 gnd.n1155 19.3944
R7749 gnd.n4011 gnd.n1155 19.3944
R7750 gnd.n4011 gnd.n4010 19.3944
R7751 gnd.n4010 gnd.n4009 19.3944
R7752 gnd.n4009 gnd.n1173 19.3944
R7753 gnd.n3999 gnd.n1173 19.3944
R7754 gnd.n3999 gnd.n3998 19.3944
R7755 gnd.n3998 gnd.n3997 19.3944
R7756 gnd.n3997 gnd.n1191 19.3944
R7757 gnd.n3987 gnd.n1191 19.3944
R7758 gnd.n3987 gnd.n3986 19.3944
R7759 gnd.n3986 gnd.n3985 19.3944
R7760 gnd.n3985 gnd.n1211 19.3944
R7761 gnd.n3975 gnd.n1211 19.3944
R7762 gnd.n3975 gnd.n3974 19.3944
R7763 gnd.n3974 gnd.n3973 19.3944
R7764 gnd.n3973 gnd.n1229 19.3944
R7765 gnd.n3963 gnd.n1229 19.3944
R7766 gnd.n3963 gnd.n3962 19.3944
R7767 gnd.n3962 gnd.n3961 19.3944
R7768 gnd.n3961 gnd.n1249 19.3944
R7769 gnd.n3951 gnd.n1249 19.3944
R7770 gnd.n3951 gnd.n3950 19.3944
R7771 gnd.n3950 gnd.n3949 19.3944
R7772 gnd.n3949 gnd.n1267 19.3944
R7773 gnd.n3939 gnd.n1267 19.3944
R7774 gnd.n3939 gnd.n3938 19.3944
R7775 gnd.n3938 gnd.n3937 19.3944
R7776 gnd.n3937 gnd.n1287 19.3944
R7777 gnd.n3927 gnd.n1287 19.3944
R7778 gnd.n3927 gnd.n3926 19.3944
R7779 gnd.n3926 gnd.n3925 19.3944
R7780 gnd.n3925 gnd.n1307 19.3944
R7781 gnd.n3915 gnd.n1307 19.3944
R7782 gnd.n3915 gnd.n3914 19.3944
R7783 gnd.n3914 gnd.n3913 19.3944
R7784 gnd.n3913 gnd.n1328 19.3944
R7785 gnd.n2309 gnd.n2306 19.3944
R7786 gnd.n2309 gnd.n2303 19.3944
R7787 gnd.n2313 gnd.n2303 19.3944
R7788 gnd.n2313 gnd.n2301 19.3944
R7789 gnd.n2568 gnd.n2301 19.3944
R7790 gnd.n2568 gnd.n2299 19.3944
R7791 gnd.n2595 gnd.n2299 19.3944
R7792 gnd.n2595 gnd.n2594 19.3944
R7793 gnd.n2594 gnd.n2593 19.3944
R7794 gnd.n2593 gnd.n2574 19.3944
R7795 gnd.n2588 gnd.n2574 19.3944
R7796 gnd.n2588 gnd.n2587 19.3944
R7797 gnd.n2587 gnd.n2586 19.3944
R7798 gnd.n2586 gnd.n2581 19.3944
R7799 gnd.n2581 gnd.n2093 19.3944
R7800 gnd.n2682 gnd.n2093 19.3944
R7801 gnd.n2682 gnd.n2091 19.3944
R7802 gnd.n2688 gnd.n2091 19.3944
R7803 gnd.n2688 gnd.n2687 19.3944
R7804 gnd.n2687 gnd.n2068 19.3944
R7805 gnd.n2712 gnd.n2068 19.3944
R7806 gnd.n2712 gnd.n2066 19.3944
R7807 gnd.n2718 gnd.n2066 19.3944
R7808 gnd.n2718 gnd.n2717 19.3944
R7809 gnd.n2717 gnd.n2043 19.3944
R7810 gnd.n2742 gnd.n2043 19.3944
R7811 gnd.n2742 gnd.n2041 19.3944
R7812 gnd.n2748 gnd.n2041 19.3944
R7813 gnd.n2748 gnd.n2747 19.3944
R7814 gnd.n2747 gnd.n2018 19.3944
R7815 gnd.n2775 gnd.n2018 19.3944
R7816 gnd.n2775 gnd.n2016 19.3944
R7817 gnd.n2793 gnd.n2016 19.3944
R7818 gnd.n2793 gnd.n2792 19.3944
R7819 gnd.n2792 gnd.n2791 19.3944
R7820 gnd.n2791 gnd.n2781 19.3944
R7821 gnd.n2787 gnd.n2781 19.3944
R7822 gnd.n2787 gnd.n2786 19.3944
R7823 gnd.n2786 gnd.n1988 19.3944
R7824 gnd.n2927 gnd.n1988 19.3944
R7825 gnd.n2927 gnd.n1986 19.3944
R7826 gnd.n2933 gnd.n1986 19.3944
R7827 gnd.n2933 gnd.n2932 19.3944
R7828 gnd.n2932 gnd.n1960 19.3944
R7829 gnd.n2969 gnd.n1960 19.3944
R7830 gnd.n2969 gnd.n1958 19.3944
R7831 gnd.n2973 gnd.n1958 19.3944
R7832 gnd.n2973 gnd.n1937 19.3944
R7833 gnd.n3013 gnd.n1937 19.3944
R7834 gnd.n3013 gnd.n1935 19.3944
R7835 gnd.n3017 gnd.n1935 19.3944
R7836 gnd.n3017 gnd.n1919 19.3944
R7837 gnd.n3069 gnd.n1919 19.3944
R7838 gnd.n3069 gnd.n1917 19.3944
R7839 gnd.n3073 gnd.n1917 19.3944
R7840 gnd.n3073 gnd.n1897 19.3944
R7841 gnd.n3097 gnd.n1897 19.3944
R7842 gnd.n3097 gnd.n1895 19.3944
R7843 gnd.n3103 gnd.n1895 19.3944
R7844 gnd.n3103 gnd.n3102 19.3944
R7845 gnd.n3102 gnd.n1865 19.3944
R7846 gnd.n3142 gnd.n1865 19.3944
R7847 gnd.n3142 gnd.n1863 19.3944
R7848 gnd.n3146 gnd.n1863 19.3944
R7849 gnd.n3146 gnd.n1841 19.3944
R7850 gnd.n3183 gnd.n1841 19.3944
R7851 gnd.n3183 gnd.n1839 19.3944
R7852 gnd.n3187 gnd.n1839 19.3944
R7853 gnd.n3187 gnd.n1824 19.3944
R7854 gnd.n3242 gnd.n1824 19.3944
R7855 gnd.n3242 gnd.n1822 19.3944
R7856 gnd.n3246 gnd.n1822 19.3944
R7857 gnd.n3246 gnd.n1803 19.3944
R7858 gnd.n3269 gnd.n1803 19.3944
R7859 gnd.n3269 gnd.n1801 19.3944
R7860 gnd.n3275 gnd.n1801 19.3944
R7861 gnd.n3275 gnd.n3274 19.3944
R7862 gnd.n3274 gnd.n1774 19.3944
R7863 gnd.n3316 gnd.n1774 19.3944
R7864 gnd.n3316 gnd.n1772 19.3944
R7865 gnd.n3320 gnd.n1772 19.3944
R7866 gnd.n3320 gnd.n1751 19.3944
R7867 gnd.n3357 gnd.n1751 19.3944
R7868 gnd.n3357 gnd.n1749 19.3944
R7869 gnd.n3361 gnd.n1749 19.3944
R7870 gnd.n3361 gnd.n1735 19.3944
R7871 gnd.n3399 gnd.n1735 19.3944
R7872 gnd.n3399 gnd.n1733 19.3944
R7873 gnd.n3403 gnd.n1733 19.3944
R7874 gnd.n3403 gnd.n1643 19.3944
R7875 gnd.n3546 gnd.n1643 19.3944
R7876 gnd.n3546 gnd.n1641 19.3944
R7877 gnd.n3550 gnd.n1641 19.3944
R7878 gnd.n3550 gnd.n1630 19.3944
R7879 gnd.n3566 gnd.n1630 19.3944
R7880 gnd.n3566 gnd.n1628 19.3944
R7881 gnd.n3570 gnd.n1628 19.3944
R7882 gnd.n3570 gnd.n1619 19.3944
R7883 gnd.n3588 gnd.n1619 19.3944
R7884 gnd.n3588 gnd.n1617 19.3944
R7885 gnd.n3592 gnd.n1617 19.3944
R7886 gnd.n3592 gnd.n1606 19.3944
R7887 gnd.n3608 gnd.n1606 19.3944
R7888 gnd.n3608 gnd.n1604 19.3944
R7889 gnd.n3612 gnd.n1604 19.3944
R7890 gnd.n3612 gnd.n1593 19.3944
R7891 gnd.n3628 gnd.n1593 19.3944
R7892 gnd.n3628 gnd.n1591 19.3944
R7893 gnd.n3632 gnd.n1591 19.3944
R7894 gnd.n3632 gnd.n1579 19.3944
R7895 gnd.n3648 gnd.n1579 19.3944
R7896 gnd.n3648 gnd.n1577 19.3944
R7897 gnd.n3658 gnd.n1577 19.3944
R7898 gnd.n3658 gnd.n3657 19.3944
R7899 gnd.n3657 gnd.n3656 19.3944
R7900 gnd.n3656 gnd.n493 19.3944
R7901 gnd.n6336 gnd.n493 19.3944
R7902 gnd.n6336 gnd.n6335 19.3944
R7903 gnd.n6335 gnd.n6334 19.3944
R7904 gnd.n6334 gnd.n497 19.3944
R7905 gnd.n499 gnd.n497 19.3944
R7906 gnd.n508 gnd.n499 19.3944
R7907 gnd.n6320 gnd.n508 19.3944
R7908 gnd.n6320 gnd.n6319 19.3944
R7909 gnd.n6319 gnd.n6318 19.3944
R7910 gnd.n6318 gnd.n515 19.3944
R7911 gnd.n6314 gnd.n515 19.3944
R7912 gnd.n6314 gnd.n6313 19.3944
R7913 gnd.n6100 gnd.n645 19.3944
R7914 gnd.n6100 gnd.n641 19.3944
R7915 gnd.n6106 gnd.n641 19.3944
R7916 gnd.n6106 gnd.n639 19.3944
R7917 gnd.n6110 gnd.n639 19.3944
R7918 gnd.n6110 gnd.n635 19.3944
R7919 gnd.n6116 gnd.n635 19.3944
R7920 gnd.n6116 gnd.n633 19.3944
R7921 gnd.n6120 gnd.n633 19.3944
R7922 gnd.n6120 gnd.n629 19.3944
R7923 gnd.n6126 gnd.n629 19.3944
R7924 gnd.n6126 gnd.n627 19.3944
R7925 gnd.n6130 gnd.n627 19.3944
R7926 gnd.n6130 gnd.n623 19.3944
R7927 gnd.n6136 gnd.n623 19.3944
R7928 gnd.n6136 gnd.n621 19.3944
R7929 gnd.n6140 gnd.n621 19.3944
R7930 gnd.n6140 gnd.n617 19.3944
R7931 gnd.n6146 gnd.n617 19.3944
R7932 gnd.n6146 gnd.n615 19.3944
R7933 gnd.n6150 gnd.n615 19.3944
R7934 gnd.n6150 gnd.n611 19.3944
R7935 gnd.n6156 gnd.n611 19.3944
R7936 gnd.n6156 gnd.n609 19.3944
R7937 gnd.n6160 gnd.n609 19.3944
R7938 gnd.n6160 gnd.n605 19.3944
R7939 gnd.n6166 gnd.n605 19.3944
R7940 gnd.n6166 gnd.n603 19.3944
R7941 gnd.n6170 gnd.n603 19.3944
R7942 gnd.n6170 gnd.n599 19.3944
R7943 gnd.n6176 gnd.n599 19.3944
R7944 gnd.n6176 gnd.n597 19.3944
R7945 gnd.n6180 gnd.n597 19.3944
R7946 gnd.n6180 gnd.n593 19.3944
R7947 gnd.n6186 gnd.n593 19.3944
R7948 gnd.n6186 gnd.n591 19.3944
R7949 gnd.n6190 gnd.n591 19.3944
R7950 gnd.n6190 gnd.n587 19.3944
R7951 gnd.n6196 gnd.n587 19.3944
R7952 gnd.n6196 gnd.n585 19.3944
R7953 gnd.n6200 gnd.n585 19.3944
R7954 gnd.n6200 gnd.n581 19.3944
R7955 gnd.n6206 gnd.n581 19.3944
R7956 gnd.n6206 gnd.n579 19.3944
R7957 gnd.n6210 gnd.n579 19.3944
R7958 gnd.n6210 gnd.n575 19.3944
R7959 gnd.n6216 gnd.n575 19.3944
R7960 gnd.n6216 gnd.n573 19.3944
R7961 gnd.n6220 gnd.n573 19.3944
R7962 gnd.n6220 gnd.n569 19.3944
R7963 gnd.n6226 gnd.n569 19.3944
R7964 gnd.n6226 gnd.n567 19.3944
R7965 gnd.n6230 gnd.n567 19.3944
R7966 gnd.n6230 gnd.n563 19.3944
R7967 gnd.n6236 gnd.n563 19.3944
R7968 gnd.n6236 gnd.n561 19.3944
R7969 gnd.n6240 gnd.n561 19.3944
R7970 gnd.n6240 gnd.n557 19.3944
R7971 gnd.n6246 gnd.n557 19.3944
R7972 gnd.n6246 gnd.n555 19.3944
R7973 gnd.n6250 gnd.n555 19.3944
R7974 gnd.n6250 gnd.n551 19.3944
R7975 gnd.n6256 gnd.n551 19.3944
R7976 gnd.n6256 gnd.n549 19.3944
R7977 gnd.n6260 gnd.n549 19.3944
R7978 gnd.n6260 gnd.n545 19.3944
R7979 gnd.n6266 gnd.n545 19.3944
R7980 gnd.n6266 gnd.n543 19.3944
R7981 gnd.n6270 gnd.n543 19.3944
R7982 gnd.n6270 gnd.n539 19.3944
R7983 gnd.n6276 gnd.n539 19.3944
R7984 gnd.n6276 gnd.n537 19.3944
R7985 gnd.n6280 gnd.n537 19.3944
R7986 gnd.n6280 gnd.n533 19.3944
R7987 gnd.n6286 gnd.n533 19.3944
R7988 gnd.n6286 gnd.n531 19.3944
R7989 gnd.n6290 gnd.n531 19.3944
R7990 gnd.n6290 gnd.n527 19.3944
R7991 gnd.n6296 gnd.n527 19.3944
R7992 gnd.n6296 gnd.n525 19.3944
R7993 gnd.n6302 gnd.n525 19.3944
R7994 gnd.n6302 gnd.n6301 19.3944
R7995 gnd.n6301 gnd.n521 19.3944
R7996 gnd.n6310 gnd.n521 19.3944
R7997 gnd.n5776 gnd.n837 19.3944
R7998 gnd.n5780 gnd.n837 19.3944
R7999 gnd.n5780 gnd.n833 19.3944
R8000 gnd.n5786 gnd.n833 19.3944
R8001 gnd.n5786 gnd.n831 19.3944
R8002 gnd.n5790 gnd.n831 19.3944
R8003 gnd.n5790 gnd.n827 19.3944
R8004 gnd.n5796 gnd.n827 19.3944
R8005 gnd.n5796 gnd.n825 19.3944
R8006 gnd.n5800 gnd.n825 19.3944
R8007 gnd.n5800 gnd.n821 19.3944
R8008 gnd.n5806 gnd.n821 19.3944
R8009 gnd.n5806 gnd.n819 19.3944
R8010 gnd.n5810 gnd.n819 19.3944
R8011 gnd.n5810 gnd.n815 19.3944
R8012 gnd.n5816 gnd.n815 19.3944
R8013 gnd.n5816 gnd.n813 19.3944
R8014 gnd.n5820 gnd.n813 19.3944
R8015 gnd.n5820 gnd.n809 19.3944
R8016 gnd.n5826 gnd.n809 19.3944
R8017 gnd.n5826 gnd.n807 19.3944
R8018 gnd.n5830 gnd.n807 19.3944
R8019 gnd.n5830 gnd.n803 19.3944
R8020 gnd.n5836 gnd.n803 19.3944
R8021 gnd.n5836 gnd.n801 19.3944
R8022 gnd.n5840 gnd.n801 19.3944
R8023 gnd.n5840 gnd.n797 19.3944
R8024 gnd.n5846 gnd.n797 19.3944
R8025 gnd.n5846 gnd.n795 19.3944
R8026 gnd.n5850 gnd.n795 19.3944
R8027 gnd.n5850 gnd.n791 19.3944
R8028 gnd.n5856 gnd.n791 19.3944
R8029 gnd.n5856 gnd.n789 19.3944
R8030 gnd.n5860 gnd.n789 19.3944
R8031 gnd.n5860 gnd.n785 19.3944
R8032 gnd.n5866 gnd.n785 19.3944
R8033 gnd.n5866 gnd.n783 19.3944
R8034 gnd.n5870 gnd.n783 19.3944
R8035 gnd.n5870 gnd.n779 19.3944
R8036 gnd.n5876 gnd.n779 19.3944
R8037 gnd.n5876 gnd.n777 19.3944
R8038 gnd.n5880 gnd.n777 19.3944
R8039 gnd.n5880 gnd.n773 19.3944
R8040 gnd.n5886 gnd.n773 19.3944
R8041 gnd.n5886 gnd.n771 19.3944
R8042 gnd.n5890 gnd.n771 19.3944
R8043 gnd.n5890 gnd.n767 19.3944
R8044 gnd.n5896 gnd.n767 19.3944
R8045 gnd.n5896 gnd.n765 19.3944
R8046 gnd.n5900 gnd.n765 19.3944
R8047 gnd.n5900 gnd.n761 19.3944
R8048 gnd.n5906 gnd.n761 19.3944
R8049 gnd.n5906 gnd.n759 19.3944
R8050 gnd.n5910 gnd.n759 19.3944
R8051 gnd.n5910 gnd.n755 19.3944
R8052 gnd.n5916 gnd.n755 19.3944
R8053 gnd.n5916 gnd.n753 19.3944
R8054 gnd.n5920 gnd.n753 19.3944
R8055 gnd.n5920 gnd.n749 19.3944
R8056 gnd.n5926 gnd.n749 19.3944
R8057 gnd.n5926 gnd.n747 19.3944
R8058 gnd.n5930 gnd.n747 19.3944
R8059 gnd.n5930 gnd.n743 19.3944
R8060 gnd.n5936 gnd.n743 19.3944
R8061 gnd.n5936 gnd.n741 19.3944
R8062 gnd.n5940 gnd.n741 19.3944
R8063 gnd.n5940 gnd.n737 19.3944
R8064 gnd.n5946 gnd.n737 19.3944
R8065 gnd.n5946 gnd.n735 19.3944
R8066 gnd.n5950 gnd.n735 19.3944
R8067 gnd.n5950 gnd.n731 19.3944
R8068 gnd.n5956 gnd.n731 19.3944
R8069 gnd.n5956 gnd.n729 19.3944
R8070 gnd.n5960 gnd.n729 19.3944
R8071 gnd.n5960 gnd.n725 19.3944
R8072 gnd.n5966 gnd.n725 19.3944
R8073 gnd.n5966 gnd.n723 19.3944
R8074 gnd.n5970 gnd.n723 19.3944
R8075 gnd.n5970 gnd.n719 19.3944
R8076 gnd.n5976 gnd.n719 19.3944
R8077 gnd.n5976 gnd.n717 19.3944
R8078 gnd.n5980 gnd.n717 19.3944
R8079 gnd.n5980 gnd.n713 19.3944
R8080 gnd.n5986 gnd.n713 19.3944
R8081 gnd.n5986 gnd.n711 19.3944
R8082 gnd.n5990 gnd.n711 19.3944
R8083 gnd.n5990 gnd.n707 19.3944
R8084 gnd.n5996 gnd.n707 19.3944
R8085 gnd.n5996 gnd.n705 19.3944
R8086 gnd.n6000 gnd.n705 19.3944
R8087 gnd.n6000 gnd.n701 19.3944
R8088 gnd.n6006 gnd.n701 19.3944
R8089 gnd.n6006 gnd.n699 19.3944
R8090 gnd.n6010 gnd.n699 19.3944
R8091 gnd.n6010 gnd.n695 19.3944
R8092 gnd.n6016 gnd.n695 19.3944
R8093 gnd.n6016 gnd.n693 19.3944
R8094 gnd.n6020 gnd.n693 19.3944
R8095 gnd.n6020 gnd.n689 19.3944
R8096 gnd.n6026 gnd.n689 19.3944
R8097 gnd.n6026 gnd.n687 19.3944
R8098 gnd.n6030 gnd.n687 19.3944
R8099 gnd.n6030 gnd.n683 19.3944
R8100 gnd.n6036 gnd.n683 19.3944
R8101 gnd.n6036 gnd.n681 19.3944
R8102 gnd.n6040 gnd.n681 19.3944
R8103 gnd.n6040 gnd.n677 19.3944
R8104 gnd.n6046 gnd.n677 19.3944
R8105 gnd.n6046 gnd.n675 19.3944
R8106 gnd.n6050 gnd.n675 19.3944
R8107 gnd.n6050 gnd.n671 19.3944
R8108 gnd.n6056 gnd.n671 19.3944
R8109 gnd.n6056 gnd.n669 19.3944
R8110 gnd.n6060 gnd.n669 19.3944
R8111 gnd.n6060 gnd.n665 19.3944
R8112 gnd.n6066 gnd.n665 19.3944
R8113 gnd.n6066 gnd.n663 19.3944
R8114 gnd.n6070 gnd.n663 19.3944
R8115 gnd.n6070 gnd.n659 19.3944
R8116 gnd.n6076 gnd.n659 19.3944
R8117 gnd.n6076 gnd.n657 19.3944
R8118 gnd.n6080 gnd.n657 19.3944
R8119 gnd.n6080 gnd.n653 19.3944
R8120 gnd.n6086 gnd.n653 19.3944
R8121 gnd.n6086 gnd.n651 19.3944
R8122 gnd.n6090 gnd.n651 19.3944
R8123 gnd.n6090 gnd.n647 19.3944
R8124 gnd.n6096 gnd.n647 19.3944
R8125 gnd.n5770 gnd.n842 19.3944
R8126 gnd.n5770 gnd.n5769 19.3944
R8127 gnd.n5769 gnd.n5768 19.3944
R8128 gnd.n5768 gnd.n846 19.3944
R8129 gnd.n5762 gnd.n846 19.3944
R8130 gnd.n5762 gnd.n5761 19.3944
R8131 gnd.n5761 gnd.n5760 19.3944
R8132 gnd.n5760 gnd.n854 19.3944
R8133 gnd.n5754 gnd.n854 19.3944
R8134 gnd.n5754 gnd.n5753 19.3944
R8135 gnd.n5753 gnd.n5752 19.3944
R8136 gnd.n5752 gnd.n862 19.3944
R8137 gnd.n5746 gnd.n862 19.3944
R8138 gnd.n5746 gnd.n5745 19.3944
R8139 gnd.n5745 gnd.n5744 19.3944
R8140 gnd.n5744 gnd.n870 19.3944
R8141 gnd.n5738 gnd.n870 19.3944
R8142 gnd.n5738 gnd.n5737 19.3944
R8143 gnd.n5737 gnd.n5736 19.3944
R8144 gnd.n5736 gnd.n878 19.3944
R8145 gnd.n5730 gnd.n878 19.3944
R8146 gnd.n5730 gnd.n5729 19.3944
R8147 gnd.n5729 gnd.n5728 19.3944
R8148 gnd.n5728 gnd.n886 19.3944
R8149 gnd.n5722 gnd.n886 19.3944
R8150 gnd.n5722 gnd.n5721 19.3944
R8151 gnd.n5721 gnd.n5720 19.3944
R8152 gnd.n5720 gnd.n894 19.3944
R8153 gnd.n5714 gnd.n894 19.3944
R8154 gnd.n5714 gnd.n5713 19.3944
R8155 gnd.n5713 gnd.n5712 19.3944
R8156 gnd.n5712 gnd.n902 19.3944
R8157 gnd.n5706 gnd.n902 19.3944
R8158 gnd.n5706 gnd.n5705 19.3944
R8159 gnd.n5705 gnd.n5704 19.3944
R8160 gnd.n5704 gnd.n910 19.3944
R8161 gnd.n5698 gnd.n910 19.3944
R8162 gnd.n5698 gnd.n5697 19.3944
R8163 gnd.n5697 gnd.n5696 19.3944
R8164 gnd.n5696 gnd.n918 19.3944
R8165 gnd.n5690 gnd.n918 19.3944
R8166 gnd.n5690 gnd.n5689 19.3944
R8167 gnd.n5689 gnd.n5688 19.3944
R8168 gnd.n5688 gnd.n926 19.3944
R8169 gnd.n5682 gnd.n926 19.3944
R8170 gnd.n5682 gnd.n5681 19.3944
R8171 gnd.n5681 gnd.n5680 19.3944
R8172 gnd.n5680 gnd.n934 19.3944
R8173 gnd.n5674 gnd.n934 19.3944
R8174 gnd.n5674 gnd.n5673 19.3944
R8175 gnd.n5673 gnd.n5672 19.3944
R8176 gnd.n5672 gnd.n942 19.3944
R8177 gnd.n5666 gnd.n942 19.3944
R8178 gnd.n5666 gnd.n5665 19.3944
R8179 gnd.n5665 gnd.n5664 19.3944
R8180 gnd.n5664 gnd.n950 19.3944
R8181 gnd.n5658 gnd.n950 19.3944
R8182 gnd.n5658 gnd.n5657 19.3944
R8183 gnd.n5657 gnd.n5656 19.3944
R8184 gnd.n5656 gnd.n958 19.3944
R8185 gnd.n5650 gnd.n958 19.3944
R8186 gnd.n5650 gnd.n5649 19.3944
R8187 gnd.n5649 gnd.n5648 19.3944
R8188 gnd.n5648 gnd.n966 19.3944
R8189 gnd.n5642 gnd.n966 19.3944
R8190 gnd.n5642 gnd.n5641 19.3944
R8191 gnd.n5641 gnd.n5640 19.3944
R8192 gnd.n5640 gnd.n974 19.3944
R8193 gnd.n5634 gnd.n974 19.3944
R8194 gnd.n5634 gnd.n5633 19.3944
R8195 gnd.n5633 gnd.n5632 19.3944
R8196 gnd.n5632 gnd.n982 19.3944
R8197 gnd.n5626 gnd.n982 19.3944
R8198 gnd.n5626 gnd.n5625 19.3944
R8199 gnd.n5625 gnd.n5624 19.3944
R8200 gnd.n5624 gnd.n990 19.3944
R8201 gnd.n5618 gnd.n990 19.3944
R8202 gnd.n5618 gnd.n5617 19.3944
R8203 gnd.n5617 gnd.n5616 19.3944
R8204 gnd.n5616 gnd.n998 19.3944
R8205 gnd.n5610 gnd.n998 19.3944
R8206 gnd.n5610 gnd.n5609 19.3944
R8207 gnd.n5609 gnd.n5608 19.3944
R8208 gnd.n5608 gnd.n1006 19.3944
R8209 gnd.n2668 gnd.n2106 19.3944
R8210 gnd.n2668 gnd.n2107 19.3944
R8211 gnd.n2107 gnd.n2084 19.3944
R8212 gnd.n2693 gnd.n2084 19.3944
R8213 gnd.n2693 gnd.n2081 19.3944
R8214 gnd.n2698 gnd.n2081 19.3944
R8215 gnd.n2698 gnd.n2082 19.3944
R8216 gnd.n2082 gnd.n2059 19.3944
R8217 gnd.n2723 gnd.n2059 19.3944
R8218 gnd.n2723 gnd.n2056 19.3944
R8219 gnd.n2728 gnd.n2056 19.3944
R8220 gnd.n2728 gnd.n2057 19.3944
R8221 gnd.n2057 gnd.n2033 19.3944
R8222 gnd.n2753 gnd.n2033 19.3944
R8223 gnd.n2753 gnd.n2030 19.3944
R8224 gnd.n2758 gnd.n2030 19.3944
R8225 gnd.n2758 gnd.n2031 19.3944
R8226 gnd.n2031 gnd.n2009 19.3944
R8227 gnd.n2798 gnd.n2009 19.3944
R8228 gnd.n2798 gnd.n2006 19.3944
R8229 gnd.n2803 gnd.n2006 19.3944
R8230 gnd.n2803 gnd.n2007 19.3944
R8231 gnd.n2007 gnd.n1477 19.3944
R8232 gnd.n3776 gnd.n1477 19.3944
R8233 gnd.n3776 gnd.n1478 19.3944
R8234 gnd.n3772 gnd.n1478 19.3944
R8235 gnd.n3772 gnd.n3771 19.3944
R8236 gnd.n3771 gnd.n3770 19.3944
R8237 gnd.n3770 gnd.n1484 19.3944
R8238 gnd.n3766 gnd.n1484 19.3944
R8239 gnd.n3766 gnd.n3765 19.3944
R8240 gnd.n3765 gnd.n3764 19.3944
R8241 gnd.n3764 gnd.n1489 19.3944
R8242 gnd.n3760 gnd.n1489 19.3944
R8243 gnd.n3760 gnd.n3759 19.3944
R8244 gnd.n3759 gnd.n3758 19.3944
R8245 gnd.n3758 gnd.n1494 19.3944
R8246 gnd.n3754 gnd.n1494 19.3944
R8247 gnd.n3754 gnd.n3753 19.3944
R8248 gnd.n3753 gnd.n3752 19.3944
R8249 gnd.n3752 gnd.n1499 19.3944
R8250 gnd.n3748 gnd.n1499 19.3944
R8251 gnd.n3748 gnd.n3747 19.3944
R8252 gnd.n3747 gnd.n3746 19.3944
R8253 gnd.n3746 gnd.n1504 19.3944
R8254 gnd.n3742 gnd.n1504 19.3944
R8255 gnd.n3742 gnd.n3741 19.3944
R8256 gnd.n3741 gnd.n3740 19.3944
R8257 gnd.n3740 gnd.n1509 19.3944
R8258 gnd.n3736 gnd.n1509 19.3944
R8259 gnd.n3736 gnd.n3735 19.3944
R8260 gnd.n3735 gnd.n3734 19.3944
R8261 gnd.n3734 gnd.n1514 19.3944
R8262 gnd.n3730 gnd.n1514 19.3944
R8263 gnd.n3730 gnd.n3729 19.3944
R8264 gnd.n3729 gnd.n3728 19.3944
R8265 gnd.n3728 gnd.n1519 19.3944
R8266 gnd.n3724 gnd.n1519 19.3944
R8267 gnd.n3724 gnd.n3723 19.3944
R8268 gnd.n3723 gnd.n3722 19.3944
R8269 gnd.n3722 gnd.n1524 19.3944
R8270 gnd.n3718 gnd.n1524 19.3944
R8271 gnd.n3718 gnd.n3717 19.3944
R8272 gnd.n3717 gnd.n3716 19.3944
R8273 gnd.n3716 gnd.n1529 19.3944
R8274 gnd.n3712 gnd.n1529 19.3944
R8275 gnd.n3712 gnd.n3711 19.3944
R8276 gnd.n3711 gnd.n3710 19.3944
R8277 gnd.n3710 gnd.n1534 19.3944
R8278 gnd.n3706 gnd.n1534 19.3944
R8279 gnd.n3706 gnd.n3705 19.3944
R8280 gnd.n3705 gnd.n3704 19.3944
R8281 gnd.n3704 gnd.n1539 19.3944
R8282 gnd.n3700 gnd.n1539 19.3944
R8283 gnd.n3700 gnd.n3699 19.3944
R8284 gnd.n3699 gnd.n3698 19.3944
R8285 gnd.n3698 gnd.n1544 19.3944
R8286 gnd.n3694 gnd.n1544 19.3944
R8287 gnd.n3694 gnd.n3693 19.3944
R8288 gnd.n3693 gnd.n3692 19.3944
R8289 gnd.n3692 gnd.n1549 19.3944
R8290 gnd.n3688 gnd.n1549 19.3944
R8291 gnd.n3688 gnd.n3687 19.3944
R8292 gnd.n3687 gnd.n3686 19.3944
R8293 gnd.n3686 gnd.n1554 19.3944
R8294 gnd.n3682 gnd.n1554 19.3944
R8295 gnd.n3682 gnd.n3681 19.3944
R8296 gnd.n3681 gnd.n3680 19.3944
R8297 gnd.n3680 gnd.n1559 19.3944
R8298 gnd.n3676 gnd.n1559 19.3944
R8299 gnd.n3676 gnd.n3675 19.3944
R8300 gnd.n3675 gnd.n3674 19.3944
R8301 gnd.n3674 gnd.n1564 19.3944
R8302 gnd.n3670 gnd.n1564 19.3944
R8303 gnd.n3670 gnd.n3669 19.3944
R8304 gnd.n3669 gnd.n3668 19.3944
R8305 gnd.n3668 gnd.n1569 19.3944
R8306 gnd.n3664 gnd.n1569 19.3944
R8307 gnd.n3664 gnd.n3663 19.3944
R8308 gnd.n3663 gnd.n461 19.3944
R8309 gnd.n6353 gnd.n461 19.3944
R8310 gnd.n6350 gnd.n6349 19.3944
R8311 gnd.n6349 gnd.n6348 19.3944
R8312 gnd.n6348 gnd.n466 19.3944
R8313 gnd.n6344 gnd.n466 19.3944
R8314 gnd.n6344 gnd.n6343 19.3944
R8315 gnd.n6343 gnd.n391 19.3944
R8316 gnd.n6415 gnd.n391 19.3944
R8317 gnd.n6415 gnd.n6414 19.3944
R8318 gnd.n6414 gnd.n6413 19.3944
R8319 gnd.n6413 gnd.n395 19.3944
R8320 gnd.n6406 gnd.n395 19.3944
R8321 gnd.n6406 gnd.n6405 19.3944
R8322 gnd.n6405 gnd.n405 19.3944
R8323 gnd.n6398 gnd.n405 19.3944
R8324 gnd.n6398 gnd.n6397 19.3944
R8325 gnd.n6397 gnd.n415 19.3944
R8326 gnd.n6390 gnd.n415 19.3944
R8327 gnd.n6390 gnd.n6389 19.3944
R8328 gnd.n6389 gnd.n423 19.3944
R8329 gnd.n6382 gnd.n423 19.3944
R8330 gnd.n6382 gnd.n6381 19.3944
R8331 gnd.n6381 gnd.n433 19.3944
R8332 gnd.n6374 gnd.n433 19.3944
R8333 gnd.n6374 gnd.n6373 19.3944
R8334 gnd.n6363 gnd.n449 19.3944
R8335 gnd.n6363 gnd.n6362 19.3944
R8336 gnd.n6362 gnd.n452 19.3944
R8337 gnd.n5606 gnd.n5605 19.3895
R8338 gnd.n4991 gnd.t182 18.8012
R8339 gnd.n4976 gnd.t2 18.8012
R8340 gnd.n4835 gnd.n4834 18.4825
R8341 gnd.n6482 gnd.n6481 18.4247
R8342 gnd.n3854 gnd.n3853 18.4247
R8343 gnd.n6370 gnd.n6369 18.2308
R8344 gnd.n6785 gnd.n6737 18.2308
R8345 gnd.n2603 gnd.n2602 18.2308
R8346 gnd.n2456 gnd.n2455 18.2308
R8347 gnd.t179 gnd.n4515 18.1639
R8348 gnd.n3935 gnd.n1291 18.1639
R8349 gnd.n6605 gnd.n229 18.1639
R8350 gnd.n3783 gnd.n3782 17.6395
R8351 gnd.n3541 gnd.n3540 17.6395
R8352 gnd.n4543 gnd.t189 17.5266
R8353 gnd.n4942 gnd.t66 16.8893
R8354 gnd.n4033 gnd.t227 16.8893
R8355 gnd.t28 gnd.n1302 16.8893
R8356 gnd.n3911 gnd.t231 16.8893
R8357 gnd.n6540 gnd.t215 16.8893
R8358 gnd.n516 gnd.t50 16.8893
R8359 gnd.n7053 gnd.t205 16.8893
R8360 gnd.n6965 gnd.n6962 16.6793
R8361 gnd.n6464 gnd.n6461 16.6793
R8362 gnd.n4084 gnd.n4081 16.6793
R8363 gnd.n2240 gnd.n2214 16.6793
R8364 gnd.n4770 gnd.t302 16.2519
R8365 gnd.n4470 gnd.t177 16.2519
R8366 gnd.n2810 gnd.n2809 16.0975
R8367 gnd.n1699 gnd.n1698 16.0975
R8368 gnd.n3785 gnd.n3784 16.0975
R8369 gnd.n1693 gnd.n1692 16.0975
R8370 gnd.n2584 gnd.n2583 15.9333
R8371 gnd.n2583 gnd.n2102 15.9333
R8372 gnd.n2670 gnd.n2102 15.9333
R8373 gnd.n2670 gnd.n2103 15.9333
R8374 gnd.n2680 gnd.n2095 15.9333
R8375 gnd.n2680 gnd.n2679 15.9333
R8376 gnd.n2679 gnd.n2086 15.9333
R8377 gnd.n2691 gnd.n2086 15.9333
R8378 gnd.n2691 gnd.n2690 15.9333
R8379 gnd.n2690 gnd.n2088 15.9333
R8380 gnd.n2088 gnd.n2077 15.9333
R8381 gnd.n2700 gnd.n2077 15.9333
R8382 gnd.n2700 gnd.n2078 15.9333
R8383 gnd.n2710 gnd.n2070 15.9333
R8384 gnd.n2710 gnd.n2709 15.9333
R8385 gnd.n2709 gnd.n2061 15.9333
R8386 gnd.n2721 gnd.n2061 15.9333
R8387 gnd.n2721 gnd.n2720 15.9333
R8388 gnd.n2720 gnd.n2063 15.9333
R8389 gnd.n2063 gnd.n2052 15.9333
R8390 gnd.n2730 gnd.n2052 15.9333
R8391 gnd.n2053 gnd.n2045 15.9333
R8392 gnd.n2740 gnd.n2045 15.9333
R8393 gnd.n2740 gnd.n2739 15.9333
R8394 gnd.n2739 gnd.n2035 15.9333
R8395 gnd.n2751 gnd.n2035 15.9333
R8396 gnd.n2751 gnd.n2750 15.9333
R8397 gnd.n2750 gnd.n2037 15.9333
R8398 gnd.n2039 gnd.n2037 15.9333
R8399 gnd.n2760 gnd.n2027 15.9333
R8400 gnd.n2027 gnd.n2020 15.9333
R8401 gnd.n2773 gnd.n2020 15.9333
R8402 gnd.n2773 gnd.n2772 15.9333
R8403 gnd.n2772 gnd.n2011 15.9333
R8404 gnd.n2796 gnd.n2011 15.9333
R8405 gnd.n2796 gnd.n2795 15.9333
R8406 gnd.n2795 gnd.n2013 15.9333
R8407 gnd.n2805 gnd.n2002 15.9333
R8408 gnd.n2805 gnd.n2003 15.9333
R8409 gnd.n2003 gnd.n1413 15.9333
R8410 gnd.n2876 gnd.n1445 15.9333
R8411 gnd.n3778 gnd.n1474 15.9333
R8412 gnd.n2917 gnd.n2916 15.9333
R8413 gnd.n2908 gnd.n1982 15.9333
R8414 gnd.n2977 gnd.n2975 15.9333
R8415 gnd.n3019 gnd.n1933 15.9333
R8416 gnd.n3067 gnd.n1921 15.9333
R8417 gnd.n3077 gnd.n3075 15.9333
R8418 gnd.n3087 gnd.n3086 15.9333
R8419 gnd.n3037 gnd.n1891 15.9333
R8420 gnd.n3148 gnd.n1859 15.9333
R8421 gnd.n3148 gnd.n1861 15.9333
R8422 gnd.n3240 gnd.n1826 15.9333
R8423 gnd.n3249 gnd.n3248 15.9333
R8424 gnd.n3259 gnd.n3258 15.9333
R8425 gnd.n3210 gnd.n3209 15.9333
R8426 gnd.n3199 gnd.n1794 15.9333
R8427 gnd.n3322 gnd.n1770 15.9333
R8428 gnd.n3397 gnd.n1738 15.9333
R8429 gnd.n3406 gnd.n3405 15.9333
R8430 gnd.n3416 gnd.n1723 15.9333
R8431 gnd.n1671 gnd.n1646 15.9333
R8432 gnd.n3552 gnd.n1639 15.9333
R8433 gnd.n3554 gnd.n3552 15.9333
R8434 gnd.n3554 gnd.n3553 15.9333
R8435 gnd.n3564 gnd.n1633 15.9333
R8436 gnd.n3564 gnd.n3563 15.9333
R8437 gnd.n3563 gnd.n3562 15.9333
R8438 gnd.n3562 gnd.n1626 15.9333
R8439 gnd.n3572 gnd.n1626 15.9333
R8440 gnd.n3576 gnd.n3572 15.9333
R8441 gnd.n3576 gnd.n3575 15.9333
R8442 gnd.n3575 gnd.n3574 15.9333
R8443 gnd.n3586 gnd.n3585 15.9333
R8444 gnd.n3585 gnd.n3584 15.9333
R8445 gnd.n3584 gnd.n1615 15.9333
R8446 gnd.n3594 gnd.n1615 15.9333
R8447 gnd.n3596 gnd.n3594 15.9333
R8448 gnd.n3596 gnd.n3595 15.9333
R8449 gnd.n3595 gnd.n1609 15.9333
R8450 gnd.n3606 gnd.n1609 15.9333
R8451 gnd.n3605 gnd.n3604 15.9333
R8452 gnd.n3604 gnd.n1602 15.9333
R8453 gnd.n3614 gnd.n1602 15.9333
R8454 gnd.n3616 gnd.n3614 15.9333
R8455 gnd.n3616 gnd.n3615 15.9333
R8456 gnd.n3615 gnd.n1596 15.9333
R8457 gnd.n3626 gnd.n1596 15.9333
R8458 gnd.n3626 gnd.n3625 15.9333
R8459 gnd.n3624 gnd.n1589 15.9333
R8460 gnd.n3634 gnd.n1589 15.9333
R8461 gnd.n3636 gnd.n3634 15.9333
R8462 gnd.n3636 gnd.n3635 15.9333
R8463 gnd.n3635 gnd.n1582 15.9333
R8464 gnd.n3646 gnd.n1582 15.9333
R8465 gnd.n3646 gnd.n3645 15.9333
R8466 gnd.n3645 gnd.n1572 15.9333
R8467 gnd.n3661 gnd.n1572 15.9333
R8468 gnd.n3660 gnd.n1574 15.9333
R8469 gnd.n1574 gnd.n457 15.9333
R8470 gnd.n6355 gnd.n457 15.9333
R8471 gnd.n6355 gnd.n458 15.9333
R8472 gnd.n5457 gnd.n5455 15.6674
R8473 gnd.n5425 gnd.n5423 15.6674
R8474 gnd.n5393 gnd.n5391 15.6674
R8475 gnd.n5362 gnd.n5360 15.6674
R8476 gnd.n5330 gnd.n5328 15.6674
R8477 gnd.n5298 gnd.n5296 15.6674
R8478 gnd.n5266 gnd.n5264 15.6674
R8479 gnd.n5235 gnd.n5233 15.6674
R8480 gnd.n4761 gnd.t302 15.6146
R8481 gnd.t219 gnd.n4224 15.6146
R8482 gnd.t320 gnd.n4225 15.6146
R8483 gnd.n7046 gnd.n6722 15.3217
R8484 gnd.n6421 gnd.n385 15.3217
R8485 gnd.n4041 gnd.n1126 15.3217
R8486 gnd.n2294 gnd.n2202 15.3217
R8487 gnd.n3779 gnd.n1471 15.296
R8488 gnd.n2967 gnd.t95 15.296
R8489 gnd.n3048 gnd.n1914 15.296
R8490 gnd.n3095 gnd.n1899 15.296
R8491 gnd.n3221 gnd.n1818 15.296
R8492 gnd.n3267 gnd.n1805 15.296
R8493 gnd.n3355 gnd.t175 15.296
R8494 gnd.n1654 gnd.n1653 15.0827
R8495 gnd.n1457 gnd.n1452 15.0481
R8496 gnd.n1664 gnd.n1663 15.0481
R8497 gnd.n5129 gnd.t187 14.9773
R8498 gnd.n1146 gnd.t227 14.9773
R8499 gnd.n2013 gnd.t195 14.9773
R8500 gnd.t61 gnd.n1633 14.9773
R8501 gnd.t205 gnd.n154 14.9773
R8502 gnd.n2915 gnd.t239 14.6587
R8503 gnd.n2952 gnd.n1962 14.6587
R8504 gnd.n3010 gnd.n1940 14.6587
R8505 gnd.n3300 gnd.n1776 14.6587
R8506 gnd.n3354 gnd.n1754 14.6587
R8507 gnd.t235 gnd.n1731 14.6587
R8508 gnd.t38 gnd.n4267 14.34
R8509 gnd.n5207 gnd.t65 14.34
R8510 gnd.n3380 gnd.n3379 14.0214
R8511 gnd.n4917 gnd.t137 13.7027
R8512 gnd.n1299 gnd.n1291 13.7027
R8513 gnd.n6594 gnd.n229 13.7027
R8514 gnd.n4627 gnd.n4626 13.5763
R8515 gnd.n5571 gnd.n4181 13.5763
R8516 gnd.n4835 gnd.n4573 13.384
R8517 gnd.n2944 gnd.n2942 13.384
R8518 gnd.n3020 gnd.n1928 13.384
R8519 gnd.n3113 gnd.n3112 13.384
R8520 gnd.t77 gnd.n1886 13.384
R8521 gnd.t75 gnd.n3139 13.384
R8522 gnd.n3161 gnd.t153 13.384
R8523 gnd.n3189 gnd.t80 13.384
R8524 gnd.n3190 gnd.n1834 13.384
R8525 gnd.n3285 gnd.n3284 13.384
R8526 gnd.n3364 gnd.n1744 13.384
R8527 gnd.n1468 gnd.n1449 13.1884
R8528 gnd.n1463 gnd.n1462 13.1884
R8529 gnd.n1462 gnd.n1461 13.1884
R8530 gnd.n1657 gnd.n1652 13.1884
R8531 gnd.n1658 gnd.n1657 13.1884
R8532 gnd.n1464 gnd.n1451 13.146
R8533 gnd.n1460 gnd.n1451 13.146
R8534 gnd.n1656 gnd.n1655 13.146
R8535 gnd.n1656 gnd.n1651 13.146
R8536 gnd.n5458 gnd.n5454 12.8005
R8537 gnd.n5426 gnd.n5422 12.8005
R8538 gnd.n5394 gnd.n5390 12.8005
R8539 gnd.n5363 gnd.n5359 12.8005
R8540 gnd.n5331 gnd.n5327 12.8005
R8541 gnd.n5299 gnd.n5295 12.8005
R8542 gnd.n5267 gnd.n5263 12.8005
R8543 gnd.n5236 gnd.n5232 12.8005
R8544 gnd.n3004 gnd.n3003 12.7467
R8545 gnd.n3030 gnd.n1876 12.7467
R8546 gnd.n3174 gnd.n1847 12.7467
R8547 gnd.n3200 gnd.n1784 12.7467
R8548 gnd.t82 gnd.n2070 12.4281
R8549 gnd.n3625 gnd.t59 12.4281
R8550 gnd.n4626 gnd.n4621 12.4126
R8551 gnd.n5574 gnd.n5571 12.4126
R8552 gnd.n3846 gnd.n3783 12.1761
R8553 gnd.n3540 gnd.n3539 12.1761
R8554 gnd.n2909 gnd.n1991 12.1094
R8555 gnd.n3066 gnd.n1923 12.1094
R8556 gnd.n3038 gnd.n1901 12.1094
R8557 gnd.n3239 gnd.n1829 12.1094
R8558 gnd.n3211 gnd.n3208 12.1094
R8559 gnd.n3396 gnd.t314 12.1094
R8560 gnd.n5462 gnd.n5461 12.0247
R8561 gnd.n5430 gnd.n5429 12.0247
R8562 gnd.n5398 gnd.n5397 12.0247
R8563 gnd.n5367 gnd.n5366 12.0247
R8564 gnd.n5335 gnd.n5334 12.0247
R8565 gnd.n5303 gnd.n5302 12.0247
R8566 gnd.n5271 gnd.n5270 12.0247
R8567 gnd.n5240 gnd.n5239 12.0247
R8568 gnd.t40 gnd.n1159 11.7908
R8569 gnd.n2531 gnd.t28 11.7908
R8570 gnd.n2566 gnd.t231 11.7908
R8571 gnd.n6322 gnd.t215 11.7908
R8572 gnd.n6575 gnd.t50 11.7908
R8573 gnd.n142 gnd.t99 11.7908
R8574 gnd.t246 gnd.n2935 11.4721
R8575 gnd.n2965 gnd.n1964 11.4721
R8576 gnd.n2957 gnd.t18 11.4721
R8577 gnd.n2996 gnd.n1946 11.4721
R8578 gnd.n3137 gnd.n1870 11.4721
R8579 gnd.n3160 gnd.n1855 11.4721
R8580 gnd.n3312 gnd.n1779 11.4721
R8581 gnd.n3291 gnd.t147 11.4721
R8582 gnd.n3333 gnd.n1765 11.4721
R8583 gnd.n5465 gnd.n5452 11.249
R8584 gnd.n5433 gnd.n5420 11.249
R8585 gnd.n5401 gnd.n5388 11.249
R8586 gnd.n5370 gnd.n5357 11.249
R8587 gnd.n5338 gnd.n5325 11.249
R8588 gnd.n5306 gnd.n5293 11.249
R8589 gnd.n5274 gnd.n5261 11.249
R8590 gnd.n5243 gnd.n5230 11.249
R8591 gnd.n4905 gnd.t137 11.1535
R8592 gnd.t87 gnd.n1196 11.1535
R8593 gnd.n1269 gnd.t117 11.1535
R8594 gnd.n2039 gnd.t171 11.1535
R8595 gnd.n3586 gnd.t155 11.1535
R8596 gnd.n212 gnd.t36 11.1535
R8597 gnd.n104 gnd.t23 11.1535
R8598 gnd.n3088 gnd.n1905 10.8348
R8599 gnd.n1820 gnd.n1819 10.8348
R8600 gnd.n3388 gnd.n3387 10.8348
R8601 gnd.n6923 gnd.n6722 10.6672
R8602 gnd.n6424 gnd.n6421 10.6672
R8603 gnd.n4044 gnd.n4041 10.6672
R8604 gnd.n2290 gnd.n2202 10.6672
R8605 gnd.n3475 gnd.n1696 10.6151
R8606 gnd.n3475 gnd.n3474 10.6151
R8607 gnd.n3472 gnd.n1700 10.6151
R8608 gnd.n3467 gnd.n1700 10.6151
R8609 gnd.n3467 gnd.n3466 10.6151
R8610 gnd.n3466 gnd.n3465 10.6151
R8611 gnd.n3465 gnd.n1703 10.6151
R8612 gnd.n3460 gnd.n1703 10.6151
R8613 gnd.n3460 gnd.n3459 10.6151
R8614 gnd.n3459 gnd.n3458 10.6151
R8615 gnd.n3458 gnd.n1706 10.6151
R8616 gnd.n3453 gnd.n1706 10.6151
R8617 gnd.n3453 gnd.n3452 10.6151
R8618 gnd.n3452 gnd.n3451 10.6151
R8619 gnd.n3451 gnd.n1709 10.6151
R8620 gnd.n3446 gnd.n1709 10.6151
R8621 gnd.n3446 gnd.n3445 10.6151
R8622 gnd.n3445 gnd.n3444 10.6151
R8623 gnd.n3444 gnd.n1712 10.6151
R8624 gnd.n3439 gnd.n1712 10.6151
R8625 gnd.n3439 gnd.n3438 10.6151
R8626 gnd.n3438 gnd.n3437 10.6151
R8627 gnd.n3437 gnd.n1715 10.6151
R8628 gnd.n3432 gnd.n1715 10.6151
R8629 gnd.n3432 gnd.n3431 10.6151
R8630 gnd.n3431 gnd.n3430 10.6151
R8631 gnd.n3430 gnd.n1718 10.6151
R8632 gnd.n3425 gnd.n1718 10.6151
R8633 gnd.n3425 gnd.n3424 10.6151
R8634 gnd.n3424 gnd.n3423 10.6151
R8635 gnd.n2873 gnd.n1995 10.6151
R8636 gnd.n2891 gnd.n1995 10.6151
R8637 gnd.n2892 gnd.n2891 10.6151
R8638 gnd.n2913 gnd.n2892 10.6151
R8639 gnd.n2913 gnd.n2912 10.6151
R8640 gnd.n2912 gnd.n2911 10.6151
R8641 gnd.n2911 gnd.n2907 10.6151
R8642 gnd.n2907 gnd.n2906 10.6151
R8643 gnd.n2906 gnd.n2904 10.6151
R8644 gnd.n2904 gnd.n2903 10.6151
R8645 gnd.n2903 gnd.n2899 10.6151
R8646 gnd.n2899 gnd.n2898 10.6151
R8647 gnd.n2898 gnd.n2896 10.6151
R8648 gnd.n2896 gnd.n2895 10.6151
R8649 gnd.n2895 gnd.n2893 10.6151
R8650 gnd.n2893 gnd.n1944 10.6151
R8651 gnd.n2998 gnd.n1944 10.6151
R8652 gnd.n2999 gnd.n2998 10.6151
R8653 gnd.n3000 gnd.n2999 10.6151
R8654 gnd.n3000 gnd.n1930 10.6151
R8655 gnd.n3022 gnd.n1930 10.6151
R8656 gnd.n3023 gnd.n3022 10.6151
R8657 gnd.n3053 gnd.n3023 10.6151
R8658 gnd.n3053 gnd.n3052 10.6151
R8659 gnd.n3052 gnd.n3051 10.6151
R8660 gnd.n3051 gnd.n3024 10.6151
R8661 gnd.n3045 gnd.n3024 10.6151
R8662 gnd.n3045 gnd.n3044 10.6151
R8663 gnd.n3044 gnd.n3043 10.6151
R8664 gnd.n3043 gnd.n3041 10.6151
R8665 gnd.n3041 gnd.n3040 10.6151
R8666 gnd.n3040 gnd.n3036 10.6151
R8667 gnd.n3036 gnd.n3035 10.6151
R8668 gnd.n3035 gnd.n3033 10.6151
R8669 gnd.n3033 gnd.n3032 10.6151
R8670 gnd.n3032 gnd.n3028 10.6151
R8671 gnd.n3028 gnd.n3027 10.6151
R8672 gnd.n3027 gnd.n3025 10.6151
R8673 gnd.n3025 gnd.n1857 10.6151
R8674 gnd.n3150 gnd.n1857 10.6151
R8675 gnd.n3151 gnd.n3150 10.6151
R8676 gnd.n3158 gnd.n3151 10.6151
R8677 gnd.n3158 gnd.n3157 10.6151
R8678 gnd.n3157 gnd.n3156 10.6151
R8679 gnd.n3156 gnd.n1836 10.6151
R8680 gnd.n3192 gnd.n1836 10.6151
R8681 gnd.n3193 gnd.n3192 10.6151
R8682 gnd.n3226 gnd.n3193 10.6151
R8683 gnd.n3226 gnd.n3225 10.6151
R8684 gnd.n3225 gnd.n3224 10.6151
R8685 gnd.n3224 gnd.n3194 10.6151
R8686 gnd.n3218 gnd.n3194 10.6151
R8687 gnd.n3218 gnd.n3217 10.6151
R8688 gnd.n3217 gnd.n3216 10.6151
R8689 gnd.n3216 gnd.n3214 10.6151
R8690 gnd.n3214 gnd.n3213 10.6151
R8691 gnd.n3213 gnd.n3206 10.6151
R8692 gnd.n3206 gnd.n3205 10.6151
R8693 gnd.n3205 gnd.n3203 10.6151
R8694 gnd.n3203 gnd.n3202 10.6151
R8695 gnd.n3202 gnd.n3198 10.6151
R8696 gnd.n3198 gnd.n3197 10.6151
R8697 gnd.n3197 gnd.n3195 10.6151
R8698 gnd.n3195 gnd.n1767 10.6151
R8699 gnd.n3324 gnd.n1767 10.6151
R8700 gnd.n3325 gnd.n3324 10.6151
R8701 gnd.n3331 gnd.n3325 10.6151
R8702 gnd.n3331 gnd.n3330 10.6151
R8703 gnd.n3330 gnd.n3329 10.6151
R8704 gnd.n3329 gnd.n1746 10.6151
R8705 gnd.n3366 gnd.n1746 10.6151
R8706 gnd.n3367 gnd.n3366 10.6151
R8707 gnd.n3377 gnd.n3367 10.6151
R8708 gnd.n3377 gnd.n3376 10.6151
R8709 gnd.n3376 gnd.n3375 10.6151
R8710 gnd.n3375 gnd.n3368 10.6151
R8711 gnd.n3369 gnd.n3368 10.6151
R8712 gnd.n3369 gnd.n1721 10.6151
R8713 gnd.n3419 gnd.n1721 10.6151
R8714 gnd.n3420 gnd.n3419 10.6151
R8715 gnd.n2811 gnd.n1409 10.6151
R8716 gnd.n2814 gnd.n2811 10.6151
R8717 gnd.n2819 gnd.n2816 10.6151
R8718 gnd.n2820 gnd.n2819 10.6151
R8719 gnd.n2823 gnd.n2820 10.6151
R8720 gnd.n2824 gnd.n2823 10.6151
R8721 gnd.n2827 gnd.n2824 10.6151
R8722 gnd.n2828 gnd.n2827 10.6151
R8723 gnd.n2831 gnd.n2828 10.6151
R8724 gnd.n2832 gnd.n2831 10.6151
R8725 gnd.n2835 gnd.n2832 10.6151
R8726 gnd.n2836 gnd.n2835 10.6151
R8727 gnd.n2839 gnd.n2836 10.6151
R8728 gnd.n2840 gnd.n2839 10.6151
R8729 gnd.n2843 gnd.n2840 10.6151
R8730 gnd.n2844 gnd.n2843 10.6151
R8731 gnd.n2847 gnd.n2844 10.6151
R8732 gnd.n2848 gnd.n2847 10.6151
R8733 gnd.n2851 gnd.n2848 10.6151
R8734 gnd.n2852 gnd.n2851 10.6151
R8735 gnd.n2855 gnd.n2852 10.6151
R8736 gnd.n2856 gnd.n2855 10.6151
R8737 gnd.n2859 gnd.n2856 10.6151
R8738 gnd.n2860 gnd.n2859 10.6151
R8739 gnd.n2863 gnd.n2860 10.6151
R8740 gnd.n2864 gnd.n2863 10.6151
R8741 gnd.n2867 gnd.n2864 10.6151
R8742 gnd.n2868 gnd.n2867 10.6151
R8743 gnd.n2871 gnd.n2868 10.6151
R8744 gnd.n2872 gnd.n2871 10.6151
R8745 gnd.n3846 gnd.n3845 10.6151
R8746 gnd.n3845 gnd.n3844 10.6151
R8747 gnd.n3844 gnd.n3843 10.6151
R8748 gnd.n3843 gnd.n3841 10.6151
R8749 gnd.n3841 gnd.n3838 10.6151
R8750 gnd.n3838 gnd.n3837 10.6151
R8751 gnd.n3837 gnd.n3834 10.6151
R8752 gnd.n3834 gnd.n3833 10.6151
R8753 gnd.n3833 gnd.n3830 10.6151
R8754 gnd.n3830 gnd.n3829 10.6151
R8755 gnd.n3829 gnd.n3826 10.6151
R8756 gnd.n3826 gnd.n3825 10.6151
R8757 gnd.n3825 gnd.n3822 10.6151
R8758 gnd.n3822 gnd.n3821 10.6151
R8759 gnd.n3821 gnd.n3818 10.6151
R8760 gnd.n3818 gnd.n3817 10.6151
R8761 gnd.n3817 gnd.n3814 10.6151
R8762 gnd.n3814 gnd.n3813 10.6151
R8763 gnd.n3813 gnd.n3810 10.6151
R8764 gnd.n3810 gnd.n3809 10.6151
R8765 gnd.n3809 gnd.n3806 10.6151
R8766 gnd.n3806 gnd.n3805 10.6151
R8767 gnd.n3805 gnd.n3802 10.6151
R8768 gnd.n3802 gnd.n3801 10.6151
R8769 gnd.n3801 gnd.n3798 10.6151
R8770 gnd.n3798 gnd.n3797 10.6151
R8771 gnd.n3797 gnd.n3794 10.6151
R8772 gnd.n3794 gnd.n3793 10.6151
R8773 gnd.n3790 gnd.n3789 10.6151
R8774 gnd.n3789 gnd.n1410 10.6151
R8775 gnd.n3539 gnd.n3538 10.6151
R8776 gnd.n3538 gnd.n1669 10.6151
R8777 gnd.n3533 gnd.n1669 10.6151
R8778 gnd.n3533 gnd.n3532 10.6151
R8779 gnd.n3532 gnd.n3531 10.6151
R8780 gnd.n3531 gnd.n1674 10.6151
R8781 gnd.n3526 gnd.n1674 10.6151
R8782 gnd.n3526 gnd.n3525 10.6151
R8783 gnd.n3525 gnd.n3524 10.6151
R8784 gnd.n3524 gnd.n1677 10.6151
R8785 gnd.n3519 gnd.n1677 10.6151
R8786 gnd.n3519 gnd.n3518 10.6151
R8787 gnd.n3518 gnd.n3517 10.6151
R8788 gnd.n3517 gnd.n1680 10.6151
R8789 gnd.n3512 gnd.n1680 10.6151
R8790 gnd.n3512 gnd.n3511 10.6151
R8791 gnd.n3511 gnd.n3510 10.6151
R8792 gnd.n3510 gnd.n1683 10.6151
R8793 gnd.n3505 gnd.n1683 10.6151
R8794 gnd.n3505 gnd.n3504 10.6151
R8795 gnd.n3504 gnd.n3503 10.6151
R8796 gnd.n3503 gnd.n1686 10.6151
R8797 gnd.n3498 gnd.n1686 10.6151
R8798 gnd.n3498 gnd.n3497 10.6151
R8799 gnd.n3497 gnd.n3496 10.6151
R8800 gnd.n3496 gnd.n1689 10.6151
R8801 gnd.n3491 gnd.n1689 10.6151
R8802 gnd.n3491 gnd.n3490 10.6151
R8803 gnd.n3488 gnd.n1694 10.6151
R8804 gnd.n3483 gnd.n1694 10.6151
R8805 gnd.n3782 gnd.n3781 10.6151
R8806 gnd.n3781 gnd.n1469 10.6151
R8807 gnd.n2920 gnd.n1469 10.6151
R8808 gnd.n2921 gnd.n2920 10.6151
R8809 gnd.n2922 gnd.n2921 10.6151
R8810 gnd.n2922 gnd.n1980 10.6151
R8811 gnd.n2938 gnd.n1980 10.6151
R8812 gnd.n2939 gnd.n2938 10.6151
R8813 gnd.n2940 gnd.n2939 10.6151
R8814 gnd.n2940 gnd.n1967 10.6151
R8815 gnd.n2955 gnd.n1967 10.6151
R8816 gnd.n2956 gnd.n2955 10.6151
R8817 gnd.n2963 gnd.n2956 10.6151
R8818 gnd.n2963 gnd.n2962 10.6151
R8819 gnd.n2962 gnd.n2961 10.6151
R8820 gnd.n2961 gnd.n2960 10.6151
R8821 gnd.n2960 gnd.n1943 10.6151
R8822 gnd.n3008 gnd.n1943 10.6151
R8823 gnd.n3008 gnd.n3007 10.6151
R8824 gnd.n3007 gnd.n3006 10.6151
R8825 gnd.n3006 gnd.n1926 10.6151
R8826 gnd.n3059 gnd.n1926 10.6151
R8827 gnd.n3060 gnd.n3059 10.6151
R8828 gnd.n3064 gnd.n3060 10.6151
R8829 gnd.n3064 gnd.n3063 10.6151
R8830 gnd.n3063 gnd.n3062 10.6151
R8831 gnd.n3062 gnd.n1903 10.6151
R8832 gnd.n3090 gnd.n1903 10.6151
R8833 gnd.n3091 gnd.n3090 10.6151
R8834 gnd.n3092 gnd.n3091 10.6151
R8835 gnd.n3092 gnd.n1888 10.6151
R8836 gnd.n3108 gnd.n1888 10.6151
R8837 gnd.n3109 gnd.n3108 10.6151
R8838 gnd.n3110 gnd.n3109 10.6151
R8839 gnd.n3110 gnd.n1874 10.6151
R8840 gnd.n3128 gnd.n1874 10.6151
R8841 gnd.n3129 gnd.n3128 10.6151
R8842 gnd.n3135 gnd.n3129 10.6151
R8843 gnd.n3135 gnd.n3134 10.6151
R8844 gnd.n3134 gnd.n3133 10.6151
R8845 gnd.n3133 gnd.n3132 10.6151
R8846 gnd.n3132 gnd.n1846 10.6151
R8847 gnd.n3178 gnd.n1846 10.6151
R8848 gnd.n3178 gnd.n3177 10.6151
R8849 gnd.n3177 gnd.n3176 10.6151
R8850 gnd.n3176 gnd.n1832 10.6151
R8851 gnd.n3232 gnd.n1832 10.6151
R8852 gnd.n3233 gnd.n3232 10.6151
R8853 gnd.n3237 gnd.n3233 10.6151
R8854 gnd.n3237 gnd.n3236 10.6151
R8855 gnd.n3236 gnd.n3235 10.6151
R8856 gnd.n3235 gnd.n1808 10.6151
R8857 gnd.n3262 gnd.n1808 10.6151
R8858 gnd.n3263 gnd.n3262 10.6151
R8859 gnd.n3264 gnd.n3263 10.6151
R8860 gnd.n3264 gnd.n1796 10.6151
R8861 gnd.n3280 gnd.n1796 10.6151
R8862 gnd.n3281 gnd.n3280 10.6151
R8863 gnd.n3282 gnd.n3281 10.6151
R8864 gnd.n3282 gnd.n1782 10.6151
R8865 gnd.n3303 gnd.n1782 10.6151
R8866 gnd.n3304 gnd.n3303 10.6151
R8867 gnd.n3310 gnd.n3304 10.6151
R8868 gnd.n3310 gnd.n3309 10.6151
R8869 gnd.n3309 gnd.n3308 10.6151
R8870 gnd.n3308 gnd.n3307 10.6151
R8871 gnd.n3307 gnd.n1757 10.6151
R8872 gnd.n3352 gnd.n1757 10.6151
R8873 gnd.n3352 gnd.n3351 10.6151
R8874 gnd.n3351 gnd.n3350 10.6151
R8875 gnd.n3350 gnd.n1742 10.6151
R8876 gnd.n3383 gnd.n1742 10.6151
R8877 gnd.n3384 gnd.n3383 10.6151
R8878 gnd.n3394 gnd.n3384 10.6151
R8879 gnd.n3394 gnd.n3393 10.6151
R8880 gnd.n3393 gnd.n3392 10.6151
R8881 gnd.n3392 gnd.n3385 10.6151
R8882 gnd.n3386 gnd.n3385 10.6151
R8883 gnd.n3386 gnd.n1649 10.6151
R8884 gnd.n3541 gnd.n1649 10.6151
R8885 gnd.n4824 gnd.t157 10.5161
R8886 gnd.n4269 gnd.t38 10.5161
R8887 gnd.n5190 gnd.t65 10.5161
R8888 gnd.n1231 gnd.t16 10.5161
R8889 gnd.t32 gnd.n1234 10.5161
R8890 gnd.n3849 gnd.n1445 10.5161
R8891 gnd.n1672 gnd.n1671 10.5161
R8892 gnd.n6672 gnd.t0 10.5161
R8893 gnd.n6680 gnd.t7 10.5161
R8894 gnd.n5466 gnd.n5450 10.4732
R8895 gnd.n5434 gnd.n5418 10.4732
R8896 gnd.n5402 gnd.n5386 10.4732
R8897 gnd.n5371 gnd.n5355 10.4732
R8898 gnd.n5339 gnd.n5323 10.4732
R8899 gnd.n5307 gnd.n5291 10.4732
R8900 gnd.n5275 gnd.n5259 10.4732
R8901 gnd.n5244 gnd.n5228 10.4732
R8902 gnd.n1964 gnd.n1954 10.1975
R8903 gnd.t13 gnd.n3055 10.1975
R8904 gnd.n1872 gnd.n1870 10.1975
R8905 gnd.n3130 gnd.n1855 10.1975
R8906 gnd.n3278 gnd.t96 10.1975
R8907 gnd.n3305 gnd.n1765 10.1975
R8908 gnd.t187 gnd.n4286 9.87883
R8909 gnd.n1193 gnd.t46 9.87883
R8910 gnd.t42 gnd.n1272 9.87883
R8911 gnd.t20 gnd.n209 9.87883
R8912 gnd.t106 gnd.n107 9.87883
R8913 gnd.n5470 gnd.n5469 9.69747
R8914 gnd.n5438 gnd.n5437 9.69747
R8915 gnd.n5406 gnd.n5405 9.69747
R8916 gnd.n5375 gnd.n5374 9.69747
R8917 gnd.n5343 gnd.n5342 9.69747
R8918 gnd.n5311 gnd.n5310 9.69747
R8919 gnd.n5279 gnd.n5278 9.69747
R8920 gnd.n5248 gnd.n5247 9.69747
R8921 gnd.n2924 gnd.n1991 9.56018
R8922 gnd.n2995 gnd.t97 9.56018
R8923 gnd.n3094 gnd.n1901 9.56018
R8924 gnd.n3222 gnd.n1829 9.56018
R8925 gnd.t6 gnd.n3313 9.56018
R8926 gnd.n3373 gnd.t314 9.56018
R8927 gnd.n3417 gnd.t209 9.56018
R8928 gnd.n3543 gnd.n1646 9.56018
R8929 gnd.n5476 gnd.n5475 9.45567
R8930 gnd.n5444 gnd.n5443 9.45567
R8931 gnd.n5412 gnd.n5411 9.45567
R8932 gnd.n5381 gnd.n5380 9.45567
R8933 gnd.n5349 gnd.n5348 9.45567
R8934 gnd.n5317 gnd.n5316 9.45567
R8935 gnd.n5285 gnd.n5284 9.45567
R8936 gnd.n5254 gnd.n5253 9.45567
R8937 gnd.n6962 gnd.n6902 9.30959
R8938 gnd.n6461 gnd.n6460 9.30959
R8939 gnd.n4081 gnd.n4080 9.30959
R8940 gnd.n2244 gnd.n2214 9.30959
R8941 gnd.n6421 gnd.n6420 9.3005
R8942 gnd.n6424 gnd.n384 9.3005
R8943 gnd.n6425 gnd.n383 9.3005
R8944 gnd.n6428 gnd.n382 9.3005
R8945 gnd.n6429 gnd.n381 9.3005
R8946 gnd.n6432 gnd.n380 9.3005
R8947 gnd.n6433 gnd.n379 9.3005
R8948 gnd.n6436 gnd.n378 9.3005
R8949 gnd.n6437 gnd.n377 9.3005
R8950 gnd.n6440 gnd.n376 9.3005
R8951 gnd.n6441 gnd.n375 9.3005
R8952 gnd.n6444 gnd.n374 9.3005
R8953 gnd.n6445 gnd.n373 9.3005
R8954 gnd.n6448 gnd.n372 9.3005
R8955 gnd.n6449 gnd.n371 9.3005
R8956 gnd.n6452 gnd.n370 9.3005
R8957 gnd.n6453 gnd.n369 9.3005
R8958 gnd.n6456 gnd.n368 9.3005
R8959 gnd.n6457 gnd.n367 9.3005
R8960 gnd.n6460 gnd.n366 9.3005
R8961 gnd.n6464 gnd.n362 9.3005
R8962 gnd.n6465 gnd.n361 9.3005
R8963 gnd.n6468 gnd.n360 9.3005
R8964 gnd.n6469 gnd.n359 9.3005
R8965 gnd.n6472 gnd.n358 9.3005
R8966 gnd.n6473 gnd.n357 9.3005
R8967 gnd.n6476 gnd.n356 9.3005
R8968 gnd.n6477 gnd.n355 9.3005
R8969 gnd.n6480 gnd.n354 9.3005
R8970 gnd.n6482 gnd.n350 9.3005
R8971 gnd.n6485 gnd.n349 9.3005
R8972 gnd.n6486 gnd.n348 9.3005
R8973 gnd.n6489 gnd.n347 9.3005
R8974 gnd.n6490 gnd.n346 9.3005
R8975 gnd.n6493 gnd.n345 9.3005
R8976 gnd.n6494 gnd.n344 9.3005
R8977 gnd.n6497 gnd.n343 9.3005
R8978 gnd.n6499 gnd.n340 9.3005
R8979 gnd.n6502 gnd.n339 9.3005
R8980 gnd.n6503 gnd.n338 9.3005
R8981 gnd.n6506 gnd.n337 9.3005
R8982 gnd.n6507 gnd.n336 9.3005
R8983 gnd.n6510 gnd.n335 9.3005
R8984 gnd.n6511 gnd.n334 9.3005
R8985 gnd.n6514 gnd.n333 9.3005
R8986 gnd.n6515 gnd.n332 9.3005
R8987 gnd.n6518 gnd.n331 9.3005
R8988 gnd.n6519 gnd.n330 9.3005
R8989 gnd.n6522 gnd.n329 9.3005
R8990 gnd.n6523 gnd.n328 9.3005
R8991 gnd.n6526 gnd.n327 9.3005
R8992 gnd.n6527 gnd.n326 9.3005
R8993 gnd.n6528 gnd.n325 9.3005
R8994 gnd.n282 gnd.n281 9.3005
R8995 gnd.n6534 gnd.n6533 9.3005
R8996 gnd.n6461 gnd.n363 9.3005
R8997 gnd.n6419 gnd.n385 9.3005
R8998 gnd.n6538 gnd.n6537 9.3005
R8999 gnd.n6536 gnd.n280 9.3005
R9000 gnd.n253 gnd.n252 9.3005
R9001 gnd.n6568 gnd.n6567 9.3005
R9002 gnd.n6569 gnd.n251 9.3005
R9003 gnd.n6573 gnd.n6570 9.3005
R9004 gnd.n6572 gnd.n6571 9.3005
R9005 gnd.n227 gnd.n226 9.3005
R9006 gnd.n6608 gnd.n6607 9.3005
R9007 gnd.n6609 gnd.n225 9.3005
R9008 gnd.n6611 gnd.n6610 9.3005
R9009 gnd.n207 gnd.n206 9.3005
R9010 gnd.n6632 gnd.n6631 9.3005
R9011 gnd.n6633 gnd.n205 9.3005
R9012 gnd.n6637 gnd.n6634 9.3005
R9013 gnd.n6636 gnd.n6635 9.3005
R9014 gnd.n6535 gnd.n279 9.3005
R9015 gnd.n184 gnd.n183 9.3005
R9016 gnd.n6664 gnd.n6663 9.3005
R9017 gnd.n6665 gnd.n182 9.3005
R9018 gnd.n6670 gnd.n6666 9.3005
R9019 gnd.n6669 gnd.n6668 9.3005
R9020 gnd.n6667 gnd.n78 9.3005
R9021 gnd.n7105 gnd.n79 9.3005
R9022 gnd.n7104 gnd.n80 9.3005
R9023 gnd.n7103 gnd.n81 9.3005
R9024 gnd.n98 gnd.n82 9.3005
R9025 gnd.n7093 gnd.n99 9.3005
R9026 gnd.n7092 gnd.n100 9.3005
R9027 gnd.n7091 gnd.n101 9.3005
R9028 gnd.n118 gnd.n102 9.3005
R9029 gnd.n7081 gnd.n119 9.3005
R9030 gnd.n7080 gnd.n120 9.3005
R9031 gnd.n7079 gnd.n121 9.3005
R9032 gnd.n136 gnd.n122 9.3005
R9033 gnd.n7069 gnd.n137 9.3005
R9034 gnd.n7068 gnd.n138 9.3005
R9035 gnd.n7067 gnd.n139 9.3005
R9036 gnd.n156 gnd.n140 9.3005
R9037 gnd.n7057 gnd.n157 9.3005
R9038 gnd.n7056 gnd.n158 9.3005
R9039 gnd.n7055 gnd.n159 9.3005
R9040 gnd.n6866 gnd.n160 9.3005
R9041 gnd.n7111 gnd.n7110 9.3005
R9042 gnd.n7109 gnd.n69 9.3005
R9043 gnd.n6796 gnd.n71 9.3005
R9044 gnd.n6798 gnd.n6797 9.3005
R9045 gnd.n6801 gnd.n6800 9.3005
R9046 gnd.n6802 gnd.n6795 9.3005
R9047 gnd.n6805 gnd.n6803 9.3005
R9048 gnd.n6806 gnd.n6794 9.3005
R9049 gnd.n6809 gnd.n6808 9.3005
R9050 gnd.n6810 gnd.n6793 9.3005
R9051 gnd.n6813 gnd.n6811 9.3005
R9052 gnd.n6814 gnd.n6792 9.3005
R9053 gnd.n6817 gnd.n6816 9.3005
R9054 gnd.n6818 gnd.n6791 9.3005
R9055 gnd.n6821 gnd.n6819 9.3005
R9056 gnd.n6822 gnd.n6790 9.3005
R9057 gnd.n6825 gnd.n6824 9.3005
R9058 gnd.n6826 gnd.n6789 9.3005
R9059 gnd.n6829 gnd.n6827 9.3005
R9060 gnd.n6830 gnd.n6788 9.3005
R9061 gnd.n6832 gnd.n6831 9.3005
R9062 gnd.n6748 gnd.n6747 9.3005
R9063 gnd.n6750 gnd.n6749 9.3005
R9064 gnd.n6753 gnd.n6744 9.3005
R9065 gnd.n6757 gnd.n6756 9.3005
R9066 gnd.n6758 gnd.n6743 9.3005
R9067 gnd.n6760 gnd.n6759 9.3005
R9068 gnd.n6763 gnd.n6742 9.3005
R9069 gnd.n6767 gnd.n6766 9.3005
R9070 gnd.n6768 gnd.n6741 9.3005
R9071 gnd.n6770 gnd.n6769 9.3005
R9072 gnd.n6773 gnd.n6740 9.3005
R9073 gnd.n6777 gnd.n6776 9.3005
R9074 gnd.n6778 gnd.n6739 9.3005
R9075 gnd.n6780 gnd.n6779 9.3005
R9076 gnd.n6783 gnd.n6738 9.3005
R9077 gnd.n6786 gnd.n6785 9.3005
R9078 gnd.n6787 gnd.n6737 9.3005
R9079 gnd.n6834 gnd.n6833 9.3005
R9080 gnd.n6745 gnd.n6718 9.3005
R9081 gnd.n7039 gnd.n7038 9.3005
R9082 gnd.n7037 gnd.n6868 9.3005
R9083 gnd.n7036 gnd.n7035 9.3005
R9084 gnd.n7032 gnd.n6869 9.3005
R9085 gnd.n7029 gnd.n6870 9.3005
R9086 gnd.n7028 gnd.n6871 9.3005
R9087 gnd.n7025 gnd.n6872 9.3005
R9088 gnd.n7024 gnd.n6873 9.3005
R9089 gnd.n7021 gnd.n6874 9.3005
R9090 gnd.n7020 gnd.n6875 9.3005
R9091 gnd.n7017 gnd.n6876 9.3005
R9092 gnd.n7016 gnd.n6877 9.3005
R9093 gnd.n7013 gnd.n6878 9.3005
R9094 gnd.n7012 gnd.n6879 9.3005
R9095 gnd.n7009 gnd.n6880 9.3005
R9096 gnd.n7008 gnd.n6881 9.3005
R9097 gnd.n7005 gnd.n6882 9.3005
R9098 gnd.n7001 gnd.n6883 9.3005
R9099 gnd.n6998 gnd.n6884 9.3005
R9100 gnd.n6997 gnd.n6885 9.3005
R9101 gnd.n6994 gnd.n6886 9.3005
R9102 gnd.n6993 gnd.n6887 9.3005
R9103 gnd.n6990 gnd.n6888 9.3005
R9104 gnd.n6989 gnd.n6889 9.3005
R9105 gnd.n6986 gnd.n6890 9.3005
R9106 gnd.n6985 gnd.n6891 9.3005
R9107 gnd.n6982 gnd.n6892 9.3005
R9108 gnd.n6981 gnd.n6893 9.3005
R9109 gnd.n6978 gnd.n6894 9.3005
R9110 gnd.n6977 gnd.n6895 9.3005
R9111 gnd.n6974 gnd.n6896 9.3005
R9112 gnd.n6973 gnd.n6897 9.3005
R9113 gnd.n6970 gnd.n6898 9.3005
R9114 gnd.n6969 gnd.n6899 9.3005
R9115 gnd.n6966 gnd.n6900 9.3005
R9116 gnd.n6965 gnd.n6901 9.3005
R9117 gnd.n6962 gnd.n6961 9.3005
R9118 gnd.n6960 gnd.n6902 9.3005
R9119 gnd.n6959 gnd.n6958 9.3005
R9120 gnd.n6955 gnd.n6905 9.3005
R9121 gnd.n6952 gnd.n6906 9.3005
R9122 gnd.n6951 gnd.n6907 9.3005
R9123 gnd.n6948 gnd.n6908 9.3005
R9124 gnd.n6947 gnd.n6909 9.3005
R9125 gnd.n6944 gnd.n6910 9.3005
R9126 gnd.n6943 gnd.n6911 9.3005
R9127 gnd.n6940 gnd.n6912 9.3005
R9128 gnd.n6939 gnd.n6913 9.3005
R9129 gnd.n6936 gnd.n6914 9.3005
R9130 gnd.n6935 gnd.n6915 9.3005
R9131 gnd.n6932 gnd.n6916 9.3005
R9132 gnd.n6931 gnd.n6917 9.3005
R9133 gnd.n6928 gnd.n6918 9.3005
R9134 gnd.n6927 gnd.n6919 9.3005
R9135 gnd.n6924 gnd.n6920 9.3005
R9136 gnd.n6923 gnd.n6921 9.3005
R9137 gnd.n6722 gnd.n6719 9.3005
R9138 gnd.n7047 gnd.n7046 9.3005
R9139 gnd.n7040 gnd.n6867 9.3005
R9140 gnd.n505 gnd.n504 9.3005
R9141 gnd.n506 gnd.n264 9.3005
R9142 gnd.n6551 gnd.n265 9.3005
R9143 gnd.n6552 gnd.n262 9.3005
R9144 gnd.n6555 gnd.n263 9.3005
R9145 gnd.n6557 gnd.n6556 9.3005
R9146 gnd.n6558 gnd.n236 9.3005
R9147 gnd.n6596 gnd.n237 9.3005
R9148 gnd.n6597 gnd.n235 9.3005
R9149 gnd.n6599 gnd.n6598 9.3005
R9150 gnd.n6600 gnd.n218 9.3005
R9151 gnd.n6616 gnd.n219 9.3005
R9152 gnd.n6617 gnd.n216 9.3005
R9153 gnd.n6619 gnd.n217 9.3005
R9154 gnd.n6621 gnd.n6620 9.3005
R9155 gnd.n6622 gnd.n192 9.3005
R9156 gnd.n6654 gnd.n191 9.3005
R9157 gnd.n6658 gnd.n6657 9.3005
R9158 gnd.n6656 gnd.n174 9.3005
R9159 gnd.n6675 gnd.n173 9.3005
R9160 gnd.n6677 gnd.n6676 9.3005
R9161 gnd.n6678 gnd.n168 9.3005
R9162 gnd.n6684 gnd.n167 9.3005
R9163 gnd.n6687 gnd.n6685 9.3005
R9164 gnd.n6688 gnd.n90 9.3005
R9165 gnd.n6690 gnd.n91 9.3005
R9166 gnd.n6691 gnd.n92 9.3005
R9167 gnd.n6694 gnd.n6692 9.3005
R9168 gnd.n6695 gnd.n109 9.3005
R9169 gnd.n6697 gnd.n110 9.3005
R9170 gnd.n6698 gnd.n111 9.3005
R9171 gnd.n6701 gnd.n6699 9.3005
R9172 gnd.n6702 gnd.n128 9.3005
R9173 gnd.n6704 gnd.n129 9.3005
R9174 gnd.n6705 gnd.n130 9.3005
R9175 gnd.n6708 gnd.n6706 9.3005
R9176 gnd.n6709 gnd.n147 9.3005
R9177 gnd.n6711 gnd.n148 9.3005
R9178 gnd.n6712 gnd.n149 9.3005
R9179 gnd.n6715 gnd.n6713 9.3005
R9180 gnd.n6716 gnd.n166 9.3005
R9181 gnd.n7049 gnd.n6717 9.3005
R9182 gnd.n503 gnd.n388 9.3005
R9183 gnd.n6326 gnd.n505 9.3005
R9184 gnd.n6325 gnd.n506 9.3005
R9185 gnd.n265 gnd.n261 9.3005
R9186 gnd.n6563 gnd.n262 9.3005
R9187 gnd.n6562 gnd.n263 9.3005
R9188 gnd.n6561 gnd.n6557 9.3005
R9189 gnd.n6560 gnd.n6558 9.3005
R9190 gnd.n237 gnd.n234 9.3005
R9191 gnd.n6603 gnd.n235 9.3005
R9192 gnd.n6602 gnd.n6599 9.3005
R9193 gnd.n6601 gnd.n6600 9.3005
R9194 gnd.n219 gnd.n215 9.3005
R9195 gnd.n6627 gnd.n216 9.3005
R9196 gnd.n6626 gnd.n217 9.3005
R9197 gnd.n6625 gnd.n6621 9.3005
R9198 gnd.n6624 gnd.n6622 9.3005
R9199 gnd.n191 gnd.n190 9.3005
R9200 gnd.n6659 gnd.n6658 9.3005
R9201 gnd.n175 gnd.n174 9.3005
R9202 gnd.n6675 gnd.n6674 9.3005
R9203 gnd.n6676 gnd.n169 9.3005
R9204 gnd.n6682 gnd.n168 9.3005
R9205 gnd.n6684 gnd.n6683 9.3005
R9206 gnd.n6685 gnd.n89 9.3005
R9207 gnd.n7099 gnd.n90 9.3005
R9208 gnd.n7098 gnd.n91 9.3005
R9209 gnd.n7097 gnd.n92 9.3005
R9210 gnd.n6692 gnd.n93 9.3005
R9211 gnd.n7087 gnd.n109 9.3005
R9212 gnd.n7086 gnd.n110 9.3005
R9213 gnd.n7085 gnd.n111 9.3005
R9214 gnd.n6699 gnd.n112 9.3005
R9215 gnd.n7075 gnd.n128 9.3005
R9216 gnd.n7074 gnd.n129 9.3005
R9217 gnd.n7073 gnd.n130 9.3005
R9218 gnd.n6706 gnd.n131 9.3005
R9219 gnd.n7063 gnd.n147 9.3005
R9220 gnd.n7062 gnd.n148 9.3005
R9221 gnd.n7061 gnd.n149 9.3005
R9222 gnd.n6713 gnd.n150 9.3005
R9223 gnd.n7051 gnd.n166 9.3005
R9224 gnd.n7050 gnd.n7049 9.3005
R9225 gnd.n6327 gnd.n388 9.3005
R9226 gnd.n5475 gnd.n5474 9.3005
R9227 gnd.n5448 gnd.n5447 9.3005
R9228 gnd.n5469 gnd.n5468 9.3005
R9229 gnd.n5467 gnd.n5466 9.3005
R9230 gnd.n5452 gnd.n5451 9.3005
R9231 gnd.n5461 gnd.n5460 9.3005
R9232 gnd.n5459 gnd.n5458 9.3005
R9233 gnd.n5443 gnd.n5442 9.3005
R9234 gnd.n5416 gnd.n5415 9.3005
R9235 gnd.n5437 gnd.n5436 9.3005
R9236 gnd.n5435 gnd.n5434 9.3005
R9237 gnd.n5420 gnd.n5419 9.3005
R9238 gnd.n5429 gnd.n5428 9.3005
R9239 gnd.n5427 gnd.n5426 9.3005
R9240 gnd.n5411 gnd.n5410 9.3005
R9241 gnd.n5384 gnd.n5383 9.3005
R9242 gnd.n5405 gnd.n5404 9.3005
R9243 gnd.n5403 gnd.n5402 9.3005
R9244 gnd.n5388 gnd.n5387 9.3005
R9245 gnd.n5397 gnd.n5396 9.3005
R9246 gnd.n5395 gnd.n5394 9.3005
R9247 gnd.n5380 gnd.n5379 9.3005
R9248 gnd.n5353 gnd.n5352 9.3005
R9249 gnd.n5374 gnd.n5373 9.3005
R9250 gnd.n5372 gnd.n5371 9.3005
R9251 gnd.n5357 gnd.n5356 9.3005
R9252 gnd.n5366 gnd.n5365 9.3005
R9253 gnd.n5364 gnd.n5363 9.3005
R9254 gnd.n5348 gnd.n5347 9.3005
R9255 gnd.n5321 gnd.n5320 9.3005
R9256 gnd.n5342 gnd.n5341 9.3005
R9257 gnd.n5340 gnd.n5339 9.3005
R9258 gnd.n5325 gnd.n5324 9.3005
R9259 gnd.n5334 gnd.n5333 9.3005
R9260 gnd.n5332 gnd.n5331 9.3005
R9261 gnd.n5316 gnd.n5315 9.3005
R9262 gnd.n5289 gnd.n5288 9.3005
R9263 gnd.n5310 gnd.n5309 9.3005
R9264 gnd.n5308 gnd.n5307 9.3005
R9265 gnd.n5293 gnd.n5292 9.3005
R9266 gnd.n5302 gnd.n5301 9.3005
R9267 gnd.n5300 gnd.n5299 9.3005
R9268 gnd.n5284 gnd.n5283 9.3005
R9269 gnd.n5257 gnd.n5256 9.3005
R9270 gnd.n5278 gnd.n5277 9.3005
R9271 gnd.n5276 gnd.n5275 9.3005
R9272 gnd.n5261 gnd.n5260 9.3005
R9273 gnd.n5270 gnd.n5269 9.3005
R9274 gnd.n5268 gnd.n5267 9.3005
R9275 gnd.n5253 gnd.n5252 9.3005
R9276 gnd.n5226 gnd.n5225 9.3005
R9277 gnd.n5247 gnd.n5246 9.3005
R9278 gnd.n5245 gnd.n5244 9.3005
R9279 gnd.n5230 gnd.n5229 9.3005
R9280 gnd.n5239 gnd.n5238 9.3005
R9281 gnd.n5237 gnd.n5236 9.3005
R9282 gnd.n5601 gnd.n5600 9.3005
R9283 gnd.n5599 gnd.n4169 9.3005
R9284 gnd.n5598 gnd.n5597 9.3005
R9285 gnd.n5594 gnd.n4170 9.3005
R9286 gnd.n5591 gnd.n4171 9.3005
R9287 gnd.n5590 gnd.n4172 9.3005
R9288 gnd.n5587 gnd.n4173 9.3005
R9289 gnd.n5586 gnd.n4174 9.3005
R9290 gnd.n5583 gnd.n4175 9.3005
R9291 gnd.n5582 gnd.n4176 9.3005
R9292 gnd.n5579 gnd.n4177 9.3005
R9293 gnd.n5578 gnd.n4178 9.3005
R9294 gnd.n5575 gnd.n4179 9.3005
R9295 gnd.n5574 gnd.n4180 9.3005
R9296 gnd.n5571 gnd.n5570 9.3005
R9297 gnd.n5569 gnd.n4181 9.3005
R9298 gnd.n5602 gnd.n4168 9.3005
R9299 gnd.n4843 gnd.n4842 9.3005
R9300 gnd.n4547 gnd.n4546 9.3005
R9301 gnd.n4870 gnd.n4869 9.3005
R9302 gnd.n4871 gnd.n4545 9.3005
R9303 gnd.n4875 gnd.n4872 9.3005
R9304 gnd.n4874 gnd.n4873 9.3005
R9305 gnd.n4519 gnd.n4518 9.3005
R9306 gnd.n4900 gnd.n4899 9.3005
R9307 gnd.n4901 gnd.n4517 9.3005
R9308 gnd.n4903 gnd.n4902 9.3005
R9309 gnd.n4497 gnd.n4496 9.3005
R9310 gnd.n4931 gnd.n4930 9.3005
R9311 gnd.n4932 gnd.n4495 9.3005
R9312 gnd.n4940 gnd.n4933 9.3005
R9313 gnd.n4939 gnd.n4934 9.3005
R9314 gnd.n4938 gnd.n4936 9.3005
R9315 gnd.n4935 gnd.n4444 9.3005
R9316 gnd.n4988 gnd.n4445 9.3005
R9317 gnd.n4987 gnd.n4446 9.3005
R9318 gnd.n4986 gnd.n4447 9.3005
R9319 gnd.n4466 gnd.n4448 9.3005
R9320 gnd.n4468 gnd.n4467 9.3005
R9321 gnd.n4366 gnd.n4365 9.3005
R9322 gnd.n5026 gnd.n5025 9.3005
R9323 gnd.n5027 gnd.n4364 9.3005
R9324 gnd.n5031 gnd.n5028 9.3005
R9325 gnd.n5030 gnd.n5029 9.3005
R9326 gnd.n4339 gnd.n4338 9.3005
R9327 gnd.n5066 gnd.n5065 9.3005
R9328 gnd.n5067 gnd.n4337 9.3005
R9329 gnd.n5071 gnd.n5068 9.3005
R9330 gnd.n5070 gnd.n5069 9.3005
R9331 gnd.n4312 gnd.n4311 9.3005
R9332 gnd.n5111 gnd.n5110 9.3005
R9333 gnd.n5112 gnd.n4310 9.3005
R9334 gnd.n5116 gnd.n5113 9.3005
R9335 gnd.n5115 gnd.n5114 9.3005
R9336 gnd.n4284 gnd.n4283 9.3005
R9337 gnd.n5151 gnd.n5150 9.3005
R9338 gnd.n5152 gnd.n4282 9.3005
R9339 gnd.n5156 gnd.n5153 9.3005
R9340 gnd.n5155 gnd.n5154 9.3005
R9341 gnd.n4257 gnd.n4256 9.3005
R9342 gnd.n5200 gnd.n5199 9.3005
R9343 gnd.n5201 gnd.n4255 9.3005
R9344 gnd.n5205 gnd.n5202 9.3005
R9345 gnd.n5204 gnd.n5203 9.3005
R9346 gnd.n4230 gnd.n4229 9.3005
R9347 gnd.n5494 gnd.n5493 9.3005
R9348 gnd.n5495 gnd.n4228 9.3005
R9349 gnd.n5501 gnd.n5496 9.3005
R9350 gnd.n5500 gnd.n5497 9.3005
R9351 gnd.n5499 gnd.n5498 9.3005
R9352 gnd.n4844 gnd.n4841 9.3005
R9353 gnd.n4626 gnd.n4585 9.3005
R9354 gnd.n4621 gnd.n4620 9.3005
R9355 gnd.n4619 gnd.n4586 9.3005
R9356 gnd.n4618 gnd.n4617 9.3005
R9357 gnd.n4614 gnd.n4587 9.3005
R9358 gnd.n4611 gnd.n4610 9.3005
R9359 gnd.n4609 gnd.n4588 9.3005
R9360 gnd.n4608 gnd.n4607 9.3005
R9361 gnd.n4604 gnd.n4589 9.3005
R9362 gnd.n4601 gnd.n4600 9.3005
R9363 gnd.n4599 gnd.n4590 9.3005
R9364 gnd.n4598 gnd.n4597 9.3005
R9365 gnd.n4594 gnd.n4592 9.3005
R9366 gnd.n4591 gnd.n4571 9.3005
R9367 gnd.n4838 gnd.n4570 9.3005
R9368 gnd.n4840 gnd.n4839 9.3005
R9369 gnd.n4628 gnd.n4627 9.3005
R9370 gnd.n4851 gnd.n4557 9.3005
R9371 gnd.n4858 gnd.n4558 9.3005
R9372 gnd.n4860 gnd.n4859 9.3005
R9373 gnd.n4861 gnd.n4538 9.3005
R9374 gnd.n4880 gnd.n4879 9.3005
R9375 gnd.n4882 gnd.n4530 9.3005
R9376 gnd.n4889 gnd.n4532 9.3005
R9377 gnd.n4890 gnd.n4527 9.3005
R9378 gnd.n4892 gnd.n4891 9.3005
R9379 gnd.n4528 gnd.n4513 9.3005
R9380 gnd.n4908 gnd.n4511 9.3005
R9381 gnd.n4912 gnd.n4911 9.3005
R9382 gnd.n4910 gnd.n4487 9.3005
R9383 gnd.n4947 gnd.n4486 9.3005
R9384 gnd.n4950 gnd.n4949 9.3005
R9385 gnd.n4483 gnd.n4482 9.3005
R9386 gnd.n4956 gnd.n4484 9.3005
R9387 gnd.n4958 gnd.n4957 9.3005
R9388 gnd.n4960 gnd.n4481 9.3005
R9389 gnd.n4963 gnd.n4962 9.3005
R9390 gnd.n4966 gnd.n4964 9.3005
R9391 gnd.n4968 gnd.n4967 9.3005
R9392 gnd.n4974 gnd.n4969 9.3005
R9393 gnd.n4973 gnd.n4972 9.3005
R9394 gnd.n4357 gnd.n4356 9.3005
R9395 gnd.n5040 gnd.n5039 9.3005
R9396 gnd.n5041 gnd.n4350 9.3005
R9397 gnd.n5049 gnd.n4349 9.3005
R9398 gnd.n5052 gnd.n5051 9.3005
R9399 gnd.n5054 gnd.n5053 9.3005
R9400 gnd.n5057 gnd.n4332 9.3005
R9401 gnd.n5055 gnd.n4330 9.3005
R9402 gnd.n5077 gnd.n4328 9.3005
R9403 gnd.n5079 gnd.n5078 9.3005
R9404 gnd.n4302 gnd.n4301 9.3005
R9405 gnd.n5125 gnd.n5124 9.3005
R9406 gnd.n5126 gnd.n4295 9.3005
R9407 gnd.n5134 gnd.n4294 9.3005
R9408 gnd.n5137 gnd.n5136 9.3005
R9409 gnd.n5139 gnd.n5138 9.3005
R9410 gnd.n5142 gnd.n4277 9.3005
R9411 gnd.n5140 gnd.n4275 9.3005
R9412 gnd.n5162 gnd.n4273 9.3005
R9413 gnd.n5164 gnd.n5163 9.3005
R9414 gnd.n4248 gnd.n4247 9.3005
R9415 gnd.n5214 gnd.n5213 9.3005
R9416 gnd.n5215 gnd.n4241 9.3005
R9417 gnd.n5223 gnd.n4240 9.3005
R9418 gnd.n5482 gnd.n5481 9.3005
R9419 gnd.n5484 gnd.n5483 9.3005
R9420 gnd.n5485 gnd.n4221 9.3005
R9421 gnd.n5509 gnd.n5508 9.3005
R9422 gnd.n4222 gnd.n4184 9.3005
R9423 gnd.n4849 gnd.n4848 9.3005
R9424 gnd.n5565 gnd.n4185 9.3005
R9425 gnd.n5564 gnd.n4187 9.3005
R9426 gnd.n5561 gnd.n4188 9.3005
R9427 gnd.n5560 gnd.n4189 9.3005
R9428 gnd.n5557 gnd.n4190 9.3005
R9429 gnd.n5556 gnd.n4191 9.3005
R9430 gnd.n5553 gnd.n4192 9.3005
R9431 gnd.n5552 gnd.n4193 9.3005
R9432 gnd.n5549 gnd.n4194 9.3005
R9433 gnd.n5548 gnd.n4195 9.3005
R9434 gnd.n5545 gnd.n4196 9.3005
R9435 gnd.n5544 gnd.n4197 9.3005
R9436 gnd.n5541 gnd.n4198 9.3005
R9437 gnd.n5540 gnd.n4199 9.3005
R9438 gnd.n5537 gnd.n4200 9.3005
R9439 gnd.n5536 gnd.n4201 9.3005
R9440 gnd.n5533 gnd.n4202 9.3005
R9441 gnd.n5532 gnd.n4203 9.3005
R9442 gnd.n5529 gnd.n4204 9.3005
R9443 gnd.n5528 gnd.n4205 9.3005
R9444 gnd.n5525 gnd.n4206 9.3005
R9445 gnd.n5524 gnd.n4207 9.3005
R9446 gnd.n5521 gnd.n4211 9.3005
R9447 gnd.n5520 gnd.n4212 9.3005
R9448 gnd.n5517 gnd.n4213 9.3005
R9449 gnd.n5516 gnd.n4214 9.3005
R9450 gnd.n5567 gnd.n5566 9.3005
R9451 gnd.n5018 gnd.n5002 9.3005
R9452 gnd.n5017 gnd.n5003 9.3005
R9453 gnd.n5016 gnd.n5004 9.3005
R9454 gnd.n5014 gnd.n5005 9.3005
R9455 gnd.n5013 gnd.n5006 9.3005
R9456 gnd.n5011 gnd.n5007 9.3005
R9457 gnd.n5010 gnd.n5008 9.3005
R9458 gnd.n4320 gnd.n4319 9.3005
R9459 gnd.n5087 gnd.n5086 9.3005
R9460 gnd.n5088 gnd.n4318 9.3005
R9461 gnd.n5105 gnd.n5089 9.3005
R9462 gnd.n5104 gnd.n5090 9.3005
R9463 gnd.n5103 gnd.n5091 9.3005
R9464 gnd.n5101 gnd.n5092 9.3005
R9465 gnd.n5100 gnd.n5093 9.3005
R9466 gnd.n5098 gnd.n5094 9.3005
R9467 gnd.n5097 gnd.n5095 9.3005
R9468 gnd.n4264 gnd.n4263 9.3005
R9469 gnd.n5172 gnd.n5171 9.3005
R9470 gnd.n5173 gnd.n4262 9.3005
R9471 gnd.n5194 gnd.n5174 9.3005
R9472 gnd.n5193 gnd.n5175 9.3005
R9473 gnd.n5192 gnd.n5176 9.3005
R9474 gnd.n5189 gnd.n5177 9.3005
R9475 gnd.n5188 gnd.n5178 9.3005
R9476 gnd.n5186 gnd.n5179 9.3005
R9477 gnd.n5185 gnd.n5180 9.3005
R9478 gnd.n5183 gnd.n5182 9.3005
R9479 gnd.n5181 gnd.n4216 9.3005
R9480 gnd.n4759 gnd.n4758 9.3005
R9481 gnd.n4649 gnd.n4648 9.3005
R9482 gnd.n4773 gnd.n4772 9.3005
R9483 gnd.n4774 gnd.n4647 9.3005
R9484 gnd.n4776 gnd.n4775 9.3005
R9485 gnd.n4637 gnd.n4636 9.3005
R9486 gnd.n4789 gnd.n4788 9.3005
R9487 gnd.n4790 gnd.n4635 9.3005
R9488 gnd.n4822 gnd.n4791 9.3005
R9489 gnd.n4821 gnd.n4792 9.3005
R9490 gnd.n4820 gnd.n4793 9.3005
R9491 gnd.n4819 gnd.n4794 9.3005
R9492 gnd.n4816 gnd.n4795 9.3005
R9493 gnd.n4815 gnd.n4796 9.3005
R9494 gnd.n4814 gnd.n4797 9.3005
R9495 gnd.n4812 gnd.n4798 9.3005
R9496 gnd.n4811 gnd.n4799 9.3005
R9497 gnd.n4808 gnd.n4800 9.3005
R9498 gnd.n4807 gnd.n4801 9.3005
R9499 gnd.n4806 gnd.n4802 9.3005
R9500 gnd.n4804 gnd.n4803 9.3005
R9501 gnd.n4503 gnd.n4502 9.3005
R9502 gnd.n4920 gnd.n4919 9.3005
R9503 gnd.n4921 gnd.n4501 9.3005
R9504 gnd.n4925 gnd.n4922 9.3005
R9505 gnd.n4924 gnd.n4923 9.3005
R9506 gnd.n4425 gnd.n4424 9.3005
R9507 gnd.n5000 gnd.n4999 9.3005
R9508 gnd.n4757 gnd.n4658 9.3005
R9509 gnd.n4660 gnd.n4659 9.3005
R9510 gnd.n4704 gnd.n4702 9.3005
R9511 gnd.n4705 gnd.n4701 9.3005
R9512 gnd.n4708 gnd.n4697 9.3005
R9513 gnd.n4709 gnd.n4696 9.3005
R9514 gnd.n4712 gnd.n4695 9.3005
R9515 gnd.n4713 gnd.n4694 9.3005
R9516 gnd.n4716 gnd.n4693 9.3005
R9517 gnd.n4717 gnd.n4692 9.3005
R9518 gnd.n4720 gnd.n4691 9.3005
R9519 gnd.n4721 gnd.n4690 9.3005
R9520 gnd.n4724 gnd.n4689 9.3005
R9521 gnd.n4725 gnd.n4688 9.3005
R9522 gnd.n4728 gnd.n4687 9.3005
R9523 gnd.n4729 gnd.n4686 9.3005
R9524 gnd.n4732 gnd.n4685 9.3005
R9525 gnd.n4733 gnd.n4684 9.3005
R9526 gnd.n4736 gnd.n4683 9.3005
R9527 gnd.n4737 gnd.n4682 9.3005
R9528 gnd.n4740 gnd.n4681 9.3005
R9529 gnd.n4741 gnd.n4680 9.3005
R9530 gnd.n4744 gnd.n4679 9.3005
R9531 gnd.n4746 gnd.n4678 9.3005
R9532 gnd.n4747 gnd.n4677 9.3005
R9533 gnd.n4748 gnd.n4676 9.3005
R9534 gnd.n4749 gnd.n4675 9.3005
R9535 gnd.n4756 gnd.n4755 9.3005
R9536 gnd.n4765 gnd.n4764 9.3005
R9537 gnd.n4766 gnd.n4652 9.3005
R9538 gnd.n4768 gnd.n4767 9.3005
R9539 gnd.n4643 gnd.n4642 9.3005
R9540 gnd.n4781 gnd.n4780 9.3005
R9541 gnd.n4782 gnd.n4641 9.3005
R9542 gnd.n4784 gnd.n4783 9.3005
R9543 gnd.n4630 gnd.n4629 9.3005
R9544 gnd.n4827 gnd.n4826 9.3005
R9545 gnd.n4828 gnd.n4584 9.3005
R9546 gnd.n4832 gnd.n4830 9.3005
R9547 gnd.n4831 gnd.n4563 9.3005
R9548 gnd.n4850 gnd.n4562 9.3005
R9549 gnd.n4853 gnd.n4852 9.3005
R9550 gnd.n4556 gnd.n4555 9.3005
R9551 gnd.n4864 gnd.n4862 9.3005
R9552 gnd.n4863 gnd.n4537 9.3005
R9553 gnd.n4881 gnd.n4536 9.3005
R9554 gnd.n4884 gnd.n4883 9.3005
R9555 gnd.n4531 gnd.n4526 9.3005
R9556 gnd.n4894 gnd.n4893 9.3005
R9557 gnd.n4529 gnd.n4509 9.3005
R9558 gnd.n4915 gnd.n4510 9.3005
R9559 gnd.n4914 gnd.n4913 9.3005
R9560 gnd.n4512 gnd.n4488 9.3005
R9561 gnd.n4946 gnd.n4945 9.3005
R9562 gnd.n4948 gnd.n4433 9.3005
R9563 gnd.n4995 gnd.n4434 9.3005
R9564 gnd.n4994 gnd.n4435 9.3005
R9565 gnd.n4993 gnd.n4436 9.3005
R9566 gnd.n4959 gnd.n4437 9.3005
R9567 gnd.n4961 gnd.n4455 9.3005
R9568 gnd.n4981 gnd.n4456 9.3005
R9569 gnd.n4980 gnd.n4457 9.3005
R9570 gnd.n4979 gnd.n4458 9.3005
R9571 gnd.n4970 gnd.n4459 9.3005
R9572 gnd.n4971 gnd.n4358 9.3005
R9573 gnd.n5037 gnd.n5036 9.3005
R9574 gnd.n5038 gnd.n4351 9.3005
R9575 gnd.n5048 gnd.n5047 9.3005
R9576 gnd.n5050 gnd.n4347 9.3005
R9577 gnd.n5060 gnd.n4348 9.3005
R9578 gnd.n5059 gnd.n5058 9.3005
R9579 gnd.n5056 gnd.n4326 9.3005
R9580 gnd.n5082 gnd.n4327 9.3005
R9581 gnd.n5081 gnd.n5080 9.3005
R9582 gnd.n4329 gnd.n4303 9.3005
R9583 gnd.n5122 gnd.n5121 9.3005
R9584 gnd.n5123 gnd.n4296 9.3005
R9585 gnd.n5133 gnd.n5132 9.3005
R9586 gnd.n5135 gnd.n4292 9.3005
R9587 gnd.n5145 gnd.n4293 9.3005
R9588 gnd.n5144 gnd.n5143 9.3005
R9589 gnd.n5141 gnd.n4271 9.3005
R9590 gnd.n5167 gnd.n4272 9.3005
R9591 gnd.n5166 gnd.n5165 9.3005
R9592 gnd.n4274 gnd.n4249 9.3005
R9593 gnd.n5211 gnd.n5210 9.3005
R9594 gnd.n5212 gnd.n4242 9.3005
R9595 gnd.n5222 gnd.n5221 9.3005
R9596 gnd.n5480 gnd.n4238 9.3005
R9597 gnd.n5488 gnd.n4239 9.3005
R9598 gnd.n5487 gnd.n5486 9.3005
R9599 gnd.n4220 gnd.n4219 9.3005
R9600 gnd.n5511 gnd.n5510 9.3005
R9601 gnd.n4654 gnd.n4653 9.3005
R9602 gnd.n2502 gnd.n2392 9.3005
R9603 gnd.n2462 gnd.n2402 9.3005
R9604 gnd.n2465 gnd.n2464 9.3005
R9605 gnd.n2466 gnd.n2401 9.3005
R9606 gnd.n2469 gnd.n2467 9.3005
R9607 gnd.n2470 gnd.n2400 9.3005
R9608 gnd.n2473 gnd.n2472 9.3005
R9609 gnd.n2474 gnd.n2399 9.3005
R9610 gnd.n2477 gnd.n2475 9.3005
R9611 gnd.n2478 gnd.n2398 9.3005
R9612 gnd.n2481 gnd.n2480 9.3005
R9613 gnd.n2482 gnd.n2397 9.3005
R9614 gnd.n2485 gnd.n2483 9.3005
R9615 gnd.n2486 gnd.n2396 9.3005
R9616 gnd.n2489 gnd.n2488 9.3005
R9617 gnd.n2490 gnd.n2395 9.3005
R9618 gnd.n2493 gnd.n2491 9.3005
R9619 gnd.n2494 gnd.n2394 9.3005
R9620 gnd.n2497 gnd.n2496 9.3005
R9621 gnd.n2498 gnd.n2393 9.3005
R9622 gnd.n2501 gnd.n2499 9.3005
R9623 gnd.n2461 gnd.n2459 9.3005
R9624 gnd.n3854 gnd.n1405 9.3005
R9625 gnd.n3857 gnd.n1404 9.3005
R9626 gnd.n3858 gnd.n1403 9.3005
R9627 gnd.n3861 gnd.n1402 9.3005
R9628 gnd.n3862 gnd.n1401 9.3005
R9629 gnd.n3865 gnd.n1400 9.3005
R9630 gnd.n3866 gnd.n1399 9.3005
R9631 gnd.n3869 gnd.n1398 9.3005
R9632 gnd.n3871 gnd.n1395 9.3005
R9633 gnd.n3874 gnd.n1394 9.3005
R9634 gnd.n3875 gnd.n1393 9.3005
R9635 gnd.n3878 gnd.n1392 9.3005
R9636 gnd.n3879 gnd.n1391 9.3005
R9637 gnd.n3882 gnd.n1390 9.3005
R9638 gnd.n3883 gnd.n1389 9.3005
R9639 gnd.n3886 gnd.n1388 9.3005
R9640 gnd.n3887 gnd.n1387 9.3005
R9641 gnd.n3890 gnd.n1386 9.3005
R9642 gnd.n3891 gnd.n1385 9.3005
R9643 gnd.n3894 gnd.n1384 9.3005
R9644 gnd.n3895 gnd.n1383 9.3005
R9645 gnd.n3898 gnd.n1382 9.3005
R9646 gnd.n3899 gnd.n1381 9.3005
R9647 gnd.n3900 gnd.n1380 9.3005
R9648 gnd.n1337 gnd.n1336 9.3005
R9649 gnd.n3906 gnd.n3905 9.3005
R9650 gnd.n2222 gnd.n2220 9.3005
R9651 gnd.n2224 gnd.n2223 9.3005
R9652 gnd.n2227 gnd.n2217 9.3005
R9653 gnd.n2231 gnd.n2230 9.3005
R9654 gnd.n2232 gnd.n2216 9.3005
R9655 gnd.n2234 gnd.n2233 9.3005
R9656 gnd.n2237 gnd.n2215 9.3005
R9657 gnd.n2241 gnd.n2240 9.3005
R9658 gnd.n2242 gnd.n2214 9.3005
R9659 gnd.n2244 gnd.n2243 9.3005
R9660 gnd.n2247 gnd.n2211 9.3005
R9661 gnd.n2251 gnd.n2250 9.3005
R9662 gnd.n2252 gnd.n2210 9.3005
R9663 gnd.n2254 gnd.n2253 9.3005
R9664 gnd.n2257 gnd.n2209 9.3005
R9665 gnd.n2261 gnd.n2260 9.3005
R9666 gnd.n2262 gnd.n2208 9.3005
R9667 gnd.n2264 gnd.n2263 9.3005
R9668 gnd.n2267 gnd.n2207 9.3005
R9669 gnd.n2271 gnd.n2270 9.3005
R9670 gnd.n2272 gnd.n2206 9.3005
R9671 gnd.n2274 gnd.n2273 9.3005
R9672 gnd.n2277 gnd.n2205 9.3005
R9673 gnd.n2281 gnd.n2280 9.3005
R9674 gnd.n2282 gnd.n2204 9.3005
R9675 gnd.n2284 gnd.n2283 9.3005
R9676 gnd.n2287 gnd.n2203 9.3005
R9677 gnd.n2291 gnd.n2290 9.3005
R9678 gnd.n2292 gnd.n2202 9.3005
R9679 gnd.n2294 gnd.n2293 9.3005
R9680 gnd.n2221 gnd.n1406 9.3005
R9681 gnd.n3981 gnd.n1217 9.3005
R9682 gnd.n3980 gnd.n1218 9.3005
R9683 gnd.n3979 gnd.n1219 9.3005
R9684 gnd.n1236 gnd.n1220 9.3005
R9685 gnd.n3969 gnd.n1237 9.3005
R9686 gnd.n3968 gnd.n1238 9.3005
R9687 gnd.n3967 gnd.n1239 9.3005
R9688 gnd.n1255 gnd.n1240 9.3005
R9689 gnd.n3957 gnd.n1256 9.3005
R9690 gnd.n3956 gnd.n1257 9.3005
R9691 gnd.n3955 gnd.n1258 9.3005
R9692 gnd.n1274 gnd.n1259 9.3005
R9693 gnd.n3945 gnd.n1275 9.3005
R9694 gnd.n3944 gnd.n1276 9.3005
R9695 gnd.n3943 gnd.n1277 9.3005
R9696 gnd.n1293 gnd.n1278 9.3005
R9697 gnd.n3933 gnd.n1294 9.3005
R9698 gnd.n3932 gnd.n1295 9.3005
R9699 gnd.n3931 gnd.n1296 9.3005
R9700 gnd.n1314 gnd.n1297 9.3005
R9701 gnd.n3921 gnd.n1315 9.3005
R9702 gnd.n3920 gnd.n1316 9.3005
R9703 gnd.n3919 gnd.n1317 9.3005
R9704 gnd.n1334 gnd.n1318 9.3005
R9705 gnd.n3909 gnd.n1335 9.3005
R9706 gnd.n3908 gnd.n3907 9.3005
R9707 gnd.n4031 gnd.n4030 9.3005
R9708 gnd.n4029 gnd.n1141 9.3005
R9709 gnd.n4028 gnd.n4027 9.3005
R9710 gnd.n1144 gnd.n1143 9.3005
R9711 gnd.n4017 gnd.n1161 9.3005
R9712 gnd.n4016 gnd.n1162 9.3005
R9713 gnd.n4015 gnd.n1163 9.3005
R9714 gnd.n1178 gnd.n1164 9.3005
R9715 gnd.n4005 gnd.n1179 9.3005
R9716 gnd.n4004 gnd.n1180 9.3005
R9717 gnd.n4003 gnd.n1181 9.3005
R9718 gnd.n1198 gnd.n1182 9.3005
R9719 gnd.n3993 gnd.n1199 9.3005
R9720 gnd.n3992 gnd.n1200 9.3005
R9721 gnd.n3991 gnd.n1201 9.3005
R9722 gnd.n1216 gnd.n1202 9.3005
R9723 gnd.n1142 gnd.n1140 9.3005
R9724 gnd.n4041 gnd.n4040 9.3005
R9725 gnd.n4044 gnd.n1125 9.3005
R9726 gnd.n4045 gnd.n1124 9.3005
R9727 gnd.n4048 gnd.n1123 9.3005
R9728 gnd.n4049 gnd.n1122 9.3005
R9729 gnd.n4052 gnd.n1121 9.3005
R9730 gnd.n4053 gnd.n1120 9.3005
R9731 gnd.n4056 gnd.n1119 9.3005
R9732 gnd.n4057 gnd.n1118 9.3005
R9733 gnd.n4060 gnd.n1117 9.3005
R9734 gnd.n4061 gnd.n1116 9.3005
R9735 gnd.n4064 gnd.n1115 9.3005
R9736 gnd.n4065 gnd.n1114 9.3005
R9737 gnd.n4068 gnd.n1113 9.3005
R9738 gnd.n4069 gnd.n1112 9.3005
R9739 gnd.n4072 gnd.n1111 9.3005
R9740 gnd.n4073 gnd.n1110 9.3005
R9741 gnd.n4076 gnd.n1109 9.3005
R9742 gnd.n4077 gnd.n1108 9.3005
R9743 gnd.n4080 gnd.n1107 9.3005
R9744 gnd.n4084 gnd.n1103 9.3005
R9745 gnd.n4085 gnd.n1102 9.3005
R9746 gnd.n4088 gnd.n1101 9.3005
R9747 gnd.n4089 gnd.n1100 9.3005
R9748 gnd.n4092 gnd.n1099 9.3005
R9749 gnd.n4093 gnd.n1098 9.3005
R9750 gnd.n4096 gnd.n1097 9.3005
R9751 gnd.n4097 gnd.n1096 9.3005
R9752 gnd.n4100 gnd.n1095 9.3005
R9753 gnd.n4101 gnd.n1094 9.3005
R9754 gnd.n4104 gnd.n1093 9.3005
R9755 gnd.n4105 gnd.n1092 9.3005
R9756 gnd.n4108 gnd.n1091 9.3005
R9757 gnd.n4109 gnd.n1090 9.3005
R9758 gnd.n4112 gnd.n1089 9.3005
R9759 gnd.n4113 gnd.n1088 9.3005
R9760 gnd.n4116 gnd.n1087 9.3005
R9761 gnd.n4117 gnd.n1086 9.3005
R9762 gnd.n4120 gnd.n1085 9.3005
R9763 gnd.n4122 gnd.n1082 9.3005
R9764 gnd.n4125 gnd.n1081 9.3005
R9765 gnd.n4126 gnd.n1080 9.3005
R9766 gnd.n4129 gnd.n1079 9.3005
R9767 gnd.n4130 gnd.n1078 9.3005
R9768 gnd.n4133 gnd.n1077 9.3005
R9769 gnd.n4134 gnd.n1076 9.3005
R9770 gnd.n4137 gnd.n1075 9.3005
R9771 gnd.n4138 gnd.n1074 9.3005
R9772 gnd.n4141 gnd.n1073 9.3005
R9773 gnd.n4142 gnd.n1072 9.3005
R9774 gnd.n4145 gnd.n1071 9.3005
R9775 gnd.n4146 gnd.n1070 9.3005
R9776 gnd.n4149 gnd.n1069 9.3005
R9777 gnd.n4151 gnd.n1068 9.3005
R9778 gnd.n4152 gnd.n1067 9.3005
R9779 gnd.n4153 gnd.n1066 9.3005
R9780 gnd.n4154 gnd.n1065 9.3005
R9781 gnd.n4081 gnd.n1104 9.3005
R9782 gnd.n4039 gnd.n1126 9.3005
R9783 gnd.n2455 gnd.n2454 9.3005
R9784 gnd.n2453 gnd.n2407 9.3005
R9785 gnd.n2452 gnd.n2451 9.3005
R9786 gnd.n2448 gnd.n2410 9.3005
R9787 gnd.n2447 gnd.n2444 9.3005
R9788 gnd.n2443 gnd.n2411 9.3005
R9789 gnd.n2442 gnd.n2441 9.3005
R9790 gnd.n2438 gnd.n2412 9.3005
R9791 gnd.n2437 gnd.n2434 9.3005
R9792 gnd.n2433 gnd.n2413 9.3005
R9793 gnd.n2432 gnd.n2431 9.3005
R9794 gnd.n2428 gnd.n2414 9.3005
R9795 gnd.n2427 gnd.n2424 9.3005
R9796 gnd.n2423 gnd.n2415 9.3005
R9797 gnd.n2422 gnd.n2421 9.3005
R9798 gnd.n2418 gnd.n2416 9.3005
R9799 gnd.n2417 gnd.n1129 9.3005
R9800 gnd.n2456 gnd.n2403 9.3005
R9801 gnd.n2458 gnd.n2457 9.3005
R9802 gnd.n2321 gnd.n1131 9.3005
R9803 gnd.n2324 gnd.n2322 9.3005
R9804 gnd.n2325 gnd.n1152 9.3005
R9805 gnd.n2327 gnd.n1153 9.3005
R9806 gnd.n2328 gnd.n1154 9.3005
R9807 gnd.n2331 gnd.n2329 9.3005
R9808 gnd.n2332 gnd.n1170 9.3005
R9809 gnd.n2334 gnd.n1171 9.3005
R9810 gnd.n2335 gnd.n1172 9.3005
R9811 gnd.n2338 gnd.n2336 9.3005
R9812 gnd.n2339 gnd.n1188 9.3005
R9813 gnd.n2341 gnd.n1189 9.3005
R9814 gnd.n2342 gnd.n1190 9.3005
R9815 gnd.n2345 gnd.n2343 9.3005
R9816 gnd.n2346 gnd.n1208 9.3005
R9817 gnd.n2348 gnd.n1209 9.3005
R9818 gnd.n2349 gnd.n1210 9.3005
R9819 gnd.n2352 gnd.n2350 9.3005
R9820 gnd.n2353 gnd.n1226 9.3005
R9821 gnd.n2355 gnd.n1227 9.3005
R9822 gnd.n2356 gnd.n1228 9.3005
R9823 gnd.n2359 gnd.n2357 9.3005
R9824 gnd.n2360 gnd.n1246 9.3005
R9825 gnd.n2362 gnd.n1247 9.3005
R9826 gnd.n2363 gnd.n1248 9.3005
R9827 gnd.n2366 gnd.n2364 9.3005
R9828 gnd.n2367 gnd.n1264 9.3005
R9829 gnd.n2369 gnd.n1265 9.3005
R9830 gnd.n2370 gnd.n1266 9.3005
R9831 gnd.n2373 gnd.n2371 9.3005
R9832 gnd.n2374 gnd.n1284 9.3005
R9833 gnd.n2376 gnd.n1285 9.3005
R9834 gnd.n2377 gnd.n1286 9.3005
R9835 gnd.n2380 gnd.n2378 9.3005
R9836 gnd.n2381 gnd.n1304 9.3005
R9837 gnd.n2533 gnd.n1305 9.3005
R9838 gnd.n2534 gnd.n1306 9.3005
R9839 gnd.n2541 gnd.n2535 9.3005
R9840 gnd.n2540 gnd.n1325 9.3005
R9841 gnd.n2539 gnd.n1326 9.3005
R9842 gnd.n2538 gnd.n1327 9.3005
R9843 gnd.n2537 gnd.n2536 9.3005
R9844 gnd.n4037 gnd.n1130 9.3005
R9845 gnd.n1132 gnd.n1131 9.3005
R9846 gnd.n2322 gnd.n1151 9.3005
R9847 gnd.n4023 gnd.n1152 9.3005
R9848 gnd.n4022 gnd.n1153 9.3005
R9849 gnd.n4021 gnd.n1154 9.3005
R9850 gnd.n2329 gnd.n1155 9.3005
R9851 gnd.n4011 gnd.n1170 9.3005
R9852 gnd.n4010 gnd.n1171 9.3005
R9853 gnd.n4009 gnd.n1172 9.3005
R9854 gnd.n2336 gnd.n1173 9.3005
R9855 gnd.n3999 gnd.n1188 9.3005
R9856 gnd.n3998 gnd.n1189 9.3005
R9857 gnd.n3997 gnd.n1190 9.3005
R9858 gnd.n2343 gnd.n1191 9.3005
R9859 gnd.n3987 gnd.n1208 9.3005
R9860 gnd.n3986 gnd.n1209 9.3005
R9861 gnd.n3985 gnd.n1210 9.3005
R9862 gnd.n2350 gnd.n1211 9.3005
R9863 gnd.n3975 gnd.n1226 9.3005
R9864 gnd.n3974 gnd.n1227 9.3005
R9865 gnd.n3973 gnd.n1228 9.3005
R9866 gnd.n2357 gnd.n1229 9.3005
R9867 gnd.n3963 gnd.n1246 9.3005
R9868 gnd.n3962 gnd.n1247 9.3005
R9869 gnd.n3961 gnd.n1248 9.3005
R9870 gnd.n2364 gnd.n1249 9.3005
R9871 gnd.n3951 gnd.n1264 9.3005
R9872 gnd.n3950 gnd.n1265 9.3005
R9873 gnd.n3949 gnd.n1266 9.3005
R9874 gnd.n2371 gnd.n1267 9.3005
R9875 gnd.n3939 gnd.n1284 9.3005
R9876 gnd.n3938 gnd.n1285 9.3005
R9877 gnd.n3937 gnd.n1286 9.3005
R9878 gnd.n2378 gnd.n1287 9.3005
R9879 gnd.n3927 gnd.n1304 9.3005
R9880 gnd.n3926 gnd.n1305 9.3005
R9881 gnd.n3925 gnd.n1306 9.3005
R9882 gnd.n2535 gnd.n1307 9.3005
R9883 gnd.n3915 gnd.n1325 9.3005
R9884 gnd.n3914 gnd.n1326 9.3005
R9885 gnd.n3913 gnd.n1327 9.3005
R9886 gnd.n2536 gnd.n1328 9.3005
R9887 gnd.n4037 gnd.n4036 9.3005
R9888 gnd.n5777 gnd.n5776 9.3005
R9889 gnd.n5778 gnd.n837 9.3005
R9890 gnd.n5780 gnd.n5779 9.3005
R9891 gnd.n833 gnd.n832 9.3005
R9892 gnd.n5787 gnd.n5786 9.3005
R9893 gnd.n5788 gnd.n831 9.3005
R9894 gnd.n5790 gnd.n5789 9.3005
R9895 gnd.n827 gnd.n826 9.3005
R9896 gnd.n5797 gnd.n5796 9.3005
R9897 gnd.n5798 gnd.n825 9.3005
R9898 gnd.n5800 gnd.n5799 9.3005
R9899 gnd.n821 gnd.n820 9.3005
R9900 gnd.n5807 gnd.n5806 9.3005
R9901 gnd.n5808 gnd.n819 9.3005
R9902 gnd.n5810 gnd.n5809 9.3005
R9903 gnd.n815 gnd.n814 9.3005
R9904 gnd.n5817 gnd.n5816 9.3005
R9905 gnd.n5818 gnd.n813 9.3005
R9906 gnd.n5820 gnd.n5819 9.3005
R9907 gnd.n809 gnd.n808 9.3005
R9908 gnd.n5827 gnd.n5826 9.3005
R9909 gnd.n5828 gnd.n807 9.3005
R9910 gnd.n5830 gnd.n5829 9.3005
R9911 gnd.n803 gnd.n802 9.3005
R9912 gnd.n5837 gnd.n5836 9.3005
R9913 gnd.n5838 gnd.n801 9.3005
R9914 gnd.n5840 gnd.n5839 9.3005
R9915 gnd.n797 gnd.n796 9.3005
R9916 gnd.n5847 gnd.n5846 9.3005
R9917 gnd.n5848 gnd.n795 9.3005
R9918 gnd.n5850 gnd.n5849 9.3005
R9919 gnd.n791 gnd.n790 9.3005
R9920 gnd.n5857 gnd.n5856 9.3005
R9921 gnd.n5858 gnd.n789 9.3005
R9922 gnd.n5860 gnd.n5859 9.3005
R9923 gnd.n785 gnd.n784 9.3005
R9924 gnd.n5867 gnd.n5866 9.3005
R9925 gnd.n5868 gnd.n783 9.3005
R9926 gnd.n5870 gnd.n5869 9.3005
R9927 gnd.n779 gnd.n778 9.3005
R9928 gnd.n5877 gnd.n5876 9.3005
R9929 gnd.n5878 gnd.n777 9.3005
R9930 gnd.n5880 gnd.n5879 9.3005
R9931 gnd.n773 gnd.n772 9.3005
R9932 gnd.n5887 gnd.n5886 9.3005
R9933 gnd.n5888 gnd.n771 9.3005
R9934 gnd.n5890 gnd.n5889 9.3005
R9935 gnd.n767 gnd.n766 9.3005
R9936 gnd.n5897 gnd.n5896 9.3005
R9937 gnd.n5898 gnd.n765 9.3005
R9938 gnd.n5900 gnd.n5899 9.3005
R9939 gnd.n761 gnd.n760 9.3005
R9940 gnd.n5907 gnd.n5906 9.3005
R9941 gnd.n5908 gnd.n759 9.3005
R9942 gnd.n5910 gnd.n5909 9.3005
R9943 gnd.n755 gnd.n754 9.3005
R9944 gnd.n5917 gnd.n5916 9.3005
R9945 gnd.n5918 gnd.n753 9.3005
R9946 gnd.n5920 gnd.n5919 9.3005
R9947 gnd.n749 gnd.n748 9.3005
R9948 gnd.n5927 gnd.n5926 9.3005
R9949 gnd.n5928 gnd.n747 9.3005
R9950 gnd.n5930 gnd.n5929 9.3005
R9951 gnd.n743 gnd.n742 9.3005
R9952 gnd.n5937 gnd.n5936 9.3005
R9953 gnd.n5938 gnd.n741 9.3005
R9954 gnd.n5940 gnd.n5939 9.3005
R9955 gnd.n737 gnd.n736 9.3005
R9956 gnd.n5947 gnd.n5946 9.3005
R9957 gnd.n5948 gnd.n735 9.3005
R9958 gnd.n5950 gnd.n5949 9.3005
R9959 gnd.n731 gnd.n730 9.3005
R9960 gnd.n5957 gnd.n5956 9.3005
R9961 gnd.n5958 gnd.n729 9.3005
R9962 gnd.n5960 gnd.n5959 9.3005
R9963 gnd.n725 gnd.n724 9.3005
R9964 gnd.n5967 gnd.n5966 9.3005
R9965 gnd.n5968 gnd.n723 9.3005
R9966 gnd.n5970 gnd.n5969 9.3005
R9967 gnd.n719 gnd.n718 9.3005
R9968 gnd.n5977 gnd.n5976 9.3005
R9969 gnd.n5978 gnd.n717 9.3005
R9970 gnd.n5980 gnd.n5979 9.3005
R9971 gnd.n713 gnd.n712 9.3005
R9972 gnd.n5987 gnd.n5986 9.3005
R9973 gnd.n5988 gnd.n711 9.3005
R9974 gnd.n5990 gnd.n5989 9.3005
R9975 gnd.n707 gnd.n706 9.3005
R9976 gnd.n5997 gnd.n5996 9.3005
R9977 gnd.n5998 gnd.n705 9.3005
R9978 gnd.n6000 gnd.n5999 9.3005
R9979 gnd.n701 gnd.n700 9.3005
R9980 gnd.n6007 gnd.n6006 9.3005
R9981 gnd.n6008 gnd.n699 9.3005
R9982 gnd.n6010 gnd.n6009 9.3005
R9983 gnd.n695 gnd.n694 9.3005
R9984 gnd.n6017 gnd.n6016 9.3005
R9985 gnd.n6018 gnd.n693 9.3005
R9986 gnd.n6020 gnd.n6019 9.3005
R9987 gnd.n689 gnd.n688 9.3005
R9988 gnd.n6027 gnd.n6026 9.3005
R9989 gnd.n6028 gnd.n687 9.3005
R9990 gnd.n6030 gnd.n6029 9.3005
R9991 gnd.n683 gnd.n682 9.3005
R9992 gnd.n6037 gnd.n6036 9.3005
R9993 gnd.n6038 gnd.n681 9.3005
R9994 gnd.n6040 gnd.n6039 9.3005
R9995 gnd.n677 gnd.n676 9.3005
R9996 gnd.n6047 gnd.n6046 9.3005
R9997 gnd.n6048 gnd.n675 9.3005
R9998 gnd.n6050 gnd.n6049 9.3005
R9999 gnd.n671 gnd.n670 9.3005
R10000 gnd.n6057 gnd.n6056 9.3005
R10001 gnd.n6058 gnd.n669 9.3005
R10002 gnd.n6060 gnd.n6059 9.3005
R10003 gnd.n665 gnd.n664 9.3005
R10004 gnd.n6067 gnd.n6066 9.3005
R10005 gnd.n6068 gnd.n663 9.3005
R10006 gnd.n6070 gnd.n6069 9.3005
R10007 gnd.n659 gnd.n658 9.3005
R10008 gnd.n6077 gnd.n6076 9.3005
R10009 gnd.n6078 gnd.n657 9.3005
R10010 gnd.n6080 gnd.n6079 9.3005
R10011 gnd.n653 gnd.n652 9.3005
R10012 gnd.n6087 gnd.n6086 9.3005
R10013 gnd.n6088 gnd.n651 9.3005
R10014 gnd.n6090 gnd.n6089 9.3005
R10015 gnd.n647 gnd.n646 9.3005
R10016 gnd.n6097 gnd.n6096 9.3005
R10017 gnd.n6100 gnd.n6099 9.3005
R10018 gnd.n641 gnd.n640 9.3005
R10019 gnd.n6107 gnd.n6106 9.3005
R10020 gnd.n6108 gnd.n639 9.3005
R10021 gnd.n6110 gnd.n6109 9.3005
R10022 gnd.n635 gnd.n634 9.3005
R10023 gnd.n6117 gnd.n6116 9.3005
R10024 gnd.n6118 gnd.n633 9.3005
R10025 gnd.n6120 gnd.n6119 9.3005
R10026 gnd.n629 gnd.n628 9.3005
R10027 gnd.n6127 gnd.n6126 9.3005
R10028 gnd.n6128 gnd.n627 9.3005
R10029 gnd.n6130 gnd.n6129 9.3005
R10030 gnd.n623 gnd.n622 9.3005
R10031 gnd.n6137 gnd.n6136 9.3005
R10032 gnd.n6138 gnd.n621 9.3005
R10033 gnd.n6140 gnd.n6139 9.3005
R10034 gnd.n617 gnd.n616 9.3005
R10035 gnd.n6147 gnd.n6146 9.3005
R10036 gnd.n6148 gnd.n615 9.3005
R10037 gnd.n6150 gnd.n6149 9.3005
R10038 gnd.n611 gnd.n610 9.3005
R10039 gnd.n6157 gnd.n6156 9.3005
R10040 gnd.n6158 gnd.n609 9.3005
R10041 gnd.n6160 gnd.n6159 9.3005
R10042 gnd.n605 gnd.n604 9.3005
R10043 gnd.n6167 gnd.n6166 9.3005
R10044 gnd.n6168 gnd.n603 9.3005
R10045 gnd.n6170 gnd.n6169 9.3005
R10046 gnd.n599 gnd.n598 9.3005
R10047 gnd.n6177 gnd.n6176 9.3005
R10048 gnd.n6178 gnd.n597 9.3005
R10049 gnd.n6180 gnd.n6179 9.3005
R10050 gnd.n593 gnd.n592 9.3005
R10051 gnd.n6187 gnd.n6186 9.3005
R10052 gnd.n6188 gnd.n591 9.3005
R10053 gnd.n6190 gnd.n6189 9.3005
R10054 gnd.n587 gnd.n586 9.3005
R10055 gnd.n6197 gnd.n6196 9.3005
R10056 gnd.n6198 gnd.n585 9.3005
R10057 gnd.n6200 gnd.n6199 9.3005
R10058 gnd.n581 gnd.n580 9.3005
R10059 gnd.n6207 gnd.n6206 9.3005
R10060 gnd.n6208 gnd.n579 9.3005
R10061 gnd.n6210 gnd.n6209 9.3005
R10062 gnd.n575 gnd.n574 9.3005
R10063 gnd.n6217 gnd.n6216 9.3005
R10064 gnd.n6218 gnd.n573 9.3005
R10065 gnd.n6220 gnd.n6219 9.3005
R10066 gnd.n569 gnd.n568 9.3005
R10067 gnd.n6227 gnd.n6226 9.3005
R10068 gnd.n6228 gnd.n567 9.3005
R10069 gnd.n6230 gnd.n6229 9.3005
R10070 gnd.n563 gnd.n562 9.3005
R10071 gnd.n6237 gnd.n6236 9.3005
R10072 gnd.n6238 gnd.n561 9.3005
R10073 gnd.n6240 gnd.n6239 9.3005
R10074 gnd.n557 gnd.n556 9.3005
R10075 gnd.n6247 gnd.n6246 9.3005
R10076 gnd.n6248 gnd.n555 9.3005
R10077 gnd.n6250 gnd.n6249 9.3005
R10078 gnd.n551 gnd.n550 9.3005
R10079 gnd.n6257 gnd.n6256 9.3005
R10080 gnd.n6258 gnd.n549 9.3005
R10081 gnd.n6260 gnd.n6259 9.3005
R10082 gnd.n545 gnd.n544 9.3005
R10083 gnd.n6267 gnd.n6266 9.3005
R10084 gnd.n6268 gnd.n543 9.3005
R10085 gnd.n6270 gnd.n6269 9.3005
R10086 gnd.n539 gnd.n538 9.3005
R10087 gnd.n6277 gnd.n6276 9.3005
R10088 gnd.n6278 gnd.n537 9.3005
R10089 gnd.n6280 gnd.n6279 9.3005
R10090 gnd.n533 gnd.n532 9.3005
R10091 gnd.n6287 gnd.n6286 9.3005
R10092 gnd.n6288 gnd.n531 9.3005
R10093 gnd.n6290 gnd.n6289 9.3005
R10094 gnd.n527 gnd.n526 9.3005
R10095 gnd.n6297 gnd.n6296 9.3005
R10096 gnd.n6298 gnd.n525 9.3005
R10097 gnd.n6302 gnd.n6299 9.3005
R10098 gnd.n6301 gnd.n6300 9.3005
R10099 gnd.n521 gnd.n520 9.3005
R10100 gnd.n6311 gnd.n6310 9.3005
R10101 gnd.n6098 gnd.n645 9.3005
R10102 gnd.n2310 gnd.n2309 9.3005
R10103 gnd.n2311 gnd.n2303 9.3005
R10104 gnd.n2313 gnd.n2312 9.3005
R10105 gnd.n2301 gnd.n2300 9.3005
R10106 gnd.n2569 gnd.n2568 9.3005
R10107 gnd.n2570 gnd.n2299 9.3005
R10108 gnd.n2595 gnd.n2571 9.3005
R10109 gnd.n2594 gnd.n2572 9.3005
R10110 gnd.n2593 gnd.n2573 9.3005
R10111 gnd.n2576 gnd.n2574 9.3005
R10112 gnd.n2588 gnd.n2577 9.3005
R10113 gnd.n2587 gnd.n2578 9.3005
R10114 gnd.n2586 gnd.n2579 9.3005
R10115 gnd.n2581 gnd.n2580 9.3005
R10116 gnd.n2093 gnd.n2092 9.3005
R10117 gnd.n2683 gnd.n2682 9.3005
R10118 gnd.n2684 gnd.n2091 9.3005
R10119 gnd.n2688 gnd.n2685 9.3005
R10120 gnd.n2687 gnd.n2686 9.3005
R10121 gnd.n2068 gnd.n2067 9.3005
R10122 gnd.n2713 gnd.n2712 9.3005
R10123 gnd.n2714 gnd.n2066 9.3005
R10124 gnd.n2718 gnd.n2715 9.3005
R10125 gnd.n2717 gnd.n2716 9.3005
R10126 gnd.n2043 gnd.n2042 9.3005
R10127 gnd.n2743 gnd.n2742 9.3005
R10128 gnd.n2744 gnd.n2041 9.3005
R10129 gnd.n2748 gnd.n2745 9.3005
R10130 gnd.n2747 gnd.n2746 9.3005
R10131 gnd.n2018 gnd.n2017 9.3005
R10132 gnd.n2776 gnd.n2775 9.3005
R10133 gnd.n2777 gnd.n2016 9.3005
R10134 gnd.n2793 gnd.n2778 9.3005
R10135 gnd.n2792 gnd.n2779 9.3005
R10136 gnd.n2791 gnd.n2780 9.3005
R10137 gnd.n2783 gnd.n2781 9.3005
R10138 gnd.n2787 gnd.n2784 9.3005
R10139 gnd.n2786 gnd.n2785 9.3005
R10140 gnd.n1988 gnd.n1987 9.3005
R10141 gnd.n2928 gnd.n2927 9.3005
R10142 gnd.n2929 gnd.n1986 9.3005
R10143 gnd.n2933 gnd.n2930 9.3005
R10144 gnd.n2932 gnd.n2931 9.3005
R10145 gnd.n1960 gnd.n1959 9.3005
R10146 gnd.n2970 gnd.n2969 9.3005
R10147 gnd.n2971 gnd.n1958 9.3005
R10148 gnd.n2973 gnd.n2972 9.3005
R10149 gnd.n1937 gnd.n1936 9.3005
R10150 gnd.n3014 gnd.n3013 9.3005
R10151 gnd.n3015 gnd.n1935 9.3005
R10152 gnd.n3017 gnd.n3016 9.3005
R10153 gnd.n1919 gnd.n1918 9.3005
R10154 gnd.n3070 gnd.n3069 9.3005
R10155 gnd.n3071 gnd.n1917 9.3005
R10156 gnd.n3073 gnd.n3072 9.3005
R10157 gnd.n1897 gnd.n1896 9.3005
R10158 gnd.n3098 gnd.n3097 9.3005
R10159 gnd.n3099 gnd.n1895 9.3005
R10160 gnd.n3103 gnd.n3100 9.3005
R10161 gnd.n3102 gnd.n3101 9.3005
R10162 gnd.n1865 gnd.n1864 9.3005
R10163 gnd.n3143 gnd.n3142 9.3005
R10164 gnd.n3144 gnd.n1863 9.3005
R10165 gnd.n3146 gnd.n3145 9.3005
R10166 gnd.n1841 gnd.n1840 9.3005
R10167 gnd.n3184 gnd.n3183 9.3005
R10168 gnd.n3185 gnd.n1839 9.3005
R10169 gnd.n3187 gnd.n3186 9.3005
R10170 gnd.n1824 gnd.n1823 9.3005
R10171 gnd.n3243 gnd.n3242 9.3005
R10172 gnd.n3244 gnd.n1822 9.3005
R10173 gnd.n3246 gnd.n3245 9.3005
R10174 gnd.n1803 gnd.n1802 9.3005
R10175 gnd.n3270 gnd.n3269 9.3005
R10176 gnd.n3271 gnd.n1801 9.3005
R10177 gnd.n3275 gnd.n3272 9.3005
R10178 gnd.n3274 gnd.n3273 9.3005
R10179 gnd.n1774 gnd.n1773 9.3005
R10180 gnd.n3317 gnd.n3316 9.3005
R10181 gnd.n3318 gnd.n1772 9.3005
R10182 gnd.n3320 gnd.n3319 9.3005
R10183 gnd.n1751 gnd.n1750 9.3005
R10184 gnd.n3358 gnd.n3357 9.3005
R10185 gnd.n3359 gnd.n1749 9.3005
R10186 gnd.n3361 gnd.n3360 9.3005
R10187 gnd.n1735 gnd.n1734 9.3005
R10188 gnd.n3400 gnd.n3399 9.3005
R10189 gnd.n3401 gnd.n1733 9.3005
R10190 gnd.n3403 gnd.n3402 9.3005
R10191 gnd.n1643 gnd.n1642 9.3005
R10192 gnd.n3547 gnd.n3546 9.3005
R10193 gnd.n3548 gnd.n1641 9.3005
R10194 gnd.n3550 gnd.n3549 9.3005
R10195 gnd.n1630 gnd.n1629 9.3005
R10196 gnd.n3567 gnd.n3566 9.3005
R10197 gnd.n3568 gnd.n1628 9.3005
R10198 gnd.n3570 gnd.n3569 9.3005
R10199 gnd.n1619 gnd.n1618 9.3005
R10200 gnd.n3589 gnd.n3588 9.3005
R10201 gnd.n3590 gnd.n1617 9.3005
R10202 gnd.n3592 gnd.n3591 9.3005
R10203 gnd.n1606 gnd.n1605 9.3005
R10204 gnd.n3609 gnd.n3608 9.3005
R10205 gnd.n3610 gnd.n1604 9.3005
R10206 gnd.n3612 gnd.n3611 9.3005
R10207 gnd.n1593 gnd.n1592 9.3005
R10208 gnd.n3629 gnd.n3628 9.3005
R10209 gnd.n3630 gnd.n1591 9.3005
R10210 gnd.n3632 gnd.n3631 9.3005
R10211 gnd.n1579 gnd.n1578 9.3005
R10212 gnd.n3649 gnd.n3648 9.3005
R10213 gnd.n3650 gnd.n1577 9.3005
R10214 gnd.n3658 gnd.n3651 9.3005
R10215 gnd.n3657 gnd.n3652 9.3005
R10216 gnd.n3656 gnd.n3654 9.3005
R10217 gnd.n3653 gnd.n493 9.3005
R10218 gnd.n6336 gnd.n494 9.3005
R10219 gnd.n6335 gnd.n495 9.3005
R10220 gnd.n6334 gnd.n496 9.3005
R10221 gnd.n509 gnd.n497 9.3005
R10222 gnd.n510 gnd.n499 9.3005
R10223 gnd.n511 gnd.n508 9.3005
R10224 gnd.n6320 gnd.n512 9.3005
R10225 gnd.n6319 gnd.n513 9.3005
R10226 gnd.n6318 gnd.n514 9.3005
R10227 gnd.n518 gnd.n515 9.3005
R10228 gnd.n6314 gnd.n519 9.3005
R10229 gnd.n6313 gnd.n6312 9.3005
R10230 gnd.n2306 gnd.n2305 9.3005
R10231 gnd.n5608 gnd.n1005 9.3005
R10232 gnd.n5609 gnd.n1004 9.3005
R10233 gnd.n5610 gnd.n1003 9.3005
R10234 gnd.n1002 gnd.n998 9.3005
R10235 gnd.n5616 gnd.n997 9.3005
R10236 gnd.n5617 gnd.n996 9.3005
R10237 gnd.n5618 gnd.n995 9.3005
R10238 gnd.n994 gnd.n990 9.3005
R10239 gnd.n5624 gnd.n989 9.3005
R10240 gnd.n5625 gnd.n988 9.3005
R10241 gnd.n5626 gnd.n987 9.3005
R10242 gnd.n986 gnd.n982 9.3005
R10243 gnd.n5632 gnd.n981 9.3005
R10244 gnd.n5633 gnd.n980 9.3005
R10245 gnd.n5634 gnd.n979 9.3005
R10246 gnd.n978 gnd.n974 9.3005
R10247 gnd.n5640 gnd.n973 9.3005
R10248 gnd.n5641 gnd.n972 9.3005
R10249 gnd.n5642 gnd.n971 9.3005
R10250 gnd.n970 gnd.n966 9.3005
R10251 gnd.n5648 gnd.n965 9.3005
R10252 gnd.n5649 gnd.n964 9.3005
R10253 gnd.n5650 gnd.n963 9.3005
R10254 gnd.n962 gnd.n958 9.3005
R10255 gnd.n5656 gnd.n957 9.3005
R10256 gnd.n5657 gnd.n956 9.3005
R10257 gnd.n5658 gnd.n955 9.3005
R10258 gnd.n954 gnd.n950 9.3005
R10259 gnd.n5664 gnd.n949 9.3005
R10260 gnd.n5665 gnd.n948 9.3005
R10261 gnd.n5666 gnd.n947 9.3005
R10262 gnd.n946 gnd.n942 9.3005
R10263 gnd.n5672 gnd.n941 9.3005
R10264 gnd.n5673 gnd.n940 9.3005
R10265 gnd.n5674 gnd.n939 9.3005
R10266 gnd.n938 gnd.n934 9.3005
R10267 gnd.n5680 gnd.n933 9.3005
R10268 gnd.n5681 gnd.n932 9.3005
R10269 gnd.n5682 gnd.n931 9.3005
R10270 gnd.n930 gnd.n926 9.3005
R10271 gnd.n5688 gnd.n925 9.3005
R10272 gnd.n5689 gnd.n924 9.3005
R10273 gnd.n5690 gnd.n923 9.3005
R10274 gnd.n922 gnd.n918 9.3005
R10275 gnd.n5696 gnd.n917 9.3005
R10276 gnd.n5697 gnd.n916 9.3005
R10277 gnd.n5698 gnd.n915 9.3005
R10278 gnd.n914 gnd.n910 9.3005
R10279 gnd.n5704 gnd.n909 9.3005
R10280 gnd.n5705 gnd.n908 9.3005
R10281 gnd.n5706 gnd.n907 9.3005
R10282 gnd.n906 gnd.n902 9.3005
R10283 gnd.n5712 gnd.n901 9.3005
R10284 gnd.n5713 gnd.n900 9.3005
R10285 gnd.n5714 gnd.n899 9.3005
R10286 gnd.n898 gnd.n894 9.3005
R10287 gnd.n5720 gnd.n893 9.3005
R10288 gnd.n5721 gnd.n892 9.3005
R10289 gnd.n5722 gnd.n891 9.3005
R10290 gnd.n890 gnd.n886 9.3005
R10291 gnd.n5728 gnd.n885 9.3005
R10292 gnd.n5729 gnd.n884 9.3005
R10293 gnd.n5730 gnd.n883 9.3005
R10294 gnd.n882 gnd.n878 9.3005
R10295 gnd.n5736 gnd.n877 9.3005
R10296 gnd.n5737 gnd.n876 9.3005
R10297 gnd.n5738 gnd.n875 9.3005
R10298 gnd.n874 gnd.n870 9.3005
R10299 gnd.n5744 gnd.n869 9.3005
R10300 gnd.n5745 gnd.n868 9.3005
R10301 gnd.n5746 gnd.n867 9.3005
R10302 gnd.n866 gnd.n862 9.3005
R10303 gnd.n5752 gnd.n861 9.3005
R10304 gnd.n5753 gnd.n860 9.3005
R10305 gnd.n5754 gnd.n859 9.3005
R10306 gnd.n858 gnd.n854 9.3005
R10307 gnd.n5760 gnd.n853 9.3005
R10308 gnd.n5761 gnd.n852 9.3005
R10309 gnd.n5762 gnd.n851 9.3005
R10310 gnd.n850 gnd.n846 9.3005
R10311 gnd.n5768 gnd.n845 9.3005
R10312 gnd.n5769 gnd.n844 9.3005
R10313 gnd.n5770 gnd.n843 9.3005
R10314 gnd.n842 gnd.n838 9.3005
R10315 gnd.n2304 gnd.n1006 9.3005
R10316 gnd.n6359 gnd.n452 9.3005
R10317 gnd.n2673 gnd.n2672 9.3005
R10318 gnd.n2674 gnd.n2097 9.3005
R10319 gnd.n2677 gnd.n2676 9.3005
R10320 gnd.n2675 gnd.n2098 9.3005
R10321 gnd.n2075 gnd.n2074 9.3005
R10322 gnd.n2703 gnd.n2702 9.3005
R10323 gnd.n2704 gnd.n2072 9.3005
R10324 gnd.n2707 gnd.n2706 9.3005
R10325 gnd.n2705 gnd.n2073 9.3005
R10326 gnd.n2050 gnd.n2049 9.3005
R10327 gnd.n2733 gnd.n2732 9.3005
R10328 gnd.n2734 gnd.n2047 9.3005
R10329 gnd.n2737 gnd.n2736 9.3005
R10330 gnd.n2735 gnd.n2048 9.3005
R10331 gnd.n2025 gnd.n2024 9.3005
R10332 gnd.n2763 gnd.n2762 9.3005
R10333 gnd.n2764 gnd.n2022 9.3005
R10334 gnd.n2770 gnd.n2769 9.3005
R10335 gnd.n2768 gnd.n2023 9.3005
R10336 gnd.n2767 gnd.n2766 9.3005
R10337 gnd.n2765 gnd.n2001 9.3005
R10338 gnd.n1999 gnd.n1998 9.3005
R10339 gnd.n2879 gnd.n2878 9.3005
R10340 gnd.n2880 gnd.n1996 9.3005
R10341 gnd.n2886 gnd.n2885 9.3005
R10342 gnd.n2884 gnd.n1997 9.3005
R10343 gnd.n2883 gnd.n2882 9.3005
R10344 gnd.n1974 gnd.n1973 9.3005
R10345 gnd.n2947 gnd.n2946 9.3005
R10346 gnd.n2948 gnd.n1972 9.3005
R10347 gnd.n2950 gnd.n2949 9.3005
R10348 gnd.n1952 gnd.n1951 9.3005
R10349 gnd.n2980 gnd.n2979 9.3005
R10350 gnd.n2981 gnd.n1949 9.3005
R10351 gnd.n2993 gnd.n2992 9.3005
R10352 gnd.n2991 gnd.n1950 9.3005
R10353 gnd.n2990 gnd.n2989 9.3005
R10354 gnd.n2988 gnd.n2982 9.3005
R10355 gnd.n2987 gnd.n2986 9.3005
R10356 gnd.n1912 gnd.n1911 9.3005
R10357 gnd.n3080 gnd.n3079 9.3005
R10358 gnd.n3081 gnd.n1909 9.3005
R10359 gnd.n3084 gnd.n3083 9.3005
R10360 gnd.n3082 gnd.n1910 9.3005
R10361 gnd.n1882 gnd.n1881 9.3005
R10362 gnd.n3116 gnd.n3115 9.3005
R10363 gnd.n3117 gnd.n1879 9.3005
R10364 gnd.n3123 gnd.n3122 9.3005
R10365 gnd.n3121 gnd.n1880 9.3005
R10366 gnd.n3120 gnd.n3119 9.3005
R10367 gnd.n1853 gnd.n1852 9.3005
R10368 gnd.n3164 gnd.n3163 9.3005
R10369 gnd.n3165 gnd.n1850 9.3005
R10370 gnd.n3171 gnd.n3170 9.3005
R10371 gnd.n3169 gnd.n1851 9.3005
R10372 gnd.n3168 gnd.n3167 9.3005
R10373 gnd.n1816 gnd.n1815 9.3005
R10374 gnd.n3252 gnd.n3251 9.3005
R10375 gnd.n3253 gnd.n1813 9.3005
R10376 gnd.n3256 gnd.n3255 9.3005
R10377 gnd.n3254 gnd.n1814 9.3005
R10378 gnd.n1790 gnd.n1789 9.3005
R10379 gnd.n3288 gnd.n3287 9.3005
R10380 gnd.n3289 gnd.n1787 9.3005
R10381 gnd.n3297 gnd.n3296 9.3005
R10382 gnd.n3295 gnd.n1788 9.3005
R10383 gnd.n3294 gnd.n3293 9.3005
R10384 gnd.n1763 gnd.n1762 9.3005
R10385 gnd.n3338 gnd.n3337 9.3005
R10386 gnd.n3339 gnd.n1760 9.3005
R10387 gnd.n3345 gnd.n3344 9.3005
R10388 gnd.n3343 gnd.n1761 9.3005
R10389 gnd.n3342 gnd.n3341 9.3005
R10390 gnd.n1729 gnd.n1728 9.3005
R10391 gnd.n3409 gnd.n3408 9.3005
R10392 gnd.n3410 gnd.n1726 9.3005
R10393 gnd.n3413 gnd.n3412 9.3005
R10394 gnd.n3411 gnd.n1727 9.3005
R10395 gnd.n1637 gnd.n1636 9.3005
R10396 gnd.n3557 gnd.n3556 9.3005
R10397 gnd.n3558 gnd.n1635 9.3005
R10398 gnd.n3560 gnd.n3559 9.3005
R10399 gnd.n1624 gnd.n1623 9.3005
R10400 gnd.n3579 gnd.n3578 9.3005
R10401 gnd.n3580 gnd.n1622 9.3005
R10402 gnd.n3582 gnd.n3581 9.3005
R10403 gnd.n1613 gnd.n1612 9.3005
R10404 gnd.n3599 gnd.n3598 9.3005
R10405 gnd.n3600 gnd.n1611 9.3005
R10406 gnd.n3602 gnd.n3601 9.3005
R10407 gnd.n1600 gnd.n1599 9.3005
R10408 gnd.n3619 gnd.n3618 9.3005
R10409 gnd.n3620 gnd.n1598 9.3005
R10410 gnd.n3622 gnd.n3621 9.3005
R10411 gnd.n1587 gnd.n1586 9.3005
R10412 gnd.n3639 gnd.n3638 9.3005
R10413 gnd.n3640 gnd.n1584 9.3005
R10414 gnd.n3643 gnd.n3642 9.3005
R10415 gnd.n3641 gnd.n1585 9.3005
R10416 gnd.n454 gnd.n453 9.3005
R10417 gnd.n6358 gnd.n6357 9.3005
R10418 gnd.n2100 gnd.n2099 9.3005
R10419 gnd.n2556 gnd.n2548 9.3005
R10420 gnd.n2505 gnd.n2504 9.3005
R10421 gnd.n2506 gnd.n2390 9.3005
R10422 gnd.n2508 gnd.n2507 9.3005
R10423 gnd.n2509 gnd.n2389 9.3005
R10424 gnd.n2512 gnd.n2511 9.3005
R10425 gnd.n2513 gnd.n2387 9.3005
R10426 gnd.n2515 gnd.n2514 9.3005
R10427 gnd.n2516 gnd.n2386 9.3005
R10428 gnd.n2519 gnd.n2518 9.3005
R10429 gnd.n2520 gnd.n2384 9.3005
R10430 gnd.n2522 gnd.n2521 9.3005
R10431 gnd.n2523 gnd.n2383 9.3005
R10432 gnd.n2526 gnd.n2525 9.3005
R10433 gnd.n2527 gnd.n2382 9.3005
R10434 gnd.n2529 gnd.n2528 9.3005
R10435 gnd.n2320 gnd.n2319 9.3005
R10436 gnd.n2546 gnd.n2545 9.3005
R10437 gnd.n2547 gnd.n2317 9.3005
R10438 gnd.n2563 gnd.n2562 9.3005
R10439 gnd.n2561 gnd.n2318 9.3005
R10440 gnd.n2560 gnd.n2199 9.3005
R10441 gnd.n2644 gnd.n2643 9.3005
R10442 gnd.n2642 gnd.n2641 9.3005
R10443 gnd.n2145 gnd.n2144 9.3005
R10444 gnd.n2636 gnd.n2635 9.3005
R10445 gnd.n2634 gnd.n2633 9.3005
R10446 gnd.n2155 gnd.n2154 9.3005
R10447 gnd.n2628 gnd.n2627 9.3005
R10448 gnd.n2626 gnd.n2625 9.3005
R10449 gnd.n2165 gnd.n2164 9.3005
R10450 gnd.n2620 gnd.n2619 9.3005
R10451 gnd.n2618 gnd.n2617 9.3005
R10452 gnd.n2175 gnd.n2174 9.3005
R10453 gnd.n2612 gnd.n2611 9.3005
R10454 gnd.n2610 gnd.n2609 9.3005
R10455 gnd.n2185 gnd.n2184 9.3005
R10456 gnd.n2604 gnd.n2603 9.3005
R10457 gnd.n2602 gnd.n2196 9.3005
R10458 gnd.n2601 gnd.n2198 9.3005
R10459 gnd.n2140 gnd.n2135 9.3005
R10460 gnd.n2558 gnd.n2557 9.3005
R10461 gnd.n2552 gnd.n2551 9.3005
R10462 gnd.n2550 gnd.n2192 9.3005
R10463 gnd.n2606 gnd.n2605 9.3005
R10464 gnd.n2608 gnd.n2607 9.3005
R10465 gnd.n2179 gnd.n2178 9.3005
R10466 gnd.n2614 gnd.n2613 9.3005
R10467 gnd.n2616 gnd.n2615 9.3005
R10468 gnd.n2171 gnd.n2170 9.3005
R10469 gnd.n2622 gnd.n2621 9.3005
R10470 gnd.n2624 gnd.n2623 9.3005
R10471 gnd.n2159 gnd.n2158 9.3005
R10472 gnd.n2630 gnd.n2629 9.3005
R10473 gnd.n2632 gnd.n2631 9.3005
R10474 gnd.n2151 gnd.n2150 9.3005
R10475 gnd.n2638 gnd.n2637 9.3005
R10476 gnd.n2640 gnd.n2639 9.3005
R10477 gnd.n2139 gnd.n2138 9.3005
R10478 gnd.n2646 gnd.n2645 9.3005
R10479 gnd.n2648 gnd.n2647 9.3005
R10480 gnd.n2649 gnd.n2133 9.3005
R10481 gnd.n2652 gnd.n2651 9.3005
R10482 gnd.n2653 gnd.n2128 9.3005
R10483 gnd.n2655 gnd.n2654 9.3005
R10484 gnd.n2656 gnd.n2127 9.3005
R10485 gnd.n2658 gnd.n2657 9.3005
R10486 gnd.n2109 gnd.n2108 9.3005
R10487 gnd.n2664 gnd.n2663 9.3005
R10488 gnd.n2668 gnd.n2667 9.3005
R10489 gnd.n2666 gnd.n2107 9.3005
R10490 gnd.n2084 gnd.n2083 9.3005
R10491 gnd.n2694 gnd.n2693 9.3005
R10492 gnd.n2695 gnd.n2081 9.3005
R10493 gnd.n2698 gnd.n2697 9.3005
R10494 gnd.n2696 gnd.n2082 9.3005
R10495 gnd.n2059 gnd.n2058 9.3005
R10496 gnd.n2724 gnd.n2723 9.3005
R10497 gnd.n2725 gnd.n2056 9.3005
R10498 gnd.n2728 gnd.n2727 9.3005
R10499 gnd.n2726 gnd.n2057 9.3005
R10500 gnd.n2033 gnd.n2032 9.3005
R10501 gnd.n2754 gnd.n2753 9.3005
R10502 gnd.n2755 gnd.n2030 9.3005
R10503 gnd.n2758 gnd.n2757 9.3005
R10504 gnd.n2756 gnd.n2031 9.3005
R10505 gnd.n2009 gnd.n2008 9.3005
R10506 gnd.n2799 gnd.n2798 9.3005
R10507 gnd.n2800 gnd.n2006 9.3005
R10508 gnd.n2803 gnd.n2802 9.3005
R10509 gnd.n2801 gnd.n2007 9.3005
R10510 gnd.n1479 gnd.n1477 9.3005
R10511 gnd.n3776 gnd.n3775 9.3005
R10512 gnd.n3774 gnd.n1478 9.3005
R10513 gnd.n3773 gnd.n3772 9.3005
R10514 gnd.n3771 gnd.n1480 9.3005
R10515 gnd.n3770 gnd.n3769 9.3005
R10516 gnd.n3768 gnd.n1484 9.3005
R10517 gnd.n3767 gnd.n3766 9.3005
R10518 gnd.n3765 gnd.n1485 9.3005
R10519 gnd.n3764 gnd.n3763 9.3005
R10520 gnd.n3762 gnd.n1489 9.3005
R10521 gnd.n3761 gnd.n3760 9.3005
R10522 gnd.n3759 gnd.n1490 9.3005
R10523 gnd.n3758 gnd.n3757 9.3005
R10524 gnd.n3756 gnd.n1494 9.3005
R10525 gnd.n3755 gnd.n3754 9.3005
R10526 gnd.n3753 gnd.n1495 9.3005
R10527 gnd.n3752 gnd.n3751 9.3005
R10528 gnd.n3750 gnd.n1499 9.3005
R10529 gnd.n3749 gnd.n3748 9.3005
R10530 gnd.n3747 gnd.n1500 9.3005
R10531 gnd.n3746 gnd.n3745 9.3005
R10532 gnd.n3744 gnd.n1504 9.3005
R10533 gnd.n3743 gnd.n3742 9.3005
R10534 gnd.n3741 gnd.n1505 9.3005
R10535 gnd.n3740 gnd.n3739 9.3005
R10536 gnd.n3738 gnd.n1509 9.3005
R10537 gnd.n3737 gnd.n3736 9.3005
R10538 gnd.n3735 gnd.n1510 9.3005
R10539 gnd.n3734 gnd.n3733 9.3005
R10540 gnd.n3732 gnd.n1514 9.3005
R10541 gnd.n3731 gnd.n3730 9.3005
R10542 gnd.n3729 gnd.n1515 9.3005
R10543 gnd.n3728 gnd.n3727 9.3005
R10544 gnd.n3726 gnd.n1519 9.3005
R10545 gnd.n3725 gnd.n3724 9.3005
R10546 gnd.n3723 gnd.n1520 9.3005
R10547 gnd.n3722 gnd.n3721 9.3005
R10548 gnd.n3720 gnd.n1524 9.3005
R10549 gnd.n3719 gnd.n3718 9.3005
R10550 gnd.n3717 gnd.n1525 9.3005
R10551 gnd.n3716 gnd.n3715 9.3005
R10552 gnd.n3714 gnd.n1529 9.3005
R10553 gnd.n3713 gnd.n3712 9.3005
R10554 gnd.n3711 gnd.n1530 9.3005
R10555 gnd.n3710 gnd.n3709 9.3005
R10556 gnd.n3708 gnd.n1534 9.3005
R10557 gnd.n3707 gnd.n3706 9.3005
R10558 gnd.n3705 gnd.n1535 9.3005
R10559 gnd.n3704 gnd.n3703 9.3005
R10560 gnd.n3702 gnd.n1539 9.3005
R10561 gnd.n3701 gnd.n3700 9.3005
R10562 gnd.n3699 gnd.n1540 9.3005
R10563 gnd.n3698 gnd.n3697 9.3005
R10564 gnd.n3696 gnd.n1544 9.3005
R10565 gnd.n3695 gnd.n3694 9.3005
R10566 gnd.n3693 gnd.n1545 9.3005
R10567 gnd.n3692 gnd.n3691 9.3005
R10568 gnd.n3690 gnd.n1549 9.3005
R10569 gnd.n3689 gnd.n3688 9.3005
R10570 gnd.n3687 gnd.n1550 9.3005
R10571 gnd.n3686 gnd.n3685 9.3005
R10572 gnd.n3684 gnd.n1554 9.3005
R10573 gnd.n3683 gnd.n3682 9.3005
R10574 gnd.n3681 gnd.n1555 9.3005
R10575 gnd.n3680 gnd.n3679 9.3005
R10576 gnd.n3678 gnd.n1559 9.3005
R10577 gnd.n3677 gnd.n3676 9.3005
R10578 gnd.n3675 gnd.n1560 9.3005
R10579 gnd.n3674 gnd.n3673 9.3005
R10580 gnd.n3672 gnd.n1564 9.3005
R10581 gnd.n3671 gnd.n3670 9.3005
R10582 gnd.n3669 gnd.n1565 9.3005
R10583 gnd.n3668 gnd.n3667 9.3005
R10584 gnd.n3666 gnd.n1569 9.3005
R10585 gnd.n3665 gnd.n3664 9.3005
R10586 gnd.n3663 gnd.n1570 9.3005
R10587 gnd.n462 gnd.n461 9.3005
R10588 gnd.n6353 gnd.n6352 9.3005
R10589 gnd.n2665 gnd.n2106 9.3005
R10590 gnd.n6349 gnd.n463 9.3005
R10591 gnd.n6348 gnd.n6347 9.3005
R10592 gnd.n6346 gnd.n466 9.3005
R10593 gnd.n6345 gnd.n6344 9.3005
R10594 gnd.n6343 gnd.n467 9.3005
R10595 gnd.n391 gnd.n389 9.3005
R10596 gnd.n6351 gnd.n6350 9.3005
R10597 gnd.n6371 gnd.n6370 9.3005
R10598 gnd.n438 gnd.n437 9.3005
R10599 gnd.n6377 gnd.n6376 9.3005
R10600 gnd.n6379 gnd.n6378 9.3005
R10601 gnd.n430 gnd.n429 9.3005
R10602 gnd.n6385 gnd.n6384 9.3005
R10603 gnd.n6387 gnd.n6386 9.3005
R10604 gnd.n420 gnd.n419 9.3005
R10605 gnd.n6393 gnd.n6392 9.3005
R10606 gnd.n6395 gnd.n6394 9.3005
R10607 gnd.n412 gnd.n411 9.3005
R10608 gnd.n6401 gnd.n6400 9.3005
R10609 gnd.n6403 gnd.n6402 9.3005
R10610 gnd.n402 gnd.n401 9.3005
R10611 gnd.n6409 gnd.n6408 9.3005
R10612 gnd.n6411 gnd.n6410 9.3005
R10613 gnd.n398 gnd.n396 9.3005
R10614 gnd.n6369 gnd.n6365 9.3005
R10615 gnd.n448 gnd.n447 9.3005
R10616 gnd.n6416 gnd.n6415 9.3005
R10617 gnd.n6414 gnd.n390 9.3005
R10618 gnd.n6413 gnd.n6412 9.3005
R10619 gnd.n397 gnd.n395 9.3005
R10620 gnd.n6407 gnd.n6406 9.3005
R10621 gnd.n6405 gnd.n6404 9.3005
R10622 gnd.n406 gnd.n405 9.3005
R10623 gnd.n6399 gnd.n6398 9.3005
R10624 gnd.n6397 gnd.n6396 9.3005
R10625 gnd.n416 gnd.n415 9.3005
R10626 gnd.n6391 gnd.n6390 9.3005
R10627 gnd.n6389 gnd.n6388 9.3005
R10628 gnd.n424 gnd.n423 9.3005
R10629 gnd.n6383 gnd.n6382 9.3005
R10630 gnd.n6381 gnd.n6380 9.3005
R10631 gnd.n434 gnd.n433 9.3005
R10632 gnd.n6375 gnd.n6374 9.3005
R10633 gnd.n6373 gnd.n6372 9.3005
R10634 gnd.n449 gnd.n444 9.3005
R10635 gnd.n6364 gnd.n6363 9.3005
R10636 gnd.n6362 gnd.n6361 9.3005
R10637 gnd.n6543 gnd.n6542 9.3005
R10638 gnd.n6544 gnd.n269 9.3005
R10639 gnd.n6547 gnd.n6546 9.3005
R10640 gnd.n6545 gnd.n270 9.3005
R10641 gnd.n244 gnd.n243 9.3005
R10642 gnd.n6578 gnd.n6577 9.3005
R10643 gnd.n6579 gnd.n241 9.3005
R10644 gnd.n6592 gnd.n6591 9.3005
R10645 gnd.n6590 gnd.n242 9.3005
R10646 gnd.n6589 gnd.n6588 9.3005
R10647 gnd.n6587 gnd.n6580 9.3005
R10648 gnd.n6586 gnd.n6585 9.3005
R10649 gnd.n6584 gnd.n6583 9.3005
R10650 gnd.n199 gnd.n198 9.3005
R10651 gnd.n6642 gnd.n6641 9.3005
R10652 gnd.n6643 gnd.n196 9.3005
R10653 gnd.n6650 gnd.n6649 9.3005
R10654 gnd.n6648 gnd.n197 9.3005
R10655 gnd.n6647 gnd.n6646 9.3005
R10656 gnd.n6645 gnd.n67 9.3005
R10657 gnd.n272 gnd.n271 9.3005
R10658 gnd.n7112 gnd.n68 9.3005
R10659 gnd.t180 gnd.n4333 9.24152
R10660 gnd.n4235 gnd.t219 9.24152
R10661 gnd.n5503 gnd.t320 9.24152
R10662 gnd.n3347 gnd.t149 9.24152
R10663 gnd.t151 gnd.t180 8.92286
R10664 gnd.n2953 gnd.n1969 8.92286
R10665 gnd.n3003 gnd.n3002 8.92286
R10666 gnd.t25 gnd.n1923 8.92286
R10667 gnd.n1915 gnd.t48 8.92286
R10668 gnd.n3126 gnd.n1876 8.92286
R10669 gnd.n3154 gnd.n1847 8.92286
R10670 gnd.n3260 gnd.t159 8.92286
R10671 gnd.n3208 gnd.t76 8.92286
R10672 gnd.n3301 gnd.n1784 8.92286
R10673 gnd.n3327 gnd.n3326 8.92286
R10674 gnd.n5473 gnd.n5448 8.92171
R10675 gnd.n5441 gnd.n5416 8.92171
R10676 gnd.n5409 gnd.n5384 8.92171
R10677 gnd.n5378 gnd.n5353 8.92171
R10678 gnd.n5346 gnd.n5321 8.92171
R10679 gnd.n5314 gnd.n5289 8.92171
R10680 gnd.n5282 gnd.n5257 8.92171
R10681 gnd.n5251 gnd.n5226 8.92171
R10682 gnd.n1668 gnd.n1650 8.72777
R10683 gnd.n4977 gnd.t177 8.60421
R10684 gnd.n2103 gnd.t249 8.60421
R10685 gnd.t200 gnd.n2053 8.60421
R10686 gnd.t126 gnd.n1867 8.60421
R10687 gnd.n3180 gnd.t102 8.60421
R10688 gnd.n3606 gnd.t124 8.60421
R10689 gnd.t223 gnd.n3660 8.60421
R10690 gnd.n6306 gnd.n116 8.60421
R10691 gnd.n4397 gnd.n4385 8.43656
R10692 gnd.n42 gnd.n30 8.43656
R10693 gnd.n2944 gnd.n1976 8.28555
R10694 gnd.n3057 gnd.n1928 8.28555
R10695 gnd.n3113 gnd.n1884 8.28555
R10696 gnd.n3230 gnd.n1834 8.28555
R10697 gnd.n3285 gnd.n1792 8.28555
R10698 gnd.n3381 gnd.n1744 8.28555
R10699 gnd.n5474 gnd.n5446 8.14595
R10700 gnd.n5442 gnd.n5414 8.14595
R10701 gnd.n5410 gnd.n5382 8.14595
R10702 gnd.n5379 gnd.n5351 8.14595
R10703 gnd.n5347 gnd.n5319 8.14595
R10704 gnd.n5315 gnd.n5287 8.14595
R10705 gnd.n5283 gnd.n5255 8.14595
R10706 gnd.n5252 gnd.n5224 8.14595
R10707 gnd.n2392 gnd.n0 8.10675
R10708 gnd.n7113 gnd.n7112 8.10675
R10709 gnd.n5479 gnd.n5478 7.97301
R10710 gnd.t66 gnd.n4492 7.9669
R10711 gnd.n2660 gnd.n2125 7.9669
R10712 gnd.n2918 gnd.t202 7.9669
R10713 gnd.t192 gnd.t266 7.9669
R10714 gnd.n6339 gnd.n470 7.9669
R10715 gnd.n7113 gnd.n66 7.78567
R10716 gnd.n6369 gnd.n447 7.75808
R10717 gnd.n6834 gnd.n6737 7.75808
R10718 gnd.n2602 gnd.n2601 7.75808
R10719 gnd.n2457 gnd.n2456 7.75808
R10720 gnd.n2935 gnd.n1976 7.64824
R10721 gnd.n3057 gnd.n3056 7.64824
R10722 gnd.t79 gnd.n3105 7.64824
R10723 gnd.n3105 gnd.n1884 7.64824
R10724 gnd.n3230 gnd.n3229 7.64824
R10725 gnd.n3229 gnd.t27 7.64824
R10726 gnd.n3277 gnd.n1792 7.64824
R10727 gnd.n4422 gnd.n4421 7.53171
R10728 gnd.n4886 gnd.t189 7.32958
R10729 gnd.t249 gnd.n2095 7.32958
R10730 gnd.n2730 gnd.t200 7.32958
R10731 gnd.t124 gnd.n3605 7.32958
R10732 gnd.n3661 gnd.t223 7.32958
R10733 gnd.n1467 gnd.n1466 7.30353
R10734 gnd.n1667 gnd.n1666 7.30353
R10735 gnd.n4846 gnd.n4565 7.01093
R10736 gnd.n4568 gnd.n4566 7.01093
R10737 gnd.n4856 gnd.n4855 7.01093
R10738 gnd.n4867 gnd.n4549 7.01093
R10739 gnd.n4866 gnd.n4552 7.01093
R10740 gnd.n4877 gnd.n4540 7.01093
R10741 gnd.n4543 gnd.n4541 7.01093
R10742 gnd.n4887 gnd.n4886 7.01093
R10743 gnd.n4897 gnd.n4521 7.01093
R10744 gnd.n4896 gnd.n4524 7.01093
R10745 gnd.n4905 gnd.n4515 7.01093
R10746 gnd.n4917 gnd.n4505 7.01093
R10747 gnd.n4927 gnd.n4490 7.01093
R10748 gnd.n4943 gnd.n4942 7.01093
R10749 gnd.n4492 gnd.n4429 7.01093
R10750 gnd.n4997 gnd.n4430 7.01093
R10751 gnd.n4991 gnd.n4990 7.01093
R10752 gnd.n4479 gnd.n4441 7.01093
R10753 gnd.n4983 gnd.n4452 7.01093
R10754 gnd.n4470 gnd.n4465 7.01093
R10755 gnd.n4977 gnd.n4976 7.01093
R10756 gnd.n5023 gnd.n4368 7.01093
R10757 gnd.n5022 gnd.n5021 7.01093
R10758 gnd.n5034 gnd.n5033 7.01093
R10759 gnd.n4361 gnd.n4353 7.01093
R10760 gnd.n5063 gnd.n4341 7.01093
R10761 gnd.n5062 gnd.n4344 7.01093
R10762 gnd.n5073 gnd.n4333 7.01093
R10763 gnd.n4334 gnd.n4322 7.01093
R10764 gnd.n5084 gnd.n4323 7.01093
R10765 gnd.n5108 gnd.n4314 7.01093
R10766 gnd.n5107 gnd.n4305 7.01093
R10767 gnd.n5130 gnd.n5129 7.01093
R10768 gnd.n5148 gnd.n4286 7.01093
R10769 gnd.n5147 gnd.n4289 7.01093
R10770 gnd.n5158 gnd.n4278 7.01093
R10771 gnd.n4279 gnd.n4266 7.01093
R10772 gnd.n5169 gnd.n4267 7.01093
R10773 gnd.n5196 gnd.n4251 7.01093
R10774 gnd.n5208 gnd.n5207 7.01093
R10775 gnd.n5190 gnd.n4244 7.01093
R10776 gnd.n5219 gnd.n5218 7.01093
R10777 gnd.n5491 gnd.n4232 7.01093
R10778 gnd.n5490 gnd.n4235 7.01093
R10779 gnd.n5503 gnd.n4224 7.01093
R10780 gnd.n4225 gnd.n4217 7.01093
R10781 gnd.n5513 gnd.n1008 7.01093
R10782 gnd.n2901 gnd.t120 7.01093
R10783 gnd.n2953 gnd.n2952 7.01093
R10784 gnd.n3002 gnd.n1940 7.01093
R10785 gnd.n3126 gnd.n3125 7.01093
R10786 gnd.n3154 gnd.n3153 7.01093
R10787 gnd.n3301 gnd.n3300 7.01093
R10788 gnd.n3327 gnd.n1754 7.01093
R10789 gnd.n3348 gnd.t26 7.01093
R10790 gnd.n4524 gnd.t179 6.69227
R10791 gnd.n4344 gnd.t151 6.69227
R10792 gnd.n5197 gnd.t105 6.69227
R10793 gnd.t185 gnd.n1978 6.69227
R10794 gnd.n3363 gnd.t149 6.69227
R10795 gnd.n3474 gnd.n3473 6.5566
R10796 gnd.n2815 gnd.n2814 6.5566
R10797 gnd.n3790 gnd.n3786 6.5566
R10798 gnd.n3489 gnd.n3488 6.5566
R10799 gnd.n2875 gnd.n1471 6.37362
R10800 gnd.n2925 gnd.n2924 6.37362
R10801 gnd.n2900 gnd.t299 6.37362
R10802 gnd.n3011 gnd.t97 6.37362
R10803 gnd.n3049 gnd.n3048 6.37362
R10804 gnd.n3106 gnd.t79 6.37362
R10805 gnd.t27 gnd.n3228 6.37362
R10806 gnd.n3267 gnd.n3266 6.37362
R10807 gnd.n3314 gnd.t6 6.37362
R10808 gnd.n3373 gnd.n3372 6.37362
R10809 gnd.n3544 gnd.n3543 6.37362
R10810 gnd.n2550 gnd.n2191 6.20656
R10811 gnd.n449 gnd.n443 6.20656
R10812 gnd.t84 gnd.n4953 6.05496
R10813 gnd.n4954 gnd.t182 6.05496
R10814 gnd.t2 gnd.n4368 6.05496
R10815 gnd.t64 gnd.n5118 6.05496
R10816 gnd.n3125 gnd.t126 6.05496
R10817 gnd.n3153 gnd.t102 6.05496
R10818 gnd.n5476 gnd.n5446 5.81868
R10819 gnd.n5444 gnd.n5414 5.81868
R10820 gnd.n5412 gnd.n5382 5.81868
R10821 gnd.n5381 gnd.n5351 5.81868
R10822 gnd.n5349 gnd.n5319 5.81868
R10823 gnd.n5317 gnd.n5287 5.81868
R10824 gnd.n5285 gnd.n5255 5.81868
R10825 gnd.n5254 gnd.n5224 5.81868
R10826 gnd.t290 gnd.n2888 5.73631
R10827 gnd.t120 gnd.n1969 5.73631
R10828 gnd.n2977 gnd.n1954 5.73631
R10829 gnd.n2958 gnd.n2957 5.73631
R10830 gnd.n1872 gnd.n1859 5.73631
R10831 gnd.n3130 gnd.n1861 5.73631
R10832 gnd.n3291 gnd.n3290 5.73631
R10833 gnd.n3305 gnd.n1770 5.73631
R10834 gnd.n3326 gnd.t26 5.73631
R10835 gnd.n3544 gnd.t209 5.73631
R10836 gnd.n1696 gnd.n351 5.62001
R10837 gnd.n3852 gnd.n1409 5.62001
R10838 gnd.n3852 gnd.n1410 5.62001
R10839 gnd.n3483 gnd.n351 5.62001
R10840 gnd.n4705 gnd.n4700 5.4308
R10841 gnd.n5521 gnd.n4210 5.4308
R10842 gnd.n5021 gnd.t188 5.41765
R10843 gnd.t63 gnd.n5044 5.41765
R10844 gnd.t92 gnd.n4298 5.41765
R10845 gnd.n5605 gnd.n1008 5.41765
R10846 gnd.n3849 gnd.n1413 5.41765
R10847 gnd.t108 gnd.n1946 5.41765
R10848 gnd.t129 gnd.n1779 5.41765
R10849 gnd.n2876 gnd.t212 5.09899
R10850 gnd.n2889 gnd.n1474 5.09899
R10851 gnd.n2889 gnd.t290 5.09899
R10852 gnd.n2918 gnd.n2917 5.09899
R10853 gnd.n3075 gnd.n1915 5.09899
R10854 gnd.n3088 gnd.n3087 5.09899
R10855 gnd.n3248 gnd.n1820 5.09899
R10856 gnd.n3260 gnd.n3259 5.09899
R10857 gnd.t243 gnd.n3380 5.09899
R10858 gnd.n3405 gnd.t266 5.09899
R10859 gnd.n3388 gnd.n1723 5.09899
R10860 gnd.n5474 gnd.n5473 5.04292
R10861 gnd.n5442 gnd.n5441 5.04292
R10862 gnd.n5410 gnd.n5409 5.04292
R10863 gnd.n5379 gnd.n5378 5.04292
R10864 gnd.n5347 gnd.n5346 5.04292
R10865 gnd.n5315 gnd.n5314 5.04292
R10866 gnd.n5283 gnd.n5282 5.04292
R10867 gnd.n5252 gnd.n5251 5.04292
R10868 gnd.n4984 gnd.t183 4.78034
R10869 gnd.n4323 gnd.t176 4.78034
R10870 gnd.n2760 gnd.t171 4.78034
R10871 gnd.n2958 gnd.t108 4.78034
R10872 gnd.n3290 gnd.t129 4.78034
R10873 gnd.n1672 gnd.t281 4.78034
R10874 gnd.n3574 gnd.t155 4.78034
R10875 gnd.n4426 gnd.n4423 4.74817
R10876 gnd.n4476 gnd.n4374 4.74817
R10877 gnd.n4463 gnd.n4373 4.74817
R10878 gnd.n4372 gnd.n4371 4.74817
R10879 gnd.n4472 gnd.n4423 4.74817
R10880 gnd.n4473 gnd.n4374 4.74817
R10881 gnd.n4475 gnd.n4373 4.74817
R10882 gnd.n4462 gnd.n4372 4.74817
R10883 gnd.n4421 gnd.n4420 4.74296
R10884 gnd.n66 gnd.n65 4.74296
R10885 gnd.n4397 gnd.n4396 4.7074
R10886 gnd.n4409 gnd.n4408 4.7074
R10887 gnd.n42 gnd.n41 4.7074
R10888 gnd.n54 gnd.n53 4.7074
R10889 gnd.n4421 gnd.n4409 4.65959
R10890 gnd.n66 gnd.n54 4.65959
R10891 gnd.n6481 gnd.n353 4.6132
R10892 gnd.n3853 gnd.n1408 4.6132
R10893 gnd.t212 gnd.n2875 4.46168
R10894 gnd.n2966 gnd.n2965 4.46168
R10895 gnd.n2975 gnd.t18 4.46168
R10896 gnd.n2996 gnd.n2995 4.46168
R10897 gnd.n3139 gnd.n3137 4.46168
R10898 gnd.n3161 gnd.n3160 4.46168
R10899 gnd.n3313 gnd.n3312 4.46168
R10900 gnd.n3322 gnd.t147 4.46168
R10901 gnd.n3335 gnd.n3333 4.46168
R10902 gnd.n1663 gnd.n1650 4.46111
R10903 gnd.n5459 gnd.n5455 4.38594
R10904 gnd.n5427 gnd.n5423 4.38594
R10905 gnd.n5395 gnd.n5391 4.38594
R10906 gnd.n5364 gnd.n5360 4.38594
R10907 gnd.n5332 gnd.n5328 4.38594
R10908 gnd.n5300 gnd.n5296 4.38594
R10909 gnd.n5268 gnd.n5264 4.38594
R10910 gnd.n5237 gnd.n5233 4.38594
R10911 gnd.n5470 gnd.n5448 4.26717
R10912 gnd.n5438 gnd.n5416 4.26717
R10913 gnd.n5406 gnd.n5384 4.26717
R10914 gnd.n5375 gnd.n5353 4.26717
R10915 gnd.n5343 gnd.n5321 4.26717
R10916 gnd.n5311 gnd.n5289 4.26717
R10917 gnd.n5279 gnd.n5257 4.26717
R10918 gnd.n5248 gnd.n5226 4.26717
R10919 gnd.n4928 gnd.t181 4.14303
R10920 gnd.n5158 gnd.t178 4.14303
R10921 gnd.n5478 gnd.n5477 4.08274
R10922 gnd.n3473 gnd.n3472 4.05904
R10923 gnd.n2816 gnd.n2815 4.05904
R10924 gnd.n3793 gnd.n3786 4.05904
R10925 gnd.n3490 gnd.n3489 4.05904
R10926 gnd.n19 gnd.n9 3.99943
R10927 gnd.n3903 gnd.n1350 3.82437
R10928 gnd.n2909 gnd.n2908 3.82437
R10929 gnd.n3056 gnd.t13 3.82437
R10930 gnd.n3067 gnd.n3066 3.82437
R10931 gnd.n3038 gnd.n3037 3.82437
R10932 gnd.n3240 gnd.n3239 3.82437
R10933 gnd.n3211 gnd.n3210 3.82437
R10934 gnd.t96 gnd.n3277 3.82437
R10935 gnd.n3397 gnd.n3396 3.82437
R10936 gnd.n6530 gnd.n284 3.82437
R10937 gnd.n5001 gnd.n4422 3.81325
R10938 gnd.n4409 gnd.n4397 3.72967
R10939 gnd.n54 gnd.n42 3.72967
R10940 gnd.n5478 gnd.n5350 3.70378
R10941 gnd.n19 gnd.n18 3.60163
R10942 gnd.n2078 gnd.t82 3.50571
R10943 gnd.t59 gnd.n3624 3.50571
R10944 gnd.n5469 gnd.n5450 3.49141
R10945 gnd.n5437 gnd.n5418 3.49141
R10946 gnd.n5405 gnd.n5386 3.49141
R10947 gnd.n5374 gnd.n5355 3.49141
R10948 gnd.n5342 gnd.n5323 3.49141
R10949 gnd.n5310 gnd.n5291 3.49141
R10950 gnd.n5278 gnd.n5259 3.49141
R10951 gnd.n5247 gnd.n5228 3.49141
R10952 gnd.n7004 gnd.n7001 3.29747
R10953 gnd.n7005 gnd.n7004 3.29747
R10954 gnd.n6499 gnd.n6498 3.29747
R10955 gnd.n6498 gnd.n6497 3.29747
R10956 gnd.n4122 gnd.n4121 3.29747
R10957 gnd.n4121 gnd.n4120 3.29747
R10958 gnd.n3871 gnd.n3870 3.29747
R10959 gnd.n3870 gnd.n3869 3.29747
R10960 gnd.n3929 gnd.n1302 3.18706
R10961 gnd.n2531 gnd.n1309 3.18706
R10962 gnd.n3923 gnd.n1312 3.18706
R10963 gnd.n2543 gnd.n1320 3.18706
R10964 gnd.n3917 gnd.n1323 3.18706
R10965 gnd.n2566 gnd.n2565 3.18706
R10966 gnd.n3911 gnd.n1332 3.18706
R10967 gnd.n2598 gnd.n2597 3.18706
R10968 gnd.n2901 gnd.n2900 3.18706
R10969 gnd.t327 gnd.n3094 3.18706
R10970 gnd.n3030 gnd.n3029 3.18706
R10971 gnd.n3174 gnd.n3173 3.18706
R10972 gnd.n3222 gnd.t121 3.18706
R10973 gnd.n3348 gnd.n3347 3.18706
R10974 gnd.n6330 gnd.n6329 3.18706
R10975 gnd.n6540 gnd.n274 3.18706
R10976 gnd.n6323 gnd.n6322 3.18706
R10977 gnd.n6549 gnd.n267 3.18706
R10978 gnd.n6565 gnd.n255 3.18706
R10979 gnd.n6553 gnd.n258 3.18706
R10980 gnd.n6575 gnd.n246 3.18706
R10981 gnd.n516 gnd.n239 3.18706
R10982 gnd.n4507 gnd.t181 2.8684
R10983 gnd.n2888 gnd.t202 2.8684
R10984 gnd.t299 gnd.t185 2.8684
R10985 gnd.n3387 gnd.t192 2.8684
R10986 gnd.n4410 gnd.t163 2.82907
R10987 gnd.n4410 gnd.t194 2.82907
R10988 gnd.n4412 gnd.t144 2.82907
R10989 gnd.n4412 gnd.t141 2.82907
R10990 gnd.n4414 gnd.t142 2.82907
R10991 gnd.n4414 gnd.t199 2.82907
R10992 gnd.n4416 gnd.t333 2.82907
R10993 gnd.n4416 gnd.t164 2.82907
R10994 gnd.n4418 gnd.t161 2.82907
R10995 gnd.n4418 gnd.t47 2.82907
R10996 gnd.n4375 gnd.t43 2.82907
R10997 gnd.n4375 gnd.t170 2.82907
R10998 gnd.n4377 gnd.t132 2.82907
R10999 gnd.n4377 gnd.t118 2.82907
R11000 gnd.n4379 gnd.t98 2.82907
R11001 gnd.n4379 gnd.t34 2.82907
R11002 gnd.n4381 gnd.t88 2.82907
R11003 gnd.n4381 gnd.t131 2.82907
R11004 gnd.n4383 gnd.t166 2.82907
R11005 gnd.n4383 gnd.t86 2.82907
R11006 gnd.n4386 gnd.t104 2.82907
R11007 gnd.n4386 gnd.t135 2.82907
R11008 gnd.n4388 gnd.t45 2.82907
R11009 gnd.n4388 gnd.t165 2.82907
R11010 gnd.n4390 gnd.t17 2.82907
R11011 gnd.n4390 gnd.t325 2.82907
R11012 gnd.n4392 gnd.t331 2.82907
R11013 gnd.n4392 gnd.t31 2.82907
R11014 gnd.n4394 gnd.t5 2.82907
R11015 gnd.n4394 gnd.t330 2.82907
R11016 gnd.n4398 gnd.t134 2.82907
R11017 gnd.n4398 gnd.t71 2.82907
R11018 gnd.n4400 gnd.t190 2.82907
R11019 gnd.n4400 gnd.t324 2.82907
R11020 gnd.n4402 gnd.t329 2.82907
R11021 gnd.n4402 gnd.t33 2.82907
R11022 gnd.n4404 gnd.t111 2.82907
R11023 gnd.n4404 gnd.t160 2.82907
R11024 gnd.n4406 gnd.t49 2.82907
R11025 gnd.n4406 gnd.t174 2.82907
R11026 gnd.n63 gnd.t328 2.82907
R11027 gnd.n63 gnd.t191 2.82907
R11028 gnd.n61 gnd.t169 2.82907
R11029 gnd.n61 gnd.t24 2.82907
R11030 gnd.n59 gnd.t78 2.82907
R11031 gnd.n59 gnd.t8 2.82907
R11032 gnd.n57 gnd.t154 2.82907
R11033 gnd.n57 gnd.t143 2.82907
R11034 gnd.n55 gnd.t136 2.82907
R11035 gnd.n55 gnd.t22 2.82907
R11036 gnd.n28 gnd.t323 2.82907
R11037 gnd.n28 gnd.t54 2.82907
R11038 gnd.n26 gnd.t68 2.82907
R11039 gnd.n26 gnd.t81 2.82907
R11040 gnd.n24 gnd.t101 2.82907
R11041 gnd.n24 gnd.t119 2.82907
R11042 gnd.n22 gnd.t112 2.82907
R11043 gnd.n22 gnd.t69 2.82907
R11044 gnd.n20 gnd.t332 2.82907
R11045 gnd.n20 gnd.t72 2.82907
R11046 gnd.n39 gnd.t107 2.82907
R11047 gnd.n39 gnd.t10 2.82907
R11048 gnd.n37 gnd.t146 2.82907
R11049 gnd.n37 gnd.t94 2.82907
R11050 gnd.n35 gnd.t1 2.82907
R11051 gnd.n35 gnd.t74 2.82907
R11052 gnd.n33 gnd.t56 2.82907
R11053 gnd.n33 gnd.t53 2.82907
R11054 gnd.n31 gnd.t197 2.82907
R11055 gnd.n31 gnd.t21 2.82907
R11056 gnd.n51 gnd.t148 2.82907
R11057 gnd.n51 gnd.t90 2.82907
R11058 gnd.n49 gnd.t168 2.82907
R11059 gnd.n49 gnd.t55 2.82907
R11060 gnd.n47 gnd.t198 2.82907
R11061 gnd.n47 gnd.t145 2.82907
R11062 gnd.n45 gnd.t37 2.82907
R11063 gnd.n45 gnd.t89 2.82907
R11064 gnd.n43 gnd.t58 2.82907
R11065 gnd.n43 gnd.t167 2.82907
R11066 gnd.n5466 gnd.n5465 2.71565
R11067 gnd.n5434 gnd.n5433 2.71565
R11068 gnd.n5402 gnd.n5401 2.71565
R11069 gnd.n5371 gnd.n5370 2.71565
R11070 gnd.n5339 gnd.n5338 2.71565
R11071 gnd.n5307 gnd.n5306 2.71565
R11072 gnd.n5275 gnd.n5274 2.71565
R11073 gnd.n5244 gnd.n5243 2.71565
R11074 gnd.n2936 gnd.t246 2.54975
R11075 gnd.n2942 gnd.n1978 2.54975
R11076 gnd.n3020 gnd.n3019 2.54975
R11077 gnd.n3112 gnd.n1886 2.54975
R11078 gnd.n3029 gnd.t77 2.54975
R11079 gnd.n3140 gnd.t75 2.54975
R11080 gnd.n3181 gnd.t153 2.54975
R11081 gnd.n3173 gnd.t80 2.54975
R11082 gnd.n3190 gnd.n3189 2.54975
R11083 gnd.n3284 gnd.n1794 2.54975
R11084 gnd.n3364 gnd.n3363 2.54975
R11085 gnd.n3381 gnd.t243 2.54975
R11086 gnd.n5001 gnd.n4423 2.27742
R11087 gnd.n5001 gnd.n4374 2.27742
R11088 gnd.n5001 gnd.n4373 2.27742
R11089 gnd.n5001 gnd.n4372 2.27742
R11090 gnd.n4855 gnd.t262 2.23109
R11091 gnd.n4478 gnd.t183 2.23109
R11092 gnd.n3095 gnd.t14 2.23109
R11093 gnd.t114 gnd.n3221 2.23109
R11094 gnd.n5462 gnd.n5452 1.93989
R11095 gnd.n5430 gnd.n5420 1.93989
R11096 gnd.n5398 gnd.n5388 1.93989
R11097 gnd.n5367 gnd.n5357 1.93989
R11098 gnd.n5335 gnd.n5325 1.93989
R11099 gnd.n5303 gnd.n5293 1.93989
R11100 gnd.n5271 gnd.n5261 1.93989
R11101 gnd.n5240 gnd.n5230 1.93989
R11102 gnd.n2936 gnd.n1982 1.91244
R11103 gnd.n3004 gnd.t19 1.91244
R11104 gnd.t48 gnd.n1905 1.91244
R11105 gnd.n3106 gnd.n1891 1.91244
R11106 gnd.n3228 gnd.n1826 1.91244
R11107 gnd.n1819 gnd.t159 1.91244
R11108 gnd.n3200 gnd.t35 1.91244
R11109 gnd.n3379 gnd.n1738 1.91244
R11110 gnd.t139 gnd.n4866 1.59378
R11111 gnd.n5045 gnd.t63 1.59378
R11112 gnd.n4307 gnd.t92 1.59378
R11113 gnd.t122 gnd.n1921 1.59378
R11114 gnd.n3209 gnd.t11 1.59378
R11115 gnd.n2967 gnd.n1962 1.27512
R11116 gnd.n3011 gnd.n3010 1.27512
R11117 gnd.t19 gnd.n1933 1.27512
R11118 gnd.n3140 gnd.n1867 1.27512
R11119 gnd.n3181 gnd.n3180 1.27512
R11120 gnd.t35 gnd.n3199 1.27512
R11121 gnd.n3314 gnd.n1776 1.27512
R11122 gnd.n3355 gnd.n3354 1.27512
R11123 gnd.n4708 gnd.n4700 1.16414
R11124 gnd.n5524 gnd.n4210 1.16414
R11125 gnd.n5461 gnd.n5454 1.16414
R11126 gnd.n5429 gnd.n5422 1.16414
R11127 gnd.n5397 gnd.n5390 1.16414
R11128 gnd.n5366 gnd.n5359 1.16414
R11129 gnd.n5334 gnd.n5327 1.16414
R11130 gnd.n5302 gnd.n5295 1.16414
R11131 gnd.n5270 gnd.n5263 1.16414
R11132 gnd.n5239 gnd.n5232 1.16414
R11133 gnd.n6481 gnd.n6480 0.970197
R11134 gnd.n3853 gnd.n1406 0.970197
R11135 gnd.n5445 gnd.n5413 0.962709
R11136 gnd.n5477 gnd.n5445 0.962709
R11137 gnd.n5318 gnd.n5286 0.962709
R11138 gnd.n5350 gnd.n5318 0.962709
R11139 gnd.n4954 gnd.t84 0.956468
R11140 gnd.n5119 gnd.t64 0.956468
R11141 gnd.n4007 gnd.t4 0.956468
R11142 gnd.n3935 gnd.t70 0.956468
R11143 gnd.t195 gnd.n2002 0.956468
R11144 gnd.t14 gnd.t327 0.956468
R11145 gnd.t121 gnd.t114 0.956468
R11146 gnd.n3553 gnd.t61 0.956468
R11147 gnd.n6605 gnd.t57 0.956468
R11148 gnd.n7077 gnd.t9 0.956468
R11149 gnd.n2 gnd.n1 0.672012
R11150 gnd.n3 gnd.n2 0.672012
R11151 gnd.n4 gnd.n3 0.672012
R11152 gnd.n5 gnd.n4 0.672012
R11153 gnd.n6 gnd.n5 0.672012
R11154 gnd.n7 gnd.n6 0.672012
R11155 gnd.n8 gnd.n7 0.672012
R11156 gnd.n9 gnd.n8 0.672012
R11157 gnd.n11 gnd.n10 0.672012
R11158 gnd.n12 gnd.n11 0.672012
R11159 gnd.n13 gnd.n12 0.672012
R11160 gnd.n14 gnd.n13 0.672012
R11161 gnd.n15 gnd.n14 0.672012
R11162 gnd.n16 gnd.n15 0.672012
R11163 gnd.n17 gnd.n16 0.672012
R11164 gnd.n18 gnd.n17 0.672012
R11165 gnd.n3779 gnd.n3778 0.637812
R11166 gnd.n2916 gnd.n2915 0.637812
R11167 gnd.n2925 gnd.t239 0.637812
R11168 gnd.t95 gnd.n2966 0.637812
R11169 gnd.n3049 gnd.t25 0.637812
R11170 gnd.n3077 gnd.n1914 0.637812
R11171 gnd.n3086 gnd.n1899 0.637812
R11172 gnd.n3249 gnd.n1818 0.637812
R11173 gnd.n3258 gnd.n1805 0.637812
R11174 gnd.n3266 gnd.t76 0.637812
R11175 gnd.n3335 gnd.t175 0.637812
R11176 gnd.n3372 gnd.t235 0.637812
R11177 gnd.n3406 gnd.n1731 0.637812
R11178 gnd.n3417 gnd.n3416 0.637812
R11179 gnd.t281 gnd.n1639 0.637812
R11180 gnd gnd.n0 0.624033
R11181 gnd.n4420 gnd.n4419 0.573776
R11182 gnd.n4419 gnd.n4417 0.573776
R11183 gnd.n4417 gnd.n4415 0.573776
R11184 gnd.n4415 gnd.n4413 0.573776
R11185 gnd.n4413 gnd.n4411 0.573776
R11186 gnd.n4385 gnd.n4384 0.573776
R11187 gnd.n4384 gnd.n4382 0.573776
R11188 gnd.n4382 gnd.n4380 0.573776
R11189 gnd.n4380 gnd.n4378 0.573776
R11190 gnd.n4378 gnd.n4376 0.573776
R11191 gnd.n4396 gnd.n4395 0.573776
R11192 gnd.n4395 gnd.n4393 0.573776
R11193 gnd.n4393 gnd.n4391 0.573776
R11194 gnd.n4391 gnd.n4389 0.573776
R11195 gnd.n4389 gnd.n4387 0.573776
R11196 gnd.n4408 gnd.n4407 0.573776
R11197 gnd.n4407 gnd.n4405 0.573776
R11198 gnd.n4405 gnd.n4403 0.573776
R11199 gnd.n4403 gnd.n4401 0.573776
R11200 gnd.n4401 gnd.n4399 0.573776
R11201 gnd.n58 gnd.n56 0.573776
R11202 gnd.n60 gnd.n58 0.573776
R11203 gnd.n62 gnd.n60 0.573776
R11204 gnd.n64 gnd.n62 0.573776
R11205 gnd.n65 gnd.n64 0.573776
R11206 gnd.n23 gnd.n21 0.573776
R11207 gnd.n25 gnd.n23 0.573776
R11208 gnd.n27 gnd.n25 0.573776
R11209 gnd.n29 gnd.n27 0.573776
R11210 gnd.n30 gnd.n29 0.573776
R11211 gnd.n34 gnd.n32 0.573776
R11212 gnd.n36 gnd.n34 0.573776
R11213 gnd.n38 gnd.n36 0.573776
R11214 gnd.n40 gnd.n38 0.573776
R11215 gnd.n41 gnd.n40 0.573776
R11216 gnd.n46 gnd.n44 0.573776
R11217 gnd.n48 gnd.n46 0.573776
R11218 gnd.n50 gnd.n48 0.573776
R11219 gnd.n52 gnd.n50 0.573776
R11220 gnd.n53 gnd.n52 0.573776
R11221 gnd.n6833 gnd.n6832 0.532512
R11222 gnd.n2459 gnd.n2458 0.532512
R11223 gnd.n6867 gnd.n6866 0.497451
R11224 gnd.n3907 gnd.n3906 0.497451
R11225 gnd.n6535 gnd.n6534 0.497451
R11226 gnd.n1142 gnd.n1065 0.497451
R11227 gnd.n5181 gnd.n4214 0.486781
R11228 gnd.n4757 gnd.n4756 0.48678
R11229 gnd.n5498 gnd.n4168 0.480683
R11230 gnd.n4841 gnd.n4840 0.480683
R11231 gnd.n7114 gnd.n7113 0.4705
R11232 gnd.n6359 gnd.n6358 0.451719
R11233 gnd.n2548 gnd.n2099 0.451719
R11234 gnd.n2665 gnd.n2664 0.451719
R11235 gnd.n6352 gnd.n6351 0.451719
R11236 gnd.n5777 gnd.n838 0.416659
R11237 gnd.n6098 gnd.n6097 0.416659
R11238 gnd.n6312 gnd.n6311 0.416659
R11239 gnd.n2305 gnd.n2304 0.416659
R11240 gnd.n2606 gnd.n2191 0.388379
R11241 gnd.n5458 gnd.n5457 0.388379
R11242 gnd.n5426 gnd.n5425 0.388379
R11243 gnd.n5394 gnd.n5393 0.388379
R11244 gnd.n5363 gnd.n5362 0.388379
R11245 gnd.n5331 gnd.n5330 0.388379
R11246 gnd.n5299 gnd.n5298 0.388379
R11247 gnd.n5267 gnd.n5266 0.388379
R11248 gnd.n5236 gnd.n5235 0.388379
R11249 gnd.n6373 gnd.n443 0.388379
R11250 gnd.n7114 gnd.n19 0.374463
R11251 gnd gnd.n7114 0.367492
R11252 gnd.n4269 gnd.t105 0.319156
R11253 gnd.n3983 gnd.t30 0.319156
R11254 gnd.n3959 gnd.t44 0.319156
R11255 gnd.n3055 gnd.t122 0.319156
R11256 gnd.n3278 gnd.t11 0.319156
R11257 gnd.n6652 gnd.t52 0.319156
R11258 gnd.n7101 gnd.t67 0.319156
R11259 gnd.n4675 gnd.n4653 0.311721
R11260 gnd.n2560 gnd.n2559 0.302329
R11261 gnd.n6360 gnd.n271 0.302329
R11262 gnd.n7048 gnd.n6718 0.293183
R11263 gnd.n4038 gnd.n1129 0.293183
R11264 gnd.n5569 gnd.n5568 0.268793
R11265 gnd.n6419 gnd.n6418 0.258122
R11266 gnd.n7048 gnd.n7047 0.258122
R11267 gnd.n2293 gnd.n2134 0.258122
R11268 gnd.n4039 gnd.n4038 0.258122
R11269 gnd.n5568 gnd.n5567 0.241354
R11270 gnd.n353 gnd.n350 0.229039
R11271 gnd.n354 gnd.n353 0.229039
R11272 gnd.n1408 gnd.n1405 0.229039
R11273 gnd.n2221 gnd.n1408 0.229039
R11274 gnd.n4829 gnd.n4628 0.206293
R11275 gnd.n5475 gnd.n5447 0.155672
R11276 gnd.n5468 gnd.n5447 0.155672
R11277 gnd.n5468 gnd.n5467 0.155672
R11278 gnd.n5467 gnd.n5451 0.155672
R11279 gnd.n5460 gnd.n5451 0.155672
R11280 gnd.n5460 gnd.n5459 0.155672
R11281 gnd.n5443 gnd.n5415 0.155672
R11282 gnd.n5436 gnd.n5415 0.155672
R11283 gnd.n5436 gnd.n5435 0.155672
R11284 gnd.n5435 gnd.n5419 0.155672
R11285 gnd.n5428 gnd.n5419 0.155672
R11286 gnd.n5428 gnd.n5427 0.155672
R11287 gnd.n5411 gnd.n5383 0.155672
R11288 gnd.n5404 gnd.n5383 0.155672
R11289 gnd.n5404 gnd.n5403 0.155672
R11290 gnd.n5403 gnd.n5387 0.155672
R11291 gnd.n5396 gnd.n5387 0.155672
R11292 gnd.n5396 gnd.n5395 0.155672
R11293 gnd.n5380 gnd.n5352 0.155672
R11294 gnd.n5373 gnd.n5352 0.155672
R11295 gnd.n5373 gnd.n5372 0.155672
R11296 gnd.n5372 gnd.n5356 0.155672
R11297 gnd.n5365 gnd.n5356 0.155672
R11298 gnd.n5365 gnd.n5364 0.155672
R11299 gnd.n5348 gnd.n5320 0.155672
R11300 gnd.n5341 gnd.n5320 0.155672
R11301 gnd.n5341 gnd.n5340 0.155672
R11302 gnd.n5340 gnd.n5324 0.155672
R11303 gnd.n5333 gnd.n5324 0.155672
R11304 gnd.n5333 gnd.n5332 0.155672
R11305 gnd.n5316 gnd.n5288 0.155672
R11306 gnd.n5309 gnd.n5288 0.155672
R11307 gnd.n5309 gnd.n5308 0.155672
R11308 gnd.n5308 gnd.n5292 0.155672
R11309 gnd.n5301 gnd.n5292 0.155672
R11310 gnd.n5301 gnd.n5300 0.155672
R11311 gnd.n5284 gnd.n5256 0.155672
R11312 gnd.n5277 gnd.n5256 0.155672
R11313 gnd.n5277 gnd.n5276 0.155672
R11314 gnd.n5276 gnd.n5260 0.155672
R11315 gnd.n5269 gnd.n5260 0.155672
R11316 gnd.n5269 gnd.n5268 0.155672
R11317 gnd.n5253 gnd.n5225 0.155672
R11318 gnd.n5246 gnd.n5225 0.155672
R11319 gnd.n5246 gnd.n5245 0.155672
R11320 gnd.n5245 gnd.n5229 0.155672
R11321 gnd.n5238 gnd.n5229 0.155672
R11322 gnd.n5238 gnd.n5237 0.155672
R11323 gnd.n6534 gnd.n281 0.152939
R11324 gnd.n325 gnd.n281 0.152939
R11325 gnd.n326 gnd.n325 0.152939
R11326 gnd.n327 gnd.n326 0.152939
R11327 gnd.n328 gnd.n327 0.152939
R11328 gnd.n329 gnd.n328 0.152939
R11329 gnd.n330 gnd.n329 0.152939
R11330 gnd.n331 gnd.n330 0.152939
R11331 gnd.n332 gnd.n331 0.152939
R11332 gnd.n333 gnd.n332 0.152939
R11333 gnd.n334 gnd.n333 0.152939
R11334 gnd.n335 gnd.n334 0.152939
R11335 gnd.n336 gnd.n335 0.152939
R11336 gnd.n337 gnd.n336 0.152939
R11337 gnd.n338 gnd.n337 0.152939
R11338 gnd.n339 gnd.n338 0.152939
R11339 gnd.n340 gnd.n339 0.152939
R11340 gnd.n343 gnd.n340 0.152939
R11341 gnd.n344 gnd.n343 0.152939
R11342 gnd.n345 gnd.n344 0.152939
R11343 gnd.n346 gnd.n345 0.152939
R11344 gnd.n347 gnd.n346 0.152939
R11345 gnd.n348 gnd.n347 0.152939
R11346 gnd.n349 gnd.n348 0.152939
R11347 gnd.n350 gnd.n349 0.152939
R11348 gnd.n355 gnd.n354 0.152939
R11349 gnd.n356 gnd.n355 0.152939
R11350 gnd.n357 gnd.n356 0.152939
R11351 gnd.n358 gnd.n357 0.152939
R11352 gnd.n359 gnd.n358 0.152939
R11353 gnd.n360 gnd.n359 0.152939
R11354 gnd.n361 gnd.n360 0.152939
R11355 gnd.n362 gnd.n361 0.152939
R11356 gnd.n363 gnd.n362 0.152939
R11357 gnd.n366 gnd.n363 0.152939
R11358 gnd.n367 gnd.n366 0.152939
R11359 gnd.n368 gnd.n367 0.152939
R11360 gnd.n369 gnd.n368 0.152939
R11361 gnd.n370 gnd.n369 0.152939
R11362 gnd.n371 gnd.n370 0.152939
R11363 gnd.n372 gnd.n371 0.152939
R11364 gnd.n373 gnd.n372 0.152939
R11365 gnd.n374 gnd.n373 0.152939
R11366 gnd.n375 gnd.n374 0.152939
R11367 gnd.n376 gnd.n375 0.152939
R11368 gnd.n377 gnd.n376 0.152939
R11369 gnd.n378 gnd.n377 0.152939
R11370 gnd.n379 gnd.n378 0.152939
R11371 gnd.n380 gnd.n379 0.152939
R11372 gnd.n381 gnd.n380 0.152939
R11373 gnd.n382 gnd.n381 0.152939
R11374 gnd.n383 gnd.n382 0.152939
R11375 gnd.n384 gnd.n383 0.152939
R11376 gnd.n6420 gnd.n384 0.152939
R11377 gnd.n6420 gnd.n6419 0.152939
R11378 gnd.n6537 gnd.n6535 0.152939
R11379 gnd.n6537 gnd.n6536 0.152939
R11380 gnd.n6536 gnd.n252 0.152939
R11381 gnd.n6568 gnd.n252 0.152939
R11382 gnd.n6569 gnd.n6568 0.152939
R11383 gnd.n6570 gnd.n6569 0.152939
R11384 gnd.n6571 gnd.n6570 0.152939
R11385 gnd.n6571 gnd.n226 0.152939
R11386 gnd.n6608 gnd.n226 0.152939
R11387 gnd.n6609 gnd.n6608 0.152939
R11388 gnd.n6610 gnd.n6609 0.152939
R11389 gnd.n6610 gnd.n206 0.152939
R11390 gnd.n6632 gnd.n206 0.152939
R11391 gnd.n6633 gnd.n6632 0.152939
R11392 gnd.n6634 gnd.n6633 0.152939
R11393 gnd.n6635 gnd.n6634 0.152939
R11394 gnd.n99 gnd.n98 0.152939
R11395 gnd.n100 gnd.n99 0.152939
R11396 gnd.n101 gnd.n100 0.152939
R11397 gnd.n118 gnd.n101 0.152939
R11398 gnd.n119 gnd.n118 0.152939
R11399 gnd.n120 gnd.n119 0.152939
R11400 gnd.n121 gnd.n120 0.152939
R11401 gnd.n136 gnd.n121 0.152939
R11402 gnd.n137 gnd.n136 0.152939
R11403 gnd.n138 gnd.n137 0.152939
R11404 gnd.n139 gnd.n138 0.152939
R11405 gnd.n156 gnd.n139 0.152939
R11406 gnd.n157 gnd.n156 0.152939
R11407 gnd.n158 gnd.n157 0.152939
R11408 gnd.n159 gnd.n158 0.152939
R11409 gnd.n6866 gnd.n159 0.152939
R11410 gnd.n7111 gnd.n69 0.152939
R11411 gnd.n6796 gnd.n69 0.152939
R11412 gnd.n6797 gnd.n6796 0.152939
R11413 gnd.n6801 gnd.n6797 0.152939
R11414 gnd.n6802 gnd.n6801 0.152939
R11415 gnd.n6803 gnd.n6802 0.152939
R11416 gnd.n6803 gnd.n6794 0.152939
R11417 gnd.n6809 gnd.n6794 0.152939
R11418 gnd.n6810 gnd.n6809 0.152939
R11419 gnd.n6811 gnd.n6810 0.152939
R11420 gnd.n6811 gnd.n6792 0.152939
R11421 gnd.n6817 gnd.n6792 0.152939
R11422 gnd.n6818 gnd.n6817 0.152939
R11423 gnd.n6819 gnd.n6818 0.152939
R11424 gnd.n6819 gnd.n6790 0.152939
R11425 gnd.n6825 gnd.n6790 0.152939
R11426 gnd.n6826 gnd.n6825 0.152939
R11427 gnd.n6827 gnd.n6826 0.152939
R11428 gnd.n6827 gnd.n6788 0.152939
R11429 gnd.n6832 gnd.n6788 0.152939
R11430 gnd.n6748 gnd.n6718 0.152939
R11431 gnd.n6749 gnd.n6748 0.152939
R11432 gnd.n6749 gnd.n6744 0.152939
R11433 gnd.n6757 gnd.n6744 0.152939
R11434 gnd.n6758 gnd.n6757 0.152939
R11435 gnd.n6759 gnd.n6758 0.152939
R11436 gnd.n6759 gnd.n6742 0.152939
R11437 gnd.n6767 gnd.n6742 0.152939
R11438 gnd.n6768 gnd.n6767 0.152939
R11439 gnd.n6769 gnd.n6768 0.152939
R11440 gnd.n6769 gnd.n6740 0.152939
R11441 gnd.n6777 gnd.n6740 0.152939
R11442 gnd.n6778 gnd.n6777 0.152939
R11443 gnd.n6779 gnd.n6778 0.152939
R11444 gnd.n6779 gnd.n6738 0.152939
R11445 gnd.n6786 gnd.n6738 0.152939
R11446 gnd.n6787 gnd.n6786 0.152939
R11447 gnd.n6833 gnd.n6787 0.152939
R11448 gnd.n7038 gnd.n6867 0.152939
R11449 gnd.n7038 gnd.n7037 0.152939
R11450 gnd.n7037 gnd.n7036 0.152939
R11451 gnd.n7036 gnd.n6869 0.152939
R11452 gnd.n6870 gnd.n6869 0.152939
R11453 gnd.n6871 gnd.n6870 0.152939
R11454 gnd.n6872 gnd.n6871 0.152939
R11455 gnd.n6873 gnd.n6872 0.152939
R11456 gnd.n6874 gnd.n6873 0.152939
R11457 gnd.n6875 gnd.n6874 0.152939
R11458 gnd.n6876 gnd.n6875 0.152939
R11459 gnd.n6877 gnd.n6876 0.152939
R11460 gnd.n6878 gnd.n6877 0.152939
R11461 gnd.n6879 gnd.n6878 0.152939
R11462 gnd.n6880 gnd.n6879 0.152939
R11463 gnd.n6881 gnd.n6880 0.152939
R11464 gnd.n6882 gnd.n6881 0.152939
R11465 gnd.n6883 gnd.n6882 0.152939
R11466 gnd.n6884 gnd.n6883 0.152939
R11467 gnd.n6885 gnd.n6884 0.152939
R11468 gnd.n6886 gnd.n6885 0.152939
R11469 gnd.n6887 gnd.n6886 0.152939
R11470 gnd.n6888 gnd.n6887 0.152939
R11471 gnd.n6889 gnd.n6888 0.152939
R11472 gnd.n6890 gnd.n6889 0.152939
R11473 gnd.n6891 gnd.n6890 0.152939
R11474 gnd.n6892 gnd.n6891 0.152939
R11475 gnd.n6893 gnd.n6892 0.152939
R11476 gnd.n6894 gnd.n6893 0.152939
R11477 gnd.n6895 gnd.n6894 0.152939
R11478 gnd.n6896 gnd.n6895 0.152939
R11479 gnd.n6897 gnd.n6896 0.152939
R11480 gnd.n6898 gnd.n6897 0.152939
R11481 gnd.n6899 gnd.n6898 0.152939
R11482 gnd.n6900 gnd.n6899 0.152939
R11483 gnd.n6901 gnd.n6900 0.152939
R11484 gnd.n6961 gnd.n6901 0.152939
R11485 gnd.n6961 gnd.n6960 0.152939
R11486 gnd.n6960 gnd.n6959 0.152939
R11487 gnd.n6959 gnd.n6905 0.152939
R11488 gnd.n6906 gnd.n6905 0.152939
R11489 gnd.n6907 gnd.n6906 0.152939
R11490 gnd.n6908 gnd.n6907 0.152939
R11491 gnd.n6909 gnd.n6908 0.152939
R11492 gnd.n6910 gnd.n6909 0.152939
R11493 gnd.n6911 gnd.n6910 0.152939
R11494 gnd.n6912 gnd.n6911 0.152939
R11495 gnd.n6913 gnd.n6912 0.152939
R11496 gnd.n6914 gnd.n6913 0.152939
R11497 gnd.n6915 gnd.n6914 0.152939
R11498 gnd.n6916 gnd.n6915 0.152939
R11499 gnd.n6917 gnd.n6916 0.152939
R11500 gnd.n6918 gnd.n6917 0.152939
R11501 gnd.n6919 gnd.n6918 0.152939
R11502 gnd.n6920 gnd.n6919 0.152939
R11503 gnd.n6921 gnd.n6920 0.152939
R11504 gnd.n6921 gnd.n6719 0.152939
R11505 gnd.n7047 gnd.n6719 0.152939
R11506 gnd.n5600 gnd.n4168 0.152939
R11507 gnd.n5600 gnd.n5599 0.152939
R11508 gnd.n5599 gnd.n5598 0.152939
R11509 gnd.n5598 gnd.n4170 0.152939
R11510 gnd.n4171 gnd.n4170 0.152939
R11511 gnd.n4172 gnd.n4171 0.152939
R11512 gnd.n4173 gnd.n4172 0.152939
R11513 gnd.n4174 gnd.n4173 0.152939
R11514 gnd.n4175 gnd.n4174 0.152939
R11515 gnd.n4176 gnd.n4175 0.152939
R11516 gnd.n4177 gnd.n4176 0.152939
R11517 gnd.n4178 gnd.n4177 0.152939
R11518 gnd.n4179 gnd.n4178 0.152939
R11519 gnd.n4180 gnd.n4179 0.152939
R11520 gnd.n5570 gnd.n4180 0.152939
R11521 gnd.n5570 gnd.n5569 0.152939
R11522 gnd.n4842 gnd.n4841 0.152939
R11523 gnd.n4842 gnd.n4546 0.152939
R11524 gnd.n4870 gnd.n4546 0.152939
R11525 gnd.n4871 gnd.n4870 0.152939
R11526 gnd.n4872 gnd.n4871 0.152939
R11527 gnd.n4873 gnd.n4872 0.152939
R11528 gnd.n4873 gnd.n4518 0.152939
R11529 gnd.n4900 gnd.n4518 0.152939
R11530 gnd.n4901 gnd.n4900 0.152939
R11531 gnd.n4902 gnd.n4901 0.152939
R11532 gnd.n4902 gnd.n4496 0.152939
R11533 gnd.n4931 gnd.n4496 0.152939
R11534 gnd.n4932 gnd.n4931 0.152939
R11535 gnd.n4933 gnd.n4932 0.152939
R11536 gnd.n4934 gnd.n4933 0.152939
R11537 gnd.n4936 gnd.n4934 0.152939
R11538 gnd.n4936 gnd.n4935 0.152939
R11539 gnd.n4935 gnd.n4445 0.152939
R11540 gnd.n4446 gnd.n4445 0.152939
R11541 gnd.n4447 gnd.n4446 0.152939
R11542 gnd.n4466 gnd.n4447 0.152939
R11543 gnd.n4467 gnd.n4466 0.152939
R11544 gnd.n4467 gnd.n4365 0.152939
R11545 gnd.n5026 gnd.n4365 0.152939
R11546 gnd.n5027 gnd.n5026 0.152939
R11547 gnd.n5028 gnd.n5027 0.152939
R11548 gnd.n5029 gnd.n5028 0.152939
R11549 gnd.n5029 gnd.n4338 0.152939
R11550 gnd.n5066 gnd.n4338 0.152939
R11551 gnd.n5067 gnd.n5066 0.152939
R11552 gnd.n5068 gnd.n5067 0.152939
R11553 gnd.n5069 gnd.n5068 0.152939
R11554 gnd.n5069 gnd.n4311 0.152939
R11555 gnd.n5111 gnd.n4311 0.152939
R11556 gnd.n5112 gnd.n5111 0.152939
R11557 gnd.n5113 gnd.n5112 0.152939
R11558 gnd.n5114 gnd.n5113 0.152939
R11559 gnd.n5114 gnd.n4283 0.152939
R11560 gnd.n5151 gnd.n4283 0.152939
R11561 gnd.n5152 gnd.n5151 0.152939
R11562 gnd.n5153 gnd.n5152 0.152939
R11563 gnd.n5154 gnd.n5153 0.152939
R11564 gnd.n5154 gnd.n4256 0.152939
R11565 gnd.n5200 gnd.n4256 0.152939
R11566 gnd.n5201 gnd.n5200 0.152939
R11567 gnd.n5202 gnd.n5201 0.152939
R11568 gnd.n5203 gnd.n5202 0.152939
R11569 gnd.n5203 gnd.n4229 0.152939
R11570 gnd.n5494 gnd.n4229 0.152939
R11571 gnd.n5495 gnd.n5494 0.152939
R11572 gnd.n5496 gnd.n5495 0.152939
R11573 gnd.n5497 gnd.n5496 0.152939
R11574 gnd.n5498 gnd.n5497 0.152939
R11575 gnd.n4840 gnd.n4570 0.152939
R11576 gnd.n4591 gnd.n4570 0.152939
R11577 gnd.n4592 gnd.n4591 0.152939
R11578 gnd.n4598 gnd.n4592 0.152939
R11579 gnd.n4599 gnd.n4598 0.152939
R11580 gnd.n4600 gnd.n4599 0.152939
R11581 gnd.n4600 gnd.n4589 0.152939
R11582 gnd.n4608 gnd.n4589 0.152939
R11583 gnd.n4609 gnd.n4608 0.152939
R11584 gnd.n4610 gnd.n4609 0.152939
R11585 gnd.n4610 gnd.n4587 0.152939
R11586 gnd.n4618 gnd.n4587 0.152939
R11587 gnd.n4619 gnd.n4618 0.152939
R11588 gnd.n4620 gnd.n4619 0.152939
R11589 gnd.n4620 gnd.n4585 0.152939
R11590 gnd.n4628 gnd.n4585 0.152939
R11591 gnd.n5567 gnd.n4185 0.152939
R11592 gnd.n4187 gnd.n4185 0.152939
R11593 gnd.n4188 gnd.n4187 0.152939
R11594 gnd.n4189 gnd.n4188 0.152939
R11595 gnd.n4190 gnd.n4189 0.152939
R11596 gnd.n4191 gnd.n4190 0.152939
R11597 gnd.n4192 gnd.n4191 0.152939
R11598 gnd.n4193 gnd.n4192 0.152939
R11599 gnd.n4194 gnd.n4193 0.152939
R11600 gnd.n4195 gnd.n4194 0.152939
R11601 gnd.n4196 gnd.n4195 0.152939
R11602 gnd.n4197 gnd.n4196 0.152939
R11603 gnd.n4198 gnd.n4197 0.152939
R11604 gnd.n4199 gnd.n4198 0.152939
R11605 gnd.n4200 gnd.n4199 0.152939
R11606 gnd.n4201 gnd.n4200 0.152939
R11607 gnd.n4202 gnd.n4201 0.152939
R11608 gnd.n4203 gnd.n4202 0.152939
R11609 gnd.n4204 gnd.n4203 0.152939
R11610 gnd.n4205 gnd.n4204 0.152939
R11611 gnd.n4206 gnd.n4205 0.152939
R11612 gnd.n4207 gnd.n4206 0.152939
R11613 gnd.n4211 gnd.n4207 0.152939
R11614 gnd.n4212 gnd.n4211 0.152939
R11615 gnd.n4213 gnd.n4212 0.152939
R11616 gnd.n4214 gnd.n4213 0.152939
R11617 gnd.n5003 gnd.n5002 0.152939
R11618 gnd.n5004 gnd.n5003 0.152939
R11619 gnd.n5005 gnd.n5004 0.152939
R11620 gnd.n5006 gnd.n5005 0.152939
R11621 gnd.n5007 gnd.n5006 0.152939
R11622 gnd.n5008 gnd.n5007 0.152939
R11623 gnd.n5008 gnd.n4319 0.152939
R11624 gnd.n5087 gnd.n4319 0.152939
R11625 gnd.n5088 gnd.n5087 0.152939
R11626 gnd.n5089 gnd.n5088 0.152939
R11627 gnd.n5090 gnd.n5089 0.152939
R11628 gnd.n5091 gnd.n5090 0.152939
R11629 gnd.n5092 gnd.n5091 0.152939
R11630 gnd.n5093 gnd.n5092 0.152939
R11631 gnd.n5094 gnd.n5093 0.152939
R11632 gnd.n5095 gnd.n5094 0.152939
R11633 gnd.n5095 gnd.n4263 0.152939
R11634 gnd.n5172 gnd.n4263 0.152939
R11635 gnd.n5173 gnd.n5172 0.152939
R11636 gnd.n5174 gnd.n5173 0.152939
R11637 gnd.n5175 gnd.n5174 0.152939
R11638 gnd.n5176 gnd.n5175 0.152939
R11639 gnd.n5177 gnd.n5176 0.152939
R11640 gnd.n5178 gnd.n5177 0.152939
R11641 gnd.n5179 gnd.n5178 0.152939
R11642 gnd.n5180 gnd.n5179 0.152939
R11643 gnd.n5182 gnd.n5180 0.152939
R11644 gnd.n5182 gnd.n5181 0.152939
R11645 gnd.n4758 gnd.n4757 0.152939
R11646 gnd.n4758 gnd.n4648 0.152939
R11647 gnd.n4773 gnd.n4648 0.152939
R11648 gnd.n4774 gnd.n4773 0.152939
R11649 gnd.n4775 gnd.n4774 0.152939
R11650 gnd.n4775 gnd.n4636 0.152939
R11651 gnd.n4789 gnd.n4636 0.152939
R11652 gnd.n4790 gnd.n4789 0.152939
R11653 gnd.n4791 gnd.n4790 0.152939
R11654 gnd.n4792 gnd.n4791 0.152939
R11655 gnd.n4793 gnd.n4792 0.152939
R11656 gnd.n4794 gnd.n4793 0.152939
R11657 gnd.n4795 gnd.n4794 0.152939
R11658 gnd.n4796 gnd.n4795 0.152939
R11659 gnd.n4797 gnd.n4796 0.152939
R11660 gnd.n4798 gnd.n4797 0.152939
R11661 gnd.n4799 gnd.n4798 0.152939
R11662 gnd.n4800 gnd.n4799 0.152939
R11663 gnd.n4801 gnd.n4800 0.152939
R11664 gnd.n4802 gnd.n4801 0.152939
R11665 gnd.n4803 gnd.n4802 0.152939
R11666 gnd.n4803 gnd.n4502 0.152939
R11667 gnd.n4920 gnd.n4502 0.152939
R11668 gnd.n4921 gnd.n4920 0.152939
R11669 gnd.n4922 gnd.n4921 0.152939
R11670 gnd.n4923 gnd.n4922 0.152939
R11671 gnd.n4923 gnd.n4424 0.152939
R11672 gnd.n5000 gnd.n4424 0.152939
R11673 gnd.n4676 gnd.n4675 0.152939
R11674 gnd.n4677 gnd.n4676 0.152939
R11675 gnd.n4678 gnd.n4677 0.152939
R11676 gnd.n4679 gnd.n4678 0.152939
R11677 gnd.n4680 gnd.n4679 0.152939
R11678 gnd.n4681 gnd.n4680 0.152939
R11679 gnd.n4682 gnd.n4681 0.152939
R11680 gnd.n4683 gnd.n4682 0.152939
R11681 gnd.n4684 gnd.n4683 0.152939
R11682 gnd.n4685 gnd.n4684 0.152939
R11683 gnd.n4686 gnd.n4685 0.152939
R11684 gnd.n4687 gnd.n4686 0.152939
R11685 gnd.n4688 gnd.n4687 0.152939
R11686 gnd.n4689 gnd.n4688 0.152939
R11687 gnd.n4690 gnd.n4689 0.152939
R11688 gnd.n4691 gnd.n4690 0.152939
R11689 gnd.n4692 gnd.n4691 0.152939
R11690 gnd.n4693 gnd.n4692 0.152939
R11691 gnd.n4694 gnd.n4693 0.152939
R11692 gnd.n4695 gnd.n4694 0.152939
R11693 gnd.n4696 gnd.n4695 0.152939
R11694 gnd.n4697 gnd.n4696 0.152939
R11695 gnd.n4701 gnd.n4697 0.152939
R11696 gnd.n4702 gnd.n4701 0.152939
R11697 gnd.n4702 gnd.n4659 0.152939
R11698 gnd.n4756 gnd.n4659 0.152939
R11699 gnd.n2459 gnd.n2402 0.152939
R11700 gnd.n2465 gnd.n2402 0.152939
R11701 gnd.n2466 gnd.n2465 0.152939
R11702 gnd.n2467 gnd.n2466 0.152939
R11703 gnd.n2467 gnd.n2400 0.152939
R11704 gnd.n2473 gnd.n2400 0.152939
R11705 gnd.n2474 gnd.n2473 0.152939
R11706 gnd.n2475 gnd.n2474 0.152939
R11707 gnd.n2475 gnd.n2398 0.152939
R11708 gnd.n2481 gnd.n2398 0.152939
R11709 gnd.n2482 gnd.n2481 0.152939
R11710 gnd.n2483 gnd.n2482 0.152939
R11711 gnd.n2483 gnd.n2396 0.152939
R11712 gnd.n2489 gnd.n2396 0.152939
R11713 gnd.n2490 gnd.n2489 0.152939
R11714 gnd.n2491 gnd.n2490 0.152939
R11715 gnd.n2491 gnd.n2394 0.152939
R11716 gnd.n2497 gnd.n2394 0.152939
R11717 gnd.n2498 gnd.n2497 0.152939
R11718 gnd.n2499 gnd.n2498 0.152939
R11719 gnd.n3906 gnd.n1336 0.152939
R11720 gnd.n1380 gnd.n1336 0.152939
R11721 gnd.n1381 gnd.n1380 0.152939
R11722 gnd.n1382 gnd.n1381 0.152939
R11723 gnd.n1383 gnd.n1382 0.152939
R11724 gnd.n1384 gnd.n1383 0.152939
R11725 gnd.n1385 gnd.n1384 0.152939
R11726 gnd.n1386 gnd.n1385 0.152939
R11727 gnd.n1387 gnd.n1386 0.152939
R11728 gnd.n1388 gnd.n1387 0.152939
R11729 gnd.n1389 gnd.n1388 0.152939
R11730 gnd.n1390 gnd.n1389 0.152939
R11731 gnd.n1391 gnd.n1390 0.152939
R11732 gnd.n1392 gnd.n1391 0.152939
R11733 gnd.n1393 gnd.n1392 0.152939
R11734 gnd.n1394 gnd.n1393 0.152939
R11735 gnd.n1395 gnd.n1394 0.152939
R11736 gnd.n1398 gnd.n1395 0.152939
R11737 gnd.n1399 gnd.n1398 0.152939
R11738 gnd.n1400 gnd.n1399 0.152939
R11739 gnd.n1401 gnd.n1400 0.152939
R11740 gnd.n1402 gnd.n1401 0.152939
R11741 gnd.n1403 gnd.n1402 0.152939
R11742 gnd.n1404 gnd.n1403 0.152939
R11743 gnd.n1405 gnd.n1404 0.152939
R11744 gnd.n2222 gnd.n2221 0.152939
R11745 gnd.n2223 gnd.n2222 0.152939
R11746 gnd.n2223 gnd.n2217 0.152939
R11747 gnd.n2231 gnd.n2217 0.152939
R11748 gnd.n2232 gnd.n2231 0.152939
R11749 gnd.n2233 gnd.n2232 0.152939
R11750 gnd.n2233 gnd.n2215 0.152939
R11751 gnd.n2241 gnd.n2215 0.152939
R11752 gnd.n2242 gnd.n2241 0.152939
R11753 gnd.n2243 gnd.n2242 0.152939
R11754 gnd.n2243 gnd.n2211 0.152939
R11755 gnd.n2251 gnd.n2211 0.152939
R11756 gnd.n2252 gnd.n2251 0.152939
R11757 gnd.n2253 gnd.n2252 0.152939
R11758 gnd.n2253 gnd.n2209 0.152939
R11759 gnd.n2261 gnd.n2209 0.152939
R11760 gnd.n2262 gnd.n2261 0.152939
R11761 gnd.n2263 gnd.n2262 0.152939
R11762 gnd.n2263 gnd.n2207 0.152939
R11763 gnd.n2271 gnd.n2207 0.152939
R11764 gnd.n2272 gnd.n2271 0.152939
R11765 gnd.n2273 gnd.n2272 0.152939
R11766 gnd.n2273 gnd.n2205 0.152939
R11767 gnd.n2281 gnd.n2205 0.152939
R11768 gnd.n2282 gnd.n2281 0.152939
R11769 gnd.n2283 gnd.n2282 0.152939
R11770 gnd.n2283 gnd.n2203 0.152939
R11771 gnd.n2291 gnd.n2203 0.152939
R11772 gnd.n2292 gnd.n2291 0.152939
R11773 gnd.n2293 gnd.n2292 0.152939
R11774 gnd.n1258 gnd.n1257 0.152939
R11775 gnd.n1274 gnd.n1258 0.152939
R11776 gnd.n1275 gnd.n1274 0.152939
R11777 gnd.n1276 gnd.n1275 0.152939
R11778 gnd.n1277 gnd.n1276 0.152939
R11779 gnd.n1293 gnd.n1277 0.152939
R11780 gnd.n1294 gnd.n1293 0.152939
R11781 gnd.n1295 gnd.n1294 0.152939
R11782 gnd.n1296 gnd.n1295 0.152939
R11783 gnd.n1314 gnd.n1296 0.152939
R11784 gnd.n1315 gnd.n1314 0.152939
R11785 gnd.n1316 gnd.n1315 0.152939
R11786 gnd.n1317 gnd.n1316 0.152939
R11787 gnd.n1334 gnd.n1317 0.152939
R11788 gnd.n1335 gnd.n1334 0.152939
R11789 gnd.n3907 gnd.n1335 0.152939
R11790 gnd.n4030 gnd.n1142 0.152939
R11791 gnd.n4030 gnd.n4029 0.152939
R11792 gnd.n4029 gnd.n4028 0.152939
R11793 gnd.n4028 gnd.n1143 0.152939
R11794 gnd.n1161 gnd.n1143 0.152939
R11795 gnd.n1162 gnd.n1161 0.152939
R11796 gnd.n1163 gnd.n1162 0.152939
R11797 gnd.n1178 gnd.n1163 0.152939
R11798 gnd.n1179 gnd.n1178 0.152939
R11799 gnd.n1180 gnd.n1179 0.152939
R11800 gnd.n1181 gnd.n1180 0.152939
R11801 gnd.n1198 gnd.n1181 0.152939
R11802 gnd.n1199 gnd.n1198 0.152939
R11803 gnd.n1200 gnd.n1199 0.152939
R11804 gnd.n1201 gnd.n1200 0.152939
R11805 gnd.n1216 gnd.n1201 0.152939
R11806 gnd.n1066 gnd.n1065 0.152939
R11807 gnd.n1067 gnd.n1066 0.152939
R11808 gnd.n1068 gnd.n1067 0.152939
R11809 gnd.n1069 gnd.n1068 0.152939
R11810 gnd.n1070 gnd.n1069 0.152939
R11811 gnd.n1071 gnd.n1070 0.152939
R11812 gnd.n1072 gnd.n1071 0.152939
R11813 gnd.n1073 gnd.n1072 0.152939
R11814 gnd.n1074 gnd.n1073 0.152939
R11815 gnd.n1075 gnd.n1074 0.152939
R11816 gnd.n1076 gnd.n1075 0.152939
R11817 gnd.n1077 gnd.n1076 0.152939
R11818 gnd.n1078 gnd.n1077 0.152939
R11819 gnd.n1079 gnd.n1078 0.152939
R11820 gnd.n1080 gnd.n1079 0.152939
R11821 gnd.n1081 gnd.n1080 0.152939
R11822 gnd.n1082 gnd.n1081 0.152939
R11823 gnd.n1085 gnd.n1082 0.152939
R11824 gnd.n1086 gnd.n1085 0.152939
R11825 gnd.n1087 gnd.n1086 0.152939
R11826 gnd.n1088 gnd.n1087 0.152939
R11827 gnd.n1089 gnd.n1088 0.152939
R11828 gnd.n1090 gnd.n1089 0.152939
R11829 gnd.n1091 gnd.n1090 0.152939
R11830 gnd.n1092 gnd.n1091 0.152939
R11831 gnd.n1093 gnd.n1092 0.152939
R11832 gnd.n1094 gnd.n1093 0.152939
R11833 gnd.n1095 gnd.n1094 0.152939
R11834 gnd.n1096 gnd.n1095 0.152939
R11835 gnd.n1097 gnd.n1096 0.152939
R11836 gnd.n1098 gnd.n1097 0.152939
R11837 gnd.n1099 gnd.n1098 0.152939
R11838 gnd.n1100 gnd.n1099 0.152939
R11839 gnd.n1101 gnd.n1100 0.152939
R11840 gnd.n1102 gnd.n1101 0.152939
R11841 gnd.n1103 gnd.n1102 0.152939
R11842 gnd.n1104 gnd.n1103 0.152939
R11843 gnd.n1107 gnd.n1104 0.152939
R11844 gnd.n1108 gnd.n1107 0.152939
R11845 gnd.n1109 gnd.n1108 0.152939
R11846 gnd.n1110 gnd.n1109 0.152939
R11847 gnd.n1111 gnd.n1110 0.152939
R11848 gnd.n1112 gnd.n1111 0.152939
R11849 gnd.n1113 gnd.n1112 0.152939
R11850 gnd.n1114 gnd.n1113 0.152939
R11851 gnd.n1115 gnd.n1114 0.152939
R11852 gnd.n1116 gnd.n1115 0.152939
R11853 gnd.n1117 gnd.n1116 0.152939
R11854 gnd.n1118 gnd.n1117 0.152939
R11855 gnd.n1119 gnd.n1118 0.152939
R11856 gnd.n1120 gnd.n1119 0.152939
R11857 gnd.n1121 gnd.n1120 0.152939
R11858 gnd.n1122 gnd.n1121 0.152939
R11859 gnd.n1123 gnd.n1122 0.152939
R11860 gnd.n1124 gnd.n1123 0.152939
R11861 gnd.n1125 gnd.n1124 0.152939
R11862 gnd.n4040 gnd.n1125 0.152939
R11863 gnd.n4040 gnd.n4039 0.152939
R11864 gnd.n2416 gnd.n1129 0.152939
R11865 gnd.n2422 gnd.n2416 0.152939
R11866 gnd.n2423 gnd.n2422 0.152939
R11867 gnd.n2424 gnd.n2423 0.152939
R11868 gnd.n2424 gnd.n2414 0.152939
R11869 gnd.n2432 gnd.n2414 0.152939
R11870 gnd.n2433 gnd.n2432 0.152939
R11871 gnd.n2434 gnd.n2433 0.152939
R11872 gnd.n2434 gnd.n2412 0.152939
R11873 gnd.n2442 gnd.n2412 0.152939
R11874 gnd.n2443 gnd.n2442 0.152939
R11875 gnd.n2444 gnd.n2443 0.152939
R11876 gnd.n2444 gnd.n2410 0.152939
R11877 gnd.n2452 gnd.n2410 0.152939
R11878 gnd.n2453 gnd.n2452 0.152939
R11879 gnd.n2454 gnd.n2453 0.152939
R11880 gnd.n2454 gnd.n2403 0.152939
R11881 gnd.n2458 gnd.n2403 0.152939
R11882 gnd.n5778 gnd.n5777 0.152939
R11883 gnd.n5779 gnd.n5778 0.152939
R11884 gnd.n5779 gnd.n832 0.152939
R11885 gnd.n5787 gnd.n832 0.152939
R11886 gnd.n5788 gnd.n5787 0.152939
R11887 gnd.n5789 gnd.n5788 0.152939
R11888 gnd.n5789 gnd.n826 0.152939
R11889 gnd.n5797 gnd.n826 0.152939
R11890 gnd.n5798 gnd.n5797 0.152939
R11891 gnd.n5799 gnd.n5798 0.152939
R11892 gnd.n5799 gnd.n820 0.152939
R11893 gnd.n5807 gnd.n820 0.152939
R11894 gnd.n5808 gnd.n5807 0.152939
R11895 gnd.n5809 gnd.n5808 0.152939
R11896 gnd.n5809 gnd.n814 0.152939
R11897 gnd.n5817 gnd.n814 0.152939
R11898 gnd.n5818 gnd.n5817 0.152939
R11899 gnd.n5819 gnd.n5818 0.152939
R11900 gnd.n5819 gnd.n808 0.152939
R11901 gnd.n5827 gnd.n808 0.152939
R11902 gnd.n5828 gnd.n5827 0.152939
R11903 gnd.n5829 gnd.n5828 0.152939
R11904 gnd.n5829 gnd.n802 0.152939
R11905 gnd.n5837 gnd.n802 0.152939
R11906 gnd.n5838 gnd.n5837 0.152939
R11907 gnd.n5839 gnd.n5838 0.152939
R11908 gnd.n5839 gnd.n796 0.152939
R11909 gnd.n5847 gnd.n796 0.152939
R11910 gnd.n5848 gnd.n5847 0.152939
R11911 gnd.n5849 gnd.n5848 0.152939
R11912 gnd.n5849 gnd.n790 0.152939
R11913 gnd.n5857 gnd.n790 0.152939
R11914 gnd.n5858 gnd.n5857 0.152939
R11915 gnd.n5859 gnd.n5858 0.152939
R11916 gnd.n5859 gnd.n784 0.152939
R11917 gnd.n5867 gnd.n784 0.152939
R11918 gnd.n5868 gnd.n5867 0.152939
R11919 gnd.n5869 gnd.n5868 0.152939
R11920 gnd.n5869 gnd.n778 0.152939
R11921 gnd.n5877 gnd.n778 0.152939
R11922 gnd.n5878 gnd.n5877 0.152939
R11923 gnd.n5879 gnd.n5878 0.152939
R11924 gnd.n5879 gnd.n772 0.152939
R11925 gnd.n5887 gnd.n772 0.152939
R11926 gnd.n5888 gnd.n5887 0.152939
R11927 gnd.n5889 gnd.n5888 0.152939
R11928 gnd.n5889 gnd.n766 0.152939
R11929 gnd.n5897 gnd.n766 0.152939
R11930 gnd.n5898 gnd.n5897 0.152939
R11931 gnd.n5899 gnd.n5898 0.152939
R11932 gnd.n5899 gnd.n760 0.152939
R11933 gnd.n5907 gnd.n760 0.152939
R11934 gnd.n5908 gnd.n5907 0.152939
R11935 gnd.n5909 gnd.n5908 0.152939
R11936 gnd.n5909 gnd.n754 0.152939
R11937 gnd.n5917 gnd.n754 0.152939
R11938 gnd.n5918 gnd.n5917 0.152939
R11939 gnd.n5919 gnd.n5918 0.152939
R11940 gnd.n5919 gnd.n748 0.152939
R11941 gnd.n5927 gnd.n748 0.152939
R11942 gnd.n5928 gnd.n5927 0.152939
R11943 gnd.n5929 gnd.n5928 0.152939
R11944 gnd.n5929 gnd.n742 0.152939
R11945 gnd.n5937 gnd.n742 0.152939
R11946 gnd.n5938 gnd.n5937 0.152939
R11947 gnd.n5939 gnd.n5938 0.152939
R11948 gnd.n5939 gnd.n736 0.152939
R11949 gnd.n5947 gnd.n736 0.152939
R11950 gnd.n5948 gnd.n5947 0.152939
R11951 gnd.n5949 gnd.n5948 0.152939
R11952 gnd.n5949 gnd.n730 0.152939
R11953 gnd.n5957 gnd.n730 0.152939
R11954 gnd.n5958 gnd.n5957 0.152939
R11955 gnd.n5959 gnd.n5958 0.152939
R11956 gnd.n5959 gnd.n724 0.152939
R11957 gnd.n5967 gnd.n724 0.152939
R11958 gnd.n5968 gnd.n5967 0.152939
R11959 gnd.n5969 gnd.n5968 0.152939
R11960 gnd.n5969 gnd.n718 0.152939
R11961 gnd.n5977 gnd.n718 0.152939
R11962 gnd.n5978 gnd.n5977 0.152939
R11963 gnd.n5979 gnd.n5978 0.152939
R11964 gnd.n5979 gnd.n712 0.152939
R11965 gnd.n5987 gnd.n712 0.152939
R11966 gnd.n5988 gnd.n5987 0.152939
R11967 gnd.n5989 gnd.n5988 0.152939
R11968 gnd.n5989 gnd.n706 0.152939
R11969 gnd.n5997 gnd.n706 0.152939
R11970 gnd.n5998 gnd.n5997 0.152939
R11971 gnd.n5999 gnd.n5998 0.152939
R11972 gnd.n5999 gnd.n700 0.152939
R11973 gnd.n6007 gnd.n700 0.152939
R11974 gnd.n6008 gnd.n6007 0.152939
R11975 gnd.n6009 gnd.n6008 0.152939
R11976 gnd.n6009 gnd.n694 0.152939
R11977 gnd.n6017 gnd.n694 0.152939
R11978 gnd.n6018 gnd.n6017 0.152939
R11979 gnd.n6019 gnd.n6018 0.152939
R11980 gnd.n6019 gnd.n688 0.152939
R11981 gnd.n6027 gnd.n688 0.152939
R11982 gnd.n6028 gnd.n6027 0.152939
R11983 gnd.n6029 gnd.n6028 0.152939
R11984 gnd.n6029 gnd.n682 0.152939
R11985 gnd.n6037 gnd.n682 0.152939
R11986 gnd.n6038 gnd.n6037 0.152939
R11987 gnd.n6039 gnd.n6038 0.152939
R11988 gnd.n6039 gnd.n676 0.152939
R11989 gnd.n6047 gnd.n676 0.152939
R11990 gnd.n6048 gnd.n6047 0.152939
R11991 gnd.n6049 gnd.n6048 0.152939
R11992 gnd.n6049 gnd.n670 0.152939
R11993 gnd.n6057 gnd.n670 0.152939
R11994 gnd.n6058 gnd.n6057 0.152939
R11995 gnd.n6059 gnd.n6058 0.152939
R11996 gnd.n6059 gnd.n664 0.152939
R11997 gnd.n6067 gnd.n664 0.152939
R11998 gnd.n6068 gnd.n6067 0.152939
R11999 gnd.n6069 gnd.n6068 0.152939
R12000 gnd.n6069 gnd.n658 0.152939
R12001 gnd.n6077 gnd.n658 0.152939
R12002 gnd.n6078 gnd.n6077 0.152939
R12003 gnd.n6079 gnd.n6078 0.152939
R12004 gnd.n6079 gnd.n652 0.152939
R12005 gnd.n6087 gnd.n652 0.152939
R12006 gnd.n6088 gnd.n6087 0.152939
R12007 gnd.n6089 gnd.n6088 0.152939
R12008 gnd.n6089 gnd.n646 0.152939
R12009 gnd.n6097 gnd.n646 0.152939
R12010 gnd.n6099 gnd.n6098 0.152939
R12011 gnd.n6099 gnd.n640 0.152939
R12012 gnd.n6107 gnd.n640 0.152939
R12013 gnd.n6108 gnd.n6107 0.152939
R12014 gnd.n6109 gnd.n6108 0.152939
R12015 gnd.n6109 gnd.n634 0.152939
R12016 gnd.n6117 gnd.n634 0.152939
R12017 gnd.n6118 gnd.n6117 0.152939
R12018 gnd.n6119 gnd.n6118 0.152939
R12019 gnd.n6119 gnd.n628 0.152939
R12020 gnd.n6127 gnd.n628 0.152939
R12021 gnd.n6128 gnd.n6127 0.152939
R12022 gnd.n6129 gnd.n6128 0.152939
R12023 gnd.n6129 gnd.n622 0.152939
R12024 gnd.n6137 gnd.n622 0.152939
R12025 gnd.n6138 gnd.n6137 0.152939
R12026 gnd.n6139 gnd.n6138 0.152939
R12027 gnd.n6139 gnd.n616 0.152939
R12028 gnd.n6147 gnd.n616 0.152939
R12029 gnd.n6148 gnd.n6147 0.152939
R12030 gnd.n6149 gnd.n6148 0.152939
R12031 gnd.n6149 gnd.n610 0.152939
R12032 gnd.n6157 gnd.n610 0.152939
R12033 gnd.n6158 gnd.n6157 0.152939
R12034 gnd.n6159 gnd.n6158 0.152939
R12035 gnd.n6159 gnd.n604 0.152939
R12036 gnd.n6167 gnd.n604 0.152939
R12037 gnd.n6168 gnd.n6167 0.152939
R12038 gnd.n6169 gnd.n6168 0.152939
R12039 gnd.n6169 gnd.n598 0.152939
R12040 gnd.n6177 gnd.n598 0.152939
R12041 gnd.n6178 gnd.n6177 0.152939
R12042 gnd.n6179 gnd.n6178 0.152939
R12043 gnd.n6179 gnd.n592 0.152939
R12044 gnd.n6187 gnd.n592 0.152939
R12045 gnd.n6188 gnd.n6187 0.152939
R12046 gnd.n6189 gnd.n6188 0.152939
R12047 gnd.n6189 gnd.n586 0.152939
R12048 gnd.n6197 gnd.n586 0.152939
R12049 gnd.n6198 gnd.n6197 0.152939
R12050 gnd.n6199 gnd.n6198 0.152939
R12051 gnd.n6199 gnd.n580 0.152939
R12052 gnd.n6207 gnd.n580 0.152939
R12053 gnd.n6208 gnd.n6207 0.152939
R12054 gnd.n6209 gnd.n6208 0.152939
R12055 gnd.n6209 gnd.n574 0.152939
R12056 gnd.n6217 gnd.n574 0.152939
R12057 gnd.n6218 gnd.n6217 0.152939
R12058 gnd.n6219 gnd.n6218 0.152939
R12059 gnd.n6219 gnd.n568 0.152939
R12060 gnd.n6227 gnd.n568 0.152939
R12061 gnd.n6228 gnd.n6227 0.152939
R12062 gnd.n6229 gnd.n6228 0.152939
R12063 gnd.n6229 gnd.n562 0.152939
R12064 gnd.n6237 gnd.n562 0.152939
R12065 gnd.n6238 gnd.n6237 0.152939
R12066 gnd.n6239 gnd.n6238 0.152939
R12067 gnd.n6239 gnd.n556 0.152939
R12068 gnd.n6247 gnd.n556 0.152939
R12069 gnd.n6248 gnd.n6247 0.152939
R12070 gnd.n6249 gnd.n6248 0.152939
R12071 gnd.n6249 gnd.n550 0.152939
R12072 gnd.n6257 gnd.n550 0.152939
R12073 gnd.n6258 gnd.n6257 0.152939
R12074 gnd.n6259 gnd.n6258 0.152939
R12075 gnd.n6259 gnd.n544 0.152939
R12076 gnd.n6267 gnd.n544 0.152939
R12077 gnd.n6268 gnd.n6267 0.152939
R12078 gnd.n6269 gnd.n6268 0.152939
R12079 gnd.n6269 gnd.n538 0.152939
R12080 gnd.n6277 gnd.n538 0.152939
R12081 gnd.n6278 gnd.n6277 0.152939
R12082 gnd.n6279 gnd.n6278 0.152939
R12083 gnd.n6279 gnd.n532 0.152939
R12084 gnd.n6287 gnd.n532 0.152939
R12085 gnd.n6288 gnd.n6287 0.152939
R12086 gnd.n6289 gnd.n6288 0.152939
R12087 gnd.n6289 gnd.n526 0.152939
R12088 gnd.n6297 gnd.n526 0.152939
R12089 gnd.n6298 gnd.n6297 0.152939
R12090 gnd.n6299 gnd.n6298 0.152939
R12091 gnd.n6300 gnd.n6299 0.152939
R12092 gnd.n6300 gnd.n520 0.152939
R12093 gnd.n6311 gnd.n520 0.152939
R12094 gnd.n2310 gnd.n2305 0.152939
R12095 gnd.n2311 gnd.n2310 0.152939
R12096 gnd.n2312 gnd.n2311 0.152939
R12097 gnd.n2312 gnd.n2300 0.152939
R12098 gnd.n2569 gnd.n2300 0.152939
R12099 gnd.n2570 gnd.n2569 0.152939
R12100 gnd.n2571 gnd.n2570 0.152939
R12101 gnd.n2572 gnd.n2571 0.152939
R12102 gnd.n2573 gnd.n2572 0.152939
R12103 gnd.n2576 gnd.n2573 0.152939
R12104 gnd.n2577 gnd.n2576 0.152939
R12105 gnd.n2578 gnd.n2577 0.152939
R12106 gnd.n2579 gnd.n2578 0.152939
R12107 gnd.n2580 gnd.n2579 0.152939
R12108 gnd.n2580 gnd.n2092 0.152939
R12109 gnd.n2683 gnd.n2092 0.152939
R12110 gnd.n2684 gnd.n2683 0.152939
R12111 gnd.n2685 gnd.n2684 0.152939
R12112 gnd.n2686 gnd.n2685 0.152939
R12113 gnd.n2686 gnd.n2067 0.152939
R12114 gnd.n2713 gnd.n2067 0.152939
R12115 gnd.n2714 gnd.n2713 0.152939
R12116 gnd.n2715 gnd.n2714 0.152939
R12117 gnd.n2716 gnd.n2715 0.152939
R12118 gnd.n2716 gnd.n2042 0.152939
R12119 gnd.n2743 gnd.n2042 0.152939
R12120 gnd.n2744 gnd.n2743 0.152939
R12121 gnd.n2745 gnd.n2744 0.152939
R12122 gnd.n2746 gnd.n2745 0.152939
R12123 gnd.n2746 gnd.n2017 0.152939
R12124 gnd.n2776 gnd.n2017 0.152939
R12125 gnd.n2777 gnd.n2776 0.152939
R12126 gnd.n2778 gnd.n2777 0.152939
R12127 gnd.n2779 gnd.n2778 0.152939
R12128 gnd.n2780 gnd.n2779 0.152939
R12129 gnd.n2783 gnd.n2780 0.152939
R12130 gnd.n2784 gnd.n2783 0.152939
R12131 gnd.n2785 gnd.n2784 0.152939
R12132 gnd.n2785 gnd.n1987 0.152939
R12133 gnd.n2928 gnd.n1987 0.152939
R12134 gnd.n2929 gnd.n2928 0.152939
R12135 gnd.n2930 gnd.n2929 0.152939
R12136 gnd.n2931 gnd.n2930 0.152939
R12137 gnd.n2931 gnd.n1959 0.152939
R12138 gnd.n2970 gnd.n1959 0.152939
R12139 gnd.n2971 gnd.n2970 0.152939
R12140 gnd.n2972 gnd.n2971 0.152939
R12141 gnd.n2972 gnd.n1936 0.152939
R12142 gnd.n3014 gnd.n1936 0.152939
R12143 gnd.n3015 gnd.n3014 0.152939
R12144 gnd.n3016 gnd.n3015 0.152939
R12145 gnd.n3016 gnd.n1918 0.152939
R12146 gnd.n3070 gnd.n1918 0.152939
R12147 gnd.n3071 gnd.n3070 0.152939
R12148 gnd.n3072 gnd.n3071 0.152939
R12149 gnd.n3072 gnd.n1896 0.152939
R12150 gnd.n3098 gnd.n1896 0.152939
R12151 gnd.n3099 gnd.n3098 0.152939
R12152 gnd.n3100 gnd.n3099 0.152939
R12153 gnd.n3101 gnd.n3100 0.152939
R12154 gnd.n3101 gnd.n1864 0.152939
R12155 gnd.n3143 gnd.n1864 0.152939
R12156 gnd.n3144 gnd.n3143 0.152939
R12157 gnd.n3145 gnd.n3144 0.152939
R12158 gnd.n3145 gnd.n1840 0.152939
R12159 gnd.n3184 gnd.n1840 0.152939
R12160 gnd.n3185 gnd.n3184 0.152939
R12161 gnd.n3186 gnd.n3185 0.152939
R12162 gnd.n3186 gnd.n1823 0.152939
R12163 gnd.n3243 gnd.n1823 0.152939
R12164 gnd.n3244 gnd.n3243 0.152939
R12165 gnd.n3245 gnd.n3244 0.152939
R12166 gnd.n3245 gnd.n1802 0.152939
R12167 gnd.n3270 gnd.n1802 0.152939
R12168 gnd.n3271 gnd.n3270 0.152939
R12169 gnd.n3272 gnd.n3271 0.152939
R12170 gnd.n3273 gnd.n3272 0.152939
R12171 gnd.n3273 gnd.n1773 0.152939
R12172 gnd.n3317 gnd.n1773 0.152939
R12173 gnd.n3318 gnd.n3317 0.152939
R12174 gnd.n3319 gnd.n3318 0.152939
R12175 gnd.n3319 gnd.n1750 0.152939
R12176 gnd.n3358 gnd.n1750 0.152939
R12177 gnd.n3359 gnd.n3358 0.152939
R12178 gnd.n3360 gnd.n3359 0.152939
R12179 gnd.n3360 gnd.n1734 0.152939
R12180 gnd.n3400 gnd.n1734 0.152939
R12181 gnd.n3401 gnd.n3400 0.152939
R12182 gnd.n3402 gnd.n3401 0.152939
R12183 gnd.n3402 gnd.n1642 0.152939
R12184 gnd.n3547 gnd.n1642 0.152939
R12185 gnd.n3548 gnd.n3547 0.152939
R12186 gnd.n3549 gnd.n3548 0.152939
R12187 gnd.n3549 gnd.n1629 0.152939
R12188 gnd.n3567 gnd.n1629 0.152939
R12189 gnd.n3568 gnd.n3567 0.152939
R12190 gnd.n3569 gnd.n3568 0.152939
R12191 gnd.n3569 gnd.n1618 0.152939
R12192 gnd.n3589 gnd.n1618 0.152939
R12193 gnd.n3590 gnd.n3589 0.152939
R12194 gnd.n3591 gnd.n3590 0.152939
R12195 gnd.n3591 gnd.n1605 0.152939
R12196 gnd.n3609 gnd.n1605 0.152939
R12197 gnd.n3610 gnd.n3609 0.152939
R12198 gnd.n3611 gnd.n3610 0.152939
R12199 gnd.n3611 gnd.n1592 0.152939
R12200 gnd.n3629 gnd.n1592 0.152939
R12201 gnd.n3630 gnd.n3629 0.152939
R12202 gnd.n3631 gnd.n3630 0.152939
R12203 gnd.n3631 gnd.n1578 0.152939
R12204 gnd.n3649 gnd.n1578 0.152939
R12205 gnd.n3650 gnd.n3649 0.152939
R12206 gnd.n3651 gnd.n3650 0.152939
R12207 gnd.n3652 gnd.n3651 0.152939
R12208 gnd.n3654 gnd.n3652 0.152939
R12209 gnd.n3654 gnd.n3653 0.152939
R12210 gnd.n3653 gnd.n494 0.152939
R12211 gnd.n495 gnd.n494 0.152939
R12212 gnd.n496 gnd.n495 0.152939
R12213 gnd.n509 gnd.n496 0.152939
R12214 gnd.n510 gnd.n509 0.152939
R12215 gnd.n511 gnd.n510 0.152939
R12216 gnd.n512 gnd.n511 0.152939
R12217 gnd.n513 gnd.n512 0.152939
R12218 gnd.n514 gnd.n513 0.152939
R12219 gnd.n518 gnd.n514 0.152939
R12220 gnd.n519 gnd.n518 0.152939
R12221 gnd.n6312 gnd.n519 0.152939
R12222 gnd.n843 gnd.n838 0.152939
R12223 gnd.n844 gnd.n843 0.152939
R12224 gnd.n845 gnd.n844 0.152939
R12225 gnd.n850 gnd.n845 0.152939
R12226 gnd.n851 gnd.n850 0.152939
R12227 gnd.n852 gnd.n851 0.152939
R12228 gnd.n853 gnd.n852 0.152939
R12229 gnd.n858 gnd.n853 0.152939
R12230 gnd.n859 gnd.n858 0.152939
R12231 gnd.n860 gnd.n859 0.152939
R12232 gnd.n861 gnd.n860 0.152939
R12233 gnd.n866 gnd.n861 0.152939
R12234 gnd.n867 gnd.n866 0.152939
R12235 gnd.n868 gnd.n867 0.152939
R12236 gnd.n869 gnd.n868 0.152939
R12237 gnd.n874 gnd.n869 0.152939
R12238 gnd.n875 gnd.n874 0.152939
R12239 gnd.n876 gnd.n875 0.152939
R12240 gnd.n877 gnd.n876 0.152939
R12241 gnd.n882 gnd.n877 0.152939
R12242 gnd.n883 gnd.n882 0.152939
R12243 gnd.n884 gnd.n883 0.152939
R12244 gnd.n885 gnd.n884 0.152939
R12245 gnd.n890 gnd.n885 0.152939
R12246 gnd.n891 gnd.n890 0.152939
R12247 gnd.n892 gnd.n891 0.152939
R12248 gnd.n893 gnd.n892 0.152939
R12249 gnd.n898 gnd.n893 0.152939
R12250 gnd.n899 gnd.n898 0.152939
R12251 gnd.n900 gnd.n899 0.152939
R12252 gnd.n901 gnd.n900 0.152939
R12253 gnd.n906 gnd.n901 0.152939
R12254 gnd.n907 gnd.n906 0.152939
R12255 gnd.n908 gnd.n907 0.152939
R12256 gnd.n909 gnd.n908 0.152939
R12257 gnd.n914 gnd.n909 0.152939
R12258 gnd.n915 gnd.n914 0.152939
R12259 gnd.n916 gnd.n915 0.152939
R12260 gnd.n917 gnd.n916 0.152939
R12261 gnd.n922 gnd.n917 0.152939
R12262 gnd.n923 gnd.n922 0.152939
R12263 gnd.n924 gnd.n923 0.152939
R12264 gnd.n925 gnd.n924 0.152939
R12265 gnd.n930 gnd.n925 0.152939
R12266 gnd.n931 gnd.n930 0.152939
R12267 gnd.n932 gnd.n931 0.152939
R12268 gnd.n933 gnd.n932 0.152939
R12269 gnd.n938 gnd.n933 0.152939
R12270 gnd.n939 gnd.n938 0.152939
R12271 gnd.n940 gnd.n939 0.152939
R12272 gnd.n941 gnd.n940 0.152939
R12273 gnd.n946 gnd.n941 0.152939
R12274 gnd.n947 gnd.n946 0.152939
R12275 gnd.n948 gnd.n947 0.152939
R12276 gnd.n949 gnd.n948 0.152939
R12277 gnd.n954 gnd.n949 0.152939
R12278 gnd.n955 gnd.n954 0.152939
R12279 gnd.n956 gnd.n955 0.152939
R12280 gnd.n957 gnd.n956 0.152939
R12281 gnd.n962 gnd.n957 0.152939
R12282 gnd.n963 gnd.n962 0.152939
R12283 gnd.n964 gnd.n963 0.152939
R12284 gnd.n965 gnd.n964 0.152939
R12285 gnd.n970 gnd.n965 0.152939
R12286 gnd.n971 gnd.n970 0.152939
R12287 gnd.n972 gnd.n971 0.152939
R12288 gnd.n973 gnd.n972 0.152939
R12289 gnd.n978 gnd.n973 0.152939
R12290 gnd.n979 gnd.n978 0.152939
R12291 gnd.n980 gnd.n979 0.152939
R12292 gnd.n981 gnd.n980 0.152939
R12293 gnd.n986 gnd.n981 0.152939
R12294 gnd.n987 gnd.n986 0.152939
R12295 gnd.n988 gnd.n987 0.152939
R12296 gnd.n989 gnd.n988 0.152939
R12297 gnd.n994 gnd.n989 0.152939
R12298 gnd.n995 gnd.n994 0.152939
R12299 gnd.n996 gnd.n995 0.152939
R12300 gnd.n997 gnd.n996 0.152939
R12301 gnd.n1002 gnd.n997 0.152939
R12302 gnd.n1003 gnd.n1002 0.152939
R12303 gnd.n1004 gnd.n1003 0.152939
R12304 gnd.n1005 gnd.n1004 0.152939
R12305 gnd.n2304 gnd.n1005 0.152939
R12306 gnd.n2673 gnd.n2099 0.152939
R12307 gnd.n2674 gnd.n2673 0.152939
R12308 gnd.n2676 gnd.n2674 0.152939
R12309 gnd.n2676 gnd.n2675 0.152939
R12310 gnd.n2675 gnd.n2074 0.152939
R12311 gnd.n2703 gnd.n2074 0.152939
R12312 gnd.n2704 gnd.n2703 0.152939
R12313 gnd.n2706 gnd.n2704 0.152939
R12314 gnd.n2706 gnd.n2705 0.152939
R12315 gnd.n2705 gnd.n2049 0.152939
R12316 gnd.n2733 gnd.n2049 0.152939
R12317 gnd.n2734 gnd.n2733 0.152939
R12318 gnd.n2736 gnd.n2734 0.152939
R12319 gnd.n2736 gnd.n2735 0.152939
R12320 gnd.n2735 gnd.n2024 0.152939
R12321 gnd.n2763 gnd.n2024 0.152939
R12322 gnd.n2764 gnd.n2763 0.152939
R12323 gnd.n2769 gnd.n2764 0.152939
R12324 gnd.n2769 gnd.n2768 0.152939
R12325 gnd.n2768 gnd.n2767 0.152939
R12326 gnd.n2767 gnd.n2765 0.152939
R12327 gnd.n2765 gnd.n1998 0.152939
R12328 gnd.n2879 gnd.n1998 0.152939
R12329 gnd.n2880 gnd.n2879 0.152939
R12330 gnd.n2885 gnd.n2880 0.152939
R12331 gnd.n2885 gnd.n2884 0.152939
R12332 gnd.n2884 gnd.n2883 0.152939
R12333 gnd.n2883 gnd.n1973 0.152939
R12334 gnd.n2947 gnd.n1973 0.152939
R12335 gnd.n2948 gnd.n2947 0.152939
R12336 gnd.n2949 gnd.n2948 0.152939
R12337 gnd.n2949 gnd.n1951 0.152939
R12338 gnd.n2980 gnd.n1951 0.152939
R12339 gnd.n2981 gnd.n2980 0.152939
R12340 gnd.n2992 gnd.n2981 0.152939
R12341 gnd.n2992 gnd.n2991 0.152939
R12342 gnd.n2991 gnd.n2990 0.152939
R12343 gnd.n2990 gnd.n2982 0.152939
R12344 gnd.n2986 gnd.n2982 0.152939
R12345 gnd.n2986 gnd.n1911 0.152939
R12346 gnd.n3080 gnd.n1911 0.152939
R12347 gnd.n3081 gnd.n3080 0.152939
R12348 gnd.n3083 gnd.n3081 0.152939
R12349 gnd.n3083 gnd.n3082 0.152939
R12350 gnd.n3082 gnd.n1881 0.152939
R12351 gnd.n3116 gnd.n1881 0.152939
R12352 gnd.n3117 gnd.n3116 0.152939
R12353 gnd.n3122 gnd.n3117 0.152939
R12354 gnd.n3122 gnd.n3121 0.152939
R12355 gnd.n3121 gnd.n3120 0.152939
R12356 gnd.n3120 gnd.n1852 0.152939
R12357 gnd.n3164 gnd.n1852 0.152939
R12358 gnd.n3165 gnd.n3164 0.152939
R12359 gnd.n3170 gnd.n3165 0.152939
R12360 gnd.n3170 gnd.n3169 0.152939
R12361 gnd.n3169 gnd.n3168 0.152939
R12362 gnd.n3168 gnd.n1815 0.152939
R12363 gnd.n3252 gnd.n1815 0.152939
R12364 gnd.n3253 gnd.n3252 0.152939
R12365 gnd.n3255 gnd.n3253 0.152939
R12366 gnd.n3255 gnd.n3254 0.152939
R12367 gnd.n3254 gnd.n1789 0.152939
R12368 gnd.n3288 gnd.n1789 0.152939
R12369 gnd.n3289 gnd.n3288 0.152939
R12370 gnd.n3296 gnd.n3289 0.152939
R12371 gnd.n3296 gnd.n3295 0.152939
R12372 gnd.n3295 gnd.n3294 0.152939
R12373 gnd.n3294 gnd.n1762 0.152939
R12374 gnd.n3338 gnd.n1762 0.152939
R12375 gnd.n3339 gnd.n3338 0.152939
R12376 gnd.n3344 gnd.n3339 0.152939
R12377 gnd.n3344 gnd.n3343 0.152939
R12378 gnd.n3343 gnd.n3342 0.152939
R12379 gnd.n3342 gnd.n1728 0.152939
R12380 gnd.n3409 gnd.n1728 0.152939
R12381 gnd.n3410 gnd.n3409 0.152939
R12382 gnd.n3412 gnd.n3410 0.152939
R12383 gnd.n3412 gnd.n3411 0.152939
R12384 gnd.n3411 gnd.n1636 0.152939
R12385 gnd.n3557 gnd.n1636 0.152939
R12386 gnd.n3558 gnd.n3557 0.152939
R12387 gnd.n3559 gnd.n3558 0.152939
R12388 gnd.n3559 gnd.n1623 0.152939
R12389 gnd.n3579 gnd.n1623 0.152939
R12390 gnd.n3580 gnd.n3579 0.152939
R12391 gnd.n3581 gnd.n3580 0.152939
R12392 gnd.n3581 gnd.n1612 0.152939
R12393 gnd.n3599 gnd.n1612 0.152939
R12394 gnd.n3600 gnd.n3599 0.152939
R12395 gnd.n3601 gnd.n3600 0.152939
R12396 gnd.n3601 gnd.n1599 0.152939
R12397 gnd.n3619 gnd.n1599 0.152939
R12398 gnd.n3620 gnd.n3619 0.152939
R12399 gnd.n3621 gnd.n3620 0.152939
R12400 gnd.n3621 gnd.n1586 0.152939
R12401 gnd.n3639 gnd.n1586 0.152939
R12402 gnd.n3640 gnd.n3639 0.152939
R12403 gnd.n3642 gnd.n3640 0.152939
R12404 gnd.n3642 gnd.n3641 0.152939
R12405 gnd.n3641 gnd.n453 0.152939
R12406 gnd.n6358 gnd.n453 0.152939
R12407 gnd.n2506 gnd.n2505 0.152939
R12408 gnd.n2507 gnd.n2506 0.152939
R12409 gnd.n2507 gnd.n2389 0.152939
R12410 gnd.n2512 gnd.n2389 0.152939
R12411 gnd.n2513 gnd.n2512 0.152939
R12412 gnd.n2514 gnd.n2513 0.152939
R12413 gnd.n2514 gnd.n2386 0.152939
R12414 gnd.n2519 gnd.n2386 0.152939
R12415 gnd.n2520 gnd.n2519 0.152939
R12416 gnd.n2521 gnd.n2520 0.152939
R12417 gnd.n2521 gnd.n2383 0.152939
R12418 gnd.n2526 gnd.n2383 0.152939
R12419 gnd.n2527 gnd.n2526 0.152939
R12420 gnd.n2528 gnd.n2527 0.152939
R12421 gnd.n2528 gnd.n2319 0.152939
R12422 gnd.n2546 gnd.n2319 0.152939
R12423 gnd.n2547 gnd.n2546 0.152939
R12424 gnd.n2562 gnd.n2547 0.152939
R12425 gnd.n2562 gnd.n2561 0.152939
R12426 gnd.n2561 gnd.n2560 0.152939
R12427 gnd.n2664 gnd.n2108 0.152939
R12428 gnd.n2657 gnd.n2108 0.152939
R12429 gnd.n2657 gnd.n2656 0.152939
R12430 gnd.n2656 gnd.n2655 0.152939
R12431 gnd.n2655 gnd.n2128 0.152939
R12432 gnd.n2651 gnd.n2128 0.152939
R12433 gnd.n2667 gnd.n2665 0.152939
R12434 gnd.n2667 gnd.n2666 0.152939
R12435 gnd.n2666 gnd.n2083 0.152939
R12436 gnd.n2694 gnd.n2083 0.152939
R12437 gnd.n2695 gnd.n2694 0.152939
R12438 gnd.n2697 gnd.n2695 0.152939
R12439 gnd.n2697 gnd.n2696 0.152939
R12440 gnd.n2696 gnd.n2058 0.152939
R12441 gnd.n2724 gnd.n2058 0.152939
R12442 gnd.n2725 gnd.n2724 0.152939
R12443 gnd.n2727 gnd.n2725 0.152939
R12444 gnd.n2727 gnd.n2726 0.152939
R12445 gnd.n2726 gnd.n2032 0.152939
R12446 gnd.n2754 gnd.n2032 0.152939
R12447 gnd.n2755 gnd.n2754 0.152939
R12448 gnd.n2757 gnd.n2755 0.152939
R12449 gnd.n2757 gnd.n2756 0.152939
R12450 gnd.n2756 gnd.n2008 0.152939
R12451 gnd.n2799 gnd.n2008 0.152939
R12452 gnd.n2800 gnd.n2799 0.152939
R12453 gnd.n2802 gnd.n2800 0.152939
R12454 gnd.n2802 gnd.n2801 0.152939
R12455 gnd.n2801 gnd.n1479 0.152939
R12456 gnd.n3775 gnd.n1479 0.152939
R12457 gnd.n3775 gnd.n3774 0.152939
R12458 gnd.n3774 gnd.n3773 0.152939
R12459 gnd.n3773 gnd.n1480 0.152939
R12460 gnd.n3769 gnd.n1480 0.152939
R12461 gnd.n3769 gnd.n3768 0.152939
R12462 gnd.n3768 gnd.n3767 0.152939
R12463 gnd.n3767 gnd.n1485 0.152939
R12464 gnd.n3763 gnd.n1485 0.152939
R12465 gnd.n3763 gnd.n3762 0.152939
R12466 gnd.n3762 gnd.n3761 0.152939
R12467 gnd.n3761 gnd.n1490 0.152939
R12468 gnd.n3757 gnd.n1490 0.152939
R12469 gnd.n3757 gnd.n3756 0.152939
R12470 gnd.n3756 gnd.n3755 0.152939
R12471 gnd.n3755 gnd.n1495 0.152939
R12472 gnd.n3751 gnd.n1495 0.152939
R12473 gnd.n3751 gnd.n3750 0.152939
R12474 gnd.n3750 gnd.n3749 0.152939
R12475 gnd.n3749 gnd.n1500 0.152939
R12476 gnd.n3745 gnd.n1500 0.152939
R12477 gnd.n3745 gnd.n3744 0.152939
R12478 gnd.n3744 gnd.n3743 0.152939
R12479 gnd.n3743 gnd.n1505 0.152939
R12480 gnd.n3739 gnd.n1505 0.152939
R12481 gnd.n3739 gnd.n3738 0.152939
R12482 gnd.n3738 gnd.n3737 0.152939
R12483 gnd.n3737 gnd.n1510 0.152939
R12484 gnd.n3733 gnd.n1510 0.152939
R12485 gnd.n3733 gnd.n3732 0.152939
R12486 gnd.n3732 gnd.n3731 0.152939
R12487 gnd.n3731 gnd.n1515 0.152939
R12488 gnd.n3727 gnd.n1515 0.152939
R12489 gnd.n3727 gnd.n3726 0.152939
R12490 gnd.n3726 gnd.n3725 0.152939
R12491 gnd.n3725 gnd.n1520 0.152939
R12492 gnd.n3721 gnd.n1520 0.152939
R12493 gnd.n3721 gnd.n3720 0.152939
R12494 gnd.n3720 gnd.n3719 0.152939
R12495 gnd.n3719 gnd.n1525 0.152939
R12496 gnd.n3715 gnd.n1525 0.152939
R12497 gnd.n3715 gnd.n3714 0.152939
R12498 gnd.n3714 gnd.n3713 0.152939
R12499 gnd.n3713 gnd.n1530 0.152939
R12500 gnd.n3709 gnd.n1530 0.152939
R12501 gnd.n3709 gnd.n3708 0.152939
R12502 gnd.n3708 gnd.n3707 0.152939
R12503 gnd.n3707 gnd.n1535 0.152939
R12504 gnd.n3703 gnd.n1535 0.152939
R12505 gnd.n3703 gnd.n3702 0.152939
R12506 gnd.n3702 gnd.n3701 0.152939
R12507 gnd.n3701 gnd.n1540 0.152939
R12508 gnd.n3697 gnd.n1540 0.152939
R12509 gnd.n3697 gnd.n3696 0.152939
R12510 gnd.n3696 gnd.n3695 0.152939
R12511 gnd.n3695 gnd.n1545 0.152939
R12512 gnd.n3691 gnd.n1545 0.152939
R12513 gnd.n3691 gnd.n3690 0.152939
R12514 gnd.n3690 gnd.n3689 0.152939
R12515 gnd.n3689 gnd.n1550 0.152939
R12516 gnd.n3685 gnd.n1550 0.152939
R12517 gnd.n3685 gnd.n3684 0.152939
R12518 gnd.n3684 gnd.n3683 0.152939
R12519 gnd.n3683 gnd.n1555 0.152939
R12520 gnd.n3679 gnd.n1555 0.152939
R12521 gnd.n3679 gnd.n3678 0.152939
R12522 gnd.n3678 gnd.n3677 0.152939
R12523 gnd.n3677 gnd.n1560 0.152939
R12524 gnd.n3673 gnd.n1560 0.152939
R12525 gnd.n3673 gnd.n3672 0.152939
R12526 gnd.n3672 gnd.n3671 0.152939
R12527 gnd.n3671 gnd.n1565 0.152939
R12528 gnd.n3667 gnd.n1565 0.152939
R12529 gnd.n3667 gnd.n3666 0.152939
R12530 gnd.n3666 gnd.n3665 0.152939
R12531 gnd.n3665 gnd.n1570 0.152939
R12532 gnd.n1570 gnd.n462 0.152939
R12533 gnd.n6352 gnd.n462 0.152939
R12534 gnd.n6351 gnd.n463 0.152939
R12535 gnd.n6347 gnd.n463 0.152939
R12536 gnd.n6347 gnd.n6346 0.152939
R12537 gnd.n6346 gnd.n6345 0.152939
R12538 gnd.n6345 gnd.n467 0.152939
R12539 gnd.n467 gnd.n389 0.152939
R12540 gnd.n6543 gnd.n271 0.152939
R12541 gnd.n6544 gnd.n6543 0.152939
R12542 gnd.n6546 gnd.n6544 0.152939
R12543 gnd.n6546 gnd.n6545 0.152939
R12544 gnd.n6545 gnd.n243 0.152939
R12545 gnd.n6578 gnd.n243 0.152939
R12546 gnd.n6579 gnd.n6578 0.152939
R12547 gnd.n6591 gnd.n6579 0.152939
R12548 gnd.n6591 gnd.n6590 0.152939
R12549 gnd.n6590 gnd.n6589 0.152939
R12550 gnd.n6589 gnd.n6580 0.152939
R12551 gnd.n6585 gnd.n6580 0.152939
R12552 gnd.n6585 gnd.n6584 0.152939
R12553 gnd.n6584 gnd.n198 0.152939
R12554 gnd.n6642 gnd.n198 0.152939
R12555 gnd.n6643 gnd.n6642 0.152939
R12556 gnd.n6649 gnd.n6643 0.152939
R12557 gnd.n6649 gnd.n6648 0.152939
R12558 gnd.n6648 gnd.n6647 0.152939
R12559 gnd.n6647 gnd.n67 0.152939
R12560 gnd.n7112 gnd.n7111 0.145814
R12561 gnd.n2499 gnd.n2392 0.145814
R12562 gnd.n2505 gnd.n2392 0.145814
R12563 gnd.n7112 gnd.n67 0.145814
R12564 gnd.n2651 gnd.n2650 0.128549
R12565 gnd.n6417 gnd.n389 0.128549
R12566 gnd.n4422 gnd.n0 0.127478
R12567 gnd.n5002 gnd.n5001 0.0767195
R12568 gnd.n5001 gnd.n5000 0.0767195
R12569 gnd.n2650 gnd.n2134 0.063
R12570 gnd.n6418 gnd.n6417 0.063
R12571 gnd.n6418 gnd.n388 0.0538288
R12572 gnd.n7049 gnd.n7048 0.0538288
R12573 gnd.n4038 gnd.n4037 0.0538288
R12574 gnd.n2536 gnd.n2134 0.0538288
R12575 gnd.n5568 gnd.n4184 0.0477147
R12576 gnd.n4765 gnd.n4653 0.0442063
R12577 gnd.n4766 gnd.n4765 0.0442063
R12578 gnd.n4767 gnd.n4766 0.0442063
R12579 gnd.n4767 gnd.n4642 0.0442063
R12580 gnd.n4781 gnd.n4642 0.0442063
R12581 gnd.n4782 gnd.n4781 0.0442063
R12582 gnd.n4783 gnd.n4782 0.0442063
R12583 gnd.n4783 gnd.n4629 0.0442063
R12584 gnd.n4827 gnd.n4629 0.0442063
R12585 gnd.n4828 gnd.n4827 0.0442063
R12586 gnd.n505 gnd.n388 0.0344674
R12587 gnd.n506 gnd.n505 0.0344674
R12588 gnd.n506 gnd.n265 0.0344674
R12589 gnd.n265 gnd.n262 0.0344674
R12590 gnd.n263 gnd.n262 0.0344674
R12591 gnd.n6557 gnd.n263 0.0344674
R12592 gnd.n6558 gnd.n6557 0.0344674
R12593 gnd.n6558 gnd.n237 0.0344674
R12594 gnd.n237 gnd.n235 0.0344674
R12595 gnd.n6599 gnd.n235 0.0344674
R12596 gnd.n6600 gnd.n6599 0.0344674
R12597 gnd.n6600 gnd.n219 0.0344674
R12598 gnd.n219 gnd.n216 0.0344674
R12599 gnd.n217 gnd.n216 0.0344674
R12600 gnd.n6621 gnd.n217 0.0344674
R12601 gnd.n6622 gnd.n6621 0.0344674
R12602 gnd.n6622 gnd.n191 0.0344674
R12603 gnd.n6658 gnd.n191 0.0344674
R12604 gnd.n6658 gnd.n174 0.0344674
R12605 gnd.n6675 gnd.n174 0.0344674
R12606 gnd.n6676 gnd.n6675 0.0344674
R12607 gnd.n6676 gnd.n168 0.0344674
R12608 gnd.n6684 gnd.n168 0.0344674
R12609 gnd.n6685 gnd.n6684 0.0344674
R12610 gnd.n6685 gnd.n90 0.0344674
R12611 gnd.n91 gnd.n90 0.0344674
R12612 gnd.n92 gnd.n91 0.0344674
R12613 gnd.n6692 gnd.n92 0.0344674
R12614 gnd.n6692 gnd.n109 0.0344674
R12615 gnd.n110 gnd.n109 0.0344674
R12616 gnd.n111 gnd.n110 0.0344674
R12617 gnd.n6699 gnd.n111 0.0344674
R12618 gnd.n6699 gnd.n128 0.0344674
R12619 gnd.n129 gnd.n128 0.0344674
R12620 gnd.n130 gnd.n129 0.0344674
R12621 gnd.n6706 gnd.n130 0.0344674
R12622 gnd.n6706 gnd.n147 0.0344674
R12623 gnd.n148 gnd.n147 0.0344674
R12624 gnd.n149 gnd.n148 0.0344674
R12625 gnd.n6713 gnd.n149 0.0344674
R12626 gnd.n6713 gnd.n166 0.0344674
R12627 gnd.n7049 gnd.n166 0.0344674
R12628 gnd.n4830 gnd.n4563 0.0344674
R12629 gnd.n4037 gnd.n1131 0.0344674
R12630 gnd.n2322 gnd.n1131 0.0344674
R12631 gnd.n2322 gnd.n1152 0.0344674
R12632 gnd.n1153 gnd.n1152 0.0344674
R12633 gnd.n1154 gnd.n1153 0.0344674
R12634 gnd.n2329 gnd.n1154 0.0344674
R12635 gnd.n2329 gnd.n1170 0.0344674
R12636 gnd.n1171 gnd.n1170 0.0344674
R12637 gnd.n1172 gnd.n1171 0.0344674
R12638 gnd.n2336 gnd.n1172 0.0344674
R12639 gnd.n2336 gnd.n1188 0.0344674
R12640 gnd.n1189 gnd.n1188 0.0344674
R12641 gnd.n1190 gnd.n1189 0.0344674
R12642 gnd.n2343 gnd.n1190 0.0344674
R12643 gnd.n2343 gnd.n1208 0.0344674
R12644 gnd.n1209 gnd.n1208 0.0344674
R12645 gnd.n1210 gnd.n1209 0.0344674
R12646 gnd.n2350 gnd.n1210 0.0344674
R12647 gnd.n2350 gnd.n1226 0.0344674
R12648 gnd.n1227 gnd.n1226 0.0344674
R12649 gnd.n1228 gnd.n1227 0.0344674
R12650 gnd.n2357 gnd.n1228 0.0344674
R12651 gnd.n2357 gnd.n1246 0.0344674
R12652 gnd.n1247 gnd.n1246 0.0344674
R12653 gnd.n1248 gnd.n1247 0.0344674
R12654 gnd.n2364 gnd.n1248 0.0344674
R12655 gnd.n2364 gnd.n1264 0.0344674
R12656 gnd.n1265 gnd.n1264 0.0344674
R12657 gnd.n1266 gnd.n1265 0.0344674
R12658 gnd.n2371 gnd.n1266 0.0344674
R12659 gnd.n2371 gnd.n1284 0.0344674
R12660 gnd.n1285 gnd.n1284 0.0344674
R12661 gnd.n1286 gnd.n1285 0.0344674
R12662 gnd.n2378 gnd.n1286 0.0344674
R12663 gnd.n2378 gnd.n1304 0.0344674
R12664 gnd.n1305 gnd.n1304 0.0344674
R12665 gnd.n1306 gnd.n1305 0.0344674
R12666 gnd.n2535 gnd.n1306 0.0344674
R12667 gnd.n2535 gnd.n1325 0.0344674
R12668 gnd.n1326 gnd.n1325 0.0344674
R12669 gnd.n1327 gnd.n1326 0.0344674
R12670 gnd.n2536 gnd.n1327 0.0344674
R12671 gnd.n2649 gnd.n2648 0.0343753
R12672 gnd.n6416 gnd.n390 0.0343753
R12673 gnd.n2559 gnd.n2558 0.0296328
R12674 gnd.n6361 gnd.n6360 0.0296328
R12675 gnd.n4850 gnd.n4849 0.0269946
R12676 gnd.n4852 gnd.n4851 0.0269946
R12677 gnd.n4558 gnd.n4556 0.0269946
R12678 gnd.n4862 gnd.n4860 0.0269946
R12679 gnd.n4861 gnd.n4537 0.0269946
R12680 gnd.n4881 gnd.n4880 0.0269946
R12681 gnd.n4883 gnd.n4882 0.0269946
R12682 gnd.n4532 gnd.n4531 0.0269946
R12683 gnd.n4893 gnd.n4527 0.0269946
R12684 gnd.n4892 gnd.n4529 0.0269946
R12685 gnd.n4528 gnd.n4510 0.0269946
R12686 gnd.n4913 gnd.n4511 0.0269946
R12687 gnd.n4912 gnd.n4512 0.0269946
R12688 gnd.n4946 gnd.n4487 0.0269946
R12689 gnd.n4948 gnd.n4947 0.0269946
R12690 gnd.n4949 gnd.n4434 0.0269946
R12691 gnd.n4482 gnd.n4435 0.0269946
R12692 gnd.n4484 gnd.n4436 0.0269946
R12693 gnd.n4959 gnd.n4958 0.0269946
R12694 gnd.n4961 gnd.n4960 0.0269946
R12695 gnd.n4962 gnd.n4456 0.0269946
R12696 gnd.n4964 gnd.n4457 0.0269946
R12697 gnd.n4967 gnd.n4458 0.0269946
R12698 gnd.n4970 gnd.n4969 0.0269946
R12699 gnd.n4972 gnd.n4971 0.0269946
R12700 gnd.n5037 gnd.n4357 0.0269946
R12701 gnd.n5039 gnd.n5038 0.0269946
R12702 gnd.n5048 gnd.n4350 0.0269946
R12703 gnd.n5050 gnd.n5049 0.0269946
R12704 gnd.n5051 gnd.n4348 0.0269946
R12705 gnd.n5058 gnd.n5054 0.0269946
R12706 gnd.n5057 gnd.n5056 0.0269946
R12707 gnd.n5055 gnd.n4327 0.0269946
R12708 gnd.n5080 gnd.n4328 0.0269946
R12709 gnd.n5079 gnd.n4329 0.0269946
R12710 gnd.n5122 gnd.n4302 0.0269946
R12711 gnd.n5124 gnd.n5123 0.0269946
R12712 gnd.n5133 gnd.n4295 0.0269946
R12713 gnd.n5135 gnd.n5134 0.0269946
R12714 gnd.n5136 gnd.n4293 0.0269946
R12715 gnd.n5143 gnd.n5139 0.0269946
R12716 gnd.n5142 gnd.n5141 0.0269946
R12717 gnd.n5140 gnd.n4272 0.0269946
R12718 gnd.n5165 gnd.n4273 0.0269946
R12719 gnd.n5164 gnd.n4274 0.0269946
R12720 gnd.n5211 gnd.n4248 0.0269946
R12721 gnd.n5213 gnd.n5212 0.0269946
R12722 gnd.n5222 gnd.n4241 0.0269946
R12723 gnd.n5481 gnd.n4239 0.0269946
R12724 gnd.n5486 gnd.n5484 0.0269946
R12725 gnd.n5485 gnd.n4220 0.0269946
R12726 gnd.n5510 gnd.n5509 0.0269946
R12727 gnd.n2645 gnd.n2135 0.022519
R12728 gnd.n2644 gnd.n2139 0.022519
R12729 gnd.n2641 gnd.n2640 0.022519
R12730 gnd.n2637 gnd.n2145 0.022519
R12731 gnd.n2636 gnd.n2151 0.022519
R12732 gnd.n2633 gnd.n2632 0.022519
R12733 gnd.n2629 gnd.n2155 0.022519
R12734 gnd.n2628 gnd.n2159 0.022519
R12735 gnd.n2625 gnd.n2624 0.022519
R12736 gnd.n2621 gnd.n2165 0.022519
R12737 gnd.n2620 gnd.n2171 0.022519
R12738 gnd.n2617 gnd.n2616 0.022519
R12739 gnd.n2613 gnd.n2175 0.022519
R12740 gnd.n2612 gnd.n2179 0.022519
R12741 gnd.n2609 gnd.n2608 0.022519
R12742 gnd.n2605 gnd.n2185 0.022519
R12743 gnd.n2604 gnd.n2192 0.022519
R12744 gnd.n2551 gnd.n2196 0.022519
R12745 gnd.n2558 gnd.n2198 0.022519
R12746 gnd.n6412 gnd.n396 0.022519
R12747 gnd.n6411 gnd.n397 0.022519
R12748 gnd.n6408 gnd.n6407 0.022519
R12749 gnd.n6404 gnd.n402 0.022519
R12750 gnd.n6403 gnd.n406 0.022519
R12751 gnd.n6400 gnd.n6399 0.022519
R12752 gnd.n6396 gnd.n412 0.022519
R12753 gnd.n6395 gnd.n416 0.022519
R12754 gnd.n6392 gnd.n6391 0.022519
R12755 gnd.n6388 gnd.n420 0.022519
R12756 gnd.n6387 gnd.n424 0.022519
R12757 gnd.n6384 gnd.n6383 0.022519
R12758 gnd.n6380 gnd.n430 0.022519
R12759 gnd.n6379 gnd.n434 0.022519
R12760 gnd.n6376 gnd.n6375 0.022519
R12761 gnd.n6372 gnd.n438 0.022519
R12762 gnd.n6371 gnd.n444 0.022519
R12763 gnd.n6365 gnd.n6364 0.022519
R12764 gnd.n6361 gnd.n448 0.022519
R12765 gnd.n6360 gnd.n6359 0.0218415
R12766 gnd.n2559 gnd.n2548 0.0218415
R12767 gnd.n4830 gnd.n4829 0.0202011
R12768 gnd.n4829 gnd.n4828 0.0148637
R12769 gnd.n5479 gnd.n5223 0.0144266
R12770 gnd.n5480 gnd.n5479 0.0130679
R12771 gnd.n2648 gnd.n2135 0.0123564
R12772 gnd.n2645 gnd.n2644 0.0123564
R12773 gnd.n2641 gnd.n2139 0.0123564
R12774 gnd.n2640 gnd.n2145 0.0123564
R12775 gnd.n2637 gnd.n2636 0.0123564
R12776 gnd.n2633 gnd.n2151 0.0123564
R12777 gnd.n2632 gnd.n2155 0.0123564
R12778 gnd.n2629 gnd.n2628 0.0123564
R12779 gnd.n2625 gnd.n2159 0.0123564
R12780 gnd.n2624 gnd.n2165 0.0123564
R12781 gnd.n2621 gnd.n2620 0.0123564
R12782 gnd.n2617 gnd.n2171 0.0123564
R12783 gnd.n2616 gnd.n2175 0.0123564
R12784 gnd.n2613 gnd.n2612 0.0123564
R12785 gnd.n2609 gnd.n2179 0.0123564
R12786 gnd.n2608 gnd.n2185 0.0123564
R12787 gnd.n2605 gnd.n2604 0.0123564
R12788 gnd.n2196 gnd.n2192 0.0123564
R12789 gnd.n2551 gnd.n2198 0.0123564
R12790 gnd.n396 gnd.n390 0.0123564
R12791 gnd.n6412 gnd.n6411 0.0123564
R12792 gnd.n6408 gnd.n397 0.0123564
R12793 gnd.n6407 gnd.n402 0.0123564
R12794 gnd.n6404 gnd.n6403 0.0123564
R12795 gnd.n6400 gnd.n406 0.0123564
R12796 gnd.n6399 gnd.n412 0.0123564
R12797 gnd.n6396 gnd.n6395 0.0123564
R12798 gnd.n6392 gnd.n416 0.0123564
R12799 gnd.n6391 gnd.n420 0.0123564
R12800 gnd.n6388 gnd.n6387 0.0123564
R12801 gnd.n6384 gnd.n424 0.0123564
R12802 gnd.n6383 gnd.n430 0.0123564
R12803 gnd.n6380 gnd.n6379 0.0123564
R12804 gnd.n6376 gnd.n434 0.0123564
R12805 gnd.n6375 gnd.n438 0.0123564
R12806 gnd.n6372 gnd.n6371 0.0123564
R12807 gnd.n6365 gnd.n444 0.0123564
R12808 gnd.n6364 gnd.n448 0.0123564
R12809 gnd.n4849 gnd.n4563 0.00797283
R12810 gnd.n4851 gnd.n4850 0.00797283
R12811 gnd.n4852 gnd.n4558 0.00797283
R12812 gnd.n4860 gnd.n4556 0.00797283
R12813 gnd.n4862 gnd.n4861 0.00797283
R12814 gnd.n4880 gnd.n4537 0.00797283
R12815 gnd.n4882 gnd.n4881 0.00797283
R12816 gnd.n4883 gnd.n4532 0.00797283
R12817 gnd.n4531 gnd.n4527 0.00797283
R12818 gnd.n4893 gnd.n4892 0.00797283
R12819 gnd.n4529 gnd.n4528 0.00797283
R12820 gnd.n4511 gnd.n4510 0.00797283
R12821 gnd.n4913 gnd.n4912 0.00797283
R12822 gnd.n4512 gnd.n4487 0.00797283
R12823 gnd.n4947 gnd.n4946 0.00797283
R12824 gnd.n4949 gnd.n4948 0.00797283
R12825 gnd.n4482 gnd.n4434 0.00797283
R12826 gnd.n4484 gnd.n4435 0.00797283
R12827 gnd.n4958 gnd.n4436 0.00797283
R12828 gnd.n4960 gnd.n4959 0.00797283
R12829 gnd.n4962 gnd.n4961 0.00797283
R12830 gnd.n4964 gnd.n4456 0.00797283
R12831 gnd.n4967 gnd.n4457 0.00797283
R12832 gnd.n4969 gnd.n4458 0.00797283
R12833 gnd.n4972 gnd.n4970 0.00797283
R12834 gnd.n4971 gnd.n4357 0.00797283
R12835 gnd.n5039 gnd.n5037 0.00797283
R12836 gnd.n5038 gnd.n4350 0.00797283
R12837 gnd.n5049 gnd.n5048 0.00797283
R12838 gnd.n5051 gnd.n5050 0.00797283
R12839 gnd.n5054 gnd.n4348 0.00797283
R12840 gnd.n5058 gnd.n5057 0.00797283
R12841 gnd.n5056 gnd.n5055 0.00797283
R12842 gnd.n4328 gnd.n4327 0.00797283
R12843 gnd.n5080 gnd.n5079 0.00797283
R12844 gnd.n4329 gnd.n4302 0.00797283
R12845 gnd.n5124 gnd.n5122 0.00797283
R12846 gnd.n5123 gnd.n4295 0.00797283
R12847 gnd.n5134 gnd.n5133 0.00797283
R12848 gnd.n5136 gnd.n5135 0.00797283
R12849 gnd.n5139 gnd.n4293 0.00797283
R12850 gnd.n5143 gnd.n5142 0.00797283
R12851 gnd.n5141 gnd.n5140 0.00797283
R12852 gnd.n4273 gnd.n4272 0.00797283
R12853 gnd.n5165 gnd.n5164 0.00797283
R12854 gnd.n4274 gnd.n4248 0.00797283
R12855 gnd.n5213 gnd.n5211 0.00797283
R12856 gnd.n5212 gnd.n4241 0.00797283
R12857 gnd.n5223 gnd.n5222 0.00797283
R12858 gnd.n5481 gnd.n5480 0.00797283
R12859 gnd.n5484 gnd.n4239 0.00797283
R12860 gnd.n5486 gnd.n5485 0.00797283
R12861 gnd.n5509 gnd.n4220 0.00797283
R12862 gnd.n5510 gnd.n4184 0.00797283
R12863 gnd.n2650 gnd.n2649 0.00592005
R12864 gnd.n6417 gnd.n6416 0.00592005
R12865 gnd.n6635 gnd.n183 0.00417647
R12866 gnd.n6664 gnd.n183 0.00417647
R12867 gnd.n6665 gnd.n6664 0.00417647
R12868 gnd.n6666 gnd.n6665 0.00417647
R12869 gnd.n6668 gnd.n6666 0.00417647
R12870 gnd.n6668 gnd.n6667 0.00417647
R12871 gnd.n6667 gnd.n79 0.00417647
R12872 gnd.n80 gnd.n79 0.00417647
R12873 gnd.n81 gnd.n80 0.00417647
R12874 gnd.n98 gnd.n81 0.00417647
R12875 gnd.n1217 gnd.n1216 0.00417647
R12876 gnd.n1218 gnd.n1217 0.00417647
R12877 gnd.n1219 gnd.n1218 0.00417647
R12878 gnd.n1236 gnd.n1219 0.00417647
R12879 gnd.n1237 gnd.n1236 0.00417647
R12880 gnd.n1238 gnd.n1237 0.00417647
R12881 gnd.n1239 gnd.n1238 0.00417647
R12882 gnd.n1255 gnd.n1239 0.00417647
R12883 gnd.n1256 gnd.n1255 0.00417647
R12884 gnd.n1257 gnd.n1256 0.00417647
R12885 commonsourceibias.n25 commonsourceibias.t34 230.006
R12886 commonsourceibias.n91 commonsourceibias.t95 230.006
R12887 commonsourceibias.n218 commonsourceibias.t117 230.006
R12888 commonsourceibias.n154 commonsourceibias.t97 230.006
R12889 commonsourceibias.n322 commonsourceibias.t4 230.006
R12890 commonsourceibias.n281 commonsourceibias.t70 230.006
R12891 commonsourceibias.n483 commonsourceibias.t55 230.006
R12892 commonsourceibias.n419 commonsourceibias.t80 230.006
R12893 commonsourceibias.n70 commonsourceibias.t16 207.983
R12894 commonsourceibias.n136 commonsourceibias.t56 207.983
R12895 commonsourceibias.n263 commonsourceibias.t111 207.983
R12896 commonsourceibias.n199 commonsourceibias.t89 207.983
R12897 commonsourceibias.n368 commonsourceibias.t26 207.983
R12898 commonsourceibias.n402 commonsourceibias.t114 207.983
R12899 commonsourceibias.n529 commonsourceibias.t51 207.983
R12900 commonsourceibias.n465 commonsourceibias.t74 207.983
R12901 commonsourceibias.n10 commonsourceibias.t30 168.701
R12902 commonsourceibias.n63 commonsourceibias.t2 168.701
R12903 commonsourceibias.n57 commonsourceibias.t22 168.701
R12904 commonsourceibias.n16 commonsourceibias.t42 168.701
R12905 commonsourceibias.n49 commonsourceibias.t18 168.701
R12906 commonsourceibias.n43 commonsourceibias.t32 168.701
R12907 commonsourceibias.n19 commonsourceibias.t40 168.701
R12908 commonsourceibias.n21 commonsourceibias.t24 168.701
R12909 commonsourceibias.n23 commonsourceibias.t44 168.701
R12910 commonsourceibias.n26 commonsourceibias.t6 168.701
R12911 commonsourceibias.n1 commonsourceibias.t109 168.701
R12912 commonsourceibias.n129 commonsourceibias.t69 168.701
R12913 commonsourceibias.n123 commonsourceibias.t119 168.701
R12914 commonsourceibias.n7 commonsourceibias.t85 168.701
R12915 commonsourceibias.n115 commonsourceibias.t54 168.701
R12916 commonsourceibias.n109 commonsourceibias.t100 168.701
R12917 commonsourceibias.n85 commonsourceibias.t87 168.701
R12918 commonsourceibias.n87 commonsourceibias.t115 168.701
R12919 commonsourceibias.n89 commonsourceibias.t79 168.701
R12920 commonsourceibias.n92 commonsourceibias.t66 168.701
R12921 commonsourceibias.n219 commonsourceibias.t75 168.701
R12922 commonsourceibias.n216 commonsourceibias.t59 168.701
R12923 commonsourceibias.n214 commonsourceibias.t49 168.701
R12924 commonsourceibias.n212 commonsourceibias.t84 168.701
R12925 commonsourceibias.n236 commonsourceibias.t93 168.701
R12926 commonsourceibias.n242 commonsourceibias.t52 168.701
R12927 commonsourceibias.n209 commonsourceibias.t118 168.701
R12928 commonsourceibias.n250 commonsourceibias.t104 168.701
R12929 commonsourceibias.n256 commonsourceibias.t60 168.701
R12930 commonsourceibias.n203 commonsourceibias.t50 168.701
R12931 commonsourceibias.n139 commonsourceibias.t106 168.701
R12932 commonsourceibias.n192 commonsourceibias.t101 168.701
R12933 commonsourceibias.n186 commonsourceibias.t88 168.701
R12934 commonsourceibias.n145 commonsourceibias.t105 168.701
R12935 commonsourceibias.n178 commonsourceibias.t99 168.701
R12936 commonsourceibias.n172 commonsourceibias.t86 168.701
R12937 commonsourceibias.n148 commonsourceibias.t108 168.701
R12938 commonsourceibias.n150 commonsourceibias.t98 168.701
R12939 commonsourceibias.n152 commonsourceibias.t112 168.701
R12940 commonsourceibias.n155 commonsourceibias.t107 168.701
R12941 commonsourceibias.n323 commonsourceibias.t14 168.701
R12942 commonsourceibias.n320 commonsourceibias.t12 168.701
R12943 commonsourceibias.n318 commonsourceibias.t38 168.701
R12944 commonsourceibias.n316 commonsourceibias.t8 168.701
R12945 commonsourceibias.n340 commonsourceibias.t0 168.701
R12946 commonsourceibias.n346 commonsourceibias.t28 168.701
R12947 commonsourceibias.n348 commonsourceibias.t10 168.701
R12948 commonsourceibias.n355 commonsourceibias.t36 168.701
R12949 commonsourceibias.n361 commonsourceibias.t20 168.701
R12950 commonsourceibias.n308 commonsourceibias.t46 168.701
R12951 commonsourceibias.n267 commonsourceibias.t78 168.701
R12952 commonsourceibias.n395 commonsourceibias.t53 168.701
R12953 commonsourceibias.n389 commonsourceibias.t94 168.701
R12954 commonsourceibias.n382 commonsourceibias.t64 168.701
R12955 commonsourceibias.n380 commonsourceibias.t113 168.701
R12956 commonsourceibias.n282 commonsourceibias.t58 168.701
R12957 commonsourceibias.n279 commonsourceibias.t63 168.701
R12958 commonsourceibias.n277 commonsourceibias.t92 168.701
R12959 commonsourceibias.n275 commonsourceibias.t65 168.701
R12960 commonsourceibias.n299 commonsourceibias.t76 168.701
R12961 commonsourceibias.n484 commonsourceibias.t68 168.701
R12962 commonsourceibias.n481 commonsourceibias.t72 168.701
R12963 commonsourceibias.n479 commonsourceibias.t61 168.701
R12964 commonsourceibias.n477 commonsourceibias.t110 168.701
R12965 commonsourceibias.n501 commonsourceibias.t77 168.701
R12966 commonsourceibias.n507 commonsourceibias.t67 168.701
R12967 commonsourceibias.n509 commonsourceibias.t57 168.701
R12968 commonsourceibias.n516 commonsourceibias.t48 168.701
R12969 commonsourceibias.n522 commonsourceibias.t71 168.701
R12970 commonsourceibias.n469 commonsourceibias.t62 168.701
R12971 commonsourceibias.n420 commonsourceibias.t116 168.701
R12972 commonsourceibias.n417 commonsourceibias.t102 168.701
R12973 commonsourceibias.n415 commonsourceibias.t81 168.701
R12974 commonsourceibias.n413 commonsourceibias.t96 168.701
R12975 commonsourceibias.n437 commonsourceibias.t103 168.701
R12976 commonsourceibias.n443 commonsourceibias.t82 168.701
R12977 commonsourceibias.n445 commonsourceibias.t90 168.701
R12978 commonsourceibias.n452 commonsourceibias.t73 168.701
R12979 commonsourceibias.n458 commonsourceibias.t83 168.701
R12980 commonsourceibias.n405 commonsourceibias.t91 168.701
R12981 commonsourceibias.n27 commonsourceibias.n24 161.3
R12982 commonsourceibias.n29 commonsourceibias.n28 161.3
R12983 commonsourceibias.n31 commonsourceibias.n30 161.3
R12984 commonsourceibias.n32 commonsourceibias.n22 161.3
R12985 commonsourceibias.n34 commonsourceibias.n33 161.3
R12986 commonsourceibias.n36 commonsourceibias.n35 161.3
R12987 commonsourceibias.n37 commonsourceibias.n20 161.3
R12988 commonsourceibias.n39 commonsourceibias.n38 161.3
R12989 commonsourceibias.n41 commonsourceibias.n40 161.3
R12990 commonsourceibias.n42 commonsourceibias.n18 161.3
R12991 commonsourceibias.n45 commonsourceibias.n44 161.3
R12992 commonsourceibias.n46 commonsourceibias.n17 161.3
R12993 commonsourceibias.n48 commonsourceibias.n47 161.3
R12994 commonsourceibias.n50 commonsourceibias.n15 161.3
R12995 commonsourceibias.n52 commonsourceibias.n51 161.3
R12996 commonsourceibias.n53 commonsourceibias.n14 161.3
R12997 commonsourceibias.n55 commonsourceibias.n54 161.3
R12998 commonsourceibias.n56 commonsourceibias.n13 161.3
R12999 commonsourceibias.n59 commonsourceibias.n58 161.3
R13000 commonsourceibias.n60 commonsourceibias.n12 161.3
R13001 commonsourceibias.n62 commonsourceibias.n61 161.3
R13002 commonsourceibias.n64 commonsourceibias.n11 161.3
R13003 commonsourceibias.n66 commonsourceibias.n65 161.3
R13004 commonsourceibias.n68 commonsourceibias.n67 161.3
R13005 commonsourceibias.n69 commonsourceibias.n9 161.3
R13006 commonsourceibias.n93 commonsourceibias.n90 161.3
R13007 commonsourceibias.n95 commonsourceibias.n94 161.3
R13008 commonsourceibias.n97 commonsourceibias.n96 161.3
R13009 commonsourceibias.n98 commonsourceibias.n88 161.3
R13010 commonsourceibias.n100 commonsourceibias.n99 161.3
R13011 commonsourceibias.n102 commonsourceibias.n101 161.3
R13012 commonsourceibias.n103 commonsourceibias.n86 161.3
R13013 commonsourceibias.n105 commonsourceibias.n104 161.3
R13014 commonsourceibias.n107 commonsourceibias.n106 161.3
R13015 commonsourceibias.n108 commonsourceibias.n84 161.3
R13016 commonsourceibias.n111 commonsourceibias.n110 161.3
R13017 commonsourceibias.n112 commonsourceibias.n8 161.3
R13018 commonsourceibias.n114 commonsourceibias.n113 161.3
R13019 commonsourceibias.n116 commonsourceibias.n6 161.3
R13020 commonsourceibias.n118 commonsourceibias.n117 161.3
R13021 commonsourceibias.n119 commonsourceibias.n5 161.3
R13022 commonsourceibias.n121 commonsourceibias.n120 161.3
R13023 commonsourceibias.n122 commonsourceibias.n4 161.3
R13024 commonsourceibias.n125 commonsourceibias.n124 161.3
R13025 commonsourceibias.n126 commonsourceibias.n3 161.3
R13026 commonsourceibias.n128 commonsourceibias.n127 161.3
R13027 commonsourceibias.n130 commonsourceibias.n2 161.3
R13028 commonsourceibias.n132 commonsourceibias.n131 161.3
R13029 commonsourceibias.n134 commonsourceibias.n133 161.3
R13030 commonsourceibias.n135 commonsourceibias.n0 161.3
R13031 commonsourceibias.n262 commonsourceibias.n202 161.3
R13032 commonsourceibias.n261 commonsourceibias.n260 161.3
R13033 commonsourceibias.n259 commonsourceibias.n258 161.3
R13034 commonsourceibias.n257 commonsourceibias.n204 161.3
R13035 commonsourceibias.n255 commonsourceibias.n254 161.3
R13036 commonsourceibias.n253 commonsourceibias.n205 161.3
R13037 commonsourceibias.n252 commonsourceibias.n251 161.3
R13038 commonsourceibias.n249 commonsourceibias.n206 161.3
R13039 commonsourceibias.n248 commonsourceibias.n247 161.3
R13040 commonsourceibias.n246 commonsourceibias.n207 161.3
R13041 commonsourceibias.n245 commonsourceibias.n244 161.3
R13042 commonsourceibias.n243 commonsourceibias.n208 161.3
R13043 commonsourceibias.n241 commonsourceibias.n240 161.3
R13044 commonsourceibias.n239 commonsourceibias.n210 161.3
R13045 commonsourceibias.n238 commonsourceibias.n237 161.3
R13046 commonsourceibias.n235 commonsourceibias.n211 161.3
R13047 commonsourceibias.n234 commonsourceibias.n233 161.3
R13048 commonsourceibias.n232 commonsourceibias.n231 161.3
R13049 commonsourceibias.n230 commonsourceibias.n213 161.3
R13050 commonsourceibias.n229 commonsourceibias.n228 161.3
R13051 commonsourceibias.n227 commonsourceibias.n226 161.3
R13052 commonsourceibias.n225 commonsourceibias.n215 161.3
R13053 commonsourceibias.n224 commonsourceibias.n223 161.3
R13054 commonsourceibias.n222 commonsourceibias.n221 161.3
R13055 commonsourceibias.n220 commonsourceibias.n217 161.3
R13056 commonsourceibias.n156 commonsourceibias.n153 161.3
R13057 commonsourceibias.n158 commonsourceibias.n157 161.3
R13058 commonsourceibias.n160 commonsourceibias.n159 161.3
R13059 commonsourceibias.n161 commonsourceibias.n151 161.3
R13060 commonsourceibias.n163 commonsourceibias.n162 161.3
R13061 commonsourceibias.n165 commonsourceibias.n164 161.3
R13062 commonsourceibias.n166 commonsourceibias.n149 161.3
R13063 commonsourceibias.n168 commonsourceibias.n167 161.3
R13064 commonsourceibias.n170 commonsourceibias.n169 161.3
R13065 commonsourceibias.n171 commonsourceibias.n147 161.3
R13066 commonsourceibias.n174 commonsourceibias.n173 161.3
R13067 commonsourceibias.n175 commonsourceibias.n146 161.3
R13068 commonsourceibias.n177 commonsourceibias.n176 161.3
R13069 commonsourceibias.n179 commonsourceibias.n144 161.3
R13070 commonsourceibias.n181 commonsourceibias.n180 161.3
R13071 commonsourceibias.n182 commonsourceibias.n143 161.3
R13072 commonsourceibias.n184 commonsourceibias.n183 161.3
R13073 commonsourceibias.n185 commonsourceibias.n142 161.3
R13074 commonsourceibias.n188 commonsourceibias.n187 161.3
R13075 commonsourceibias.n189 commonsourceibias.n141 161.3
R13076 commonsourceibias.n191 commonsourceibias.n190 161.3
R13077 commonsourceibias.n193 commonsourceibias.n140 161.3
R13078 commonsourceibias.n195 commonsourceibias.n194 161.3
R13079 commonsourceibias.n197 commonsourceibias.n196 161.3
R13080 commonsourceibias.n198 commonsourceibias.n138 161.3
R13081 commonsourceibias.n367 commonsourceibias.n307 161.3
R13082 commonsourceibias.n366 commonsourceibias.n365 161.3
R13083 commonsourceibias.n364 commonsourceibias.n363 161.3
R13084 commonsourceibias.n362 commonsourceibias.n309 161.3
R13085 commonsourceibias.n360 commonsourceibias.n359 161.3
R13086 commonsourceibias.n358 commonsourceibias.n310 161.3
R13087 commonsourceibias.n357 commonsourceibias.n356 161.3
R13088 commonsourceibias.n354 commonsourceibias.n311 161.3
R13089 commonsourceibias.n353 commonsourceibias.n352 161.3
R13090 commonsourceibias.n351 commonsourceibias.n312 161.3
R13091 commonsourceibias.n350 commonsourceibias.n349 161.3
R13092 commonsourceibias.n347 commonsourceibias.n313 161.3
R13093 commonsourceibias.n345 commonsourceibias.n344 161.3
R13094 commonsourceibias.n343 commonsourceibias.n314 161.3
R13095 commonsourceibias.n342 commonsourceibias.n341 161.3
R13096 commonsourceibias.n339 commonsourceibias.n315 161.3
R13097 commonsourceibias.n338 commonsourceibias.n337 161.3
R13098 commonsourceibias.n336 commonsourceibias.n335 161.3
R13099 commonsourceibias.n334 commonsourceibias.n317 161.3
R13100 commonsourceibias.n333 commonsourceibias.n332 161.3
R13101 commonsourceibias.n331 commonsourceibias.n330 161.3
R13102 commonsourceibias.n329 commonsourceibias.n319 161.3
R13103 commonsourceibias.n328 commonsourceibias.n327 161.3
R13104 commonsourceibias.n326 commonsourceibias.n325 161.3
R13105 commonsourceibias.n324 commonsourceibias.n321 161.3
R13106 commonsourceibias.n301 commonsourceibias.n300 161.3
R13107 commonsourceibias.n298 commonsourceibias.n274 161.3
R13108 commonsourceibias.n297 commonsourceibias.n296 161.3
R13109 commonsourceibias.n295 commonsourceibias.n294 161.3
R13110 commonsourceibias.n293 commonsourceibias.n276 161.3
R13111 commonsourceibias.n292 commonsourceibias.n291 161.3
R13112 commonsourceibias.n290 commonsourceibias.n289 161.3
R13113 commonsourceibias.n288 commonsourceibias.n278 161.3
R13114 commonsourceibias.n287 commonsourceibias.n286 161.3
R13115 commonsourceibias.n285 commonsourceibias.n284 161.3
R13116 commonsourceibias.n283 commonsourceibias.n280 161.3
R13117 commonsourceibias.n377 commonsourceibias.n273 161.3
R13118 commonsourceibias.n401 commonsourceibias.n266 161.3
R13119 commonsourceibias.n400 commonsourceibias.n399 161.3
R13120 commonsourceibias.n398 commonsourceibias.n397 161.3
R13121 commonsourceibias.n396 commonsourceibias.n268 161.3
R13122 commonsourceibias.n394 commonsourceibias.n393 161.3
R13123 commonsourceibias.n392 commonsourceibias.n269 161.3
R13124 commonsourceibias.n391 commonsourceibias.n390 161.3
R13125 commonsourceibias.n388 commonsourceibias.n270 161.3
R13126 commonsourceibias.n387 commonsourceibias.n386 161.3
R13127 commonsourceibias.n385 commonsourceibias.n271 161.3
R13128 commonsourceibias.n384 commonsourceibias.n383 161.3
R13129 commonsourceibias.n381 commonsourceibias.n272 161.3
R13130 commonsourceibias.n379 commonsourceibias.n378 161.3
R13131 commonsourceibias.n528 commonsourceibias.n468 161.3
R13132 commonsourceibias.n527 commonsourceibias.n526 161.3
R13133 commonsourceibias.n525 commonsourceibias.n524 161.3
R13134 commonsourceibias.n523 commonsourceibias.n470 161.3
R13135 commonsourceibias.n521 commonsourceibias.n520 161.3
R13136 commonsourceibias.n519 commonsourceibias.n471 161.3
R13137 commonsourceibias.n518 commonsourceibias.n517 161.3
R13138 commonsourceibias.n515 commonsourceibias.n472 161.3
R13139 commonsourceibias.n514 commonsourceibias.n513 161.3
R13140 commonsourceibias.n512 commonsourceibias.n473 161.3
R13141 commonsourceibias.n511 commonsourceibias.n510 161.3
R13142 commonsourceibias.n508 commonsourceibias.n474 161.3
R13143 commonsourceibias.n506 commonsourceibias.n505 161.3
R13144 commonsourceibias.n504 commonsourceibias.n475 161.3
R13145 commonsourceibias.n503 commonsourceibias.n502 161.3
R13146 commonsourceibias.n500 commonsourceibias.n476 161.3
R13147 commonsourceibias.n499 commonsourceibias.n498 161.3
R13148 commonsourceibias.n497 commonsourceibias.n496 161.3
R13149 commonsourceibias.n495 commonsourceibias.n478 161.3
R13150 commonsourceibias.n494 commonsourceibias.n493 161.3
R13151 commonsourceibias.n492 commonsourceibias.n491 161.3
R13152 commonsourceibias.n490 commonsourceibias.n480 161.3
R13153 commonsourceibias.n489 commonsourceibias.n488 161.3
R13154 commonsourceibias.n487 commonsourceibias.n486 161.3
R13155 commonsourceibias.n485 commonsourceibias.n482 161.3
R13156 commonsourceibias.n464 commonsourceibias.n404 161.3
R13157 commonsourceibias.n463 commonsourceibias.n462 161.3
R13158 commonsourceibias.n461 commonsourceibias.n460 161.3
R13159 commonsourceibias.n459 commonsourceibias.n406 161.3
R13160 commonsourceibias.n457 commonsourceibias.n456 161.3
R13161 commonsourceibias.n455 commonsourceibias.n407 161.3
R13162 commonsourceibias.n454 commonsourceibias.n453 161.3
R13163 commonsourceibias.n451 commonsourceibias.n408 161.3
R13164 commonsourceibias.n450 commonsourceibias.n449 161.3
R13165 commonsourceibias.n448 commonsourceibias.n409 161.3
R13166 commonsourceibias.n447 commonsourceibias.n446 161.3
R13167 commonsourceibias.n444 commonsourceibias.n410 161.3
R13168 commonsourceibias.n442 commonsourceibias.n441 161.3
R13169 commonsourceibias.n440 commonsourceibias.n411 161.3
R13170 commonsourceibias.n439 commonsourceibias.n438 161.3
R13171 commonsourceibias.n436 commonsourceibias.n412 161.3
R13172 commonsourceibias.n435 commonsourceibias.n434 161.3
R13173 commonsourceibias.n433 commonsourceibias.n432 161.3
R13174 commonsourceibias.n431 commonsourceibias.n414 161.3
R13175 commonsourceibias.n430 commonsourceibias.n429 161.3
R13176 commonsourceibias.n428 commonsourceibias.n427 161.3
R13177 commonsourceibias.n426 commonsourceibias.n416 161.3
R13178 commonsourceibias.n425 commonsourceibias.n424 161.3
R13179 commonsourceibias.n423 commonsourceibias.n422 161.3
R13180 commonsourceibias.n421 commonsourceibias.n418 161.3
R13181 commonsourceibias.n80 commonsourceibias.n78 81.5057
R13182 commonsourceibias.n304 commonsourceibias.n302 81.5057
R13183 commonsourceibias.n80 commonsourceibias.n79 80.9324
R13184 commonsourceibias.n82 commonsourceibias.n81 80.9324
R13185 commonsourceibias.n77 commonsourceibias.n76 80.9324
R13186 commonsourceibias.n75 commonsourceibias.n74 80.9324
R13187 commonsourceibias.n73 commonsourceibias.n72 80.9324
R13188 commonsourceibias.n371 commonsourceibias.n370 80.9324
R13189 commonsourceibias.n373 commonsourceibias.n372 80.9324
R13190 commonsourceibias.n375 commonsourceibias.n374 80.9324
R13191 commonsourceibias.n306 commonsourceibias.n305 80.9324
R13192 commonsourceibias.n304 commonsourceibias.n303 80.9324
R13193 commonsourceibias.n71 commonsourceibias.n70 80.6037
R13194 commonsourceibias.n137 commonsourceibias.n136 80.6037
R13195 commonsourceibias.n264 commonsourceibias.n263 80.6037
R13196 commonsourceibias.n200 commonsourceibias.n199 80.6037
R13197 commonsourceibias.n369 commonsourceibias.n368 80.6037
R13198 commonsourceibias.n403 commonsourceibias.n402 80.6037
R13199 commonsourceibias.n530 commonsourceibias.n529 80.6037
R13200 commonsourceibias.n466 commonsourceibias.n465 80.6037
R13201 commonsourceibias.n65 commonsourceibias.n64 56.5617
R13202 commonsourceibias.n51 commonsourceibias.n50 56.5617
R13203 commonsourceibias.n42 commonsourceibias.n41 56.5617
R13204 commonsourceibias.n28 commonsourceibias.n27 56.5617
R13205 commonsourceibias.n131 commonsourceibias.n130 56.5617
R13206 commonsourceibias.n117 commonsourceibias.n116 56.5617
R13207 commonsourceibias.n108 commonsourceibias.n107 56.5617
R13208 commonsourceibias.n94 commonsourceibias.n93 56.5617
R13209 commonsourceibias.n221 commonsourceibias.n220 56.5617
R13210 commonsourceibias.n235 commonsourceibias.n234 56.5617
R13211 commonsourceibias.n244 commonsourceibias.n243 56.5617
R13212 commonsourceibias.n258 commonsourceibias.n257 56.5617
R13213 commonsourceibias.n194 commonsourceibias.n193 56.5617
R13214 commonsourceibias.n180 commonsourceibias.n179 56.5617
R13215 commonsourceibias.n171 commonsourceibias.n170 56.5617
R13216 commonsourceibias.n157 commonsourceibias.n156 56.5617
R13217 commonsourceibias.n325 commonsourceibias.n324 56.5617
R13218 commonsourceibias.n339 commonsourceibias.n338 56.5617
R13219 commonsourceibias.n349 commonsourceibias.n347 56.5617
R13220 commonsourceibias.n363 commonsourceibias.n362 56.5617
R13221 commonsourceibias.n397 commonsourceibias.n396 56.5617
R13222 commonsourceibias.n383 commonsourceibias.n381 56.5617
R13223 commonsourceibias.n284 commonsourceibias.n283 56.5617
R13224 commonsourceibias.n298 commonsourceibias.n297 56.5617
R13225 commonsourceibias.n486 commonsourceibias.n485 56.5617
R13226 commonsourceibias.n500 commonsourceibias.n499 56.5617
R13227 commonsourceibias.n510 commonsourceibias.n508 56.5617
R13228 commonsourceibias.n524 commonsourceibias.n523 56.5617
R13229 commonsourceibias.n422 commonsourceibias.n421 56.5617
R13230 commonsourceibias.n436 commonsourceibias.n435 56.5617
R13231 commonsourceibias.n446 commonsourceibias.n444 56.5617
R13232 commonsourceibias.n460 commonsourceibias.n459 56.5617
R13233 commonsourceibias.n56 commonsourceibias.n55 56.0773
R13234 commonsourceibias.n37 commonsourceibias.n36 56.0773
R13235 commonsourceibias.n122 commonsourceibias.n121 56.0773
R13236 commonsourceibias.n103 commonsourceibias.n102 56.0773
R13237 commonsourceibias.n230 commonsourceibias.n229 56.0773
R13238 commonsourceibias.n249 commonsourceibias.n248 56.0773
R13239 commonsourceibias.n185 commonsourceibias.n184 56.0773
R13240 commonsourceibias.n166 commonsourceibias.n165 56.0773
R13241 commonsourceibias.n334 commonsourceibias.n333 56.0773
R13242 commonsourceibias.n354 commonsourceibias.n353 56.0773
R13243 commonsourceibias.n388 commonsourceibias.n387 56.0773
R13244 commonsourceibias.n293 commonsourceibias.n292 56.0773
R13245 commonsourceibias.n495 commonsourceibias.n494 56.0773
R13246 commonsourceibias.n515 commonsourceibias.n514 56.0773
R13247 commonsourceibias.n431 commonsourceibias.n430 56.0773
R13248 commonsourceibias.n451 commonsourceibias.n450 56.0773
R13249 commonsourceibias.n70 commonsourceibias.n69 46.0096
R13250 commonsourceibias.n136 commonsourceibias.n135 46.0096
R13251 commonsourceibias.n263 commonsourceibias.n262 46.0096
R13252 commonsourceibias.n199 commonsourceibias.n198 46.0096
R13253 commonsourceibias.n368 commonsourceibias.n367 46.0096
R13254 commonsourceibias.n402 commonsourceibias.n401 46.0096
R13255 commonsourceibias.n529 commonsourceibias.n528 46.0096
R13256 commonsourceibias.n465 commonsourceibias.n464 46.0096
R13257 commonsourceibias.n58 commonsourceibias.n12 41.5458
R13258 commonsourceibias.n33 commonsourceibias.n32 41.5458
R13259 commonsourceibias.n124 commonsourceibias.n3 41.5458
R13260 commonsourceibias.n99 commonsourceibias.n98 41.5458
R13261 commonsourceibias.n226 commonsourceibias.n225 41.5458
R13262 commonsourceibias.n251 commonsourceibias.n205 41.5458
R13263 commonsourceibias.n187 commonsourceibias.n141 41.5458
R13264 commonsourceibias.n162 commonsourceibias.n161 41.5458
R13265 commonsourceibias.n330 commonsourceibias.n329 41.5458
R13266 commonsourceibias.n356 commonsourceibias.n310 41.5458
R13267 commonsourceibias.n390 commonsourceibias.n269 41.5458
R13268 commonsourceibias.n289 commonsourceibias.n288 41.5458
R13269 commonsourceibias.n491 commonsourceibias.n490 41.5458
R13270 commonsourceibias.n517 commonsourceibias.n471 41.5458
R13271 commonsourceibias.n427 commonsourceibias.n426 41.5458
R13272 commonsourceibias.n453 commonsourceibias.n407 41.5458
R13273 commonsourceibias.n48 commonsourceibias.n17 40.577
R13274 commonsourceibias.n44 commonsourceibias.n17 40.577
R13275 commonsourceibias.n114 commonsourceibias.n8 40.577
R13276 commonsourceibias.n110 commonsourceibias.n8 40.577
R13277 commonsourceibias.n237 commonsourceibias.n210 40.577
R13278 commonsourceibias.n241 commonsourceibias.n210 40.577
R13279 commonsourceibias.n177 commonsourceibias.n146 40.577
R13280 commonsourceibias.n173 commonsourceibias.n146 40.577
R13281 commonsourceibias.n341 commonsourceibias.n314 40.577
R13282 commonsourceibias.n345 commonsourceibias.n314 40.577
R13283 commonsourceibias.n379 commonsourceibias.n273 40.577
R13284 commonsourceibias.n300 commonsourceibias.n273 40.577
R13285 commonsourceibias.n502 commonsourceibias.n475 40.577
R13286 commonsourceibias.n506 commonsourceibias.n475 40.577
R13287 commonsourceibias.n438 commonsourceibias.n411 40.577
R13288 commonsourceibias.n442 commonsourceibias.n411 40.577
R13289 commonsourceibias.n62 commonsourceibias.n12 39.6083
R13290 commonsourceibias.n32 commonsourceibias.n31 39.6083
R13291 commonsourceibias.n128 commonsourceibias.n3 39.6083
R13292 commonsourceibias.n98 commonsourceibias.n97 39.6083
R13293 commonsourceibias.n225 commonsourceibias.n224 39.6083
R13294 commonsourceibias.n255 commonsourceibias.n205 39.6083
R13295 commonsourceibias.n191 commonsourceibias.n141 39.6083
R13296 commonsourceibias.n161 commonsourceibias.n160 39.6083
R13297 commonsourceibias.n329 commonsourceibias.n328 39.6083
R13298 commonsourceibias.n360 commonsourceibias.n310 39.6083
R13299 commonsourceibias.n394 commonsourceibias.n269 39.6083
R13300 commonsourceibias.n288 commonsourceibias.n287 39.6083
R13301 commonsourceibias.n490 commonsourceibias.n489 39.6083
R13302 commonsourceibias.n521 commonsourceibias.n471 39.6083
R13303 commonsourceibias.n426 commonsourceibias.n425 39.6083
R13304 commonsourceibias.n457 commonsourceibias.n407 39.6083
R13305 commonsourceibias.n26 commonsourceibias.n25 33.0515
R13306 commonsourceibias.n92 commonsourceibias.n91 33.0515
R13307 commonsourceibias.n155 commonsourceibias.n154 33.0515
R13308 commonsourceibias.n219 commonsourceibias.n218 33.0515
R13309 commonsourceibias.n323 commonsourceibias.n322 33.0515
R13310 commonsourceibias.n282 commonsourceibias.n281 33.0515
R13311 commonsourceibias.n484 commonsourceibias.n483 33.0515
R13312 commonsourceibias.n420 commonsourceibias.n419 33.0515
R13313 commonsourceibias.n25 commonsourceibias.n24 28.5514
R13314 commonsourceibias.n91 commonsourceibias.n90 28.5514
R13315 commonsourceibias.n218 commonsourceibias.n217 28.5514
R13316 commonsourceibias.n154 commonsourceibias.n153 28.5514
R13317 commonsourceibias.n322 commonsourceibias.n321 28.5514
R13318 commonsourceibias.n281 commonsourceibias.n280 28.5514
R13319 commonsourceibias.n483 commonsourceibias.n482 28.5514
R13320 commonsourceibias.n419 commonsourceibias.n418 28.5514
R13321 commonsourceibias.n69 commonsourceibias.n68 26.0455
R13322 commonsourceibias.n135 commonsourceibias.n134 26.0455
R13323 commonsourceibias.n262 commonsourceibias.n261 26.0455
R13324 commonsourceibias.n198 commonsourceibias.n197 26.0455
R13325 commonsourceibias.n367 commonsourceibias.n366 26.0455
R13326 commonsourceibias.n401 commonsourceibias.n400 26.0455
R13327 commonsourceibias.n528 commonsourceibias.n527 26.0455
R13328 commonsourceibias.n464 commonsourceibias.n463 26.0455
R13329 commonsourceibias.n55 commonsourceibias.n14 25.0767
R13330 commonsourceibias.n38 commonsourceibias.n37 25.0767
R13331 commonsourceibias.n121 commonsourceibias.n5 25.0767
R13332 commonsourceibias.n104 commonsourceibias.n103 25.0767
R13333 commonsourceibias.n231 commonsourceibias.n230 25.0767
R13334 commonsourceibias.n248 commonsourceibias.n207 25.0767
R13335 commonsourceibias.n184 commonsourceibias.n143 25.0767
R13336 commonsourceibias.n167 commonsourceibias.n166 25.0767
R13337 commonsourceibias.n335 commonsourceibias.n334 25.0767
R13338 commonsourceibias.n353 commonsourceibias.n312 25.0767
R13339 commonsourceibias.n387 commonsourceibias.n271 25.0767
R13340 commonsourceibias.n294 commonsourceibias.n293 25.0767
R13341 commonsourceibias.n496 commonsourceibias.n495 25.0767
R13342 commonsourceibias.n514 commonsourceibias.n473 25.0767
R13343 commonsourceibias.n432 commonsourceibias.n431 25.0767
R13344 commonsourceibias.n450 commonsourceibias.n409 25.0767
R13345 commonsourceibias.n51 commonsourceibias.n16 24.3464
R13346 commonsourceibias.n41 commonsourceibias.n19 24.3464
R13347 commonsourceibias.n117 commonsourceibias.n7 24.3464
R13348 commonsourceibias.n107 commonsourceibias.n85 24.3464
R13349 commonsourceibias.n234 commonsourceibias.n212 24.3464
R13350 commonsourceibias.n244 commonsourceibias.n209 24.3464
R13351 commonsourceibias.n180 commonsourceibias.n145 24.3464
R13352 commonsourceibias.n170 commonsourceibias.n148 24.3464
R13353 commonsourceibias.n338 commonsourceibias.n316 24.3464
R13354 commonsourceibias.n349 commonsourceibias.n348 24.3464
R13355 commonsourceibias.n383 commonsourceibias.n382 24.3464
R13356 commonsourceibias.n297 commonsourceibias.n275 24.3464
R13357 commonsourceibias.n499 commonsourceibias.n477 24.3464
R13358 commonsourceibias.n510 commonsourceibias.n509 24.3464
R13359 commonsourceibias.n435 commonsourceibias.n413 24.3464
R13360 commonsourceibias.n446 commonsourceibias.n445 24.3464
R13361 commonsourceibias.n65 commonsourceibias.n10 23.8546
R13362 commonsourceibias.n27 commonsourceibias.n26 23.8546
R13363 commonsourceibias.n131 commonsourceibias.n1 23.8546
R13364 commonsourceibias.n93 commonsourceibias.n92 23.8546
R13365 commonsourceibias.n220 commonsourceibias.n219 23.8546
R13366 commonsourceibias.n258 commonsourceibias.n203 23.8546
R13367 commonsourceibias.n194 commonsourceibias.n139 23.8546
R13368 commonsourceibias.n156 commonsourceibias.n155 23.8546
R13369 commonsourceibias.n324 commonsourceibias.n323 23.8546
R13370 commonsourceibias.n363 commonsourceibias.n308 23.8546
R13371 commonsourceibias.n397 commonsourceibias.n267 23.8546
R13372 commonsourceibias.n283 commonsourceibias.n282 23.8546
R13373 commonsourceibias.n485 commonsourceibias.n484 23.8546
R13374 commonsourceibias.n524 commonsourceibias.n469 23.8546
R13375 commonsourceibias.n421 commonsourceibias.n420 23.8546
R13376 commonsourceibias.n460 commonsourceibias.n405 23.8546
R13377 commonsourceibias.n64 commonsourceibias.n63 16.9689
R13378 commonsourceibias.n28 commonsourceibias.n23 16.9689
R13379 commonsourceibias.n130 commonsourceibias.n129 16.9689
R13380 commonsourceibias.n94 commonsourceibias.n89 16.9689
R13381 commonsourceibias.n221 commonsourceibias.n216 16.9689
R13382 commonsourceibias.n257 commonsourceibias.n256 16.9689
R13383 commonsourceibias.n193 commonsourceibias.n192 16.9689
R13384 commonsourceibias.n157 commonsourceibias.n152 16.9689
R13385 commonsourceibias.n325 commonsourceibias.n320 16.9689
R13386 commonsourceibias.n362 commonsourceibias.n361 16.9689
R13387 commonsourceibias.n396 commonsourceibias.n395 16.9689
R13388 commonsourceibias.n284 commonsourceibias.n279 16.9689
R13389 commonsourceibias.n486 commonsourceibias.n481 16.9689
R13390 commonsourceibias.n523 commonsourceibias.n522 16.9689
R13391 commonsourceibias.n422 commonsourceibias.n417 16.9689
R13392 commonsourceibias.n459 commonsourceibias.n458 16.9689
R13393 commonsourceibias.n50 commonsourceibias.n49 16.477
R13394 commonsourceibias.n43 commonsourceibias.n42 16.477
R13395 commonsourceibias.n116 commonsourceibias.n115 16.477
R13396 commonsourceibias.n109 commonsourceibias.n108 16.477
R13397 commonsourceibias.n236 commonsourceibias.n235 16.477
R13398 commonsourceibias.n243 commonsourceibias.n242 16.477
R13399 commonsourceibias.n179 commonsourceibias.n178 16.477
R13400 commonsourceibias.n172 commonsourceibias.n171 16.477
R13401 commonsourceibias.n340 commonsourceibias.n339 16.477
R13402 commonsourceibias.n347 commonsourceibias.n346 16.477
R13403 commonsourceibias.n381 commonsourceibias.n380 16.477
R13404 commonsourceibias.n299 commonsourceibias.n298 16.477
R13405 commonsourceibias.n501 commonsourceibias.n500 16.477
R13406 commonsourceibias.n508 commonsourceibias.n507 16.477
R13407 commonsourceibias.n437 commonsourceibias.n436 16.477
R13408 commonsourceibias.n444 commonsourceibias.n443 16.477
R13409 commonsourceibias.n57 commonsourceibias.n56 15.9852
R13410 commonsourceibias.n36 commonsourceibias.n21 15.9852
R13411 commonsourceibias.n123 commonsourceibias.n122 15.9852
R13412 commonsourceibias.n102 commonsourceibias.n87 15.9852
R13413 commonsourceibias.n229 commonsourceibias.n214 15.9852
R13414 commonsourceibias.n250 commonsourceibias.n249 15.9852
R13415 commonsourceibias.n186 commonsourceibias.n185 15.9852
R13416 commonsourceibias.n165 commonsourceibias.n150 15.9852
R13417 commonsourceibias.n333 commonsourceibias.n318 15.9852
R13418 commonsourceibias.n355 commonsourceibias.n354 15.9852
R13419 commonsourceibias.n389 commonsourceibias.n388 15.9852
R13420 commonsourceibias.n292 commonsourceibias.n277 15.9852
R13421 commonsourceibias.n494 commonsourceibias.n479 15.9852
R13422 commonsourceibias.n516 commonsourceibias.n515 15.9852
R13423 commonsourceibias.n430 commonsourceibias.n415 15.9852
R13424 commonsourceibias.n452 commonsourceibias.n451 15.9852
R13425 commonsourceibias.n73 commonsourceibias.n71 13.2057
R13426 commonsourceibias.n371 commonsourceibias.n369 13.2057
R13427 commonsourceibias.n532 commonsourceibias.n265 10.4122
R13428 commonsourceibias.n112 commonsourceibias.n83 9.50363
R13429 commonsourceibias.n377 commonsourceibias.n376 9.50363
R13430 commonsourceibias.n201 commonsourceibias.n137 8.7339
R13431 commonsourceibias.n467 commonsourceibias.n403 8.7339
R13432 commonsourceibias.n58 commonsourceibias.n57 8.60764
R13433 commonsourceibias.n33 commonsourceibias.n21 8.60764
R13434 commonsourceibias.n124 commonsourceibias.n123 8.60764
R13435 commonsourceibias.n99 commonsourceibias.n87 8.60764
R13436 commonsourceibias.n226 commonsourceibias.n214 8.60764
R13437 commonsourceibias.n251 commonsourceibias.n250 8.60764
R13438 commonsourceibias.n187 commonsourceibias.n186 8.60764
R13439 commonsourceibias.n162 commonsourceibias.n150 8.60764
R13440 commonsourceibias.n330 commonsourceibias.n318 8.60764
R13441 commonsourceibias.n356 commonsourceibias.n355 8.60764
R13442 commonsourceibias.n390 commonsourceibias.n389 8.60764
R13443 commonsourceibias.n289 commonsourceibias.n277 8.60764
R13444 commonsourceibias.n491 commonsourceibias.n479 8.60764
R13445 commonsourceibias.n517 commonsourceibias.n516 8.60764
R13446 commonsourceibias.n427 commonsourceibias.n415 8.60764
R13447 commonsourceibias.n453 commonsourceibias.n452 8.60764
R13448 commonsourceibias.n532 commonsourceibias.n531 8.46921
R13449 commonsourceibias.n49 commonsourceibias.n48 8.11581
R13450 commonsourceibias.n44 commonsourceibias.n43 8.11581
R13451 commonsourceibias.n115 commonsourceibias.n114 8.11581
R13452 commonsourceibias.n110 commonsourceibias.n109 8.11581
R13453 commonsourceibias.n237 commonsourceibias.n236 8.11581
R13454 commonsourceibias.n242 commonsourceibias.n241 8.11581
R13455 commonsourceibias.n178 commonsourceibias.n177 8.11581
R13456 commonsourceibias.n173 commonsourceibias.n172 8.11581
R13457 commonsourceibias.n341 commonsourceibias.n340 8.11581
R13458 commonsourceibias.n346 commonsourceibias.n345 8.11581
R13459 commonsourceibias.n380 commonsourceibias.n379 8.11581
R13460 commonsourceibias.n300 commonsourceibias.n299 8.11581
R13461 commonsourceibias.n502 commonsourceibias.n501 8.11581
R13462 commonsourceibias.n507 commonsourceibias.n506 8.11581
R13463 commonsourceibias.n438 commonsourceibias.n437 8.11581
R13464 commonsourceibias.n443 commonsourceibias.n442 8.11581
R13465 commonsourceibias.n63 commonsourceibias.n62 7.62397
R13466 commonsourceibias.n31 commonsourceibias.n23 7.62397
R13467 commonsourceibias.n129 commonsourceibias.n128 7.62397
R13468 commonsourceibias.n97 commonsourceibias.n89 7.62397
R13469 commonsourceibias.n224 commonsourceibias.n216 7.62397
R13470 commonsourceibias.n256 commonsourceibias.n255 7.62397
R13471 commonsourceibias.n192 commonsourceibias.n191 7.62397
R13472 commonsourceibias.n160 commonsourceibias.n152 7.62397
R13473 commonsourceibias.n328 commonsourceibias.n320 7.62397
R13474 commonsourceibias.n361 commonsourceibias.n360 7.62397
R13475 commonsourceibias.n395 commonsourceibias.n394 7.62397
R13476 commonsourceibias.n287 commonsourceibias.n279 7.62397
R13477 commonsourceibias.n489 commonsourceibias.n481 7.62397
R13478 commonsourceibias.n522 commonsourceibias.n521 7.62397
R13479 commonsourceibias.n425 commonsourceibias.n417 7.62397
R13480 commonsourceibias.n458 commonsourceibias.n457 7.62397
R13481 commonsourceibias.n265 commonsourceibias.n264 5.00473
R13482 commonsourceibias.n201 commonsourceibias.n200 5.00473
R13483 commonsourceibias.n531 commonsourceibias.n530 5.00473
R13484 commonsourceibias.n467 commonsourceibias.n466 5.00473
R13485 commonsourceibias commonsourceibias.n532 3.87639
R13486 commonsourceibias.n265 commonsourceibias.n201 3.72967
R13487 commonsourceibias.n531 commonsourceibias.n467 3.72967
R13488 commonsourceibias.n78 commonsourceibias.t7 2.82907
R13489 commonsourceibias.n78 commonsourceibias.t35 2.82907
R13490 commonsourceibias.n79 commonsourceibias.t25 2.82907
R13491 commonsourceibias.n79 commonsourceibias.t45 2.82907
R13492 commonsourceibias.n81 commonsourceibias.t33 2.82907
R13493 commonsourceibias.n81 commonsourceibias.t41 2.82907
R13494 commonsourceibias.n76 commonsourceibias.t43 2.82907
R13495 commonsourceibias.n76 commonsourceibias.t19 2.82907
R13496 commonsourceibias.n74 commonsourceibias.t3 2.82907
R13497 commonsourceibias.n74 commonsourceibias.t23 2.82907
R13498 commonsourceibias.n72 commonsourceibias.t17 2.82907
R13499 commonsourceibias.n72 commonsourceibias.t31 2.82907
R13500 commonsourceibias.n370 commonsourceibias.t47 2.82907
R13501 commonsourceibias.n370 commonsourceibias.t27 2.82907
R13502 commonsourceibias.n372 commonsourceibias.t37 2.82907
R13503 commonsourceibias.n372 commonsourceibias.t21 2.82907
R13504 commonsourceibias.n374 commonsourceibias.t29 2.82907
R13505 commonsourceibias.n374 commonsourceibias.t11 2.82907
R13506 commonsourceibias.n305 commonsourceibias.t9 2.82907
R13507 commonsourceibias.n305 commonsourceibias.t1 2.82907
R13508 commonsourceibias.n303 commonsourceibias.t13 2.82907
R13509 commonsourceibias.n303 commonsourceibias.t39 2.82907
R13510 commonsourceibias.n302 commonsourceibias.t5 2.82907
R13511 commonsourceibias.n302 commonsourceibias.t15 2.82907
R13512 commonsourceibias.n68 commonsourceibias.n10 0.738255
R13513 commonsourceibias.n134 commonsourceibias.n1 0.738255
R13514 commonsourceibias.n261 commonsourceibias.n203 0.738255
R13515 commonsourceibias.n197 commonsourceibias.n139 0.738255
R13516 commonsourceibias.n366 commonsourceibias.n308 0.738255
R13517 commonsourceibias.n400 commonsourceibias.n267 0.738255
R13518 commonsourceibias.n527 commonsourceibias.n469 0.738255
R13519 commonsourceibias.n463 commonsourceibias.n405 0.738255
R13520 commonsourceibias.n75 commonsourceibias.n73 0.573776
R13521 commonsourceibias.n77 commonsourceibias.n75 0.573776
R13522 commonsourceibias.n82 commonsourceibias.n80 0.573776
R13523 commonsourceibias.n306 commonsourceibias.n304 0.573776
R13524 commonsourceibias.n375 commonsourceibias.n373 0.573776
R13525 commonsourceibias.n373 commonsourceibias.n371 0.573776
R13526 commonsourceibias.n83 commonsourceibias.n77 0.287138
R13527 commonsourceibias.n83 commonsourceibias.n82 0.287138
R13528 commonsourceibias.n376 commonsourceibias.n306 0.287138
R13529 commonsourceibias.n376 commonsourceibias.n375 0.287138
R13530 commonsourceibias.n71 commonsourceibias.n9 0.285035
R13531 commonsourceibias.n137 commonsourceibias.n0 0.285035
R13532 commonsourceibias.n264 commonsourceibias.n202 0.285035
R13533 commonsourceibias.n200 commonsourceibias.n138 0.285035
R13534 commonsourceibias.n369 commonsourceibias.n307 0.285035
R13535 commonsourceibias.n403 commonsourceibias.n266 0.285035
R13536 commonsourceibias.n530 commonsourceibias.n468 0.285035
R13537 commonsourceibias.n466 commonsourceibias.n404 0.285035
R13538 commonsourceibias.n16 commonsourceibias.n14 0.246418
R13539 commonsourceibias.n38 commonsourceibias.n19 0.246418
R13540 commonsourceibias.n7 commonsourceibias.n5 0.246418
R13541 commonsourceibias.n104 commonsourceibias.n85 0.246418
R13542 commonsourceibias.n231 commonsourceibias.n212 0.246418
R13543 commonsourceibias.n209 commonsourceibias.n207 0.246418
R13544 commonsourceibias.n145 commonsourceibias.n143 0.246418
R13545 commonsourceibias.n167 commonsourceibias.n148 0.246418
R13546 commonsourceibias.n335 commonsourceibias.n316 0.246418
R13547 commonsourceibias.n348 commonsourceibias.n312 0.246418
R13548 commonsourceibias.n382 commonsourceibias.n271 0.246418
R13549 commonsourceibias.n294 commonsourceibias.n275 0.246418
R13550 commonsourceibias.n496 commonsourceibias.n477 0.246418
R13551 commonsourceibias.n509 commonsourceibias.n473 0.246418
R13552 commonsourceibias.n432 commonsourceibias.n413 0.246418
R13553 commonsourceibias.n445 commonsourceibias.n409 0.246418
R13554 commonsourceibias.n67 commonsourceibias.n9 0.189894
R13555 commonsourceibias.n67 commonsourceibias.n66 0.189894
R13556 commonsourceibias.n66 commonsourceibias.n11 0.189894
R13557 commonsourceibias.n61 commonsourceibias.n11 0.189894
R13558 commonsourceibias.n61 commonsourceibias.n60 0.189894
R13559 commonsourceibias.n60 commonsourceibias.n59 0.189894
R13560 commonsourceibias.n59 commonsourceibias.n13 0.189894
R13561 commonsourceibias.n54 commonsourceibias.n13 0.189894
R13562 commonsourceibias.n54 commonsourceibias.n53 0.189894
R13563 commonsourceibias.n53 commonsourceibias.n52 0.189894
R13564 commonsourceibias.n52 commonsourceibias.n15 0.189894
R13565 commonsourceibias.n47 commonsourceibias.n15 0.189894
R13566 commonsourceibias.n47 commonsourceibias.n46 0.189894
R13567 commonsourceibias.n46 commonsourceibias.n45 0.189894
R13568 commonsourceibias.n45 commonsourceibias.n18 0.189894
R13569 commonsourceibias.n40 commonsourceibias.n18 0.189894
R13570 commonsourceibias.n40 commonsourceibias.n39 0.189894
R13571 commonsourceibias.n39 commonsourceibias.n20 0.189894
R13572 commonsourceibias.n35 commonsourceibias.n20 0.189894
R13573 commonsourceibias.n35 commonsourceibias.n34 0.189894
R13574 commonsourceibias.n34 commonsourceibias.n22 0.189894
R13575 commonsourceibias.n30 commonsourceibias.n22 0.189894
R13576 commonsourceibias.n30 commonsourceibias.n29 0.189894
R13577 commonsourceibias.n29 commonsourceibias.n24 0.189894
R13578 commonsourceibias.n111 commonsourceibias.n84 0.189894
R13579 commonsourceibias.n106 commonsourceibias.n84 0.189894
R13580 commonsourceibias.n106 commonsourceibias.n105 0.189894
R13581 commonsourceibias.n105 commonsourceibias.n86 0.189894
R13582 commonsourceibias.n101 commonsourceibias.n86 0.189894
R13583 commonsourceibias.n101 commonsourceibias.n100 0.189894
R13584 commonsourceibias.n100 commonsourceibias.n88 0.189894
R13585 commonsourceibias.n96 commonsourceibias.n88 0.189894
R13586 commonsourceibias.n96 commonsourceibias.n95 0.189894
R13587 commonsourceibias.n95 commonsourceibias.n90 0.189894
R13588 commonsourceibias.n133 commonsourceibias.n0 0.189894
R13589 commonsourceibias.n133 commonsourceibias.n132 0.189894
R13590 commonsourceibias.n132 commonsourceibias.n2 0.189894
R13591 commonsourceibias.n127 commonsourceibias.n2 0.189894
R13592 commonsourceibias.n127 commonsourceibias.n126 0.189894
R13593 commonsourceibias.n126 commonsourceibias.n125 0.189894
R13594 commonsourceibias.n125 commonsourceibias.n4 0.189894
R13595 commonsourceibias.n120 commonsourceibias.n4 0.189894
R13596 commonsourceibias.n120 commonsourceibias.n119 0.189894
R13597 commonsourceibias.n119 commonsourceibias.n118 0.189894
R13598 commonsourceibias.n118 commonsourceibias.n6 0.189894
R13599 commonsourceibias.n113 commonsourceibias.n6 0.189894
R13600 commonsourceibias.n260 commonsourceibias.n202 0.189894
R13601 commonsourceibias.n260 commonsourceibias.n259 0.189894
R13602 commonsourceibias.n259 commonsourceibias.n204 0.189894
R13603 commonsourceibias.n254 commonsourceibias.n204 0.189894
R13604 commonsourceibias.n254 commonsourceibias.n253 0.189894
R13605 commonsourceibias.n253 commonsourceibias.n252 0.189894
R13606 commonsourceibias.n252 commonsourceibias.n206 0.189894
R13607 commonsourceibias.n247 commonsourceibias.n206 0.189894
R13608 commonsourceibias.n247 commonsourceibias.n246 0.189894
R13609 commonsourceibias.n246 commonsourceibias.n245 0.189894
R13610 commonsourceibias.n245 commonsourceibias.n208 0.189894
R13611 commonsourceibias.n240 commonsourceibias.n208 0.189894
R13612 commonsourceibias.n240 commonsourceibias.n239 0.189894
R13613 commonsourceibias.n239 commonsourceibias.n238 0.189894
R13614 commonsourceibias.n238 commonsourceibias.n211 0.189894
R13615 commonsourceibias.n233 commonsourceibias.n211 0.189894
R13616 commonsourceibias.n233 commonsourceibias.n232 0.189894
R13617 commonsourceibias.n232 commonsourceibias.n213 0.189894
R13618 commonsourceibias.n228 commonsourceibias.n213 0.189894
R13619 commonsourceibias.n228 commonsourceibias.n227 0.189894
R13620 commonsourceibias.n227 commonsourceibias.n215 0.189894
R13621 commonsourceibias.n223 commonsourceibias.n215 0.189894
R13622 commonsourceibias.n223 commonsourceibias.n222 0.189894
R13623 commonsourceibias.n222 commonsourceibias.n217 0.189894
R13624 commonsourceibias.n196 commonsourceibias.n138 0.189894
R13625 commonsourceibias.n196 commonsourceibias.n195 0.189894
R13626 commonsourceibias.n195 commonsourceibias.n140 0.189894
R13627 commonsourceibias.n190 commonsourceibias.n140 0.189894
R13628 commonsourceibias.n190 commonsourceibias.n189 0.189894
R13629 commonsourceibias.n189 commonsourceibias.n188 0.189894
R13630 commonsourceibias.n188 commonsourceibias.n142 0.189894
R13631 commonsourceibias.n183 commonsourceibias.n142 0.189894
R13632 commonsourceibias.n183 commonsourceibias.n182 0.189894
R13633 commonsourceibias.n182 commonsourceibias.n181 0.189894
R13634 commonsourceibias.n181 commonsourceibias.n144 0.189894
R13635 commonsourceibias.n176 commonsourceibias.n144 0.189894
R13636 commonsourceibias.n176 commonsourceibias.n175 0.189894
R13637 commonsourceibias.n175 commonsourceibias.n174 0.189894
R13638 commonsourceibias.n174 commonsourceibias.n147 0.189894
R13639 commonsourceibias.n169 commonsourceibias.n147 0.189894
R13640 commonsourceibias.n169 commonsourceibias.n168 0.189894
R13641 commonsourceibias.n168 commonsourceibias.n149 0.189894
R13642 commonsourceibias.n164 commonsourceibias.n149 0.189894
R13643 commonsourceibias.n164 commonsourceibias.n163 0.189894
R13644 commonsourceibias.n163 commonsourceibias.n151 0.189894
R13645 commonsourceibias.n159 commonsourceibias.n151 0.189894
R13646 commonsourceibias.n159 commonsourceibias.n158 0.189894
R13647 commonsourceibias.n158 commonsourceibias.n153 0.189894
R13648 commonsourceibias.n326 commonsourceibias.n321 0.189894
R13649 commonsourceibias.n327 commonsourceibias.n326 0.189894
R13650 commonsourceibias.n327 commonsourceibias.n319 0.189894
R13651 commonsourceibias.n331 commonsourceibias.n319 0.189894
R13652 commonsourceibias.n332 commonsourceibias.n331 0.189894
R13653 commonsourceibias.n332 commonsourceibias.n317 0.189894
R13654 commonsourceibias.n336 commonsourceibias.n317 0.189894
R13655 commonsourceibias.n337 commonsourceibias.n336 0.189894
R13656 commonsourceibias.n337 commonsourceibias.n315 0.189894
R13657 commonsourceibias.n342 commonsourceibias.n315 0.189894
R13658 commonsourceibias.n343 commonsourceibias.n342 0.189894
R13659 commonsourceibias.n344 commonsourceibias.n343 0.189894
R13660 commonsourceibias.n344 commonsourceibias.n313 0.189894
R13661 commonsourceibias.n350 commonsourceibias.n313 0.189894
R13662 commonsourceibias.n351 commonsourceibias.n350 0.189894
R13663 commonsourceibias.n352 commonsourceibias.n351 0.189894
R13664 commonsourceibias.n352 commonsourceibias.n311 0.189894
R13665 commonsourceibias.n357 commonsourceibias.n311 0.189894
R13666 commonsourceibias.n358 commonsourceibias.n357 0.189894
R13667 commonsourceibias.n359 commonsourceibias.n358 0.189894
R13668 commonsourceibias.n359 commonsourceibias.n309 0.189894
R13669 commonsourceibias.n364 commonsourceibias.n309 0.189894
R13670 commonsourceibias.n365 commonsourceibias.n364 0.189894
R13671 commonsourceibias.n365 commonsourceibias.n307 0.189894
R13672 commonsourceibias.n285 commonsourceibias.n280 0.189894
R13673 commonsourceibias.n286 commonsourceibias.n285 0.189894
R13674 commonsourceibias.n286 commonsourceibias.n278 0.189894
R13675 commonsourceibias.n290 commonsourceibias.n278 0.189894
R13676 commonsourceibias.n291 commonsourceibias.n290 0.189894
R13677 commonsourceibias.n291 commonsourceibias.n276 0.189894
R13678 commonsourceibias.n295 commonsourceibias.n276 0.189894
R13679 commonsourceibias.n296 commonsourceibias.n295 0.189894
R13680 commonsourceibias.n296 commonsourceibias.n274 0.189894
R13681 commonsourceibias.n301 commonsourceibias.n274 0.189894
R13682 commonsourceibias.n378 commonsourceibias.n272 0.189894
R13683 commonsourceibias.n384 commonsourceibias.n272 0.189894
R13684 commonsourceibias.n385 commonsourceibias.n384 0.189894
R13685 commonsourceibias.n386 commonsourceibias.n385 0.189894
R13686 commonsourceibias.n386 commonsourceibias.n270 0.189894
R13687 commonsourceibias.n391 commonsourceibias.n270 0.189894
R13688 commonsourceibias.n392 commonsourceibias.n391 0.189894
R13689 commonsourceibias.n393 commonsourceibias.n392 0.189894
R13690 commonsourceibias.n393 commonsourceibias.n268 0.189894
R13691 commonsourceibias.n398 commonsourceibias.n268 0.189894
R13692 commonsourceibias.n399 commonsourceibias.n398 0.189894
R13693 commonsourceibias.n399 commonsourceibias.n266 0.189894
R13694 commonsourceibias.n487 commonsourceibias.n482 0.189894
R13695 commonsourceibias.n488 commonsourceibias.n487 0.189894
R13696 commonsourceibias.n488 commonsourceibias.n480 0.189894
R13697 commonsourceibias.n492 commonsourceibias.n480 0.189894
R13698 commonsourceibias.n493 commonsourceibias.n492 0.189894
R13699 commonsourceibias.n493 commonsourceibias.n478 0.189894
R13700 commonsourceibias.n497 commonsourceibias.n478 0.189894
R13701 commonsourceibias.n498 commonsourceibias.n497 0.189894
R13702 commonsourceibias.n498 commonsourceibias.n476 0.189894
R13703 commonsourceibias.n503 commonsourceibias.n476 0.189894
R13704 commonsourceibias.n504 commonsourceibias.n503 0.189894
R13705 commonsourceibias.n505 commonsourceibias.n504 0.189894
R13706 commonsourceibias.n505 commonsourceibias.n474 0.189894
R13707 commonsourceibias.n511 commonsourceibias.n474 0.189894
R13708 commonsourceibias.n512 commonsourceibias.n511 0.189894
R13709 commonsourceibias.n513 commonsourceibias.n512 0.189894
R13710 commonsourceibias.n513 commonsourceibias.n472 0.189894
R13711 commonsourceibias.n518 commonsourceibias.n472 0.189894
R13712 commonsourceibias.n519 commonsourceibias.n518 0.189894
R13713 commonsourceibias.n520 commonsourceibias.n519 0.189894
R13714 commonsourceibias.n520 commonsourceibias.n470 0.189894
R13715 commonsourceibias.n525 commonsourceibias.n470 0.189894
R13716 commonsourceibias.n526 commonsourceibias.n525 0.189894
R13717 commonsourceibias.n526 commonsourceibias.n468 0.189894
R13718 commonsourceibias.n423 commonsourceibias.n418 0.189894
R13719 commonsourceibias.n424 commonsourceibias.n423 0.189894
R13720 commonsourceibias.n424 commonsourceibias.n416 0.189894
R13721 commonsourceibias.n428 commonsourceibias.n416 0.189894
R13722 commonsourceibias.n429 commonsourceibias.n428 0.189894
R13723 commonsourceibias.n429 commonsourceibias.n414 0.189894
R13724 commonsourceibias.n433 commonsourceibias.n414 0.189894
R13725 commonsourceibias.n434 commonsourceibias.n433 0.189894
R13726 commonsourceibias.n434 commonsourceibias.n412 0.189894
R13727 commonsourceibias.n439 commonsourceibias.n412 0.189894
R13728 commonsourceibias.n440 commonsourceibias.n439 0.189894
R13729 commonsourceibias.n441 commonsourceibias.n440 0.189894
R13730 commonsourceibias.n441 commonsourceibias.n410 0.189894
R13731 commonsourceibias.n447 commonsourceibias.n410 0.189894
R13732 commonsourceibias.n448 commonsourceibias.n447 0.189894
R13733 commonsourceibias.n449 commonsourceibias.n448 0.189894
R13734 commonsourceibias.n449 commonsourceibias.n408 0.189894
R13735 commonsourceibias.n454 commonsourceibias.n408 0.189894
R13736 commonsourceibias.n455 commonsourceibias.n454 0.189894
R13737 commonsourceibias.n456 commonsourceibias.n455 0.189894
R13738 commonsourceibias.n456 commonsourceibias.n406 0.189894
R13739 commonsourceibias.n461 commonsourceibias.n406 0.189894
R13740 commonsourceibias.n462 commonsourceibias.n461 0.189894
R13741 commonsourceibias.n462 commonsourceibias.n404 0.189894
R13742 commonsourceibias.n112 commonsourceibias.n111 0.170955
R13743 commonsourceibias.n113 commonsourceibias.n112 0.170955
R13744 commonsourceibias.n377 commonsourceibias.n301 0.170955
R13745 commonsourceibias.n378 commonsourceibias.n377 0.170955
R13746 a_n5644_8799.n94 a_n5644_8799.t69 485.149
R13747 a_n5644_8799.n101 a_n5644_8799.t72 485.149
R13748 a_n5644_8799.n109 a_n5644_8799.t38 485.149
R13749 a_n5644_8799.n70 a_n5644_8799.t53 485.149
R13750 a_n5644_8799.n77 a_n5644_8799.t58 485.149
R13751 a_n5644_8799.n85 a_n5644_8799.t39 485.149
R13752 a_n5644_8799.n24 a_n5644_8799.t60 485.135
R13753 a_n5644_8799.n98 a_n5644_8799.t59 464.166
R13754 a_n5644_8799.n92 a_n5644_8799.t46 464.166
R13755 a_n5644_8799.n97 a_n5644_8799.t76 464.166
R13756 a_n5644_8799.n96 a_n5644_8799.t61 464.166
R13757 a_n5644_8799.n93 a_n5644_8799.t51 464.166
R13758 a_n5644_8799.n95 a_n5644_8799.t78 464.166
R13759 a_n5644_8799.n29 a_n5644_8799.t64 485.135
R13760 a_n5644_8799.n105 a_n5644_8799.t63 464.166
R13761 a_n5644_8799.n99 a_n5644_8799.t55 464.166
R13762 a_n5644_8799.n104 a_n5644_8799.t80 464.166
R13763 a_n5644_8799.n103 a_n5644_8799.t67 464.166
R13764 a_n5644_8799.n100 a_n5644_8799.t56 464.166
R13765 a_n5644_8799.n102 a_n5644_8799.t36 464.166
R13766 a_n5644_8799.n34 a_n5644_8799.t82 485.135
R13767 a_n5644_8799.n113 a_n5644_8799.t44 464.166
R13768 a_n5644_8799.n107 a_n5644_8799.t65 464.166
R13769 a_n5644_8799.n112 a_n5644_8799.t37 464.166
R13770 a_n5644_8799.n111 a_n5644_8799.t73 464.166
R13771 a_n5644_8799.n108 a_n5644_8799.t50 464.166
R13772 a_n5644_8799.n110 a_n5644_8799.t70 464.166
R13773 a_n5644_8799.n71 a_n5644_8799.t62 464.166
R13774 a_n5644_8799.n72 a_n5644_8799.t77 464.166
R13775 a_n5644_8799.n73 a_n5644_8799.t42 464.166
R13776 a_n5644_8799.n74 a_n5644_8799.t52 464.166
R13777 a_n5644_8799.n69 a_n5644_8799.t75 464.166
R13778 a_n5644_8799.n75 a_n5644_8799.t41 464.166
R13779 a_n5644_8799.n78 a_n5644_8799.t68 464.166
R13780 a_n5644_8799.n79 a_n5644_8799.t81 464.166
R13781 a_n5644_8799.n80 a_n5644_8799.t49 464.166
R13782 a_n5644_8799.n81 a_n5644_8799.t57 464.166
R13783 a_n5644_8799.n76 a_n5644_8799.t79 464.166
R13784 a_n5644_8799.n82 a_n5644_8799.t45 464.166
R13785 a_n5644_8799.n86 a_n5644_8799.t71 464.166
R13786 a_n5644_8799.n87 a_n5644_8799.t48 464.166
R13787 a_n5644_8799.n88 a_n5644_8799.t74 464.166
R13788 a_n5644_8799.n89 a_n5644_8799.t54 464.166
R13789 a_n5644_8799.n84 a_n5644_8799.t66 464.166
R13790 a_n5644_8799.n90 a_n5644_8799.t43 464.166
R13791 a_n5644_8799.n16 a_n5644_8799.n28 72.3034
R13792 a_n5644_8799.n28 a_n5644_8799.n93 16.6962
R13793 a_n5644_8799.n27 a_n5644_8799.n16 77.6622
R13794 a_n5644_8799.n96 a_n5644_8799.n27 5.97853
R13795 a_n5644_8799.n26 a_n5644_8799.n15 77.6622
R13796 a_n5644_8799.n15 a_n5644_8799.n25 72.3034
R13797 a_n5644_8799.n98 a_n5644_8799.n24 20.9683
R13798 a_n5644_8799.n17 a_n5644_8799.n24 70.1674
R13799 a_n5644_8799.n13 a_n5644_8799.n33 72.3034
R13800 a_n5644_8799.n33 a_n5644_8799.n100 16.6962
R13801 a_n5644_8799.n32 a_n5644_8799.n13 77.6622
R13802 a_n5644_8799.n103 a_n5644_8799.n32 5.97853
R13803 a_n5644_8799.n31 a_n5644_8799.n12 77.6622
R13804 a_n5644_8799.n12 a_n5644_8799.n30 72.3034
R13805 a_n5644_8799.n105 a_n5644_8799.n29 20.9683
R13806 a_n5644_8799.n14 a_n5644_8799.n29 70.1674
R13807 a_n5644_8799.n10 a_n5644_8799.n38 72.3034
R13808 a_n5644_8799.n38 a_n5644_8799.n108 16.6962
R13809 a_n5644_8799.n37 a_n5644_8799.n10 77.6622
R13810 a_n5644_8799.n111 a_n5644_8799.n37 5.97853
R13811 a_n5644_8799.n36 a_n5644_8799.n9 77.6622
R13812 a_n5644_8799.n9 a_n5644_8799.n35 72.3034
R13813 a_n5644_8799.n113 a_n5644_8799.n34 20.9683
R13814 a_n5644_8799.n11 a_n5644_8799.n34 70.1674
R13815 a_n5644_8799.n7 a_n5644_8799.n43 70.1674
R13816 a_n5644_8799.n75 a_n5644_8799.n43 20.9683
R13817 a_n5644_8799.n42 a_n5644_8799.n7 72.3034
R13818 a_n5644_8799.n42 a_n5644_8799.n69 16.6962
R13819 a_n5644_8799.n6 a_n5644_8799.n41 77.6622
R13820 a_n5644_8799.n74 a_n5644_8799.n41 5.97853
R13821 a_n5644_8799.n40 a_n5644_8799.n6 77.6622
R13822 a_n5644_8799.n39 a_n5644_8799.n72 16.6962
R13823 a_n5644_8799.n39 a_n5644_8799.n8 72.3034
R13824 a_n5644_8799.n4 a_n5644_8799.n48 70.1674
R13825 a_n5644_8799.n82 a_n5644_8799.n48 20.9683
R13826 a_n5644_8799.n47 a_n5644_8799.n4 72.3034
R13827 a_n5644_8799.n47 a_n5644_8799.n76 16.6962
R13828 a_n5644_8799.n3 a_n5644_8799.n46 77.6622
R13829 a_n5644_8799.n81 a_n5644_8799.n46 5.97853
R13830 a_n5644_8799.n45 a_n5644_8799.n3 77.6622
R13831 a_n5644_8799.n44 a_n5644_8799.n79 16.6962
R13832 a_n5644_8799.n44 a_n5644_8799.n5 72.3034
R13833 a_n5644_8799.n1 a_n5644_8799.n53 70.1674
R13834 a_n5644_8799.n90 a_n5644_8799.n53 20.9683
R13835 a_n5644_8799.n52 a_n5644_8799.n1 72.3034
R13836 a_n5644_8799.n52 a_n5644_8799.n84 16.6962
R13837 a_n5644_8799.n0 a_n5644_8799.n51 77.6622
R13838 a_n5644_8799.n89 a_n5644_8799.n51 5.97853
R13839 a_n5644_8799.n50 a_n5644_8799.n0 77.6622
R13840 a_n5644_8799.n49 a_n5644_8799.n87 16.6962
R13841 a_n5644_8799.n49 a_n5644_8799.n2 72.3034
R13842 a_n5644_8799.n21 a_n5644_8799.n54 98.9633
R13843 a_n5644_8799.n22 a_n5644_8799.n119 98.9631
R13844 a_n5644_8799.n22 a_n5644_8799.n118 98.6055
R13845 a_n5644_8799.n21 a_n5644_8799.n56 98.6055
R13846 a_n5644_8799.n21 a_n5644_8799.n55 98.6055
R13847 a_n5644_8799.n120 a_n5644_8799.n22 98.6054
R13848 a_n5644_8799.n19 a_n5644_8799.n57 81.2902
R13849 a_n5644_8799.n23 a_n5644_8799.n63 81.2902
R13850 a_n5644_8799.n18 a_n5644_8799.n60 81.2902
R13851 a_n5644_8799.n20 a_n5644_8799.n66 80.9324
R13852 a_n5644_8799.n20 a_n5644_8799.n67 80.9324
R13853 a_n5644_8799.n19 a_n5644_8799.n68 80.9324
R13854 a_n5644_8799.n19 a_n5644_8799.n59 80.9324
R13855 a_n5644_8799.n19 a_n5644_8799.n58 80.9324
R13856 a_n5644_8799.n23 a_n5644_8799.n64 80.9324
R13857 a_n5644_8799.n18 a_n5644_8799.n65 80.9324
R13858 a_n5644_8799.n18 a_n5644_8799.n62 80.9324
R13859 a_n5644_8799.n18 a_n5644_8799.n61 80.9324
R13860 a_n5644_8799.n16 a_n5644_8799.n94 70.4033
R13861 a_n5644_8799.n13 a_n5644_8799.n101 70.4033
R13862 a_n5644_8799.n10 a_n5644_8799.n109 70.4033
R13863 a_n5644_8799.n70 a_n5644_8799.n8 70.4033
R13864 a_n5644_8799.n77 a_n5644_8799.n5 70.4033
R13865 a_n5644_8799.n85 a_n5644_8799.n2 70.4033
R13866 a_n5644_8799.n97 a_n5644_8799.n96 48.2005
R13867 a_n5644_8799.n104 a_n5644_8799.n103 48.2005
R13868 a_n5644_8799.n112 a_n5644_8799.n111 48.2005
R13869 a_n5644_8799.n74 a_n5644_8799.n73 48.2005
R13870 a_n5644_8799.t40 a_n5644_8799.n43 485.135
R13871 a_n5644_8799.n81 a_n5644_8799.n80 48.2005
R13872 a_n5644_8799.t47 a_n5644_8799.n48 485.135
R13873 a_n5644_8799.n89 a_n5644_8799.n88 48.2005
R13874 a_n5644_8799.t83 a_n5644_8799.n53 485.135
R13875 a_n5644_8799.n25 a_n5644_8799.n92 16.6962
R13876 a_n5644_8799.n95 a_n5644_8799.n28 27.6507
R13877 a_n5644_8799.n30 a_n5644_8799.n99 16.6962
R13878 a_n5644_8799.n102 a_n5644_8799.n33 27.6507
R13879 a_n5644_8799.n35 a_n5644_8799.n107 16.6962
R13880 a_n5644_8799.n110 a_n5644_8799.n38 27.6507
R13881 a_n5644_8799.n75 a_n5644_8799.n42 27.6507
R13882 a_n5644_8799.n82 a_n5644_8799.n47 27.6507
R13883 a_n5644_8799.n90 a_n5644_8799.n52 27.6507
R13884 a_n5644_8799.n26 a_n5644_8799.n92 41.7634
R13885 a_n5644_8799.n31 a_n5644_8799.n99 41.7634
R13886 a_n5644_8799.n36 a_n5644_8799.n107 41.7634
R13887 a_n5644_8799.n72 a_n5644_8799.n40 41.7634
R13888 a_n5644_8799.n79 a_n5644_8799.n45 41.7634
R13889 a_n5644_8799.n87 a_n5644_8799.n50 41.7634
R13890 a_n5644_8799.n20 a_n5644_8799.n18 32.5134
R13891 a_n5644_8799.n95 a_n5644_8799.n94 20.9576
R13892 a_n5644_8799.n102 a_n5644_8799.n101 20.9576
R13893 a_n5644_8799.n110 a_n5644_8799.n109 20.9576
R13894 a_n5644_8799.n71 a_n5644_8799.n70 20.9576
R13895 a_n5644_8799.n78 a_n5644_8799.n77 20.9576
R13896 a_n5644_8799.n86 a_n5644_8799.n85 20.9576
R13897 a_n5644_8799.n26 a_n5644_8799.n97 5.97853
R13898 a_n5644_8799.n27 a_n5644_8799.n93 41.7634
R13899 a_n5644_8799.n31 a_n5644_8799.n104 5.97853
R13900 a_n5644_8799.n32 a_n5644_8799.n100 41.7634
R13901 a_n5644_8799.n36 a_n5644_8799.n112 5.97853
R13902 a_n5644_8799.n37 a_n5644_8799.n108 41.7634
R13903 a_n5644_8799.n73 a_n5644_8799.n40 5.97853
R13904 a_n5644_8799.n69 a_n5644_8799.n41 41.7634
R13905 a_n5644_8799.n80 a_n5644_8799.n45 5.97853
R13906 a_n5644_8799.n76 a_n5644_8799.n46 41.7634
R13907 a_n5644_8799.n88 a_n5644_8799.n50 5.97853
R13908 a_n5644_8799.n84 a_n5644_8799.n51 41.7634
R13909 a_n5644_8799.n22 a_n5644_8799.n117 31.0347
R13910 a_n5644_8799.n116 a_n5644_8799.n19 12.3339
R13911 a_n5644_8799.n117 a_n5644_8799.n116 11.4887
R13912 a_n5644_8799.n98 a_n5644_8799.n25 27.6507
R13913 a_n5644_8799.n105 a_n5644_8799.n30 27.6507
R13914 a_n5644_8799.n113 a_n5644_8799.n35 27.6507
R13915 a_n5644_8799.n39 a_n5644_8799.n71 27.6507
R13916 a_n5644_8799.n44 a_n5644_8799.n78 27.6507
R13917 a_n5644_8799.n49 a_n5644_8799.n86 27.6507
R13918 a_n5644_8799.n117 a_n5644_8799.n21 18.1305
R13919 a_n5644_8799.n106 a_n5644_8799.n17 9.05164
R13920 a_n5644_8799.n83 a_n5644_8799.n7 9.05164
R13921 a_n5644_8799.n115 a_n5644_8799.n91 6.86452
R13922 a_n5644_8799.n115 a_n5644_8799.n114 6.51829
R13923 a_n5644_8799.n106 a_n5644_8799.n14 4.94368
R13924 a_n5644_8799.n114 a_n5644_8799.n11 4.94368
R13925 a_n5644_8799.n83 a_n5644_8799.n4 4.94368
R13926 a_n5644_8799.n91 a_n5644_8799.n1 4.94368
R13927 a_n5644_8799.n114 a_n5644_8799.n106 4.10845
R13928 a_n5644_8799.n91 a_n5644_8799.n83 4.10845
R13929 a_n5644_8799.n119 a_n5644_8799.t30 3.61217
R13930 a_n5644_8799.n119 a_n5644_8799.t12 3.61217
R13931 a_n5644_8799.n118 a_n5644_8799.t9 3.61217
R13932 a_n5644_8799.n118 a_n5644_8799.t10 3.61217
R13933 a_n5644_8799.n56 a_n5644_8799.t19 3.61217
R13934 a_n5644_8799.n56 a_n5644_8799.t18 3.61217
R13935 a_n5644_8799.n55 a_n5644_8799.t15 3.61217
R13936 a_n5644_8799.n55 a_n5644_8799.t20 3.61217
R13937 a_n5644_8799.n54 a_n5644_8799.t13 3.61217
R13938 a_n5644_8799.n54 a_n5644_8799.t32 3.61217
R13939 a_n5644_8799.n120 a_n5644_8799.t11 3.61217
R13940 a_n5644_8799.t7 a_n5644_8799.n120 3.61217
R13941 a_n5644_8799.n116 a_n5644_8799.n115 3.4105
R13942 a_n5644_8799.n66 a_n5644_8799.t28 2.82907
R13943 a_n5644_8799.n66 a_n5644_8799.t5 2.82907
R13944 a_n5644_8799.n67 a_n5644_8799.t0 2.82907
R13945 a_n5644_8799.n67 a_n5644_8799.t35 2.82907
R13946 a_n5644_8799.n68 a_n5644_8799.t21 2.82907
R13947 a_n5644_8799.n68 a_n5644_8799.t31 2.82907
R13948 a_n5644_8799.n59 a_n5644_8799.t25 2.82907
R13949 a_n5644_8799.n59 a_n5644_8799.t24 2.82907
R13950 a_n5644_8799.n58 a_n5644_8799.t6 2.82907
R13951 a_n5644_8799.n58 a_n5644_8799.t16 2.82907
R13952 a_n5644_8799.n57 a_n5644_8799.t27 2.82907
R13953 a_n5644_8799.n57 a_n5644_8799.t26 2.82907
R13954 a_n5644_8799.n63 a_n5644_8799.t14 2.82907
R13955 a_n5644_8799.n63 a_n5644_8799.t23 2.82907
R13956 a_n5644_8799.n64 a_n5644_8799.t34 2.82907
R13957 a_n5644_8799.n64 a_n5644_8799.t29 2.82907
R13958 a_n5644_8799.n65 a_n5644_8799.t4 2.82907
R13959 a_n5644_8799.n65 a_n5644_8799.t8 2.82907
R13960 a_n5644_8799.n62 a_n5644_8799.t3 2.82907
R13961 a_n5644_8799.n62 a_n5644_8799.t1 2.82907
R13962 a_n5644_8799.n61 a_n5644_8799.t2 2.82907
R13963 a_n5644_8799.n61 a_n5644_8799.t17 2.82907
R13964 a_n5644_8799.n60 a_n5644_8799.t33 2.82907
R13965 a_n5644_8799.n60 a_n5644_8799.t22 2.82907
R13966 a_n5644_8799.n19 a_n5644_8799.n20 1.43153
R13967 a_n5644_8799.n16 a_n5644_8799.n15 1.13686
R13968 a_n5644_8799.n13 a_n5644_8799.n12 1.13686
R13969 a_n5644_8799.n10 a_n5644_8799.n9 1.13686
R13970 a_n5644_8799.n7 a_n5644_8799.n6 1.13686
R13971 a_n5644_8799.n4 a_n5644_8799.n3 1.13686
R13972 a_n5644_8799.n1 a_n5644_8799.n0 1.13686
R13973 a_n5644_8799.n18 a_n5644_8799.n23 1.07378
R13974 a_n5644_8799.n0 a_n5644_8799.n2 0.568682
R13975 a_n5644_8799.n3 a_n5644_8799.n5 0.568682
R13976 a_n5644_8799.n6 a_n5644_8799.n8 0.568682
R13977 a_n5644_8799.n9 a_n5644_8799.n11 0.568682
R13978 a_n5644_8799.n12 a_n5644_8799.n14 0.568682
R13979 a_n5644_8799.n15 a_n5644_8799.n17 0.568682
R13980 CSoutput.n19 CSoutput.t137 184.661
R13981 CSoutput.n78 CSoutput.n77 165.8
R13982 CSoutput.n76 CSoutput.n0 165.8
R13983 CSoutput.n75 CSoutput.n74 165.8
R13984 CSoutput.n73 CSoutput.n72 165.8
R13985 CSoutput.n71 CSoutput.n2 165.8
R13986 CSoutput.n69 CSoutput.n68 165.8
R13987 CSoutput.n67 CSoutput.n3 165.8
R13988 CSoutput.n66 CSoutput.n65 165.8
R13989 CSoutput.n63 CSoutput.n4 165.8
R13990 CSoutput.n61 CSoutput.n60 165.8
R13991 CSoutput.n59 CSoutput.n5 165.8
R13992 CSoutput.n58 CSoutput.n57 165.8
R13993 CSoutput.n55 CSoutput.n6 165.8
R13994 CSoutput.n54 CSoutput.n53 165.8
R13995 CSoutput.n52 CSoutput.n51 165.8
R13996 CSoutput.n50 CSoutput.n8 165.8
R13997 CSoutput.n48 CSoutput.n47 165.8
R13998 CSoutput.n46 CSoutput.n9 165.8
R13999 CSoutput.n45 CSoutput.n44 165.8
R14000 CSoutput.n42 CSoutput.n10 165.8
R14001 CSoutput.n41 CSoutput.n40 165.8
R14002 CSoutput.n39 CSoutput.n38 165.8
R14003 CSoutput.n37 CSoutput.n12 165.8
R14004 CSoutput.n35 CSoutput.n34 165.8
R14005 CSoutput.n33 CSoutput.n13 165.8
R14006 CSoutput.n32 CSoutput.n31 165.8
R14007 CSoutput.n29 CSoutput.n14 165.8
R14008 CSoutput.n28 CSoutput.n27 165.8
R14009 CSoutput.n26 CSoutput.n25 165.8
R14010 CSoutput.n24 CSoutput.n16 165.8
R14011 CSoutput.n22 CSoutput.n21 165.8
R14012 CSoutput.n20 CSoutput.n17 165.8
R14013 CSoutput.n77 CSoutput.t138 162.194
R14014 CSoutput.n18 CSoutput.t126 120.501
R14015 CSoutput.n23 CSoutput.t128 120.501
R14016 CSoutput.n15 CSoutput.t139 120.501
R14017 CSoutput.n30 CSoutput.t129 120.501
R14018 CSoutput.n36 CSoutput.t130 120.501
R14019 CSoutput.n11 CSoutput.t124 120.501
R14020 CSoutput.n43 CSoutput.t136 120.501
R14021 CSoutput.n49 CSoutput.t133 120.501
R14022 CSoutput.n7 CSoutput.t127 120.501
R14023 CSoutput.n56 CSoutput.t123 120.501
R14024 CSoutput.n62 CSoutput.t134 120.501
R14025 CSoutput.n64 CSoutput.t135 120.501
R14026 CSoutput.n70 CSoutput.t125 120.501
R14027 CSoutput.n1 CSoutput.t120 120.501
R14028 CSoutput.n270 CSoutput.n268 103.469
R14029 CSoutput.n262 CSoutput.n260 103.469
R14030 CSoutput.n255 CSoutput.n253 103.469
R14031 CSoutput.n96 CSoutput.n94 103.469
R14032 CSoutput.n88 CSoutput.n86 103.469
R14033 CSoutput.n81 CSoutput.n79 103.469
R14034 CSoutput.n272 CSoutput.n271 103.111
R14035 CSoutput.n270 CSoutput.n269 103.111
R14036 CSoutput.n266 CSoutput.n265 103.111
R14037 CSoutput.n264 CSoutput.n263 103.111
R14038 CSoutput.n262 CSoutput.n261 103.111
R14039 CSoutput.n259 CSoutput.n258 103.111
R14040 CSoutput.n257 CSoutput.n256 103.111
R14041 CSoutput.n255 CSoutput.n254 103.111
R14042 CSoutput.n96 CSoutput.n95 103.111
R14043 CSoutput.n98 CSoutput.n97 103.111
R14044 CSoutput.n100 CSoutput.n99 103.111
R14045 CSoutput.n88 CSoutput.n87 103.111
R14046 CSoutput.n90 CSoutput.n89 103.111
R14047 CSoutput.n92 CSoutput.n91 103.111
R14048 CSoutput.n81 CSoutput.n80 103.111
R14049 CSoutput.n83 CSoutput.n82 103.111
R14050 CSoutput.n85 CSoutput.n84 103.111
R14051 CSoutput.n274 CSoutput.n273 103.111
R14052 CSoutput.n302 CSoutput.n300 81.5057
R14053 CSoutput.n290 CSoutput.n288 81.5057
R14054 CSoutput.n279 CSoutput.n277 81.5057
R14055 CSoutput.n338 CSoutput.n336 81.5057
R14056 CSoutput.n326 CSoutput.n324 81.5057
R14057 CSoutput.n315 CSoutput.n313 81.5057
R14058 CSoutput.n310 CSoutput.n309 80.9324
R14059 CSoutput.n308 CSoutput.n307 80.9324
R14060 CSoutput.n306 CSoutput.n305 80.9324
R14061 CSoutput.n304 CSoutput.n303 80.9324
R14062 CSoutput.n302 CSoutput.n301 80.9324
R14063 CSoutput.n298 CSoutput.n297 80.9324
R14064 CSoutput.n296 CSoutput.n295 80.9324
R14065 CSoutput.n294 CSoutput.n293 80.9324
R14066 CSoutput.n292 CSoutput.n291 80.9324
R14067 CSoutput.n290 CSoutput.n289 80.9324
R14068 CSoutput.n287 CSoutput.n286 80.9324
R14069 CSoutput.n285 CSoutput.n284 80.9324
R14070 CSoutput.n283 CSoutput.n282 80.9324
R14071 CSoutput.n281 CSoutput.n280 80.9324
R14072 CSoutput.n279 CSoutput.n278 80.9324
R14073 CSoutput.n338 CSoutput.n337 80.9324
R14074 CSoutput.n340 CSoutput.n339 80.9324
R14075 CSoutput.n342 CSoutput.n341 80.9324
R14076 CSoutput.n344 CSoutput.n343 80.9324
R14077 CSoutput.n346 CSoutput.n345 80.9324
R14078 CSoutput.n326 CSoutput.n325 80.9324
R14079 CSoutput.n328 CSoutput.n327 80.9324
R14080 CSoutput.n330 CSoutput.n329 80.9324
R14081 CSoutput.n332 CSoutput.n331 80.9324
R14082 CSoutput.n334 CSoutput.n333 80.9324
R14083 CSoutput.n315 CSoutput.n314 80.9324
R14084 CSoutput.n317 CSoutput.n316 80.9324
R14085 CSoutput.n319 CSoutput.n318 80.9324
R14086 CSoutput.n321 CSoutput.n320 80.9324
R14087 CSoutput.n323 CSoutput.n322 80.9324
R14088 CSoutput.n25 CSoutput.n24 48.1486
R14089 CSoutput.n69 CSoutput.n3 48.1486
R14090 CSoutput.n38 CSoutput.n37 48.1486
R14091 CSoutput.n42 CSoutput.n41 48.1486
R14092 CSoutput.n51 CSoutput.n50 48.1486
R14093 CSoutput.n55 CSoutput.n54 48.1486
R14094 CSoutput.n22 CSoutput.n17 46.462
R14095 CSoutput.n72 CSoutput.n71 46.462
R14096 CSoutput.n20 CSoutput.n19 44.9055
R14097 CSoutput.n29 CSoutput.n28 43.7635
R14098 CSoutput.n65 CSoutput.n63 43.7635
R14099 CSoutput.n35 CSoutput.n13 41.7396
R14100 CSoutput.n57 CSoutput.n5 41.7396
R14101 CSoutput.n44 CSoutput.n9 37.0171
R14102 CSoutput.n48 CSoutput.n9 37.0171
R14103 CSoutput.n76 CSoutput.n75 34.9932
R14104 CSoutput.n31 CSoutput.n13 32.2947
R14105 CSoutput.n61 CSoutput.n5 32.2947
R14106 CSoutput.n30 CSoutput.n29 29.6014
R14107 CSoutput.n63 CSoutput.n62 29.6014
R14108 CSoutput.n19 CSoutput.n18 28.4085
R14109 CSoutput.n18 CSoutput.n17 25.1176
R14110 CSoutput.n72 CSoutput.n1 25.1176
R14111 CSoutput.n43 CSoutput.n42 22.0922
R14112 CSoutput.n50 CSoutput.n49 22.0922
R14113 CSoutput.n77 CSoutput.n76 21.8586
R14114 CSoutput.n37 CSoutput.n36 18.9681
R14115 CSoutput.n56 CSoutput.n55 18.9681
R14116 CSoutput.n25 CSoutput.n15 17.6292
R14117 CSoutput.n64 CSoutput.n3 17.6292
R14118 CSoutput.n24 CSoutput.n23 15.844
R14119 CSoutput.n70 CSoutput.n69 15.844
R14120 CSoutput.n38 CSoutput.n11 14.5051
R14121 CSoutput.n54 CSoutput.n7 14.5051
R14122 CSoutput.n349 CSoutput.n78 11.4982
R14123 CSoutput.n41 CSoutput.n11 11.3811
R14124 CSoutput.n51 CSoutput.n7 11.3811
R14125 CSoutput.n23 CSoutput.n22 10.0422
R14126 CSoutput.n71 CSoutput.n70 10.0422
R14127 CSoutput.n267 CSoutput.n259 9.25285
R14128 CSoutput.n93 CSoutput.n85 9.25285
R14129 CSoutput.n312 CSoutput.n276 9.07337
R14130 CSoutput.n299 CSoutput.n287 8.98182
R14131 CSoutput.n335 CSoutput.n323 8.98182
R14132 CSoutput.n28 CSoutput.n15 8.25698
R14133 CSoutput.n65 CSoutput.n64 8.25698
R14134 CSoutput.n276 CSoutput.n275 7.12641
R14135 CSoutput.n102 CSoutput.n101 7.12641
R14136 CSoutput.n36 CSoutput.n35 6.91809
R14137 CSoutput.n57 CSoutput.n56 6.91809
R14138 CSoutput.n312 CSoutput.n311 6.02792
R14139 CSoutput.n348 CSoutput.n347 6.02792
R14140 CSoutput.n349 CSoutput.n102 5.48093
R14141 CSoutput.n311 CSoutput.n310 5.25266
R14142 CSoutput.n299 CSoutput.n298 5.25266
R14143 CSoutput.n347 CSoutput.n346 5.25266
R14144 CSoutput.n335 CSoutput.n334 5.25266
R14145 CSoutput.n275 CSoutput.n274 5.1449
R14146 CSoutput.n267 CSoutput.n266 5.1449
R14147 CSoutput.n101 CSoutput.n100 5.1449
R14148 CSoutput.n93 CSoutput.n92 5.1449
R14149 CSoutput.n193 CSoutput.n146 4.5005
R14150 CSoutput.n162 CSoutput.n146 4.5005
R14151 CSoutput.n157 CSoutput.n141 4.5005
R14152 CSoutput.n157 CSoutput.n143 4.5005
R14153 CSoutput.n157 CSoutput.n140 4.5005
R14154 CSoutput.n157 CSoutput.n144 4.5005
R14155 CSoutput.n157 CSoutput.n139 4.5005
R14156 CSoutput.n157 CSoutput.t140 4.5005
R14157 CSoutput.n157 CSoutput.n138 4.5005
R14158 CSoutput.n157 CSoutput.n145 4.5005
R14159 CSoutput.n157 CSoutput.n146 4.5005
R14160 CSoutput.n155 CSoutput.n141 4.5005
R14161 CSoutput.n155 CSoutput.n143 4.5005
R14162 CSoutput.n155 CSoutput.n140 4.5005
R14163 CSoutput.n155 CSoutput.n144 4.5005
R14164 CSoutput.n155 CSoutput.n139 4.5005
R14165 CSoutput.n155 CSoutput.t140 4.5005
R14166 CSoutput.n155 CSoutput.n138 4.5005
R14167 CSoutput.n155 CSoutput.n145 4.5005
R14168 CSoutput.n155 CSoutput.n146 4.5005
R14169 CSoutput.n154 CSoutput.n141 4.5005
R14170 CSoutput.n154 CSoutput.n143 4.5005
R14171 CSoutput.n154 CSoutput.n140 4.5005
R14172 CSoutput.n154 CSoutput.n144 4.5005
R14173 CSoutput.n154 CSoutput.n139 4.5005
R14174 CSoutput.n154 CSoutput.t140 4.5005
R14175 CSoutput.n154 CSoutput.n138 4.5005
R14176 CSoutput.n154 CSoutput.n145 4.5005
R14177 CSoutput.n154 CSoutput.n146 4.5005
R14178 CSoutput.n239 CSoutput.n141 4.5005
R14179 CSoutput.n239 CSoutput.n143 4.5005
R14180 CSoutput.n239 CSoutput.n140 4.5005
R14181 CSoutput.n239 CSoutput.n144 4.5005
R14182 CSoutput.n239 CSoutput.n139 4.5005
R14183 CSoutput.n239 CSoutput.t140 4.5005
R14184 CSoutput.n239 CSoutput.n138 4.5005
R14185 CSoutput.n239 CSoutput.n145 4.5005
R14186 CSoutput.n239 CSoutput.n146 4.5005
R14187 CSoutput.n237 CSoutput.n141 4.5005
R14188 CSoutput.n237 CSoutput.n143 4.5005
R14189 CSoutput.n237 CSoutput.n140 4.5005
R14190 CSoutput.n237 CSoutput.n144 4.5005
R14191 CSoutput.n237 CSoutput.n139 4.5005
R14192 CSoutput.n237 CSoutput.t140 4.5005
R14193 CSoutput.n237 CSoutput.n138 4.5005
R14194 CSoutput.n237 CSoutput.n145 4.5005
R14195 CSoutput.n235 CSoutput.n141 4.5005
R14196 CSoutput.n235 CSoutput.n143 4.5005
R14197 CSoutput.n235 CSoutput.n140 4.5005
R14198 CSoutput.n235 CSoutput.n144 4.5005
R14199 CSoutput.n235 CSoutput.n139 4.5005
R14200 CSoutput.n235 CSoutput.t140 4.5005
R14201 CSoutput.n235 CSoutput.n138 4.5005
R14202 CSoutput.n235 CSoutput.n145 4.5005
R14203 CSoutput.n165 CSoutput.n141 4.5005
R14204 CSoutput.n165 CSoutput.n143 4.5005
R14205 CSoutput.n165 CSoutput.n140 4.5005
R14206 CSoutput.n165 CSoutput.n144 4.5005
R14207 CSoutput.n165 CSoutput.n139 4.5005
R14208 CSoutput.n165 CSoutput.t140 4.5005
R14209 CSoutput.n165 CSoutput.n138 4.5005
R14210 CSoutput.n165 CSoutput.n145 4.5005
R14211 CSoutput.n165 CSoutput.n146 4.5005
R14212 CSoutput.n164 CSoutput.n141 4.5005
R14213 CSoutput.n164 CSoutput.n143 4.5005
R14214 CSoutput.n164 CSoutput.n140 4.5005
R14215 CSoutput.n164 CSoutput.n144 4.5005
R14216 CSoutput.n164 CSoutput.n139 4.5005
R14217 CSoutput.n164 CSoutput.t140 4.5005
R14218 CSoutput.n164 CSoutput.n138 4.5005
R14219 CSoutput.n164 CSoutput.n145 4.5005
R14220 CSoutput.n164 CSoutput.n146 4.5005
R14221 CSoutput.n168 CSoutput.n141 4.5005
R14222 CSoutput.n168 CSoutput.n143 4.5005
R14223 CSoutput.n168 CSoutput.n140 4.5005
R14224 CSoutput.n168 CSoutput.n144 4.5005
R14225 CSoutput.n168 CSoutput.n139 4.5005
R14226 CSoutput.n168 CSoutput.t140 4.5005
R14227 CSoutput.n168 CSoutput.n138 4.5005
R14228 CSoutput.n168 CSoutput.n145 4.5005
R14229 CSoutput.n168 CSoutput.n146 4.5005
R14230 CSoutput.n167 CSoutput.n141 4.5005
R14231 CSoutput.n167 CSoutput.n143 4.5005
R14232 CSoutput.n167 CSoutput.n140 4.5005
R14233 CSoutput.n167 CSoutput.n144 4.5005
R14234 CSoutput.n167 CSoutput.n139 4.5005
R14235 CSoutput.n167 CSoutput.t140 4.5005
R14236 CSoutput.n167 CSoutput.n138 4.5005
R14237 CSoutput.n167 CSoutput.n145 4.5005
R14238 CSoutput.n167 CSoutput.n146 4.5005
R14239 CSoutput.n150 CSoutput.n141 4.5005
R14240 CSoutput.n150 CSoutput.n143 4.5005
R14241 CSoutput.n150 CSoutput.n140 4.5005
R14242 CSoutput.n150 CSoutput.n144 4.5005
R14243 CSoutput.n150 CSoutput.n139 4.5005
R14244 CSoutput.n150 CSoutput.t140 4.5005
R14245 CSoutput.n150 CSoutput.n138 4.5005
R14246 CSoutput.n150 CSoutput.n145 4.5005
R14247 CSoutput.n150 CSoutput.n146 4.5005
R14248 CSoutput.n242 CSoutput.n141 4.5005
R14249 CSoutput.n242 CSoutput.n143 4.5005
R14250 CSoutput.n242 CSoutput.n140 4.5005
R14251 CSoutput.n242 CSoutput.n144 4.5005
R14252 CSoutput.n242 CSoutput.n139 4.5005
R14253 CSoutput.n242 CSoutput.t140 4.5005
R14254 CSoutput.n242 CSoutput.n138 4.5005
R14255 CSoutput.n242 CSoutput.n145 4.5005
R14256 CSoutput.n242 CSoutput.n146 4.5005
R14257 CSoutput.n229 CSoutput.n200 4.5005
R14258 CSoutput.n229 CSoutput.n206 4.5005
R14259 CSoutput.n187 CSoutput.n176 4.5005
R14260 CSoutput.n187 CSoutput.n178 4.5005
R14261 CSoutput.n187 CSoutput.n175 4.5005
R14262 CSoutput.n187 CSoutput.n179 4.5005
R14263 CSoutput.n187 CSoutput.n174 4.5005
R14264 CSoutput.n187 CSoutput.t132 4.5005
R14265 CSoutput.n187 CSoutput.n173 4.5005
R14266 CSoutput.n187 CSoutput.n180 4.5005
R14267 CSoutput.n229 CSoutput.n187 4.5005
R14268 CSoutput.n208 CSoutput.n176 4.5005
R14269 CSoutput.n208 CSoutput.n178 4.5005
R14270 CSoutput.n208 CSoutput.n175 4.5005
R14271 CSoutput.n208 CSoutput.n179 4.5005
R14272 CSoutput.n208 CSoutput.n174 4.5005
R14273 CSoutput.n208 CSoutput.t132 4.5005
R14274 CSoutput.n208 CSoutput.n173 4.5005
R14275 CSoutput.n208 CSoutput.n180 4.5005
R14276 CSoutput.n229 CSoutput.n208 4.5005
R14277 CSoutput.n186 CSoutput.n176 4.5005
R14278 CSoutput.n186 CSoutput.n178 4.5005
R14279 CSoutput.n186 CSoutput.n175 4.5005
R14280 CSoutput.n186 CSoutput.n179 4.5005
R14281 CSoutput.n186 CSoutput.n174 4.5005
R14282 CSoutput.n186 CSoutput.t132 4.5005
R14283 CSoutput.n186 CSoutput.n173 4.5005
R14284 CSoutput.n186 CSoutput.n180 4.5005
R14285 CSoutput.n229 CSoutput.n186 4.5005
R14286 CSoutput.n210 CSoutput.n176 4.5005
R14287 CSoutput.n210 CSoutput.n178 4.5005
R14288 CSoutput.n210 CSoutput.n175 4.5005
R14289 CSoutput.n210 CSoutput.n179 4.5005
R14290 CSoutput.n210 CSoutput.n174 4.5005
R14291 CSoutput.n210 CSoutput.t132 4.5005
R14292 CSoutput.n210 CSoutput.n173 4.5005
R14293 CSoutput.n210 CSoutput.n180 4.5005
R14294 CSoutput.n229 CSoutput.n210 4.5005
R14295 CSoutput.n176 CSoutput.n171 4.5005
R14296 CSoutput.n178 CSoutput.n171 4.5005
R14297 CSoutput.n175 CSoutput.n171 4.5005
R14298 CSoutput.n179 CSoutput.n171 4.5005
R14299 CSoutput.n174 CSoutput.n171 4.5005
R14300 CSoutput.t132 CSoutput.n171 4.5005
R14301 CSoutput.n173 CSoutput.n171 4.5005
R14302 CSoutput.n180 CSoutput.n171 4.5005
R14303 CSoutput.n232 CSoutput.n176 4.5005
R14304 CSoutput.n232 CSoutput.n178 4.5005
R14305 CSoutput.n232 CSoutput.n175 4.5005
R14306 CSoutput.n232 CSoutput.n179 4.5005
R14307 CSoutput.n232 CSoutput.n174 4.5005
R14308 CSoutput.n232 CSoutput.t132 4.5005
R14309 CSoutput.n232 CSoutput.n173 4.5005
R14310 CSoutput.n232 CSoutput.n180 4.5005
R14311 CSoutput.n230 CSoutput.n176 4.5005
R14312 CSoutput.n230 CSoutput.n178 4.5005
R14313 CSoutput.n230 CSoutput.n175 4.5005
R14314 CSoutput.n230 CSoutput.n179 4.5005
R14315 CSoutput.n230 CSoutput.n174 4.5005
R14316 CSoutput.n230 CSoutput.t132 4.5005
R14317 CSoutput.n230 CSoutput.n173 4.5005
R14318 CSoutput.n230 CSoutput.n180 4.5005
R14319 CSoutput.n230 CSoutput.n229 4.5005
R14320 CSoutput.n212 CSoutput.n176 4.5005
R14321 CSoutput.n212 CSoutput.n178 4.5005
R14322 CSoutput.n212 CSoutput.n175 4.5005
R14323 CSoutput.n212 CSoutput.n179 4.5005
R14324 CSoutput.n212 CSoutput.n174 4.5005
R14325 CSoutput.n212 CSoutput.t132 4.5005
R14326 CSoutput.n212 CSoutput.n173 4.5005
R14327 CSoutput.n212 CSoutput.n180 4.5005
R14328 CSoutput.n229 CSoutput.n212 4.5005
R14329 CSoutput.n184 CSoutput.n176 4.5005
R14330 CSoutput.n184 CSoutput.n178 4.5005
R14331 CSoutput.n184 CSoutput.n175 4.5005
R14332 CSoutput.n184 CSoutput.n179 4.5005
R14333 CSoutput.n184 CSoutput.n174 4.5005
R14334 CSoutput.n184 CSoutput.t132 4.5005
R14335 CSoutput.n184 CSoutput.n173 4.5005
R14336 CSoutput.n184 CSoutput.n180 4.5005
R14337 CSoutput.n229 CSoutput.n184 4.5005
R14338 CSoutput.n214 CSoutput.n176 4.5005
R14339 CSoutput.n214 CSoutput.n178 4.5005
R14340 CSoutput.n214 CSoutput.n175 4.5005
R14341 CSoutput.n214 CSoutput.n179 4.5005
R14342 CSoutput.n214 CSoutput.n174 4.5005
R14343 CSoutput.n214 CSoutput.t132 4.5005
R14344 CSoutput.n214 CSoutput.n173 4.5005
R14345 CSoutput.n214 CSoutput.n180 4.5005
R14346 CSoutput.n229 CSoutput.n214 4.5005
R14347 CSoutput.n183 CSoutput.n176 4.5005
R14348 CSoutput.n183 CSoutput.n178 4.5005
R14349 CSoutput.n183 CSoutput.n175 4.5005
R14350 CSoutput.n183 CSoutput.n179 4.5005
R14351 CSoutput.n183 CSoutput.n174 4.5005
R14352 CSoutput.n183 CSoutput.t132 4.5005
R14353 CSoutput.n183 CSoutput.n173 4.5005
R14354 CSoutput.n183 CSoutput.n180 4.5005
R14355 CSoutput.n229 CSoutput.n183 4.5005
R14356 CSoutput.n228 CSoutput.n176 4.5005
R14357 CSoutput.n228 CSoutput.n178 4.5005
R14358 CSoutput.n228 CSoutput.n175 4.5005
R14359 CSoutput.n228 CSoutput.n179 4.5005
R14360 CSoutput.n228 CSoutput.n174 4.5005
R14361 CSoutput.n228 CSoutput.t132 4.5005
R14362 CSoutput.n228 CSoutput.n173 4.5005
R14363 CSoutput.n228 CSoutput.n180 4.5005
R14364 CSoutput.n229 CSoutput.n228 4.5005
R14365 CSoutput.n227 CSoutput.n112 4.5005
R14366 CSoutput.n128 CSoutput.n112 4.5005
R14367 CSoutput.n123 CSoutput.n107 4.5005
R14368 CSoutput.n123 CSoutput.n109 4.5005
R14369 CSoutput.n123 CSoutput.n106 4.5005
R14370 CSoutput.n123 CSoutput.n110 4.5005
R14371 CSoutput.n123 CSoutput.n105 4.5005
R14372 CSoutput.n123 CSoutput.t131 4.5005
R14373 CSoutput.n123 CSoutput.n104 4.5005
R14374 CSoutput.n123 CSoutput.n111 4.5005
R14375 CSoutput.n123 CSoutput.n112 4.5005
R14376 CSoutput.n121 CSoutput.n107 4.5005
R14377 CSoutput.n121 CSoutput.n109 4.5005
R14378 CSoutput.n121 CSoutput.n106 4.5005
R14379 CSoutput.n121 CSoutput.n110 4.5005
R14380 CSoutput.n121 CSoutput.n105 4.5005
R14381 CSoutput.n121 CSoutput.t131 4.5005
R14382 CSoutput.n121 CSoutput.n104 4.5005
R14383 CSoutput.n121 CSoutput.n111 4.5005
R14384 CSoutput.n121 CSoutput.n112 4.5005
R14385 CSoutput.n120 CSoutput.n107 4.5005
R14386 CSoutput.n120 CSoutput.n109 4.5005
R14387 CSoutput.n120 CSoutput.n106 4.5005
R14388 CSoutput.n120 CSoutput.n110 4.5005
R14389 CSoutput.n120 CSoutput.n105 4.5005
R14390 CSoutput.n120 CSoutput.t131 4.5005
R14391 CSoutput.n120 CSoutput.n104 4.5005
R14392 CSoutput.n120 CSoutput.n111 4.5005
R14393 CSoutput.n120 CSoutput.n112 4.5005
R14394 CSoutput.n249 CSoutput.n107 4.5005
R14395 CSoutput.n249 CSoutput.n109 4.5005
R14396 CSoutput.n249 CSoutput.n106 4.5005
R14397 CSoutput.n249 CSoutput.n110 4.5005
R14398 CSoutput.n249 CSoutput.n105 4.5005
R14399 CSoutput.n249 CSoutput.t131 4.5005
R14400 CSoutput.n249 CSoutput.n104 4.5005
R14401 CSoutput.n249 CSoutput.n111 4.5005
R14402 CSoutput.n249 CSoutput.n112 4.5005
R14403 CSoutput.n247 CSoutput.n107 4.5005
R14404 CSoutput.n247 CSoutput.n109 4.5005
R14405 CSoutput.n247 CSoutput.n106 4.5005
R14406 CSoutput.n247 CSoutput.n110 4.5005
R14407 CSoutput.n247 CSoutput.n105 4.5005
R14408 CSoutput.n247 CSoutput.t131 4.5005
R14409 CSoutput.n247 CSoutput.n104 4.5005
R14410 CSoutput.n247 CSoutput.n111 4.5005
R14411 CSoutput.n245 CSoutput.n107 4.5005
R14412 CSoutput.n245 CSoutput.n109 4.5005
R14413 CSoutput.n245 CSoutput.n106 4.5005
R14414 CSoutput.n245 CSoutput.n110 4.5005
R14415 CSoutput.n245 CSoutput.n105 4.5005
R14416 CSoutput.n245 CSoutput.t131 4.5005
R14417 CSoutput.n245 CSoutput.n104 4.5005
R14418 CSoutput.n245 CSoutput.n111 4.5005
R14419 CSoutput.n131 CSoutput.n107 4.5005
R14420 CSoutput.n131 CSoutput.n109 4.5005
R14421 CSoutput.n131 CSoutput.n106 4.5005
R14422 CSoutput.n131 CSoutput.n110 4.5005
R14423 CSoutput.n131 CSoutput.n105 4.5005
R14424 CSoutput.n131 CSoutput.t131 4.5005
R14425 CSoutput.n131 CSoutput.n104 4.5005
R14426 CSoutput.n131 CSoutput.n111 4.5005
R14427 CSoutput.n131 CSoutput.n112 4.5005
R14428 CSoutput.n130 CSoutput.n107 4.5005
R14429 CSoutput.n130 CSoutput.n109 4.5005
R14430 CSoutput.n130 CSoutput.n106 4.5005
R14431 CSoutput.n130 CSoutput.n110 4.5005
R14432 CSoutput.n130 CSoutput.n105 4.5005
R14433 CSoutput.n130 CSoutput.t131 4.5005
R14434 CSoutput.n130 CSoutput.n104 4.5005
R14435 CSoutput.n130 CSoutput.n111 4.5005
R14436 CSoutput.n130 CSoutput.n112 4.5005
R14437 CSoutput.n134 CSoutput.n107 4.5005
R14438 CSoutput.n134 CSoutput.n109 4.5005
R14439 CSoutput.n134 CSoutput.n106 4.5005
R14440 CSoutput.n134 CSoutput.n110 4.5005
R14441 CSoutput.n134 CSoutput.n105 4.5005
R14442 CSoutput.n134 CSoutput.t131 4.5005
R14443 CSoutput.n134 CSoutput.n104 4.5005
R14444 CSoutput.n134 CSoutput.n111 4.5005
R14445 CSoutput.n134 CSoutput.n112 4.5005
R14446 CSoutput.n133 CSoutput.n107 4.5005
R14447 CSoutput.n133 CSoutput.n109 4.5005
R14448 CSoutput.n133 CSoutput.n106 4.5005
R14449 CSoutput.n133 CSoutput.n110 4.5005
R14450 CSoutput.n133 CSoutput.n105 4.5005
R14451 CSoutput.n133 CSoutput.t131 4.5005
R14452 CSoutput.n133 CSoutput.n104 4.5005
R14453 CSoutput.n133 CSoutput.n111 4.5005
R14454 CSoutput.n133 CSoutput.n112 4.5005
R14455 CSoutput.n116 CSoutput.n107 4.5005
R14456 CSoutput.n116 CSoutput.n109 4.5005
R14457 CSoutput.n116 CSoutput.n106 4.5005
R14458 CSoutput.n116 CSoutput.n110 4.5005
R14459 CSoutput.n116 CSoutput.n105 4.5005
R14460 CSoutput.n116 CSoutput.t131 4.5005
R14461 CSoutput.n116 CSoutput.n104 4.5005
R14462 CSoutput.n116 CSoutput.n111 4.5005
R14463 CSoutput.n116 CSoutput.n112 4.5005
R14464 CSoutput.n252 CSoutput.n107 4.5005
R14465 CSoutput.n252 CSoutput.n109 4.5005
R14466 CSoutput.n252 CSoutput.n106 4.5005
R14467 CSoutput.n252 CSoutput.n110 4.5005
R14468 CSoutput.n252 CSoutput.n105 4.5005
R14469 CSoutput.n252 CSoutput.t131 4.5005
R14470 CSoutput.n252 CSoutput.n104 4.5005
R14471 CSoutput.n252 CSoutput.n111 4.5005
R14472 CSoutput.n252 CSoutput.n112 4.5005
R14473 CSoutput.n275 CSoutput.n267 4.10845
R14474 CSoutput.n101 CSoutput.n93 4.10845
R14475 CSoutput.n273 CSoutput.t109 4.06363
R14476 CSoutput.n273 CSoutput.t118 4.06363
R14477 CSoutput.n271 CSoutput.t101 4.06363
R14478 CSoutput.n271 CSoutput.t116 4.06363
R14479 CSoutput.n269 CSoutput.t93 4.06363
R14480 CSoutput.n269 CSoutput.t73 4.06363
R14481 CSoutput.n268 CSoutput.t102 4.06363
R14482 CSoutput.n268 CSoutput.t103 4.06363
R14483 CSoutput.n265 CSoutput.t72 4.06363
R14484 CSoutput.n265 CSoutput.t104 4.06363
R14485 CSoutput.n263 CSoutput.t94 4.06363
R14486 CSoutput.n263 CSoutput.t78 4.06363
R14487 CSoutput.n261 CSoutput.t79 4.06363
R14488 CSoutput.n261 CSoutput.t81 4.06363
R14489 CSoutput.n260 CSoutput.t98 4.06363
R14490 CSoutput.n260 CSoutput.t99 4.06363
R14491 CSoutput.n258 CSoutput.t117 4.06363
R14492 CSoutput.n258 CSoutput.t107 4.06363
R14493 CSoutput.n256 CSoutput.t91 4.06363
R14494 CSoutput.n256 CSoutput.t111 4.06363
R14495 CSoutput.n254 CSoutput.t97 4.06363
R14496 CSoutput.n254 CSoutput.t108 4.06363
R14497 CSoutput.n253 CSoutput.t88 4.06363
R14498 CSoutput.n253 CSoutput.t84 4.06363
R14499 CSoutput.n94 CSoutput.t76 4.06363
R14500 CSoutput.n94 CSoutput.t77 4.06363
R14501 CSoutput.n95 CSoutput.t115 4.06363
R14502 CSoutput.n95 CSoutput.t74 4.06363
R14503 CSoutput.n97 CSoutput.t110 4.06363
R14504 CSoutput.n97 CSoutput.t75 4.06363
R14505 CSoutput.n99 CSoutput.t114 4.06363
R14506 CSoutput.n99 CSoutput.t100 4.06363
R14507 CSoutput.n86 CSoutput.t83 4.06363
R14508 CSoutput.n86 CSoutput.t92 4.06363
R14509 CSoutput.n87 CSoutput.t87 4.06363
R14510 CSoutput.n87 CSoutput.t82 4.06363
R14511 CSoutput.n89 CSoutput.t89 4.06363
R14512 CSoutput.n89 CSoutput.t112 4.06363
R14513 CSoutput.n91 CSoutput.t86 4.06363
R14514 CSoutput.n91 CSoutput.t119 4.06363
R14515 CSoutput.n79 CSoutput.t85 4.06363
R14516 CSoutput.n79 CSoutput.t96 4.06363
R14517 CSoutput.n80 CSoutput.t80 4.06363
R14518 CSoutput.n80 CSoutput.t95 4.06363
R14519 CSoutput.n82 CSoutput.t113 4.06363
R14520 CSoutput.n82 CSoutput.t90 4.06363
R14521 CSoutput.n84 CSoutput.t106 4.06363
R14522 CSoutput.n84 CSoutput.t105 4.06363
R14523 CSoutput.n44 CSoutput.n43 3.79402
R14524 CSoutput.n49 CSoutput.n48 3.79402
R14525 CSoutput.n311 CSoutput.n299 3.72967
R14526 CSoutput.n347 CSoutput.n335 3.72967
R14527 CSoutput.n349 CSoutput.n348 3.57343
R14528 CSoutput.n348 CSoutput.n312 3.04641
R14529 CSoutput.n309 CSoutput.t44 2.82907
R14530 CSoutput.n309 CSoutput.t2 2.82907
R14531 CSoutput.n307 CSoutput.t70 2.82907
R14532 CSoutput.n307 CSoutput.t60 2.82907
R14533 CSoutput.n305 CSoutput.t26 2.82907
R14534 CSoutput.n305 CSoutput.t35 2.82907
R14535 CSoutput.n303 CSoutput.t1 2.82907
R14536 CSoutput.n303 CSoutput.t67 2.82907
R14537 CSoutput.n301 CSoutput.t59 2.82907
R14538 CSoutput.n301 CSoutput.t15 2.82907
R14539 CSoutput.n300 CSoutput.t8 2.82907
R14540 CSoutput.n300 CSoutput.t69 2.82907
R14541 CSoutput.n297 CSoutput.t12 2.82907
R14542 CSoutput.n297 CSoutput.t22 2.82907
R14543 CSoutput.n295 CSoutput.t21 2.82907
R14544 CSoutput.n295 CSoutput.t7 2.82907
R14545 CSoutput.n293 CSoutput.t33 2.82907
R14546 CSoutput.n293 CSoutput.t11 2.82907
R14547 CSoutput.n291 CSoutput.t14 2.82907
R14548 CSoutput.n291 CSoutput.t20 2.82907
R14549 CSoutput.n289 CSoutput.t18 2.82907
R14550 CSoutput.n289 CSoutput.t31 2.82907
R14551 CSoutput.n288 CSoutput.t30 2.82907
R14552 CSoutput.n288 CSoutput.t13 2.82907
R14553 CSoutput.n286 CSoutput.t53 2.82907
R14554 CSoutput.n286 CSoutput.t24 2.82907
R14555 CSoutput.n284 CSoutput.t4 2.82907
R14556 CSoutput.n284 CSoutput.t40 2.82907
R14557 CSoutput.n282 CSoutput.t19 2.82907
R14558 CSoutput.n282 CSoutput.t32 2.82907
R14559 CSoutput.n280 CSoutput.t34 2.82907
R14560 CSoutput.n280 CSoutput.t65 2.82907
R14561 CSoutput.n278 CSoutput.t50 2.82907
R14562 CSoutput.n278 CSoutput.t0 2.82907
R14563 CSoutput.n277 CSoutput.t63 2.82907
R14564 CSoutput.n277 CSoutput.t10 2.82907
R14565 CSoutput.n336 CSoutput.t57 2.82907
R14566 CSoutput.n336 CSoutput.t68 2.82907
R14567 CSoutput.n337 CSoutput.t71 2.82907
R14568 CSoutput.n337 CSoutput.t48 2.82907
R14569 CSoutput.n339 CSoutput.t52 2.82907
R14570 CSoutput.n339 CSoutput.t62 2.82907
R14571 CSoutput.n341 CSoutput.t9 2.82907
R14572 CSoutput.n341 CSoutput.t42 2.82907
R14573 CSoutput.n343 CSoutput.t47 2.82907
R14574 CSoutput.n343 CSoutput.t58 2.82907
R14575 CSoutput.n345 CSoutput.t64 2.82907
R14576 CSoutput.n345 CSoutput.t51 2.82907
R14577 CSoutput.n324 CSoutput.t28 2.82907
R14578 CSoutput.n324 CSoutput.t45 2.82907
R14579 CSoutput.n325 CSoutput.t46 2.82907
R14580 CSoutput.n325 CSoutput.t36 2.82907
R14581 CSoutput.n327 CSoutput.t37 2.82907
R14582 CSoutput.n327 CSoutput.t29 2.82907
R14583 CSoutput.n329 CSoutput.t23 2.82907
R14584 CSoutput.n329 CSoutput.t16 2.82907
R14585 CSoutput.n331 CSoutput.t17 2.82907
R14586 CSoutput.n331 CSoutput.t38 2.82907
R14587 CSoutput.n333 CSoutput.t39 2.82907
R14588 CSoutput.n333 CSoutput.t3 2.82907
R14589 CSoutput.n313 CSoutput.t41 2.82907
R14590 CSoutput.n313 CSoutput.t5 2.82907
R14591 CSoutput.n314 CSoutput.t25 2.82907
R14592 CSoutput.n314 CSoutput.t66 2.82907
R14593 CSoutput.n316 CSoutput.t6 2.82907
R14594 CSoutput.n316 CSoutput.t55 2.82907
R14595 CSoutput.n318 CSoutput.t54 2.82907
R14596 CSoutput.n318 CSoutput.t43 2.82907
R14597 CSoutput.n320 CSoutput.t56 2.82907
R14598 CSoutput.n320 CSoutput.t27 2.82907
R14599 CSoutput.n322 CSoutput.t49 2.82907
R14600 CSoutput.n322 CSoutput.t61 2.82907
R14601 CSoutput.n75 CSoutput.n1 2.45513
R14602 CSoutput.n193 CSoutput.n191 2.251
R14603 CSoutput.n193 CSoutput.n190 2.251
R14604 CSoutput.n193 CSoutput.n189 2.251
R14605 CSoutput.n193 CSoutput.n188 2.251
R14606 CSoutput.n162 CSoutput.n161 2.251
R14607 CSoutput.n162 CSoutput.n160 2.251
R14608 CSoutput.n162 CSoutput.n159 2.251
R14609 CSoutput.n162 CSoutput.n158 2.251
R14610 CSoutput.n235 CSoutput.n234 2.251
R14611 CSoutput.n200 CSoutput.n198 2.251
R14612 CSoutput.n200 CSoutput.n197 2.251
R14613 CSoutput.n200 CSoutput.n196 2.251
R14614 CSoutput.n218 CSoutput.n200 2.251
R14615 CSoutput.n206 CSoutput.n205 2.251
R14616 CSoutput.n206 CSoutput.n204 2.251
R14617 CSoutput.n206 CSoutput.n203 2.251
R14618 CSoutput.n206 CSoutput.n202 2.251
R14619 CSoutput.n232 CSoutput.n172 2.251
R14620 CSoutput.n227 CSoutput.n225 2.251
R14621 CSoutput.n227 CSoutput.n224 2.251
R14622 CSoutput.n227 CSoutput.n223 2.251
R14623 CSoutput.n227 CSoutput.n222 2.251
R14624 CSoutput.n128 CSoutput.n127 2.251
R14625 CSoutput.n128 CSoutput.n126 2.251
R14626 CSoutput.n128 CSoutput.n125 2.251
R14627 CSoutput.n128 CSoutput.n124 2.251
R14628 CSoutput.n245 CSoutput.n244 2.251
R14629 CSoutput.n162 CSoutput.n142 2.2505
R14630 CSoutput.n157 CSoutput.n142 2.2505
R14631 CSoutput.n155 CSoutput.n142 2.2505
R14632 CSoutput.n154 CSoutput.n142 2.2505
R14633 CSoutput.n239 CSoutput.n142 2.2505
R14634 CSoutput.n237 CSoutput.n142 2.2505
R14635 CSoutput.n235 CSoutput.n142 2.2505
R14636 CSoutput.n165 CSoutput.n142 2.2505
R14637 CSoutput.n164 CSoutput.n142 2.2505
R14638 CSoutput.n168 CSoutput.n142 2.2505
R14639 CSoutput.n167 CSoutput.n142 2.2505
R14640 CSoutput.n150 CSoutput.n142 2.2505
R14641 CSoutput.n242 CSoutput.n142 2.2505
R14642 CSoutput.n242 CSoutput.n241 2.2505
R14643 CSoutput.n206 CSoutput.n177 2.2505
R14644 CSoutput.n187 CSoutput.n177 2.2505
R14645 CSoutput.n208 CSoutput.n177 2.2505
R14646 CSoutput.n186 CSoutput.n177 2.2505
R14647 CSoutput.n210 CSoutput.n177 2.2505
R14648 CSoutput.n177 CSoutput.n171 2.2505
R14649 CSoutput.n232 CSoutput.n177 2.2505
R14650 CSoutput.n230 CSoutput.n177 2.2505
R14651 CSoutput.n212 CSoutput.n177 2.2505
R14652 CSoutput.n184 CSoutput.n177 2.2505
R14653 CSoutput.n214 CSoutput.n177 2.2505
R14654 CSoutput.n183 CSoutput.n177 2.2505
R14655 CSoutput.n228 CSoutput.n177 2.2505
R14656 CSoutput.n228 CSoutput.n181 2.2505
R14657 CSoutput.n128 CSoutput.n108 2.2505
R14658 CSoutput.n123 CSoutput.n108 2.2505
R14659 CSoutput.n121 CSoutput.n108 2.2505
R14660 CSoutput.n120 CSoutput.n108 2.2505
R14661 CSoutput.n249 CSoutput.n108 2.2505
R14662 CSoutput.n247 CSoutput.n108 2.2505
R14663 CSoutput.n245 CSoutput.n108 2.2505
R14664 CSoutput.n131 CSoutput.n108 2.2505
R14665 CSoutput.n130 CSoutput.n108 2.2505
R14666 CSoutput.n134 CSoutput.n108 2.2505
R14667 CSoutput.n133 CSoutput.n108 2.2505
R14668 CSoutput.n116 CSoutput.n108 2.2505
R14669 CSoutput.n252 CSoutput.n108 2.2505
R14670 CSoutput.n252 CSoutput.n251 2.2505
R14671 CSoutput.n170 CSoutput.n163 2.25024
R14672 CSoutput.n170 CSoutput.n156 2.25024
R14673 CSoutput.n238 CSoutput.n170 2.25024
R14674 CSoutput.n170 CSoutput.n166 2.25024
R14675 CSoutput.n170 CSoutput.n169 2.25024
R14676 CSoutput.n170 CSoutput.n137 2.25024
R14677 CSoutput.n220 CSoutput.n217 2.25024
R14678 CSoutput.n220 CSoutput.n216 2.25024
R14679 CSoutput.n220 CSoutput.n215 2.25024
R14680 CSoutput.n220 CSoutput.n182 2.25024
R14681 CSoutput.n220 CSoutput.n219 2.25024
R14682 CSoutput.n221 CSoutput.n220 2.25024
R14683 CSoutput.n136 CSoutput.n129 2.25024
R14684 CSoutput.n136 CSoutput.n122 2.25024
R14685 CSoutput.n248 CSoutput.n136 2.25024
R14686 CSoutput.n136 CSoutput.n132 2.25024
R14687 CSoutput.n136 CSoutput.n135 2.25024
R14688 CSoutput.n136 CSoutput.n103 2.25024
R14689 CSoutput.n276 CSoutput.n102 1.95131
R14690 CSoutput.n237 CSoutput.n147 1.50111
R14691 CSoutput.n185 CSoutput.n171 1.50111
R14692 CSoutput.n247 CSoutput.n113 1.50111
R14693 CSoutput.n193 CSoutput.n192 1.501
R14694 CSoutput.n200 CSoutput.n199 1.501
R14695 CSoutput.n227 CSoutput.n226 1.501
R14696 CSoutput.n241 CSoutput.n152 1.12536
R14697 CSoutput.n241 CSoutput.n153 1.12536
R14698 CSoutput.n241 CSoutput.n240 1.12536
R14699 CSoutput.n201 CSoutput.n181 1.12536
R14700 CSoutput.n207 CSoutput.n181 1.12536
R14701 CSoutput.n209 CSoutput.n181 1.12536
R14702 CSoutput.n251 CSoutput.n118 1.12536
R14703 CSoutput.n251 CSoutput.n119 1.12536
R14704 CSoutput.n251 CSoutput.n250 1.12536
R14705 CSoutput.n241 CSoutput.n148 1.12536
R14706 CSoutput.n241 CSoutput.n149 1.12536
R14707 CSoutput.n241 CSoutput.n151 1.12536
R14708 CSoutput.n231 CSoutput.n181 1.12536
R14709 CSoutput.n211 CSoutput.n181 1.12536
R14710 CSoutput.n213 CSoutput.n181 1.12536
R14711 CSoutput.n251 CSoutput.n114 1.12536
R14712 CSoutput.n251 CSoutput.n115 1.12536
R14713 CSoutput.n251 CSoutput.n117 1.12536
R14714 CSoutput.n31 CSoutput.n30 0.669944
R14715 CSoutput.n62 CSoutput.n61 0.669944
R14716 CSoutput.n304 CSoutput.n302 0.573776
R14717 CSoutput.n306 CSoutput.n304 0.573776
R14718 CSoutput.n308 CSoutput.n306 0.573776
R14719 CSoutput.n310 CSoutput.n308 0.573776
R14720 CSoutput.n292 CSoutput.n290 0.573776
R14721 CSoutput.n294 CSoutput.n292 0.573776
R14722 CSoutput.n296 CSoutput.n294 0.573776
R14723 CSoutput.n298 CSoutput.n296 0.573776
R14724 CSoutput.n281 CSoutput.n279 0.573776
R14725 CSoutput.n283 CSoutput.n281 0.573776
R14726 CSoutput.n285 CSoutput.n283 0.573776
R14727 CSoutput.n287 CSoutput.n285 0.573776
R14728 CSoutput.n346 CSoutput.n344 0.573776
R14729 CSoutput.n344 CSoutput.n342 0.573776
R14730 CSoutput.n342 CSoutput.n340 0.573776
R14731 CSoutput.n340 CSoutput.n338 0.573776
R14732 CSoutput.n334 CSoutput.n332 0.573776
R14733 CSoutput.n332 CSoutput.n330 0.573776
R14734 CSoutput.n330 CSoutput.n328 0.573776
R14735 CSoutput.n328 CSoutput.n326 0.573776
R14736 CSoutput.n323 CSoutput.n321 0.573776
R14737 CSoutput.n321 CSoutput.n319 0.573776
R14738 CSoutput.n319 CSoutput.n317 0.573776
R14739 CSoutput.n317 CSoutput.n315 0.573776
R14740 CSoutput.n349 CSoutput.n252 0.53442
R14741 CSoutput.n272 CSoutput.n270 0.358259
R14742 CSoutput.n274 CSoutput.n272 0.358259
R14743 CSoutput.n264 CSoutput.n262 0.358259
R14744 CSoutput.n266 CSoutput.n264 0.358259
R14745 CSoutput.n257 CSoutput.n255 0.358259
R14746 CSoutput.n259 CSoutput.n257 0.358259
R14747 CSoutput.n100 CSoutput.n98 0.358259
R14748 CSoutput.n98 CSoutput.n96 0.358259
R14749 CSoutput.n92 CSoutput.n90 0.358259
R14750 CSoutput.n90 CSoutput.n88 0.358259
R14751 CSoutput.n85 CSoutput.n83 0.358259
R14752 CSoutput.n83 CSoutput.n81 0.358259
R14753 CSoutput.n21 CSoutput.n20 0.169105
R14754 CSoutput.n21 CSoutput.n16 0.169105
R14755 CSoutput.n26 CSoutput.n16 0.169105
R14756 CSoutput.n27 CSoutput.n26 0.169105
R14757 CSoutput.n27 CSoutput.n14 0.169105
R14758 CSoutput.n32 CSoutput.n14 0.169105
R14759 CSoutput.n33 CSoutput.n32 0.169105
R14760 CSoutput.n34 CSoutput.n33 0.169105
R14761 CSoutput.n34 CSoutput.n12 0.169105
R14762 CSoutput.n39 CSoutput.n12 0.169105
R14763 CSoutput.n40 CSoutput.n39 0.169105
R14764 CSoutput.n40 CSoutput.n10 0.169105
R14765 CSoutput.n45 CSoutput.n10 0.169105
R14766 CSoutput.n46 CSoutput.n45 0.169105
R14767 CSoutput.n47 CSoutput.n46 0.169105
R14768 CSoutput.n47 CSoutput.n8 0.169105
R14769 CSoutput.n52 CSoutput.n8 0.169105
R14770 CSoutput.n53 CSoutput.n52 0.169105
R14771 CSoutput.n53 CSoutput.n6 0.169105
R14772 CSoutput.n58 CSoutput.n6 0.169105
R14773 CSoutput.n59 CSoutput.n58 0.169105
R14774 CSoutput.n60 CSoutput.n59 0.169105
R14775 CSoutput.n60 CSoutput.n4 0.169105
R14776 CSoutput.n66 CSoutput.n4 0.169105
R14777 CSoutput.n67 CSoutput.n66 0.169105
R14778 CSoutput.n68 CSoutput.n67 0.169105
R14779 CSoutput.n68 CSoutput.n2 0.169105
R14780 CSoutput.n73 CSoutput.n2 0.169105
R14781 CSoutput.n74 CSoutput.n73 0.169105
R14782 CSoutput.n74 CSoutput.n0 0.169105
R14783 CSoutput.n78 CSoutput.n0 0.169105
R14784 CSoutput.n195 CSoutput.n194 0.0910737
R14785 CSoutput.n246 CSoutput.n243 0.0723685
R14786 CSoutput.n200 CSoutput.n195 0.0522944
R14787 CSoutput.n243 CSoutput.n242 0.0499135
R14788 CSoutput.n194 CSoutput.n193 0.0499135
R14789 CSoutput.n228 CSoutput.n227 0.0464294
R14790 CSoutput.n236 CSoutput.n233 0.0391444
R14791 CSoutput.n195 CSoutput.t141 0.023435
R14792 CSoutput.n243 CSoutput.t121 0.02262
R14793 CSoutput.n194 CSoutput.t122 0.02262
R14794 CSoutput CSoutput.n349 0.0052
R14795 CSoutput.n165 CSoutput.n148 0.00365111
R14796 CSoutput.n168 CSoutput.n149 0.00365111
R14797 CSoutput.n151 CSoutput.n150 0.00365111
R14798 CSoutput.n193 CSoutput.n152 0.00365111
R14799 CSoutput.n157 CSoutput.n153 0.00365111
R14800 CSoutput.n240 CSoutput.n154 0.00365111
R14801 CSoutput.n231 CSoutput.n230 0.00365111
R14802 CSoutput.n211 CSoutput.n184 0.00365111
R14803 CSoutput.n213 CSoutput.n183 0.00365111
R14804 CSoutput.n201 CSoutput.n200 0.00365111
R14805 CSoutput.n207 CSoutput.n187 0.00365111
R14806 CSoutput.n209 CSoutput.n186 0.00365111
R14807 CSoutput.n131 CSoutput.n114 0.00365111
R14808 CSoutput.n134 CSoutput.n115 0.00365111
R14809 CSoutput.n117 CSoutput.n116 0.00365111
R14810 CSoutput.n227 CSoutput.n118 0.00365111
R14811 CSoutput.n123 CSoutput.n119 0.00365111
R14812 CSoutput.n250 CSoutput.n120 0.00365111
R14813 CSoutput.n162 CSoutput.n152 0.00340054
R14814 CSoutput.n155 CSoutput.n153 0.00340054
R14815 CSoutput.n240 CSoutput.n239 0.00340054
R14816 CSoutput.n235 CSoutput.n148 0.00340054
R14817 CSoutput.n164 CSoutput.n149 0.00340054
R14818 CSoutput.n167 CSoutput.n151 0.00340054
R14819 CSoutput.n206 CSoutput.n201 0.00340054
R14820 CSoutput.n208 CSoutput.n207 0.00340054
R14821 CSoutput.n210 CSoutput.n209 0.00340054
R14822 CSoutput.n232 CSoutput.n231 0.00340054
R14823 CSoutput.n212 CSoutput.n211 0.00340054
R14824 CSoutput.n214 CSoutput.n213 0.00340054
R14825 CSoutput.n128 CSoutput.n118 0.00340054
R14826 CSoutput.n121 CSoutput.n119 0.00340054
R14827 CSoutput.n250 CSoutput.n249 0.00340054
R14828 CSoutput.n245 CSoutput.n114 0.00340054
R14829 CSoutput.n130 CSoutput.n115 0.00340054
R14830 CSoutput.n133 CSoutput.n117 0.00340054
R14831 CSoutput.n163 CSoutput.n157 0.00252698
R14832 CSoutput.n156 CSoutput.n154 0.00252698
R14833 CSoutput.n238 CSoutput.n237 0.00252698
R14834 CSoutput.n166 CSoutput.n164 0.00252698
R14835 CSoutput.n169 CSoutput.n167 0.00252698
R14836 CSoutput.n242 CSoutput.n137 0.00252698
R14837 CSoutput.n163 CSoutput.n162 0.00252698
R14838 CSoutput.n156 CSoutput.n155 0.00252698
R14839 CSoutput.n239 CSoutput.n238 0.00252698
R14840 CSoutput.n166 CSoutput.n165 0.00252698
R14841 CSoutput.n169 CSoutput.n168 0.00252698
R14842 CSoutput.n150 CSoutput.n137 0.00252698
R14843 CSoutput.n217 CSoutput.n187 0.00252698
R14844 CSoutput.n216 CSoutput.n186 0.00252698
R14845 CSoutput.n215 CSoutput.n171 0.00252698
R14846 CSoutput.n212 CSoutput.n182 0.00252698
R14847 CSoutput.n219 CSoutput.n214 0.00252698
R14848 CSoutput.n228 CSoutput.n221 0.00252698
R14849 CSoutput.n217 CSoutput.n206 0.00252698
R14850 CSoutput.n216 CSoutput.n208 0.00252698
R14851 CSoutput.n215 CSoutput.n210 0.00252698
R14852 CSoutput.n230 CSoutput.n182 0.00252698
R14853 CSoutput.n219 CSoutput.n184 0.00252698
R14854 CSoutput.n221 CSoutput.n183 0.00252698
R14855 CSoutput.n129 CSoutput.n123 0.00252698
R14856 CSoutput.n122 CSoutput.n120 0.00252698
R14857 CSoutput.n248 CSoutput.n247 0.00252698
R14858 CSoutput.n132 CSoutput.n130 0.00252698
R14859 CSoutput.n135 CSoutput.n133 0.00252698
R14860 CSoutput.n252 CSoutput.n103 0.00252698
R14861 CSoutput.n129 CSoutput.n128 0.00252698
R14862 CSoutput.n122 CSoutput.n121 0.00252698
R14863 CSoutput.n249 CSoutput.n248 0.00252698
R14864 CSoutput.n132 CSoutput.n131 0.00252698
R14865 CSoutput.n135 CSoutput.n134 0.00252698
R14866 CSoutput.n116 CSoutput.n103 0.00252698
R14867 CSoutput.n237 CSoutput.n236 0.0020275
R14868 CSoutput.n236 CSoutput.n235 0.0020275
R14869 CSoutput.n233 CSoutput.n171 0.0020275
R14870 CSoutput.n233 CSoutput.n232 0.0020275
R14871 CSoutput.n247 CSoutput.n246 0.0020275
R14872 CSoutput.n246 CSoutput.n245 0.0020275
R14873 CSoutput.n147 CSoutput.n146 0.00166668
R14874 CSoutput.n229 CSoutput.n185 0.00166668
R14875 CSoutput.n113 CSoutput.n112 0.00166668
R14876 CSoutput.n251 CSoutput.n113 0.00133328
R14877 CSoutput.n185 CSoutput.n181 0.00133328
R14878 CSoutput.n241 CSoutput.n147 0.00133328
R14879 CSoutput.n244 CSoutput.n136 0.001
R14880 CSoutput.n222 CSoutput.n136 0.001
R14881 CSoutput.n124 CSoutput.n104 0.001
R14882 CSoutput.n223 CSoutput.n104 0.001
R14883 CSoutput.n125 CSoutput.n105 0.001
R14884 CSoutput.n224 CSoutput.n105 0.001
R14885 CSoutput.n126 CSoutput.n106 0.001
R14886 CSoutput.n225 CSoutput.n106 0.001
R14887 CSoutput.n127 CSoutput.n107 0.001
R14888 CSoutput.n226 CSoutput.n107 0.001
R14889 CSoutput.n220 CSoutput.n172 0.001
R14890 CSoutput.n220 CSoutput.n218 0.001
R14891 CSoutput.n202 CSoutput.n173 0.001
R14892 CSoutput.n196 CSoutput.n173 0.001
R14893 CSoutput.n203 CSoutput.n174 0.001
R14894 CSoutput.n197 CSoutput.n174 0.001
R14895 CSoutput.n204 CSoutput.n175 0.001
R14896 CSoutput.n198 CSoutput.n175 0.001
R14897 CSoutput.n205 CSoutput.n176 0.001
R14898 CSoutput.n199 CSoutput.n176 0.001
R14899 CSoutput.n234 CSoutput.n170 0.001
R14900 CSoutput.n188 CSoutput.n170 0.001
R14901 CSoutput.n158 CSoutput.n138 0.001
R14902 CSoutput.n189 CSoutput.n138 0.001
R14903 CSoutput.n159 CSoutput.n139 0.001
R14904 CSoutput.n190 CSoutput.n139 0.001
R14905 CSoutput.n160 CSoutput.n140 0.001
R14906 CSoutput.n191 CSoutput.n140 0.001
R14907 CSoutput.n161 CSoutput.n141 0.001
R14908 CSoutput.n192 CSoutput.n141 0.001
R14909 CSoutput.n192 CSoutput.n142 0.001
R14910 CSoutput.n191 CSoutput.n143 0.001
R14911 CSoutput.n190 CSoutput.n144 0.001
R14912 CSoutput.n189 CSoutput.t140 0.001
R14913 CSoutput.n188 CSoutput.n145 0.001
R14914 CSoutput.n161 CSoutput.n143 0.001
R14915 CSoutput.n160 CSoutput.n144 0.001
R14916 CSoutput.n159 CSoutput.t140 0.001
R14917 CSoutput.n158 CSoutput.n145 0.001
R14918 CSoutput.n234 CSoutput.n146 0.001
R14919 CSoutput.n199 CSoutput.n177 0.001
R14920 CSoutput.n198 CSoutput.n178 0.001
R14921 CSoutput.n197 CSoutput.n179 0.001
R14922 CSoutput.n196 CSoutput.t132 0.001
R14923 CSoutput.n218 CSoutput.n180 0.001
R14924 CSoutput.n205 CSoutput.n178 0.001
R14925 CSoutput.n204 CSoutput.n179 0.001
R14926 CSoutput.n203 CSoutput.t132 0.001
R14927 CSoutput.n202 CSoutput.n180 0.001
R14928 CSoutput.n229 CSoutput.n172 0.001
R14929 CSoutput.n226 CSoutput.n108 0.001
R14930 CSoutput.n225 CSoutput.n109 0.001
R14931 CSoutput.n224 CSoutput.n110 0.001
R14932 CSoutput.n223 CSoutput.t131 0.001
R14933 CSoutput.n222 CSoutput.n111 0.001
R14934 CSoutput.n127 CSoutput.n109 0.001
R14935 CSoutput.n126 CSoutput.n110 0.001
R14936 CSoutput.n125 CSoutput.t131 0.001
R14937 CSoutput.n124 CSoutput.n111 0.001
R14938 CSoutput.n244 CSoutput.n112 0.001
R14939 vdd.n291 vdd.n255 756.745
R14940 vdd.n244 vdd.n208 756.745
R14941 vdd.n201 vdd.n165 756.745
R14942 vdd.n154 vdd.n118 756.745
R14943 vdd.n112 vdd.n76 756.745
R14944 vdd.n65 vdd.n29 756.745
R14945 vdd.n1106 vdd.n1070 756.745
R14946 vdd.n1153 vdd.n1117 756.745
R14947 vdd.n1016 vdd.n980 756.745
R14948 vdd.n1063 vdd.n1027 756.745
R14949 vdd.n927 vdd.n891 756.745
R14950 vdd.n974 vdd.n938 756.745
R14951 vdd.n1791 vdd.t88 640.208
R14952 vdd.n755 vdd.t73 640.208
R14953 vdd.n1765 vdd.t114 640.208
R14954 vdd.n747 vdd.t105 640.208
R14955 vdd.n2536 vdd.t56 640.208
R14956 vdd.n2256 vdd.t96 640.208
R14957 vdd.n622 vdd.t77 640.208
R14958 vdd.n2253 vdd.t81 640.208
R14959 vdd.n589 vdd.t85 640.208
R14960 vdd.n817 vdd.t92 640.208
R14961 vdd.n1320 vdd.t52 592.009
R14962 vdd.n1358 vdd.t99 592.009
R14963 vdd.n1254 vdd.t102 592.009
R14964 vdd.n1947 vdd.t48 592.009
R14965 vdd.n1584 vdd.t60 592.009
R14966 vdd.n1544 vdd.t67 592.009
R14967 vdd.n2908 vdd.t111 592.009
R14968 vdd.n405 vdd.t63 592.009
R14969 vdd.n365 vdd.t70 592.009
R14970 vdd.n557 vdd.t41 592.009
R14971 vdd.n2804 vdd.t45 592.009
R14972 vdd.n2711 vdd.t108 592.009
R14973 vdd.n292 vdd.n291 585
R14974 vdd.n290 vdd.n257 585
R14975 vdd.n289 vdd.n288 585
R14976 vdd.n260 vdd.n258 585
R14977 vdd.n283 vdd.n282 585
R14978 vdd.n281 vdd.n280 585
R14979 vdd.n264 vdd.n263 585
R14980 vdd.n275 vdd.n274 585
R14981 vdd.n273 vdd.n272 585
R14982 vdd.n268 vdd.n267 585
R14983 vdd.n245 vdd.n244 585
R14984 vdd.n243 vdd.n210 585
R14985 vdd.n242 vdd.n241 585
R14986 vdd.n213 vdd.n211 585
R14987 vdd.n236 vdd.n235 585
R14988 vdd.n234 vdd.n233 585
R14989 vdd.n217 vdd.n216 585
R14990 vdd.n228 vdd.n227 585
R14991 vdd.n226 vdd.n225 585
R14992 vdd.n221 vdd.n220 585
R14993 vdd.n202 vdd.n201 585
R14994 vdd.n200 vdd.n167 585
R14995 vdd.n199 vdd.n198 585
R14996 vdd.n170 vdd.n168 585
R14997 vdd.n193 vdd.n192 585
R14998 vdd.n191 vdd.n190 585
R14999 vdd.n174 vdd.n173 585
R15000 vdd.n185 vdd.n184 585
R15001 vdd.n183 vdd.n182 585
R15002 vdd.n178 vdd.n177 585
R15003 vdd.n155 vdd.n154 585
R15004 vdd.n153 vdd.n120 585
R15005 vdd.n152 vdd.n151 585
R15006 vdd.n123 vdd.n121 585
R15007 vdd.n146 vdd.n145 585
R15008 vdd.n144 vdd.n143 585
R15009 vdd.n127 vdd.n126 585
R15010 vdd.n138 vdd.n137 585
R15011 vdd.n136 vdd.n135 585
R15012 vdd.n131 vdd.n130 585
R15013 vdd.n113 vdd.n112 585
R15014 vdd.n111 vdd.n78 585
R15015 vdd.n110 vdd.n109 585
R15016 vdd.n81 vdd.n79 585
R15017 vdd.n104 vdd.n103 585
R15018 vdd.n102 vdd.n101 585
R15019 vdd.n85 vdd.n84 585
R15020 vdd.n96 vdd.n95 585
R15021 vdd.n94 vdd.n93 585
R15022 vdd.n89 vdd.n88 585
R15023 vdd.n66 vdd.n65 585
R15024 vdd.n64 vdd.n31 585
R15025 vdd.n63 vdd.n62 585
R15026 vdd.n34 vdd.n32 585
R15027 vdd.n57 vdd.n56 585
R15028 vdd.n55 vdd.n54 585
R15029 vdd.n38 vdd.n37 585
R15030 vdd.n49 vdd.n48 585
R15031 vdd.n47 vdd.n46 585
R15032 vdd.n42 vdd.n41 585
R15033 vdd.n1107 vdd.n1106 585
R15034 vdd.n1105 vdd.n1072 585
R15035 vdd.n1104 vdd.n1103 585
R15036 vdd.n1075 vdd.n1073 585
R15037 vdd.n1098 vdd.n1097 585
R15038 vdd.n1096 vdd.n1095 585
R15039 vdd.n1079 vdd.n1078 585
R15040 vdd.n1090 vdd.n1089 585
R15041 vdd.n1088 vdd.n1087 585
R15042 vdd.n1083 vdd.n1082 585
R15043 vdd.n1154 vdd.n1153 585
R15044 vdd.n1152 vdd.n1119 585
R15045 vdd.n1151 vdd.n1150 585
R15046 vdd.n1122 vdd.n1120 585
R15047 vdd.n1145 vdd.n1144 585
R15048 vdd.n1143 vdd.n1142 585
R15049 vdd.n1126 vdd.n1125 585
R15050 vdd.n1137 vdd.n1136 585
R15051 vdd.n1135 vdd.n1134 585
R15052 vdd.n1130 vdd.n1129 585
R15053 vdd.n1017 vdd.n1016 585
R15054 vdd.n1015 vdd.n982 585
R15055 vdd.n1014 vdd.n1013 585
R15056 vdd.n985 vdd.n983 585
R15057 vdd.n1008 vdd.n1007 585
R15058 vdd.n1006 vdd.n1005 585
R15059 vdd.n989 vdd.n988 585
R15060 vdd.n1000 vdd.n999 585
R15061 vdd.n998 vdd.n997 585
R15062 vdd.n993 vdd.n992 585
R15063 vdd.n1064 vdd.n1063 585
R15064 vdd.n1062 vdd.n1029 585
R15065 vdd.n1061 vdd.n1060 585
R15066 vdd.n1032 vdd.n1030 585
R15067 vdd.n1055 vdd.n1054 585
R15068 vdd.n1053 vdd.n1052 585
R15069 vdd.n1036 vdd.n1035 585
R15070 vdd.n1047 vdd.n1046 585
R15071 vdd.n1045 vdd.n1044 585
R15072 vdd.n1040 vdd.n1039 585
R15073 vdd.n928 vdd.n927 585
R15074 vdd.n926 vdd.n893 585
R15075 vdd.n925 vdd.n924 585
R15076 vdd.n896 vdd.n894 585
R15077 vdd.n919 vdd.n918 585
R15078 vdd.n917 vdd.n916 585
R15079 vdd.n900 vdd.n899 585
R15080 vdd.n911 vdd.n910 585
R15081 vdd.n909 vdd.n908 585
R15082 vdd.n904 vdd.n903 585
R15083 vdd.n975 vdd.n974 585
R15084 vdd.n973 vdd.n940 585
R15085 vdd.n972 vdd.n971 585
R15086 vdd.n943 vdd.n941 585
R15087 vdd.n966 vdd.n965 585
R15088 vdd.n964 vdd.n963 585
R15089 vdd.n947 vdd.n946 585
R15090 vdd.n958 vdd.n957 585
R15091 vdd.n956 vdd.n955 585
R15092 vdd.n951 vdd.n950 585
R15093 vdd.n3024 vdd.n330 515.122
R15094 vdd.n2906 vdd.n328 515.122
R15095 vdd.n515 vdd.n478 515.122
R15096 vdd.n2842 vdd.n479 515.122
R15097 vdd.n1942 vdd.n865 515.122
R15098 vdd.n1945 vdd.n1944 515.122
R15099 vdd.n1227 vdd.n1191 515.122
R15100 vdd.n1423 vdd.n1192 515.122
R15101 vdd.n269 vdd.t141 329.043
R15102 vdd.n222 vdd.t152 329.043
R15103 vdd.n179 vdd.t137 329.043
R15104 vdd.n132 vdd.t147 329.043
R15105 vdd.n90 vdd.t178 329.043
R15106 vdd.n43 vdd.t120 329.043
R15107 vdd.n1084 vdd.t176 329.043
R15108 vdd.n1131 vdd.t162 329.043
R15109 vdd.n994 vdd.t168 329.043
R15110 vdd.n1041 vdd.t155 329.043
R15111 vdd.n905 vdd.t118 329.043
R15112 vdd.n952 vdd.t177 329.043
R15113 vdd.n1320 vdd.t55 319.788
R15114 vdd.n1358 vdd.t101 319.788
R15115 vdd.n1254 vdd.t104 319.788
R15116 vdd.n1947 vdd.t50 319.788
R15117 vdd.n1584 vdd.t61 319.788
R15118 vdd.n1544 vdd.t68 319.788
R15119 vdd.n2908 vdd.t112 319.788
R15120 vdd.n405 vdd.t65 319.788
R15121 vdd.n365 vdd.t71 319.788
R15122 vdd.n557 vdd.t44 319.788
R15123 vdd.n2804 vdd.t47 319.788
R15124 vdd.n2711 vdd.t110 319.788
R15125 vdd.n1321 vdd.t54 303.69
R15126 vdd.n1359 vdd.t100 303.69
R15127 vdd.n1255 vdd.t103 303.69
R15128 vdd.n1948 vdd.t51 303.69
R15129 vdd.n1585 vdd.t62 303.69
R15130 vdd.n1545 vdd.t69 303.69
R15131 vdd.n2909 vdd.t113 303.69
R15132 vdd.n406 vdd.t66 303.69
R15133 vdd.n366 vdd.t72 303.69
R15134 vdd.n558 vdd.t43 303.69
R15135 vdd.n2805 vdd.t46 303.69
R15136 vdd.n2712 vdd.t109 303.69
R15137 vdd.n2479 vdd.n703 297.074
R15138 vdd.n2672 vdd.n599 297.074
R15139 vdd.n2609 vdd.n596 297.074
R15140 vdd.n2402 vdd.n704 297.074
R15141 vdd.n2217 vdd.n744 297.074
R15142 vdd.n2148 vdd.n2147 297.074
R15143 vdd.n1894 vdd.n840 297.074
R15144 vdd.n1990 vdd.n838 297.074
R15145 vdd.n2588 vdd.n597 297.074
R15146 vdd.n2675 vdd.n2674 297.074
R15147 vdd.n2251 vdd.n705 297.074
R15148 vdd.n2477 vdd.n706 297.074
R15149 vdd.n2145 vdd.n753 297.074
R15150 vdd.n751 vdd.n726 297.074
R15151 vdd.n1831 vdd.n841 297.074
R15152 vdd.n1988 vdd.n842 297.074
R15153 vdd.n2590 vdd.n597 185
R15154 vdd.n2673 vdd.n597 185
R15155 vdd.n2592 vdd.n2591 185
R15156 vdd.n2591 vdd.n595 185
R15157 vdd.n2593 vdd.n629 185
R15158 vdd.n2603 vdd.n629 185
R15159 vdd.n2594 vdd.n638 185
R15160 vdd.n638 vdd.n636 185
R15161 vdd.n2596 vdd.n2595 185
R15162 vdd.n2597 vdd.n2596 185
R15163 vdd.n2549 vdd.n637 185
R15164 vdd.n637 vdd.n633 185
R15165 vdd.n2548 vdd.n2547 185
R15166 vdd.n2547 vdd.n2546 185
R15167 vdd.n640 vdd.n639 185
R15168 vdd.n641 vdd.n640 185
R15169 vdd.n2539 vdd.n2538 185
R15170 vdd.n2540 vdd.n2539 185
R15171 vdd.n2535 vdd.n650 185
R15172 vdd.n650 vdd.n647 185
R15173 vdd.n2534 vdd.n2533 185
R15174 vdd.n2533 vdd.n2532 185
R15175 vdd.n652 vdd.n651 185
R15176 vdd.n660 vdd.n652 185
R15177 vdd.n2525 vdd.n2524 185
R15178 vdd.n2526 vdd.n2525 185
R15179 vdd.n2523 vdd.n661 185
R15180 vdd.n2374 vdd.n661 185
R15181 vdd.n2522 vdd.n2521 185
R15182 vdd.n2521 vdd.n2520 185
R15183 vdd.n663 vdd.n662 185
R15184 vdd.n664 vdd.n663 185
R15185 vdd.n2513 vdd.n2512 185
R15186 vdd.n2514 vdd.n2513 185
R15187 vdd.n2511 vdd.n673 185
R15188 vdd.n673 vdd.n670 185
R15189 vdd.n2510 vdd.n2509 185
R15190 vdd.n2509 vdd.n2508 185
R15191 vdd.n675 vdd.n674 185
R15192 vdd.n683 vdd.n675 185
R15193 vdd.n2501 vdd.n2500 185
R15194 vdd.n2502 vdd.n2501 185
R15195 vdd.n2499 vdd.n684 185
R15196 vdd.n690 vdd.n684 185
R15197 vdd.n2498 vdd.n2497 185
R15198 vdd.n2497 vdd.n2496 185
R15199 vdd.n686 vdd.n685 185
R15200 vdd.n687 vdd.n686 185
R15201 vdd.n2489 vdd.n2488 185
R15202 vdd.n2490 vdd.n2489 185
R15203 vdd.n2487 vdd.n696 185
R15204 vdd.n2395 vdd.n696 185
R15205 vdd.n2486 vdd.n2485 185
R15206 vdd.n2485 vdd.n2484 185
R15207 vdd.n698 vdd.n697 185
R15208 vdd.t190 vdd.n698 185
R15209 vdd.n2477 vdd.n2476 185
R15210 vdd.n2478 vdd.n2477 185
R15211 vdd.n2475 vdd.n706 185
R15212 vdd.n2474 vdd.n2473 185
R15213 vdd.n708 vdd.n707 185
R15214 vdd.n2260 vdd.n2259 185
R15215 vdd.n2262 vdd.n2261 185
R15216 vdd.n2264 vdd.n2263 185
R15217 vdd.n2266 vdd.n2265 185
R15218 vdd.n2268 vdd.n2267 185
R15219 vdd.n2270 vdd.n2269 185
R15220 vdd.n2272 vdd.n2271 185
R15221 vdd.n2274 vdd.n2273 185
R15222 vdd.n2276 vdd.n2275 185
R15223 vdd.n2278 vdd.n2277 185
R15224 vdd.n2280 vdd.n2279 185
R15225 vdd.n2282 vdd.n2281 185
R15226 vdd.n2284 vdd.n2283 185
R15227 vdd.n2286 vdd.n2285 185
R15228 vdd.n2288 vdd.n2287 185
R15229 vdd.n2290 vdd.n2289 185
R15230 vdd.n2292 vdd.n2291 185
R15231 vdd.n2294 vdd.n2293 185
R15232 vdd.n2296 vdd.n2295 185
R15233 vdd.n2298 vdd.n2297 185
R15234 vdd.n2300 vdd.n2299 185
R15235 vdd.n2302 vdd.n2301 185
R15236 vdd.n2304 vdd.n2303 185
R15237 vdd.n2306 vdd.n2305 185
R15238 vdd.n2308 vdd.n2307 185
R15239 vdd.n2310 vdd.n2309 185
R15240 vdd.n2312 vdd.n2311 185
R15241 vdd.n2314 vdd.n2313 185
R15242 vdd.n2316 vdd.n2315 185
R15243 vdd.n2318 vdd.n2317 185
R15244 vdd.n2320 vdd.n2319 185
R15245 vdd.n2321 vdd.n2251 185
R15246 vdd.n2471 vdd.n2251 185
R15247 vdd.n2676 vdd.n2675 185
R15248 vdd.n2677 vdd.n588 185
R15249 vdd.n2679 vdd.n2678 185
R15250 vdd.n2681 vdd.n586 185
R15251 vdd.n2683 vdd.n2682 185
R15252 vdd.n2684 vdd.n585 185
R15253 vdd.n2686 vdd.n2685 185
R15254 vdd.n2688 vdd.n583 185
R15255 vdd.n2690 vdd.n2689 185
R15256 vdd.n2691 vdd.n582 185
R15257 vdd.n2693 vdd.n2692 185
R15258 vdd.n2695 vdd.n580 185
R15259 vdd.n2697 vdd.n2696 185
R15260 vdd.n2698 vdd.n579 185
R15261 vdd.n2700 vdd.n2699 185
R15262 vdd.n2702 vdd.n578 185
R15263 vdd.n2703 vdd.n576 185
R15264 vdd.n2706 vdd.n2705 185
R15265 vdd.n577 vdd.n575 185
R15266 vdd.n2562 vdd.n2561 185
R15267 vdd.n2564 vdd.n2563 185
R15268 vdd.n2566 vdd.n2558 185
R15269 vdd.n2568 vdd.n2567 185
R15270 vdd.n2569 vdd.n2557 185
R15271 vdd.n2571 vdd.n2570 185
R15272 vdd.n2573 vdd.n2555 185
R15273 vdd.n2575 vdd.n2574 185
R15274 vdd.n2576 vdd.n2554 185
R15275 vdd.n2578 vdd.n2577 185
R15276 vdd.n2580 vdd.n2552 185
R15277 vdd.n2582 vdd.n2581 185
R15278 vdd.n2583 vdd.n2551 185
R15279 vdd.n2585 vdd.n2584 185
R15280 vdd.n2587 vdd.n2550 185
R15281 vdd.n2589 vdd.n2588 185
R15282 vdd.n2588 vdd.n484 185
R15283 vdd.n2674 vdd.n592 185
R15284 vdd.n2674 vdd.n2673 185
R15285 vdd.n2326 vdd.n594 185
R15286 vdd.n595 vdd.n594 185
R15287 vdd.n2327 vdd.n628 185
R15288 vdd.n2603 vdd.n628 185
R15289 vdd.n2329 vdd.n2328 185
R15290 vdd.n2328 vdd.n636 185
R15291 vdd.n2330 vdd.n635 185
R15292 vdd.n2597 vdd.n635 185
R15293 vdd.n2332 vdd.n2331 185
R15294 vdd.n2331 vdd.n633 185
R15295 vdd.n2333 vdd.n643 185
R15296 vdd.n2546 vdd.n643 185
R15297 vdd.n2335 vdd.n2334 185
R15298 vdd.n2334 vdd.n641 185
R15299 vdd.n2336 vdd.n649 185
R15300 vdd.n2540 vdd.n649 185
R15301 vdd.n2338 vdd.n2337 185
R15302 vdd.n2337 vdd.n647 185
R15303 vdd.n2339 vdd.n654 185
R15304 vdd.n2532 vdd.n654 185
R15305 vdd.n2341 vdd.n2340 185
R15306 vdd.n2340 vdd.n660 185
R15307 vdd.n2342 vdd.n659 185
R15308 vdd.n2526 vdd.n659 185
R15309 vdd.n2376 vdd.n2375 185
R15310 vdd.n2375 vdd.n2374 185
R15311 vdd.n2377 vdd.n666 185
R15312 vdd.n2520 vdd.n666 185
R15313 vdd.n2379 vdd.n2378 185
R15314 vdd.n2378 vdd.n664 185
R15315 vdd.n2380 vdd.n672 185
R15316 vdd.n2514 vdd.n672 185
R15317 vdd.n2382 vdd.n2381 185
R15318 vdd.n2381 vdd.n670 185
R15319 vdd.n2383 vdd.n677 185
R15320 vdd.n2508 vdd.n677 185
R15321 vdd.n2385 vdd.n2384 185
R15322 vdd.n2384 vdd.n683 185
R15323 vdd.n2386 vdd.n682 185
R15324 vdd.n2502 vdd.n682 185
R15325 vdd.n2388 vdd.n2387 185
R15326 vdd.n2387 vdd.n690 185
R15327 vdd.n2389 vdd.n689 185
R15328 vdd.n2496 vdd.n689 185
R15329 vdd.n2391 vdd.n2390 185
R15330 vdd.n2390 vdd.n687 185
R15331 vdd.n2392 vdd.n695 185
R15332 vdd.n2490 vdd.n695 185
R15333 vdd.n2394 vdd.n2393 185
R15334 vdd.n2395 vdd.n2394 185
R15335 vdd.n2325 vdd.n700 185
R15336 vdd.n2484 vdd.n700 185
R15337 vdd.n2324 vdd.n2323 185
R15338 vdd.n2323 vdd.t190 185
R15339 vdd.n2322 vdd.n705 185
R15340 vdd.n2478 vdd.n705 185
R15341 vdd.n1942 vdd.n1941 185
R15342 vdd.n1943 vdd.n1942 185
R15343 vdd.n866 vdd.n864 185
R15344 vdd.n1508 vdd.n864 185
R15345 vdd.n1511 vdd.n1510 185
R15346 vdd.n1510 vdd.n1509 185
R15347 vdd.n869 vdd.n868 185
R15348 vdd.n870 vdd.n869 185
R15349 vdd.n1497 vdd.n1496 185
R15350 vdd.n1498 vdd.n1497 185
R15351 vdd.n878 vdd.n877 185
R15352 vdd.n1489 vdd.n877 185
R15353 vdd.n1492 vdd.n1491 185
R15354 vdd.n1491 vdd.n1490 185
R15355 vdd.n881 vdd.n880 185
R15356 vdd.n888 vdd.n881 185
R15357 vdd.n1480 vdd.n1479 185
R15358 vdd.n1481 vdd.n1480 185
R15359 vdd.n890 vdd.n889 185
R15360 vdd.n889 vdd.n887 185
R15361 vdd.n1475 vdd.n1474 185
R15362 vdd.n1474 vdd.n1473 185
R15363 vdd.n1163 vdd.n1162 185
R15364 vdd.n1164 vdd.n1163 185
R15365 vdd.n1464 vdd.n1463 185
R15366 vdd.n1465 vdd.n1464 185
R15367 vdd.n1171 vdd.n1170 185
R15368 vdd.n1455 vdd.n1170 185
R15369 vdd.n1458 vdd.n1457 185
R15370 vdd.n1457 vdd.n1456 185
R15371 vdd.n1174 vdd.n1173 185
R15372 vdd.n1180 vdd.n1174 185
R15373 vdd.n1446 vdd.n1445 185
R15374 vdd.n1447 vdd.n1446 185
R15375 vdd.n1182 vdd.n1181 185
R15376 vdd.n1438 vdd.n1181 185
R15377 vdd.n1441 vdd.n1440 185
R15378 vdd.n1440 vdd.n1439 185
R15379 vdd.n1185 vdd.n1184 185
R15380 vdd.n1186 vdd.n1185 185
R15381 vdd.n1429 vdd.n1428 185
R15382 vdd.n1430 vdd.n1429 185
R15383 vdd.n1193 vdd.n1192 185
R15384 vdd.n1228 vdd.n1192 185
R15385 vdd.n1424 vdd.n1423 185
R15386 vdd.n1196 vdd.n1195 185
R15387 vdd.n1420 vdd.n1419 185
R15388 vdd.n1421 vdd.n1420 185
R15389 vdd.n1230 vdd.n1229 185
R15390 vdd.n1415 vdd.n1232 185
R15391 vdd.n1414 vdd.n1233 185
R15392 vdd.n1413 vdd.n1234 185
R15393 vdd.n1236 vdd.n1235 185
R15394 vdd.n1409 vdd.n1238 185
R15395 vdd.n1408 vdd.n1239 185
R15396 vdd.n1407 vdd.n1240 185
R15397 vdd.n1242 vdd.n1241 185
R15398 vdd.n1403 vdd.n1244 185
R15399 vdd.n1402 vdd.n1245 185
R15400 vdd.n1401 vdd.n1246 185
R15401 vdd.n1248 vdd.n1247 185
R15402 vdd.n1397 vdd.n1250 185
R15403 vdd.n1396 vdd.n1251 185
R15404 vdd.n1395 vdd.n1252 185
R15405 vdd.n1256 vdd.n1253 185
R15406 vdd.n1391 vdd.n1258 185
R15407 vdd.n1390 vdd.n1259 185
R15408 vdd.n1389 vdd.n1260 185
R15409 vdd.n1262 vdd.n1261 185
R15410 vdd.n1385 vdd.n1264 185
R15411 vdd.n1384 vdd.n1265 185
R15412 vdd.n1383 vdd.n1266 185
R15413 vdd.n1268 vdd.n1267 185
R15414 vdd.n1379 vdd.n1270 185
R15415 vdd.n1378 vdd.n1271 185
R15416 vdd.n1377 vdd.n1272 185
R15417 vdd.n1274 vdd.n1273 185
R15418 vdd.n1373 vdd.n1276 185
R15419 vdd.n1372 vdd.n1277 185
R15420 vdd.n1371 vdd.n1278 185
R15421 vdd.n1280 vdd.n1279 185
R15422 vdd.n1367 vdd.n1282 185
R15423 vdd.n1366 vdd.n1283 185
R15424 vdd.n1365 vdd.n1284 185
R15425 vdd.n1286 vdd.n1285 185
R15426 vdd.n1361 vdd.n1288 185
R15427 vdd.n1360 vdd.n1357 185
R15428 vdd.n1356 vdd.n1289 185
R15429 vdd.n1291 vdd.n1290 185
R15430 vdd.n1352 vdd.n1293 185
R15431 vdd.n1351 vdd.n1294 185
R15432 vdd.n1350 vdd.n1295 185
R15433 vdd.n1297 vdd.n1296 185
R15434 vdd.n1346 vdd.n1299 185
R15435 vdd.n1345 vdd.n1300 185
R15436 vdd.n1344 vdd.n1301 185
R15437 vdd.n1303 vdd.n1302 185
R15438 vdd.n1340 vdd.n1305 185
R15439 vdd.n1339 vdd.n1306 185
R15440 vdd.n1338 vdd.n1307 185
R15441 vdd.n1309 vdd.n1308 185
R15442 vdd.n1334 vdd.n1311 185
R15443 vdd.n1333 vdd.n1312 185
R15444 vdd.n1332 vdd.n1313 185
R15445 vdd.n1315 vdd.n1314 185
R15446 vdd.n1328 vdd.n1317 185
R15447 vdd.n1327 vdd.n1318 185
R15448 vdd.n1326 vdd.n1319 185
R15449 vdd.n1323 vdd.n1227 185
R15450 vdd.n1421 vdd.n1227 185
R15451 vdd.n1946 vdd.n1945 185
R15452 vdd.n1950 vdd.n859 185
R15453 vdd.n1613 vdd.n858 185
R15454 vdd.n1616 vdd.n1615 185
R15455 vdd.n1618 vdd.n1617 185
R15456 vdd.n1621 vdd.n1620 185
R15457 vdd.n1623 vdd.n1622 185
R15458 vdd.n1625 vdd.n1611 185
R15459 vdd.n1627 vdd.n1626 185
R15460 vdd.n1628 vdd.n1605 185
R15461 vdd.n1630 vdd.n1629 185
R15462 vdd.n1632 vdd.n1603 185
R15463 vdd.n1634 vdd.n1633 185
R15464 vdd.n1635 vdd.n1598 185
R15465 vdd.n1637 vdd.n1636 185
R15466 vdd.n1639 vdd.n1596 185
R15467 vdd.n1641 vdd.n1640 185
R15468 vdd.n1642 vdd.n1592 185
R15469 vdd.n1644 vdd.n1643 185
R15470 vdd.n1646 vdd.n1589 185
R15471 vdd.n1648 vdd.n1647 185
R15472 vdd.n1590 vdd.n1583 185
R15473 vdd.n1652 vdd.n1587 185
R15474 vdd.n1653 vdd.n1579 185
R15475 vdd.n1655 vdd.n1654 185
R15476 vdd.n1657 vdd.n1577 185
R15477 vdd.n1659 vdd.n1658 185
R15478 vdd.n1660 vdd.n1572 185
R15479 vdd.n1662 vdd.n1661 185
R15480 vdd.n1664 vdd.n1570 185
R15481 vdd.n1666 vdd.n1665 185
R15482 vdd.n1667 vdd.n1565 185
R15483 vdd.n1669 vdd.n1668 185
R15484 vdd.n1671 vdd.n1563 185
R15485 vdd.n1673 vdd.n1672 185
R15486 vdd.n1674 vdd.n1558 185
R15487 vdd.n1676 vdd.n1675 185
R15488 vdd.n1678 vdd.n1556 185
R15489 vdd.n1680 vdd.n1679 185
R15490 vdd.n1681 vdd.n1552 185
R15491 vdd.n1683 vdd.n1682 185
R15492 vdd.n1685 vdd.n1549 185
R15493 vdd.n1687 vdd.n1686 185
R15494 vdd.n1550 vdd.n1543 185
R15495 vdd.n1691 vdd.n1547 185
R15496 vdd.n1692 vdd.n1539 185
R15497 vdd.n1694 vdd.n1693 185
R15498 vdd.n1696 vdd.n1537 185
R15499 vdd.n1698 vdd.n1697 185
R15500 vdd.n1699 vdd.n1532 185
R15501 vdd.n1701 vdd.n1700 185
R15502 vdd.n1703 vdd.n1530 185
R15503 vdd.n1705 vdd.n1704 185
R15504 vdd.n1706 vdd.n1525 185
R15505 vdd.n1708 vdd.n1707 185
R15506 vdd.n1710 vdd.n1524 185
R15507 vdd.n1711 vdd.n1521 185
R15508 vdd.n1714 vdd.n1713 185
R15509 vdd.n1523 vdd.n1519 185
R15510 vdd.n1931 vdd.n1517 185
R15511 vdd.n1933 vdd.n1932 185
R15512 vdd.n1935 vdd.n1515 185
R15513 vdd.n1937 vdd.n1936 185
R15514 vdd.n1938 vdd.n865 185
R15515 vdd.n1944 vdd.n862 185
R15516 vdd.n1944 vdd.n1943 185
R15517 vdd.n873 vdd.n861 185
R15518 vdd.n1508 vdd.n861 185
R15519 vdd.n1507 vdd.n1506 185
R15520 vdd.n1509 vdd.n1507 185
R15521 vdd.n872 vdd.n871 185
R15522 vdd.n871 vdd.n870 185
R15523 vdd.n1500 vdd.n1499 185
R15524 vdd.n1499 vdd.n1498 185
R15525 vdd.n876 vdd.n875 185
R15526 vdd.n1489 vdd.n876 185
R15527 vdd.n1488 vdd.n1487 185
R15528 vdd.n1490 vdd.n1488 185
R15529 vdd.n883 vdd.n882 185
R15530 vdd.n888 vdd.n882 185
R15531 vdd.n1483 vdd.n1482 185
R15532 vdd.n1482 vdd.n1481 185
R15533 vdd.n886 vdd.n885 185
R15534 vdd.n887 vdd.n886 185
R15535 vdd.n1472 vdd.n1471 185
R15536 vdd.n1473 vdd.n1472 185
R15537 vdd.n1166 vdd.n1165 185
R15538 vdd.n1165 vdd.n1164 185
R15539 vdd.n1467 vdd.n1466 185
R15540 vdd.n1466 vdd.n1465 185
R15541 vdd.n1169 vdd.n1168 185
R15542 vdd.n1455 vdd.n1169 185
R15543 vdd.n1454 vdd.n1453 185
R15544 vdd.n1456 vdd.n1454 185
R15545 vdd.n1176 vdd.n1175 185
R15546 vdd.n1180 vdd.n1175 185
R15547 vdd.n1449 vdd.n1448 185
R15548 vdd.n1448 vdd.n1447 185
R15549 vdd.n1179 vdd.n1178 185
R15550 vdd.n1438 vdd.n1179 185
R15551 vdd.n1437 vdd.n1436 185
R15552 vdd.n1439 vdd.n1437 185
R15553 vdd.n1188 vdd.n1187 185
R15554 vdd.n1187 vdd.n1186 185
R15555 vdd.n1432 vdd.n1431 185
R15556 vdd.n1431 vdd.n1430 185
R15557 vdd.n1191 vdd.n1190 185
R15558 vdd.n1228 vdd.n1191 185
R15559 vdd.n746 vdd.n744 185
R15560 vdd.n2146 vdd.n744 185
R15561 vdd.n2068 vdd.n763 185
R15562 vdd.n763 vdd.t188 185
R15563 vdd.n2070 vdd.n2069 185
R15564 vdd.n2071 vdd.n2070 185
R15565 vdd.n2067 vdd.n762 185
R15566 vdd.n1770 vdd.n762 185
R15567 vdd.n2066 vdd.n2065 185
R15568 vdd.n2065 vdd.n2064 185
R15569 vdd.n765 vdd.n764 185
R15570 vdd.n766 vdd.n765 185
R15571 vdd.n2055 vdd.n2054 185
R15572 vdd.n2056 vdd.n2055 185
R15573 vdd.n2053 vdd.n776 185
R15574 vdd.n776 vdd.n773 185
R15575 vdd.n2052 vdd.n2051 185
R15576 vdd.n2051 vdd.n2050 185
R15577 vdd.n778 vdd.n777 185
R15578 vdd.n779 vdd.n778 185
R15579 vdd.n2043 vdd.n2042 185
R15580 vdd.n2044 vdd.n2043 185
R15581 vdd.n2041 vdd.n787 185
R15582 vdd.n792 vdd.n787 185
R15583 vdd.n2040 vdd.n2039 185
R15584 vdd.n2039 vdd.n2038 185
R15585 vdd.n789 vdd.n788 185
R15586 vdd.n798 vdd.n789 185
R15587 vdd.n2031 vdd.n2030 185
R15588 vdd.n2032 vdd.n2031 185
R15589 vdd.n2029 vdd.n799 185
R15590 vdd.n1871 vdd.n799 185
R15591 vdd.n2028 vdd.n2027 185
R15592 vdd.n2027 vdd.n2026 185
R15593 vdd.n801 vdd.n800 185
R15594 vdd.n802 vdd.n801 185
R15595 vdd.n2019 vdd.n2018 185
R15596 vdd.n2020 vdd.n2019 185
R15597 vdd.n2017 vdd.n811 185
R15598 vdd.n811 vdd.n808 185
R15599 vdd.n2016 vdd.n2015 185
R15600 vdd.n2015 vdd.n2014 185
R15601 vdd.n813 vdd.n812 185
R15602 vdd.n823 vdd.n813 185
R15603 vdd.n2006 vdd.n2005 185
R15604 vdd.n2007 vdd.n2006 185
R15605 vdd.n2004 vdd.n824 185
R15606 vdd.n824 vdd.n820 185
R15607 vdd.n2003 vdd.n2002 185
R15608 vdd.n2002 vdd.n2001 185
R15609 vdd.n826 vdd.n825 185
R15610 vdd.n827 vdd.n826 185
R15611 vdd.n1994 vdd.n1993 185
R15612 vdd.n1995 vdd.n1994 185
R15613 vdd.n1992 vdd.n836 185
R15614 vdd.n836 vdd.n833 185
R15615 vdd.n1991 vdd.n1990 185
R15616 vdd.n1990 vdd.n1989 185
R15617 vdd.n838 vdd.n837 185
R15618 vdd.n1726 vdd.n1725 185
R15619 vdd.n1727 vdd.n1723 185
R15620 vdd.n1723 vdd.n839 185
R15621 vdd.n1729 vdd.n1728 185
R15622 vdd.n1731 vdd.n1722 185
R15623 vdd.n1734 vdd.n1733 185
R15624 vdd.n1735 vdd.n1721 185
R15625 vdd.n1737 vdd.n1736 185
R15626 vdd.n1739 vdd.n1720 185
R15627 vdd.n1742 vdd.n1741 185
R15628 vdd.n1743 vdd.n1719 185
R15629 vdd.n1745 vdd.n1744 185
R15630 vdd.n1747 vdd.n1718 185
R15631 vdd.n1750 vdd.n1749 185
R15632 vdd.n1751 vdd.n1717 185
R15633 vdd.n1753 vdd.n1752 185
R15634 vdd.n1755 vdd.n1716 185
R15635 vdd.n1928 vdd.n1756 185
R15636 vdd.n1927 vdd.n1926 185
R15637 vdd.n1924 vdd.n1757 185
R15638 vdd.n1922 vdd.n1921 185
R15639 vdd.n1920 vdd.n1758 185
R15640 vdd.n1919 vdd.n1918 185
R15641 vdd.n1916 vdd.n1759 185
R15642 vdd.n1914 vdd.n1913 185
R15643 vdd.n1912 vdd.n1760 185
R15644 vdd.n1911 vdd.n1910 185
R15645 vdd.n1908 vdd.n1761 185
R15646 vdd.n1906 vdd.n1905 185
R15647 vdd.n1904 vdd.n1762 185
R15648 vdd.n1903 vdd.n1902 185
R15649 vdd.n1900 vdd.n1763 185
R15650 vdd.n1898 vdd.n1897 185
R15651 vdd.n1896 vdd.n1764 185
R15652 vdd.n1895 vdd.n1894 185
R15653 vdd.n2149 vdd.n2148 185
R15654 vdd.n2151 vdd.n2150 185
R15655 vdd.n2153 vdd.n2152 185
R15656 vdd.n2156 vdd.n2155 185
R15657 vdd.n2158 vdd.n2157 185
R15658 vdd.n2160 vdd.n2159 185
R15659 vdd.n2162 vdd.n2161 185
R15660 vdd.n2164 vdd.n2163 185
R15661 vdd.n2166 vdd.n2165 185
R15662 vdd.n2168 vdd.n2167 185
R15663 vdd.n2170 vdd.n2169 185
R15664 vdd.n2172 vdd.n2171 185
R15665 vdd.n2174 vdd.n2173 185
R15666 vdd.n2176 vdd.n2175 185
R15667 vdd.n2178 vdd.n2177 185
R15668 vdd.n2180 vdd.n2179 185
R15669 vdd.n2182 vdd.n2181 185
R15670 vdd.n2184 vdd.n2183 185
R15671 vdd.n2186 vdd.n2185 185
R15672 vdd.n2188 vdd.n2187 185
R15673 vdd.n2190 vdd.n2189 185
R15674 vdd.n2192 vdd.n2191 185
R15675 vdd.n2194 vdd.n2193 185
R15676 vdd.n2196 vdd.n2195 185
R15677 vdd.n2198 vdd.n2197 185
R15678 vdd.n2200 vdd.n2199 185
R15679 vdd.n2202 vdd.n2201 185
R15680 vdd.n2204 vdd.n2203 185
R15681 vdd.n2206 vdd.n2205 185
R15682 vdd.n2208 vdd.n2207 185
R15683 vdd.n2210 vdd.n2209 185
R15684 vdd.n2212 vdd.n2211 185
R15685 vdd.n2214 vdd.n2213 185
R15686 vdd.n2215 vdd.n745 185
R15687 vdd.n2217 vdd.n2216 185
R15688 vdd.n2218 vdd.n2217 185
R15689 vdd.n2147 vdd.n749 185
R15690 vdd.n2147 vdd.n2146 185
R15691 vdd.n1768 vdd.n750 185
R15692 vdd.t188 vdd.n750 185
R15693 vdd.n1769 vdd.n760 185
R15694 vdd.n2071 vdd.n760 185
R15695 vdd.n1772 vdd.n1771 185
R15696 vdd.n1771 vdd.n1770 185
R15697 vdd.n1773 vdd.n767 185
R15698 vdd.n2064 vdd.n767 185
R15699 vdd.n1775 vdd.n1774 185
R15700 vdd.n1774 vdd.n766 185
R15701 vdd.n1776 vdd.n774 185
R15702 vdd.n2056 vdd.n774 185
R15703 vdd.n1778 vdd.n1777 185
R15704 vdd.n1777 vdd.n773 185
R15705 vdd.n1779 vdd.n780 185
R15706 vdd.n2050 vdd.n780 185
R15707 vdd.n1781 vdd.n1780 185
R15708 vdd.n1780 vdd.n779 185
R15709 vdd.n1782 vdd.n785 185
R15710 vdd.n2044 vdd.n785 185
R15711 vdd.n1784 vdd.n1783 185
R15712 vdd.n1783 vdd.n792 185
R15713 vdd.n1785 vdd.n790 185
R15714 vdd.n2038 vdd.n790 185
R15715 vdd.n1787 vdd.n1786 185
R15716 vdd.n1786 vdd.n798 185
R15717 vdd.n1788 vdd.n796 185
R15718 vdd.n2032 vdd.n796 185
R15719 vdd.n1873 vdd.n1872 185
R15720 vdd.n1872 vdd.n1871 185
R15721 vdd.n1874 vdd.n803 185
R15722 vdd.n2026 vdd.n803 185
R15723 vdd.n1876 vdd.n1875 185
R15724 vdd.n1875 vdd.n802 185
R15725 vdd.n1877 vdd.n809 185
R15726 vdd.n2020 vdd.n809 185
R15727 vdd.n1879 vdd.n1878 185
R15728 vdd.n1878 vdd.n808 185
R15729 vdd.n1880 vdd.n814 185
R15730 vdd.n2014 vdd.n814 185
R15731 vdd.n1882 vdd.n1881 185
R15732 vdd.n1881 vdd.n823 185
R15733 vdd.n1883 vdd.n821 185
R15734 vdd.n2007 vdd.n821 185
R15735 vdd.n1885 vdd.n1884 185
R15736 vdd.n1884 vdd.n820 185
R15737 vdd.n1886 vdd.n828 185
R15738 vdd.n2001 vdd.n828 185
R15739 vdd.n1888 vdd.n1887 185
R15740 vdd.n1887 vdd.n827 185
R15741 vdd.n1889 vdd.n834 185
R15742 vdd.n1995 vdd.n834 185
R15743 vdd.n1891 vdd.n1890 185
R15744 vdd.n1890 vdd.n833 185
R15745 vdd.n1892 vdd.n840 185
R15746 vdd.n1989 vdd.n840 185
R15747 vdd.n3024 vdd.n3023 185
R15748 vdd.n3025 vdd.n3024 185
R15749 vdd.n325 vdd.n324 185
R15750 vdd.n3026 vdd.n325 185
R15751 vdd.n3029 vdd.n3028 185
R15752 vdd.n3028 vdd.n3027 185
R15753 vdd.n3030 vdd.n319 185
R15754 vdd.n319 vdd.n318 185
R15755 vdd.n3032 vdd.n3031 185
R15756 vdd.n3033 vdd.n3032 185
R15757 vdd.n314 vdd.n313 185
R15758 vdd.n3034 vdd.n314 185
R15759 vdd.n3037 vdd.n3036 185
R15760 vdd.n3036 vdd.n3035 185
R15761 vdd.n3038 vdd.n309 185
R15762 vdd.n309 vdd.n308 185
R15763 vdd.n3040 vdd.n3039 185
R15764 vdd.n3041 vdd.n3040 185
R15765 vdd.n303 vdd.n301 185
R15766 vdd.n3042 vdd.n303 185
R15767 vdd.n3045 vdd.n3044 185
R15768 vdd.n3044 vdd.n3043 185
R15769 vdd.n302 vdd.n300 185
R15770 vdd.n304 vdd.n302 185
R15771 vdd.n2881 vdd.n2880 185
R15772 vdd.n2882 vdd.n2881 185
R15773 vdd.n458 vdd.n457 185
R15774 vdd.n457 vdd.n456 185
R15775 vdd.n2876 vdd.n2875 185
R15776 vdd.n2875 vdd.n2874 185
R15777 vdd.n461 vdd.n460 185
R15778 vdd.n467 vdd.n461 185
R15779 vdd.n2865 vdd.n2864 185
R15780 vdd.n2866 vdd.n2865 185
R15781 vdd.n469 vdd.n468 185
R15782 vdd.n2857 vdd.n468 185
R15783 vdd.n2860 vdd.n2859 185
R15784 vdd.n2859 vdd.n2858 185
R15785 vdd.n472 vdd.n471 185
R15786 vdd.n473 vdd.n472 185
R15787 vdd.n2848 vdd.n2847 185
R15788 vdd.n2849 vdd.n2848 185
R15789 vdd.n480 vdd.n479 185
R15790 vdd.n516 vdd.n479 185
R15791 vdd.n2843 vdd.n2842 185
R15792 vdd.n483 vdd.n482 185
R15793 vdd.n2839 vdd.n2838 185
R15794 vdd.n2840 vdd.n2839 185
R15795 vdd.n518 vdd.n517 185
R15796 vdd.n522 vdd.n521 185
R15797 vdd.n2834 vdd.n523 185
R15798 vdd.n2833 vdd.n2832 185
R15799 vdd.n2831 vdd.n2830 185
R15800 vdd.n2829 vdd.n2828 185
R15801 vdd.n2827 vdd.n2826 185
R15802 vdd.n2825 vdd.n2824 185
R15803 vdd.n2823 vdd.n2822 185
R15804 vdd.n2821 vdd.n2820 185
R15805 vdd.n2819 vdd.n2818 185
R15806 vdd.n2817 vdd.n2816 185
R15807 vdd.n2815 vdd.n2814 185
R15808 vdd.n2813 vdd.n2812 185
R15809 vdd.n2811 vdd.n2810 185
R15810 vdd.n2809 vdd.n2808 185
R15811 vdd.n2807 vdd.n2806 185
R15812 vdd.n2798 vdd.n536 185
R15813 vdd.n2800 vdd.n2799 185
R15814 vdd.n2797 vdd.n2796 185
R15815 vdd.n2795 vdd.n2794 185
R15816 vdd.n2793 vdd.n2792 185
R15817 vdd.n2791 vdd.n2790 185
R15818 vdd.n2789 vdd.n2788 185
R15819 vdd.n2787 vdd.n2786 185
R15820 vdd.n2785 vdd.n2784 185
R15821 vdd.n2783 vdd.n2782 185
R15822 vdd.n2781 vdd.n2780 185
R15823 vdd.n2779 vdd.n2778 185
R15824 vdd.n2777 vdd.n2776 185
R15825 vdd.n2775 vdd.n2774 185
R15826 vdd.n2773 vdd.n2772 185
R15827 vdd.n2771 vdd.n2770 185
R15828 vdd.n2769 vdd.n2768 185
R15829 vdd.n2767 vdd.n2766 185
R15830 vdd.n2765 vdd.n2764 185
R15831 vdd.n2763 vdd.n2762 185
R15832 vdd.n2761 vdd.n2760 185
R15833 vdd.n2759 vdd.n2758 185
R15834 vdd.n2752 vdd.n556 185
R15835 vdd.n2754 vdd.n2753 185
R15836 vdd.n2751 vdd.n2750 185
R15837 vdd.n2749 vdd.n2748 185
R15838 vdd.n2747 vdd.n2746 185
R15839 vdd.n2745 vdd.n2744 185
R15840 vdd.n2743 vdd.n2742 185
R15841 vdd.n2741 vdd.n2740 185
R15842 vdd.n2739 vdd.n2738 185
R15843 vdd.n2737 vdd.n2736 185
R15844 vdd.n2735 vdd.n2734 185
R15845 vdd.n2733 vdd.n2732 185
R15846 vdd.n2731 vdd.n2730 185
R15847 vdd.n2729 vdd.n2728 185
R15848 vdd.n2727 vdd.n2726 185
R15849 vdd.n2725 vdd.n2724 185
R15850 vdd.n2723 vdd.n2722 185
R15851 vdd.n2721 vdd.n2720 185
R15852 vdd.n2719 vdd.n2718 185
R15853 vdd.n2717 vdd.n2716 185
R15854 vdd.n2715 vdd.n2714 185
R15855 vdd.n2710 vdd.n515 185
R15856 vdd.n2840 vdd.n515 185
R15857 vdd.n2907 vdd.n2906 185
R15858 vdd.n2911 vdd.n440 185
R15859 vdd.n2913 vdd.n2912 185
R15860 vdd.n2915 vdd.n438 185
R15861 vdd.n2917 vdd.n2916 185
R15862 vdd.n2918 vdd.n433 185
R15863 vdd.n2920 vdd.n2919 185
R15864 vdd.n2922 vdd.n431 185
R15865 vdd.n2924 vdd.n2923 185
R15866 vdd.n2925 vdd.n426 185
R15867 vdd.n2927 vdd.n2926 185
R15868 vdd.n2929 vdd.n424 185
R15869 vdd.n2931 vdd.n2930 185
R15870 vdd.n2932 vdd.n419 185
R15871 vdd.n2934 vdd.n2933 185
R15872 vdd.n2936 vdd.n417 185
R15873 vdd.n2938 vdd.n2937 185
R15874 vdd.n2939 vdd.n413 185
R15875 vdd.n2941 vdd.n2940 185
R15876 vdd.n2943 vdd.n410 185
R15877 vdd.n2945 vdd.n2944 185
R15878 vdd.n411 vdd.n404 185
R15879 vdd.n2949 vdd.n408 185
R15880 vdd.n2950 vdd.n400 185
R15881 vdd.n2952 vdd.n2951 185
R15882 vdd.n2954 vdd.n398 185
R15883 vdd.n2956 vdd.n2955 185
R15884 vdd.n2957 vdd.n393 185
R15885 vdd.n2959 vdd.n2958 185
R15886 vdd.n2961 vdd.n391 185
R15887 vdd.n2963 vdd.n2962 185
R15888 vdd.n2964 vdd.n386 185
R15889 vdd.n2966 vdd.n2965 185
R15890 vdd.n2968 vdd.n384 185
R15891 vdd.n2970 vdd.n2969 185
R15892 vdd.n2971 vdd.n379 185
R15893 vdd.n2973 vdd.n2972 185
R15894 vdd.n2975 vdd.n377 185
R15895 vdd.n2977 vdd.n2976 185
R15896 vdd.n2978 vdd.n373 185
R15897 vdd.n2980 vdd.n2979 185
R15898 vdd.n2982 vdd.n370 185
R15899 vdd.n2984 vdd.n2983 185
R15900 vdd.n371 vdd.n364 185
R15901 vdd.n2988 vdd.n368 185
R15902 vdd.n2989 vdd.n360 185
R15903 vdd.n2991 vdd.n2990 185
R15904 vdd.n2993 vdd.n358 185
R15905 vdd.n2995 vdd.n2994 185
R15906 vdd.n2996 vdd.n353 185
R15907 vdd.n2998 vdd.n2997 185
R15908 vdd.n3000 vdd.n351 185
R15909 vdd.n3002 vdd.n3001 185
R15910 vdd.n3003 vdd.n346 185
R15911 vdd.n3005 vdd.n3004 185
R15912 vdd.n3007 vdd.n344 185
R15913 vdd.n3009 vdd.n3008 185
R15914 vdd.n3010 vdd.n338 185
R15915 vdd.n3012 vdd.n3011 185
R15916 vdd.n3014 vdd.n337 185
R15917 vdd.n3015 vdd.n336 185
R15918 vdd.n3018 vdd.n3017 185
R15919 vdd.n3019 vdd.n334 185
R15920 vdd.n3020 vdd.n330 185
R15921 vdd.n2902 vdd.n328 185
R15922 vdd.n3025 vdd.n328 185
R15923 vdd.n2901 vdd.n327 185
R15924 vdd.n3026 vdd.n327 185
R15925 vdd.n2900 vdd.n326 185
R15926 vdd.n3027 vdd.n326 185
R15927 vdd.n446 vdd.n445 185
R15928 vdd.n445 vdd.n318 185
R15929 vdd.n2896 vdd.n317 185
R15930 vdd.n3033 vdd.n317 185
R15931 vdd.n2895 vdd.n316 185
R15932 vdd.n3034 vdd.n316 185
R15933 vdd.n2894 vdd.n315 185
R15934 vdd.n3035 vdd.n315 185
R15935 vdd.n449 vdd.n448 185
R15936 vdd.n448 vdd.n308 185
R15937 vdd.n2890 vdd.n307 185
R15938 vdd.n3041 vdd.n307 185
R15939 vdd.n2889 vdd.n306 185
R15940 vdd.n3042 vdd.n306 185
R15941 vdd.n2888 vdd.n305 185
R15942 vdd.n3043 vdd.n305 185
R15943 vdd.n455 vdd.n451 185
R15944 vdd.n455 vdd.n304 185
R15945 vdd.n2884 vdd.n2883 185
R15946 vdd.n2883 vdd.n2882 185
R15947 vdd.n454 vdd.n453 185
R15948 vdd.n456 vdd.n454 185
R15949 vdd.n2873 vdd.n2872 185
R15950 vdd.n2874 vdd.n2873 185
R15951 vdd.n463 vdd.n462 185
R15952 vdd.n467 vdd.n462 185
R15953 vdd.n2868 vdd.n2867 185
R15954 vdd.n2867 vdd.n2866 185
R15955 vdd.n466 vdd.n465 185
R15956 vdd.n2857 vdd.n466 185
R15957 vdd.n2856 vdd.n2855 185
R15958 vdd.n2858 vdd.n2856 185
R15959 vdd.n475 vdd.n474 185
R15960 vdd.n474 vdd.n473 185
R15961 vdd.n2851 vdd.n2850 185
R15962 vdd.n2850 vdd.n2849 185
R15963 vdd.n478 vdd.n477 185
R15964 vdd.n516 vdd.n478 185
R15965 vdd.n703 vdd.n702 185
R15966 vdd.n2469 vdd.n2468 185
R15967 vdd.n2467 vdd.n2252 185
R15968 vdd.n2471 vdd.n2252 185
R15969 vdd.n2466 vdd.n2465 185
R15970 vdd.n2464 vdd.n2463 185
R15971 vdd.n2462 vdd.n2461 185
R15972 vdd.n2460 vdd.n2459 185
R15973 vdd.n2458 vdd.n2457 185
R15974 vdd.n2456 vdd.n2455 185
R15975 vdd.n2454 vdd.n2453 185
R15976 vdd.n2452 vdd.n2451 185
R15977 vdd.n2450 vdd.n2449 185
R15978 vdd.n2448 vdd.n2447 185
R15979 vdd.n2446 vdd.n2445 185
R15980 vdd.n2444 vdd.n2443 185
R15981 vdd.n2442 vdd.n2441 185
R15982 vdd.n2440 vdd.n2439 185
R15983 vdd.n2438 vdd.n2437 185
R15984 vdd.n2436 vdd.n2435 185
R15985 vdd.n2434 vdd.n2433 185
R15986 vdd.n2432 vdd.n2431 185
R15987 vdd.n2430 vdd.n2429 185
R15988 vdd.n2428 vdd.n2427 185
R15989 vdd.n2426 vdd.n2425 185
R15990 vdd.n2424 vdd.n2423 185
R15991 vdd.n2422 vdd.n2421 185
R15992 vdd.n2420 vdd.n2419 185
R15993 vdd.n2418 vdd.n2417 185
R15994 vdd.n2416 vdd.n2415 185
R15995 vdd.n2414 vdd.n2413 185
R15996 vdd.n2412 vdd.n2411 185
R15997 vdd.n2410 vdd.n2409 185
R15998 vdd.n2407 vdd.n2406 185
R15999 vdd.n2405 vdd.n2404 185
R16000 vdd.n2403 vdd.n2402 185
R16001 vdd.n2609 vdd.n2608 185
R16002 vdd.n2611 vdd.n624 185
R16003 vdd.n2613 vdd.n2612 185
R16004 vdd.n2615 vdd.n621 185
R16005 vdd.n2617 vdd.n2616 185
R16006 vdd.n2619 vdd.n619 185
R16007 vdd.n2621 vdd.n2620 185
R16008 vdd.n2622 vdd.n618 185
R16009 vdd.n2624 vdd.n2623 185
R16010 vdd.n2626 vdd.n616 185
R16011 vdd.n2628 vdd.n2627 185
R16012 vdd.n2629 vdd.n615 185
R16013 vdd.n2631 vdd.n2630 185
R16014 vdd.n2633 vdd.n613 185
R16015 vdd.n2635 vdd.n2634 185
R16016 vdd.n2636 vdd.n612 185
R16017 vdd.n2638 vdd.n2637 185
R16018 vdd.n2640 vdd.n520 185
R16019 vdd.n2642 vdd.n2641 185
R16020 vdd.n2644 vdd.n610 185
R16021 vdd.n2646 vdd.n2645 185
R16022 vdd.n2647 vdd.n609 185
R16023 vdd.n2649 vdd.n2648 185
R16024 vdd.n2651 vdd.n607 185
R16025 vdd.n2653 vdd.n2652 185
R16026 vdd.n2654 vdd.n606 185
R16027 vdd.n2656 vdd.n2655 185
R16028 vdd.n2658 vdd.n604 185
R16029 vdd.n2660 vdd.n2659 185
R16030 vdd.n2661 vdd.n603 185
R16031 vdd.n2663 vdd.n2662 185
R16032 vdd.n2665 vdd.n602 185
R16033 vdd.n2666 vdd.n601 185
R16034 vdd.n2669 vdd.n2668 185
R16035 vdd.n2670 vdd.n599 185
R16036 vdd.n599 vdd.n484 185
R16037 vdd.n2607 vdd.n596 185
R16038 vdd.n2673 vdd.n596 185
R16039 vdd.n2606 vdd.n2605 185
R16040 vdd.n2605 vdd.n595 185
R16041 vdd.n2604 vdd.n626 185
R16042 vdd.n2604 vdd.n2603 185
R16043 vdd.n2358 vdd.n627 185
R16044 vdd.n636 vdd.n627 185
R16045 vdd.n2359 vdd.n634 185
R16046 vdd.n2597 vdd.n634 185
R16047 vdd.n2361 vdd.n2360 185
R16048 vdd.n2360 vdd.n633 185
R16049 vdd.n2362 vdd.n642 185
R16050 vdd.n2546 vdd.n642 185
R16051 vdd.n2364 vdd.n2363 185
R16052 vdd.n2363 vdd.n641 185
R16053 vdd.n2365 vdd.n648 185
R16054 vdd.n2540 vdd.n648 185
R16055 vdd.n2367 vdd.n2366 185
R16056 vdd.n2366 vdd.n647 185
R16057 vdd.n2368 vdd.n653 185
R16058 vdd.n2532 vdd.n653 185
R16059 vdd.n2370 vdd.n2369 185
R16060 vdd.n2369 vdd.n660 185
R16061 vdd.n2371 vdd.n658 185
R16062 vdd.n2526 vdd.n658 185
R16063 vdd.n2373 vdd.n2372 185
R16064 vdd.n2374 vdd.n2373 185
R16065 vdd.n2357 vdd.n665 185
R16066 vdd.n2520 vdd.n665 185
R16067 vdd.n2356 vdd.n2355 185
R16068 vdd.n2355 vdd.n664 185
R16069 vdd.n2354 vdd.n671 185
R16070 vdd.n2514 vdd.n671 185
R16071 vdd.n2353 vdd.n2352 185
R16072 vdd.n2352 vdd.n670 185
R16073 vdd.n2351 vdd.n676 185
R16074 vdd.n2508 vdd.n676 185
R16075 vdd.n2350 vdd.n2349 185
R16076 vdd.n2349 vdd.n683 185
R16077 vdd.n2348 vdd.n681 185
R16078 vdd.n2502 vdd.n681 185
R16079 vdd.n2347 vdd.n2346 185
R16080 vdd.n2346 vdd.n690 185
R16081 vdd.n2345 vdd.n688 185
R16082 vdd.n2496 vdd.n688 185
R16083 vdd.n2344 vdd.n2343 185
R16084 vdd.n2343 vdd.n687 185
R16085 vdd.n2255 vdd.n694 185
R16086 vdd.n2490 vdd.n694 185
R16087 vdd.n2397 vdd.n2396 185
R16088 vdd.n2396 vdd.n2395 185
R16089 vdd.n2398 vdd.n699 185
R16090 vdd.n2484 vdd.n699 185
R16091 vdd.n2400 vdd.n2399 185
R16092 vdd.n2399 vdd.t190 185
R16093 vdd.n2401 vdd.n704 185
R16094 vdd.n2478 vdd.n704 185
R16095 vdd.n2480 vdd.n2479 185
R16096 vdd.n2479 vdd.n2478 185
R16097 vdd.n2481 vdd.n701 185
R16098 vdd.n701 vdd.t190 185
R16099 vdd.n2483 vdd.n2482 185
R16100 vdd.n2484 vdd.n2483 185
R16101 vdd.n693 vdd.n692 185
R16102 vdd.n2395 vdd.n693 185
R16103 vdd.n2492 vdd.n2491 185
R16104 vdd.n2491 vdd.n2490 185
R16105 vdd.n2493 vdd.n691 185
R16106 vdd.n691 vdd.n687 185
R16107 vdd.n2495 vdd.n2494 185
R16108 vdd.n2496 vdd.n2495 185
R16109 vdd.n680 vdd.n679 185
R16110 vdd.n690 vdd.n680 185
R16111 vdd.n2504 vdd.n2503 185
R16112 vdd.n2503 vdd.n2502 185
R16113 vdd.n2505 vdd.n678 185
R16114 vdd.n683 vdd.n678 185
R16115 vdd.n2507 vdd.n2506 185
R16116 vdd.n2508 vdd.n2507 185
R16117 vdd.n669 vdd.n668 185
R16118 vdd.n670 vdd.n669 185
R16119 vdd.n2516 vdd.n2515 185
R16120 vdd.n2515 vdd.n2514 185
R16121 vdd.n2517 vdd.n667 185
R16122 vdd.n667 vdd.n664 185
R16123 vdd.n2519 vdd.n2518 185
R16124 vdd.n2520 vdd.n2519 185
R16125 vdd.n657 vdd.n656 185
R16126 vdd.n2374 vdd.n657 185
R16127 vdd.n2528 vdd.n2527 185
R16128 vdd.n2527 vdd.n2526 185
R16129 vdd.n2529 vdd.n655 185
R16130 vdd.n660 vdd.n655 185
R16131 vdd.n2531 vdd.n2530 185
R16132 vdd.n2532 vdd.n2531 185
R16133 vdd.n646 vdd.n645 185
R16134 vdd.n647 vdd.n646 185
R16135 vdd.n2542 vdd.n2541 185
R16136 vdd.n2541 vdd.n2540 185
R16137 vdd.n2543 vdd.n644 185
R16138 vdd.n644 vdd.n641 185
R16139 vdd.n2545 vdd.n2544 185
R16140 vdd.n2546 vdd.n2545 185
R16141 vdd.n632 vdd.n631 185
R16142 vdd.n633 vdd.n632 185
R16143 vdd.n2599 vdd.n2598 185
R16144 vdd.n2598 vdd.n2597 185
R16145 vdd.n2600 vdd.n630 185
R16146 vdd.n636 vdd.n630 185
R16147 vdd.n2602 vdd.n2601 185
R16148 vdd.n2603 vdd.n2602 185
R16149 vdd.n600 vdd.n598 185
R16150 vdd.n598 vdd.n595 185
R16151 vdd.n2672 vdd.n2671 185
R16152 vdd.n2673 vdd.n2672 185
R16153 vdd.n2145 vdd.n2144 185
R16154 vdd.n2146 vdd.n2145 185
R16155 vdd.n754 vdd.n752 185
R16156 vdd.n752 vdd.t188 185
R16157 vdd.n2060 vdd.n761 185
R16158 vdd.n2071 vdd.n761 185
R16159 vdd.n2061 vdd.n770 185
R16160 vdd.n1770 vdd.n770 185
R16161 vdd.n2063 vdd.n2062 185
R16162 vdd.n2064 vdd.n2063 185
R16163 vdd.n2059 vdd.n769 185
R16164 vdd.n769 vdd.n766 185
R16165 vdd.n2058 vdd.n2057 185
R16166 vdd.n2057 vdd.n2056 185
R16167 vdd.n772 vdd.n771 185
R16168 vdd.n773 vdd.n772 185
R16169 vdd.n2049 vdd.n2048 185
R16170 vdd.n2050 vdd.n2049 185
R16171 vdd.n2047 vdd.n782 185
R16172 vdd.n782 vdd.n779 185
R16173 vdd.n2046 vdd.n2045 185
R16174 vdd.n2045 vdd.n2044 185
R16175 vdd.n784 vdd.n783 185
R16176 vdd.n792 vdd.n784 185
R16177 vdd.n2037 vdd.n2036 185
R16178 vdd.n2038 vdd.n2037 185
R16179 vdd.n2035 vdd.n793 185
R16180 vdd.n798 vdd.n793 185
R16181 vdd.n2034 vdd.n2033 185
R16182 vdd.n2033 vdd.n2032 185
R16183 vdd.n795 vdd.n794 185
R16184 vdd.n1871 vdd.n795 185
R16185 vdd.n2025 vdd.n2024 185
R16186 vdd.n2026 vdd.n2025 185
R16187 vdd.n2023 vdd.n805 185
R16188 vdd.n805 vdd.n802 185
R16189 vdd.n2022 vdd.n2021 185
R16190 vdd.n2021 vdd.n2020 185
R16191 vdd.n807 vdd.n806 185
R16192 vdd.n808 vdd.n807 185
R16193 vdd.n2013 vdd.n2012 185
R16194 vdd.n2014 vdd.n2013 185
R16195 vdd.n2010 vdd.n816 185
R16196 vdd.n823 vdd.n816 185
R16197 vdd.n2009 vdd.n2008 185
R16198 vdd.n2008 vdd.n2007 185
R16199 vdd.n819 vdd.n818 185
R16200 vdd.n820 vdd.n819 185
R16201 vdd.n2000 vdd.n1999 185
R16202 vdd.n2001 vdd.n2000 185
R16203 vdd.n1998 vdd.n830 185
R16204 vdd.n830 vdd.n827 185
R16205 vdd.n1997 vdd.n1996 185
R16206 vdd.n1996 vdd.n1995 185
R16207 vdd.n832 vdd.n831 185
R16208 vdd.n833 vdd.n832 185
R16209 vdd.n1988 vdd.n1987 185
R16210 vdd.n1989 vdd.n1988 185
R16211 vdd.n2076 vdd.n726 185
R16212 vdd.n2218 vdd.n726 185
R16213 vdd.n2078 vdd.n2077 185
R16214 vdd.n2080 vdd.n2079 185
R16215 vdd.n2082 vdd.n2081 185
R16216 vdd.n2084 vdd.n2083 185
R16217 vdd.n2086 vdd.n2085 185
R16218 vdd.n2088 vdd.n2087 185
R16219 vdd.n2090 vdd.n2089 185
R16220 vdd.n2092 vdd.n2091 185
R16221 vdd.n2094 vdd.n2093 185
R16222 vdd.n2096 vdd.n2095 185
R16223 vdd.n2098 vdd.n2097 185
R16224 vdd.n2100 vdd.n2099 185
R16225 vdd.n2102 vdd.n2101 185
R16226 vdd.n2104 vdd.n2103 185
R16227 vdd.n2106 vdd.n2105 185
R16228 vdd.n2108 vdd.n2107 185
R16229 vdd.n2110 vdd.n2109 185
R16230 vdd.n2112 vdd.n2111 185
R16231 vdd.n2114 vdd.n2113 185
R16232 vdd.n2116 vdd.n2115 185
R16233 vdd.n2118 vdd.n2117 185
R16234 vdd.n2120 vdd.n2119 185
R16235 vdd.n2122 vdd.n2121 185
R16236 vdd.n2124 vdd.n2123 185
R16237 vdd.n2126 vdd.n2125 185
R16238 vdd.n2128 vdd.n2127 185
R16239 vdd.n2130 vdd.n2129 185
R16240 vdd.n2132 vdd.n2131 185
R16241 vdd.n2134 vdd.n2133 185
R16242 vdd.n2136 vdd.n2135 185
R16243 vdd.n2138 vdd.n2137 185
R16244 vdd.n2140 vdd.n2139 185
R16245 vdd.n2142 vdd.n2141 185
R16246 vdd.n2143 vdd.n753 185
R16247 vdd.n2075 vdd.n751 185
R16248 vdd.n2146 vdd.n751 185
R16249 vdd.n2074 vdd.n2073 185
R16250 vdd.n2073 vdd.t188 185
R16251 vdd.n2072 vdd.n758 185
R16252 vdd.n2072 vdd.n2071 185
R16253 vdd.n1852 vdd.n759 185
R16254 vdd.n1770 vdd.n759 185
R16255 vdd.n1853 vdd.n768 185
R16256 vdd.n2064 vdd.n768 185
R16257 vdd.n1855 vdd.n1854 185
R16258 vdd.n1854 vdd.n766 185
R16259 vdd.n1856 vdd.n775 185
R16260 vdd.n2056 vdd.n775 185
R16261 vdd.n1858 vdd.n1857 185
R16262 vdd.n1857 vdd.n773 185
R16263 vdd.n1859 vdd.n781 185
R16264 vdd.n2050 vdd.n781 185
R16265 vdd.n1861 vdd.n1860 185
R16266 vdd.n1860 vdd.n779 185
R16267 vdd.n1862 vdd.n786 185
R16268 vdd.n2044 vdd.n786 185
R16269 vdd.n1864 vdd.n1863 185
R16270 vdd.n1863 vdd.n792 185
R16271 vdd.n1865 vdd.n791 185
R16272 vdd.n2038 vdd.n791 185
R16273 vdd.n1867 vdd.n1866 185
R16274 vdd.n1866 vdd.n798 185
R16275 vdd.n1868 vdd.n797 185
R16276 vdd.n2032 vdd.n797 185
R16277 vdd.n1870 vdd.n1869 185
R16278 vdd.n1871 vdd.n1870 185
R16279 vdd.n1851 vdd.n804 185
R16280 vdd.n2026 vdd.n804 185
R16281 vdd.n1850 vdd.n1849 185
R16282 vdd.n1849 vdd.n802 185
R16283 vdd.n1848 vdd.n810 185
R16284 vdd.n2020 vdd.n810 185
R16285 vdd.n1847 vdd.n1846 185
R16286 vdd.n1846 vdd.n808 185
R16287 vdd.n1845 vdd.n815 185
R16288 vdd.n2014 vdd.n815 185
R16289 vdd.n1844 vdd.n1843 185
R16290 vdd.n1843 vdd.n823 185
R16291 vdd.n1842 vdd.n822 185
R16292 vdd.n2007 vdd.n822 185
R16293 vdd.n1841 vdd.n1840 185
R16294 vdd.n1840 vdd.n820 185
R16295 vdd.n1839 vdd.n829 185
R16296 vdd.n2001 vdd.n829 185
R16297 vdd.n1838 vdd.n1837 185
R16298 vdd.n1837 vdd.n827 185
R16299 vdd.n1836 vdd.n835 185
R16300 vdd.n1995 vdd.n835 185
R16301 vdd.n1835 vdd.n1834 185
R16302 vdd.n1834 vdd.n833 185
R16303 vdd.n1833 vdd.n841 185
R16304 vdd.n1989 vdd.n841 185
R16305 vdd.n1986 vdd.n842 185
R16306 vdd.n1985 vdd.n1984 185
R16307 vdd.n1982 vdd.n843 185
R16308 vdd.n1980 vdd.n1979 185
R16309 vdd.n1978 vdd.n844 185
R16310 vdd.n1977 vdd.n1976 185
R16311 vdd.n1974 vdd.n845 185
R16312 vdd.n1972 vdd.n1971 185
R16313 vdd.n1970 vdd.n846 185
R16314 vdd.n1969 vdd.n1968 185
R16315 vdd.n1966 vdd.n847 185
R16316 vdd.n1964 vdd.n1963 185
R16317 vdd.n1962 vdd.n848 185
R16318 vdd.n1961 vdd.n1960 185
R16319 vdd.n1958 vdd.n849 185
R16320 vdd.n1956 vdd.n1955 185
R16321 vdd.n1954 vdd.n850 185
R16322 vdd.n1953 vdd.n852 185
R16323 vdd.n1798 vdd.n853 185
R16324 vdd.n1801 vdd.n1800 185
R16325 vdd.n1803 vdd.n1802 185
R16326 vdd.n1805 vdd.n1797 185
R16327 vdd.n1808 vdd.n1807 185
R16328 vdd.n1809 vdd.n1796 185
R16329 vdd.n1811 vdd.n1810 185
R16330 vdd.n1813 vdd.n1795 185
R16331 vdd.n1816 vdd.n1815 185
R16332 vdd.n1817 vdd.n1794 185
R16333 vdd.n1819 vdd.n1818 185
R16334 vdd.n1821 vdd.n1793 185
R16335 vdd.n1824 vdd.n1823 185
R16336 vdd.n1825 vdd.n1790 185
R16337 vdd.n1828 vdd.n1827 185
R16338 vdd.n1830 vdd.n1789 185
R16339 vdd.n1832 vdd.n1831 185
R16340 vdd.n1831 vdd.n839 185
R16341 vdd.n291 vdd.n290 171.744
R16342 vdd.n290 vdd.n289 171.744
R16343 vdd.n289 vdd.n258 171.744
R16344 vdd.n282 vdd.n258 171.744
R16345 vdd.n282 vdd.n281 171.744
R16346 vdd.n281 vdd.n263 171.744
R16347 vdd.n274 vdd.n263 171.744
R16348 vdd.n274 vdd.n273 171.744
R16349 vdd.n273 vdd.n267 171.744
R16350 vdd.n244 vdd.n243 171.744
R16351 vdd.n243 vdd.n242 171.744
R16352 vdd.n242 vdd.n211 171.744
R16353 vdd.n235 vdd.n211 171.744
R16354 vdd.n235 vdd.n234 171.744
R16355 vdd.n234 vdd.n216 171.744
R16356 vdd.n227 vdd.n216 171.744
R16357 vdd.n227 vdd.n226 171.744
R16358 vdd.n226 vdd.n220 171.744
R16359 vdd.n201 vdd.n200 171.744
R16360 vdd.n200 vdd.n199 171.744
R16361 vdd.n199 vdd.n168 171.744
R16362 vdd.n192 vdd.n168 171.744
R16363 vdd.n192 vdd.n191 171.744
R16364 vdd.n191 vdd.n173 171.744
R16365 vdd.n184 vdd.n173 171.744
R16366 vdd.n184 vdd.n183 171.744
R16367 vdd.n183 vdd.n177 171.744
R16368 vdd.n154 vdd.n153 171.744
R16369 vdd.n153 vdd.n152 171.744
R16370 vdd.n152 vdd.n121 171.744
R16371 vdd.n145 vdd.n121 171.744
R16372 vdd.n145 vdd.n144 171.744
R16373 vdd.n144 vdd.n126 171.744
R16374 vdd.n137 vdd.n126 171.744
R16375 vdd.n137 vdd.n136 171.744
R16376 vdd.n136 vdd.n130 171.744
R16377 vdd.n112 vdd.n111 171.744
R16378 vdd.n111 vdd.n110 171.744
R16379 vdd.n110 vdd.n79 171.744
R16380 vdd.n103 vdd.n79 171.744
R16381 vdd.n103 vdd.n102 171.744
R16382 vdd.n102 vdd.n84 171.744
R16383 vdd.n95 vdd.n84 171.744
R16384 vdd.n95 vdd.n94 171.744
R16385 vdd.n94 vdd.n88 171.744
R16386 vdd.n65 vdd.n64 171.744
R16387 vdd.n64 vdd.n63 171.744
R16388 vdd.n63 vdd.n32 171.744
R16389 vdd.n56 vdd.n32 171.744
R16390 vdd.n56 vdd.n55 171.744
R16391 vdd.n55 vdd.n37 171.744
R16392 vdd.n48 vdd.n37 171.744
R16393 vdd.n48 vdd.n47 171.744
R16394 vdd.n47 vdd.n41 171.744
R16395 vdd.n1106 vdd.n1105 171.744
R16396 vdd.n1105 vdd.n1104 171.744
R16397 vdd.n1104 vdd.n1073 171.744
R16398 vdd.n1097 vdd.n1073 171.744
R16399 vdd.n1097 vdd.n1096 171.744
R16400 vdd.n1096 vdd.n1078 171.744
R16401 vdd.n1089 vdd.n1078 171.744
R16402 vdd.n1089 vdd.n1088 171.744
R16403 vdd.n1088 vdd.n1082 171.744
R16404 vdd.n1153 vdd.n1152 171.744
R16405 vdd.n1152 vdd.n1151 171.744
R16406 vdd.n1151 vdd.n1120 171.744
R16407 vdd.n1144 vdd.n1120 171.744
R16408 vdd.n1144 vdd.n1143 171.744
R16409 vdd.n1143 vdd.n1125 171.744
R16410 vdd.n1136 vdd.n1125 171.744
R16411 vdd.n1136 vdd.n1135 171.744
R16412 vdd.n1135 vdd.n1129 171.744
R16413 vdd.n1016 vdd.n1015 171.744
R16414 vdd.n1015 vdd.n1014 171.744
R16415 vdd.n1014 vdd.n983 171.744
R16416 vdd.n1007 vdd.n983 171.744
R16417 vdd.n1007 vdd.n1006 171.744
R16418 vdd.n1006 vdd.n988 171.744
R16419 vdd.n999 vdd.n988 171.744
R16420 vdd.n999 vdd.n998 171.744
R16421 vdd.n998 vdd.n992 171.744
R16422 vdd.n1063 vdd.n1062 171.744
R16423 vdd.n1062 vdd.n1061 171.744
R16424 vdd.n1061 vdd.n1030 171.744
R16425 vdd.n1054 vdd.n1030 171.744
R16426 vdd.n1054 vdd.n1053 171.744
R16427 vdd.n1053 vdd.n1035 171.744
R16428 vdd.n1046 vdd.n1035 171.744
R16429 vdd.n1046 vdd.n1045 171.744
R16430 vdd.n1045 vdd.n1039 171.744
R16431 vdd.n927 vdd.n926 171.744
R16432 vdd.n926 vdd.n925 171.744
R16433 vdd.n925 vdd.n894 171.744
R16434 vdd.n918 vdd.n894 171.744
R16435 vdd.n918 vdd.n917 171.744
R16436 vdd.n917 vdd.n899 171.744
R16437 vdd.n910 vdd.n899 171.744
R16438 vdd.n910 vdd.n909 171.744
R16439 vdd.n909 vdd.n903 171.744
R16440 vdd.n974 vdd.n973 171.744
R16441 vdd.n973 vdd.n972 171.744
R16442 vdd.n972 vdd.n941 171.744
R16443 vdd.n965 vdd.n941 171.744
R16444 vdd.n965 vdd.n964 171.744
R16445 vdd.n964 vdd.n946 171.744
R16446 vdd.n957 vdd.n946 171.744
R16447 vdd.n957 vdd.n956 171.744
R16448 vdd.n956 vdd.n950 171.744
R16449 vdd.n3017 vdd.n334 146.341
R16450 vdd.n3015 vdd.n3014 146.341
R16451 vdd.n3012 vdd.n338 146.341
R16452 vdd.n3008 vdd.n3007 146.341
R16453 vdd.n3005 vdd.n346 146.341
R16454 vdd.n3001 vdd.n3000 146.341
R16455 vdd.n2998 vdd.n353 146.341
R16456 vdd.n2994 vdd.n2993 146.341
R16457 vdd.n2991 vdd.n360 146.341
R16458 vdd.n371 vdd.n368 146.341
R16459 vdd.n2983 vdd.n2982 146.341
R16460 vdd.n2980 vdd.n373 146.341
R16461 vdd.n2976 vdd.n2975 146.341
R16462 vdd.n2973 vdd.n379 146.341
R16463 vdd.n2969 vdd.n2968 146.341
R16464 vdd.n2966 vdd.n386 146.341
R16465 vdd.n2962 vdd.n2961 146.341
R16466 vdd.n2959 vdd.n393 146.341
R16467 vdd.n2955 vdd.n2954 146.341
R16468 vdd.n2952 vdd.n400 146.341
R16469 vdd.n411 vdd.n408 146.341
R16470 vdd.n2944 vdd.n2943 146.341
R16471 vdd.n2941 vdd.n413 146.341
R16472 vdd.n2937 vdd.n2936 146.341
R16473 vdd.n2934 vdd.n419 146.341
R16474 vdd.n2930 vdd.n2929 146.341
R16475 vdd.n2927 vdd.n426 146.341
R16476 vdd.n2923 vdd.n2922 146.341
R16477 vdd.n2920 vdd.n433 146.341
R16478 vdd.n2916 vdd.n2915 146.341
R16479 vdd.n2913 vdd.n440 146.341
R16480 vdd.n2850 vdd.n478 146.341
R16481 vdd.n2850 vdd.n474 146.341
R16482 vdd.n2856 vdd.n474 146.341
R16483 vdd.n2856 vdd.n466 146.341
R16484 vdd.n2867 vdd.n466 146.341
R16485 vdd.n2867 vdd.n462 146.341
R16486 vdd.n2873 vdd.n462 146.341
R16487 vdd.n2873 vdd.n454 146.341
R16488 vdd.n2883 vdd.n454 146.341
R16489 vdd.n2883 vdd.n455 146.341
R16490 vdd.n455 vdd.n305 146.341
R16491 vdd.n306 vdd.n305 146.341
R16492 vdd.n307 vdd.n306 146.341
R16493 vdd.n448 vdd.n307 146.341
R16494 vdd.n448 vdd.n315 146.341
R16495 vdd.n316 vdd.n315 146.341
R16496 vdd.n317 vdd.n316 146.341
R16497 vdd.n445 vdd.n317 146.341
R16498 vdd.n445 vdd.n326 146.341
R16499 vdd.n327 vdd.n326 146.341
R16500 vdd.n328 vdd.n327 146.341
R16501 vdd.n2839 vdd.n483 146.341
R16502 vdd.n2839 vdd.n517 146.341
R16503 vdd.n523 vdd.n522 146.341
R16504 vdd.n2832 vdd.n2831 146.341
R16505 vdd.n2828 vdd.n2827 146.341
R16506 vdd.n2824 vdd.n2823 146.341
R16507 vdd.n2820 vdd.n2819 146.341
R16508 vdd.n2816 vdd.n2815 146.341
R16509 vdd.n2812 vdd.n2811 146.341
R16510 vdd.n2808 vdd.n2807 146.341
R16511 vdd.n2799 vdd.n2798 146.341
R16512 vdd.n2796 vdd.n2795 146.341
R16513 vdd.n2792 vdd.n2791 146.341
R16514 vdd.n2788 vdd.n2787 146.341
R16515 vdd.n2784 vdd.n2783 146.341
R16516 vdd.n2780 vdd.n2779 146.341
R16517 vdd.n2776 vdd.n2775 146.341
R16518 vdd.n2772 vdd.n2771 146.341
R16519 vdd.n2768 vdd.n2767 146.341
R16520 vdd.n2764 vdd.n2763 146.341
R16521 vdd.n2760 vdd.n2759 146.341
R16522 vdd.n2753 vdd.n2752 146.341
R16523 vdd.n2750 vdd.n2749 146.341
R16524 vdd.n2746 vdd.n2745 146.341
R16525 vdd.n2742 vdd.n2741 146.341
R16526 vdd.n2738 vdd.n2737 146.341
R16527 vdd.n2734 vdd.n2733 146.341
R16528 vdd.n2730 vdd.n2729 146.341
R16529 vdd.n2726 vdd.n2725 146.341
R16530 vdd.n2722 vdd.n2721 146.341
R16531 vdd.n2718 vdd.n2717 146.341
R16532 vdd.n2714 vdd.n515 146.341
R16533 vdd.n2848 vdd.n479 146.341
R16534 vdd.n2848 vdd.n472 146.341
R16535 vdd.n2859 vdd.n472 146.341
R16536 vdd.n2859 vdd.n468 146.341
R16537 vdd.n2865 vdd.n468 146.341
R16538 vdd.n2865 vdd.n461 146.341
R16539 vdd.n2875 vdd.n461 146.341
R16540 vdd.n2875 vdd.n457 146.341
R16541 vdd.n2881 vdd.n457 146.341
R16542 vdd.n2881 vdd.n302 146.341
R16543 vdd.n3044 vdd.n302 146.341
R16544 vdd.n3044 vdd.n303 146.341
R16545 vdd.n3040 vdd.n303 146.341
R16546 vdd.n3040 vdd.n309 146.341
R16547 vdd.n3036 vdd.n309 146.341
R16548 vdd.n3036 vdd.n314 146.341
R16549 vdd.n3032 vdd.n314 146.341
R16550 vdd.n3032 vdd.n319 146.341
R16551 vdd.n3028 vdd.n319 146.341
R16552 vdd.n3028 vdd.n325 146.341
R16553 vdd.n3024 vdd.n325 146.341
R16554 vdd.n1936 vdd.n1935 146.341
R16555 vdd.n1933 vdd.n1517 146.341
R16556 vdd.n1713 vdd.n1523 146.341
R16557 vdd.n1711 vdd.n1710 146.341
R16558 vdd.n1708 vdd.n1525 146.341
R16559 vdd.n1704 vdd.n1703 146.341
R16560 vdd.n1701 vdd.n1532 146.341
R16561 vdd.n1697 vdd.n1696 146.341
R16562 vdd.n1694 vdd.n1539 146.341
R16563 vdd.n1550 vdd.n1547 146.341
R16564 vdd.n1686 vdd.n1685 146.341
R16565 vdd.n1683 vdd.n1552 146.341
R16566 vdd.n1679 vdd.n1678 146.341
R16567 vdd.n1676 vdd.n1558 146.341
R16568 vdd.n1672 vdd.n1671 146.341
R16569 vdd.n1669 vdd.n1565 146.341
R16570 vdd.n1665 vdd.n1664 146.341
R16571 vdd.n1662 vdd.n1572 146.341
R16572 vdd.n1658 vdd.n1657 146.341
R16573 vdd.n1655 vdd.n1579 146.341
R16574 vdd.n1590 vdd.n1587 146.341
R16575 vdd.n1647 vdd.n1646 146.341
R16576 vdd.n1644 vdd.n1592 146.341
R16577 vdd.n1640 vdd.n1639 146.341
R16578 vdd.n1637 vdd.n1598 146.341
R16579 vdd.n1633 vdd.n1632 146.341
R16580 vdd.n1630 vdd.n1605 146.341
R16581 vdd.n1626 vdd.n1625 146.341
R16582 vdd.n1623 vdd.n1620 146.341
R16583 vdd.n1618 vdd.n1615 146.341
R16584 vdd.n1613 vdd.n859 146.341
R16585 vdd.n1431 vdd.n1191 146.341
R16586 vdd.n1431 vdd.n1187 146.341
R16587 vdd.n1437 vdd.n1187 146.341
R16588 vdd.n1437 vdd.n1179 146.341
R16589 vdd.n1448 vdd.n1179 146.341
R16590 vdd.n1448 vdd.n1175 146.341
R16591 vdd.n1454 vdd.n1175 146.341
R16592 vdd.n1454 vdd.n1169 146.341
R16593 vdd.n1466 vdd.n1169 146.341
R16594 vdd.n1466 vdd.n1165 146.341
R16595 vdd.n1472 vdd.n1165 146.341
R16596 vdd.n1472 vdd.n886 146.341
R16597 vdd.n1482 vdd.n886 146.341
R16598 vdd.n1482 vdd.n882 146.341
R16599 vdd.n1488 vdd.n882 146.341
R16600 vdd.n1488 vdd.n876 146.341
R16601 vdd.n1499 vdd.n876 146.341
R16602 vdd.n1499 vdd.n871 146.341
R16603 vdd.n1507 vdd.n871 146.341
R16604 vdd.n1507 vdd.n861 146.341
R16605 vdd.n1944 vdd.n861 146.341
R16606 vdd.n1420 vdd.n1196 146.341
R16607 vdd.n1420 vdd.n1229 146.341
R16608 vdd.n1233 vdd.n1232 146.341
R16609 vdd.n1235 vdd.n1234 146.341
R16610 vdd.n1239 vdd.n1238 146.341
R16611 vdd.n1241 vdd.n1240 146.341
R16612 vdd.n1245 vdd.n1244 146.341
R16613 vdd.n1247 vdd.n1246 146.341
R16614 vdd.n1251 vdd.n1250 146.341
R16615 vdd.n1253 vdd.n1252 146.341
R16616 vdd.n1259 vdd.n1258 146.341
R16617 vdd.n1261 vdd.n1260 146.341
R16618 vdd.n1265 vdd.n1264 146.341
R16619 vdd.n1267 vdd.n1266 146.341
R16620 vdd.n1271 vdd.n1270 146.341
R16621 vdd.n1273 vdd.n1272 146.341
R16622 vdd.n1277 vdd.n1276 146.341
R16623 vdd.n1279 vdd.n1278 146.341
R16624 vdd.n1283 vdd.n1282 146.341
R16625 vdd.n1285 vdd.n1284 146.341
R16626 vdd.n1357 vdd.n1288 146.341
R16627 vdd.n1290 vdd.n1289 146.341
R16628 vdd.n1294 vdd.n1293 146.341
R16629 vdd.n1296 vdd.n1295 146.341
R16630 vdd.n1300 vdd.n1299 146.341
R16631 vdd.n1302 vdd.n1301 146.341
R16632 vdd.n1306 vdd.n1305 146.341
R16633 vdd.n1308 vdd.n1307 146.341
R16634 vdd.n1312 vdd.n1311 146.341
R16635 vdd.n1314 vdd.n1313 146.341
R16636 vdd.n1318 vdd.n1317 146.341
R16637 vdd.n1319 vdd.n1227 146.341
R16638 vdd.n1429 vdd.n1192 146.341
R16639 vdd.n1429 vdd.n1185 146.341
R16640 vdd.n1440 vdd.n1185 146.341
R16641 vdd.n1440 vdd.n1181 146.341
R16642 vdd.n1446 vdd.n1181 146.341
R16643 vdd.n1446 vdd.n1174 146.341
R16644 vdd.n1457 vdd.n1174 146.341
R16645 vdd.n1457 vdd.n1170 146.341
R16646 vdd.n1464 vdd.n1170 146.341
R16647 vdd.n1464 vdd.n1163 146.341
R16648 vdd.n1474 vdd.n1163 146.341
R16649 vdd.n1474 vdd.n889 146.341
R16650 vdd.n1480 vdd.n889 146.341
R16651 vdd.n1480 vdd.n881 146.341
R16652 vdd.n1491 vdd.n881 146.341
R16653 vdd.n1491 vdd.n877 146.341
R16654 vdd.n1497 vdd.n877 146.341
R16655 vdd.n1497 vdd.n869 146.341
R16656 vdd.n1510 vdd.n869 146.341
R16657 vdd.n1510 vdd.n864 146.341
R16658 vdd.n1942 vdd.n864 146.341
R16659 vdd.n863 vdd.n839 141.707
R16660 vdd.n2840 vdd.n484 141.707
R16661 vdd.n1791 vdd.t91 127.284
R16662 vdd.n755 vdd.t75 127.284
R16663 vdd.n1765 vdd.t116 127.284
R16664 vdd.n747 vdd.t106 127.284
R16665 vdd.n2536 vdd.t58 127.284
R16666 vdd.n2536 vdd.t59 127.284
R16667 vdd.n2256 vdd.t98 127.284
R16668 vdd.n622 vdd.t79 127.284
R16669 vdd.n2253 vdd.t84 127.284
R16670 vdd.n589 vdd.t86 127.284
R16671 vdd.n817 vdd.t94 127.284
R16672 vdd.n817 vdd.t95 127.284
R16673 vdd.n22 vdd.n20 117.314
R16674 vdd.n17 vdd.n15 117.314
R16675 vdd.n27 vdd.n26 116.927
R16676 vdd.n24 vdd.n23 116.927
R16677 vdd.n22 vdd.n21 116.927
R16678 vdd.n17 vdd.n16 116.927
R16679 vdd.n19 vdd.n18 116.927
R16680 vdd.n27 vdd.n25 116.927
R16681 vdd.n1792 vdd.t90 111.188
R16682 vdd.n756 vdd.t76 111.188
R16683 vdd.n1766 vdd.t115 111.188
R16684 vdd.n748 vdd.t107 111.188
R16685 vdd.n2257 vdd.t97 111.188
R16686 vdd.n623 vdd.t80 111.188
R16687 vdd.n2254 vdd.t83 111.188
R16688 vdd.n590 vdd.t87 111.188
R16689 vdd.n2479 vdd.n701 99.5127
R16690 vdd.n2483 vdd.n701 99.5127
R16691 vdd.n2483 vdd.n693 99.5127
R16692 vdd.n2491 vdd.n693 99.5127
R16693 vdd.n2491 vdd.n691 99.5127
R16694 vdd.n2495 vdd.n691 99.5127
R16695 vdd.n2495 vdd.n680 99.5127
R16696 vdd.n2503 vdd.n680 99.5127
R16697 vdd.n2503 vdd.n678 99.5127
R16698 vdd.n2507 vdd.n678 99.5127
R16699 vdd.n2507 vdd.n669 99.5127
R16700 vdd.n2515 vdd.n669 99.5127
R16701 vdd.n2515 vdd.n667 99.5127
R16702 vdd.n2519 vdd.n667 99.5127
R16703 vdd.n2519 vdd.n657 99.5127
R16704 vdd.n2527 vdd.n657 99.5127
R16705 vdd.n2527 vdd.n655 99.5127
R16706 vdd.n2531 vdd.n655 99.5127
R16707 vdd.n2531 vdd.n646 99.5127
R16708 vdd.n2541 vdd.n646 99.5127
R16709 vdd.n2541 vdd.n644 99.5127
R16710 vdd.n2545 vdd.n644 99.5127
R16711 vdd.n2545 vdd.n632 99.5127
R16712 vdd.n2598 vdd.n632 99.5127
R16713 vdd.n2598 vdd.n630 99.5127
R16714 vdd.n2602 vdd.n630 99.5127
R16715 vdd.n2602 vdd.n598 99.5127
R16716 vdd.n2672 vdd.n598 99.5127
R16717 vdd.n2668 vdd.n599 99.5127
R16718 vdd.n2666 vdd.n2665 99.5127
R16719 vdd.n2663 vdd.n603 99.5127
R16720 vdd.n2659 vdd.n2658 99.5127
R16721 vdd.n2656 vdd.n606 99.5127
R16722 vdd.n2652 vdd.n2651 99.5127
R16723 vdd.n2649 vdd.n609 99.5127
R16724 vdd.n2645 vdd.n2644 99.5127
R16725 vdd.n2642 vdd.n2640 99.5127
R16726 vdd.n2638 vdd.n612 99.5127
R16727 vdd.n2634 vdd.n2633 99.5127
R16728 vdd.n2631 vdd.n615 99.5127
R16729 vdd.n2627 vdd.n2626 99.5127
R16730 vdd.n2624 vdd.n618 99.5127
R16731 vdd.n2620 vdd.n2619 99.5127
R16732 vdd.n2617 vdd.n621 99.5127
R16733 vdd.n2612 vdd.n2611 99.5127
R16734 vdd.n2399 vdd.n704 99.5127
R16735 vdd.n2399 vdd.n699 99.5127
R16736 vdd.n2396 vdd.n699 99.5127
R16737 vdd.n2396 vdd.n694 99.5127
R16738 vdd.n2343 vdd.n694 99.5127
R16739 vdd.n2343 vdd.n688 99.5127
R16740 vdd.n2346 vdd.n688 99.5127
R16741 vdd.n2346 vdd.n681 99.5127
R16742 vdd.n2349 vdd.n681 99.5127
R16743 vdd.n2349 vdd.n676 99.5127
R16744 vdd.n2352 vdd.n676 99.5127
R16745 vdd.n2352 vdd.n671 99.5127
R16746 vdd.n2355 vdd.n671 99.5127
R16747 vdd.n2355 vdd.n665 99.5127
R16748 vdd.n2373 vdd.n665 99.5127
R16749 vdd.n2373 vdd.n658 99.5127
R16750 vdd.n2369 vdd.n658 99.5127
R16751 vdd.n2369 vdd.n653 99.5127
R16752 vdd.n2366 vdd.n653 99.5127
R16753 vdd.n2366 vdd.n648 99.5127
R16754 vdd.n2363 vdd.n648 99.5127
R16755 vdd.n2363 vdd.n642 99.5127
R16756 vdd.n2360 vdd.n642 99.5127
R16757 vdd.n2360 vdd.n634 99.5127
R16758 vdd.n634 vdd.n627 99.5127
R16759 vdd.n2604 vdd.n627 99.5127
R16760 vdd.n2605 vdd.n2604 99.5127
R16761 vdd.n2605 vdd.n596 99.5127
R16762 vdd.n2469 vdd.n2252 99.5127
R16763 vdd.n2465 vdd.n2252 99.5127
R16764 vdd.n2463 vdd.n2462 99.5127
R16765 vdd.n2459 vdd.n2458 99.5127
R16766 vdd.n2455 vdd.n2454 99.5127
R16767 vdd.n2451 vdd.n2450 99.5127
R16768 vdd.n2447 vdd.n2446 99.5127
R16769 vdd.n2443 vdd.n2442 99.5127
R16770 vdd.n2439 vdd.n2438 99.5127
R16771 vdd.n2435 vdd.n2434 99.5127
R16772 vdd.n2431 vdd.n2430 99.5127
R16773 vdd.n2427 vdd.n2426 99.5127
R16774 vdd.n2423 vdd.n2422 99.5127
R16775 vdd.n2419 vdd.n2418 99.5127
R16776 vdd.n2415 vdd.n2414 99.5127
R16777 vdd.n2411 vdd.n2410 99.5127
R16778 vdd.n2406 vdd.n2405 99.5127
R16779 vdd.n2217 vdd.n745 99.5127
R16780 vdd.n2213 vdd.n2212 99.5127
R16781 vdd.n2209 vdd.n2208 99.5127
R16782 vdd.n2205 vdd.n2204 99.5127
R16783 vdd.n2201 vdd.n2200 99.5127
R16784 vdd.n2197 vdd.n2196 99.5127
R16785 vdd.n2193 vdd.n2192 99.5127
R16786 vdd.n2189 vdd.n2188 99.5127
R16787 vdd.n2185 vdd.n2184 99.5127
R16788 vdd.n2181 vdd.n2180 99.5127
R16789 vdd.n2177 vdd.n2176 99.5127
R16790 vdd.n2173 vdd.n2172 99.5127
R16791 vdd.n2169 vdd.n2168 99.5127
R16792 vdd.n2165 vdd.n2164 99.5127
R16793 vdd.n2161 vdd.n2160 99.5127
R16794 vdd.n2157 vdd.n2156 99.5127
R16795 vdd.n2152 vdd.n2151 99.5127
R16796 vdd.n1890 vdd.n840 99.5127
R16797 vdd.n1890 vdd.n834 99.5127
R16798 vdd.n1887 vdd.n834 99.5127
R16799 vdd.n1887 vdd.n828 99.5127
R16800 vdd.n1884 vdd.n828 99.5127
R16801 vdd.n1884 vdd.n821 99.5127
R16802 vdd.n1881 vdd.n821 99.5127
R16803 vdd.n1881 vdd.n814 99.5127
R16804 vdd.n1878 vdd.n814 99.5127
R16805 vdd.n1878 vdd.n809 99.5127
R16806 vdd.n1875 vdd.n809 99.5127
R16807 vdd.n1875 vdd.n803 99.5127
R16808 vdd.n1872 vdd.n803 99.5127
R16809 vdd.n1872 vdd.n796 99.5127
R16810 vdd.n1786 vdd.n796 99.5127
R16811 vdd.n1786 vdd.n790 99.5127
R16812 vdd.n1783 vdd.n790 99.5127
R16813 vdd.n1783 vdd.n785 99.5127
R16814 vdd.n1780 vdd.n785 99.5127
R16815 vdd.n1780 vdd.n780 99.5127
R16816 vdd.n1777 vdd.n780 99.5127
R16817 vdd.n1777 vdd.n774 99.5127
R16818 vdd.n1774 vdd.n774 99.5127
R16819 vdd.n1774 vdd.n767 99.5127
R16820 vdd.n1771 vdd.n767 99.5127
R16821 vdd.n1771 vdd.n760 99.5127
R16822 vdd.n760 vdd.n750 99.5127
R16823 vdd.n2147 vdd.n750 99.5127
R16824 vdd.n1725 vdd.n1723 99.5127
R16825 vdd.n1729 vdd.n1723 99.5127
R16826 vdd.n1733 vdd.n1731 99.5127
R16827 vdd.n1737 vdd.n1721 99.5127
R16828 vdd.n1741 vdd.n1739 99.5127
R16829 vdd.n1745 vdd.n1719 99.5127
R16830 vdd.n1749 vdd.n1747 99.5127
R16831 vdd.n1753 vdd.n1717 99.5127
R16832 vdd.n1756 vdd.n1755 99.5127
R16833 vdd.n1926 vdd.n1924 99.5127
R16834 vdd.n1922 vdd.n1758 99.5127
R16835 vdd.n1918 vdd.n1916 99.5127
R16836 vdd.n1914 vdd.n1760 99.5127
R16837 vdd.n1910 vdd.n1908 99.5127
R16838 vdd.n1906 vdd.n1762 99.5127
R16839 vdd.n1902 vdd.n1900 99.5127
R16840 vdd.n1898 vdd.n1764 99.5127
R16841 vdd.n1990 vdd.n836 99.5127
R16842 vdd.n1994 vdd.n836 99.5127
R16843 vdd.n1994 vdd.n826 99.5127
R16844 vdd.n2002 vdd.n826 99.5127
R16845 vdd.n2002 vdd.n824 99.5127
R16846 vdd.n2006 vdd.n824 99.5127
R16847 vdd.n2006 vdd.n813 99.5127
R16848 vdd.n2015 vdd.n813 99.5127
R16849 vdd.n2015 vdd.n811 99.5127
R16850 vdd.n2019 vdd.n811 99.5127
R16851 vdd.n2019 vdd.n801 99.5127
R16852 vdd.n2027 vdd.n801 99.5127
R16853 vdd.n2027 vdd.n799 99.5127
R16854 vdd.n2031 vdd.n799 99.5127
R16855 vdd.n2031 vdd.n789 99.5127
R16856 vdd.n2039 vdd.n789 99.5127
R16857 vdd.n2039 vdd.n787 99.5127
R16858 vdd.n2043 vdd.n787 99.5127
R16859 vdd.n2043 vdd.n778 99.5127
R16860 vdd.n2051 vdd.n778 99.5127
R16861 vdd.n2051 vdd.n776 99.5127
R16862 vdd.n2055 vdd.n776 99.5127
R16863 vdd.n2055 vdd.n765 99.5127
R16864 vdd.n2065 vdd.n765 99.5127
R16865 vdd.n2065 vdd.n762 99.5127
R16866 vdd.n2070 vdd.n762 99.5127
R16867 vdd.n2070 vdd.n763 99.5127
R16868 vdd.n763 vdd.n744 99.5127
R16869 vdd.n2588 vdd.n2587 99.5127
R16870 vdd.n2585 vdd.n2551 99.5127
R16871 vdd.n2581 vdd.n2580 99.5127
R16872 vdd.n2578 vdd.n2554 99.5127
R16873 vdd.n2574 vdd.n2573 99.5127
R16874 vdd.n2571 vdd.n2557 99.5127
R16875 vdd.n2567 vdd.n2566 99.5127
R16876 vdd.n2564 vdd.n2561 99.5127
R16877 vdd.n2705 vdd.n577 99.5127
R16878 vdd.n2703 vdd.n2702 99.5127
R16879 vdd.n2700 vdd.n579 99.5127
R16880 vdd.n2696 vdd.n2695 99.5127
R16881 vdd.n2693 vdd.n582 99.5127
R16882 vdd.n2689 vdd.n2688 99.5127
R16883 vdd.n2686 vdd.n585 99.5127
R16884 vdd.n2682 vdd.n2681 99.5127
R16885 vdd.n2679 vdd.n588 99.5127
R16886 vdd.n2323 vdd.n705 99.5127
R16887 vdd.n2323 vdd.n700 99.5127
R16888 vdd.n2394 vdd.n700 99.5127
R16889 vdd.n2394 vdd.n695 99.5127
R16890 vdd.n2390 vdd.n695 99.5127
R16891 vdd.n2390 vdd.n689 99.5127
R16892 vdd.n2387 vdd.n689 99.5127
R16893 vdd.n2387 vdd.n682 99.5127
R16894 vdd.n2384 vdd.n682 99.5127
R16895 vdd.n2384 vdd.n677 99.5127
R16896 vdd.n2381 vdd.n677 99.5127
R16897 vdd.n2381 vdd.n672 99.5127
R16898 vdd.n2378 vdd.n672 99.5127
R16899 vdd.n2378 vdd.n666 99.5127
R16900 vdd.n2375 vdd.n666 99.5127
R16901 vdd.n2375 vdd.n659 99.5127
R16902 vdd.n2340 vdd.n659 99.5127
R16903 vdd.n2340 vdd.n654 99.5127
R16904 vdd.n2337 vdd.n654 99.5127
R16905 vdd.n2337 vdd.n649 99.5127
R16906 vdd.n2334 vdd.n649 99.5127
R16907 vdd.n2334 vdd.n643 99.5127
R16908 vdd.n2331 vdd.n643 99.5127
R16909 vdd.n2331 vdd.n635 99.5127
R16910 vdd.n2328 vdd.n635 99.5127
R16911 vdd.n2328 vdd.n628 99.5127
R16912 vdd.n628 vdd.n594 99.5127
R16913 vdd.n2674 vdd.n594 99.5127
R16914 vdd.n2473 vdd.n708 99.5127
R16915 vdd.n2261 vdd.n2260 99.5127
R16916 vdd.n2265 vdd.n2264 99.5127
R16917 vdd.n2269 vdd.n2268 99.5127
R16918 vdd.n2273 vdd.n2272 99.5127
R16919 vdd.n2277 vdd.n2276 99.5127
R16920 vdd.n2281 vdd.n2280 99.5127
R16921 vdd.n2285 vdd.n2284 99.5127
R16922 vdd.n2289 vdd.n2288 99.5127
R16923 vdd.n2293 vdd.n2292 99.5127
R16924 vdd.n2297 vdd.n2296 99.5127
R16925 vdd.n2301 vdd.n2300 99.5127
R16926 vdd.n2305 vdd.n2304 99.5127
R16927 vdd.n2309 vdd.n2308 99.5127
R16928 vdd.n2313 vdd.n2312 99.5127
R16929 vdd.n2317 vdd.n2316 99.5127
R16930 vdd.n2319 vdd.n2251 99.5127
R16931 vdd.n2477 vdd.n698 99.5127
R16932 vdd.n2485 vdd.n698 99.5127
R16933 vdd.n2485 vdd.n696 99.5127
R16934 vdd.n2489 vdd.n696 99.5127
R16935 vdd.n2489 vdd.n686 99.5127
R16936 vdd.n2497 vdd.n686 99.5127
R16937 vdd.n2497 vdd.n684 99.5127
R16938 vdd.n2501 vdd.n684 99.5127
R16939 vdd.n2501 vdd.n675 99.5127
R16940 vdd.n2509 vdd.n675 99.5127
R16941 vdd.n2509 vdd.n673 99.5127
R16942 vdd.n2513 vdd.n673 99.5127
R16943 vdd.n2513 vdd.n663 99.5127
R16944 vdd.n2521 vdd.n663 99.5127
R16945 vdd.n2521 vdd.n661 99.5127
R16946 vdd.n2525 vdd.n661 99.5127
R16947 vdd.n2525 vdd.n652 99.5127
R16948 vdd.n2533 vdd.n652 99.5127
R16949 vdd.n2533 vdd.n650 99.5127
R16950 vdd.n2539 vdd.n650 99.5127
R16951 vdd.n2539 vdd.n640 99.5127
R16952 vdd.n2547 vdd.n640 99.5127
R16953 vdd.n2547 vdd.n637 99.5127
R16954 vdd.n2596 vdd.n637 99.5127
R16955 vdd.n2596 vdd.n638 99.5127
R16956 vdd.n638 vdd.n629 99.5127
R16957 vdd.n2591 vdd.n629 99.5127
R16958 vdd.n2591 vdd.n597 99.5127
R16959 vdd.n2141 vdd.n2140 99.5127
R16960 vdd.n2137 vdd.n2136 99.5127
R16961 vdd.n2133 vdd.n2132 99.5127
R16962 vdd.n2129 vdd.n2128 99.5127
R16963 vdd.n2125 vdd.n2124 99.5127
R16964 vdd.n2121 vdd.n2120 99.5127
R16965 vdd.n2117 vdd.n2116 99.5127
R16966 vdd.n2113 vdd.n2112 99.5127
R16967 vdd.n2109 vdd.n2108 99.5127
R16968 vdd.n2105 vdd.n2104 99.5127
R16969 vdd.n2101 vdd.n2100 99.5127
R16970 vdd.n2097 vdd.n2096 99.5127
R16971 vdd.n2093 vdd.n2092 99.5127
R16972 vdd.n2089 vdd.n2088 99.5127
R16973 vdd.n2085 vdd.n2084 99.5127
R16974 vdd.n2081 vdd.n2080 99.5127
R16975 vdd.n2077 vdd.n726 99.5127
R16976 vdd.n1834 vdd.n841 99.5127
R16977 vdd.n1834 vdd.n835 99.5127
R16978 vdd.n1837 vdd.n835 99.5127
R16979 vdd.n1837 vdd.n829 99.5127
R16980 vdd.n1840 vdd.n829 99.5127
R16981 vdd.n1840 vdd.n822 99.5127
R16982 vdd.n1843 vdd.n822 99.5127
R16983 vdd.n1843 vdd.n815 99.5127
R16984 vdd.n1846 vdd.n815 99.5127
R16985 vdd.n1846 vdd.n810 99.5127
R16986 vdd.n1849 vdd.n810 99.5127
R16987 vdd.n1849 vdd.n804 99.5127
R16988 vdd.n1870 vdd.n804 99.5127
R16989 vdd.n1870 vdd.n797 99.5127
R16990 vdd.n1866 vdd.n797 99.5127
R16991 vdd.n1866 vdd.n791 99.5127
R16992 vdd.n1863 vdd.n791 99.5127
R16993 vdd.n1863 vdd.n786 99.5127
R16994 vdd.n1860 vdd.n786 99.5127
R16995 vdd.n1860 vdd.n781 99.5127
R16996 vdd.n1857 vdd.n781 99.5127
R16997 vdd.n1857 vdd.n775 99.5127
R16998 vdd.n1854 vdd.n775 99.5127
R16999 vdd.n1854 vdd.n768 99.5127
R17000 vdd.n768 vdd.n759 99.5127
R17001 vdd.n2072 vdd.n759 99.5127
R17002 vdd.n2073 vdd.n2072 99.5127
R17003 vdd.n2073 vdd.n751 99.5127
R17004 vdd.n1984 vdd.n1982 99.5127
R17005 vdd.n1980 vdd.n844 99.5127
R17006 vdd.n1976 vdd.n1974 99.5127
R17007 vdd.n1972 vdd.n846 99.5127
R17008 vdd.n1968 vdd.n1966 99.5127
R17009 vdd.n1964 vdd.n848 99.5127
R17010 vdd.n1960 vdd.n1958 99.5127
R17011 vdd.n1956 vdd.n850 99.5127
R17012 vdd.n1798 vdd.n852 99.5127
R17013 vdd.n1803 vdd.n1800 99.5127
R17014 vdd.n1807 vdd.n1805 99.5127
R17015 vdd.n1811 vdd.n1796 99.5127
R17016 vdd.n1815 vdd.n1813 99.5127
R17017 vdd.n1819 vdd.n1794 99.5127
R17018 vdd.n1823 vdd.n1821 99.5127
R17019 vdd.n1828 vdd.n1790 99.5127
R17020 vdd.n1831 vdd.n1830 99.5127
R17021 vdd.n1988 vdd.n832 99.5127
R17022 vdd.n1996 vdd.n832 99.5127
R17023 vdd.n1996 vdd.n830 99.5127
R17024 vdd.n2000 vdd.n830 99.5127
R17025 vdd.n2000 vdd.n819 99.5127
R17026 vdd.n2008 vdd.n819 99.5127
R17027 vdd.n2008 vdd.n816 99.5127
R17028 vdd.n2013 vdd.n816 99.5127
R17029 vdd.n2013 vdd.n807 99.5127
R17030 vdd.n2021 vdd.n807 99.5127
R17031 vdd.n2021 vdd.n805 99.5127
R17032 vdd.n2025 vdd.n805 99.5127
R17033 vdd.n2025 vdd.n795 99.5127
R17034 vdd.n2033 vdd.n795 99.5127
R17035 vdd.n2033 vdd.n793 99.5127
R17036 vdd.n2037 vdd.n793 99.5127
R17037 vdd.n2037 vdd.n784 99.5127
R17038 vdd.n2045 vdd.n784 99.5127
R17039 vdd.n2045 vdd.n782 99.5127
R17040 vdd.n2049 vdd.n782 99.5127
R17041 vdd.n2049 vdd.n772 99.5127
R17042 vdd.n2057 vdd.n772 99.5127
R17043 vdd.n2057 vdd.n769 99.5127
R17044 vdd.n2063 vdd.n769 99.5127
R17045 vdd.n2063 vdd.n770 99.5127
R17046 vdd.n770 vdd.n761 99.5127
R17047 vdd.n761 vdd.n752 99.5127
R17048 vdd.n2145 vdd.n752 99.5127
R17049 vdd.n9 vdd.n7 98.9633
R17050 vdd.n2 vdd.n0 98.9633
R17051 vdd.n9 vdd.n8 98.6055
R17052 vdd.n11 vdd.n10 98.6055
R17053 vdd.n13 vdd.n12 98.6055
R17054 vdd.n6 vdd.n5 98.6055
R17055 vdd.n4 vdd.n3 98.6055
R17056 vdd.n2 vdd.n1 98.6055
R17057 vdd.t141 vdd.n267 85.8723
R17058 vdd.t152 vdd.n220 85.8723
R17059 vdd.t137 vdd.n177 85.8723
R17060 vdd.t147 vdd.n130 85.8723
R17061 vdd.t178 vdd.n88 85.8723
R17062 vdd.t120 vdd.n41 85.8723
R17063 vdd.t176 vdd.n1082 85.8723
R17064 vdd.t162 vdd.n1129 85.8723
R17065 vdd.t168 vdd.n992 85.8723
R17066 vdd.t155 vdd.n1039 85.8723
R17067 vdd.t118 vdd.n903 85.8723
R17068 vdd.t177 vdd.n950 85.8723
R17069 vdd.n2537 vdd.n2536 78.546
R17070 vdd.n2011 vdd.n817 78.546
R17071 vdd.n254 vdd.n253 75.1835
R17072 vdd.n252 vdd.n251 75.1835
R17073 vdd.n250 vdd.n249 75.1835
R17074 vdd.n164 vdd.n163 75.1835
R17075 vdd.n162 vdd.n161 75.1835
R17076 vdd.n160 vdd.n159 75.1835
R17077 vdd.n75 vdd.n74 75.1835
R17078 vdd.n73 vdd.n72 75.1835
R17079 vdd.n71 vdd.n70 75.1835
R17080 vdd.n1112 vdd.n1111 75.1835
R17081 vdd.n1114 vdd.n1113 75.1835
R17082 vdd.n1116 vdd.n1115 75.1835
R17083 vdd.n1022 vdd.n1021 75.1835
R17084 vdd.n1024 vdd.n1023 75.1835
R17085 vdd.n1026 vdd.n1025 75.1835
R17086 vdd.n933 vdd.n932 75.1835
R17087 vdd.n935 vdd.n934 75.1835
R17088 vdd.n937 vdd.n936 75.1835
R17089 vdd.n2472 vdd.n2471 72.8958
R17090 vdd.n2471 vdd.n2235 72.8958
R17091 vdd.n2471 vdd.n2236 72.8958
R17092 vdd.n2471 vdd.n2237 72.8958
R17093 vdd.n2471 vdd.n2238 72.8958
R17094 vdd.n2471 vdd.n2239 72.8958
R17095 vdd.n2471 vdd.n2240 72.8958
R17096 vdd.n2471 vdd.n2241 72.8958
R17097 vdd.n2471 vdd.n2242 72.8958
R17098 vdd.n2471 vdd.n2243 72.8958
R17099 vdd.n2471 vdd.n2244 72.8958
R17100 vdd.n2471 vdd.n2245 72.8958
R17101 vdd.n2471 vdd.n2246 72.8958
R17102 vdd.n2471 vdd.n2247 72.8958
R17103 vdd.n2471 vdd.n2248 72.8958
R17104 vdd.n2471 vdd.n2249 72.8958
R17105 vdd.n2471 vdd.n2250 72.8958
R17106 vdd.n593 vdd.n484 72.8958
R17107 vdd.n2680 vdd.n484 72.8958
R17108 vdd.n587 vdd.n484 72.8958
R17109 vdd.n2687 vdd.n484 72.8958
R17110 vdd.n584 vdd.n484 72.8958
R17111 vdd.n2694 vdd.n484 72.8958
R17112 vdd.n581 vdd.n484 72.8958
R17113 vdd.n2701 vdd.n484 72.8958
R17114 vdd.n2704 vdd.n484 72.8958
R17115 vdd.n2560 vdd.n484 72.8958
R17116 vdd.n2565 vdd.n484 72.8958
R17117 vdd.n2559 vdd.n484 72.8958
R17118 vdd.n2572 vdd.n484 72.8958
R17119 vdd.n2556 vdd.n484 72.8958
R17120 vdd.n2579 vdd.n484 72.8958
R17121 vdd.n2553 vdd.n484 72.8958
R17122 vdd.n2586 vdd.n484 72.8958
R17123 vdd.n1724 vdd.n839 72.8958
R17124 vdd.n1730 vdd.n839 72.8958
R17125 vdd.n1732 vdd.n839 72.8958
R17126 vdd.n1738 vdd.n839 72.8958
R17127 vdd.n1740 vdd.n839 72.8958
R17128 vdd.n1746 vdd.n839 72.8958
R17129 vdd.n1748 vdd.n839 72.8958
R17130 vdd.n1754 vdd.n839 72.8958
R17131 vdd.n1925 vdd.n839 72.8958
R17132 vdd.n1923 vdd.n839 72.8958
R17133 vdd.n1917 vdd.n839 72.8958
R17134 vdd.n1915 vdd.n839 72.8958
R17135 vdd.n1909 vdd.n839 72.8958
R17136 vdd.n1907 vdd.n839 72.8958
R17137 vdd.n1901 vdd.n839 72.8958
R17138 vdd.n1899 vdd.n839 72.8958
R17139 vdd.n1893 vdd.n839 72.8958
R17140 vdd.n2218 vdd.n727 72.8958
R17141 vdd.n2218 vdd.n728 72.8958
R17142 vdd.n2218 vdd.n729 72.8958
R17143 vdd.n2218 vdd.n730 72.8958
R17144 vdd.n2218 vdd.n731 72.8958
R17145 vdd.n2218 vdd.n732 72.8958
R17146 vdd.n2218 vdd.n733 72.8958
R17147 vdd.n2218 vdd.n734 72.8958
R17148 vdd.n2218 vdd.n735 72.8958
R17149 vdd.n2218 vdd.n736 72.8958
R17150 vdd.n2218 vdd.n737 72.8958
R17151 vdd.n2218 vdd.n738 72.8958
R17152 vdd.n2218 vdd.n739 72.8958
R17153 vdd.n2218 vdd.n740 72.8958
R17154 vdd.n2218 vdd.n741 72.8958
R17155 vdd.n2218 vdd.n742 72.8958
R17156 vdd.n2218 vdd.n743 72.8958
R17157 vdd.n2471 vdd.n2470 72.8958
R17158 vdd.n2471 vdd.n2219 72.8958
R17159 vdd.n2471 vdd.n2220 72.8958
R17160 vdd.n2471 vdd.n2221 72.8958
R17161 vdd.n2471 vdd.n2222 72.8958
R17162 vdd.n2471 vdd.n2223 72.8958
R17163 vdd.n2471 vdd.n2224 72.8958
R17164 vdd.n2471 vdd.n2225 72.8958
R17165 vdd.n2471 vdd.n2226 72.8958
R17166 vdd.n2471 vdd.n2227 72.8958
R17167 vdd.n2471 vdd.n2228 72.8958
R17168 vdd.n2471 vdd.n2229 72.8958
R17169 vdd.n2471 vdd.n2230 72.8958
R17170 vdd.n2471 vdd.n2231 72.8958
R17171 vdd.n2471 vdd.n2232 72.8958
R17172 vdd.n2471 vdd.n2233 72.8958
R17173 vdd.n2471 vdd.n2234 72.8958
R17174 vdd.n2610 vdd.n484 72.8958
R17175 vdd.n625 vdd.n484 72.8958
R17176 vdd.n2618 vdd.n484 72.8958
R17177 vdd.n620 vdd.n484 72.8958
R17178 vdd.n2625 vdd.n484 72.8958
R17179 vdd.n617 vdd.n484 72.8958
R17180 vdd.n2632 vdd.n484 72.8958
R17181 vdd.n614 vdd.n484 72.8958
R17182 vdd.n2639 vdd.n484 72.8958
R17183 vdd.n2643 vdd.n484 72.8958
R17184 vdd.n611 vdd.n484 72.8958
R17185 vdd.n2650 vdd.n484 72.8958
R17186 vdd.n608 vdd.n484 72.8958
R17187 vdd.n2657 vdd.n484 72.8958
R17188 vdd.n605 vdd.n484 72.8958
R17189 vdd.n2664 vdd.n484 72.8958
R17190 vdd.n2667 vdd.n484 72.8958
R17191 vdd.n2218 vdd.n725 72.8958
R17192 vdd.n2218 vdd.n724 72.8958
R17193 vdd.n2218 vdd.n723 72.8958
R17194 vdd.n2218 vdd.n722 72.8958
R17195 vdd.n2218 vdd.n721 72.8958
R17196 vdd.n2218 vdd.n720 72.8958
R17197 vdd.n2218 vdd.n719 72.8958
R17198 vdd.n2218 vdd.n718 72.8958
R17199 vdd.n2218 vdd.n717 72.8958
R17200 vdd.n2218 vdd.n716 72.8958
R17201 vdd.n2218 vdd.n715 72.8958
R17202 vdd.n2218 vdd.n714 72.8958
R17203 vdd.n2218 vdd.n713 72.8958
R17204 vdd.n2218 vdd.n712 72.8958
R17205 vdd.n2218 vdd.n711 72.8958
R17206 vdd.n2218 vdd.n710 72.8958
R17207 vdd.n2218 vdd.n709 72.8958
R17208 vdd.n1983 vdd.n839 72.8958
R17209 vdd.n1981 vdd.n839 72.8958
R17210 vdd.n1975 vdd.n839 72.8958
R17211 vdd.n1973 vdd.n839 72.8958
R17212 vdd.n1967 vdd.n839 72.8958
R17213 vdd.n1965 vdd.n839 72.8958
R17214 vdd.n1959 vdd.n839 72.8958
R17215 vdd.n1957 vdd.n839 72.8958
R17216 vdd.n851 vdd.n839 72.8958
R17217 vdd.n1799 vdd.n839 72.8958
R17218 vdd.n1804 vdd.n839 72.8958
R17219 vdd.n1806 vdd.n839 72.8958
R17220 vdd.n1812 vdd.n839 72.8958
R17221 vdd.n1814 vdd.n839 72.8958
R17222 vdd.n1820 vdd.n839 72.8958
R17223 vdd.n1822 vdd.n839 72.8958
R17224 vdd.n1829 vdd.n839 72.8958
R17225 vdd.n1422 vdd.n1421 66.2847
R17226 vdd.n1421 vdd.n1197 66.2847
R17227 vdd.n1421 vdd.n1198 66.2847
R17228 vdd.n1421 vdd.n1199 66.2847
R17229 vdd.n1421 vdd.n1200 66.2847
R17230 vdd.n1421 vdd.n1201 66.2847
R17231 vdd.n1421 vdd.n1202 66.2847
R17232 vdd.n1421 vdd.n1203 66.2847
R17233 vdd.n1421 vdd.n1204 66.2847
R17234 vdd.n1421 vdd.n1205 66.2847
R17235 vdd.n1421 vdd.n1206 66.2847
R17236 vdd.n1421 vdd.n1207 66.2847
R17237 vdd.n1421 vdd.n1208 66.2847
R17238 vdd.n1421 vdd.n1209 66.2847
R17239 vdd.n1421 vdd.n1210 66.2847
R17240 vdd.n1421 vdd.n1211 66.2847
R17241 vdd.n1421 vdd.n1212 66.2847
R17242 vdd.n1421 vdd.n1213 66.2847
R17243 vdd.n1421 vdd.n1214 66.2847
R17244 vdd.n1421 vdd.n1215 66.2847
R17245 vdd.n1421 vdd.n1216 66.2847
R17246 vdd.n1421 vdd.n1217 66.2847
R17247 vdd.n1421 vdd.n1218 66.2847
R17248 vdd.n1421 vdd.n1219 66.2847
R17249 vdd.n1421 vdd.n1220 66.2847
R17250 vdd.n1421 vdd.n1221 66.2847
R17251 vdd.n1421 vdd.n1222 66.2847
R17252 vdd.n1421 vdd.n1223 66.2847
R17253 vdd.n1421 vdd.n1224 66.2847
R17254 vdd.n1421 vdd.n1225 66.2847
R17255 vdd.n1421 vdd.n1226 66.2847
R17256 vdd.n863 vdd.n860 66.2847
R17257 vdd.n1614 vdd.n863 66.2847
R17258 vdd.n1619 vdd.n863 66.2847
R17259 vdd.n1624 vdd.n863 66.2847
R17260 vdd.n1612 vdd.n863 66.2847
R17261 vdd.n1631 vdd.n863 66.2847
R17262 vdd.n1604 vdd.n863 66.2847
R17263 vdd.n1638 vdd.n863 66.2847
R17264 vdd.n1597 vdd.n863 66.2847
R17265 vdd.n1645 vdd.n863 66.2847
R17266 vdd.n1591 vdd.n863 66.2847
R17267 vdd.n1586 vdd.n863 66.2847
R17268 vdd.n1656 vdd.n863 66.2847
R17269 vdd.n1578 vdd.n863 66.2847
R17270 vdd.n1663 vdd.n863 66.2847
R17271 vdd.n1571 vdd.n863 66.2847
R17272 vdd.n1670 vdd.n863 66.2847
R17273 vdd.n1564 vdd.n863 66.2847
R17274 vdd.n1677 vdd.n863 66.2847
R17275 vdd.n1557 vdd.n863 66.2847
R17276 vdd.n1684 vdd.n863 66.2847
R17277 vdd.n1551 vdd.n863 66.2847
R17278 vdd.n1546 vdd.n863 66.2847
R17279 vdd.n1695 vdd.n863 66.2847
R17280 vdd.n1538 vdd.n863 66.2847
R17281 vdd.n1702 vdd.n863 66.2847
R17282 vdd.n1531 vdd.n863 66.2847
R17283 vdd.n1709 vdd.n863 66.2847
R17284 vdd.n1712 vdd.n863 66.2847
R17285 vdd.n1522 vdd.n863 66.2847
R17286 vdd.n1934 vdd.n863 66.2847
R17287 vdd.n1516 vdd.n863 66.2847
R17288 vdd.n2841 vdd.n2840 66.2847
R17289 vdd.n2840 vdd.n485 66.2847
R17290 vdd.n2840 vdd.n486 66.2847
R17291 vdd.n2840 vdd.n487 66.2847
R17292 vdd.n2840 vdd.n488 66.2847
R17293 vdd.n2840 vdd.n489 66.2847
R17294 vdd.n2840 vdd.n490 66.2847
R17295 vdd.n2840 vdd.n491 66.2847
R17296 vdd.n2840 vdd.n492 66.2847
R17297 vdd.n2840 vdd.n493 66.2847
R17298 vdd.n2840 vdd.n494 66.2847
R17299 vdd.n2840 vdd.n495 66.2847
R17300 vdd.n2840 vdd.n496 66.2847
R17301 vdd.n2840 vdd.n497 66.2847
R17302 vdd.n2840 vdd.n498 66.2847
R17303 vdd.n2840 vdd.n499 66.2847
R17304 vdd.n2840 vdd.n500 66.2847
R17305 vdd.n2840 vdd.n501 66.2847
R17306 vdd.n2840 vdd.n502 66.2847
R17307 vdd.n2840 vdd.n503 66.2847
R17308 vdd.n2840 vdd.n504 66.2847
R17309 vdd.n2840 vdd.n505 66.2847
R17310 vdd.n2840 vdd.n506 66.2847
R17311 vdd.n2840 vdd.n507 66.2847
R17312 vdd.n2840 vdd.n508 66.2847
R17313 vdd.n2840 vdd.n509 66.2847
R17314 vdd.n2840 vdd.n510 66.2847
R17315 vdd.n2840 vdd.n511 66.2847
R17316 vdd.n2840 vdd.n512 66.2847
R17317 vdd.n2840 vdd.n513 66.2847
R17318 vdd.n2840 vdd.n514 66.2847
R17319 vdd.n2905 vdd.n329 66.2847
R17320 vdd.n2914 vdd.n329 66.2847
R17321 vdd.n439 vdd.n329 66.2847
R17322 vdd.n2921 vdd.n329 66.2847
R17323 vdd.n432 vdd.n329 66.2847
R17324 vdd.n2928 vdd.n329 66.2847
R17325 vdd.n425 vdd.n329 66.2847
R17326 vdd.n2935 vdd.n329 66.2847
R17327 vdd.n418 vdd.n329 66.2847
R17328 vdd.n2942 vdd.n329 66.2847
R17329 vdd.n412 vdd.n329 66.2847
R17330 vdd.n407 vdd.n329 66.2847
R17331 vdd.n2953 vdd.n329 66.2847
R17332 vdd.n399 vdd.n329 66.2847
R17333 vdd.n2960 vdd.n329 66.2847
R17334 vdd.n392 vdd.n329 66.2847
R17335 vdd.n2967 vdd.n329 66.2847
R17336 vdd.n385 vdd.n329 66.2847
R17337 vdd.n2974 vdd.n329 66.2847
R17338 vdd.n378 vdd.n329 66.2847
R17339 vdd.n2981 vdd.n329 66.2847
R17340 vdd.n372 vdd.n329 66.2847
R17341 vdd.n367 vdd.n329 66.2847
R17342 vdd.n2992 vdd.n329 66.2847
R17343 vdd.n359 vdd.n329 66.2847
R17344 vdd.n2999 vdd.n329 66.2847
R17345 vdd.n352 vdd.n329 66.2847
R17346 vdd.n3006 vdd.n329 66.2847
R17347 vdd.n345 vdd.n329 66.2847
R17348 vdd.n3013 vdd.n329 66.2847
R17349 vdd.n3016 vdd.n329 66.2847
R17350 vdd.n333 vdd.n329 66.2847
R17351 vdd.n334 vdd.n333 52.4337
R17352 vdd.n3016 vdd.n3015 52.4337
R17353 vdd.n3013 vdd.n3012 52.4337
R17354 vdd.n3008 vdd.n345 52.4337
R17355 vdd.n3006 vdd.n3005 52.4337
R17356 vdd.n3001 vdd.n352 52.4337
R17357 vdd.n2999 vdd.n2998 52.4337
R17358 vdd.n2994 vdd.n359 52.4337
R17359 vdd.n2992 vdd.n2991 52.4337
R17360 vdd.n368 vdd.n367 52.4337
R17361 vdd.n2983 vdd.n372 52.4337
R17362 vdd.n2981 vdd.n2980 52.4337
R17363 vdd.n2976 vdd.n378 52.4337
R17364 vdd.n2974 vdd.n2973 52.4337
R17365 vdd.n2969 vdd.n385 52.4337
R17366 vdd.n2967 vdd.n2966 52.4337
R17367 vdd.n2962 vdd.n392 52.4337
R17368 vdd.n2960 vdd.n2959 52.4337
R17369 vdd.n2955 vdd.n399 52.4337
R17370 vdd.n2953 vdd.n2952 52.4337
R17371 vdd.n408 vdd.n407 52.4337
R17372 vdd.n2944 vdd.n412 52.4337
R17373 vdd.n2942 vdd.n2941 52.4337
R17374 vdd.n2937 vdd.n418 52.4337
R17375 vdd.n2935 vdd.n2934 52.4337
R17376 vdd.n2930 vdd.n425 52.4337
R17377 vdd.n2928 vdd.n2927 52.4337
R17378 vdd.n2923 vdd.n432 52.4337
R17379 vdd.n2921 vdd.n2920 52.4337
R17380 vdd.n2916 vdd.n439 52.4337
R17381 vdd.n2914 vdd.n2913 52.4337
R17382 vdd.n2906 vdd.n2905 52.4337
R17383 vdd.n2842 vdd.n2841 52.4337
R17384 vdd.n517 vdd.n485 52.4337
R17385 vdd.n523 vdd.n486 52.4337
R17386 vdd.n2831 vdd.n487 52.4337
R17387 vdd.n2827 vdd.n488 52.4337
R17388 vdd.n2823 vdd.n489 52.4337
R17389 vdd.n2819 vdd.n490 52.4337
R17390 vdd.n2815 vdd.n491 52.4337
R17391 vdd.n2811 vdd.n492 52.4337
R17392 vdd.n2807 vdd.n493 52.4337
R17393 vdd.n2799 vdd.n494 52.4337
R17394 vdd.n2795 vdd.n495 52.4337
R17395 vdd.n2791 vdd.n496 52.4337
R17396 vdd.n2787 vdd.n497 52.4337
R17397 vdd.n2783 vdd.n498 52.4337
R17398 vdd.n2779 vdd.n499 52.4337
R17399 vdd.n2775 vdd.n500 52.4337
R17400 vdd.n2771 vdd.n501 52.4337
R17401 vdd.n2767 vdd.n502 52.4337
R17402 vdd.n2763 vdd.n503 52.4337
R17403 vdd.n2759 vdd.n504 52.4337
R17404 vdd.n2753 vdd.n505 52.4337
R17405 vdd.n2749 vdd.n506 52.4337
R17406 vdd.n2745 vdd.n507 52.4337
R17407 vdd.n2741 vdd.n508 52.4337
R17408 vdd.n2737 vdd.n509 52.4337
R17409 vdd.n2733 vdd.n510 52.4337
R17410 vdd.n2729 vdd.n511 52.4337
R17411 vdd.n2725 vdd.n512 52.4337
R17412 vdd.n2721 vdd.n513 52.4337
R17413 vdd.n2717 vdd.n514 52.4337
R17414 vdd.n1936 vdd.n1516 52.4337
R17415 vdd.n1934 vdd.n1933 52.4337
R17416 vdd.n1523 vdd.n1522 52.4337
R17417 vdd.n1712 vdd.n1711 52.4337
R17418 vdd.n1709 vdd.n1708 52.4337
R17419 vdd.n1704 vdd.n1531 52.4337
R17420 vdd.n1702 vdd.n1701 52.4337
R17421 vdd.n1697 vdd.n1538 52.4337
R17422 vdd.n1695 vdd.n1694 52.4337
R17423 vdd.n1547 vdd.n1546 52.4337
R17424 vdd.n1686 vdd.n1551 52.4337
R17425 vdd.n1684 vdd.n1683 52.4337
R17426 vdd.n1679 vdd.n1557 52.4337
R17427 vdd.n1677 vdd.n1676 52.4337
R17428 vdd.n1672 vdd.n1564 52.4337
R17429 vdd.n1670 vdd.n1669 52.4337
R17430 vdd.n1665 vdd.n1571 52.4337
R17431 vdd.n1663 vdd.n1662 52.4337
R17432 vdd.n1658 vdd.n1578 52.4337
R17433 vdd.n1656 vdd.n1655 52.4337
R17434 vdd.n1587 vdd.n1586 52.4337
R17435 vdd.n1647 vdd.n1591 52.4337
R17436 vdd.n1645 vdd.n1644 52.4337
R17437 vdd.n1640 vdd.n1597 52.4337
R17438 vdd.n1638 vdd.n1637 52.4337
R17439 vdd.n1633 vdd.n1604 52.4337
R17440 vdd.n1631 vdd.n1630 52.4337
R17441 vdd.n1626 vdd.n1612 52.4337
R17442 vdd.n1624 vdd.n1623 52.4337
R17443 vdd.n1619 vdd.n1618 52.4337
R17444 vdd.n1614 vdd.n1613 52.4337
R17445 vdd.n1945 vdd.n860 52.4337
R17446 vdd.n1423 vdd.n1422 52.4337
R17447 vdd.n1229 vdd.n1197 52.4337
R17448 vdd.n1233 vdd.n1198 52.4337
R17449 vdd.n1235 vdd.n1199 52.4337
R17450 vdd.n1239 vdd.n1200 52.4337
R17451 vdd.n1241 vdd.n1201 52.4337
R17452 vdd.n1245 vdd.n1202 52.4337
R17453 vdd.n1247 vdd.n1203 52.4337
R17454 vdd.n1251 vdd.n1204 52.4337
R17455 vdd.n1253 vdd.n1205 52.4337
R17456 vdd.n1259 vdd.n1206 52.4337
R17457 vdd.n1261 vdd.n1207 52.4337
R17458 vdd.n1265 vdd.n1208 52.4337
R17459 vdd.n1267 vdd.n1209 52.4337
R17460 vdd.n1271 vdd.n1210 52.4337
R17461 vdd.n1273 vdd.n1211 52.4337
R17462 vdd.n1277 vdd.n1212 52.4337
R17463 vdd.n1279 vdd.n1213 52.4337
R17464 vdd.n1283 vdd.n1214 52.4337
R17465 vdd.n1285 vdd.n1215 52.4337
R17466 vdd.n1357 vdd.n1216 52.4337
R17467 vdd.n1290 vdd.n1217 52.4337
R17468 vdd.n1294 vdd.n1218 52.4337
R17469 vdd.n1296 vdd.n1219 52.4337
R17470 vdd.n1300 vdd.n1220 52.4337
R17471 vdd.n1302 vdd.n1221 52.4337
R17472 vdd.n1306 vdd.n1222 52.4337
R17473 vdd.n1308 vdd.n1223 52.4337
R17474 vdd.n1312 vdd.n1224 52.4337
R17475 vdd.n1314 vdd.n1225 52.4337
R17476 vdd.n1318 vdd.n1226 52.4337
R17477 vdd.n1422 vdd.n1196 52.4337
R17478 vdd.n1232 vdd.n1197 52.4337
R17479 vdd.n1234 vdd.n1198 52.4337
R17480 vdd.n1238 vdd.n1199 52.4337
R17481 vdd.n1240 vdd.n1200 52.4337
R17482 vdd.n1244 vdd.n1201 52.4337
R17483 vdd.n1246 vdd.n1202 52.4337
R17484 vdd.n1250 vdd.n1203 52.4337
R17485 vdd.n1252 vdd.n1204 52.4337
R17486 vdd.n1258 vdd.n1205 52.4337
R17487 vdd.n1260 vdd.n1206 52.4337
R17488 vdd.n1264 vdd.n1207 52.4337
R17489 vdd.n1266 vdd.n1208 52.4337
R17490 vdd.n1270 vdd.n1209 52.4337
R17491 vdd.n1272 vdd.n1210 52.4337
R17492 vdd.n1276 vdd.n1211 52.4337
R17493 vdd.n1278 vdd.n1212 52.4337
R17494 vdd.n1282 vdd.n1213 52.4337
R17495 vdd.n1284 vdd.n1214 52.4337
R17496 vdd.n1288 vdd.n1215 52.4337
R17497 vdd.n1289 vdd.n1216 52.4337
R17498 vdd.n1293 vdd.n1217 52.4337
R17499 vdd.n1295 vdd.n1218 52.4337
R17500 vdd.n1299 vdd.n1219 52.4337
R17501 vdd.n1301 vdd.n1220 52.4337
R17502 vdd.n1305 vdd.n1221 52.4337
R17503 vdd.n1307 vdd.n1222 52.4337
R17504 vdd.n1311 vdd.n1223 52.4337
R17505 vdd.n1313 vdd.n1224 52.4337
R17506 vdd.n1317 vdd.n1225 52.4337
R17507 vdd.n1319 vdd.n1226 52.4337
R17508 vdd.n860 vdd.n859 52.4337
R17509 vdd.n1615 vdd.n1614 52.4337
R17510 vdd.n1620 vdd.n1619 52.4337
R17511 vdd.n1625 vdd.n1624 52.4337
R17512 vdd.n1612 vdd.n1605 52.4337
R17513 vdd.n1632 vdd.n1631 52.4337
R17514 vdd.n1604 vdd.n1598 52.4337
R17515 vdd.n1639 vdd.n1638 52.4337
R17516 vdd.n1597 vdd.n1592 52.4337
R17517 vdd.n1646 vdd.n1645 52.4337
R17518 vdd.n1591 vdd.n1590 52.4337
R17519 vdd.n1586 vdd.n1579 52.4337
R17520 vdd.n1657 vdd.n1656 52.4337
R17521 vdd.n1578 vdd.n1572 52.4337
R17522 vdd.n1664 vdd.n1663 52.4337
R17523 vdd.n1571 vdd.n1565 52.4337
R17524 vdd.n1671 vdd.n1670 52.4337
R17525 vdd.n1564 vdd.n1558 52.4337
R17526 vdd.n1678 vdd.n1677 52.4337
R17527 vdd.n1557 vdd.n1552 52.4337
R17528 vdd.n1685 vdd.n1684 52.4337
R17529 vdd.n1551 vdd.n1550 52.4337
R17530 vdd.n1546 vdd.n1539 52.4337
R17531 vdd.n1696 vdd.n1695 52.4337
R17532 vdd.n1538 vdd.n1532 52.4337
R17533 vdd.n1703 vdd.n1702 52.4337
R17534 vdd.n1531 vdd.n1525 52.4337
R17535 vdd.n1710 vdd.n1709 52.4337
R17536 vdd.n1713 vdd.n1712 52.4337
R17537 vdd.n1522 vdd.n1517 52.4337
R17538 vdd.n1935 vdd.n1934 52.4337
R17539 vdd.n1516 vdd.n865 52.4337
R17540 vdd.n2841 vdd.n483 52.4337
R17541 vdd.n522 vdd.n485 52.4337
R17542 vdd.n2832 vdd.n486 52.4337
R17543 vdd.n2828 vdd.n487 52.4337
R17544 vdd.n2824 vdd.n488 52.4337
R17545 vdd.n2820 vdd.n489 52.4337
R17546 vdd.n2816 vdd.n490 52.4337
R17547 vdd.n2812 vdd.n491 52.4337
R17548 vdd.n2808 vdd.n492 52.4337
R17549 vdd.n2798 vdd.n493 52.4337
R17550 vdd.n2796 vdd.n494 52.4337
R17551 vdd.n2792 vdd.n495 52.4337
R17552 vdd.n2788 vdd.n496 52.4337
R17553 vdd.n2784 vdd.n497 52.4337
R17554 vdd.n2780 vdd.n498 52.4337
R17555 vdd.n2776 vdd.n499 52.4337
R17556 vdd.n2772 vdd.n500 52.4337
R17557 vdd.n2768 vdd.n501 52.4337
R17558 vdd.n2764 vdd.n502 52.4337
R17559 vdd.n2760 vdd.n503 52.4337
R17560 vdd.n2752 vdd.n504 52.4337
R17561 vdd.n2750 vdd.n505 52.4337
R17562 vdd.n2746 vdd.n506 52.4337
R17563 vdd.n2742 vdd.n507 52.4337
R17564 vdd.n2738 vdd.n508 52.4337
R17565 vdd.n2734 vdd.n509 52.4337
R17566 vdd.n2730 vdd.n510 52.4337
R17567 vdd.n2726 vdd.n511 52.4337
R17568 vdd.n2722 vdd.n512 52.4337
R17569 vdd.n2718 vdd.n513 52.4337
R17570 vdd.n2714 vdd.n514 52.4337
R17571 vdd.n2905 vdd.n440 52.4337
R17572 vdd.n2915 vdd.n2914 52.4337
R17573 vdd.n439 vdd.n433 52.4337
R17574 vdd.n2922 vdd.n2921 52.4337
R17575 vdd.n432 vdd.n426 52.4337
R17576 vdd.n2929 vdd.n2928 52.4337
R17577 vdd.n425 vdd.n419 52.4337
R17578 vdd.n2936 vdd.n2935 52.4337
R17579 vdd.n418 vdd.n413 52.4337
R17580 vdd.n2943 vdd.n2942 52.4337
R17581 vdd.n412 vdd.n411 52.4337
R17582 vdd.n407 vdd.n400 52.4337
R17583 vdd.n2954 vdd.n2953 52.4337
R17584 vdd.n399 vdd.n393 52.4337
R17585 vdd.n2961 vdd.n2960 52.4337
R17586 vdd.n392 vdd.n386 52.4337
R17587 vdd.n2968 vdd.n2967 52.4337
R17588 vdd.n385 vdd.n379 52.4337
R17589 vdd.n2975 vdd.n2974 52.4337
R17590 vdd.n378 vdd.n373 52.4337
R17591 vdd.n2982 vdd.n2981 52.4337
R17592 vdd.n372 vdd.n371 52.4337
R17593 vdd.n367 vdd.n360 52.4337
R17594 vdd.n2993 vdd.n2992 52.4337
R17595 vdd.n359 vdd.n353 52.4337
R17596 vdd.n3000 vdd.n2999 52.4337
R17597 vdd.n352 vdd.n346 52.4337
R17598 vdd.n3007 vdd.n3006 52.4337
R17599 vdd.n345 vdd.n338 52.4337
R17600 vdd.n3014 vdd.n3013 52.4337
R17601 vdd.n3017 vdd.n3016 52.4337
R17602 vdd.n333 vdd.n330 52.4337
R17603 vdd.t38 vdd.t36 51.4683
R17604 vdd.n250 vdd.n248 42.0461
R17605 vdd.n160 vdd.n158 42.0461
R17606 vdd.n71 vdd.n69 42.0461
R17607 vdd.n1112 vdd.n1110 42.0461
R17608 vdd.n1022 vdd.n1020 42.0461
R17609 vdd.n933 vdd.n931 42.0461
R17610 vdd.n296 vdd.n295 41.6884
R17611 vdd.n206 vdd.n205 41.6884
R17612 vdd.n117 vdd.n116 41.6884
R17613 vdd.n1158 vdd.n1157 41.6884
R17614 vdd.n1068 vdd.n1067 41.6884
R17615 vdd.n979 vdd.n978 41.6884
R17616 vdd.n1322 vdd.n1321 41.1157
R17617 vdd.n1360 vdd.n1359 41.1157
R17618 vdd.n1256 vdd.n1255 41.1157
R17619 vdd.n2910 vdd.n2909 41.1157
R17620 vdd.n2949 vdd.n406 41.1157
R17621 vdd.n2988 vdd.n366 41.1157
R17622 vdd.n2667 vdd.n2666 39.2114
R17623 vdd.n2664 vdd.n2663 39.2114
R17624 vdd.n2659 vdd.n605 39.2114
R17625 vdd.n2657 vdd.n2656 39.2114
R17626 vdd.n2652 vdd.n608 39.2114
R17627 vdd.n2650 vdd.n2649 39.2114
R17628 vdd.n2645 vdd.n611 39.2114
R17629 vdd.n2643 vdd.n2642 39.2114
R17630 vdd.n2639 vdd.n2638 39.2114
R17631 vdd.n2634 vdd.n614 39.2114
R17632 vdd.n2632 vdd.n2631 39.2114
R17633 vdd.n2627 vdd.n617 39.2114
R17634 vdd.n2625 vdd.n2624 39.2114
R17635 vdd.n2620 vdd.n620 39.2114
R17636 vdd.n2618 vdd.n2617 39.2114
R17637 vdd.n2612 vdd.n625 39.2114
R17638 vdd.n2610 vdd.n2609 39.2114
R17639 vdd.n2470 vdd.n703 39.2114
R17640 vdd.n2465 vdd.n2219 39.2114
R17641 vdd.n2462 vdd.n2220 39.2114
R17642 vdd.n2458 vdd.n2221 39.2114
R17643 vdd.n2454 vdd.n2222 39.2114
R17644 vdd.n2450 vdd.n2223 39.2114
R17645 vdd.n2446 vdd.n2224 39.2114
R17646 vdd.n2442 vdd.n2225 39.2114
R17647 vdd.n2438 vdd.n2226 39.2114
R17648 vdd.n2434 vdd.n2227 39.2114
R17649 vdd.n2430 vdd.n2228 39.2114
R17650 vdd.n2426 vdd.n2229 39.2114
R17651 vdd.n2422 vdd.n2230 39.2114
R17652 vdd.n2418 vdd.n2231 39.2114
R17653 vdd.n2414 vdd.n2232 39.2114
R17654 vdd.n2410 vdd.n2233 39.2114
R17655 vdd.n2405 vdd.n2234 39.2114
R17656 vdd.n2213 vdd.n743 39.2114
R17657 vdd.n2209 vdd.n742 39.2114
R17658 vdd.n2205 vdd.n741 39.2114
R17659 vdd.n2201 vdd.n740 39.2114
R17660 vdd.n2197 vdd.n739 39.2114
R17661 vdd.n2193 vdd.n738 39.2114
R17662 vdd.n2189 vdd.n737 39.2114
R17663 vdd.n2185 vdd.n736 39.2114
R17664 vdd.n2181 vdd.n735 39.2114
R17665 vdd.n2177 vdd.n734 39.2114
R17666 vdd.n2173 vdd.n733 39.2114
R17667 vdd.n2169 vdd.n732 39.2114
R17668 vdd.n2165 vdd.n731 39.2114
R17669 vdd.n2161 vdd.n730 39.2114
R17670 vdd.n2157 vdd.n729 39.2114
R17671 vdd.n2152 vdd.n728 39.2114
R17672 vdd.n2148 vdd.n727 39.2114
R17673 vdd.n1724 vdd.n838 39.2114
R17674 vdd.n1730 vdd.n1729 39.2114
R17675 vdd.n1733 vdd.n1732 39.2114
R17676 vdd.n1738 vdd.n1737 39.2114
R17677 vdd.n1741 vdd.n1740 39.2114
R17678 vdd.n1746 vdd.n1745 39.2114
R17679 vdd.n1749 vdd.n1748 39.2114
R17680 vdd.n1754 vdd.n1753 39.2114
R17681 vdd.n1925 vdd.n1756 39.2114
R17682 vdd.n1924 vdd.n1923 39.2114
R17683 vdd.n1917 vdd.n1758 39.2114
R17684 vdd.n1916 vdd.n1915 39.2114
R17685 vdd.n1909 vdd.n1760 39.2114
R17686 vdd.n1908 vdd.n1907 39.2114
R17687 vdd.n1901 vdd.n1762 39.2114
R17688 vdd.n1900 vdd.n1899 39.2114
R17689 vdd.n1893 vdd.n1764 39.2114
R17690 vdd.n2586 vdd.n2585 39.2114
R17691 vdd.n2581 vdd.n2553 39.2114
R17692 vdd.n2579 vdd.n2578 39.2114
R17693 vdd.n2574 vdd.n2556 39.2114
R17694 vdd.n2572 vdd.n2571 39.2114
R17695 vdd.n2567 vdd.n2559 39.2114
R17696 vdd.n2565 vdd.n2564 39.2114
R17697 vdd.n2560 vdd.n577 39.2114
R17698 vdd.n2704 vdd.n2703 39.2114
R17699 vdd.n2701 vdd.n2700 39.2114
R17700 vdd.n2696 vdd.n581 39.2114
R17701 vdd.n2694 vdd.n2693 39.2114
R17702 vdd.n2689 vdd.n584 39.2114
R17703 vdd.n2687 vdd.n2686 39.2114
R17704 vdd.n2682 vdd.n587 39.2114
R17705 vdd.n2680 vdd.n2679 39.2114
R17706 vdd.n2675 vdd.n593 39.2114
R17707 vdd.n2472 vdd.n706 39.2114
R17708 vdd.n2235 vdd.n708 39.2114
R17709 vdd.n2261 vdd.n2236 39.2114
R17710 vdd.n2265 vdd.n2237 39.2114
R17711 vdd.n2269 vdd.n2238 39.2114
R17712 vdd.n2273 vdd.n2239 39.2114
R17713 vdd.n2277 vdd.n2240 39.2114
R17714 vdd.n2281 vdd.n2241 39.2114
R17715 vdd.n2285 vdd.n2242 39.2114
R17716 vdd.n2289 vdd.n2243 39.2114
R17717 vdd.n2293 vdd.n2244 39.2114
R17718 vdd.n2297 vdd.n2245 39.2114
R17719 vdd.n2301 vdd.n2246 39.2114
R17720 vdd.n2305 vdd.n2247 39.2114
R17721 vdd.n2309 vdd.n2248 39.2114
R17722 vdd.n2313 vdd.n2249 39.2114
R17723 vdd.n2317 vdd.n2250 39.2114
R17724 vdd.n2473 vdd.n2472 39.2114
R17725 vdd.n2260 vdd.n2235 39.2114
R17726 vdd.n2264 vdd.n2236 39.2114
R17727 vdd.n2268 vdd.n2237 39.2114
R17728 vdd.n2272 vdd.n2238 39.2114
R17729 vdd.n2276 vdd.n2239 39.2114
R17730 vdd.n2280 vdd.n2240 39.2114
R17731 vdd.n2284 vdd.n2241 39.2114
R17732 vdd.n2288 vdd.n2242 39.2114
R17733 vdd.n2292 vdd.n2243 39.2114
R17734 vdd.n2296 vdd.n2244 39.2114
R17735 vdd.n2300 vdd.n2245 39.2114
R17736 vdd.n2304 vdd.n2246 39.2114
R17737 vdd.n2308 vdd.n2247 39.2114
R17738 vdd.n2312 vdd.n2248 39.2114
R17739 vdd.n2316 vdd.n2249 39.2114
R17740 vdd.n2319 vdd.n2250 39.2114
R17741 vdd.n593 vdd.n588 39.2114
R17742 vdd.n2681 vdd.n2680 39.2114
R17743 vdd.n587 vdd.n585 39.2114
R17744 vdd.n2688 vdd.n2687 39.2114
R17745 vdd.n584 vdd.n582 39.2114
R17746 vdd.n2695 vdd.n2694 39.2114
R17747 vdd.n581 vdd.n579 39.2114
R17748 vdd.n2702 vdd.n2701 39.2114
R17749 vdd.n2705 vdd.n2704 39.2114
R17750 vdd.n2561 vdd.n2560 39.2114
R17751 vdd.n2566 vdd.n2565 39.2114
R17752 vdd.n2559 vdd.n2557 39.2114
R17753 vdd.n2573 vdd.n2572 39.2114
R17754 vdd.n2556 vdd.n2554 39.2114
R17755 vdd.n2580 vdd.n2579 39.2114
R17756 vdd.n2553 vdd.n2551 39.2114
R17757 vdd.n2587 vdd.n2586 39.2114
R17758 vdd.n1725 vdd.n1724 39.2114
R17759 vdd.n1731 vdd.n1730 39.2114
R17760 vdd.n1732 vdd.n1721 39.2114
R17761 vdd.n1739 vdd.n1738 39.2114
R17762 vdd.n1740 vdd.n1719 39.2114
R17763 vdd.n1747 vdd.n1746 39.2114
R17764 vdd.n1748 vdd.n1717 39.2114
R17765 vdd.n1755 vdd.n1754 39.2114
R17766 vdd.n1926 vdd.n1925 39.2114
R17767 vdd.n1923 vdd.n1922 39.2114
R17768 vdd.n1918 vdd.n1917 39.2114
R17769 vdd.n1915 vdd.n1914 39.2114
R17770 vdd.n1910 vdd.n1909 39.2114
R17771 vdd.n1907 vdd.n1906 39.2114
R17772 vdd.n1902 vdd.n1901 39.2114
R17773 vdd.n1899 vdd.n1898 39.2114
R17774 vdd.n1894 vdd.n1893 39.2114
R17775 vdd.n2151 vdd.n727 39.2114
R17776 vdd.n2156 vdd.n728 39.2114
R17777 vdd.n2160 vdd.n729 39.2114
R17778 vdd.n2164 vdd.n730 39.2114
R17779 vdd.n2168 vdd.n731 39.2114
R17780 vdd.n2172 vdd.n732 39.2114
R17781 vdd.n2176 vdd.n733 39.2114
R17782 vdd.n2180 vdd.n734 39.2114
R17783 vdd.n2184 vdd.n735 39.2114
R17784 vdd.n2188 vdd.n736 39.2114
R17785 vdd.n2192 vdd.n737 39.2114
R17786 vdd.n2196 vdd.n738 39.2114
R17787 vdd.n2200 vdd.n739 39.2114
R17788 vdd.n2204 vdd.n740 39.2114
R17789 vdd.n2208 vdd.n741 39.2114
R17790 vdd.n2212 vdd.n742 39.2114
R17791 vdd.n745 vdd.n743 39.2114
R17792 vdd.n2470 vdd.n2469 39.2114
R17793 vdd.n2463 vdd.n2219 39.2114
R17794 vdd.n2459 vdd.n2220 39.2114
R17795 vdd.n2455 vdd.n2221 39.2114
R17796 vdd.n2451 vdd.n2222 39.2114
R17797 vdd.n2447 vdd.n2223 39.2114
R17798 vdd.n2443 vdd.n2224 39.2114
R17799 vdd.n2439 vdd.n2225 39.2114
R17800 vdd.n2435 vdd.n2226 39.2114
R17801 vdd.n2431 vdd.n2227 39.2114
R17802 vdd.n2427 vdd.n2228 39.2114
R17803 vdd.n2423 vdd.n2229 39.2114
R17804 vdd.n2419 vdd.n2230 39.2114
R17805 vdd.n2415 vdd.n2231 39.2114
R17806 vdd.n2411 vdd.n2232 39.2114
R17807 vdd.n2406 vdd.n2233 39.2114
R17808 vdd.n2402 vdd.n2234 39.2114
R17809 vdd.n2611 vdd.n2610 39.2114
R17810 vdd.n625 vdd.n621 39.2114
R17811 vdd.n2619 vdd.n2618 39.2114
R17812 vdd.n620 vdd.n618 39.2114
R17813 vdd.n2626 vdd.n2625 39.2114
R17814 vdd.n617 vdd.n615 39.2114
R17815 vdd.n2633 vdd.n2632 39.2114
R17816 vdd.n614 vdd.n612 39.2114
R17817 vdd.n2640 vdd.n2639 39.2114
R17818 vdd.n2644 vdd.n2643 39.2114
R17819 vdd.n611 vdd.n609 39.2114
R17820 vdd.n2651 vdd.n2650 39.2114
R17821 vdd.n608 vdd.n606 39.2114
R17822 vdd.n2658 vdd.n2657 39.2114
R17823 vdd.n605 vdd.n603 39.2114
R17824 vdd.n2665 vdd.n2664 39.2114
R17825 vdd.n2668 vdd.n2667 39.2114
R17826 vdd.n753 vdd.n709 39.2114
R17827 vdd.n2140 vdd.n710 39.2114
R17828 vdd.n2136 vdd.n711 39.2114
R17829 vdd.n2132 vdd.n712 39.2114
R17830 vdd.n2128 vdd.n713 39.2114
R17831 vdd.n2124 vdd.n714 39.2114
R17832 vdd.n2120 vdd.n715 39.2114
R17833 vdd.n2116 vdd.n716 39.2114
R17834 vdd.n2112 vdd.n717 39.2114
R17835 vdd.n2108 vdd.n718 39.2114
R17836 vdd.n2104 vdd.n719 39.2114
R17837 vdd.n2100 vdd.n720 39.2114
R17838 vdd.n2096 vdd.n721 39.2114
R17839 vdd.n2092 vdd.n722 39.2114
R17840 vdd.n2088 vdd.n723 39.2114
R17841 vdd.n2084 vdd.n724 39.2114
R17842 vdd.n2080 vdd.n725 39.2114
R17843 vdd.n1983 vdd.n842 39.2114
R17844 vdd.n1982 vdd.n1981 39.2114
R17845 vdd.n1975 vdd.n844 39.2114
R17846 vdd.n1974 vdd.n1973 39.2114
R17847 vdd.n1967 vdd.n846 39.2114
R17848 vdd.n1966 vdd.n1965 39.2114
R17849 vdd.n1959 vdd.n848 39.2114
R17850 vdd.n1958 vdd.n1957 39.2114
R17851 vdd.n851 vdd.n850 39.2114
R17852 vdd.n1799 vdd.n1798 39.2114
R17853 vdd.n1804 vdd.n1803 39.2114
R17854 vdd.n1807 vdd.n1806 39.2114
R17855 vdd.n1812 vdd.n1811 39.2114
R17856 vdd.n1815 vdd.n1814 39.2114
R17857 vdd.n1820 vdd.n1819 39.2114
R17858 vdd.n1823 vdd.n1822 39.2114
R17859 vdd.n1829 vdd.n1828 39.2114
R17860 vdd.n2077 vdd.n725 39.2114
R17861 vdd.n2081 vdd.n724 39.2114
R17862 vdd.n2085 vdd.n723 39.2114
R17863 vdd.n2089 vdd.n722 39.2114
R17864 vdd.n2093 vdd.n721 39.2114
R17865 vdd.n2097 vdd.n720 39.2114
R17866 vdd.n2101 vdd.n719 39.2114
R17867 vdd.n2105 vdd.n718 39.2114
R17868 vdd.n2109 vdd.n717 39.2114
R17869 vdd.n2113 vdd.n716 39.2114
R17870 vdd.n2117 vdd.n715 39.2114
R17871 vdd.n2121 vdd.n714 39.2114
R17872 vdd.n2125 vdd.n713 39.2114
R17873 vdd.n2129 vdd.n712 39.2114
R17874 vdd.n2133 vdd.n711 39.2114
R17875 vdd.n2137 vdd.n710 39.2114
R17876 vdd.n2141 vdd.n709 39.2114
R17877 vdd.n1984 vdd.n1983 39.2114
R17878 vdd.n1981 vdd.n1980 39.2114
R17879 vdd.n1976 vdd.n1975 39.2114
R17880 vdd.n1973 vdd.n1972 39.2114
R17881 vdd.n1968 vdd.n1967 39.2114
R17882 vdd.n1965 vdd.n1964 39.2114
R17883 vdd.n1960 vdd.n1959 39.2114
R17884 vdd.n1957 vdd.n1956 39.2114
R17885 vdd.n852 vdd.n851 39.2114
R17886 vdd.n1800 vdd.n1799 39.2114
R17887 vdd.n1805 vdd.n1804 39.2114
R17888 vdd.n1806 vdd.n1796 39.2114
R17889 vdd.n1813 vdd.n1812 39.2114
R17890 vdd.n1814 vdd.n1794 39.2114
R17891 vdd.n1821 vdd.n1820 39.2114
R17892 vdd.n1822 vdd.n1790 39.2114
R17893 vdd.n1830 vdd.n1829 39.2114
R17894 vdd.n1949 vdd.n1948 37.2369
R17895 vdd.n1652 vdd.n1585 37.2369
R17896 vdd.n1691 vdd.n1545 37.2369
R17897 vdd.n2758 vdd.n558 37.2369
R17898 vdd.n2806 vdd.n2805 37.2369
R17899 vdd.n2713 vdd.n2712 37.2369
R17900 vdd.n1991 vdd.n837 31.6883
R17901 vdd.n2216 vdd.n746 31.6883
R17902 vdd.n2149 vdd.n749 31.6883
R17903 vdd.n1895 vdd.n1892 31.6883
R17904 vdd.n2403 vdd.n2401 31.6883
R17905 vdd.n2608 vdd.n2607 31.6883
R17906 vdd.n2480 vdd.n702 31.6883
R17907 vdd.n2671 vdd.n2670 31.6883
R17908 vdd.n2590 vdd.n2589 31.6883
R17909 vdd.n2676 vdd.n592 31.6883
R17910 vdd.n2322 vdd.n2321 31.6883
R17911 vdd.n2476 vdd.n2475 31.6883
R17912 vdd.n1987 vdd.n1986 31.6883
R17913 vdd.n2144 vdd.n2143 31.6883
R17914 vdd.n2076 vdd.n2075 31.6883
R17915 vdd.n1833 vdd.n1832 31.6883
R17916 vdd.n1826 vdd.n1792 30.449
R17917 vdd.n757 vdd.n756 30.449
R17918 vdd.n1767 vdd.n1766 30.449
R17919 vdd.n2154 vdd.n748 30.449
R17920 vdd.n2258 vdd.n2257 30.449
R17921 vdd.n2614 vdd.n623 30.449
R17922 vdd.n2408 vdd.n2254 30.449
R17923 vdd.n591 vdd.n590 30.449
R17924 vdd.n1421 vdd.n1228 22.6735
R17925 vdd.n1943 vdd.n863 22.6735
R17926 vdd.n2840 vdd.n516 22.6735
R17927 vdd.n3025 vdd.n329 22.6735
R17928 vdd.n1432 vdd.n1190 19.3944
R17929 vdd.n1432 vdd.n1188 19.3944
R17930 vdd.n1436 vdd.n1188 19.3944
R17931 vdd.n1436 vdd.n1178 19.3944
R17932 vdd.n1449 vdd.n1178 19.3944
R17933 vdd.n1449 vdd.n1176 19.3944
R17934 vdd.n1453 vdd.n1176 19.3944
R17935 vdd.n1453 vdd.n1168 19.3944
R17936 vdd.n1467 vdd.n1168 19.3944
R17937 vdd.n1467 vdd.n1166 19.3944
R17938 vdd.n1471 vdd.n1166 19.3944
R17939 vdd.n1471 vdd.n885 19.3944
R17940 vdd.n1483 vdd.n885 19.3944
R17941 vdd.n1483 vdd.n883 19.3944
R17942 vdd.n1487 vdd.n883 19.3944
R17943 vdd.n1487 vdd.n875 19.3944
R17944 vdd.n1500 vdd.n875 19.3944
R17945 vdd.n1500 vdd.n872 19.3944
R17946 vdd.n1506 vdd.n872 19.3944
R17947 vdd.n1506 vdd.n873 19.3944
R17948 vdd.n873 vdd.n862 19.3944
R17949 vdd.n1356 vdd.n1291 19.3944
R17950 vdd.n1352 vdd.n1291 19.3944
R17951 vdd.n1352 vdd.n1351 19.3944
R17952 vdd.n1351 vdd.n1350 19.3944
R17953 vdd.n1350 vdd.n1297 19.3944
R17954 vdd.n1346 vdd.n1297 19.3944
R17955 vdd.n1346 vdd.n1345 19.3944
R17956 vdd.n1345 vdd.n1344 19.3944
R17957 vdd.n1344 vdd.n1303 19.3944
R17958 vdd.n1340 vdd.n1303 19.3944
R17959 vdd.n1340 vdd.n1339 19.3944
R17960 vdd.n1339 vdd.n1338 19.3944
R17961 vdd.n1338 vdd.n1309 19.3944
R17962 vdd.n1334 vdd.n1309 19.3944
R17963 vdd.n1334 vdd.n1333 19.3944
R17964 vdd.n1333 vdd.n1332 19.3944
R17965 vdd.n1332 vdd.n1315 19.3944
R17966 vdd.n1328 vdd.n1315 19.3944
R17967 vdd.n1328 vdd.n1327 19.3944
R17968 vdd.n1327 vdd.n1326 19.3944
R17969 vdd.n1391 vdd.n1390 19.3944
R17970 vdd.n1390 vdd.n1389 19.3944
R17971 vdd.n1389 vdd.n1262 19.3944
R17972 vdd.n1385 vdd.n1262 19.3944
R17973 vdd.n1385 vdd.n1384 19.3944
R17974 vdd.n1384 vdd.n1383 19.3944
R17975 vdd.n1383 vdd.n1268 19.3944
R17976 vdd.n1379 vdd.n1268 19.3944
R17977 vdd.n1379 vdd.n1378 19.3944
R17978 vdd.n1378 vdd.n1377 19.3944
R17979 vdd.n1377 vdd.n1274 19.3944
R17980 vdd.n1373 vdd.n1274 19.3944
R17981 vdd.n1373 vdd.n1372 19.3944
R17982 vdd.n1372 vdd.n1371 19.3944
R17983 vdd.n1371 vdd.n1280 19.3944
R17984 vdd.n1367 vdd.n1280 19.3944
R17985 vdd.n1367 vdd.n1366 19.3944
R17986 vdd.n1366 vdd.n1365 19.3944
R17987 vdd.n1365 vdd.n1286 19.3944
R17988 vdd.n1361 vdd.n1286 19.3944
R17989 vdd.n1424 vdd.n1195 19.3944
R17990 vdd.n1419 vdd.n1195 19.3944
R17991 vdd.n1419 vdd.n1230 19.3944
R17992 vdd.n1415 vdd.n1230 19.3944
R17993 vdd.n1415 vdd.n1414 19.3944
R17994 vdd.n1414 vdd.n1413 19.3944
R17995 vdd.n1413 vdd.n1236 19.3944
R17996 vdd.n1409 vdd.n1236 19.3944
R17997 vdd.n1409 vdd.n1408 19.3944
R17998 vdd.n1408 vdd.n1407 19.3944
R17999 vdd.n1407 vdd.n1242 19.3944
R18000 vdd.n1403 vdd.n1242 19.3944
R18001 vdd.n1403 vdd.n1402 19.3944
R18002 vdd.n1402 vdd.n1401 19.3944
R18003 vdd.n1401 vdd.n1248 19.3944
R18004 vdd.n1397 vdd.n1248 19.3944
R18005 vdd.n1397 vdd.n1396 19.3944
R18006 vdd.n1396 vdd.n1395 19.3944
R18007 vdd.n1648 vdd.n1583 19.3944
R18008 vdd.n1648 vdd.n1589 19.3944
R18009 vdd.n1643 vdd.n1589 19.3944
R18010 vdd.n1643 vdd.n1642 19.3944
R18011 vdd.n1642 vdd.n1641 19.3944
R18012 vdd.n1641 vdd.n1596 19.3944
R18013 vdd.n1636 vdd.n1596 19.3944
R18014 vdd.n1636 vdd.n1635 19.3944
R18015 vdd.n1635 vdd.n1634 19.3944
R18016 vdd.n1634 vdd.n1603 19.3944
R18017 vdd.n1629 vdd.n1603 19.3944
R18018 vdd.n1629 vdd.n1628 19.3944
R18019 vdd.n1628 vdd.n1627 19.3944
R18020 vdd.n1627 vdd.n1611 19.3944
R18021 vdd.n1622 vdd.n1611 19.3944
R18022 vdd.n1622 vdd.n1621 19.3944
R18023 vdd.n1617 vdd.n1616 19.3944
R18024 vdd.n1950 vdd.n858 19.3944
R18025 vdd.n1687 vdd.n1543 19.3944
R18026 vdd.n1687 vdd.n1549 19.3944
R18027 vdd.n1682 vdd.n1549 19.3944
R18028 vdd.n1682 vdd.n1681 19.3944
R18029 vdd.n1681 vdd.n1680 19.3944
R18030 vdd.n1680 vdd.n1556 19.3944
R18031 vdd.n1675 vdd.n1556 19.3944
R18032 vdd.n1675 vdd.n1674 19.3944
R18033 vdd.n1674 vdd.n1673 19.3944
R18034 vdd.n1673 vdd.n1563 19.3944
R18035 vdd.n1668 vdd.n1563 19.3944
R18036 vdd.n1668 vdd.n1667 19.3944
R18037 vdd.n1667 vdd.n1666 19.3944
R18038 vdd.n1666 vdd.n1570 19.3944
R18039 vdd.n1661 vdd.n1570 19.3944
R18040 vdd.n1661 vdd.n1660 19.3944
R18041 vdd.n1660 vdd.n1659 19.3944
R18042 vdd.n1659 vdd.n1577 19.3944
R18043 vdd.n1654 vdd.n1577 19.3944
R18044 vdd.n1654 vdd.n1653 19.3944
R18045 vdd.n1938 vdd.n1937 19.3944
R18046 vdd.n1937 vdd.n1515 19.3944
R18047 vdd.n1932 vdd.n1931 19.3944
R18048 vdd.n1714 vdd.n1519 19.3944
R18049 vdd.n1714 vdd.n1521 19.3944
R18050 vdd.n1524 vdd.n1521 19.3944
R18051 vdd.n1707 vdd.n1524 19.3944
R18052 vdd.n1707 vdd.n1706 19.3944
R18053 vdd.n1706 vdd.n1705 19.3944
R18054 vdd.n1705 vdd.n1530 19.3944
R18055 vdd.n1700 vdd.n1530 19.3944
R18056 vdd.n1700 vdd.n1699 19.3944
R18057 vdd.n1699 vdd.n1698 19.3944
R18058 vdd.n1698 vdd.n1537 19.3944
R18059 vdd.n1693 vdd.n1537 19.3944
R18060 vdd.n1693 vdd.n1692 19.3944
R18061 vdd.n1428 vdd.n1193 19.3944
R18062 vdd.n1428 vdd.n1184 19.3944
R18063 vdd.n1441 vdd.n1184 19.3944
R18064 vdd.n1441 vdd.n1182 19.3944
R18065 vdd.n1445 vdd.n1182 19.3944
R18066 vdd.n1445 vdd.n1173 19.3944
R18067 vdd.n1458 vdd.n1173 19.3944
R18068 vdd.n1458 vdd.n1171 19.3944
R18069 vdd.n1463 vdd.n1171 19.3944
R18070 vdd.n1463 vdd.n1162 19.3944
R18071 vdd.n1475 vdd.n1162 19.3944
R18072 vdd.n1475 vdd.n890 19.3944
R18073 vdd.n1479 vdd.n890 19.3944
R18074 vdd.n1479 vdd.n880 19.3944
R18075 vdd.n1492 vdd.n880 19.3944
R18076 vdd.n1492 vdd.n878 19.3944
R18077 vdd.n1496 vdd.n878 19.3944
R18078 vdd.n1496 vdd.n868 19.3944
R18079 vdd.n1511 vdd.n868 19.3944
R18080 vdd.n1511 vdd.n866 19.3944
R18081 vdd.n1941 vdd.n866 19.3944
R18082 vdd.n2851 vdd.n477 19.3944
R18083 vdd.n2851 vdd.n475 19.3944
R18084 vdd.n2855 vdd.n475 19.3944
R18085 vdd.n2855 vdd.n465 19.3944
R18086 vdd.n2868 vdd.n465 19.3944
R18087 vdd.n2868 vdd.n463 19.3944
R18088 vdd.n2872 vdd.n463 19.3944
R18089 vdd.n2872 vdd.n453 19.3944
R18090 vdd.n2884 vdd.n453 19.3944
R18091 vdd.n2884 vdd.n451 19.3944
R18092 vdd.n2888 vdd.n451 19.3944
R18093 vdd.n2889 vdd.n2888 19.3944
R18094 vdd.n2890 vdd.n2889 19.3944
R18095 vdd.n2890 vdd.n449 19.3944
R18096 vdd.n2894 vdd.n449 19.3944
R18097 vdd.n2895 vdd.n2894 19.3944
R18098 vdd.n2896 vdd.n2895 19.3944
R18099 vdd.n2896 vdd.n446 19.3944
R18100 vdd.n2900 vdd.n446 19.3944
R18101 vdd.n2901 vdd.n2900 19.3944
R18102 vdd.n2902 vdd.n2901 19.3944
R18103 vdd.n2945 vdd.n404 19.3944
R18104 vdd.n2945 vdd.n410 19.3944
R18105 vdd.n2940 vdd.n410 19.3944
R18106 vdd.n2940 vdd.n2939 19.3944
R18107 vdd.n2939 vdd.n2938 19.3944
R18108 vdd.n2938 vdd.n417 19.3944
R18109 vdd.n2933 vdd.n417 19.3944
R18110 vdd.n2933 vdd.n2932 19.3944
R18111 vdd.n2932 vdd.n2931 19.3944
R18112 vdd.n2931 vdd.n424 19.3944
R18113 vdd.n2926 vdd.n424 19.3944
R18114 vdd.n2926 vdd.n2925 19.3944
R18115 vdd.n2925 vdd.n2924 19.3944
R18116 vdd.n2924 vdd.n431 19.3944
R18117 vdd.n2919 vdd.n431 19.3944
R18118 vdd.n2919 vdd.n2918 19.3944
R18119 vdd.n2918 vdd.n2917 19.3944
R18120 vdd.n2917 vdd.n438 19.3944
R18121 vdd.n2912 vdd.n438 19.3944
R18122 vdd.n2912 vdd.n2911 19.3944
R18123 vdd.n2984 vdd.n364 19.3944
R18124 vdd.n2984 vdd.n370 19.3944
R18125 vdd.n2979 vdd.n370 19.3944
R18126 vdd.n2979 vdd.n2978 19.3944
R18127 vdd.n2978 vdd.n2977 19.3944
R18128 vdd.n2977 vdd.n377 19.3944
R18129 vdd.n2972 vdd.n377 19.3944
R18130 vdd.n2972 vdd.n2971 19.3944
R18131 vdd.n2971 vdd.n2970 19.3944
R18132 vdd.n2970 vdd.n384 19.3944
R18133 vdd.n2965 vdd.n384 19.3944
R18134 vdd.n2965 vdd.n2964 19.3944
R18135 vdd.n2964 vdd.n2963 19.3944
R18136 vdd.n2963 vdd.n391 19.3944
R18137 vdd.n2958 vdd.n391 19.3944
R18138 vdd.n2958 vdd.n2957 19.3944
R18139 vdd.n2957 vdd.n2956 19.3944
R18140 vdd.n2956 vdd.n398 19.3944
R18141 vdd.n2951 vdd.n398 19.3944
R18142 vdd.n2951 vdd.n2950 19.3944
R18143 vdd.n3020 vdd.n3019 19.3944
R18144 vdd.n3019 vdd.n3018 19.3944
R18145 vdd.n3018 vdd.n336 19.3944
R18146 vdd.n337 vdd.n336 19.3944
R18147 vdd.n3011 vdd.n337 19.3944
R18148 vdd.n3011 vdd.n3010 19.3944
R18149 vdd.n3010 vdd.n3009 19.3944
R18150 vdd.n3009 vdd.n344 19.3944
R18151 vdd.n3004 vdd.n344 19.3944
R18152 vdd.n3004 vdd.n3003 19.3944
R18153 vdd.n3003 vdd.n3002 19.3944
R18154 vdd.n3002 vdd.n351 19.3944
R18155 vdd.n2997 vdd.n351 19.3944
R18156 vdd.n2997 vdd.n2996 19.3944
R18157 vdd.n2996 vdd.n2995 19.3944
R18158 vdd.n2995 vdd.n358 19.3944
R18159 vdd.n2990 vdd.n358 19.3944
R18160 vdd.n2990 vdd.n2989 19.3944
R18161 vdd.n2847 vdd.n480 19.3944
R18162 vdd.n2847 vdd.n471 19.3944
R18163 vdd.n2860 vdd.n471 19.3944
R18164 vdd.n2860 vdd.n469 19.3944
R18165 vdd.n2864 vdd.n469 19.3944
R18166 vdd.n2864 vdd.n460 19.3944
R18167 vdd.n2876 vdd.n460 19.3944
R18168 vdd.n2876 vdd.n458 19.3944
R18169 vdd.n2880 vdd.n458 19.3944
R18170 vdd.n2880 vdd.n300 19.3944
R18171 vdd.n3045 vdd.n300 19.3944
R18172 vdd.n3045 vdd.n301 19.3944
R18173 vdd.n3039 vdd.n301 19.3944
R18174 vdd.n3039 vdd.n3038 19.3944
R18175 vdd.n3038 vdd.n3037 19.3944
R18176 vdd.n3037 vdd.n313 19.3944
R18177 vdd.n3031 vdd.n313 19.3944
R18178 vdd.n3031 vdd.n3030 19.3944
R18179 vdd.n3030 vdd.n3029 19.3944
R18180 vdd.n3029 vdd.n324 19.3944
R18181 vdd.n3023 vdd.n324 19.3944
R18182 vdd.n2800 vdd.n536 19.3944
R18183 vdd.n2800 vdd.n2797 19.3944
R18184 vdd.n2797 vdd.n2794 19.3944
R18185 vdd.n2794 vdd.n2793 19.3944
R18186 vdd.n2793 vdd.n2790 19.3944
R18187 vdd.n2790 vdd.n2789 19.3944
R18188 vdd.n2789 vdd.n2786 19.3944
R18189 vdd.n2786 vdd.n2785 19.3944
R18190 vdd.n2785 vdd.n2782 19.3944
R18191 vdd.n2782 vdd.n2781 19.3944
R18192 vdd.n2781 vdd.n2778 19.3944
R18193 vdd.n2778 vdd.n2777 19.3944
R18194 vdd.n2777 vdd.n2774 19.3944
R18195 vdd.n2774 vdd.n2773 19.3944
R18196 vdd.n2773 vdd.n2770 19.3944
R18197 vdd.n2770 vdd.n2769 19.3944
R18198 vdd.n2769 vdd.n2766 19.3944
R18199 vdd.n2766 vdd.n2765 19.3944
R18200 vdd.n2765 vdd.n2762 19.3944
R18201 vdd.n2762 vdd.n2761 19.3944
R18202 vdd.n2843 vdd.n482 19.3944
R18203 vdd.n2838 vdd.n482 19.3944
R18204 vdd.n521 vdd.n518 19.3944
R18205 vdd.n2834 vdd.n2833 19.3944
R18206 vdd.n2833 vdd.n2830 19.3944
R18207 vdd.n2830 vdd.n2829 19.3944
R18208 vdd.n2829 vdd.n2826 19.3944
R18209 vdd.n2826 vdd.n2825 19.3944
R18210 vdd.n2825 vdd.n2822 19.3944
R18211 vdd.n2822 vdd.n2821 19.3944
R18212 vdd.n2821 vdd.n2818 19.3944
R18213 vdd.n2818 vdd.n2817 19.3944
R18214 vdd.n2817 vdd.n2814 19.3944
R18215 vdd.n2814 vdd.n2813 19.3944
R18216 vdd.n2813 vdd.n2810 19.3944
R18217 vdd.n2810 vdd.n2809 19.3944
R18218 vdd.n2754 vdd.n556 19.3944
R18219 vdd.n2754 vdd.n2751 19.3944
R18220 vdd.n2751 vdd.n2748 19.3944
R18221 vdd.n2748 vdd.n2747 19.3944
R18222 vdd.n2747 vdd.n2744 19.3944
R18223 vdd.n2744 vdd.n2743 19.3944
R18224 vdd.n2743 vdd.n2740 19.3944
R18225 vdd.n2740 vdd.n2739 19.3944
R18226 vdd.n2739 vdd.n2736 19.3944
R18227 vdd.n2736 vdd.n2735 19.3944
R18228 vdd.n2735 vdd.n2732 19.3944
R18229 vdd.n2732 vdd.n2731 19.3944
R18230 vdd.n2731 vdd.n2728 19.3944
R18231 vdd.n2728 vdd.n2727 19.3944
R18232 vdd.n2727 vdd.n2724 19.3944
R18233 vdd.n2724 vdd.n2723 19.3944
R18234 vdd.n2720 vdd.n2719 19.3944
R18235 vdd.n2716 vdd.n2715 19.3944
R18236 vdd.n1360 vdd.n1356 19.0066
R18237 vdd.n1652 vdd.n1583 19.0066
R18238 vdd.n2949 vdd.n404 19.0066
R18239 vdd.n2758 vdd.n556 19.0066
R18240 vdd.n1792 vdd.n1791 16.0975
R18241 vdd.n756 vdd.n755 16.0975
R18242 vdd.n1321 vdd.n1320 16.0975
R18243 vdd.n1359 vdd.n1358 16.0975
R18244 vdd.n1255 vdd.n1254 16.0975
R18245 vdd.n1948 vdd.n1947 16.0975
R18246 vdd.n1585 vdd.n1584 16.0975
R18247 vdd.n1545 vdd.n1544 16.0975
R18248 vdd.n1766 vdd.n1765 16.0975
R18249 vdd.n748 vdd.n747 16.0975
R18250 vdd.n2257 vdd.n2256 16.0975
R18251 vdd.n2909 vdd.n2908 16.0975
R18252 vdd.n406 vdd.n405 16.0975
R18253 vdd.n366 vdd.n365 16.0975
R18254 vdd.n558 vdd.n557 16.0975
R18255 vdd.n2805 vdd.n2804 16.0975
R18256 vdd.n623 vdd.n622 16.0975
R18257 vdd.n2254 vdd.n2253 16.0975
R18258 vdd.n2712 vdd.n2711 16.0975
R18259 vdd.n590 vdd.n589 16.0975
R18260 vdd.t36 vdd.n2218 15.4182
R18261 vdd.n2471 vdd.t38 15.4182
R18262 vdd.n28 vdd.n27 14.5458
R18263 vdd.n1989 vdd.n839 14.5112
R18264 vdd.n2673 vdd.n484 14.5112
R18265 vdd.n292 vdd.n257 13.1884
R18266 vdd.n245 vdd.n210 13.1884
R18267 vdd.n202 vdd.n167 13.1884
R18268 vdd.n155 vdd.n120 13.1884
R18269 vdd.n113 vdd.n78 13.1884
R18270 vdd.n66 vdd.n31 13.1884
R18271 vdd.n1107 vdd.n1072 13.1884
R18272 vdd.n1154 vdd.n1119 13.1884
R18273 vdd.n1017 vdd.n982 13.1884
R18274 vdd.n1064 vdd.n1029 13.1884
R18275 vdd.n928 vdd.n893 13.1884
R18276 vdd.n975 vdd.n940 13.1884
R18277 vdd.n1391 vdd.n1256 12.9944
R18278 vdd.n1395 vdd.n1256 12.9944
R18279 vdd.n1691 vdd.n1543 12.9944
R18280 vdd.n1692 vdd.n1691 12.9944
R18281 vdd.n2988 vdd.n364 12.9944
R18282 vdd.n2989 vdd.n2988 12.9944
R18283 vdd.n2806 vdd.n536 12.9944
R18284 vdd.n2809 vdd.n2806 12.9944
R18285 vdd.n293 vdd.n255 12.8005
R18286 vdd.n288 vdd.n259 12.8005
R18287 vdd.n246 vdd.n208 12.8005
R18288 vdd.n241 vdd.n212 12.8005
R18289 vdd.n203 vdd.n165 12.8005
R18290 vdd.n198 vdd.n169 12.8005
R18291 vdd.n156 vdd.n118 12.8005
R18292 vdd.n151 vdd.n122 12.8005
R18293 vdd.n114 vdd.n76 12.8005
R18294 vdd.n109 vdd.n80 12.8005
R18295 vdd.n67 vdd.n29 12.8005
R18296 vdd.n62 vdd.n33 12.8005
R18297 vdd.n1108 vdd.n1070 12.8005
R18298 vdd.n1103 vdd.n1074 12.8005
R18299 vdd.n1155 vdd.n1117 12.8005
R18300 vdd.n1150 vdd.n1121 12.8005
R18301 vdd.n1018 vdd.n980 12.8005
R18302 vdd.n1013 vdd.n984 12.8005
R18303 vdd.n1065 vdd.n1027 12.8005
R18304 vdd.n1060 vdd.n1031 12.8005
R18305 vdd.n929 vdd.n891 12.8005
R18306 vdd.n924 vdd.n895 12.8005
R18307 vdd.n976 vdd.n938 12.8005
R18308 vdd.n971 vdd.n942 12.8005
R18309 vdd.n287 vdd.n260 12.0247
R18310 vdd.n240 vdd.n213 12.0247
R18311 vdd.n197 vdd.n170 12.0247
R18312 vdd.n150 vdd.n123 12.0247
R18313 vdd.n108 vdd.n81 12.0247
R18314 vdd.n61 vdd.n34 12.0247
R18315 vdd.n1102 vdd.n1075 12.0247
R18316 vdd.n1149 vdd.n1122 12.0247
R18317 vdd.n1012 vdd.n985 12.0247
R18318 vdd.n1059 vdd.n1032 12.0247
R18319 vdd.n923 vdd.n896 12.0247
R18320 vdd.n970 vdd.n943 12.0247
R18321 vdd.n1430 vdd.n1186 11.337
R18322 vdd.n1439 vdd.n1186 11.337
R18323 vdd.n1439 vdd.n1438 11.337
R18324 vdd.n1447 vdd.n1180 11.337
R18325 vdd.n1456 vdd.n1455 11.337
R18326 vdd.n1473 vdd.n1164 11.337
R18327 vdd.n1481 vdd.n887 11.337
R18328 vdd.n1490 vdd.n1489 11.337
R18329 vdd.n1498 vdd.n870 11.337
R18330 vdd.n1509 vdd.n870 11.337
R18331 vdd.n1509 vdd.n1508 11.337
R18332 vdd.n2849 vdd.n473 11.337
R18333 vdd.n2858 vdd.n473 11.337
R18334 vdd.n2858 vdd.n2857 11.337
R18335 vdd.n2866 vdd.n467 11.337
R18336 vdd.n2882 vdd.n456 11.337
R18337 vdd.n3043 vdd.n304 11.337
R18338 vdd.n3041 vdd.n308 11.337
R18339 vdd.n3035 vdd.n3034 11.337
R18340 vdd.n3033 vdd.n318 11.337
R18341 vdd.n3027 vdd.n318 11.337
R18342 vdd.n3027 vdd.n3026 11.337
R18343 vdd.n284 vdd.n283 11.249
R18344 vdd.n237 vdd.n236 11.249
R18345 vdd.n194 vdd.n193 11.249
R18346 vdd.n147 vdd.n146 11.249
R18347 vdd.n105 vdd.n104 11.249
R18348 vdd.n58 vdd.n57 11.249
R18349 vdd.n1099 vdd.n1098 11.249
R18350 vdd.n1146 vdd.n1145 11.249
R18351 vdd.n1009 vdd.n1008 11.249
R18352 vdd.n1056 vdd.n1055 11.249
R18353 vdd.n920 vdd.n919 11.249
R18354 vdd.n967 vdd.n966 11.249
R18355 vdd.n2146 vdd.t16 11.1103
R18356 vdd.n2478 vdd.t192 11.1103
R18357 vdd.n1228 vdd.t53 10.7702
R18358 vdd.t64 vdd.n3025 10.7702
R18359 vdd.n269 vdd.n268 10.7238
R18360 vdd.n222 vdd.n221 10.7238
R18361 vdd.n179 vdd.n178 10.7238
R18362 vdd.n132 vdd.n131 10.7238
R18363 vdd.n90 vdd.n89 10.7238
R18364 vdd.n43 vdd.n42 10.7238
R18365 vdd.n1084 vdd.n1083 10.7238
R18366 vdd.n1131 vdd.n1130 10.7238
R18367 vdd.n994 vdd.n993 10.7238
R18368 vdd.n1041 vdd.n1040 10.7238
R18369 vdd.n905 vdd.n904 10.7238
R18370 vdd.n952 vdd.n951 10.7238
R18371 vdd.n1992 vdd.n1991 10.6151
R18372 vdd.n1993 vdd.n1992 10.6151
R18373 vdd.n1993 vdd.n825 10.6151
R18374 vdd.n2003 vdd.n825 10.6151
R18375 vdd.n2004 vdd.n2003 10.6151
R18376 vdd.n2005 vdd.n2004 10.6151
R18377 vdd.n2005 vdd.n812 10.6151
R18378 vdd.n2016 vdd.n812 10.6151
R18379 vdd.n2017 vdd.n2016 10.6151
R18380 vdd.n2018 vdd.n2017 10.6151
R18381 vdd.n2018 vdd.n800 10.6151
R18382 vdd.n2028 vdd.n800 10.6151
R18383 vdd.n2029 vdd.n2028 10.6151
R18384 vdd.n2030 vdd.n2029 10.6151
R18385 vdd.n2030 vdd.n788 10.6151
R18386 vdd.n2040 vdd.n788 10.6151
R18387 vdd.n2041 vdd.n2040 10.6151
R18388 vdd.n2042 vdd.n2041 10.6151
R18389 vdd.n2042 vdd.n777 10.6151
R18390 vdd.n2052 vdd.n777 10.6151
R18391 vdd.n2053 vdd.n2052 10.6151
R18392 vdd.n2054 vdd.n2053 10.6151
R18393 vdd.n2054 vdd.n764 10.6151
R18394 vdd.n2066 vdd.n764 10.6151
R18395 vdd.n2067 vdd.n2066 10.6151
R18396 vdd.n2069 vdd.n2067 10.6151
R18397 vdd.n2069 vdd.n2068 10.6151
R18398 vdd.n2068 vdd.n746 10.6151
R18399 vdd.n2216 vdd.n2215 10.6151
R18400 vdd.n2215 vdd.n2214 10.6151
R18401 vdd.n2214 vdd.n2211 10.6151
R18402 vdd.n2211 vdd.n2210 10.6151
R18403 vdd.n2210 vdd.n2207 10.6151
R18404 vdd.n2207 vdd.n2206 10.6151
R18405 vdd.n2206 vdd.n2203 10.6151
R18406 vdd.n2203 vdd.n2202 10.6151
R18407 vdd.n2202 vdd.n2199 10.6151
R18408 vdd.n2199 vdd.n2198 10.6151
R18409 vdd.n2198 vdd.n2195 10.6151
R18410 vdd.n2195 vdd.n2194 10.6151
R18411 vdd.n2194 vdd.n2191 10.6151
R18412 vdd.n2191 vdd.n2190 10.6151
R18413 vdd.n2190 vdd.n2187 10.6151
R18414 vdd.n2187 vdd.n2186 10.6151
R18415 vdd.n2186 vdd.n2183 10.6151
R18416 vdd.n2183 vdd.n2182 10.6151
R18417 vdd.n2182 vdd.n2179 10.6151
R18418 vdd.n2179 vdd.n2178 10.6151
R18419 vdd.n2178 vdd.n2175 10.6151
R18420 vdd.n2175 vdd.n2174 10.6151
R18421 vdd.n2174 vdd.n2171 10.6151
R18422 vdd.n2171 vdd.n2170 10.6151
R18423 vdd.n2170 vdd.n2167 10.6151
R18424 vdd.n2167 vdd.n2166 10.6151
R18425 vdd.n2166 vdd.n2163 10.6151
R18426 vdd.n2163 vdd.n2162 10.6151
R18427 vdd.n2162 vdd.n2159 10.6151
R18428 vdd.n2159 vdd.n2158 10.6151
R18429 vdd.n2158 vdd.n2155 10.6151
R18430 vdd.n2153 vdd.n2150 10.6151
R18431 vdd.n2150 vdd.n2149 10.6151
R18432 vdd.n1892 vdd.n1891 10.6151
R18433 vdd.n1891 vdd.n1889 10.6151
R18434 vdd.n1889 vdd.n1888 10.6151
R18435 vdd.n1888 vdd.n1886 10.6151
R18436 vdd.n1886 vdd.n1885 10.6151
R18437 vdd.n1885 vdd.n1883 10.6151
R18438 vdd.n1883 vdd.n1882 10.6151
R18439 vdd.n1882 vdd.n1880 10.6151
R18440 vdd.n1880 vdd.n1879 10.6151
R18441 vdd.n1879 vdd.n1877 10.6151
R18442 vdd.n1877 vdd.n1876 10.6151
R18443 vdd.n1876 vdd.n1874 10.6151
R18444 vdd.n1874 vdd.n1873 10.6151
R18445 vdd.n1873 vdd.n1788 10.6151
R18446 vdd.n1788 vdd.n1787 10.6151
R18447 vdd.n1787 vdd.n1785 10.6151
R18448 vdd.n1785 vdd.n1784 10.6151
R18449 vdd.n1784 vdd.n1782 10.6151
R18450 vdd.n1782 vdd.n1781 10.6151
R18451 vdd.n1781 vdd.n1779 10.6151
R18452 vdd.n1779 vdd.n1778 10.6151
R18453 vdd.n1778 vdd.n1776 10.6151
R18454 vdd.n1776 vdd.n1775 10.6151
R18455 vdd.n1775 vdd.n1773 10.6151
R18456 vdd.n1773 vdd.n1772 10.6151
R18457 vdd.n1772 vdd.n1769 10.6151
R18458 vdd.n1769 vdd.n1768 10.6151
R18459 vdd.n1768 vdd.n749 10.6151
R18460 vdd.n1726 vdd.n837 10.6151
R18461 vdd.n1727 vdd.n1726 10.6151
R18462 vdd.n1728 vdd.n1727 10.6151
R18463 vdd.n1728 vdd.n1722 10.6151
R18464 vdd.n1734 vdd.n1722 10.6151
R18465 vdd.n1735 vdd.n1734 10.6151
R18466 vdd.n1736 vdd.n1735 10.6151
R18467 vdd.n1736 vdd.n1720 10.6151
R18468 vdd.n1742 vdd.n1720 10.6151
R18469 vdd.n1743 vdd.n1742 10.6151
R18470 vdd.n1744 vdd.n1743 10.6151
R18471 vdd.n1744 vdd.n1718 10.6151
R18472 vdd.n1750 vdd.n1718 10.6151
R18473 vdd.n1751 vdd.n1750 10.6151
R18474 vdd.n1752 vdd.n1751 10.6151
R18475 vdd.n1752 vdd.n1716 10.6151
R18476 vdd.n1928 vdd.n1716 10.6151
R18477 vdd.n1928 vdd.n1927 10.6151
R18478 vdd.n1927 vdd.n1757 10.6151
R18479 vdd.n1921 vdd.n1757 10.6151
R18480 vdd.n1921 vdd.n1920 10.6151
R18481 vdd.n1920 vdd.n1919 10.6151
R18482 vdd.n1919 vdd.n1759 10.6151
R18483 vdd.n1913 vdd.n1759 10.6151
R18484 vdd.n1913 vdd.n1912 10.6151
R18485 vdd.n1912 vdd.n1911 10.6151
R18486 vdd.n1911 vdd.n1761 10.6151
R18487 vdd.n1905 vdd.n1761 10.6151
R18488 vdd.n1905 vdd.n1904 10.6151
R18489 vdd.n1904 vdd.n1903 10.6151
R18490 vdd.n1903 vdd.n1763 10.6151
R18491 vdd.n1897 vdd.n1896 10.6151
R18492 vdd.n1896 vdd.n1895 10.6151
R18493 vdd.n2401 vdd.n2400 10.6151
R18494 vdd.n2400 vdd.n2398 10.6151
R18495 vdd.n2398 vdd.n2397 10.6151
R18496 vdd.n2397 vdd.n2255 10.6151
R18497 vdd.n2344 vdd.n2255 10.6151
R18498 vdd.n2345 vdd.n2344 10.6151
R18499 vdd.n2347 vdd.n2345 10.6151
R18500 vdd.n2348 vdd.n2347 10.6151
R18501 vdd.n2350 vdd.n2348 10.6151
R18502 vdd.n2351 vdd.n2350 10.6151
R18503 vdd.n2353 vdd.n2351 10.6151
R18504 vdd.n2354 vdd.n2353 10.6151
R18505 vdd.n2356 vdd.n2354 10.6151
R18506 vdd.n2357 vdd.n2356 10.6151
R18507 vdd.n2372 vdd.n2357 10.6151
R18508 vdd.n2372 vdd.n2371 10.6151
R18509 vdd.n2371 vdd.n2370 10.6151
R18510 vdd.n2370 vdd.n2368 10.6151
R18511 vdd.n2368 vdd.n2367 10.6151
R18512 vdd.n2367 vdd.n2365 10.6151
R18513 vdd.n2365 vdd.n2364 10.6151
R18514 vdd.n2364 vdd.n2362 10.6151
R18515 vdd.n2362 vdd.n2361 10.6151
R18516 vdd.n2361 vdd.n2359 10.6151
R18517 vdd.n2359 vdd.n2358 10.6151
R18518 vdd.n2358 vdd.n626 10.6151
R18519 vdd.n2606 vdd.n626 10.6151
R18520 vdd.n2607 vdd.n2606 10.6151
R18521 vdd.n2468 vdd.n702 10.6151
R18522 vdd.n2468 vdd.n2467 10.6151
R18523 vdd.n2467 vdd.n2466 10.6151
R18524 vdd.n2466 vdd.n2464 10.6151
R18525 vdd.n2464 vdd.n2461 10.6151
R18526 vdd.n2461 vdd.n2460 10.6151
R18527 vdd.n2460 vdd.n2457 10.6151
R18528 vdd.n2457 vdd.n2456 10.6151
R18529 vdd.n2456 vdd.n2453 10.6151
R18530 vdd.n2453 vdd.n2452 10.6151
R18531 vdd.n2452 vdd.n2449 10.6151
R18532 vdd.n2449 vdd.n2448 10.6151
R18533 vdd.n2448 vdd.n2445 10.6151
R18534 vdd.n2445 vdd.n2444 10.6151
R18535 vdd.n2444 vdd.n2441 10.6151
R18536 vdd.n2441 vdd.n2440 10.6151
R18537 vdd.n2440 vdd.n2437 10.6151
R18538 vdd.n2437 vdd.n2436 10.6151
R18539 vdd.n2436 vdd.n2433 10.6151
R18540 vdd.n2433 vdd.n2432 10.6151
R18541 vdd.n2432 vdd.n2429 10.6151
R18542 vdd.n2429 vdd.n2428 10.6151
R18543 vdd.n2428 vdd.n2425 10.6151
R18544 vdd.n2425 vdd.n2424 10.6151
R18545 vdd.n2424 vdd.n2421 10.6151
R18546 vdd.n2421 vdd.n2420 10.6151
R18547 vdd.n2420 vdd.n2417 10.6151
R18548 vdd.n2417 vdd.n2416 10.6151
R18549 vdd.n2416 vdd.n2413 10.6151
R18550 vdd.n2413 vdd.n2412 10.6151
R18551 vdd.n2412 vdd.n2409 10.6151
R18552 vdd.n2407 vdd.n2404 10.6151
R18553 vdd.n2404 vdd.n2403 10.6151
R18554 vdd.n2481 vdd.n2480 10.6151
R18555 vdd.n2482 vdd.n2481 10.6151
R18556 vdd.n2482 vdd.n692 10.6151
R18557 vdd.n2492 vdd.n692 10.6151
R18558 vdd.n2493 vdd.n2492 10.6151
R18559 vdd.n2494 vdd.n2493 10.6151
R18560 vdd.n2494 vdd.n679 10.6151
R18561 vdd.n2504 vdd.n679 10.6151
R18562 vdd.n2505 vdd.n2504 10.6151
R18563 vdd.n2506 vdd.n2505 10.6151
R18564 vdd.n2506 vdd.n668 10.6151
R18565 vdd.n2516 vdd.n668 10.6151
R18566 vdd.n2517 vdd.n2516 10.6151
R18567 vdd.n2518 vdd.n2517 10.6151
R18568 vdd.n2518 vdd.n656 10.6151
R18569 vdd.n2528 vdd.n656 10.6151
R18570 vdd.n2529 vdd.n2528 10.6151
R18571 vdd.n2530 vdd.n2529 10.6151
R18572 vdd.n2530 vdd.n645 10.6151
R18573 vdd.n2542 vdd.n645 10.6151
R18574 vdd.n2543 vdd.n2542 10.6151
R18575 vdd.n2544 vdd.n2543 10.6151
R18576 vdd.n2544 vdd.n631 10.6151
R18577 vdd.n2599 vdd.n631 10.6151
R18578 vdd.n2600 vdd.n2599 10.6151
R18579 vdd.n2601 vdd.n2600 10.6151
R18580 vdd.n2601 vdd.n600 10.6151
R18581 vdd.n2671 vdd.n600 10.6151
R18582 vdd.n2670 vdd.n2669 10.6151
R18583 vdd.n2669 vdd.n601 10.6151
R18584 vdd.n602 vdd.n601 10.6151
R18585 vdd.n2662 vdd.n602 10.6151
R18586 vdd.n2662 vdd.n2661 10.6151
R18587 vdd.n2661 vdd.n2660 10.6151
R18588 vdd.n2660 vdd.n604 10.6151
R18589 vdd.n2655 vdd.n604 10.6151
R18590 vdd.n2655 vdd.n2654 10.6151
R18591 vdd.n2654 vdd.n2653 10.6151
R18592 vdd.n2653 vdd.n607 10.6151
R18593 vdd.n2648 vdd.n607 10.6151
R18594 vdd.n2648 vdd.n2647 10.6151
R18595 vdd.n2647 vdd.n2646 10.6151
R18596 vdd.n2646 vdd.n610 10.6151
R18597 vdd.n2641 vdd.n610 10.6151
R18598 vdd.n2641 vdd.n520 10.6151
R18599 vdd.n2637 vdd.n520 10.6151
R18600 vdd.n2637 vdd.n2636 10.6151
R18601 vdd.n2636 vdd.n2635 10.6151
R18602 vdd.n2635 vdd.n613 10.6151
R18603 vdd.n2630 vdd.n613 10.6151
R18604 vdd.n2630 vdd.n2629 10.6151
R18605 vdd.n2629 vdd.n2628 10.6151
R18606 vdd.n2628 vdd.n616 10.6151
R18607 vdd.n2623 vdd.n616 10.6151
R18608 vdd.n2623 vdd.n2622 10.6151
R18609 vdd.n2622 vdd.n2621 10.6151
R18610 vdd.n2621 vdd.n619 10.6151
R18611 vdd.n2616 vdd.n619 10.6151
R18612 vdd.n2616 vdd.n2615 10.6151
R18613 vdd.n2613 vdd.n624 10.6151
R18614 vdd.n2608 vdd.n624 10.6151
R18615 vdd.n2589 vdd.n2550 10.6151
R18616 vdd.n2584 vdd.n2550 10.6151
R18617 vdd.n2584 vdd.n2583 10.6151
R18618 vdd.n2583 vdd.n2582 10.6151
R18619 vdd.n2582 vdd.n2552 10.6151
R18620 vdd.n2577 vdd.n2552 10.6151
R18621 vdd.n2577 vdd.n2576 10.6151
R18622 vdd.n2576 vdd.n2575 10.6151
R18623 vdd.n2575 vdd.n2555 10.6151
R18624 vdd.n2570 vdd.n2555 10.6151
R18625 vdd.n2570 vdd.n2569 10.6151
R18626 vdd.n2569 vdd.n2568 10.6151
R18627 vdd.n2568 vdd.n2558 10.6151
R18628 vdd.n2563 vdd.n2558 10.6151
R18629 vdd.n2563 vdd.n2562 10.6151
R18630 vdd.n2562 vdd.n575 10.6151
R18631 vdd.n2706 vdd.n575 10.6151
R18632 vdd.n2706 vdd.n576 10.6151
R18633 vdd.n578 vdd.n576 10.6151
R18634 vdd.n2699 vdd.n578 10.6151
R18635 vdd.n2699 vdd.n2698 10.6151
R18636 vdd.n2698 vdd.n2697 10.6151
R18637 vdd.n2697 vdd.n580 10.6151
R18638 vdd.n2692 vdd.n580 10.6151
R18639 vdd.n2692 vdd.n2691 10.6151
R18640 vdd.n2691 vdd.n2690 10.6151
R18641 vdd.n2690 vdd.n583 10.6151
R18642 vdd.n2685 vdd.n583 10.6151
R18643 vdd.n2685 vdd.n2684 10.6151
R18644 vdd.n2684 vdd.n2683 10.6151
R18645 vdd.n2683 vdd.n586 10.6151
R18646 vdd.n2678 vdd.n2677 10.6151
R18647 vdd.n2677 vdd.n2676 10.6151
R18648 vdd.n2324 vdd.n2322 10.6151
R18649 vdd.n2325 vdd.n2324 10.6151
R18650 vdd.n2393 vdd.n2325 10.6151
R18651 vdd.n2393 vdd.n2392 10.6151
R18652 vdd.n2392 vdd.n2391 10.6151
R18653 vdd.n2391 vdd.n2389 10.6151
R18654 vdd.n2389 vdd.n2388 10.6151
R18655 vdd.n2388 vdd.n2386 10.6151
R18656 vdd.n2386 vdd.n2385 10.6151
R18657 vdd.n2385 vdd.n2383 10.6151
R18658 vdd.n2383 vdd.n2382 10.6151
R18659 vdd.n2382 vdd.n2380 10.6151
R18660 vdd.n2380 vdd.n2379 10.6151
R18661 vdd.n2379 vdd.n2377 10.6151
R18662 vdd.n2377 vdd.n2376 10.6151
R18663 vdd.n2376 vdd.n2342 10.6151
R18664 vdd.n2342 vdd.n2341 10.6151
R18665 vdd.n2341 vdd.n2339 10.6151
R18666 vdd.n2339 vdd.n2338 10.6151
R18667 vdd.n2338 vdd.n2336 10.6151
R18668 vdd.n2336 vdd.n2335 10.6151
R18669 vdd.n2335 vdd.n2333 10.6151
R18670 vdd.n2333 vdd.n2332 10.6151
R18671 vdd.n2332 vdd.n2330 10.6151
R18672 vdd.n2330 vdd.n2329 10.6151
R18673 vdd.n2329 vdd.n2327 10.6151
R18674 vdd.n2327 vdd.n2326 10.6151
R18675 vdd.n2326 vdd.n592 10.6151
R18676 vdd.n2475 vdd.n2474 10.6151
R18677 vdd.n2474 vdd.n707 10.6151
R18678 vdd.n2259 vdd.n707 10.6151
R18679 vdd.n2262 vdd.n2259 10.6151
R18680 vdd.n2263 vdd.n2262 10.6151
R18681 vdd.n2266 vdd.n2263 10.6151
R18682 vdd.n2267 vdd.n2266 10.6151
R18683 vdd.n2270 vdd.n2267 10.6151
R18684 vdd.n2271 vdd.n2270 10.6151
R18685 vdd.n2274 vdd.n2271 10.6151
R18686 vdd.n2275 vdd.n2274 10.6151
R18687 vdd.n2278 vdd.n2275 10.6151
R18688 vdd.n2279 vdd.n2278 10.6151
R18689 vdd.n2282 vdd.n2279 10.6151
R18690 vdd.n2283 vdd.n2282 10.6151
R18691 vdd.n2286 vdd.n2283 10.6151
R18692 vdd.n2287 vdd.n2286 10.6151
R18693 vdd.n2290 vdd.n2287 10.6151
R18694 vdd.n2291 vdd.n2290 10.6151
R18695 vdd.n2294 vdd.n2291 10.6151
R18696 vdd.n2295 vdd.n2294 10.6151
R18697 vdd.n2298 vdd.n2295 10.6151
R18698 vdd.n2299 vdd.n2298 10.6151
R18699 vdd.n2302 vdd.n2299 10.6151
R18700 vdd.n2303 vdd.n2302 10.6151
R18701 vdd.n2306 vdd.n2303 10.6151
R18702 vdd.n2307 vdd.n2306 10.6151
R18703 vdd.n2310 vdd.n2307 10.6151
R18704 vdd.n2311 vdd.n2310 10.6151
R18705 vdd.n2314 vdd.n2311 10.6151
R18706 vdd.n2315 vdd.n2314 10.6151
R18707 vdd.n2320 vdd.n2318 10.6151
R18708 vdd.n2321 vdd.n2320 10.6151
R18709 vdd.n2476 vdd.n697 10.6151
R18710 vdd.n2486 vdd.n697 10.6151
R18711 vdd.n2487 vdd.n2486 10.6151
R18712 vdd.n2488 vdd.n2487 10.6151
R18713 vdd.n2488 vdd.n685 10.6151
R18714 vdd.n2498 vdd.n685 10.6151
R18715 vdd.n2499 vdd.n2498 10.6151
R18716 vdd.n2500 vdd.n2499 10.6151
R18717 vdd.n2500 vdd.n674 10.6151
R18718 vdd.n2510 vdd.n674 10.6151
R18719 vdd.n2511 vdd.n2510 10.6151
R18720 vdd.n2512 vdd.n2511 10.6151
R18721 vdd.n2512 vdd.n662 10.6151
R18722 vdd.n2522 vdd.n662 10.6151
R18723 vdd.n2523 vdd.n2522 10.6151
R18724 vdd.n2524 vdd.n2523 10.6151
R18725 vdd.n2524 vdd.n651 10.6151
R18726 vdd.n2534 vdd.n651 10.6151
R18727 vdd.n2535 vdd.n2534 10.6151
R18728 vdd.n2538 vdd.n2535 10.6151
R18729 vdd.n2548 vdd.n639 10.6151
R18730 vdd.n2549 vdd.n2548 10.6151
R18731 vdd.n2595 vdd.n2549 10.6151
R18732 vdd.n2595 vdd.n2594 10.6151
R18733 vdd.n2594 vdd.n2593 10.6151
R18734 vdd.n2593 vdd.n2592 10.6151
R18735 vdd.n2592 vdd.n2590 10.6151
R18736 vdd.n1987 vdd.n831 10.6151
R18737 vdd.n1997 vdd.n831 10.6151
R18738 vdd.n1998 vdd.n1997 10.6151
R18739 vdd.n1999 vdd.n1998 10.6151
R18740 vdd.n1999 vdd.n818 10.6151
R18741 vdd.n2009 vdd.n818 10.6151
R18742 vdd.n2010 vdd.n2009 10.6151
R18743 vdd.n2012 vdd.n806 10.6151
R18744 vdd.n2022 vdd.n806 10.6151
R18745 vdd.n2023 vdd.n2022 10.6151
R18746 vdd.n2024 vdd.n2023 10.6151
R18747 vdd.n2024 vdd.n794 10.6151
R18748 vdd.n2034 vdd.n794 10.6151
R18749 vdd.n2035 vdd.n2034 10.6151
R18750 vdd.n2036 vdd.n2035 10.6151
R18751 vdd.n2036 vdd.n783 10.6151
R18752 vdd.n2046 vdd.n783 10.6151
R18753 vdd.n2047 vdd.n2046 10.6151
R18754 vdd.n2048 vdd.n2047 10.6151
R18755 vdd.n2048 vdd.n771 10.6151
R18756 vdd.n2058 vdd.n771 10.6151
R18757 vdd.n2059 vdd.n2058 10.6151
R18758 vdd.n2062 vdd.n2059 10.6151
R18759 vdd.n2062 vdd.n2061 10.6151
R18760 vdd.n2061 vdd.n2060 10.6151
R18761 vdd.n2060 vdd.n754 10.6151
R18762 vdd.n2144 vdd.n754 10.6151
R18763 vdd.n2143 vdd.n2142 10.6151
R18764 vdd.n2142 vdd.n2139 10.6151
R18765 vdd.n2139 vdd.n2138 10.6151
R18766 vdd.n2138 vdd.n2135 10.6151
R18767 vdd.n2135 vdd.n2134 10.6151
R18768 vdd.n2134 vdd.n2131 10.6151
R18769 vdd.n2131 vdd.n2130 10.6151
R18770 vdd.n2130 vdd.n2127 10.6151
R18771 vdd.n2127 vdd.n2126 10.6151
R18772 vdd.n2126 vdd.n2123 10.6151
R18773 vdd.n2123 vdd.n2122 10.6151
R18774 vdd.n2122 vdd.n2119 10.6151
R18775 vdd.n2119 vdd.n2118 10.6151
R18776 vdd.n2118 vdd.n2115 10.6151
R18777 vdd.n2115 vdd.n2114 10.6151
R18778 vdd.n2114 vdd.n2111 10.6151
R18779 vdd.n2111 vdd.n2110 10.6151
R18780 vdd.n2110 vdd.n2107 10.6151
R18781 vdd.n2107 vdd.n2106 10.6151
R18782 vdd.n2106 vdd.n2103 10.6151
R18783 vdd.n2103 vdd.n2102 10.6151
R18784 vdd.n2102 vdd.n2099 10.6151
R18785 vdd.n2099 vdd.n2098 10.6151
R18786 vdd.n2098 vdd.n2095 10.6151
R18787 vdd.n2095 vdd.n2094 10.6151
R18788 vdd.n2094 vdd.n2091 10.6151
R18789 vdd.n2091 vdd.n2090 10.6151
R18790 vdd.n2090 vdd.n2087 10.6151
R18791 vdd.n2087 vdd.n2086 10.6151
R18792 vdd.n2086 vdd.n2083 10.6151
R18793 vdd.n2083 vdd.n2082 10.6151
R18794 vdd.n2079 vdd.n2078 10.6151
R18795 vdd.n2078 vdd.n2076 10.6151
R18796 vdd.n1835 vdd.n1833 10.6151
R18797 vdd.n1836 vdd.n1835 10.6151
R18798 vdd.n1838 vdd.n1836 10.6151
R18799 vdd.n1839 vdd.n1838 10.6151
R18800 vdd.n1841 vdd.n1839 10.6151
R18801 vdd.n1842 vdd.n1841 10.6151
R18802 vdd.n1844 vdd.n1842 10.6151
R18803 vdd.n1845 vdd.n1844 10.6151
R18804 vdd.n1847 vdd.n1845 10.6151
R18805 vdd.n1848 vdd.n1847 10.6151
R18806 vdd.n1850 vdd.n1848 10.6151
R18807 vdd.n1851 vdd.n1850 10.6151
R18808 vdd.n1869 vdd.n1851 10.6151
R18809 vdd.n1869 vdd.n1868 10.6151
R18810 vdd.n1868 vdd.n1867 10.6151
R18811 vdd.n1867 vdd.n1865 10.6151
R18812 vdd.n1865 vdd.n1864 10.6151
R18813 vdd.n1864 vdd.n1862 10.6151
R18814 vdd.n1862 vdd.n1861 10.6151
R18815 vdd.n1861 vdd.n1859 10.6151
R18816 vdd.n1859 vdd.n1858 10.6151
R18817 vdd.n1858 vdd.n1856 10.6151
R18818 vdd.n1856 vdd.n1855 10.6151
R18819 vdd.n1855 vdd.n1853 10.6151
R18820 vdd.n1853 vdd.n1852 10.6151
R18821 vdd.n1852 vdd.n758 10.6151
R18822 vdd.n2074 vdd.n758 10.6151
R18823 vdd.n2075 vdd.n2074 10.6151
R18824 vdd.n1986 vdd.n1985 10.6151
R18825 vdd.n1985 vdd.n843 10.6151
R18826 vdd.n1979 vdd.n843 10.6151
R18827 vdd.n1979 vdd.n1978 10.6151
R18828 vdd.n1978 vdd.n1977 10.6151
R18829 vdd.n1977 vdd.n845 10.6151
R18830 vdd.n1971 vdd.n845 10.6151
R18831 vdd.n1971 vdd.n1970 10.6151
R18832 vdd.n1970 vdd.n1969 10.6151
R18833 vdd.n1969 vdd.n847 10.6151
R18834 vdd.n1963 vdd.n847 10.6151
R18835 vdd.n1963 vdd.n1962 10.6151
R18836 vdd.n1962 vdd.n1961 10.6151
R18837 vdd.n1961 vdd.n849 10.6151
R18838 vdd.n1955 vdd.n849 10.6151
R18839 vdd.n1955 vdd.n1954 10.6151
R18840 vdd.n1954 vdd.n1953 10.6151
R18841 vdd.n1953 vdd.n853 10.6151
R18842 vdd.n1801 vdd.n853 10.6151
R18843 vdd.n1802 vdd.n1801 10.6151
R18844 vdd.n1802 vdd.n1797 10.6151
R18845 vdd.n1808 vdd.n1797 10.6151
R18846 vdd.n1809 vdd.n1808 10.6151
R18847 vdd.n1810 vdd.n1809 10.6151
R18848 vdd.n1810 vdd.n1795 10.6151
R18849 vdd.n1816 vdd.n1795 10.6151
R18850 vdd.n1817 vdd.n1816 10.6151
R18851 vdd.n1818 vdd.n1817 10.6151
R18852 vdd.n1818 vdd.n1793 10.6151
R18853 vdd.n1824 vdd.n1793 10.6151
R18854 vdd.n1825 vdd.n1824 10.6151
R18855 vdd.n1827 vdd.n1789 10.6151
R18856 vdd.n1832 vdd.n1789 10.6151
R18857 vdd.n280 vdd.n262 10.4732
R18858 vdd.n233 vdd.n215 10.4732
R18859 vdd.n190 vdd.n172 10.4732
R18860 vdd.n143 vdd.n125 10.4732
R18861 vdd.n101 vdd.n83 10.4732
R18862 vdd.n54 vdd.n36 10.4732
R18863 vdd.n1095 vdd.n1077 10.4732
R18864 vdd.n1142 vdd.n1124 10.4732
R18865 vdd.n1005 vdd.n987 10.4732
R18866 vdd.n1052 vdd.n1034 10.4732
R18867 vdd.n916 vdd.n898 10.4732
R18868 vdd.n963 vdd.n945 10.4732
R18869 vdd.t125 vdd.n888 10.3167
R18870 vdd.n2874 vdd.t145 10.3167
R18871 vdd.n1465 vdd.t121 10.09
R18872 vdd.n3042 vdd.t158 10.09
R18873 vdd.n279 vdd.n264 9.69747
R18874 vdd.n232 vdd.n217 9.69747
R18875 vdd.n189 vdd.n174 9.69747
R18876 vdd.n142 vdd.n127 9.69747
R18877 vdd.n100 vdd.n85 9.69747
R18878 vdd.n53 vdd.n38 9.69747
R18879 vdd.n1094 vdd.n1079 9.69747
R18880 vdd.n1141 vdd.n1126 9.69747
R18881 vdd.n1004 vdd.n989 9.69747
R18882 vdd.n1051 vdd.n1036 9.69747
R18883 vdd.n915 vdd.n900 9.69747
R18884 vdd.n962 vdd.n947 9.69747
R18885 vdd.n1929 vdd.n1928 9.67831
R18886 vdd.n2836 vdd.n520 9.67831
R18887 vdd.n2707 vdd.n2706 9.67831
R18888 vdd.n1953 vdd.n1952 9.67831
R18889 vdd.n295 vdd.n294 9.45567
R18890 vdd.n248 vdd.n247 9.45567
R18891 vdd.n205 vdd.n204 9.45567
R18892 vdd.n158 vdd.n157 9.45567
R18893 vdd.n116 vdd.n115 9.45567
R18894 vdd.n69 vdd.n68 9.45567
R18895 vdd.n1110 vdd.n1109 9.45567
R18896 vdd.n1157 vdd.n1156 9.45567
R18897 vdd.n1020 vdd.n1019 9.45567
R18898 vdd.n1067 vdd.n1066 9.45567
R18899 vdd.n931 vdd.n930 9.45567
R18900 vdd.n978 vdd.n977 9.45567
R18901 vdd.n1689 vdd.n1543 9.3005
R18902 vdd.n1688 vdd.n1687 9.3005
R18903 vdd.n1549 vdd.n1548 9.3005
R18904 vdd.n1682 vdd.n1553 9.3005
R18905 vdd.n1681 vdd.n1554 9.3005
R18906 vdd.n1680 vdd.n1555 9.3005
R18907 vdd.n1559 vdd.n1556 9.3005
R18908 vdd.n1675 vdd.n1560 9.3005
R18909 vdd.n1674 vdd.n1561 9.3005
R18910 vdd.n1673 vdd.n1562 9.3005
R18911 vdd.n1566 vdd.n1563 9.3005
R18912 vdd.n1668 vdd.n1567 9.3005
R18913 vdd.n1667 vdd.n1568 9.3005
R18914 vdd.n1666 vdd.n1569 9.3005
R18915 vdd.n1573 vdd.n1570 9.3005
R18916 vdd.n1661 vdd.n1574 9.3005
R18917 vdd.n1660 vdd.n1575 9.3005
R18918 vdd.n1659 vdd.n1576 9.3005
R18919 vdd.n1580 vdd.n1577 9.3005
R18920 vdd.n1654 vdd.n1581 9.3005
R18921 vdd.n1653 vdd.n1582 9.3005
R18922 vdd.n1652 vdd.n1651 9.3005
R18923 vdd.n1650 vdd.n1583 9.3005
R18924 vdd.n1649 vdd.n1648 9.3005
R18925 vdd.n1589 vdd.n1588 9.3005
R18926 vdd.n1643 vdd.n1593 9.3005
R18927 vdd.n1642 vdd.n1594 9.3005
R18928 vdd.n1641 vdd.n1595 9.3005
R18929 vdd.n1599 vdd.n1596 9.3005
R18930 vdd.n1636 vdd.n1600 9.3005
R18931 vdd.n1635 vdd.n1601 9.3005
R18932 vdd.n1634 vdd.n1602 9.3005
R18933 vdd.n1606 vdd.n1603 9.3005
R18934 vdd.n1629 vdd.n1607 9.3005
R18935 vdd.n1628 vdd.n1608 9.3005
R18936 vdd.n1627 vdd.n1609 9.3005
R18937 vdd.n1611 vdd.n1610 9.3005
R18938 vdd.n1622 vdd.n854 9.3005
R18939 vdd.n1691 vdd.n1690 9.3005
R18940 vdd.n1715 vdd.n1714 9.3005
R18941 vdd.n1521 vdd.n1520 9.3005
R18942 vdd.n1526 vdd.n1524 9.3005
R18943 vdd.n1707 vdd.n1527 9.3005
R18944 vdd.n1706 vdd.n1528 9.3005
R18945 vdd.n1705 vdd.n1529 9.3005
R18946 vdd.n1533 vdd.n1530 9.3005
R18947 vdd.n1700 vdd.n1534 9.3005
R18948 vdd.n1699 vdd.n1535 9.3005
R18949 vdd.n1698 vdd.n1536 9.3005
R18950 vdd.n1540 vdd.n1537 9.3005
R18951 vdd.n1693 vdd.n1541 9.3005
R18952 vdd.n1692 vdd.n1542 9.3005
R18953 vdd.n1937 vdd.n1514 9.3005
R18954 vdd.n1939 vdd.n1938 9.3005
R18955 vdd.n1476 vdd.n1475 9.3005
R18956 vdd.n1477 vdd.n890 9.3005
R18957 vdd.n1479 vdd.n1478 9.3005
R18958 vdd.n880 vdd.n879 9.3005
R18959 vdd.n1493 vdd.n1492 9.3005
R18960 vdd.n1494 vdd.n878 9.3005
R18961 vdd.n1496 vdd.n1495 9.3005
R18962 vdd.n868 vdd.n867 9.3005
R18963 vdd.n1512 vdd.n1511 9.3005
R18964 vdd.n1513 vdd.n866 9.3005
R18965 vdd.n1941 vdd.n1940 9.3005
R18966 vdd.n271 vdd.n270 9.3005
R18967 vdd.n266 vdd.n265 9.3005
R18968 vdd.n277 vdd.n276 9.3005
R18969 vdd.n279 vdd.n278 9.3005
R18970 vdd.n262 vdd.n261 9.3005
R18971 vdd.n285 vdd.n284 9.3005
R18972 vdd.n287 vdd.n286 9.3005
R18973 vdd.n259 vdd.n256 9.3005
R18974 vdd.n294 vdd.n293 9.3005
R18975 vdd.n224 vdd.n223 9.3005
R18976 vdd.n219 vdd.n218 9.3005
R18977 vdd.n230 vdd.n229 9.3005
R18978 vdd.n232 vdd.n231 9.3005
R18979 vdd.n215 vdd.n214 9.3005
R18980 vdd.n238 vdd.n237 9.3005
R18981 vdd.n240 vdd.n239 9.3005
R18982 vdd.n212 vdd.n209 9.3005
R18983 vdd.n247 vdd.n246 9.3005
R18984 vdd.n181 vdd.n180 9.3005
R18985 vdd.n176 vdd.n175 9.3005
R18986 vdd.n187 vdd.n186 9.3005
R18987 vdd.n189 vdd.n188 9.3005
R18988 vdd.n172 vdd.n171 9.3005
R18989 vdd.n195 vdd.n194 9.3005
R18990 vdd.n197 vdd.n196 9.3005
R18991 vdd.n169 vdd.n166 9.3005
R18992 vdd.n204 vdd.n203 9.3005
R18993 vdd.n134 vdd.n133 9.3005
R18994 vdd.n129 vdd.n128 9.3005
R18995 vdd.n140 vdd.n139 9.3005
R18996 vdd.n142 vdd.n141 9.3005
R18997 vdd.n125 vdd.n124 9.3005
R18998 vdd.n148 vdd.n147 9.3005
R18999 vdd.n150 vdd.n149 9.3005
R19000 vdd.n122 vdd.n119 9.3005
R19001 vdd.n157 vdd.n156 9.3005
R19002 vdd.n92 vdd.n91 9.3005
R19003 vdd.n87 vdd.n86 9.3005
R19004 vdd.n98 vdd.n97 9.3005
R19005 vdd.n100 vdd.n99 9.3005
R19006 vdd.n83 vdd.n82 9.3005
R19007 vdd.n106 vdd.n105 9.3005
R19008 vdd.n108 vdd.n107 9.3005
R19009 vdd.n80 vdd.n77 9.3005
R19010 vdd.n115 vdd.n114 9.3005
R19011 vdd.n45 vdd.n44 9.3005
R19012 vdd.n40 vdd.n39 9.3005
R19013 vdd.n51 vdd.n50 9.3005
R19014 vdd.n53 vdd.n52 9.3005
R19015 vdd.n36 vdd.n35 9.3005
R19016 vdd.n59 vdd.n58 9.3005
R19017 vdd.n61 vdd.n60 9.3005
R19018 vdd.n33 vdd.n30 9.3005
R19019 vdd.n68 vdd.n67 9.3005
R19020 vdd.n2758 vdd.n2757 9.3005
R19021 vdd.n2761 vdd.n555 9.3005
R19022 vdd.n2762 vdd.n554 9.3005
R19023 vdd.n2765 vdd.n553 9.3005
R19024 vdd.n2766 vdd.n552 9.3005
R19025 vdd.n2769 vdd.n551 9.3005
R19026 vdd.n2770 vdd.n550 9.3005
R19027 vdd.n2773 vdd.n549 9.3005
R19028 vdd.n2774 vdd.n548 9.3005
R19029 vdd.n2777 vdd.n547 9.3005
R19030 vdd.n2778 vdd.n546 9.3005
R19031 vdd.n2781 vdd.n545 9.3005
R19032 vdd.n2782 vdd.n544 9.3005
R19033 vdd.n2785 vdd.n543 9.3005
R19034 vdd.n2786 vdd.n542 9.3005
R19035 vdd.n2789 vdd.n541 9.3005
R19036 vdd.n2790 vdd.n540 9.3005
R19037 vdd.n2793 vdd.n539 9.3005
R19038 vdd.n2794 vdd.n538 9.3005
R19039 vdd.n2797 vdd.n537 9.3005
R19040 vdd.n2801 vdd.n2800 9.3005
R19041 vdd.n2802 vdd.n536 9.3005
R19042 vdd.n2806 vdd.n2803 9.3005
R19043 vdd.n2809 vdd.n535 9.3005
R19044 vdd.n2810 vdd.n534 9.3005
R19045 vdd.n2813 vdd.n533 9.3005
R19046 vdd.n2814 vdd.n532 9.3005
R19047 vdd.n2817 vdd.n531 9.3005
R19048 vdd.n2818 vdd.n530 9.3005
R19049 vdd.n2821 vdd.n529 9.3005
R19050 vdd.n2822 vdd.n528 9.3005
R19051 vdd.n2825 vdd.n527 9.3005
R19052 vdd.n2826 vdd.n526 9.3005
R19053 vdd.n2829 vdd.n525 9.3005
R19054 vdd.n2830 vdd.n524 9.3005
R19055 vdd.n2833 vdd.n519 9.3005
R19056 vdd.n482 vdd.n481 9.3005
R19057 vdd.n2844 vdd.n2843 9.3005
R19058 vdd.n2847 vdd.n2846 9.3005
R19059 vdd.n471 vdd.n470 9.3005
R19060 vdd.n2861 vdd.n2860 9.3005
R19061 vdd.n2862 vdd.n469 9.3005
R19062 vdd.n2864 vdd.n2863 9.3005
R19063 vdd.n460 vdd.n459 9.3005
R19064 vdd.n2877 vdd.n2876 9.3005
R19065 vdd.n2878 vdd.n458 9.3005
R19066 vdd.n2880 vdd.n2879 9.3005
R19067 vdd.n300 vdd.n298 9.3005
R19068 vdd.n2845 vdd.n480 9.3005
R19069 vdd.n3046 vdd.n3045 9.3005
R19070 vdd.n301 vdd.n299 9.3005
R19071 vdd.n3039 vdd.n310 9.3005
R19072 vdd.n3038 vdd.n311 9.3005
R19073 vdd.n3037 vdd.n312 9.3005
R19074 vdd.n320 vdd.n313 9.3005
R19075 vdd.n3031 vdd.n321 9.3005
R19076 vdd.n3030 vdd.n322 9.3005
R19077 vdd.n3029 vdd.n323 9.3005
R19078 vdd.n331 vdd.n324 9.3005
R19079 vdd.n3023 vdd.n3022 9.3005
R19080 vdd.n3019 vdd.n332 9.3005
R19081 vdd.n3018 vdd.n335 9.3005
R19082 vdd.n339 vdd.n336 9.3005
R19083 vdd.n340 vdd.n337 9.3005
R19084 vdd.n3011 vdd.n341 9.3005
R19085 vdd.n3010 vdd.n342 9.3005
R19086 vdd.n3009 vdd.n343 9.3005
R19087 vdd.n347 vdd.n344 9.3005
R19088 vdd.n3004 vdd.n348 9.3005
R19089 vdd.n3003 vdd.n349 9.3005
R19090 vdd.n3002 vdd.n350 9.3005
R19091 vdd.n354 vdd.n351 9.3005
R19092 vdd.n2997 vdd.n355 9.3005
R19093 vdd.n2996 vdd.n356 9.3005
R19094 vdd.n2995 vdd.n357 9.3005
R19095 vdd.n361 vdd.n358 9.3005
R19096 vdd.n2990 vdd.n362 9.3005
R19097 vdd.n2989 vdd.n363 9.3005
R19098 vdd.n2988 vdd.n2987 9.3005
R19099 vdd.n2986 vdd.n364 9.3005
R19100 vdd.n2985 vdd.n2984 9.3005
R19101 vdd.n370 vdd.n369 9.3005
R19102 vdd.n2979 vdd.n374 9.3005
R19103 vdd.n2978 vdd.n375 9.3005
R19104 vdd.n2977 vdd.n376 9.3005
R19105 vdd.n380 vdd.n377 9.3005
R19106 vdd.n2972 vdd.n381 9.3005
R19107 vdd.n2971 vdd.n382 9.3005
R19108 vdd.n2970 vdd.n383 9.3005
R19109 vdd.n387 vdd.n384 9.3005
R19110 vdd.n2965 vdd.n388 9.3005
R19111 vdd.n2964 vdd.n389 9.3005
R19112 vdd.n2963 vdd.n390 9.3005
R19113 vdd.n394 vdd.n391 9.3005
R19114 vdd.n2958 vdd.n395 9.3005
R19115 vdd.n2957 vdd.n396 9.3005
R19116 vdd.n2956 vdd.n397 9.3005
R19117 vdd.n401 vdd.n398 9.3005
R19118 vdd.n2951 vdd.n402 9.3005
R19119 vdd.n2950 vdd.n403 9.3005
R19120 vdd.n2949 vdd.n2948 9.3005
R19121 vdd.n2947 vdd.n404 9.3005
R19122 vdd.n2946 vdd.n2945 9.3005
R19123 vdd.n410 vdd.n409 9.3005
R19124 vdd.n2940 vdd.n414 9.3005
R19125 vdd.n2939 vdd.n415 9.3005
R19126 vdd.n2938 vdd.n416 9.3005
R19127 vdd.n420 vdd.n417 9.3005
R19128 vdd.n2933 vdd.n421 9.3005
R19129 vdd.n2932 vdd.n422 9.3005
R19130 vdd.n2931 vdd.n423 9.3005
R19131 vdd.n427 vdd.n424 9.3005
R19132 vdd.n2926 vdd.n428 9.3005
R19133 vdd.n2925 vdd.n429 9.3005
R19134 vdd.n2924 vdd.n430 9.3005
R19135 vdd.n434 vdd.n431 9.3005
R19136 vdd.n2919 vdd.n435 9.3005
R19137 vdd.n2918 vdd.n436 9.3005
R19138 vdd.n2917 vdd.n437 9.3005
R19139 vdd.n441 vdd.n438 9.3005
R19140 vdd.n2912 vdd.n442 9.3005
R19141 vdd.n2911 vdd.n443 9.3005
R19142 vdd.n2907 vdd.n2904 9.3005
R19143 vdd.n3021 vdd.n3020 9.3005
R19144 vdd.n2852 vdd.n2851 9.3005
R19145 vdd.n2853 vdd.n475 9.3005
R19146 vdd.n2855 vdd.n2854 9.3005
R19147 vdd.n465 vdd.n464 9.3005
R19148 vdd.n2869 vdd.n2868 9.3005
R19149 vdd.n2870 vdd.n463 9.3005
R19150 vdd.n2872 vdd.n2871 9.3005
R19151 vdd.n453 vdd.n452 9.3005
R19152 vdd.n2885 vdd.n2884 9.3005
R19153 vdd.n2886 vdd.n451 9.3005
R19154 vdd.n2888 vdd.n2887 9.3005
R19155 vdd.n2889 vdd.n450 9.3005
R19156 vdd.n2891 vdd.n2890 9.3005
R19157 vdd.n2892 vdd.n449 9.3005
R19158 vdd.n2894 vdd.n2893 9.3005
R19159 vdd.n2895 vdd.n447 9.3005
R19160 vdd.n2897 vdd.n2896 9.3005
R19161 vdd.n2898 vdd.n446 9.3005
R19162 vdd.n2900 vdd.n2899 9.3005
R19163 vdd.n2901 vdd.n444 9.3005
R19164 vdd.n2903 vdd.n2902 9.3005
R19165 vdd.n477 vdd.n476 9.3005
R19166 vdd.n2710 vdd.n2709 9.3005
R19167 vdd.n2715 vdd.n2708 9.3005
R19168 vdd.n2724 vdd.n572 9.3005
R19169 vdd.n2727 vdd.n571 9.3005
R19170 vdd.n2728 vdd.n570 9.3005
R19171 vdd.n2731 vdd.n569 9.3005
R19172 vdd.n2732 vdd.n568 9.3005
R19173 vdd.n2735 vdd.n567 9.3005
R19174 vdd.n2736 vdd.n566 9.3005
R19175 vdd.n2739 vdd.n565 9.3005
R19176 vdd.n2740 vdd.n564 9.3005
R19177 vdd.n2743 vdd.n563 9.3005
R19178 vdd.n2744 vdd.n562 9.3005
R19179 vdd.n2747 vdd.n561 9.3005
R19180 vdd.n2748 vdd.n560 9.3005
R19181 vdd.n2751 vdd.n559 9.3005
R19182 vdd.n2755 vdd.n2754 9.3005
R19183 vdd.n2756 vdd.n556 9.3005
R19184 vdd.n1951 vdd.n1950 9.3005
R19185 vdd.n1946 vdd.n857 9.3005
R19186 vdd.n1433 vdd.n1432 9.3005
R19187 vdd.n1434 vdd.n1188 9.3005
R19188 vdd.n1436 vdd.n1435 9.3005
R19189 vdd.n1178 vdd.n1177 9.3005
R19190 vdd.n1450 vdd.n1449 9.3005
R19191 vdd.n1451 vdd.n1176 9.3005
R19192 vdd.n1453 vdd.n1452 9.3005
R19193 vdd.n1168 vdd.n1167 9.3005
R19194 vdd.n1468 vdd.n1467 9.3005
R19195 vdd.n1469 vdd.n1166 9.3005
R19196 vdd.n1471 vdd.n1470 9.3005
R19197 vdd.n885 vdd.n884 9.3005
R19198 vdd.n1484 vdd.n1483 9.3005
R19199 vdd.n1485 vdd.n883 9.3005
R19200 vdd.n1487 vdd.n1486 9.3005
R19201 vdd.n875 vdd.n874 9.3005
R19202 vdd.n1501 vdd.n1500 9.3005
R19203 vdd.n1502 vdd.n872 9.3005
R19204 vdd.n1506 vdd.n1505 9.3005
R19205 vdd.n1504 vdd.n873 9.3005
R19206 vdd.n1503 vdd.n862 9.3005
R19207 vdd.n1190 vdd.n1189 9.3005
R19208 vdd.n1326 vdd.n1325 9.3005
R19209 vdd.n1327 vdd.n1316 9.3005
R19210 vdd.n1329 vdd.n1328 9.3005
R19211 vdd.n1330 vdd.n1315 9.3005
R19212 vdd.n1332 vdd.n1331 9.3005
R19213 vdd.n1333 vdd.n1310 9.3005
R19214 vdd.n1335 vdd.n1334 9.3005
R19215 vdd.n1336 vdd.n1309 9.3005
R19216 vdd.n1338 vdd.n1337 9.3005
R19217 vdd.n1339 vdd.n1304 9.3005
R19218 vdd.n1341 vdd.n1340 9.3005
R19219 vdd.n1342 vdd.n1303 9.3005
R19220 vdd.n1344 vdd.n1343 9.3005
R19221 vdd.n1345 vdd.n1298 9.3005
R19222 vdd.n1347 vdd.n1346 9.3005
R19223 vdd.n1348 vdd.n1297 9.3005
R19224 vdd.n1350 vdd.n1349 9.3005
R19225 vdd.n1351 vdd.n1292 9.3005
R19226 vdd.n1353 vdd.n1352 9.3005
R19227 vdd.n1354 vdd.n1291 9.3005
R19228 vdd.n1356 vdd.n1355 9.3005
R19229 vdd.n1360 vdd.n1287 9.3005
R19230 vdd.n1362 vdd.n1361 9.3005
R19231 vdd.n1363 vdd.n1286 9.3005
R19232 vdd.n1365 vdd.n1364 9.3005
R19233 vdd.n1366 vdd.n1281 9.3005
R19234 vdd.n1368 vdd.n1367 9.3005
R19235 vdd.n1369 vdd.n1280 9.3005
R19236 vdd.n1371 vdd.n1370 9.3005
R19237 vdd.n1372 vdd.n1275 9.3005
R19238 vdd.n1374 vdd.n1373 9.3005
R19239 vdd.n1375 vdd.n1274 9.3005
R19240 vdd.n1377 vdd.n1376 9.3005
R19241 vdd.n1378 vdd.n1269 9.3005
R19242 vdd.n1380 vdd.n1379 9.3005
R19243 vdd.n1381 vdd.n1268 9.3005
R19244 vdd.n1383 vdd.n1382 9.3005
R19245 vdd.n1384 vdd.n1263 9.3005
R19246 vdd.n1386 vdd.n1385 9.3005
R19247 vdd.n1387 vdd.n1262 9.3005
R19248 vdd.n1389 vdd.n1388 9.3005
R19249 vdd.n1390 vdd.n1257 9.3005
R19250 vdd.n1392 vdd.n1391 9.3005
R19251 vdd.n1393 vdd.n1256 9.3005
R19252 vdd.n1395 vdd.n1394 9.3005
R19253 vdd.n1396 vdd.n1249 9.3005
R19254 vdd.n1398 vdd.n1397 9.3005
R19255 vdd.n1399 vdd.n1248 9.3005
R19256 vdd.n1401 vdd.n1400 9.3005
R19257 vdd.n1402 vdd.n1243 9.3005
R19258 vdd.n1404 vdd.n1403 9.3005
R19259 vdd.n1405 vdd.n1242 9.3005
R19260 vdd.n1407 vdd.n1406 9.3005
R19261 vdd.n1408 vdd.n1237 9.3005
R19262 vdd.n1410 vdd.n1409 9.3005
R19263 vdd.n1411 vdd.n1236 9.3005
R19264 vdd.n1413 vdd.n1412 9.3005
R19265 vdd.n1414 vdd.n1231 9.3005
R19266 vdd.n1416 vdd.n1415 9.3005
R19267 vdd.n1417 vdd.n1230 9.3005
R19268 vdd.n1419 vdd.n1418 9.3005
R19269 vdd.n1195 vdd.n1194 9.3005
R19270 vdd.n1425 vdd.n1424 9.3005
R19271 vdd.n1324 vdd.n1323 9.3005
R19272 vdd.n1428 vdd.n1427 9.3005
R19273 vdd.n1184 vdd.n1183 9.3005
R19274 vdd.n1442 vdd.n1441 9.3005
R19275 vdd.n1443 vdd.n1182 9.3005
R19276 vdd.n1445 vdd.n1444 9.3005
R19277 vdd.n1173 vdd.n1172 9.3005
R19278 vdd.n1459 vdd.n1458 9.3005
R19279 vdd.n1460 vdd.n1171 9.3005
R19280 vdd.n1463 vdd.n1462 9.3005
R19281 vdd.n1461 vdd.n1162 9.3005
R19282 vdd.n1426 vdd.n1193 9.3005
R19283 vdd.n1086 vdd.n1085 9.3005
R19284 vdd.n1081 vdd.n1080 9.3005
R19285 vdd.n1092 vdd.n1091 9.3005
R19286 vdd.n1094 vdd.n1093 9.3005
R19287 vdd.n1077 vdd.n1076 9.3005
R19288 vdd.n1100 vdd.n1099 9.3005
R19289 vdd.n1102 vdd.n1101 9.3005
R19290 vdd.n1074 vdd.n1071 9.3005
R19291 vdd.n1109 vdd.n1108 9.3005
R19292 vdd.n1133 vdd.n1132 9.3005
R19293 vdd.n1128 vdd.n1127 9.3005
R19294 vdd.n1139 vdd.n1138 9.3005
R19295 vdd.n1141 vdd.n1140 9.3005
R19296 vdd.n1124 vdd.n1123 9.3005
R19297 vdd.n1147 vdd.n1146 9.3005
R19298 vdd.n1149 vdd.n1148 9.3005
R19299 vdd.n1121 vdd.n1118 9.3005
R19300 vdd.n1156 vdd.n1155 9.3005
R19301 vdd.n996 vdd.n995 9.3005
R19302 vdd.n991 vdd.n990 9.3005
R19303 vdd.n1002 vdd.n1001 9.3005
R19304 vdd.n1004 vdd.n1003 9.3005
R19305 vdd.n987 vdd.n986 9.3005
R19306 vdd.n1010 vdd.n1009 9.3005
R19307 vdd.n1012 vdd.n1011 9.3005
R19308 vdd.n984 vdd.n981 9.3005
R19309 vdd.n1019 vdd.n1018 9.3005
R19310 vdd.n1043 vdd.n1042 9.3005
R19311 vdd.n1038 vdd.n1037 9.3005
R19312 vdd.n1049 vdd.n1048 9.3005
R19313 vdd.n1051 vdd.n1050 9.3005
R19314 vdd.n1034 vdd.n1033 9.3005
R19315 vdd.n1057 vdd.n1056 9.3005
R19316 vdd.n1059 vdd.n1058 9.3005
R19317 vdd.n1031 vdd.n1028 9.3005
R19318 vdd.n1066 vdd.n1065 9.3005
R19319 vdd.n907 vdd.n906 9.3005
R19320 vdd.n902 vdd.n901 9.3005
R19321 vdd.n913 vdd.n912 9.3005
R19322 vdd.n915 vdd.n914 9.3005
R19323 vdd.n898 vdd.n897 9.3005
R19324 vdd.n921 vdd.n920 9.3005
R19325 vdd.n923 vdd.n922 9.3005
R19326 vdd.n895 vdd.n892 9.3005
R19327 vdd.n930 vdd.n929 9.3005
R19328 vdd.n954 vdd.n953 9.3005
R19329 vdd.n949 vdd.n948 9.3005
R19330 vdd.n960 vdd.n959 9.3005
R19331 vdd.n962 vdd.n961 9.3005
R19332 vdd.n945 vdd.n944 9.3005
R19333 vdd.n968 vdd.n967 9.3005
R19334 vdd.n970 vdd.n969 9.3005
R19335 vdd.n942 vdd.n939 9.3005
R19336 vdd.n977 vdd.n976 9.3005
R19337 vdd.n1438 vdd.t154 8.95635
R19338 vdd.t136 vdd.n3033 8.95635
R19339 vdd.n276 vdd.n275 8.92171
R19340 vdd.n229 vdd.n228 8.92171
R19341 vdd.n186 vdd.n185 8.92171
R19342 vdd.n139 vdd.n138 8.92171
R19343 vdd.n97 vdd.n96 8.92171
R19344 vdd.n50 vdd.n49 8.92171
R19345 vdd.n1091 vdd.n1090 8.92171
R19346 vdd.n1138 vdd.n1137 8.92171
R19347 vdd.n1001 vdd.n1000 8.92171
R19348 vdd.n1048 vdd.n1047 8.92171
R19349 vdd.n912 vdd.n911 8.92171
R19350 vdd.n959 vdd.n958 8.92171
R19351 vdd.n207 vdd.n117 8.81535
R19352 vdd.n1069 vdd.n979 8.81535
R19353 vdd.n1465 vdd.t132 8.72962
R19354 vdd.t134 vdd.n3042 8.72962
R19355 vdd.n888 vdd.t170 8.50289
R19356 vdd.n1943 vdd.t49 8.50289
R19357 vdd.n516 vdd.t42 8.50289
R19358 vdd.n2874 vdd.t148 8.50289
R19359 vdd.n28 vdd.n14 8.42249
R19360 vdd.n3048 vdd.n3047 8.16225
R19361 vdd.n1161 vdd.n1160 8.16225
R19362 vdd.n272 vdd.n266 8.14595
R19363 vdd.n225 vdd.n219 8.14595
R19364 vdd.n182 vdd.n176 8.14595
R19365 vdd.n135 vdd.n129 8.14595
R19366 vdd.n93 vdd.n87 8.14595
R19367 vdd.n46 vdd.n40 8.14595
R19368 vdd.n1087 vdd.n1081 8.14595
R19369 vdd.n1134 vdd.n1128 8.14595
R19370 vdd.n997 vdd.n991 8.14595
R19371 vdd.n1044 vdd.n1038 8.14595
R19372 vdd.n908 vdd.n902 8.14595
R19373 vdd.n955 vdd.n949 8.14595
R19374 vdd.n2537 vdd.n639 8.11757
R19375 vdd.n2011 vdd.n2010 8.11757
R19376 vdd.n1989 vdd.n833 7.70933
R19377 vdd.n1995 vdd.n833 7.70933
R19378 vdd.n2001 vdd.n827 7.70933
R19379 vdd.n2001 vdd.n820 7.70933
R19380 vdd.n2007 vdd.n820 7.70933
R19381 vdd.n2007 vdd.n823 7.70933
R19382 vdd.n2014 vdd.n808 7.70933
R19383 vdd.n2020 vdd.n808 7.70933
R19384 vdd.n2026 vdd.n802 7.70933
R19385 vdd.n2032 vdd.n798 7.70933
R19386 vdd.n2038 vdd.n792 7.70933
R19387 vdd.n2050 vdd.n779 7.70933
R19388 vdd.n2056 vdd.n773 7.70933
R19389 vdd.n2056 vdd.n766 7.70933
R19390 vdd.n2064 vdd.n766 7.70933
R19391 vdd.n2071 vdd.t188 7.70933
R19392 vdd.n2146 vdd.t188 7.70933
R19393 vdd.n2478 vdd.t190 7.70933
R19394 vdd.n2484 vdd.t190 7.70933
R19395 vdd.n2490 vdd.n687 7.70933
R19396 vdd.n2496 vdd.n687 7.70933
R19397 vdd.n2496 vdd.n690 7.70933
R19398 vdd.n2502 vdd.n683 7.70933
R19399 vdd.n2514 vdd.n670 7.70933
R19400 vdd.n2520 vdd.n664 7.70933
R19401 vdd.n2526 vdd.n660 7.70933
R19402 vdd.n2532 vdd.n647 7.70933
R19403 vdd.n2540 vdd.n647 7.70933
R19404 vdd.n2546 vdd.n641 7.70933
R19405 vdd.n2546 vdd.n633 7.70933
R19406 vdd.n2597 vdd.n633 7.70933
R19407 vdd.n2597 vdd.n636 7.70933
R19408 vdd.n2603 vdd.n595 7.70933
R19409 vdd.n2673 vdd.n595 7.70933
R19410 vdd.n271 vdd.n268 7.3702
R19411 vdd.n224 vdd.n221 7.3702
R19412 vdd.n181 vdd.n178 7.3702
R19413 vdd.n134 vdd.n131 7.3702
R19414 vdd.n92 vdd.n89 7.3702
R19415 vdd.n45 vdd.n42 7.3702
R19416 vdd.n1086 vdd.n1083 7.3702
R19417 vdd.n1133 vdd.n1130 7.3702
R19418 vdd.n996 vdd.n993 7.3702
R19419 vdd.n1043 vdd.n1040 7.3702
R19420 vdd.n907 vdd.n904 7.3702
R19421 vdd.n954 vdd.n951 7.3702
R19422 vdd.n1361 vdd.n1360 6.98232
R19423 vdd.n1653 vdd.n1652 6.98232
R19424 vdd.n2950 vdd.n2949 6.98232
R19425 vdd.n2761 vdd.n2758 6.98232
R19426 vdd.n1498 vdd.t117 6.68904
R19427 vdd.n2857 vdd.t119 6.68904
R19428 vdd.t156 vdd.n887 6.46231
R19429 vdd.n2882 vdd.t123 6.46231
R19430 vdd.n1456 vdd.t138 6.23558
R19431 vdd.t127 vdd.n308 6.23558
R19432 vdd.n3048 vdd.n297 6.22547
R19433 vdd.n1160 vdd.n1159 6.22547
R19434 vdd.n2026 vdd.t29 6.00885
R19435 vdd.n2526 vdd.t187 6.00885
R19436 vdd.n823 vdd.t93 5.89549
R19437 vdd.t57 vdd.n641 5.89549
R19438 vdd.n272 vdd.n271 5.81868
R19439 vdd.n225 vdd.n224 5.81868
R19440 vdd.n182 vdd.n181 5.81868
R19441 vdd.n135 vdd.n134 5.81868
R19442 vdd.n93 vdd.n92 5.81868
R19443 vdd.n46 vdd.n45 5.81868
R19444 vdd.n1087 vdd.n1086 5.81868
R19445 vdd.n1134 vdd.n1133 5.81868
R19446 vdd.n997 vdd.n996 5.81868
R19447 vdd.n1044 vdd.n1043 5.81868
R19448 vdd.n908 vdd.n907 5.81868
R19449 vdd.n955 vdd.n954 5.81868
R19450 vdd.t89 vdd.n827 5.78212
R19451 vdd.n1770 vdd.t74 5.78212
R19452 vdd.n2395 vdd.t82 5.78212
R19453 vdd.n636 vdd.t78 5.78212
R19454 vdd.n2154 vdd.n2153 5.77611
R19455 vdd.n1897 vdd.n1767 5.77611
R19456 vdd.n2408 vdd.n2407 5.77611
R19457 vdd.n2614 vdd.n2613 5.77611
R19458 vdd.n2678 vdd.n591 5.77611
R19459 vdd.n2318 vdd.n2258 5.77611
R19460 vdd.n2079 vdd.n757 5.77611
R19461 vdd.n1827 vdd.n1826 5.77611
R19462 vdd.n1323 vdd.n1322 5.62474
R19463 vdd.n1949 vdd.n1946 5.62474
R19464 vdd.n2910 vdd.n2907 5.62474
R19465 vdd.n2713 vdd.n2710 5.62474
R19466 vdd.t25 vdd.n779 5.44203
R19467 vdd.n683 vdd.t18 5.44203
R19468 vdd.n1180 vdd.t138 5.10193
R19469 vdd.t24 vdd.n802 5.10193
R19470 vdd.n792 vdd.t196 5.10193
R19471 vdd.t197 vdd.n670 5.10193
R19472 vdd.n660 vdd.t34 5.10193
R19473 vdd.n3035 vdd.t127 5.10193
R19474 vdd.n275 vdd.n266 5.04292
R19475 vdd.n228 vdd.n219 5.04292
R19476 vdd.n185 vdd.n176 5.04292
R19477 vdd.n138 vdd.n129 5.04292
R19478 vdd.n96 vdd.n87 5.04292
R19479 vdd.n49 vdd.n40 5.04292
R19480 vdd.n1090 vdd.n1081 5.04292
R19481 vdd.n1137 vdd.n1128 5.04292
R19482 vdd.n1000 vdd.n991 5.04292
R19483 vdd.n1047 vdd.n1038 5.04292
R19484 vdd.n911 vdd.n902 5.04292
R19485 vdd.n958 vdd.n949 5.04292
R19486 vdd.n1473 vdd.t156 4.8752
R19487 vdd.t20 vdd.t185 4.8752
R19488 vdd.t30 vdd.t198 4.8752
R19489 vdd.t194 vdd.t33 4.8752
R19490 vdd.t27 vdd.t35 4.8752
R19491 vdd.t123 vdd.n304 4.8752
R19492 vdd.n2155 vdd.n2154 4.83952
R19493 vdd.n1767 vdd.n1763 4.83952
R19494 vdd.n2409 vdd.n2408 4.83952
R19495 vdd.n2615 vdd.n2614 4.83952
R19496 vdd.n591 vdd.n586 4.83952
R19497 vdd.n2315 vdd.n2258 4.83952
R19498 vdd.n2082 vdd.n757 4.83952
R19499 vdd.n1826 vdd.n1825 4.83952
R19500 vdd.n1621 vdd.n855 4.74817
R19501 vdd.n1616 vdd.n856 4.74817
R19502 vdd.n1518 vdd.n1515 4.74817
R19503 vdd.n1930 vdd.n1519 4.74817
R19504 vdd.n1932 vdd.n1518 4.74817
R19505 vdd.n1931 vdd.n1930 4.74817
R19506 vdd.n2838 vdd.n2837 4.74817
R19507 vdd.n2835 vdd.n2834 4.74817
R19508 vdd.n2835 vdd.n521 4.74817
R19509 vdd.n2837 vdd.n518 4.74817
R19510 vdd.n2720 vdd.n573 4.74817
R19511 vdd.n2716 vdd.n574 4.74817
R19512 vdd.n2719 vdd.n574 4.74817
R19513 vdd.n2723 vdd.n573 4.74817
R19514 vdd.n1617 vdd.n855 4.74817
R19515 vdd.n858 vdd.n856 4.74817
R19516 vdd.n297 vdd.n296 4.7074
R19517 vdd.n207 vdd.n206 4.7074
R19518 vdd.n1159 vdd.n1158 4.7074
R19519 vdd.n1069 vdd.n1068 4.7074
R19520 vdd.n1489 vdd.t117 4.64847
R19521 vdd.n2866 vdd.t119 4.64847
R19522 vdd.n2032 vdd.t21 4.53511
R19523 vdd.n2520 vdd.t183 4.53511
R19524 vdd.n2064 vdd.t181 4.30838
R19525 vdd.n2490 vdd.t31 4.30838
R19526 vdd.n276 vdd.n264 4.26717
R19527 vdd.n229 vdd.n217 4.26717
R19528 vdd.n186 vdd.n174 4.26717
R19529 vdd.n139 vdd.n127 4.26717
R19530 vdd.n97 vdd.n85 4.26717
R19531 vdd.n50 vdd.n38 4.26717
R19532 vdd.n1091 vdd.n1079 4.26717
R19533 vdd.n1138 vdd.n1126 4.26717
R19534 vdd.n1001 vdd.n989 4.26717
R19535 vdd.n1048 vdd.n1036 4.26717
R19536 vdd.n912 vdd.n900 4.26717
R19537 vdd.n959 vdd.n947 4.26717
R19538 vdd.n297 vdd.n207 4.10845
R19539 vdd.n1159 vdd.n1069 4.10845
R19540 vdd.n253 vdd.t164 4.06363
R19541 vdd.n253 vdd.t128 4.06363
R19542 vdd.n251 vdd.t130 4.06363
R19543 vdd.n251 vdd.t151 4.06363
R19544 vdd.n249 vdd.t153 4.06363
R19545 vdd.n249 vdd.t169 4.06363
R19546 vdd.n163 vdd.t159 4.06363
R19547 vdd.n163 vdd.t180 4.06363
R19548 vdd.n161 vdd.t124 4.06363
R19549 vdd.n161 vdd.t143 4.06363
R19550 vdd.n159 vdd.t149 4.06363
R19551 vdd.n159 vdd.t160 4.06363
R19552 vdd.n74 vdd.t165 4.06363
R19553 vdd.n74 vdd.t140 4.06363
R19554 vdd.n72 vdd.t179 4.06363
R19555 vdd.n72 vdd.t135 4.06363
R19556 vdd.n70 vdd.t172 4.06363
R19557 vdd.n70 vdd.t146 4.06363
R19558 vdd.n1111 vdd.t131 4.06363
R19559 vdd.n1111 vdd.t175 4.06363
R19560 vdd.n1113 vdd.t174 4.06363
R19561 vdd.n1113 vdd.t163 4.06363
R19562 vdd.n1115 vdd.t150 4.06363
R19563 vdd.n1115 vdd.t129 4.06363
R19564 vdd.n1021 vdd.t126 4.06363
R19565 vdd.n1021 vdd.t171 4.06363
R19566 vdd.n1023 vdd.t166 4.06363
R19567 vdd.n1023 vdd.t157 4.06363
R19568 vdd.n1025 vdd.t142 4.06363
R19569 vdd.n1025 vdd.t122 4.06363
R19570 vdd.n932 vdd.t144 4.06363
R19571 vdd.n932 vdd.t173 4.06363
R19572 vdd.n934 vdd.t133 4.06363
R19573 vdd.n934 vdd.t161 4.06363
R19574 vdd.n936 vdd.t139 4.06363
R19575 vdd.n936 vdd.t167 4.06363
R19576 vdd.n26 vdd.t3 3.9605
R19577 vdd.n26 vdd.t11 3.9605
R19578 vdd.n23 vdd.t13 3.9605
R19579 vdd.n23 vdd.t6 3.9605
R19580 vdd.n21 vdd.t4 3.9605
R19581 vdd.n21 vdd.t2 3.9605
R19582 vdd.n20 vdd.t12 3.9605
R19583 vdd.n20 vdd.t1 3.9605
R19584 vdd.n15 vdd.t5 3.9605
R19585 vdd.n15 vdd.t9 3.9605
R19586 vdd.n16 vdd.t7 3.9605
R19587 vdd.n16 vdd.t10 3.9605
R19588 vdd.n18 vdd.t14 3.9605
R19589 vdd.n18 vdd.t0 3.9605
R19590 vdd.n25 vdd.t8 3.9605
R19591 vdd.n25 vdd.t15 3.9605
R19592 vdd.n7 vdd.t28 3.61217
R19593 vdd.n7 vdd.t184 3.61217
R19594 vdd.n8 vdd.t195 3.61217
R19595 vdd.n8 vdd.t19 3.61217
R19596 vdd.n10 vdd.t191 3.61217
R19597 vdd.n10 vdd.t32 3.61217
R19598 vdd.n12 vdd.t39 3.61217
R19599 vdd.n12 vdd.t193 3.61217
R19600 vdd.n5 vdd.t17 3.61217
R19601 vdd.n5 vdd.t37 3.61217
R19602 vdd.n3 vdd.t182 3.61217
R19603 vdd.n3 vdd.t189 3.61217
R19604 vdd.n1 vdd.t26 3.61217
R19605 vdd.n1 vdd.t199 3.61217
R19606 vdd.n0 vdd.t22 3.61217
R19607 vdd.n0 vdd.t186 3.61217
R19608 vdd.n280 vdd.n279 3.49141
R19609 vdd.n233 vdd.n232 3.49141
R19610 vdd.n190 vdd.n189 3.49141
R19611 vdd.n143 vdd.n142 3.49141
R19612 vdd.n101 vdd.n100 3.49141
R19613 vdd.n54 vdd.n53 3.49141
R19614 vdd.n1095 vdd.n1094 3.49141
R19615 vdd.n1142 vdd.n1141 3.49141
R19616 vdd.n1005 vdd.n1004 3.49141
R19617 vdd.n1052 vdd.n1051 3.49141
R19618 vdd.n916 vdd.n915 3.49141
R19619 vdd.n963 vdd.n962 3.49141
R19620 vdd.n1770 vdd.t181 3.40145
R19621 vdd.n2218 vdd.t16 3.40145
R19622 vdd.n2471 vdd.t192 3.40145
R19623 vdd.n2395 vdd.t31 3.40145
R19624 vdd.n1871 vdd.t21 3.17472
R19625 vdd.n2374 vdd.t183 3.17472
R19626 vdd.n1490 vdd.t170 2.83463
R19627 vdd.n1508 vdd.t49 2.83463
R19628 vdd.n2849 vdd.t42 2.83463
R19629 vdd.n467 vdd.t148 2.83463
R19630 vdd.n283 vdd.n262 2.71565
R19631 vdd.n236 vdd.n215 2.71565
R19632 vdd.n193 vdd.n172 2.71565
R19633 vdd.n146 vdd.n125 2.71565
R19634 vdd.n104 vdd.n83 2.71565
R19635 vdd.n57 vdd.n36 2.71565
R19636 vdd.n1098 vdd.n1077 2.71565
R19637 vdd.n1145 vdd.n1124 2.71565
R19638 vdd.n1008 vdd.n987 2.71565
R19639 vdd.n1055 vdd.n1034 2.71565
R19640 vdd.n919 vdd.n898 2.71565
R19641 vdd.n966 vdd.n945 2.71565
R19642 vdd.t132 vdd.n1164 2.6079
R19643 vdd.n2020 vdd.t24 2.6079
R19644 vdd.n2044 vdd.t196 2.6079
R19645 vdd.n2508 vdd.t197 2.6079
R19646 vdd.n2532 vdd.t34 2.6079
R19647 vdd.n3043 vdd.t134 2.6079
R19648 vdd.n2538 vdd.n2537 2.49806
R19649 vdd.n2012 vdd.n2011 2.49806
R19650 vdd.n270 vdd.n269 2.4129
R19651 vdd.n223 vdd.n222 2.4129
R19652 vdd.n180 vdd.n179 2.4129
R19653 vdd.n133 vdd.n132 2.4129
R19654 vdd.n91 vdd.n90 2.4129
R19655 vdd.n44 vdd.n43 2.4129
R19656 vdd.n1085 vdd.n1084 2.4129
R19657 vdd.n1132 vdd.n1131 2.4129
R19658 vdd.n995 vdd.n994 2.4129
R19659 vdd.n1042 vdd.n1041 2.4129
R19660 vdd.n906 vdd.n905 2.4129
R19661 vdd.n953 vdd.n952 2.4129
R19662 vdd.n1447 vdd.t154 2.38117
R19663 vdd.n3034 vdd.t136 2.38117
R19664 vdd.n1929 vdd.n1518 2.27742
R19665 vdd.n1930 vdd.n1929 2.27742
R19666 vdd.n2836 vdd.n2835 2.27742
R19667 vdd.n2837 vdd.n2836 2.27742
R19668 vdd.n2707 vdd.n574 2.27742
R19669 vdd.n2707 vdd.n573 2.27742
R19670 vdd.n1952 vdd.n855 2.27742
R19671 vdd.n1952 vdd.n856 2.27742
R19672 vdd.n2044 vdd.t25 2.2678
R19673 vdd.n2508 vdd.t18 2.2678
R19674 vdd.t198 vdd.n773 2.04107
R19675 vdd.n690 vdd.t194 2.04107
R19676 vdd.n284 vdd.n260 1.93989
R19677 vdd.n237 vdd.n213 1.93989
R19678 vdd.n194 vdd.n170 1.93989
R19679 vdd.n147 vdd.n123 1.93989
R19680 vdd.n105 vdd.n81 1.93989
R19681 vdd.n58 vdd.n34 1.93989
R19682 vdd.n1099 vdd.n1075 1.93989
R19683 vdd.n1146 vdd.n1122 1.93989
R19684 vdd.n1009 vdd.n985 1.93989
R19685 vdd.n1056 vdd.n1032 1.93989
R19686 vdd.n920 vdd.n896 1.93989
R19687 vdd.n967 vdd.n943 1.93989
R19688 vdd.n1995 vdd.t89 1.92771
R19689 vdd.n2071 vdd.t74 1.92771
R19690 vdd.n2484 vdd.t82 1.92771
R19691 vdd.n2603 vdd.t78 1.92771
R19692 vdd.n1871 vdd.t29 1.70098
R19693 vdd.n798 vdd.t20 1.70098
R19694 vdd.t35 vdd.n664 1.70098
R19695 vdd.n2374 vdd.t187 1.70098
R19696 vdd.n1455 vdd.t121 1.24752
R19697 vdd.t158 vdd.n3041 1.24752
R19698 vdd.n295 vdd.n255 1.16414
R19699 vdd.n288 vdd.n287 1.16414
R19700 vdd.n248 vdd.n208 1.16414
R19701 vdd.n241 vdd.n240 1.16414
R19702 vdd.n205 vdd.n165 1.16414
R19703 vdd.n198 vdd.n197 1.16414
R19704 vdd.n158 vdd.n118 1.16414
R19705 vdd.n151 vdd.n150 1.16414
R19706 vdd.n116 vdd.n76 1.16414
R19707 vdd.n109 vdd.n108 1.16414
R19708 vdd.n69 vdd.n29 1.16414
R19709 vdd.n62 vdd.n61 1.16414
R19710 vdd.n1110 vdd.n1070 1.16414
R19711 vdd.n1103 vdd.n1102 1.16414
R19712 vdd.n1157 vdd.n1117 1.16414
R19713 vdd.n1150 vdd.n1149 1.16414
R19714 vdd.n1020 vdd.n980 1.16414
R19715 vdd.n1013 vdd.n1012 1.16414
R19716 vdd.n1067 vdd.n1027 1.16414
R19717 vdd.n1060 vdd.n1059 1.16414
R19718 vdd.n931 vdd.n891 1.16414
R19719 vdd.n924 vdd.n923 1.16414
R19720 vdd.n978 vdd.n938 1.16414
R19721 vdd.n971 vdd.n970 1.16414
R19722 vdd.n2038 vdd.t185 1.13415
R19723 vdd.n2514 vdd.t27 1.13415
R19724 vdd.n1481 vdd.t125 1.02079
R19725 vdd.t93 vdd.t23 1.02079
R19726 vdd.t40 vdd.t57 1.02079
R19727 vdd.t145 vdd.n456 1.02079
R19728 vdd.n1326 vdd.n1322 0.970197
R19729 vdd.n1950 vdd.n1949 0.970197
R19730 vdd.n2911 vdd.n2910 0.970197
R19731 vdd.n2715 vdd.n2713 0.970197
R19732 vdd.n2014 vdd.t23 0.794056
R19733 vdd.n2050 vdd.t30 0.794056
R19734 vdd.n2502 vdd.t33 0.794056
R19735 vdd.n2540 vdd.t40 0.794056
R19736 vdd.n1160 vdd.n28 0.74827
R19737 vdd vdd.n3048 0.740437
R19738 vdd.n1430 vdd.t53 0.567326
R19739 vdd.n3026 vdd.t64 0.567326
R19740 vdd.n1940 vdd.n1939 0.537085
R19741 vdd.n2845 vdd.n2844 0.537085
R19742 vdd.n3022 vdd.n3021 0.537085
R19743 vdd.n2904 vdd.n2903 0.537085
R19744 vdd.n2709 vdd.n476 0.537085
R19745 vdd.n1503 vdd.n857 0.537085
R19746 vdd.n1324 vdd.n1189 0.537085
R19747 vdd.n1426 vdd.n1425 0.537085
R19748 vdd.n4 vdd.n2 0.459552
R19749 vdd.n11 vdd.n9 0.459552
R19750 vdd.n293 vdd.n292 0.388379
R19751 vdd.n259 vdd.n257 0.388379
R19752 vdd.n246 vdd.n245 0.388379
R19753 vdd.n212 vdd.n210 0.388379
R19754 vdd.n203 vdd.n202 0.388379
R19755 vdd.n169 vdd.n167 0.388379
R19756 vdd.n156 vdd.n155 0.388379
R19757 vdd.n122 vdd.n120 0.388379
R19758 vdd.n114 vdd.n113 0.388379
R19759 vdd.n80 vdd.n78 0.388379
R19760 vdd.n67 vdd.n66 0.388379
R19761 vdd.n33 vdd.n31 0.388379
R19762 vdd.n1108 vdd.n1107 0.388379
R19763 vdd.n1074 vdd.n1072 0.388379
R19764 vdd.n1155 vdd.n1154 0.388379
R19765 vdd.n1121 vdd.n1119 0.388379
R19766 vdd.n1018 vdd.n1017 0.388379
R19767 vdd.n984 vdd.n982 0.388379
R19768 vdd.n1065 vdd.n1064 0.388379
R19769 vdd.n1031 vdd.n1029 0.388379
R19770 vdd.n929 vdd.n928 0.388379
R19771 vdd.n895 vdd.n893 0.388379
R19772 vdd.n976 vdd.n975 0.388379
R19773 vdd.n942 vdd.n940 0.388379
R19774 vdd.n19 vdd.n17 0.387128
R19775 vdd.n24 vdd.n22 0.387128
R19776 vdd.n6 vdd.n4 0.358259
R19777 vdd.n13 vdd.n11 0.358259
R19778 vdd.n252 vdd.n250 0.358259
R19779 vdd.n254 vdd.n252 0.358259
R19780 vdd.n296 vdd.n254 0.358259
R19781 vdd.n162 vdd.n160 0.358259
R19782 vdd.n164 vdd.n162 0.358259
R19783 vdd.n206 vdd.n164 0.358259
R19784 vdd.n73 vdd.n71 0.358259
R19785 vdd.n75 vdd.n73 0.358259
R19786 vdd.n117 vdd.n75 0.358259
R19787 vdd.n1158 vdd.n1116 0.358259
R19788 vdd.n1116 vdd.n1114 0.358259
R19789 vdd.n1114 vdd.n1112 0.358259
R19790 vdd.n1068 vdd.n1026 0.358259
R19791 vdd.n1026 vdd.n1024 0.358259
R19792 vdd.n1024 vdd.n1022 0.358259
R19793 vdd.n979 vdd.n937 0.358259
R19794 vdd.n937 vdd.n935 0.358259
R19795 vdd.n935 vdd.n933 0.358259
R19796 vdd.n14 vdd.n6 0.334552
R19797 vdd.n14 vdd.n13 0.334552
R19798 vdd.n27 vdd.n19 0.21707
R19799 vdd.n27 vdd.n24 0.21707
R19800 vdd.n294 vdd.n256 0.155672
R19801 vdd.n286 vdd.n256 0.155672
R19802 vdd.n286 vdd.n285 0.155672
R19803 vdd.n285 vdd.n261 0.155672
R19804 vdd.n278 vdd.n261 0.155672
R19805 vdd.n278 vdd.n277 0.155672
R19806 vdd.n277 vdd.n265 0.155672
R19807 vdd.n270 vdd.n265 0.155672
R19808 vdd.n247 vdd.n209 0.155672
R19809 vdd.n239 vdd.n209 0.155672
R19810 vdd.n239 vdd.n238 0.155672
R19811 vdd.n238 vdd.n214 0.155672
R19812 vdd.n231 vdd.n214 0.155672
R19813 vdd.n231 vdd.n230 0.155672
R19814 vdd.n230 vdd.n218 0.155672
R19815 vdd.n223 vdd.n218 0.155672
R19816 vdd.n204 vdd.n166 0.155672
R19817 vdd.n196 vdd.n166 0.155672
R19818 vdd.n196 vdd.n195 0.155672
R19819 vdd.n195 vdd.n171 0.155672
R19820 vdd.n188 vdd.n171 0.155672
R19821 vdd.n188 vdd.n187 0.155672
R19822 vdd.n187 vdd.n175 0.155672
R19823 vdd.n180 vdd.n175 0.155672
R19824 vdd.n157 vdd.n119 0.155672
R19825 vdd.n149 vdd.n119 0.155672
R19826 vdd.n149 vdd.n148 0.155672
R19827 vdd.n148 vdd.n124 0.155672
R19828 vdd.n141 vdd.n124 0.155672
R19829 vdd.n141 vdd.n140 0.155672
R19830 vdd.n140 vdd.n128 0.155672
R19831 vdd.n133 vdd.n128 0.155672
R19832 vdd.n115 vdd.n77 0.155672
R19833 vdd.n107 vdd.n77 0.155672
R19834 vdd.n107 vdd.n106 0.155672
R19835 vdd.n106 vdd.n82 0.155672
R19836 vdd.n99 vdd.n82 0.155672
R19837 vdd.n99 vdd.n98 0.155672
R19838 vdd.n98 vdd.n86 0.155672
R19839 vdd.n91 vdd.n86 0.155672
R19840 vdd.n68 vdd.n30 0.155672
R19841 vdd.n60 vdd.n30 0.155672
R19842 vdd.n60 vdd.n59 0.155672
R19843 vdd.n59 vdd.n35 0.155672
R19844 vdd.n52 vdd.n35 0.155672
R19845 vdd.n52 vdd.n51 0.155672
R19846 vdd.n51 vdd.n39 0.155672
R19847 vdd.n44 vdd.n39 0.155672
R19848 vdd.n1109 vdd.n1071 0.155672
R19849 vdd.n1101 vdd.n1071 0.155672
R19850 vdd.n1101 vdd.n1100 0.155672
R19851 vdd.n1100 vdd.n1076 0.155672
R19852 vdd.n1093 vdd.n1076 0.155672
R19853 vdd.n1093 vdd.n1092 0.155672
R19854 vdd.n1092 vdd.n1080 0.155672
R19855 vdd.n1085 vdd.n1080 0.155672
R19856 vdd.n1156 vdd.n1118 0.155672
R19857 vdd.n1148 vdd.n1118 0.155672
R19858 vdd.n1148 vdd.n1147 0.155672
R19859 vdd.n1147 vdd.n1123 0.155672
R19860 vdd.n1140 vdd.n1123 0.155672
R19861 vdd.n1140 vdd.n1139 0.155672
R19862 vdd.n1139 vdd.n1127 0.155672
R19863 vdd.n1132 vdd.n1127 0.155672
R19864 vdd.n1019 vdd.n981 0.155672
R19865 vdd.n1011 vdd.n981 0.155672
R19866 vdd.n1011 vdd.n1010 0.155672
R19867 vdd.n1010 vdd.n986 0.155672
R19868 vdd.n1003 vdd.n986 0.155672
R19869 vdd.n1003 vdd.n1002 0.155672
R19870 vdd.n1002 vdd.n990 0.155672
R19871 vdd.n995 vdd.n990 0.155672
R19872 vdd.n1066 vdd.n1028 0.155672
R19873 vdd.n1058 vdd.n1028 0.155672
R19874 vdd.n1058 vdd.n1057 0.155672
R19875 vdd.n1057 vdd.n1033 0.155672
R19876 vdd.n1050 vdd.n1033 0.155672
R19877 vdd.n1050 vdd.n1049 0.155672
R19878 vdd.n1049 vdd.n1037 0.155672
R19879 vdd.n1042 vdd.n1037 0.155672
R19880 vdd.n930 vdd.n892 0.155672
R19881 vdd.n922 vdd.n892 0.155672
R19882 vdd.n922 vdd.n921 0.155672
R19883 vdd.n921 vdd.n897 0.155672
R19884 vdd.n914 vdd.n897 0.155672
R19885 vdd.n914 vdd.n913 0.155672
R19886 vdd.n913 vdd.n901 0.155672
R19887 vdd.n906 vdd.n901 0.155672
R19888 vdd.n977 vdd.n939 0.155672
R19889 vdd.n969 vdd.n939 0.155672
R19890 vdd.n969 vdd.n968 0.155672
R19891 vdd.n968 vdd.n944 0.155672
R19892 vdd.n961 vdd.n944 0.155672
R19893 vdd.n961 vdd.n960 0.155672
R19894 vdd.n960 vdd.n948 0.155672
R19895 vdd.n953 vdd.n948 0.155672
R19896 vdd.n1715 vdd.n1520 0.152939
R19897 vdd.n1526 vdd.n1520 0.152939
R19898 vdd.n1527 vdd.n1526 0.152939
R19899 vdd.n1528 vdd.n1527 0.152939
R19900 vdd.n1529 vdd.n1528 0.152939
R19901 vdd.n1533 vdd.n1529 0.152939
R19902 vdd.n1534 vdd.n1533 0.152939
R19903 vdd.n1535 vdd.n1534 0.152939
R19904 vdd.n1536 vdd.n1535 0.152939
R19905 vdd.n1540 vdd.n1536 0.152939
R19906 vdd.n1541 vdd.n1540 0.152939
R19907 vdd.n1542 vdd.n1541 0.152939
R19908 vdd.n1690 vdd.n1542 0.152939
R19909 vdd.n1690 vdd.n1689 0.152939
R19910 vdd.n1689 vdd.n1688 0.152939
R19911 vdd.n1688 vdd.n1548 0.152939
R19912 vdd.n1553 vdd.n1548 0.152939
R19913 vdd.n1554 vdd.n1553 0.152939
R19914 vdd.n1555 vdd.n1554 0.152939
R19915 vdd.n1559 vdd.n1555 0.152939
R19916 vdd.n1560 vdd.n1559 0.152939
R19917 vdd.n1561 vdd.n1560 0.152939
R19918 vdd.n1562 vdd.n1561 0.152939
R19919 vdd.n1566 vdd.n1562 0.152939
R19920 vdd.n1567 vdd.n1566 0.152939
R19921 vdd.n1568 vdd.n1567 0.152939
R19922 vdd.n1569 vdd.n1568 0.152939
R19923 vdd.n1573 vdd.n1569 0.152939
R19924 vdd.n1574 vdd.n1573 0.152939
R19925 vdd.n1575 vdd.n1574 0.152939
R19926 vdd.n1576 vdd.n1575 0.152939
R19927 vdd.n1580 vdd.n1576 0.152939
R19928 vdd.n1581 vdd.n1580 0.152939
R19929 vdd.n1582 vdd.n1581 0.152939
R19930 vdd.n1651 vdd.n1582 0.152939
R19931 vdd.n1651 vdd.n1650 0.152939
R19932 vdd.n1650 vdd.n1649 0.152939
R19933 vdd.n1649 vdd.n1588 0.152939
R19934 vdd.n1593 vdd.n1588 0.152939
R19935 vdd.n1594 vdd.n1593 0.152939
R19936 vdd.n1595 vdd.n1594 0.152939
R19937 vdd.n1599 vdd.n1595 0.152939
R19938 vdd.n1600 vdd.n1599 0.152939
R19939 vdd.n1601 vdd.n1600 0.152939
R19940 vdd.n1602 vdd.n1601 0.152939
R19941 vdd.n1606 vdd.n1602 0.152939
R19942 vdd.n1607 vdd.n1606 0.152939
R19943 vdd.n1608 vdd.n1607 0.152939
R19944 vdd.n1609 vdd.n1608 0.152939
R19945 vdd.n1610 vdd.n1609 0.152939
R19946 vdd.n1610 vdd.n854 0.152939
R19947 vdd.n1939 vdd.n1514 0.152939
R19948 vdd.n1477 vdd.n1476 0.152939
R19949 vdd.n1478 vdd.n1477 0.152939
R19950 vdd.n1478 vdd.n879 0.152939
R19951 vdd.n1493 vdd.n879 0.152939
R19952 vdd.n1494 vdd.n1493 0.152939
R19953 vdd.n1495 vdd.n1494 0.152939
R19954 vdd.n1495 vdd.n867 0.152939
R19955 vdd.n1512 vdd.n867 0.152939
R19956 vdd.n1513 vdd.n1512 0.152939
R19957 vdd.n1940 vdd.n1513 0.152939
R19958 vdd.n524 vdd.n519 0.152939
R19959 vdd.n525 vdd.n524 0.152939
R19960 vdd.n526 vdd.n525 0.152939
R19961 vdd.n527 vdd.n526 0.152939
R19962 vdd.n528 vdd.n527 0.152939
R19963 vdd.n529 vdd.n528 0.152939
R19964 vdd.n530 vdd.n529 0.152939
R19965 vdd.n531 vdd.n530 0.152939
R19966 vdd.n532 vdd.n531 0.152939
R19967 vdd.n533 vdd.n532 0.152939
R19968 vdd.n534 vdd.n533 0.152939
R19969 vdd.n535 vdd.n534 0.152939
R19970 vdd.n2803 vdd.n535 0.152939
R19971 vdd.n2803 vdd.n2802 0.152939
R19972 vdd.n2802 vdd.n2801 0.152939
R19973 vdd.n2801 vdd.n537 0.152939
R19974 vdd.n538 vdd.n537 0.152939
R19975 vdd.n539 vdd.n538 0.152939
R19976 vdd.n540 vdd.n539 0.152939
R19977 vdd.n541 vdd.n540 0.152939
R19978 vdd.n542 vdd.n541 0.152939
R19979 vdd.n543 vdd.n542 0.152939
R19980 vdd.n544 vdd.n543 0.152939
R19981 vdd.n545 vdd.n544 0.152939
R19982 vdd.n546 vdd.n545 0.152939
R19983 vdd.n547 vdd.n546 0.152939
R19984 vdd.n548 vdd.n547 0.152939
R19985 vdd.n549 vdd.n548 0.152939
R19986 vdd.n550 vdd.n549 0.152939
R19987 vdd.n551 vdd.n550 0.152939
R19988 vdd.n552 vdd.n551 0.152939
R19989 vdd.n553 vdd.n552 0.152939
R19990 vdd.n554 vdd.n553 0.152939
R19991 vdd.n555 vdd.n554 0.152939
R19992 vdd.n2757 vdd.n555 0.152939
R19993 vdd.n2757 vdd.n2756 0.152939
R19994 vdd.n2756 vdd.n2755 0.152939
R19995 vdd.n2755 vdd.n559 0.152939
R19996 vdd.n560 vdd.n559 0.152939
R19997 vdd.n561 vdd.n560 0.152939
R19998 vdd.n562 vdd.n561 0.152939
R19999 vdd.n563 vdd.n562 0.152939
R20000 vdd.n564 vdd.n563 0.152939
R20001 vdd.n565 vdd.n564 0.152939
R20002 vdd.n566 vdd.n565 0.152939
R20003 vdd.n567 vdd.n566 0.152939
R20004 vdd.n568 vdd.n567 0.152939
R20005 vdd.n569 vdd.n568 0.152939
R20006 vdd.n570 vdd.n569 0.152939
R20007 vdd.n571 vdd.n570 0.152939
R20008 vdd.n572 vdd.n571 0.152939
R20009 vdd.n2844 vdd.n481 0.152939
R20010 vdd.n2846 vdd.n2845 0.152939
R20011 vdd.n2846 vdd.n470 0.152939
R20012 vdd.n2861 vdd.n470 0.152939
R20013 vdd.n2862 vdd.n2861 0.152939
R20014 vdd.n2863 vdd.n2862 0.152939
R20015 vdd.n2863 vdd.n459 0.152939
R20016 vdd.n2877 vdd.n459 0.152939
R20017 vdd.n2878 vdd.n2877 0.152939
R20018 vdd.n2879 vdd.n2878 0.152939
R20019 vdd.n2879 vdd.n298 0.152939
R20020 vdd.n3046 vdd.n299 0.152939
R20021 vdd.n310 vdd.n299 0.152939
R20022 vdd.n311 vdd.n310 0.152939
R20023 vdd.n312 vdd.n311 0.152939
R20024 vdd.n320 vdd.n312 0.152939
R20025 vdd.n321 vdd.n320 0.152939
R20026 vdd.n322 vdd.n321 0.152939
R20027 vdd.n323 vdd.n322 0.152939
R20028 vdd.n331 vdd.n323 0.152939
R20029 vdd.n3022 vdd.n331 0.152939
R20030 vdd.n3021 vdd.n332 0.152939
R20031 vdd.n335 vdd.n332 0.152939
R20032 vdd.n339 vdd.n335 0.152939
R20033 vdd.n340 vdd.n339 0.152939
R20034 vdd.n341 vdd.n340 0.152939
R20035 vdd.n342 vdd.n341 0.152939
R20036 vdd.n343 vdd.n342 0.152939
R20037 vdd.n347 vdd.n343 0.152939
R20038 vdd.n348 vdd.n347 0.152939
R20039 vdd.n349 vdd.n348 0.152939
R20040 vdd.n350 vdd.n349 0.152939
R20041 vdd.n354 vdd.n350 0.152939
R20042 vdd.n355 vdd.n354 0.152939
R20043 vdd.n356 vdd.n355 0.152939
R20044 vdd.n357 vdd.n356 0.152939
R20045 vdd.n361 vdd.n357 0.152939
R20046 vdd.n362 vdd.n361 0.152939
R20047 vdd.n363 vdd.n362 0.152939
R20048 vdd.n2987 vdd.n363 0.152939
R20049 vdd.n2987 vdd.n2986 0.152939
R20050 vdd.n2986 vdd.n2985 0.152939
R20051 vdd.n2985 vdd.n369 0.152939
R20052 vdd.n374 vdd.n369 0.152939
R20053 vdd.n375 vdd.n374 0.152939
R20054 vdd.n376 vdd.n375 0.152939
R20055 vdd.n380 vdd.n376 0.152939
R20056 vdd.n381 vdd.n380 0.152939
R20057 vdd.n382 vdd.n381 0.152939
R20058 vdd.n383 vdd.n382 0.152939
R20059 vdd.n387 vdd.n383 0.152939
R20060 vdd.n388 vdd.n387 0.152939
R20061 vdd.n389 vdd.n388 0.152939
R20062 vdd.n390 vdd.n389 0.152939
R20063 vdd.n394 vdd.n390 0.152939
R20064 vdd.n395 vdd.n394 0.152939
R20065 vdd.n396 vdd.n395 0.152939
R20066 vdd.n397 vdd.n396 0.152939
R20067 vdd.n401 vdd.n397 0.152939
R20068 vdd.n402 vdd.n401 0.152939
R20069 vdd.n403 vdd.n402 0.152939
R20070 vdd.n2948 vdd.n403 0.152939
R20071 vdd.n2948 vdd.n2947 0.152939
R20072 vdd.n2947 vdd.n2946 0.152939
R20073 vdd.n2946 vdd.n409 0.152939
R20074 vdd.n414 vdd.n409 0.152939
R20075 vdd.n415 vdd.n414 0.152939
R20076 vdd.n416 vdd.n415 0.152939
R20077 vdd.n420 vdd.n416 0.152939
R20078 vdd.n421 vdd.n420 0.152939
R20079 vdd.n422 vdd.n421 0.152939
R20080 vdd.n423 vdd.n422 0.152939
R20081 vdd.n427 vdd.n423 0.152939
R20082 vdd.n428 vdd.n427 0.152939
R20083 vdd.n429 vdd.n428 0.152939
R20084 vdd.n430 vdd.n429 0.152939
R20085 vdd.n434 vdd.n430 0.152939
R20086 vdd.n435 vdd.n434 0.152939
R20087 vdd.n436 vdd.n435 0.152939
R20088 vdd.n437 vdd.n436 0.152939
R20089 vdd.n441 vdd.n437 0.152939
R20090 vdd.n442 vdd.n441 0.152939
R20091 vdd.n443 vdd.n442 0.152939
R20092 vdd.n2904 vdd.n443 0.152939
R20093 vdd.n2852 vdd.n476 0.152939
R20094 vdd.n2853 vdd.n2852 0.152939
R20095 vdd.n2854 vdd.n2853 0.152939
R20096 vdd.n2854 vdd.n464 0.152939
R20097 vdd.n2869 vdd.n464 0.152939
R20098 vdd.n2870 vdd.n2869 0.152939
R20099 vdd.n2871 vdd.n2870 0.152939
R20100 vdd.n2871 vdd.n452 0.152939
R20101 vdd.n2885 vdd.n452 0.152939
R20102 vdd.n2886 vdd.n2885 0.152939
R20103 vdd.n2887 vdd.n2886 0.152939
R20104 vdd.n2887 vdd.n450 0.152939
R20105 vdd.n2891 vdd.n450 0.152939
R20106 vdd.n2892 vdd.n2891 0.152939
R20107 vdd.n2893 vdd.n2892 0.152939
R20108 vdd.n2893 vdd.n447 0.152939
R20109 vdd.n2897 vdd.n447 0.152939
R20110 vdd.n2898 vdd.n2897 0.152939
R20111 vdd.n2899 vdd.n2898 0.152939
R20112 vdd.n2899 vdd.n444 0.152939
R20113 vdd.n2903 vdd.n444 0.152939
R20114 vdd.n2709 vdd.n2708 0.152939
R20115 vdd.n1951 vdd.n857 0.152939
R20116 vdd.n1433 vdd.n1189 0.152939
R20117 vdd.n1434 vdd.n1433 0.152939
R20118 vdd.n1435 vdd.n1434 0.152939
R20119 vdd.n1435 vdd.n1177 0.152939
R20120 vdd.n1450 vdd.n1177 0.152939
R20121 vdd.n1451 vdd.n1450 0.152939
R20122 vdd.n1452 vdd.n1451 0.152939
R20123 vdd.n1452 vdd.n1167 0.152939
R20124 vdd.n1468 vdd.n1167 0.152939
R20125 vdd.n1469 vdd.n1468 0.152939
R20126 vdd.n1470 vdd.n1469 0.152939
R20127 vdd.n1470 vdd.n884 0.152939
R20128 vdd.n1484 vdd.n884 0.152939
R20129 vdd.n1485 vdd.n1484 0.152939
R20130 vdd.n1486 vdd.n1485 0.152939
R20131 vdd.n1486 vdd.n874 0.152939
R20132 vdd.n1501 vdd.n874 0.152939
R20133 vdd.n1502 vdd.n1501 0.152939
R20134 vdd.n1505 vdd.n1502 0.152939
R20135 vdd.n1505 vdd.n1504 0.152939
R20136 vdd.n1504 vdd.n1503 0.152939
R20137 vdd.n1425 vdd.n1194 0.152939
R20138 vdd.n1418 vdd.n1194 0.152939
R20139 vdd.n1418 vdd.n1417 0.152939
R20140 vdd.n1417 vdd.n1416 0.152939
R20141 vdd.n1416 vdd.n1231 0.152939
R20142 vdd.n1412 vdd.n1231 0.152939
R20143 vdd.n1412 vdd.n1411 0.152939
R20144 vdd.n1411 vdd.n1410 0.152939
R20145 vdd.n1410 vdd.n1237 0.152939
R20146 vdd.n1406 vdd.n1237 0.152939
R20147 vdd.n1406 vdd.n1405 0.152939
R20148 vdd.n1405 vdd.n1404 0.152939
R20149 vdd.n1404 vdd.n1243 0.152939
R20150 vdd.n1400 vdd.n1243 0.152939
R20151 vdd.n1400 vdd.n1399 0.152939
R20152 vdd.n1399 vdd.n1398 0.152939
R20153 vdd.n1398 vdd.n1249 0.152939
R20154 vdd.n1394 vdd.n1249 0.152939
R20155 vdd.n1394 vdd.n1393 0.152939
R20156 vdd.n1393 vdd.n1392 0.152939
R20157 vdd.n1392 vdd.n1257 0.152939
R20158 vdd.n1388 vdd.n1257 0.152939
R20159 vdd.n1388 vdd.n1387 0.152939
R20160 vdd.n1387 vdd.n1386 0.152939
R20161 vdd.n1386 vdd.n1263 0.152939
R20162 vdd.n1382 vdd.n1263 0.152939
R20163 vdd.n1382 vdd.n1381 0.152939
R20164 vdd.n1381 vdd.n1380 0.152939
R20165 vdd.n1380 vdd.n1269 0.152939
R20166 vdd.n1376 vdd.n1269 0.152939
R20167 vdd.n1376 vdd.n1375 0.152939
R20168 vdd.n1375 vdd.n1374 0.152939
R20169 vdd.n1374 vdd.n1275 0.152939
R20170 vdd.n1370 vdd.n1275 0.152939
R20171 vdd.n1370 vdd.n1369 0.152939
R20172 vdd.n1369 vdd.n1368 0.152939
R20173 vdd.n1368 vdd.n1281 0.152939
R20174 vdd.n1364 vdd.n1281 0.152939
R20175 vdd.n1364 vdd.n1363 0.152939
R20176 vdd.n1363 vdd.n1362 0.152939
R20177 vdd.n1362 vdd.n1287 0.152939
R20178 vdd.n1355 vdd.n1287 0.152939
R20179 vdd.n1355 vdd.n1354 0.152939
R20180 vdd.n1354 vdd.n1353 0.152939
R20181 vdd.n1353 vdd.n1292 0.152939
R20182 vdd.n1349 vdd.n1292 0.152939
R20183 vdd.n1349 vdd.n1348 0.152939
R20184 vdd.n1348 vdd.n1347 0.152939
R20185 vdd.n1347 vdd.n1298 0.152939
R20186 vdd.n1343 vdd.n1298 0.152939
R20187 vdd.n1343 vdd.n1342 0.152939
R20188 vdd.n1342 vdd.n1341 0.152939
R20189 vdd.n1341 vdd.n1304 0.152939
R20190 vdd.n1337 vdd.n1304 0.152939
R20191 vdd.n1337 vdd.n1336 0.152939
R20192 vdd.n1336 vdd.n1335 0.152939
R20193 vdd.n1335 vdd.n1310 0.152939
R20194 vdd.n1331 vdd.n1310 0.152939
R20195 vdd.n1331 vdd.n1330 0.152939
R20196 vdd.n1330 vdd.n1329 0.152939
R20197 vdd.n1329 vdd.n1316 0.152939
R20198 vdd.n1325 vdd.n1316 0.152939
R20199 vdd.n1325 vdd.n1324 0.152939
R20200 vdd.n1427 vdd.n1426 0.152939
R20201 vdd.n1427 vdd.n1183 0.152939
R20202 vdd.n1442 vdd.n1183 0.152939
R20203 vdd.n1443 vdd.n1442 0.152939
R20204 vdd.n1444 vdd.n1443 0.152939
R20205 vdd.n1444 vdd.n1172 0.152939
R20206 vdd.n1459 vdd.n1172 0.152939
R20207 vdd.n1460 vdd.n1459 0.152939
R20208 vdd.n1462 vdd.n1460 0.152939
R20209 vdd.n1462 vdd.n1461 0.152939
R20210 vdd.n1929 vdd.n1514 0.110256
R20211 vdd.n2836 vdd.n481 0.110256
R20212 vdd.n2708 vdd.n2707 0.110256
R20213 vdd.n1952 vdd.n1951 0.110256
R20214 vdd.n1476 vdd.n1161 0.0695946
R20215 vdd.n3047 vdd.n298 0.0695946
R20216 vdd.n3047 vdd.n3046 0.0695946
R20217 vdd.n1461 vdd.n1161 0.0695946
R20218 vdd.n1929 vdd.n1715 0.0431829
R20219 vdd.n1952 vdd.n854 0.0431829
R20220 vdd.n2836 vdd.n519 0.0431829
R20221 vdd.n2707 vdd.n572 0.0431829
R20222 vdd vdd.n28 0.00833333
R20223 a_n1986_13878.n83 a_n1986_13878.t64 512.366
R20224 a_n1986_13878.n82 a_n1986_13878.t55 512.366
R20225 a_n1986_13878.n81 a_n1986_13878.t49 512.366
R20226 a_n1986_13878.n85 a_n1986_13878.t72 512.366
R20227 a_n1986_13878.n84 a_n1986_13878.t61 512.366
R20228 a_n1986_13878.n80 a_n1986_13878.t60 512.366
R20229 a_n1986_13878.n87 a_n1986_13878.t68 512.366
R20230 a_n1986_13878.n86 a_n1986_13878.t53 512.366
R20231 a_n1986_13878.n79 a_n1986_13878.t54 512.366
R20232 a_n1986_13878.n89 a_n1986_13878.t57 512.366
R20233 a_n1986_13878.n88 a_n1986_13878.t66 512.366
R20234 a_n1986_13878.n78 a_n1986_13878.t48 512.366
R20235 a_n1986_13878.n21 a_n1986_13878.t75 539.01
R20236 a_n1986_13878.n70 a_n1986_13878.t58 512.366
R20237 a_n1986_13878.n69 a_n1986_13878.t62 512.366
R20238 a_n1986_13878.n67 a_n1986_13878.t52 512.366
R20239 a_n1986_13878.n68 a_n1986_13878.t67 512.366
R20240 a_n1986_13878.n17 a_n1986_13878.t23 539.01
R20241 a_n1986_13878.n73 a_n1986_13878.t21 512.366
R20242 a_n1986_13878.n72 a_n1986_13878.t25 512.366
R20243 a_n1986_13878.n54 a_n1986_13878.t19 512.366
R20244 a_n1986_13878.n71 a_n1986_13878.t17 512.366
R20245 a_n1986_13878.n11 a_n1986_13878.t13 539.01
R20246 a_n1986_13878.n94 a_n1986_13878.t15 512.366
R20247 a_n1986_13878.n95 a_n1986_13878.t29 512.366
R20248 a_n1986_13878.n52 a_n1986_13878.t27 512.366
R20249 a_n1986_13878.n96 a_n1986_13878.t33 512.366
R20250 a_n1986_13878.n15 a_n1986_13878.t70 539.01
R20251 a_n1986_13878.n91 a_n1986_13878.t71 512.366
R20252 a_n1986_13878.n92 a_n1986_13878.t50 512.366
R20253 a_n1986_13878.n53 a_n1986_13878.t56 512.366
R20254 a_n1986_13878.n93 a_n1986_13878.t65 512.366
R20255 a_n1986_13878.n0 a_n1986_13878.n50 70.1674
R20256 a_n1986_13878.n2 a_n1986_13878.n48 70.1674
R20257 a_n1986_13878.n4 a_n1986_13878.n46 70.1674
R20258 a_n1986_13878.n6 a_n1986_13878.n44 70.1674
R20259 a_n1986_13878.n33 a_n1986_13878.n19 70.3058
R20260 a_n1986_13878.n51 a_n1986_13878.n29 70.3058
R20261 a_n1986_13878.n20 a_n1986_13878.n31 70.1674
R20262 a_n1986_13878.n31 a_n1986_13878.n67 20.9683
R20263 a_n1986_13878.n30 a_n1986_13878.n20 75.0448
R20264 a_n1986_13878.n69 a_n1986_13878.n30 11.2134
R20265 a_n1986_13878.n18 a_n1986_13878.n21 44.8194
R20266 a_n1986_13878.n29 a_n1986_13878.n36 70.1674
R20267 a_n1986_13878.n36 a_n1986_13878.n54 20.9683
R20268 a_n1986_13878.n35 a_n1986_13878.n34 75.0448
R20269 a_n1986_13878.n72 a_n1986_13878.n35 11.2134
R20270 a_n1986_13878.n16 a_n1986_13878.n17 44.8194
R20271 a_n1986_13878.n8 a_n1986_13878.n42 70.3058
R20272 a_n1986_13878.n12 a_n1986_13878.n39 70.3058
R20273 a_n1986_13878.n38 a_n1986_13878.n13 70.1674
R20274 a_n1986_13878.n38 a_n1986_13878.n53 20.9683
R20275 a_n1986_13878.n13 a_n1986_13878.n37 75.0448
R20276 a_n1986_13878.n92 a_n1986_13878.n37 11.2134
R20277 a_n1986_13878.n14 a_n1986_13878.n15 44.8194
R20278 a_n1986_13878.n41 a_n1986_13878.n9 70.1674
R20279 a_n1986_13878.n41 a_n1986_13878.n52 20.9683
R20280 a_n1986_13878.n9 a_n1986_13878.n40 75.0448
R20281 a_n1986_13878.n95 a_n1986_13878.n40 11.2134
R20282 a_n1986_13878.n10 a_n1986_13878.n11 44.8194
R20283 a_n1986_13878.n44 a_n1986_13878.n78 20.9683
R20284 a_n1986_13878.n43 a_n1986_13878.n7 75.0448
R20285 a_n1986_13878.n88 a_n1986_13878.n43 11.2134
R20286 a_n1986_13878.n7 a_n1986_13878.n89 161.3
R20287 a_n1986_13878.n46 a_n1986_13878.n79 20.9683
R20288 a_n1986_13878.n45 a_n1986_13878.n5 75.0448
R20289 a_n1986_13878.n86 a_n1986_13878.n45 11.2134
R20290 a_n1986_13878.n5 a_n1986_13878.n87 161.3
R20291 a_n1986_13878.n48 a_n1986_13878.n80 20.9683
R20292 a_n1986_13878.n47 a_n1986_13878.n3 75.0448
R20293 a_n1986_13878.n84 a_n1986_13878.n47 11.2134
R20294 a_n1986_13878.n3 a_n1986_13878.n85 161.3
R20295 a_n1986_13878.n50 a_n1986_13878.n81 20.9683
R20296 a_n1986_13878.n49 a_n1986_13878.n1 75.0448
R20297 a_n1986_13878.n82 a_n1986_13878.n49 11.2134
R20298 a_n1986_13878.n1 a_n1986_13878.n83 161.3
R20299 a_n1986_13878.n27 a_n1986_13878.n64 81.2902
R20300 a_n1986_13878.n28 a_n1986_13878.n58 81.2902
R20301 a_n1986_13878.n22 a_n1986_13878.n55 81.2902
R20302 a_n1986_13878.n27 a_n1986_13878.n65 80.9324
R20303 a_n1986_13878.n24 a_n1986_13878.n66 80.9324
R20304 a_n1986_13878.n24 a_n1986_13878.n63 80.9324
R20305 a_n1986_13878.n24 a_n1986_13878.n62 80.9324
R20306 a_n1986_13878.n23 a_n1986_13878.n61 80.9324
R20307 a_n1986_13878.n28 a_n1986_13878.n59 80.9324
R20308 a_n1986_13878.n22 a_n1986_13878.n60 80.9324
R20309 a_n1986_13878.n22 a_n1986_13878.n57 80.9324
R20310 a_n1986_13878.n22 a_n1986_13878.n56 80.9324
R20311 a_n1986_13878.n25 a_n1986_13878.t32 74.6477
R20312 a_n1986_13878.t14 a_n1986_13878.n100 74.6477
R20313 a_n1986_13878.n76 a_n1986_13878.t24 74.2899
R20314 a_n1986_13878.n26 a_n1986_13878.t36 74.2897
R20315 a_n1986_13878.n26 a_n1986_13878.n98 70.6783
R20316 a_n1986_13878.n100 a_n1986_13878.n99 70.6783
R20317 a_n1986_13878.n25 a_n1986_13878.n74 70.6783
R20318 a_n1986_13878.n25 a_n1986_13878.n75 70.6783
R20319 a_n1986_13878.n83 a_n1986_13878.n82 48.2005
R20320 a_n1986_13878.t69 a_n1986_13878.n50 533.335
R20321 a_n1986_13878.n85 a_n1986_13878.n84 48.2005
R20322 a_n1986_13878.t74 a_n1986_13878.n48 533.335
R20323 a_n1986_13878.n87 a_n1986_13878.n86 48.2005
R20324 a_n1986_13878.t63 a_n1986_13878.n46 533.335
R20325 a_n1986_13878.n89 a_n1986_13878.n88 48.2005
R20326 a_n1986_13878.t59 a_n1986_13878.n44 533.335
R20327 a_n1986_13878.n70 a_n1986_13878.n69 48.2005
R20328 a_n1986_13878.n68 a_n1986_13878.n31 20.9683
R20329 a_n1986_13878.n73 a_n1986_13878.n72 48.2005
R20330 a_n1986_13878.n71 a_n1986_13878.n36 20.9683
R20331 a_n1986_13878.n95 a_n1986_13878.n94 48.2005
R20332 a_n1986_13878.n96 a_n1986_13878.n41 20.9683
R20333 a_n1986_13878.n92 a_n1986_13878.n91 48.2005
R20334 a_n1986_13878.n93 a_n1986_13878.n38 20.9683
R20335 a_n1986_13878.n33 a_n1986_13878.t73 533.058
R20336 a_n1986_13878.n51 a_n1986_13878.t31 533.058
R20337 a_n1986_13878.t35 a_n1986_13878.n42 533.058
R20338 a_n1986_13878.t51 a_n1986_13878.n39 533.058
R20339 a_n1986_13878.n23 a_n1986_13878.n22 31.7747
R20340 a_n1986_13878.n49 a_n1986_13878.n81 35.3134
R20341 a_n1986_13878.n47 a_n1986_13878.n80 35.3134
R20342 a_n1986_13878.n45 a_n1986_13878.n79 35.3134
R20343 a_n1986_13878.n43 a_n1986_13878.n78 35.3134
R20344 a_n1986_13878.n30 a_n1986_13878.n67 35.3134
R20345 a_n1986_13878.n35 a_n1986_13878.n54 35.3134
R20346 a_n1986_13878.n52 a_n1986_13878.n40 35.3134
R20347 a_n1986_13878.n53 a_n1986_13878.n37 35.3134
R20348 a_n1986_13878.n29 a_n1986_13878.n24 23.891
R20349 a_n1986_13878.n14 a_n1986_13878.n90 12.046
R20350 a_n1986_13878.n19 a_n1986_13878.n32 11.8414
R20351 a_n1986_13878.n77 a_n1986_13878.n16 10.5365
R20352 a_n1986_13878.n26 a_n1986_13878.n97 9.50122
R20353 a_n1986_13878.n90 a_n1986_13878.n7 7.47588
R20354 a_n1986_13878.n0 a_n1986_13878.n32 7.47588
R20355 a_n1986_13878.n97 a_n1986_13878.n8 6.70126
R20356 a_n1986_13878.n77 a_n1986_13878.n76 5.65783
R20357 a_n1986_13878.n97 a_n1986_13878.n32 5.3452
R20358 a_n1986_13878.n29 a_n1986_13878.n18 3.95126
R20359 a_n1986_13878.n10 a_n1986_13878.n12 3.95126
R20360 a_n1986_13878.n98 a_n1986_13878.t28 3.61217
R20361 a_n1986_13878.n98 a_n1986_13878.t34 3.61217
R20362 a_n1986_13878.n99 a_n1986_13878.t16 3.61217
R20363 a_n1986_13878.n99 a_n1986_13878.t30 3.61217
R20364 a_n1986_13878.n74 a_n1986_13878.t20 3.61217
R20365 a_n1986_13878.n74 a_n1986_13878.t18 3.61217
R20366 a_n1986_13878.n75 a_n1986_13878.t22 3.61217
R20367 a_n1986_13878.n75 a_n1986_13878.t26 3.61217
R20368 a_n1986_13878.n64 a_n1986_13878.t47 2.82907
R20369 a_n1986_13878.n64 a_n1986_13878.t3 2.82907
R20370 a_n1986_13878.n65 a_n1986_13878.t44 2.82907
R20371 a_n1986_13878.n65 a_n1986_13878.t5 2.82907
R20372 a_n1986_13878.n66 a_n1986_13878.t40 2.82907
R20373 a_n1986_13878.n66 a_n1986_13878.t1 2.82907
R20374 a_n1986_13878.n63 a_n1986_13878.t11 2.82907
R20375 a_n1986_13878.n63 a_n1986_13878.t10 2.82907
R20376 a_n1986_13878.n62 a_n1986_13878.t45 2.82907
R20377 a_n1986_13878.n62 a_n1986_13878.t9 2.82907
R20378 a_n1986_13878.n61 a_n1986_13878.t12 2.82907
R20379 a_n1986_13878.n61 a_n1986_13878.t7 2.82907
R20380 a_n1986_13878.n58 a_n1986_13878.t43 2.82907
R20381 a_n1986_13878.n58 a_n1986_13878.t41 2.82907
R20382 a_n1986_13878.n59 a_n1986_13878.t38 2.82907
R20383 a_n1986_13878.n59 a_n1986_13878.t37 2.82907
R20384 a_n1986_13878.n60 a_n1986_13878.t8 2.82907
R20385 a_n1986_13878.n60 a_n1986_13878.t0 2.82907
R20386 a_n1986_13878.n57 a_n1986_13878.t42 2.82907
R20387 a_n1986_13878.n57 a_n1986_13878.t4 2.82907
R20388 a_n1986_13878.n56 a_n1986_13878.t2 2.82907
R20389 a_n1986_13878.n56 a_n1986_13878.t46 2.82907
R20390 a_n1986_13878.n55 a_n1986_13878.t39 2.82907
R20391 a_n1986_13878.n55 a_n1986_13878.t6 2.82907
R20392 a_n1986_13878.n90 a_n1986_13878.n77 1.30542
R20393 a_n1986_13878.n4 a_n1986_13878.n3 1.04595
R20394 a_n1986_13878.n21 a_n1986_13878.n70 13.657
R20395 a_n1986_13878.n68 a_n1986_13878.n33 21.4216
R20396 a_n1986_13878.n17 a_n1986_13878.n73 13.657
R20397 a_n1986_13878.n71 a_n1986_13878.n51 21.4216
R20398 a_n1986_13878.n94 a_n1986_13878.n11 13.657
R20399 a_n1986_13878.n42 a_n1986_13878.n96 21.4216
R20400 a_n1986_13878.n91 a_n1986_13878.n15 13.657
R20401 a_n1986_13878.n39 a_n1986_13878.n93 21.4216
R20402 a_n1986_13878.n22 a_n1986_13878.n28 1.07378
R20403 a_n1986_13878.n20 a_n1986_13878.n18 0.758076
R20404 a_n1986_13878.n20 a_n1986_13878.n19 0.758076
R20405 a_n1986_13878.n34 a_n1986_13878.n16 0.758076
R20406 a_n1986_13878.n14 a_n1986_13878.n13 0.758076
R20407 a_n1986_13878.n13 a_n1986_13878.n12 0.758076
R20408 a_n1986_13878.n10 a_n1986_13878.n9 0.758076
R20409 a_n1986_13878.n9 a_n1986_13878.n8 0.758076
R20410 a_n1986_13878.n7 a_n1986_13878.n6 0.758076
R20411 a_n1986_13878.n5 a_n1986_13878.n4 0.758076
R20412 a_n1986_13878.n3 a_n1986_13878.n2 0.758076
R20413 a_n1986_13878.n1 a_n1986_13878.n0 0.758076
R20414 a_n1986_13878.n34 a_n1986_13878.n29 0.720197
R20415 a_n1986_13878.n24 a_n1986_13878.n27 0.716017
R20416 a_n1986_13878.n100 a_n1986_13878.n26 0.716017
R20417 a_n1986_13878.n76 a_n1986_13878.n25 0.716017
R20418 a_n1986_13878.n24 a_n1986_13878.n23 0.716017
R20419 a_n1986_13878.n6 a_n1986_13878.n5 0.67853
R20420 a_n1986_13878.n2 a_n1986_13878.n1 0.67853
R20421 a_n1986_8322.n6 a_n1986_8322.t6 74.6477
R20422 a_n1986_8322.n1 a_n1986_8322.t13 74.6477
R20423 a_n1986_8322.t22 a_n1986_8322.n18 74.6476
R20424 a_n1986_8322.n14 a_n1986_8322.t15 74.2899
R20425 a_n1986_8322.n7 a_n1986_8322.t4 74.2899
R20426 a_n1986_8322.n8 a_n1986_8322.t7 74.2899
R20427 a_n1986_8322.n11 a_n1986_8322.t8 74.2899
R20428 a_n1986_8322.n4 a_n1986_8322.t12 74.2899
R20429 a_n1986_8322.n18 a_n1986_8322.n17 70.6783
R20430 a_n1986_8322.n16 a_n1986_8322.n15 70.6783
R20431 a_n1986_8322.n6 a_n1986_8322.n5 70.6783
R20432 a_n1986_8322.n10 a_n1986_8322.n9 70.6783
R20433 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R20434 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R20435 a_n1986_8322.n12 a_n1986_8322.n4 22.7556
R20436 a_n1986_8322.n13 a_n1986_8322.t0 9.94227
R20437 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R20438 a_n1986_8322.n14 a_n1986_8322.n13 5.83671
R20439 a_n1986_8322.n13 a_n1986_8322.n12 5.3452
R20440 a_n1986_8322.n17 a_n1986_8322.t20 3.61217
R20441 a_n1986_8322.n17 a_n1986_8322.t17 3.61217
R20442 a_n1986_8322.n15 a_n1986_8322.t14 3.61217
R20443 a_n1986_8322.n15 a_n1986_8322.t23 3.61217
R20444 a_n1986_8322.n5 a_n1986_8322.t10 3.61217
R20445 a_n1986_8322.n5 a_n1986_8322.t9 3.61217
R20446 a_n1986_8322.n9 a_n1986_8322.t5 3.61217
R20447 a_n1986_8322.n9 a_n1986_8322.t11 3.61217
R20448 a_n1986_8322.n0 a_n1986_8322.t21 3.61217
R20449 a_n1986_8322.n0 a_n1986_8322.t16 3.61217
R20450 a_n1986_8322.n2 a_n1986_8322.t19 3.61217
R20451 a_n1986_8322.n2 a_n1986_8322.t18 3.61217
R20452 a_n1986_8322.n11 a_n1986_8322.n10 0.358259
R20453 a_n1986_8322.n10 a_n1986_8322.n8 0.358259
R20454 a_n1986_8322.n7 a_n1986_8322.n6 0.358259
R20455 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R20456 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R20457 a_n1986_8322.n16 a_n1986_8322.n14 0.358259
R20458 a_n1986_8322.n18 a_n1986_8322.n16 0.358259
R20459 a_n1986_8322.n8 a_n1986_8322.n7 0.101793
R20460 a_n1986_8322.t3 a_n1986_8322.t2 0.0788333
R20461 a_n1986_8322.t1 a_n1986_8322.t3 0.0631667
R20462 a_n1986_8322.t0 a_n1986_8322.t1 0.0471944
R20463 a_n1986_8322.t0 a_n1986_8322.t2 0.0453889
R20464 a_n1808_13878.n5 a_n1808_13878.n3 98.9633
R20465 a_n1808_13878.n2 a_n1808_13878.n0 98.7517
R20466 a_n1808_13878.n2 a_n1808_13878.n1 98.6055
R20467 a_n1808_13878.n5 a_n1808_13878.n4 98.6055
R20468 a_n1808_13878.n17 a_n1808_13878.n16 98.6054
R20469 a_n1808_13878.n7 a_n1808_13878.n6 98.6054
R20470 a_n1808_13878.n9 a_n1808_13878.t13 74.6477
R20471 a_n1808_13878.n14 a_n1808_13878.t14 74.2899
R20472 a_n1808_13878.n11 a_n1808_13878.t15 74.2899
R20473 a_n1808_13878.n10 a_n1808_13878.t12 74.2899
R20474 a_n1808_13878.n13 a_n1808_13878.n12 70.6783
R20475 a_n1808_13878.n9 a_n1808_13878.n8 70.6783
R20476 a_n1808_13878.n16 a_n1808_13878.n15 13.5694
R20477 a_n1808_13878.n15 a_n1808_13878.n7 11.5762
R20478 a_n1808_13878.n15 a_n1808_13878.n14 6.2408
R20479 a_n1808_13878.n1 a_n1808_13878.t6 3.61217
R20480 a_n1808_13878.n1 a_n1808_13878.t1 3.61217
R20481 a_n1808_13878.n0 a_n1808_13878.t0 3.61217
R20482 a_n1808_13878.n0 a_n1808_13878.t2 3.61217
R20483 a_n1808_13878.n6 a_n1808_13878.t7 3.61217
R20484 a_n1808_13878.n6 a_n1808_13878.t8 3.61217
R20485 a_n1808_13878.n4 a_n1808_13878.t10 3.61217
R20486 a_n1808_13878.n4 a_n1808_13878.t3 3.61217
R20487 a_n1808_13878.n3 a_n1808_13878.t5 3.61217
R20488 a_n1808_13878.n3 a_n1808_13878.t9 3.61217
R20489 a_n1808_13878.n12 a_n1808_13878.t18 3.61217
R20490 a_n1808_13878.n12 a_n1808_13878.t19 3.61217
R20491 a_n1808_13878.n8 a_n1808_13878.t16 3.61217
R20492 a_n1808_13878.n8 a_n1808_13878.t17 3.61217
R20493 a_n1808_13878.n17 a_n1808_13878.t4 3.61217
R20494 a_n1808_13878.t11 a_n1808_13878.n17 3.61217
R20495 a_n1808_13878.n7 a_n1808_13878.n5 0.358259
R20496 a_n1808_13878.n10 a_n1808_13878.n9 0.358259
R20497 a_n1808_13878.n13 a_n1808_13878.n11 0.358259
R20498 a_n1808_13878.n14 a_n1808_13878.n13 0.358259
R20499 a_n1808_13878.n16 a_n1808_13878.n2 0.146627
R20500 a_n1808_13878.n11 a_n1808_13878.n10 0.101793
R20501 diffpairibias.n0 diffpairibias.t27 436.822
R20502 diffpairibias.n27 diffpairibias.t24 435.479
R20503 diffpairibias.n26 diffpairibias.t21 435.479
R20504 diffpairibias.n25 diffpairibias.t22 435.479
R20505 diffpairibias.n24 diffpairibias.t26 435.479
R20506 diffpairibias.n23 diffpairibias.t20 435.479
R20507 diffpairibias.n0 diffpairibias.t23 435.479
R20508 diffpairibias.n1 diffpairibias.t28 435.479
R20509 diffpairibias.n2 diffpairibias.t25 435.479
R20510 diffpairibias.n3 diffpairibias.t29 435.479
R20511 diffpairibias.n13 diffpairibias.t14 377.536
R20512 diffpairibias.n13 diffpairibias.t0 376.193
R20513 diffpairibias.n14 diffpairibias.t10 376.193
R20514 diffpairibias.n15 diffpairibias.t12 376.193
R20515 diffpairibias.n16 diffpairibias.t6 376.193
R20516 diffpairibias.n17 diffpairibias.t2 376.193
R20517 diffpairibias.n18 diffpairibias.t16 376.193
R20518 diffpairibias.n19 diffpairibias.t4 376.193
R20519 diffpairibias.n20 diffpairibias.t18 376.193
R20520 diffpairibias.n21 diffpairibias.t8 376.193
R20521 diffpairibias.n4 diffpairibias.t15 113.368
R20522 diffpairibias.n4 diffpairibias.t1 112.698
R20523 diffpairibias.n5 diffpairibias.t11 112.698
R20524 diffpairibias.n6 diffpairibias.t13 112.698
R20525 diffpairibias.n7 diffpairibias.t7 112.698
R20526 diffpairibias.n8 diffpairibias.t3 112.698
R20527 diffpairibias.n9 diffpairibias.t17 112.698
R20528 diffpairibias.n10 diffpairibias.t5 112.698
R20529 diffpairibias.n11 diffpairibias.t19 112.698
R20530 diffpairibias.n12 diffpairibias.t9 112.698
R20531 diffpairibias.n22 diffpairibias.n21 4.77242
R20532 diffpairibias.n22 diffpairibias.n12 4.30807
R20533 diffpairibias.n23 diffpairibias.n22 4.13945
R20534 diffpairibias.n21 diffpairibias.n20 1.34352
R20535 diffpairibias.n20 diffpairibias.n19 1.34352
R20536 diffpairibias.n19 diffpairibias.n18 1.34352
R20537 diffpairibias.n18 diffpairibias.n17 1.34352
R20538 diffpairibias.n17 diffpairibias.n16 1.34352
R20539 diffpairibias.n16 diffpairibias.n15 1.34352
R20540 diffpairibias.n15 diffpairibias.n14 1.34352
R20541 diffpairibias.n14 diffpairibias.n13 1.34352
R20542 diffpairibias.n3 diffpairibias.n2 1.34352
R20543 diffpairibias.n2 diffpairibias.n1 1.34352
R20544 diffpairibias.n1 diffpairibias.n0 1.34352
R20545 diffpairibias.n24 diffpairibias.n23 1.34352
R20546 diffpairibias.n25 diffpairibias.n24 1.34352
R20547 diffpairibias.n26 diffpairibias.n25 1.34352
R20548 diffpairibias.n27 diffpairibias.n26 1.34352
R20549 diffpairibias.n28 diffpairibias.n27 0.862419
R20550 diffpairibias diffpairibias.n28 0.684875
R20551 diffpairibias.n12 diffpairibias.n11 0.672012
R20552 diffpairibias.n11 diffpairibias.n10 0.672012
R20553 diffpairibias.n10 diffpairibias.n9 0.672012
R20554 diffpairibias.n9 diffpairibias.n8 0.672012
R20555 diffpairibias.n8 diffpairibias.n7 0.672012
R20556 diffpairibias.n7 diffpairibias.n6 0.672012
R20557 diffpairibias.n6 diffpairibias.n5 0.672012
R20558 diffpairibias.n5 diffpairibias.n4 0.672012
R20559 diffpairibias.n28 diffpairibias.n3 0.190907
R20560 a_n3827_n3924.n51 a_n3827_n3924.t13 214.994
R20561 a_n3827_n3924.t20 a_n3827_n3924.n58 214.994
R20562 a_n3827_n3924.n51 a_n3827_n3924.t17 214.321
R20563 a_n3827_n3924.n53 a_n3827_n3924.t12 214.321
R20564 a_n3827_n3924.n54 a_n3827_n3924.t15 214.321
R20565 a_n3827_n3924.n55 a_n3827_n3924.t11 214.321
R20566 a_n3827_n3924.n56 a_n3827_n3924.t16 214.321
R20567 a_n3827_n3924.n57 a_n3827_n3924.t19 214.321
R20568 a_n3827_n3924.n0 a_n3827_n3924.t18 214.321
R20569 a_n3827_n3924.n58 a_n3827_n3924.t14 214.321
R20570 a_n3827_n3924.n14 a_n3827_n3924.t45 55.8337
R20571 a_n3827_n3924.n13 a_n3827_n3924.t21 55.8337
R20572 a_n3827_n3924.n2 a_n3827_n3924.t31 55.8337
R20573 a_n3827_n3924.n25 a_n3827_n3924.t5 55.8335
R20574 a_n3827_n3924.n49 a_n3827_n3924.t38 55.8335
R20575 a_n3827_n3924.n38 a_n3827_n3924.t36 55.8335
R20576 a_n3827_n3924.n37 a_n3827_n3924.t41 55.8335
R20577 a_n3827_n3924.n26 a_n3827_n3924.t55 55.8335
R20578 a_n3827_n3924.n24 a_n3827_n3924.n23 53.0052
R20579 a_n3827_n3924.n22 a_n3827_n3924.n21 53.0052
R20580 a_n3827_n3924.n20 a_n3827_n3924.n19 53.0052
R20581 a_n3827_n3924.n18 a_n3827_n3924.n17 53.0052
R20582 a_n3827_n3924.n16 a_n3827_n3924.n15 53.0052
R20583 a_n3827_n3924.n12 a_n3827_n3924.n11 53.0052
R20584 a_n3827_n3924.n10 a_n3827_n3924.n9 53.0052
R20585 a_n3827_n3924.n8 a_n3827_n3924.n7 53.0052
R20586 a_n3827_n3924.n6 a_n3827_n3924.n5 53.0052
R20587 a_n3827_n3924.n4 a_n3827_n3924.n3 53.0052
R20588 a_n3827_n3924.n48 a_n3827_n3924.n47 53.0051
R20589 a_n3827_n3924.n46 a_n3827_n3924.n45 53.0051
R20590 a_n3827_n3924.n44 a_n3827_n3924.n43 53.0051
R20591 a_n3827_n3924.n42 a_n3827_n3924.n41 53.0051
R20592 a_n3827_n3924.n40 a_n3827_n3924.n39 53.0051
R20593 a_n3827_n3924.n36 a_n3827_n3924.n35 53.0051
R20594 a_n3827_n3924.n34 a_n3827_n3924.n33 53.0051
R20595 a_n3827_n3924.n32 a_n3827_n3924.n31 53.0051
R20596 a_n3827_n3924.n30 a_n3827_n3924.n29 53.0051
R20597 a_n3827_n3924.n28 a_n3827_n3924.n27 53.0051
R20598 a_n3827_n3924.n2 a_n3827_n3924.n1 12.1555
R20599 a_n3827_n3924.n50 a_n3827_n3924.n25 12.1555
R20600 a_n3827_n3924.n26 a_n3827_n3924.n1 5.07593
R20601 a_n3827_n3924.n50 a_n3827_n3924.n49 5.07593
R20602 a_n3827_n3924.n47 a_n3827_n3924.t34 2.82907
R20603 a_n3827_n3924.n47 a_n3827_n3924.t50 2.82907
R20604 a_n3827_n3924.n45 a_n3827_n3924.t7 2.82907
R20605 a_n3827_n3924.n45 a_n3827_n3924.t35 2.82907
R20606 a_n3827_n3924.n43 a_n3827_n3924.t22 2.82907
R20607 a_n3827_n3924.n43 a_n3827_n3924.t27 2.82907
R20608 a_n3827_n3924.n41 a_n3827_n3924.t53 2.82907
R20609 a_n3827_n3924.n41 a_n3827_n3924.t49 2.82907
R20610 a_n3827_n3924.n39 a_n3827_n3924.t25 2.82907
R20611 a_n3827_n3924.n39 a_n3827_n3924.t10 2.82907
R20612 a_n3827_n3924.n35 a_n3827_n3924.t47 2.82907
R20613 a_n3827_n3924.n35 a_n3827_n3924.t23 2.82907
R20614 a_n3827_n3924.n33 a_n3827_n3924.t9 2.82907
R20615 a_n3827_n3924.n33 a_n3827_n3924.t56 2.82907
R20616 a_n3827_n3924.n31 a_n3827_n3924.t1 2.82907
R20617 a_n3827_n3924.n31 a_n3827_n3924.t4 2.82907
R20618 a_n3827_n3924.n29 a_n3827_n3924.t33 2.82907
R20619 a_n3827_n3924.n29 a_n3827_n3924.t3 2.82907
R20620 a_n3827_n3924.n27 a_n3827_n3924.t40 2.82907
R20621 a_n3827_n3924.n27 a_n3827_n3924.t2 2.82907
R20622 a_n3827_n3924.n23 a_n3827_n3924.t57 2.82907
R20623 a_n3827_n3924.n23 a_n3827_n3924.t46 2.82907
R20624 a_n3827_n3924.n21 a_n3827_n3924.t48 2.82907
R20625 a_n3827_n3924.n21 a_n3827_n3924.t0 2.82907
R20626 a_n3827_n3924.n19 a_n3827_n3924.t42 2.82907
R20627 a_n3827_n3924.n19 a_n3827_n3924.t39 2.82907
R20628 a_n3827_n3924.n17 a_n3827_n3924.t32 2.82907
R20629 a_n3827_n3924.n17 a_n3827_n3924.t43 2.82907
R20630 a_n3827_n3924.n15 a_n3827_n3924.t44 2.82907
R20631 a_n3827_n3924.n15 a_n3827_n3924.t6 2.82907
R20632 a_n3827_n3924.n11 a_n3827_n3924.t24 2.82907
R20633 a_n3827_n3924.n11 a_n3827_n3924.t54 2.82907
R20634 a_n3827_n3924.n9 a_n3827_n3924.t8 2.82907
R20635 a_n3827_n3924.n9 a_n3827_n3924.t51 2.82907
R20636 a_n3827_n3924.n7 a_n3827_n3924.t29 2.82907
R20637 a_n3827_n3924.n7 a_n3827_n3924.t37 2.82907
R20638 a_n3827_n3924.n5 a_n3827_n3924.t28 2.82907
R20639 a_n3827_n3924.n5 a_n3827_n3924.t30 2.82907
R20640 a_n3827_n3924.n3 a_n3827_n3924.t26 2.82907
R20641 a_n3827_n3924.n3 a_n3827_n3924.t52 2.82907
R20642 a_n3827_n3924.n0 a_n3827_n3924.n1 1.95694
R20643 a_n3827_n3924.n52 a_n3827_n3924.n50 1.95694
R20644 a_n3827_n3924.n58 a_n3827_n3924.n0 0.672012
R20645 a_n3827_n3924.n57 a_n3827_n3924.n56 0.672012
R20646 a_n3827_n3924.n56 a_n3827_n3924.n55 0.672012
R20647 a_n3827_n3924.n55 a_n3827_n3924.n54 0.672012
R20648 a_n3827_n3924.n54 a_n3827_n3924.n53 0.672012
R20649 a_n3827_n3924.n0 a_n3827_n3924.n57 0.672012
R20650 a_n3827_n3924.n53 a_n3827_n3924.n52 0.501227
R20651 a_n3827_n3924.n4 a_n3827_n3924.n2 0.358259
R20652 a_n3827_n3924.n6 a_n3827_n3924.n4 0.358259
R20653 a_n3827_n3924.n8 a_n3827_n3924.n6 0.358259
R20654 a_n3827_n3924.n10 a_n3827_n3924.n8 0.358259
R20655 a_n3827_n3924.n12 a_n3827_n3924.n10 0.358259
R20656 a_n3827_n3924.n13 a_n3827_n3924.n12 0.358259
R20657 a_n3827_n3924.n16 a_n3827_n3924.n14 0.358259
R20658 a_n3827_n3924.n18 a_n3827_n3924.n16 0.358259
R20659 a_n3827_n3924.n20 a_n3827_n3924.n18 0.358259
R20660 a_n3827_n3924.n22 a_n3827_n3924.n20 0.358259
R20661 a_n3827_n3924.n24 a_n3827_n3924.n22 0.358259
R20662 a_n3827_n3924.n25 a_n3827_n3924.n24 0.358259
R20663 a_n3827_n3924.n28 a_n3827_n3924.n26 0.358259
R20664 a_n3827_n3924.n30 a_n3827_n3924.n28 0.358259
R20665 a_n3827_n3924.n32 a_n3827_n3924.n30 0.358259
R20666 a_n3827_n3924.n34 a_n3827_n3924.n32 0.358259
R20667 a_n3827_n3924.n36 a_n3827_n3924.n34 0.358259
R20668 a_n3827_n3924.n37 a_n3827_n3924.n36 0.358259
R20669 a_n3827_n3924.n40 a_n3827_n3924.n38 0.358259
R20670 a_n3827_n3924.n42 a_n3827_n3924.n40 0.358259
R20671 a_n3827_n3924.n44 a_n3827_n3924.n42 0.358259
R20672 a_n3827_n3924.n46 a_n3827_n3924.n44 0.358259
R20673 a_n3827_n3924.n48 a_n3827_n3924.n46 0.358259
R20674 a_n3827_n3924.n49 a_n3827_n3924.n48 0.358259
R20675 a_n3827_n3924.n14 a_n3827_n3924.n13 0.235414
R20676 a_n3827_n3924.n38 a_n3827_n3924.n37 0.235414
R20677 a_n3827_n3924.n52 a_n3827_n3924.n51 0.171285
R20678 minus.n45 minus.t26 442.325
R20679 minus.n9 minus.t12 442.325
R20680 minus.n66 minus.t15 415.966
R20681 minus.n64 minus.t28 415.966
R20682 minus.n63 minus.t21 415.966
R20683 minus.n37 minus.t14 415.966
R20684 minus.n57 minus.t23 415.966
R20685 minus.n56 minus.t11 415.966
R20686 minus.n40 minus.t5 415.966
R20687 minus.n51 minus.t17 415.966
R20688 minus.n49 minus.t10 415.966
R20689 minus.n43 minus.t25 415.966
R20690 minus.n44 minus.t7 415.966
R20691 minus.n8 minus.t18 415.966
R20692 minus.n7 minus.t8 415.966
R20693 minus.n13 minus.t13 415.966
R20694 minus.n5 minus.t24 415.966
R20695 minus.n18 minus.t19 415.966
R20696 minus.n20 minus.t22 415.966
R20697 minus.n3 minus.t6 415.966
R20698 minus.n25 minus.t20 415.966
R20699 minus.n1 minus.t27 415.966
R20700 minus.n30 minus.t16 415.966
R20701 minus.n32 minus.t9 415.966
R20702 minus.n72 minus.t3 243.255
R20703 minus.n71 minus.n69 224.169
R20704 minus.n71 minus.n70 223.454
R20705 minus.n46 minus.n43 161.3
R20706 minus.n48 minus.n47 161.3
R20707 minus.n49 minus.n42 161.3
R20708 minus.n50 minus.n41 161.3
R20709 minus.n52 minus.n51 161.3
R20710 minus.n53 minus.n40 161.3
R20711 minus.n55 minus.n54 161.3
R20712 minus.n56 minus.n39 161.3
R20713 minus.n57 minus.n38 161.3
R20714 minus.n59 minus.n58 161.3
R20715 minus.n60 minus.n37 161.3
R20716 minus.n62 minus.n61 161.3
R20717 minus.n63 minus.n36 161.3
R20718 minus.n64 minus.n35 161.3
R20719 minus.n65 minus.n34 161.3
R20720 minus.n67 minus.n66 161.3
R20721 minus.n33 minus.n32 161.3
R20722 minus.n31 minus.n0 161.3
R20723 minus.n30 minus.n29 161.3
R20724 minus.n28 minus.n1 161.3
R20725 minus.n27 minus.n26 161.3
R20726 minus.n25 minus.n2 161.3
R20727 minus.n24 minus.n23 161.3
R20728 minus.n22 minus.n3 161.3
R20729 minus.n21 minus.n20 161.3
R20730 minus.n19 minus.n4 161.3
R20731 minus.n18 minus.n17 161.3
R20732 minus.n16 minus.n5 161.3
R20733 minus.n15 minus.n14 161.3
R20734 minus.n13 minus.n6 161.3
R20735 minus.n12 minus.n11 161.3
R20736 minus.n10 minus.n7 161.3
R20737 minus.n64 minus.n63 48.2005
R20738 minus.n57 minus.n56 48.2005
R20739 minus.n51 minus.n40 48.2005
R20740 minus.n44 minus.n43 48.2005
R20741 minus.n8 minus.n7 48.2005
R20742 minus.n18 minus.n5 48.2005
R20743 minus.n20 minus.n3 48.2005
R20744 minus.n30 minus.n1 48.2005
R20745 minus.n58 minus.n37 47.4702
R20746 minus.n50 minus.n49 47.4702
R20747 minus.n14 minus.n13 47.4702
R20748 minus.n25 minus.n24 47.4702
R20749 minus.n66 minus.n65 46.0096
R20750 minus.n32 minus.n31 46.0096
R20751 minus.n10 minus.n9 45.0871
R20752 minus.n46 minus.n45 45.0871
R20753 minus.n68 minus.n67 31.2713
R20754 minus.n62 minus.n37 25.5611
R20755 minus.n49 minus.n48 25.5611
R20756 minus.n13 minus.n12 25.5611
R20757 minus.n26 minus.n25 25.5611
R20758 minus.n56 minus.n55 24.1005
R20759 minus.n55 minus.n40 24.1005
R20760 minus.n19 minus.n18 24.1005
R20761 minus.n20 minus.n19 24.1005
R20762 minus.n63 minus.n62 22.6399
R20763 minus.n48 minus.n43 22.6399
R20764 minus.n12 minus.n7 22.6399
R20765 minus.n26 minus.n1 22.6399
R20766 minus.n70 minus.t2 19.8005
R20767 minus.n70 minus.t0 19.8005
R20768 minus.n69 minus.t1 19.8005
R20769 minus.n69 minus.t4 19.8005
R20770 minus.n45 minus.n44 14.1472
R20771 minus.n9 minus.n8 14.1472
R20772 minus.n68 minus.n33 11.9418
R20773 minus minus.n73 11.5306
R20774 minus.n73 minus.n72 4.80222
R20775 minus.n65 minus.n64 2.19141
R20776 minus.n31 minus.n30 2.19141
R20777 minus.n73 minus.n68 0.972091
R20778 minus.n58 minus.n57 0.730803
R20779 minus.n51 minus.n50 0.730803
R20780 minus.n14 minus.n5 0.730803
R20781 minus.n24 minus.n3 0.730803
R20782 minus.n72 minus.n71 0.716017
R20783 minus.n67 minus.n34 0.189894
R20784 minus.n35 minus.n34 0.189894
R20785 minus.n36 minus.n35 0.189894
R20786 minus.n61 minus.n36 0.189894
R20787 minus.n61 minus.n60 0.189894
R20788 minus.n60 minus.n59 0.189894
R20789 minus.n59 minus.n38 0.189894
R20790 minus.n39 minus.n38 0.189894
R20791 minus.n54 minus.n39 0.189894
R20792 minus.n54 minus.n53 0.189894
R20793 minus.n53 minus.n52 0.189894
R20794 minus.n52 minus.n41 0.189894
R20795 minus.n42 minus.n41 0.189894
R20796 minus.n47 minus.n42 0.189894
R20797 minus.n47 minus.n46 0.189894
R20798 minus.n11 minus.n10 0.189894
R20799 minus.n11 minus.n6 0.189894
R20800 minus.n15 minus.n6 0.189894
R20801 minus.n16 minus.n15 0.189894
R20802 minus.n17 minus.n16 0.189894
R20803 minus.n17 minus.n4 0.189894
R20804 minus.n21 minus.n4 0.189894
R20805 minus.n22 minus.n21 0.189894
R20806 minus.n23 minus.n22 0.189894
R20807 minus.n23 minus.n2 0.189894
R20808 minus.n27 minus.n2 0.189894
R20809 minus.n28 minus.n27 0.189894
R20810 minus.n29 minus.n28 0.189894
R20811 minus.n29 minus.n0 0.189894
R20812 minus.n33 minus.n0 0.189894
R20813 plus.n43 plus.t25 442.325
R20814 plus.n11 plus.t12 442.325
R20815 plus.n42 plus.t5 415.966
R20816 plus.n41 plus.t20 415.966
R20817 plus.n47 plus.t26 415.966
R20818 plus.n39 plus.t11 415.966
R20819 plus.n52 plus.t6 415.966
R20820 plus.n54 plus.t10 415.966
R20821 plus.n37 plus.t19 415.966
R20822 plus.n59 plus.t8 415.966
R20823 plus.n35 plus.t16 415.966
R20824 plus.n64 plus.t28 415.966
R20825 plus.n66 plus.t21 415.966
R20826 plus.n32 plus.t23 415.966
R20827 plus.n30 plus.t13 415.966
R20828 plus.n29 plus.t27 415.966
R20829 plus.n3 plus.t22 415.966
R20830 plus.n23 plus.t7 415.966
R20831 plus.n22 plus.t18 415.966
R20832 plus.n6 plus.t14 415.966
R20833 plus.n17 plus.t24 415.966
R20834 plus.n15 plus.t17 415.966
R20835 plus.n9 plus.t9 415.966
R20836 plus.n10 plus.t15 415.966
R20837 plus.n70 plus.t3 243.97
R20838 plus.n70 plus.n69 223.454
R20839 plus.n72 plus.n71 223.454
R20840 plus.n67 plus.n66 161.3
R20841 plus.n65 plus.n34 161.3
R20842 plus.n64 plus.n63 161.3
R20843 plus.n62 plus.n35 161.3
R20844 plus.n61 plus.n60 161.3
R20845 plus.n59 plus.n36 161.3
R20846 plus.n58 plus.n57 161.3
R20847 plus.n56 plus.n37 161.3
R20848 plus.n55 plus.n54 161.3
R20849 plus.n53 plus.n38 161.3
R20850 plus.n52 plus.n51 161.3
R20851 plus.n50 plus.n39 161.3
R20852 plus.n49 plus.n48 161.3
R20853 plus.n47 plus.n40 161.3
R20854 plus.n46 plus.n45 161.3
R20855 plus.n44 plus.n41 161.3
R20856 plus.n12 plus.n9 161.3
R20857 plus.n14 plus.n13 161.3
R20858 plus.n15 plus.n8 161.3
R20859 plus.n16 plus.n7 161.3
R20860 plus.n18 plus.n17 161.3
R20861 plus.n19 plus.n6 161.3
R20862 plus.n21 plus.n20 161.3
R20863 plus.n22 plus.n5 161.3
R20864 plus.n23 plus.n4 161.3
R20865 plus.n25 plus.n24 161.3
R20866 plus.n26 plus.n3 161.3
R20867 plus.n28 plus.n27 161.3
R20868 plus.n29 plus.n2 161.3
R20869 plus.n30 plus.n1 161.3
R20870 plus.n31 plus.n0 161.3
R20871 plus.n33 plus.n32 161.3
R20872 plus.n42 plus.n41 48.2005
R20873 plus.n52 plus.n39 48.2005
R20874 plus.n54 plus.n37 48.2005
R20875 plus.n64 plus.n35 48.2005
R20876 plus.n30 plus.n29 48.2005
R20877 plus.n23 plus.n22 48.2005
R20878 plus.n17 plus.n6 48.2005
R20879 plus.n10 plus.n9 48.2005
R20880 plus.n48 plus.n47 47.4702
R20881 plus.n59 plus.n58 47.4702
R20882 plus.n24 plus.n3 47.4702
R20883 plus.n16 plus.n15 47.4702
R20884 plus.n66 plus.n65 46.0096
R20885 plus.n32 plus.n31 46.0096
R20886 plus.n44 plus.n43 45.0871
R20887 plus.n12 plus.n11 45.0871
R20888 plus.n68 plus.n67 31.0554
R20889 plus.n47 plus.n46 25.5611
R20890 plus.n60 plus.n59 25.5611
R20891 plus.n28 plus.n3 25.5611
R20892 plus.n15 plus.n14 25.5611
R20893 plus.n53 plus.n52 24.1005
R20894 plus.n54 plus.n53 24.1005
R20895 plus.n22 plus.n21 24.1005
R20896 plus.n21 plus.n6 24.1005
R20897 plus.n46 plus.n41 22.6399
R20898 plus.n60 plus.n35 22.6399
R20899 plus.n29 plus.n28 22.6399
R20900 plus.n14 plus.n9 22.6399
R20901 plus.n69 plus.t4 19.8005
R20902 plus.n69 plus.t1 19.8005
R20903 plus.n71 plus.t0 19.8005
R20904 plus.n71 plus.t2 19.8005
R20905 plus plus.n73 14.3678
R20906 plus.n43 plus.n42 14.1472
R20907 plus.n11 plus.n10 14.1472
R20908 plus.n68 plus.n33 11.7259
R20909 plus.n73 plus.n72 5.40567
R20910 plus.n65 plus.n64 2.19141
R20911 plus.n31 plus.n30 2.19141
R20912 plus.n73 plus.n68 1.188
R20913 plus.n48 plus.n39 0.730803
R20914 plus.n58 plus.n37 0.730803
R20915 plus.n24 plus.n23 0.730803
R20916 plus.n17 plus.n16 0.730803
R20917 plus.n72 plus.n70 0.716017
R20918 plus.n45 plus.n44 0.189894
R20919 plus.n45 plus.n40 0.189894
R20920 plus.n49 plus.n40 0.189894
R20921 plus.n50 plus.n49 0.189894
R20922 plus.n51 plus.n50 0.189894
R20923 plus.n51 plus.n38 0.189894
R20924 plus.n55 plus.n38 0.189894
R20925 plus.n56 plus.n55 0.189894
R20926 plus.n57 plus.n56 0.189894
R20927 plus.n57 plus.n36 0.189894
R20928 plus.n61 plus.n36 0.189894
R20929 plus.n62 plus.n61 0.189894
R20930 plus.n63 plus.n62 0.189894
R20931 plus.n63 plus.n34 0.189894
R20932 plus.n67 plus.n34 0.189894
R20933 plus.n33 plus.n0 0.189894
R20934 plus.n1 plus.n0 0.189894
R20935 plus.n2 plus.n1 0.189894
R20936 plus.n27 plus.n2 0.189894
R20937 plus.n27 plus.n26 0.189894
R20938 plus.n26 plus.n25 0.189894
R20939 plus.n25 plus.n4 0.189894
R20940 plus.n5 plus.n4 0.189894
R20941 plus.n20 plus.n5 0.189894
R20942 plus.n20 plus.n19 0.189894
R20943 plus.n19 plus.n18 0.189894
R20944 plus.n18 plus.n7 0.189894
R20945 plus.n8 plus.n7 0.189894
R20946 plus.n13 plus.n8 0.189894
R20947 plus.n13 plus.n12 0.189894
R20948 outputibias.n27 outputibias.n1 289.615
R20949 outputibias.n58 outputibias.n32 289.615
R20950 outputibias.n90 outputibias.n64 289.615
R20951 outputibias.n122 outputibias.n96 289.615
R20952 outputibias.n28 outputibias.n27 185
R20953 outputibias.n26 outputibias.n25 185
R20954 outputibias.n5 outputibias.n4 185
R20955 outputibias.n20 outputibias.n19 185
R20956 outputibias.n18 outputibias.n17 185
R20957 outputibias.n9 outputibias.n8 185
R20958 outputibias.n12 outputibias.n11 185
R20959 outputibias.n59 outputibias.n58 185
R20960 outputibias.n57 outputibias.n56 185
R20961 outputibias.n36 outputibias.n35 185
R20962 outputibias.n51 outputibias.n50 185
R20963 outputibias.n49 outputibias.n48 185
R20964 outputibias.n40 outputibias.n39 185
R20965 outputibias.n43 outputibias.n42 185
R20966 outputibias.n91 outputibias.n90 185
R20967 outputibias.n89 outputibias.n88 185
R20968 outputibias.n68 outputibias.n67 185
R20969 outputibias.n83 outputibias.n82 185
R20970 outputibias.n81 outputibias.n80 185
R20971 outputibias.n72 outputibias.n71 185
R20972 outputibias.n75 outputibias.n74 185
R20973 outputibias.n123 outputibias.n122 185
R20974 outputibias.n121 outputibias.n120 185
R20975 outputibias.n100 outputibias.n99 185
R20976 outputibias.n115 outputibias.n114 185
R20977 outputibias.n113 outputibias.n112 185
R20978 outputibias.n104 outputibias.n103 185
R20979 outputibias.n107 outputibias.n106 185
R20980 outputibias.n0 outputibias.t10 178.945
R20981 outputibias.n133 outputibias.t8 177.018
R20982 outputibias.n132 outputibias.t11 177.018
R20983 outputibias.n0 outputibias.t9 177.018
R20984 outputibias.t7 outputibias.n10 147.661
R20985 outputibias.t1 outputibias.n41 147.661
R20986 outputibias.t3 outputibias.n73 147.661
R20987 outputibias.t5 outputibias.n105 147.661
R20988 outputibias.n128 outputibias.t6 132.363
R20989 outputibias.n128 outputibias.t0 130.436
R20990 outputibias.n129 outputibias.t2 130.436
R20991 outputibias.n130 outputibias.t4 130.436
R20992 outputibias.n27 outputibias.n26 104.615
R20993 outputibias.n26 outputibias.n4 104.615
R20994 outputibias.n19 outputibias.n4 104.615
R20995 outputibias.n19 outputibias.n18 104.615
R20996 outputibias.n18 outputibias.n8 104.615
R20997 outputibias.n11 outputibias.n8 104.615
R20998 outputibias.n58 outputibias.n57 104.615
R20999 outputibias.n57 outputibias.n35 104.615
R21000 outputibias.n50 outputibias.n35 104.615
R21001 outputibias.n50 outputibias.n49 104.615
R21002 outputibias.n49 outputibias.n39 104.615
R21003 outputibias.n42 outputibias.n39 104.615
R21004 outputibias.n90 outputibias.n89 104.615
R21005 outputibias.n89 outputibias.n67 104.615
R21006 outputibias.n82 outputibias.n67 104.615
R21007 outputibias.n82 outputibias.n81 104.615
R21008 outputibias.n81 outputibias.n71 104.615
R21009 outputibias.n74 outputibias.n71 104.615
R21010 outputibias.n122 outputibias.n121 104.615
R21011 outputibias.n121 outputibias.n99 104.615
R21012 outputibias.n114 outputibias.n99 104.615
R21013 outputibias.n114 outputibias.n113 104.615
R21014 outputibias.n113 outputibias.n103 104.615
R21015 outputibias.n106 outputibias.n103 104.615
R21016 outputibias.n63 outputibias.n31 95.6354
R21017 outputibias.n63 outputibias.n62 94.6732
R21018 outputibias.n95 outputibias.n94 94.6732
R21019 outputibias.n127 outputibias.n126 94.6732
R21020 outputibias.n11 outputibias.t7 52.3082
R21021 outputibias.n42 outputibias.t1 52.3082
R21022 outputibias.n74 outputibias.t3 52.3082
R21023 outputibias.n106 outputibias.t5 52.3082
R21024 outputibias.n12 outputibias.n10 15.6674
R21025 outputibias.n43 outputibias.n41 15.6674
R21026 outputibias.n75 outputibias.n73 15.6674
R21027 outputibias.n107 outputibias.n105 15.6674
R21028 outputibias.n13 outputibias.n9 12.8005
R21029 outputibias.n44 outputibias.n40 12.8005
R21030 outputibias.n76 outputibias.n72 12.8005
R21031 outputibias.n108 outputibias.n104 12.8005
R21032 outputibias.n17 outputibias.n16 12.0247
R21033 outputibias.n48 outputibias.n47 12.0247
R21034 outputibias.n80 outputibias.n79 12.0247
R21035 outputibias.n112 outputibias.n111 12.0247
R21036 outputibias.n20 outputibias.n7 11.249
R21037 outputibias.n51 outputibias.n38 11.249
R21038 outputibias.n83 outputibias.n70 11.249
R21039 outputibias.n115 outputibias.n102 11.249
R21040 outputibias.n21 outputibias.n5 10.4732
R21041 outputibias.n52 outputibias.n36 10.4732
R21042 outputibias.n84 outputibias.n68 10.4732
R21043 outputibias.n116 outputibias.n100 10.4732
R21044 outputibias.n25 outputibias.n24 9.69747
R21045 outputibias.n56 outputibias.n55 9.69747
R21046 outputibias.n88 outputibias.n87 9.69747
R21047 outputibias.n120 outputibias.n119 9.69747
R21048 outputibias.n31 outputibias.n30 9.45567
R21049 outputibias.n62 outputibias.n61 9.45567
R21050 outputibias.n94 outputibias.n93 9.45567
R21051 outputibias.n126 outputibias.n125 9.45567
R21052 outputibias.n30 outputibias.n29 9.3005
R21053 outputibias.n3 outputibias.n2 9.3005
R21054 outputibias.n24 outputibias.n23 9.3005
R21055 outputibias.n22 outputibias.n21 9.3005
R21056 outputibias.n7 outputibias.n6 9.3005
R21057 outputibias.n16 outputibias.n15 9.3005
R21058 outputibias.n14 outputibias.n13 9.3005
R21059 outputibias.n61 outputibias.n60 9.3005
R21060 outputibias.n34 outputibias.n33 9.3005
R21061 outputibias.n55 outputibias.n54 9.3005
R21062 outputibias.n53 outputibias.n52 9.3005
R21063 outputibias.n38 outputibias.n37 9.3005
R21064 outputibias.n47 outputibias.n46 9.3005
R21065 outputibias.n45 outputibias.n44 9.3005
R21066 outputibias.n93 outputibias.n92 9.3005
R21067 outputibias.n66 outputibias.n65 9.3005
R21068 outputibias.n87 outputibias.n86 9.3005
R21069 outputibias.n85 outputibias.n84 9.3005
R21070 outputibias.n70 outputibias.n69 9.3005
R21071 outputibias.n79 outputibias.n78 9.3005
R21072 outputibias.n77 outputibias.n76 9.3005
R21073 outputibias.n125 outputibias.n124 9.3005
R21074 outputibias.n98 outputibias.n97 9.3005
R21075 outputibias.n119 outputibias.n118 9.3005
R21076 outputibias.n117 outputibias.n116 9.3005
R21077 outputibias.n102 outputibias.n101 9.3005
R21078 outputibias.n111 outputibias.n110 9.3005
R21079 outputibias.n109 outputibias.n108 9.3005
R21080 outputibias.n28 outputibias.n3 8.92171
R21081 outputibias.n59 outputibias.n34 8.92171
R21082 outputibias.n91 outputibias.n66 8.92171
R21083 outputibias.n123 outputibias.n98 8.92171
R21084 outputibias.n29 outputibias.n1 8.14595
R21085 outputibias.n60 outputibias.n32 8.14595
R21086 outputibias.n92 outputibias.n64 8.14595
R21087 outputibias.n124 outputibias.n96 8.14595
R21088 outputibias.n31 outputibias.n1 5.81868
R21089 outputibias.n62 outputibias.n32 5.81868
R21090 outputibias.n94 outputibias.n64 5.81868
R21091 outputibias.n126 outputibias.n96 5.81868
R21092 outputibias.n131 outputibias.n130 5.20947
R21093 outputibias.n29 outputibias.n28 5.04292
R21094 outputibias.n60 outputibias.n59 5.04292
R21095 outputibias.n92 outputibias.n91 5.04292
R21096 outputibias.n124 outputibias.n123 5.04292
R21097 outputibias.n131 outputibias.n127 4.42209
R21098 outputibias.n14 outputibias.n10 4.38594
R21099 outputibias.n45 outputibias.n41 4.38594
R21100 outputibias.n77 outputibias.n73 4.38594
R21101 outputibias.n109 outputibias.n105 4.38594
R21102 outputibias.n132 outputibias.n131 4.28454
R21103 outputibias.n25 outputibias.n3 4.26717
R21104 outputibias.n56 outputibias.n34 4.26717
R21105 outputibias.n88 outputibias.n66 4.26717
R21106 outputibias.n120 outputibias.n98 4.26717
R21107 outputibias.n24 outputibias.n5 3.49141
R21108 outputibias.n55 outputibias.n36 3.49141
R21109 outputibias.n87 outputibias.n68 3.49141
R21110 outputibias.n119 outputibias.n100 3.49141
R21111 outputibias.n21 outputibias.n20 2.71565
R21112 outputibias.n52 outputibias.n51 2.71565
R21113 outputibias.n84 outputibias.n83 2.71565
R21114 outputibias.n116 outputibias.n115 2.71565
R21115 outputibias.n17 outputibias.n7 1.93989
R21116 outputibias.n48 outputibias.n38 1.93989
R21117 outputibias.n80 outputibias.n70 1.93989
R21118 outputibias.n112 outputibias.n102 1.93989
R21119 outputibias.n130 outputibias.n129 1.9266
R21120 outputibias.n129 outputibias.n128 1.9266
R21121 outputibias.n133 outputibias.n132 1.92658
R21122 outputibias.n134 outputibias.n133 1.29913
R21123 outputibias.n16 outputibias.n9 1.16414
R21124 outputibias.n47 outputibias.n40 1.16414
R21125 outputibias.n79 outputibias.n72 1.16414
R21126 outputibias.n111 outputibias.n104 1.16414
R21127 outputibias.n127 outputibias.n95 0.962709
R21128 outputibias.n95 outputibias.n63 0.962709
R21129 outputibias.n13 outputibias.n12 0.388379
R21130 outputibias.n44 outputibias.n43 0.388379
R21131 outputibias.n76 outputibias.n75 0.388379
R21132 outputibias.n108 outputibias.n107 0.388379
R21133 outputibias.n134 outputibias.n0 0.337251
R21134 outputibias outputibias.n134 0.302375
R21135 outputibias.n30 outputibias.n2 0.155672
R21136 outputibias.n23 outputibias.n2 0.155672
R21137 outputibias.n23 outputibias.n22 0.155672
R21138 outputibias.n22 outputibias.n6 0.155672
R21139 outputibias.n15 outputibias.n6 0.155672
R21140 outputibias.n15 outputibias.n14 0.155672
R21141 outputibias.n61 outputibias.n33 0.155672
R21142 outputibias.n54 outputibias.n33 0.155672
R21143 outputibias.n54 outputibias.n53 0.155672
R21144 outputibias.n53 outputibias.n37 0.155672
R21145 outputibias.n46 outputibias.n37 0.155672
R21146 outputibias.n46 outputibias.n45 0.155672
R21147 outputibias.n93 outputibias.n65 0.155672
R21148 outputibias.n86 outputibias.n65 0.155672
R21149 outputibias.n86 outputibias.n85 0.155672
R21150 outputibias.n85 outputibias.n69 0.155672
R21151 outputibias.n78 outputibias.n69 0.155672
R21152 outputibias.n78 outputibias.n77 0.155672
R21153 outputibias.n125 outputibias.n97 0.155672
R21154 outputibias.n118 outputibias.n97 0.155672
R21155 outputibias.n118 outputibias.n117 0.155672
R21156 outputibias.n117 outputibias.n101 0.155672
R21157 outputibias.n110 outputibias.n101 0.155672
R21158 outputibias.n110 outputibias.n109 0.155672
R21159 output.n41 output.n15 289.615
R21160 output.n72 output.n46 289.615
R21161 output.n104 output.n78 289.615
R21162 output.n136 output.n110 289.615
R21163 output.n77 output.n45 197.26
R21164 output.n77 output.n76 196.298
R21165 output.n109 output.n108 196.298
R21166 output.n141 output.n140 196.298
R21167 output.n42 output.n41 185
R21168 output.n40 output.n39 185
R21169 output.n19 output.n18 185
R21170 output.n34 output.n33 185
R21171 output.n32 output.n31 185
R21172 output.n23 output.n22 185
R21173 output.n26 output.n25 185
R21174 output.n73 output.n72 185
R21175 output.n71 output.n70 185
R21176 output.n50 output.n49 185
R21177 output.n65 output.n64 185
R21178 output.n63 output.n62 185
R21179 output.n54 output.n53 185
R21180 output.n57 output.n56 185
R21181 output.n105 output.n104 185
R21182 output.n103 output.n102 185
R21183 output.n82 output.n81 185
R21184 output.n97 output.n96 185
R21185 output.n95 output.n94 185
R21186 output.n86 output.n85 185
R21187 output.n89 output.n88 185
R21188 output.n137 output.n136 185
R21189 output.n135 output.n134 185
R21190 output.n114 output.n113 185
R21191 output.n129 output.n128 185
R21192 output.n127 output.n126 185
R21193 output.n118 output.n117 185
R21194 output.n121 output.n120 185
R21195 output.t17 output.n24 147.661
R21196 output.t18 output.n55 147.661
R21197 output.t19 output.n87 147.661
R21198 output.t16 output.n119 147.661
R21199 output.n41 output.n40 104.615
R21200 output.n40 output.n18 104.615
R21201 output.n33 output.n18 104.615
R21202 output.n33 output.n32 104.615
R21203 output.n32 output.n22 104.615
R21204 output.n25 output.n22 104.615
R21205 output.n72 output.n71 104.615
R21206 output.n71 output.n49 104.615
R21207 output.n64 output.n49 104.615
R21208 output.n64 output.n63 104.615
R21209 output.n63 output.n53 104.615
R21210 output.n56 output.n53 104.615
R21211 output.n104 output.n103 104.615
R21212 output.n103 output.n81 104.615
R21213 output.n96 output.n81 104.615
R21214 output.n96 output.n95 104.615
R21215 output.n95 output.n85 104.615
R21216 output.n88 output.n85 104.615
R21217 output.n136 output.n135 104.615
R21218 output.n135 output.n113 104.615
R21219 output.n128 output.n113 104.615
R21220 output.n128 output.n127 104.615
R21221 output.n127 output.n117 104.615
R21222 output.n120 output.n117 104.615
R21223 output.n1 output.t1 77.056
R21224 output.n14 output.t2 76.6694
R21225 output.n1 output.n0 72.7095
R21226 output.n3 output.n2 72.7095
R21227 output.n5 output.n4 72.7095
R21228 output.n7 output.n6 72.7095
R21229 output.n9 output.n8 72.7095
R21230 output.n11 output.n10 72.7095
R21231 output.n13 output.n12 72.7095
R21232 output.n25 output.t17 52.3082
R21233 output.n56 output.t18 52.3082
R21234 output.n88 output.t19 52.3082
R21235 output.n120 output.t16 52.3082
R21236 output.n26 output.n24 15.6674
R21237 output.n57 output.n55 15.6674
R21238 output.n89 output.n87 15.6674
R21239 output.n121 output.n119 15.6674
R21240 output.n27 output.n23 12.8005
R21241 output.n58 output.n54 12.8005
R21242 output.n90 output.n86 12.8005
R21243 output.n122 output.n118 12.8005
R21244 output.n31 output.n30 12.0247
R21245 output.n62 output.n61 12.0247
R21246 output.n94 output.n93 12.0247
R21247 output.n126 output.n125 12.0247
R21248 output.n34 output.n21 11.249
R21249 output.n65 output.n52 11.249
R21250 output.n97 output.n84 11.249
R21251 output.n129 output.n116 11.249
R21252 output.n35 output.n19 10.4732
R21253 output.n66 output.n50 10.4732
R21254 output.n98 output.n82 10.4732
R21255 output.n130 output.n114 10.4732
R21256 output.n39 output.n38 9.69747
R21257 output.n70 output.n69 9.69747
R21258 output.n102 output.n101 9.69747
R21259 output.n134 output.n133 9.69747
R21260 output.n45 output.n44 9.45567
R21261 output.n76 output.n75 9.45567
R21262 output.n108 output.n107 9.45567
R21263 output.n140 output.n139 9.45567
R21264 output.n44 output.n43 9.3005
R21265 output.n17 output.n16 9.3005
R21266 output.n38 output.n37 9.3005
R21267 output.n36 output.n35 9.3005
R21268 output.n21 output.n20 9.3005
R21269 output.n30 output.n29 9.3005
R21270 output.n28 output.n27 9.3005
R21271 output.n75 output.n74 9.3005
R21272 output.n48 output.n47 9.3005
R21273 output.n69 output.n68 9.3005
R21274 output.n67 output.n66 9.3005
R21275 output.n52 output.n51 9.3005
R21276 output.n61 output.n60 9.3005
R21277 output.n59 output.n58 9.3005
R21278 output.n107 output.n106 9.3005
R21279 output.n80 output.n79 9.3005
R21280 output.n101 output.n100 9.3005
R21281 output.n99 output.n98 9.3005
R21282 output.n84 output.n83 9.3005
R21283 output.n93 output.n92 9.3005
R21284 output.n91 output.n90 9.3005
R21285 output.n139 output.n138 9.3005
R21286 output.n112 output.n111 9.3005
R21287 output.n133 output.n132 9.3005
R21288 output.n131 output.n130 9.3005
R21289 output.n116 output.n115 9.3005
R21290 output.n125 output.n124 9.3005
R21291 output.n123 output.n122 9.3005
R21292 output.n42 output.n17 8.92171
R21293 output.n73 output.n48 8.92171
R21294 output.n105 output.n80 8.92171
R21295 output.n137 output.n112 8.92171
R21296 output output.n141 8.15037
R21297 output.n43 output.n15 8.14595
R21298 output.n74 output.n46 8.14595
R21299 output.n106 output.n78 8.14595
R21300 output.n138 output.n110 8.14595
R21301 output.n45 output.n15 5.81868
R21302 output.n76 output.n46 5.81868
R21303 output.n108 output.n78 5.81868
R21304 output.n140 output.n110 5.81868
R21305 output.n43 output.n42 5.04292
R21306 output.n74 output.n73 5.04292
R21307 output.n106 output.n105 5.04292
R21308 output.n138 output.n137 5.04292
R21309 output.n28 output.n24 4.38594
R21310 output.n59 output.n55 4.38594
R21311 output.n91 output.n87 4.38594
R21312 output.n123 output.n119 4.38594
R21313 output.n39 output.n17 4.26717
R21314 output.n70 output.n48 4.26717
R21315 output.n102 output.n80 4.26717
R21316 output.n134 output.n112 4.26717
R21317 output.n0 output.t12 3.9605
R21318 output.n0 output.t15 3.9605
R21319 output.n2 output.t5 3.9605
R21320 output.n2 output.t4 3.9605
R21321 output.n4 output.t10 3.9605
R21322 output.n4 output.t14 3.9605
R21323 output.n6 output.t3 3.9605
R21324 output.n6 output.t6 3.9605
R21325 output.n8 output.t7 3.9605
R21326 output.n8 output.t13 3.9605
R21327 output.n10 output.t0 3.9605
R21328 output.n10 output.t8 3.9605
R21329 output.n12 output.t11 3.9605
R21330 output.n12 output.t9 3.9605
R21331 output.n38 output.n19 3.49141
R21332 output.n69 output.n50 3.49141
R21333 output.n101 output.n82 3.49141
R21334 output.n133 output.n114 3.49141
R21335 output.n35 output.n34 2.71565
R21336 output.n66 output.n65 2.71565
R21337 output.n98 output.n97 2.71565
R21338 output.n130 output.n129 2.71565
R21339 output.n31 output.n21 1.93989
R21340 output.n62 output.n52 1.93989
R21341 output.n94 output.n84 1.93989
R21342 output.n126 output.n116 1.93989
R21343 output.n30 output.n23 1.16414
R21344 output.n61 output.n54 1.16414
R21345 output.n93 output.n86 1.16414
R21346 output.n125 output.n118 1.16414
R21347 output.n141 output.n109 0.962709
R21348 output.n109 output.n77 0.962709
R21349 output.n27 output.n26 0.388379
R21350 output.n58 output.n57 0.388379
R21351 output.n90 output.n89 0.388379
R21352 output.n122 output.n121 0.388379
R21353 output.n14 output.n13 0.387128
R21354 output.n13 output.n11 0.387128
R21355 output.n11 output.n9 0.387128
R21356 output.n9 output.n7 0.387128
R21357 output.n7 output.n5 0.387128
R21358 output.n5 output.n3 0.387128
R21359 output.n3 output.n1 0.387128
R21360 output.n44 output.n16 0.155672
R21361 output.n37 output.n16 0.155672
R21362 output.n37 output.n36 0.155672
R21363 output.n36 output.n20 0.155672
R21364 output.n29 output.n20 0.155672
R21365 output.n29 output.n28 0.155672
R21366 output.n75 output.n47 0.155672
R21367 output.n68 output.n47 0.155672
R21368 output.n68 output.n67 0.155672
R21369 output.n67 output.n51 0.155672
R21370 output.n60 output.n51 0.155672
R21371 output.n60 output.n59 0.155672
R21372 output.n107 output.n79 0.155672
R21373 output.n100 output.n79 0.155672
R21374 output.n100 output.n99 0.155672
R21375 output.n99 output.n83 0.155672
R21376 output.n92 output.n83 0.155672
R21377 output.n92 output.n91 0.155672
R21378 output.n139 output.n111 0.155672
R21379 output.n132 output.n111 0.155672
R21380 output.n132 output.n131 0.155672
R21381 output.n131 output.n115 0.155672
R21382 output.n124 output.n115 0.155672
R21383 output.n124 output.n123 0.155672
R21384 output output.n14 0.126227
C0 minus diffpairibias 2.98e-19
C1 commonsourceibias output 0.006808f
C2 CSoutput minus 2.75386f
C3 vdd plus 0.065528f
C4 commonsourceibias outputibias 0.003832f
C5 plus diffpairibias 2.75e-19
C6 vdd commonsourceibias 0.004218f
C7 CSoutput plus 0.852171f
C8 commonsourceibias diffpairibias 0.064336f
C9 CSoutput commonsourceibias 42.3358f
C10 minus plus 9.09051f
C11 minus commonsourceibias 0.331305f
C12 plus commonsourceibias 0.276969f
C13 output outputibias 2.34152f
C14 vdd output 7.23429f
C15 CSoutput output 6.13881f
C16 CSoutput outputibias 0.032386f
C17 vdd CSoutput 67.6707f
C18 diffpairibias gnd 60.00273f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.14503p
C22 plus gnd 33.159603f
C23 minus gnd 27.49461f
C24 CSoutput gnd 0.108289p
C25 vdd gnd 0.345061p
C26 output.t1 gnd 0.464308f
C27 output.t12 gnd 0.044422f
C28 output.t15 gnd 0.044422f
C29 output.n0 gnd 0.364624f
C30 output.n1 gnd 0.614102f
C31 output.t5 gnd 0.044422f
C32 output.t4 gnd 0.044422f
C33 output.n2 gnd 0.364624f
C34 output.n3 gnd 0.350265f
C35 output.t10 gnd 0.044422f
C36 output.t14 gnd 0.044422f
C37 output.n4 gnd 0.364624f
C38 output.n5 gnd 0.350265f
C39 output.t3 gnd 0.044422f
C40 output.t6 gnd 0.044422f
C41 output.n6 gnd 0.364624f
C42 output.n7 gnd 0.350265f
C43 output.t7 gnd 0.044422f
C44 output.t13 gnd 0.044422f
C45 output.n8 gnd 0.364624f
C46 output.n9 gnd 0.350265f
C47 output.t0 gnd 0.044422f
C48 output.t8 gnd 0.044422f
C49 output.n10 gnd 0.364624f
C50 output.n11 gnd 0.350265f
C51 output.t11 gnd 0.044422f
C52 output.t9 gnd 0.044422f
C53 output.n12 gnd 0.364624f
C54 output.n13 gnd 0.350265f
C55 output.t2 gnd 0.462979f
C56 output.n14 gnd 0.28994f
C57 output.n15 gnd 0.015803f
C58 output.n16 gnd 0.011243f
C59 output.n17 gnd 0.006041f
C60 output.n18 gnd 0.01428f
C61 output.n19 gnd 0.006397f
C62 output.n20 gnd 0.011243f
C63 output.n21 gnd 0.006041f
C64 output.n22 gnd 0.01428f
C65 output.n23 gnd 0.006397f
C66 output.n24 gnd 0.048111f
C67 output.t17 gnd 0.023274f
C68 output.n25 gnd 0.01071f
C69 output.n26 gnd 0.008435f
C70 output.n27 gnd 0.006041f
C71 output.n28 gnd 0.267512f
C72 output.n29 gnd 0.011243f
C73 output.n30 gnd 0.006041f
C74 output.n31 gnd 0.006397f
C75 output.n32 gnd 0.01428f
C76 output.n33 gnd 0.01428f
C77 output.n34 gnd 0.006397f
C78 output.n35 gnd 0.006041f
C79 output.n36 gnd 0.011243f
C80 output.n37 gnd 0.011243f
C81 output.n38 gnd 0.006041f
C82 output.n39 gnd 0.006397f
C83 output.n40 gnd 0.01428f
C84 output.n41 gnd 0.030913f
C85 output.n42 gnd 0.006397f
C86 output.n43 gnd 0.006041f
C87 output.n44 gnd 0.025987f
C88 output.n45 gnd 0.097665f
C89 output.n46 gnd 0.015803f
C90 output.n47 gnd 0.011243f
C91 output.n48 gnd 0.006041f
C92 output.n49 gnd 0.01428f
C93 output.n50 gnd 0.006397f
C94 output.n51 gnd 0.011243f
C95 output.n52 gnd 0.006041f
C96 output.n53 gnd 0.01428f
C97 output.n54 gnd 0.006397f
C98 output.n55 gnd 0.048111f
C99 output.t18 gnd 0.023274f
C100 output.n56 gnd 0.01071f
C101 output.n57 gnd 0.008435f
C102 output.n58 gnd 0.006041f
C103 output.n59 gnd 0.267512f
C104 output.n60 gnd 0.011243f
C105 output.n61 gnd 0.006041f
C106 output.n62 gnd 0.006397f
C107 output.n63 gnd 0.01428f
C108 output.n64 gnd 0.01428f
C109 output.n65 gnd 0.006397f
C110 output.n66 gnd 0.006041f
C111 output.n67 gnd 0.011243f
C112 output.n68 gnd 0.011243f
C113 output.n69 gnd 0.006041f
C114 output.n70 gnd 0.006397f
C115 output.n71 gnd 0.01428f
C116 output.n72 gnd 0.030913f
C117 output.n73 gnd 0.006397f
C118 output.n74 gnd 0.006041f
C119 output.n75 gnd 0.025987f
C120 output.n76 gnd 0.09306f
C121 output.n77 gnd 1.65264f
C122 output.n78 gnd 0.015803f
C123 output.n79 gnd 0.011243f
C124 output.n80 gnd 0.006041f
C125 output.n81 gnd 0.01428f
C126 output.n82 gnd 0.006397f
C127 output.n83 gnd 0.011243f
C128 output.n84 gnd 0.006041f
C129 output.n85 gnd 0.01428f
C130 output.n86 gnd 0.006397f
C131 output.n87 gnd 0.048111f
C132 output.t19 gnd 0.023274f
C133 output.n88 gnd 0.01071f
C134 output.n89 gnd 0.008435f
C135 output.n90 gnd 0.006041f
C136 output.n91 gnd 0.267512f
C137 output.n92 gnd 0.011243f
C138 output.n93 gnd 0.006041f
C139 output.n94 gnd 0.006397f
C140 output.n95 gnd 0.01428f
C141 output.n96 gnd 0.01428f
C142 output.n97 gnd 0.006397f
C143 output.n98 gnd 0.006041f
C144 output.n99 gnd 0.011243f
C145 output.n100 gnd 0.011243f
C146 output.n101 gnd 0.006041f
C147 output.n102 gnd 0.006397f
C148 output.n103 gnd 0.01428f
C149 output.n104 gnd 0.030913f
C150 output.n105 gnd 0.006397f
C151 output.n106 gnd 0.006041f
C152 output.n107 gnd 0.025987f
C153 output.n108 gnd 0.09306f
C154 output.n109 gnd 0.713089f
C155 output.n110 gnd 0.015803f
C156 output.n111 gnd 0.011243f
C157 output.n112 gnd 0.006041f
C158 output.n113 gnd 0.01428f
C159 output.n114 gnd 0.006397f
C160 output.n115 gnd 0.011243f
C161 output.n116 gnd 0.006041f
C162 output.n117 gnd 0.01428f
C163 output.n118 gnd 0.006397f
C164 output.n119 gnd 0.048111f
C165 output.t16 gnd 0.023274f
C166 output.n120 gnd 0.01071f
C167 output.n121 gnd 0.008435f
C168 output.n122 gnd 0.006041f
C169 output.n123 gnd 0.267512f
C170 output.n124 gnd 0.011243f
C171 output.n125 gnd 0.006041f
C172 output.n126 gnd 0.006397f
C173 output.n127 gnd 0.01428f
C174 output.n128 gnd 0.01428f
C175 output.n129 gnd 0.006397f
C176 output.n130 gnd 0.006041f
C177 output.n131 gnd 0.011243f
C178 output.n132 gnd 0.011243f
C179 output.n133 gnd 0.006041f
C180 output.n134 gnd 0.006397f
C181 output.n135 gnd 0.01428f
C182 output.n136 gnd 0.030913f
C183 output.n137 gnd 0.006397f
C184 output.n138 gnd 0.006041f
C185 output.n139 gnd 0.025987f
C186 output.n140 gnd 0.09306f
C187 output.n141 gnd 1.67353f
C188 outputibias.t9 gnd 0.11477f
C189 outputibias.t10 gnd 0.115567f
C190 outputibias.n0 gnd 0.130108f
C191 outputibias.n1 gnd 0.001372f
C192 outputibias.n2 gnd 9.76e-19
C193 outputibias.n3 gnd 5.24e-19
C194 outputibias.n4 gnd 0.001239f
C195 outputibias.n5 gnd 5.55e-19
C196 outputibias.n6 gnd 9.76e-19
C197 outputibias.n7 gnd 5.24e-19
C198 outputibias.n8 gnd 0.001239f
C199 outputibias.n9 gnd 5.55e-19
C200 outputibias.n10 gnd 0.004176f
C201 outputibias.t7 gnd 0.00202f
C202 outputibias.n11 gnd 9.3e-19
C203 outputibias.n12 gnd 7.32e-19
C204 outputibias.n13 gnd 5.24e-19
C205 outputibias.n14 gnd 0.02322f
C206 outputibias.n15 gnd 9.76e-19
C207 outputibias.n16 gnd 5.24e-19
C208 outputibias.n17 gnd 5.55e-19
C209 outputibias.n18 gnd 0.001239f
C210 outputibias.n19 gnd 0.001239f
C211 outputibias.n20 gnd 5.55e-19
C212 outputibias.n21 gnd 5.24e-19
C213 outputibias.n22 gnd 9.76e-19
C214 outputibias.n23 gnd 9.76e-19
C215 outputibias.n24 gnd 5.24e-19
C216 outputibias.n25 gnd 5.55e-19
C217 outputibias.n26 gnd 0.001239f
C218 outputibias.n27 gnd 0.002683f
C219 outputibias.n28 gnd 5.55e-19
C220 outputibias.n29 gnd 5.24e-19
C221 outputibias.n30 gnd 0.002256f
C222 outputibias.n31 gnd 0.005781f
C223 outputibias.n32 gnd 0.001372f
C224 outputibias.n33 gnd 9.76e-19
C225 outputibias.n34 gnd 5.24e-19
C226 outputibias.n35 gnd 0.001239f
C227 outputibias.n36 gnd 5.55e-19
C228 outputibias.n37 gnd 9.76e-19
C229 outputibias.n38 gnd 5.24e-19
C230 outputibias.n39 gnd 0.001239f
C231 outputibias.n40 gnd 5.55e-19
C232 outputibias.n41 gnd 0.004176f
C233 outputibias.t1 gnd 0.00202f
C234 outputibias.n42 gnd 9.3e-19
C235 outputibias.n43 gnd 7.32e-19
C236 outputibias.n44 gnd 5.24e-19
C237 outputibias.n45 gnd 0.02322f
C238 outputibias.n46 gnd 9.76e-19
C239 outputibias.n47 gnd 5.24e-19
C240 outputibias.n48 gnd 5.55e-19
C241 outputibias.n49 gnd 0.001239f
C242 outputibias.n50 gnd 0.001239f
C243 outputibias.n51 gnd 5.55e-19
C244 outputibias.n52 gnd 5.24e-19
C245 outputibias.n53 gnd 9.76e-19
C246 outputibias.n54 gnd 9.76e-19
C247 outputibias.n55 gnd 5.24e-19
C248 outputibias.n56 gnd 5.55e-19
C249 outputibias.n57 gnd 0.001239f
C250 outputibias.n58 gnd 0.002683f
C251 outputibias.n59 gnd 5.55e-19
C252 outputibias.n60 gnd 5.24e-19
C253 outputibias.n61 gnd 0.002256f
C254 outputibias.n62 gnd 0.005197f
C255 outputibias.n63 gnd 0.121892f
C256 outputibias.n64 gnd 0.001372f
C257 outputibias.n65 gnd 9.76e-19
C258 outputibias.n66 gnd 5.24e-19
C259 outputibias.n67 gnd 0.001239f
C260 outputibias.n68 gnd 5.55e-19
C261 outputibias.n69 gnd 9.76e-19
C262 outputibias.n70 gnd 5.24e-19
C263 outputibias.n71 gnd 0.001239f
C264 outputibias.n72 gnd 5.55e-19
C265 outputibias.n73 gnd 0.004176f
C266 outputibias.t3 gnd 0.00202f
C267 outputibias.n74 gnd 9.3e-19
C268 outputibias.n75 gnd 7.32e-19
C269 outputibias.n76 gnd 5.24e-19
C270 outputibias.n77 gnd 0.02322f
C271 outputibias.n78 gnd 9.76e-19
C272 outputibias.n79 gnd 5.24e-19
C273 outputibias.n80 gnd 5.55e-19
C274 outputibias.n81 gnd 0.001239f
C275 outputibias.n82 gnd 0.001239f
C276 outputibias.n83 gnd 5.55e-19
C277 outputibias.n84 gnd 5.24e-19
C278 outputibias.n85 gnd 9.76e-19
C279 outputibias.n86 gnd 9.76e-19
C280 outputibias.n87 gnd 5.24e-19
C281 outputibias.n88 gnd 5.55e-19
C282 outputibias.n89 gnd 0.001239f
C283 outputibias.n90 gnd 0.002683f
C284 outputibias.n91 gnd 5.55e-19
C285 outputibias.n92 gnd 5.24e-19
C286 outputibias.n93 gnd 0.002256f
C287 outputibias.n94 gnd 0.005197f
C288 outputibias.n95 gnd 0.064513f
C289 outputibias.n96 gnd 0.001372f
C290 outputibias.n97 gnd 9.76e-19
C291 outputibias.n98 gnd 5.24e-19
C292 outputibias.n99 gnd 0.001239f
C293 outputibias.n100 gnd 5.55e-19
C294 outputibias.n101 gnd 9.76e-19
C295 outputibias.n102 gnd 5.24e-19
C296 outputibias.n103 gnd 0.001239f
C297 outputibias.n104 gnd 5.55e-19
C298 outputibias.n105 gnd 0.004176f
C299 outputibias.t5 gnd 0.00202f
C300 outputibias.n106 gnd 9.3e-19
C301 outputibias.n107 gnd 7.32e-19
C302 outputibias.n108 gnd 5.24e-19
C303 outputibias.n109 gnd 0.02322f
C304 outputibias.n110 gnd 9.76e-19
C305 outputibias.n111 gnd 5.24e-19
C306 outputibias.n112 gnd 5.55e-19
C307 outputibias.n113 gnd 0.001239f
C308 outputibias.n114 gnd 0.001239f
C309 outputibias.n115 gnd 5.55e-19
C310 outputibias.n116 gnd 5.24e-19
C311 outputibias.n117 gnd 9.76e-19
C312 outputibias.n118 gnd 9.76e-19
C313 outputibias.n119 gnd 5.24e-19
C314 outputibias.n120 gnd 5.55e-19
C315 outputibias.n121 gnd 0.001239f
C316 outputibias.n122 gnd 0.002683f
C317 outputibias.n123 gnd 5.55e-19
C318 outputibias.n124 gnd 5.24e-19
C319 outputibias.n125 gnd 0.002256f
C320 outputibias.n126 gnd 0.005197f
C321 outputibias.n127 gnd 0.084814f
C322 outputibias.t4 gnd 0.108319f
C323 outputibias.t2 gnd 0.108319f
C324 outputibias.t0 gnd 0.108319f
C325 outputibias.t6 gnd 0.109238f
C326 outputibias.n128 gnd 0.134674f
C327 outputibias.n129 gnd 0.07244f
C328 outputibias.n130 gnd 0.079818f
C329 outputibias.n131 gnd 0.164901f
C330 outputibias.t11 gnd 0.11477f
C331 outputibias.n132 gnd 0.067481f
C332 outputibias.t8 gnd 0.11477f
C333 outputibias.n133 gnd 0.065115f
C334 outputibias.n134 gnd 0.029159f
C335 plus.n0 gnd 0.023974f
C336 plus.t23 gnd 0.242206f
C337 plus.n1 gnd 0.023974f
C338 plus.t13 gnd 0.242206f
C339 plus.n2 gnd 0.023974f
C340 plus.t27 gnd 0.242206f
C341 plus.t22 gnd 0.242206f
C342 plus.n3 gnd 0.111979f
C343 plus.n4 gnd 0.023974f
C344 plus.t7 gnd 0.242206f
C345 plus.n5 gnd 0.023974f
C346 plus.t18 gnd 0.242206f
C347 plus.t14 gnd 0.242206f
C348 plus.n6 gnd 0.111906f
C349 plus.n7 gnd 0.023974f
C350 plus.t24 gnd 0.242206f
C351 plus.n8 gnd 0.023974f
C352 plus.t17 gnd 0.242206f
C353 plus.t9 gnd 0.242206f
C354 plus.n9 gnd 0.111758f
C355 plus.t12 gnd 0.248727f
C356 plus.t15 gnd 0.242206f
C357 plus.n10 gnd 0.114594f
C358 plus.n11 gnd 0.103731f
C359 plus.n12 gnd 0.097344f
C360 plus.n13 gnd 0.023974f
C361 plus.n14 gnd 0.00544f
C362 plus.n15 gnd 0.111979f
C363 plus.n16 gnd 0.00544f
C364 plus.n17 gnd 0.109541f
C365 plus.n18 gnd 0.023974f
C366 plus.n19 gnd 0.023974f
C367 plus.n20 gnd 0.023974f
C368 plus.n21 gnd 0.00544f
C369 plus.n22 gnd 0.111906f
C370 plus.n23 gnd 0.109541f
C371 plus.n24 gnd 0.00544f
C372 plus.n25 gnd 0.023974f
C373 plus.n26 gnd 0.023974f
C374 plus.n27 gnd 0.023974f
C375 plus.n28 gnd 0.00544f
C376 plus.n29 gnd 0.111758f
C377 plus.n30 gnd 0.109688f
C378 plus.n31 gnd 0.00544f
C379 plus.n32 gnd 0.109245f
C380 plus.n33 gnd 0.262859f
C381 plus.n34 gnd 0.023974f
C382 plus.t16 gnd 0.242206f
C383 plus.n35 gnd 0.111758f
C384 plus.t28 gnd 0.242206f
C385 plus.n36 gnd 0.023974f
C386 plus.t19 gnd 0.242206f
C387 plus.n37 gnd 0.109541f
C388 plus.n38 gnd 0.023974f
C389 plus.t11 gnd 0.242206f
C390 plus.n39 gnd 0.109541f
C391 plus.t6 gnd 0.242206f
C392 plus.n40 gnd 0.023974f
C393 plus.t20 gnd 0.242206f
C394 plus.n41 gnd 0.111758f
C395 plus.t25 gnd 0.248727f
C396 plus.t5 gnd 0.242206f
C397 plus.n42 gnd 0.114594f
C398 plus.n43 gnd 0.103731f
C399 plus.n44 gnd 0.097344f
C400 plus.n45 gnd 0.023974f
C401 plus.n46 gnd 0.00544f
C402 plus.t26 gnd 0.242206f
C403 plus.n47 gnd 0.111979f
C404 plus.n48 gnd 0.00544f
C405 plus.n49 gnd 0.023974f
C406 plus.n50 gnd 0.023974f
C407 plus.n51 gnd 0.023974f
C408 plus.n52 gnd 0.111906f
C409 plus.n53 gnd 0.00544f
C410 plus.t10 gnd 0.242206f
C411 plus.n54 gnd 0.111906f
C412 plus.n55 gnd 0.023974f
C413 plus.n56 gnd 0.023974f
C414 plus.n57 gnd 0.023974f
C415 plus.n58 gnd 0.00544f
C416 plus.t8 gnd 0.242206f
C417 plus.n59 gnd 0.111979f
C418 plus.n60 gnd 0.00544f
C419 plus.n61 gnd 0.023974f
C420 plus.n62 gnd 0.023974f
C421 plus.n63 gnd 0.023974f
C422 plus.n64 gnd 0.109688f
C423 plus.n65 gnd 0.00544f
C424 plus.t21 gnd 0.242206f
C425 plus.n66 gnd 0.109245f
C426 plus.n67 gnd 0.717857f
C427 plus.n68 gnd 1.0941f
C428 plus.t3 gnd 0.041386f
C429 plus.t4 gnd 0.00739f
C430 plus.t1 gnd 0.00739f
C431 plus.n69 gnd 0.023968f
C432 plus.n70 gnd 0.18607f
C433 plus.t0 gnd 0.00739f
C434 plus.t2 gnd 0.00739f
C435 plus.n71 gnd 0.023968f
C436 plus.n72 gnd 0.139668f
C437 plus.n73 gnd 2.65334f
C438 minus.n0 gnd 0.033094f
C439 minus.t27 gnd 0.33435f
C440 minus.n1 gnd 0.154274f
C441 minus.n2 gnd 0.033094f
C442 minus.t6 gnd 0.33435f
C443 minus.n3 gnd 0.151214f
C444 minus.n4 gnd 0.033094f
C445 minus.t24 gnd 0.33435f
C446 minus.n5 gnd 0.151214f
C447 minus.n6 gnd 0.033094f
C448 minus.t8 gnd 0.33435f
C449 minus.n7 gnd 0.154274f
C450 minus.t12 gnd 0.343352f
C451 minus.t18 gnd 0.33435f
C452 minus.n8 gnd 0.15819f
C453 minus.n9 gnd 0.143194f
C454 minus.n10 gnd 0.134377f
C455 minus.n11 gnd 0.033094f
C456 minus.n12 gnd 0.00751f
C457 minus.t13 gnd 0.33435f
C458 minus.n13 gnd 0.154581f
C459 minus.n14 gnd 0.00751f
C460 minus.n15 gnd 0.033094f
C461 minus.n16 gnd 0.033094f
C462 minus.n17 gnd 0.033094f
C463 minus.t19 gnd 0.33435f
C464 minus.n18 gnd 0.154479f
C465 minus.n19 gnd 0.00751f
C466 minus.t22 gnd 0.33435f
C467 minus.n20 gnd 0.154479f
C468 minus.n21 gnd 0.033094f
C469 minus.n22 gnd 0.033094f
C470 minus.n23 gnd 0.033094f
C471 minus.n24 gnd 0.00751f
C472 minus.t20 gnd 0.33435f
C473 minus.n25 gnd 0.154581f
C474 minus.n26 gnd 0.00751f
C475 minus.n27 gnd 0.033094f
C476 minus.n28 gnd 0.033094f
C477 minus.n29 gnd 0.033094f
C478 minus.t16 gnd 0.33435f
C479 minus.n30 gnd 0.151418f
C480 minus.n31 gnd 0.00751f
C481 minus.t9 gnd 0.33435f
C482 minus.n32 gnd 0.150806f
C483 minus.n33 gnd 0.371412f
C484 minus.n34 gnd 0.033094f
C485 minus.t15 gnd 0.33435f
C486 minus.t28 gnd 0.33435f
C487 minus.n35 gnd 0.033094f
C488 minus.t21 gnd 0.33435f
C489 minus.n36 gnd 0.033094f
C490 minus.t14 gnd 0.33435f
C491 minus.n37 gnd 0.154581f
C492 minus.n38 gnd 0.033094f
C493 minus.t23 gnd 0.33435f
C494 minus.t11 gnd 0.33435f
C495 minus.n39 gnd 0.033094f
C496 minus.t5 gnd 0.33435f
C497 minus.n40 gnd 0.154479f
C498 minus.n41 gnd 0.033094f
C499 minus.t17 gnd 0.33435f
C500 minus.t10 gnd 0.33435f
C501 minus.n42 gnd 0.033094f
C502 minus.t25 gnd 0.33435f
C503 minus.n43 gnd 0.154274f
C504 minus.t26 gnd 0.343352f
C505 minus.t7 gnd 0.33435f
C506 minus.n44 gnd 0.15819f
C507 minus.n45 gnd 0.143194f
C508 minus.n46 gnd 0.134377f
C509 minus.n47 gnd 0.033094f
C510 minus.n48 gnd 0.00751f
C511 minus.n49 gnd 0.154581f
C512 minus.n50 gnd 0.00751f
C513 minus.n51 gnd 0.151214f
C514 minus.n52 gnd 0.033094f
C515 minus.n53 gnd 0.033094f
C516 minus.n54 gnd 0.033094f
C517 minus.n55 gnd 0.00751f
C518 minus.n56 gnd 0.154479f
C519 minus.n57 gnd 0.151214f
C520 minus.n58 gnd 0.00751f
C521 minus.n59 gnd 0.033094f
C522 minus.n60 gnd 0.033094f
C523 minus.n61 gnd 0.033094f
C524 minus.n62 gnd 0.00751f
C525 minus.n63 gnd 0.154274f
C526 minus.n64 gnd 0.151418f
C527 minus.n65 gnd 0.00751f
C528 minus.n66 gnd 0.150806f
C529 minus.n67 gnd 1.00426f
C530 minus.n68 gnd 1.52338f
C531 minus.t1 gnd 0.010202f
C532 minus.t4 gnd 0.010202f
C533 minus.n69 gnd 0.033547f
C534 minus.t2 gnd 0.010202f
C535 minus.t0 gnd 0.010202f
C536 minus.n70 gnd 0.033087f
C537 minus.n71 gnd 0.282383f
C538 minus.t3 gnd 0.056783f
C539 minus.n72 gnd 0.154094f
C540 minus.n73 gnd 2.07222f
C541 a_n3827_n3924.n0 gnd 1.10033f
C542 a_n3827_n3924.n1 gnd 0.958536f
C543 a_n3827_n3924.t31 gnd 1.06719f
C544 a_n3827_n3924.n2 gnd 0.920943f
C545 a_n3827_n3924.t26 gnd 0.102682f
C546 a_n3827_n3924.t52 gnd 0.102682f
C547 a_n3827_n3924.n3 gnd 0.838616f
C548 a_n3827_n3924.n4 gnd 0.340114f
C549 a_n3827_n3924.t28 gnd 0.102682f
C550 a_n3827_n3924.t30 gnd 0.102682f
C551 a_n3827_n3924.n5 gnd 0.838616f
C552 a_n3827_n3924.n6 gnd 0.340114f
C553 a_n3827_n3924.t29 gnd 0.102682f
C554 a_n3827_n3924.t37 gnd 0.102682f
C555 a_n3827_n3924.n7 gnd 0.838616f
C556 a_n3827_n3924.n8 gnd 0.340114f
C557 a_n3827_n3924.t8 gnd 0.102682f
C558 a_n3827_n3924.t51 gnd 0.102682f
C559 a_n3827_n3924.n9 gnd 0.838616f
C560 a_n3827_n3924.n10 gnd 0.340114f
C561 a_n3827_n3924.t24 gnd 0.102682f
C562 a_n3827_n3924.t54 gnd 0.102682f
C563 a_n3827_n3924.n11 gnd 0.838616f
C564 a_n3827_n3924.n12 gnd 0.340114f
C565 a_n3827_n3924.t21 gnd 1.06719f
C566 a_n3827_n3924.n13 gnd 0.362194f
C567 a_n3827_n3924.t45 gnd 1.06719f
C568 a_n3827_n3924.n14 gnd 0.362194f
C569 a_n3827_n3924.t44 gnd 0.102682f
C570 a_n3827_n3924.t6 gnd 0.102682f
C571 a_n3827_n3924.n15 gnd 0.838616f
C572 a_n3827_n3924.n16 gnd 0.340114f
C573 a_n3827_n3924.t32 gnd 0.102682f
C574 a_n3827_n3924.t43 gnd 0.102682f
C575 a_n3827_n3924.n17 gnd 0.838616f
C576 a_n3827_n3924.n18 gnd 0.340114f
C577 a_n3827_n3924.t42 gnd 0.102682f
C578 a_n3827_n3924.t39 gnd 0.102682f
C579 a_n3827_n3924.n19 gnd 0.838616f
C580 a_n3827_n3924.n20 gnd 0.340114f
C581 a_n3827_n3924.t48 gnd 0.102682f
C582 a_n3827_n3924.t0 gnd 0.102682f
C583 a_n3827_n3924.n21 gnd 0.838616f
C584 a_n3827_n3924.n22 gnd 0.340114f
C585 a_n3827_n3924.t57 gnd 0.102682f
C586 a_n3827_n3924.t46 gnd 0.102682f
C587 a_n3827_n3924.n23 gnd 0.838616f
C588 a_n3827_n3924.n24 gnd 0.340114f
C589 a_n3827_n3924.t5 gnd 1.06718f
C590 a_n3827_n3924.n25 gnd 0.920947f
C591 a_n3827_n3924.t55 gnd 1.06718f
C592 a_n3827_n3924.n26 gnd 0.58539f
C593 a_n3827_n3924.t40 gnd 0.102682f
C594 a_n3827_n3924.t2 gnd 0.102682f
C595 a_n3827_n3924.n27 gnd 0.838615f
C596 a_n3827_n3924.n28 gnd 0.340116f
C597 a_n3827_n3924.t33 gnd 0.102682f
C598 a_n3827_n3924.t3 gnd 0.102682f
C599 a_n3827_n3924.n29 gnd 0.838615f
C600 a_n3827_n3924.n30 gnd 0.340116f
C601 a_n3827_n3924.t1 gnd 0.102682f
C602 a_n3827_n3924.t4 gnd 0.102682f
C603 a_n3827_n3924.n31 gnd 0.838615f
C604 a_n3827_n3924.n32 gnd 0.340116f
C605 a_n3827_n3924.t9 gnd 0.102682f
C606 a_n3827_n3924.t56 gnd 0.102682f
C607 a_n3827_n3924.n33 gnd 0.838615f
C608 a_n3827_n3924.n34 gnd 0.340116f
C609 a_n3827_n3924.t47 gnd 0.102682f
C610 a_n3827_n3924.t23 gnd 0.102682f
C611 a_n3827_n3924.n35 gnd 0.838615f
C612 a_n3827_n3924.n36 gnd 0.340116f
C613 a_n3827_n3924.t41 gnd 1.06718f
C614 a_n3827_n3924.n37 gnd 0.362198f
C615 a_n3827_n3924.t36 gnd 1.06718f
C616 a_n3827_n3924.n38 gnd 0.362198f
C617 a_n3827_n3924.t25 gnd 0.102682f
C618 a_n3827_n3924.t10 gnd 0.102682f
C619 a_n3827_n3924.n39 gnd 0.838615f
C620 a_n3827_n3924.n40 gnd 0.340116f
C621 a_n3827_n3924.t53 gnd 0.102682f
C622 a_n3827_n3924.t49 gnd 0.102682f
C623 a_n3827_n3924.n41 gnd 0.838615f
C624 a_n3827_n3924.n42 gnd 0.340116f
C625 a_n3827_n3924.t22 gnd 0.102682f
C626 a_n3827_n3924.t27 gnd 0.102682f
C627 a_n3827_n3924.n43 gnd 0.838615f
C628 a_n3827_n3924.n44 gnd 0.340116f
C629 a_n3827_n3924.t7 gnd 0.102682f
C630 a_n3827_n3924.t35 gnd 0.102682f
C631 a_n3827_n3924.n45 gnd 0.838615f
C632 a_n3827_n3924.n46 gnd 0.340116f
C633 a_n3827_n3924.t34 gnd 0.102682f
C634 a_n3827_n3924.t50 gnd 0.102682f
C635 a_n3827_n3924.n47 gnd 0.838615f
C636 a_n3827_n3924.n48 gnd 0.340116f
C637 a_n3827_n3924.t38 gnd 1.06718f
C638 a_n3827_n3924.n49 gnd 0.58539f
C639 a_n3827_n3924.n50 gnd 0.958536f
C640 a_n3827_n3924.t13 gnd 1.32959f
C641 a_n3827_n3924.t17 gnd 1.32595f
C642 a_n3827_n3924.n51 gnd 1.82937f
C643 a_n3827_n3924.n52 gnd 0.504753f
C644 a_n3827_n3924.t12 gnd 1.32595f
C645 a_n3827_n3924.n53 gnd 0.844057f
C646 a_n3827_n3924.t15 gnd 1.32595f
C647 a_n3827_n3924.n54 gnd 0.933892f
C648 a_n3827_n3924.t11 gnd 1.32595f
C649 a_n3827_n3924.n55 gnd 0.933892f
C650 a_n3827_n3924.t16 gnd 1.32595f
C651 a_n3827_n3924.n56 gnd 0.933892f
C652 a_n3827_n3924.t19 gnd 1.32595f
C653 a_n3827_n3924.n57 gnd 0.918983f
C654 a_n3827_n3924.t18 gnd 1.32595f
C655 a_n3827_n3924.t14 gnd 1.32595f
C656 a_n3827_n3924.n58 gnd 1.5379f
C657 a_n3827_n3924.t20 gnd 1.32785f
C658 diffpairibias.t27 gnd 0.090128f
C659 diffpairibias.t23 gnd 0.08996f
C660 diffpairibias.n0 gnd 0.105991f
C661 diffpairibias.t28 gnd 0.08996f
C662 diffpairibias.n1 gnd 0.051736f
C663 diffpairibias.t25 gnd 0.08996f
C664 diffpairibias.n2 gnd 0.051736f
C665 diffpairibias.t29 gnd 0.08996f
C666 diffpairibias.n3 gnd 0.041084f
C667 diffpairibias.t15 gnd 0.086371f
C668 diffpairibias.t1 gnd 0.085993f
C669 diffpairibias.n4 gnd 0.13579f
C670 diffpairibias.t11 gnd 0.085993f
C671 diffpairibias.n5 gnd 0.072463f
C672 diffpairibias.t13 gnd 0.085993f
C673 diffpairibias.n6 gnd 0.072463f
C674 diffpairibias.t7 gnd 0.085993f
C675 diffpairibias.n7 gnd 0.072463f
C676 diffpairibias.t3 gnd 0.085993f
C677 diffpairibias.n8 gnd 0.072463f
C678 diffpairibias.t17 gnd 0.085993f
C679 diffpairibias.n9 gnd 0.072463f
C680 diffpairibias.t5 gnd 0.085993f
C681 diffpairibias.n10 gnd 0.072463f
C682 diffpairibias.t19 gnd 0.085993f
C683 diffpairibias.n11 gnd 0.072463f
C684 diffpairibias.t9 gnd 0.085993f
C685 diffpairibias.n12 gnd 0.102883f
C686 diffpairibias.t14 gnd 0.086899f
C687 diffpairibias.t0 gnd 0.086748f
C688 diffpairibias.n13 gnd 0.094648f
C689 diffpairibias.t10 gnd 0.086748f
C690 diffpairibias.n14 gnd 0.052262f
C691 diffpairibias.t12 gnd 0.086748f
C692 diffpairibias.n15 gnd 0.052262f
C693 diffpairibias.t6 gnd 0.086748f
C694 diffpairibias.n16 gnd 0.052262f
C695 diffpairibias.t2 gnd 0.086748f
C696 diffpairibias.n17 gnd 0.052262f
C697 diffpairibias.t16 gnd 0.086748f
C698 diffpairibias.n18 gnd 0.052262f
C699 diffpairibias.t4 gnd 0.086748f
C700 diffpairibias.n19 gnd 0.052262f
C701 diffpairibias.t18 gnd 0.086748f
C702 diffpairibias.n20 gnd 0.052262f
C703 diffpairibias.t8 gnd 0.086748f
C704 diffpairibias.n21 gnd 0.061849f
C705 diffpairibias.n22 gnd 0.233513f
C706 diffpairibias.t20 gnd 0.08996f
C707 diffpairibias.n23 gnd 0.051747f
C708 diffpairibias.t26 gnd 0.08996f
C709 diffpairibias.n24 gnd 0.051736f
C710 diffpairibias.t22 gnd 0.08996f
C711 diffpairibias.n25 gnd 0.051736f
C712 diffpairibias.t21 gnd 0.08996f
C713 diffpairibias.n26 gnd 0.051736f
C714 diffpairibias.t24 gnd 0.08996f
C715 diffpairibias.n27 gnd 0.04729f
C716 diffpairibias.n28 gnd 0.047711f
C717 a_n1808_13878.t4 gnd 0.185683f
C718 a_n1808_13878.t0 gnd 0.185683f
C719 a_n1808_13878.t2 gnd 0.185683f
C720 a_n1808_13878.n0 gnd 1.46364f
C721 a_n1808_13878.t6 gnd 0.185683f
C722 a_n1808_13878.t1 gnd 0.185683f
C723 a_n1808_13878.n1 gnd 1.46209f
C724 a_n1808_13878.n2 gnd 2.04299f
C725 a_n1808_13878.t5 gnd 0.185683f
C726 a_n1808_13878.t9 gnd 0.185683f
C727 a_n1808_13878.n3 gnd 1.46451f
C728 a_n1808_13878.t10 gnd 0.185683f
C729 a_n1808_13878.t3 gnd 0.185683f
C730 a_n1808_13878.n4 gnd 1.46209f
C731 a_n1808_13878.n5 gnd 1.31424f
C732 a_n1808_13878.t7 gnd 0.185683f
C733 a_n1808_13878.t8 gnd 0.185683f
C734 a_n1808_13878.n6 gnd 1.46209f
C735 a_n1808_13878.n7 gnd 1.80499f
C736 a_n1808_13878.t13 gnd 1.73864f
C737 a_n1808_13878.t16 gnd 0.185683f
C738 a_n1808_13878.t17 gnd 0.185683f
C739 a_n1808_13878.n8 gnd 1.30795f
C740 a_n1808_13878.n9 gnd 1.46144f
C741 a_n1808_13878.t12 gnd 1.73518f
C742 a_n1808_13878.n10 gnd 0.735417f
C743 a_n1808_13878.t15 gnd 1.73518f
C744 a_n1808_13878.n11 gnd 0.735417f
C745 a_n1808_13878.t18 gnd 0.185683f
C746 a_n1808_13878.t19 gnd 0.185683f
C747 a_n1808_13878.n12 gnd 1.30795f
C748 a_n1808_13878.n13 gnd 0.742539f
C749 a_n1808_13878.t14 gnd 1.73518f
C750 a_n1808_13878.n14 gnd 1.73174f
C751 a_n1808_13878.n15 gnd 2.52099f
C752 a_n1808_13878.n16 gnd 3.70273f
C753 a_n1808_13878.n17 gnd 1.46209f
C754 a_n1808_13878.t11 gnd 0.185683f
C755 a_n1986_8322.t2 gnd 38.652897f
C756 a_n1986_8322.t0 gnd 28.1251f
C757 a_n1986_8322.t3 gnd 19.258501f
C758 a_n1986_8322.t1 gnd 38.652897f
C759 a_n1986_8322.t13 gnd 0.875352f
C760 a_n1986_8322.t21 gnd 0.093486f
C761 a_n1986_8322.t16 gnd 0.093486f
C762 a_n1986_8322.n0 gnd 0.658513f
C763 a_n1986_8322.n1 gnd 0.735791f
C764 a_n1986_8322.t19 gnd 0.093486f
C765 a_n1986_8322.t18 gnd 0.093486f
C766 a_n1986_8322.n2 gnd 0.658513f
C767 a_n1986_8322.n3 gnd 0.373846f
C768 a_n1986_8322.t12 gnd 0.873609f
C769 a_n1986_8322.n4 gnd 1.39826f
C770 a_n1986_8322.t6 gnd 0.875352f
C771 a_n1986_8322.t10 gnd 0.093486f
C772 a_n1986_8322.t9 gnd 0.093486f
C773 a_n1986_8322.n5 gnd 0.658513f
C774 a_n1986_8322.n6 gnd 0.735791f
C775 a_n1986_8322.t4 gnd 0.873609f
C776 a_n1986_8322.n7 gnd 0.37026f
C777 a_n1986_8322.t7 gnd 0.873609f
C778 a_n1986_8322.n8 gnd 0.37026f
C779 a_n1986_8322.t5 gnd 0.093486f
C780 a_n1986_8322.t11 gnd 0.093486f
C781 a_n1986_8322.n9 gnd 0.658513f
C782 a_n1986_8322.n10 gnd 0.373846f
C783 a_n1986_8322.t8 gnd 0.873609f
C784 a_n1986_8322.n11 gnd 0.871879f
C785 a_n1986_8322.n12 gnd 1.58991f
C786 a_n1986_8322.n13 gnd 3.44798f
C787 a_n1986_8322.t15 gnd 0.873609f
C788 a_n1986_8322.n14 gnd 0.766135f
C789 a_n1986_8322.t14 gnd 0.093486f
C790 a_n1986_8322.t23 gnd 0.093486f
C791 a_n1986_8322.n15 gnd 0.658513f
C792 a_n1986_8322.n16 gnd 0.373846f
C793 a_n1986_8322.t20 gnd 0.093486f
C794 a_n1986_8322.t17 gnd 0.093486f
C795 a_n1986_8322.n17 gnd 0.658513f
C796 a_n1986_8322.n18 gnd 0.735789f
C797 a_n1986_8322.t22 gnd 0.875354f
C798 a_n1986_13878.n0 gnd 0.543543f
C799 a_n1986_13878.n1 gnd 0.211712f
C800 a_n1986_13878.n2 gnd 0.15593f
C801 a_n1986_13878.n3 gnd 0.245072f
C802 a_n1986_13878.n4 gnd 0.18929f
C803 a_n1986_13878.n5 gnd 0.211712f
C804 a_n1986_13878.n6 gnd 0.15593f
C805 a_n1986_13878.n7 gnd 0.599325f
C806 a_n1986_13878.n8 gnd 0.446674f
C807 a_n1986_13878.n9 gnd 0.223128f
C808 a_n1986_13878.n10 gnd 0.50886f
C809 a_n1986_13878.n11 gnd 0.291913f
C810 a_n1986_13878.n12 gnd 0.453077f
C811 a_n1986_13878.n13 gnd 0.223128f
C812 a_n1986_13878.n14 gnd 0.755878f
C813 a_n1986_13878.n15 gnd 0.291913f
C814 a_n1986_13878.n16 gnd 0.66047f
C815 a_n1986_13878.n17 gnd 0.291913f
C816 a_n1986_13878.n18 gnd 0.50886f
C817 a_n1986_13878.n19 gnd 0.686545f
C818 a_n1986_13878.n20 gnd 0.223128f
C819 a_n1986_13878.n21 gnd 0.291913f
C820 a_n1986_13878.n22 gnd 3.60937f
C821 a_n1986_13878.n23 gnd 2.74915f
C822 a_n1986_13878.n24 gnd 3.87242f
C823 a_n1986_13878.n25 gnd 1.83699f
C824 a_n1986_13878.n26 gnd 1.97943f
C825 a_n1986_13878.n27 gnd 0.751202f
C826 a_n1986_13878.n28 gnd 0.751204f
C827 a_n1986_13878.n29 gnd 3.32125f
C828 a_n1986_13878.n30 gnd 0.008639f
C829 a_n1986_13878.n32 gnd 1.38299f
C830 a_n1986_13878.n33 gnd 0.295172f
C831 a_n1986_13878.n34 gnd 0.111564f
C832 a_n1986_13878.n35 gnd 0.008639f
C833 a_n1986_13878.n37 gnd 0.008639f
C834 a_n1986_13878.n39 gnd 0.295172f
C835 a_n1986_13878.n40 gnd 0.008639f
C836 a_n1986_13878.n42 gnd 0.295172f
C837 a_n1986_13878.n43 gnd 0.008639f
C838 a_n1986_13878.n44 gnd 0.294752f
C839 a_n1986_13878.n45 gnd 0.008639f
C840 a_n1986_13878.n46 gnd 0.294752f
C841 a_n1986_13878.n47 gnd 0.008639f
C842 a_n1986_13878.n48 gnd 0.294752f
C843 a_n1986_13878.n49 gnd 0.008639f
C844 a_n1986_13878.n50 gnd 0.294752f
C845 a_n1986_13878.n51 gnd 0.295172f
C846 a_n1986_13878.t27 gnd 0.719888f
C847 a_n1986_13878.n52 gnd 0.316509f
C848 a_n1986_13878.t33 gnd 0.719888f
C849 a_n1986_13878.t15 gnd 0.719888f
C850 a_n1986_13878.t56 gnd 0.719888f
C851 a_n1986_13878.n53 gnd 0.316509f
C852 a_n1986_13878.t65 gnd 0.719888f
C853 a_n1986_13878.t71 gnd 0.719888f
C854 a_n1986_13878.t23 gnd 0.73505f
C855 a_n1986_13878.t21 gnd 0.719888f
C856 a_n1986_13878.t25 gnd 0.719888f
C857 a_n1986_13878.t19 gnd 0.719888f
C858 a_n1986_13878.n54 gnd 0.316509f
C859 a_n1986_13878.t17 gnd 0.719888f
C860 a_n1986_13878.t31 gnd 0.731791f
C861 a_n1986_13878.t39 gnd 0.120372f
C862 a_n1986_13878.t6 gnd 0.120372f
C863 a_n1986_13878.n55 gnd 1.06535f
C864 a_n1986_13878.t2 gnd 0.120372f
C865 a_n1986_13878.t46 gnd 0.120372f
C866 a_n1986_13878.n56 gnd 1.06365f
C867 a_n1986_13878.t42 gnd 0.120372f
C868 a_n1986_13878.t4 gnd 0.120372f
C869 a_n1986_13878.n57 gnd 1.06365f
C870 a_n1986_13878.t43 gnd 0.120372f
C871 a_n1986_13878.t41 gnd 0.120372f
C872 a_n1986_13878.n58 gnd 1.06535f
C873 a_n1986_13878.t38 gnd 0.120372f
C874 a_n1986_13878.t37 gnd 0.120372f
C875 a_n1986_13878.n59 gnd 1.06365f
C876 a_n1986_13878.t8 gnd 0.120372f
C877 a_n1986_13878.t0 gnd 0.120372f
C878 a_n1986_13878.n60 gnd 1.06365f
C879 a_n1986_13878.t12 gnd 0.120372f
C880 a_n1986_13878.t7 gnd 0.120372f
C881 a_n1986_13878.n61 gnd 1.06365f
C882 a_n1986_13878.t45 gnd 0.120372f
C883 a_n1986_13878.t9 gnd 0.120372f
C884 a_n1986_13878.n62 gnd 1.06365f
C885 a_n1986_13878.t11 gnd 0.120372f
C886 a_n1986_13878.t10 gnd 0.120372f
C887 a_n1986_13878.n63 gnd 1.06365f
C888 a_n1986_13878.t47 gnd 0.120372f
C889 a_n1986_13878.t3 gnd 0.120372f
C890 a_n1986_13878.n64 gnd 1.06535f
C891 a_n1986_13878.t44 gnd 0.120372f
C892 a_n1986_13878.t5 gnd 0.120372f
C893 a_n1986_13878.n65 gnd 1.06365f
C894 a_n1986_13878.t40 gnd 0.120372f
C895 a_n1986_13878.t1 gnd 0.120372f
C896 a_n1986_13878.n66 gnd 1.06365f
C897 a_n1986_13878.t75 gnd 0.73505f
C898 a_n1986_13878.t58 gnd 0.719888f
C899 a_n1986_13878.t62 gnd 0.719888f
C900 a_n1986_13878.t52 gnd 0.719888f
C901 a_n1986_13878.n67 gnd 0.316509f
C902 a_n1986_13878.t67 gnd 0.719888f
C903 a_n1986_13878.t73 gnd 0.731791f
C904 a_n1986_13878.n68 gnd 0.319213f
C905 a_n1986_13878.n69 gnd 0.312489f
C906 a_n1986_13878.n70 gnd 0.319212f
C907 a_n1986_13878.n71 gnd 0.319213f
C908 a_n1986_13878.n72 gnd 0.312489f
C909 a_n1986_13878.n73 gnd 0.319212f
C910 a_n1986_13878.t32 gnd 1.44913f
C911 a_n1986_13878.t20 gnd 0.154764f
C912 a_n1986_13878.t18 gnd 0.154764f
C913 a_n1986_13878.n74 gnd 1.09016f
C914 a_n1986_13878.t22 gnd 0.154764f
C915 a_n1986_13878.t26 gnd 0.154764f
C916 a_n1986_13878.n75 gnd 1.09016f
C917 a_n1986_13878.t24 gnd 1.44625f
C918 a_n1986_13878.n76 gnd 1.18267f
C919 a_n1986_13878.n77 gnd 0.813122f
C920 a_n1986_13878.t57 gnd 0.719888f
C921 a_n1986_13878.t66 gnd 0.719888f
C922 a_n1986_13878.t48 gnd 0.719888f
C923 a_n1986_13878.n78 gnd 0.316509f
C924 a_n1986_13878.t68 gnd 0.719888f
C925 a_n1986_13878.t53 gnd 0.719888f
C926 a_n1986_13878.t54 gnd 0.719888f
C927 a_n1986_13878.n79 gnd 0.316509f
C928 a_n1986_13878.t72 gnd 0.719888f
C929 a_n1986_13878.t61 gnd 0.719888f
C930 a_n1986_13878.t60 gnd 0.719888f
C931 a_n1986_13878.n80 gnd 0.316509f
C932 a_n1986_13878.t64 gnd 0.719888f
C933 a_n1986_13878.t55 gnd 0.719888f
C934 a_n1986_13878.t49 gnd 0.719888f
C935 a_n1986_13878.n81 gnd 0.316509f
C936 a_n1986_13878.t69 gnd 0.731951f
C937 a_n1986_13878.n82 gnd 0.312489f
C938 a_n1986_13878.n83 gnd 0.306815f
C939 a_n1986_13878.t74 gnd 0.731951f
C940 a_n1986_13878.n84 gnd 0.312489f
C941 a_n1986_13878.n85 gnd 0.306815f
C942 a_n1986_13878.t63 gnd 0.731951f
C943 a_n1986_13878.n86 gnd 0.312489f
C944 a_n1986_13878.n87 gnd 0.306815f
C945 a_n1986_13878.t59 gnd 0.731951f
C946 a_n1986_13878.n88 gnd 0.312489f
C947 a_n1986_13878.n89 gnd 0.306815f
C948 a_n1986_13878.n90 gnd 1.03979f
C949 a_n1986_13878.t70 gnd 0.73505f
C950 a_n1986_13878.n91 gnd 0.319212f
C951 a_n1986_13878.t50 gnd 0.719888f
C952 a_n1986_13878.n92 gnd 0.312489f
C953 a_n1986_13878.n93 gnd 0.319213f
C954 a_n1986_13878.t51 gnd 0.731791f
C955 a_n1986_13878.t13 gnd 0.73505f
C956 a_n1986_13878.n94 gnd 0.319212f
C957 a_n1986_13878.t29 gnd 0.719888f
C958 a_n1986_13878.n95 gnd 0.312489f
C959 a_n1986_13878.n96 gnd 0.319213f
C960 a_n1986_13878.t35 gnd 0.731791f
C961 a_n1986_13878.n97 gnd 1.16971f
C962 a_n1986_13878.t36 gnd 1.44624f
C963 a_n1986_13878.t28 gnd 0.154764f
C964 a_n1986_13878.t34 gnd 0.154764f
C965 a_n1986_13878.n98 gnd 1.09016f
C966 a_n1986_13878.t16 gnd 0.154764f
C967 a_n1986_13878.t30 gnd 0.154764f
C968 a_n1986_13878.n99 gnd 1.09016f
C969 a_n1986_13878.n100 gnd 1.21809f
C970 a_n1986_13878.t14 gnd 1.44913f
C971 vdd.t22 gnd 0.032948f
C972 vdd.t186 gnd 0.032948f
C973 vdd.n0 gnd 0.259864f
C974 vdd.t26 gnd 0.032948f
C975 vdd.t199 gnd 0.032948f
C976 vdd.n1 gnd 0.259435f
C977 vdd.n2 gnd 0.239248f
C978 vdd.t182 gnd 0.032948f
C979 vdd.t189 gnd 0.032948f
C980 vdd.n3 gnd 0.259435f
C981 vdd.n4 gnd 0.120997f
C982 vdd.t17 gnd 0.032948f
C983 vdd.t37 gnd 0.032948f
C984 vdd.n5 gnd 0.259435f
C985 vdd.n6 gnd 0.113533f
C986 vdd.t28 gnd 0.032948f
C987 vdd.t184 gnd 0.032948f
C988 vdd.n7 gnd 0.259864f
C989 vdd.t195 gnd 0.032948f
C990 vdd.t19 gnd 0.032948f
C991 vdd.n8 gnd 0.259435f
C992 vdd.n9 gnd 0.239248f
C993 vdd.t191 gnd 0.032948f
C994 vdd.t32 gnd 0.032948f
C995 vdd.n10 gnd 0.259435f
C996 vdd.n11 gnd 0.120997f
C997 vdd.t39 gnd 0.032948f
C998 vdd.t193 gnd 0.032948f
C999 vdd.n12 gnd 0.259435f
C1000 vdd.n13 gnd 0.113533f
C1001 vdd.n14 gnd 0.080266f
C1002 vdd.t5 gnd 0.018304f
C1003 vdd.t9 gnd 0.018304f
C1004 vdd.n15 gnd 0.168483f
C1005 vdd.t7 gnd 0.018304f
C1006 vdd.t10 gnd 0.018304f
C1007 vdd.n16 gnd 0.16799f
C1008 vdd.n17 gnd 0.292355f
C1009 vdd.t14 gnd 0.018304f
C1010 vdd.t0 gnd 0.018304f
C1011 vdd.n18 gnd 0.16799f
C1012 vdd.n19 gnd 0.120951f
C1013 vdd.t12 gnd 0.018304f
C1014 vdd.t1 gnd 0.018304f
C1015 vdd.n20 gnd 0.168483f
C1016 vdd.t4 gnd 0.018304f
C1017 vdd.t2 gnd 0.018304f
C1018 vdd.n21 gnd 0.16799f
C1019 vdd.n22 gnd 0.292355f
C1020 vdd.t13 gnd 0.018304f
C1021 vdd.t6 gnd 0.018304f
C1022 vdd.n23 gnd 0.16799f
C1023 vdd.n24 gnd 0.120951f
C1024 vdd.t8 gnd 0.018304f
C1025 vdd.t15 gnd 0.018304f
C1026 vdd.n25 gnd 0.16799f
C1027 vdd.t3 gnd 0.018304f
C1028 vdd.t11 gnd 0.018304f
C1029 vdd.n26 gnd 0.16799f
C1030 vdd.n27 gnd 18.392f
C1031 vdd.n28 gnd 6.85872f
C1032 vdd.n29 gnd 0.004992f
C1033 vdd.n30 gnd 0.004633f
C1034 vdd.n31 gnd 0.002563f
C1035 vdd.n32 gnd 0.005884f
C1036 vdd.n33 gnd 0.002489f
C1037 vdd.n34 gnd 0.002636f
C1038 vdd.n35 gnd 0.004633f
C1039 vdd.n36 gnd 0.002489f
C1040 vdd.n37 gnd 0.005884f
C1041 vdd.n38 gnd 0.002636f
C1042 vdd.n39 gnd 0.004633f
C1043 vdd.n40 gnd 0.002489f
C1044 vdd.n41 gnd 0.004413f
C1045 vdd.n42 gnd 0.004426f
C1046 vdd.t120 gnd 0.012641f
C1047 vdd.n43 gnd 0.028127f
C1048 vdd.n44 gnd 0.146377f
C1049 vdd.n45 gnd 0.002489f
C1050 vdd.n46 gnd 0.002636f
C1051 vdd.n47 gnd 0.005884f
C1052 vdd.n48 gnd 0.005884f
C1053 vdd.n49 gnd 0.002636f
C1054 vdd.n50 gnd 0.002489f
C1055 vdd.n51 gnd 0.004633f
C1056 vdd.n52 gnd 0.004633f
C1057 vdd.n53 gnd 0.002489f
C1058 vdd.n54 gnd 0.002636f
C1059 vdd.n55 gnd 0.005884f
C1060 vdd.n56 gnd 0.005884f
C1061 vdd.n57 gnd 0.002636f
C1062 vdd.n58 gnd 0.002489f
C1063 vdd.n59 gnd 0.004633f
C1064 vdd.n60 gnd 0.004633f
C1065 vdd.n61 gnd 0.002489f
C1066 vdd.n62 gnd 0.002636f
C1067 vdd.n63 gnd 0.005884f
C1068 vdd.n64 gnd 0.005884f
C1069 vdd.n65 gnd 0.013911f
C1070 vdd.n66 gnd 0.002563f
C1071 vdd.n67 gnd 0.002489f
C1072 vdd.n68 gnd 0.011974f
C1073 vdd.n69 gnd 0.008359f
C1074 vdd.t172 gnd 0.029287f
C1075 vdd.t146 gnd 0.029287f
C1076 vdd.n70 gnd 0.201279f
C1077 vdd.n71 gnd 0.158275f
C1078 vdd.t179 gnd 0.029287f
C1079 vdd.t135 gnd 0.029287f
C1080 vdd.n72 gnd 0.201279f
C1081 vdd.n73 gnd 0.127727f
C1082 vdd.t165 gnd 0.029287f
C1083 vdd.t140 gnd 0.029287f
C1084 vdd.n74 gnd 0.201279f
C1085 vdd.n75 gnd 0.127727f
C1086 vdd.n76 gnd 0.004992f
C1087 vdd.n77 gnd 0.004633f
C1088 vdd.n78 gnd 0.002563f
C1089 vdd.n79 gnd 0.005884f
C1090 vdd.n80 gnd 0.002489f
C1091 vdd.n81 gnd 0.002636f
C1092 vdd.n82 gnd 0.004633f
C1093 vdd.n83 gnd 0.002489f
C1094 vdd.n84 gnd 0.005884f
C1095 vdd.n85 gnd 0.002636f
C1096 vdd.n86 gnd 0.004633f
C1097 vdd.n87 gnd 0.002489f
C1098 vdd.n88 gnd 0.004413f
C1099 vdd.n89 gnd 0.004426f
C1100 vdd.t178 gnd 0.012641f
C1101 vdd.n90 gnd 0.028127f
C1102 vdd.n91 gnd 0.146377f
C1103 vdd.n92 gnd 0.002489f
C1104 vdd.n93 gnd 0.002636f
C1105 vdd.n94 gnd 0.005884f
C1106 vdd.n95 gnd 0.005884f
C1107 vdd.n96 gnd 0.002636f
C1108 vdd.n97 gnd 0.002489f
C1109 vdd.n98 gnd 0.004633f
C1110 vdd.n99 gnd 0.004633f
C1111 vdd.n100 gnd 0.002489f
C1112 vdd.n101 gnd 0.002636f
C1113 vdd.n102 gnd 0.005884f
C1114 vdd.n103 gnd 0.005884f
C1115 vdd.n104 gnd 0.002636f
C1116 vdd.n105 gnd 0.002489f
C1117 vdd.n106 gnd 0.004633f
C1118 vdd.n107 gnd 0.004633f
C1119 vdd.n108 gnd 0.002489f
C1120 vdd.n109 gnd 0.002636f
C1121 vdd.n110 gnd 0.005884f
C1122 vdd.n111 gnd 0.005884f
C1123 vdd.n112 gnd 0.013911f
C1124 vdd.n113 gnd 0.002563f
C1125 vdd.n114 gnd 0.002489f
C1126 vdd.n115 gnd 0.011974f
C1127 vdd.n116 gnd 0.008097f
C1128 vdd.n117 gnd 0.09503f
C1129 vdd.n118 gnd 0.004992f
C1130 vdd.n119 gnd 0.004633f
C1131 vdd.n120 gnd 0.002563f
C1132 vdd.n121 gnd 0.005884f
C1133 vdd.n122 gnd 0.002489f
C1134 vdd.n123 gnd 0.002636f
C1135 vdd.n124 gnd 0.004633f
C1136 vdd.n125 gnd 0.002489f
C1137 vdd.n126 gnd 0.005884f
C1138 vdd.n127 gnd 0.002636f
C1139 vdd.n128 gnd 0.004633f
C1140 vdd.n129 gnd 0.002489f
C1141 vdd.n130 gnd 0.004413f
C1142 vdd.n131 gnd 0.004426f
C1143 vdd.t147 gnd 0.012641f
C1144 vdd.n132 gnd 0.028127f
C1145 vdd.n133 gnd 0.146377f
C1146 vdd.n134 gnd 0.002489f
C1147 vdd.n135 gnd 0.002636f
C1148 vdd.n136 gnd 0.005884f
C1149 vdd.n137 gnd 0.005884f
C1150 vdd.n138 gnd 0.002636f
C1151 vdd.n139 gnd 0.002489f
C1152 vdd.n140 gnd 0.004633f
C1153 vdd.n141 gnd 0.004633f
C1154 vdd.n142 gnd 0.002489f
C1155 vdd.n143 gnd 0.002636f
C1156 vdd.n144 gnd 0.005884f
C1157 vdd.n145 gnd 0.005884f
C1158 vdd.n146 gnd 0.002636f
C1159 vdd.n147 gnd 0.002489f
C1160 vdd.n148 gnd 0.004633f
C1161 vdd.n149 gnd 0.004633f
C1162 vdd.n150 gnd 0.002489f
C1163 vdd.n151 gnd 0.002636f
C1164 vdd.n152 gnd 0.005884f
C1165 vdd.n153 gnd 0.005884f
C1166 vdd.n154 gnd 0.013911f
C1167 vdd.n155 gnd 0.002563f
C1168 vdd.n156 gnd 0.002489f
C1169 vdd.n157 gnd 0.011974f
C1170 vdd.n158 gnd 0.008359f
C1171 vdd.t149 gnd 0.029287f
C1172 vdd.t160 gnd 0.029287f
C1173 vdd.n159 gnd 0.201279f
C1174 vdd.n160 gnd 0.158275f
C1175 vdd.t124 gnd 0.029287f
C1176 vdd.t143 gnd 0.029287f
C1177 vdd.n161 gnd 0.201279f
C1178 vdd.n162 gnd 0.127727f
C1179 vdd.t159 gnd 0.029287f
C1180 vdd.t180 gnd 0.029287f
C1181 vdd.n163 gnd 0.201279f
C1182 vdd.n164 gnd 0.127727f
C1183 vdd.n165 gnd 0.004992f
C1184 vdd.n166 gnd 0.004633f
C1185 vdd.n167 gnd 0.002563f
C1186 vdd.n168 gnd 0.005884f
C1187 vdd.n169 gnd 0.002489f
C1188 vdd.n170 gnd 0.002636f
C1189 vdd.n171 gnd 0.004633f
C1190 vdd.n172 gnd 0.002489f
C1191 vdd.n173 gnd 0.005884f
C1192 vdd.n174 gnd 0.002636f
C1193 vdd.n175 gnd 0.004633f
C1194 vdd.n176 gnd 0.002489f
C1195 vdd.n177 gnd 0.004413f
C1196 vdd.n178 gnd 0.004426f
C1197 vdd.t137 gnd 0.012641f
C1198 vdd.n179 gnd 0.028127f
C1199 vdd.n180 gnd 0.146377f
C1200 vdd.n181 gnd 0.002489f
C1201 vdd.n182 gnd 0.002636f
C1202 vdd.n183 gnd 0.005884f
C1203 vdd.n184 gnd 0.005884f
C1204 vdd.n185 gnd 0.002636f
C1205 vdd.n186 gnd 0.002489f
C1206 vdd.n187 gnd 0.004633f
C1207 vdd.n188 gnd 0.004633f
C1208 vdd.n189 gnd 0.002489f
C1209 vdd.n190 gnd 0.002636f
C1210 vdd.n191 gnd 0.005884f
C1211 vdd.n192 gnd 0.005884f
C1212 vdd.n193 gnd 0.002636f
C1213 vdd.n194 gnd 0.002489f
C1214 vdd.n195 gnd 0.004633f
C1215 vdd.n196 gnd 0.004633f
C1216 vdd.n197 gnd 0.002489f
C1217 vdd.n198 gnd 0.002636f
C1218 vdd.n199 gnd 0.005884f
C1219 vdd.n200 gnd 0.005884f
C1220 vdd.n201 gnd 0.013911f
C1221 vdd.n202 gnd 0.002563f
C1222 vdd.n203 gnd 0.002489f
C1223 vdd.n204 gnd 0.011974f
C1224 vdd.n205 gnd 0.008097f
C1225 vdd.n206 gnd 0.056533f
C1226 vdd.n207 gnd 0.203704f
C1227 vdd.n208 gnd 0.004992f
C1228 vdd.n209 gnd 0.004633f
C1229 vdd.n210 gnd 0.002563f
C1230 vdd.n211 gnd 0.005884f
C1231 vdd.n212 gnd 0.002489f
C1232 vdd.n213 gnd 0.002636f
C1233 vdd.n214 gnd 0.004633f
C1234 vdd.n215 gnd 0.002489f
C1235 vdd.n216 gnd 0.005884f
C1236 vdd.n217 gnd 0.002636f
C1237 vdd.n218 gnd 0.004633f
C1238 vdd.n219 gnd 0.002489f
C1239 vdd.n220 gnd 0.004413f
C1240 vdd.n221 gnd 0.004426f
C1241 vdd.t152 gnd 0.012641f
C1242 vdd.n222 gnd 0.028127f
C1243 vdd.n223 gnd 0.146377f
C1244 vdd.n224 gnd 0.002489f
C1245 vdd.n225 gnd 0.002636f
C1246 vdd.n226 gnd 0.005884f
C1247 vdd.n227 gnd 0.005884f
C1248 vdd.n228 gnd 0.002636f
C1249 vdd.n229 gnd 0.002489f
C1250 vdd.n230 gnd 0.004633f
C1251 vdd.n231 gnd 0.004633f
C1252 vdd.n232 gnd 0.002489f
C1253 vdd.n233 gnd 0.002636f
C1254 vdd.n234 gnd 0.005884f
C1255 vdd.n235 gnd 0.005884f
C1256 vdd.n236 gnd 0.002636f
C1257 vdd.n237 gnd 0.002489f
C1258 vdd.n238 gnd 0.004633f
C1259 vdd.n239 gnd 0.004633f
C1260 vdd.n240 gnd 0.002489f
C1261 vdd.n241 gnd 0.002636f
C1262 vdd.n242 gnd 0.005884f
C1263 vdd.n243 gnd 0.005884f
C1264 vdd.n244 gnd 0.013911f
C1265 vdd.n245 gnd 0.002563f
C1266 vdd.n246 gnd 0.002489f
C1267 vdd.n247 gnd 0.011974f
C1268 vdd.n248 gnd 0.008359f
C1269 vdd.t153 gnd 0.029287f
C1270 vdd.t169 gnd 0.029287f
C1271 vdd.n249 gnd 0.201279f
C1272 vdd.n250 gnd 0.158275f
C1273 vdd.t130 gnd 0.029287f
C1274 vdd.t151 gnd 0.029287f
C1275 vdd.n251 gnd 0.201279f
C1276 vdd.n252 gnd 0.127727f
C1277 vdd.t164 gnd 0.029287f
C1278 vdd.t128 gnd 0.029287f
C1279 vdd.n253 gnd 0.201279f
C1280 vdd.n254 gnd 0.127727f
C1281 vdd.n255 gnd 0.004992f
C1282 vdd.n256 gnd 0.004633f
C1283 vdd.n257 gnd 0.002563f
C1284 vdd.n258 gnd 0.005884f
C1285 vdd.n259 gnd 0.002489f
C1286 vdd.n260 gnd 0.002636f
C1287 vdd.n261 gnd 0.004633f
C1288 vdd.n262 gnd 0.002489f
C1289 vdd.n263 gnd 0.005884f
C1290 vdd.n264 gnd 0.002636f
C1291 vdd.n265 gnd 0.004633f
C1292 vdd.n266 gnd 0.002489f
C1293 vdd.n267 gnd 0.004413f
C1294 vdd.n268 gnd 0.004426f
C1295 vdd.t141 gnd 0.012641f
C1296 vdd.n269 gnd 0.028127f
C1297 vdd.n270 gnd 0.146377f
C1298 vdd.n271 gnd 0.002489f
C1299 vdd.n272 gnd 0.002636f
C1300 vdd.n273 gnd 0.005884f
C1301 vdd.n274 gnd 0.005884f
C1302 vdd.n275 gnd 0.002636f
C1303 vdd.n276 gnd 0.002489f
C1304 vdd.n277 gnd 0.004633f
C1305 vdd.n278 gnd 0.004633f
C1306 vdd.n279 gnd 0.002489f
C1307 vdd.n280 gnd 0.002636f
C1308 vdd.n281 gnd 0.005884f
C1309 vdd.n282 gnd 0.005884f
C1310 vdd.n283 gnd 0.002636f
C1311 vdd.n284 gnd 0.002489f
C1312 vdd.n285 gnd 0.004633f
C1313 vdd.n286 gnd 0.004633f
C1314 vdd.n287 gnd 0.002489f
C1315 vdd.n288 gnd 0.002636f
C1316 vdd.n289 gnd 0.005884f
C1317 vdd.n290 gnd 0.005884f
C1318 vdd.n291 gnd 0.013911f
C1319 vdd.n292 gnd 0.002563f
C1320 vdd.n293 gnd 0.002489f
C1321 vdd.n294 gnd 0.011974f
C1322 vdd.n295 gnd 0.008097f
C1323 vdd.n296 gnd 0.056533f
C1324 vdd.n297 gnd 0.220485f
C1325 vdd.n298 gnd 0.006991f
C1326 vdd.n299 gnd 0.009097f
C1327 vdd.n300 gnd 0.007322f
C1328 vdd.n301 gnd 0.007322f
C1329 vdd.n302 gnd 0.009097f
C1330 vdd.n303 gnd 0.009097f
C1331 vdd.n304 gnd 0.664689f
C1332 vdd.n305 gnd 0.009097f
C1333 vdd.n306 gnd 0.009097f
C1334 vdd.n307 gnd 0.009097f
C1335 vdd.n308 gnd 0.720467f
C1336 vdd.n309 gnd 0.009097f
C1337 vdd.n310 gnd 0.009097f
C1338 vdd.n311 gnd 0.009097f
C1339 vdd.n312 gnd 0.009097f
C1340 vdd.n313 gnd 0.007322f
C1341 vdd.n314 gnd 0.009097f
C1342 vdd.t127 gnd 0.464817f
C1343 vdd.n315 gnd 0.009097f
C1344 vdd.n316 gnd 0.009097f
C1345 vdd.n317 gnd 0.009097f
C1346 vdd.n318 gnd 0.929634f
C1347 vdd.n319 gnd 0.009097f
C1348 vdd.n320 gnd 0.009097f
C1349 vdd.n321 gnd 0.009097f
C1350 vdd.n322 gnd 0.009097f
C1351 vdd.n323 gnd 0.009097f
C1352 vdd.n324 gnd 0.007322f
C1353 vdd.n325 gnd 0.009097f
C1354 vdd.n326 gnd 0.009097f
C1355 vdd.n327 gnd 0.009097f
C1356 vdd.n328 gnd 0.022169f
C1357 vdd.n329 gnd 2.22183f
C1358 vdd.n330 gnd 0.022678f
C1359 vdd.n331 gnd 0.009097f
C1360 vdd.n332 gnd 0.009097f
C1361 vdd.n334 gnd 0.009097f
C1362 vdd.n335 gnd 0.009097f
C1363 vdd.n336 gnd 0.007322f
C1364 vdd.n337 gnd 0.007322f
C1365 vdd.n338 gnd 0.009097f
C1366 vdd.n339 gnd 0.009097f
C1367 vdd.n340 gnd 0.009097f
C1368 vdd.n341 gnd 0.009097f
C1369 vdd.n342 gnd 0.009097f
C1370 vdd.n343 gnd 0.009097f
C1371 vdd.n344 gnd 0.007322f
C1372 vdd.n346 gnd 0.009097f
C1373 vdd.n347 gnd 0.009097f
C1374 vdd.n348 gnd 0.009097f
C1375 vdd.n349 gnd 0.009097f
C1376 vdd.n350 gnd 0.009097f
C1377 vdd.n351 gnd 0.007322f
C1378 vdd.n353 gnd 0.009097f
C1379 vdd.n354 gnd 0.009097f
C1380 vdd.n355 gnd 0.009097f
C1381 vdd.n356 gnd 0.009097f
C1382 vdd.n357 gnd 0.009097f
C1383 vdd.n358 gnd 0.007322f
C1384 vdd.n360 gnd 0.009097f
C1385 vdd.n361 gnd 0.009097f
C1386 vdd.n362 gnd 0.009097f
C1387 vdd.n363 gnd 0.009097f
C1388 vdd.n364 gnd 0.006114f
C1389 vdd.t72 gnd 0.111913f
C1390 vdd.t71 gnd 0.119604f
C1391 vdd.t70 gnd 0.146157f
C1392 vdd.n365 gnd 0.187352f
C1393 vdd.n366 gnd 0.158142f
C1394 vdd.n368 gnd 0.009097f
C1395 vdd.n369 gnd 0.009097f
C1396 vdd.n370 gnd 0.007322f
C1397 vdd.n371 gnd 0.009097f
C1398 vdd.n373 gnd 0.009097f
C1399 vdd.n374 gnd 0.009097f
C1400 vdd.n375 gnd 0.009097f
C1401 vdd.n376 gnd 0.009097f
C1402 vdd.n377 gnd 0.007322f
C1403 vdd.n379 gnd 0.009097f
C1404 vdd.n380 gnd 0.009097f
C1405 vdd.n381 gnd 0.009097f
C1406 vdd.n382 gnd 0.009097f
C1407 vdd.n383 gnd 0.009097f
C1408 vdd.n384 gnd 0.007322f
C1409 vdd.n386 gnd 0.009097f
C1410 vdd.n387 gnd 0.009097f
C1411 vdd.n388 gnd 0.009097f
C1412 vdd.n389 gnd 0.009097f
C1413 vdd.n390 gnd 0.009097f
C1414 vdd.n391 gnd 0.007322f
C1415 vdd.n393 gnd 0.009097f
C1416 vdd.n394 gnd 0.009097f
C1417 vdd.n395 gnd 0.009097f
C1418 vdd.n396 gnd 0.009097f
C1419 vdd.n397 gnd 0.009097f
C1420 vdd.n398 gnd 0.007322f
C1421 vdd.n400 gnd 0.009097f
C1422 vdd.n401 gnd 0.009097f
C1423 vdd.n402 gnd 0.009097f
C1424 vdd.n403 gnd 0.009097f
C1425 vdd.n404 gnd 0.007248f
C1426 vdd.t66 gnd 0.111913f
C1427 vdd.t65 gnd 0.119604f
C1428 vdd.t63 gnd 0.146157f
C1429 vdd.n405 gnd 0.187352f
C1430 vdd.n406 gnd 0.158142f
C1431 vdd.n408 gnd 0.009097f
C1432 vdd.n409 gnd 0.009097f
C1433 vdd.n410 gnd 0.007322f
C1434 vdd.n411 gnd 0.009097f
C1435 vdd.n413 gnd 0.009097f
C1436 vdd.n414 gnd 0.009097f
C1437 vdd.n415 gnd 0.009097f
C1438 vdd.n416 gnd 0.009097f
C1439 vdd.n417 gnd 0.007322f
C1440 vdd.n419 gnd 0.009097f
C1441 vdd.n420 gnd 0.009097f
C1442 vdd.n421 gnd 0.009097f
C1443 vdd.n422 gnd 0.009097f
C1444 vdd.n423 gnd 0.009097f
C1445 vdd.n424 gnd 0.007322f
C1446 vdd.n426 gnd 0.009097f
C1447 vdd.n427 gnd 0.009097f
C1448 vdd.n428 gnd 0.009097f
C1449 vdd.n429 gnd 0.009097f
C1450 vdd.n430 gnd 0.009097f
C1451 vdd.n431 gnd 0.007322f
C1452 vdd.n433 gnd 0.009097f
C1453 vdd.n434 gnd 0.009097f
C1454 vdd.n435 gnd 0.009097f
C1455 vdd.n436 gnd 0.009097f
C1456 vdd.n437 gnd 0.009097f
C1457 vdd.n438 gnd 0.007322f
C1458 vdd.n440 gnd 0.009097f
C1459 vdd.n441 gnd 0.009097f
C1460 vdd.n442 gnd 0.009097f
C1461 vdd.n443 gnd 0.009097f
C1462 vdd.n444 gnd 0.009097f
C1463 vdd.n445 gnd 0.009097f
C1464 vdd.n446 gnd 0.007322f
C1465 vdd.n447 gnd 0.009097f
C1466 vdd.n448 gnd 0.009097f
C1467 vdd.n449 gnd 0.007322f
C1468 vdd.n450 gnd 0.009097f
C1469 vdd.n451 gnd 0.007322f
C1470 vdd.n452 gnd 0.009097f
C1471 vdd.n453 gnd 0.007322f
C1472 vdd.n454 gnd 0.009097f
C1473 vdd.n455 gnd 0.009097f
C1474 vdd.n456 gnd 0.506651f
C1475 vdd.t123 gnd 0.464817f
C1476 vdd.n457 gnd 0.009097f
C1477 vdd.n458 gnd 0.007322f
C1478 vdd.n459 gnd 0.009097f
C1479 vdd.n460 gnd 0.007322f
C1480 vdd.n461 gnd 0.009097f
C1481 vdd.t148 gnd 0.464817f
C1482 vdd.n462 gnd 0.009097f
C1483 vdd.n463 gnd 0.007322f
C1484 vdd.n464 gnd 0.009097f
C1485 vdd.n465 gnd 0.007322f
C1486 vdd.n466 gnd 0.009097f
C1487 vdd.t119 gnd 0.464817f
C1488 vdd.n467 gnd 0.581022f
C1489 vdd.n468 gnd 0.009097f
C1490 vdd.n469 gnd 0.007322f
C1491 vdd.n470 gnd 0.009097f
C1492 vdd.n471 gnd 0.007322f
C1493 vdd.n472 gnd 0.009097f
C1494 vdd.n473 gnd 0.929634f
C1495 vdd.n474 gnd 0.009097f
C1496 vdd.n475 gnd 0.007322f
C1497 vdd.n476 gnd 0.022169f
C1498 vdd.n477 gnd 0.006077f
C1499 vdd.n478 gnd 0.022169f
C1500 vdd.t42 gnd 0.464817f
C1501 vdd.n479 gnd 0.022169f
C1502 vdd.n480 gnd 0.006077f
C1503 vdd.n481 gnd 0.007823f
C1504 vdd.n482 gnd 0.007322f
C1505 vdd.n483 gnd 0.009097f
C1506 vdd.n484 gnd 6.40518f
C1507 vdd.n515 gnd 0.022678f
C1508 vdd.n516 gnd 1.27825f
C1509 vdd.n517 gnd 0.009097f
C1510 vdd.n518 gnd 0.007322f
C1511 vdd.n519 gnd 0.005822f
C1512 vdd.n520 gnd 0.014864f
C1513 vdd.n521 gnd 0.007322f
C1514 vdd.n522 gnd 0.009097f
C1515 vdd.n523 gnd 0.009097f
C1516 vdd.n524 gnd 0.009097f
C1517 vdd.n525 gnd 0.009097f
C1518 vdd.n526 gnd 0.009097f
C1519 vdd.n527 gnd 0.009097f
C1520 vdd.n528 gnd 0.009097f
C1521 vdd.n529 gnd 0.009097f
C1522 vdd.n530 gnd 0.009097f
C1523 vdd.n531 gnd 0.009097f
C1524 vdd.n532 gnd 0.009097f
C1525 vdd.n533 gnd 0.009097f
C1526 vdd.n534 gnd 0.009097f
C1527 vdd.n535 gnd 0.009097f
C1528 vdd.n536 gnd 0.006114f
C1529 vdd.n537 gnd 0.009097f
C1530 vdd.n538 gnd 0.009097f
C1531 vdd.n539 gnd 0.009097f
C1532 vdd.n540 gnd 0.009097f
C1533 vdd.n541 gnd 0.009097f
C1534 vdd.n542 gnd 0.009097f
C1535 vdd.n543 gnd 0.009097f
C1536 vdd.n544 gnd 0.009097f
C1537 vdd.n545 gnd 0.009097f
C1538 vdd.n546 gnd 0.009097f
C1539 vdd.n547 gnd 0.009097f
C1540 vdd.n548 gnd 0.009097f
C1541 vdd.n549 gnd 0.009097f
C1542 vdd.n550 gnd 0.009097f
C1543 vdd.n551 gnd 0.009097f
C1544 vdd.n552 gnd 0.009097f
C1545 vdd.n553 gnd 0.009097f
C1546 vdd.n554 gnd 0.009097f
C1547 vdd.n555 gnd 0.009097f
C1548 vdd.n556 gnd 0.007248f
C1549 vdd.t43 gnd 0.111913f
C1550 vdd.t44 gnd 0.119604f
C1551 vdd.t41 gnd 0.146157f
C1552 vdd.n557 gnd 0.187352f
C1553 vdd.n558 gnd 0.15741f
C1554 vdd.n559 gnd 0.009097f
C1555 vdd.n560 gnd 0.009097f
C1556 vdd.n561 gnd 0.009097f
C1557 vdd.n562 gnd 0.009097f
C1558 vdd.n563 gnd 0.009097f
C1559 vdd.n564 gnd 0.009097f
C1560 vdd.n565 gnd 0.009097f
C1561 vdd.n566 gnd 0.009097f
C1562 vdd.n567 gnd 0.009097f
C1563 vdd.n568 gnd 0.009097f
C1564 vdd.n569 gnd 0.009097f
C1565 vdd.n570 gnd 0.009097f
C1566 vdd.n571 gnd 0.009097f
C1567 vdd.n572 gnd 0.005822f
C1568 vdd.n575 gnd 0.006186f
C1569 vdd.n576 gnd 0.006186f
C1570 vdd.n577 gnd 0.006186f
C1571 vdd.n578 gnd 0.006186f
C1572 vdd.n579 gnd 0.006186f
C1573 vdd.n580 gnd 0.006186f
C1574 vdd.n582 gnd 0.006186f
C1575 vdd.n583 gnd 0.006186f
C1576 vdd.n585 gnd 0.006186f
C1577 vdd.n586 gnd 0.004503f
C1578 vdd.n588 gnd 0.006186f
C1579 vdd.t87 gnd 0.249964f
C1580 vdd.t86 gnd 0.255869f
C1581 vdd.t85 gnd 0.163186f
C1582 vdd.n589 gnd 0.088193f
C1583 vdd.n590 gnd 0.050026f
C1584 vdd.n591 gnd 0.00884f
C1585 vdd.n592 gnd 0.014457f
C1586 vdd.n594 gnd 0.006186f
C1587 vdd.n595 gnd 0.632151f
C1588 vdd.n596 gnd 0.013704f
C1589 vdd.n597 gnd 0.013704f
C1590 vdd.n598 gnd 0.006186f
C1591 vdd.n599 gnd 0.014678f
C1592 vdd.n600 gnd 0.006186f
C1593 vdd.n601 gnd 0.006186f
C1594 vdd.n602 gnd 0.006186f
C1595 vdd.n603 gnd 0.006186f
C1596 vdd.n604 gnd 0.006186f
C1597 vdd.n606 gnd 0.006186f
C1598 vdd.n607 gnd 0.006186f
C1599 vdd.n609 gnd 0.006186f
C1600 vdd.n610 gnd 0.006186f
C1601 vdd.n612 gnd 0.006186f
C1602 vdd.n613 gnd 0.006186f
C1603 vdd.n615 gnd 0.006186f
C1604 vdd.n616 gnd 0.006186f
C1605 vdd.n618 gnd 0.006186f
C1606 vdd.n619 gnd 0.006186f
C1607 vdd.n621 gnd 0.006186f
C1608 vdd.t80 gnd 0.249964f
C1609 vdd.t79 gnd 0.255869f
C1610 vdd.t77 gnd 0.163186f
C1611 vdd.n622 gnd 0.088193f
C1612 vdd.n623 gnd 0.050026f
C1613 vdd.n624 gnd 0.006186f
C1614 vdd.n626 gnd 0.006186f
C1615 vdd.n627 gnd 0.006186f
C1616 vdd.t78 gnd 0.316076f
C1617 vdd.n628 gnd 0.006186f
C1618 vdd.n629 gnd 0.006186f
C1619 vdd.n630 gnd 0.006186f
C1620 vdd.n631 gnd 0.006186f
C1621 vdd.n632 gnd 0.006186f
C1622 vdd.n633 gnd 0.632151f
C1623 vdd.n634 gnd 0.006186f
C1624 vdd.n635 gnd 0.006186f
C1625 vdd.n636 gnd 0.553133f
C1626 vdd.n637 gnd 0.006186f
C1627 vdd.n638 gnd 0.006186f
C1628 vdd.n639 gnd 0.005458f
C1629 vdd.n640 gnd 0.006186f
C1630 vdd.n641 gnd 0.557781f
C1631 vdd.n642 gnd 0.006186f
C1632 vdd.n643 gnd 0.006186f
C1633 vdd.n644 gnd 0.006186f
C1634 vdd.n645 gnd 0.006186f
C1635 vdd.n646 gnd 0.006186f
C1636 vdd.n647 gnd 0.632151f
C1637 vdd.n648 gnd 0.006186f
C1638 vdd.n649 gnd 0.006186f
C1639 vdd.t57 gnd 0.283539f
C1640 vdd.t40 gnd 0.074371f
C1641 vdd.n650 gnd 0.006186f
C1642 vdd.n651 gnd 0.006186f
C1643 vdd.n652 gnd 0.006186f
C1644 vdd.t34 gnd 0.316076f
C1645 vdd.n653 gnd 0.006186f
C1646 vdd.n654 gnd 0.006186f
C1647 vdd.n655 gnd 0.006186f
C1648 vdd.n656 gnd 0.006186f
C1649 vdd.n657 gnd 0.006186f
C1650 vdd.t187 gnd 0.316076f
C1651 vdd.n658 gnd 0.006186f
C1652 vdd.n659 gnd 0.006186f
C1653 vdd.n660 gnd 0.525243f
C1654 vdd.n661 gnd 0.006186f
C1655 vdd.n662 gnd 0.006186f
C1656 vdd.n663 gnd 0.006186f
C1657 vdd.n664 gnd 0.385798f
C1658 vdd.n665 gnd 0.006186f
C1659 vdd.n666 gnd 0.006186f
C1660 vdd.t183 gnd 0.316076f
C1661 vdd.n667 gnd 0.006186f
C1662 vdd.n668 gnd 0.006186f
C1663 vdd.n669 gnd 0.006186f
C1664 vdd.n670 gnd 0.525243f
C1665 vdd.n671 gnd 0.006186f
C1666 vdd.n672 gnd 0.006186f
C1667 vdd.t35 gnd 0.269594f
C1668 vdd.t27 gnd 0.246353f
C1669 vdd.n673 gnd 0.006186f
C1670 vdd.n674 gnd 0.006186f
C1671 vdd.n675 gnd 0.006186f
C1672 vdd.t18 gnd 0.316076f
C1673 vdd.n676 gnd 0.006186f
C1674 vdd.n677 gnd 0.006186f
C1675 vdd.t197 gnd 0.316076f
C1676 vdd.n678 gnd 0.006186f
C1677 vdd.n679 gnd 0.006186f
C1678 vdd.n680 gnd 0.006186f
C1679 vdd.t33 gnd 0.232409f
C1680 vdd.n681 gnd 0.006186f
C1681 vdd.n682 gnd 0.006186f
C1682 vdd.n683 gnd 0.539188f
C1683 vdd.n684 gnd 0.006186f
C1684 vdd.n685 gnd 0.006186f
C1685 vdd.n686 gnd 0.006186f
C1686 vdd.n687 gnd 0.632151f
C1687 vdd.n688 gnd 0.006186f
C1688 vdd.n689 gnd 0.006186f
C1689 vdd.t194 gnd 0.283539f
C1690 vdd.n690 gnd 0.399743f
C1691 vdd.n691 gnd 0.006186f
C1692 vdd.n692 gnd 0.006186f
C1693 vdd.n693 gnd 0.006186f
C1694 vdd.t31 gnd 0.316076f
C1695 vdd.n694 gnd 0.006186f
C1696 vdd.n695 gnd 0.006186f
C1697 vdd.n696 gnd 0.006186f
C1698 vdd.n697 gnd 0.006186f
C1699 vdd.n698 gnd 0.006186f
C1700 vdd.t190 gnd 0.632151f
C1701 vdd.n699 gnd 0.006186f
C1702 vdd.n700 gnd 0.006186f
C1703 vdd.t82 gnd 0.316076f
C1704 vdd.n701 gnd 0.006186f
C1705 vdd.n702 gnd 0.014678f
C1706 vdd.n703 gnd 0.014678f
C1707 vdd.t192 gnd 0.594966f
C1708 vdd.n704 gnd 0.013704f
C1709 vdd.n705 gnd 0.013704f
C1710 vdd.n706 gnd 0.014678f
C1711 vdd.n707 gnd 0.006186f
C1712 vdd.n708 gnd 0.006186f
C1713 vdd.t16 gnd 0.594966f
C1714 vdd.n726 gnd 0.014678f
C1715 vdd.n744 gnd 0.013704f
C1716 vdd.n745 gnd 0.006186f
C1717 vdd.n746 gnd 0.013704f
C1718 vdd.t107 gnd 0.249964f
C1719 vdd.t106 gnd 0.255869f
C1720 vdd.t105 gnd 0.163186f
C1721 vdd.n747 gnd 0.088193f
C1722 vdd.n748 gnd 0.050026f
C1723 vdd.n749 gnd 0.014457f
C1724 vdd.n750 gnd 0.006186f
C1725 vdd.t188 gnd 0.632151f
C1726 vdd.n751 gnd 0.013704f
C1727 vdd.n752 gnd 0.006186f
C1728 vdd.n753 gnd 0.014678f
C1729 vdd.n754 gnd 0.006186f
C1730 vdd.t76 gnd 0.249964f
C1731 vdd.t75 gnd 0.255869f
C1732 vdd.t73 gnd 0.163186f
C1733 vdd.n755 gnd 0.088193f
C1734 vdd.n756 gnd 0.050026f
C1735 vdd.n757 gnd 0.00884f
C1736 vdd.n758 gnd 0.006186f
C1737 vdd.n759 gnd 0.006186f
C1738 vdd.t74 gnd 0.316076f
C1739 vdd.n760 gnd 0.006186f
C1740 vdd.n761 gnd 0.006186f
C1741 vdd.n762 gnd 0.006186f
C1742 vdd.n763 gnd 0.006186f
C1743 vdd.n764 gnd 0.006186f
C1744 vdd.n765 gnd 0.006186f
C1745 vdd.n766 gnd 0.632151f
C1746 vdd.n767 gnd 0.006186f
C1747 vdd.n768 gnd 0.006186f
C1748 vdd.t181 gnd 0.316076f
C1749 vdd.n769 gnd 0.006186f
C1750 vdd.n770 gnd 0.006186f
C1751 vdd.n771 gnd 0.006186f
C1752 vdd.n772 gnd 0.006186f
C1753 vdd.n773 gnd 0.399743f
C1754 vdd.n774 gnd 0.006186f
C1755 vdd.n775 gnd 0.006186f
C1756 vdd.n776 gnd 0.006186f
C1757 vdd.n777 gnd 0.006186f
C1758 vdd.n778 gnd 0.006186f
C1759 vdd.n779 gnd 0.539188f
C1760 vdd.n780 gnd 0.006186f
C1761 vdd.n781 gnd 0.006186f
C1762 vdd.t198 gnd 0.283539f
C1763 vdd.t30 gnd 0.232409f
C1764 vdd.n782 gnd 0.006186f
C1765 vdd.n783 gnd 0.006186f
C1766 vdd.n784 gnd 0.006186f
C1767 vdd.t196 gnd 0.316076f
C1768 vdd.n785 gnd 0.006186f
C1769 vdd.n786 gnd 0.006186f
C1770 vdd.t25 gnd 0.316076f
C1771 vdd.n787 gnd 0.006186f
C1772 vdd.n788 gnd 0.006186f
C1773 vdd.n789 gnd 0.006186f
C1774 vdd.t185 gnd 0.246353f
C1775 vdd.n790 gnd 0.006186f
C1776 vdd.n791 gnd 0.006186f
C1777 vdd.n792 gnd 0.525243f
C1778 vdd.n793 gnd 0.006186f
C1779 vdd.n794 gnd 0.006186f
C1780 vdd.n795 gnd 0.006186f
C1781 vdd.t21 gnd 0.316076f
C1782 vdd.n796 gnd 0.006186f
C1783 vdd.n797 gnd 0.006186f
C1784 vdd.t20 gnd 0.269594f
C1785 vdd.n798 gnd 0.385798f
C1786 vdd.n799 gnd 0.006186f
C1787 vdd.n800 gnd 0.006186f
C1788 vdd.n801 gnd 0.006186f
C1789 vdd.n802 gnd 0.525243f
C1790 vdd.n803 gnd 0.006186f
C1791 vdd.n804 gnd 0.006186f
C1792 vdd.t29 gnd 0.316076f
C1793 vdd.n805 gnd 0.006186f
C1794 vdd.n806 gnd 0.006186f
C1795 vdd.n807 gnd 0.006186f
C1796 vdd.n808 gnd 0.632151f
C1797 vdd.n809 gnd 0.006186f
C1798 vdd.n810 gnd 0.006186f
C1799 vdd.t24 gnd 0.316076f
C1800 vdd.n811 gnd 0.006186f
C1801 vdd.n812 gnd 0.006186f
C1802 vdd.n813 gnd 0.006186f
C1803 vdd.t23 gnd 0.074371f
C1804 vdd.n814 gnd 0.006186f
C1805 vdd.n815 gnd 0.006186f
C1806 vdd.n816 gnd 0.006186f
C1807 vdd.t94 gnd 0.255869f
C1808 vdd.t92 gnd 0.163186f
C1809 vdd.t95 gnd 0.255869f
C1810 vdd.n817 gnd 0.143809f
C1811 vdd.n818 gnd 0.006186f
C1812 vdd.n819 gnd 0.006186f
C1813 vdd.n820 gnd 0.632151f
C1814 vdd.n821 gnd 0.006186f
C1815 vdd.n822 gnd 0.006186f
C1816 vdd.t93 gnd 0.283539f
C1817 vdd.n823 gnd 0.557781f
C1818 vdd.n824 gnd 0.006186f
C1819 vdd.n825 gnd 0.006186f
C1820 vdd.n826 gnd 0.006186f
C1821 vdd.n827 gnd 0.553133f
C1822 vdd.n828 gnd 0.006186f
C1823 vdd.n829 gnd 0.006186f
C1824 vdd.n830 gnd 0.006186f
C1825 vdd.n831 gnd 0.006186f
C1826 vdd.n832 gnd 0.006186f
C1827 vdd.n833 gnd 0.632151f
C1828 vdd.n834 gnd 0.006186f
C1829 vdd.n835 gnd 0.006186f
C1830 vdd.t89 gnd 0.316076f
C1831 vdd.n836 gnd 0.006186f
C1832 vdd.n837 gnd 0.014678f
C1833 vdd.n838 gnd 0.014678f
C1834 vdd.n839 gnd 6.40518f
C1835 vdd.n840 gnd 0.013704f
C1836 vdd.n841 gnd 0.013704f
C1837 vdd.n842 gnd 0.014678f
C1838 vdd.n843 gnd 0.006186f
C1839 vdd.n844 gnd 0.006186f
C1840 vdd.n845 gnd 0.006186f
C1841 vdd.n846 gnd 0.006186f
C1842 vdd.n847 gnd 0.006186f
C1843 vdd.n848 gnd 0.006186f
C1844 vdd.n849 gnd 0.006186f
C1845 vdd.n850 gnd 0.006186f
C1846 vdd.n852 gnd 0.006186f
C1847 vdd.n853 gnd 0.006186f
C1848 vdd.n854 gnd 0.005822f
C1849 vdd.n857 gnd 0.022678f
C1850 vdd.n858 gnd 0.007322f
C1851 vdd.n859 gnd 0.009097f
C1852 vdd.n861 gnd 0.009097f
C1853 vdd.n862 gnd 0.006077f
C1854 vdd.t49 gnd 0.464817f
C1855 vdd.n863 gnd 6.73985f
C1856 vdd.n864 gnd 0.009097f
C1857 vdd.n865 gnd 0.022678f
C1858 vdd.n866 gnd 0.007322f
C1859 vdd.n867 gnd 0.009097f
C1860 vdd.n868 gnd 0.007322f
C1861 vdd.n869 gnd 0.009097f
C1862 vdd.n870 gnd 0.929634f
C1863 vdd.n871 gnd 0.009097f
C1864 vdd.n872 gnd 0.007322f
C1865 vdd.n873 gnd 0.007322f
C1866 vdd.n874 gnd 0.009097f
C1867 vdd.n875 gnd 0.007322f
C1868 vdd.n876 gnd 0.009097f
C1869 vdd.t117 gnd 0.464817f
C1870 vdd.n877 gnd 0.009097f
C1871 vdd.n878 gnd 0.007322f
C1872 vdd.n879 gnd 0.009097f
C1873 vdd.n880 gnd 0.007322f
C1874 vdd.n881 gnd 0.009097f
C1875 vdd.t170 gnd 0.464817f
C1876 vdd.n882 gnd 0.009097f
C1877 vdd.n883 gnd 0.007322f
C1878 vdd.n884 gnd 0.009097f
C1879 vdd.n885 gnd 0.007322f
C1880 vdd.n886 gnd 0.009097f
C1881 vdd.n887 gnd 0.729763f
C1882 vdd.n888 gnd 0.771597f
C1883 vdd.t125 gnd 0.464817f
C1884 vdd.n889 gnd 0.009097f
C1885 vdd.n890 gnd 0.007322f
C1886 vdd.n891 gnd 0.004992f
C1887 vdd.n892 gnd 0.004633f
C1888 vdd.n893 gnd 0.002563f
C1889 vdd.n894 gnd 0.005884f
C1890 vdd.n895 gnd 0.002489f
C1891 vdd.n896 gnd 0.002636f
C1892 vdd.n897 gnd 0.004633f
C1893 vdd.n898 gnd 0.002489f
C1894 vdd.n899 gnd 0.005884f
C1895 vdd.n900 gnd 0.002636f
C1896 vdd.n901 gnd 0.004633f
C1897 vdd.n902 gnd 0.002489f
C1898 vdd.n903 gnd 0.004413f
C1899 vdd.n904 gnd 0.004426f
C1900 vdd.t118 gnd 0.012641f
C1901 vdd.n905 gnd 0.028127f
C1902 vdd.n906 gnd 0.146377f
C1903 vdd.n907 gnd 0.002489f
C1904 vdd.n908 gnd 0.002636f
C1905 vdd.n909 gnd 0.005884f
C1906 vdd.n910 gnd 0.005884f
C1907 vdd.n911 gnd 0.002636f
C1908 vdd.n912 gnd 0.002489f
C1909 vdd.n913 gnd 0.004633f
C1910 vdd.n914 gnd 0.004633f
C1911 vdd.n915 gnd 0.002489f
C1912 vdd.n916 gnd 0.002636f
C1913 vdd.n917 gnd 0.005884f
C1914 vdd.n918 gnd 0.005884f
C1915 vdd.n919 gnd 0.002636f
C1916 vdd.n920 gnd 0.002489f
C1917 vdd.n921 gnd 0.004633f
C1918 vdd.n922 gnd 0.004633f
C1919 vdd.n923 gnd 0.002489f
C1920 vdd.n924 gnd 0.002636f
C1921 vdd.n925 gnd 0.005884f
C1922 vdd.n926 gnd 0.005884f
C1923 vdd.n927 gnd 0.013911f
C1924 vdd.n928 gnd 0.002563f
C1925 vdd.n929 gnd 0.002489f
C1926 vdd.n930 gnd 0.011974f
C1927 vdd.n931 gnd 0.008359f
C1928 vdd.t144 gnd 0.029287f
C1929 vdd.t173 gnd 0.029287f
C1930 vdd.n932 gnd 0.201279f
C1931 vdd.n933 gnd 0.158275f
C1932 vdd.t133 gnd 0.029287f
C1933 vdd.t161 gnd 0.029287f
C1934 vdd.n934 gnd 0.201279f
C1935 vdd.n935 gnd 0.127727f
C1936 vdd.t139 gnd 0.029287f
C1937 vdd.t167 gnd 0.029287f
C1938 vdd.n936 gnd 0.201279f
C1939 vdd.n937 gnd 0.127727f
C1940 vdd.n938 gnd 0.004992f
C1941 vdd.n939 gnd 0.004633f
C1942 vdd.n940 gnd 0.002563f
C1943 vdd.n941 gnd 0.005884f
C1944 vdd.n942 gnd 0.002489f
C1945 vdd.n943 gnd 0.002636f
C1946 vdd.n944 gnd 0.004633f
C1947 vdd.n945 gnd 0.002489f
C1948 vdd.n946 gnd 0.005884f
C1949 vdd.n947 gnd 0.002636f
C1950 vdd.n948 gnd 0.004633f
C1951 vdd.n949 gnd 0.002489f
C1952 vdd.n950 gnd 0.004413f
C1953 vdd.n951 gnd 0.004426f
C1954 vdd.t177 gnd 0.012641f
C1955 vdd.n952 gnd 0.028127f
C1956 vdd.n953 gnd 0.146377f
C1957 vdd.n954 gnd 0.002489f
C1958 vdd.n955 gnd 0.002636f
C1959 vdd.n956 gnd 0.005884f
C1960 vdd.n957 gnd 0.005884f
C1961 vdd.n958 gnd 0.002636f
C1962 vdd.n959 gnd 0.002489f
C1963 vdd.n960 gnd 0.004633f
C1964 vdd.n961 gnd 0.004633f
C1965 vdd.n962 gnd 0.002489f
C1966 vdd.n963 gnd 0.002636f
C1967 vdd.n964 gnd 0.005884f
C1968 vdd.n965 gnd 0.005884f
C1969 vdd.n966 gnd 0.002636f
C1970 vdd.n967 gnd 0.002489f
C1971 vdd.n968 gnd 0.004633f
C1972 vdd.n969 gnd 0.004633f
C1973 vdd.n970 gnd 0.002489f
C1974 vdd.n971 gnd 0.002636f
C1975 vdd.n972 gnd 0.005884f
C1976 vdd.n973 gnd 0.005884f
C1977 vdd.n974 gnd 0.013911f
C1978 vdd.n975 gnd 0.002563f
C1979 vdd.n976 gnd 0.002489f
C1980 vdd.n977 gnd 0.011974f
C1981 vdd.n978 gnd 0.008097f
C1982 vdd.n979 gnd 0.09503f
C1983 vdd.n980 gnd 0.004992f
C1984 vdd.n981 gnd 0.004633f
C1985 vdd.n982 gnd 0.002563f
C1986 vdd.n983 gnd 0.005884f
C1987 vdd.n984 gnd 0.002489f
C1988 vdd.n985 gnd 0.002636f
C1989 vdd.n986 gnd 0.004633f
C1990 vdd.n987 gnd 0.002489f
C1991 vdd.n988 gnd 0.005884f
C1992 vdd.n989 gnd 0.002636f
C1993 vdd.n990 gnd 0.004633f
C1994 vdd.n991 gnd 0.002489f
C1995 vdd.n992 gnd 0.004413f
C1996 vdd.n993 gnd 0.004426f
C1997 vdd.t168 gnd 0.012641f
C1998 vdd.n994 gnd 0.028127f
C1999 vdd.n995 gnd 0.146377f
C2000 vdd.n996 gnd 0.002489f
C2001 vdd.n997 gnd 0.002636f
C2002 vdd.n998 gnd 0.005884f
C2003 vdd.n999 gnd 0.005884f
C2004 vdd.n1000 gnd 0.002636f
C2005 vdd.n1001 gnd 0.002489f
C2006 vdd.n1002 gnd 0.004633f
C2007 vdd.n1003 gnd 0.004633f
C2008 vdd.n1004 gnd 0.002489f
C2009 vdd.n1005 gnd 0.002636f
C2010 vdd.n1006 gnd 0.005884f
C2011 vdd.n1007 gnd 0.005884f
C2012 vdd.n1008 gnd 0.002636f
C2013 vdd.n1009 gnd 0.002489f
C2014 vdd.n1010 gnd 0.004633f
C2015 vdd.n1011 gnd 0.004633f
C2016 vdd.n1012 gnd 0.002489f
C2017 vdd.n1013 gnd 0.002636f
C2018 vdd.n1014 gnd 0.005884f
C2019 vdd.n1015 gnd 0.005884f
C2020 vdd.n1016 gnd 0.013911f
C2021 vdd.n1017 gnd 0.002563f
C2022 vdd.n1018 gnd 0.002489f
C2023 vdd.n1019 gnd 0.011974f
C2024 vdd.n1020 gnd 0.008359f
C2025 vdd.t126 gnd 0.029287f
C2026 vdd.t171 gnd 0.029287f
C2027 vdd.n1021 gnd 0.201279f
C2028 vdd.n1022 gnd 0.158275f
C2029 vdd.t166 gnd 0.029287f
C2030 vdd.t157 gnd 0.029287f
C2031 vdd.n1023 gnd 0.201279f
C2032 vdd.n1024 gnd 0.127727f
C2033 vdd.t142 gnd 0.029287f
C2034 vdd.t122 gnd 0.029287f
C2035 vdd.n1025 gnd 0.201279f
C2036 vdd.n1026 gnd 0.127727f
C2037 vdd.n1027 gnd 0.004992f
C2038 vdd.n1028 gnd 0.004633f
C2039 vdd.n1029 gnd 0.002563f
C2040 vdd.n1030 gnd 0.005884f
C2041 vdd.n1031 gnd 0.002489f
C2042 vdd.n1032 gnd 0.002636f
C2043 vdd.n1033 gnd 0.004633f
C2044 vdd.n1034 gnd 0.002489f
C2045 vdd.n1035 gnd 0.005884f
C2046 vdd.n1036 gnd 0.002636f
C2047 vdd.n1037 gnd 0.004633f
C2048 vdd.n1038 gnd 0.002489f
C2049 vdd.n1039 gnd 0.004413f
C2050 vdd.n1040 gnd 0.004426f
C2051 vdd.t155 gnd 0.012641f
C2052 vdd.n1041 gnd 0.028127f
C2053 vdd.n1042 gnd 0.146377f
C2054 vdd.n1043 gnd 0.002489f
C2055 vdd.n1044 gnd 0.002636f
C2056 vdd.n1045 gnd 0.005884f
C2057 vdd.n1046 gnd 0.005884f
C2058 vdd.n1047 gnd 0.002636f
C2059 vdd.n1048 gnd 0.002489f
C2060 vdd.n1049 gnd 0.004633f
C2061 vdd.n1050 gnd 0.004633f
C2062 vdd.n1051 gnd 0.002489f
C2063 vdd.n1052 gnd 0.002636f
C2064 vdd.n1053 gnd 0.005884f
C2065 vdd.n1054 gnd 0.005884f
C2066 vdd.n1055 gnd 0.002636f
C2067 vdd.n1056 gnd 0.002489f
C2068 vdd.n1057 gnd 0.004633f
C2069 vdd.n1058 gnd 0.004633f
C2070 vdd.n1059 gnd 0.002489f
C2071 vdd.n1060 gnd 0.002636f
C2072 vdd.n1061 gnd 0.005884f
C2073 vdd.n1062 gnd 0.005884f
C2074 vdd.n1063 gnd 0.013911f
C2075 vdd.n1064 gnd 0.002563f
C2076 vdd.n1065 gnd 0.002489f
C2077 vdd.n1066 gnd 0.011974f
C2078 vdd.n1067 gnd 0.008097f
C2079 vdd.n1068 gnd 0.056533f
C2080 vdd.n1069 gnd 0.203704f
C2081 vdd.n1070 gnd 0.004992f
C2082 vdd.n1071 gnd 0.004633f
C2083 vdd.n1072 gnd 0.002563f
C2084 vdd.n1073 gnd 0.005884f
C2085 vdd.n1074 gnd 0.002489f
C2086 vdd.n1075 gnd 0.002636f
C2087 vdd.n1076 gnd 0.004633f
C2088 vdd.n1077 gnd 0.002489f
C2089 vdd.n1078 gnd 0.005884f
C2090 vdd.n1079 gnd 0.002636f
C2091 vdd.n1080 gnd 0.004633f
C2092 vdd.n1081 gnd 0.002489f
C2093 vdd.n1082 gnd 0.004413f
C2094 vdd.n1083 gnd 0.004426f
C2095 vdd.t176 gnd 0.012641f
C2096 vdd.n1084 gnd 0.028127f
C2097 vdd.n1085 gnd 0.146377f
C2098 vdd.n1086 gnd 0.002489f
C2099 vdd.n1087 gnd 0.002636f
C2100 vdd.n1088 gnd 0.005884f
C2101 vdd.n1089 gnd 0.005884f
C2102 vdd.n1090 gnd 0.002636f
C2103 vdd.n1091 gnd 0.002489f
C2104 vdd.n1092 gnd 0.004633f
C2105 vdd.n1093 gnd 0.004633f
C2106 vdd.n1094 gnd 0.002489f
C2107 vdd.n1095 gnd 0.002636f
C2108 vdd.n1096 gnd 0.005884f
C2109 vdd.n1097 gnd 0.005884f
C2110 vdd.n1098 gnd 0.002636f
C2111 vdd.n1099 gnd 0.002489f
C2112 vdd.n1100 gnd 0.004633f
C2113 vdd.n1101 gnd 0.004633f
C2114 vdd.n1102 gnd 0.002489f
C2115 vdd.n1103 gnd 0.002636f
C2116 vdd.n1104 gnd 0.005884f
C2117 vdd.n1105 gnd 0.005884f
C2118 vdd.n1106 gnd 0.013911f
C2119 vdd.n1107 gnd 0.002563f
C2120 vdd.n1108 gnd 0.002489f
C2121 vdd.n1109 gnd 0.011974f
C2122 vdd.n1110 gnd 0.008359f
C2123 vdd.t131 gnd 0.029287f
C2124 vdd.t175 gnd 0.029287f
C2125 vdd.n1111 gnd 0.201279f
C2126 vdd.n1112 gnd 0.158275f
C2127 vdd.t174 gnd 0.029287f
C2128 vdd.t163 gnd 0.029287f
C2129 vdd.n1113 gnd 0.201279f
C2130 vdd.n1114 gnd 0.127727f
C2131 vdd.t150 gnd 0.029287f
C2132 vdd.t129 gnd 0.029287f
C2133 vdd.n1115 gnd 0.201279f
C2134 vdd.n1116 gnd 0.127727f
C2135 vdd.n1117 gnd 0.004992f
C2136 vdd.n1118 gnd 0.004633f
C2137 vdd.n1119 gnd 0.002563f
C2138 vdd.n1120 gnd 0.005884f
C2139 vdd.n1121 gnd 0.002489f
C2140 vdd.n1122 gnd 0.002636f
C2141 vdd.n1123 gnd 0.004633f
C2142 vdd.n1124 gnd 0.002489f
C2143 vdd.n1125 gnd 0.005884f
C2144 vdd.n1126 gnd 0.002636f
C2145 vdd.n1127 gnd 0.004633f
C2146 vdd.n1128 gnd 0.002489f
C2147 vdd.n1129 gnd 0.004413f
C2148 vdd.n1130 gnd 0.004426f
C2149 vdd.t162 gnd 0.012641f
C2150 vdd.n1131 gnd 0.028127f
C2151 vdd.n1132 gnd 0.146377f
C2152 vdd.n1133 gnd 0.002489f
C2153 vdd.n1134 gnd 0.002636f
C2154 vdd.n1135 gnd 0.005884f
C2155 vdd.n1136 gnd 0.005884f
C2156 vdd.n1137 gnd 0.002636f
C2157 vdd.n1138 gnd 0.002489f
C2158 vdd.n1139 gnd 0.004633f
C2159 vdd.n1140 gnd 0.004633f
C2160 vdd.n1141 gnd 0.002489f
C2161 vdd.n1142 gnd 0.002636f
C2162 vdd.n1143 gnd 0.005884f
C2163 vdd.n1144 gnd 0.005884f
C2164 vdd.n1145 gnd 0.002636f
C2165 vdd.n1146 gnd 0.002489f
C2166 vdd.n1147 gnd 0.004633f
C2167 vdd.n1148 gnd 0.004633f
C2168 vdd.n1149 gnd 0.002489f
C2169 vdd.n1150 gnd 0.002636f
C2170 vdd.n1151 gnd 0.005884f
C2171 vdd.n1152 gnd 0.005884f
C2172 vdd.n1153 gnd 0.013911f
C2173 vdd.n1154 gnd 0.002563f
C2174 vdd.n1155 gnd 0.002489f
C2175 vdd.n1156 gnd 0.011974f
C2176 vdd.n1157 gnd 0.008097f
C2177 vdd.n1158 gnd 0.056533f
C2178 vdd.n1159 gnd 0.220485f
C2179 vdd.n1160 gnd 1.85301f
C2180 vdd.n1161 gnd 0.536555f
C2181 vdd.n1162 gnd 0.007322f
C2182 vdd.n1163 gnd 0.009097f
C2183 vdd.n1164 gnd 0.571725f
C2184 vdd.n1165 gnd 0.009097f
C2185 vdd.n1166 gnd 0.007322f
C2186 vdd.n1167 gnd 0.009097f
C2187 vdd.n1168 gnd 0.007322f
C2188 vdd.n1169 gnd 0.009097f
C2189 vdd.t121 gnd 0.464817f
C2190 vdd.t132 gnd 0.464817f
C2191 vdd.n1170 gnd 0.009097f
C2192 vdd.n1171 gnd 0.007322f
C2193 vdd.n1172 gnd 0.009097f
C2194 vdd.n1173 gnd 0.007322f
C2195 vdd.n1174 gnd 0.009097f
C2196 vdd.t138 gnd 0.464817f
C2197 vdd.n1175 gnd 0.009097f
C2198 vdd.n1176 gnd 0.007322f
C2199 vdd.n1177 gnd 0.009097f
C2200 vdd.n1178 gnd 0.007322f
C2201 vdd.n1179 gnd 0.009097f
C2202 vdd.t154 gnd 0.464817f
C2203 vdd.n1180 gnd 0.673985f
C2204 vdd.n1181 gnd 0.009097f
C2205 vdd.n1182 gnd 0.007322f
C2206 vdd.n1183 gnd 0.009097f
C2207 vdd.n1184 gnd 0.007322f
C2208 vdd.n1185 gnd 0.009097f
C2209 vdd.n1186 gnd 0.929634f
C2210 vdd.n1187 gnd 0.009097f
C2211 vdd.n1188 gnd 0.007322f
C2212 vdd.n1189 gnd 0.022169f
C2213 vdd.n1190 gnd 0.006077f
C2214 vdd.n1191 gnd 0.022169f
C2215 vdd.t53 gnd 0.464817f
C2216 vdd.n1192 gnd 0.022169f
C2217 vdd.n1193 gnd 0.006077f
C2218 vdd.n1194 gnd 0.009097f
C2219 vdd.n1195 gnd 0.007322f
C2220 vdd.n1196 gnd 0.009097f
C2221 vdd.n1227 gnd 0.022678f
C2222 vdd.n1228 gnd 1.37121f
C2223 vdd.n1229 gnd 0.009097f
C2224 vdd.n1230 gnd 0.007322f
C2225 vdd.n1231 gnd 0.009097f
C2226 vdd.n1232 gnd 0.009097f
C2227 vdd.n1233 gnd 0.009097f
C2228 vdd.n1234 gnd 0.009097f
C2229 vdd.n1235 gnd 0.009097f
C2230 vdd.n1236 gnd 0.007322f
C2231 vdd.n1237 gnd 0.009097f
C2232 vdd.n1238 gnd 0.009097f
C2233 vdd.n1239 gnd 0.009097f
C2234 vdd.n1240 gnd 0.009097f
C2235 vdd.n1241 gnd 0.009097f
C2236 vdd.n1242 gnd 0.007322f
C2237 vdd.n1243 gnd 0.009097f
C2238 vdd.n1244 gnd 0.009097f
C2239 vdd.n1245 gnd 0.009097f
C2240 vdd.n1246 gnd 0.009097f
C2241 vdd.n1247 gnd 0.009097f
C2242 vdd.n1248 gnd 0.007322f
C2243 vdd.n1249 gnd 0.009097f
C2244 vdd.n1250 gnd 0.009097f
C2245 vdd.n1251 gnd 0.009097f
C2246 vdd.n1252 gnd 0.009097f
C2247 vdd.n1253 gnd 0.009097f
C2248 vdd.t103 gnd 0.111913f
C2249 vdd.t104 gnd 0.119604f
C2250 vdd.t102 gnd 0.146157f
C2251 vdd.n1254 gnd 0.187352f
C2252 vdd.n1255 gnd 0.158142f
C2253 vdd.n1256 gnd 0.015668f
C2254 vdd.n1257 gnd 0.009097f
C2255 vdd.n1258 gnd 0.009097f
C2256 vdd.n1259 gnd 0.009097f
C2257 vdd.n1260 gnd 0.009097f
C2258 vdd.n1261 gnd 0.009097f
C2259 vdd.n1262 gnd 0.007322f
C2260 vdd.n1263 gnd 0.009097f
C2261 vdd.n1264 gnd 0.009097f
C2262 vdd.n1265 gnd 0.009097f
C2263 vdd.n1266 gnd 0.009097f
C2264 vdd.n1267 gnd 0.009097f
C2265 vdd.n1268 gnd 0.007322f
C2266 vdd.n1269 gnd 0.009097f
C2267 vdd.n1270 gnd 0.009097f
C2268 vdd.n1271 gnd 0.009097f
C2269 vdd.n1272 gnd 0.009097f
C2270 vdd.n1273 gnd 0.009097f
C2271 vdd.n1274 gnd 0.007322f
C2272 vdd.n1275 gnd 0.009097f
C2273 vdd.n1276 gnd 0.009097f
C2274 vdd.n1277 gnd 0.009097f
C2275 vdd.n1278 gnd 0.009097f
C2276 vdd.n1279 gnd 0.009097f
C2277 vdd.n1280 gnd 0.007322f
C2278 vdd.n1281 gnd 0.009097f
C2279 vdd.n1282 gnd 0.009097f
C2280 vdd.n1283 gnd 0.009097f
C2281 vdd.n1284 gnd 0.009097f
C2282 vdd.n1285 gnd 0.009097f
C2283 vdd.n1286 gnd 0.007322f
C2284 vdd.n1287 gnd 0.009097f
C2285 vdd.n1288 gnd 0.009097f
C2286 vdd.n1289 gnd 0.009097f
C2287 vdd.n1290 gnd 0.009097f
C2288 vdd.n1291 gnd 0.007322f
C2289 vdd.n1292 gnd 0.009097f
C2290 vdd.n1293 gnd 0.009097f
C2291 vdd.n1294 gnd 0.009097f
C2292 vdd.n1295 gnd 0.009097f
C2293 vdd.n1296 gnd 0.009097f
C2294 vdd.n1297 gnd 0.007322f
C2295 vdd.n1298 gnd 0.009097f
C2296 vdd.n1299 gnd 0.009097f
C2297 vdd.n1300 gnd 0.009097f
C2298 vdd.n1301 gnd 0.009097f
C2299 vdd.n1302 gnd 0.009097f
C2300 vdd.n1303 gnd 0.007322f
C2301 vdd.n1304 gnd 0.009097f
C2302 vdd.n1305 gnd 0.009097f
C2303 vdd.n1306 gnd 0.009097f
C2304 vdd.n1307 gnd 0.009097f
C2305 vdd.n1308 gnd 0.009097f
C2306 vdd.n1309 gnd 0.007322f
C2307 vdd.n1310 gnd 0.009097f
C2308 vdd.n1311 gnd 0.009097f
C2309 vdd.n1312 gnd 0.009097f
C2310 vdd.n1313 gnd 0.009097f
C2311 vdd.n1314 gnd 0.009097f
C2312 vdd.n1315 gnd 0.007322f
C2313 vdd.n1316 gnd 0.009097f
C2314 vdd.n1317 gnd 0.009097f
C2315 vdd.n1318 gnd 0.009097f
C2316 vdd.n1319 gnd 0.009097f
C2317 vdd.t54 gnd 0.111913f
C2318 vdd.t55 gnd 0.119604f
C2319 vdd.t52 gnd 0.146157f
C2320 vdd.n1320 gnd 0.187352f
C2321 vdd.n1321 gnd 0.158142f
C2322 vdd.n1322 gnd 0.012008f
C2323 vdd.n1323 gnd 0.003478f
C2324 vdd.n1324 gnd 0.022678f
C2325 vdd.n1325 gnd 0.009097f
C2326 vdd.n1326 gnd 0.003844f
C2327 vdd.n1327 gnd 0.007322f
C2328 vdd.n1328 gnd 0.007322f
C2329 vdd.n1329 gnd 0.009097f
C2330 vdd.n1330 gnd 0.009097f
C2331 vdd.n1331 gnd 0.009097f
C2332 vdd.n1332 gnd 0.007322f
C2333 vdd.n1333 gnd 0.007322f
C2334 vdd.n1334 gnd 0.007322f
C2335 vdd.n1335 gnd 0.009097f
C2336 vdd.n1336 gnd 0.009097f
C2337 vdd.n1337 gnd 0.009097f
C2338 vdd.n1338 gnd 0.007322f
C2339 vdd.n1339 gnd 0.007322f
C2340 vdd.n1340 gnd 0.007322f
C2341 vdd.n1341 gnd 0.009097f
C2342 vdd.n1342 gnd 0.009097f
C2343 vdd.n1343 gnd 0.009097f
C2344 vdd.n1344 gnd 0.007322f
C2345 vdd.n1345 gnd 0.007322f
C2346 vdd.n1346 gnd 0.007322f
C2347 vdd.n1347 gnd 0.009097f
C2348 vdd.n1348 gnd 0.009097f
C2349 vdd.n1349 gnd 0.009097f
C2350 vdd.n1350 gnd 0.007322f
C2351 vdd.n1351 gnd 0.007322f
C2352 vdd.n1352 gnd 0.007322f
C2353 vdd.n1353 gnd 0.009097f
C2354 vdd.n1354 gnd 0.009097f
C2355 vdd.n1355 gnd 0.009097f
C2356 vdd.n1356 gnd 0.007248f
C2357 vdd.n1357 gnd 0.009097f
C2358 vdd.t100 gnd 0.111913f
C2359 vdd.t101 gnd 0.119604f
C2360 vdd.t99 gnd 0.146157f
C2361 vdd.n1358 gnd 0.187352f
C2362 vdd.n1359 gnd 0.158142f
C2363 vdd.n1360 gnd 0.015668f
C2364 vdd.n1361 gnd 0.004979f
C2365 vdd.n1362 gnd 0.009097f
C2366 vdd.n1363 gnd 0.009097f
C2367 vdd.n1364 gnd 0.009097f
C2368 vdd.n1365 gnd 0.007322f
C2369 vdd.n1366 gnd 0.007322f
C2370 vdd.n1367 gnd 0.007322f
C2371 vdd.n1368 gnd 0.009097f
C2372 vdd.n1369 gnd 0.009097f
C2373 vdd.n1370 gnd 0.009097f
C2374 vdd.n1371 gnd 0.007322f
C2375 vdd.n1372 gnd 0.007322f
C2376 vdd.n1373 gnd 0.007322f
C2377 vdd.n1374 gnd 0.009097f
C2378 vdd.n1375 gnd 0.009097f
C2379 vdd.n1376 gnd 0.009097f
C2380 vdd.n1377 gnd 0.007322f
C2381 vdd.n1378 gnd 0.007322f
C2382 vdd.n1379 gnd 0.007322f
C2383 vdd.n1380 gnd 0.009097f
C2384 vdd.n1381 gnd 0.009097f
C2385 vdd.n1382 gnd 0.009097f
C2386 vdd.n1383 gnd 0.007322f
C2387 vdd.n1384 gnd 0.007322f
C2388 vdd.n1385 gnd 0.007322f
C2389 vdd.n1386 gnd 0.009097f
C2390 vdd.n1387 gnd 0.009097f
C2391 vdd.n1388 gnd 0.009097f
C2392 vdd.n1389 gnd 0.007322f
C2393 vdd.n1390 gnd 0.007322f
C2394 vdd.n1391 gnd 0.006114f
C2395 vdd.n1392 gnd 0.009097f
C2396 vdd.n1393 gnd 0.009097f
C2397 vdd.n1394 gnd 0.009097f
C2398 vdd.n1395 gnd 0.006114f
C2399 vdd.n1396 gnd 0.007322f
C2400 vdd.n1397 gnd 0.007322f
C2401 vdd.n1398 gnd 0.009097f
C2402 vdd.n1399 gnd 0.009097f
C2403 vdd.n1400 gnd 0.009097f
C2404 vdd.n1401 gnd 0.007322f
C2405 vdd.n1402 gnd 0.007322f
C2406 vdd.n1403 gnd 0.007322f
C2407 vdd.n1404 gnd 0.009097f
C2408 vdd.n1405 gnd 0.009097f
C2409 vdd.n1406 gnd 0.009097f
C2410 vdd.n1407 gnd 0.007322f
C2411 vdd.n1408 gnd 0.007322f
C2412 vdd.n1409 gnd 0.007322f
C2413 vdd.n1410 gnd 0.009097f
C2414 vdd.n1411 gnd 0.009097f
C2415 vdd.n1412 gnd 0.009097f
C2416 vdd.n1413 gnd 0.007322f
C2417 vdd.n1414 gnd 0.007322f
C2418 vdd.n1415 gnd 0.007322f
C2419 vdd.n1416 gnd 0.009097f
C2420 vdd.n1417 gnd 0.009097f
C2421 vdd.n1418 gnd 0.009097f
C2422 vdd.n1419 gnd 0.007322f
C2423 vdd.n1420 gnd 0.009097f
C2424 vdd.n1421 gnd 2.22183f
C2425 vdd.n1423 gnd 0.022678f
C2426 vdd.n1424 gnd 0.006077f
C2427 vdd.n1425 gnd 0.022678f
C2428 vdd.n1426 gnd 0.022169f
C2429 vdd.n1427 gnd 0.009097f
C2430 vdd.n1428 gnd 0.007322f
C2431 vdd.n1429 gnd 0.009097f
C2432 vdd.n1430 gnd 0.488058f
C2433 vdd.n1431 gnd 0.009097f
C2434 vdd.n1432 gnd 0.007322f
C2435 vdd.n1433 gnd 0.009097f
C2436 vdd.n1434 gnd 0.009097f
C2437 vdd.n1435 gnd 0.009097f
C2438 vdd.n1436 gnd 0.007322f
C2439 vdd.n1437 gnd 0.009097f
C2440 vdd.n1438 gnd 0.832023f
C2441 vdd.n1439 gnd 0.929634f
C2442 vdd.n1440 gnd 0.009097f
C2443 vdd.n1441 gnd 0.007322f
C2444 vdd.n1442 gnd 0.009097f
C2445 vdd.n1443 gnd 0.009097f
C2446 vdd.n1444 gnd 0.009097f
C2447 vdd.n1445 gnd 0.007322f
C2448 vdd.n1446 gnd 0.009097f
C2449 vdd.n1447 gnd 0.562429f
C2450 vdd.n1448 gnd 0.009097f
C2451 vdd.n1449 gnd 0.007322f
C2452 vdd.n1450 gnd 0.009097f
C2453 vdd.n1451 gnd 0.009097f
C2454 vdd.n1452 gnd 0.009097f
C2455 vdd.n1453 gnd 0.007322f
C2456 vdd.n1454 gnd 0.009097f
C2457 vdd.n1455 gnd 0.515947f
C2458 vdd.n1456 gnd 0.720467f
C2459 vdd.n1457 gnd 0.009097f
C2460 vdd.n1458 gnd 0.007322f
C2461 vdd.n1459 gnd 0.009097f
C2462 vdd.n1460 gnd 0.009097f
C2463 vdd.n1461 gnd 0.006991f
C2464 vdd.n1462 gnd 0.009097f
C2465 vdd.n1463 gnd 0.007322f
C2466 vdd.n1464 gnd 0.009097f
C2467 vdd.n1465 gnd 0.771597f
C2468 vdd.n1466 gnd 0.009097f
C2469 vdd.n1467 gnd 0.007322f
C2470 vdd.n1468 gnd 0.009097f
C2471 vdd.n1469 gnd 0.009097f
C2472 vdd.n1470 gnd 0.009097f
C2473 vdd.n1471 gnd 0.007322f
C2474 vdd.n1472 gnd 0.009097f
C2475 vdd.t156 gnd 0.464817f
C2476 vdd.n1473 gnd 0.664689f
C2477 vdd.n1474 gnd 0.009097f
C2478 vdd.n1475 gnd 0.007322f
C2479 vdd.n1476 gnd 0.006991f
C2480 vdd.n1477 gnd 0.009097f
C2481 vdd.n1478 gnd 0.009097f
C2482 vdd.n1479 gnd 0.007322f
C2483 vdd.n1480 gnd 0.009097f
C2484 vdd.n1481 gnd 0.506651f
C2485 vdd.n1482 gnd 0.009097f
C2486 vdd.n1483 gnd 0.007322f
C2487 vdd.n1484 gnd 0.009097f
C2488 vdd.n1485 gnd 0.009097f
C2489 vdd.n1486 gnd 0.009097f
C2490 vdd.n1487 gnd 0.007322f
C2491 vdd.n1488 gnd 0.009097f
C2492 vdd.n1489 gnd 0.655392f
C2493 vdd.n1490 gnd 0.581022f
C2494 vdd.n1491 gnd 0.009097f
C2495 vdd.n1492 gnd 0.007322f
C2496 vdd.n1493 gnd 0.009097f
C2497 vdd.n1494 gnd 0.009097f
C2498 vdd.n1495 gnd 0.009097f
C2499 vdd.n1496 gnd 0.007322f
C2500 vdd.n1497 gnd 0.009097f
C2501 vdd.n1498 gnd 0.739059f
C2502 vdd.n1499 gnd 0.009097f
C2503 vdd.n1500 gnd 0.007322f
C2504 vdd.n1501 gnd 0.009097f
C2505 vdd.n1502 gnd 0.009097f
C2506 vdd.n1503 gnd 0.022169f
C2507 vdd.n1504 gnd 0.009097f
C2508 vdd.n1505 gnd 0.009097f
C2509 vdd.n1506 gnd 0.007322f
C2510 vdd.n1507 gnd 0.009097f
C2511 vdd.n1508 gnd 0.581022f
C2512 vdd.n1509 gnd 0.929634f
C2513 vdd.n1510 gnd 0.009097f
C2514 vdd.n1511 gnd 0.007322f
C2515 vdd.n1512 gnd 0.009097f
C2516 vdd.n1513 gnd 0.009097f
C2517 vdd.n1514 gnd 0.007823f
C2518 vdd.n1515 gnd 0.007322f
C2519 vdd.n1517 gnd 0.009097f
C2520 vdd.n1519 gnd 0.007322f
C2521 vdd.n1520 gnd 0.009097f
C2522 vdd.n1521 gnd 0.007322f
C2523 vdd.n1523 gnd 0.009097f
C2524 vdd.n1524 gnd 0.007322f
C2525 vdd.n1525 gnd 0.009097f
C2526 vdd.n1526 gnd 0.009097f
C2527 vdd.n1527 gnd 0.009097f
C2528 vdd.n1528 gnd 0.009097f
C2529 vdd.n1529 gnd 0.009097f
C2530 vdd.n1530 gnd 0.007322f
C2531 vdd.n1532 gnd 0.009097f
C2532 vdd.n1533 gnd 0.009097f
C2533 vdd.n1534 gnd 0.009097f
C2534 vdd.n1535 gnd 0.009097f
C2535 vdd.n1536 gnd 0.009097f
C2536 vdd.n1537 gnd 0.007322f
C2537 vdd.n1539 gnd 0.009097f
C2538 vdd.n1540 gnd 0.009097f
C2539 vdd.n1541 gnd 0.009097f
C2540 vdd.n1542 gnd 0.009097f
C2541 vdd.n1543 gnd 0.006114f
C2542 vdd.t69 gnd 0.111913f
C2543 vdd.t68 gnd 0.119604f
C2544 vdd.t67 gnd 0.146157f
C2545 vdd.n1544 gnd 0.187352f
C2546 vdd.n1545 gnd 0.15741f
C2547 vdd.n1547 gnd 0.009097f
C2548 vdd.n1548 gnd 0.009097f
C2549 vdd.n1549 gnd 0.007322f
C2550 vdd.n1550 gnd 0.009097f
C2551 vdd.n1552 gnd 0.009097f
C2552 vdd.n1553 gnd 0.009097f
C2553 vdd.n1554 gnd 0.009097f
C2554 vdd.n1555 gnd 0.009097f
C2555 vdd.n1556 gnd 0.007322f
C2556 vdd.n1558 gnd 0.009097f
C2557 vdd.n1559 gnd 0.009097f
C2558 vdd.n1560 gnd 0.009097f
C2559 vdd.n1561 gnd 0.009097f
C2560 vdd.n1562 gnd 0.009097f
C2561 vdd.n1563 gnd 0.007322f
C2562 vdd.n1565 gnd 0.009097f
C2563 vdd.n1566 gnd 0.009097f
C2564 vdd.n1567 gnd 0.009097f
C2565 vdd.n1568 gnd 0.009097f
C2566 vdd.n1569 gnd 0.009097f
C2567 vdd.n1570 gnd 0.007322f
C2568 vdd.n1572 gnd 0.009097f
C2569 vdd.n1573 gnd 0.009097f
C2570 vdd.n1574 gnd 0.009097f
C2571 vdd.n1575 gnd 0.009097f
C2572 vdd.n1576 gnd 0.009097f
C2573 vdd.n1577 gnd 0.007322f
C2574 vdd.n1579 gnd 0.009097f
C2575 vdd.n1580 gnd 0.009097f
C2576 vdd.n1581 gnd 0.009097f
C2577 vdd.n1582 gnd 0.009097f
C2578 vdd.n1583 gnd 0.007248f
C2579 vdd.t62 gnd 0.111913f
C2580 vdd.t61 gnd 0.119604f
C2581 vdd.t60 gnd 0.146157f
C2582 vdd.n1584 gnd 0.187352f
C2583 vdd.n1585 gnd 0.15741f
C2584 vdd.n1587 gnd 0.009097f
C2585 vdd.n1588 gnd 0.009097f
C2586 vdd.n1589 gnd 0.007322f
C2587 vdd.n1590 gnd 0.009097f
C2588 vdd.n1592 gnd 0.009097f
C2589 vdd.n1593 gnd 0.009097f
C2590 vdd.n1594 gnd 0.009097f
C2591 vdd.n1595 gnd 0.009097f
C2592 vdd.n1596 gnd 0.007322f
C2593 vdd.n1598 gnd 0.009097f
C2594 vdd.n1599 gnd 0.009097f
C2595 vdd.n1600 gnd 0.009097f
C2596 vdd.n1601 gnd 0.009097f
C2597 vdd.n1602 gnd 0.009097f
C2598 vdd.n1603 gnd 0.007322f
C2599 vdd.n1605 gnd 0.009097f
C2600 vdd.n1606 gnd 0.009097f
C2601 vdd.n1607 gnd 0.009097f
C2602 vdd.n1608 gnd 0.009097f
C2603 vdd.n1609 gnd 0.009097f
C2604 vdd.n1610 gnd 0.009097f
C2605 vdd.n1611 gnd 0.007322f
C2606 vdd.n1613 gnd 0.009097f
C2607 vdd.n1615 gnd 0.009097f
C2608 vdd.n1616 gnd 0.007322f
C2609 vdd.n1617 gnd 0.007322f
C2610 vdd.n1618 gnd 0.009097f
C2611 vdd.n1620 gnd 0.009097f
C2612 vdd.n1621 gnd 0.007322f
C2613 vdd.n1622 gnd 0.007322f
C2614 vdd.n1623 gnd 0.009097f
C2615 vdd.n1625 gnd 0.009097f
C2616 vdd.n1626 gnd 0.009097f
C2617 vdd.n1627 gnd 0.007322f
C2618 vdd.n1628 gnd 0.007322f
C2619 vdd.n1629 gnd 0.007322f
C2620 vdd.n1630 gnd 0.009097f
C2621 vdd.n1632 gnd 0.009097f
C2622 vdd.n1633 gnd 0.009097f
C2623 vdd.n1634 gnd 0.007322f
C2624 vdd.n1635 gnd 0.007322f
C2625 vdd.n1636 gnd 0.007322f
C2626 vdd.n1637 gnd 0.009097f
C2627 vdd.n1639 gnd 0.009097f
C2628 vdd.n1640 gnd 0.009097f
C2629 vdd.n1641 gnd 0.007322f
C2630 vdd.n1642 gnd 0.007322f
C2631 vdd.n1643 gnd 0.007322f
C2632 vdd.n1644 gnd 0.009097f
C2633 vdd.n1646 gnd 0.009097f
C2634 vdd.n1647 gnd 0.009097f
C2635 vdd.n1648 gnd 0.007322f
C2636 vdd.n1649 gnd 0.009097f
C2637 vdd.n1650 gnd 0.009097f
C2638 vdd.n1651 gnd 0.009097f
C2639 vdd.n1652 gnd 0.014936f
C2640 vdd.n1653 gnd 0.004979f
C2641 vdd.n1654 gnd 0.007322f
C2642 vdd.n1655 gnd 0.009097f
C2643 vdd.n1657 gnd 0.009097f
C2644 vdd.n1658 gnd 0.009097f
C2645 vdd.n1659 gnd 0.007322f
C2646 vdd.n1660 gnd 0.007322f
C2647 vdd.n1661 gnd 0.007322f
C2648 vdd.n1662 gnd 0.009097f
C2649 vdd.n1664 gnd 0.009097f
C2650 vdd.n1665 gnd 0.009097f
C2651 vdd.n1666 gnd 0.007322f
C2652 vdd.n1667 gnd 0.007322f
C2653 vdd.n1668 gnd 0.007322f
C2654 vdd.n1669 gnd 0.009097f
C2655 vdd.n1671 gnd 0.009097f
C2656 vdd.n1672 gnd 0.009097f
C2657 vdd.n1673 gnd 0.007322f
C2658 vdd.n1674 gnd 0.007322f
C2659 vdd.n1675 gnd 0.007322f
C2660 vdd.n1676 gnd 0.009097f
C2661 vdd.n1678 gnd 0.009097f
C2662 vdd.n1679 gnd 0.009097f
C2663 vdd.n1680 gnd 0.007322f
C2664 vdd.n1681 gnd 0.007322f
C2665 vdd.n1682 gnd 0.007322f
C2666 vdd.n1683 gnd 0.009097f
C2667 vdd.n1685 gnd 0.009097f
C2668 vdd.n1686 gnd 0.009097f
C2669 vdd.n1687 gnd 0.007322f
C2670 vdd.n1688 gnd 0.009097f
C2671 vdd.n1689 gnd 0.009097f
C2672 vdd.n1690 gnd 0.009097f
C2673 vdd.n1691 gnd 0.014936f
C2674 vdd.n1692 gnd 0.006114f
C2675 vdd.n1693 gnd 0.007322f
C2676 vdd.n1694 gnd 0.009097f
C2677 vdd.n1696 gnd 0.009097f
C2678 vdd.n1697 gnd 0.009097f
C2679 vdd.n1698 gnd 0.007322f
C2680 vdd.n1699 gnd 0.007322f
C2681 vdd.n1700 gnd 0.007322f
C2682 vdd.n1701 gnd 0.009097f
C2683 vdd.n1703 gnd 0.009097f
C2684 vdd.n1704 gnd 0.009097f
C2685 vdd.n1705 gnd 0.007322f
C2686 vdd.n1706 gnd 0.007322f
C2687 vdd.n1707 gnd 0.007322f
C2688 vdd.n1708 gnd 0.009097f
C2689 vdd.n1710 gnd 0.009097f
C2690 vdd.n1711 gnd 0.009097f
C2691 vdd.n1713 gnd 0.009097f
C2692 vdd.n1714 gnd 0.007322f
C2693 vdd.n1715 gnd 0.005822f
C2694 vdd.n1716 gnd 0.006186f
C2695 vdd.n1717 gnd 0.006186f
C2696 vdd.n1718 gnd 0.006186f
C2697 vdd.n1719 gnd 0.006186f
C2698 vdd.n1720 gnd 0.006186f
C2699 vdd.n1721 gnd 0.006186f
C2700 vdd.n1722 gnd 0.006186f
C2701 vdd.n1723 gnd 0.006186f
C2702 vdd.n1725 gnd 0.006186f
C2703 vdd.n1726 gnd 0.006186f
C2704 vdd.n1727 gnd 0.006186f
C2705 vdd.n1728 gnd 0.006186f
C2706 vdd.n1729 gnd 0.006186f
C2707 vdd.n1731 gnd 0.006186f
C2708 vdd.n1733 gnd 0.006186f
C2709 vdd.n1734 gnd 0.006186f
C2710 vdd.n1735 gnd 0.006186f
C2711 vdd.n1736 gnd 0.006186f
C2712 vdd.n1737 gnd 0.006186f
C2713 vdd.n1739 gnd 0.006186f
C2714 vdd.n1741 gnd 0.006186f
C2715 vdd.n1742 gnd 0.006186f
C2716 vdd.n1743 gnd 0.006186f
C2717 vdd.n1744 gnd 0.006186f
C2718 vdd.n1745 gnd 0.006186f
C2719 vdd.n1747 gnd 0.006186f
C2720 vdd.n1749 gnd 0.006186f
C2721 vdd.n1750 gnd 0.006186f
C2722 vdd.n1751 gnd 0.006186f
C2723 vdd.n1752 gnd 0.006186f
C2724 vdd.n1753 gnd 0.006186f
C2725 vdd.n1755 gnd 0.006186f
C2726 vdd.n1756 gnd 0.006186f
C2727 vdd.n1757 gnd 0.006186f
C2728 vdd.n1758 gnd 0.006186f
C2729 vdd.n1759 gnd 0.006186f
C2730 vdd.n1760 gnd 0.006186f
C2731 vdd.n1761 gnd 0.006186f
C2732 vdd.n1762 gnd 0.006186f
C2733 vdd.n1763 gnd 0.004503f
C2734 vdd.n1764 gnd 0.006186f
C2735 vdd.t115 gnd 0.249964f
C2736 vdd.t116 gnd 0.255869f
C2737 vdd.t114 gnd 0.163186f
C2738 vdd.n1765 gnd 0.088193f
C2739 vdd.n1766 gnd 0.050026f
C2740 vdd.n1767 gnd 0.00884f
C2741 vdd.n1768 gnd 0.006186f
C2742 vdd.n1769 gnd 0.006186f
C2743 vdd.n1770 gnd 0.376502f
C2744 vdd.n1771 gnd 0.006186f
C2745 vdd.n1772 gnd 0.006186f
C2746 vdd.n1773 gnd 0.006186f
C2747 vdd.n1774 gnd 0.006186f
C2748 vdd.n1775 gnd 0.006186f
C2749 vdd.n1776 gnd 0.006186f
C2750 vdd.n1777 gnd 0.006186f
C2751 vdd.n1778 gnd 0.006186f
C2752 vdd.n1779 gnd 0.006186f
C2753 vdd.n1780 gnd 0.006186f
C2754 vdd.n1781 gnd 0.006186f
C2755 vdd.n1782 gnd 0.006186f
C2756 vdd.n1783 gnd 0.006186f
C2757 vdd.n1784 gnd 0.006186f
C2758 vdd.n1785 gnd 0.006186f
C2759 vdd.n1786 gnd 0.006186f
C2760 vdd.n1787 gnd 0.006186f
C2761 vdd.n1788 gnd 0.006186f
C2762 vdd.n1789 gnd 0.006186f
C2763 vdd.n1790 gnd 0.006186f
C2764 vdd.t90 gnd 0.249964f
C2765 vdd.t91 gnd 0.255869f
C2766 vdd.t88 gnd 0.163186f
C2767 vdd.n1791 gnd 0.088193f
C2768 vdd.n1792 gnd 0.050026f
C2769 vdd.n1793 gnd 0.006186f
C2770 vdd.n1794 gnd 0.006186f
C2771 vdd.n1795 gnd 0.006186f
C2772 vdd.n1796 gnd 0.006186f
C2773 vdd.n1797 gnd 0.006186f
C2774 vdd.n1798 gnd 0.006186f
C2775 vdd.n1800 gnd 0.006186f
C2776 vdd.n1801 gnd 0.006186f
C2777 vdd.n1802 gnd 0.006186f
C2778 vdd.n1803 gnd 0.006186f
C2779 vdd.n1805 gnd 0.006186f
C2780 vdd.n1807 gnd 0.006186f
C2781 vdd.n1808 gnd 0.006186f
C2782 vdd.n1809 gnd 0.006186f
C2783 vdd.n1810 gnd 0.006186f
C2784 vdd.n1811 gnd 0.006186f
C2785 vdd.n1813 gnd 0.006186f
C2786 vdd.n1815 gnd 0.006186f
C2787 vdd.n1816 gnd 0.006186f
C2788 vdd.n1817 gnd 0.006186f
C2789 vdd.n1818 gnd 0.006186f
C2790 vdd.n1819 gnd 0.006186f
C2791 vdd.n1821 gnd 0.006186f
C2792 vdd.n1823 gnd 0.006186f
C2793 vdd.n1824 gnd 0.006186f
C2794 vdd.n1825 gnd 0.004503f
C2795 vdd.n1826 gnd 0.00884f
C2796 vdd.n1827 gnd 0.004776f
C2797 vdd.n1828 gnd 0.006186f
C2798 vdd.n1830 gnd 0.006186f
C2799 vdd.n1831 gnd 0.014678f
C2800 vdd.n1832 gnd 0.014678f
C2801 vdd.n1833 gnd 0.013704f
C2802 vdd.n1834 gnd 0.006186f
C2803 vdd.n1835 gnd 0.006186f
C2804 vdd.n1836 gnd 0.006186f
C2805 vdd.n1837 gnd 0.006186f
C2806 vdd.n1838 gnd 0.006186f
C2807 vdd.n1839 gnd 0.006186f
C2808 vdd.n1840 gnd 0.006186f
C2809 vdd.n1841 gnd 0.006186f
C2810 vdd.n1842 gnd 0.006186f
C2811 vdd.n1843 gnd 0.006186f
C2812 vdd.n1844 gnd 0.006186f
C2813 vdd.n1845 gnd 0.006186f
C2814 vdd.n1846 gnd 0.006186f
C2815 vdd.n1847 gnd 0.006186f
C2816 vdd.n1848 gnd 0.006186f
C2817 vdd.n1849 gnd 0.006186f
C2818 vdd.n1850 gnd 0.006186f
C2819 vdd.n1851 gnd 0.006186f
C2820 vdd.n1852 gnd 0.006186f
C2821 vdd.n1853 gnd 0.006186f
C2822 vdd.n1854 gnd 0.006186f
C2823 vdd.n1855 gnd 0.006186f
C2824 vdd.n1856 gnd 0.006186f
C2825 vdd.n1857 gnd 0.006186f
C2826 vdd.n1858 gnd 0.006186f
C2827 vdd.n1859 gnd 0.006186f
C2828 vdd.n1860 gnd 0.006186f
C2829 vdd.n1861 gnd 0.006186f
C2830 vdd.n1862 gnd 0.006186f
C2831 vdd.n1863 gnd 0.006186f
C2832 vdd.n1864 gnd 0.006186f
C2833 vdd.n1865 gnd 0.006186f
C2834 vdd.n1866 gnd 0.006186f
C2835 vdd.n1867 gnd 0.006186f
C2836 vdd.n1868 gnd 0.006186f
C2837 vdd.n1869 gnd 0.006186f
C2838 vdd.n1870 gnd 0.006186f
C2839 vdd.n1871 gnd 0.199871f
C2840 vdd.n1872 gnd 0.006186f
C2841 vdd.n1873 gnd 0.006186f
C2842 vdd.n1874 gnd 0.006186f
C2843 vdd.n1875 gnd 0.006186f
C2844 vdd.n1876 gnd 0.006186f
C2845 vdd.n1877 gnd 0.006186f
C2846 vdd.n1878 gnd 0.006186f
C2847 vdd.n1879 gnd 0.006186f
C2848 vdd.n1880 gnd 0.006186f
C2849 vdd.n1881 gnd 0.006186f
C2850 vdd.n1882 gnd 0.006186f
C2851 vdd.n1883 gnd 0.006186f
C2852 vdd.n1884 gnd 0.006186f
C2853 vdd.n1885 gnd 0.006186f
C2854 vdd.n1886 gnd 0.006186f
C2855 vdd.n1887 gnd 0.006186f
C2856 vdd.n1888 gnd 0.006186f
C2857 vdd.n1889 gnd 0.006186f
C2858 vdd.n1890 gnd 0.006186f
C2859 vdd.n1891 gnd 0.006186f
C2860 vdd.n1892 gnd 0.013704f
C2861 vdd.n1894 gnd 0.014678f
C2862 vdd.n1895 gnd 0.014678f
C2863 vdd.n1896 gnd 0.006186f
C2864 vdd.n1897 gnd 0.004776f
C2865 vdd.n1898 gnd 0.006186f
C2866 vdd.n1900 gnd 0.006186f
C2867 vdd.n1902 gnd 0.006186f
C2868 vdd.n1903 gnd 0.006186f
C2869 vdd.n1904 gnd 0.006186f
C2870 vdd.n1905 gnd 0.006186f
C2871 vdd.n1906 gnd 0.006186f
C2872 vdd.n1908 gnd 0.006186f
C2873 vdd.n1910 gnd 0.006186f
C2874 vdd.n1911 gnd 0.006186f
C2875 vdd.n1912 gnd 0.006186f
C2876 vdd.n1913 gnd 0.006186f
C2877 vdd.n1914 gnd 0.006186f
C2878 vdd.n1916 gnd 0.006186f
C2879 vdd.n1918 gnd 0.006186f
C2880 vdd.n1919 gnd 0.006186f
C2881 vdd.n1920 gnd 0.006186f
C2882 vdd.n1921 gnd 0.006186f
C2883 vdd.n1922 gnd 0.006186f
C2884 vdd.n1924 gnd 0.006186f
C2885 vdd.n1926 gnd 0.006186f
C2886 vdd.n1927 gnd 0.006186f
C2887 vdd.n1928 gnd 0.018451f
C2888 vdd.n1929 gnd 0.546958f
C2889 vdd.n1931 gnd 0.007322f
C2890 vdd.n1932 gnd 0.007322f
C2891 vdd.n1933 gnd 0.009097f
C2892 vdd.n1935 gnd 0.009097f
C2893 vdd.n1936 gnd 0.009097f
C2894 vdd.n1937 gnd 0.007322f
C2895 vdd.n1938 gnd 0.006077f
C2896 vdd.n1939 gnd 0.022678f
C2897 vdd.n1940 gnd 0.022169f
C2898 vdd.n1941 gnd 0.006077f
C2899 vdd.n1942 gnd 0.022169f
C2900 vdd.n1943 gnd 1.27825f
C2901 vdd.n1944 gnd 0.022169f
C2902 vdd.n1945 gnd 0.022678f
C2903 vdd.n1946 gnd 0.003478f
C2904 vdd.t51 gnd 0.111913f
C2905 vdd.t50 gnd 0.119604f
C2906 vdd.t48 gnd 0.146157f
C2907 vdd.n1947 gnd 0.187352f
C2908 vdd.n1948 gnd 0.15741f
C2909 vdd.n1949 gnd 0.011275f
C2910 vdd.n1950 gnd 0.003844f
C2911 vdd.n1951 gnd 0.007823f
C2912 vdd.n1952 gnd 0.546958f
C2913 vdd.n1953 gnd 0.018451f
C2914 vdd.n1954 gnd 0.006186f
C2915 vdd.n1955 gnd 0.006186f
C2916 vdd.n1956 gnd 0.006186f
C2917 vdd.n1958 gnd 0.006186f
C2918 vdd.n1960 gnd 0.006186f
C2919 vdd.n1961 gnd 0.006186f
C2920 vdd.n1962 gnd 0.006186f
C2921 vdd.n1963 gnd 0.006186f
C2922 vdd.n1964 gnd 0.006186f
C2923 vdd.n1966 gnd 0.006186f
C2924 vdd.n1968 gnd 0.006186f
C2925 vdd.n1969 gnd 0.006186f
C2926 vdd.n1970 gnd 0.006186f
C2927 vdd.n1971 gnd 0.006186f
C2928 vdd.n1972 gnd 0.006186f
C2929 vdd.n1974 gnd 0.006186f
C2930 vdd.n1976 gnd 0.006186f
C2931 vdd.n1977 gnd 0.006186f
C2932 vdd.n1978 gnd 0.006186f
C2933 vdd.n1979 gnd 0.006186f
C2934 vdd.n1980 gnd 0.006186f
C2935 vdd.n1982 gnd 0.006186f
C2936 vdd.n1984 gnd 0.006186f
C2937 vdd.n1985 gnd 0.006186f
C2938 vdd.n1986 gnd 0.014678f
C2939 vdd.n1987 gnd 0.013704f
C2940 vdd.n1988 gnd 0.013704f
C2941 vdd.n1989 gnd 0.911042f
C2942 vdd.n1990 gnd 0.013704f
C2943 vdd.n1991 gnd 0.013704f
C2944 vdd.n1992 gnd 0.006186f
C2945 vdd.n1993 gnd 0.006186f
C2946 vdd.n1994 gnd 0.006186f
C2947 vdd.n1995 gnd 0.395095f
C2948 vdd.n1996 gnd 0.006186f
C2949 vdd.n1997 gnd 0.006186f
C2950 vdd.n1998 gnd 0.006186f
C2951 vdd.n1999 gnd 0.006186f
C2952 vdd.n2000 gnd 0.006186f
C2953 vdd.n2001 gnd 0.632151f
C2954 vdd.n2002 gnd 0.006186f
C2955 vdd.n2003 gnd 0.006186f
C2956 vdd.n2004 gnd 0.006186f
C2957 vdd.n2005 gnd 0.006186f
C2958 vdd.n2006 gnd 0.006186f
C2959 vdd.n2007 gnd 0.632151f
C2960 vdd.n2008 gnd 0.006186f
C2961 vdd.n2009 gnd 0.006186f
C2962 vdd.n2010 gnd 0.005458f
C2963 vdd.n2011 gnd 0.017919f
C2964 vdd.n2012 gnd 0.003821f
C2965 vdd.n2013 gnd 0.006186f
C2966 vdd.n2014 gnd 0.348613f
C2967 vdd.n2015 gnd 0.006186f
C2968 vdd.n2016 gnd 0.006186f
C2969 vdd.n2017 gnd 0.006186f
C2970 vdd.n2018 gnd 0.006186f
C2971 vdd.n2019 gnd 0.006186f
C2972 vdd.n2020 gnd 0.422984f
C2973 vdd.n2021 gnd 0.006186f
C2974 vdd.n2022 gnd 0.006186f
C2975 vdd.n2023 gnd 0.006186f
C2976 vdd.n2024 gnd 0.006186f
C2977 vdd.n2025 gnd 0.006186f
C2978 vdd.n2026 gnd 0.562429f
C2979 vdd.n2027 gnd 0.006186f
C2980 vdd.n2028 gnd 0.006186f
C2981 vdd.n2029 gnd 0.006186f
C2982 vdd.n2030 gnd 0.006186f
C2983 vdd.n2031 gnd 0.006186f
C2984 vdd.n2032 gnd 0.502003f
C2985 vdd.n2033 gnd 0.006186f
C2986 vdd.n2034 gnd 0.006186f
C2987 vdd.n2035 gnd 0.006186f
C2988 vdd.n2036 gnd 0.006186f
C2989 vdd.n2037 gnd 0.006186f
C2990 vdd.n2038 gnd 0.362557f
C2991 vdd.n2039 gnd 0.006186f
C2992 vdd.n2040 gnd 0.006186f
C2993 vdd.n2041 gnd 0.006186f
C2994 vdd.n2042 gnd 0.006186f
C2995 vdd.n2043 gnd 0.006186f
C2996 vdd.n2044 gnd 0.199871f
C2997 vdd.n2045 gnd 0.006186f
C2998 vdd.n2046 gnd 0.006186f
C2999 vdd.n2047 gnd 0.006186f
C3000 vdd.n2048 gnd 0.006186f
C3001 vdd.n2049 gnd 0.006186f
C3002 vdd.n2050 gnd 0.348613f
C3003 vdd.n2051 gnd 0.006186f
C3004 vdd.n2052 gnd 0.006186f
C3005 vdd.n2053 gnd 0.006186f
C3006 vdd.n2054 gnd 0.006186f
C3007 vdd.n2055 gnd 0.006186f
C3008 vdd.n2056 gnd 0.632151f
C3009 vdd.n2057 gnd 0.006186f
C3010 vdd.n2058 gnd 0.006186f
C3011 vdd.n2059 gnd 0.006186f
C3012 vdd.n2060 gnd 0.006186f
C3013 vdd.n2061 gnd 0.006186f
C3014 vdd.n2062 gnd 0.006186f
C3015 vdd.n2063 gnd 0.006186f
C3016 vdd.n2064 gnd 0.492706f
C3017 vdd.n2065 gnd 0.006186f
C3018 vdd.n2066 gnd 0.006186f
C3019 vdd.n2067 gnd 0.006186f
C3020 vdd.n2068 gnd 0.006186f
C3021 vdd.n2069 gnd 0.006186f
C3022 vdd.n2070 gnd 0.006186f
C3023 vdd.n2071 gnd 0.395095f
C3024 vdd.n2072 gnd 0.006186f
C3025 vdd.n2073 gnd 0.006186f
C3026 vdd.n2074 gnd 0.006186f
C3027 vdd.n2075 gnd 0.014457f
C3028 vdd.n2076 gnd 0.013924f
C3029 vdd.n2077 gnd 0.006186f
C3030 vdd.n2078 gnd 0.006186f
C3031 vdd.n2079 gnd 0.004776f
C3032 vdd.n2080 gnd 0.006186f
C3033 vdd.n2081 gnd 0.006186f
C3034 vdd.n2082 gnd 0.004503f
C3035 vdd.n2083 gnd 0.006186f
C3036 vdd.n2084 gnd 0.006186f
C3037 vdd.n2085 gnd 0.006186f
C3038 vdd.n2086 gnd 0.006186f
C3039 vdd.n2087 gnd 0.006186f
C3040 vdd.n2088 gnd 0.006186f
C3041 vdd.n2089 gnd 0.006186f
C3042 vdd.n2090 gnd 0.006186f
C3043 vdd.n2091 gnd 0.006186f
C3044 vdd.n2092 gnd 0.006186f
C3045 vdd.n2093 gnd 0.006186f
C3046 vdd.n2094 gnd 0.006186f
C3047 vdd.n2095 gnd 0.006186f
C3048 vdd.n2096 gnd 0.006186f
C3049 vdd.n2097 gnd 0.006186f
C3050 vdd.n2098 gnd 0.006186f
C3051 vdd.n2099 gnd 0.006186f
C3052 vdd.n2100 gnd 0.006186f
C3053 vdd.n2101 gnd 0.006186f
C3054 vdd.n2102 gnd 0.006186f
C3055 vdd.n2103 gnd 0.006186f
C3056 vdd.n2104 gnd 0.006186f
C3057 vdd.n2105 gnd 0.006186f
C3058 vdd.n2106 gnd 0.006186f
C3059 vdd.n2107 gnd 0.006186f
C3060 vdd.n2108 gnd 0.006186f
C3061 vdd.n2109 gnd 0.006186f
C3062 vdd.n2110 gnd 0.006186f
C3063 vdd.n2111 gnd 0.006186f
C3064 vdd.n2112 gnd 0.006186f
C3065 vdd.n2113 gnd 0.006186f
C3066 vdd.n2114 gnd 0.006186f
C3067 vdd.n2115 gnd 0.006186f
C3068 vdd.n2116 gnd 0.006186f
C3069 vdd.n2117 gnd 0.006186f
C3070 vdd.n2118 gnd 0.006186f
C3071 vdd.n2119 gnd 0.006186f
C3072 vdd.n2120 gnd 0.006186f
C3073 vdd.n2121 gnd 0.006186f
C3074 vdd.n2122 gnd 0.006186f
C3075 vdd.n2123 gnd 0.006186f
C3076 vdd.n2124 gnd 0.006186f
C3077 vdd.n2125 gnd 0.006186f
C3078 vdd.n2126 gnd 0.006186f
C3079 vdd.n2127 gnd 0.006186f
C3080 vdd.n2128 gnd 0.006186f
C3081 vdd.n2129 gnd 0.006186f
C3082 vdd.n2130 gnd 0.006186f
C3083 vdd.n2131 gnd 0.006186f
C3084 vdd.n2132 gnd 0.006186f
C3085 vdd.n2133 gnd 0.006186f
C3086 vdd.n2134 gnd 0.006186f
C3087 vdd.n2135 gnd 0.006186f
C3088 vdd.n2136 gnd 0.006186f
C3089 vdd.n2137 gnd 0.006186f
C3090 vdd.n2138 gnd 0.006186f
C3091 vdd.n2139 gnd 0.006186f
C3092 vdd.n2140 gnd 0.006186f
C3093 vdd.n2141 gnd 0.006186f
C3094 vdd.n2142 gnd 0.006186f
C3095 vdd.n2143 gnd 0.014678f
C3096 vdd.n2144 gnd 0.013704f
C3097 vdd.n2145 gnd 0.013704f
C3098 vdd.n2146 gnd 0.771597f
C3099 vdd.n2147 gnd 0.013704f
C3100 vdd.n2148 gnd 0.014678f
C3101 vdd.n2149 gnd 0.013924f
C3102 vdd.n2150 gnd 0.006186f
C3103 vdd.n2151 gnd 0.006186f
C3104 vdd.n2152 gnd 0.006186f
C3105 vdd.n2153 gnd 0.004776f
C3106 vdd.n2154 gnd 0.00884f
C3107 vdd.n2155 gnd 0.004503f
C3108 vdd.n2156 gnd 0.006186f
C3109 vdd.n2157 gnd 0.006186f
C3110 vdd.n2158 gnd 0.006186f
C3111 vdd.n2159 gnd 0.006186f
C3112 vdd.n2160 gnd 0.006186f
C3113 vdd.n2161 gnd 0.006186f
C3114 vdd.n2162 gnd 0.006186f
C3115 vdd.n2163 gnd 0.006186f
C3116 vdd.n2164 gnd 0.006186f
C3117 vdd.n2165 gnd 0.006186f
C3118 vdd.n2166 gnd 0.006186f
C3119 vdd.n2167 gnd 0.006186f
C3120 vdd.n2168 gnd 0.006186f
C3121 vdd.n2169 gnd 0.006186f
C3122 vdd.n2170 gnd 0.006186f
C3123 vdd.n2171 gnd 0.006186f
C3124 vdd.n2172 gnd 0.006186f
C3125 vdd.n2173 gnd 0.006186f
C3126 vdd.n2174 gnd 0.006186f
C3127 vdd.n2175 gnd 0.006186f
C3128 vdd.n2176 gnd 0.006186f
C3129 vdd.n2177 gnd 0.006186f
C3130 vdd.n2178 gnd 0.006186f
C3131 vdd.n2179 gnd 0.006186f
C3132 vdd.n2180 gnd 0.006186f
C3133 vdd.n2181 gnd 0.006186f
C3134 vdd.n2182 gnd 0.006186f
C3135 vdd.n2183 gnd 0.006186f
C3136 vdd.n2184 gnd 0.006186f
C3137 vdd.n2185 gnd 0.006186f
C3138 vdd.n2186 gnd 0.006186f
C3139 vdd.n2187 gnd 0.006186f
C3140 vdd.n2188 gnd 0.006186f
C3141 vdd.n2189 gnd 0.006186f
C3142 vdd.n2190 gnd 0.006186f
C3143 vdd.n2191 gnd 0.006186f
C3144 vdd.n2192 gnd 0.006186f
C3145 vdd.n2193 gnd 0.006186f
C3146 vdd.n2194 gnd 0.006186f
C3147 vdd.n2195 gnd 0.006186f
C3148 vdd.n2196 gnd 0.006186f
C3149 vdd.n2197 gnd 0.006186f
C3150 vdd.n2198 gnd 0.006186f
C3151 vdd.n2199 gnd 0.006186f
C3152 vdd.n2200 gnd 0.006186f
C3153 vdd.n2201 gnd 0.006186f
C3154 vdd.n2202 gnd 0.006186f
C3155 vdd.n2203 gnd 0.006186f
C3156 vdd.n2204 gnd 0.006186f
C3157 vdd.n2205 gnd 0.006186f
C3158 vdd.n2206 gnd 0.006186f
C3159 vdd.n2207 gnd 0.006186f
C3160 vdd.n2208 gnd 0.006186f
C3161 vdd.n2209 gnd 0.006186f
C3162 vdd.n2210 gnd 0.006186f
C3163 vdd.n2211 gnd 0.006186f
C3164 vdd.n2212 gnd 0.006186f
C3165 vdd.n2213 gnd 0.006186f
C3166 vdd.n2214 gnd 0.006186f
C3167 vdd.n2215 gnd 0.006186f
C3168 vdd.n2216 gnd 0.014678f
C3169 vdd.n2217 gnd 0.014678f
C3170 vdd.n2218 gnd 0.771597f
C3171 vdd.t36 gnd 2.74242f
C3172 vdd.t38 gnd 2.74242f
C3173 vdd.n2251 gnd 0.014678f
C3174 vdd.n2252 gnd 0.006186f
C3175 vdd.t83 gnd 0.249964f
C3176 vdd.t84 gnd 0.255869f
C3177 vdd.t81 gnd 0.163186f
C3178 vdd.n2253 gnd 0.088193f
C3179 vdd.n2254 gnd 0.050026f
C3180 vdd.n2255 gnd 0.006186f
C3181 vdd.t97 gnd 0.249964f
C3182 vdd.t98 gnd 0.255869f
C3183 vdd.t96 gnd 0.163186f
C3184 vdd.n2256 gnd 0.088193f
C3185 vdd.n2257 gnd 0.050026f
C3186 vdd.n2258 gnd 0.00884f
C3187 vdd.n2259 gnd 0.006186f
C3188 vdd.n2260 gnd 0.006186f
C3189 vdd.n2261 gnd 0.006186f
C3190 vdd.n2262 gnd 0.006186f
C3191 vdd.n2263 gnd 0.006186f
C3192 vdd.n2264 gnd 0.006186f
C3193 vdd.n2265 gnd 0.006186f
C3194 vdd.n2266 gnd 0.006186f
C3195 vdd.n2267 gnd 0.006186f
C3196 vdd.n2268 gnd 0.006186f
C3197 vdd.n2269 gnd 0.006186f
C3198 vdd.n2270 gnd 0.006186f
C3199 vdd.n2271 gnd 0.006186f
C3200 vdd.n2272 gnd 0.006186f
C3201 vdd.n2273 gnd 0.006186f
C3202 vdd.n2274 gnd 0.006186f
C3203 vdd.n2275 gnd 0.006186f
C3204 vdd.n2276 gnd 0.006186f
C3205 vdd.n2277 gnd 0.006186f
C3206 vdd.n2278 gnd 0.006186f
C3207 vdd.n2279 gnd 0.006186f
C3208 vdd.n2280 gnd 0.006186f
C3209 vdd.n2281 gnd 0.006186f
C3210 vdd.n2282 gnd 0.006186f
C3211 vdd.n2283 gnd 0.006186f
C3212 vdd.n2284 gnd 0.006186f
C3213 vdd.n2285 gnd 0.006186f
C3214 vdd.n2286 gnd 0.006186f
C3215 vdd.n2287 gnd 0.006186f
C3216 vdd.n2288 gnd 0.006186f
C3217 vdd.n2289 gnd 0.006186f
C3218 vdd.n2290 gnd 0.006186f
C3219 vdd.n2291 gnd 0.006186f
C3220 vdd.n2292 gnd 0.006186f
C3221 vdd.n2293 gnd 0.006186f
C3222 vdd.n2294 gnd 0.006186f
C3223 vdd.n2295 gnd 0.006186f
C3224 vdd.n2296 gnd 0.006186f
C3225 vdd.n2297 gnd 0.006186f
C3226 vdd.n2298 gnd 0.006186f
C3227 vdd.n2299 gnd 0.006186f
C3228 vdd.n2300 gnd 0.006186f
C3229 vdd.n2301 gnd 0.006186f
C3230 vdd.n2302 gnd 0.006186f
C3231 vdd.n2303 gnd 0.006186f
C3232 vdd.n2304 gnd 0.006186f
C3233 vdd.n2305 gnd 0.006186f
C3234 vdd.n2306 gnd 0.006186f
C3235 vdd.n2307 gnd 0.006186f
C3236 vdd.n2308 gnd 0.006186f
C3237 vdd.n2309 gnd 0.006186f
C3238 vdd.n2310 gnd 0.006186f
C3239 vdd.n2311 gnd 0.006186f
C3240 vdd.n2312 gnd 0.006186f
C3241 vdd.n2313 gnd 0.006186f
C3242 vdd.n2314 gnd 0.006186f
C3243 vdd.n2315 gnd 0.004503f
C3244 vdd.n2316 gnd 0.006186f
C3245 vdd.n2317 gnd 0.006186f
C3246 vdd.n2318 gnd 0.004776f
C3247 vdd.n2319 gnd 0.006186f
C3248 vdd.n2320 gnd 0.006186f
C3249 vdd.n2321 gnd 0.014678f
C3250 vdd.n2322 gnd 0.013704f
C3251 vdd.n2323 gnd 0.006186f
C3252 vdd.n2324 gnd 0.006186f
C3253 vdd.n2325 gnd 0.006186f
C3254 vdd.n2326 gnd 0.006186f
C3255 vdd.n2327 gnd 0.006186f
C3256 vdd.n2328 gnd 0.006186f
C3257 vdd.n2329 gnd 0.006186f
C3258 vdd.n2330 gnd 0.006186f
C3259 vdd.n2331 gnd 0.006186f
C3260 vdd.n2332 gnd 0.006186f
C3261 vdd.n2333 gnd 0.006186f
C3262 vdd.n2334 gnd 0.006186f
C3263 vdd.n2335 gnd 0.006186f
C3264 vdd.n2336 gnd 0.006186f
C3265 vdd.n2337 gnd 0.006186f
C3266 vdd.n2338 gnd 0.006186f
C3267 vdd.n2339 gnd 0.006186f
C3268 vdd.n2340 gnd 0.006186f
C3269 vdd.n2341 gnd 0.006186f
C3270 vdd.n2342 gnd 0.006186f
C3271 vdd.n2343 gnd 0.006186f
C3272 vdd.n2344 gnd 0.006186f
C3273 vdd.n2345 gnd 0.006186f
C3274 vdd.n2346 gnd 0.006186f
C3275 vdd.n2347 gnd 0.006186f
C3276 vdd.n2348 gnd 0.006186f
C3277 vdd.n2349 gnd 0.006186f
C3278 vdd.n2350 gnd 0.006186f
C3279 vdd.n2351 gnd 0.006186f
C3280 vdd.n2352 gnd 0.006186f
C3281 vdd.n2353 gnd 0.006186f
C3282 vdd.n2354 gnd 0.006186f
C3283 vdd.n2355 gnd 0.006186f
C3284 vdd.n2356 gnd 0.006186f
C3285 vdd.n2357 gnd 0.006186f
C3286 vdd.n2358 gnd 0.006186f
C3287 vdd.n2359 gnd 0.006186f
C3288 vdd.n2360 gnd 0.006186f
C3289 vdd.n2361 gnd 0.006186f
C3290 vdd.n2362 gnd 0.006186f
C3291 vdd.n2363 gnd 0.006186f
C3292 vdd.n2364 gnd 0.006186f
C3293 vdd.n2365 gnd 0.006186f
C3294 vdd.n2366 gnd 0.006186f
C3295 vdd.n2367 gnd 0.006186f
C3296 vdd.n2368 gnd 0.006186f
C3297 vdd.n2369 gnd 0.006186f
C3298 vdd.n2370 gnd 0.006186f
C3299 vdd.n2371 gnd 0.006186f
C3300 vdd.n2372 gnd 0.006186f
C3301 vdd.n2373 gnd 0.006186f
C3302 vdd.n2374 gnd 0.199871f
C3303 vdd.n2375 gnd 0.006186f
C3304 vdd.n2376 gnd 0.006186f
C3305 vdd.n2377 gnd 0.006186f
C3306 vdd.n2378 gnd 0.006186f
C3307 vdd.n2379 gnd 0.006186f
C3308 vdd.n2380 gnd 0.006186f
C3309 vdd.n2381 gnd 0.006186f
C3310 vdd.n2382 gnd 0.006186f
C3311 vdd.n2383 gnd 0.006186f
C3312 vdd.n2384 gnd 0.006186f
C3313 vdd.n2385 gnd 0.006186f
C3314 vdd.n2386 gnd 0.006186f
C3315 vdd.n2387 gnd 0.006186f
C3316 vdd.n2388 gnd 0.006186f
C3317 vdd.n2389 gnd 0.006186f
C3318 vdd.n2390 gnd 0.006186f
C3319 vdd.n2391 gnd 0.006186f
C3320 vdd.n2392 gnd 0.006186f
C3321 vdd.n2393 gnd 0.006186f
C3322 vdd.n2394 gnd 0.006186f
C3323 vdd.n2395 gnd 0.376502f
C3324 vdd.n2396 gnd 0.006186f
C3325 vdd.n2397 gnd 0.006186f
C3326 vdd.n2398 gnd 0.006186f
C3327 vdd.n2399 gnd 0.006186f
C3328 vdd.n2400 gnd 0.006186f
C3329 vdd.n2401 gnd 0.013704f
C3330 vdd.n2402 gnd 0.014678f
C3331 vdd.n2403 gnd 0.014678f
C3332 vdd.n2404 gnd 0.006186f
C3333 vdd.n2405 gnd 0.006186f
C3334 vdd.n2406 gnd 0.006186f
C3335 vdd.n2407 gnd 0.004776f
C3336 vdd.n2408 gnd 0.00884f
C3337 vdd.n2409 gnd 0.004503f
C3338 vdd.n2410 gnd 0.006186f
C3339 vdd.n2411 gnd 0.006186f
C3340 vdd.n2412 gnd 0.006186f
C3341 vdd.n2413 gnd 0.006186f
C3342 vdd.n2414 gnd 0.006186f
C3343 vdd.n2415 gnd 0.006186f
C3344 vdd.n2416 gnd 0.006186f
C3345 vdd.n2417 gnd 0.006186f
C3346 vdd.n2418 gnd 0.006186f
C3347 vdd.n2419 gnd 0.006186f
C3348 vdd.n2420 gnd 0.006186f
C3349 vdd.n2421 gnd 0.006186f
C3350 vdd.n2422 gnd 0.006186f
C3351 vdd.n2423 gnd 0.006186f
C3352 vdd.n2424 gnd 0.006186f
C3353 vdd.n2425 gnd 0.006186f
C3354 vdd.n2426 gnd 0.006186f
C3355 vdd.n2427 gnd 0.006186f
C3356 vdd.n2428 gnd 0.006186f
C3357 vdd.n2429 gnd 0.006186f
C3358 vdd.n2430 gnd 0.006186f
C3359 vdd.n2431 gnd 0.006186f
C3360 vdd.n2432 gnd 0.006186f
C3361 vdd.n2433 gnd 0.006186f
C3362 vdd.n2434 gnd 0.006186f
C3363 vdd.n2435 gnd 0.006186f
C3364 vdd.n2436 gnd 0.006186f
C3365 vdd.n2437 gnd 0.006186f
C3366 vdd.n2438 gnd 0.006186f
C3367 vdd.n2439 gnd 0.006186f
C3368 vdd.n2440 gnd 0.006186f
C3369 vdd.n2441 gnd 0.006186f
C3370 vdd.n2442 gnd 0.006186f
C3371 vdd.n2443 gnd 0.006186f
C3372 vdd.n2444 gnd 0.006186f
C3373 vdd.n2445 gnd 0.006186f
C3374 vdd.n2446 gnd 0.006186f
C3375 vdd.n2447 gnd 0.006186f
C3376 vdd.n2448 gnd 0.006186f
C3377 vdd.n2449 gnd 0.006186f
C3378 vdd.n2450 gnd 0.006186f
C3379 vdd.n2451 gnd 0.006186f
C3380 vdd.n2452 gnd 0.006186f
C3381 vdd.n2453 gnd 0.006186f
C3382 vdd.n2454 gnd 0.006186f
C3383 vdd.n2455 gnd 0.006186f
C3384 vdd.n2456 gnd 0.006186f
C3385 vdd.n2457 gnd 0.006186f
C3386 vdd.n2458 gnd 0.006186f
C3387 vdd.n2459 gnd 0.006186f
C3388 vdd.n2460 gnd 0.006186f
C3389 vdd.n2461 gnd 0.006186f
C3390 vdd.n2462 gnd 0.006186f
C3391 vdd.n2463 gnd 0.006186f
C3392 vdd.n2464 gnd 0.006186f
C3393 vdd.n2465 gnd 0.006186f
C3394 vdd.n2466 gnd 0.006186f
C3395 vdd.n2467 gnd 0.006186f
C3396 vdd.n2468 gnd 0.006186f
C3397 vdd.n2469 gnd 0.006186f
C3398 vdd.n2471 gnd 0.771597f
C3399 vdd.n2473 gnd 0.006186f
C3400 vdd.n2474 gnd 0.006186f
C3401 vdd.n2475 gnd 0.014678f
C3402 vdd.n2476 gnd 0.013704f
C3403 vdd.n2477 gnd 0.013704f
C3404 vdd.n2478 gnd 0.771597f
C3405 vdd.n2479 gnd 0.013704f
C3406 vdd.n2480 gnd 0.013704f
C3407 vdd.n2481 gnd 0.006186f
C3408 vdd.n2482 gnd 0.006186f
C3409 vdd.n2483 gnd 0.006186f
C3410 vdd.n2484 gnd 0.395095f
C3411 vdd.n2485 gnd 0.006186f
C3412 vdd.n2486 gnd 0.006186f
C3413 vdd.n2487 gnd 0.006186f
C3414 vdd.n2488 gnd 0.006186f
C3415 vdd.n2489 gnd 0.006186f
C3416 vdd.n2490 gnd 0.492706f
C3417 vdd.n2491 gnd 0.006186f
C3418 vdd.n2492 gnd 0.006186f
C3419 vdd.n2493 gnd 0.006186f
C3420 vdd.n2494 gnd 0.006186f
C3421 vdd.n2495 gnd 0.006186f
C3422 vdd.n2496 gnd 0.632151f
C3423 vdd.n2497 gnd 0.006186f
C3424 vdd.n2498 gnd 0.006186f
C3425 vdd.n2499 gnd 0.006186f
C3426 vdd.n2500 gnd 0.006186f
C3427 vdd.n2501 gnd 0.006186f
C3428 vdd.n2502 gnd 0.348613f
C3429 vdd.n2503 gnd 0.006186f
C3430 vdd.n2504 gnd 0.006186f
C3431 vdd.n2505 gnd 0.006186f
C3432 vdd.n2506 gnd 0.006186f
C3433 vdd.n2507 gnd 0.006186f
C3434 vdd.n2508 gnd 0.199871f
C3435 vdd.n2509 gnd 0.006186f
C3436 vdd.n2510 gnd 0.006186f
C3437 vdd.n2511 gnd 0.006186f
C3438 vdd.n2512 gnd 0.006186f
C3439 vdd.n2513 gnd 0.006186f
C3440 vdd.n2514 gnd 0.362557f
C3441 vdd.n2515 gnd 0.006186f
C3442 vdd.n2516 gnd 0.006186f
C3443 vdd.n2517 gnd 0.006186f
C3444 vdd.n2518 gnd 0.006186f
C3445 vdd.n2519 gnd 0.006186f
C3446 vdd.n2520 gnd 0.502003f
C3447 vdd.n2521 gnd 0.006186f
C3448 vdd.n2522 gnd 0.006186f
C3449 vdd.n2523 gnd 0.006186f
C3450 vdd.n2524 gnd 0.006186f
C3451 vdd.n2525 gnd 0.006186f
C3452 vdd.n2526 gnd 0.562429f
C3453 vdd.n2527 gnd 0.006186f
C3454 vdd.n2528 gnd 0.006186f
C3455 vdd.n2529 gnd 0.006186f
C3456 vdd.n2530 gnd 0.006186f
C3457 vdd.n2531 gnd 0.006186f
C3458 vdd.n2532 gnd 0.422984f
C3459 vdd.n2533 gnd 0.006186f
C3460 vdd.n2534 gnd 0.006186f
C3461 vdd.n2535 gnd 0.006186f
C3462 vdd.t58 gnd 0.255869f
C3463 vdd.t56 gnd 0.163186f
C3464 vdd.t59 gnd 0.255869f
C3465 vdd.n2536 gnd 0.143809f
C3466 vdd.n2537 gnd 0.017919f
C3467 vdd.n2538 gnd 0.003821f
C3468 vdd.n2539 gnd 0.006186f
C3469 vdd.n2540 gnd 0.348613f
C3470 vdd.n2541 gnd 0.006186f
C3471 vdd.n2542 gnd 0.006186f
C3472 vdd.n2543 gnd 0.006186f
C3473 vdd.n2544 gnd 0.006186f
C3474 vdd.n2545 gnd 0.006186f
C3475 vdd.n2546 gnd 0.632151f
C3476 vdd.n2547 gnd 0.006186f
C3477 vdd.n2548 gnd 0.006186f
C3478 vdd.n2549 gnd 0.006186f
C3479 vdd.n2550 gnd 0.006186f
C3480 vdd.n2551 gnd 0.006186f
C3481 vdd.n2552 gnd 0.006186f
C3482 vdd.n2554 gnd 0.006186f
C3483 vdd.n2555 gnd 0.006186f
C3484 vdd.n2557 gnd 0.006186f
C3485 vdd.n2558 gnd 0.006186f
C3486 vdd.n2561 gnd 0.006186f
C3487 vdd.n2562 gnd 0.006186f
C3488 vdd.n2563 gnd 0.006186f
C3489 vdd.n2564 gnd 0.006186f
C3490 vdd.n2566 gnd 0.006186f
C3491 vdd.n2567 gnd 0.006186f
C3492 vdd.n2568 gnd 0.006186f
C3493 vdd.n2569 gnd 0.006186f
C3494 vdd.n2570 gnd 0.006186f
C3495 vdd.n2571 gnd 0.006186f
C3496 vdd.n2573 gnd 0.006186f
C3497 vdd.n2574 gnd 0.006186f
C3498 vdd.n2575 gnd 0.006186f
C3499 vdd.n2576 gnd 0.006186f
C3500 vdd.n2577 gnd 0.006186f
C3501 vdd.n2578 gnd 0.006186f
C3502 vdd.n2580 gnd 0.006186f
C3503 vdd.n2581 gnd 0.006186f
C3504 vdd.n2582 gnd 0.006186f
C3505 vdd.n2583 gnd 0.006186f
C3506 vdd.n2584 gnd 0.006186f
C3507 vdd.n2585 gnd 0.006186f
C3508 vdd.n2587 gnd 0.006186f
C3509 vdd.n2588 gnd 0.014678f
C3510 vdd.n2589 gnd 0.014678f
C3511 vdd.n2590 gnd 0.013704f
C3512 vdd.n2591 gnd 0.006186f
C3513 vdd.n2592 gnd 0.006186f
C3514 vdd.n2593 gnd 0.006186f
C3515 vdd.n2594 gnd 0.006186f
C3516 vdd.n2595 gnd 0.006186f
C3517 vdd.n2596 gnd 0.006186f
C3518 vdd.n2597 gnd 0.632151f
C3519 vdd.n2598 gnd 0.006186f
C3520 vdd.n2599 gnd 0.006186f
C3521 vdd.n2600 gnd 0.006186f
C3522 vdd.n2601 gnd 0.006186f
C3523 vdd.n2602 gnd 0.006186f
C3524 vdd.n2603 gnd 0.395095f
C3525 vdd.n2604 gnd 0.006186f
C3526 vdd.n2605 gnd 0.006186f
C3527 vdd.n2606 gnd 0.006186f
C3528 vdd.n2607 gnd 0.014457f
C3529 vdd.n2608 gnd 0.013924f
C3530 vdd.n2609 gnd 0.014678f
C3531 vdd.n2611 gnd 0.006186f
C3532 vdd.n2612 gnd 0.006186f
C3533 vdd.n2613 gnd 0.004776f
C3534 vdd.n2614 gnd 0.00884f
C3535 vdd.n2615 gnd 0.004503f
C3536 vdd.n2616 gnd 0.006186f
C3537 vdd.n2617 gnd 0.006186f
C3538 vdd.n2619 gnd 0.006186f
C3539 vdd.n2620 gnd 0.006186f
C3540 vdd.n2621 gnd 0.006186f
C3541 vdd.n2622 gnd 0.006186f
C3542 vdd.n2623 gnd 0.006186f
C3543 vdd.n2624 gnd 0.006186f
C3544 vdd.n2626 gnd 0.006186f
C3545 vdd.n2627 gnd 0.006186f
C3546 vdd.n2628 gnd 0.006186f
C3547 vdd.n2629 gnd 0.006186f
C3548 vdd.n2630 gnd 0.006186f
C3549 vdd.n2631 gnd 0.006186f
C3550 vdd.n2633 gnd 0.006186f
C3551 vdd.n2634 gnd 0.006186f
C3552 vdd.n2635 gnd 0.006186f
C3553 vdd.n2636 gnd 0.006186f
C3554 vdd.n2637 gnd 0.006186f
C3555 vdd.n2638 gnd 0.006186f
C3556 vdd.n2640 gnd 0.006186f
C3557 vdd.n2641 gnd 0.006186f
C3558 vdd.n2642 gnd 0.006186f
C3559 vdd.n2644 gnd 0.006186f
C3560 vdd.n2645 gnd 0.006186f
C3561 vdd.n2646 gnd 0.006186f
C3562 vdd.n2647 gnd 0.006186f
C3563 vdd.n2648 gnd 0.006186f
C3564 vdd.n2649 gnd 0.006186f
C3565 vdd.n2651 gnd 0.006186f
C3566 vdd.n2652 gnd 0.006186f
C3567 vdd.n2653 gnd 0.006186f
C3568 vdd.n2654 gnd 0.006186f
C3569 vdd.n2655 gnd 0.006186f
C3570 vdd.n2656 gnd 0.006186f
C3571 vdd.n2658 gnd 0.006186f
C3572 vdd.n2659 gnd 0.006186f
C3573 vdd.n2660 gnd 0.006186f
C3574 vdd.n2661 gnd 0.006186f
C3575 vdd.n2662 gnd 0.006186f
C3576 vdd.n2663 gnd 0.006186f
C3577 vdd.n2665 gnd 0.006186f
C3578 vdd.n2666 gnd 0.006186f
C3579 vdd.n2668 gnd 0.006186f
C3580 vdd.n2669 gnd 0.006186f
C3581 vdd.n2670 gnd 0.014678f
C3582 vdd.n2671 gnd 0.013704f
C3583 vdd.n2672 gnd 0.013704f
C3584 vdd.n2673 gnd 0.911042f
C3585 vdd.n2674 gnd 0.013704f
C3586 vdd.n2675 gnd 0.014678f
C3587 vdd.n2676 gnd 0.013924f
C3588 vdd.n2677 gnd 0.006186f
C3589 vdd.n2678 gnd 0.004776f
C3590 vdd.n2679 gnd 0.006186f
C3591 vdd.n2681 gnd 0.006186f
C3592 vdd.n2682 gnd 0.006186f
C3593 vdd.n2683 gnd 0.006186f
C3594 vdd.n2684 gnd 0.006186f
C3595 vdd.n2685 gnd 0.006186f
C3596 vdd.n2686 gnd 0.006186f
C3597 vdd.n2688 gnd 0.006186f
C3598 vdd.n2689 gnd 0.006186f
C3599 vdd.n2690 gnd 0.006186f
C3600 vdd.n2691 gnd 0.006186f
C3601 vdd.n2692 gnd 0.006186f
C3602 vdd.n2693 gnd 0.006186f
C3603 vdd.n2695 gnd 0.006186f
C3604 vdd.n2696 gnd 0.006186f
C3605 vdd.n2697 gnd 0.006186f
C3606 vdd.n2698 gnd 0.006186f
C3607 vdd.n2699 gnd 0.006186f
C3608 vdd.n2700 gnd 0.006186f
C3609 vdd.n2702 gnd 0.006186f
C3610 vdd.n2703 gnd 0.006186f
C3611 vdd.n2705 gnd 0.006186f
C3612 vdd.n2706 gnd 0.014864f
C3613 vdd.n2707 gnd 0.550544f
C3614 vdd.n2708 gnd 0.007823f
C3615 vdd.n2709 gnd 0.022678f
C3616 vdd.n2710 gnd 0.003478f
C3617 vdd.t109 gnd 0.111913f
C3618 vdd.t110 gnd 0.119604f
C3619 vdd.t108 gnd 0.146157f
C3620 vdd.n2711 gnd 0.187352f
C3621 vdd.n2712 gnd 0.15741f
C3622 vdd.n2713 gnd 0.011275f
C3623 vdd.n2714 gnd 0.009097f
C3624 vdd.n2715 gnd 0.003844f
C3625 vdd.n2716 gnd 0.007322f
C3626 vdd.n2717 gnd 0.009097f
C3627 vdd.n2718 gnd 0.009097f
C3628 vdd.n2719 gnd 0.007322f
C3629 vdd.n2720 gnd 0.007322f
C3630 vdd.n2721 gnd 0.009097f
C3631 vdd.n2722 gnd 0.009097f
C3632 vdd.n2723 gnd 0.007322f
C3633 vdd.n2724 gnd 0.007322f
C3634 vdd.n2725 gnd 0.009097f
C3635 vdd.n2726 gnd 0.009097f
C3636 vdd.n2727 gnd 0.007322f
C3637 vdd.n2728 gnd 0.007322f
C3638 vdd.n2729 gnd 0.009097f
C3639 vdd.n2730 gnd 0.009097f
C3640 vdd.n2731 gnd 0.007322f
C3641 vdd.n2732 gnd 0.007322f
C3642 vdd.n2733 gnd 0.009097f
C3643 vdd.n2734 gnd 0.009097f
C3644 vdd.n2735 gnd 0.007322f
C3645 vdd.n2736 gnd 0.007322f
C3646 vdd.n2737 gnd 0.009097f
C3647 vdd.n2738 gnd 0.009097f
C3648 vdd.n2739 gnd 0.007322f
C3649 vdd.n2740 gnd 0.007322f
C3650 vdd.n2741 gnd 0.009097f
C3651 vdd.n2742 gnd 0.009097f
C3652 vdd.n2743 gnd 0.007322f
C3653 vdd.n2744 gnd 0.007322f
C3654 vdd.n2745 gnd 0.009097f
C3655 vdd.n2746 gnd 0.009097f
C3656 vdd.n2747 gnd 0.007322f
C3657 vdd.n2748 gnd 0.007322f
C3658 vdd.n2749 gnd 0.009097f
C3659 vdd.n2750 gnd 0.009097f
C3660 vdd.n2751 gnd 0.007322f
C3661 vdd.n2752 gnd 0.009097f
C3662 vdd.n2753 gnd 0.009097f
C3663 vdd.n2754 gnd 0.007322f
C3664 vdd.n2755 gnd 0.009097f
C3665 vdd.n2756 gnd 0.009097f
C3666 vdd.n2757 gnd 0.009097f
C3667 vdd.n2758 gnd 0.014936f
C3668 vdd.n2759 gnd 0.009097f
C3669 vdd.n2760 gnd 0.009097f
C3670 vdd.n2761 gnd 0.004979f
C3671 vdd.n2762 gnd 0.007322f
C3672 vdd.n2763 gnd 0.009097f
C3673 vdd.n2764 gnd 0.009097f
C3674 vdd.n2765 gnd 0.007322f
C3675 vdd.n2766 gnd 0.007322f
C3676 vdd.n2767 gnd 0.009097f
C3677 vdd.n2768 gnd 0.009097f
C3678 vdd.n2769 gnd 0.007322f
C3679 vdd.n2770 gnd 0.007322f
C3680 vdd.n2771 gnd 0.009097f
C3681 vdd.n2772 gnd 0.009097f
C3682 vdd.n2773 gnd 0.007322f
C3683 vdd.n2774 gnd 0.007322f
C3684 vdd.n2775 gnd 0.009097f
C3685 vdd.n2776 gnd 0.009097f
C3686 vdd.n2777 gnd 0.007322f
C3687 vdd.n2778 gnd 0.007322f
C3688 vdd.n2779 gnd 0.009097f
C3689 vdd.n2780 gnd 0.009097f
C3690 vdd.n2781 gnd 0.007322f
C3691 vdd.n2782 gnd 0.007322f
C3692 vdd.n2783 gnd 0.009097f
C3693 vdd.n2784 gnd 0.009097f
C3694 vdd.n2785 gnd 0.007322f
C3695 vdd.n2786 gnd 0.007322f
C3696 vdd.n2787 gnd 0.009097f
C3697 vdd.n2788 gnd 0.009097f
C3698 vdd.n2789 gnd 0.007322f
C3699 vdd.n2790 gnd 0.007322f
C3700 vdd.n2791 gnd 0.009097f
C3701 vdd.n2792 gnd 0.009097f
C3702 vdd.n2793 gnd 0.007322f
C3703 vdd.n2794 gnd 0.007322f
C3704 vdd.n2795 gnd 0.009097f
C3705 vdd.n2796 gnd 0.009097f
C3706 vdd.n2797 gnd 0.007322f
C3707 vdd.n2798 gnd 0.009097f
C3708 vdd.n2799 gnd 0.009097f
C3709 vdd.n2800 gnd 0.007322f
C3710 vdd.n2801 gnd 0.009097f
C3711 vdd.n2802 gnd 0.009097f
C3712 vdd.n2803 gnd 0.009097f
C3713 vdd.t46 gnd 0.111913f
C3714 vdd.t47 gnd 0.119604f
C3715 vdd.t45 gnd 0.146157f
C3716 vdd.n2804 gnd 0.187352f
C3717 vdd.n2805 gnd 0.15741f
C3718 vdd.n2806 gnd 0.014936f
C3719 vdd.n2807 gnd 0.009097f
C3720 vdd.n2808 gnd 0.009097f
C3721 vdd.n2809 gnd 0.006114f
C3722 vdd.n2810 gnd 0.007322f
C3723 vdd.n2811 gnd 0.009097f
C3724 vdd.n2812 gnd 0.009097f
C3725 vdd.n2813 gnd 0.007322f
C3726 vdd.n2814 gnd 0.007322f
C3727 vdd.n2815 gnd 0.009097f
C3728 vdd.n2816 gnd 0.009097f
C3729 vdd.n2817 gnd 0.007322f
C3730 vdd.n2818 gnd 0.007322f
C3731 vdd.n2819 gnd 0.009097f
C3732 vdd.n2820 gnd 0.009097f
C3733 vdd.n2821 gnd 0.007322f
C3734 vdd.n2822 gnd 0.007322f
C3735 vdd.n2823 gnd 0.009097f
C3736 vdd.n2824 gnd 0.009097f
C3737 vdd.n2825 gnd 0.007322f
C3738 vdd.n2826 gnd 0.007322f
C3739 vdd.n2827 gnd 0.009097f
C3740 vdd.n2828 gnd 0.009097f
C3741 vdd.n2829 gnd 0.007322f
C3742 vdd.n2830 gnd 0.007322f
C3743 vdd.n2831 gnd 0.009097f
C3744 vdd.n2832 gnd 0.009097f
C3745 vdd.n2833 gnd 0.007322f
C3746 vdd.n2834 gnd 0.007322f
C3747 vdd.n2836 gnd 0.550544f
C3748 vdd.n2838 gnd 0.007322f
C3749 vdd.n2839 gnd 0.009097f
C3750 vdd.n2840 gnd 6.73985f
C3751 vdd.n2842 gnd 0.022678f
C3752 vdd.n2843 gnd 0.006077f
C3753 vdd.n2844 gnd 0.022678f
C3754 vdd.n2845 gnd 0.022169f
C3755 vdd.n2846 gnd 0.009097f
C3756 vdd.n2847 gnd 0.007322f
C3757 vdd.n2848 gnd 0.009097f
C3758 vdd.n2849 gnd 0.581022f
C3759 vdd.n2850 gnd 0.009097f
C3760 vdd.n2851 gnd 0.007322f
C3761 vdd.n2852 gnd 0.009097f
C3762 vdd.n2853 gnd 0.009097f
C3763 vdd.n2854 gnd 0.009097f
C3764 vdd.n2855 gnd 0.007322f
C3765 vdd.n2856 gnd 0.009097f
C3766 vdd.n2857 gnd 0.739059f
C3767 vdd.n2858 gnd 0.929634f
C3768 vdd.n2859 gnd 0.009097f
C3769 vdd.n2860 gnd 0.007322f
C3770 vdd.n2861 gnd 0.009097f
C3771 vdd.n2862 gnd 0.009097f
C3772 vdd.n2863 gnd 0.009097f
C3773 vdd.n2864 gnd 0.007322f
C3774 vdd.n2865 gnd 0.009097f
C3775 vdd.n2866 gnd 0.655392f
C3776 vdd.n2867 gnd 0.009097f
C3777 vdd.n2868 gnd 0.007322f
C3778 vdd.n2869 gnd 0.009097f
C3779 vdd.n2870 gnd 0.009097f
C3780 vdd.n2871 gnd 0.009097f
C3781 vdd.n2872 gnd 0.007322f
C3782 vdd.n2873 gnd 0.009097f
C3783 vdd.t145 gnd 0.464817f
C3784 vdd.n2874 gnd 0.771597f
C3785 vdd.n2875 gnd 0.009097f
C3786 vdd.n2876 gnd 0.007322f
C3787 vdd.n2877 gnd 0.009097f
C3788 vdd.n2878 gnd 0.009097f
C3789 vdd.n2879 gnd 0.009097f
C3790 vdd.n2880 gnd 0.007322f
C3791 vdd.n2881 gnd 0.009097f
C3792 vdd.n2882 gnd 0.729763f
C3793 vdd.n2883 gnd 0.009097f
C3794 vdd.n2884 gnd 0.007322f
C3795 vdd.n2885 gnd 0.009097f
C3796 vdd.n2886 gnd 0.009097f
C3797 vdd.n2887 gnd 0.009097f
C3798 vdd.n2888 gnd 0.007322f
C3799 vdd.n2889 gnd 0.007322f
C3800 vdd.n2890 gnd 0.007322f
C3801 vdd.n2891 gnd 0.009097f
C3802 vdd.n2892 gnd 0.009097f
C3803 vdd.n2893 gnd 0.009097f
C3804 vdd.n2894 gnd 0.007322f
C3805 vdd.n2895 gnd 0.007322f
C3806 vdd.n2896 gnd 0.007322f
C3807 vdd.n2897 gnd 0.009097f
C3808 vdd.n2898 gnd 0.009097f
C3809 vdd.n2899 gnd 0.009097f
C3810 vdd.n2900 gnd 0.007322f
C3811 vdd.n2901 gnd 0.007322f
C3812 vdd.n2902 gnd 0.006077f
C3813 vdd.n2903 gnd 0.022169f
C3814 vdd.n2904 gnd 0.022678f
C3815 vdd.n2906 gnd 0.022678f
C3816 vdd.n2907 gnd 0.003478f
C3817 vdd.t113 gnd 0.111913f
C3818 vdd.t112 gnd 0.119604f
C3819 vdd.t111 gnd 0.146157f
C3820 vdd.n2908 gnd 0.187352f
C3821 vdd.n2909 gnd 0.158142f
C3822 vdd.n2910 gnd 0.012008f
C3823 vdd.n2911 gnd 0.003844f
C3824 vdd.n2912 gnd 0.007322f
C3825 vdd.n2913 gnd 0.009097f
C3826 vdd.n2915 gnd 0.009097f
C3827 vdd.n2916 gnd 0.009097f
C3828 vdd.n2917 gnd 0.007322f
C3829 vdd.n2918 gnd 0.007322f
C3830 vdd.n2919 gnd 0.007322f
C3831 vdd.n2920 gnd 0.009097f
C3832 vdd.n2922 gnd 0.009097f
C3833 vdd.n2923 gnd 0.009097f
C3834 vdd.n2924 gnd 0.007322f
C3835 vdd.n2925 gnd 0.007322f
C3836 vdd.n2926 gnd 0.007322f
C3837 vdd.n2927 gnd 0.009097f
C3838 vdd.n2929 gnd 0.009097f
C3839 vdd.n2930 gnd 0.009097f
C3840 vdd.n2931 gnd 0.007322f
C3841 vdd.n2932 gnd 0.007322f
C3842 vdd.n2933 gnd 0.007322f
C3843 vdd.n2934 gnd 0.009097f
C3844 vdd.n2936 gnd 0.009097f
C3845 vdd.n2937 gnd 0.009097f
C3846 vdd.n2938 gnd 0.007322f
C3847 vdd.n2939 gnd 0.007322f
C3848 vdd.n2940 gnd 0.007322f
C3849 vdd.n2941 gnd 0.009097f
C3850 vdd.n2943 gnd 0.009097f
C3851 vdd.n2944 gnd 0.009097f
C3852 vdd.n2945 gnd 0.007322f
C3853 vdd.n2946 gnd 0.009097f
C3854 vdd.n2947 gnd 0.009097f
C3855 vdd.n2948 gnd 0.009097f
C3856 vdd.n2949 gnd 0.015668f
C3857 vdd.n2950 gnd 0.004979f
C3858 vdd.n2951 gnd 0.007322f
C3859 vdd.n2952 gnd 0.009097f
C3860 vdd.n2954 gnd 0.009097f
C3861 vdd.n2955 gnd 0.009097f
C3862 vdd.n2956 gnd 0.007322f
C3863 vdd.n2957 gnd 0.007322f
C3864 vdd.n2958 gnd 0.007322f
C3865 vdd.n2959 gnd 0.009097f
C3866 vdd.n2961 gnd 0.009097f
C3867 vdd.n2962 gnd 0.009097f
C3868 vdd.n2963 gnd 0.007322f
C3869 vdd.n2964 gnd 0.007322f
C3870 vdd.n2965 gnd 0.007322f
C3871 vdd.n2966 gnd 0.009097f
C3872 vdd.n2968 gnd 0.009097f
C3873 vdd.n2969 gnd 0.009097f
C3874 vdd.n2970 gnd 0.007322f
C3875 vdd.n2971 gnd 0.007322f
C3876 vdd.n2972 gnd 0.007322f
C3877 vdd.n2973 gnd 0.009097f
C3878 vdd.n2975 gnd 0.009097f
C3879 vdd.n2976 gnd 0.009097f
C3880 vdd.n2977 gnd 0.007322f
C3881 vdd.n2978 gnd 0.007322f
C3882 vdd.n2979 gnd 0.007322f
C3883 vdd.n2980 gnd 0.009097f
C3884 vdd.n2982 gnd 0.009097f
C3885 vdd.n2983 gnd 0.009097f
C3886 vdd.n2984 gnd 0.007322f
C3887 vdd.n2985 gnd 0.009097f
C3888 vdd.n2986 gnd 0.009097f
C3889 vdd.n2987 gnd 0.009097f
C3890 vdd.n2988 gnd 0.015668f
C3891 vdd.n2989 gnd 0.006114f
C3892 vdd.n2990 gnd 0.007322f
C3893 vdd.n2991 gnd 0.009097f
C3894 vdd.n2993 gnd 0.009097f
C3895 vdd.n2994 gnd 0.009097f
C3896 vdd.n2995 gnd 0.007322f
C3897 vdd.n2996 gnd 0.007322f
C3898 vdd.n2997 gnd 0.007322f
C3899 vdd.n2998 gnd 0.009097f
C3900 vdd.n3000 gnd 0.009097f
C3901 vdd.n3001 gnd 0.009097f
C3902 vdd.n3002 gnd 0.007322f
C3903 vdd.n3003 gnd 0.007322f
C3904 vdd.n3004 gnd 0.007322f
C3905 vdd.n3005 gnd 0.009097f
C3906 vdd.n3007 gnd 0.009097f
C3907 vdd.n3008 gnd 0.009097f
C3908 vdd.n3009 gnd 0.007322f
C3909 vdd.n3010 gnd 0.007322f
C3910 vdd.n3011 gnd 0.007322f
C3911 vdd.n3012 gnd 0.009097f
C3912 vdd.n3014 gnd 0.009097f
C3913 vdd.n3015 gnd 0.009097f
C3914 vdd.n3017 gnd 0.009097f
C3915 vdd.n3018 gnd 0.007322f
C3916 vdd.n3019 gnd 0.007322f
C3917 vdd.n3020 gnd 0.006077f
C3918 vdd.n3021 gnd 0.022678f
C3919 vdd.n3022 gnd 0.022169f
C3920 vdd.n3023 gnd 0.006077f
C3921 vdd.n3024 gnd 0.022169f
C3922 vdd.n3025 gnd 1.37121f
C3923 vdd.t64 gnd 0.464817f
C3924 vdd.n3026 gnd 0.488058f
C3925 vdd.n3027 gnd 0.929634f
C3926 vdd.n3028 gnd 0.009097f
C3927 vdd.n3029 gnd 0.007322f
C3928 vdd.n3030 gnd 0.007322f
C3929 vdd.n3031 gnd 0.007322f
C3930 vdd.n3032 gnd 0.009097f
C3931 vdd.n3033 gnd 0.832023f
C3932 vdd.t136 gnd 0.464817f
C3933 vdd.n3034 gnd 0.562429f
C3934 vdd.n3035 gnd 0.673985f
C3935 vdd.n3036 gnd 0.009097f
C3936 vdd.n3037 gnd 0.007322f
C3937 vdd.n3038 gnd 0.007322f
C3938 vdd.n3039 gnd 0.007322f
C3939 vdd.n3040 gnd 0.009097f
C3940 vdd.n3041 gnd 0.515947f
C3941 vdd.t158 gnd 0.464817f
C3942 vdd.n3042 gnd 0.771597f
C3943 vdd.t134 gnd 0.464817f
C3944 vdd.n3043 gnd 0.571725f
C3945 vdd.n3044 gnd 0.009097f
C3946 vdd.n3045 gnd 0.007322f
C3947 vdd.n3046 gnd 0.006991f
C3948 vdd.n3047 gnd 0.536555f
C3949 vdd.n3048 gnd 1.84238f
C3950 CSoutput.n0 gnd 0.037129f
C3951 CSoutput.t120 gnd 0.245601f
C3952 CSoutput.n1 gnd 0.110901f
C3953 CSoutput.n2 gnd 0.037129f
C3954 CSoutput.t125 gnd 0.245601f
C3955 CSoutput.n3 gnd 0.029428f
C3956 CSoutput.n4 gnd 0.037129f
C3957 CSoutput.t134 gnd 0.245601f
C3958 CSoutput.n5 gnd 0.025376f
C3959 CSoutput.n6 gnd 0.037129f
C3960 CSoutput.t123 gnd 0.245601f
C3961 CSoutput.t127 gnd 0.245601f
C3962 CSoutput.n7 gnd 0.109692f
C3963 CSoutput.n8 gnd 0.037129f
C3964 CSoutput.t133 gnd 0.245601f
C3965 CSoutput.n9 gnd 0.024194f
C3966 CSoutput.n10 gnd 0.037129f
C3967 CSoutput.t136 gnd 0.245601f
C3968 CSoutput.t124 gnd 0.245601f
C3969 CSoutput.n11 gnd 0.109692f
C3970 CSoutput.n12 gnd 0.037129f
C3971 CSoutput.t130 gnd 0.245601f
C3972 CSoutput.n13 gnd 0.025376f
C3973 CSoutput.n14 gnd 0.037129f
C3974 CSoutput.t129 gnd 0.245601f
C3975 CSoutput.t139 gnd 0.245601f
C3976 CSoutput.n15 gnd 0.109692f
C3977 CSoutput.n16 gnd 0.037129f
C3978 CSoutput.t128 gnd 0.245601f
C3979 CSoutput.n17 gnd 0.027103f
C3980 CSoutput.t137 gnd 0.293499f
C3981 CSoutput.t126 gnd 0.245601f
C3982 CSoutput.n18 gnd 0.140034f
C3983 CSoutput.n19 gnd 0.135882f
C3984 CSoutput.n20 gnd 0.157639f
C3985 CSoutput.n21 gnd 0.037129f
C3986 CSoutput.n22 gnd 0.030988f
C3987 CSoutput.n23 gnd 0.109692f
C3988 CSoutput.n24 gnd 0.029872f
C3989 CSoutput.n25 gnd 0.029428f
C3990 CSoutput.n26 gnd 0.037129f
C3991 CSoutput.n27 gnd 0.037129f
C3992 CSoutput.n28 gnd 0.03075f
C3993 CSoutput.n29 gnd 0.026108f
C3994 CSoutput.n30 gnd 0.112134f
C3995 CSoutput.n31 gnd 0.026467f
C3996 CSoutput.n32 gnd 0.037129f
C3997 CSoutput.n33 gnd 0.037129f
C3998 CSoutput.n34 gnd 0.037129f
C3999 CSoutput.n35 gnd 0.030423f
C4000 CSoutput.n36 gnd 0.109692f
C4001 CSoutput.n37 gnd 0.029095f
C4002 CSoutput.n38 gnd 0.030205f
C4003 CSoutput.n39 gnd 0.037129f
C4004 CSoutput.n40 gnd 0.037129f
C4005 CSoutput.n41 gnd 0.030982f
C4006 CSoutput.n42 gnd 0.028318f
C4007 CSoutput.n43 gnd 0.109692f
C4008 CSoutput.n44 gnd 0.029035f
C4009 CSoutput.n45 gnd 0.037129f
C4010 CSoutput.n46 gnd 0.037129f
C4011 CSoutput.n47 gnd 0.037129f
C4012 CSoutput.n48 gnd 0.029035f
C4013 CSoutput.n49 gnd 0.109692f
C4014 CSoutput.n50 gnd 0.028318f
C4015 CSoutput.n51 gnd 0.030982f
C4016 CSoutput.n52 gnd 0.037129f
C4017 CSoutput.n53 gnd 0.037129f
C4018 CSoutput.n54 gnd 0.030205f
C4019 CSoutput.n55 gnd 0.029095f
C4020 CSoutput.n56 gnd 0.109692f
C4021 CSoutput.n57 gnd 0.030423f
C4022 CSoutput.n58 gnd 0.037129f
C4023 CSoutput.n59 gnd 0.037129f
C4024 CSoutput.n60 gnd 0.037129f
C4025 CSoutput.n61 gnd 0.026467f
C4026 CSoutput.n62 gnd 0.112134f
C4027 CSoutput.n63 gnd 0.026108f
C4028 CSoutput.t135 gnd 0.245601f
C4029 CSoutput.n64 gnd 0.109692f
C4030 CSoutput.n65 gnd 0.03075f
C4031 CSoutput.n66 gnd 0.037129f
C4032 CSoutput.n67 gnd 0.037129f
C4033 CSoutput.n68 gnd 0.037129f
C4034 CSoutput.n69 gnd 0.029872f
C4035 CSoutput.n70 gnd 0.109692f
C4036 CSoutput.n71 gnd 0.030988f
C4037 CSoutput.n72 gnd 0.027103f
C4038 CSoutput.n73 gnd 0.037129f
C4039 CSoutput.n74 gnd 0.037129f
C4040 CSoutput.n75 gnd 0.028107f
C4041 CSoutput.n76 gnd 0.016693f
C4042 CSoutput.t138 gnd 0.27595f
C4043 CSoutput.n77 gnd 0.137081f
C4044 CSoutput.n78 gnd 0.560791f
C4045 CSoutput.t85 gnd 0.046313f
C4046 CSoutput.t96 gnd 0.046313f
C4047 CSoutput.n79 gnd 0.358573f
C4048 CSoutput.t80 gnd 0.046313f
C4049 CSoutput.t95 gnd 0.046313f
C4050 CSoutput.n80 gnd 0.357933f
C4051 CSoutput.n81 gnd 0.363302f
C4052 CSoutput.t113 gnd 0.046313f
C4053 CSoutput.t90 gnd 0.046313f
C4054 CSoutput.n82 gnd 0.357933f
C4055 CSoutput.n83 gnd 0.17902f
C4056 CSoutput.t106 gnd 0.046313f
C4057 CSoutput.t105 gnd 0.046313f
C4058 CSoutput.n84 gnd 0.357933f
C4059 CSoutput.n85 gnd 0.328281f
C4060 CSoutput.t83 gnd 0.046313f
C4061 CSoutput.t92 gnd 0.046313f
C4062 CSoutput.n86 gnd 0.358573f
C4063 CSoutput.t87 gnd 0.046313f
C4064 CSoutput.t82 gnd 0.046313f
C4065 CSoutput.n87 gnd 0.357933f
C4066 CSoutput.n88 gnd 0.363302f
C4067 CSoutput.t89 gnd 0.046313f
C4068 CSoutput.t112 gnd 0.046313f
C4069 CSoutput.n89 gnd 0.357933f
C4070 CSoutput.n90 gnd 0.17902f
C4071 CSoutput.t86 gnd 0.046313f
C4072 CSoutput.t119 gnd 0.046313f
C4073 CSoutput.n91 gnd 0.357933f
C4074 CSoutput.n92 gnd 0.266964f
C4075 CSoutput.n93 gnd 0.336639f
C4076 CSoutput.t76 gnd 0.046313f
C4077 CSoutput.t77 gnd 0.046313f
C4078 CSoutput.n94 gnd 0.358573f
C4079 CSoutput.t115 gnd 0.046313f
C4080 CSoutput.t74 gnd 0.046313f
C4081 CSoutput.n95 gnd 0.357933f
C4082 CSoutput.n96 gnd 0.363302f
C4083 CSoutput.t110 gnd 0.046313f
C4084 CSoutput.t75 gnd 0.046313f
C4085 CSoutput.n97 gnd 0.357933f
C4086 CSoutput.n98 gnd 0.17902f
C4087 CSoutput.t114 gnd 0.046313f
C4088 CSoutput.t100 gnd 0.046313f
C4089 CSoutput.n99 gnd 0.357933f
C4090 CSoutput.n100 gnd 0.266964f
C4091 CSoutput.n101 gnd 0.376277f
C4092 CSoutput.n102 gnd 6.73022f
C4093 CSoutput.n104 gnd 0.656807f
C4094 CSoutput.n105 gnd 0.492605f
C4095 CSoutput.n106 gnd 0.656807f
C4096 CSoutput.n107 gnd 0.656807f
C4097 CSoutput.n108 gnd 1.76833f
C4098 CSoutput.n109 gnd 0.656807f
C4099 CSoutput.n110 gnd 0.656807f
C4100 CSoutput.t131 gnd 0.821008f
C4101 CSoutput.n111 gnd 0.656807f
C4102 CSoutput.n112 gnd 0.656807f
C4103 CSoutput.n116 gnd 0.656807f
C4104 CSoutput.n120 gnd 0.656807f
C4105 CSoutput.n121 gnd 0.656807f
C4106 CSoutput.n123 gnd 0.656807f
C4107 CSoutput.n128 gnd 0.656807f
C4108 CSoutput.n130 gnd 0.656807f
C4109 CSoutput.n131 gnd 0.656807f
C4110 CSoutput.n133 gnd 0.656807f
C4111 CSoutput.n134 gnd 0.656807f
C4112 CSoutput.n136 gnd 0.656807f
C4113 CSoutput.t121 gnd 10.9752f
C4114 CSoutput.n138 gnd 0.656807f
C4115 CSoutput.n139 gnd 0.492605f
C4116 CSoutput.n140 gnd 0.656807f
C4117 CSoutput.n141 gnd 0.656807f
C4118 CSoutput.n142 gnd 1.76833f
C4119 CSoutput.n143 gnd 0.656807f
C4120 CSoutput.n144 gnd 0.656807f
C4121 CSoutput.t140 gnd 0.821008f
C4122 CSoutput.n145 gnd 0.656807f
C4123 CSoutput.n146 gnd 0.656807f
C4124 CSoutput.n150 gnd 0.656807f
C4125 CSoutput.n154 gnd 0.656807f
C4126 CSoutput.n155 gnd 0.656807f
C4127 CSoutput.n157 gnd 0.656807f
C4128 CSoutput.n162 gnd 0.656807f
C4129 CSoutput.n164 gnd 0.656807f
C4130 CSoutput.n165 gnd 0.656807f
C4131 CSoutput.n167 gnd 0.656807f
C4132 CSoutput.n168 gnd 0.656807f
C4133 CSoutput.n170 gnd 0.656807f
C4134 CSoutput.n171 gnd 0.492605f
C4135 CSoutput.n173 gnd 0.656807f
C4136 CSoutput.n174 gnd 0.492605f
C4137 CSoutput.n175 gnd 0.656807f
C4138 CSoutput.n176 gnd 0.656807f
C4139 CSoutput.n177 gnd 1.76833f
C4140 CSoutput.n178 gnd 0.656807f
C4141 CSoutput.n179 gnd 0.656807f
C4142 CSoutput.t132 gnd 0.821008f
C4143 CSoutput.n180 gnd 0.656807f
C4144 CSoutput.n181 gnd 1.76833f
C4145 CSoutput.n183 gnd 0.656807f
C4146 CSoutput.n184 gnd 0.656807f
C4147 CSoutput.n186 gnd 0.656807f
C4148 CSoutput.n187 gnd 0.656807f
C4149 CSoutput.t141 gnd 10.7963f
C4150 CSoutput.t122 gnd 10.9752f
C4151 CSoutput.n193 gnd 2.0605f
C4152 CSoutput.n194 gnd 8.39372f
C4153 CSoutput.n195 gnd 8.74495f
C4154 CSoutput.n200 gnd 2.23207f
C4155 CSoutput.n206 gnd 0.656807f
C4156 CSoutput.n208 gnd 0.656807f
C4157 CSoutput.n210 gnd 0.656807f
C4158 CSoutput.n212 gnd 0.656807f
C4159 CSoutput.n214 gnd 0.656807f
C4160 CSoutput.n220 gnd 0.656807f
C4161 CSoutput.n227 gnd 1.20499f
C4162 CSoutput.n228 gnd 1.20499f
C4163 CSoutput.n229 gnd 0.656807f
C4164 CSoutput.n230 gnd 0.656807f
C4165 CSoutput.n232 gnd 0.492605f
C4166 CSoutput.n233 gnd 0.421872f
C4167 CSoutput.n235 gnd 0.492605f
C4168 CSoutput.n236 gnd 0.421872f
C4169 CSoutput.n237 gnd 0.492605f
C4170 CSoutput.n239 gnd 0.656807f
C4171 CSoutput.n241 gnd 1.76833f
C4172 CSoutput.n242 gnd 2.0605f
C4173 CSoutput.n243 gnd 7.72006f
C4174 CSoutput.n245 gnd 0.492605f
C4175 CSoutput.n246 gnd 1.2675f
C4176 CSoutput.n247 gnd 0.492605f
C4177 CSoutput.n249 gnd 0.656807f
C4178 CSoutput.n251 gnd 1.76833f
C4179 CSoutput.n252 gnd 3.8517f
C4180 CSoutput.t88 gnd 0.046313f
C4181 CSoutput.t84 gnd 0.046313f
C4182 CSoutput.n253 gnd 0.358573f
C4183 CSoutput.t97 gnd 0.046313f
C4184 CSoutput.t108 gnd 0.046313f
C4185 CSoutput.n254 gnd 0.357933f
C4186 CSoutput.n255 gnd 0.363302f
C4187 CSoutput.t91 gnd 0.046313f
C4188 CSoutput.t111 gnd 0.046313f
C4189 CSoutput.n256 gnd 0.357933f
C4190 CSoutput.n257 gnd 0.17902f
C4191 CSoutput.t117 gnd 0.046313f
C4192 CSoutput.t107 gnd 0.046313f
C4193 CSoutput.n258 gnd 0.357933f
C4194 CSoutput.n259 gnd 0.328281f
C4195 CSoutput.t98 gnd 0.046313f
C4196 CSoutput.t99 gnd 0.046313f
C4197 CSoutput.n260 gnd 0.358573f
C4198 CSoutput.t79 gnd 0.046313f
C4199 CSoutput.t81 gnd 0.046313f
C4200 CSoutput.n261 gnd 0.357933f
C4201 CSoutput.n262 gnd 0.363302f
C4202 CSoutput.t94 gnd 0.046313f
C4203 CSoutput.t78 gnd 0.046313f
C4204 CSoutput.n263 gnd 0.357933f
C4205 CSoutput.n264 gnd 0.17902f
C4206 CSoutput.t72 gnd 0.046313f
C4207 CSoutput.t104 gnd 0.046313f
C4208 CSoutput.n265 gnd 0.357933f
C4209 CSoutput.n266 gnd 0.266964f
C4210 CSoutput.n267 gnd 0.336639f
C4211 CSoutput.t102 gnd 0.046313f
C4212 CSoutput.t103 gnd 0.046313f
C4213 CSoutput.n268 gnd 0.358573f
C4214 CSoutput.t93 gnd 0.046313f
C4215 CSoutput.t73 gnd 0.046313f
C4216 CSoutput.n269 gnd 0.357933f
C4217 CSoutput.n270 gnd 0.363302f
C4218 CSoutput.t101 gnd 0.046313f
C4219 CSoutput.t116 gnd 0.046313f
C4220 CSoutput.n271 gnd 0.357933f
C4221 CSoutput.n272 gnd 0.17902f
C4222 CSoutput.t109 gnd 0.046313f
C4223 CSoutput.t118 gnd 0.046313f
C4224 CSoutput.n273 gnd 0.357932f
C4225 CSoutput.n274 gnd 0.266965f
C4226 CSoutput.n275 gnd 0.376277f
C4227 CSoutput.n276 gnd 9.68117f
C4228 CSoutput.t63 gnd 0.040524f
C4229 CSoutput.t10 gnd 0.040524f
C4230 CSoutput.n277 gnd 0.359284f
C4231 CSoutput.t50 gnd 0.040524f
C4232 CSoutput.t0 gnd 0.040524f
C4233 CSoutput.n278 gnd 0.358085f
C4234 CSoutput.n279 gnd 0.333669f
C4235 CSoutput.t34 gnd 0.040524f
C4236 CSoutput.t65 gnd 0.040524f
C4237 CSoutput.n280 gnd 0.358085f
C4238 CSoutput.n281 gnd 0.164483f
C4239 CSoutput.t19 gnd 0.040524f
C4240 CSoutput.t32 gnd 0.040524f
C4241 CSoutput.n282 gnd 0.358085f
C4242 CSoutput.n283 gnd 0.164483f
C4243 CSoutput.t4 gnd 0.040524f
C4244 CSoutput.t40 gnd 0.040524f
C4245 CSoutput.n284 gnd 0.358085f
C4246 CSoutput.n285 gnd 0.164483f
C4247 CSoutput.t53 gnd 0.040524f
C4248 CSoutput.t24 gnd 0.040524f
C4249 CSoutput.n286 gnd 0.358085f
C4250 CSoutput.n287 gnd 0.30338f
C4251 CSoutput.t30 gnd 0.040524f
C4252 CSoutput.t13 gnd 0.040524f
C4253 CSoutput.n288 gnd 0.359284f
C4254 CSoutput.t18 gnd 0.040524f
C4255 CSoutput.t31 gnd 0.040524f
C4256 CSoutput.n289 gnd 0.358085f
C4257 CSoutput.n290 gnd 0.333669f
C4258 CSoutput.t14 gnd 0.040524f
C4259 CSoutput.t20 gnd 0.040524f
C4260 CSoutput.n291 gnd 0.358085f
C4261 CSoutput.n292 gnd 0.164483f
C4262 CSoutput.t33 gnd 0.040524f
C4263 CSoutput.t11 gnd 0.040524f
C4264 CSoutput.n293 gnd 0.358085f
C4265 CSoutput.n294 gnd 0.164483f
C4266 CSoutput.t21 gnd 0.040524f
C4267 CSoutput.t7 gnd 0.040524f
C4268 CSoutput.n295 gnd 0.358085f
C4269 CSoutput.n296 gnd 0.164483f
C4270 CSoutput.t12 gnd 0.040524f
C4271 CSoutput.t22 gnd 0.040524f
C4272 CSoutput.n297 gnd 0.358085f
C4273 CSoutput.n298 gnd 0.24972f
C4274 CSoutput.n299 gnd 0.314975f
C4275 CSoutput.t8 gnd 0.040524f
C4276 CSoutput.t69 gnd 0.040524f
C4277 CSoutput.n300 gnd 0.359284f
C4278 CSoutput.t59 gnd 0.040524f
C4279 CSoutput.t15 gnd 0.040524f
C4280 CSoutput.n301 gnd 0.358085f
C4281 CSoutput.n302 gnd 0.333669f
C4282 CSoutput.t1 gnd 0.040524f
C4283 CSoutput.t67 gnd 0.040524f
C4284 CSoutput.n303 gnd 0.358085f
C4285 CSoutput.n304 gnd 0.164483f
C4286 CSoutput.t26 gnd 0.040524f
C4287 CSoutput.t35 gnd 0.040524f
C4288 CSoutput.n305 gnd 0.358085f
C4289 CSoutput.n306 gnd 0.164483f
C4290 CSoutput.t70 gnd 0.040524f
C4291 CSoutput.t60 gnd 0.040524f
C4292 CSoutput.n307 gnd 0.358085f
C4293 CSoutput.n308 gnd 0.164483f
C4294 CSoutput.t44 gnd 0.040524f
C4295 CSoutput.t2 gnd 0.040524f
C4296 CSoutput.n309 gnd 0.358085f
C4297 CSoutput.n310 gnd 0.24972f
C4298 CSoutput.n311 gnd 0.338234f
C4299 CSoutput.n312 gnd 10.3298f
C4300 CSoutput.t41 gnd 0.040524f
C4301 CSoutput.t5 gnd 0.040524f
C4302 CSoutput.n313 gnd 0.359284f
C4303 CSoutput.t25 gnd 0.040524f
C4304 CSoutput.t66 gnd 0.040524f
C4305 CSoutput.n314 gnd 0.358085f
C4306 CSoutput.n315 gnd 0.333669f
C4307 CSoutput.t6 gnd 0.040524f
C4308 CSoutput.t55 gnd 0.040524f
C4309 CSoutput.n316 gnd 0.358085f
C4310 CSoutput.n317 gnd 0.164483f
C4311 CSoutput.t54 gnd 0.040524f
C4312 CSoutput.t43 gnd 0.040524f
C4313 CSoutput.n318 gnd 0.358085f
C4314 CSoutput.n319 gnd 0.164483f
C4315 CSoutput.t56 gnd 0.040524f
C4316 CSoutput.t27 gnd 0.040524f
C4317 CSoutput.n320 gnd 0.358085f
C4318 CSoutput.n321 gnd 0.164483f
C4319 CSoutput.t49 gnd 0.040524f
C4320 CSoutput.t61 gnd 0.040524f
C4321 CSoutput.n322 gnd 0.358085f
C4322 CSoutput.n323 gnd 0.30338f
C4323 CSoutput.t28 gnd 0.040524f
C4324 CSoutput.t45 gnd 0.040524f
C4325 CSoutput.n324 gnd 0.359284f
C4326 CSoutput.t46 gnd 0.040524f
C4327 CSoutput.t36 gnd 0.040524f
C4328 CSoutput.n325 gnd 0.358085f
C4329 CSoutput.n326 gnd 0.333669f
C4330 CSoutput.t37 gnd 0.040524f
C4331 CSoutput.t29 gnd 0.040524f
C4332 CSoutput.n327 gnd 0.358085f
C4333 CSoutput.n328 gnd 0.164483f
C4334 CSoutput.t23 gnd 0.040524f
C4335 CSoutput.t16 gnd 0.040524f
C4336 CSoutput.n329 gnd 0.358085f
C4337 CSoutput.n330 gnd 0.164483f
C4338 CSoutput.t17 gnd 0.040524f
C4339 CSoutput.t38 gnd 0.040524f
C4340 CSoutput.n331 gnd 0.358085f
C4341 CSoutput.n332 gnd 0.164483f
C4342 CSoutput.t39 gnd 0.040524f
C4343 CSoutput.t3 gnd 0.040524f
C4344 CSoutput.n333 gnd 0.358085f
C4345 CSoutput.n334 gnd 0.24972f
C4346 CSoutput.n335 gnd 0.314975f
C4347 CSoutput.t57 gnd 0.040524f
C4348 CSoutput.t68 gnd 0.040524f
C4349 CSoutput.n336 gnd 0.359284f
C4350 CSoutput.t71 gnd 0.040524f
C4351 CSoutput.t48 gnd 0.040524f
C4352 CSoutput.n337 gnd 0.358085f
C4353 CSoutput.n338 gnd 0.333669f
C4354 CSoutput.t52 gnd 0.040524f
C4355 CSoutput.t62 gnd 0.040524f
C4356 CSoutput.n339 gnd 0.358085f
C4357 CSoutput.n340 gnd 0.164483f
C4358 CSoutput.t9 gnd 0.040524f
C4359 CSoutput.t42 gnd 0.040524f
C4360 CSoutput.n341 gnd 0.358085f
C4361 CSoutput.n342 gnd 0.164483f
C4362 CSoutput.t47 gnd 0.040524f
C4363 CSoutput.t58 gnd 0.040524f
C4364 CSoutput.n343 gnd 0.358085f
C4365 CSoutput.n344 gnd 0.164483f
C4366 CSoutput.t64 gnd 0.040524f
C4367 CSoutput.t51 gnd 0.040524f
C4368 CSoutput.n345 gnd 0.358085f
C4369 CSoutput.n346 gnd 0.24972f
C4370 CSoutput.n347 gnd 0.338234f
C4371 CSoutput.n348 gnd 5.8275f
C4372 CSoutput.n349 gnd 11.424901f
C4373 a_n5644_8799.n0 gnd 0.213234f
C4374 a_n5644_8799.n1 gnd 0.293964f
C4375 a_n5644_8799.n2 gnd 0.223034f
C4376 a_n5644_8799.n3 gnd 0.213234f
C4377 a_n5644_8799.n4 gnd 0.293964f
C4378 a_n5644_8799.n5 gnd 0.223034f
C4379 a_n5644_8799.n6 gnd 0.213234f
C4380 a_n5644_8799.n7 gnd 0.463262f
C4381 a_n5644_8799.n8 gnd 0.223034f
C4382 a_n5644_8799.n9 gnd 0.213234f
C4383 a_n5644_8799.n10 gnd 0.329651f
C4384 a_n5644_8799.n11 gnd 0.187347f
C4385 a_n5644_8799.n12 gnd 0.213234f
C4386 a_n5644_8799.n13 gnd 0.329651f
C4387 a_n5644_8799.n14 gnd 0.187347f
C4388 a_n5644_8799.n15 gnd 0.213234f
C4389 a_n5644_8799.n16 gnd 0.329651f
C4390 a_n5644_8799.n17 gnd 0.356645f
C4391 a_n5644_8799.n18 gnd 3.49946f
C4392 a_n5644_8799.n19 gnd 1.78434f
C4393 a_n5644_8799.n20 gnd 3.03595f
C4394 a_n5644_8799.n21 gnd 2.90994f
C4395 a_n5644_8799.n22 gnd 4.07258f
C4396 a_n5644_8799.n23 gnd 0.717892f
C4397 a_n5644_8799.n24 gnd 0.256713f
C4398 a_n5644_8799.n25 gnd 0.004793f
C4399 a_n5644_8799.n26 gnd 0.010365f
C4400 a_n5644_8799.n27 gnd 0.010365f
C4401 a_n5644_8799.n28 gnd 0.004793f
C4402 a_n5644_8799.n29 gnd 0.256713f
C4403 a_n5644_8799.n30 gnd 0.004793f
C4404 a_n5644_8799.n31 gnd 0.010365f
C4405 a_n5644_8799.n32 gnd 0.010365f
C4406 a_n5644_8799.n33 gnd 0.004793f
C4407 a_n5644_8799.n34 gnd 0.256713f
C4408 a_n5644_8799.n35 gnd 0.004793f
C4409 a_n5644_8799.n36 gnd 0.010365f
C4410 a_n5644_8799.n37 gnd 0.010365f
C4411 a_n5644_8799.n38 gnd 0.004793f
C4412 a_n5644_8799.n39 gnd 0.004793f
C4413 a_n5644_8799.n40 gnd 0.010365f
C4414 a_n5644_8799.n41 gnd 0.010365f
C4415 a_n5644_8799.n42 gnd 0.004793f
C4416 a_n5644_8799.n43 gnd 0.256713f
C4417 a_n5644_8799.n44 gnd 0.004793f
C4418 a_n5644_8799.n45 gnd 0.010365f
C4419 a_n5644_8799.n46 gnd 0.010365f
C4420 a_n5644_8799.n47 gnd 0.004793f
C4421 a_n5644_8799.n48 gnd 0.256713f
C4422 a_n5644_8799.n49 gnd 0.004793f
C4423 a_n5644_8799.n50 gnd 0.010365f
C4424 a_n5644_8799.n51 gnd 0.010365f
C4425 a_n5644_8799.n52 gnd 0.004793f
C4426 a_n5644_8799.n53 gnd 0.256713f
C4427 a_n5644_8799.t11 gnd 0.147901f
C4428 a_n5644_8799.t13 gnd 0.147901f
C4429 a_n5644_8799.t32 gnd 0.147901f
C4430 a_n5644_8799.n54 gnd 1.16652f
C4431 a_n5644_8799.t15 gnd 0.147901f
C4432 a_n5644_8799.t20 gnd 0.147901f
C4433 a_n5644_8799.n55 gnd 1.1646f
C4434 a_n5644_8799.t19 gnd 0.147901f
C4435 a_n5644_8799.t18 gnd 0.147901f
C4436 a_n5644_8799.n56 gnd 1.1646f
C4437 a_n5644_8799.t27 gnd 0.115034f
C4438 a_n5644_8799.t26 gnd 0.115034f
C4439 a_n5644_8799.n57 gnd 1.0181f
C4440 a_n5644_8799.t6 gnd 0.115034f
C4441 a_n5644_8799.t16 gnd 0.115034f
C4442 a_n5644_8799.n58 gnd 1.01648f
C4443 a_n5644_8799.t25 gnd 0.115034f
C4444 a_n5644_8799.t24 gnd 0.115034f
C4445 a_n5644_8799.n59 gnd 1.01648f
C4446 a_n5644_8799.t33 gnd 0.115034f
C4447 a_n5644_8799.t22 gnd 0.115034f
C4448 a_n5644_8799.n60 gnd 1.0181f
C4449 a_n5644_8799.t2 gnd 0.115034f
C4450 a_n5644_8799.t17 gnd 0.115034f
C4451 a_n5644_8799.n61 gnd 1.01648f
C4452 a_n5644_8799.t3 gnd 0.115034f
C4453 a_n5644_8799.t1 gnd 0.115034f
C4454 a_n5644_8799.n62 gnd 1.01648f
C4455 a_n5644_8799.t14 gnd 0.115034f
C4456 a_n5644_8799.t23 gnd 0.115034f
C4457 a_n5644_8799.n63 gnd 1.0181f
C4458 a_n5644_8799.t34 gnd 0.115034f
C4459 a_n5644_8799.t29 gnd 0.115034f
C4460 a_n5644_8799.n64 gnd 1.01648f
C4461 a_n5644_8799.t4 gnd 0.115034f
C4462 a_n5644_8799.t8 gnd 0.115034f
C4463 a_n5644_8799.n65 gnd 1.01648f
C4464 a_n5644_8799.t28 gnd 0.115034f
C4465 a_n5644_8799.t5 gnd 0.115034f
C4466 a_n5644_8799.n66 gnd 1.01648f
C4467 a_n5644_8799.t0 gnd 0.115034f
C4468 a_n5644_8799.t35 gnd 0.115034f
C4469 a_n5644_8799.n67 gnd 1.01648f
C4470 a_n5644_8799.t21 gnd 0.115034f
C4471 a_n5644_8799.t31 gnd 0.115034f
C4472 a_n5644_8799.n68 gnd 1.01648f
C4473 a_n5644_8799.t75 gnd 0.613267f
C4474 a_n5644_8799.n69 gnd 0.275628f
C4475 a_n5644_8799.t42 gnd 0.613267f
C4476 a_n5644_8799.t62 gnd 0.613267f
C4477 a_n5644_8799.t53 gnd 0.624874f
C4478 a_n5644_8799.n70 gnd 0.257091f
C4479 a_n5644_8799.n71 gnd 0.278079f
C4480 a_n5644_8799.t77 gnd 0.613267f
C4481 a_n5644_8799.n72 gnd 0.275628f
C4482 a_n5644_8799.n73 gnd 0.271103f
C4483 a_n5644_8799.t52 gnd 0.613267f
C4484 a_n5644_8799.n74 gnd 0.271103f
C4485 a_n5644_8799.t41 gnd 0.613267f
C4486 a_n5644_8799.n75 gnd 0.278079f
C4487 a_n5644_8799.t40 gnd 0.624864f
C4488 a_n5644_8799.t79 gnd 0.613267f
C4489 a_n5644_8799.n76 gnd 0.275628f
C4490 a_n5644_8799.t49 gnd 0.613267f
C4491 a_n5644_8799.t68 gnd 0.613267f
C4492 a_n5644_8799.t58 gnd 0.624874f
C4493 a_n5644_8799.n77 gnd 0.257091f
C4494 a_n5644_8799.n78 gnd 0.278079f
C4495 a_n5644_8799.t81 gnd 0.613267f
C4496 a_n5644_8799.n79 gnd 0.275628f
C4497 a_n5644_8799.n80 gnd 0.271103f
C4498 a_n5644_8799.t57 gnd 0.613267f
C4499 a_n5644_8799.n81 gnd 0.271103f
C4500 a_n5644_8799.t45 gnd 0.613267f
C4501 a_n5644_8799.n82 gnd 0.278079f
C4502 a_n5644_8799.t47 gnd 0.624864f
C4503 a_n5644_8799.n83 gnd 0.922333f
C4504 a_n5644_8799.t66 gnd 0.613267f
C4505 a_n5644_8799.n84 gnd 0.275628f
C4506 a_n5644_8799.t74 gnd 0.613267f
C4507 a_n5644_8799.t71 gnd 0.613267f
C4508 a_n5644_8799.t39 gnd 0.624874f
C4509 a_n5644_8799.n85 gnd 0.257091f
C4510 a_n5644_8799.n86 gnd 0.278079f
C4511 a_n5644_8799.t48 gnd 0.613267f
C4512 a_n5644_8799.n87 gnd 0.275628f
C4513 a_n5644_8799.n88 gnd 0.271103f
C4514 a_n5644_8799.t54 gnd 0.613267f
C4515 a_n5644_8799.n89 gnd 0.271103f
C4516 a_n5644_8799.t43 gnd 0.613267f
C4517 a_n5644_8799.n90 gnd 0.278079f
C4518 a_n5644_8799.t83 gnd 0.624864f
C4519 a_n5644_8799.n91 gnd 1.49112f
C4520 a_n5644_8799.t60 gnd 0.624864f
C4521 a_n5644_8799.t59 gnd 0.613267f
C4522 a_n5644_8799.t46 gnd 0.613267f
C4523 a_n5644_8799.n92 gnd 0.275628f
C4524 a_n5644_8799.t76 gnd 0.613267f
C4525 a_n5644_8799.t61 gnd 0.613267f
C4526 a_n5644_8799.t51 gnd 0.613267f
C4527 a_n5644_8799.n93 gnd 0.275628f
C4528 a_n5644_8799.t69 gnd 0.624874f
C4529 a_n5644_8799.n94 gnd 0.257091f
C4530 a_n5644_8799.t78 gnd 0.613267f
C4531 a_n5644_8799.n95 gnd 0.278079f
C4532 a_n5644_8799.n96 gnd 0.271103f
C4533 a_n5644_8799.n97 gnd 0.271103f
C4534 a_n5644_8799.n98 gnd 0.278079f
C4535 a_n5644_8799.t64 gnd 0.624864f
C4536 a_n5644_8799.t63 gnd 0.613267f
C4537 a_n5644_8799.t55 gnd 0.613267f
C4538 a_n5644_8799.n99 gnd 0.275628f
C4539 a_n5644_8799.t80 gnd 0.613267f
C4540 a_n5644_8799.t67 gnd 0.613267f
C4541 a_n5644_8799.t56 gnd 0.613267f
C4542 a_n5644_8799.n100 gnd 0.275628f
C4543 a_n5644_8799.t72 gnd 0.624874f
C4544 a_n5644_8799.n101 gnd 0.257091f
C4545 a_n5644_8799.t36 gnd 0.613267f
C4546 a_n5644_8799.n102 gnd 0.278079f
C4547 a_n5644_8799.n103 gnd 0.271103f
C4548 a_n5644_8799.n104 gnd 0.271103f
C4549 a_n5644_8799.n105 gnd 0.278079f
C4550 a_n5644_8799.n106 gnd 0.922333f
C4551 a_n5644_8799.t82 gnd 0.624864f
C4552 a_n5644_8799.t44 gnd 0.613267f
C4553 a_n5644_8799.t65 gnd 0.613267f
C4554 a_n5644_8799.n107 gnd 0.275628f
C4555 a_n5644_8799.t37 gnd 0.613267f
C4556 a_n5644_8799.t73 gnd 0.613267f
C4557 a_n5644_8799.t50 gnd 0.613267f
C4558 a_n5644_8799.n108 gnd 0.275628f
C4559 a_n5644_8799.t38 gnd 0.624874f
C4560 a_n5644_8799.n109 gnd 0.257091f
C4561 a_n5644_8799.t70 gnd 0.613267f
C4562 a_n5644_8799.n110 gnd 0.278079f
C4563 a_n5644_8799.n111 gnd 0.271103f
C4564 a_n5644_8799.n112 gnd 0.271103f
C4565 a_n5644_8799.n113 gnd 0.278079f
C4566 a_n5644_8799.n114 gnd 1.1661f
C4567 a_n5644_8799.n115 gnd 12.562f
C4568 a_n5644_8799.n116 gnd 4.48823f
C4569 a_n5644_8799.n117 gnd 5.8395f
C4570 a_n5644_8799.t9 gnd 0.147901f
C4571 a_n5644_8799.t10 gnd 0.147901f
C4572 a_n5644_8799.n118 gnd 1.1646f
C4573 a_n5644_8799.t30 gnd 0.147901f
C4574 a_n5644_8799.t12 gnd 0.147901f
C4575 a_n5644_8799.n119 gnd 1.16652f
C4576 a_n5644_8799.n120 gnd 1.1646f
C4577 a_n5644_8799.t7 gnd 0.147901f
C4578 commonsourceibias.n0 gnd 0.012299f
C4579 commonsourceibias.t56 gnd 0.18623f
C4580 commonsourceibias.t109 gnd 0.172196f
C4581 commonsourceibias.n1 gnd 0.068706f
C4582 commonsourceibias.n2 gnd 0.009217f
C4583 commonsourceibias.t69 gnd 0.172196f
C4584 commonsourceibias.n3 gnd 0.007456f
C4585 commonsourceibias.n4 gnd 0.009217f
C4586 commonsourceibias.t119 gnd 0.172196f
C4587 commonsourceibias.n5 gnd 0.008898f
C4588 commonsourceibias.n6 gnd 0.009217f
C4589 commonsourceibias.t85 gnd 0.172196f
C4590 commonsourceibias.n7 gnd 0.068706f
C4591 commonsourceibias.t54 gnd 0.172196f
C4592 commonsourceibias.n8 gnd 0.007444f
C4593 commonsourceibias.n9 gnd 0.012299f
C4594 commonsourceibias.t16 gnd 0.18623f
C4595 commonsourceibias.t30 gnd 0.172196f
C4596 commonsourceibias.n10 gnd 0.068706f
C4597 commonsourceibias.n11 gnd 0.009217f
C4598 commonsourceibias.t2 gnd 0.172196f
C4599 commonsourceibias.n12 gnd 0.007456f
C4600 commonsourceibias.n13 gnd 0.009217f
C4601 commonsourceibias.t22 gnd 0.172196f
C4602 commonsourceibias.n14 gnd 0.008898f
C4603 commonsourceibias.n15 gnd 0.009217f
C4604 commonsourceibias.t42 gnd 0.172196f
C4605 commonsourceibias.n16 gnd 0.068706f
C4606 commonsourceibias.t18 gnd 0.172196f
C4607 commonsourceibias.n17 gnd 0.007444f
C4608 commonsourceibias.n18 gnd 0.009217f
C4609 commonsourceibias.t32 gnd 0.172196f
C4610 commonsourceibias.t40 gnd 0.172196f
C4611 commonsourceibias.n19 gnd 0.068706f
C4612 commonsourceibias.n20 gnd 0.009217f
C4613 commonsourceibias.t24 gnd 0.172196f
C4614 commonsourceibias.n21 gnd 0.068706f
C4615 commonsourceibias.n22 gnd 0.009217f
C4616 commonsourceibias.t44 gnd 0.172196f
C4617 commonsourceibias.n23 gnd 0.068706f
C4618 commonsourceibias.n24 gnd 0.046399f
C4619 commonsourceibias.t6 gnd 0.172196f
C4620 commonsourceibias.t34 gnd 0.194303f
C4621 commonsourceibias.n25 gnd 0.079733f
C4622 commonsourceibias.n26 gnd 0.082545f
C4623 commonsourceibias.n27 gnd 0.01136f
C4624 commonsourceibias.n28 gnd 0.012567f
C4625 commonsourceibias.n29 gnd 0.009217f
C4626 commonsourceibias.n30 gnd 0.009217f
C4627 commonsourceibias.n31 gnd 0.012485f
C4628 commonsourceibias.n32 gnd 0.007456f
C4629 commonsourceibias.n33 gnd 0.01264f
C4630 commonsourceibias.n34 gnd 0.009217f
C4631 commonsourceibias.n35 gnd 0.009217f
C4632 commonsourceibias.n36 gnd 0.012717f
C4633 commonsourceibias.n37 gnd 0.010966f
C4634 commonsourceibias.n38 gnd 0.008898f
C4635 commonsourceibias.n39 gnd 0.009217f
C4636 commonsourceibias.n40 gnd 0.009217f
C4637 commonsourceibias.n41 gnd 0.011274f
C4638 commonsourceibias.n42 gnd 0.012653f
C4639 commonsourceibias.n43 gnd 0.068706f
C4640 commonsourceibias.n44 gnd 0.012568f
C4641 commonsourceibias.n45 gnd 0.009217f
C4642 commonsourceibias.n46 gnd 0.009217f
C4643 commonsourceibias.n47 gnd 0.009217f
C4644 commonsourceibias.n48 gnd 0.012568f
C4645 commonsourceibias.n49 gnd 0.068706f
C4646 commonsourceibias.n50 gnd 0.012653f
C4647 commonsourceibias.n51 gnd 0.011274f
C4648 commonsourceibias.n52 gnd 0.009217f
C4649 commonsourceibias.n53 gnd 0.009217f
C4650 commonsourceibias.n54 gnd 0.009217f
C4651 commonsourceibias.n55 gnd 0.010966f
C4652 commonsourceibias.n56 gnd 0.012717f
C4653 commonsourceibias.n57 gnd 0.068706f
C4654 commonsourceibias.n58 gnd 0.01264f
C4655 commonsourceibias.n59 gnd 0.009217f
C4656 commonsourceibias.n60 gnd 0.009217f
C4657 commonsourceibias.n61 gnd 0.009217f
C4658 commonsourceibias.n62 gnd 0.012485f
C4659 commonsourceibias.n63 gnd 0.068706f
C4660 commonsourceibias.n64 gnd 0.012567f
C4661 commonsourceibias.n65 gnd 0.01136f
C4662 commonsourceibias.n66 gnd 0.009217f
C4663 commonsourceibias.n67 gnd 0.009217f
C4664 commonsourceibias.n68 gnd 0.009349f
C4665 commonsourceibias.n69 gnd 0.009666f
C4666 commonsourceibias.n70 gnd 0.082208f
C4667 commonsourceibias.n71 gnd 0.091197f
C4668 commonsourceibias.t17 gnd 0.019889f
C4669 commonsourceibias.t31 gnd 0.019889f
C4670 commonsourceibias.n72 gnd 0.175743f
C4671 commonsourceibias.n73 gnd 0.151855f
C4672 commonsourceibias.t3 gnd 0.019889f
C4673 commonsourceibias.t23 gnd 0.019889f
C4674 commonsourceibias.n74 gnd 0.175743f
C4675 commonsourceibias.n75 gnd 0.080726f
C4676 commonsourceibias.t43 gnd 0.019889f
C4677 commonsourceibias.t19 gnd 0.019889f
C4678 commonsourceibias.n76 gnd 0.175743f
C4679 commonsourceibias.n77 gnd 0.067443f
C4680 commonsourceibias.t7 gnd 0.019889f
C4681 commonsourceibias.t35 gnd 0.019889f
C4682 commonsourceibias.n78 gnd 0.176331f
C4683 commonsourceibias.t25 gnd 0.019889f
C4684 commonsourceibias.t45 gnd 0.019889f
C4685 commonsourceibias.n79 gnd 0.175743f
C4686 commonsourceibias.n80 gnd 0.16376f
C4687 commonsourceibias.t33 gnd 0.019889f
C4688 commonsourceibias.t41 gnd 0.019889f
C4689 commonsourceibias.n81 gnd 0.175743f
C4690 commonsourceibias.n82 gnd 0.067443f
C4691 commonsourceibias.n83 gnd 0.081666f
C4692 commonsourceibias.n84 gnd 0.009217f
C4693 commonsourceibias.t100 gnd 0.172196f
C4694 commonsourceibias.t87 gnd 0.172196f
C4695 commonsourceibias.n85 gnd 0.068706f
C4696 commonsourceibias.n86 gnd 0.009217f
C4697 commonsourceibias.t115 gnd 0.172196f
C4698 commonsourceibias.n87 gnd 0.068706f
C4699 commonsourceibias.n88 gnd 0.009217f
C4700 commonsourceibias.t79 gnd 0.172196f
C4701 commonsourceibias.n89 gnd 0.068706f
C4702 commonsourceibias.n90 gnd 0.046399f
C4703 commonsourceibias.t66 gnd 0.172196f
C4704 commonsourceibias.t95 gnd 0.194303f
C4705 commonsourceibias.n91 gnd 0.079733f
C4706 commonsourceibias.n92 gnd 0.082545f
C4707 commonsourceibias.n93 gnd 0.01136f
C4708 commonsourceibias.n94 gnd 0.012567f
C4709 commonsourceibias.n95 gnd 0.009217f
C4710 commonsourceibias.n96 gnd 0.009217f
C4711 commonsourceibias.n97 gnd 0.012485f
C4712 commonsourceibias.n98 gnd 0.007456f
C4713 commonsourceibias.n99 gnd 0.01264f
C4714 commonsourceibias.n100 gnd 0.009217f
C4715 commonsourceibias.n101 gnd 0.009217f
C4716 commonsourceibias.n102 gnd 0.012717f
C4717 commonsourceibias.n103 gnd 0.010966f
C4718 commonsourceibias.n104 gnd 0.008898f
C4719 commonsourceibias.n105 gnd 0.009217f
C4720 commonsourceibias.n106 gnd 0.009217f
C4721 commonsourceibias.n107 gnd 0.011274f
C4722 commonsourceibias.n108 gnd 0.012653f
C4723 commonsourceibias.n109 gnd 0.068706f
C4724 commonsourceibias.n110 gnd 0.012568f
C4725 commonsourceibias.n111 gnd 0.009172f
C4726 commonsourceibias.n112 gnd 0.066626f
C4727 commonsourceibias.n113 gnd 0.009172f
C4728 commonsourceibias.n114 gnd 0.012568f
C4729 commonsourceibias.n115 gnd 0.068706f
C4730 commonsourceibias.n116 gnd 0.012653f
C4731 commonsourceibias.n117 gnd 0.011274f
C4732 commonsourceibias.n118 gnd 0.009217f
C4733 commonsourceibias.n119 gnd 0.009217f
C4734 commonsourceibias.n120 gnd 0.009217f
C4735 commonsourceibias.n121 gnd 0.010966f
C4736 commonsourceibias.n122 gnd 0.012717f
C4737 commonsourceibias.n123 gnd 0.068706f
C4738 commonsourceibias.n124 gnd 0.01264f
C4739 commonsourceibias.n125 gnd 0.009217f
C4740 commonsourceibias.n126 gnd 0.009217f
C4741 commonsourceibias.n127 gnd 0.009217f
C4742 commonsourceibias.n128 gnd 0.012485f
C4743 commonsourceibias.n129 gnd 0.068706f
C4744 commonsourceibias.n130 gnd 0.012567f
C4745 commonsourceibias.n131 gnd 0.01136f
C4746 commonsourceibias.n132 gnd 0.009217f
C4747 commonsourceibias.n133 gnd 0.009217f
C4748 commonsourceibias.n134 gnd 0.009349f
C4749 commonsourceibias.n135 gnd 0.009666f
C4750 commonsourceibias.n136 gnd 0.082208f
C4751 commonsourceibias.n137 gnd 0.05322f
C4752 commonsourceibias.n138 gnd 0.012299f
C4753 commonsourceibias.t89 gnd 0.18623f
C4754 commonsourceibias.t106 gnd 0.172196f
C4755 commonsourceibias.n139 gnd 0.068706f
C4756 commonsourceibias.n140 gnd 0.009217f
C4757 commonsourceibias.t101 gnd 0.172196f
C4758 commonsourceibias.n141 gnd 0.007456f
C4759 commonsourceibias.n142 gnd 0.009217f
C4760 commonsourceibias.t88 gnd 0.172196f
C4761 commonsourceibias.n143 gnd 0.008898f
C4762 commonsourceibias.n144 gnd 0.009217f
C4763 commonsourceibias.t105 gnd 0.172196f
C4764 commonsourceibias.n145 gnd 0.068706f
C4765 commonsourceibias.t99 gnd 0.172196f
C4766 commonsourceibias.n146 gnd 0.007444f
C4767 commonsourceibias.n147 gnd 0.009217f
C4768 commonsourceibias.t86 gnd 0.172196f
C4769 commonsourceibias.t108 gnd 0.172196f
C4770 commonsourceibias.n148 gnd 0.068706f
C4771 commonsourceibias.n149 gnd 0.009217f
C4772 commonsourceibias.t98 gnd 0.172196f
C4773 commonsourceibias.n150 gnd 0.068706f
C4774 commonsourceibias.n151 gnd 0.009217f
C4775 commonsourceibias.t112 gnd 0.172196f
C4776 commonsourceibias.n152 gnd 0.068706f
C4777 commonsourceibias.n153 gnd 0.046399f
C4778 commonsourceibias.t107 gnd 0.172196f
C4779 commonsourceibias.t97 gnd 0.194303f
C4780 commonsourceibias.n154 gnd 0.079733f
C4781 commonsourceibias.n155 gnd 0.082545f
C4782 commonsourceibias.n156 gnd 0.01136f
C4783 commonsourceibias.n157 gnd 0.012567f
C4784 commonsourceibias.n158 gnd 0.009217f
C4785 commonsourceibias.n159 gnd 0.009217f
C4786 commonsourceibias.n160 gnd 0.012485f
C4787 commonsourceibias.n161 gnd 0.007456f
C4788 commonsourceibias.n162 gnd 0.01264f
C4789 commonsourceibias.n163 gnd 0.009217f
C4790 commonsourceibias.n164 gnd 0.009217f
C4791 commonsourceibias.n165 gnd 0.012717f
C4792 commonsourceibias.n166 gnd 0.010966f
C4793 commonsourceibias.n167 gnd 0.008898f
C4794 commonsourceibias.n168 gnd 0.009217f
C4795 commonsourceibias.n169 gnd 0.009217f
C4796 commonsourceibias.n170 gnd 0.011274f
C4797 commonsourceibias.n171 gnd 0.012653f
C4798 commonsourceibias.n172 gnd 0.068706f
C4799 commonsourceibias.n173 gnd 0.012568f
C4800 commonsourceibias.n174 gnd 0.009217f
C4801 commonsourceibias.n175 gnd 0.009217f
C4802 commonsourceibias.n176 gnd 0.009217f
C4803 commonsourceibias.n177 gnd 0.012568f
C4804 commonsourceibias.n178 gnd 0.068706f
C4805 commonsourceibias.n179 gnd 0.012653f
C4806 commonsourceibias.n180 gnd 0.011274f
C4807 commonsourceibias.n181 gnd 0.009217f
C4808 commonsourceibias.n182 gnd 0.009217f
C4809 commonsourceibias.n183 gnd 0.009217f
C4810 commonsourceibias.n184 gnd 0.010966f
C4811 commonsourceibias.n185 gnd 0.012717f
C4812 commonsourceibias.n186 gnd 0.068706f
C4813 commonsourceibias.n187 gnd 0.01264f
C4814 commonsourceibias.n188 gnd 0.009217f
C4815 commonsourceibias.n189 gnd 0.009217f
C4816 commonsourceibias.n190 gnd 0.009217f
C4817 commonsourceibias.n191 gnd 0.012485f
C4818 commonsourceibias.n192 gnd 0.068706f
C4819 commonsourceibias.n193 gnd 0.012567f
C4820 commonsourceibias.n194 gnd 0.01136f
C4821 commonsourceibias.n195 gnd 0.009217f
C4822 commonsourceibias.n196 gnd 0.009217f
C4823 commonsourceibias.n197 gnd 0.009349f
C4824 commonsourceibias.n198 gnd 0.009666f
C4825 commonsourceibias.n199 gnd 0.082208f
C4826 commonsourceibias.n200 gnd 0.027976f
C4827 commonsourceibias.n201 gnd 0.147064f
C4828 commonsourceibias.n202 gnd 0.012299f
C4829 commonsourceibias.t50 gnd 0.172196f
C4830 commonsourceibias.n203 gnd 0.068706f
C4831 commonsourceibias.n204 gnd 0.009217f
C4832 commonsourceibias.t60 gnd 0.172196f
C4833 commonsourceibias.n205 gnd 0.007456f
C4834 commonsourceibias.n206 gnd 0.009217f
C4835 commonsourceibias.t104 gnd 0.172196f
C4836 commonsourceibias.n207 gnd 0.008898f
C4837 commonsourceibias.n208 gnd 0.009217f
C4838 commonsourceibias.t118 gnd 0.172196f
C4839 commonsourceibias.n209 gnd 0.068706f
C4840 commonsourceibias.t52 gnd 0.172196f
C4841 commonsourceibias.n210 gnd 0.007444f
C4842 commonsourceibias.n211 gnd 0.009217f
C4843 commonsourceibias.t93 gnd 0.172196f
C4844 commonsourceibias.t84 gnd 0.172196f
C4845 commonsourceibias.n212 gnd 0.068706f
C4846 commonsourceibias.n213 gnd 0.009217f
C4847 commonsourceibias.t49 gnd 0.172196f
C4848 commonsourceibias.n214 gnd 0.068706f
C4849 commonsourceibias.n215 gnd 0.009217f
C4850 commonsourceibias.t59 gnd 0.172196f
C4851 commonsourceibias.n216 gnd 0.068706f
C4852 commonsourceibias.n217 gnd 0.046399f
C4853 commonsourceibias.t75 gnd 0.172196f
C4854 commonsourceibias.t117 gnd 0.194303f
C4855 commonsourceibias.n218 gnd 0.079733f
C4856 commonsourceibias.n219 gnd 0.082545f
C4857 commonsourceibias.n220 gnd 0.01136f
C4858 commonsourceibias.n221 gnd 0.012567f
C4859 commonsourceibias.n222 gnd 0.009217f
C4860 commonsourceibias.n223 gnd 0.009217f
C4861 commonsourceibias.n224 gnd 0.012485f
C4862 commonsourceibias.n225 gnd 0.007456f
C4863 commonsourceibias.n226 gnd 0.01264f
C4864 commonsourceibias.n227 gnd 0.009217f
C4865 commonsourceibias.n228 gnd 0.009217f
C4866 commonsourceibias.n229 gnd 0.012717f
C4867 commonsourceibias.n230 gnd 0.010966f
C4868 commonsourceibias.n231 gnd 0.008898f
C4869 commonsourceibias.n232 gnd 0.009217f
C4870 commonsourceibias.n233 gnd 0.009217f
C4871 commonsourceibias.n234 gnd 0.011274f
C4872 commonsourceibias.n235 gnd 0.012653f
C4873 commonsourceibias.n236 gnd 0.068706f
C4874 commonsourceibias.n237 gnd 0.012568f
C4875 commonsourceibias.n238 gnd 0.009217f
C4876 commonsourceibias.n239 gnd 0.009217f
C4877 commonsourceibias.n240 gnd 0.009217f
C4878 commonsourceibias.n241 gnd 0.012568f
C4879 commonsourceibias.n242 gnd 0.068706f
C4880 commonsourceibias.n243 gnd 0.012653f
C4881 commonsourceibias.n244 gnd 0.011274f
C4882 commonsourceibias.n245 gnd 0.009217f
C4883 commonsourceibias.n246 gnd 0.009217f
C4884 commonsourceibias.n247 gnd 0.009217f
C4885 commonsourceibias.n248 gnd 0.010966f
C4886 commonsourceibias.n249 gnd 0.012717f
C4887 commonsourceibias.n250 gnd 0.068706f
C4888 commonsourceibias.n251 gnd 0.01264f
C4889 commonsourceibias.n252 gnd 0.009217f
C4890 commonsourceibias.n253 gnd 0.009217f
C4891 commonsourceibias.n254 gnd 0.009217f
C4892 commonsourceibias.n255 gnd 0.012485f
C4893 commonsourceibias.n256 gnd 0.068706f
C4894 commonsourceibias.n257 gnd 0.012567f
C4895 commonsourceibias.n258 gnd 0.01136f
C4896 commonsourceibias.n259 gnd 0.009217f
C4897 commonsourceibias.n260 gnd 0.009217f
C4898 commonsourceibias.n261 gnd 0.009349f
C4899 commonsourceibias.n262 gnd 0.009666f
C4900 commonsourceibias.t111 gnd 0.18623f
C4901 commonsourceibias.n263 gnd 0.082208f
C4902 commonsourceibias.n264 gnd 0.027976f
C4903 commonsourceibias.n265 gnd 0.517265f
C4904 commonsourceibias.n266 gnd 0.012299f
C4905 commonsourceibias.t114 gnd 0.18623f
C4906 commonsourceibias.t78 gnd 0.172196f
C4907 commonsourceibias.n267 gnd 0.068706f
C4908 commonsourceibias.n268 gnd 0.009217f
C4909 commonsourceibias.t53 gnd 0.172196f
C4910 commonsourceibias.n269 gnd 0.007456f
C4911 commonsourceibias.n270 gnd 0.009217f
C4912 commonsourceibias.t94 gnd 0.172196f
C4913 commonsourceibias.n271 gnd 0.008898f
C4914 commonsourceibias.n272 gnd 0.009217f
C4915 commonsourceibias.t113 gnd 0.172196f
C4916 commonsourceibias.n273 gnd 0.007444f
C4917 commonsourceibias.n274 gnd 0.009217f
C4918 commonsourceibias.t76 gnd 0.172196f
C4919 commonsourceibias.t65 gnd 0.172196f
C4920 commonsourceibias.n275 gnd 0.068706f
C4921 commonsourceibias.n276 gnd 0.009217f
C4922 commonsourceibias.t92 gnd 0.172196f
C4923 commonsourceibias.n277 gnd 0.068706f
C4924 commonsourceibias.n278 gnd 0.009217f
C4925 commonsourceibias.t63 gnd 0.172196f
C4926 commonsourceibias.n279 gnd 0.068706f
C4927 commonsourceibias.n280 gnd 0.046399f
C4928 commonsourceibias.t58 gnd 0.172196f
C4929 commonsourceibias.t70 gnd 0.194303f
C4930 commonsourceibias.n281 gnd 0.079733f
C4931 commonsourceibias.n282 gnd 0.082545f
C4932 commonsourceibias.n283 gnd 0.01136f
C4933 commonsourceibias.n284 gnd 0.012567f
C4934 commonsourceibias.n285 gnd 0.009217f
C4935 commonsourceibias.n286 gnd 0.009217f
C4936 commonsourceibias.n287 gnd 0.012485f
C4937 commonsourceibias.n288 gnd 0.007456f
C4938 commonsourceibias.n289 gnd 0.01264f
C4939 commonsourceibias.n290 gnd 0.009217f
C4940 commonsourceibias.n291 gnd 0.009217f
C4941 commonsourceibias.n292 gnd 0.012717f
C4942 commonsourceibias.n293 gnd 0.010966f
C4943 commonsourceibias.n294 gnd 0.008898f
C4944 commonsourceibias.n295 gnd 0.009217f
C4945 commonsourceibias.n296 gnd 0.009217f
C4946 commonsourceibias.n297 gnd 0.011274f
C4947 commonsourceibias.n298 gnd 0.012653f
C4948 commonsourceibias.n299 gnd 0.068706f
C4949 commonsourceibias.n300 gnd 0.012568f
C4950 commonsourceibias.n301 gnd 0.009172f
C4951 commonsourceibias.t5 gnd 0.019889f
C4952 commonsourceibias.t15 gnd 0.019889f
C4953 commonsourceibias.n302 gnd 0.176331f
C4954 commonsourceibias.t13 gnd 0.019889f
C4955 commonsourceibias.t39 gnd 0.019889f
C4956 commonsourceibias.n303 gnd 0.175743f
C4957 commonsourceibias.n304 gnd 0.16376f
C4958 commonsourceibias.t9 gnd 0.019889f
C4959 commonsourceibias.t1 gnd 0.019889f
C4960 commonsourceibias.n305 gnd 0.175743f
C4961 commonsourceibias.n306 gnd 0.067443f
C4962 commonsourceibias.n307 gnd 0.012299f
C4963 commonsourceibias.t46 gnd 0.172196f
C4964 commonsourceibias.n308 gnd 0.068706f
C4965 commonsourceibias.n309 gnd 0.009217f
C4966 commonsourceibias.t20 gnd 0.172196f
C4967 commonsourceibias.n310 gnd 0.007456f
C4968 commonsourceibias.n311 gnd 0.009217f
C4969 commonsourceibias.t36 gnd 0.172196f
C4970 commonsourceibias.n312 gnd 0.008898f
C4971 commonsourceibias.n313 gnd 0.009217f
C4972 commonsourceibias.t28 gnd 0.172196f
C4973 commonsourceibias.n314 gnd 0.007444f
C4974 commonsourceibias.n315 gnd 0.009217f
C4975 commonsourceibias.t0 gnd 0.172196f
C4976 commonsourceibias.t8 gnd 0.172196f
C4977 commonsourceibias.n316 gnd 0.068706f
C4978 commonsourceibias.n317 gnd 0.009217f
C4979 commonsourceibias.t38 gnd 0.172196f
C4980 commonsourceibias.n318 gnd 0.068706f
C4981 commonsourceibias.n319 gnd 0.009217f
C4982 commonsourceibias.t12 gnd 0.172196f
C4983 commonsourceibias.n320 gnd 0.068706f
C4984 commonsourceibias.n321 gnd 0.046399f
C4985 commonsourceibias.t14 gnd 0.172196f
C4986 commonsourceibias.t4 gnd 0.194303f
C4987 commonsourceibias.n322 gnd 0.079733f
C4988 commonsourceibias.n323 gnd 0.082545f
C4989 commonsourceibias.n324 gnd 0.01136f
C4990 commonsourceibias.n325 gnd 0.012567f
C4991 commonsourceibias.n326 gnd 0.009217f
C4992 commonsourceibias.n327 gnd 0.009217f
C4993 commonsourceibias.n328 gnd 0.012485f
C4994 commonsourceibias.n329 gnd 0.007456f
C4995 commonsourceibias.n330 gnd 0.01264f
C4996 commonsourceibias.n331 gnd 0.009217f
C4997 commonsourceibias.n332 gnd 0.009217f
C4998 commonsourceibias.n333 gnd 0.012717f
C4999 commonsourceibias.n334 gnd 0.010966f
C5000 commonsourceibias.n335 gnd 0.008898f
C5001 commonsourceibias.n336 gnd 0.009217f
C5002 commonsourceibias.n337 gnd 0.009217f
C5003 commonsourceibias.n338 gnd 0.011274f
C5004 commonsourceibias.n339 gnd 0.012653f
C5005 commonsourceibias.n340 gnd 0.068706f
C5006 commonsourceibias.n341 gnd 0.012568f
C5007 commonsourceibias.n342 gnd 0.009217f
C5008 commonsourceibias.n343 gnd 0.009217f
C5009 commonsourceibias.n344 gnd 0.009217f
C5010 commonsourceibias.n345 gnd 0.012568f
C5011 commonsourceibias.n346 gnd 0.068706f
C5012 commonsourceibias.n347 gnd 0.012653f
C5013 commonsourceibias.t10 gnd 0.172196f
C5014 commonsourceibias.n348 gnd 0.068706f
C5015 commonsourceibias.n349 gnd 0.011274f
C5016 commonsourceibias.n350 gnd 0.009217f
C5017 commonsourceibias.n351 gnd 0.009217f
C5018 commonsourceibias.n352 gnd 0.009217f
C5019 commonsourceibias.n353 gnd 0.010966f
C5020 commonsourceibias.n354 gnd 0.012717f
C5021 commonsourceibias.n355 gnd 0.068706f
C5022 commonsourceibias.n356 gnd 0.01264f
C5023 commonsourceibias.n357 gnd 0.009217f
C5024 commonsourceibias.n358 gnd 0.009217f
C5025 commonsourceibias.n359 gnd 0.009217f
C5026 commonsourceibias.n360 gnd 0.012485f
C5027 commonsourceibias.n361 gnd 0.068706f
C5028 commonsourceibias.n362 gnd 0.012567f
C5029 commonsourceibias.n363 gnd 0.01136f
C5030 commonsourceibias.n364 gnd 0.009217f
C5031 commonsourceibias.n365 gnd 0.009217f
C5032 commonsourceibias.n366 gnd 0.009349f
C5033 commonsourceibias.n367 gnd 0.009666f
C5034 commonsourceibias.t26 gnd 0.18623f
C5035 commonsourceibias.n368 gnd 0.082208f
C5036 commonsourceibias.n369 gnd 0.091197f
C5037 commonsourceibias.t47 gnd 0.019889f
C5038 commonsourceibias.t27 gnd 0.019889f
C5039 commonsourceibias.n370 gnd 0.175743f
C5040 commonsourceibias.n371 gnd 0.151855f
C5041 commonsourceibias.t37 gnd 0.019889f
C5042 commonsourceibias.t21 gnd 0.019889f
C5043 commonsourceibias.n372 gnd 0.175743f
C5044 commonsourceibias.n373 gnd 0.080726f
C5045 commonsourceibias.t29 gnd 0.019889f
C5046 commonsourceibias.t11 gnd 0.019889f
C5047 commonsourceibias.n374 gnd 0.175743f
C5048 commonsourceibias.n375 gnd 0.067443f
C5049 commonsourceibias.n376 gnd 0.081666f
C5050 commonsourceibias.n377 gnd 0.066626f
C5051 commonsourceibias.n378 gnd 0.009172f
C5052 commonsourceibias.n379 gnd 0.012568f
C5053 commonsourceibias.n380 gnd 0.068706f
C5054 commonsourceibias.n381 gnd 0.012653f
C5055 commonsourceibias.t64 gnd 0.172196f
C5056 commonsourceibias.n382 gnd 0.068706f
C5057 commonsourceibias.n383 gnd 0.011274f
C5058 commonsourceibias.n384 gnd 0.009217f
C5059 commonsourceibias.n385 gnd 0.009217f
C5060 commonsourceibias.n386 gnd 0.009217f
C5061 commonsourceibias.n387 gnd 0.010966f
C5062 commonsourceibias.n388 gnd 0.012717f
C5063 commonsourceibias.n389 gnd 0.068706f
C5064 commonsourceibias.n390 gnd 0.01264f
C5065 commonsourceibias.n391 gnd 0.009217f
C5066 commonsourceibias.n392 gnd 0.009217f
C5067 commonsourceibias.n393 gnd 0.009217f
C5068 commonsourceibias.n394 gnd 0.012485f
C5069 commonsourceibias.n395 gnd 0.068706f
C5070 commonsourceibias.n396 gnd 0.012567f
C5071 commonsourceibias.n397 gnd 0.01136f
C5072 commonsourceibias.n398 gnd 0.009217f
C5073 commonsourceibias.n399 gnd 0.009217f
C5074 commonsourceibias.n400 gnd 0.009349f
C5075 commonsourceibias.n401 gnd 0.009666f
C5076 commonsourceibias.n402 gnd 0.082208f
C5077 commonsourceibias.n403 gnd 0.05322f
C5078 commonsourceibias.n404 gnd 0.012299f
C5079 commonsourceibias.t91 gnd 0.172196f
C5080 commonsourceibias.n405 gnd 0.068706f
C5081 commonsourceibias.n406 gnd 0.009217f
C5082 commonsourceibias.t83 gnd 0.172196f
C5083 commonsourceibias.n407 gnd 0.007456f
C5084 commonsourceibias.n408 gnd 0.009217f
C5085 commonsourceibias.t73 gnd 0.172196f
C5086 commonsourceibias.n409 gnd 0.008898f
C5087 commonsourceibias.n410 gnd 0.009217f
C5088 commonsourceibias.t82 gnd 0.172196f
C5089 commonsourceibias.n411 gnd 0.007444f
C5090 commonsourceibias.n412 gnd 0.009217f
C5091 commonsourceibias.t103 gnd 0.172196f
C5092 commonsourceibias.t96 gnd 0.172196f
C5093 commonsourceibias.n413 gnd 0.068706f
C5094 commonsourceibias.n414 gnd 0.009217f
C5095 commonsourceibias.t81 gnd 0.172196f
C5096 commonsourceibias.n415 gnd 0.068706f
C5097 commonsourceibias.n416 gnd 0.009217f
C5098 commonsourceibias.t102 gnd 0.172196f
C5099 commonsourceibias.n417 gnd 0.068706f
C5100 commonsourceibias.n418 gnd 0.046399f
C5101 commonsourceibias.t116 gnd 0.172196f
C5102 commonsourceibias.t80 gnd 0.194303f
C5103 commonsourceibias.n419 gnd 0.079733f
C5104 commonsourceibias.n420 gnd 0.082545f
C5105 commonsourceibias.n421 gnd 0.01136f
C5106 commonsourceibias.n422 gnd 0.012567f
C5107 commonsourceibias.n423 gnd 0.009217f
C5108 commonsourceibias.n424 gnd 0.009217f
C5109 commonsourceibias.n425 gnd 0.012485f
C5110 commonsourceibias.n426 gnd 0.007456f
C5111 commonsourceibias.n427 gnd 0.01264f
C5112 commonsourceibias.n428 gnd 0.009217f
C5113 commonsourceibias.n429 gnd 0.009217f
C5114 commonsourceibias.n430 gnd 0.012717f
C5115 commonsourceibias.n431 gnd 0.010966f
C5116 commonsourceibias.n432 gnd 0.008898f
C5117 commonsourceibias.n433 gnd 0.009217f
C5118 commonsourceibias.n434 gnd 0.009217f
C5119 commonsourceibias.n435 gnd 0.011274f
C5120 commonsourceibias.n436 gnd 0.012653f
C5121 commonsourceibias.n437 gnd 0.068706f
C5122 commonsourceibias.n438 gnd 0.012568f
C5123 commonsourceibias.n439 gnd 0.009217f
C5124 commonsourceibias.n440 gnd 0.009217f
C5125 commonsourceibias.n441 gnd 0.009217f
C5126 commonsourceibias.n442 gnd 0.012568f
C5127 commonsourceibias.n443 gnd 0.068706f
C5128 commonsourceibias.n444 gnd 0.012653f
C5129 commonsourceibias.t90 gnd 0.172196f
C5130 commonsourceibias.n445 gnd 0.068706f
C5131 commonsourceibias.n446 gnd 0.011274f
C5132 commonsourceibias.n447 gnd 0.009217f
C5133 commonsourceibias.n448 gnd 0.009217f
C5134 commonsourceibias.n449 gnd 0.009217f
C5135 commonsourceibias.n450 gnd 0.010966f
C5136 commonsourceibias.n451 gnd 0.012717f
C5137 commonsourceibias.n452 gnd 0.068706f
C5138 commonsourceibias.n453 gnd 0.01264f
C5139 commonsourceibias.n454 gnd 0.009217f
C5140 commonsourceibias.n455 gnd 0.009217f
C5141 commonsourceibias.n456 gnd 0.009217f
C5142 commonsourceibias.n457 gnd 0.012485f
C5143 commonsourceibias.n458 gnd 0.068706f
C5144 commonsourceibias.n459 gnd 0.012567f
C5145 commonsourceibias.n460 gnd 0.01136f
C5146 commonsourceibias.n461 gnd 0.009217f
C5147 commonsourceibias.n462 gnd 0.009217f
C5148 commonsourceibias.n463 gnd 0.009349f
C5149 commonsourceibias.n464 gnd 0.009666f
C5150 commonsourceibias.t74 gnd 0.18623f
C5151 commonsourceibias.n465 gnd 0.082208f
C5152 commonsourceibias.n466 gnd 0.027976f
C5153 commonsourceibias.n467 gnd 0.147064f
C5154 commonsourceibias.n468 gnd 0.012299f
C5155 commonsourceibias.t62 gnd 0.172196f
C5156 commonsourceibias.n469 gnd 0.068706f
C5157 commonsourceibias.n470 gnd 0.009217f
C5158 commonsourceibias.t71 gnd 0.172196f
C5159 commonsourceibias.n471 gnd 0.007456f
C5160 commonsourceibias.n472 gnd 0.009217f
C5161 commonsourceibias.t48 gnd 0.172196f
C5162 commonsourceibias.n473 gnd 0.008898f
C5163 commonsourceibias.n474 gnd 0.009217f
C5164 commonsourceibias.t67 gnd 0.172196f
C5165 commonsourceibias.n475 gnd 0.007444f
C5166 commonsourceibias.n476 gnd 0.009217f
C5167 commonsourceibias.t77 gnd 0.172196f
C5168 commonsourceibias.t110 gnd 0.172196f
C5169 commonsourceibias.n477 gnd 0.068706f
C5170 commonsourceibias.n478 gnd 0.009217f
C5171 commonsourceibias.t61 gnd 0.172196f
C5172 commonsourceibias.n479 gnd 0.068706f
C5173 commonsourceibias.n480 gnd 0.009217f
C5174 commonsourceibias.t72 gnd 0.172196f
C5175 commonsourceibias.n481 gnd 0.068706f
C5176 commonsourceibias.n482 gnd 0.046399f
C5177 commonsourceibias.t68 gnd 0.172196f
C5178 commonsourceibias.t55 gnd 0.194303f
C5179 commonsourceibias.n483 gnd 0.079733f
C5180 commonsourceibias.n484 gnd 0.082545f
C5181 commonsourceibias.n485 gnd 0.01136f
C5182 commonsourceibias.n486 gnd 0.012567f
C5183 commonsourceibias.n487 gnd 0.009217f
C5184 commonsourceibias.n488 gnd 0.009217f
C5185 commonsourceibias.n489 gnd 0.012485f
C5186 commonsourceibias.n490 gnd 0.007456f
C5187 commonsourceibias.n491 gnd 0.01264f
C5188 commonsourceibias.n492 gnd 0.009217f
C5189 commonsourceibias.n493 gnd 0.009217f
C5190 commonsourceibias.n494 gnd 0.012717f
C5191 commonsourceibias.n495 gnd 0.010966f
C5192 commonsourceibias.n496 gnd 0.008898f
C5193 commonsourceibias.n497 gnd 0.009217f
C5194 commonsourceibias.n498 gnd 0.009217f
C5195 commonsourceibias.n499 gnd 0.011274f
C5196 commonsourceibias.n500 gnd 0.012653f
C5197 commonsourceibias.n501 gnd 0.068706f
C5198 commonsourceibias.n502 gnd 0.012568f
C5199 commonsourceibias.n503 gnd 0.009217f
C5200 commonsourceibias.n504 gnd 0.009217f
C5201 commonsourceibias.n505 gnd 0.009217f
C5202 commonsourceibias.n506 gnd 0.012568f
C5203 commonsourceibias.n507 gnd 0.068706f
C5204 commonsourceibias.n508 gnd 0.012653f
C5205 commonsourceibias.t57 gnd 0.172196f
C5206 commonsourceibias.n509 gnd 0.068706f
C5207 commonsourceibias.n510 gnd 0.011274f
C5208 commonsourceibias.n511 gnd 0.009217f
C5209 commonsourceibias.n512 gnd 0.009217f
C5210 commonsourceibias.n513 gnd 0.009217f
C5211 commonsourceibias.n514 gnd 0.010966f
C5212 commonsourceibias.n515 gnd 0.012717f
C5213 commonsourceibias.n516 gnd 0.068706f
C5214 commonsourceibias.n517 gnd 0.01264f
C5215 commonsourceibias.n518 gnd 0.009217f
C5216 commonsourceibias.n519 gnd 0.009217f
C5217 commonsourceibias.n520 gnd 0.009217f
C5218 commonsourceibias.n521 gnd 0.012485f
C5219 commonsourceibias.n522 gnd 0.068706f
C5220 commonsourceibias.n523 gnd 0.012567f
C5221 commonsourceibias.n524 gnd 0.01136f
C5222 commonsourceibias.n525 gnd 0.009217f
C5223 commonsourceibias.n526 gnd 0.009217f
C5224 commonsourceibias.n527 gnd 0.009349f
C5225 commonsourceibias.n528 gnd 0.009666f
C5226 commonsourceibias.t51 gnd 0.18623f
C5227 commonsourceibias.n529 gnd 0.082208f
C5228 commonsourceibias.n530 gnd 0.027976f
C5229 commonsourceibias.n531 gnd 0.194274f
C5230 commonsourceibias.n532 gnd 5.09694f
.ends

