* NGSPICE file created from opamp.ext - technology: sky130A

.subckt opamp CSoutput output vdd plus minus commonsourceibias outputibias diffpairibias
+ gnd
X0 gnd.t312 gnd.t309 gnd.t311 gnd.t310 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X1 gnd.t324 commonsourceibias.t46 commonsourceibias.t47 gnd.t123 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X2 vdd.t129 vdd.t127 vdd.t128 vdd.t115 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X3 vdd.t190 a_n6308_8799.t36 CSoutput.t143 vdd.t187 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X4 a_n1986_8322.t23 a_n2848_n452.t48 vdd.t160 vdd.t159 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X5 a_n1808_13878.t11 a_n2848_n452.t24 a_n2848_n452.t25 vdd.t9 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X6 a_n6308_8799.t11 plus.t5 a_n3827_n3924.t38 gnd.t110 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X7 commonsourceibias.t45 commonsourceibias.t44 gnd.t135 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 a_n3827_n3924.t37 plus.t6 a_n6308_8799.t28 gnd.t85 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X9 a_n3827_n3924.t0 diffpairibias.t20 gnd.t2 gnd.t1 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X10 a_n2848_n452.t33 a_n2848_n452.t32 a_n1808_13878.t10 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X11 a_n1808_13878.t9 a_n2848_n452.t30 a_n2848_n452.t31 vdd.t34 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X12 vdd.t126 vdd.t124 vdd.t125 vdd.t98 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X13 CSoutput.t142 a_n6308_8799.t37 vdd.t191 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X14 a_n1808_13878.t19 a_n2848_n452.t49 vdd.t162 vdd.t161 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X15 vdd.t123 vdd.t121 vdd.t122 vdd.t115 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X16 vdd.t120 vdd.t118 vdd.t119 vdd.t66 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X17 CSoutput.t141 a_n6308_8799.t38 vdd.t148 vdd.t147 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X18 gnd.t63 commonsourceibias.t42 commonsourceibias.t43 gnd.t62 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X19 gnd.t84 commonsourceibias.t48 CSoutput.t71 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X20 commonsourceibias.t41 commonsourceibias.t40 gnd.t120 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X21 CSoutput.t140 a_n6308_8799.t39 vdd.t150 vdd.t149 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X22 output.t3 outputibias.t8 gnd.t332 gnd.t331 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X23 gnd.t308 gnd.t306 gnd.t307 gnd.t243 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X24 a_n1986_8322.t15 a_n2848_n452.t50 a_n6308_8799.t7 vdd.t151 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X25 a_n2848_n452.t46 minus.t5 a_n3827_n3924.t55 gnd.t315 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X26 a_n6308_8799.t30 plus.t7 a_n3827_n3924.t36 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X27 plus.t4 gnd.t303 gnd.t305 gnd.t304 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X28 a_n2848_n452.t8 minus.t6 a_n3827_n3924.t10 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X29 commonsourceibias.t39 commonsourceibias.t38 gnd.t187 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X30 gnd.t319 commonsourceibias.t49 CSoutput.t70 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X31 CSoutput.t69 commonsourceibias.t50 gnd.t325 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 gnd.t302 gnd.t299 gnd.t301 gnd.t300 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X33 CSoutput.t139 a_n6308_8799.t40 vdd.t24 vdd.t23 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X34 vdd.t26 a_n6308_8799.t41 CSoutput.t138 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X35 a_n3827_n3924.t35 plus.t8 a_n6308_8799.t33 gnd.t92 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X36 gnd.t101 commonsourceibias.t36 commonsourceibias.t37 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X37 a_n6308_8799.t8 a_n2848_n452.t51 a_n1986_8322.t14 vdd.t9 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X38 CSoutput.t137 a_n6308_8799.t42 vdd.t43 vdd.t42 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X39 vdd.t45 a_n6308_8799.t43 CSoutput.t136 vdd.t44 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X40 a_n3827_n3924.t9 minus.t7 a_n2848_n452.t7 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X41 a_n3827_n3924.t51 diffpairibias.t21 gnd.t154 gnd.t153 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X42 commonsourceibias.t35 commonsourceibias.t34 gnd.t125 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X43 vdd.t117 vdd.t114 vdd.t116 vdd.t115 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X44 CSoutput.t135 a_n6308_8799.t44 vdd.t31 vdd.t30 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X45 CSoutput.t134 a_n6308_8799.t45 vdd.t33 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X46 vdd.t113 vdd.t111 vdd.t112 vdd.t55 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X47 CSoutput.t68 commonsourceibias.t51 gnd.t320 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X48 gnd.t100 commonsourceibias.t32 commonsourceibias.t33 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X49 output.t19 CSoutput.t144 vdd.t189 gnd.t147 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X50 gnd.t298 gnd.t296 gnd.t297 gnd.t232 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X51 output.t2 outputibias.t9 gnd.t12 gnd.t11 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X52 CSoutput.t133 a_n6308_8799.t46 vdd.t204 vdd.t149 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X53 a_n3827_n3924.t34 plus.t9 a_n6308_8799.t12 gnd.t91 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X54 a_n1808_13878.t8 a_n2848_n452.t18 a_n2848_n452.t19 vdd.t38 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X55 vdd.t205 a_n6308_8799.t47 CSoutput.t132 vdd.t44 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X56 a_n3827_n3924.t33 plus.t10 a_n6308_8799.t19 gnd.t93 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X57 a_n3827_n3924.t47 minus.t8 a_n2848_n452.t42 gnd.t111 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X58 diffpairibias.t19 diffpairibias.t18 gnd.t137 gnd.t136 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X59 a_n2848_n452.t29 a_n2848_n452.t28 a_n1808_13878.t7 vdd.t146 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X60 CSoutput.t131 a_n6308_8799.t48 vdd.t133 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X61 vdd.t110 vdd.t108 vdd.t109 vdd.t83 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X62 CSoutput.t67 commonsourceibias.t52 gnd.t179 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X63 gnd.t295 gnd.t293 gnd.t294 gnd.t207 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X64 CSoutput.t66 commonsourceibias.t53 gnd.t142 gnd.t132 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X65 diffpairibias.t17 diffpairibias.t16 gnd.t317 gnd.t316 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X66 gnd.t292 gnd.t290 gnd.t291 gnd.t207 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X67 CSoutput.t145 a_n1986_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X68 vdd.t134 a_n6308_8799.t49 CSoutput.t130 vdd.t44 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X69 CSoutput.t65 commonsourceibias.t54 gnd.t327 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X70 vdd.t194 a_n6308_8799.t50 CSoutput.t129 vdd.t28 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X71 CSoutput.t128 a_n6308_8799.t51 vdd.t195 vdd.t42 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X72 a_n3827_n3924.t3 minus.t9 a_n2848_n452.t2 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X73 a_n3827_n3924.t32 plus.t11 a_n6308_8799.t9 gnd.t29 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X74 gnd.t169 commonsourceibias.t55 CSoutput.t64 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X75 vdd.t206 a_n6308_8799.t52 CSoutput.t127 vdd.t178 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X76 gnd.t27 commonsourceibias.t56 CSoutput.t63 gnd.t26 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X77 a_n6308_8799.t14 plus.t12 a_n3827_n3924.t31 gnd.t89 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X78 CSoutput.t62 commonsourceibias.t57 gnd.t170 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X79 CSoutput.t146 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X80 gnd.t289 gnd.t287 gnd.t288 gnd.t243 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X81 CSoutput.t126 a_n6308_8799.t53 vdd.t207 vdd.t30 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X82 CSoutput.t125 a_n6308_8799.t54 vdd.t36 vdd.t35 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X83 output.t18 CSoutput.t147 vdd.t8 gnd.t23 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X84 a_n3827_n3924.t45 diffpairibias.t22 gnd.t95 gnd.t94 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X85 CSoutput.t124 a_n6308_8799.t55 vdd.t37 vdd.t35 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 a_n3827_n3924.t30 plus.t13 a_n6308_8799.t10 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X87 CSoutput.t61 commonsourceibias.t58 gnd.t174 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 vdd.t136 a_n6308_8799.t56 CSoutput.t123 vdd.t39 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X89 outputibias.t7 outputibias.t6 gnd.t150 gnd.t149 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X90 a_n2848_n452.t23 a_n2848_n452.t22 a_n1808_13878.t6 vdd.t151 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X91 CSoutput.t60 commonsourceibias.t59 gnd.t191 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X92 gnd.t72 commonsourceibias.t60 CSoutput.t59 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X93 commonsourceibias.t31 commonsourceibias.t30 gnd.t35 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 a_n2848_n452.t11 a_n2848_n452.t10 a_n1808_13878.t5 vdd.t15 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X95 vdd.t137 a_n6308_8799.t57 CSoutput.t122 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X96 vdd.t139 a_n6308_8799.t58 CSoutput.t121 vdd.t138 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X97 a_n6308_8799.t6 a_n2848_n452.t52 a_n1986_8322.t13 vdd.t143 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X98 gnd.t286 gnd.t284 gnd.t285 gnd.t236 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X99 vdd.t140 a_n6308_8799.t59 CSoutput.t120 vdd.t39 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X100 a_n2848_n452.t6 minus.t10 a_n3827_n3924.t8 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X101 diffpairibias.t15 diffpairibias.t14 gnd.t97 gnd.t96 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X102 outputibias.t5 outputibias.t4 gnd.t74 gnd.t73 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X103 vdd.t202 a_n6308_8799.t60 CSoutput.t119 vdd.t46 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X104 CSoutput.t118 a_n6308_8799.t61 vdd.t203 vdd.t48 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X105 vdd.t141 a_n6308_8799.t62 CSoutput.t117 vdd.t28 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X106 vdd.t107 vdd.t105 vdd.t106 vdd.t91 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X107 CSoutput.t58 commonsourceibias.t61 gnd.t129 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 gnd.t88 commonsourceibias.t28 commonsourceibias.t29 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X109 vdd.t104 vdd.t101 vdd.t103 vdd.t102 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X110 gnd.t183 commonsourceibias.t62 CSoutput.t57 gnd.t123 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X111 output.t17 CSoutput.t148 vdd.t10 gnd.t38 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X112 a_n3827_n3924.t52 diffpairibias.t23 gnd.t159 gnd.t158 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X113 vdd.t100 vdd.t97 vdd.t99 vdd.t98 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X114 gnd.t283 gnd.t281 minus.t4 gnd.t282 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X115 gnd.t280 gnd.t278 gnd.t279 gnd.t222 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X116 vdd.t11 CSoutput.t149 output.t16 gnd.t39 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X117 vdd.t145 a_n2848_n452.t53 a_n1986_8322.t22 vdd.t144 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X118 vdd.t96 vdd.t94 vdd.t95 vdd.t87 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X119 commonsourceibias.t27 commonsourceibias.t26 gnd.t143 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X120 gnd.t37 commonsourceibias.t63 CSoutput.t56 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X121 CSoutput.t116 a_n6308_8799.t63 vdd.t142 vdd.t35 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X122 a_n1986_8322.t21 a_n2848_n452.t54 vdd.t164 vdd.t163 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X123 gnd.t277 gnd.t275 gnd.t276 gnd.t194 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X124 gnd.t335 commonsourceibias.t24 commonsourceibias.t25 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X125 gnd.t274 gnd.t272 gnd.t273 gnd.t236 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X126 vdd.t40 a_n6308_8799.t64 CSoutput.t115 vdd.t39 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X127 vdd.t12 CSoutput.t150 output.t15 gnd.t40 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X128 vdd.t166 a_n2848_n452.t55 a_n1808_13878.t18 vdd.t165 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X129 gnd.t271 gnd.t269 plus.t3 gnd.t270 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X130 CSoutput.t55 commonsourceibias.t64 gnd.t122 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X131 a_n2848_n452.t9 minus.t11 a_n3827_n3924.t11 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X132 a_n6308_8799.t31 plus.t14 a_n3827_n3924.t29 gnd.t145 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X133 gnd.t146 commonsourceibias.t65 CSoutput.t54 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X134 commonsourceibias.t23 commonsourceibias.t22 gnd.t156 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X135 vdd.t93 vdd.t90 vdd.t92 vdd.t91 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X136 a_n6308_8799.t13 plus.t15 a_n3827_n3924.t28 gnd.t90 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X137 a_n2848_n452.t45 minus.t12 a_n3827_n3924.t54 gnd.t164 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X138 diffpairibias.t13 diffpairibias.t12 gnd.t33 gnd.t32 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X139 vdd.t89 vdd.t86 vdd.t88 vdd.t87 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X140 vdd.t41 a_n6308_8799.t65 CSoutput.t114 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X141 a_n6308_8799.t29 a_n2848_n452.t56 a_n1986_8322.t12 vdd.t219 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X142 a_n1986_8322.t20 a_n2848_n452.t57 vdd.t221 vdd.t220 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X143 vdd.t85 vdd.t82 vdd.t84 vdd.t83 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X144 vdd.t47 a_n6308_8799.t66 CSoutput.t113 vdd.t46 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X145 a_n2848_n452.t15 a_n2848_n452.t14 a_n1808_13878.t4 vdd.t132 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X146 gnd.t10 commonsourceibias.t66 CSoutput.t53 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X147 a_n3827_n3924.t7 minus.t13 a_n2848_n452.t5 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X148 gnd.t321 commonsourceibias.t67 CSoutput.t52 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X149 CSoutput.t112 a_n6308_8799.t67 vdd.t49 vdd.t48 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X150 a_n6308_8799.t32 a_n2848_n452.t58 a_n1986_8322.t11 vdd.t34 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X151 vdd.t0 CSoutput.t151 output.t14 gnd.t3 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X152 a_n1808_13878.t3 a_n2848_n452.t26 a_n2848_n452.t27 vdd.t143 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X153 a_n3827_n3924.t27 plus.t16 a_n6308_8799.t26 gnd.t314 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X154 a_n2848_n452.t44 minus.t14 a_n3827_n3924.t53 gnd.t110 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X155 output.t13 CSoutput.t152 vdd.t1 gnd.t4 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X156 gnd.t268 gnd.t266 gnd.t267 gnd.t243 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X157 CSoutput.t51 commonsourceibias.t68 gnd.t160 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X158 vdd.t227 a_n2848_n452.t59 a_n1986_8322.t19 vdd.t226 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X159 gnd.t330 commonsourceibias.t69 CSoutput.t50 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X160 output.t12 CSoutput.t153 vdd.t2 gnd.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X161 gnd.t20 commonsourceibias.t70 CSoutput.t49 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X162 a_n3827_n3924.t49 diffpairibias.t24 gnd.t117 gnd.t116 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X163 CSoutput.t111 a_n6308_8799.t68 vdd.t20 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X164 a_n6308_8799.t3 plus.t17 a_n3827_n3924.t26 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X165 a_n3827_n3924.t12 diffpairibias.t25 gnd.t66 gnd.t65 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X166 vdd.t22 a_n6308_8799.t69 CSoutput.t110 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X167 gnd.t265 gnd.t263 gnd.t264 gnd.t194 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X168 a_n6308_8799.t4 plus.t18 a_n3827_n3924.t25 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X169 vdd.t224 a_n6308_8799.t70 CSoutput.t109 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X170 minus.t3 gnd.t260 gnd.t262 gnd.t261 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X171 CSoutput.t48 commonsourceibias.t71 gnd.t133 gnd.t132 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X172 gnd.t259 gnd.t256 gnd.t258 gnd.t257 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X173 gnd.t255 gnd.t253 gnd.t254 gnd.t207 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X174 gnd.t186 commonsourceibias.t72 CSoutput.t47 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X175 diffpairibias.t11 diffpairibias.t10 gnd.t166 gnd.t165 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X176 a_n2848_n452.t35 minus.t15 a_n3827_n3924.t14 gnd.t78 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X177 vdd.t135 CSoutput.t154 output.t11 gnd.t71 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X178 CSoutput.t108 a_n6308_8799.t71 vdd.t225 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X179 a_n3827_n3924.t24 plus.t19 a_n6308_8799.t23 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X180 gnd.t151 commonsourceibias.t73 CSoutput.t46 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X181 CSoutput.t45 commonsourceibias.t74 gnd.t334 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X182 CSoutput.t107 a_n6308_8799.t72 vdd.t209 vdd.t208 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X183 vdd.t81 vdd.t79 vdd.t80 vdd.t62 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X184 a_n1808_13878.t17 a_n2848_n452.t60 vdd.t171 vdd.t170 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X185 vdd.t173 a_n2848_n452.t61 a_n1808_13878.t16 vdd.t172 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X186 gnd.t178 commonsourceibias.t75 CSoutput.t44 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X187 diffpairibias.t9 diffpairibias.t8 gnd.t168 gnd.t167 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X188 CSoutput.t155 a_n1986_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X189 gnd.t230 gnd.t228 gnd.t229 gnd.t194 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X190 a_n3827_n3924.t13 minus.t16 a_n2848_n452.t34 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X191 commonsourceibias.t21 commonsourceibias.t20 gnd.t176 gnd.t132 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X192 diffpairibias.t7 diffpairibias.t6 gnd.t139 gnd.t138 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X193 CSoutput.t106 a_n6308_8799.t73 vdd.t210 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X194 vdd.t27 a_n6308_8799.t74 CSoutput.t105 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X195 a_n3827_n3924.t44 minus.t17 a_n2848_n452.t41 gnd.t93 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X196 a_n3827_n3924.t23 plus.t20 a_n6308_8799.t27 gnd.t111 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X197 CSoutput.t156 a_n1986_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X198 output.t1 outputibias.t10 gnd.t109 gnd.t108 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X199 CSoutput.t43 commonsourceibias.t76 gnd.t181 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X200 a_n1986_8322.t10 a_n2848_n452.t62 a_n6308_8799.t2 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X201 a_n3827_n3924.t39 minus.t18 a_n2848_n452.t36 gnd.t85 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X202 gnd.t252 gnd.t250 gnd.t251 gnd.t236 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X203 commonsourceibias.t19 commonsourceibias.t18 gnd.t313 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X204 vdd.t29 a_n6308_8799.t75 CSoutput.t104 vdd.t28 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X205 CSoutput.t103 a_n6308_8799.t76 vdd.t5 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X206 gnd.t249 gnd.t246 gnd.t248 gnd.t247 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X207 vdd.t7 a_n6308_8799.t77 CSoutput.t102 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X208 vdd.t18 a_n2848_n452.t63 a_n1986_8322.t18 vdd.t17 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X209 CSoutput.t42 commonsourceibias.t77 gnd.t163 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X210 output.t0 outputibias.t11 gnd.t25 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X211 gnd.t124 commonsourceibias.t78 CSoutput.t41 gnd.t123 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X212 CSoutput.t40 commonsourceibias.t79 gnd.t171 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X213 output.t10 CSoutput.t157 vdd.t51 gnd.t57 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X214 gnd.t180 commonsourceibias.t16 commonsourceibias.t17 gnd.t26 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X215 gnd.t131 commonsourceibias.t80 CSoutput.t39 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X216 a_n1808_13878.t15 a_n2848_n452.t64 vdd.t131 vdd.t130 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X217 gnd.t245 gnd.t242 gnd.t244 gnd.t243 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X218 CSoutput.t38 commonsourceibias.t81 gnd.t61 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X219 gnd.t329 commonsourceibias.t82 CSoutput.t37 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X220 CSoutput.t36 commonsourceibias.t83 gnd.t157 gnd.t132 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X221 minus.t2 gnd.t239 gnd.t241 gnd.t240 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X222 commonsourceibias.t15 commonsourceibias.t14 gnd.t44 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X223 a_n3827_n3924.t6 diffpairibias.t26 gnd.t31 gnd.t30 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X224 vdd.t211 a_n6308_8799.t78 CSoutput.t101 vdd.t138 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X225 vdd.t78 vdd.t76 vdd.t77 vdd.t66 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X226 CSoutput.t100 a_n6308_8799.t79 vdd.t212 vdd.t208 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X227 CSoutput.t35 commonsourceibias.t84 gnd.t80 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X228 gnd.t152 commonsourceibias.t85 CSoutput.t34 gnd.t62 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X229 a_n6308_8799.t34 plus.t21 a_n3827_n3924.t22 gnd.t315 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X230 a_n2848_n452.t1 minus.t19 a_n3827_n3924.t2 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X231 CSoutput.t99 a_n6308_8799.t80 vdd.t186 vdd.t23 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X232 a_n3827_n3924.t5 minus.t20 a_n2848_n452.t4 gnd.t29 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X233 vdd.t75 vdd.t73 vdd.t74 vdd.t62 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X234 gnd.t53 commonsourceibias.t86 CSoutput.t33 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 CSoutput.t32 commonsourceibias.t87 gnd.t318 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X236 a_n1986_8322.t9 a_n2848_n452.t65 a_n6308_8799.t5 vdd.t132 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X237 vdd.t185 a_n2848_n452.t66 a_n1986_8322.t17 vdd.t184 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X238 vdd.t188 a_n6308_8799.t81 CSoutput.t98 vdd.t187 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X239 CSoutput.t97 a_n6308_8799.t82 vdd.t222 vdd.t208 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X240 CSoutput.t31 commonsourceibias.t88 gnd.t184 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X241 gnd.t173 commonsourceibias.t89 CSoutput.t30 gnd.t26 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X242 CSoutput.t96 a_n6308_8799.t83 vdd.t223 vdd.t152 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X243 a_n3827_n3924.t1 minus.t21 a_n2848_n452.t0 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X244 gnd.t238 gnd.t235 gnd.t237 gnd.t236 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X245 vdd.t167 a_n6308_8799.t84 CSoutput.t95 vdd.t154 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X246 vdd.t169 a_n6308_8799.t85 CSoutput.t94 vdd.t168 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X247 a_n3827_n3924.t43 minus.t22 a_n2848_n452.t40 gnd.t92 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X248 diffpairibias.t5 diffpairibias.t4 gnd.t68 gnd.t67 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X249 CSoutput.t29 commonsourceibias.t90 gnd.t190 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X250 gnd.t134 commonsourceibias.t91 CSoutput.t28 gnd.t123 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X251 vdd.t72 vdd.t69 vdd.t71 vdd.t70 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X252 CSoutput.t27 commonsourceibias.t92 gnd.t144 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X253 a_n1808_13878.t2 a_n2848_n452.t16 a_n2848_n452.t17 vdd.t174 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X254 gnd.t188 commonsourceibias.t93 CSoutput.t26 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X255 vdd.t52 CSoutput.t158 output.t9 gnd.t58 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X256 a_n3827_n3924.t57 diffpairibias.t27 gnd.t323 gnd.t322 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X257 a_n1986_8322.t8 a_n2848_n452.t67 a_n6308_8799.t16 vdd.t146 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X258 gnd.t161 commonsourceibias.t94 CSoutput.t25 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X259 CSoutput.t24 commonsourceibias.t95 gnd.t126 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X260 gnd.t234 gnd.t231 gnd.t233 gnd.t232 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X261 gnd.t127 commonsourceibias.t12 commonsourceibias.t13 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X262 outputibias.t3 outputibias.t2 gnd.t7 gnd.t6 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X263 gnd.t326 commonsourceibias.t96 CSoutput.t23 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X264 vdd.t217 a_n6308_8799.t86 CSoutput.t93 vdd.t154 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X265 CSoutput.t92 a_n6308_8799.t87 vdd.t218 vdd.t48 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X266 a_n3827_n3924.t42 minus.t23 a_n2848_n452.t39 gnd.t91 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X267 vdd.t192 a_n6308_8799.t88 CSoutput.t91 vdd.t138 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X268 CSoutput.t90 a_n6308_8799.t89 vdd.t193 vdd.t23 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X269 a_n1986_8322.t16 a_n2848_n452.t68 vdd.t197 vdd.t196 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X270 vdd.t68 vdd.t65 vdd.t67 vdd.t66 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X271 CSoutput.t22 commonsourceibias.t97 gnd.t76 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X272 gnd.t115 commonsourceibias.t98 CSoutput.t21 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X273 CSoutput.t20 commonsourceibias.t99 gnd.t141 gnd.t140 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X274 gnd.t162 commonsourceibias.t100 CSoutput.t19 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X275 gnd.t227 gnd.t225 plus.t2 gnd.t226 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X276 gnd.t15 commonsourceibias.t101 CSoutput.t18 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X277 gnd.t224 gnd.t221 gnd.t223 gnd.t222 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X278 commonsourceibias.t11 commonsourceibias.t10 gnd.t175 gnd.t121 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X279 gnd.t46 commonsourceibias.t8 commonsourceibias.t9 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X280 vdd.t199 a_n2848_n452.t69 a_n1808_13878.t14 vdd.t198 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X281 output.t8 CSoutput.t159 vdd.t53 gnd.t59 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X282 CSoutput.t89 a_n6308_8799.t90 vdd.t153 vdd.t152 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X283 vdd.t155 a_n6308_8799.t91 CSoutput.t88 vdd.t154 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X284 gnd.t177 commonsourceibias.t102 CSoutput.t17 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X285 CSoutput.t16 commonsourceibias.t103 gnd.t192 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X286 vdd.t182 a_n6308_8799.t92 CSoutput.t87 vdd.t168 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X287 vdd.t64 vdd.t61 vdd.t63 vdd.t62 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X288 a_n1986_8322.t7 a_n2848_n452.t70 a_n6308_8799.t21 vdd.t3 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X289 a_n3827_n3924.t21 plus.t22 a_n6308_8799.t15 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X290 gnd.t47 commonsourceibias.t6 commonsourceibias.t7 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X291 vdd.t60 vdd.t58 vdd.t59 vdd.t55 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X292 a_n6308_8799.t22 a_n2848_n452.t71 a_n1986_8322.t6 vdd.t174 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X293 a_n1808_13878.t13 a_n2848_n452.t72 vdd.t201 vdd.t200 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X294 vdd.t183 a_n6308_8799.t93 CSoutput.t86 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X295 CSoutput.t85 a_n6308_8799.t94 vdd.t215 vdd.t30 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X296 gnd.t220 gnd.t218 minus.t1 gnd.t219 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X297 CSoutput.t15 commonsourceibias.t104 gnd.t333 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X298 a_n2848_n452.t38 minus.t24 a_n3827_n3924.t41 gnd.t90 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X299 a_n6308_8799.t35 plus.t23 a_n3827_n3924.t20 gnd.t164 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X300 vdd.t156 CSoutput.t160 output.t7 gnd.t102 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X301 output.t6 CSoutput.t161 vdd.t157 gnd.t103 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X302 a_n2848_n452.t37 minus.t25 a_n3827_n3924.t40 gnd.t89 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X303 gnd.t128 commonsourceibias.t105 CSoutput.t14 gnd.t62 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X304 CSoutput.t13 commonsourceibias.t106 gnd.t182 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X305 gnd.t81 commonsourceibias.t4 commonsourceibias.t5 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X306 gnd.t82 commonsourceibias.t2 commonsourceibias.t3 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X307 CSoutput.t84 a_n6308_8799.t95 vdd.t216 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X308 a_n1808_13878.t1 a_n2848_n452.t20 a_n2848_n452.t21 vdd.t219 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X309 gnd.t130 commonsourceibias.t107 CSoutput.t12 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X310 CSoutput.t11 commonsourceibias.t108 gnd.t107 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X311 a_n3827_n3924.t56 minus.t26 a_n2848_n452.t47 gnd.t314 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X312 a_n3827_n3924.t46 diffpairibias.t28 gnd.t106 gnd.t105 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X313 a_n6308_8799.t0 plus.t24 a_n3827_n3924.t19 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X314 vdd.t158 CSoutput.t162 output.t5 gnd.t104 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X315 CSoutput.t83 a_n6308_8799.t96 vdd.t228 vdd.t147 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X316 gnd.t217 gnd.t214 gnd.t216 gnd.t215 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X317 vdd.t229 a_n6308_8799.t97 CSoutput.t82 vdd.t178 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X318 CSoutput.t10 commonsourceibias.t109 gnd.t64 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X319 gnd.t148 commonsourceibias.t110 CSoutput.t9 gnd.t45 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X320 diffpairibias.t3 diffpairibias.t2 gnd.t18 gnd.t17 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X321 gnd.t213 gnd.t210 gnd.t212 gnd.t211 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X322 a_n6308_8799.t20 a_n2848_n452.t73 a_n1986_8322.t5 vdd.t38 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X323 a_n2848_n452.t13 a_n2848_n452.t12 a_n1808_13878.t0 vdd.t3 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X324 gnd.t205 gnd.t203 plus.t1 gnd.t204 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X325 a_n2848_n452.t3 minus.t27 a_n3827_n3924.t4 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X326 vdd.t213 a_n6308_8799.t98 CSoutput.t81 vdd.t187 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X327 gnd.t155 commonsourceibias.t111 CSoutput.t8 gnd.t26 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X328 vdd.t50 CSoutput.t163 output.t4 gnd.t56 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X329 CSoutput.t164 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X330 gnd.t209 gnd.t206 gnd.t208 gnd.t207 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X331 vdd.t57 vdd.t54 vdd.t56 vdd.t55 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X332 vdd.t214 a_n6308_8799.t99 CSoutput.t80 vdd.t46 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X333 CSoutput.t7 commonsourceibias.t112 gnd.t55 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X334 diffpairibias.t1 diffpairibias.t0 gnd.t119 gnd.t118 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X335 CSoutput.t79 a_n6308_8799.t100 vdd.t230 vdd.t152 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X336 outputibias.t1 outputibias.t0 gnd.t49 gnd.t48 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X337 CSoutput.t165 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X338 plus.t0 gnd.t200 gnd.t202 gnd.t201 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X339 gnd.t22 commonsourceibias.t113 CSoutput.t6 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X340 gnd.t199 gnd.t197 minus.t0 gnd.t198 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X341 a_n6308_8799.t17 plus.t25 a_n3827_n3924.t18 gnd.t78 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X342 gnd.t196 gnd.t193 gnd.t195 gnd.t194 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X343 vdd.t14 a_n2848_n452.t74 a_n1808_13878.t12 vdd.t13 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X344 CSoutput.t78 a_n6308_8799.t101 vdd.t231 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X345 a_n6308_8799.t25 plus.t26 a_n3827_n3924.t17 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X346 a_n2848_n452.t43 minus.t28 a_n3827_n3924.t50 gnd.t145 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X347 CSoutput.t77 a_n6308_8799.t102 vdd.t180 vdd.t149 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X348 vdd.t181 a_n6308_8799.t103 CSoutput.t76 vdd.t168 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X349 CSoutput.t5 commonsourceibias.t114 gnd.t70 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X350 gnd.t185 commonsourceibias.t115 CSoutput.t4 gnd.t114 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X351 commonsourceibias.t1 commonsourceibias.t0 gnd.t87 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X352 CSoutput.t75 a_n6308_8799.t104 vdd.t177 vdd.t147 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X353 CSoutput.t3 commonsourceibias.t116 gnd.t189 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X354 vdd.t179 a_n6308_8799.t105 CSoutput.t74 vdd.t178 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X355 a_n1986_8322.t4 a_n2848_n452.t75 a_n6308_8799.t1 vdd.t15 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X356 a_n3827_n3924.t16 plus.t27 a_n6308_8799.t24 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X357 vdd.t175 a_n6308_8799.t106 CSoutput.t73 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X358 CSoutput.t72 a_n6308_8799.t107 vdd.t176 vdd.t42 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X359 CSoutput.t2 commonsourceibias.t117 gnd.t172 gnd.t75 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X360 gnd.t328 commonsourceibias.t118 CSoutput.t1 gnd.t62 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X361 CSoutput.t0 commonsourceibias.t119 gnd.t99 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X362 a_n3827_n3924.t15 plus.t28 a_n6308_8799.t18 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X363 a_n3827_n3924.t48 diffpairibias.t29 gnd.t113 gnd.t112 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
R0 gnd.n6527 gnd.n381 1056.13
R1 gnd.n5975 gnd.n5928 939.716
R2 gnd.n6881 gnd.n166 838.452
R3 gnd.n6992 gnd.n6891 838.452
R4 gnd.n2889 gnd.n2765 838.452
R5 gnd.n5194 gnd.n5193 838.452
R6 gnd.n2475 gnd.n2463 838.452
R7 gnd.n3926 gnd.n3925 838.452
R8 gnd.n3727 gnd.n2192 838.452
R9 gnd.n5806 gnd.n2265 838.452
R10 gnd.n7198 gnd.n162 783.196
R11 gnd.n7202 gnd.n7201 783.196
R12 gnd.n2888 gnd.n2887 783.196
R13 gnd.n5395 gnd.n2807 783.196
R14 gnd.n5675 gnd.n2468 783.196
R15 gnd.n3617 gnd.n3616 783.196
R16 gnd.n2268 gnd.n2267 783.196
R17 gnd.n5926 gnd.n2196 783.196
R18 gnd.n5990 gnd.n778 766.379
R19 gnd.n2153 gnd.n775 766.379
R20 gnd.n1465 gnd.n1368 766.379
R21 gnd.n1461 gnd.n1366 766.379
R22 gnd.n5974 gnd.n772 756.769
R23 gnd.n5985 gnd.n5984 756.769
R24 gnd.n1558 gnd.n1275 756.769
R25 gnd.n1556 gnd.n1278 756.769
R26 gnd.n3987 gnd.n3414 711.122
R27 gnd.n5050 gnd.n2903 711.122
R28 gnd.n3991 gnd.n3393 711.122
R29 gnd.n5410 gnd.n2730 711.122
R30 gnd.n6169 gnd.n594 689.5
R31 gnd.n6526 gnd.n382 689.5
R32 gnd.n6738 gnd.n6737 689.5
R33 gnd.n3634 gnd.n762 689.5
R34 gnd.n597 gnd.n594 585
R35 gnd.n6167 gnd.n594 585
R36 gnd.n6165 gnd.n6164 585
R37 gnd.n6166 gnd.n6165 585
R38 gnd.n6163 gnd.n596 585
R39 gnd.n596 gnd.n595 585
R40 gnd.n6162 gnd.n6161 585
R41 gnd.n6161 gnd.n6160 585
R42 gnd.n602 gnd.n601 585
R43 gnd.n6159 gnd.n602 585
R44 gnd.n6157 gnd.n6156 585
R45 gnd.n6158 gnd.n6157 585
R46 gnd.n6155 gnd.n604 585
R47 gnd.n604 gnd.n603 585
R48 gnd.n6154 gnd.n6153 585
R49 gnd.n6153 gnd.n6152 585
R50 gnd.n610 gnd.n609 585
R51 gnd.n6151 gnd.n610 585
R52 gnd.n6149 gnd.n6148 585
R53 gnd.n6150 gnd.n6149 585
R54 gnd.n6147 gnd.n612 585
R55 gnd.n612 gnd.n611 585
R56 gnd.n6146 gnd.n6145 585
R57 gnd.n6145 gnd.n6144 585
R58 gnd.n618 gnd.n617 585
R59 gnd.n6143 gnd.n618 585
R60 gnd.n6141 gnd.n6140 585
R61 gnd.n6142 gnd.n6141 585
R62 gnd.n6139 gnd.n620 585
R63 gnd.n620 gnd.n619 585
R64 gnd.n6138 gnd.n6137 585
R65 gnd.n6137 gnd.n6136 585
R66 gnd.n626 gnd.n625 585
R67 gnd.n6135 gnd.n626 585
R68 gnd.n6133 gnd.n6132 585
R69 gnd.n6134 gnd.n6133 585
R70 gnd.n6131 gnd.n628 585
R71 gnd.n628 gnd.n627 585
R72 gnd.n6130 gnd.n6129 585
R73 gnd.n6129 gnd.n6128 585
R74 gnd.n634 gnd.n633 585
R75 gnd.n6127 gnd.n634 585
R76 gnd.n6125 gnd.n6124 585
R77 gnd.n6126 gnd.n6125 585
R78 gnd.n6123 gnd.n636 585
R79 gnd.n636 gnd.n635 585
R80 gnd.n6122 gnd.n6121 585
R81 gnd.n6121 gnd.n6120 585
R82 gnd.n642 gnd.n641 585
R83 gnd.n6119 gnd.n642 585
R84 gnd.n6117 gnd.n6116 585
R85 gnd.n6118 gnd.n6117 585
R86 gnd.n6115 gnd.n644 585
R87 gnd.n644 gnd.n643 585
R88 gnd.n6114 gnd.n6113 585
R89 gnd.n6113 gnd.n6112 585
R90 gnd.n650 gnd.n649 585
R91 gnd.n6111 gnd.n650 585
R92 gnd.n6109 gnd.n6108 585
R93 gnd.n6110 gnd.n6109 585
R94 gnd.n6107 gnd.n652 585
R95 gnd.n652 gnd.n651 585
R96 gnd.n6106 gnd.n6105 585
R97 gnd.n6105 gnd.n6104 585
R98 gnd.n658 gnd.n657 585
R99 gnd.n6103 gnd.n658 585
R100 gnd.n6101 gnd.n6100 585
R101 gnd.n6102 gnd.n6101 585
R102 gnd.n6099 gnd.n660 585
R103 gnd.n660 gnd.n659 585
R104 gnd.n6098 gnd.n6097 585
R105 gnd.n6097 gnd.n6096 585
R106 gnd.n666 gnd.n665 585
R107 gnd.n6095 gnd.n666 585
R108 gnd.n6093 gnd.n6092 585
R109 gnd.n6094 gnd.n6093 585
R110 gnd.n6091 gnd.n668 585
R111 gnd.n668 gnd.n667 585
R112 gnd.n6090 gnd.n6089 585
R113 gnd.n6089 gnd.n6088 585
R114 gnd.n674 gnd.n673 585
R115 gnd.n6087 gnd.n674 585
R116 gnd.n6085 gnd.n6084 585
R117 gnd.n6086 gnd.n6085 585
R118 gnd.n6083 gnd.n676 585
R119 gnd.n676 gnd.n675 585
R120 gnd.n6082 gnd.n6081 585
R121 gnd.n6081 gnd.n6080 585
R122 gnd.n682 gnd.n681 585
R123 gnd.n6079 gnd.n682 585
R124 gnd.n6077 gnd.n6076 585
R125 gnd.n6078 gnd.n6077 585
R126 gnd.n6075 gnd.n684 585
R127 gnd.n684 gnd.n683 585
R128 gnd.n6074 gnd.n6073 585
R129 gnd.n6073 gnd.n6072 585
R130 gnd.n690 gnd.n689 585
R131 gnd.n6071 gnd.n690 585
R132 gnd.n6069 gnd.n6068 585
R133 gnd.n6070 gnd.n6069 585
R134 gnd.n6067 gnd.n692 585
R135 gnd.n692 gnd.n691 585
R136 gnd.n6066 gnd.n6065 585
R137 gnd.n6065 gnd.n6064 585
R138 gnd.n698 gnd.n697 585
R139 gnd.n6063 gnd.n698 585
R140 gnd.n6061 gnd.n6060 585
R141 gnd.n6062 gnd.n6061 585
R142 gnd.n6059 gnd.n700 585
R143 gnd.n700 gnd.n699 585
R144 gnd.n6058 gnd.n6057 585
R145 gnd.n6057 gnd.n6056 585
R146 gnd.n706 gnd.n705 585
R147 gnd.n6055 gnd.n706 585
R148 gnd.n6053 gnd.n6052 585
R149 gnd.n6054 gnd.n6053 585
R150 gnd.n6051 gnd.n708 585
R151 gnd.n708 gnd.n707 585
R152 gnd.n6050 gnd.n6049 585
R153 gnd.n6049 gnd.n6048 585
R154 gnd.n714 gnd.n713 585
R155 gnd.n6047 gnd.n714 585
R156 gnd.n6045 gnd.n6044 585
R157 gnd.n6046 gnd.n6045 585
R158 gnd.n6043 gnd.n716 585
R159 gnd.n716 gnd.n715 585
R160 gnd.n6042 gnd.n6041 585
R161 gnd.n6041 gnd.n6040 585
R162 gnd.n722 gnd.n721 585
R163 gnd.n6039 gnd.n722 585
R164 gnd.n6037 gnd.n6036 585
R165 gnd.n6038 gnd.n6037 585
R166 gnd.n6035 gnd.n724 585
R167 gnd.n724 gnd.n723 585
R168 gnd.n6034 gnd.n6033 585
R169 gnd.n6033 gnd.n6032 585
R170 gnd.n730 gnd.n729 585
R171 gnd.n6031 gnd.n730 585
R172 gnd.n6029 gnd.n6028 585
R173 gnd.n6030 gnd.n6029 585
R174 gnd.n6027 gnd.n732 585
R175 gnd.n732 gnd.n731 585
R176 gnd.n6026 gnd.n6025 585
R177 gnd.n6025 gnd.n6024 585
R178 gnd.n738 gnd.n737 585
R179 gnd.n6023 gnd.n738 585
R180 gnd.n6021 gnd.n6020 585
R181 gnd.n6022 gnd.n6021 585
R182 gnd.n6019 gnd.n740 585
R183 gnd.n740 gnd.n739 585
R184 gnd.n6018 gnd.n6017 585
R185 gnd.n6017 gnd.n6016 585
R186 gnd.n746 gnd.n745 585
R187 gnd.n6015 gnd.n746 585
R188 gnd.n6013 gnd.n6012 585
R189 gnd.n6014 gnd.n6013 585
R190 gnd.n6011 gnd.n748 585
R191 gnd.n748 gnd.n747 585
R192 gnd.n6010 gnd.n6009 585
R193 gnd.n6009 gnd.n6008 585
R194 gnd.n754 gnd.n753 585
R195 gnd.n6007 gnd.n754 585
R196 gnd.n6005 gnd.n6004 585
R197 gnd.n6006 gnd.n6005 585
R198 gnd.n6003 gnd.n756 585
R199 gnd.n756 gnd.n755 585
R200 gnd.n6002 gnd.n6001 585
R201 gnd.n6001 gnd.n6000 585
R202 gnd.n6170 gnd.n6169 585
R203 gnd.n6169 gnd.n6168 585
R204 gnd.n592 gnd.n591 585
R205 gnd.n591 gnd.n590 585
R206 gnd.n6175 gnd.n6174 585
R207 gnd.n6176 gnd.n6175 585
R208 gnd.n589 gnd.n588 585
R209 gnd.n6177 gnd.n589 585
R210 gnd.n6180 gnd.n6179 585
R211 gnd.n6179 gnd.n6178 585
R212 gnd.n586 gnd.n585 585
R213 gnd.n585 gnd.n584 585
R214 gnd.n6185 gnd.n6184 585
R215 gnd.n6186 gnd.n6185 585
R216 gnd.n583 gnd.n582 585
R217 gnd.n6187 gnd.n583 585
R218 gnd.n6190 gnd.n6189 585
R219 gnd.n6189 gnd.n6188 585
R220 gnd.n580 gnd.n579 585
R221 gnd.n579 gnd.n578 585
R222 gnd.n6195 gnd.n6194 585
R223 gnd.n6196 gnd.n6195 585
R224 gnd.n577 gnd.n576 585
R225 gnd.n6197 gnd.n577 585
R226 gnd.n6200 gnd.n6199 585
R227 gnd.n6199 gnd.n6198 585
R228 gnd.n574 gnd.n573 585
R229 gnd.n573 gnd.n572 585
R230 gnd.n6205 gnd.n6204 585
R231 gnd.n6206 gnd.n6205 585
R232 gnd.n571 gnd.n570 585
R233 gnd.n6207 gnd.n571 585
R234 gnd.n6210 gnd.n6209 585
R235 gnd.n6209 gnd.n6208 585
R236 gnd.n568 gnd.n567 585
R237 gnd.n567 gnd.n566 585
R238 gnd.n6215 gnd.n6214 585
R239 gnd.n6216 gnd.n6215 585
R240 gnd.n565 gnd.n564 585
R241 gnd.n6217 gnd.n565 585
R242 gnd.n6220 gnd.n6219 585
R243 gnd.n6219 gnd.n6218 585
R244 gnd.n562 gnd.n561 585
R245 gnd.n561 gnd.n560 585
R246 gnd.n6225 gnd.n6224 585
R247 gnd.n6226 gnd.n6225 585
R248 gnd.n559 gnd.n558 585
R249 gnd.n6227 gnd.n559 585
R250 gnd.n6230 gnd.n6229 585
R251 gnd.n6229 gnd.n6228 585
R252 gnd.n556 gnd.n555 585
R253 gnd.n555 gnd.n554 585
R254 gnd.n6235 gnd.n6234 585
R255 gnd.n6236 gnd.n6235 585
R256 gnd.n553 gnd.n552 585
R257 gnd.n6237 gnd.n553 585
R258 gnd.n6240 gnd.n6239 585
R259 gnd.n6239 gnd.n6238 585
R260 gnd.n550 gnd.n549 585
R261 gnd.n549 gnd.n548 585
R262 gnd.n6245 gnd.n6244 585
R263 gnd.n6246 gnd.n6245 585
R264 gnd.n547 gnd.n546 585
R265 gnd.n6247 gnd.n547 585
R266 gnd.n6250 gnd.n6249 585
R267 gnd.n6249 gnd.n6248 585
R268 gnd.n544 gnd.n543 585
R269 gnd.n543 gnd.n542 585
R270 gnd.n6255 gnd.n6254 585
R271 gnd.n6256 gnd.n6255 585
R272 gnd.n541 gnd.n540 585
R273 gnd.n6257 gnd.n541 585
R274 gnd.n6260 gnd.n6259 585
R275 gnd.n6259 gnd.n6258 585
R276 gnd.n538 gnd.n537 585
R277 gnd.n537 gnd.n536 585
R278 gnd.n6265 gnd.n6264 585
R279 gnd.n6266 gnd.n6265 585
R280 gnd.n535 gnd.n534 585
R281 gnd.n6267 gnd.n535 585
R282 gnd.n6270 gnd.n6269 585
R283 gnd.n6269 gnd.n6268 585
R284 gnd.n532 gnd.n531 585
R285 gnd.n531 gnd.n530 585
R286 gnd.n6275 gnd.n6274 585
R287 gnd.n6276 gnd.n6275 585
R288 gnd.n529 gnd.n528 585
R289 gnd.n6277 gnd.n529 585
R290 gnd.n6280 gnd.n6279 585
R291 gnd.n6279 gnd.n6278 585
R292 gnd.n526 gnd.n525 585
R293 gnd.n525 gnd.n524 585
R294 gnd.n6285 gnd.n6284 585
R295 gnd.n6286 gnd.n6285 585
R296 gnd.n523 gnd.n522 585
R297 gnd.n6287 gnd.n523 585
R298 gnd.n6290 gnd.n6289 585
R299 gnd.n6289 gnd.n6288 585
R300 gnd.n520 gnd.n519 585
R301 gnd.n519 gnd.n518 585
R302 gnd.n6295 gnd.n6294 585
R303 gnd.n6296 gnd.n6295 585
R304 gnd.n517 gnd.n516 585
R305 gnd.n6297 gnd.n517 585
R306 gnd.n6300 gnd.n6299 585
R307 gnd.n6299 gnd.n6298 585
R308 gnd.n514 gnd.n513 585
R309 gnd.n513 gnd.n512 585
R310 gnd.n6305 gnd.n6304 585
R311 gnd.n6306 gnd.n6305 585
R312 gnd.n511 gnd.n510 585
R313 gnd.n6307 gnd.n511 585
R314 gnd.n6310 gnd.n6309 585
R315 gnd.n6309 gnd.n6308 585
R316 gnd.n508 gnd.n507 585
R317 gnd.n507 gnd.n506 585
R318 gnd.n6315 gnd.n6314 585
R319 gnd.n6316 gnd.n6315 585
R320 gnd.n505 gnd.n504 585
R321 gnd.n6317 gnd.n505 585
R322 gnd.n6320 gnd.n6319 585
R323 gnd.n6319 gnd.n6318 585
R324 gnd.n502 gnd.n501 585
R325 gnd.n501 gnd.n500 585
R326 gnd.n6325 gnd.n6324 585
R327 gnd.n6326 gnd.n6325 585
R328 gnd.n499 gnd.n498 585
R329 gnd.n6327 gnd.n499 585
R330 gnd.n6330 gnd.n6329 585
R331 gnd.n6329 gnd.n6328 585
R332 gnd.n496 gnd.n495 585
R333 gnd.n495 gnd.n494 585
R334 gnd.n6335 gnd.n6334 585
R335 gnd.n6336 gnd.n6335 585
R336 gnd.n493 gnd.n492 585
R337 gnd.n6337 gnd.n493 585
R338 gnd.n6340 gnd.n6339 585
R339 gnd.n6339 gnd.n6338 585
R340 gnd.n490 gnd.n489 585
R341 gnd.n489 gnd.n488 585
R342 gnd.n6345 gnd.n6344 585
R343 gnd.n6346 gnd.n6345 585
R344 gnd.n487 gnd.n486 585
R345 gnd.n6347 gnd.n487 585
R346 gnd.n6350 gnd.n6349 585
R347 gnd.n6349 gnd.n6348 585
R348 gnd.n484 gnd.n483 585
R349 gnd.n483 gnd.n482 585
R350 gnd.n6355 gnd.n6354 585
R351 gnd.n6356 gnd.n6355 585
R352 gnd.n481 gnd.n480 585
R353 gnd.n6357 gnd.n481 585
R354 gnd.n6360 gnd.n6359 585
R355 gnd.n6359 gnd.n6358 585
R356 gnd.n478 gnd.n477 585
R357 gnd.n477 gnd.n476 585
R358 gnd.n6365 gnd.n6364 585
R359 gnd.n6366 gnd.n6365 585
R360 gnd.n475 gnd.n474 585
R361 gnd.n6367 gnd.n475 585
R362 gnd.n6370 gnd.n6369 585
R363 gnd.n6369 gnd.n6368 585
R364 gnd.n472 gnd.n471 585
R365 gnd.n471 gnd.n470 585
R366 gnd.n6375 gnd.n6374 585
R367 gnd.n6376 gnd.n6375 585
R368 gnd.n469 gnd.n468 585
R369 gnd.n6377 gnd.n469 585
R370 gnd.n6380 gnd.n6379 585
R371 gnd.n6379 gnd.n6378 585
R372 gnd.n466 gnd.n465 585
R373 gnd.n465 gnd.n464 585
R374 gnd.n6385 gnd.n6384 585
R375 gnd.n6386 gnd.n6385 585
R376 gnd.n463 gnd.n462 585
R377 gnd.n6387 gnd.n463 585
R378 gnd.n6390 gnd.n6389 585
R379 gnd.n6389 gnd.n6388 585
R380 gnd.n460 gnd.n459 585
R381 gnd.n459 gnd.n458 585
R382 gnd.n6395 gnd.n6394 585
R383 gnd.n6396 gnd.n6395 585
R384 gnd.n457 gnd.n456 585
R385 gnd.n6397 gnd.n457 585
R386 gnd.n6400 gnd.n6399 585
R387 gnd.n6399 gnd.n6398 585
R388 gnd.n454 gnd.n453 585
R389 gnd.n453 gnd.n452 585
R390 gnd.n6405 gnd.n6404 585
R391 gnd.n6406 gnd.n6405 585
R392 gnd.n451 gnd.n450 585
R393 gnd.n6407 gnd.n451 585
R394 gnd.n6410 gnd.n6409 585
R395 gnd.n6409 gnd.n6408 585
R396 gnd.n448 gnd.n447 585
R397 gnd.n447 gnd.n446 585
R398 gnd.n6415 gnd.n6414 585
R399 gnd.n6416 gnd.n6415 585
R400 gnd.n445 gnd.n444 585
R401 gnd.n6417 gnd.n445 585
R402 gnd.n6420 gnd.n6419 585
R403 gnd.n6419 gnd.n6418 585
R404 gnd.n442 gnd.n441 585
R405 gnd.n441 gnd.n440 585
R406 gnd.n6425 gnd.n6424 585
R407 gnd.n6426 gnd.n6425 585
R408 gnd.n439 gnd.n438 585
R409 gnd.n6427 gnd.n439 585
R410 gnd.n6430 gnd.n6429 585
R411 gnd.n6429 gnd.n6428 585
R412 gnd.n436 gnd.n435 585
R413 gnd.n435 gnd.n434 585
R414 gnd.n6435 gnd.n6434 585
R415 gnd.n6436 gnd.n6435 585
R416 gnd.n433 gnd.n432 585
R417 gnd.n6437 gnd.n433 585
R418 gnd.n6440 gnd.n6439 585
R419 gnd.n6439 gnd.n6438 585
R420 gnd.n430 gnd.n429 585
R421 gnd.n429 gnd.n428 585
R422 gnd.n6445 gnd.n6444 585
R423 gnd.n6446 gnd.n6445 585
R424 gnd.n427 gnd.n426 585
R425 gnd.n6447 gnd.n427 585
R426 gnd.n6450 gnd.n6449 585
R427 gnd.n6449 gnd.n6448 585
R428 gnd.n424 gnd.n423 585
R429 gnd.n423 gnd.n422 585
R430 gnd.n6455 gnd.n6454 585
R431 gnd.n6456 gnd.n6455 585
R432 gnd.n421 gnd.n420 585
R433 gnd.n6457 gnd.n421 585
R434 gnd.n6460 gnd.n6459 585
R435 gnd.n6459 gnd.n6458 585
R436 gnd.n418 gnd.n417 585
R437 gnd.n417 gnd.n416 585
R438 gnd.n6465 gnd.n6464 585
R439 gnd.n6466 gnd.n6465 585
R440 gnd.n415 gnd.n414 585
R441 gnd.n6467 gnd.n415 585
R442 gnd.n6470 gnd.n6469 585
R443 gnd.n6469 gnd.n6468 585
R444 gnd.n412 gnd.n411 585
R445 gnd.n411 gnd.n410 585
R446 gnd.n6475 gnd.n6474 585
R447 gnd.n6476 gnd.n6475 585
R448 gnd.n409 gnd.n408 585
R449 gnd.n6477 gnd.n409 585
R450 gnd.n6480 gnd.n6479 585
R451 gnd.n6479 gnd.n6478 585
R452 gnd.n406 gnd.n405 585
R453 gnd.n405 gnd.n404 585
R454 gnd.n6485 gnd.n6484 585
R455 gnd.n6486 gnd.n6485 585
R456 gnd.n403 gnd.n402 585
R457 gnd.n6487 gnd.n403 585
R458 gnd.n6490 gnd.n6489 585
R459 gnd.n6489 gnd.n6488 585
R460 gnd.n400 gnd.n399 585
R461 gnd.n399 gnd.n398 585
R462 gnd.n6495 gnd.n6494 585
R463 gnd.n6496 gnd.n6495 585
R464 gnd.n397 gnd.n396 585
R465 gnd.n6497 gnd.n397 585
R466 gnd.n6500 gnd.n6499 585
R467 gnd.n6499 gnd.n6498 585
R468 gnd.n394 gnd.n393 585
R469 gnd.n393 gnd.n392 585
R470 gnd.n6505 gnd.n6504 585
R471 gnd.n6506 gnd.n6505 585
R472 gnd.n391 gnd.n390 585
R473 gnd.n6507 gnd.n391 585
R474 gnd.n6510 gnd.n6509 585
R475 gnd.n6509 gnd.n6508 585
R476 gnd.n388 gnd.n387 585
R477 gnd.n387 gnd.n386 585
R478 gnd.n6516 gnd.n6515 585
R479 gnd.n6517 gnd.n6516 585
R480 gnd.n385 gnd.n384 585
R481 gnd.n6518 gnd.n385 585
R482 gnd.n6521 gnd.n6520 585
R483 gnd.n6520 gnd.n6519 585
R484 gnd.n6522 gnd.n382 585
R485 gnd.n382 gnd.n381 585
R486 gnd.n257 gnd.n256 585
R487 gnd.n6729 gnd.n256 585
R488 gnd.n6732 gnd.n6731 585
R489 gnd.n6731 gnd.n6730 585
R490 gnd.n260 gnd.n259 585
R491 gnd.n6728 gnd.n260 585
R492 gnd.n6726 gnd.n6725 585
R493 gnd.n6727 gnd.n6726 585
R494 gnd.n263 gnd.n262 585
R495 gnd.n262 gnd.n261 585
R496 gnd.n6721 gnd.n6720 585
R497 gnd.n6720 gnd.n6719 585
R498 gnd.n266 gnd.n265 585
R499 gnd.n6718 gnd.n266 585
R500 gnd.n6716 gnd.n6715 585
R501 gnd.n6717 gnd.n6716 585
R502 gnd.n269 gnd.n268 585
R503 gnd.n268 gnd.n267 585
R504 gnd.n6711 gnd.n6710 585
R505 gnd.n6710 gnd.n6709 585
R506 gnd.n272 gnd.n271 585
R507 gnd.n6708 gnd.n272 585
R508 gnd.n6706 gnd.n6705 585
R509 gnd.n6707 gnd.n6706 585
R510 gnd.n275 gnd.n274 585
R511 gnd.n274 gnd.n273 585
R512 gnd.n6701 gnd.n6700 585
R513 gnd.n6700 gnd.n6699 585
R514 gnd.n278 gnd.n277 585
R515 gnd.n6698 gnd.n278 585
R516 gnd.n6696 gnd.n6695 585
R517 gnd.n6697 gnd.n6696 585
R518 gnd.n281 gnd.n280 585
R519 gnd.n280 gnd.n279 585
R520 gnd.n6691 gnd.n6690 585
R521 gnd.n6690 gnd.n6689 585
R522 gnd.n284 gnd.n283 585
R523 gnd.n6688 gnd.n284 585
R524 gnd.n6686 gnd.n6685 585
R525 gnd.n6687 gnd.n6686 585
R526 gnd.n287 gnd.n286 585
R527 gnd.n286 gnd.n285 585
R528 gnd.n6681 gnd.n6680 585
R529 gnd.n6680 gnd.n6679 585
R530 gnd.n290 gnd.n289 585
R531 gnd.n6678 gnd.n290 585
R532 gnd.n6676 gnd.n6675 585
R533 gnd.n6677 gnd.n6676 585
R534 gnd.n293 gnd.n292 585
R535 gnd.n292 gnd.n291 585
R536 gnd.n6671 gnd.n6670 585
R537 gnd.n6670 gnd.n6669 585
R538 gnd.n296 gnd.n295 585
R539 gnd.n6668 gnd.n296 585
R540 gnd.n6666 gnd.n6665 585
R541 gnd.n6667 gnd.n6666 585
R542 gnd.n299 gnd.n298 585
R543 gnd.n298 gnd.n297 585
R544 gnd.n6661 gnd.n6660 585
R545 gnd.n6660 gnd.n6659 585
R546 gnd.n302 gnd.n301 585
R547 gnd.n6658 gnd.n302 585
R548 gnd.n6656 gnd.n6655 585
R549 gnd.n6657 gnd.n6656 585
R550 gnd.n305 gnd.n304 585
R551 gnd.n304 gnd.n303 585
R552 gnd.n6651 gnd.n6650 585
R553 gnd.n6650 gnd.n6649 585
R554 gnd.n308 gnd.n307 585
R555 gnd.n6648 gnd.n308 585
R556 gnd.n6646 gnd.n6645 585
R557 gnd.n6647 gnd.n6646 585
R558 gnd.n311 gnd.n310 585
R559 gnd.n310 gnd.n309 585
R560 gnd.n6641 gnd.n6640 585
R561 gnd.n6640 gnd.n6639 585
R562 gnd.n314 gnd.n313 585
R563 gnd.n6638 gnd.n314 585
R564 gnd.n6636 gnd.n6635 585
R565 gnd.n6637 gnd.n6636 585
R566 gnd.n317 gnd.n316 585
R567 gnd.n316 gnd.n315 585
R568 gnd.n6631 gnd.n6630 585
R569 gnd.n6630 gnd.n6629 585
R570 gnd.n320 gnd.n319 585
R571 gnd.n6628 gnd.n320 585
R572 gnd.n6626 gnd.n6625 585
R573 gnd.n6627 gnd.n6626 585
R574 gnd.n323 gnd.n322 585
R575 gnd.n322 gnd.n321 585
R576 gnd.n6621 gnd.n6620 585
R577 gnd.n6620 gnd.n6619 585
R578 gnd.n326 gnd.n325 585
R579 gnd.n6618 gnd.n326 585
R580 gnd.n6616 gnd.n6615 585
R581 gnd.n6617 gnd.n6616 585
R582 gnd.n329 gnd.n328 585
R583 gnd.n328 gnd.n327 585
R584 gnd.n6611 gnd.n6610 585
R585 gnd.n6610 gnd.n6609 585
R586 gnd.n332 gnd.n331 585
R587 gnd.n6608 gnd.n332 585
R588 gnd.n6606 gnd.n6605 585
R589 gnd.n6607 gnd.n6606 585
R590 gnd.n335 gnd.n334 585
R591 gnd.n334 gnd.n333 585
R592 gnd.n6601 gnd.n6600 585
R593 gnd.n6600 gnd.n6599 585
R594 gnd.n338 gnd.n337 585
R595 gnd.n6598 gnd.n338 585
R596 gnd.n6596 gnd.n6595 585
R597 gnd.n6597 gnd.n6596 585
R598 gnd.n341 gnd.n340 585
R599 gnd.n340 gnd.n339 585
R600 gnd.n6591 gnd.n6590 585
R601 gnd.n6590 gnd.n6589 585
R602 gnd.n344 gnd.n343 585
R603 gnd.n6588 gnd.n344 585
R604 gnd.n6586 gnd.n6585 585
R605 gnd.n6587 gnd.n6586 585
R606 gnd.n347 gnd.n346 585
R607 gnd.n346 gnd.n345 585
R608 gnd.n6581 gnd.n6580 585
R609 gnd.n6580 gnd.n6579 585
R610 gnd.n350 gnd.n349 585
R611 gnd.n6578 gnd.n350 585
R612 gnd.n6576 gnd.n6575 585
R613 gnd.n6577 gnd.n6576 585
R614 gnd.n353 gnd.n352 585
R615 gnd.n352 gnd.n351 585
R616 gnd.n6571 gnd.n6570 585
R617 gnd.n6570 gnd.n6569 585
R618 gnd.n356 gnd.n355 585
R619 gnd.n6568 gnd.n356 585
R620 gnd.n6566 gnd.n6565 585
R621 gnd.n6567 gnd.n6566 585
R622 gnd.n359 gnd.n358 585
R623 gnd.n358 gnd.n357 585
R624 gnd.n6561 gnd.n6560 585
R625 gnd.n6560 gnd.n6559 585
R626 gnd.n362 gnd.n361 585
R627 gnd.n6558 gnd.n362 585
R628 gnd.n6556 gnd.n6555 585
R629 gnd.n6557 gnd.n6556 585
R630 gnd.n365 gnd.n364 585
R631 gnd.n364 gnd.n363 585
R632 gnd.n6551 gnd.n6550 585
R633 gnd.n6550 gnd.n6549 585
R634 gnd.n368 gnd.n367 585
R635 gnd.n6548 gnd.n368 585
R636 gnd.n6546 gnd.n6545 585
R637 gnd.n6547 gnd.n6546 585
R638 gnd.n371 gnd.n370 585
R639 gnd.n370 gnd.n369 585
R640 gnd.n6541 gnd.n6540 585
R641 gnd.n6540 gnd.n6539 585
R642 gnd.n374 gnd.n373 585
R643 gnd.n6538 gnd.n374 585
R644 gnd.n6536 gnd.n6535 585
R645 gnd.n6537 gnd.n6536 585
R646 gnd.n377 gnd.n376 585
R647 gnd.n376 gnd.n375 585
R648 gnd.n6531 gnd.n6530 585
R649 gnd.n6530 gnd.n6529 585
R650 gnd.n380 gnd.n379 585
R651 gnd.n6528 gnd.n380 585
R652 gnd.n6526 gnd.n6525 585
R653 gnd.n6527 gnd.n6526 585
R654 gnd.n2463 gnd.n2462 585
R655 gnd.n3924 gnd.n2463 585
R656 gnd.n5684 gnd.n5683 585
R657 gnd.n5683 gnd.n5682 585
R658 gnd.n5685 gnd.n2458 585
R659 gnd.n3863 gnd.n2458 585
R660 gnd.n5687 gnd.n5686 585
R661 gnd.n5688 gnd.n5687 585
R662 gnd.n2442 gnd.n2441 585
R663 gnd.n3854 gnd.n2442 585
R664 gnd.n5696 gnd.n5695 585
R665 gnd.n5695 gnd.n5694 585
R666 gnd.n5697 gnd.n2437 585
R667 gnd.n3849 gnd.n2437 585
R668 gnd.n5699 gnd.n5698 585
R669 gnd.n5700 gnd.n5699 585
R670 gnd.n2422 gnd.n2421 585
R671 gnd.n3845 gnd.n2422 585
R672 gnd.n5708 gnd.n5707 585
R673 gnd.n5707 gnd.n5706 585
R674 gnd.n5709 gnd.n2417 585
R675 gnd.n3883 gnd.n2417 585
R676 gnd.n5711 gnd.n5710 585
R677 gnd.n5712 gnd.n5711 585
R678 gnd.n2401 gnd.n2400 585
R679 gnd.n3838 gnd.n2401 585
R680 gnd.n5720 gnd.n5719 585
R681 gnd.n5719 gnd.n5718 585
R682 gnd.n5721 gnd.n2396 585
R683 gnd.n3830 gnd.n2396 585
R684 gnd.n5723 gnd.n5722 585
R685 gnd.n5724 gnd.n5723 585
R686 gnd.n2382 gnd.n2381 585
R687 gnd.n2385 gnd.n2382 585
R688 gnd.n5732 gnd.n5731 585
R689 gnd.n5731 gnd.n5730 585
R690 gnd.n5733 gnd.n2377 585
R691 gnd.n2377 gnd.n2376 585
R692 gnd.n5735 gnd.n5734 585
R693 gnd.n5736 gnd.n5735 585
R694 gnd.n2362 gnd.n2361 585
R695 gnd.n2366 gnd.n2362 585
R696 gnd.n5744 gnd.n5743 585
R697 gnd.n5743 gnd.n5742 585
R698 gnd.n5745 gnd.n2357 585
R699 gnd.n2363 gnd.n2357 585
R700 gnd.n5747 gnd.n5746 585
R701 gnd.n5748 gnd.n5747 585
R702 gnd.n2344 gnd.n2343 585
R703 gnd.n2354 gnd.n2344 585
R704 gnd.n5756 gnd.n5755 585
R705 gnd.n5755 gnd.n5754 585
R706 gnd.n5757 gnd.n2339 585
R707 gnd.n2339 gnd.n2338 585
R708 gnd.n5759 gnd.n5758 585
R709 gnd.n5760 gnd.n5759 585
R710 gnd.n2324 gnd.n2323 585
R711 gnd.n2328 gnd.n2324 585
R712 gnd.n5768 gnd.n5767 585
R713 gnd.n5767 gnd.n5766 585
R714 gnd.n5769 gnd.n2319 585
R715 gnd.n2325 gnd.n2319 585
R716 gnd.n5771 gnd.n5770 585
R717 gnd.n5772 gnd.n5771 585
R718 gnd.n2306 gnd.n2305 585
R719 gnd.n2316 gnd.n2306 585
R720 gnd.n5780 gnd.n5779 585
R721 gnd.n5779 gnd.n5778 585
R722 gnd.n5781 gnd.n2301 585
R723 gnd.n2301 gnd.n2300 585
R724 gnd.n5783 gnd.n5782 585
R725 gnd.n5784 gnd.n5783 585
R726 gnd.n2288 gnd.n2287 585
R727 gnd.n2291 gnd.n2288 585
R728 gnd.n5792 gnd.n5791 585
R729 gnd.n5791 gnd.n5790 585
R730 gnd.n5793 gnd.n2282 585
R731 gnd.n2282 gnd.n2281 585
R732 gnd.n5795 gnd.n5794 585
R733 gnd.n5796 gnd.n5795 585
R734 gnd.n2283 gnd.n2266 585
R735 gnd.n2278 gnd.n2266 585
R736 gnd.n5805 gnd.n2264 585
R737 gnd.n5805 gnd.n5804 585
R738 gnd.n5807 gnd.n5806 585
R739 gnd.n5806 gnd.n2193 585
R740 gnd.n3685 gnd.n2265 585
R741 gnd.n3687 gnd.n3686 585
R742 gnd.n3689 gnd.n3688 585
R743 gnd.n3693 gnd.n3683 585
R744 gnd.n3695 gnd.n3694 585
R745 gnd.n3697 gnd.n3696 585
R746 gnd.n3699 gnd.n3698 585
R747 gnd.n3703 gnd.n3681 585
R748 gnd.n3705 gnd.n3704 585
R749 gnd.n3707 gnd.n3706 585
R750 gnd.n3709 gnd.n3708 585
R751 gnd.n3713 gnd.n3679 585
R752 gnd.n3715 gnd.n3714 585
R753 gnd.n3717 gnd.n3716 585
R754 gnd.n3719 gnd.n3718 585
R755 gnd.n3676 gnd.n3675 585
R756 gnd.n3723 gnd.n3677 585
R757 gnd.n3724 gnd.n3672 585
R758 gnd.n3725 gnd.n2192 585
R759 gnd.n5928 gnd.n2192 585
R760 gnd.n3927 gnd.n3926 585
R761 gnd.n3928 gnd.n3512 585
R762 gnd.n3929 gnd.n3508 585
R763 gnd.n3499 gnd.n3498 585
R764 gnd.n3936 gnd.n3497 585
R765 gnd.n3937 gnd.n3496 585
R766 gnd.n3495 gnd.n3489 585
R767 gnd.n3944 gnd.n3488 585
R768 gnd.n3945 gnd.n3487 585
R769 gnd.n3479 gnd.n3478 585
R770 gnd.n3952 gnd.n3477 585
R771 gnd.n3953 gnd.n3476 585
R772 gnd.n3475 gnd.n3469 585
R773 gnd.n3960 gnd.n3468 585
R774 gnd.n3961 gnd.n3467 585
R775 gnd.n3459 gnd.n3458 585
R776 gnd.n3968 gnd.n3457 585
R777 gnd.n3969 gnd.n3456 585
R778 gnd.n3455 gnd.n2475 585
R779 gnd.n5674 gnd.n2475 585
R780 gnd.n3925 gnd.n3520 585
R781 gnd.n3925 gnd.n3924 585
R782 gnd.n3865 gnd.n2466 585
R783 gnd.n5682 gnd.n2466 585
R784 gnd.n3869 gnd.n3864 585
R785 gnd.n3864 gnd.n3863 585
R786 gnd.n3870 gnd.n2456 585
R787 gnd.n5688 gnd.n2456 585
R788 gnd.n3871 gnd.n3651 585
R789 gnd.n3854 gnd.n3651 585
R790 gnd.n3649 gnd.n2445 585
R791 gnd.n5694 gnd.n2445 585
R792 gnd.n3875 gnd.n3648 585
R793 gnd.n3849 gnd.n3648 585
R794 gnd.n3876 gnd.n2435 585
R795 gnd.n5700 gnd.n2435 585
R796 gnd.n3877 gnd.n3647 585
R797 gnd.n3845 gnd.n3647 585
R798 gnd.n3644 gnd.n2424 585
R799 gnd.n5706 gnd.n2424 585
R800 gnd.n3882 gnd.n3881 585
R801 gnd.n3883 gnd.n3882 585
R802 gnd.n3643 gnd.n2415 585
R803 gnd.n5712 gnd.n2415 585
R804 gnd.n3837 gnd.n3836 585
R805 gnd.n3838 gnd.n3837 585
R806 gnd.n3654 gnd.n2404 585
R807 gnd.n5718 gnd.n2404 585
R808 gnd.n3832 gnd.n3831 585
R809 gnd.n3831 gnd.n3830 585
R810 gnd.n3780 gnd.n2395 585
R811 gnd.n5724 gnd.n2395 585
R812 gnd.n3779 gnd.n3657 585
R813 gnd.n3657 gnd.n2385 585
R814 gnd.n3656 gnd.n2384 585
R815 gnd.n5730 gnd.n2384 585
R816 gnd.n3775 gnd.n3774 585
R817 gnd.n3774 gnd.n2376 585
R818 gnd.n3773 gnd.n2375 585
R819 gnd.n5736 gnd.n2375 585
R820 gnd.n3772 gnd.n3660 585
R821 gnd.n3660 gnd.n2366 585
R822 gnd.n3659 gnd.n2365 585
R823 gnd.n5742 gnd.n2365 585
R824 gnd.n3768 gnd.n3767 585
R825 gnd.n3767 gnd.n2363 585
R826 gnd.n3766 gnd.n2356 585
R827 gnd.n5748 gnd.n2356 585
R828 gnd.n3765 gnd.n3764 585
R829 gnd.n3764 gnd.n2354 585
R830 gnd.n3662 gnd.n2346 585
R831 gnd.n5754 gnd.n2346 585
R832 gnd.n3760 gnd.n3759 585
R833 gnd.n3759 gnd.n2338 585
R834 gnd.n3758 gnd.n2337 585
R835 gnd.n5760 gnd.n2337 585
R836 gnd.n3757 gnd.n3756 585
R837 gnd.n3756 gnd.n2328 585
R838 gnd.n3664 gnd.n2327 585
R839 gnd.n5766 gnd.n2327 585
R840 gnd.n3752 gnd.n3751 585
R841 gnd.n3751 gnd.n2325 585
R842 gnd.n3750 gnd.n2318 585
R843 gnd.n5772 gnd.n2318 585
R844 gnd.n3749 gnd.n3748 585
R845 gnd.n3748 gnd.n2316 585
R846 gnd.n3666 gnd.n2308 585
R847 gnd.n5778 gnd.n2308 585
R848 gnd.n3744 gnd.n3743 585
R849 gnd.n3743 gnd.n2300 585
R850 gnd.n3742 gnd.n2299 585
R851 gnd.n5784 gnd.n2299 585
R852 gnd.n3741 gnd.n3740 585
R853 gnd.n3740 gnd.n2291 585
R854 gnd.n3668 gnd.n2290 585
R855 gnd.n5790 gnd.n2290 585
R856 gnd.n3736 gnd.n3735 585
R857 gnd.n3735 gnd.n2281 585
R858 gnd.n3734 gnd.n2280 585
R859 gnd.n5796 gnd.n2280 585
R860 gnd.n3733 gnd.n3732 585
R861 gnd.n3732 gnd.n2278 585
R862 gnd.n3670 gnd.n2270 585
R863 gnd.n5804 gnd.n2270 585
R864 gnd.n3728 gnd.n3727 585
R865 gnd.n3727 gnd.n2193 585
R866 gnd.n5990 gnd.n5989 585
R867 gnd.n5991 gnd.n5990 585
R868 gnd.n779 gnd.n777 585
R869 gnd.n777 gnd.n773 585
R870 gnd.n2144 gnd.n2143 585
R871 gnd.n2145 gnd.n2144 585
R872 gnd.n887 gnd.n886 585
R873 gnd.n886 gnd.n763 585
R874 gnd.n2133 gnd.n2132 585
R875 gnd.n2134 gnd.n2133 585
R876 gnd.n897 gnd.n896 585
R877 gnd.n902 gnd.n896 585
R878 gnd.n1854 gnd.n914 585
R879 gnd.n914 gnd.n901 585
R880 gnd.n1856 gnd.n1855 585
R881 gnd.n1857 gnd.n1856 585
R882 gnd.n915 gnd.n913 585
R883 gnd.n913 gnd.n909 585
R884 gnd.n1845 gnd.n1844 585
R885 gnd.n1846 gnd.n1845 585
R886 gnd.n922 gnd.n921 585
R887 gnd.n927 gnd.n921 585
R888 gnd.n1823 gnd.n940 585
R889 gnd.n940 gnd.n926 585
R890 gnd.n1825 gnd.n1824 585
R891 gnd.n1826 gnd.n1825 585
R892 gnd.n941 gnd.n939 585
R893 gnd.n939 gnd.n935 585
R894 gnd.n1814 gnd.n1813 585
R895 gnd.n1815 gnd.n1814 585
R896 gnd.n948 gnd.n947 585
R897 gnd.n952 gnd.n947 585
R898 gnd.n1792 gnd.n964 585
R899 gnd.n1097 gnd.n964 585
R900 gnd.n1794 gnd.n1793 585
R901 gnd.n1795 gnd.n1794 585
R902 gnd.n965 gnd.n963 585
R903 gnd.n963 gnd.n960 585
R904 gnd.n1783 gnd.n1782 585
R905 gnd.n1784 gnd.n1783 585
R906 gnd.n972 gnd.n971 585
R907 gnd.n977 gnd.n971 585
R908 gnd.n1761 gnd.n990 585
R909 gnd.n990 gnd.n976 585
R910 gnd.n1763 gnd.n1762 585
R911 gnd.n1764 gnd.n1763 585
R912 gnd.n991 gnd.n989 585
R913 gnd.n989 gnd.n985 585
R914 gnd.n1752 gnd.n1751 585
R915 gnd.n1753 gnd.n1752 585
R916 gnd.n999 gnd.n998 585
R917 gnd.n1004 gnd.n998 585
R918 gnd.n1730 gnd.n1016 585
R919 gnd.n1016 gnd.n1003 585
R920 gnd.n1732 gnd.n1731 585
R921 gnd.n1733 gnd.n1732 585
R922 gnd.n1017 gnd.n1015 585
R923 gnd.n1015 gnd.n1011 585
R924 gnd.n1721 gnd.n1720 585
R925 gnd.n1722 gnd.n1721 585
R926 gnd.n1024 gnd.n1023 585
R927 gnd.n1122 gnd.n1023 585
R928 gnd.n1699 gnd.n1039 585
R929 gnd.n1039 gnd.n1028 585
R930 gnd.n1701 gnd.n1700 585
R931 gnd.n1702 gnd.n1701 585
R932 gnd.n1040 gnd.n1038 585
R933 gnd.n1691 gnd.n1038 585
R934 gnd.n1191 gnd.n1190 585
R935 gnd.n1191 gnd.n1045 585
R936 gnd.n1678 gnd.n1677 585
R937 gnd.n1677 gnd.n1676 585
R938 gnd.n1679 gnd.n1183 585
R939 gnd.n1656 gnd.n1183 585
R940 gnd.n1681 gnd.n1680 585
R941 gnd.n1682 gnd.n1681 585
R942 gnd.n1184 gnd.n1182 585
R943 gnd.n1664 gnd.n1182 585
R944 gnd.n1648 gnd.n1647 585
R945 gnd.n1647 gnd.n1201 585
R946 gnd.n1646 gnd.n1206 585
R947 gnd.n1646 gnd.n1645 585
R948 gnd.n1631 gnd.n1207 585
R949 gnd.n1215 gnd.n1207 585
R950 gnd.n1633 gnd.n1632 585
R951 gnd.n1634 gnd.n1633 585
R952 gnd.n1218 gnd.n1217 585
R953 gnd.n1225 gnd.n1217 585
R954 gnd.n1606 gnd.n1605 585
R955 gnd.n1607 gnd.n1606 585
R956 gnd.n1237 gnd.n1236 585
R957 gnd.n1236 gnd.n1232 585
R958 gnd.n1596 gnd.n1595 585
R959 gnd.n1597 gnd.n1596 585
R960 gnd.n1247 gnd.n1246 585
R961 gnd.n1252 gnd.n1246 585
R962 gnd.n1574 gnd.n1265 585
R963 gnd.n1265 gnd.n1251 585
R964 gnd.n1576 gnd.n1575 585
R965 gnd.n1577 gnd.n1576 585
R966 gnd.n1266 gnd.n1264 585
R967 gnd.n1264 gnd.n1260 585
R968 gnd.n1565 gnd.n1564 585
R969 gnd.n1566 gnd.n1565 585
R970 gnd.n1273 gnd.n1272 585
R971 gnd.n1277 gnd.n1272 585
R972 gnd.n1542 gnd.n1294 585
R973 gnd.n1294 gnd.n1276 585
R974 gnd.n1544 gnd.n1543 585
R975 gnd.n1545 gnd.n1544 585
R976 gnd.n1295 gnd.n1293 585
R977 gnd.n1293 gnd.n1284 585
R978 gnd.n1537 gnd.n1536 585
R979 gnd.n1536 gnd.n1535 585
R980 gnd.n1342 gnd.n1341 585
R981 gnd.n1343 gnd.n1342 585
R982 gnd.n1496 gnd.n1495 585
R983 gnd.n1497 gnd.n1496 585
R984 gnd.n1352 gnd.n1351 585
R985 gnd.n1351 gnd.n1350 585
R986 gnd.n1491 gnd.n1490 585
R987 gnd.n1490 gnd.n1489 585
R988 gnd.n1355 gnd.n1354 585
R989 gnd.n1356 gnd.n1355 585
R990 gnd.n1480 gnd.n1479 585
R991 gnd.n1481 gnd.n1480 585
R992 gnd.n1363 gnd.n1362 585
R993 gnd.n1472 gnd.n1362 585
R994 gnd.n1475 gnd.n1474 585
R995 gnd.n1474 gnd.n1473 585
R996 gnd.n1366 gnd.n1365 585
R997 gnd.n1367 gnd.n1366 585
R998 gnd.n1461 gnd.n1460 585
R999 gnd.n1459 gnd.n1385 585
R1000 gnd.n1458 gnd.n1384 585
R1001 gnd.n1463 gnd.n1384 585
R1002 gnd.n1457 gnd.n1456 585
R1003 gnd.n1455 gnd.n1454 585
R1004 gnd.n1453 gnd.n1452 585
R1005 gnd.n1451 gnd.n1450 585
R1006 gnd.n1449 gnd.n1448 585
R1007 gnd.n1447 gnd.n1446 585
R1008 gnd.n1445 gnd.n1444 585
R1009 gnd.n1443 gnd.n1442 585
R1010 gnd.n1441 gnd.n1440 585
R1011 gnd.n1439 gnd.n1438 585
R1012 gnd.n1437 gnd.n1436 585
R1013 gnd.n1435 gnd.n1434 585
R1014 gnd.n1433 gnd.n1432 585
R1015 gnd.n1431 gnd.n1430 585
R1016 gnd.n1429 gnd.n1428 585
R1017 gnd.n1427 gnd.n1426 585
R1018 gnd.n1425 gnd.n1424 585
R1019 gnd.n1423 gnd.n1422 585
R1020 gnd.n1421 gnd.n1420 585
R1021 gnd.n1419 gnd.n1418 585
R1022 gnd.n1417 gnd.n1416 585
R1023 gnd.n1415 gnd.n1414 585
R1024 gnd.n1372 gnd.n1371 585
R1025 gnd.n1466 gnd.n1465 585
R1026 gnd.n2153 gnd.n2152 585
R1027 gnd.n803 gnd.n802 585
R1028 gnd.n879 gnd.n878 585
R1029 gnd.n877 gnd.n876 585
R1030 gnd.n875 gnd.n874 585
R1031 gnd.n868 gnd.n808 585
R1032 gnd.n870 gnd.n869 585
R1033 gnd.n867 gnd.n866 585
R1034 gnd.n865 gnd.n864 585
R1035 gnd.n858 gnd.n810 585
R1036 gnd.n860 gnd.n859 585
R1037 gnd.n857 gnd.n856 585
R1038 gnd.n855 gnd.n854 585
R1039 gnd.n848 gnd.n812 585
R1040 gnd.n850 gnd.n849 585
R1041 gnd.n847 gnd.n846 585
R1042 gnd.n845 gnd.n844 585
R1043 gnd.n838 gnd.n814 585
R1044 gnd.n840 gnd.n839 585
R1045 gnd.n837 gnd.n836 585
R1046 gnd.n835 gnd.n834 585
R1047 gnd.n828 gnd.n816 585
R1048 gnd.n830 gnd.n829 585
R1049 gnd.n827 gnd.n826 585
R1050 gnd.n825 gnd.n824 585
R1051 gnd.n819 gnd.n818 585
R1052 gnd.n820 gnd.n778 585
R1053 gnd.n5975 gnd.n778 585
R1054 gnd.n2149 gnd.n775 585
R1055 gnd.n5991 gnd.n775 585
R1056 gnd.n2148 gnd.n2147 585
R1057 gnd.n2147 gnd.n773 585
R1058 gnd.n2146 gnd.n883 585
R1059 gnd.n2146 gnd.n2145 585
R1060 gnd.n1076 gnd.n884 585
R1061 gnd.n884 gnd.n763 585
R1062 gnd.n1077 gnd.n895 585
R1063 gnd.n2134 gnd.n895 585
R1064 gnd.n1079 gnd.n1078 585
R1065 gnd.n1079 gnd.n902 585
R1066 gnd.n1081 gnd.n1080 585
R1067 gnd.n1080 gnd.n901 585
R1068 gnd.n1082 gnd.n911 585
R1069 gnd.n1857 gnd.n911 585
R1070 gnd.n1084 gnd.n1083 585
R1071 gnd.n1083 gnd.n909 585
R1072 gnd.n1085 gnd.n920 585
R1073 gnd.n1846 gnd.n920 585
R1074 gnd.n1087 gnd.n1086 585
R1075 gnd.n1087 gnd.n927 585
R1076 gnd.n1089 gnd.n1088 585
R1077 gnd.n1088 gnd.n926 585
R1078 gnd.n1090 gnd.n937 585
R1079 gnd.n1826 gnd.n937 585
R1080 gnd.n1092 gnd.n1091 585
R1081 gnd.n1091 gnd.n935 585
R1082 gnd.n1093 gnd.n946 585
R1083 gnd.n1815 gnd.n946 585
R1084 gnd.n1095 gnd.n1094 585
R1085 gnd.n1095 gnd.n952 585
R1086 gnd.n1099 gnd.n1098 585
R1087 gnd.n1098 gnd.n1097 585
R1088 gnd.n1100 gnd.n962 585
R1089 gnd.n1795 gnd.n962 585
R1090 gnd.n1102 gnd.n1101 585
R1091 gnd.n1101 gnd.n960 585
R1092 gnd.n1103 gnd.n970 585
R1093 gnd.n1784 gnd.n970 585
R1094 gnd.n1105 gnd.n1104 585
R1095 gnd.n1105 gnd.n977 585
R1096 gnd.n1107 gnd.n1106 585
R1097 gnd.n1106 gnd.n976 585
R1098 gnd.n1108 gnd.n987 585
R1099 gnd.n1764 gnd.n987 585
R1100 gnd.n1110 gnd.n1109 585
R1101 gnd.n1109 gnd.n985 585
R1102 gnd.n1111 gnd.n997 585
R1103 gnd.n1753 gnd.n997 585
R1104 gnd.n1113 gnd.n1112 585
R1105 gnd.n1113 gnd.n1004 585
R1106 gnd.n1115 gnd.n1114 585
R1107 gnd.n1114 gnd.n1003 585
R1108 gnd.n1116 gnd.n1013 585
R1109 gnd.n1733 gnd.n1013 585
R1110 gnd.n1118 gnd.n1117 585
R1111 gnd.n1117 gnd.n1011 585
R1112 gnd.n1119 gnd.n1022 585
R1113 gnd.n1722 gnd.n1022 585
R1114 gnd.n1124 gnd.n1123 585
R1115 gnd.n1123 gnd.n1122 585
R1116 gnd.n1120 gnd.n1048 585
R1117 gnd.n1120 gnd.n1028 585
R1118 gnd.n1688 gnd.n1036 585
R1119 gnd.n1702 gnd.n1036 585
R1120 gnd.n1690 gnd.n1689 585
R1121 gnd.n1691 gnd.n1690 585
R1122 gnd.n1192 gnd.n1046 585
R1123 gnd.n1046 gnd.n1045 585
R1124 gnd.n1194 gnd.n1193 585
R1125 gnd.n1676 gnd.n1194 585
R1126 gnd.n1179 gnd.n1177 585
R1127 gnd.n1656 gnd.n1179 585
R1128 gnd.n1684 gnd.n1683 585
R1129 gnd.n1683 gnd.n1682 585
R1130 gnd.n1178 gnd.n1176 585
R1131 gnd.n1664 gnd.n1178 585
R1132 gnd.n1641 gnd.n1210 585
R1133 gnd.n1210 gnd.n1201 585
R1134 gnd.n1643 gnd.n1642 585
R1135 gnd.n1645 gnd.n1643 585
R1136 gnd.n1211 gnd.n1209 585
R1137 gnd.n1215 gnd.n1209 585
R1138 gnd.n1636 gnd.n1635 585
R1139 gnd.n1635 gnd.n1634 585
R1140 gnd.n1214 gnd.n1213 585
R1141 gnd.n1225 gnd.n1214 585
R1142 gnd.n1515 gnd.n1234 585
R1143 gnd.n1607 gnd.n1234 585
R1144 gnd.n1517 gnd.n1516 585
R1145 gnd.n1516 gnd.n1232 585
R1146 gnd.n1518 gnd.n1245 585
R1147 gnd.n1597 gnd.n1245 585
R1148 gnd.n1520 gnd.n1519 585
R1149 gnd.n1520 gnd.n1252 585
R1150 gnd.n1522 gnd.n1521 585
R1151 gnd.n1521 gnd.n1251 585
R1152 gnd.n1523 gnd.n1262 585
R1153 gnd.n1577 gnd.n1262 585
R1154 gnd.n1525 gnd.n1524 585
R1155 gnd.n1524 gnd.n1260 585
R1156 gnd.n1526 gnd.n1271 585
R1157 gnd.n1566 gnd.n1271 585
R1158 gnd.n1528 gnd.n1527 585
R1159 gnd.n1528 gnd.n1277 585
R1160 gnd.n1530 gnd.n1529 585
R1161 gnd.n1529 gnd.n1276 585
R1162 gnd.n1531 gnd.n1292 585
R1163 gnd.n1545 gnd.n1292 585
R1164 gnd.n1532 gnd.n1345 585
R1165 gnd.n1345 gnd.n1284 585
R1166 gnd.n1534 gnd.n1533 585
R1167 gnd.n1535 gnd.n1534 585
R1168 gnd.n1346 gnd.n1344 585
R1169 gnd.n1344 gnd.n1343 585
R1170 gnd.n1499 gnd.n1498 585
R1171 gnd.n1498 gnd.n1497 585
R1172 gnd.n1349 gnd.n1348 585
R1173 gnd.n1350 gnd.n1349 585
R1174 gnd.n1488 gnd.n1487 585
R1175 gnd.n1489 gnd.n1488 585
R1176 gnd.n1358 gnd.n1357 585
R1177 gnd.n1357 gnd.n1356 585
R1178 gnd.n1483 gnd.n1482 585
R1179 gnd.n1482 gnd.n1481 585
R1180 gnd.n1361 gnd.n1360 585
R1181 gnd.n1472 gnd.n1361 585
R1182 gnd.n1471 gnd.n1470 585
R1183 gnd.n1473 gnd.n1471 585
R1184 gnd.n1369 gnd.n1368 585
R1185 gnd.n1368 gnd.n1367 585
R1186 gnd.n7207 gnd.n166 585
R1187 gnd.n166 gnd.n165 585
R1188 gnd.n7209 gnd.n7208 585
R1189 gnd.n7210 gnd.n7209 585
R1190 gnd.n152 gnd.n151 585
R1191 gnd.n155 gnd.n152 585
R1192 gnd.n7218 gnd.n7217 585
R1193 gnd.n7217 gnd.n7216 585
R1194 gnd.n7219 gnd.n147 585
R1195 gnd.n147 gnd.n146 585
R1196 gnd.n7221 gnd.n7220 585
R1197 gnd.n7222 gnd.n7221 585
R1198 gnd.n132 gnd.n131 585
R1199 gnd.n143 gnd.n132 585
R1200 gnd.n7230 gnd.n7229 585
R1201 gnd.n7229 gnd.n7228 585
R1202 gnd.n7231 gnd.n127 585
R1203 gnd.n127 gnd.n126 585
R1204 gnd.n7233 gnd.n7232 585
R1205 gnd.n7234 gnd.n7233 585
R1206 gnd.n113 gnd.n112 585
R1207 gnd.n116 gnd.n113 585
R1208 gnd.n7242 gnd.n7241 585
R1209 gnd.n7241 gnd.n7240 585
R1210 gnd.n7243 gnd.n108 585
R1211 gnd.n108 gnd.n107 585
R1212 gnd.n7245 gnd.n7244 585
R1213 gnd.n7246 gnd.n7245 585
R1214 gnd.n94 gnd.n93 585
R1215 gnd.n104 gnd.n94 585
R1216 gnd.n7254 gnd.n7253 585
R1217 gnd.n7253 gnd.n7252 585
R1218 gnd.n7255 gnd.n88 585
R1219 gnd.n88 gnd.n86 585
R1220 gnd.n7257 gnd.n7256 585
R1221 gnd.n7258 gnd.n7257 585
R1222 gnd.n89 gnd.n87 585
R1223 gnd.n87 gnd.n74 585
R1224 gnd.n6840 gnd.n75 585
R1225 gnd.n7264 gnd.n75 585
R1226 gnd.n6839 gnd.n6838 585
R1227 gnd.n6838 gnd.n6837 585
R1228 gnd.n171 gnd.n170 585
R1229 gnd.n172 gnd.n171 585
R1230 gnd.n6831 gnd.n6830 585
R1231 gnd.n6830 gnd.n6829 585
R1232 gnd.n177 gnd.n176 585
R1233 gnd.n189 gnd.n177 585
R1234 gnd.n6817 gnd.n6816 585
R1235 gnd.n6818 gnd.n6817 585
R1236 gnd.n191 gnd.n190 585
R1237 gnd.n6809 gnd.n190 585
R1238 gnd.n6781 gnd.n6780 585
R1239 gnd.n6780 gnd.n195 585
R1240 gnd.n6782 gnd.n204 585
R1241 gnd.n6796 gnd.n204 585
R1242 gnd.n6783 gnd.n216 585
R1243 gnd.n6774 gnd.n216 585
R1244 gnd.n6785 gnd.n6784 585
R1245 gnd.n6786 gnd.n6785 585
R1246 gnd.n217 gnd.n215 585
R1247 gnd.n6770 gnd.n215 585
R1248 gnd.n6746 gnd.n6745 585
R1249 gnd.n6745 gnd.n6744 585
R1250 gnd.n6747 gnd.n232 585
R1251 gnd.n6761 gnd.n232 585
R1252 gnd.n6748 gnd.n244 585
R1253 gnd.n5102 gnd.n244 585
R1254 gnd.n6750 gnd.n6749 585
R1255 gnd.n6751 gnd.n6750 585
R1256 gnd.n245 gnd.n243 585
R1257 gnd.n5170 gnd.n243 585
R1258 gnd.n5175 gnd.n5097 585
R1259 gnd.n5128 gnd.n5097 585
R1260 gnd.n5177 gnd.n5176 585
R1261 gnd.n5178 gnd.n5177 585
R1262 gnd.n5098 gnd.n5096 585
R1263 gnd.n5160 gnd.n5096 585
R1264 gnd.n5154 gnd.n5076 585
R1265 gnd.n5184 gnd.n5076 585
R1266 gnd.n5153 gnd.n5152 585
R1267 gnd.n5152 gnd.n5072 585
R1268 gnd.n5151 gnd.n2884 585
R1269 gnd.n2890 gnd.n2884 585
R1270 gnd.n5193 gnd.n2885 585
R1271 gnd.n5193 gnd.n5192 585
R1272 gnd.n5195 gnd.n5194 585
R1273 gnd.n5273 gnd.n5196 585
R1274 gnd.n5272 gnd.n5197 585
R1275 gnd.n5204 gnd.n5198 585
R1276 gnd.n5265 gnd.n5205 585
R1277 gnd.n5264 gnd.n5206 585
R1278 gnd.n5208 gnd.n5207 585
R1279 gnd.n5257 gnd.n5216 585
R1280 gnd.n5256 gnd.n5217 585
R1281 gnd.n5224 gnd.n5218 585
R1282 gnd.n5249 gnd.n5225 585
R1283 gnd.n5248 gnd.n5226 585
R1284 gnd.n5228 gnd.n5227 585
R1285 gnd.n5241 gnd.n5236 585
R1286 gnd.n5240 gnd.n5237 585
R1287 gnd.n2802 gnd.n2755 585
R1288 gnd.n5403 gnd.n2756 585
R1289 gnd.n5402 gnd.n5399 585
R1290 gnd.n2765 gnd.n2757 585
R1291 gnd.n5397 gnd.n2765 585
R1292 gnd.n6992 gnd.n6991 585
R1293 gnd.n6894 gnd.n6890 585
R1294 gnd.n6942 gnd.n6941 585
R1295 gnd.n6940 gnd.n6939 585
R1296 gnd.n6938 gnd.n6937 585
R1297 gnd.n6931 gnd.n6896 585
R1298 gnd.n6933 gnd.n6932 585
R1299 gnd.n6930 gnd.n6929 585
R1300 gnd.n6928 gnd.n6927 585
R1301 gnd.n6921 gnd.n6898 585
R1302 gnd.n6923 gnd.n6922 585
R1303 gnd.n6920 gnd.n6919 585
R1304 gnd.n6918 gnd.n6917 585
R1305 gnd.n6911 gnd.n6900 585
R1306 gnd.n6913 gnd.n6912 585
R1307 gnd.n6910 gnd.n6909 585
R1308 gnd.n6908 gnd.n6907 585
R1309 gnd.n6904 gnd.n6903 585
R1310 gnd.n6902 gnd.n6881 585
R1311 gnd.n7199 gnd.n6881 585
R1312 gnd.n6988 gnd.n6891 585
R1313 gnd.n6891 gnd.n165 585
R1314 gnd.n6987 gnd.n164 585
R1315 gnd.n7210 gnd.n164 585
R1316 gnd.n6986 gnd.n6985 585
R1317 gnd.n6985 gnd.n155 585
R1318 gnd.n6946 gnd.n154 585
R1319 gnd.n7216 gnd.n154 585
R1320 gnd.n6981 gnd.n6980 585
R1321 gnd.n6980 gnd.n146 585
R1322 gnd.n6979 gnd.n145 585
R1323 gnd.n7222 gnd.n145 585
R1324 gnd.n6978 gnd.n6977 585
R1325 gnd.n6977 gnd.n143 585
R1326 gnd.n6948 gnd.n134 585
R1327 gnd.n7228 gnd.n134 585
R1328 gnd.n6973 gnd.n6972 585
R1329 gnd.n6972 gnd.n126 585
R1330 gnd.n6971 gnd.n125 585
R1331 gnd.n7234 gnd.n125 585
R1332 gnd.n6970 gnd.n6969 585
R1333 gnd.n6969 gnd.n116 585
R1334 gnd.n6950 gnd.n115 585
R1335 gnd.n7240 gnd.n115 585
R1336 gnd.n6965 gnd.n6964 585
R1337 gnd.n6964 gnd.n107 585
R1338 gnd.n6963 gnd.n106 585
R1339 gnd.n7246 gnd.n106 585
R1340 gnd.n6962 gnd.n6961 585
R1341 gnd.n6961 gnd.n104 585
R1342 gnd.n6952 gnd.n96 585
R1343 gnd.n7252 gnd.n96 585
R1344 gnd.n6957 gnd.n6956 585
R1345 gnd.n6956 gnd.n86 585
R1346 gnd.n6955 gnd.n85 585
R1347 gnd.n7258 gnd.n85 585
R1348 gnd.n72 gnd.n71 585
R1349 gnd.n74 gnd.n72 585
R1350 gnd.n7266 gnd.n7265 585
R1351 gnd.n7265 gnd.n7264 585
R1352 gnd.n7267 gnd.n70 585
R1353 gnd.n6837 gnd.n70 585
R1354 gnd.n179 gnd.n68 585
R1355 gnd.n179 gnd.n172 585
R1356 gnd.n6802 gnd.n180 585
R1357 gnd.n6829 gnd.n180 585
R1358 gnd.n6803 gnd.n6801 585
R1359 gnd.n6801 gnd.n189 585
R1360 gnd.n198 gnd.n188 585
R1361 gnd.n6818 gnd.n188 585
R1362 gnd.n6808 gnd.n6807 585
R1363 gnd.n6809 gnd.n6808 585
R1364 gnd.n197 gnd.n196 585
R1365 gnd.n196 gnd.n195 585
R1366 gnd.n6798 gnd.n6797 585
R1367 gnd.n6797 gnd.n6796 585
R1368 gnd.n201 gnd.n200 585
R1369 gnd.n6774 gnd.n201 585
R1370 gnd.n225 gnd.n213 585
R1371 gnd.n6786 gnd.n213 585
R1372 gnd.n6769 gnd.n6768 585
R1373 gnd.n6770 gnd.n6769 585
R1374 gnd.n224 gnd.n223 585
R1375 gnd.n6744 gnd.n223 585
R1376 gnd.n6763 gnd.n6762 585
R1377 gnd.n6762 gnd.n6761 585
R1378 gnd.n228 gnd.n227 585
R1379 gnd.n5102 gnd.n228 585
R1380 gnd.n5131 gnd.n241 585
R1381 gnd.n6751 gnd.n241 585
R1382 gnd.n5169 gnd.n5168 585
R1383 gnd.n5170 gnd.n5169 585
R1384 gnd.n5130 gnd.n5129 585
R1385 gnd.n5129 gnd.n5128 585
R1386 gnd.n5163 gnd.n5094 585
R1387 gnd.n5178 gnd.n5094 585
R1388 gnd.n5162 gnd.n5161 585
R1389 gnd.n5161 gnd.n5160 585
R1390 gnd.n5142 gnd.n5074 585
R1391 gnd.n5184 gnd.n5074 585
R1392 gnd.n5136 gnd.n5133 585
R1393 gnd.n5136 gnd.n5072 585
R1394 gnd.n5138 gnd.n5137 585
R1395 gnd.n5137 gnd.n2890 585
R1396 gnd.n5135 gnd.n2889 585
R1397 gnd.n5192 gnd.n2889 585
R1398 gnd.n772 gnd.n771 585
R1399 gnd.n776 gnd.n772 585
R1400 gnd.n5994 gnd.n5993 585
R1401 gnd.n5993 gnd.n5992 585
R1402 gnd.n5995 gnd.n766 585
R1403 gnd.n885 gnd.n766 585
R1404 gnd.n5997 gnd.n5996 585
R1405 gnd.n5998 gnd.n5997 585
R1406 gnd.n767 gnd.n765 585
R1407 gnd.n2135 gnd.n765 585
R1408 gnd.n1866 gnd.n904 585
R1409 gnd.n904 gnd.n894 585
R1410 gnd.n1868 gnd.n1867 585
R1411 gnd.n1869 gnd.n1868 585
R1412 gnd.n905 gnd.n903 585
R1413 gnd.n912 gnd.n903 585
R1414 gnd.n1860 gnd.n1859 585
R1415 gnd.n1859 gnd.n1858 585
R1416 gnd.n908 gnd.n907 585
R1417 gnd.n1847 gnd.n908 585
R1418 gnd.n1834 gnd.n930 585
R1419 gnd.n930 gnd.n929 585
R1420 gnd.n1836 gnd.n1835 585
R1421 gnd.n1837 gnd.n1836 585
R1422 gnd.n931 gnd.n928 585
R1423 gnd.n938 gnd.n928 585
R1424 gnd.n1829 gnd.n1828 585
R1425 gnd.n1828 gnd.n1827 585
R1426 gnd.n934 gnd.n933 585
R1427 gnd.n1816 gnd.n934 585
R1428 gnd.n1803 gnd.n955 585
R1429 gnd.n955 gnd.n954 585
R1430 gnd.n1805 gnd.n1804 585
R1431 gnd.n1806 gnd.n1805 585
R1432 gnd.n956 gnd.n953 585
R1433 gnd.n1096 gnd.n953 585
R1434 gnd.n1798 gnd.n1797 585
R1435 gnd.n1797 gnd.n1796 585
R1436 gnd.n959 gnd.n958 585
R1437 gnd.n1785 gnd.n959 585
R1438 gnd.n1772 gnd.n980 585
R1439 gnd.n980 gnd.n979 585
R1440 gnd.n1774 gnd.n1773 585
R1441 gnd.n1775 gnd.n1774 585
R1442 gnd.n981 gnd.n978 585
R1443 gnd.n988 gnd.n978 585
R1444 gnd.n1767 gnd.n1766 585
R1445 gnd.n1766 gnd.n1765 585
R1446 gnd.n984 gnd.n983 585
R1447 gnd.n1754 gnd.n984 585
R1448 gnd.n1741 gnd.n1006 585
R1449 gnd.n1006 gnd.n996 585
R1450 gnd.n1743 gnd.n1742 585
R1451 gnd.n1744 gnd.n1743 585
R1452 gnd.n1007 gnd.n1005 585
R1453 gnd.n1014 gnd.n1005 585
R1454 gnd.n1736 gnd.n1735 585
R1455 gnd.n1735 gnd.n1734 585
R1456 gnd.n1010 gnd.n1009 585
R1457 gnd.n1723 gnd.n1010 585
R1458 gnd.n1710 gnd.n1030 585
R1459 gnd.n1121 gnd.n1030 585
R1460 gnd.n1712 gnd.n1711 585
R1461 gnd.n1713 gnd.n1712 585
R1462 gnd.n1031 gnd.n1029 585
R1463 gnd.n1037 gnd.n1029 585
R1464 gnd.n1705 gnd.n1704 585
R1465 gnd.n1704 gnd.n1703 585
R1466 gnd.n1034 gnd.n1033 585
R1467 gnd.n1692 gnd.n1034 585
R1468 gnd.n1674 gnd.n1673 585
R1469 gnd.n1675 gnd.n1674 585
R1470 gnd.n1196 gnd.n1195 585
R1471 gnd.n1657 gnd.n1195 585
R1472 gnd.n1669 gnd.n1668 585
R1473 gnd.n1668 gnd.n1181 585
R1474 gnd.n1667 gnd.n1198 585
R1475 gnd.n1667 gnd.n1180 585
R1476 gnd.n1666 gnd.n1200 585
R1477 gnd.n1666 gnd.n1665 585
R1478 gnd.n1618 gnd.n1199 585
R1479 gnd.n1644 gnd.n1199 585
R1480 gnd.n1620 gnd.n1619 585
R1481 gnd.n1619 gnd.n1208 585
R1482 gnd.n1621 gnd.n1227 585
R1483 gnd.n1227 gnd.n1216 585
R1484 gnd.n1623 gnd.n1622 585
R1485 gnd.n1624 gnd.n1623 585
R1486 gnd.n1228 gnd.n1226 585
R1487 gnd.n1235 gnd.n1226 585
R1488 gnd.n1610 gnd.n1609 585
R1489 gnd.n1609 gnd.n1608 585
R1490 gnd.n1231 gnd.n1230 585
R1491 gnd.n1598 gnd.n1231 585
R1492 gnd.n1585 gnd.n1255 585
R1493 gnd.n1255 gnd.n1254 585
R1494 gnd.n1587 gnd.n1586 585
R1495 gnd.n1588 gnd.n1587 585
R1496 gnd.n1256 gnd.n1253 585
R1497 gnd.n1263 gnd.n1253 585
R1498 gnd.n1580 gnd.n1579 585
R1499 gnd.n1579 gnd.n1578 585
R1500 gnd.n1259 gnd.n1258 585
R1501 gnd.n1567 gnd.n1259 585
R1502 gnd.n1554 gnd.n1280 585
R1503 gnd.n1280 gnd.n1279 585
R1504 gnd.n1556 gnd.n1555 585
R1505 gnd.n1557 gnd.n1556 585
R1506 gnd.n1550 gnd.n1278 585
R1507 gnd.n1549 gnd.n1548 585
R1508 gnd.n1283 gnd.n1282 585
R1509 gnd.n1546 gnd.n1283 585
R1510 gnd.n1305 gnd.n1304 585
R1511 gnd.n1308 gnd.n1307 585
R1512 gnd.n1306 gnd.n1301 585
R1513 gnd.n1313 gnd.n1312 585
R1514 gnd.n1315 gnd.n1314 585
R1515 gnd.n1318 gnd.n1317 585
R1516 gnd.n1316 gnd.n1299 585
R1517 gnd.n1323 gnd.n1322 585
R1518 gnd.n1325 gnd.n1324 585
R1519 gnd.n1328 gnd.n1327 585
R1520 gnd.n1326 gnd.n1297 585
R1521 gnd.n1333 gnd.n1332 585
R1522 gnd.n1337 gnd.n1334 585
R1523 gnd.n1338 gnd.n1275 585
R1524 gnd.n5984 gnd.n5983 585
R1525 gnd.n5977 gnd.n786 585
R1526 gnd.n5979 gnd.n5978 585
R1527 gnd.n789 gnd.n788 585
R1528 gnd.n5949 gnd.n5948 585
R1529 gnd.n5951 gnd.n5950 585
R1530 gnd.n5953 gnd.n5952 585
R1531 gnd.n5955 gnd.n5954 585
R1532 gnd.n5957 gnd.n5956 585
R1533 gnd.n5959 gnd.n5958 585
R1534 gnd.n5961 gnd.n5960 585
R1535 gnd.n5963 gnd.n5962 585
R1536 gnd.n5965 gnd.n5964 585
R1537 gnd.n5968 gnd.n5967 585
R1538 gnd.n5966 gnd.n5938 585
R1539 gnd.n5972 gnd.n5935 585
R1540 gnd.n5974 gnd.n5973 585
R1541 gnd.n5975 gnd.n5974 585
R1542 gnd.n5986 gnd.n5985 585
R1543 gnd.n5985 gnd.n776 585
R1544 gnd.n782 gnd.n774 585
R1545 gnd.n5992 gnd.n774 585
R1546 gnd.n2140 gnd.n2139 585
R1547 gnd.n2139 gnd.n885 585
R1548 gnd.n2138 gnd.n764 585
R1549 gnd.n5998 gnd.n764 585
R1550 gnd.n2137 gnd.n2136 585
R1551 gnd.n2136 gnd.n2135 585
R1552 gnd.n893 gnd.n890 585
R1553 gnd.n894 gnd.n893 585
R1554 gnd.n1871 gnd.n1870 585
R1555 gnd.n1870 gnd.n1869 585
R1556 gnd.n900 gnd.n899 585
R1557 gnd.n912 gnd.n900 585
R1558 gnd.n1850 gnd.n910 585
R1559 gnd.n1858 gnd.n910 585
R1560 gnd.n1849 gnd.n1848 585
R1561 gnd.n1848 gnd.n1847 585
R1562 gnd.n919 gnd.n917 585
R1563 gnd.n929 gnd.n919 585
R1564 gnd.n1839 gnd.n1838 585
R1565 gnd.n1838 gnd.n1837 585
R1566 gnd.n925 gnd.n924 585
R1567 gnd.n938 gnd.n925 585
R1568 gnd.n1819 gnd.n936 585
R1569 gnd.n1827 gnd.n936 585
R1570 gnd.n1818 gnd.n1817 585
R1571 gnd.n1817 gnd.n1816 585
R1572 gnd.n945 gnd.n943 585
R1573 gnd.n954 gnd.n945 585
R1574 gnd.n1808 gnd.n1807 585
R1575 gnd.n1807 gnd.n1806 585
R1576 gnd.n951 gnd.n950 585
R1577 gnd.n1096 gnd.n951 585
R1578 gnd.n1788 gnd.n961 585
R1579 gnd.n1796 gnd.n961 585
R1580 gnd.n1787 gnd.n1786 585
R1581 gnd.n1786 gnd.n1785 585
R1582 gnd.n969 gnd.n967 585
R1583 gnd.n979 gnd.n969 585
R1584 gnd.n1777 gnd.n1776 585
R1585 gnd.n1776 gnd.n1775 585
R1586 gnd.n975 gnd.n974 585
R1587 gnd.n988 gnd.n975 585
R1588 gnd.n1757 gnd.n986 585
R1589 gnd.n1765 gnd.n986 585
R1590 gnd.n1756 gnd.n1755 585
R1591 gnd.n1755 gnd.n1754 585
R1592 gnd.n995 gnd.n993 585
R1593 gnd.n996 gnd.n995 585
R1594 gnd.n1746 gnd.n1745 585
R1595 gnd.n1745 gnd.n1744 585
R1596 gnd.n1002 gnd.n1001 585
R1597 gnd.n1014 gnd.n1002 585
R1598 gnd.n1726 gnd.n1012 585
R1599 gnd.n1734 gnd.n1012 585
R1600 gnd.n1725 gnd.n1724 585
R1601 gnd.n1724 gnd.n1723 585
R1602 gnd.n1021 gnd.n1019 585
R1603 gnd.n1121 gnd.n1021 585
R1604 gnd.n1715 gnd.n1714 585
R1605 gnd.n1714 gnd.n1713 585
R1606 gnd.n1027 gnd.n1026 585
R1607 gnd.n1037 gnd.n1027 585
R1608 gnd.n1695 gnd.n1035 585
R1609 gnd.n1703 gnd.n1035 585
R1610 gnd.n1694 gnd.n1693 585
R1611 gnd.n1693 gnd.n1692 585
R1612 gnd.n1044 gnd.n1042 585
R1613 gnd.n1675 gnd.n1044 585
R1614 gnd.n1658 gnd.n1655 585
R1615 gnd.n1658 gnd.n1657 585
R1616 gnd.n1660 gnd.n1659 585
R1617 gnd.n1659 gnd.n1181 585
R1618 gnd.n1661 gnd.n1203 585
R1619 gnd.n1203 gnd.n1180 585
R1620 gnd.n1663 gnd.n1662 585
R1621 gnd.n1665 gnd.n1663 585
R1622 gnd.n1204 gnd.n1202 585
R1623 gnd.n1644 gnd.n1202 585
R1624 gnd.n1628 gnd.n1627 585
R1625 gnd.n1627 gnd.n1208 585
R1626 gnd.n1626 gnd.n1222 585
R1627 gnd.n1626 gnd.n1216 585
R1628 gnd.n1625 gnd.n1224 585
R1629 gnd.n1625 gnd.n1624 585
R1630 gnd.n1602 gnd.n1223 585
R1631 gnd.n1235 gnd.n1223 585
R1632 gnd.n1601 gnd.n1233 585
R1633 gnd.n1608 gnd.n1233 585
R1634 gnd.n1600 gnd.n1599 585
R1635 gnd.n1599 gnd.n1598 585
R1636 gnd.n1244 gnd.n1241 585
R1637 gnd.n1254 gnd.n1244 585
R1638 gnd.n1590 gnd.n1589 585
R1639 gnd.n1589 gnd.n1588 585
R1640 gnd.n1250 gnd.n1249 585
R1641 gnd.n1263 gnd.n1250 585
R1642 gnd.n1570 gnd.n1261 585
R1643 gnd.n1578 gnd.n1261 585
R1644 gnd.n1569 gnd.n1568 585
R1645 gnd.n1568 gnd.n1567 585
R1646 gnd.n1270 gnd.n1268 585
R1647 gnd.n1279 gnd.n1270 585
R1648 gnd.n1559 gnd.n1558 585
R1649 gnd.n1558 gnd.n1557 585
R1650 gnd.n4909 gnd.n4908 585
R1651 gnd.n4910 gnd.n4909 585
R1652 gnd.n4820 gnd.n2977 585
R1653 gnd.n2983 gnd.n2977 585
R1654 gnd.n4819 gnd.n4818 585
R1655 gnd.n4818 gnd.n4817 585
R1656 gnd.n2980 gnd.n2979 585
R1657 gnd.n2991 gnd.n2980 585
R1658 gnd.n4805 gnd.n4804 585
R1659 gnd.n4806 gnd.n4805 585
R1660 gnd.n4803 gnd.n2992 585
R1661 gnd.n4798 gnd.n2992 585
R1662 gnd.n4802 gnd.n4801 585
R1663 gnd.n4801 gnd.n4800 585
R1664 gnd.n2994 gnd.n2993 585
R1665 gnd.n2995 gnd.n2994 585
R1666 gnd.n4785 gnd.n4784 585
R1667 gnd.n4786 gnd.n4785 585
R1668 gnd.n4783 gnd.n3001 585
R1669 gnd.n4779 gnd.n3001 585
R1670 gnd.n4782 gnd.n4781 585
R1671 gnd.n4781 gnd.n4780 585
R1672 gnd.n3003 gnd.n3002 585
R1673 gnd.n4733 gnd.n3003 585
R1674 gnd.n4771 gnd.n4770 585
R1675 gnd.n4772 gnd.n4771 585
R1676 gnd.n4769 gnd.n3010 585
R1677 gnd.n3010 gnd.n3009 585
R1678 gnd.n4768 gnd.n4767 585
R1679 gnd.n4767 gnd.n4766 585
R1680 gnd.n3012 gnd.n3011 585
R1681 gnd.n4697 gnd.n3012 585
R1682 gnd.n4711 gnd.n4710 585
R1683 gnd.n4710 gnd.n3036 585
R1684 gnd.n4712 gnd.n3048 585
R1685 gnd.n3048 gnd.n3035 585
R1686 gnd.n4714 gnd.n4713 585
R1687 gnd.n4715 gnd.n4714 585
R1688 gnd.n4709 gnd.n3047 585
R1689 gnd.n3047 gnd.n3043 585
R1690 gnd.n4708 gnd.n4707 585
R1691 gnd.n4707 gnd.n4706 585
R1692 gnd.n3050 gnd.n3049 585
R1693 gnd.n3056 gnd.n3050 585
R1694 gnd.n4689 gnd.n4688 585
R1695 gnd.n4690 gnd.n4689 585
R1696 gnd.n4687 gnd.n3059 585
R1697 gnd.n3064 gnd.n3059 585
R1698 gnd.n4686 gnd.n4685 585
R1699 gnd.n4685 gnd.n4684 585
R1700 gnd.n3061 gnd.n3060 585
R1701 gnd.n3074 gnd.n3061 585
R1702 gnd.n4671 gnd.n4670 585
R1703 gnd.n4672 gnd.n4671 585
R1704 gnd.n4669 gnd.n3075 585
R1705 gnd.n3075 gnd.n3071 585
R1706 gnd.n4668 gnd.n4667 585
R1707 gnd.n4667 gnd.n4666 585
R1708 gnd.n3077 gnd.n3076 585
R1709 gnd.n3078 gnd.n3077 585
R1710 gnd.n4623 gnd.n4622 585
R1711 gnd.n4623 gnd.n3087 585
R1712 gnd.n4625 gnd.n4624 585
R1713 gnd.n4624 gnd.n3086 585
R1714 gnd.n4626 gnd.n3100 585
R1715 gnd.n4611 gnd.n3100 585
R1716 gnd.n4628 gnd.n4627 585
R1717 gnd.n4629 gnd.n4628 585
R1718 gnd.n4621 gnd.n3099 585
R1719 gnd.n3099 gnd.n3095 585
R1720 gnd.n4620 gnd.n4619 585
R1721 gnd.n4619 gnd.n4618 585
R1722 gnd.n3102 gnd.n3101 585
R1723 gnd.n3108 gnd.n3102 585
R1724 gnd.n4593 gnd.n4592 585
R1725 gnd.n4594 gnd.n4593 585
R1726 gnd.n4591 gnd.n3110 585
R1727 gnd.n3117 gnd.n3110 585
R1728 gnd.n4590 gnd.n4589 585
R1729 gnd.n4589 gnd.n4588 585
R1730 gnd.n3112 gnd.n3111 585
R1731 gnd.n4463 gnd.n3112 585
R1732 gnd.n4575 gnd.n4574 585
R1733 gnd.n4576 gnd.n4575 585
R1734 gnd.n4573 gnd.n3127 585
R1735 gnd.n3127 gnd.n3124 585
R1736 gnd.n4572 gnd.n4571 585
R1737 gnd.n4571 gnd.n4570 585
R1738 gnd.n3129 gnd.n3128 585
R1739 gnd.n4460 gnd.n3129 585
R1740 gnd.n4530 gnd.n4529 585
R1741 gnd.n4530 gnd.n3139 585
R1742 gnd.n4532 gnd.n4531 585
R1743 gnd.n4531 gnd.n3138 585
R1744 gnd.n4533 gnd.n3151 585
R1745 gnd.n4475 gnd.n3151 585
R1746 gnd.n4535 gnd.n4534 585
R1747 gnd.n4536 gnd.n4535 585
R1748 gnd.n4528 gnd.n3150 585
R1749 gnd.n3150 gnd.n3147 585
R1750 gnd.n4527 gnd.n4526 585
R1751 gnd.n4526 gnd.n4525 585
R1752 gnd.n3153 gnd.n3152 585
R1753 gnd.n3154 gnd.n3153 585
R1754 gnd.n4498 gnd.n4497 585
R1755 gnd.n4498 gnd.n3163 585
R1756 gnd.n4500 gnd.n4499 585
R1757 gnd.n4499 gnd.n3162 585
R1758 gnd.n4501 gnd.n3177 585
R1759 gnd.n4486 gnd.n3177 585
R1760 gnd.n4503 gnd.n4502 585
R1761 gnd.n4504 gnd.n4503 585
R1762 gnd.n4496 gnd.n3176 585
R1763 gnd.n3176 gnd.n3172 585
R1764 gnd.n4495 gnd.n4494 585
R1765 gnd.n4494 gnd.n4493 585
R1766 gnd.n3179 gnd.n3178 585
R1767 gnd.n3187 gnd.n3179 585
R1768 gnd.n4452 gnd.n4451 585
R1769 gnd.n4453 gnd.n4452 585
R1770 gnd.n4450 gnd.n3189 585
R1771 gnd.n3189 gnd.n3186 585
R1772 gnd.n4449 gnd.n4448 585
R1773 gnd.n4448 gnd.n4447 585
R1774 gnd.n3191 gnd.n3190 585
R1775 gnd.n4319 gnd.n3191 585
R1776 gnd.n4433 gnd.n4432 585
R1777 gnd.n4434 gnd.n4433 585
R1778 gnd.n4431 gnd.n3204 585
R1779 gnd.n3204 gnd.n3201 585
R1780 gnd.n4430 gnd.n4429 585
R1781 gnd.n4429 gnd.n4428 585
R1782 gnd.n3206 gnd.n3205 585
R1783 gnd.n4316 gnd.n3206 585
R1784 gnd.n4388 gnd.n4387 585
R1785 gnd.n4388 gnd.n3215 585
R1786 gnd.n4390 gnd.n4389 585
R1787 gnd.n4389 gnd.n3214 585
R1788 gnd.n4391 gnd.n3226 585
R1789 gnd.n4332 gnd.n3226 585
R1790 gnd.n4393 gnd.n4392 585
R1791 gnd.n4394 gnd.n4393 585
R1792 gnd.n4386 gnd.n3225 585
R1793 gnd.n3225 gnd.n3222 585
R1794 gnd.n4385 gnd.n4384 585
R1795 gnd.n4384 gnd.n4383 585
R1796 gnd.n3228 gnd.n3227 585
R1797 gnd.n4312 gnd.n3228 585
R1798 gnd.n4356 gnd.n4355 585
R1799 gnd.n4356 gnd.n3237 585
R1800 gnd.n4358 gnd.n4357 585
R1801 gnd.n4357 gnd.n3236 585
R1802 gnd.n4359 gnd.n3249 585
R1803 gnd.n4344 gnd.n3249 585
R1804 gnd.n4361 gnd.n4360 585
R1805 gnd.n4362 gnd.n4361 585
R1806 gnd.n4354 gnd.n3248 585
R1807 gnd.n3248 gnd.n3245 585
R1808 gnd.n4353 gnd.n4352 585
R1809 gnd.n4352 gnd.n4351 585
R1810 gnd.n3251 gnd.n3250 585
R1811 gnd.n3258 gnd.n3251 585
R1812 gnd.n4305 gnd.n4304 585
R1813 gnd.n4306 gnd.n4305 585
R1814 gnd.n4303 gnd.n3261 585
R1815 gnd.n3261 gnd.n3257 585
R1816 gnd.n4302 gnd.n4301 585
R1817 gnd.n4301 gnd.n4300 585
R1818 gnd.n3263 gnd.n3262 585
R1819 gnd.n3275 gnd.n3263 585
R1820 gnd.n4287 gnd.n4286 585
R1821 gnd.n4288 gnd.n4287 585
R1822 gnd.n4285 gnd.n3276 585
R1823 gnd.n4279 gnd.n3276 585
R1824 gnd.n4284 gnd.n4283 585
R1825 gnd.n4283 gnd.n4282 585
R1826 gnd.n3278 gnd.n3277 585
R1827 gnd.n4269 gnd.n3278 585
R1828 gnd.n4255 gnd.n4254 585
R1829 gnd.n4254 gnd.n3283 585
R1830 gnd.n4256 gnd.n3294 585
R1831 gnd.n4221 gnd.n3294 585
R1832 gnd.n4258 gnd.n4257 585
R1833 gnd.n4259 gnd.n4258 585
R1834 gnd.n4253 gnd.n3293 585
R1835 gnd.n3293 gnd.n3290 585
R1836 gnd.n4252 gnd.n4251 585
R1837 gnd.n4251 gnd.n4250 585
R1838 gnd.n3296 gnd.n3295 585
R1839 gnd.n4212 gnd.n3296 585
R1840 gnd.n4210 gnd.n4209 585
R1841 gnd.n4211 gnd.n4210 585
R1842 gnd.n4208 gnd.n3307 585
R1843 gnd.n3313 gnd.n3307 585
R1844 gnd.n4207 gnd.n4206 585
R1845 gnd.n4206 gnd.n4205 585
R1846 gnd.n3309 gnd.n3308 585
R1847 gnd.n3310 gnd.n3309 585
R1848 gnd.n4189 gnd.n4188 585
R1849 gnd.n4190 gnd.n4189 585
R1850 gnd.n4187 gnd.n3325 585
R1851 gnd.n3325 gnd.n3320 585
R1852 gnd.n4186 gnd.n4185 585
R1853 gnd.n4185 gnd.n4184 585
R1854 gnd.n3327 gnd.n3326 585
R1855 gnd.n3333 gnd.n3327 585
R1856 gnd.n4170 gnd.n4169 585
R1857 gnd.n4171 gnd.n4170 585
R1858 gnd.n4168 gnd.n3339 585
R1859 gnd.n4163 gnd.n3339 585
R1860 gnd.n4167 gnd.n4166 585
R1861 gnd.n4166 gnd.n4165 585
R1862 gnd.n3341 gnd.n3340 585
R1863 gnd.n4137 gnd.n3341 585
R1864 gnd.n4139 gnd.n4138 585
R1865 gnd.n4140 gnd.n4139 585
R1866 gnd.n2604 gnd.n2603 585
R1867 gnd.n4061 gnd.n2604 585
R1868 gnd.n5552 gnd.n5551 585
R1869 gnd.n5551 gnd.n5550 585
R1870 gnd.n5553 gnd.n2582 585
R1871 gnd.n2605 gnd.n2582 585
R1872 gnd.n5618 gnd.n5617 585
R1873 gnd.n5616 gnd.n2581 585
R1874 gnd.n5615 gnd.n2580 585
R1875 gnd.n5620 gnd.n2580 585
R1876 gnd.n5614 gnd.n5613 585
R1877 gnd.n5612 gnd.n5611 585
R1878 gnd.n5610 gnd.n5609 585
R1879 gnd.n5608 gnd.n5607 585
R1880 gnd.n5606 gnd.n5605 585
R1881 gnd.n5604 gnd.n5603 585
R1882 gnd.n5602 gnd.n5601 585
R1883 gnd.n5600 gnd.n5599 585
R1884 gnd.n5598 gnd.n5597 585
R1885 gnd.n5596 gnd.n5595 585
R1886 gnd.n5594 gnd.n5593 585
R1887 gnd.n5592 gnd.n5591 585
R1888 gnd.n5590 gnd.n5589 585
R1889 gnd.n5588 gnd.n5587 585
R1890 gnd.n5586 gnd.n5585 585
R1891 gnd.n5584 gnd.n5583 585
R1892 gnd.n5582 gnd.n5581 585
R1893 gnd.n5580 gnd.n5579 585
R1894 gnd.n5578 gnd.n5577 585
R1895 gnd.n5576 gnd.n5575 585
R1896 gnd.n5574 gnd.n5573 585
R1897 gnd.n5572 gnd.n5571 585
R1898 gnd.n5570 gnd.n5569 585
R1899 gnd.n5568 gnd.n5567 585
R1900 gnd.n5566 gnd.n5565 585
R1901 gnd.n5564 gnd.n5563 585
R1902 gnd.n5562 gnd.n5561 585
R1903 gnd.n5560 gnd.n5559 585
R1904 gnd.n5558 gnd.n2545 585
R1905 gnd.n5623 gnd.n5622 585
R1906 gnd.n2547 gnd.n2544 585
R1907 gnd.n4066 gnd.n4065 585
R1908 gnd.n4068 gnd.n4067 585
R1909 gnd.n4071 gnd.n4070 585
R1910 gnd.n4073 gnd.n4072 585
R1911 gnd.n4075 gnd.n4074 585
R1912 gnd.n4077 gnd.n4076 585
R1913 gnd.n4079 gnd.n4078 585
R1914 gnd.n4081 gnd.n4080 585
R1915 gnd.n4083 gnd.n4082 585
R1916 gnd.n4085 gnd.n4084 585
R1917 gnd.n4087 gnd.n4086 585
R1918 gnd.n4089 gnd.n4088 585
R1919 gnd.n4091 gnd.n4090 585
R1920 gnd.n4093 gnd.n4092 585
R1921 gnd.n4095 gnd.n4094 585
R1922 gnd.n4097 gnd.n4096 585
R1923 gnd.n4099 gnd.n4098 585
R1924 gnd.n4101 gnd.n4100 585
R1925 gnd.n4103 gnd.n4102 585
R1926 gnd.n4105 gnd.n4104 585
R1927 gnd.n4107 gnd.n4106 585
R1928 gnd.n4109 gnd.n4108 585
R1929 gnd.n4111 gnd.n4110 585
R1930 gnd.n4113 gnd.n4112 585
R1931 gnd.n4115 gnd.n4114 585
R1932 gnd.n4117 gnd.n4116 585
R1933 gnd.n4119 gnd.n4118 585
R1934 gnd.n4121 gnd.n4120 585
R1935 gnd.n4123 gnd.n4122 585
R1936 gnd.n4125 gnd.n4124 585
R1937 gnd.n4127 gnd.n4126 585
R1938 gnd.n4913 gnd.n4912 585
R1939 gnd.n4915 gnd.n4914 585
R1940 gnd.n4917 gnd.n4916 585
R1941 gnd.n4919 gnd.n4918 585
R1942 gnd.n4921 gnd.n4920 585
R1943 gnd.n4923 gnd.n4922 585
R1944 gnd.n4925 gnd.n4924 585
R1945 gnd.n4927 gnd.n4926 585
R1946 gnd.n4929 gnd.n4928 585
R1947 gnd.n4931 gnd.n4930 585
R1948 gnd.n4933 gnd.n4932 585
R1949 gnd.n4935 gnd.n4934 585
R1950 gnd.n4937 gnd.n4936 585
R1951 gnd.n4939 gnd.n4938 585
R1952 gnd.n4941 gnd.n4940 585
R1953 gnd.n4943 gnd.n4942 585
R1954 gnd.n4945 gnd.n4944 585
R1955 gnd.n4947 gnd.n4946 585
R1956 gnd.n4949 gnd.n4948 585
R1957 gnd.n4951 gnd.n4950 585
R1958 gnd.n4953 gnd.n4952 585
R1959 gnd.n4955 gnd.n4954 585
R1960 gnd.n4957 gnd.n4956 585
R1961 gnd.n4959 gnd.n4958 585
R1962 gnd.n4961 gnd.n4960 585
R1963 gnd.n4963 gnd.n4962 585
R1964 gnd.n4965 gnd.n4964 585
R1965 gnd.n4967 gnd.n4966 585
R1966 gnd.n4969 gnd.n4968 585
R1967 gnd.n4972 gnd.n4971 585
R1968 gnd.n4974 gnd.n4973 585
R1969 gnd.n4976 gnd.n4975 585
R1970 gnd.n4978 gnd.n4977 585
R1971 gnd.n4842 gnd.n2836 585
R1972 gnd.n4844 gnd.n4843 585
R1973 gnd.n4846 gnd.n4845 585
R1974 gnd.n4848 gnd.n4847 585
R1975 gnd.n4851 gnd.n4850 585
R1976 gnd.n4853 gnd.n4852 585
R1977 gnd.n4855 gnd.n4854 585
R1978 gnd.n4857 gnd.n4856 585
R1979 gnd.n4859 gnd.n4858 585
R1980 gnd.n4861 gnd.n4860 585
R1981 gnd.n4863 gnd.n4862 585
R1982 gnd.n4865 gnd.n4864 585
R1983 gnd.n4867 gnd.n4866 585
R1984 gnd.n4869 gnd.n4868 585
R1985 gnd.n4871 gnd.n4870 585
R1986 gnd.n4873 gnd.n4872 585
R1987 gnd.n4875 gnd.n4874 585
R1988 gnd.n4877 gnd.n4876 585
R1989 gnd.n4879 gnd.n4878 585
R1990 gnd.n4881 gnd.n4880 585
R1991 gnd.n4883 gnd.n4882 585
R1992 gnd.n4885 gnd.n4884 585
R1993 gnd.n4887 gnd.n4886 585
R1994 gnd.n4889 gnd.n4888 585
R1995 gnd.n4891 gnd.n4890 585
R1996 gnd.n4893 gnd.n4892 585
R1997 gnd.n4895 gnd.n4894 585
R1998 gnd.n4897 gnd.n4896 585
R1999 gnd.n4899 gnd.n4898 585
R2000 gnd.n4901 gnd.n4900 585
R2001 gnd.n4903 gnd.n4902 585
R2002 gnd.n4905 gnd.n4904 585
R2003 gnd.n4906 gnd.n2978 585
R2004 gnd.n4911 gnd.n2975 585
R2005 gnd.n4911 gnd.n4910 585
R2006 gnd.n4791 gnd.n2976 585
R2007 gnd.n2983 gnd.n2976 585
R2008 gnd.n4792 gnd.n2981 585
R2009 gnd.n4817 gnd.n2981 585
R2010 gnd.n4794 gnd.n4793 585
R2011 gnd.n4793 gnd.n2991 585
R2012 gnd.n4795 gnd.n2990 585
R2013 gnd.n4806 gnd.n2990 585
R2014 gnd.n4797 gnd.n4796 585
R2015 gnd.n4798 gnd.n4797 585
R2016 gnd.n4790 gnd.n2996 585
R2017 gnd.n4800 gnd.n2996 585
R2018 gnd.n4789 gnd.n4788 585
R2019 gnd.n4788 gnd.n2995 585
R2020 gnd.n4787 gnd.n2998 585
R2021 gnd.n4787 gnd.n4786 585
R2022 gnd.n4776 gnd.n2999 585
R2023 gnd.n4779 gnd.n2999 585
R2024 gnd.n4778 gnd.n4777 585
R2025 gnd.n4780 gnd.n4778 585
R2026 gnd.n4775 gnd.n3006 585
R2027 gnd.n4733 gnd.n3006 585
R2028 gnd.n4774 gnd.n4773 585
R2029 gnd.n4773 gnd.n4772 585
R2030 gnd.n3008 gnd.n3007 585
R2031 gnd.n3009 gnd.n3008 585
R2032 gnd.n4695 gnd.n3014 585
R2033 gnd.n4766 gnd.n3014 585
R2034 gnd.n4698 gnd.n4696 585
R2035 gnd.n4698 gnd.n4697 585
R2036 gnd.n4699 gnd.n4694 585
R2037 gnd.n4699 gnd.n3036 585
R2038 gnd.n4701 gnd.n4700 585
R2039 gnd.n4700 gnd.n3035 585
R2040 gnd.n4702 gnd.n3045 585
R2041 gnd.n4715 gnd.n3045 585
R2042 gnd.n4703 gnd.n3053 585
R2043 gnd.n3053 gnd.n3043 585
R2044 gnd.n4705 gnd.n4704 585
R2045 gnd.n4706 gnd.n4705 585
R2046 gnd.n4693 gnd.n3052 585
R2047 gnd.n3056 gnd.n3052 585
R2048 gnd.n4692 gnd.n4691 585
R2049 gnd.n4691 gnd.n4690 585
R2050 gnd.n3055 gnd.n3054 585
R2051 gnd.n3064 gnd.n3055 585
R2052 gnd.n4600 gnd.n3062 585
R2053 gnd.n4684 gnd.n3062 585
R2054 gnd.n4602 gnd.n4601 585
R2055 gnd.n4601 gnd.n3074 585
R2056 gnd.n4603 gnd.n3073 585
R2057 gnd.n4672 gnd.n3073 585
R2058 gnd.n4605 gnd.n4604 585
R2059 gnd.n4604 gnd.n3071 585
R2060 gnd.n4606 gnd.n3079 585
R2061 gnd.n4666 gnd.n3079 585
R2062 gnd.n4607 gnd.n4599 585
R2063 gnd.n4599 gnd.n3078 585
R2064 gnd.n4609 gnd.n4608 585
R2065 gnd.n4609 gnd.n3087 585
R2066 gnd.n4610 gnd.n4598 585
R2067 gnd.n4610 gnd.n3086 585
R2068 gnd.n4613 gnd.n4612 585
R2069 gnd.n4612 gnd.n4611 585
R2070 gnd.n4614 gnd.n3097 585
R2071 gnd.n4629 gnd.n3097 585
R2072 gnd.n4615 gnd.n3105 585
R2073 gnd.n3105 gnd.n3095 585
R2074 gnd.n4617 gnd.n4616 585
R2075 gnd.n4618 gnd.n4617 585
R2076 gnd.n4597 gnd.n3104 585
R2077 gnd.n3108 gnd.n3104 585
R2078 gnd.n4596 gnd.n4595 585
R2079 gnd.n4595 gnd.n4594 585
R2080 gnd.n3107 gnd.n3106 585
R2081 gnd.n3117 gnd.n3107 585
R2082 gnd.n4462 gnd.n3115 585
R2083 gnd.n4588 gnd.n3115 585
R2084 gnd.n4465 gnd.n4464 585
R2085 gnd.n4464 gnd.n4463 585
R2086 gnd.n4466 gnd.n3126 585
R2087 gnd.n4576 gnd.n3126 585
R2088 gnd.n4468 gnd.n4467 585
R2089 gnd.n4467 gnd.n3124 585
R2090 gnd.n4469 gnd.n3131 585
R2091 gnd.n4570 gnd.n3131 585
R2092 gnd.n4470 gnd.n4461 585
R2093 gnd.n4461 gnd.n4460 585
R2094 gnd.n4472 gnd.n4471 585
R2095 gnd.n4472 gnd.n3139 585
R2096 gnd.n4473 gnd.n4459 585
R2097 gnd.n4473 gnd.n3138 585
R2098 gnd.n4477 gnd.n4476 585
R2099 gnd.n4476 gnd.n4475 585
R2100 gnd.n4478 gnd.n3149 585
R2101 gnd.n4536 gnd.n3149 585
R2102 gnd.n4480 gnd.n4479 585
R2103 gnd.n4479 gnd.n3147 585
R2104 gnd.n4481 gnd.n3155 585
R2105 gnd.n4525 gnd.n3155 585
R2106 gnd.n4482 gnd.n4458 585
R2107 gnd.n4458 gnd.n3154 585
R2108 gnd.n4484 gnd.n4483 585
R2109 gnd.n4484 gnd.n3163 585
R2110 gnd.n4485 gnd.n4457 585
R2111 gnd.n4485 gnd.n3162 585
R2112 gnd.n4488 gnd.n4487 585
R2113 gnd.n4487 gnd.n4486 585
R2114 gnd.n4489 gnd.n3174 585
R2115 gnd.n4504 gnd.n3174 585
R2116 gnd.n4490 gnd.n3183 585
R2117 gnd.n3183 gnd.n3172 585
R2118 gnd.n4492 gnd.n4491 585
R2119 gnd.n4493 gnd.n4492 585
R2120 gnd.n4456 gnd.n3182 585
R2121 gnd.n3187 gnd.n3182 585
R2122 gnd.n4455 gnd.n4454 585
R2123 gnd.n4454 gnd.n4453 585
R2124 gnd.n3185 gnd.n3184 585
R2125 gnd.n3186 gnd.n3185 585
R2126 gnd.n4318 gnd.n3193 585
R2127 gnd.n4447 gnd.n3193 585
R2128 gnd.n4321 gnd.n4320 585
R2129 gnd.n4320 gnd.n4319 585
R2130 gnd.n4322 gnd.n3203 585
R2131 gnd.n4434 gnd.n3203 585
R2132 gnd.n4324 gnd.n4323 585
R2133 gnd.n4323 gnd.n3201 585
R2134 gnd.n4325 gnd.n3207 585
R2135 gnd.n4428 gnd.n3207 585
R2136 gnd.n4326 gnd.n4317 585
R2137 gnd.n4317 gnd.n4316 585
R2138 gnd.n4328 gnd.n4327 585
R2139 gnd.n4328 gnd.n3215 585
R2140 gnd.n4329 gnd.n4314 585
R2141 gnd.n4329 gnd.n3214 585
R2142 gnd.n4334 gnd.n4333 585
R2143 gnd.n4333 gnd.n4332 585
R2144 gnd.n4335 gnd.n3224 585
R2145 gnd.n4394 gnd.n3224 585
R2146 gnd.n4337 gnd.n4336 585
R2147 gnd.n4336 gnd.n3222 585
R2148 gnd.n4338 gnd.n3229 585
R2149 gnd.n4383 gnd.n3229 585
R2150 gnd.n4339 gnd.n4313 585
R2151 gnd.n4313 gnd.n4312 585
R2152 gnd.n4341 gnd.n4340 585
R2153 gnd.n4341 gnd.n3237 585
R2154 gnd.n4342 gnd.n4310 585
R2155 gnd.n4342 gnd.n3236 585
R2156 gnd.n4346 gnd.n4345 585
R2157 gnd.n4345 gnd.n4344 585
R2158 gnd.n4347 gnd.n3247 585
R2159 gnd.n4362 gnd.n3247 585
R2160 gnd.n4348 gnd.n3254 585
R2161 gnd.n3254 gnd.n3245 585
R2162 gnd.n4350 gnd.n4349 585
R2163 gnd.n4351 gnd.n4350 585
R2164 gnd.n4309 gnd.n3253 585
R2165 gnd.n3258 gnd.n3253 585
R2166 gnd.n4308 gnd.n4307 585
R2167 gnd.n4307 gnd.n4306 585
R2168 gnd.n3256 gnd.n3255 585
R2169 gnd.n3257 gnd.n3256 585
R2170 gnd.n4273 gnd.n3265 585
R2171 gnd.n4300 gnd.n3265 585
R2172 gnd.n4275 gnd.n4274 585
R2173 gnd.n4274 gnd.n3275 585
R2174 gnd.n4276 gnd.n3274 585
R2175 gnd.n4288 gnd.n3274 585
R2176 gnd.n4278 gnd.n4277 585
R2177 gnd.n4279 gnd.n4278 585
R2178 gnd.n4272 gnd.n3279 585
R2179 gnd.n4282 gnd.n3279 585
R2180 gnd.n4271 gnd.n4270 585
R2181 gnd.n4270 gnd.n4269 585
R2182 gnd.n3282 gnd.n3281 585
R2183 gnd.n3283 gnd.n3282 585
R2184 gnd.n4220 gnd.n4219 585
R2185 gnd.n4221 gnd.n4220 585
R2186 gnd.n4218 gnd.n3292 585
R2187 gnd.n4259 gnd.n3292 585
R2188 gnd.n4217 gnd.n4216 585
R2189 gnd.n4216 gnd.n3290 585
R2190 gnd.n4215 gnd.n3298 585
R2191 gnd.n4250 gnd.n3298 585
R2192 gnd.n4214 gnd.n4213 585
R2193 gnd.n4213 gnd.n4212 585
R2194 gnd.n3305 gnd.n3304 585
R2195 gnd.n4211 gnd.n3305 585
R2196 gnd.n4176 gnd.n4175 585
R2197 gnd.n4175 gnd.n3313 585
R2198 gnd.n4177 gnd.n3311 585
R2199 gnd.n4205 gnd.n3311 585
R2200 gnd.n4179 gnd.n4178 585
R2201 gnd.n4178 gnd.n3310 585
R2202 gnd.n4180 gnd.n3322 585
R2203 gnd.n4190 gnd.n3322 585
R2204 gnd.n4181 gnd.n3330 585
R2205 gnd.n3330 gnd.n3320 585
R2206 gnd.n4183 gnd.n4182 585
R2207 gnd.n4184 gnd.n4183 585
R2208 gnd.n4174 gnd.n3329 585
R2209 gnd.n3333 gnd.n3329 585
R2210 gnd.n4173 gnd.n4172 585
R2211 gnd.n4172 gnd.n4171 585
R2212 gnd.n3332 gnd.n3331 585
R2213 gnd.n4163 gnd.n3332 585
R2214 gnd.n4134 gnd.n3342 585
R2215 gnd.n4165 gnd.n3342 585
R2216 gnd.n4136 gnd.n4135 585
R2217 gnd.n4137 gnd.n4136 585
R2218 gnd.n4133 gnd.n4062 585
R2219 gnd.n4140 gnd.n4062 585
R2220 gnd.n4132 gnd.n4131 585
R2221 gnd.n4131 gnd.n4061 585
R2222 gnd.n4130 gnd.n2606 585
R2223 gnd.n5550 gnd.n2606 585
R2224 gnd.n4129 gnd.n4128 585
R2225 gnd.n4128 gnd.n2605 585
R2226 gnd.n5679 gnd.n2468 585
R2227 gnd.n3924 gnd.n2468 585
R2228 gnd.n5681 gnd.n5680 585
R2229 gnd.n5682 gnd.n5681 585
R2230 gnd.n2453 gnd.n2452 585
R2231 gnd.n3863 gnd.n2453 585
R2232 gnd.n5690 gnd.n5689 585
R2233 gnd.n5689 gnd.n5688 585
R2234 gnd.n5691 gnd.n2447 585
R2235 gnd.n3854 gnd.n2447 585
R2236 gnd.n5693 gnd.n5692 585
R2237 gnd.n5694 gnd.n5693 585
R2238 gnd.n2432 gnd.n2431 585
R2239 gnd.n3849 gnd.n2432 585
R2240 gnd.n5702 gnd.n5701 585
R2241 gnd.n5701 gnd.n5700 585
R2242 gnd.n5703 gnd.n2426 585
R2243 gnd.n3845 gnd.n2426 585
R2244 gnd.n5705 gnd.n5704 585
R2245 gnd.n5706 gnd.n5705 585
R2246 gnd.n2412 gnd.n2411 585
R2247 gnd.n3883 gnd.n2412 585
R2248 gnd.n5714 gnd.n5713 585
R2249 gnd.n5713 gnd.n5712 585
R2250 gnd.n5715 gnd.n2406 585
R2251 gnd.n3838 gnd.n2406 585
R2252 gnd.n5717 gnd.n5716 585
R2253 gnd.n5718 gnd.n5717 585
R2254 gnd.n2392 gnd.n2391 585
R2255 gnd.n3830 gnd.n2392 585
R2256 gnd.n5726 gnd.n5725 585
R2257 gnd.n5725 gnd.n5724 585
R2258 gnd.n5727 gnd.n2386 585
R2259 gnd.n2386 gnd.n2385 585
R2260 gnd.n5729 gnd.n5728 585
R2261 gnd.n5730 gnd.n5729 585
R2262 gnd.n2373 gnd.n2372 585
R2263 gnd.n2376 gnd.n2373 585
R2264 gnd.n5738 gnd.n5737 585
R2265 gnd.n5737 gnd.n5736 585
R2266 gnd.n5739 gnd.n2367 585
R2267 gnd.n2367 gnd.n2366 585
R2268 gnd.n5741 gnd.n5740 585
R2269 gnd.n5742 gnd.n5741 585
R2270 gnd.n2353 gnd.n2352 585
R2271 gnd.n2363 gnd.n2353 585
R2272 gnd.n5750 gnd.n5749 585
R2273 gnd.n5749 gnd.n5748 585
R2274 gnd.n5751 gnd.n2347 585
R2275 gnd.n2354 gnd.n2347 585
R2276 gnd.n5753 gnd.n5752 585
R2277 gnd.n5754 gnd.n5753 585
R2278 gnd.n2335 gnd.n2334 585
R2279 gnd.n2338 gnd.n2335 585
R2280 gnd.n5762 gnd.n5761 585
R2281 gnd.n5761 gnd.n5760 585
R2282 gnd.n5763 gnd.n2329 585
R2283 gnd.n2329 gnd.n2328 585
R2284 gnd.n5765 gnd.n5764 585
R2285 gnd.n5766 gnd.n5765 585
R2286 gnd.n2315 gnd.n2314 585
R2287 gnd.n2325 gnd.n2315 585
R2288 gnd.n5774 gnd.n5773 585
R2289 gnd.n5773 gnd.n5772 585
R2290 gnd.n5775 gnd.n2309 585
R2291 gnd.n2316 gnd.n2309 585
R2292 gnd.n5777 gnd.n5776 585
R2293 gnd.n5778 gnd.n5777 585
R2294 gnd.n2297 gnd.n2296 585
R2295 gnd.n2300 gnd.n2297 585
R2296 gnd.n5786 gnd.n5785 585
R2297 gnd.n5785 gnd.n5784 585
R2298 gnd.n5787 gnd.n2292 585
R2299 gnd.n2292 gnd.n2291 585
R2300 gnd.n5789 gnd.n5788 585
R2301 gnd.n5790 gnd.n5789 585
R2302 gnd.n2277 gnd.n2276 585
R2303 gnd.n2281 gnd.n2277 585
R2304 gnd.n5798 gnd.n5797 585
R2305 gnd.n5797 gnd.n5796 585
R2306 gnd.n2273 gnd.n2271 585
R2307 gnd.n2278 gnd.n2271 585
R2308 gnd.n5803 gnd.n5802 585
R2309 gnd.n5804 gnd.n5803 585
R2310 gnd.n2272 gnd.n2196 585
R2311 gnd.n2196 gnd.n2193 585
R2312 gnd.n5926 gnd.n5925 585
R2313 gnd.n5924 gnd.n2195 585
R2314 gnd.n5923 gnd.n2194 585
R2315 gnd.n5928 gnd.n2194 585
R2316 gnd.n5922 gnd.n5921 585
R2317 gnd.n5920 gnd.n5919 585
R2318 gnd.n5918 gnd.n5917 585
R2319 gnd.n5916 gnd.n5915 585
R2320 gnd.n5914 gnd.n5913 585
R2321 gnd.n5912 gnd.n5911 585
R2322 gnd.n5910 gnd.n5909 585
R2323 gnd.n5908 gnd.n5907 585
R2324 gnd.n5906 gnd.n5905 585
R2325 gnd.n5904 gnd.n5903 585
R2326 gnd.n5902 gnd.n5901 585
R2327 gnd.n5900 gnd.n5899 585
R2328 gnd.n5898 gnd.n5897 585
R2329 gnd.n5896 gnd.n5895 585
R2330 gnd.n5894 gnd.n5893 585
R2331 gnd.n5891 gnd.n5890 585
R2332 gnd.n5889 gnd.n5888 585
R2333 gnd.n5887 gnd.n5886 585
R2334 gnd.n5885 gnd.n5884 585
R2335 gnd.n5883 gnd.n5882 585
R2336 gnd.n5881 gnd.n5880 585
R2337 gnd.n5879 gnd.n5878 585
R2338 gnd.n5877 gnd.n5876 585
R2339 gnd.n5875 gnd.n5874 585
R2340 gnd.n5873 gnd.n5872 585
R2341 gnd.n5871 gnd.n5870 585
R2342 gnd.n5869 gnd.n5868 585
R2343 gnd.n5867 gnd.n5866 585
R2344 gnd.n5865 gnd.n5864 585
R2345 gnd.n5863 gnd.n5862 585
R2346 gnd.n5861 gnd.n5860 585
R2347 gnd.n5859 gnd.n5858 585
R2348 gnd.n5857 gnd.n5856 585
R2349 gnd.n5855 gnd.n5854 585
R2350 gnd.n5853 gnd.n5852 585
R2351 gnd.n5851 gnd.n5850 585
R2352 gnd.n5849 gnd.n5848 585
R2353 gnd.n5847 gnd.n5846 585
R2354 gnd.n5845 gnd.n5844 585
R2355 gnd.n5843 gnd.n5842 585
R2356 gnd.n5841 gnd.n5840 585
R2357 gnd.n5839 gnd.n5838 585
R2358 gnd.n5837 gnd.n5836 585
R2359 gnd.n5835 gnd.n5834 585
R2360 gnd.n5833 gnd.n5832 585
R2361 gnd.n5831 gnd.n5830 585
R2362 gnd.n5829 gnd.n5828 585
R2363 gnd.n5827 gnd.n5826 585
R2364 gnd.n5825 gnd.n5824 585
R2365 gnd.n5823 gnd.n5822 585
R2366 gnd.n5821 gnd.n5820 585
R2367 gnd.n5819 gnd.n5818 585
R2368 gnd.n5817 gnd.n5816 585
R2369 gnd.n5815 gnd.n5814 585
R2370 gnd.n5813 gnd.n5812 585
R2371 gnd.n2267 gnd.n2258 585
R2372 gnd.n3616 gnd.n3615 585
R2373 gnd.n3609 gnd.n3523 585
R2374 gnd.n3611 gnd.n3610 585
R2375 gnd.n3608 gnd.n3607 585
R2376 gnd.n3606 gnd.n3605 585
R2377 gnd.n3599 gnd.n3525 585
R2378 gnd.n3601 gnd.n3600 585
R2379 gnd.n3598 gnd.n3597 585
R2380 gnd.n3596 gnd.n3595 585
R2381 gnd.n3589 gnd.n3527 585
R2382 gnd.n3591 gnd.n3590 585
R2383 gnd.n3588 gnd.n3587 585
R2384 gnd.n3586 gnd.n3585 585
R2385 gnd.n3579 gnd.n3529 585
R2386 gnd.n3581 gnd.n3580 585
R2387 gnd.n3578 gnd.n3577 585
R2388 gnd.n3576 gnd.n3575 585
R2389 gnd.n3569 gnd.n3531 585
R2390 gnd.n3571 gnd.n3570 585
R2391 gnd.n3568 gnd.n3567 585
R2392 gnd.n3566 gnd.n3565 585
R2393 gnd.n3559 gnd.n3535 585
R2394 gnd.n3561 gnd.n3560 585
R2395 gnd.n3558 gnd.n3557 585
R2396 gnd.n3556 gnd.n3555 585
R2397 gnd.n3549 gnd.n3537 585
R2398 gnd.n3551 gnd.n3550 585
R2399 gnd.n3548 gnd.n3547 585
R2400 gnd.n3546 gnd.n3545 585
R2401 gnd.n3541 gnd.n3540 585
R2402 gnd.n3539 gnd.n2541 585
R2403 gnd.n5626 gnd.n5625 585
R2404 gnd.n5628 gnd.n5627 585
R2405 gnd.n5630 gnd.n5629 585
R2406 gnd.n5632 gnd.n5631 585
R2407 gnd.n5634 gnd.n5633 585
R2408 gnd.n5636 gnd.n5635 585
R2409 gnd.n5638 gnd.n5637 585
R2410 gnd.n5640 gnd.n5639 585
R2411 gnd.n5643 gnd.n5642 585
R2412 gnd.n5645 gnd.n5644 585
R2413 gnd.n5647 gnd.n5646 585
R2414 gnd.n5649 gnd.n5648 585
R2415 gnd.n5651 gnd.n5650 585
R2416 gnd.n5653 gnd.n5652 585
R2417 gnd.n5655 gnd.n5654 585
R2418 gnd.n5657 gnd.n5656 585
R2419 gnd.n5659 gnd.n5658 585
R2420 gnd.n5661 gnd.n5660 585
R2421 gnd.n5663 gnd.n5662 585
R2422 gnd.n5665 gnd.n5664 585
R2423 gnd.n5667 gnd.n5666 585
R2424 gnd.n5669 gnd.n5668 585
R2425 gnd.n5670 gnd.n2514 585
R2426 gnd.n5672 gnd.n5671 585
R2427 gnd.n2473 gnd.n2472 585
R2428 gnd.n5676 gnd.n5675 585
R2429 gnd.n5675 gnd.n5674 585
R2430 gnd.n3859 gnd.n3617 585
R2431 gnd.n3924 gnd.n3617 585
R2432 gnd.n3860 gnd.n2465 585
R2433 gnd.n5682 gnd.n2465 585
R2434 gnd.n3862 gnd.n3861 585
R2435 gnd.n3863 gnd.n3862 585
R2436 gnd.n3857 gnd.n2455 585
R2437 gnd.n5688 gnd.n2455 585
R2438 gnd.n3856 gnd.n3855 585
R2439 gnd.n3855 gnd.n3854 585
R2440 gnd.n3852 gnd.n2444 585
R2441 gnd.n5694 gnd.n2444 585
R2442 gnd.n3851 gnd.n3850 585
R2443 gnd.n3850 gnd.n3849 585
R2444 gnd.n3848 gnd.n2434 585
R2445 gnd.n5700 gnd.n2434 585
R2446 gnd.n3847 gnd.n3846 585
R2447 gnd.n3846 gnd.n3845 585
R2448 gnd.n3843 gnd.n2423 585
R2449 gnd.n5706 gnd.n2423 585
R2450 gnd.n3842 gnd.n3642 585
R2451 gnd.n3883 gnd.n3642 585
R2452 gnd.n3841 gnd.n2414 585
R2453 gnd.n5712 gnd.n2414 585
R2454 gnd.n3840 gnd.n3839 585
R2455 gnd.n3839 gnd.n3838 585
R2456 gnd.n3652 gnd.n2403 585
R2457 gnd.n5718 gnd.n2403 585
R2458 gnd.n3829 gnd.n3828 585
R2459 gnd.n3830 gnd.n3829 585
R2460 gnd.n3827 gnd.n2394 585
R2461 gnd.n5724 gnd.n2394 585
R2462 gnd.n3826 gnd.n3825 585
R2463 gnd.n3825 gnd.n2385 585
R2464 gnd.n3823 gnd.n2383 585
R2465 gnd.n5730 gnd.n2383 585
R2466 gnd.n3822 gnd.n3821 585
R2467 gnd.n3821 gnd.n2376 585
R2468 gnd.n3820 gnd.n2374 585
R2469 gnd.n5736 gnd.n2374 585
R2470 gnd.n3819 gnd.n3818 585
R2471 gnd.n3818 gnd.n2366 585
R2472 gnd.n3816 gnd.n2364 585
R2473 gnd.n5742 gnd.n2364 585
R2474 gnd.n3815 gnd.n3814 585
R2475 gnd.n3814 gnd.n2363 585
R2476 gnd.n3813 gnd.n2355 585
R2477 gnd.n5748 gnd.n2355 585
R2478 gnd.n3812 gnd.n3811 585
R2479 gnd.n3811 gnd.n2354 585
R2480 gnd.n3809 gnd.n2345 585
R2481 gnd.n5754 gnd.n2345 585
R2482 gnd.n3808 gnd.n3807 585
R2483 gnd.n3807 gnd.n2338 585
R2484 gnd.n3806 gnd.n2336 585
R2485 gnd.n5760 gnd.n2336 585
R2486 gnd.n3805 gnd.n3804 585
R2487 gnd.n3804 gnd.n2328 585
R2488 gnd.n3802 gnd.n2326 585
R2489 gnd.n5766 gnd.n2326 585
R2490 gnd.n3801 gnd.n3800 585
R2491 gnd.n3800 gnd.n2325 585
R2492 gnd.n3799 gnd.n2317 585
R2493 gnd.n5772 gnd.n2317 585
R2494 gnd.n3798 gnd.n3797 585
R2495 gnd.n3797 gnd.n2316 585
R2496 gnd.n3795 gnd.n2307 585
R2497 gnd.n5778 gnd.n2307 585
R2498 gnd.n3794 gnd.n3793 585
R2499 gnd.n3793 gnd.n2300 585
R2500 gnd.n3792 gnd.n2298 585
R2501 gnd.n5784 gnd.n2298 585
R2502 gnd.n3791 gnd.n3790 585
R2503 gnd.n3790 gnd.n2291 585
R2504 gnd.n3788 gnd.n2289 585
R2505 gnd.n5790 gnd.n2289 585
R2506 gnd.n3787 gnd.n3786 585
R2507 gnd.n3786 gnd.n2281 585
R2508 gnd.n3785 gnd.n2279 585
R2509 gnd.n5796 gnd.n2279 585
R2510 gnd.n3784 gnd.n3783 585
R2511 gnd.n3783 gnd.n2278 585
R2512 gnd.n3781 gnd.n2269 585
R2513 gnd.n5804 gnd.n2269 585
R2514 gnd.n2268 gnd.n2262 585
R2515 gnd.n2268 gnd.n2193 585
R2516 gnd.n162 gnd.n161 585
R2517 gnd.n165 gnd.n162 585
R2518 gnd.n7212 gnd.n7211 585
R2519 gnd.n7211 gnd.n7210 585
R2520 gnd.n7213 gnd.n156 585
R2521 gnd.n156 gnd.n155 585
R2522 gnd.n7215 gnd.n7214 585
R2523 gnd.n7216 gnd.n7215 585
R2524 gnd.n142 gnd.n141 585
R2525 gnd.n146 gnd.n142 585
R2526 gnd.n7224 gnd.n7223 585
R2527 gnd.n7223 gnd.n7222 585
R2528 gnd.n7225 gnd.n136 585
R2529 gnd.n143 gnd.n136 585
R2530 gnd.n7227 gnd.n7226 585
R2531 gnd.n7228 gnd.n7227 585
R2532 gnd.n123 gnd.n122 585
R2533 gnd.n126 gnd.n123 585
R2534 gnd.n7236 gnd.n7235 585
R2535 gnd.n7235 gnd.n7234 585
R2536 gnd.n7237 gnd.n117 585
R2537 gnd.n117 gnd.n116 585
R2538 gnd.n7239 gnd.n7238 585
R2539 gnd.n7240 gnd.n7239 585
R2540 gnd.n103 gnd.n102 585
R2541 gnd.n107 gnd.n103 585
R2542 gnd.n7248 gnd.n7247 585
R2543 gnd.n7247 gnd.n7246 585
R2544 gnd.n7249 gnd.n97 585
R2545 gnd.n104 gnd.n97 585
R2546 gnd.n7251 gnd.n7250 585
R2547 gnd.n7252 gnd.n7251 585
R2548 gnd.n83 gnd.n82 585
R2549 gnd.n86 gnd.n83 585
R2550 gnd.n7260 gnd.n7259 585
R2551 gnd.n7259 gnd.n7258 585
R2552 gnd.n7261 gnd.n77 585
R2553 gnd.n77 gnd.n74 585
R2554 gnd.n7263 gnd.n7262 585
R2555 gnd.n7264 gnd.n7263 585
R2556 gnd.n78 gnd.n76 585
R2557 gnd.n6837 gnd.n76 585
R2558 gnd.n6826 gnd.n182 585
R2559 gnd.n182 gnd.n172 585
R2560 gnd.n6828 gnd.n6827 585
R2561 gnd.n6829 gnd.n6828 585
R2562 gnd.n183 gnd.n181 585
R2563 gnd.n189 gnd.n181 585
R2564 gnd.n6820 gnd.n6819 585
R2565 gnd.n6819 gnd.n6818 585
R2566 gnd.n186 gnd.n185 585
R2567 gnd.n6809 gnd.n186 585
R2568 gnd.n6793 gnd.n206 585
R2569 gnd.n206 gnd.n195 585
R2570 gnd.n6795 gnd.n6794 585
R2571 gnd.n6796 gnd.n6795 585
R2572 gnd.n207 gnd.n205 585
R2573 gnd.n6774 gnd.n205 585
R2574 gnd.n6788 gnd.n6787 585
R2575 gnd.n6787 gnd.n6786 585
R2576 gnd.n210 gnd.n209 585
R2577 gnd.n6770 gnd.n210 585
R2578 gnd.n6758 gnd.n234 585
R2579 gnd.n6744 gnd.n234 585
R2580 gnd.n6760 gnd.n6759 585
R2581 gnd.n6761 gnd.n6760 585
R2582 gnd.n235 gnd.n233 585
R2583 gnd.n5102 gnd.n233 585
R2584 gnd.n6753 gnd.n6752 585
R2585 gnd.n6752 gnd.n6751 585
R2586 gnd.n238 gnd.n237 585
R2587 gnd.n5170 gnd.n238 585
R2588 gnd.n5091 gnd.n5090 585
R2589 gnd.n5128 gnd.n5091 585
R2590 gnd.n5180 gnd.n5179 585
R2591 gnd.n5179 gnd.n5178 585
R2592 gnd.n5181 gnd.n5078 585
R2593 gnd.n5160 gnd.n5078 585
R2594 gnd.n5183 gnd.n5182 585
R2595 gnd.n5184 gnd.n5183 585
R2596 gnd.n5079 gnd.n5077 585
R2597 gnd.n5077 gnd.n5072 585
R2598 gnd.n5083 gnd.n5082 585
R2599 gnd.n5082 gnd.n2890 585
R2600 gnd.n5081 gnd.n2807 585
R2601 gnd.n5192 gnd.n2807 585
R2602 gnd.n5395 gnd.n5394 585
R2603 gnd.n5393 gnd.n2806 585
R2604 gnd.n5392 gnd.n2805 585
R2605 gnd.n5397 gnd.n2805 585
R2606 gnd.n5391 gnd.n5390 585
R2607 gnd.n5389 gnd.n5388 585
R2608 gnd.n5387 gnd.n5386 585
R2609 gnd.n5385 gnd.n5384 585
R2610 gnd.n5383 gnd.n5382 585
R2611 gnd.n5381 gnd.n5380 585
R2612 gnd.n5379 gnd.n5378 585
R2613 gnd.n5377 gnd.n5376 585
R2614 gnd.n5375 gnd.n5374 585
R2615 gnd.n5373 gnd.n5372 585
R2616 gnd.n5371 gnd.n5370 585
R2617 gnd.n5369 gnd.n5368 585
R2618 gnd.n5367 gnd.n5366 585
R2619 gnd.n5365 gnd.n5364 585
R2620 gnd.n5363 gnd.n5362 585
R2621 gnd.n5360 gnd.n5359 585
R2622 gnd.n5358 gnd.n5357 585
R2623 gnd.n5356 gnd.n5355 585
R2624 gnd.n5354 gnd.n5353 585
R2625 gnd.n5352 gnd.n5351 585
R2626 gnd.n5350 gnd.n5349 585
R2627 gnd.n5348 gnd.n5347 585
R2628 gnd.n5346 gnd.n5345 585
R2629 gnd.n5343 gnd.n5342 585
R2630 gnd.n5341 gnd.n5340 585
R2631 gnd.n5339 gnd.n5338 585
R2632 gnd.n5337 gnd.n5336 585
R2633 gnd.n5335 gnd.n5334 585
R2634 gnd.n5333 gnd.n5332 585
R2635 gnd.n5331 gnd.n5330 585
R2636 gnd.n5329 gnd.n5328 585
R2637 gnd.n5327 gnd.n5326 585
R2638 gnd.n5325 gnd.n5324 585
R2639 gnd.n5323 gnd.n5322 585
R2640 gnd.n5321 gnd.n5320 585
R2641 gnd.n5319 gnd.n5318 585
R2642 gnd.n5317 gnd.n5316 585
R2643 gnd.n5315 gnd.n5314 585
R2644 gnd.n5313 gnd.n5312 585
R2645 gnd.n5311 gnd.n5310 585
R2646 gnd.n5309 gnd.n5308 585
R2647 gnd.n5307 gnd.n5306 585
R2648 gnd.n5305 gnd.n5304 585
R2649 gnd.n5303 gnd.n5302 585
R2650 gnd.n5301 gnd.n5300 585
R2651 gnd.n5299 gnd.n5298 585
R2652 gnd.n5297 gnd.n5296 585
R2653 gnd.n5295 gnd.n5294 585
R2654 gnd.n5293 gnd.n5292 585
R2655 gnd.n5291 gnd.n5290 585
R2656 gnd.n5289 gnd.n5288 585
R2657 gnd.n5287 gnd.n5286 585
R2658 gnd.n5285 gnd.n5284 585
R2659 gnd.n2887 gnd.n2870 585
R2660 gnd.n7203 gnd.n7202 585
R2661 gnd.n6880 gnd.n6879 585
R2662 gnd.n7080 gnd.n7079 585
R2663 gnd.n7082 gnd.n7081 585
R2664 gnd.n7084 gnd.n7083 585
R2665 gnd.n7086 gnd.n7085 585
R2666 gnd.n7088 gnd.n7087 585
R2667 gnd.n7090 gnd.n7089 585
R2668 gnd.n7092 gnd.n7091 585
R2669 gnd.n7094 gnd.n7093 585
R2670 gnd.n7096 gnd.n7095 585
R2671 gnd.n7098 gnd.n7097 585
R2672 gnd.n7100 gnd.n7099 585
R2673 gnd.n7102 gnd.n7101 585
R2674 gnd.n7104 gnd.n7103 585
R2675 gnd.n7106 gnd.n7105 585
R2676 gnd.n7108 gnd.n7107 585
R2677 gnd.n7110 gnd.n7109 585
R2678 gnd.n7112 gnd.n7111 585
R2679 gnd.n7115 gnd.n7114 585
R2680 gnd.n7113 gnd.n7059 585
R2681 gnd.n7120 gnd.n7119 585
R2682 gnd.n7122 gnd.n7121 585
R2683 gnd.n7124 gnd.n7123 585
R2684 gnd.n7126 gnd.n7125 585
R2685 gnd.n7128 gnd.n7127 585
R2686 gnd.n7130 gnd.n7129 585
R2687 gnd.n7132 gnd.n7131 585
R2688 gnd.n7134 gnd.n7133 585
R2689 gnd.n7136 gnd.n7135 585
R2690 gnd.n7138 gnd.n7137 585
R2691 gnd.n7140 gnd.n7139 585
R2692 gnd.n7142 gnd.n7141 585
R2693 gnd.n7144 gnd.n7143 585
R2694 gnd.n7146 gnd.n7145 585
R2695 gnd.n7148 gnd.n7147 585
R2696 gnd.n7150 gnd.n7149 585
R2697 gnd.n7152 gnd.n7151 585
R2698 gnd.n7154 gnd.n7153 585
R2699 gnd.n7156 gnd.n7155 585
R2700 gnd.n7158 gnd.n7157 585
R2701 gnd.n7163 gnd.n7162 585
R2702 gnd.n7165 gnd.n7164 585
R2703 gnd.n7167 gnd.n7166 585
R2704 gnd.n7169 gnd.n7168 585
R2705 gnd.n7171 gnd.n7170 585
R2706 gnd.n7173 gnd.n7172 585
R2707 gnd.n7175 gnd.n7174 585
R2708 gnd.n7177 gnd.n7176 585
R2709 gnd.n7179 gnd.n7178 585
R2710 gnd.n7181 gnd.n7180 585
R2711 gnd.n7183 gnd.n7182 585
R2712 gnd.n7185 gnd.n7184 585
R2713 gnd.n7187 gnd.n7186 585
R2714 gnd.n7189 gnd.n7188 585
R2715 gnd.n7192 gnd.n7191 585
R2716 gnd.n7190 gnd.n7025 585
R2717 gnd.n7196 gnd.n7022 585
R2718 gnd.n7198 gnd.n7197 585
R2719 gnd.n7199 gnd.n7198 585
R2720 gnd.n7201 gnd.n6874 585
R2721 gnd.n7201 gnd.n165 585
R2722 gnd.n6873 gnd.n163 585
R2723 gnd.n7210 gnd.n163 585
R2724 gnd.n6872 gnd.n6871 585
R2725 gnd.n6871 gnd.n155 585
R2726 gnd.n6869 gnd.n153 585
R2727 gnd.n7216 gnd.n153 585
R2728 gnd.n6868 gnd.n6867 585
R2729 gnd.n6867 gnd.n146 585
R2730 gnd.n6866 gnd.n144 585
R2731 gnd.n7222 gnd.n144 585
R2732 gnd.n6865 gnd.n6864 585
R2733 gnd.n6864 gnd.n143 585
R2734 gnd.n6862 gnd.n133 585
R2735 gnd.n7228 gnd.n133 585
R2736 gnd.n6861 gnd.n6860 585
R2737 gnd.n6860 gnd.n126 585
R2738 gnd.n6859 gnd.n124 585
R2739 gnd.n7234 gnd.n124 585
R2740 gnd.n6858 gnd.n6857 585
R2741 gnd.n6857 gnd.n116 585
R2742 gnd.n6855 gnd.n114 585
R2743 gnd.n7240 gnd.n114 585
R2744 gnd.n6854 gnd.n6853 585
R2745 gnd.n6853 gnd.n107 585
R2746 gnd.n6852 gnd.n105 585
R2747 gnd.n7246 gnd.n105 585
R2748 gnd.n6851 gnd.n6850 585
R2749 gnd.n6850 gnd.n104 585
R2750 gnd.n6848 gnd.n95 585
R2751 gnd.n7252 gnd.n95 585
R2752 gnd.n6847 gnd.n6846 585
R2753 gnd.n6846 gnd.n86 585
R2754 gnd.n6845 gnd.n84 585
R2755 gnd.n7258 gnd.n84 585
R2756 gnd.n6844 gnd.n6843 585
R2757 gnd.n6843 gnd.n74 585
R2758 gnd.n168 gnd.n73 585
R2759 gnd.n7264 gnd.n73 585
R2760 gnd.n6836 gnd.n6835 585
R2761 gnd.n6837 gnd.n6836 585
R2762 gnd.n6834 gnd.n173 585
R2763 gnd.n173 gnd.n172 585
R2764 gnd.n178 gnd.n174 585
R2765 gnd.n6829 gnd.n178 585
R2766 gnd.n6813 gnd.n6812 585
R2767 gnd.n6812 gnd.n189 585
R2768 gnd.n6814 gnd.n187 585
R2769 gnd.n6818 gnd.n187 585
R2770 gnd.n6811 gnd.n6810 585
R2771 gnd.n6810 gnd.n6809 585
R2772 gnd.n194 gnd.n193 585
R2773 gnd.n195 gnd.n194 585
R2774 gnd.n6777 gnd.n202 585
R2775 gnd.n6796 gnd.n202 585
R2776 gnd.n6776 gnd.n6775 585
R2777 gnd.n6775 gnd.n6774 585
R2778 gnd.n6773 gnd.n212 585
R2779 gnd.n6786 gnd.n212 585
R2780 gnd.n6772 gnd.n6771 585
R2781 gnd.n6771 gnd.n6770 585
R2782 gnd.n222 gnd.n220 585
R2783 gnd.n6744 gnd.n222 585
R2784 gnd.n5101 gnd.n230 585
R2785 gnd.n6761 gnd.n230 585
R2786 gnd.n5104 gnd.n5103 585
R2787 gnd.n5103 gnd.n5102 585
R2788 gnd.n5105 gnd.n240 585
R2789 gnd.n6751 gnd.n240 585
R2790 gnd.n5172 gnd.n5171 585
R2791 gnd.n5171 gnd.n5170 585
R2792 gnd.n5106 gnd.n5100 585
R2793 gnd.n5128 gnd.n5106 585
R2794 gnd.n5157 gnd.n5093 585
R2795 gnd.n5178 gnd.n5093 585
R2796 gnd.n5159 gnd.n5158 585
R2797 gnd.n5160 gnd.n5159 585
R2798 gnd.n5143 gnd.n5073 585
R2799 gnd.n5184 gnd.n5073 585
R2800 gnd.n5148 gnd.n5147 585
R2801 gnd.n5147 gnd.n5072 585
R2802 gnd.n5149 gnd.n5146 585
R2803 gnd.n5146 gnd.n2890 585
R2804 gnd.n5145 gnd.n2888 585
R2805 gnd.n5192 gnd.n2888 585
R2806 gnd.n762 gnd.n761 585
R2807 gnd.n2393 gnd.n762 585
R2808 gnd.n6737 gnd.n6736 585
R2809 gnd.n6737 gnd.n203 585
R2810 gnd.n6739 gnd.n6738 585
R2811 gnd.n6738 gnd.n214 585
R2812 gnd.n6740 gnd.n251 585
R2813 gnd.n251 gnd.n211 585
R2814 gnd.n6742 gnd.n6741 585
R2815 gnd.n6743 gnd.n6742 585
R2816 gnd.n252 gnd.n250 585
R2817 gnd.n250 gnd.n231 585
R2818 gnd.n5121 gnd.n5120 585
R2819 gnd.n5121 gnd.n229 585
R2820 gnd.n5123 gnd.n5122 585
R2821 gnd.n5122 gnd.n242 585
R2822 gnd.n5124 gnd.n5108 585
R2823 gnd.n5108 gnd.n239 585
R2824 gnd.n5126 gnd.n5125 585
R2825 gnd.n5127 gnd.n5126 585
R2826 gnd.n5109 gnd.n5107 585
R2827 gnd.n5107 gnd.n5095 585
R2828 gnd.n5112 gnd.n5111 585
R2829 gnd.n5111 gnd.n5092 585
R2830 gnd.n5070 gnd.n5069 585
R2831 gnd.n5075 gnd.n5070 585
R2832 gnd.n5187 gnd.n5186 585
R2833 gnd.n5186 gnd.n5185 585
R2834 gnd.n5188 gnd.n2892 585
R2835 gnd.n5071 gnd.n2892 585
R2836 gnd.n5190 gnd.n5189 585
R2837 gnd.n5191 gnd.n5190 585
R2838 gnd.n2893 gnd.n2891 585
R2839 gnd.n2891 gnd.n2886 585
R2840 gnd.n5063 gnd.n5062 585
R2841 gnd.n5062 gnd.n2804 585
R2842 gnd.n5061 gnd.n2895 585
R2843 gnd.n5061 gnd.n2766 585
R2844 gnd.n5060 gnd.n5058 585
R2845 gnd.n5060 gnd.n5059 585
R2846 gnd.n2897 gnd.n2896 585
R2847 gnd.n2896 gnd.n2746 585
R2848 gnd.n5054 gnd.n5053 585
R2849 gnd.n5053 gnd.n2732 585
R2850 gnd.n5052 gnd.n2899 585
R2851 gnd.n5052 gnd.n5051 585
R2852 gnd.n5022 gnd.n2900 585
R2853 gnd.n2901 gnd.n2900 585
R2854 gnd.n5024 gnd.n5023 585
R2855 gnd.n5025 gnd.n5024 585
R2856 gnd.n2910 gnd.n2909 585
R2857 gnd.n2909 gnd.n2908 585
R2858 gnd.n5017 gnd.n5016 585
R2859 gnd.n5016 gnd.n5015 585
R2860 gnd.n2913 gnd.n2912 585
R2861 gnd.n2914 gnd.n2913 585
R2862 gnd.n5005 gnd.n5004 585
R2863 gnd.n5006 gnd.n5005 585
R2864 gnd.n2921 gnd.n2920 585
R2865 gnd.n4996 gnd.n2920 585
R2866 gnd.n5000 gnd.n4999 585
R2867 gnd.n4999 gnd.n4998 585
R2868 gnd.n2924 gnd.n2923 585
R2869 gnd.n2925 gnd.n2924 585
R2870 gnd.n4987 gnd.n4986 585
R2871 gnd.n4988 gnd.n4987 585
R2872 gnd.n2933 gnd.n2932 585
R2873 gnd.n2932 gnd.n2931 585
R2874 gnd.n4982 gnd.n4981 585
R2875 gnd.n4981 gnd.n4980 585
R2876 gnd.n2936 gnd.n2935 585
R2877 gnd.n2937 gnd.n2936 585
R2878 gnd.n4815 gnd.n4814 585
R2879 gnd.n4816 gnd.n4815 585
R2880 gnd.n2985 gnd.n2984 585
R2881 gnd.n4741 gnd.n2984 585
R2882 gnd.n4810 gnd.n4809 585
R2883 gnd.n4809 gnd.n4808 585
R2884 gnd.n2988 gnd.n2987 585
R2885 gnd.n4799 gnd.n2988 585
R2886 gnd.n4758 gnd.n3025 585
R2887 gnd.n4758 gnd.n4757 585
R2888 gnd.n4759 gnd.n3022 585
R2889 gnd.n4759 gnd.n3000 585
R2890 gnd.n4761 gnd.n4760 585
R2891 gnd.n4760 gnd.n3005 585
R2892 gnd.n4762 gnd.n3017 585
R2893 gnd.n4734 gnd.n3017 585
R2894 gnd.n4764 gnd.n4763 585
R2895 gnd.n4765 gnd.n4764 585
R2896 gnd.n3018 gnd.n3016 585
R2897 gnd.n3016 gnd.n3013 585
R2898 gnd.n4724 gnd.n4723 585
R2899 gnd.n4725 gnd.n4724 585
R2900 gnd.n3039 gnd.n3038 585
R2901 gnd.n3046 gnd.n3038 585
R2902 gnd.n4718 gnd.n4717 585
R2903 gnd.n4717 gnd.n4716 585
R2904 gnd.n3042 gnd.n3041 585
R2905 gnd.n3051 gnd.n3042 585
R2906 gnd.n4680 gnd.n3066 585
R2907 gnd.n3066 gnd.n3058 585
R2908 gnd.n4682 gnd.n4681 585
R2909 gnd.n4683 gnd.n4682 585
R2910 gnd.n3067 gnd.n3065 585
R2911 gnd.n4647 gnd.n3065 585
R2912 gnd.n4675 gnd.n4674 585
R2913 gnd.n4674 gnd.n4673 585
R2914 gnd.n3070 gnd.n3069 585
R2915 gnd.n4665 gnd.n3070 585
R2916 gnd.n4638 gnd.n3090 585
R2917 gnd.n3090 gnd.n3089 585
R2918 gnd.n4640 gnd.n4639 585
R2919 gnd.n4641 gnd.n4640 585
R2920 gnd.n3091 gnd.n3088 585
R2921 gnd.n3098 gnd.n3088 585
R2922 gnd.n4633 gnd.n4632 585
R2923 gnd.n4632 gnd.n4631 585
R2924 gnd.n3094 gnd.n3093 585
R2925 gnd.n3103 gnd.n3094 585
R2926 gnd.n4584 gnd.n3119 585
R2927 gnd.n3119 gnd.n3109 585
R2928 gnd.n4586 gnd.n4585 585
R2929 gnd.n4587 gnd.n4586 585
R2930 gnd.n3120 gnd.n3118 585
R2931 gnd.n3118 gnd.n3114 585
R2932 gnd.n4579 gnd.n4578 585
R2933 gnd.n4578 gnd.n4577 585
R2934 gnd.n3123 gnd.n3122 585
R2935 gnd.n4569 gnd.n3123 585
R2936 gnd.n4544 gnd.n3142 585
R2937 gnd.n3142 gnd.n3130 585
R2938 gnd.n4546 gnd.n4545 585
R2939 gnd.n4547 gnd.n4546 585
R2940 gnd.n3143 gnd.n3141 585
R2941 gnd.n4474 gnd.n3141 585
R2942 gnd.n4539 gnd.n4538 585
R2943 gnd.n4538 gnd.n4537 585
R2944 gnd.n3146 gnd.n3145 585
R2945 gnd.n4524 gnd.n3146 585
R2946 gnd.n4512 gnd.n3167 585
R2947 gnd.n3167 gnd.n3166 585
R2948 gnd.n4514 gnd.n4513 585
R2949 gnd.n4515 gnd.n4514 585
R2950 gnd.n3168 gnd.n3164 585
R2951 gnd.n3175 gnd.n3164 585
R2952 gnd.n4507 gnd.n4506 585
R2953 gnd.n4506 gnd.n4505 585
R2954 gnd.n3171 gnd.n3170 585
R2955 gnd.n3181 gnd.n3171 585
R2956 gnd.n4443 gnd.n3196 585
R2957 gnd.n3196 gnd.n3188 585
R2958 gnd.n4445 gnd.n4444 585
R2959 gnd.n4446 gnd.n4445 585
R2960 gnd.n3197 gnd.n3195 585
R2961 gnd.n3195 gnd.n3192 585
R2962 gnd.n4438 gnd.n4437 585
R2963 gnd.n4437 gnd.n4436 585
R2964 gnd.n3200 gnd.n3199 585
R2965 gnd.n4427 gnd.n3200 585
R2966 gnd.n4402 gnd.n3217 585
R2967 gnd.n4315 gnd.n3217 585
R2968 gnd.n4404 gnd.n4403 585
R2969 gnd.n4405 gnd.n4404 585
R2970 gnd.n3218 gnd.n3216 585
R2971 gnd.n4331 gnd.n3216 585
R2972 gnd.n4397 gnd.n4396 585
R2973 gnd.n4396 gnd.n4395 585
R2974 gnd.n3221 gnd.n3220 585
R2975 gnd.n4382 gnd.n3221 585
R2976 gnd.n4370 gnd.n3240 585
R2977 gnd.n4311 gnd.n3240 585
R2978 gnd.n4372 gnd.n4371 585
R2979 gnd.n4373 gnd.n4372 585
R2980 gnd.n3241 gnd.n3239 585
R2981 gnd.n4343 gnd.n3239 585
R2982 gnd.n4365 gnd.n4364 585
R2983 gnd.n4364 gnd.n4363 585
R2984 gnd.n3244 gnd.n3243 585
R2985 gnd.n3252 gnd.n3244 585
R2986 gnd.n4296 gnd.n3268 585
R2987 gnd.n3268 gnd.n3260 585
R2988 gnd.n4298 gnd.n4297 585
R2989 gnd.n4299 gnd.n4298 585
R2990 gnd.n3269 gnd.n3267 585
R2991 gnd.n3267 gnd.n3264 585
R2992 gnd.n4291 gnd.n4290 585
R2993 gnd.n4290 gnd.n4289 585
R2994 gnd.n3272 gnd.n3271 585
R2995 gnd.n4281 gnd.n3272 585
R2996 gnd.n4267 gnd.n4266 585
R2997 gnd.n4268 gnd.n4267 585
R2998 gnd.n3286 gnd.n3285 585
R2999 gnd.n4222 gnd.n3285 585
R3000 gnd.n4262 gnd.n4261 585
R3001 gnd.n4261 gnd.n4260 585
R3002 gnd.n3289 gnd.n3288 585
R3003 gnd.n4249 gnd.n3289 585
R3004 gnd.n4200 gnd.n4199 585
R3005 gnd.n4199 gnd.n3297 585
R3006 gnd.n4201 gnd.n3315 585
R3007 gnd.n3315 gnd.n3306 585
R3008 gnd.n4203 gnd.n4202 585
R3009 gnd.n4204 gnd.n4203 585
R3010 gnd.n3316 gnd.n3314 585
R3011 gnd.n3324 gnd.n3314 585
R3012 gnd.n4193 gnd.n4192 585
R3013 gnd.n4192 gnd.n4191 585
R3014 gnd.n3319 gnd.n3318 585
R3015 gnd.n3328 gnd.n3319 585
R3016 gnd.n3337 gnd.n3336 585
R3017 gnd.n3338 gnd.n3337 585
R3018 gnd.n2616 gnd.n2615 585
R3019 gnd.n4164 gnd.n2616 585
R3020 gnd.n5545 gnd.n5544 585
R3021 gnd.n5544 gnd.n5543 585
R3022 gnd.n5546 gnd.n2610 585
R3023 gnd.n4141 gnd.n2610 585
R3024 gnd.n5548 gnd.n5547 585
R3025 gnd.n5549 gnd.n5548 585
R3026 gnd.n2611 gnd.n2609 585
R3027 gnd.n4029 gnd.n2609 585
R3028 gnd.n4050 gnd.n3356 585
R3029 gnd.n3356 gnd.n2579 585
R3030 gnd.n4052 gnd.n4051 585
R3031 gnd.n4053 gnd.n4052 585
R3032 gnd.n3357 gnd.n3355 585
R3033 gnd.n3355 gnd.n3353 585
R3034 gnd.n4044 gnd.n4043 585
R3035 gnd.n4043 gnd.n4042 585
R3036 gnd.n3360 gnd.n3359 585
R3037 gnd.n3361 gnd.n3360 585
R3038 gnd.n4021 gnd.n4020 585
R3039 gnd.n4022 gnd.n4021 585
R3040 gnd.n3372 gnd.n3371 585
R3041 gnd.n3378 gnd.n3371 585
R3042 gnd.n4016 gnd.n4015 585
R3043 gnd.n4015 gnd.n4014 585
R3044 gnd.n3375 gnd.n3374 585
R3045 gnd.n3376 gnd.n3375 585
R3046 gnd.n4005 gnd.n4004 585
R3047 gnd.n4006 gnd.n4005 585
R3048 gnd.n3387 gnd.n3386 585
R3049 gnd.n3386 gnd.n3384 585
R3050 gnd.n4000 gnd.n3999 585
R3051 gnd.n3999 gnd.n3998 585
R3052 gnd.n3390 gnd.n3389 585
R3053 gnd.n3391 gnd.n3390 585
R3054 gnd.n3913 gnd.n3909 585
R3055 gnd.n3909 gnd.n3411 585
R3056 gnd.n3915 gnd.n3914 585
R3057 gnd.n3915 gnd.n3398 585
R3058 gnd.n3917 gnd.n3908 585
R3059 gnd.n3917 gnd.n3916 585
R3060 gnd.n3919 gnd.n3918 585
R3061 gnd.n3918 gnd.n2485 585
R3062 gnd.n3920 gnd.n3619 585
R3063 gnd.n3619 gnd.n2474 585
R3064 gnd.n3922 gnd.n3921 585
R3065 gnd.n3923 gnd.n3922 585
R3066 gnd.n3620 gnd.n3618 585
R3067 gnd.n3618 gnd.n2467 585
R3068 gnd.n3902 gnd.n3901 585
R3069 gnd.n3901 gnd.n2464 585
R3070 gnd.n3900 gnd.n3622 585
R3071 gnd.n3900 gnd.n2457 585
R3072 gnd.n3899 gnd.n3898 585
R3073 gnd.n3899 gnd.n2454 585
R3074 gnd.n3624 gnd.n3623 585
R3075 gnd.n3623 gnd.n2446 585
R3076 gnd.n3894 gnd.n3893 585
R3077 gnd.n3893 gnd.n2443 585
R3078 gnd.n3892 gnd.n3626 585
R3079 gnd.n3892 gnd.n2436 585
R3080 gnd.n3891 gnd.n3890 585
R3081 gnd.n3891 gnd.n2433 585
R3082 gnd.n3628 gnd.n3627 585
R3083 gnd.n3627 gnd.n2425 585
R3084 gnd.n3886 gnd.n3885 585
R3085 gnd.n3885 gnd.n3884 585
R3086 gnd.n3641 gnd.n3630 585
R3087 gnd.n3641 gnd.n2416 585
R3088 gnd.n3640 gnd.n3639 585
R3089 gnd.n3640 gnd.n2413 585
R3090 gnd.n3632 gnd.n3631 585
R3091 gnd.n3631 gnd.n2405 585
R3092 gnd.n3635 gnd.n3634 585
R3093 gnd.n3634 gnd.n2402 585
R3094 gnd.n5050 gnd.n5049 585
R3095 gnd.n5051 gnd.n5050 585
R3096 gnd.n2904 gnd.n2902 585
R3097 gnd.n2902 gnd.n2901 585
R3098 gnd.n5027 gnd.n5026 585
R3099 gnd.n5026 gnd.n5025 585
R3100 gnd.n2907 gnd.n2906 585
R3101 gnd.n2908 gnd.n2907 585
R3102 gnd.n5013 gnd.n5012 585
R3103 gnd.n5015 gnd.n5013 585
R3104 gnd.n2916 gnd.n2915 585
R3105 gnd.n2915 gnd.n2914 585
R3106 gnd.n5008 gnd.n5007 585
R3107 gnd.n5007 gnd.n5006 585
R3108 gnd.n2919 gnd.n2918 585
R3109 gnd.n4996 gnd.n2919 585
R3110 gnd.n4995 gnd.n4994 585
R3111 gnd.n4998 gnd.n4995 585
R3112 gnd.n2927 gnd.n2926 585
R3113 gnd.n2926 gnd.n2925 585
R3114 gnd.n4990 gnd.n4989 585
R3115 gnd.n4989 gnd.n4988 585
R3116 gnd.n2930 gnd.n2929 585
R3117 gnd.n2931 gnd.n2930 585
R3118 gnd.n4745 gnd.n2938 585
R3119 gnd.n4980 gnd.n2938 585
R3120 gnd.n4744 gnd.n4743 585
R3121 gnd.n4743 gnd.n2937 585
R3122 gnd.n4749 gnd.n2982 585
R3123 gnd.n4816 gnd.n2982 585
R3124 gnd.n4750 gnd.n4742 585
R3125 gnd.n4742 gnd.n4741 585
R3126 gnd.n4751 gnd.n2989 585
R3127 gnd.n4808 gnd.n2989 585
R3128 gnd.n3028 gnd.n2997 585
R3129 gnd.n4799 gnd.n2997 585
R3130 gnd.n4756 gnd.n4755 585
R3131 gnd.n4757 gnd.n4756 585
R3132 gnd.n3027 gnd.n3026 585
R3133 gnd.n3026 gnd.n3000 585
R3134 gnd.n4737 gnd.n4736 585
R3135 gnd.n4736 gnd.n3005 585
R3136 gnd.n4735 gnd.n4732 585
R3137 gnd.n4735 gnd.n4734 585
R3138 gnd.n4731 gnd.n3015 585
R3139 gnd.n4765 gnd.n3015 585
R3140 gnd.n3034 gnd.n3030 585
R3141 gnd.n3034 gnd.n3013 585
R3142 gnd.n4727 gnd.n4726 585
R3143 gnd.n4726 gnd.n4725 585
R3144 gnd.n3033 gnd.n3032 585
R3145 gnd.n3046 gnd.n3033 585
R3146 gnd.n4652 gnd.n3044 585
R3147 gnd.n4716 gnd.n3044 585
R3148 gnd.n4651 gnd.n4650 585
R3149 gnd.n4650 gnd.n3051 585
R3150 gnd.n4656 gnd.n4649 585
R3151 gnd.n4649 gnd.n3058 585
R3152 gnd.n4657 gnd.n3063 585
R3153 gnd.n4683 gnd.n3063 585
R3154 gnd.n4658 gnd.n4648 585
R3155 gnd.n4648 gnd.n4647 585
R3156 gnd.n3082 gnd.n3072 585
R3157 gnd.n4673 gnd.n3072 585
R3158 gnd.n4663 gnd.n4662 585
R3159 gnd.n4665 gnd.n4663 585
R3160 gnd.n3081 gnd.n3080 585
R3161 gnd.n3089 gnd.n3080 585
R3162 gnd.n4643 gnd.n4642 585
R3163 gnd.n4642 gnd.n4641 585
R3164 gnd.n3085 gnd.n3084 585
R3165 gnd.n3098 gnd.n3085 585
R3166 gnd.n4557 gnd.n3096 585
R3167 gnd.n4631 gnd.n3096 585
R3168 gnd.n4556 gnd.n4555 585
R3169 gnd.n4555 gnd.n3103 585
R3170 gnd.n4561 gnd.n4554 585
R3171 gnd.n4554 gnd.n3109 585
R3172 gnd.n4562 gnd.n3116 585
R3173 gnd.n4587 gnd.n3116 585
R3174 gnd.n4563 gnd.n4553 585
R3175 gnd.n4553 gnd.n3114 585
R3176 gnd.n3134 gnd.n3125 585
R3177 gnd.n4577 gnd.n3125 585
R3178 gnd.n4568 gnd.n4567 585
R3179 gnd.n4569 gnd.n4568 585
R3180 gnd.n3133 gnd.n3132 585
R3181 gnd.n3132 gnd.n3130 585
R3182 gnd.n4549 gnd.n4548 585
R3183 gnd.n4548 gnd.n4547 585
R3184 gnd.n3137 gnd.n3136 585
R3185 gnd.n4474 gnd.n3137 585
R3186 gnd.n3158 gnd.n3148 585
R3187 gnd.n4537 gnd.n3148 585
R3188 gnd.n4523 gnd.n4522 585
R3189 gnd.n4524 gnd.n4523 585
R3190 gnd.n3157 gnd.n3156 585
R3191 gnd.n3166 gnd.n3156 585
R3192 gnd.n4517 gnd.n4516 585
R3193 gnd.n4516 gnd.n4515 585
R3194 gnd.n3161 gnd.n3160 585
R3195 gnd.n3175 gnd.n3161 585
R3196 gnd.n4415 gnd.n3173 585
R3197 gnd.n4505 gnd.n3173 585
R3198 gnd.n4414 gnd.n4413 585
R3199 gnd.n4413 gnd.n3181 585
R3200 gnd.n4419 gnd.n4412 585
R3201 gnd.n4412 gnd.n3188 585
R3202 gnd.n4420 gnd.n3194 585
R3203 gnd.n4446 gnd.n3194 585
R3204 gnd.n4421 gnd.n4411 585
R3205 gnd.n4411 gnd.n3192 585
R3206 gnd.n3210 gnd.n3202 585
R3207 gnd.n4436 gnd.n3202 585
R3208 gnd.n4426 gnd.n4425 585
R3209 gnd.n4427 gnd.n4426 585
R3210 gnd.n3209 gnd.n3208 585
R3211 gnd.n4315 gnd.n3208 585
R3212 gnd.n4407 gnd.n4406 585
R3213 gnd.n4406 gnd.n4405 585
R3214 gnd.n3213 gnd.n3212 585
R3215 gnd.n4331 gnd.n3213 585
R3216 gnd.n3232 gnd.n3223 585
R3217 gnd.n4395 gnd.n3223 585
R3218 gnd.n4381 gnd.n4380 585
R3219 gnd.n4382 gnd.n4381 585
R3220 gnd.n3231 gnd.n3230 585
R3221 gnd.n4311 gnd.n3230 585
R3222 gnd.n4375 gnd.n4374 585
R3223 gnd.n4374 gnd.n4373 585
R3224 gnd.n3235 gnd.n3234 585
R3225 gnd.n4343 gnd.n3235 585
R3226 gnd.n4230 gnd.n3246 585
R3227 gnd.n4363 gnd.n3246 585
R3228 gnd.n4229 gnd.n4228 585
R3229 gnd.n4228 gnd.n3252 585
R3230 gnd.n4234 gnd.n4227 585
R3231 gnd.n4227 gnd.n3260 585
R3232 gnd.n4235 gnd.n3266 585
R3233 gnd.n4299 gnd.n3266 585
R3234 gnd.n4236 gnd.n4226 585
R3235 gnd.n4226 gnd.n3264 585
R3236 gnd.n4224 gnd.n3273 585
R3237 gnd.n4289 gnd.n3273 585
R3238 gnd.n4240 gnd.n3280 585
R3239 gnd.n4281 gnd.n3280 585
R3240 gnd.n4241 gnd.n3284 585
R3241 gnd.n4268 gnd.n3284 585
R3242 gnd.n4242 gnd.n4223 585
R3243 gnd.n4223 gnd.n4222 585
R3244 gnd.n3301 gnd.n3291 585
R3245 gnd.n4260 gnd.n3291 585
R3246 gnd.n4247 gnd.n4246 585
R3247 gnd.n4249 gnd.n4247 585
R3248 gnd.n3300 gnd.n3299 585
R3249 gnd.n3299 gnd.n3297 585
R3250 gnd.n4151 gnd.n4150 585
R3251 gnd.n4150 gnd.n3306 585
R3252 gnd.n4149 gnd.n3312 585
R3253 gnd.n4204 gnd.n3312 585
R3254 gnd.n4155 gnd.n4148 585
R3255 gnd.n4148 gnd.n3324 585
R3256 gnd.n4156 gnd.n3321 585
R3257 gnd.n4191 gnd.n3321 585
R3258 gnd.n4157 gnd.n4147 585
R3259 gnd.n4147 gnd.n3328 585
R3260 gnd.n3345 gnd.n3343 585
R3261 gnd.n3343 gnd.n3338 585
R3262 gnd.n4162 gnd.n4161 585
R3263 gnd.n4164 gnd.n4162 585
R3264 gnd.n3344 gnd.n2617 585
R3265 gnd.n5543 gnd.n2617 585
R3266 gnd.n4143 gnd.n4142 585
R3267 gnd.n4142 gnd.n4141 585
R3268 gnd.n4060 gnd.n2607 585
R3269 gnd.n5549 gnd.n2607 585
R3270 gnd.n4059 gnd.n3348 585
R3271 gnd.n4029 gnd.n3348 585
R3272 gnd.n3352 gnd.n3347 585
R3273 gnd.n3352 gnd.n2579 585
R3274 gnd.n4055 gnd.n4054 585
R3275 gnd.n4054 gnd.n4053 585
R3276 gnd.n3351 gnd.n3350 585
R3277 gnd.n3353 gnd.n3351 585
R3278 gnd.n3424 gnd.n3362 585
R3279 gnd.n4042 gnd.n3362 585
R3280 gnd.n3425 gnd.n3423 585
R3281 gnd.n3423 gnd.n3361 585
R3282 gnd.n3421 gnd.n3370 585
R3283 gnd.n4022 gnd.n3370 585
R3284 gnd.n3429 gnd.n3420 585
R3285 gnd.n3420 gnd.n3378 585
R3286 gnd.n3430 gnd.n3377 585
R3287 gnd.n4014 gnd.n3377 585
R3288 gnd.n3431 gnd.n3419 585
R3289 gnd.n3419 gnd.n3376 585
R3290 gnd.n3417 gnd.n3385 585
R3291 gnd.n4006 gnd.n3385 585
R3292 gnd.n3435 gnd.n3416 585
R3293 gnd.n3416 gnd.n3384 585
R3294 gnd.n3436 gnd.n3392 585
R3295 gnd.n3998 gnd.n3392 585
R3296 gnd.n3437 gnd.n3414 585
R3297 gnd.n3414 gnd.n3391 585
R3298 gnd.n3987 gnd.n3986 585
R3299 gnd.n3985 gnd.n3413 585
R3300 gnd.n3440 gnd.n3412 585
R3301 gnd.n3989 gnd.n3412 585
R3302 gnd.n3981 gnd.n3442 585
R3303 gnd.n3980 gnd.n3443 585
R3304 gnd.n3979 gnd.n3444 585
R3305 gnd.n3448 gnd.n3445 585
R3306 gnd.n3974 gnd.n3449 585
R3307 gnd.n3973 gnd.n3450 585
R3308 gnd.n3972 gnd.n3451 585
R3309 gnd.n3461 gnd.n3452 585
R3310 gnd.n3965 gnd.n3462 585
R3311 gnd.n3964 gnd.n3463 585
R3312 gnd.n3465 gnd.n3464 585
R3313 gnd.n3957 gnd.n3471 585
R3314 gnd.n3956 gnd.n3472 585
R3315 gnd.n3481 gnd.n3473 585
R3316 gnd.n3949 gnd.n3482 585
R3317 gnd.n3948 gnd.n3483 585
R3318 gnd.n3485 gnd.n3484 585
R3319 gnd.n3941 gnd.n3491 585
R3320 gnd.n3940 gnd.n3492 585
R3321 gnd.n3501 gnd.n3493 585
R3322 gnd.n3933 gnd.n3502 585
R3323 gnd.n3932 gnd.n3503 585
R3324 gnd.n3514 gnd.n3513 585
R3325 gnd.n3516 gnd.n3515 585
R3326 gnd.n3397 gnd.n3396 585
R3327 gnd.n3992 gnd.n3991 585
R3328 gnd.n2730 gnd.n2727 585
R3329 gnd.n5051 gnd.n2730 585
R3330 gnd.n5415 gnd.n2726 585
R3331 gnd.n2901 gnd.n2726 585
R3332 gnd.n5416 gnd.n2725 585
R3333 gnd.n5025 gnd.n2725 585
R3334 gnd.n5417 gnd.n2724 585
R3335 gnd.n2908 gnd.n2724 585
R3336 gnd.n5014 gnd.n2722 585
R3337 gnd.n5015 gnd.n5014 585
R3338 gnd.n5421 gnd.n2721 585
R3339 gnd.n2914 gnd.n2721 585
R3340 gnd.n5422 gnd.n2720 585
R3341 gnd.n5006 gnd.n2720 585
R3342 gnd.n5423 gnd.n2719 585
R3343 gnd.n4996 gnd.n2719 585
R3344 gnd.n4997 gnd.n2717 585
R3345 gnd.n4998 gnd.n4997 585
R3346 gnd.n5427 gnd.n2716 585
R3347 gnd.n2925 gnd.n2716 585
R3348 gnd.n5428 gnd.n2715 585
R3349 gnd.n4988 gnd.n2715 585
R3350 gnd.n5429 gnd.n2714 585
R3351 gnd.n2931 gnd.n2714 585
R3352 gnd.n4979 gnd.n2712 585
R3353 gnd.n4980 gnd.n4979 585
R3354 gnd.n5433 gnd.n2711 585
R3355 gnd.n2937 gnd.n2711 585
R3356 gnd.n5434 gnd.n2710 585
R3357 gnd.n4816 gnd.n2710 585
R3358 gnd.n5435 gnd.n2709 585
R3359 gnd.n4741 gnd.n2709 585
R3360 gnd.n4807 gnd.n2707 585
R3361 gnd.n4808 gnd.n4807 585
R3362 gnd.n5439 gnd.n2706 585
R3363 gnd.n4799 gnd.n2706 585
R3364 gnd.n5440 gnd.n2705 585
R3365 gnd.n4757 gnd.n2705 585
R3366 gnd.n5441 gnd.n2704 585
R3367 gnd.n3000 gnd.n2704 585
R3368 gnd.n3004 gnd.n2702 585
R3369 gnd.n3005 gnd.n3004 585
R3370 gnd.n5445 gnd.n2701 585
R3371 gnd.n4734 gnd.n2701 585
R3372 gnd.n5446 gnd.n2700 585
R3373 gnd.n4765 gnd.n2700 585
R3374 gnd.n5447 gnd.n2699 585
R3375 gnd.n3013 gnd.n2699 585
R3376 gnd.n3037 gnd.n2697 585
R3377 gnd.n4725 gnd.n3037 585
R3378 gnd.n5451 gnd.n2696 585
R3379 gnd.n3046 gnd.n2696 585
R3380 gnd.n5452 gnd.n2695 585
R3381 gnd.n4716 gnd.n2695 585
R3382 gnd.n5453 gnd.n2694 585
R3383 gnd.n3051 gnd.n2694 585
R3384 gnd.n3057 gnd.n2692 585
R3385 gnd.n3058 gnd.n3057 585
R3386 gnd.n5457 gnd.n2691 585
R3387 gnd.n4683 gnd.n2691 585
R3388 gnd.n5458 gnd.n2690 585
R3389 gnd.n4647 gnd.n2690 585
R3390 gnd.n5459 gnd.n2689 585
R3391 gnd.n4673 gnd.n2689 585
R3392 gnd.n4664 gnd.n2687 585
R3393 gnd.n4665 gnd.n4664 585
R3394 gnd.n5463 gnd.n2686 585
R3395 gnd.n3089 gnd.n2686 585
R3396 gnd.n5464 gnd.n2685 585
R3397 gnd.n4641 gnd.n2685 585
R3398 gnd.n5465 gnd.n2684 585
R3399 gnd.n3098 gnd.n2684 585
R3400 gnd.n4630 gnd.n2682 585
R3401 gnd.n4631 gnd.n4630 585
R3402 gnd.n5469 gnd.n2681 585
R3403 gnd.n3103 gnd.n2681 585
R3404 gnd.n5470 gnd.n2680 585
R3405 gnd.n3109 gnd.n2680 585
R3406 gnd.n5471 gnd.n2679 585
R3407 gnd.n4587 gnd.n2679 585
R3408 gnd.n3113 gnd.n2677 585
R3409 gnd.n3114 gnd.n3113 585
R3410 gnd.n5475 gnd.n2676 585
R3411 gnd.n4577 gnd.n2676 585
R3412 gnd.n5476 gnd.n2675 585
R3413 gnd.n4569 gnd.n2675 585
R3414 gnd.n5477 gnd.n2674 585
R3415 gnd.n3130 gnd.n2674 585
R3416 gnd.n3140 gnd.n2672 585
R3417 gnd.n4547 gnd.n3140 585
R3418 gnd.n5481 gnd.n2671 585
R3419 gnd.n4474 gnd.n2671 585
R3420 gnd.n5482 gnd.n2670 585
R3421 gnd.n4537 gnd.n2670 585
R3422 gnd.n5483 gnd.n2669 585
R3423 gnd.n4524 gnd.n2669 585
R3424 gnd.n3165 gnd.n2667 585
R3425 gnd.n3166 gnd.n3165 585
R3426 gnd.n5487 gnd.n2666 585
R3427 gnd.n4515 gnd.n2666 585
R3428 gnd.n5488 gnd.n2665 585
R3429 gnd.n3175 gnd.n2665 585
R3430 gnd.n5489 gnd.n2664 585
R3431 gnd.n4505 gnd.n2664 585
R3432 gnd.n3180 gnd.n2662 585
R3433 gnd.n3181 gnd.n3180 585
R3434 gnd.n5493 gnd.n2661 585
R3435 gnd.n3188 gnd.n2661 585
R3436 gnd.n5494 gnd.n2660 585
R3437 gnd.n4446 gnd.n2660 585
R3438 gnd.n5495 gnd.n2659 585
R3439 gnd.n3192 gnd.n2659 585
R3440 gnd.n4435 gnd.n2657 585
R3441 gnd.n4436 gnd.n4435 585
R3442 gnd.n5499 gnd.n2656 585
R3443 gnd.n4427 gnd.n2656 585
R3444 gnd.n5500 gnd.n2655 585
R3445 gnd.n4315 gnd.n2655 585
R3446 gnd.n5501 gnd.n2654 585
R3447 gnd.n4405 gnd.n2654 585
R3448 gnd.n4330 gnd.n2652 585
R3449 gnd.n4331 gnd.n4330 585
R3450 gnd.n5505 gnd.n2651 585
R3451 gnd.n4395 gnd.n2651 585
R3452 gnd.n5506 gnd.n2650 585
R3453 gnd.n4382 gnd.n2650 585
R3454 gnd.n5507 gnd.n2649 585
R3455 gnd.n4311 gnd.n2649 585
R3456 gnd.n3238 gnd.n2647 585
R3457 gnd.n4373 gnd.n3238 585
R3458 gnd.n5511 gnd.n2646 585
R3459 gnd.n4343 gnd.n2646 585
R3460 gnd.n5512 gnd.n2645 585
R3461 gnd.n4363 gnd.n2645 585
R3462 gnd.n5513 gnd.n2644 585
R3463 gnd.n3252 gnd.n2644 585
R3464 gnd.n3259 gnd.n2642 585
R3465 gnd.n3260 gnd.n3259 585
R3466 gnd.n5517 gnd.n2641 585
R3467 gnd.n4299 gnd.n2641 585
R3468 gnd.n5518 gnd.n2640 585
R3469 gnd.n3264 gnd.n2640 585
R3470 gnd.n5519 gnd.n2639 585
R3471 gnd.n4289 gnd.n2639 585
R3472 gnd.n4280 gnd.n2637 585
R3473 gnd.n4281 gnd.n4280 585
R3474 gnd.n5523 gnd.n2636 585
R3475 gnd.n4268 gnd.n2636 585
R3476 gnd.n5524 gnd.n2635 585
R3477 gnd.n4222 gnd.n2635 585
R3478 gnd.n5525 gnd.n2634 585
R3479 gnd.n4260 gnd.n2634 585
R3480 gnd.n4248 gnd.n2632 585
R3481 gnd.n4249 gnd.n4248 585
R3482 gnd.n5529 gnd.n2631 585
R3483 gnd.n3297 gnd.n2631 585
R3484 gnd.n5530 gnd.n2630 585
R3485 gnd.n3306 gnd.n2630 585
R3486 gnd.n5531 gnd.n2629 585
R3487 gnd.n4204 gnd.n2629 585
R3488 gnd.n3323 gnd.n2627 585
R3489 gnd.n3324 gnd.n3323 585
R3490 gnd.n5535 gnd.n2626 585
R3491 gnd.n4191 gnd.n2626 585
R3492 gnd.n5536 gnd.n2625 585
R3493 gnd.n3328 gnd.n2625 585
R3494 gnd.n5537 gnd.n2624 585
R3495 gnd.n3338 gnd.n2624 585
R3496 gnd.n2621 gnd.n2619 585
R3497 gnd.n4164 gnd.n2619 585
R3498 gnd.n5542 gnd.n5541 585
R3499 gnd.n5543 gnd.n5542 585
R3500 gnd.n2620 gnd.n2618 585
R3501 gnd.n4141 gnd.n2618 585
R3502 gnd.n4031 gnd.n2608 585
R3503 gnd.n5549 gnd.n2608 585
R3504 gnd.n4034 gnd.n4030 585
R3505 gnd.n4030 gnd.n4029 585
R3506 gnd.n4035 gnd.n4028 585
R3507 gnd.n4028 gnd.n2579 585
R3508 gnd.n4036 gnd.n3354 585
R3509 gnd.n4053 gnd.n3354 585
R3510 gnd.n3366 gnd.n3364 585
R3511 gnd.n3364 gnd.n3353 585
R3512 gnd.n4041 gnd.n4040 585
R3513 gnd.n4042 gnd.n4041 585
R3514 gnd.n3365 gnd.n3363 585
R3515 gnd.n3363 gnd.n3361 585
R3516 gnd.n4024 gnd.n4023 585
R3517 gnd.n4023 gnd.n4022 585
R3518 gnd.n3369 gnd.n3368 585
R3519 gnd.n3378 gnd.n3369 585
R3520 gnd.n4013 gnd.n4012 585
R3521 gnd.n4014 gnd.n4013 585
R3522 gnd.n3380 gnd.n3379 585
R3523 gnd.n3379 gnd.n3376 585
R3524 gnd.n4008 gnd.n4007 585
R3525 gnd.n4007 gnd.n4006 585
R3526 gnd.n3383 gnd.n3382 585
R3527 gnd.n3384 gnd.n3383 585
R3528 gnd.n3997 gnd.n3996 585
R3529 gnd.n3998 gnd.n3997 585
R3530 gnd.n3394 gnd.n3393 585
R3531 gnd.n3393 gnd.n3391 585
R3532 gnd.n5407 gnd.n5406 585
R3533 gnd.n5408 gnd.n5407 585
R3534 gnd.n2749 gnd.n2747 585
R3535 gnd.n5234 gnd.n5233 585
R3536 gnd.n5244 gnd.n5232 585
R3537 gnd.n5245 gnd.n5231 585
R3538 gnd.n5230 gnd.n5222 585
R3539 gnd.n5252 gnd.n5221 585
R3540 gnd.n5253 gnd.n5220 585
R3541 gnd.n5214 gnd.n5213 585
R3542 gnd.n5260 gnd.n5212 585
R3543 gnd.n5261 gnd.n5211 585
R3544 gnd.n5210 gnd.n5202 585
R3545 gnd.n5268 gnd.n5201 585
R3546 gnd.n5269 gnd.n5200 585
R3547 gnd.n2881 gnd.n2880 585
R3548 gnd.n5276 gnd.n2879 585
R3549 gnd.n5277 gnd.n2878 585
R3550 gnd.n5278 gnd.n2877 585
R3551 gnd.n5037 gnd.n2876 585
R3552 gnd.n5039 gnd.n5038 585
R3553 gnd.n5040 gnd.n5036 585
R3554 gnd.n5035 gnd.n5033 585
R3555 gnd.n5044 gnd.n5032 585
R3556 gnd.n5045 gnd.n5031 585
R3557 gnd.n5046 gnd.n2903 585
R3558 gnd.n5411 gnd.n5410 585
R3559 gnd.n2731 gnd.n2729 585
R3560 gnd.n2762 gnd.n2761 585
R3561 gnd.n2760 gnd.n2748 585
R3562 gnd.n4909 gnd.n2978 506.916
R3563 gnd.n4912 gnd.n4911 506.916
R3564 gnd.n4128 gnd.n4127 506.916
R3565 gnd.n5618 gnd.n2582 506.916
R3566 gnd.n6168 gnd.n6167 396.406
R3567 gnd.n4063 gnd.t296 389.64
R3568 gnd.n2973 gnd.t221 389.64
R3569 gnd.n5555 gnd.t231 389.64
R3570 gnd.n4840 gnd.t278 389.64
R3571 gnd.n3504 gnd.t246 371.625
R3572 gnd.n5400 gnd.t206 371.625
R3573 gnd.n6877 gnd.t228 371.625
R3574 gnd.n7060 gnd.t263 371.625
R3575 gnd.n7159 gnd.t275 371.625
R3576 gnd.n2826 gnd.t290 371.625
R3577 gnd.n2849 gnd.t293 371.625
R3578 gnd.n2871 gnd.t253 371.625
R3579 gnd.n6892 gnd.t193 371.625
R3580 gnd.n3509 gnd.t242 371.625
R3581 gnd.n3673 gnd.t235 371.625
R3582 gnd.n2215 gnd.t250 371.625
R3583 gnd.n2237 gnd.t272 371.625
R3584 gnd.n2259 gnd.t284 371.625
R3585 gnd.n2531 gnd.t266 371.625
R3586 gnd.n3521 gnd.t287 371.625
R3587 gnd.n3533 gnd.t306 371.625
R3588 gnd.n2750 gnd.t214 371.625
R3589 gnd.n1335 gnd.t256 323.425
R3590 gnd.n784 gnd.t309 323.425
R3591 gnd.n2123 gnd.n2097 289.615
R3592 gnd.n2091 gnd.n2065 289.615
R3593 gnd.n2059 gnd.n2033 289.615
R3594 gnd.n2028 gnd.n2002 289.615
R3595 gnd.n1996 gnd.n1970 289.615
R3596 gnd.n1964 gnd.n1938 289.615
R3597 gnd.n1932 gnd.n1906 289.615
R3598 gnd.n1901 gnd.n1875 289.615
R3599 gnd.n1409 gnd.t299 279.217
R3600 gnd.n805 gnd.t210 279.217
R3601 gnd.n2589 gnd.t271 260.649
R3602 gnd.n4832 gnd.t283 260.649
R3603 gnd.n5620 gnd.n5619 256.663
R3604 gnd.n5620 gnd.n2548 256.663
R3605 gnd.n5620 gnd.n2549 256.663
R3606 gnd.n5620 gnd.n2550 256.663
R3607 gnd.n5620 gnd.n2551 256.663
R3608 gnd.n5620 gnd.n2552 256.663
R3609 gnd.n5620 gnd.n2553 256.663
R3610 gnd.n5620 gnd.n2554 256.663
R3611 gnd.n5620 gnd.n2555 256.663
R3612 gnd.n5620 gnd.n2556 256.663
R3613 gnd.n5620 gnd.n2557 256.663
R3614 gnd.n5620 gnd.n2558 256.663
R3615 gnd.n5620 gnd.n2559 256.663
R3616 gnd.n5620 gnd.n2560 256.663
R3617 gnd.n5620 gnd.n2561 256.663
R3618 gnd.n5620 gnd.n2562 256.663
R3619 gnd.n5623 gnd.n2546 256.663
R3620 gnd.n5621 gnd.n5620 256.663
R3621 gnd.n5620 gnd.n2563 256.663
R3622 gnd.n5620 gnd.n2564 256.663
R3623 gnd.n5620 gnd.n2565 256.663
R3624 gnd.n5620 gnd.n2566 256.663
R3625 gnd.n5620 gnd.n2567 256.663
R3626 gnd.n5620 gnd.n2568 256.663
R3627 gnd.n5620 gnd.n2569 256.663
R3628 gnd.n5620 gnd.n2570 256.663
R3629 gnd.n5620 gnd.n2571 256.663
R3630 gnd.n5620 gnd.n2572 256.663
R3631 gnd.n5620 gnd.n2573 256.663
R3632 gnd.n5620 gnd.n2574 256.663
R3633 gnd.n5620 gnd.n2575 256.663
R3634 gnd.n5620 gnd.n2576 256.663
R3635 gnd.n5620 gnd.n2577 256.663
R3636 gnd.n5620 gnd.n2578 256.663
R3637 gnd.n4978 gnd.n2956 256.663
R3638 gnd.n4978 gnd.n2957 256.663
R3639 gnd.n4978 gnd.n2958 256.663
R3640 gnd.n4978 gnd.n2959 256.663
R3641 gnd.n4978 gnd.n2960 256.663
R3642 gnd.n4978 gnd.n2961 256.663
R3643 gnd.n4978 gnd.n2962 256.663
R3644 gnd.n4978 gnd.n2963 256.663
R3645 gnd.n4978 gnd.n2964 256.663
R3646 gnd.n4978 gnd.n2965 256.663
R3647 gnd.n4978 gnd.n2966 256.663
R3648 gnd.n4978 gnd.n2967 256.663
R3649 gnd.n4978 gnd.n2968 256.663
R3650 gnd.n4978 gnd.n2969 256.663
R3651 gnd.n4978 gnd.n2970 256.663
R3652 gnd.n4978 gnd.n2971 256.663
R3653 gnd.n2972 gnd.n2836 256.663
R3654 gnd.n4978 gnd.n2955 256.663
R3655 gnd.n4978 gnd.n2954 256.663
R3656 gnd.n4978 gnd.n2953 256.663
R3657 gnd.n4978 gnd.n2952 256.663
R3658 gnd.n4978 gnd.n2951 256.663
R3659 gnd.n4978 gnd.n2950 256.663
R3660 gnd.n4978 gnd.n2949 256.663
R3661 gnd.n4978 gnd.n2948 256.663
R3662 gnd.n4978 gnd.n2947 256.663
R3663 gnd.n4978 gnd.n2946 256.663
R3664 gnd.n4978 gnd.n2945 256.663
R3665 gnd.n4978 gnd.n2944 256.663
R3666 gnd.n4978 gnd.n2943 256.663
R3667 gnd.n4978 gnd.n2942 256.663
R3668 gnd.n4978 gnd.n2941 256.663
R3669 gnd.n4978 gnd.n2940 256.663
R3670 gnd.n4978 gnd.n2939 256.663
R3671 gnd.n5928 gnd.n2183 242.672
R3672 gnd.n5928 gnd.n2184 242.672
R3673 gnd.n5928 gnd.n2185 242.672
R3674 gnd.n5928 gnd.n2186 242.672
R3675 gnd.n5928 gnd.n2187 242.672
R3676 gnd.n5928 gnd.n2188 242.672
R3677 gnd.n5928 gnd.n2189 242.672
R3678 gnd.n5928 gnd.n2190 242.672
R3679 gnd.n5928 gnd.n2191 242.672
R3680 gnd.n5674 gnd.n2484 242.672
R3681 gnd.n5674 gnd.n2483 242.672
R3682 gnd.n5674 gnd.n2482 242.672
R3683 gnd.n5674 gnd.n2481 242.672
R3684 gnd.n5674 gnd.n2480 242.672
R3685 gnd.n5674 gnd.n2479 242.672
R3686 gnd.n5674 gnd.n2478 242.672
R3687 gnd.n5674 gnd.n2477 242.672
R3688 gnd.n5674 gnd.n2476 242.672
R3689 gnd.n1463 gnd.n1462 242.672
R3690 gnd.n1463 gnd.n1373 242.672
R3691 gnd.n1463 gnd.n1374 242.672
R3692 gnd.n1463 gnd.n1375 242.672
R3693 gnd.n1463 gnd.n1376 242.672
R3694 gnd.n1463 gnd.n1377 242.672
R3695 gnd.n1463 gnd.n1378 242.672
R3696 gnd.n1463 gnd.n1379 242.672
R3697 gnd.n1463 gnd.n1380 242.672
R3698 gnd.n1463 gnd.n1381 242.672
R3699 gnd.n1463 gnd.n1382 242.672
R3700 gnd.n1463 gnd.n1383 242.672
R3701 gnd.n1464 gnd.n1463 242.672
R3702 gnd.n5975 gnd.n2154 242.672
R3703 gnd.n5975 gnd.n801 242.672
R3704 gnd.n5975 gnd.n800 242.672
R3705 gnd.n5975 gnd.n799 242.672
R3706 gnd.n5975 gnd.n798 242.672
R3707 gnd.n5975 gnd.n797 242.672
R3708 gnd.n5975 gnd.n796 242.672
R3709 gnd.n5975 gnd.n795 242.672
R3710 gnd.n5975 gnd.n794 242.672
R3711 gnd.n5975 gnd.n793 242.672
R3712 gnd.n5975 gnd.n792 242.672
R3713 gnd.n5975 gnd.n791 242.672
R3714 gnd.n5975 gnd.n790 242.672
R3715 gnd.n5397 gnd.n2795 242.672
R3716 gnd.n5397 gnd.n2796 242.672
R3717 gnd.n5397 gnd.n2797 242.672
R3718 gnd.n5397 gnd.n2798 242.672
R3719 gnd.n5397 gnd.n2799 242.672
R3720 gnd.n5397 gnd.n2800 242.672
R3721 gnd.n5397 gnd.n2801 242.672
R3722 gnd.n5397 gnd.n2803 242.672
R3723 gnd.n5398 gnd.n5397 242.672
R3724 gnd.n7199 gnd.n6993 242.672
R3725 gnd.n7199 gnd.n6889 242.672
R3726 gnd.n7199 gnd.n6888 242.672
R3727 gnd.n7199 gnd.n6887 242.672
R3728 gnd.n7199 gnd.n6886 242.672
R3729 gnd.n7199 gnd.n6885 242.672
R3730 gnd.n7199 gnd.n6884 242.672
R3731 gnd.n7199 gnd.n6883 242.672
R3732 gnd.n7199 gnd.n6882 242.672
R3733 gnd.n1547 gnd.n1546 242.672
R3734 gnd.n1546 gnd.n1285 242.672
R3735 gnd.n1546 gnd.n1286 242.672
R3736 gnd.n1546 gnd.n1287 242.672
R3737 gnd.n1546 gnd.n1288 242.672
R3738 gnd.n1546 gnd.n1289 242.672
R3739 gnd.n1546 gnd.n1290 242.672
R3740 gnd.n1546 gnd.n1291 242.672
R3741 gnd.n5975 gnd.n783 242.672
R3742 gnd.n5976 gnd.n5975 242.672
R3743 gnd.n5975 gnd.n5929 242.672
R3744 gnd.n5975 gnd.n5930 242.672
R3745 gnd.n5975 gnd.n5931 242.672
R3746 gnd.n5975 gnd.n5932 242.672
R3747 gnd.n5975 gnd.n5933 242.672
R3748 gnd.n5975 gnd.n5934 242.672
R3749 gnd.n5928 gnd.n5927 242.672
R3750 gnd.n5928 gnd.n2155 242.672
R3751 gnd.n5928 gnd.n2156 242.672
R3752 gnd.n5928 gnd.n2157 242.672
R3753 gnd.n5928 gnd.n2158 242.672
R3754 gnd.n5928 gnd.n2159 242.672
R3755 gnd.n5928 gnd.n2160 242.672
R3756 gnd.n5928 gnd.n2161 242.672
R3757 gnd.n5928 gnd.n2162 242.672
R3758 gnd.n5928 gnd.n2163 242.672
R3759 gnd.n5928 gnd.n2164 242.672
R3760 gnd.n5928 gnd.n2165 242.672
R3761 gnd.n5928 gnd.n2166 242.672
R3762 gnd.n5928 gnd.n2167 242.672
R3763 gnd.n5928 gnd.n2168 242.672
R3764 gnd.n5928 gnd.n2169 242.672
R3765 gnd.n5928 gnd.n2170 242.672
R3766 gnd.n5928 gnd.n2171 242.672
R3767 gnd.n5928 gnd.n2172 242.672
R3768 gnd.n5928 gnd.n2173 242.672
R3769 gnd.n5928 gnd.n2174 242.672
R3770 gnd.n5928 gnd.n2175 242.672
R3771 gnd.n5928 gnd.n2176 242.672
R3772 gnd.n5928 gnd.n2177 242.672
R3773 gnd.n5928 gnd.n2178 242.672
R3774 gnd.n5928 gnd.n2179 242.672
R3775 gnd.n5928 gnd.n2180 242.672
R3776 gnd.n5928 gnd.n2181 242.672
R3777 gnd.n5928 gnd.n2182 242.672
R3778 gnd.n5674 gnd.n2486 242.672
R3779 gnd.n5674 gnd.n2487 242.672
R3780 gnd.n5674 gnd.n2488 242.672
R3781 gnd.n5674 gnd.n2489 242.672
R3782 gnd.n5674 gnd.n2490 242.672
R3783 gnd.n5674 gnd.n2491 242.672
R3784 gnd.n5674 gnd.n2492 242.672
R3785 gnd.n5674 gnd.n2493 242.672
R3786 gnd.n5674 gnd.n2494 242.672
R3787 gnd.n5674 gnd.n2495 242.672
R3788 gnd.n5674 gnd.n2496 242.672
R3789 gnd.n5674 gnd.n2497 242.672
R3790 gnd.n5674 gnd.n2498 242.672
R3791 gnd.n5674 gnd.n2499 242.672
R3792 gnd.n5674 gnd.n2500 242.672
R3793 gnd.n5674 gnd.n2501 242.672
R3794 gnd.n5624 gnd.n2542 242.672
R3795 gnd.n5674 gnd.n2502 242.672
R3796 gnd.n5674 gnd.n2503 242.672
R3797 gnd.n5674 gnd.n2504 242.672
R3798 gnd.n5674 gnd.n2505 242.672
R3799 gnd.n5674 gnd.n2506 242.672
R3800 gnd.n5674 gnd.n2507 242.672
R3801 gnd.n5674 gnd.n2508 242.672
R3802 gnd.n5674 gnd.n2509 242.672
R3803 gnd.n5674 gnd.n2510 242.672
R3804 gnd.n5674 gnd.n2511 242.672
R3805 gnd.n5674 gnd.n2512 242.672
R3806 gnd.n5674 gnd.n2513 242.672
R3807 gnd.n5674 gnd.n5673 242.672
R3808 gnd.n5397 gnd.n5396 242.672
R3809 gnd.n5397 gnd.n2767 242.672
R3810 gnd.n5397 gnd.n2768 242.672
R3811 gnd.n5397 gnd.n2769 242.672
R3812 gnd.n5397 gnd.n2770 242.672
R3813 gnd.n5397 gnd.n2771 242.672
R3814 gnd.n5397 gnd.n2772 242.672
R3815 gnd.n5397 gnd.n2773 242.672
R3816 gnd.n5397 gnd.n2774 242.672
R3817 gnd.n5397 gnd.n2775 242.672
R3818 gnd.n5397 gnd.n2776 242.672
R3819 gnd.n5397 gnd.n2777 242.672
R3820 gnd.n5397 gnd.n2778 242.672
R3821 gnd.n5344 gnd.n2837 242.672
R3822 gnd.n5397 gnd.n2779 242.672
R3823 gnd.n5397 gnd.n2780 242.672
R3824 gnd.n5397 gnd.n2781 242.672
R3825 gnd.n5397 gnd.n2782 242.672
R3826 gnd.n5397 gnd.n2783 242.672
R3827 gnd.n5397 gnd.n2784 242.672
R3828 gnd.n5397 gnd.n2785 242.672
R3829 gnd.n5397 gnd.n2786 242.672
R3830 gnd.n5397 gnd.n2787 242.672
R3831 gnd.n5397 gnd.n2788 242.672
R3832 gnd.n5397 gnd.n2789 242.672
R3833 gnd.n5397 gnd.n2790 242.672
R3834 gnd.n5397 gnd.n2791 242.672
R3835 gnd.n5397 gnd.n2792 242.672
R3836 gnd.n5397 gnd.n2793 242.672
R3837 gnd.n5397 gnd.n2794 242.672
R3838 gnd.n7200 gnd.n7199 242.672
R3839 gnd.n7199 gnd.n6994 242.672
R3840 gnd.n7199 gnd.n6995 242.672
R3841 gnd.n7199 gnd.n6996 242.672
R3842 gnd.n7199 gnd.n6997 242.672
R3843 gnd.n7199 gnd.n6998 242.672
R3844 gnd.n7199 gnd.n6999 242.672
R3845 gnd.n7199 gnd.n7000 242.672
R3846 gnd.n7199 gnd.n7001 242.672
R3847 gnd.n7199 gnd.n7002 242.672
R3848 gnd.n7199 gnd.n7003 242.672
R3849 gnd.n7199 gnd.n7004 242.672
R3850 gnd.n7199 gnd.n7005 242.672
R3851 gnd.n7199 gnd.n7006 242.672
R3852 gnd.n7199 gnd.n7007 242.672
R3853 gnd.n7199 gnd.n7008 242.672
R3854 gnd.n7199 gnd.n7009 242.672
R3855 gnd.n7199 gnd.n7010 242.672
R3856 gnd.n7199 gnd.n7011 242.672
R3857 gnd.n7199 gnd.n7012 242.672
R3858 gnd.n7199 gnd.n7013 242.672
R3859 gnd.n7199 gnd.n7014 242.672
R3860 gnd.n7199 gnd.n7015 242.672
R3861 gnd.n7199 gnd.n7016 242.672
R3862 gnd.n7199 gnd.n7017 242.672
R3863 gnd.n7199 gnd.n7018 242.672
R3864 gnd.n7199 gnd.n7019 242.672
R3865 gnd.n7199 gnd.n7020 242.672
R3866 gnd.n7199 gnd.n7021 242.672
R3867 gnd.n3989 gnd.n3988 242.672
R3868 gnd.n3989 gnd.n3399 242.672
R3869 gnd.n3989 gnd.n3400 242.672
R3870 gnd.n3989 gnd.n3401 242.672
R3871 gnd.n3989 gnd.n3402 242.672
R3872 gnd.n3989 gnd.n3403 242.672
R3873 gnd.n3989 gnd.n3404 242.672
R3874 gnd.n3989 gnd.n3405 242.672
R3875 gnd.n3989 gnd.n3406 242.672
R3876 gnd.n3989 gnd.n3407 242.672
R3877 gnd.n3989 gnd.n3408 242.672
R3878 gnd.n3989 gnd.n3409 242.672
R3879 gnd.n3989 gnd.n3410 242.672
R3880 gnd.n3990 gnd.n3989 242.672
R3881 gnd.n5408 gnd.n2744 242.672
R3882 gnd.n5408 gnd.n2743 242.672
R3883 gnd.n5408 gnd.n2742 242.672
R3884 gnd.n5408 gnd.n2741 242.672
R3885 gnd.n5408 gnd.n2740 242.672
R3886 gnd.n5408 gnd.n2739 242.672
R3887 gnd.n5408 gnd.n2738 242.672
R3888 gnd.n5408 gnd.n2737 242.672
R3889 gnd.n5408 gnd.n2736 242.672
R3890 gnd.n5408 gnd.n2735 242.672
R3891 gnd.n5408 gnd.n2734 242.672
R3892 gnd.n5408 gnd.n2733 242.672
R3893 gnd.n5409 gnd.n5408 242.672
R3894 gnd.n5408 gnd.n2745 242.672
R3895 gnd.n7198 gnd.n7022 240.244
R3896 gnd.n7191 gnd.n7190 240.244
R3897 gnd.n7188 gnd.n7187 240.244
R3898 gnd.n7184 gnd.n7183 240.244
R3899 gnd.n7180 gnd.n7179 240.244
R3900 gnd.n7176 gnd.n7175 240.244
R3901 gnd.n7172 gnd.n7171 240.244
R3902 gnd.n7168 gnd.n7167 240.244
R3903 gnd.n7164 gnd.n7163 240.244
R3904 gnd.n7157 gnd.n7156 240.244
R3905 gnd.n7153 gnd.n7152 240.244
R3906 gnd.n7149 gnd.n7148 240.244
R3907 gnd.n7145 gnd.n7144 240.244
R3908 gnd.n7141 gnd.n7140 240.244
R3909 gnd.n7137 gnd.n7136 240.244
R3910 gnd.n7133 gnd.n7132 240.244
R3911 gnd.n7129 gnd.n7128 240.244
R3912 gnd.n7125 gnd.n7124 240.244
R3913 gnd.n7121 gnd.n7120 240.244
R3914 gnd.n7114 gnd.n7113 240.244
R3915 gnd.n7111 gnd.n7110 240.244
R3916 gnd.n7107 gnd.n7106 240.244
R3917 gnd.n7103 gnd.n7102 240.244
R3918 gnd.n7099 gnd.n7098 240.244
R3919 gnd.n7095 gnd.n7094 240.244
R3920 gnd.n7091 gnd.n7090 240.244
R3921 gnd.n7087 gnd.n7086 240.244
R3922 gnd.n7083 gnd.n7082 240.244
R3923 gnd.n7079 gnd.n6880 240.244
R3924 gnd.n5146 gnd.n2888 240.244
R3925 gnd.n5147 gnd.n5146 240.244
R3926 gnd.n5147 gnd.n5073 240.244
R3927 gnd.n5159 gnd.n5073 240.244
R3928 gnd.n5159 gnd.n5093 240.244
R3929 gnd.n5106 gnd.n5093 240.244
R3930 gnd.n5171 gnd.n5106 240.244
R3931 gnd.n5171 gnd.n240 240.244
R3932 gnd.n5103 gnd.n240 240.244
R3933 gnd.n5103 gnd.n230 240.244
R3934 gnd.n230 gnd.n222 240.244
R3935 gnd.n6771 gnd.n222 240.244
R3936 gnd.n6771 gnd.n212 240.244
R3937 gnd.n6775 gnd.n212 240.244
R3938 gnd.n6775 gnd.n202 240.244
R3939 gnd.n202 gnd.n194 240.244
R3940 gnd.n6810 gnd.n194 240.244
R3941 gnd.n6810 gnd.n187 240.244
R3942 gnd.n6812 gnd.n187 240.244
R3943 gnd.n6812 gnd.n178 240.244
R3944 gnd.n178 gnd.n173 240.244
R3945 gnd.n6836 gnd.n173 240.244
R3946 gnd.n6836 gnd.n73 240.244
R3947 gnd.n6843 gnd.n73 240.244
R3948 gnd.n6843 gnd.n84 240.244
R3949 gnd.n6846 gnd.n84 240.244
R3950 gnd.n6846 gnd.n95 240.244
R3951 gnd.n6850 gnd.n95 240.244
R3952 gnd.n6850 gnd.n105 240.244
R3953 gnd.n6853 gnd.n105 240.244
R3954 gnd.n6853 gnd.n114 240.244
R3955 gnd.n6857 gnd.n114 240.244
R3956 gnd.n6857 gnd.n124 240.244
R3957 gnd.n6860 gnd.n124 240.244
R3958 gnd.n6860 gnd.n133 240.244
R3959 gnd.n6864 gnd.n133 240.244
R3960 gnd.n6864 gnd.n144 240.244
R3961 gnd.n6867 gnd.n144 240.244
R3962 gnd.n6867 gnd.n153 240.244
R3963 gnd.n6871 gnd.n153 240.244
R3964 gnd.n6871 gnd.n163 240.244
R3965 gnd.n7201 gnd.n163 240.244
R3966 gnd.n2806 gnd.n2805 240.244
R3967 gnd.n5390 gnd.n2805 240.244
R3968 gnd.n5388 gnd.n5387 240.244
R3969 gnd.n5384 gnd.n5383 240.244
R3970 gnd.n5380 gnd.n5379 240.244
R3971 gnd.n5376 gnd.n5375 240.244
R3972 gnd.n5372 gnd.n5371 240.244
R3973 gnd.n5368 gnd.n5367 240.244
R3974 gnd.n5364 gnd.n5363 240.244
R3975 gnd.n5359 gnd.n5358 240.244
R3976 gnd.n5355 gnd.n5354 240.244
R3977 gnd.n5351 gnd.n5350 240.244
R3978 gnd.n5347 gnd.n5346 240.244
R3979 gnd.n5342 gnd.n5341 240.244
R3980 gnd.n5338 gnd.n5337 240.244
R3981 gnd.n5334 gnd.n5333 240.244
R3982 gnd.n5330 gnd.n5329 240.244
R3983 gnd.n5326 gnd.n5325 240.244
R3984 gnd.n5322 gnd.n5321 240.244
R3985 gnd.n5318 gnd.n5317 240.244
R3986 gnd.n5314 gnd.n5313 240.244
R3987 gnd.n5310 gnd.n5309 240.244
R3988 gnd.n5306 gnd.n5305 240.244
R3989 gnd.n5302 gnd.n5301 240.244
R3990 gnd.n5298 gnd.n5297 240.244
R3991 gnd.n5294 gnd.n5293 240.244
R3992 gnd.n5290 gnd.n5289 240.244
R3993 gnd.n5286 gnd.n5285 240.244
R3994 gnd.n5082 gnd.n2807 240.244
R3995 gnd.n5082 gnd.n5077 240.244
R3996 gnd.n5183 gnd.n5077 240.244
R3997 gnd.n5183 gnd.n5078 240.244
R3998 gnd.n5179 gnd.n5078 240.244
R3999 gnd.n5179 gnd.n5091 240.244
R4000 gnd.n5091 gnd.n238 240.244
R4001 gnd.n6752 gnd.n238 240.244
R4002 gnd.n6752 gnd.n233 240.244
R4003 gnd.n6760 gnd.n233 240.244
R4004 gnd.n6760 gnd.n234 240.244
R4005 gnd.n234 gnd.n210 240.244
R4006 gnd.n6787 gnd.n210 240.244
R4007 gnd.n6787 gnd.n205 240.244
R4008 gnd.n6795 gnd.n205 240.244
R4009 gnd.n6795 gnd.n206 240.244
R4010 gnd.n206 gnd.n186 240.244
R4011 gnd.n6819 gnd.n186 240.244
R4012 gnd.n6819 gnd.n181 240.244
R4013 gnd.n6828 gnd.n181 240.244
R4014 gnd.n6828 gnd.n182 240.244
R4015 gnd.n182 gnd.n76 240.244
R4016 gnd.n7263 gnd.n76 240.244
R4017 gnd.n7263 gnd.n77 240.244
R4018 gnd.n7259 gnd.n77 240.244
R4019 gnd.n7259 gnd.n83 240.244
R4020 gnd.n7251 gnd.n83 240.244
R4021 gnd.n7251 gnd.n97 240.244
R4022 gnd.n7247 gnd.n97 240.244
R4023 gnd.n7247 gnd.n103 240.244
R4024 gnd.n7239 gnd.n103 240.244
R4025 gnd.n7239 gnd.n117 240.244
R4026 gnd.n7235 gnd.n117 240.244
R4027 gnd.n7235 gnd.n123 240.244
R4028 gnd.n7227 gnd.n123 240.244
R4029 gnd.n7227 gnd.n136 240.244
R4030 gnd.n7223 gnd.n136 240.244
R4031 gnd.n7223 gnd.n142 240.244
R4032 gnd.n7215 gnd.n142 240.244
R4033 gnd.n7215 gnd.n156 240.244
R4034 gnd.n7211 gnd.n156 240.244
R4035 gnd.n7211 gnd.n162 240.244
R4036 gnd.n5675 gnd.n2473 240.244
R4037 gnd.n5672 gnd.n2514 240.244
R4038 gnd.n5668 gnd.n5667 240.244
R4039 gnd.n5664 gnd.n5663 240.244
R4040 gnd.n5660 gnd.n5659 240.244
R4041 gnd.n5656 gnd.n5655 240.244
R4042 gnd.n5652 gnd.n5651 240.244
R4043 gnd.n5648 gnd.n5647 240.244
R4044 gnd.n5644 gnd.n5643 240.244
R4045 gnd.n5639 gnd.n5638 240.244
R4046 gnd.n5635 gnd.n5634 240.244
R4047 gnd.n5631 gnd.n5630 240.244
R4048 gnd.n5627 gnd.n5626 240.244
R4049 gnd.n3540 gnd.n3539 240.244
R4050 gnd.n3547 gnd.n3546 240.244
R4051 gnd.n3550 gnd.n3549 240.244
R4052 gnd.n3557 gnd.n3556 240.244
R4053 gnd.n3560 gnd.n3559 240.244
R4054 gnd.n3567 gnd.n3566 240.244
R4055 gnd.n3570 gnd.n3569 240.244
R4056 gnd.n3577 gnd.n3576 240.244
R4057 gnd.n3580 gnd.n3579 240.244
R4058 gnd.n3587 gnd.n3586 240.244
R4059 gnd.n3590 gnd.n3589 240.244
R4060 gnd.n3597 gnd.n3596 240.244
R4061 gnd.n3600 gnd.n3599 240.244
R4062 gnd.n3607 gnd.n3606 240.244
R4063 gnd.n3610 gnd.n3609 240.244
R4064 gnd.n2269 gnd.n2268 240.244
R4065 gnd.n3783 gnd.n2269 240.244
R4066 gnd.n3783 gnd.n2279 240.244
R4067 gnd.n3786 gnd.n2279 240.244
R4068 gnd.n3786 gnd.n2289 240.244
R4069 gnd.n3790 gnd.n2289 240.244
R4070 gnd.n3790 gnd.n2298 240.244
R4071 gnd.n3793 gnd.n2298 240.244
R4072 gnd.n3793 gnd.n2307 240.244
R4073 gnd.n3797 gnd.n2307 240.244
R4074 gnd.n3797 gnd.n2317 240.244
R4075 gnd.n3800 gnd.n2317 240.244
R4076 gnd.n3800 gnd.n2326 240.244
R4077 gnd.n3804 gnd.n2326 240.244
R4078 gnd.n3804 gnd.n2336 240.244
R4079 gnd.n3807 gnd.n2336 240.244
R4080 gnd.n3807 gnd.n2345 240.244
R4081 gnd.n3811 gnd.n2345 240.244
R4082 gnd.n3811 gnd.n2355 240.244
R4083 gnd.n3814 gnd.n2355 240.244
R4084 gnd.n3814 gnd.n2364 240.244
R4085 gnd.n3818 gnd.n2364 240.244
R4086 gnd.n3818 gnd.n2374 240.244
R4087 gnd.n3821 gnd.n2374 240.244
R4088 gnd.n3821 gnd.n2383 240.244
R4089 gnd.n3825 gnd.n2383 240.244
R4090 gnd.n3825 gnd.n2394 240.244
R4091 gnd.n3829 gnd.n2394 240.244
R4092 gnd.n3829 gnd.n2403 240.244
R4093 gnd.n3839 gnd.n2403 240.244
R4094 gnd.n3839 gnd.n2414 240.244
R4095 gnd.n3642 gnd.n2414 240.244
R4096 gnd.n3642 gnd.n2423 240.244
R4097 gnd.n3846 gnd.n2423 240.244
R4098 gnd.n3846 gnd.n2434 240.244
R4099 gnd.n3850 gnd.n2434 240.244
R4100 gnd.n3850 gnd.n2444 240.244
R4101 gnd.n3855 gnd.n2444 240.244
R4102 gnd.n3855 gnd.n2455 240.244
R4103 gnd.n3862 gnd.n2455 240.244
R4104 gnd.n3862 gnd.n2465 240.244
R4105 gnd.n3617 gnd.n2465 240.244
R4106 gnd.n2195 gnd.n2194 240.244
R4107 gnd.n5921 gnd.n2194 240.244
R4108 gnd.n5919 gnd.n5918 240.244
R4109 gnd.n5915 gnd.n5914 240.244
R4110 gnd.n5911 gnd.n5910 240.244
R4111 gnd.n5907 gnd.n5906 240.244
R4112 gnd.n5903 gnd.n5902 240.244
R4113 gnd.n5899 gnd.n5898 240.244
R4114 gnd.n5895 gnd.n5894 240.244
R4115 gnd.n5890 gnd.n5889 240.244
R4116 gnd.n5886 gnd.n5885 240.244
R4117 gnd.n5882 gnd.n5881 240.244
R4118 gnd.n5878 gnd.n5877 240.244
R4119 gnd.n5874 gnd.n5873 240.244
R4120 gnd.n5870 gnd.n5869 240.244
R4121 gnd.n5866 gnd.n5865 240.244
R4122 gnd.n5862 gnd.n5861 240.244
R4123 gnd.n5858 gnd.n5857 240.244
R4124 gnd.n5854 gnd.n5853 240.244
R4125 gnd.n5850 gnd.n5849 240.244
R4126 gnd.n5846 gnd.n5845 240.244
R4127 gnd.n5842 gnd.n5841 240.244
R4128 gnd.n5838 gnd.n5837 240.244
R4129 gnd.n5834 gnd.n5833 240.244
R4130 gnd.n5830 gnd.n5829 240.244
R4131 gnd.n5826 gnd.n5825 240.244
R4132 gnd.n5822 gnd.n5821 240.244
R4133 gnd.n5818 gnd.n5817 240.244
R4134 gnd.n5814 gnd.n5813 240.244
R4135 gnd.n5803 gnd.n2196 240.244
R4136 gnd.n5803 gnd.n2271 240.244
R4137 gnd.n5797 gnd.n2271 240.244
R4138 gnd.n5797 gnd.n2277 240.244
R4139 gnd.n5789 gnd.n2277 240.244
R4140 gnd.n5789 gnd.n2292 240.244
R4141 gnd.n5785 gnd.n2292 240.244
R4142 gnd.n5785 gnd.n2297 240.244
R4143 gnd.n5777 gnd.n2297 240.244
R4144 gnd.n5777 gnd.n2309 240.244
R4145 gnd.n5773 gnd.n2309 240.244
R4146 gnd.n5773 gnd.n2315 240.244
R4147 gnd.n5765 gnd.n2315 240.244
R4148 gnd.n5765 gnd.n2329 240.244
R4149 gnd.n5761 gnd.n2329 240.244
R4150 gnd.n5761 gnd.n2335 240.244
R4151 gnd.n5753 gnd.n2335 240.244
R4152 gnd.n5753 gnd.n2347 240.244
R4153 gnd.n5749 gnd.n2347 240.244
R4154 gnd.n5749 gnd.n2353 240.244
R4155 gnd.n5741 gnd.n2353 240.244
R4156 gnd.n5741 gnd.n2367 240.244
R4157 gnd.n5737 gnd.n2367 240.244
R4158 gnd.n5737 gnd.n2373 240.244
R4159 gnd.n5729 gnd.n2373 240.244
R4160 gnd.n5729 gnd.n2386 240.244
R4161 gnd.n5725 gnd.n2386 240.244
R4162 gnd.n5725 gnd.n2392 240.244
R4163 gnd.n5717 gnd.n2392 240.244
R4164 gnd.n5717 gnd.n2406 240.244
R4165 gnd.n5713 gnd.n2406 240.244
R4166 gnd.n5713 gnd.n2412 240.244
R4167 gnd.n5705 gnd.n2412 240.244
R4168 gnd.n5705 gnd.n2426 240.244
R4169 gnd.n5701 gnd.n2426 240.244
R4170 gnd.n5701 gnd.n2432 240.244
R4171 gnd.n5693 gnd.n2432 240.244
R4172 gnd.n5693 gnd.n2447 240.244
R4173 gnd.n5689 gnd.n2447 240.244
R4174 gnd.n5689 gnd.n2453 240.244
R4175 gnd.n5681 gnd.n2453 240.244
R4176 gnd.n5681 gnd.n2468 240.244
R4177 gnd.n5974 gnd.n5935 240.244
R4178 gnd.n5967 gnd.n5966 240.244
R4179 gnd.n5964 gnd.n5963 240.244
R4180 gnd.n5960 gnd.n5959 240.244
R4181 gnd.n5956 gnd.n5955 240.244
R4182 gnd.n5952 gnd.n5951 240.244
R4183 gnd.n5948 gnd.n789 240.244
R4184 gnd.n5978 gnd.n5977 240.244
R4185 gnd.n1558 gnd.n1270 240.244
R4186 gnd.n1568 gnd.n1270 240.244
R4187 gnd.n1568 gnd.n1261 240.244
R4188 gnd.n1261 gnd.n1250 240.244
R4189 gnd.n1589 gnd.n1250 240.244
R4190 gnd.n1589 gnd.n1244 240.244
R4191 gnd.n1599 gnd.n1244 240.244
R4192 gnd.n1599 gnd.n1233 240.244
R4193 gnd.n1233 gnd.n1223 240.244
R4194 gnd.n1625 gnd.n1223 240.244
R4195 gnd.n1626 gnd.n1625 240.244
R4196 gnd.n1627 gnd.n1626 240.244
R4197 gnd.n1627 gnd.n1202 240.244
R4198 gnd.n1663 gnd.n1202 240.244
R4199 gnd.n1663 gnd.n1203 240.244
R4200 gnd.n1659 gnd.n1203 240.244
R4201 gnd.n1659 gnd.n1658 240.244
R4202 gnd.n1658 gnd.n1044 240.244
R4203 gnd.n1693 gnd.n1044 240.244
R4204 gnd.n1693 gnd.n1035 240.244
R4205 gnd.n1035 gnd.n1027 240.244
R4206 gnd.n1714 gnd.n1027 240.244
R4207 gnd.n1714 gnd.n1021 240.244
R4208 gnd.n1724 gnd.n1021 240.244
R4209 gnd.n1724 gnd.n1012 240.244
R4210 gnd.n1012 gnd.n1002 240.244
R4211 gnd.n1745 gnd.n1002 240.244
R4212 gnd.n1745 gnd.n995 240.244
R4213 gnd.n1755 gnd.n995 240.244
R4214 gnd.n1755 gnd.n986 240.244
R4215 gnd.n986 gnd.n975 240.244
R4216 gnd.n1776 gnd.n975 240.244
R4217 gnd.n1776 gnd.n969 240.244
R4218 gnd.n1786 gnd.n969 240.244
R4219 gnd.n1786 gnd.n961 240.244
R4220 gnd.n961 gnd.n951 240.244
R4221 gnd.n1807 gnd.n951 240.244
R4222 gnd.n1807 gnd.n945 240.244
R4223 gnd.n1817 gnd.n945 240.244
R4224 gnd.n1817 gnd.n936 240.244
R4225 gnd.n936 gnd.n925 240.244
R4226 gnd.n1838 gnd.n925 240.244
R4227 gnd.n1838 gnd.n919 240.244
R4228 gnd.n1848 gnd.n919 240.244
R4229 gnd.n1848 gnd.n910 240.244
R4230 gnd.n910 gnd.n900 240.244
R4231 gnd.n1870 gnd.n900 240.244
R4232 gnd.n1870 gnd.n893 240.244
R4233 gnd.n2136 gnd.n893 240.244
R4234 gnd.n2136 gnd.n764 240.244
R4235 gnd.n2139 gnd.n764 240.244
R4236 gnd.n2139 gnd.n774 240.244
R4237 gnd.n5985 gnd.n774 240.244
R4238 gnd.n1548 gnd.n1283 240.244
R4239 gnd.n1304 gnd.n1283 240.244
R4240 gnd.n1307 gnd.n1306 240.244
R4241 gnd.n1314 gnd.n1313 240.244
R4242 gnd.n1317 gnd.n1316 240.244
R4243 gnd.n1324 gnd.n1323 240.244
R4244 gnd.n1327 gnd.n1326 240.244
R4245 gnd.n1334 gnd.n1333 240.244
R4246 gnd.n1556 gnd.n1280 240.244
R4247 gnd.n1280 gnd.n1259 240.244
R4248 gnd.n1579 gnd.n1259 240.244
R4249 gnd.n1579 gnd.n1253 240.244
R4250 gnd.n1587 gnd.n1253 240.244
R4251 gnd.n1587 gnd.n1255 240.244
R4252 gnd.n1255 gnd.n1231 240.244
R4253 gnd.n1609 gnd.n1231 240.244
R4254 gnd.n1609 gnd.n1226 240.244
R4255 gnd.n1623 gnd.n1226 240.244
R4256 gnd.n1623 gnd.n1227 240.244
R4257 gnd.n1619 gnd.n1227 240.244
R4258 gnd.n1619 gnd.n1199 240.244
R4259 gnd.n1666 gnd.n1199 240.244
R4260 gnd.n1667 gnd.n1666 240.244
R4261 gnd.n1668 gnd.n1667 240.244
R4262 gnd.n1668 gnd.n1195 240.244
R4263 gnd.n1674 gnd.n1195 240.244
R4264 gnd.n1674 gnd.n1034 240.244
R4265 gnd.n1704 gnd.n1034 240.244
R4266 gnd.n1704 gnd.n1029 240.244
R4267 gnd.n1712 gnd.n1029 240.244
R4268 gnd.n1712 gnd.n1030 240.244
R4269 gnd.n1030 gnd.n1010 240.244
R4270 gnd.n1735 gnd.n1010 240.244
R4271 gnd.n1735 gnd.n1005 240.244
R4272 gnd.n1743 gnd.n1005 240.244
R4273 gnd.n1743 gnd.n1006 240.244
R4274 gnd.n1006 gnd.n984 240.244
R4275 gnd.n1766 gnd.n984 240.244
R4276 gnd.n1766 gnd.n978 240.244
R4277 gnd.n1774 gnd.n978 240.244
R4278 gnd.n1774 gnd.n980 240.244
R4279 gnd.n980 gnd.n959 240.244
R4280 gnd.n1797 gnd.n959 240.244
R4281 gnd.n1797 gnd.n953 240.244
R4282 gnd.n1805 gnd.n953 240.244
R4283 gnd.n1805 gnd.n955 240.244
R4284 gnd.n955 gnd.n934 240.244
R4285 gnd.n1828 gnd.n934 240.244
R4286 gnd.n1828 gnd.n928 240.244
R4287 gnd.n1836 gnd.n928 240.244
R4288 gnd.n1836 gnd.n930 240.244
R4289 gnd.n930 gnd.n908 240.244
R4290 gnd.n1859 gnd.n908 240.244
R4291 gnd.n1859 gnd.n903 240.244
R4292 gnd.n1868 gnd.n903 240.244
R4293 gnd.n1868 gnd.n904 240.244
R4294 gnd.n904 gnd.n765 240.244
R4295 gnd.n5997 gnd.n765 240.244
R4296 gnd.n5997 gnd.n766 240.244
R4297 gnd.n5993 gnd.n766 240.244
R4298 gnd.n5993 gnd.n772 240.244
R4299 gnd.n6903 gnd.n6881 240.244
R4300 gnd.n6909 gnd.n6908 240.244
R4301 gnd.n6912 gnd.n6911 240.244
R4302 gnd.n6919 gnd.n6918 240.244
R4303 gnd.n6922 gnd.n6921 240.244
R4304 gnd.n6929 gnd.n6928 240.244
R4305 gnd.n6932 gnd.n6931 240.244
R4306 gnd.n6939 gnd.n6938 240.244
R4307 gnd.n6941 gnd.n6890 240.244
R4308 gnd.n5137 gnd.n2889 240.244
R4309 gnd.n5137 gnd.n5136 240.244
R4310 gnd.n5136 gnd.n5074 240.244
R4311 gnd.n5161 gnd.n5074 240.244
R4312 gnd.n5161 gnd.n5094 240.244
R4313 gnd.n5129 gnd.n5094 240.244
R4314 gnd.n5169 gnd.n5129 240.244
R4315 gnd.n5169 gnd.n241 240.244
R4316 gnd.n241 gnd.n228 240.244
R4317 gnd.n6762 gnd.n228 240.244
R4318 gnd.n6762 gnd.n223 240.244
R4319 gnd.n6769 gnd.n223 240.244
R4320 gnd.n6769 gnd.n213 240.244
R4321 gnd.n213 gnd.n201 240.244
R4322 gnd.n6797 gnd.n201 240.244
R4323 gnd.n6797 gnd.n196 240.244
R4324 gnd.n6808 gnd.n196 240.244
R4325 gnd.n6808 gnd.n188 240.244
R4326 gnd.n6801 gnd.n188 240.244
R4327 gnd.n6801 gnd.n180 240.244
R4328 gnd.n180 gnd.n179 240.244
R4329 gnd.n179 gnd.n70 240.244
R4330 gnd.n7265 gnd.n70 240.244
R4331 gnd.n7265 gnd.n72 240.244
R4332 gnd.n85 gnd.n72 240.244
R4333 gnd.n6956 gnd.n85 240.244
R4334 gnd.n6956 gnd.n96 240.244
R4335 gnd.n6961 gnd.n96 240.244
R4336 gnd.n6961 gnd.n106 240.244
R4337 gnd.n6964 gnd.n106 240.244
R4338 gnd.n6964 gnd.n115 240.244
R4339 gnd.n6969 gnd.n115 240.244
R4340 gnd.n6969 gnd.n125 240.244
R4341 gnd.n6972 gnd.n125 240.244
R4342 gnd.n6972 gnd.n134 240.244
R4343 gnd.n6977 gnd.n134 240.244
R4344 gnd.n6977 gnd.n145 240.244
R4345 gnd.n6980 gnd.n145 240.244
R4346 gnd.n6980 gnd.n154 240.244
R4347 gnd.n6985 gnd.n154 240.244
R4348 gnd.n6985 gnd.n164 240.244
R4349 gnd.n6891 gnd.n164 240.244
R4350 gnd.n5197 gnd.n5196 240.244
R4351 gnd.n5205 gnd.n5204 240.244
R4352 gnd.n5207 gnd.n5206 240.244
R4353 gnd.n5217 gnd.n5216 240.244
R4354 gnd.n5225 gnd.n5224 240.244
R4355 gnd.n5227 gnd.n5226 240.244
R4356 gnd.n5237 gnd.n5236 240.244
R4357 gnd.n2802 gnd.n2756 240.244
R4358 gnd.n5399 gnd.n2765 240.244
R4359 gnd.n5193 gnd.n2884 240.244
R4360 gnd.n5152 gnd.n2884 240.244
R4361 gnd.n5152 gnd.n5076 240.244
R4362 gnd.n5096 gnd.n5076 240.244
R4363 gnd.n5177 gnd.n5096 240.244
R4364 gnd.n5177 gnd.n5097 240.244
R4365 gnd.n5097 gnd.n243 240.244
R4366 gnd.n6750 gnd.n243 240.244
R4367 gnd.n6750 gnd.n244 240.244
R4368 gnd.n244 gnd.n232 240.244
R4369 gnd.n6745 gnd.n232 240.244
R4370 gnd.n6745 gnd.n215 240.244
R4371 gnd.n6785 gnd.n215 240.244
R4372 gnd.n6785 gnd.n216 240.244
R4373 gnd.n216 gnd.n204 240.244
R4374 gnd.n6780 gnd.n204 240.244
R4375 gnd.n6780 gnd.n190 240.244
R4376 gnd.n6817 gnd.n190 240.244
R4377 gnd.n6817 gnd.n177 240.244
R4378 gnd.n6830 gnd.n177 240.244
R4379 gnd.n6830 gnd.n171 240.244
R4380 gnd.n6838 gnd.n171 240.244
R4381 gnd.n6838 gnd.n75 240.244
R4382 gnd.n87 gnd.n75 240.244
R4383 gnd.n7257 gnd.n87 240.244
R4384 gnd.n7257 gnd.n88 240.244
R4385 gnd.n7253 gnd.n88 240.244
R4386 gnd.n7253 gnd.n94 240.244
R4387 gnd.n7245 gnd.n94 240.244
R4388 gnd.n7245 gnd.n108 240.244
R4389 gnd.n7241 gnd.n108 240.244
R4390 gnd.n7241 gnd.n113 240.244
R4391 gnd.n7233 gnd.n113 240.244
R4392 gnd.n7233 gnd.n127 240.244
R4393 gnd.n7229 gnd.n127 240.244
R4394 gnd.n7229 gnd.n132 240.244
R4395 gnd.n7221 gnd.n132 240.244
R4396 gnd.n7221 gnd.n147 240.244
R4397 gnd.n7217 gnd.n147 240.244
R4398 gnd.n7217 gnd.n152 240.244
R4399 gnd.n7209 gnd.n152 240.244
R4400 gnd.n7209 gnd.n166 240.244
R4401 gnd.n818 gnd.n778 240.244
R4402 gnd.n826 gnd.n825 240.244
R4403 gnd.n829 gnd.n828 240.244
R4404 gnd.n836 gnd.n835 240.244
R4405 gnd.n839 gnd.n838 240.244
R4406 gnd.n846 gnd.n845 240.244
R4407 gnd.n849 gnd.n848 240.244
R4408 gnd.n856 gnd.n855 240.244
R4409 gnd.n859 gnd.n858 240.244
R4410 gnd.n866 gnd.n865 240.244
R4411 gnd.n869 gnd.n868 240.244
R4412 gnd.n876 gnd.n875 240.244
R4413 gnd.n878 gnd.n802 240.244
R4414 gnd.n1471 gnd.n1368 240.244
R4415 gnd.n1471 gnd.n1361 240.244
R4416 gnd.n1482 gnd.n1361 240.244
R4417 gnd.n1482 gnd.n1357 240.244
R4418 gnd.n1488 gnd.n1357 240.244
R4419 gnd.n1488 gnd.n1349 240.244
R4420 gnd.n1498 gnd.n1349 240.244
R4421 gnd.n1498 gnd.n1344 240.244
R4422 gnd.n1534 gnd.n1344 240.244
R4423 gnd.n1534 gnd.n1345 240.244
R4424 gnd.n1345 gnd.n1292 240.244
R4425 gnd.n1529 gnd.n1292 240.244
R4426 gnd.n1529 gnd.n1528 240.244
R4427 gnd.n1528 gnd.n1271 240.244
R4428 gnd.n1524 gnd.n1271 240.244
R4429 gnd.n1524 gnd.n1262 240.244
R4430 gnd.n1521 gnd.n1262 240.244
R4431 gnd.n1521 gnd.n1520 240.244
R4432 gnd.n1520 gnd.n1245 240.244
R4433 gnd.n1516 gnd.n1245 240.244
R4434 gnd.n1516 gnd.n1234 240.244
R4435 gnd.n1234 gnd.n1214 240.244
R4436 gnd.n1635 gnd.n1214 240.244
R4437 gnd.n1635 gnd.n1209 240.244
R4438 gnd.n1643 gnd.n1209 240.244
R4439 gnd.n1643 gnd.n1210 240.244
R4440 gnd.n1210 gnd.n1178 240.244
R4441 gnd.n1683 gnd.n1178 240.244
R4442 gnd.n1683 gnd.n1179 240.244
R4443 gnd.n1194 gnd.n1179 240.244
R4444 gnd.n1194 gnd.n1046 240.244
R4445 gnd.n1690 gnd.n1046 240.244
R4446 gnd.n1690 gnd.n1036 240.244
R4447 gnd.n1120 gnd.n1036 240.244
R4448 gnd.n1123 gnd.n1120 240.244
R4449 gnd.n1123 gnd.n1022 240.244
R4450 gnd.n1117 gnd.n1022 240.244
R4451 gnd.n1117 gnd.n1013 240.244
R4452 gnd.n1114 gnd.n1013 240.244
R4453 gnd.n1114 gnd.n1113 240.244
R4454 gnd.n1113 gnd.n997 240.244
R4455 gnd.n1109 gnd.n997 240.244
R4456 gnd.n1109 gnd.n987 240.244
R4457 gnd.n1106 gnd.n987 240.244
R4458 gnd.n1106 gnd.n1105 240.244
R4459 gnd.n1105 gnd.n970 240.244
R4460 gnd.n1101 gnd.n970 240.244
R4461 gnd.n1101 gnd.n962 240.244
R4462 gnd.n1098 gnd.n962 240.244
R4463 gnd.n1098 gnd.n1095 240.244
R4464 gnd.n1095 gnd.n946 240.244
R4465 gnd.n1091 gnd.n946 240.244
R4466 gnd.n1091 gnd.n937 240.244
R4467 gnd.n1088 gnd.n937 240.244
R4468 gnd.n1088 gnd.n1087 240.244
R4469 gnd.n1087 gnd.n920 240.244
R4470 gnd.n1083 gnd.n920 240.244
R4471 gnd.n1083 gnd.n911 240.244
R4472 gnd.n1080 gnd.n911 240.244
R4473 gnd.n1080 gnd.n1079 240.244
R4474 gnd.n1079 gnd.n895 240.244
R4475 gnd.n895 gnd.n884 240.244
R4476 gnd.n2146 gnd.n884 240.244
R4477 gnd.n2147 gnd.n2146 240.244
R4478 gnd.n2147 gnd.n775 240.244
R4479 gnd.n1385 gnd.n1384 240.244
R4480 gnd.n1456 gnd.n1384 240.244
R4481 gnd.n1454 gnd.n1453 240.244
R4482 gnd.n1450 gnd.n1449 240.244
R4483 gnd.n1446 gnd.n1445 240.244
R4484 gnd.n1442 gnd.n1441 240.244
R4485 gnd.n1438 gnd.n1437 240.244
R4486 gnd.n1434 gnd.n1433 240.244
R4487 gnd.n1430 gnd.n1429 240.244
R4488 gnd.n1426 gnd.n1425 240.244
R4489 gnd.n1422 gnd.n1421 240.244
R4490 gnd.n1418 gnd.n1417 240.244
R4491 gnd.n1414 gnd.n1372 240.244
R4492 gnd.n1474 gnd.n1366 240.244
R4493 gnd.n1474 gnd.n1362 240.244
R4494 gnd.n1480 gnd.n1362 240.244
R4495 gnd.n1480 gnd.n1355 240.244
R4496 gnd.n1490 gnd.n1355 240.244
R4497 gnd.n1490 gnd.n1351 240.244
R4498 gnd.n1496 gnd.n1351 240.244
R4499 gnd.n1496 gnd.n1342 240.244
R4500 gnd.n1536 gnd.n1342 240.244
R4501 gnd.n1536 gnd.n1293 240.244
R4502 gnd.n1544 gnd.n1293 240.244
R4503 gnd.n1544 gnd.n1294 240.244
R4504 gnd.n1294 gnd.n1272 240.244
R4505 gnd.n1565 gnd.n1272 240.244
R4506 gnd.n1565 gnd.n1264 240.244
R4507 gnd.n1576 gnd.n1264 240.244
R4508 gnd.n1576 gnd.n1265 240.244
R4509 gnd.n1265 gnd.n1246 240.244
R4510 gnd.n1596 gnd.n1246 240.244
R4511 gnd.n1596 gnd.n1236 240.244
R4512 gnd.n1606 gnd.n1236 240.244
R4513 gnd.n1606 gnd.n1217 240.244
R4514 gnd.n1633 gnd.n1217 240.244
R4515 gnd.n1633 gnd.n1207 240.244
R4516 gnd.n1646 gnd.n1207 240.244
R4517 gnd.n1647 gnd.n1646 240.244
R4518 gnd.n1647 gnd.n1182 240.244
R4519 gnd.n1681 gnd.n1182 240.244
R4520 gnd.n1681 gnd.n1183 240.244
R4521 gnd.n1677 gnd.n1183 240.244
R4522 gnd.n1677 gnd.n1191 240.244
R4523 gnd.n1191 gnd.n1038 240.244
R4524 gnd.n1701 gnd.n1038 240.244
R4525 gnd.n1701 gnd.n1039 240.244
R4526 gnd.n1039 gnd.n1023 240.244
R4527 gnd.n1721 gnd.n1023 240.244
R4528 gnd.n1721 gnd.n1015 240.244
R4529 gnd.n1732 gnd.n1015 240.244
R4530 gnd.n1732 gnd.n1016 240.244
R4531 gnd.n1016 gnd.n998 240.244
R4532 gnd.n1752 gnd.n998 240.244
R4533 gnd.n1752 gnd.n989 240.244
R4534 gnd.n1763 gnd.n989 240.244
R4535 gnd.n1763 gnd.n990 240.244
R4536 gnd.n990 gnd.n971 240.244
R4537 gnd.n1783 gnd.n971 240.244
R4538 gnd.n1783 gnd.n963 240.244
R4539 gnd.n1794 gnd.n963 240.244
R4540 gnd.n1794 gnd.n964 240.244
R4541 gnd.n964 gnd.n947 240.244
R4542 gnd.n1814 gnd.n947 240.244
R4543 gnd.n1814 gnd.n939 240.244
R4544 gnd.n1825 gnd.n939 240.244
R4545 gnd.n1825 gnd.n940 240.244
R4546 gnd.n940 gnd.n921 240.244
R4547 gnd.n1845 gnd.n921 240.244
R4548 gnd.n1845 gnd.n913 240.244
R4549 gnd.n1856 gnd.n913 240.244
R4550 gnd.n1856 gnd.n914 240.244
R4551 gnd.n914 gnd.n896 240.244
R4552 gnd.n2133 gnd.n896 240.244
R4553 gnd.n2133 gnd.n886 240.244
R4554 gnd.n2144 gnd.n886 240.244
R4555 gnd.n2144 gnd.n777 240.244
R4556 gnd.n5990 gnd.n777 240.244
R4557 gnd.n3456 gnd.n2475 240.244
R4558 gnd.n3458 gnd.n3457 240.244
R4559 gnd.n3468 gnd.n3467 240.244
R4560 gnd.n3476 gnd.n3475 240.244
R4561 gnd.n3478 gnd.n3477 240.244
R4562 gnd.n3488 gnd.n3487 240.244
R4563 gnd.n3496 gnd.n3495 240.244
R4564 gnd.n3498 gnd.n3497 240.244
R4565 gnd.n3512 gnd.n3508 240.244
R4566 gnd.n3727 gnd.n2270 240.244
R4567 gnd.n3732 gnd.n2270 240.244
R4568 gnd.n3732 gnd.n2280 240.244
R4569 gnd.n3735 gnd.n2280 240.244
R4570 gnd.n3735 gnd.n2290 240.244
R4571 gnd.n3740 gnd.n2290 240.244
R4572 gnd.n3740 gnd.n2299 240.244
R4573 gnd.n3743 gnd.n2299 240.244
R4574 gnd.n3743 gnd.n2308 240.244
R4575 gnd.n3748 gnd.n2308 240.244
R4576 gnd.n3748 gnd.n2318 240.244
R4577 gnd.n3751 gnd.n2318 240.244
R4578 gnd.n3751 gnd.n2327 240.244
R4579 gnd.n3756 gnd.n2327 240.244
R4580 gnd.n3756 gnd.n2337 240.244
R4581 gnd.n3759 gnd.n2337 240.244
R4582 gnd.n3759 gnd.n2346 240.244
R4583 gnd.n3764 gnd.n2346 240.244
R4584 gnd.n3764 gnd.n2356 240.244
R4585 gnd.n3767 gnd.n2356 240.244
R4586 gnd.n3767 gnd.n2365 240.244
R4587 gnd.n3660 gnd.n2365 240.244
R4588 gnd.n3660 gnd.n2375 240.244
R4589 gnd.n3774 gnd.n2375 240.244
R4590 gnd.n3774 gnd.n2384 240.244
R4591 gnd.n3657 gnd.n2384 240.244
R4592 gnd.n3657 gnd.n2395 240.244
R4593 gnd.n3831 gnd.n2395 240.244
R4594 gnd.n3831 gnd.n2404 240.244
R4595 gnd.n3837 gnd.n2404 240.244
R4596 gnd.n3837 gnd.n2415 240.244
R4597 gnd.n3882 gnd.n2415 240.244
R4598 gnd.n3882 gnd.n2424 240.244
R4599 gnd.n3647 gnd.n2424 240.244
R4600 gnd.n3647 gnd.n2435 240.244
R4601 gnd.n3648 gnd.n2435 240.244
R4602 gnd.n3648 gnd.n2445 240.244
R4603 gnd.n3651 gnd.n2445 240.244
R4604 gnd.n3651 gnd.n2456 240.244
R4605 gnd.n3864 gnd.n2456 240.244
R4606 gnd.n3864 gnd.n2466 240.244
R4607 gnd.n3925 gnd.n2466 240.244
R4608 gnd.n3688 gnd.n3687 240.244
R4609 gnd.n3694 gnd.n3693 240.244
R4610 gnd.n3698 gnd.n3697 240.244
R4611 gnd.n3704 gnd.n3703 240.244
R4612 gnd.n3708 gnd.n3707 240.244
R4613 gnd.n3714 gnd.n3713 240.244
R4614 gnd.n3718 gnd.n3717 240.244
R4615 gnd.n3677 gnd.n3676 240.244
R4616 gnd.n3672 gnd.n2192 240.244
R4617 gnd.n5806 gnd.n5805 240.244
R4618 gnd.n5805 gnd.n2266 240.244
R4619 gnd.n5795 gnd.n2266 240.244
R4620 gnd.n5795 gnd.n2282 240.244
R4621 gnd.n5791 gnd.n2282 240.244
R4622 gnd.n5791 gnd.n2288 240.244
R4623 gnd.n5783 gnd.n2288 240.244
R4624 gnd.n5783 gnd.n2301 240.244
R4625 gnd.n5779 gnd.n2301 240.244
R4626 gnd.n5779 gnd.n2306 240.244
R4627 gnd.n5771 gnd.n2306 240.244
R4628 gnd.n5771 gnd.n2319 240.244
R4629 gnd.n5767 gnd.n2319 240.244
R4630 gnd.n5767 gnd.n2324 240.244
R4631 gnd.n5759 gnd.n2324 240.244
R4632 gnd.n5759 gnd.n2339 240.244
R4633 gnd.n5755 gnd.n2339 240.244
R4634 gnd.n5755 gnd.n2344 240.244
R4635 gnd.n5747 gnd.n2344 240.244
R4636 gnd.n5747 gnd.n2357 240.244
R4637 gnd.n5743 gnd.n2357 240.244
R4638 gnd.n5743 gnd.n2362 240.244
R4639 gnd.n5735 gnd.n2362 240.244
R4640 gnd.n5735 gnd.n2377 240.244
R4641 gnd.n5731 gnd.n2377 240.244
R4642 gnd.n5731 gnd.n2382 240.244
R4643 gnd.n5723 gnd.n2382 240.244
R4644 gnd.n5723 gnd.n2396 240.244
R4645 gnd.n5719 gnd.n2396 240.244
R4646 gnd.n5719 gnd.n2401 240.244
R4647 gnd.n5711 gnd.n2401 240.244
R4648 gnd.n5711 gnd.n2417 240.244
R4649 gnd.n5707 gnd.n2417 240.244
R4650 gnd.n5707 gnd.n2422 240.244
R4651 gnd.n5699 gnd.n2422 240.244
R4652 gnd.n5699 gnd.n2437 240.244
R4653 gnd.n5695 gnd.n2437 240.244
R4654 gnd.n5695 gnd.n2442 240.244
R4655 gnd.n5687 gnd.n2442 240.244
R4656 gnd.n5687 gnd.n2458 240.244
R4657 gnd.n5683 gnd.n2458 240.244
R4658 gnd.n5683 gnd.n2463 240.244
R4659 gnd.n6169 gnd.n591 240.244
R4660 gnd.n6175 gnd.n591 240.244
R4661 gnd.n6175 gnd.n589 240.244
R4662 gnd.n6179 gnd.n589 240.244
R4663 gnd.n6179 gnd.n585 240.244
R4664 gnd.n6185 gnd.n585 240.244
R4665 gnd.n6185 gnd.n583 240.244
R4666 gnd.n6189 gnd.n583 240.244
R4667 gnd.n6189 gnd.n579 240.244
R4668 gnd.n6195 gnd.n579 240.244
R4669 gnd.n6195 gnd.n577 240.244
R4670 gnd.n6199 gnd.n577 240.244
R4671 gnd.n6199 gnd.n573 240.244
R4672 gnd.n6205 gnd.n573 240.244
R4673 gnd.n6205 gnd.n571 240.244
R4674 gnd.n6209 gnd.n571 240.244
R4675 gnd.n6209 gnd.n567 240.244
R4676 gnd.n6215 gnd.n567 240.244
R4677 gnd.n6215 gnd.n565 240.244
R4678 gnd.n6219 gnd.n565 240.244
R4679 gnd.n6219 gnd.n561 240.244
R4680 gnd.n6225 gnd.n561 240.244
R4681 gnd.n6225 gnd.n559 240.244
R4682 gnd.n6229 gnd.n559 240.244
R4683 gnd.n6229 gnd.n555 240.244
R4684 gnd.n6235 gnd.n555 240.244
R4685 gnd.n6235 gnd.n553 240.244
R4686 gnd.n6239 gnd.n553 240.244
R4687 gnd.n6239 gnd.n549 240.244
R4688 gnd.n6245 gnd.n549 240.244
R4689 gnd.n6245 gnd.n547 240.244
R4690 gnd.n6249 gnd.n547 240.244
R4691 gnd.n6249 gnd.n543 240.244
R4692 gnd.n6255 gnd.n543 240.244
R4693 gnd.n6255 gnd.n541 240.244
R4694 gnd.n6259 gnd.n541 240.244
R4695 gnd.n6259 gnd.n537 240.244
R4696 gnd.n6265 gnd.n537 240.244
R4697 gnd.n6265 gnd.n535 240.244
R4698 gnd.n6269 gnd.n535 240.244
R4699 gnd.n6269 gnd.n531 240.244
R4700 gnd.n6275 gnd.n531 240.244
R4701 gnd.n6275 gnd.n529 240.244
R4702 gnd.n6279 gnd.n529 240.244
R4703 gnd.n6279 gnd.n525 240.244
R4704 gnd.n6285 gnd.n525 240.244
R4705 gnd.n6285 gnd.n523 240.244
R4706 gnd.n6289 gnd.n523 240.244
R4707 gnd.n6289 gnd.n519 240.244
R4708 gnd.n6295 gnd.n519 240.244
R4709 gnd.n6295 gnd.n517 240.244
R4710 gnd.n6299 gnd.n517 240.244
R4711 gnd.n6299 gnd.n513 240.244
R4712 gnd.n6305 gnd.n513 240.244
R4713 gnd.n6305 gnd.n511 240.244
R4714 gnd.n6309 gnd.n511 240.244
R4715 gnd.n6309 gnd.n507 240.244
R4716 gnd.n6315 gnd.n507 240.244
R4717 gnd.n6315 gnd.n505 240.244
R4718 gnd.n6319 gnd.n505 240.244
R4719 gnd.n6319 gnd.n501 240.244
R4720 gnd.n6325 gnd.n501 240.244
R4721 gnd.n6325 gnd.n499 240.244
R4722 gnd.n6329 gnd.n499 240.244
R4723 gnd.n6329 gnd.n495 240.244
R4724 gnd.n6335 gnd.n495 240.244
R4725 gnd.n6335 gnd.n493 240.244
R4726 gnd.n6339 gnd.n493 240.244
R4727 gnd.n6339 gnd.n489 240.244
R4728 gnd.n6345 gnd.n489 240.244
R4729 gnd.n6345 gnd.n487 240.244
R4730 gnd.n6349 gnd.n487 240.244
R4731 gnd.n6349 gnd.n483 240.244
R4732 gnd.n6355 gnd.n483 240.244
R4733 gnd.n6355 gnd.n481 240.244
R4734 gnd.n6359 gnd.n481 240.244
R4735 gnd.n6359 gnd.n477 240.244
R4736 gnd.n6365 gnd.n477 240.244
R4737 gnd.n6365 gnd.n475 240.244
R4738 gnd.n6369 gnd.n475 240.244
R4739 gnd.n6369 gnd.n471 240.244
R4740 gnd.n6375 gnd.n471 240.244
R4741 gnd.n6375 gnd.n469 240.244
R4742 gnd.n6379 gnd.n469 240.244
R4743 gnd.n6379 gnd.n465 240.244
R4744 gnd.n6385 gnd.n465 240.244
R4745 gnd.n6385 gnd.n463 240.244
R4746 gnd.n6389 gnd.n463 240.244
R4747 gnd.n6389 gnd.n459 240.244
R4748 gnd.n6395 gnd.n459 240.244
R4749 gnd.n6395 gnd.n457 240.244
R4750 gnd.n6399 gnd.n457 240.244
R4751 gnd.n6399 gnd.n453 240.244
R4752 gnd.n6405 gnd.n453 240.244
R4753 gnd.n6405 gnd.n451 240.244
R4754 gnd.n6409 gnd.n451 240.244
R4755 gnd.n6409 gnd.n447 240.244
R4756 gnd.n6415 gnd.n447 240.244
R4757 gnd.n6415 gnd.n445 240.244
R4758 gnd.n6419 gnd.n445 240.244
R4759 gnd.n6419 gnd.n441 240.244
R4760 gnd.n6425 gnd.n441 240.244
R4761 gnd.n6425 gnd.n439 240.244
R4762 gnd.n6429 gnd.n439 240.244
R4763 gnd.n6429 gnd.n435 240.244
R4764 gnd.n6435 gnd.n435 240.244
R4765 gnd.n6435 gnd.n433 240.244
R4766 gnd.n6439 gnd.n433 240.244
R4767 gnd.n6439 gnd.n429 240.244
R4768 gnd.n6445 gnd.n429 240.244
R4769 gnd.n6445 gnd.n427 240.244
R4770 gnd.n6449 gnd.n427 240.244
R4771 gnd.n6449 gnd.n423 240.244
R4772 gnd.n6455 gnd.n423 240.244
R4773 gnd.n6455 gnd.n421 240.244
R4774 gnd.n6459 gnd.n421 240.244
R4775 gnd.n6459 gnd.n417 240.244
R4776 gnd.n6465 gnd.n417 240.244
R4777 gnd.n6465 gnd.n415 240.244
R4778 gnd.n6469 gnd.n415 240.244
R4779 gnd.n6469 gnd.n411 240.244
R4780 gnd.n6475 gnd.n411 240.244
R4781 gnd.n6475 gnd.n409 240.244
R4782 gnd.n6479 gnd.n409 240.244
R4783 gnd.n6479 gnd.n405 240.244
R4784 gnd.n6485 gnd.n405 240.244
R4785 gnd.n6485 gnd.n403 240.244
R4786 gnd.n6489 gnd.n403 240.244
R4787 gnd.n6489 gnd.n399 240.244
R4788 gnd.n6495 gnd.n399 240.244
R4789 gnd.n6495 gnd.n397 240.244
R4790 gnd.n6499 gnd.n397 240.244
R4791 gnd.n6499 gnd.n393 240.244
R4792 gnd.n6505 gnd.n393 240.244
R4793 gnd.n6505 gnd.n391 240.244
R4794 gnd.n6509 gnd.n391 240.244
R4795 gnd.n6509 gnd.n387 240.244
R4796 gnd.n6516 gnd.n387 240.244
R4797 gnd.n6516 gnd.n385 240.244
R4798 gnd.n6520 gnd.n385 240.244
R4799 gnd.n6520 gnd.n382 240.244
R4800 gnd.n6526 gnd.n380 240.244
R4801 gnd.n6530 gnd.n380 240.244
R4802 gnd.n6530 gnd.n376 240.244
R4803 gnd.n6536 gnd.n376 240.244
R4804 gnd.n6536 gnd.n374 240.244
R4805 gnd.n6540 gnd.n374 240.244
R4806 gnd.n6540 gnd.n370 240.244
R4807 gnd.n6546 gnd.n370 240.244
R4808 gnd.n6546 gnd.n368 240.244
R4809 gnd.n6550 gnd.n368 240.244
R4810 gnd.n6550 gnd.n364 240.244
R4811 gnd.n6556 gnd.n364 240.244
R4812 gnd.n6556 gnd.n362 240.244
R4813 gnd.n6560 gnd.n362 240.244
R4814 gnd.n6560 gnd.n358 240.244
R4815 gnd.n6566 gnd.n358 240.244
R4816 gnd.n6566 gnd.n356 240.244
R4817 gnd.n6570 gnd.n356 240.244
R4818 gnd.n6570 gnd.n352 240.244
R4819 gnd.n6576 gnd.n352 240.244
R4820 gnd.n6576 gnd.n350 240.244
R4821 gnd.n6580 gnd.n350 240.244
R4822 gnd.n6580 gnd.n346 240.244
R4823 gnd.n6586 gnd.n346 240.244
R4824 gnd.n6586 gnd.n344 240.244
R4825 gnd.n6590 gnd.n344 240.244
R4826 gnd.n6590 gnd.n340 240.244
R4827 gnd.n6596 gnd.n340 240.244
R4828 gnd.n6596 gnd.n338 240.244
R4829 gnd.n6600 gnd.n338 240.244
R4830 gnd.n6600 gnd.n334 240.244
R4831 gnd.n6606 gnd.n334 240.244
R4832 gnd.n6606 gnd.n332 240.244
R4833 gnd.n6610 gnd.n332 240.244
R4834 gnd.n6610 gnd.n328 240.244
R4835 gnd.n6616 gnd.n328 240.244
R4836 gnd.n6616 gnd.n326 240.244
R4837 gnd.n6620 gnd.n326 240.244
R4838 gnd.n6620 gnd.n322 240.244
R4839 gnd.n6626 gnd.n322 240.244
R4840 gnd.n6626 gnd.n320 240.244
R4841 gnd.n6630 gnd.n320 240.244
R4842 gnd.n6630 gnd.n316 240.244
R4843 gnd.n6636 gnd.n316 240.244
R4844 gnd.n6636 gnd.n314 240.244
R4845 gnd.n6640 gnd.n314 240.244
R4846 gnd.n6640 gnd.n310 240.244
R4847 gnd.n6646 gnd.n310 240.244
R4848 gnd.n6646 gnd.n308 240.244
R4849 gnd.n6650 gnd.n308 240.244
R4850 gnd.n6650 gnd.n304 240.244
R4851 gnd.n6656 gnd.n304 240.244
R4852 gnd.n6656 gnd.n302 240.244
R4853 gnd.n6660 gnd.n302 240.244
R4854 gnd.n6660 gnd.n298 240.244
R4855 gnd.n6666 gnd.n298 240.244
R4856 gnd.n6666 gnd.n296 240.244
R4857 gnd.n6670 gnd.n296 240.244
R4858 gnd.n6670 gnd.n292 240.244
R4859 gnd.n6676 gnd.n292 240.244
R4860 gnd.n6676 gnd.n290 240.244
R4861 gnd.n6680 gnd.n290 240.244
R4862 gnd.n6680 gnd.n286 240.244
R4863 gnd.n6686 gnd.n286 240.244
R4864 gnd.n6686 gnd.n284 240.244
R4865 gnd.n6690 gnd.n284 240.244
R4866 gnd.n6690 gnd.n280 240.244
R4867 gnd.n6696 gnd.n280 240.244
R4868 gnd.n6696 gnd.n278 240.244
R4869 gnd.n6700 gnd.n278 240.244
R4870 gnd.n6700 gnd.n274 240.244
R4871 gnd.n6706 gnd.n274 240.244
R4872 gnd.n6706 gnd.n272 240.244
R4873 gnd.n6710 gnd.n272 240.244
R4874 gnd.n6710 gnd.n268 240.244
R4875 gnd.n6716 gnd.n268 240.244
R4876 gnd.n6716 gnd.n266 240.244
R4877 gnd.n6720 gnd.n266 240.244
R4878 gnd.n6720 gnd.n262 240.244
R4879 gnd.n6726 gnd.n262 240.244
R4880 gnd.n6726 gnd.n260 240.244
R4881 gnd.n6731 gnd.n260 240.244
R4882 gnd.n6731 gnd.n256 240.244
R4883 gnd.n6737 gnd.n256 240.244
R4884 gnd.n3634 gnd.n3631 240.244
R4885 gnd.n3640 gnd.n3631 240.244
R4886 gnd.n3641 gnd.n3640 240.244
R4887 gnd.n3885 gnd.n3641 240.244
R4888 gnd.n3885 gnd.n3627 240.244
R4889 gnd.n3891 gnd.n3627 240.244
R4890 gnd.n3892 gnd.n3891 240.244
R4891 gnd.n3893 gnd.n3892 240.244
R4892 gnd.n3893 gnd.n3623 240.244
R4893 gnd.n3899 gnd.n3623 240.244
R4894 gnd.n3900 gnd.n3899 240.244
R4895 gnd.n3901 gnd.n3900 240.244
R4896 gnd.n3901 gnd.n3618 240.244
R4897 gnd.n3922 gnd.n3618 240.244
R4898 gnd.n3922 gnd.n3619 240.244
R4899 gnd.n3918 gnd.n3619 240.244
R4900 gnd.n3918 gnd.n3917 240.244
R4901 gnd.n3917 gnd.n3915 240.244
R4902 gnd.n3915 gnd.n3909 240.244
R4903 gnd.n3909 gnd.n3390 240.244
R4904 gnd.n3999 gnd.n3390 240.244
R4905 gnd.n3999 gnd.n3386 240.244
R4906 gnd.n4005 gnd.n3386 240.244
R4907 gnd.n4005 gnd.n3375 240.244
R4908 gnd.n4015 gnd.n3375 240.244
R4909 gnd.n4015 gnd.n3371 240.244
R4910 gnd.n4021 gnd.n3371 240.244
R4911 gnd.n4021 gnd.n3360 240.244
R4912 gnd.n4043 gnd.n3360 240.244
R4913 gnd.n4043 gnd.n3355 240.244
R4914 gnd.n4052 gnd.n3355 240.244
R4915 gnd.n4052 gnd.n3356 240.244
R4916 gnd.n3356 gnd.n2609 240.244
R4917 gnd.n5548 gnd.n2609 240.244
R4918 gnd.n5548 gnd.n2610 240.244
R4919 gnd.n5544 gnd.n2610 240.244
R4920 gnd.n5544 gnd.n2616 240.244
R4921 gnd.n3337 gnd.n2616 240.244
R4922 gnd.n3337 gnd.n3319 240.244
R4923 gnd.n4192 gnd.n3319 240.244
R4924 gnd.n4192 gnd.n3314 240.244
R4925 gnd.n4203 gnd.n3314 240.244
R4926 gnd.n4203 gnd.n3315 240.244
R4927 gnd.n4199 gnd.n3315 240.244
R4928 gnd.n4199 gnd.n3289 240.244
R4929 gnd.n4261 gnd.n3289 240.244
R4930 gnd.n4261 gnd.n3285 240.244
R4931 gnd.n4267 gnd.n3285 240.244
R4932 gnd.n4267 gnd.n3272 240.244
R4933 gnd.n4290 gnd.n3272 240.244
R4934 gnd.n4290 gnd.n3267 240.244
R4935 gnd.n4298 gnd.n3267 240.244
R4936 gnd.n4298 gnd.n3268 240.244
R4937 gnd.n3268 gnd.n3244 240.244
R4938 gnd.n4364 gnd.n3244 240.244
R4939 gnd.n4364 gnd.n3239 240.244
R4940 gnd.n4372 gnd.n3239 240.244
R4941 gnd.n4372 gnd.n3240 240.244
R4942 gnd.n3240 gnd.n3221 240.244
R4943 gnd.n4396 gnd.n3221 240.244
R4944 gnd.n4396 gnd.n3216 240.244
R4945 gnd.n4404 gnd.n3216 240.244
R4946 gnd.n4404 gnd.n3217 240.244
R4947 gnd.n3217 gnd.n3200 240.244
R4948 gnd.n4437 gnd.n3200 240.244
R4949 gnd.n4437 gnd.n3195 240.244
R4950 gnd.n4445 gnd.n3195 240.244
R4951 gnd.n4445 gnd.n3196 240.244
R4952 gnd.n3196 gnd.n3171 240.244
R4953 gnd.n4506 gnd.n3171 240.244
R4954 gnd.n4506 gnd.n3164 240.244
R4955 gnd.n4514 gnd.n3164 240.244
R4956 gnd.n4514 gnd.n3167 240.244
R4957 gnd.n3167 gnd.n3146 240.244
R4958 gnd.n4538 gnd.n3146 240.244
R4959 gnd.n4538 gnd.n3141 240.244
R4960 gnd.n4546 gnd.n3141 240.244
R4961 gnd.n4546 gnd.n3142 240.244
R4962 gnd.n3142 gnd.n3123 240.244
R4963 gnd.n4578 gnd.n3123 240.244
R4964 gnd.n4578 gnd.n3118 240.244
R4965 gnd.n4586 gnd.n3118 240.244
R4966 gnd.n4586 gnd.n3119 240.244
R4967 gnd.n3119 gnd.n3094 240.244
R4968 gnd.n4632 gnd.n3094 240.244
R4969 gnd.n4632 gnd.n3088 240.244
R4970 gnd.n4640 gnd.n3088 240.244
R4971 gnd.n4640 gnd.n3090 240.244
R4972 gnd.n3090 gnd.n3070 240.244
R4973 gnd.n4674 gnd.n3070 240.244
R4974 gnd.n4674 gnd.n3065 240.244
R4975 gnd.n4682 gnd.n3065 240.244
R4976 gnd.n4682 gnd.n3066 240.244
R4977 gnd.n3066 gnd.n3042 240.244
R4978 gnd.n4717 gnd.n3042 240.244
R4979 gnd.n4717 gnd.n3038 240.244
R4980 gnd.n4724 gnd.n3038 240.244
R4981 gnd.n4724 gnd.n3016 240.244
R4982 gnd.n4764 gnd.n3016 240.244
R4983 gnd.n4764 gnd.n3017 240.244
R4984 gnd.n4760 gnd.n3017 240.244
R4985 gnd.n4760 gnd.n4759 240.244
R4986 gnd.n4759 gnd.n4758 240.244
R4987 gnd.n4758 gnd.n2988 240.244
R4988 gnd.n4809 gnd.n2988 240.244
R4989 gnd.n4809 gnd.n2984 240.244
R4990 gnd.n4815 gnd.n2984 240.244
R4991 gnd.n4815 gnd.n2936 240.244
R4992 gnd.n4981 gnd.n2936 240.244
R4993 gnd.n4981 gnd.n2932 240.244
R4994 gnd.n4987 gnd.n2932 240.244
R4995 gnd.n4987 gnd.n2924 240.244
R4996 gnd.n4999 gnd.n2924 240.244
R4997 gnd.n4999 gnd.n2920 240.244
R4998 gnd.n5005 gnd.n2920 240.244
R4999 gnd.n5005 gnd.n2913 240.244
R5000 gnd.n5016 gnd.n2913 240.244
R5001 gnd.n5016 gnd.n2909 240.244
R5002 gnd.n5024 gnd.n2909 240.244
R5003 gnd.n5024 gnd.n2900 240.244
R5004 gnd.n5052 gnd.n2900 240.244
R5005 gnd.n5053 gnd.n5052 240.244
R5006 gnd.n5053 gnd.n2896 240.244
R5007 gnd.n5060 gnd.n2896 240.244
R5008 gnd.n5061 gnd.n5060 240.244
R5009 gnd.n5062 gnd.n5061 240.244
R5010 gnd.n5062 gnd.n2891 240.244
R5011 gnd.n5190 gnd.n2891 240.244
R5012 gnd.n5190 gnd.n2892 240.244
R5013 gnd.n5186 gnd.n2892 240.244
R5014 gnd.n5186 gnd.n5070 240.244
R5015 gnd.n5111 gnd.n5070 240.244
R5016 gnd.n5111 gnd.n5107 240.244
R5017 gnd.n5126 gnd.n5107 240.244
R5018 gnd.n5126 gnd.n5108 240.244
R5019 gnd.n5122 gnd.n5108 240.244
R5020 gnd.n5122 gnd.n5121 240.244
R5021 gnd.n5121 gnd.n250 240.244
R5022 gnd.n6742 gnd.n250 240.244
R5023 gnd.n6742 gnd.n251 240.244
R5024 gnd.n6738 gnd.n251 240.244
R5025 gnd.n6165 gnd.n594 240.244
R5026 gnd.n6165 gnd.n596 240.244
R5027 gnd.n6161 gnd.n596 240.244
R5028 gnd.n6161 gnd.n602 240.244
R5029 gnd.n6157 gnd.n602 240.244
R5030 gnd.n6157 gnd.n604 240.244
R5031 gnd.n6153 gnd.n604 240.244
R5032 gnd.n6153 gnd.n610 240.244
R5033 gnd.n6149 gnd.n610 240.244
R5034 gnd.n6149 gnd.n612 240.244
R5035 gnd.n6145 gnd.n612 240.244
R5036 gnd.n6145 gnd.n618 240.244
R5037 gnd.n6141 gnd.n618 240.244
R5038 gnd.n6141 gnd.n620 240.244
R5039 gnd.n6137 gnd.n620 240.244
R5040 gnd.n6137 gnd.n626 240.244
R5041 gnd.n6133 gnd.n626 240.244
R5042 gnd.n6133 gnd.n628 240.244
R5043 gnd.n6129 gnd.n628 240.244
R5044 gnd.n6129 gnd.n634 240.244
R5045 gnd.n6125 gnd.n634 240.244
R5046 gnd.n6125 gnd.n636 240.244
R5047 gnd.n6121 gnd.n636 240.244
R5048 gnd.n6121 gnd.n642 240.244
R5049 gnd.n6117 gnd.n642 240.244
R5050 gnd.n6117 gnd.n644 240.244
R5051 gnd.n6113 gnd.n644 240.244
R5052 gnd.n6113 gnd.n650 240.244
R5053 gnd.n6109 gnd.n650 240.244
R5054 gnd.n6109 gnd.n652 240.244
R5055 gnd.n6105 gnd.n652 240.244
R5056 gnd.n6105 gnd.n658 240.244
R5057 gnd.n6101 gnd.n658 240.244
R5058 gnd.n6101 gnd.n660 240.244
R5059 gnd.n6097 gnd.n660 240.244
R5060 gnd.n6097 gnd.n666 240.244
R5061 gnd.n6093 gnd.n666 240.244
R5062 gnd.n6093 gnd.n668 240.244
R5063 gnd.n6089 gnd.n668 240.244
R5064 gnd.n6089 gnd.n674 240.244
R5065 gnd.n6085 gnd.n674 240.244
R5066 gnd.n6085 gnd.n676 240.244
R5067 gnd.n6081 gnd.n676 240.244
R5068 gnd.n6081 gnd.n682 240.244
R5069 gnd.n6077 gnd.n682 240.244
R5070 gnd.n6077 gnd.n684 240.244
R5071 gnd.n6073 gnd.n684 240.244
R5072 gnd.n6073 gnd.n690 240.244
R5073 gnd.n6069 gnd.n690 240.244
R5074 gnd.n6069 gnd.n692 240.244
R5075 gnd.n6065 gnd.n692 240.244
R5076 gnd.n6065 gnd.n698 240.244
R5077 gnd.n6061 gnd.n698 240.244
R5078 gnd.n6061 gnd.n700 240.244
R5079 gnd.n6057 gnd.n700 240.244
R5080 gnd.n6057 gnd.n706 240.244
R5081 gnd.n6053 gnd.n706 240.244
R5082 gnd.n6053 gnd.n708 240.244
R5083 gnd.n6049 gnd.n708 240.244
R5084 gnd.n6049 gnd.n714 240.244
R5085 gnd.n6045 gnd.n714 240.244
R5086 gnd.n6045 gnd.n716 240.244
R5087 gnd.n6041 gnd.n716 240.244
R5088 gnd.n6041 gnd.n722 240.244
R5089 gnd.n6037 gnd.n722 240.244
R5090 gnd.n6037 gnd.n724 240.244
R5091 gnd.n6033 gnd.n724 240.244
R5092 gnd.n6033 gnd.n730 240.244
R5093 gnd.n6029 gnd.n730 240.244
R5094 gnd.n6029 gnd.n732 240.244
R5095 gnd.n6025 gnd.n732 240.244
R5096 gnd.n6025 gnd.n738 240.244
R5097 gnd.n6021 gnd.n738 240.244
R5098 gnd.n6021 gnd.n740 240.244
R5099 gnd.n6017 gnd.n740 240.244
R5100 gnd.n6017 gnd.n746 240.244
R5101 gnd.n6013 gnd.n746 240.244
R5102 gnd.n6013 gnd.n748 240.244
R5103 gnd.n6009 gnd.n748 240.244
R5104 gnd.n6009 gnd.n754 240.244
R5105 gnd.n6005 gnd.n754 240.244
R5106 gnd.n6005 gnd.n756 240.244
R5107 gnd.n6001 gnd.n756 240.244
R5108 gnd.n6001 gnd.n762 240.244
R5109 gnd.n3414 gnd.n3392 240.244
R5110 gnd.n3416 gnd.n3392 240.244
R5111 gnd.n3416 gnd.n3385 240.244
R5112 gnd.n3419 gnd.n3385 240.244
R5113 gnd.n3419 gnd.n3377 240.244
R5114 gnd.n3420 gnd.n3377 240.244
R5115 gnd.n3420 gnd.n3370 240.244
R5116 gnd.n3423 gnd.n3370 240.244
R5117 gnd.n3423 gnd.n3362 240.244
R5118 gnd.n3362 gnd.n3351 240.244
R5119 gnd.n4054 gnd.n3351 240.244
R5120 gnd.n4054 gnd.n3352 240.244
R5121 gnd.n3352 gnd.n3348 240.244
R5122 gnd.n3348 gnd.n2607 240.244
R5123 gnd.n4142 gnd.n2607 240.244
R5124 gnd.n4142 gnd.n2617 240.244
R5125 gnd.n4162 gnd.n2617 240.244
R5126 gnd.n4162 gnd.n3343 240.244
R5127 gnd.n4147 gnd.n3343 240.244
R5128 gnd.n4147 gnd.n3321 240.244
R5129 gnd.n4148 gnd.n3321 240.244
R5130 gnd.n4148 gnd.n3312 240.244
R5131 gnd.n4150 gnd.n3312 240.244
R5132 gnd.n4150 gnd.n3299 240.244
R5133 gnd.n4247 gnd.n3299 240.244
R5134 gnd.n4247 gnd.n3291 240.244
R5135 gnd.n4223 gnd.n3291 240.244
R5136 gnd.n4223 gnd.n3284 240.244
R5137 gnd.n3284 gnd.n3280 240.244
R5138 gnd.n3280 gnd.n3273 240.244
R5139 gnd.n4226 gnd.n3273 240.244
R5140 gnd.n4226 gnd.n3266 240.244
R5141 gnd.n4227 gnd.n3266 240.244
R5142 gnd.n4228 gnd.n4227 240.244
R5143 gnd.n4228 gnd.n3246 240.244
R5144 gnd.n3246 gnd.n3235 240.244
R5145 gnd.n4374 gnd.n3235 240.244
R5146 gnd.n4374 gnd.n3230 240.244
R5147 gnd.n4381 gnd.n3230 240.244
R5148 gnd.n4381 gnd.n3223 240.244
R5149 gnd.n3223 gnd.n3213 240.244
R5150 gnd.n4406 gnd.n3213 240.244
R5151 gnd.n4406 gnd.n3208 240.244
R5152 gnd.n4426 gnd.n3208 240.244
R5153 gnd.n4426 gnd.n3202 240.244
R5154 gnd.n4411 gnd.n3202 240.244
R5155 gnd.n4411 gnd.n3194 240.244
R5156 gnd.n4412 gnd.n3194 240.244
R5157 gnd.n4413 gnd.n4412 240.244
R5158 gnd.n4413 gnd.n3173 240.244
R5159 gnd.n3173 gnd.n3161 240.244
R5160 gnd.n4516 gnd.n3161 240.244
R5161 gnd.n4516 gnd.n3156 240.244
R5162 gnd.n4523 gnd.n3156 240.244
R5163 gnd.n4523 gnd.n3148 240.244
R5164 gnd.n3148 gnd.n3137 240.244
R5165 gnd.n4548 gnd.n3137 240.244
R5166 gnd.n4548 gnd.n3132 240.244
R5167 gnd.n4568 gnd.n3132 240.244
R5168 gnd.n4568 gnd.n3125 240.244
R5169 gnd.n4553 gnd.n3125 240.244
R5170 gnd.n4553 gnd.n3116 240.244
R5171 gnd.n4554 gnd.n3116 240.244
R5172 gnd.n4555 gnd.n4554 240.244
R5173 gnd.n4555 gnd.n3096 240.244
R5174 gnd.n3096 gnd.n3085 240.244
R5175 gnd.n4642 gnd.n3085 240.244
R5176 gnd.n4642 gnd.n3080 240.244
R5177 gnd.n4663 gnd.n3080 240.244
R5178 gnd.n4663 gnd.n3072 240.244
R5179 gnd.n4648 gnd.n3072 240.244
R5180 gnd.n4648 gnd.n3063 240.244
R5181 gnd.n4649 gnd.n3063 240.244
R5182 gnd.n4650 gnd.n4649 240.244
R5183 gnd.n4650 gnd.n3044 240.244
R5184 gnd.n3044 gnd.n3033 240.244
R5185 gnd.n4726 gnd.n3033 240.244
R5186 gnd.n4726 gnd.n3034 240.244
R5187 gnd.n3034 gnd.n3015 240.244
R5188 gnd.n4735 gnd.n3015 240.244
R5189 gnd.n4736 gnd.n4735 240.244
R5190 gnd.n4736 gnd.n3026 240.244
R5191 gnd.n4756 gnd.n3026 240.244
R5192 gnd.n4756 gnd.n2997 240.244
R5193 gnd.n2997 gnd.n2989 240.244
R5194 gnd.n4742 gnd.n2989 240.244
R5195 gnd.n4742 gnd.n2982 240.244
R5196 gnd.n4743 gnd.n2982 240.244
R5197 gnd.n4743 gnd.n2938 240.244
R5198 gnd.n2938 gnd.n2930 240.244
R5199 gnd.n4989 gnd.n2930 240.244
R5200 gnd.n4989 gnd.n2926 240.244
R5201 gnd.n4995 gnd.n2926 240.244
R5202 gnd.n4995 gnd.n2919 240.244
R5203 gnd.n5007 gnd.n2919 240.244
R5204 gnd.n5007 gnd.n2915 240.244
R5205 gnd.n5013 gnd.n2915 240.244
R5206 gnd.n5013 gnd.n2907 240.244
R5207 gnd.n5026 gnd.n2907 240.244
R5208 gnd.n5026 gnd.n2902 240.244
R5209 gnd.n5050 gnd.n2902 240.244
R5210 gnd.n3413 gnd.n3412 240.244
R5211 gnd.n3442 gnd.n3412 240.244
R5212 gnd.n3444 gnd.n3443 240.244
R5213 gnd.n3449 gnd.n3448 240.244
R5214 gnd.n3451 gnd.n3450 240.244
R5215 gnd.n3462 gnd.n3461 240.244
R5216 gnd.n3464 gnd.n3463 240.244
R5217 gnd.n3472 gnd.n3471 240.244
R5218 gnd.n3482 gnd.n3481 240.244
R5219 gnd.n3484 gnd.n3483 240.244
R5220 gnd.n3492 gnd.n3491 240.244
R5221 gnd.n3502 gnd.n3501 240.244
R5222 gnd.n3513 gnd.n3503 240.244
R5223 gnd.n3515 gnd.n3397 240.244
R5224 gnd.n3997 gnd.n3393 240.244
R5225 gnd.n3997 gnd.n3383 240.244
R5226 gnd.n4007 gnd.n3383 240.244
R5227 gnd.n4007 gnd.n3379 240.244
R5228 gnd.n4013 gnd.n3379 240.244
R5229 gnd.n4013 gnd.n3369 240.244
R5230 gnd.n4023 gnd.n3369 240.244
R5231 gnd.n4023 gnd.n3363 240.244
R5232 gnd.n4041 gnd.n3363 240.244
R5233 gnd.n4041 gnd.n3364 240.244
R5234 gnd.n3364 gnd.n3354 240.244
R5235 gnd.n4028 gnd.n3354 240.244
R5236 gnd.n4030 gnd.n4028 240.244
R5237 gnd.n4030 gnd.n2608 240.244
R5238 gnd.n2618 gnd.n2608 240.244
R5239 gnd.n5542 gnd.n2618 240.244
R5240 gnd.n5542 gnd.n2619 240.244
R5241 gnd.n2624 gnd.n2619 240.244
R5242 gnd.n2625 gnd.n2624 240.244
R5243 gnd.n2626 gnd.n2625 240.244
R5244 gnd.n3323 gnd.n2626 240.244
R5245 gnd.n3323 gnd.n2629 240.244
R5246 gnd.n2630 gnd.n2629 240.244
R5247 gnd.n2631 gnd.n2630 240.244
R5248 gnd.n4248 gnd.n2631 240.244
R5249 gnd.n4248 gnd.n2634 240.244
R5250 gnd.n2635 gnd.n2634 240.244
R5251 gnd.n2636 gnd.n2635 240.244
R5252 gnd.n4280 gnd.n2636 240.244
R5253 gnd.n4280 gnd.n2639 240.244
R5254 gnd.n2640 gnd.n2639 240.244
R5255 gnd.n2641 gnd.n2640 240.244
R5256 gnd.n3259 gnd.n2641 240.244
R5257 gnd.n3259 gnd.n2644 240.244
R5258 gnd.n2645 gnd.n2644 240.244
R5259 gnd.n2646 gnd.n2645 240.244
R5260 gnd.n3238 gnd.n2646 240.244
R5261 gnd.n3238 gnd.n2649 240.244
R5262 gnd.n2650 gnd.n2649 240.244
R5263 gnd.n2651 gnd.n2650 240.244
R5264 gnd.n4330 gnd.n2651 240.244
R5265 gnd.n4330 gnd.n2654 240.244
R5266 gnd.n2655 gnd.n2654 240.244
R5267 gnd.n2656 gnd.n2655 240.244
R5268 gnd.n4435 gnd.n2656 240.244
R5269 gnd.n4435 gnd.n2659 240.244
R5270 gnd.n2660 gnd.n2659 240.244
R5271 gnd.n2661 gnd.n2660 240.244
R5272 gnd.n3180 gnd.n2661 240.244
R5273 gnd.n3180 gnd.n2664 240.244
R5274 gnd.n2665 gnd.n2664 240.244
R5275 gnd.n2666 gnd.n2665 240.244
R5276 gnd.n3165 gnd.n2666 240.244
R5277 gnd.n3165 gnd.n2669 240.244
R5278 gnd.n2670 gnd.n2669 240.244
R5279 gnd.n2671 gnd.n2670 240.244
R5280 gnd.n3140 gnd.n2671 240.244
R5281 gnd.n3140 gnd.n2674 240.244
R5282 gnd.n2675 gnd.n2674 240.244
R5283 gnd.n2676 gnd.n2675 240.244
R5284 gnd.n3113 gnd.n2676 240.244
R5285 gnd.n3113 gnd.n2679 240.244
R5286 gnd.n2680 gnd.n2679 240.244
R5287 gnd.n2681 gnd.n2680 240.244
R5288 gnd.n4630 gnd.n2681 240.244
R5289 gnd.n4630 gnd.n2684 240.244
R5290 gnd.n2685 gnd.n2684 240.244
R5291 gnd.n2686 gnd.n2685 240.244
R5292 gnd.n4664 gnd.n2686 240.244
R5293 gnd.n4664 gnd.n2689 240.244
R5294 gnd.n2690 gnd.n2689 240.244
R5295 gnd.n2691 gnd.n2690 240.244
R5296 gnd.n3057 gnd.n2691 240.244
R5297 gnd.n3057 gnd.n2694 240.244
R5298 gnd.n2695 gnd.n2694 240.244
R5299 gnd.n2696 gnd.n2695 240.244
R5300 gnd.n3037 gnd.n2696 240.244
R5301 gnd.n3037 gnd.n2699 240.244
R5302 gnd.n2700 gnd.n2699 240.244
R5303 gnd.n2701 gnd.n2700 240.244
R5304 gnd.n3004 gnd.n2701 240.244
R5305 gnd.n3004 gnd.n2704 240.244
R5306 gnd.n2705 gnd.n2704 240.244
R5307 gnd.n2706 gnd.n2705 240.244
R5308 gnd.n4807 gnd.n2706 240.244
R5309 gnd.n4807 gnd.n2709 240.244
R5310 gnd.n2710 gnd.n2709 240.244
R5311 gnd.n2711 gnd.n2710 240.244
R5312 gnd.n4979 gnd.n2711 240.244
R5313 gnd.n4979 gnd.n2714 240.244
R5314 gnd.n2715 gnd.n2714 240.244
R5315 gnd.n2716 gnd.n2715 240.244
R5316 gnd.n4997 gnd.n2716 240.244
R5317 gnd.n4997 gnd.n2719 240.244
R5318 gnd.n2720 gnd.n2719 240.244
R5319 gnd.n2721 gnd.n2720 240.244
R5320 gnd.n5014 gnd.n2721 240.244
R5321 gnd.n5014 gnd.n2724 240.244
R5322 gnd.n2725 gnd.n2724 240.244
R5323 gnd.n2726 gnd.n2725 240.244
R5324 gnd.n2730 gnd.n2726 240.244
R5325 gnd.n5032 gnd.n5031 240.244
R5326 gnd.n5036 gnd.n5035 240.244
R5327 gnd.n5038 gnd.n5037 240.244
R5328 gnd.n2878 gnd.n2877 240.244
R5329 gnd.n2880 gnd.n2879 240.244
R5330 gnd.n5201 gnd.n5200 240.244
R5331 gnd.n5211 gnd.n5210 240.244
R5332 gnd.n5213 gnd.n5212 240.244
R5333 gnd.n5221 gnd.n5220 240.244
R5334 gnd.n5231 gnd.n5230 240.244
R5335 gnd.n5233 gnd.n5232 240.244
R5336 gnd.n5407 gnd.n2747 240.244
R5337 gnd.n5407 gnd.n2748 240.244
R5338 gnd.n2761 gnd.n2731 240.244
R5339 gnd.n2589 gnd.n2588 240.132
R5340 gnd.n4832 gnd.n4831 240.132
R5341 gnd.n6168 gnd.n590 225.874
R5342 gnd.n6176 gnd.n590 225.874
R5343 gnd.n6177 gnd.n6176 225.874
R5344 gnd.n6178 gnd.n6177 225.874
R5345 gnd.n6178 gnd.n584 225.874
R5346 gnd.n6186 gnd.n584 225.874
R5347 gnd.n6187 gnd.n6186 225.874
R5348 gnd.n6188 gnd.n6187 225.874
R5349 gnd.n6188 gnd.n578 225.874
R5350 gnd.n6196 gnd.n578 225.874
R5351 gnd.n6197 gnd.n6196 225.874
R5352 gnd.n6198 gnd.n6197 225.874
R5353 gnd.n6198 gnd.n572 225.874
R5354 gnd.n6206 gnd.n572 225.874
R5355 gnd.n6207 gnd.n6206 225.874
R5356 gnd.n6208 gnd.n6207 225.874
R5357 gnd.n6208 gnd.n566 225.874
R5358 gnd.n6216 gnd.n566 225.874
R5359 gnd.n6217 gnd.n6216 225.874
R5360 gnd.n6218 gnd.n6217 225.874
R5361 gnd.n6218 gnd.n560 225.874
R5362 gnd.n6226 gnd.n560 225.874
R5363 gnd.n6227 gnd.n6226 225.874
R5364 gnd.n6228 gnd.n6227 225.874
R5365 gnd.n6228 gnd.n554 225.874
R5366 gnd.n6236 gnd.n554 225.874
R5367 gnd.n6237 gnd.n6236 225.874
R5368 gnd.n6238 gnd.n6237 225.874
R5369 gnd.n6238 gnd.n548 225.874
R5370 gnd.n6246 gnd.n548 225.874
R5371 gnd.n6247 gnd.n6246 225.874
R5372 gnd.n6248 gnd.n6247 225.874
R5373 gnd.n6248 gnd.n542 225.874
R5374 gnd.n6256 gnd.n542 225.874
R5375 gnd.n6257 gnd.n6256 225.874
R5376 gnd.n6258 gnd.n6257 225.874
R5377 gnd.n6258 gnd.n536 225.874
R5378 gnd.n6266 gnd.n536 225.874
R5379 gnd.n6267 gnd.n6266 225.874
R5380 gnd.n6268 gnd.n6267 225.874
R5381 gnd.n6268 gnd.n530 225.874
R5382 gnd.n6276 gnd.n530 225.874
R5383 gnd.n6277 gnd.n6276 225.874
R5384 gnd.n6278 gnd.n6277 225.874
R5385 gnd.n6278 gnd.n524 225.874
R5386 gnd.n6286 gnd.n524 225.874
R5387 gnd.n6287 gnd.n6286 225.874
R5388 gnd.n6288 gnd.n6287 225.874
R5389 gnd.n6288 gnd.n518 225.874
R5390 gnd.n6296 gnd.n518 225.874
R5391 gnd.n6297 gnd.n6296 225.874
R5392 gnd.n6298 gnd.n6297 225.874
R5393 gnd.n6298 gnd.n512 225.874
R5394 gnd.n6306 gnd.n512 225.874
R5395 gnd.n6307 gnd.n6306 225.874
R5396 gnd.n6308 gnd.n6307 225.874
R5397 gnd.n6308 gnd.n506 225.874
R5398 gnd.n6316 gnd.n506 225.874
R5399 gnd.n6317 gnd.n6316 225.874
R5400 gnd.n6318 gnd.n6317 225.874
R5401 gnd.n6318 gnd.n500 225.874
R5402 gnd.n6326 gnd.n500 225.874
R5403 gnd.n6327 gnd.n6326 225.874
R5404 gnd.n6328 gnd.n6327 225.874
R5405 gnd.n6328 gnd.n494 225.874
R5406 gnd.n6336 gnd.n494 225.874
R5407 gnd.n6337 gnd.n6336 225.874
R5408 gnd.n6338 gnd.n6337 225.874
R5409 gnd.n6338 gnd.n488 225.874
R5410 gnd.n6346 gnd.n488 225.874
R5411 gnd.n6347 gnd.n6346 225.874
R5412 gnd.n6348 gnd.n6347 225.874
R5413 gnd.n6348 gnd.n482 225.874
R5414 gnd.n6356 gnd.n482 225.874
R5415 gnd.n6357 gnd.n6356 225.874
R5416 gnd.n6358 gnd.n6357 225.874
R5417 gnd.n6358 gnd.n476 225.874
R5418 gnd.n6366 gnd.n476 225.874
R5419 gnd.n6367 gnd.n6366 225.874
R5420 gnd.n6368 gnd.n6367 225.874
R5421 gnd.n6368 gnd.n470 225.874
R5422 gnd.n6376 gnd.n470 225.874
R5423 gnd.n6377 gnd.n6376 225.874
R5424 gnd.n6378 gnd.n6377 225.874
R5425 gnd.n6378 gnd.n464 225.874
R5426 gnd.n6386 gnd.n464 225.874
R5427 gnd.n6387 gnd.n6386 225.874
R5428 gnd.n6388 gnd.n6387 225.874
R5429 gnd.n6388 gnd.n458 225.874
R5430 gnd.n6396 gnd.n458 225.874
R5431 gnd.n6397 gnd.n6396 225.874
R5432 gnd.n6398 gnd.n6397 225.874
R5433 gnd.n6398 gnd.n452 225.874
R5434 gnd.n6406 gnd.n452 225.874
R5435 gnd.n6407 gnd.n6406 225.874
R5436 gnd.n6408 gnd.n6407 225.874
R5437 gnd.n6408 gnd.n446 225.874
R5438 gnd.n6416 gnd.n446 225.874
R5439 gnd.n6417 gnd.n6416 225.874
R5440 gnd.n6418 gnd.n6417 225.874
R5441 gnd.n6418 gnd.n440 225.874
R5442 gnd.n6426 gnd.n440 225.874
R5443 gnd.n6427 gnd.n6426 225.874
R5444 gnd.n6428 gnd.n6427 225.874
R5445 gnd.n6428 gnd.n434 225.874
R5446 gnd.n6436 gnd.n434 225.874
R5447 gnd.n6437 gnd.n6436 225.874
R5448 gnd.n6438 gnd.n6437 225.874
R5449 gnd.n6438 gnd.n428 225.874
R5450 gnd.n6446 gnd.n428 225.874
R5451 gnd.n6447 gnd.n6446 225.874
R5452 gnd.n6448 gnd.n6447 225.874
R5453 gnd.n6448 gnd.n422 225.874
R5454 gnd.n6456 gnd.n422 225.874
R5455 gnd.n6457 gnd.n6456 225.874
R5456 gnd.n6458 gnd.n6457 225.874
R5457 gnd.n6458 gnd.n416 225.874
R5458 gnd.n6466 gnd.n416 225.874
R5459 gnd.n6467 gnd.n6466 225.874
R5460 gnd.n6468 gnd.n6467 225.874
R5461 gnd.n6468 gnd.n410 225.874
R5462 gnd.n6476 gnd.n410 225.874
R5463 gnd.n6477 gnd.n6476 225.874
R5464 gnd.n6478 gnd.n6477 225.874
R5465 gnd.n6478 gnd.n404 225.874
R5466 gnd.n6486 gnd.n404 225.874
R5467 gnd.n6487 gnd.n6486 225.874
R5468 gnd.n6488 gnd.n6487 225.874
R5469 gnd.n6488 gnd.n398 225.874
R5470 gnd.n6496 gnd.n398 225.874
R5471 gnd.n6497 gnd.n6496 225.874
R5472 gnd.n6498 gnd.n6497 225.874
R5473 gnd.n6498 gnd.n392 225.874
R5474 gnd.n6506 gnd.n392 225.874
R5475 gnd.n6507 gnd.n6506 225.874
R5476 gnd.n6508 gnd.n6507 225.874
R5477 gnd.n6508 gnd.n386 225.874
R5478 gnd.n6517 gnd.n386 225.874
R5479 gnd.n6518 gnd.n6517 225.874
R5480 gnd.n6519 gnd.n6518 225.874
R5481 gnd.n6519 gnd.n381 225.874
R5482 gnd.n1409 gnd.t302 224.174
R5483 gnd.n805 gnd.t212 224.174
R5484 gnd.n2837 gnd.n2778 199.319
R5485 gnd.n2837 gnd.n2779 199.319
R5486 gnd.n2542 gnd.n2502 199.319
R5487 gnd.n2542 gnd.n2501 199.319
R5488 gnd.n2590 gnd.n2587 186.49
R5489 gnd.n4833 gnd.n4830 186.49
R5490 gnd.n2124 gnd.n2123 185
R5491 gnd.n2122 gnd.n2121 185
R5492 gnd.n2101 gnd.n2100 185
R5493 gnd.n2116 gnd.n2115 185
R5494 gnd.n2114 gnd.n2113 185
R5495 gnd.n2105 gnd.n2104 185
R5496 gnd.n2108 gnd.n2107 185
R5497 gnd.n2092 gnd.n2091 185
R5498 gnd.n2090 gnd.n2089 185
R5499 gnd.n2069 gnd.n2068 185
R5500 gnd.n2084 gnd.n2083 185
R5501 gnd.n2082 gnd.n2081 185
R5502 gnd.n2073 gnd.n2072 185
R5503 gnd.n2076 gnd.n2075 185
R5504 gnd.n2060 gnd.n2059 185
R5505 gnd.n2058 gnd.n2057 185
R5506 gnd.n2037 gnd.n2036 185
R5507 gnd.n2052 gnd.n2051 185
R5508 gnd.n2050 gnd.n2049 185
R5509 gnd.n2041 gnd.n2040 185
R5510 gnd.n2044 gnd.n2043 185
R5511 gnd.n2029 gnd.n2028 185
R5512 gnd.n2027 gnd.n2026 185
R5513 gnd.n2006 gnd.n2005 185
R5514 gnd.n2021 gnd.n2020 185
R5515 gnd.n2019 gnd.n2018 185
R5516 gnd.n2010 gnd.n2009 185
R5517 gnd.n2013 gnd.n2012 185
R5518 gnd.n1997 gnd.n1996 185
R5519 gnd.n1995 gnd.n1994 185
R5520 gnd.n1974 gnd.n1973 185
R5521 gnd.n1989 gnd.n1988 185
R5522 gnd.n1987 gnd.n1986 185
R5523 gnd.n1978 gnd.n1977 185
R5524 gnd.n1981 gnd.n1980 185
R5525 gnd.n1965 gnd.n1964 185
R5526 gnd.n1963 gnd.n1962 185
R5527 gnd.n1942 gnd.n1941 185
R5528 gnd.n1957 gnd.n1956 185
R5529 gnd.n1955 gnd.n1954 185
R5530 gnd.n1946 gnd.n1945 185
R5531 gnd.n1949 gnd.n1948 185
R5532 gnd.n1933 gnd.n1932 185
R5533 gnd.n1931 gnd.n1930 185
R5534 gnd.n1910 gnd.n1909 185
R5535 gnd.n1925 gnd.n1924 185
R5536 gnd.n1923 gnd.n1922 185
R5537 gnd.n1914 gnd.n1913 185
R5538 gnd.n1917 gnd.n1916 185
R5539 gnd.n1902 gnd.n1901 185
R5540 gnd.n1900 gnd.n1899 185
R5541 gnd.n1879 gnd.n1878 185
R5542 gnd.n1894 gnd.n1893 185
R5543 gnd.n1892 gnd.n1891 185
R5544 gnd.n1883 gnd.n1882 185
R5545 gnd.n1886 gnd.n1885 185
R5546 gnd.n1410 gnd.t301 178.987
R5547 gnd.n806 gnd.t213 178.987
R5548 gnd.n1 gnd.t2 170.774
R5549 gnd.n9 gnd.t323 170.103
R5550 gnd.n8 gnd.t159 170.103
R5551 gnd.n7 gnd.t106 170.103
R5552 gnd.n6 gnd.t66 170.103
R5553 gnd.n5 gnd.t113 170.103
R5554 gnd.n4 gnd.t117 170.103
R5555 gnd.n3 gnd.t154 170.103
R5556 gnd.n2 gnd.t95 170.103
R5557 gnd.n1 gnd.t31 170.103
R5558 gnd.n4904 gnd.n4903 163.367
R5559 gnd.n4900 gnd.n4899 163.367
R5560 gnd.n4896 gnd.n4895 163.367
R5561 gnd.n4892 gnd.n4891 163.367
R5562 gnd.n4888 gnd.n4887 163.367
R5563 gnd.n4884 gnd.n4883 163.367
R5564 gnd.n4880 gnd.n4879 163.367
R5565 gnd.n4876 gnd.n4875 163.367
R5566 gnd.n4872 gnd.n4871 163.367
R5567 gnd.n4868 gnd.n4867 163.367
R5568 gnd.n4864 gnd.n4863 163.367
R5569 gnd.n4860 gnd.n4859 163.367
R5570 gnd.n4856 gnd.n4855 163.367
R5571 gnd.n4852 gnd.n4851 163.367
R5572 gnd.n4847 gnd.n4846 163.367
R5573 gnd.n4843 gnd.n4842 163.367
R5574 gnd.n4977 gnd.n4976 163.367
R5575 gnd.n4973 gnd.n4972 163.367
R5576 gnd.n4968 gnd.n4967 163.367
R5577 gnd.n4964 gnd.n4963 163.367
R5578 gnd.n4960 gnd.n4959 163.367
R5579 gnd.n4956 gnd.n4955 163.367
R5580 gnd.n4952 gnd.n4951 163.367
R5581 gnd.n4948 gnd.n4947 163.367
R5582 gnd.n4944 gnd.n4943 163.367
R5583 gnd.n4940 gnd.n4939 163.367
R5584 gnd.n4936 gnd.n4935 163.367
R5585 gnd.n4932 gnd.n4931 163.367
R5586 gnd.n4928 gnd.n4927 163.367
R5587 gnd.n4924 gnd.n4923 163.367
R5588 gnd.n4920 gnd.n4919 163.367
R5589 gnd.n4916 gnd.n4915 163.367
R5590 gnd.n4128 gnd.n2606 163.367
R5591 gnd.n4131 gnd.n2606 163.367
R5592 gnd.n4131 gnd.n4062 163.367
R5593 gnd.n4136 gnd.n4062 163.367
R5594 gnd.n4136 gnd.n3342 163.367
R5595 gnd.n3342 gnd.n3332 163.367
R5596 gnd.n4172 gnd.n3332 163.367
R5597 gnd.n4172 gnd.n3329 163.367
R5598 gnd.n4183 gnd.n3329 163.367
R5599 gnd.n4183 gnd.n3330 163.367
R5600 gnd.n3330 gnd.n3322 163.367
R5601 gnd.n4178 gnd.n3322 163.367
R5602 gnd.n4178 gnd.n3311 163.367
R5603 gnd.n4175 gnd.n3311 163.367
R5604 gnd.n4175 gnd.n3305 163.367
R5605 gnd.n4213 gnd.n3305 163.367
R5606 gnd.n4213 gnd.n3298 163.367
R5607 gnd.n4216 gnd.n3298 163.367
R5608 gnd.n4216 gnd.n3292 163.367
R5609 gnd.n4220 gnd.n3292 163.367
R5610 gnd.n4220 gnd.n3282 163.367
R5611 gnd.n4270 gnd.n3282 163.367
R5612 gnd.n4270 gnd.n3279 163.367
R5613 gnd.n4278 gnd.n3279 163.367
R5614 gnd.n4278 gnd.n3274 163.367
R5615 gnd.n4274 gnd.n3274 163.367
R5616 gnd.n4274 gnd.n3265 163.367
R5617 gnd.n3265 gnd.n3256 163.367
R5618 gnd.n4307 gnd.n3256 163.367
R5619 gnd.n4307 gnd.n3253 163.367
R5620 gnd.n4350 gnd.n3253 163.367
R5621 gnd.n4350 gnd.n3254 163.367
R5622 gnd.n3254 gnd.n3247 163.367
R5623 gnd.n4345 gnd.n3247 163.367
R5624 gnd.n4345 gnd.n4342 163.367
R5625 gnd.n4342 gnd.n4341 163.367
R5626 gnd.n4341 gnd.n4313 163.367
R5627 gnd.n4313 gnd.n3229 163.367
R5628 gnd.n4336 gnd.n3229 163.367
R5629 gnd.n4336 gnd.n3224 163.367
R5630 gnd.n4333 gnd.n3224 163.367
R5631 gnd.n4333 gnd.n4329 163.367
R5632 gnd.n4329 gnd.n4328 163.367
R5633 gnd.n4328 gnd.n4317 163.367
R5634 gnd.n4317 gnd.n3207 163.367
R5635 gnd.n4323 gnd.n3207 163.367
R5636 gnd.n4323 gnd.n3203 163.367
R5637 gnd.n4320 gnd.n3203 163.367
R5638 gnd.n4320 gnd.n3193 163.367
R5639 gnd.n3193 gnd.n3185 163.367
R5640 gnd.n4454 gnd.n3185 163.367
R5641 gnd.n4454 gnd.n3182 163.367
R5642 gnd.n4492 gnd.n3182 163.367
R5643 gnd.n4492 gnd.n3183 163.367
R5644 gnd.n3183 gnd.n3174 163.367
R5645 gnd.n4487 gnd.n3174 163.367
R5646 gnd.n4487 gnd.n4485 163.367
R5647 gnd.n4485 gnd.n4484 163.367
R5648 gnd.n4484 gnd.n4458 163.367
R5649 gnd.n4458 gnd.n3155 163.367
R5650 gnd.n4479 gnd.n3155 163.367
R5651 gnd.n4479 gnd.n3149 163.367
R5652 gnd.n4476 gnd.n3149 163.367
R5653 gnd.n4476 gnd.n4473 163.367
R5654 gnd.n4473 gnd.n4472 163.367
R5655 gnd.n4472 gnd.n4461 163.367
R5656 gnd.n4461 gnd.n3131 163.367
R5657 gnd.n4467 gnd.n3131 163.367
R5658 gnd.n4467 gnd.n3126 163.367
R5659 gnd.n4464 gnd.n3126 163.367
R5660 gnd.n4464 gnd.n3115 163.367
R5661 gnd.n3115 gnd.n3107 163.367
R5662 gnd.n4595 gnd.n3107 163.367
R5663 gnd.n4595 gnd.n3104 163.367
R5664 gnd.n4617 gnd.n3104 163.367
R5665 gnd.n4617 gnd.n3105 163.367
R5666 gnd.n3105 gnd.n3097 163.367
R5667 gnd.n4612 gnd.n3097 163.367
R5668 gnd.n4612 gnd.n4610 163.367
R5669 gnd.n4610 gnd.n4609 163.367
R5670 gnd.n4609 gnd.n4599 163.367
R5671 gnd.n4599 gnd.n3079 163.367
R5672 gnd.n4604 gnd.n3079 163.367
R5673 gnd.n4604 gnd.n3073 163.367
R5674 gnd.n4601 gnd.n3073 163.367
R5675 gnd.n4601 gnd.n3062 163.367
R5676 gnd.n3062 gnd.n3055 163.367
R5677 gnd.n4691 gnd.n3055 163.367
R5678 gnd.n4691 gnd.n3052 163.367
R5679 gnd.n4705 gnd.n3052 163.367
R5680 gnd.n4705 gnd.n3053 163.367
R5681 gnd.n3053 gnd.n3045 163.367
R5682 gnd.n4700 gnd.n3045 163.367
R5683 gnd.n4700 gnd.n4699 163.367
R5684 gnd.n4699 gnd.n4698 163.367
R5685 gnd.n4698 gnd.n3014 163.367
R5686 gnd.n3014 gnd.n3008 163.367
R5687 gnd.n4773 gnd.n3008 163.367
R5688 gnd.n4773 gnd.n3006 163.367
R5689 gnd.n4778 gnd.n3006 163.367
R5690 gnd.n4778 gnd.n2999 163.367
R5691 gnd.n4787 gnd.n2999 163.367
R5692 gnd.n4788 gnd.n4787 163.367
R5693 gnd.n4788 gnd.n2996 163.367
R5694 gnd.n4797 gnd.n2996 163.367
R5695 gnd.n4797 gnd.n2990 163.367
R5696 gnd.n4793 gnd.n2990 163.367
R5697 gnd.n4793 gnd.n2981 163.367
R5698 gnd.n2981 gnd.n2976 163.367
R5699 gnd.n4911 gnd.n2976 163.367
R5700 gnd.n2581 gnd.n2580 163.367
R5701 gnd.n5613 gnd.n2580 163.367
R5702 gnd.n5611 gnd.n5610 163.367
R5703 gnd.n5607 gnd.n5606 163.367
R5704 gnd.n5603 gnd.n5602 163.367
R5705 gnd.n5599 gnd.n5598 163.367
R5706 gnd.n5595 gnd.n5594 163.367
R5707 gnd.n5591 gnd.n5590 163.367
R5708 gnd.n5587 gnd.n5586 163.367
R5709 gnd.n5583 gnd.n5582 163.367
R5710 gnd.n5579 gnd.n5578 163.367
R5711 gnd.n5575 gnd.n5574 163.367
R5712 gnd.n5571 gnd.n5570 163.367
R5713 gnd.n5567 gnd.n5566 163.367
R5714 gnd.n5563 gnd.n5562 163.367
R5715 gnd.n5559 gnd.n5558 163.367
R5716 gnd.n5622 gnd.n2547 163.367
R5717 gnd.n4067 gnd.n4066 163.367
R5718 gnd.n4072 gnd.n4071 163.367
R5719 gnd.n4076 gnd.n4075 163.367
R5720 gnd.n4080 gnd.n4079 163.367
R5721 gnd.n4084 gnd.n4083 163.367
R5722 gnd.n4088 gnd.n4087 163.367
R5723 gnd.n4092 gnd.n4091 163.367
R5724 gnd.n4096 gnd.n4095 163.367
R5725 gnd.n4100 gnd.n4099 163.367
R5726 gnd.n4104 gnd.n4103 163.367
R5727 gnd.n4108 gnd.n4107 163.367
R5728 gnd.n4112 gnd.n4111 163.367
R5729 gnd.n4116 gnd.n4115 163.367
R5730 gnd.n4120 gnd.n4119 163.367
R5731 gnd.n4124 gnd.n4123 163.367
R5732 gnd.n5551 gnd.n2582 163.367
R5733 gnd.n5551 gnd.n2604 163.367
R5734 gnd.n4139 gnd.n2604 163.367
R5735 gnd.n4139 gnd.n3341 163.367
R5736 gnd.n4166 gnd.n3341 163.367
R5737 gnd.n4166 gnd.n3339 163.367
R5738 gnd.n4170 gnd.n3339 163.367
R5739 gnd.n4170 gnd.n3327 163.367
R5740 gnd.n4185 gnd.n3327 163.367
R5741 gnd.n4185 gnd.n3325 163.367
R5742 gnd.n4189 gnd.n3325 163.367
R5743 gnd.n4189 gnd.n3309 163.367
R5744 gnd.n4206 gnd.n3309 163.367
R5745 gnd.n4206 gnd.n3307 163.367
R5746 gnd.n4210 gnd.n3307 163.367
R5747 gnd.n4210 gnd.n3296 163.367
R5748 gnd.n4251 gnd.n3296 163.367
R5749 gnd.n4251 gnd.n3293 163.367
R5750 gnd.n4258 gnd.n3293 163.367
R5751 gnd.n4258 gnd.n3294 163.367
R5752 gnd.n4254 gnd.n3294 163.367
R5753 gnd.n4254 gnd.n3278 163.367
R5754 gnd.n4283 gnd.n3278 163.367
R5755 gnd.n4283 gnd.n3276 163.367
R5756 gnd.n4287 gnd.n3276 163.367
R5757 gnd.n4287 gnd.n3263 163.367
R5758 gnd.n4301 gnd.n3263 163.367
R5759 gnd.n4301 gnd.n3261 163.367
R5760 gnd.n4305 gnd.n3261 163.367
R5761 gnd.n4305 gnd.n3251 163.367
R5762 gnd.n4352 gnd.n3251 163.367
R5763 gnd.n4352 gnd.n3248 163.367
R5764 gnd.n4361 gnd.n3248 163.367
R5765 gnd.n4361 gnd.n3249 163.367
R5766 gnd.n4357 gnd.n3249 163.367
R5767 gnd.n4357 gnd.n4356 163.367
R5768 gnd.n4356 gnd.n3228 163.367
R5769 gnd.n4384 gnd.n3228 163.367
R5770 gnd.n4384 gnd.n3225 163.367
R5771 gnd.n4393 gnd.n3225 163.367
R5772 gnd.n4393 gnd.n3226 163.367
R5773 gnd.n4389 gnd.n3226 163.367
R5774 gnd.n4389 gnd.n4388 163.367
R5775 gnd.n4388 gnd.n3206 163.367
R5776 gnd.n4429 gnd.n3206 163.367
R5777 gnd.n4429 gnd.n3204 163.367
R5778 gnd.n4433 gnd.n3204 163.367
R5779 gnd.n4433 gnd.n3191 163.367
R5780 gnd.n4448 gnd.n3191 163.367
R5781 gnd.n4448 gnd.n3189 163.367
R5782 gnd.n4452 gnd.n3189 163.367
R5783 gnd.n4452 gnd.n3179 163.367
R5784 gnd.n4494 gnd.n3179 163.367
R5785 gnd.n4494 gnd.n3176 163.367
R5786 gnd.n4503 gnd.n3176 163.367
R5787 gnd.n4503 gnd.n3177 163.367
R5788 gnd.n4499 gnd.n3177 163.367
R5789 gnd.n4499 gnd.n4498 163.367
R5790 gnd.n4498 gnd.n3153 163.367
R5791 gnd.n4526 gnd.n3153 163.367
R5792 gnd.n4526 gnd.n3150 163.367
R5793 gnd.n4535 gnd.n3150 163.367
R5794 gnd.n4535 gnd.n3151 163.367
R5795 gnd.n4531 gnd.n3151 163.367
R5796 gnd.n4531 gnd.n4530 163.367
R5797 gnd.n4530 gnd.n3129 163.367
R5798 gnd.n4571 gnd.n3129 163.367
R5799 gnd.n4571 gnd.n3127 163.367
R5800 gnd.n4575 gnd.n3127 163.367
R5801 gnd.n4575 gnd.n3112 163.367
R5802 gnd.n4589 gnd.n3112 163.367
R5803 gnd.n4589 gnd.n3110 163.367
R5804 gnd.n4593 gnd.n3110 163.367
R5805 gnd.n4593 gnd.n3102 163.367
R5806 gnd.n4619 gnd.n3102 163.367
R5807 gnd.n4619 gnd.n3099 163.367
R5808 gnd.n4628 gnd.n3099 163.367
R5809 gnd.n4628 gnd.n3100 163.367
R5810 gnd.n4624 gnd.n3100 163.367
R5811 gnd.n4624 gnd.n4623 163.367
R5812 gnd.n4623 gnd.n3077 163.367
R5813 gnd.n4667 gnd.n3077 163.367
R5814 gnd.n4667 gnd.n3075 163.367
R5815 gnd.n4671 gnd.n3075 163.367
R5816 gnd.n4671 gnd.n3061 163.367
R5817 gnd.n4685 gnd.n3061 163.367
R5818 gnd.n4685 gnd.n3059 163.367
R5819 gnd.n4689 gnd.n3059 163.367
R5820 gnd.n4689 gnd.n3050 163.367
R5821 gnd.n4707 gnd.n3050 163.367
R5822 gnd.n4707 gnd.n3047 163.367
R5823 gnd.n4714 gnd.n3047 163.367
R5824 gnd.n4714 gnd.n3048 163.367
R5825 gnd.n4710 gnd.n3048 163.367
R5826 gnd.n4710 gnd.n3012 163.367
R5827 gnd.n4767 gnd.n3012 163.367
R5828 gnd.n4767 gnd.n3010 163.367
R5829 gnd.n4771 gnd.n3010 163.367
R5830 gnd.n4771 gnd.n3003 163.367
R5831 gnd.n4781 gnd.n3003 163.367
R5832 gnd.n4781 gnd.n3001 163.367
R5833 gnd.n4785 gnd.n3001 163.367
R5834 gnd.n4785 gnd.n2994 163.367
R5835 gnd.n4801 gnd.n2994 163.367
R5836 gnd.n4801 gnd.n2992 163.367
R5837 gnd.n4805 gnd.n2992 163.367
R5838 gnd.n4805 gnd.n2980 163.367
R5839 gnd.n4818 gnd.n2980 163.367
R5840 gnd.n4818 gnd.n2977 163.367
R5841 gnd.n4909 gnd.n2977 163.367
R5842 gnd.n4839 gnd.n4838 156.462
R5843 gnd.n2064 gnd.n2032 153.042
R5844 gnd.n2128 gnd.n2127 152.079
R5845 gnd.n2096 gnd.n2095 152.079
R5846 gnd.n2064 gnd.n2063 152.079
R5847 gnd.n2595 gnd.n2594 152
R5848 gnd.n2596 gnd.n2585 152
R5849 gnd.n2598 gnd.n2597 152
R5850 gnd.n2600 gnd.n2583 152
R5851 gnd.n2602 gnd.n2601 152
R5852 gnd.n4837 gnd.n4821 152
R5853 gnd.n4829 gnd.n4822 152
R5854 gnd.n4828 gnd.n4827 152
R5855 gnd.n4826 gnd.n4823 152
R5856 gnd.n4824 gnd.t281 150.546
R5857 gnd.t109 gnd.n2106 147.661
R5858 gnd.t12 gnd.n2074 147.661
R5859 gnd.t332 gnd.n2042 147.661
R5860 gnd.t25 gnd.n2011 147.661
R5861 gnd.t150 gnd.n1979 147.661
R5862 gnd.t49 gnd.n1947 147.661
R5863 gnd.t7 gnd.n1915 147.661
R5864 gnd.t74 gnd.n1884 147.661
R5865 gnd.n2972 gnd.n2955 143.351
R5866 gnd.n2562 gnd.n2546 143.351
R5867 gnd.n5621 gnd.n2546 143.351
R5868 gnd.n2592 gnd.t203 130.484
R5869 gnd.n2601 gnd.t269 126.766
R5870 gnd.n2599 gnd.t200 126.766
R5871 gnd.n2585 gnd.t225 126.766
R5872 gnd.n2593 gnd.t303 126.766
R5873 gnd.n4825 gnd.t260 126.766
R5874 gnd.n4827 gnd.t197 126.766
R5875 gnd.n4836 gnd.t239 126.766
R5876 gnd.n4838 gnd.t218 126.766
R5877 gnd.n5344 gnd.n2836 104.897
R5878 gnd.n5624 gnd.n5623 104.897
R5879 gnd.n2123 gnd.n2122 104.615
R5880 gnd.n2122 gnd.n2100 104.615
R5881 gnd.n2115 gnd.n2100 104.615
R5882 gnd.n2115 gnd.n2114 104.615
R5883 gnd.n2114 gnd.n2104 104.615
R5884 gnd.n2107 gnd.n2104 104.615
R5885 gnd.n2091 gnd.n2090 104.615
R5886 gnd.n2090 gnd.n2068 104.615
R5887 gnd.n2083 gnd.n2068 104.615
R5888 gnd.n2083 gnd.n2082 104.615
R5889 gnd.n2082 gnd.n2072 104.615
R5890 gnd.n2075 gnd.n2072 104.615
R5891 gnd.n2059 gnd.n2058 104.615
R5892 gnd.n2058 gnd.n2036 104.615
R5893 gnd.n2051 gnd.n2036 104.615
R5894 gnd.n2051 gnd.n2050 104.615
R5895 gnd.n2050 gnd.n2040 104.615
R5896 gnd.n2043 gnd.n2040 104.615
R5897 gnd.n2028 gnd.n2027 104.615
R5898 gnd.n2027 gnd.n2005 104.615
R5899 gnd.n2020 gnd.n2005 104.615
R5900 gnd.n2020 gnd.n2019 104.615
R5901 gnd.n2019 gnd.n2009 104.615
R5902 gnd.n2012 gnd.n2009 104.615
R5903 gnd.n1996 gnd.n1995 104.615
R5904 gnd.n1995 gnd.n1973 104.615
R5905 gnd.n1988 gnd.n1973 104.615
R5906 gnd.n1988 gnd.n1987 104.615
R5907 gnd.n1987 gnd.n1977 104.615
R5908 gnd.n1980 gnd.n1977 104.615
R5909 gnd.n1964 gnd.n1963 104.615
R5910 gnd.n1963 gnd.n1941 104.615
R5911 gnd.n1956 gnd.n1941 104.615
R5912 gnd.n1956 gnd.n1955 104.615
R5913 gnd.n1955 gnd.n1945 104.615
R5914 gnd.n1948 gnd.n1945 104.615
R5915 gnd.n1932 gnd.n1931 104.615
R5916 gnd.n1931 gnd.n1909 104.615
R5917 gnd.n1924 gnd.n1909 104.615
R5918 gnd.n1924 gnd.n1923 104.615
R5919 gnd.n1923 gnd.n1913 104.615
R5920 gnd.n1916 gnd.n1913 104.615
R5921 gnd.n1901 gnd.n1900 104.615
R5922 gnd.n1900 gnd.n1878 104.615
R5923 gnd.n1893 gnd.n1878 104.615
R5924 gnd.n1893 gnd.n1892 104.615
R5925 gnd.n1892 gnd.n1882 104.615
R5926 gnd.n1885 gnd.n1882 104.615
R5927 gnd.n1335 gnd.t259 100.632
R5928 gnd.n784 gnd.t311 100.632
R5929 gnd.n6528 gnd.n6527 100.343
R5930 gnd.n6529 gnd.n6528 100.343
R5931 gnd.n6529 gnd.n375 100.343
R5932 gnd.n6537 gnd.n375 100.343
R5933 gnd.n6538 gnd.n6537 100.343
R5934 gnd.n6539 gnd.n6538 100.343
R5935 gnd.n6539 gnd.n369 100.343
R5936 gnd.n6547 gnd.n369 100.343
R5937 gnd.n6548 gnd.n6547 100.343
R5938 gnd.n6549 gnd.n6548 100.343
R5939 gnd.n6549 gnd.n363 100.343
R5940 gnd.n6557 gnd.n363 100.343
R5941 gnd.n6558 gnd.n6557 100.343
R5942 gnd.n6559 gnd.n6558 100.343
R5943 gnd.n6559 gnd.n357 100.343
R5944 gnd.n6567 gnd.n357 100.343
R5945 gnd.n6568 gnd.n6567 100.343
R5946 gnd.n6569 gnd.n6568 100.343
R5947 gnd.n6569 gnd.n351 100.343
R5948 gnd.n6577 gnd.n351 100.343
R5949 gnd.n6578 gnd.n6577 100.343
R5950 gnd.n6579 gnd.n6578 100.343
R5951 gnd.n6579 gnd.n345 100.343
R5952 gnd.n6587 gnd.n345 100.343
R5953 gnd.n6588 gnd.n6587 100.343
R5954 gnd.n6589 gnd.n6588 100.343
R5955 gnd.n6589 gnd.n339 100.343
R5956 gnd.n6597 gnd.n339 100.343
R5957 gnd.n6598 gnd.n6597 100.343
R5958 gnd.n6599 gnd.n6598 100.343
R5959 gnd.n6599 gnd.n333 100.343
R5960 gnd.n6607 gnd.n333 100.343
R5961 gnd.n6608 gnd.n6607 100.343
R5962 gnd.n6609 gnd.n6608 100.343
R5963 gnd.n6609 gnd.n327 100.343
R5964 gnd.n6617 gnd.n327 100.343
R5965 gnd.n6618 gnd.n6617 100.343
R5966 gnd.n6619 gnd.n6618 100.343
R5967 gnd.n6619 gnd.n321 100.343
R5968 gnd.n6627 gnd.n321 100.343
R5969 gnd.n6628 gnd.n6627 100.343
R5970 gnd.n6629 gnd.n6628 100.343
R5971 gnd.n6629 gnd.n315 100.343
R5972 gnd.n6637 gnd.n315 100.343
R5973 gnd.n6638 gnd.n6637 100.343
R5974 gnd.n6639 gnd.n6638 100.343
R5975 gnd.n6639 gnd.n309 100.343
R5976 gnd.n6647 gnd.n309 100.343
R5977 gnd.n6648 gnd.n6647 100.343
R5978 gnd.n6649 gnd.n6648 100.343
R5979 gnd.n6649 gnd.n303 100.343
R5980 gnd.n6657 gnd.n303 100.343
R5981 gnd.n6658 gnd.n6657 100.343
R5982 gnd.n6659 gnd.n6658 100.343
R5983 gnd.n6659 gnd.n297 100.343
R5984 gnd.n6667 gnd.n297 100.343
R5985 gnd.n6668 gnd.n6667 100.343
R5986 gnd.n6669 gnd.n6668 100.343
R5987 gnd.n6669 gnd.n291 100.343
R5988 gnd.n6677 gnd.n291 100.343
R5989 gnd.n6678 gnd.n6677 100.343
R5990 gnd.n6679 gnd.n6678 100.343
R5991 gnd.n6679 gnd.n285 100.343
R5992 gnd.n6687 gnd.n285 100.343
R5993 gnd.n6688 gnd.n6687 100.343
R5994 gnd.n6689 gnd.n6688 100.343
R5995 gnd.n6689 gnd.n279 100.343
R5996 gnd.n6697 gnd.n279 100.343
R5997 gnd.n6698 gnd.n6697 100.343
R5998 gnd.n6699 gnd.n6698 100.343
R5999 gnd.n6699 gnd.n273 100.343
R6000 gnd.n6707 gnd.n273 100.343
R6001 gnd.n6708 gnd.n6707 100.343
R6002 gnd.n6709 gnd.n6708 100.343
R6003 gnd.n6709 gnd.n267 100.343
R6004 gnd.n6717 gnd.n267 100.343
R6005 gnd.n6718 gnd.n6717 100.343
R6006 gnd.n6719 gnd.n6718 100.343
R6007 gnd.n6719 gnd.n261 100.343
R6008 gnd.n6727 gnd.n261 100.343
R6009 gnd.n6728 gnd.n6727 100.343
R6010 gnd.n6730 gnd.n6728 100.343
R6011 gnd.n6730 gnd.n6729 100.343
R6012 gnd.n7190 gnd.n7021 99.6594
R6013 gnd.n7188 gnd.n7020 99.6594
R6014 gnd.n7184 gnd.n7019 99.6594
R6015 gnd.n7180 gnd.n7018 99.6594
R6016 gnd.n7176 gnd.n7017 99.6594
R6017 gnd.n7172 gnd.n7016 99.6594
R6018 gnd.n7168 gnd.n7015 99.6594
R6019 gnd.n7164 gnd.n7014 99.6594
R6020 gnd.n7157 gnd.n7013 99.6594
R6021 gnd.n7153 gnd.n7012 99.6594
R6022 gnd.n7149 gnd.n7011 99.6594
R6023 gnd.n7145 gnd.n7010 99.6594
R6024 gnd.n7141 gnd.n7009 99.6594
R6025 gnd.n7137 gnd.n7008 99.6594
R6026 gnd.n7133 gnd.n7007 99.6594
R6027 gnd.n7129 gnd.n7006 99.6594
R6028 gnd.n7125 gnd.n7005 99.6594
R6029 gnd.n7121 gnd.n7004 99.6594
R6030 gnd.n7113 gnd.n7003 99.6594
R6031 gnd.n7111 gnd.n7002 99.6594
R6032 gnd.n7107 gnd.n7001 99.6594
R6033 gnd.n7103 gnd.n7000 99.6594
R6034 gnd.n7099 gnd.n6999 99.6594
R6035 gnd.n7095 gnd.n6998 99.6594
R6036 gnd.n7091 gnd.n6997 99.6594
R6037 gnd.n7087 gnd.n6996 99.6594
R6038 gnd.n7083 gnd.n6995 99.6594
R6039 gnd.n7079 gnd.n6994 99.6594
R6040 gnd.n7202 gnd.n7200 99.6594
R6041 gnd.n5396 gnd.n5395 99.6594
R6042 gnd.n5390 gnd.n2767 99.6594
R6043 gnd.n5387 gnd.n2768 99.6594
R6044 gnd.n5383 gnd.n2769 99.6594
R6045 gnd.n5379 gnd.n2770 99.6594
R6046 gnd.n5375 gnd.n2771 99.6594
R6047 gnd.n5371 gnd.n2772 99.6594
R6048 gnd.n5367 gnd.n2773 99.6594
R6049 gnd.n5363 gnd.n2774 99.6594
R6050 gnd.n5358 gnd.n2775 99.6594
R6051 gnd.n5354 gnd.n2776 99.6594
R6052 gnd.n5350 gnd.n2777 99.6594
R6053 gnd.n5346 gnd.n2778 99.6594
R6054 gnd.n5341 gnd.n2780 99.6594
R6055 gnd.n5337 gnd.n2781 99.6594
R6056 gnd.n5333 gnd.n2782 99.6594
R6057 gnd.n5329 gnd.n2783 99.6594
R6058 gnd.n5325 gnd.n2784 99.6594
R6059 gnd.n5321 gnd.n2785 99.6594
R6060 gnd.n5317 gnd.n2786 99.6594
R6061 gnd.n5313 gnd.n2787 99.6594
R6062 gnd.n5309 gnd.n2788 99.6594
R6063 gnd.n5305 gnd.n2789 99.6594
R6064 gnd.n5301 gnd.n2790 99.6594
R6065 gnd.n5297 gnd.n2791 99.6594
R6066 gnd.n5293 gnd.n2792 99.6594
R6067 gnd.n5289 gnd.n2793 99.6594
R6068 gnd.n5285 gnd.n2794 99.6594
R6069 gnd.n5673 gnd.n5672 99.6594
R6070 gnd.n5668 gnd.n2513 99.6594
R6071 gnd.n5664 gnd.n2512 99.6594
R6072 gnd.n5660 gnd.n2511 99.6594
R6073 gnd.n5656 gnd.n2510 99.6594
R6074 gnd.n5652 gnd.n2509 99.6594
R6075 gnd.n5648 gnd.n2508 99.6594
R6076 gnd.n5644 gnd.n2507 99.6594
R6077 gnd.n5639 gnd.n2506 99.6594
R6078 gnd.n5635 gnd.n2505 99.6594
R6079 gnd.n5631 gnd.n2504 99.6594
R6080 gnd.n5627 gnd.n2503 99.6594
R6081 gnd.n3539 gnd.n2501 99.6594
R6082 gnd.n3546 gnd.n2500 99.6594
R6083 gnd.n3550 gnd.n2499 99.6594
R6084 gnd.n3556 gnd.n2498 99.6594
R6085 gnd.n3560 gnd.n2497 99.6594
R6086 gnd.n3566 gnd.n2496 99.6594
R6087 gnd.n3570 gnd.n2495 99.6594
R6088 gnd.n3576 gnd.n2494 99.6594
R6089 gnd.n3580 gnd.n2493 99.6594
R6090 gnd.n3586 gnd.n2492 99.6594
R6091 gnd.n3590 gnd.n2491 99.6594
R6092 gnd.n3596 gnd.n2490 99.6594
R6093 gnd.n3600 gnd.n2489 99.6594
R6094 gnd.n3606 gnd.n2488 99.6594
R6095 gnd.n3610 gnd.n2487 99.6594
R6096 gnd.n3616 gnd.n2486 99.6594
R6097 gnd.n5927 gnd.n5926 99.6594
R6098 gnd.n5921 gnd.n2155 99.6594
R6099 gnd.n5918 gnd.n2156 99.6594
R6100 gnd.n5914 gnd.n2157 99.6594
R6101 gnd.n5910 gnd.n2158 99.6594
R6102 gnd.n5906 gnd.n2159 99.6594
R6103 gnd.n5902 gnd.n2160 99.6594
R6104 gnd.n5898 gnd.n2161 99.6594
R6105 gnd.n5894 gnd.n2162 99.6594
R6106 gnd.n5889 gnd.n2163 99.6594
R6107 gnd.n5885 gnd.n2164 99.6594
R6108 gnd.n5881 gnd.n2165 99.6594
R6109 gnd.n5877 gnd.n2166 99.6594
R6110 gnd.n5873 gnd.n2167 99.6594
R6111 gnd.n5869 gnd.n2168 99.6594
R6112 gnd.n5865 gnd.n2169 99.6594
R6113 gnd.n5861 gnd.n2170 99.6594
R6114 gnd.n5857 gnd.n2171 99.6594
R6115 gnd.n5853 gnd.n2172 99.6594
R6116 gnd.n5849 gnd.n2173 99.6594
R6117 gnd.n5845 gnd.n2174 99.6594
R6118 gnd.n5841 gnd.n2175 99.6594
R6119 gnd.n5837 gnd.n2176 99.6594
R6120 gnd.n5833 gnd.n2177 99.6594
R6121 gnd.n5829 gnd.n2178 99.6594
R6122 gnd.n5825 gnd.n2179 99.6594
R6123 gnd.n5821 gnd.n2180 99.6594
R6124 gnd.n5817 gnd.n2181 99.6594
R6125 gnd.n5813 gnd.n2182 99.6594
R6126 gnd.n5966 gnd.n5934 99.6594
R6127 gnd.n5964 gnd.n5933 99.6594
R6128 gnd.n5960 gnd.n5932 99.6594
R6129 gnd.n5956 gnd.n5931 99.6594
R6130 gnd.n5952 gnd.n5930 99.6594
R6131 gnd.n5948 gnd.n5929 99.6594
R6132 gnd.n5978 gnd.n5976 99.6594
R6133 gnd.n5984 gnd.n783 99.6594
R6134 gnd.n1547 gnd.n1278 99.6594
R6135 gnd.n1304 gnd.n1285 99.6594
R6136 gnd.n1306 gnd.n1286 99.6594
R6137 gnd.n1314 gnd.n1287 99.6594
R6138 gnd.n1316 gnd.n1288 99.6594
R6139 gnd.n1324 gnd.n1289 99.6594
R6140 gnd.n1326 gnd.n1290 99.6594
R6141 gnd.n1334 gnd.n1291 99.6594
R6142 gnd.n6908 gnd.n6882 99.6594
R6143 gnd.n6912 gnd.n6883 99.6594
R6144 gnd.n6918 gnd.n6884 99.6594
R6145 gnd.n6922 gnd.n6885 99.6594
R6146 gnd.n6928 gnd.n6886 99.6594
R6147 gnd.n6932 gnd.n6887 99.6594
R6148 gnd.n6938 gnd.n6888 99.6594
R6149 gnd.n6941 gnd.n6889 99.6594
R6150 gnd.n6993 gnd.n6992 99.6594
R6151 gnd.n5194 gnd.n2795 99.6594
R6152 gnd.n5197 gnd.n2796 99.6594
R6153 gnd.n5205 gnd.n2797 99.6594
R6154 gnd.n5207 gnd.n2798 99.6594
R6155 gnd.n5217 gnd.n2799 99.6594
R6156 gnd.n5225 gnd.n2800 99.6594
R6157 gnd.n5227 gnd.n2801 99.6594
R6158 gnd.n5237 gnd.n2803 99.6594
R6159 gnd.n5398 gnd.n2756 99.6594
R6160 gnd.n825 gnd.n790 99.6594
R6161 gnd.n829 gnd.n791 99.6594
R6162 gnd.n835 gnd.n792 99.6594
R6163 gnd.n839 gnd.n793 99.6594
R6164 gnd.n845 gnd.n794 99.6594
R6165 gnd.n849 gnd.n795 99.6594
R6166 gnd.n855 gnd.n796 99.6594
R6167 gnd.n859 gnd.n797 99.6594
R6168 gnd.n865 gnd.n798 99.6594
R6169 gnd.n869 gnd.n799 99.6594
R6170 gnd.n875 gnd.n800 99.6594
R6171 gnd.n878 gnd.n801 99.6594
R6172 gnd.n2154 gnd.n2153 99.6594
R6173 gnd.n1462 gnd.n1461 99.6594
R6174 gnd.n1456 gnd.n1373 99.6594
R6175 gnd.n1453 gnd.n1374 99.6594
R6176 gnd.n1449 gnd.n1375 99.6594
R6177 gnd.n1445 gnd.n1376 99.6594
R6178 gnd.n1441 gnd.n1377 99.6594
R6179 gnd.n1437 gnd.n1378 99.6594
R6180 gnd.n1433 gnd.n1379 99.6594
R6181 gnd.n1429 gnd.n1380 99.6594
R6182 gnd.n1425 gnd.n1381 99.6594
R6183 gnd.n1421 gnd.n1382 99.6594
R6184 gnd.n1417 gnd.n1383 99.6594
R6185 gnd.n1464 gnd.n1372 99.6594
R6186 gnd.n3457 gnd.n2476 99.6594
R6187 gnd.n3467 gnd.n2477 99.6594
R6188 gnd.n3475 gnd.n2478 99.6594
R6189 gnd.n3477 gnd.n2479 99.6594
R6190 gnd.n3487 gnd.n2480 99.6594
R6191 gnd.n3495 gnd.n2481 99.6594
R6192 gnd.n3497 gnd.n2482 99.6594
R6193 gnd.n3508 gnd.n2483 99.6594
R6194 gnd.n3926 gnd.n2484 99.6594
R6195 gnd.n2265 gnd.n2183 99.6594
R6196 gnd.n3688 gnd.n2184 99.6594
R6197 gnd.n3694 gnd.n2185 99.6594
R6198 gnd.n3698 gnd.n2186 99.6594
R6199 gnd.n3704 gnd.n2187 99.6594
R6200 gnd.n3708 gnd.n2188 99.6594
R6201 gnd.n3714 gnd.n2189 99.6594
R6202 gnd.n3718 gnd.n2190 99.6594
R6203 gnd.n3677 gnd.n2191 99.6594
R6204 gnd.n3687 gnd.n2183 99.6594
R6205 gnd.n3693 gnd.n2184 99.6594
R6206 gnd.n3697 gnd.n2185 99.6594
R6207 gnd.n3703 gnd.n2186 99.6594
R6208 gnd.n3707 gnd.n2187 99.6594
R6209 gnd.n3713 gnd.n2188 99.6594
R6210 gnd.n3717 gnd.n2189 99.6594
R6211 gnd.n3676 gnd.n2190 99.6594
R6212 gnd.n3672 gnd.n2191 99.6594
R6213 gnd.n3512 gnd.n2484 99.6594
R6214 gnd.n3498 gnd.n2483 99.6594
R6215 gnd.n3496 gnd.n2482 99.6594
R6216 gnd.n3488 gnd.n2481 99.6594
R6217 gnd.n3478 gnd.n2480 99.6594
R6218 gnd.n3476 gnd.n2479 99.6594
R6219 gnd.n3468 gnd.n2478 99.6594
R6220 gnd.n3458 gnd.n2477 99.6594
R6221 gnd.n3456 gnd.n2476 99.6594
R6222 gnd.n1462 gnd.n1385 99.6594
R6223 gnd.n1454 gnd.n1373 99.6594
R6224 gnd.n1450 gnd.n1374 99.6594
R6225 gnd.n1446 gnd.n1375 99.6594
R6226 gnd.n1442 gnd.n1376 99.6594
R6227 gnd.n1438 gnd.n1377 99.6594
R6228 gnd.n1434 gnd.n1378 99.6594
R6229 gnd.n1430 gnd.n1379 99.6594
R6230 gnd.n1426 gnd.n1380 99.6594
R6231 gnd.n1422 gnd.n1381 99.6594
R6232 gnd.n1418 gnd.n1382 99.6594
R6233 gnd.n1414 gnd.n1383 99.6594
R6234 gnd.n1465 gnd.n1464 99.6594
R6235 gnd.n2154 gnd.n802 99.6594
R6236 gnd.n876 gnd.n801 99.6594
R6237 gnd.n868 gnd.n800 99.6594
R6238 gnd.n866 gnd.n799 99.6594
R6239 gnd.n858 gnd.n798 99.6594
R6240 gnd.n856 gnd.n797 99.6594
R6241 gnd.n848 gnd.n796 99.6594
R6242 gnd.n846 gnd.n795 99.6594
R6243 gnd.n838 gnd.n794 99.6594
R6244 gnd.n836 gnd.n793 99.6594
R6245 gnd.n828 gnd.n792 99.6594
R6246 gnd.n826 gnd.n791 99.6594
R6247 gnd.n818 gnd.n790 99.6594
R6248 gnd.n5196 gnd.n2795 99.6594
R6249 gnd.n5204 gnd.n2796 99.6594
R6250 gnd.n5206 gnd.n2797 99.6594
R6251 gnd.n5216 gnd.n2798 99.6594
R6252 gnd.n5224 gnd.n2799 99.6594
R6253 gnd.n5226 gnd.n2800 99.6594
R6254 gnd.n5236 gnd.n2801 99.6594
R6255 gnd.n2803 gnd.n2802 99.6594
R6256 gnd.n5399 gnd.n5398 99.6594
R6257 gnd.n6993 gnd.n6890 99.6594
R6258 gnd.n6939 gnd.n6889 99.6594
R6259 gnd.n6931 gnd.n6888 99.6594
R6260 gnd.n6929 gnd.n6887 99.6594
R6261 gnd.n6921 gnd.n6886 99.6594
R6262 gnd.n6919 gnd.n6885 99.6594
R6263 gnd.n6911 gnd.n6884 99.6594
R6264 gnd.n6909 gnd.n6883 99.6594
R6265 gnd.n6903 gnd.n6882 99.6594
R6266 gnd.n1548 gnd.n1547 99.6594
R6267 gnd.n1307 gnd.n1285 99.6594
R6268 gnd.n1313 gnd.n1286 99.6594
R6269 gnd.n1317 gnd.n1287 99.6594
R6270 gnd.n1323 gnd.n1288 99.6594
R6271 gnd.n1327 gnd.n1289 99.6594
R6272 gnd.n1333 gnd.n1290 99.6594
R6273 gnd.n1291 gnd.n1275 99.6594
R6274 gnd.n5977 gnd.n783 99.6594
R6275 gnd.n5976 gnd.n789 99.6594
R6276 gnd.n5951 gnd.n5929 99.6594
R6277 gnd.n5955 gnd.n5930 99.6594
R6278 gnd.n5959 gnd.n5931 99.6594
R6279 gnd.n5963 gnd.n5932 99.6594
R6280 gnd.n5967 gnd.n5933 99.6594
R6281 gnd.n5935 gnd.n5934 99.6594
R6282 gnd.n5927 gnd.n2195 99.6594
R6283 gnd.n5919 gnd.n2155 99.6594
R6284 gnd.n5915 gnd.n2156 99.6594
R6285 gnd.n5911 gnd.n2157 99.6594
R6286 gnd.n5907 gnd.n2158 99.6594
R6287 gnd.n5903 gnd.n2159 99.6594
R6288 gnd.n5899 gnd.n2160 99.6594
R6289 gnd.n5895 gnd.n2161 99.6594
R6290 gnd.n5890 gnd.n2162 99.6594
R6291 gnd.n5886 gnd.n2163 99.6594
R6292 gnd.n5882 gnd.n2164 99.6594
R6293 gnd.n5878 gnd.n2165 99.6594
R6294 gnd.n5874 gnd.n2166 99.6594
R6295 gnd.n5870 gnd.n2167 99.6594
R6296 gnd.n5866 gnd.n2168 99.6594
R6297 gnd.n5862 gnd.n2169 99.6594
R6298 gnd.n5858 gnd.n2170 99.6594
R6299 gnd.n5854 gnd.n2171 99.6594
R6300 gnd.n5850 gnd.n2172 99.6594
R6301 gnd.n5846 gnd.n2173 99.6594
R6302 gnd.n5842 gnd.n2174 99.6594
R6303 gnd.n5838 gnd.n2175 99.6594
R6304 gnd.n5834 gnd.n2176 99.6594
R6305 gnd.n5830 gnd.n2177 99.6594
R6306 gnd.n5826 gnd.n2178 99.6594
R6307 gnd.n5822 gnd.n2179 99.6594
R6308 gnd.n5818 gnd.n2180 99.6594
R6309 gnd.n5814 gnd.n2181 99.6594
R6310 gnd.n2267 gnd.n2182 99.6594
R6311 gnd.n3609 gnd.n2486 99.6594
R6312 gnd.n3607 gnd.n2487 99.6594
R6313 gnd.n3599 gnd.n2488 99.6594
R6314 gnd.n3597 gnd.n2489 99.6594
R6315 gnd.n3589 gnd.n2490 99.6594
R6316 gnd.n3587 gnd.n2491 99.6594
R6317 gnd.n3579 gnd.n2492 99.6594
R6318 gnd.n3577 gnd.n2493 99.6594
R6319 gnd.n3569 gnd.n2494 99.6594
R6320 gnd.n3567 gnd.n2495 99.6594
R6321 gnd.n3559 gnd.n2496 99.6594
R6322 gnd.n3557 gnd.n2497 99.6594
R6323 gnd.n3549 gnd.n2498 99.6594
R6324 gnd.n3547 gnd.n2499 99.6594
R6325 gnd.n3540 gnd.n2500 99.6594
R6326 gnd.n5626 gnd.n2502 99.6594
R6327 gnd.n5630 gnd.n2503 99.6594
R6328 gnd.n5634 gnd.n2504 99.6594
R6329 gnd.n5638 gnd.n2505 99.6594
R6330 gnd.n5643 gnd.n2506 99.6594
R6331 gnd.n5647 gnd.n2507 99.6594
R6332 gnd.n5651 gnd.n2508 99.6594
R6333 gnd.n5655 gnd.n2509 99.6594
R6334 gnd.n5659 gnd.n2510 99.6594
R6335 gnd.n5663 gnd.n2511 99.6594
R6336 gnd.n5667 gnd.n2512 99.6594
R6337 gnd.n2514 gnd.n2513 99.6594
R6338 gnd.n5673 gnd.n2473 99.6594
R6339 gnd.n5396 gnd.n2806 99.6594
R6340 gnd.n5388 gnd.n2767 99.6594
R6341 gnd.n5384 gnd.n2768 99.6594
R6342 gnd.n5380 gnd.n2769 99.6594
R6343 gnd.n5376 gnd.n2770 99.6594
R6344 gnd.n5372 gnd.n2771 99.6594
R6345 gnd.n5368 gnd.n2772 99.6594
R6346 gnd.n5364 gnd.n2773 99.6594
R6347 gnd.n5359 gnd.n2774 99.6594
R6348 gnd.n5355 gnd.n2775 99.6594
R6349 gnd.n5351 gnd.n2776 99.6594
R6350 gnd.n5347 gnd.n2777 99.6594
R6351 gnd.n5342 gnd.n2779 99.6594
R6352 gnd.n5338 gnd.n2780 99.6594
R6353 gnd.n5334 gnd.n2781 99.6594
R6354 gnd.n5330 gnd.n2782 99.6594
R6355 gnd.n5326 gnd.n2783 99.6594
R6356 gnd.n5322 gnd.n2784 99.6594
R6357 gnd.n5318 gnd.n2785 99.6594
R6358 gnd.n5314 gnd.n2786 99.6594
R6359 gnd.n5310 gnd.n2787 99.6594
R6360 gnd.n5306 gnd.n2788 99.6594
R6361 gnd.n5302 gnd.n2789 99.6594
R6362 gnd.n5298 gnd.n2790 99.6594
R6363 gnd.n5294 gnd.n2791 99.6594
R6364 gnd.n5290 gnd.n2792 99.6594
R6365 gnd.n5286 gnd.n2793 99.6594
R6366 gnd.n2887 gnd.n2794 99.6594
R6367 gnd.n7200 gnd.n6880 99.6594
R6368 gnd.n7082 gnd.n6994 99.6594
R6369 gnd.n7086 gnd.n6995 99.6594
R6370 gnd.n7090 gnd.n6996 99.6594
R6371 gnd.n7094 gnd.n6997 99.6594
R6372 gnd.n7098 gnd.n6998 99.6594
R6373 gnd.n7102 gnd.n6999 99.6594
R6374 gnd.n7106 gnd.n7000 99.6594
R6375 gnd.n7110 gnd.n7001 99.6594
R6376 gnd.n7114 gnd.n7002 99.6594
R6377 gnd.n7120 gnd.n7003 99.6594
R6378 gnd.n7124 gnd.n7004 99.6594
R6379 gnd.n7128 gnd.n7005 99.6594
R6380 gnd.n7132 gnd.n7006 99.6594
R6381 gnd.n7136 gnd.n7007 99.6594
R6382 gnd.n7140 gnd.n7008 99.6594
R6383 gnd.n7144 gnd.n7009 99.6594
R6384 gnd.n7148 gnd.n7010 99.6594
R6385 gnd.n7152 gnd.n7011 99.6594
R6386 gnd.n7156 gnd.n7012 99.6594
R6387 gnd.n7163 gnd.n7013 99.6594
R6388 gnd.n7167 gnd.n7014 99.6594
R6389 gnd.n7171 gnd.n7015 99.6594
R6390 gnd.n7175 gnd.n7016 99.6594
R6391 gnd.n7179 gnd.n7017 99.6594
R6392 gnd.n7183 gnd.n7018 99.6594
R6393 gnd.n7187 gnd.n7019 99.6594
R6394 gnd.n7191 gnd.n7020 99.6594
R6395 gnd.n7022 gnd.n7021 99.6594
R6396 gnd.n3988 gnd.n3987 99.6594
R6397 gnd.n3442 gnd.n3399 99.6594
R6398 gnd.n3444 gnd.n3400 99.6594
R6399 gnd.n3449 gnd.n3401 99.6594
R6400 gnd.n3451 gnd.n3402 99.6594
R6401 gnd.n3462 gnd.n3403 99.6594
R6402 gnd.n3464 gnd.n3404 99.6594
R6403 gnd.n3472 gnd.n3405 99.6594
R6404 gnd.n3482 gnd.n3406 99.6594
R6405 gnd.n3484 gnd.n3407 99.6594
R6406 gnd.n3492 gnd.n3408 99.6594
R6407 gnd.n3502 gnd.n3409 99.6594
R6408 gnd.n3513 gnd.n3410 99.6594
R6409 gnd.n3990 gnd.n3397 99.6594
R6410 gnd.n3988 gnd.n3413 99.6594
R6411 gnd.n3443 gnd.n3399 99.6594
R6412 gnd.n3448 gnd.n3400 99.6594
R6413 gnd.n3450 gnd.n3401 99.6594
R6414 gnd.n3461 gnd.n3402 99.6594
R6415 gnd.n3463 gnd.n3403 99.6594
R6416 gnd.n3471 gnd.n3404 99.6594
R6417 gnd.n3481 gnd.n3405 99.6594
R6418 gnd.n3483 gnd.n3406 99.6594
R6419 gnd.n3491 gnd.n3407 99.6594
R6420 gnd.n3501 gnd.n3408 99.6594
R6421 gnd.n3503 gnd.n3409 99.6594
R6422 gnd.n3515 gnd.n3410 99.6594
R6423 gnd.n3991 gnd.n3990 99.6594
R6424 gnd.n5031 gnd.n2733 99.6594
R6425 gnd.n5035 gnd.n2734 99.6594
R6426 gnd.n5038 gnd.n2735 99.6594
R6427 gnd.n2877 gnd.n2736 99.6594
R6428 gnd.n2879 gnd.n2737 99.6594
R6429 gnd.n5200 gnd.n2738 99.6594
R6430 gnd.n5210 gnd.n2739 99.6594
R6431 gnd.n5212 gnd.n2740 99.6594
R6432 gnd.n5220 gnd.n2741 99.6594
R6433 gnd.n5230 gnd.n2742 99.6594
R6434 gnd.n5232 gnd.n2743 99.6594
R6435 gnd.n2747 gnd.n2744 99.6594
R6436 gnd.n2748 gnd.n2745 99.6594
R6437 gnd.n5409 gnd.n2731 99.6594
R6438 gnd.n5233 gnd.n2744 99.6594
R6439 gnd.n5231 gnd.n2743 99.6594
R6440 gnd.n5221 gnd.n2742 99.6594
R6441 gnd.n5213 gnd.n2741 99.6594
R6442 gnd.n5211 gnd.n2740 99.6594
R6443 gnd.n5201 gnd.n2739 99.6594
R6444 gnd.n2880 gnd.n2738 99.6594
R6445 gnd.n2878 gnd.n2737 99.6594
R6446 gnd.n5037 gnd.n2736 99.6594
R6447 gnd.n5036 gnd.n2735 99.6594
R6448 gnd.n5032 gnd.n2734 99.6594
R6449 gnd.n2903 gnd.n2733 99.6594
R6450 gnd.n5410 gnd.n5409 99.6594
R6451 gnd.n2761 gnd.n2745 99.6594
R6452 gnd.n3504 gnd.t249 98.63
R6453 gnd.n5400 gnd.t209 98.63
R6454 gnd.n6877 gnd.t229 98.63
R6455 gnd.n7060 gnd.t264 98.63
R6456 gnd.n7159 gnd.t276 98.63
R6457 gnd.n2826 gnd.t292 98.63
R6458 gnd.n2849 gnd.t295 98.63
R6459 gnd.n2871 gnd.t255 98.63
R6460 gnd.n6892 gnd.t195 98.63
R6461 gnd.n3509 gnd.t244 98.63
R6462 gnd.n3673 gnd.t238 98.63
R6463 gnd.n2215 gnd.t252 98.63
R6464 gnd.n2237 gnd.t274 98.63
R6465 gnd.n2259 gnd.t286 98.63
R6466 gnd.n2531 gnd.t267 98.63
R6467 gnd.n3521 gnd.t288 98.63
R6468 gnd.n3533 gnd.t307 98.63
R6469 gnd.n2750 gnd.t216 98.63
R6470 gnd.n4063 gnd.t298 96.6984
R6471 gnd.n2973 gnd.t223 96.6984
R6472 gnd.n5555 gnd.t234 96.6906
R6473 gnd.n4840 gnd.t279 96.6906
R6474 gnd.n2592 gnd.n2591 81.8399
R6475 gnd.n1336 gnd.t258 74.8376
R6476 gnd.n785 gnd.t312 74.8376
R6477 gnd.n4064 gnd.t297 72.8438
R6478 gnd.n2974 gnd.t224 72.8438
R6479 gnd.n2593 gnd.n2586 72.8411
R6480 gnd.n2599 gnd.n2584 72.8411
R6481 gnd.n4836 gnd.n4835 72.8411
R6482 gnd.n3505 gnd.t248 72.836
R6483 gnd.n5556 gnd.t233 72.836
R6484 gnd.n4841 gnd.t280 72.836
R6485 gnd.n5401 gnd.t208 72.836
R6486 gnd.n6878 gnd.t230 72.836
R6487 gnd.n7061 gnd.t265 72.836
R6488 gnd.n7160 gnd.t277 72.836
R6489 gnd.n2827 gnd.t291 72.836
R6490 gnd.n2850 gnd.t294 72.836
R6491 gnd.n2872 gnd.t254 72.836
R6492 gnd.n6893 gnd.t196 72.836
R6493 gnd.n3510 gnd.t245 72.836
R6494 gnd.n3674 gnd.t237 72.836
R6495 gnd.n2216 gnd.t251 72.836
R6496 gnd.n2238 gnd.t273 72.836
R6497 gnd.n2260 gnd.t285 72.836
R6498 gnd.n2532 gnd.t268 72.836
R6499 gnd.n3522 gnd.t289 72.836
R6500 gnd.n3534 gnd.t308 72.836
R6501 gnd.n2751 gnd.t217 72.836
R6502 gnd.n4904 gnd.n2939 71.676
R6503 gnd.n4900 gnd.n2940 71.676
R6504 gnd.n4896 gnd.n2941 71.676
R6505 gnd.n4892 gnd.n2942 71.676
R6506 gnd.n4888 gnd.n2943 71.676
R6507 gnd.n4884 gnd.n2944 71.676
R6508 gnd.n4880 gnd.n2945 71.676
R6509 gnd.n4876 gnd.n2946 71.676
R6510 gnd.n4872 gnd.n2947 71.676
R6511 gnd.n4868 gnd.n2948 71.676
R6512 gnd.n4864 gnd.n2949 71.676
R6513 gnd.n4860 gnd.n2950 71.676
R6514 gnd.n4856 gnd.n2951 71.676
R6515 gnd.n4852 gnd.n2952 71.676
R6516 gnd.n4847 gnd.n2953 71.676
R6517 gnd.n4843 gnd.n2954 71.676
R6518 gnd.n4977 gnd.n2972 71.676
R6519 gnd.n4973 gnd.n2971 71.676
R6520 gnd.n4968 gnd.n2970 71.676
R6521 gnd.n4964 gnd.n2969 71.676
R6522 gnd.n4960 gnd.n2968 71.676
R6523 gnd.n4956 gnd.n2967 71.676
R6524 gnd.n4952 gnd.n2966 71.676
R6525 gnd.n4948 gnd.n2965 71.676
R6526 gnd.n4944 gnd.n2964 71.676
R6527 gnd.n4940 gnd.n2963 71.676
R6528 gnd.n4936 gnd.n2962 71.676
R6529 gnd.n4932 gnd.n2961 71.676
R6530 gnd.n4928 gnd.n2960 71.676
R6531 gnd.n4924 gnd.n2959 71.676
R6532 gnd.n4920 gnd.n2958 71.676
R6533 gnd.n4916 gnd.n2957 71.676
R6534 gnd.n4912 gnd.n2956 71.676
R6535 gnd.n5619 gnd.n5618 71.676
R6536 gnd.n5613 gnd.n2548 71.676
R6537 gnd.n5610 gnd.n2549 71.676
R6538 gnd.n5606 gnd.n2550 71.676
R6539 gnd.n5602 gnd.n2551 71.676
R6540 gnd.n5598 gnd.n2552 71.676
R6541 gnd.n5594 gnd.n2553 71.676
R6542 gnd.n5590 gnd.n2554 71.676
R6543 gnd.n5586 gnd.n2555 71.676
R6544 gnd.n5582 gnd.n2556 71.676
R6545 gnd.n5578 gnd.n2557 71.676
R6546 gnd.n5574 gnd.n2558 71.676
R6547 gnd.n5570 gnd.n2559 71.676
R6548 gnd.n5566 gnd.n2560 71.676
R6549 gnd.n5562 gnd.n2561 71.676
R6550 gnd.n5558 gnd.n2562 71.676
R6551 gnd.n2563 gnd.n2547 71.676
R6552 gnd.n4067 gnd.n2564 71.676
R6553 gnd.n4072 gnd.n2565 71.676
R6554 gnd.n4076 gnd.n2566 71.676
R6555 gnd.n4080 gnd.n2567 71.676
R6556 gnd.n4084 gnd.n2568 71.676
R6557 gnd.n4088 gnd.n2569 71.676
R6558 gnd.n4092 gnd.n2570 71.676
R6559 gnd.n4096 gnd.n2571 71.676
R6560 gnd.n4100 gnd.n2572 71.676
R6561 gnd.n4104 gnd.n2573 71.676
R6562 gnd.n4108 gnd.n2574 71.676
R6563 gnd.n4112 gnd.n2575 71.676
R6564 gnd.n4116 gnd.n2576 71.676
R6565 gnd.n4120 gnd.n2577 71.676
R6566 gnd.n4124 gnd.n2578 71.676
R6567 gnd.n5619 gnd.n2581 71.676
R6568 gnd.n5611 gnd.n2548 71.676
R6569 gnd.n5607 gnd.n2549 71.676
R6570 gnd.n5603 gnd.n2550 71.676
R6571 gnd.n5599 gnd.n2551 71.676
R6572 gnd.n5595 gnd.n2552 71.676
R6573 gnd.n5591 gnd.n2553 71.676
R6574 gnd.n5587 gnd.n2554 71.676
R6575 gnd.n5583 gnd.n2555 71.676
R6576 gnd.n5579 gnd.n2556 71.676
R6577 gnd.n5575 gnd.n2557 71.676
R6578 gnd.n5571 gnd.n2558 71.676
R6579 gnd.n5567 gnd.n2559 71.676
R6580 gnd.n5563 gnd.n2560 71.676
R6581 gnd.n5559 gnd.n2561 71.676
R6582 gnd.n5622 gnd.n5621 71.676
R6583 gnd.n4066 gnd.n2563 71.676
R6584 gnd.n4071 gnd.n2564 71.676
R6585 gnd.n4075 gnd.n2565 71.676
R6586 gnd.n4079 gnd.n2566 71.676
R6587 gnd.n4083 gnd.n2567 71.676
R6588 gnd.n4087 gnd.n2568 71.676
R6589 gnd.n4091 gnd.n2569 71.676
R6590 gnd.n4095 gnd.n2570 71.676
R6591 gnd.n4099 gnd.n2571 71.676
R6592 gnd.n4103 gnd.n2572 71.676
R6593 gnd.n4107 gnd.n2573 71.676
R6594 gnd.n4111 gnd.n2574 71.676
R6595 gnd.n4115 gnd.n2575 71.676
R6596 gnd.n4119 gnd.n2576 71.676
R6597 gnd.n4123 gnd.n2577 71.676
R6598 gnd.n4127 gnd.n2578 71.676
R6599 gnd.n4915 gnd.n2956 71.676
R6600 gnd.n4919 gnd.n2957 71.676
R6601 gnd.n4923 gnd.n2958 71.676
R6602 gnd.n4927 gnd.n2959 71.676
R6603 gnd.n4931 gnd.n2960 71.676
R6604 gnd.n4935 gnd.n2961 71.676
R6605 gnd.n4939 gnd.n2962 71.676
R6606 gnd.n4943 gnd.n2963 71.676
R6607 gnd.n4947 gnd.n2964 71.676
R6608 gnd.n4951 gnd.n2965 71.676
R6609 gnd.n4955 gnd.n2966 71.676
R6610 gnd.n4959 gnd.n2967 71.676
R6611 gnd.n4963 gnd.n2968 71.676
R6612 gnd.n4967 gnd.n2969 71.676
R6613 gnd.n4972 gnd.n2970 71.676
R6614 gnd.n4976 gnd.n2971 71.676
R6615 gnd.n4842 gnd.n2955 71.676
R6616 gnd.n4846 gnd.n2954 71.676
R6617 gnd.n4851 gnd.n2953 71.676
R6618 gnd.n4855 gnd.n2952 71.676
R6619 gnd.n4859 gnd.n2951 71.676
R6620 gnd.n4863 gnd.n2950 71.676
R6621 gnd.n4867 gnd.n2949 71.676
R6622 gnd.n4871 gnd.n2948 71.676
R6623 gnd.n4875 gnd.n2947 71.676
R6624 gnd.n4879 gnd.n2946 71.676
R6625 gnd.n4883 gnd.n2945 71.676
R6626 gnd.n4887 gnd.n2944 71.676
R6627 gnd.n4891 gnd.n2943 71.676
R6628 gnd.n4895 gnd.n2942 71.676
R6629 gnd.n4899 gnd.n2941 71.676
R6630 gnd.n4903 gnd.n2940 71.676
R6631 gnd.n2978 gnd.n2939 71.676
R6632 gnd.n10 gnd.t168 69.1507
R6633 gnd.n18 gnd.t97 68.4792
R6634 gnd.n17 gnd.t119 68.4792
R6635 gnd.n16 gnd.t166 68.4792
R6636 gnd.n15 gnd.t33 68.4792
R6637 gnd.n14 gnd.t139 68.4792
R6638 gnd.n13 gnd.t18 68.4792
R6639 gnd.n12 gnd.t317 68.4792
R6640 gnd.n11 gnd.t68 68.4792
R6641 gnd.n10 gnd.t137 68.4792
R6642 gnd.n1463 gnd.n1367 64.369
R6643 gnd.n5928 gnd.n2193 63.0944
R6644 gnd.n7199 gnd.n165 63.0944
R6645 gnd.n6729 gnd.n135 60.2057
R6646 gnd.n4069 gnd.n4064 59.5399
R6647 gnd.n4970 gnd.n2974 59.5399
R6648 gnd.n5557 gnd.n5556 59.5399
R6649 gnd.n4849 gnd.n4841 59.5399
R6650 gnd.n5554 gnd.n2602 59.1804
R6651 gnd.n5975 gnd.n776 57.3586
R6652 gnd.n1162 gnd.t143 56.407
R6653 gnd.n1127 gnd.t320 56.407
R6654 gnd.n1138 gnd.t334 56.407
R6655 gnd.n1150 gnd.t70 56.407
R6656 gnd.n56 gnd.t180 56.407
R6657 gnd.n21 gnd.t155 56.407
R6658 gnd.n32 gnd.t173 56.407
R6659 gnd.n44 gnd.t27 56.407
R6660 gnd.n1171 gnd.t81 55.8337
R6661 gnd.n1136 gnd.t169 55.8337
R6662 gnd.n1147 gnd.t131 55.8337
R6663 gnd.n1159 gnd.t20 55.8337
R6664 gnd.n65 gnd.t125 55.8337
R6665 gnd.n30 gnd.t172 55.8337
R6666 gnd.n41 gnd.t76 55.8337
R6667 gnd.n53 gnd.t126 55.8337
R6668 gnd.n2590 gnd.n2589 54.358
R6669 gnd.n4833 gnd.n4832 54.358
R6670 gnd.n1162 gnd.n1161 53.0052
R6671 gnd.n1164 gnd.n1163 53.0052
R6672 gnd.n1166 gnd.n1165 53.0052
R6673 gnd.n1168 gnd.n1167 53.0052
R6674 gnd.n1170 gnd.n1169 53.0052
R6675 gnd.n1127 gnd.n1126 53.0052
R6676 gnd.n1129 gnd.n1128 53.0052
R6677 gnd.n1131 gnd.n1130 53.0052
R6678 gnd.n1133 gnd.n1132 53.0052
R6679 gnd.n1135 gnd.n1134 53.0052
R6680 gnd.n1138 gnd.n1137 53.0052
R6681 gnd.n1140 gnd.n1139 53.0052
R6682 gnd.n1142 gnd.n1141 53.0052
R6683 gnd.n1144 gnd.n1143 53.0052
R6684 gnd.n1146 gnd.n1145 53.0052
R6685 gnd.n1150 gnd.n1149 53.0052
R6686 gnd.n1152 gnd.n1151 53.0052
R6687 gnd.n1154 gnd.n1153 53.0052
R6688 gnd.n1156 gnd.n1155 53.0052
R6689 gnd.n1158 gnd.n1157 53.0052
R6690 gnd.n64 gnd.n63 53.0052
R6691 gnd.n62 gnd.n61 53.0052
R6692 gnd.n60 gnd.n59 53.0052
R6693 gnd.n58 gnd.n57 53.0052
R6694 gnd.n56 gnd.n55 53.0052
R6695 gnd.n29 gnd.n28 53.0052
R6696 gnd.n27 gnd.n26 53.0052
R6697 gnd.n25 gnd.n24 53.0052
R6698 gnd.n23 gnd.n22 53.0052
R6699 gnd.n21 gnd.n20 53.0052
R6700 gnd.n40 gnd.n39 53.0052
R6701 gnd.n38 gnd.n37 53.0052
R6702 gnd.n36 gnd.n35 53.0052
R6703 gnd.n34 gnd.n33 53.0052
R6704 gnd.n32 gnd.n31 53.0052
R6705 gnd.n52 gnd.n51 53.0052
R6706 gnd.n50 gnd.n49 53.0052
R6707 gnd.n48 gnd.n47 53.0052
R6708 gnd.n46 gnd.n45 53.0052
R6709 gnd.n44 gnd.n43 53.0052
R6710 gnd.n4824 gnd.n4823 52.4801
R6711 gnd.n2107 gnd.t109 52.3082
R6712 gnd.n2075 gnd.t12 52.3082
R6713 gnd.n2043 gnd.t332 52.3082
R6714 gnd.n2012 gnd.t25 52.3082
R6715 gnd.n1980 gnd.t150 52.3082
R6716 gnd.n1948 gnd.t49 52.3082
R6717 gnd.n1916 gnd.t7 52.3082
R6718 gnd.n1885 gnd.t74 52.3082
R6719 gnd.n1937 gnd.n1905 51.4173
R6720 gnd.n2001 gnd.n2000 50.455
R6721 gnd.n1969 gnd.n1968 50.455
R6722 gnd.n1937 gnd.n1936 50.455
R6723 gnd.n1410 gnd.n1409 45.1884
R6724 gnd.n806 gnd.n805 45.1884
R6725 gnd.n4907 gnd.n4839 44.3322
R6726 gnd.n2593 gnd.n2592 44.3189
R6727 gnd.n3506 gnd.n3505 42.4732
R6728 gnd.n2752 gnd.n2751 42.4732
R6729 gnd.n5402 gnd.n5401 42.2793
R6730 gnd.n6879 gnd.n6878 42.2793
R6731 gnd.n7119 gnd.n7061 42.2793
R6732 gnd.n7161 gnd.n7160 42.2793
R6733 gnd.n5361 gnd.n2827 42.2793
R6734 gnd.n5324 gnd.n2850 42.2793
R6735 gnd.n5284 gnd.n2872 42.2793
R6736 gnd.n6894 gnd.n6893 42.2793
R6737 gnd.n1411 gnd.n1410 42.2793
R6738 gnd.n807 gnd.n806 42.2793
R6739 gnd.n1337 gnd.n1336 42.2793
R6740 gnd.n786 gnd.n785 42.2793
R6741 gnd.n3928 gnd.n3510 42.2793
R6742 gnd.n3724 gnd.n3674 42.2793
R6743 gnd.n5892 gnd.n2216 42.2793
R6744 gnd.n5852 gnd.n2238 42.2793
R6745 gnd.n5812 gnd.n2260 42.2793
R6746 gnd.n5641 gnd.n2532 42.2793
R6747 gnd.n3523 gnd.n3522 42.2793
R6748 gnd.n3535 gnd.n3534 42.2793
R6749 gnd.n2591 gnd.n2590 41.6274
R6750 gnd.n4834 gnd.n4833 41.6274
R6751 gnd.n2600 gnd.n2599 40.8975
R6752 gnd.n4837 gnd.n4836 40.8975
R6753 gnd.n2599 gnd.n2598 35.055
R6754 gnd.n2594 gnd.n2593 35.055
R6755 gnd.n4826 gnd.n4825 35.055
R6756 gnd.n4836 gnd.n4822 35.055
R6757 gnd.n6167 gnd.n6166 33.9721
R6758 gnd.n6166 gnd.n595 33.9721
R6759 gnd.n6160 gnd.n595 33.9721
R6760 gnd.n6160 gnd.n6159 33.9721
R6761 gnd.n6159 gnd.n6158 33.9721
R6762 gnd.n6158 gnd.n603 33.9721
R6763 gnd.n6152 gnd.n603 33.9721
R6764 gnd.n6152 gnd.n6151 33.9721
R6765 gnd.n6151 gnd.n6150 33.9721
R6766 gnd.n6150 gnd.n611 33.9721
R6767 gnd.n6144 gnd.n611 33.9721
R6768 gnd.n6144 gnd.n6143 33.9721
R6769 gnd.n6143 gnd.n6142 33.9721
R6770 gnd.n6142 gnd.n619 33.9721
R6771 gnd.n6136 gnd.n619 33.9721
R6772 gnd.n6136 gnd.n6135 33.9721
R6773 gnd.n6135 gnd.n6134 33.9721
R6774 gnd.n6134 gnd.n627 33.9721
R6775 gnd.n6128 gnd.n627 33.9721
R6776 gnd.n6128 gnd.n6127 33.9721
R6777 gnd.n6127 gnd.n6126 33.9721
R6778 gnd.n6126 gnd.n635 33.9721
R6779 gnd.n6120 gnd.n635 33.9721
R6780 gnd.n6120 gnd.n6119 33.9721
R6781 gnd.n6119 gnd.n6118 33.9721
R6782 gnd.n6118 gnd.n643 33.9721
R6783 gnd.n6112 gnd.n643 33.9721
R6784 gnd.n6112 gnd.n6111 33.9721
R6785 gnd.n6111 gnd.n6110 33.9721
R6786 gnd.n6110 gnd.n651 33.9721
R6787 gnd.n6104 gnd.n651 33.9721
R6788 gnd.n6104 gnd.n6103 33.9721
R6789 gnd.n6103 gnd.n6102 33.9721
R6790 gnd.n6102 gnd.n659 33.9721
R6791 gnd.n6096 gnd.n659 33.9721
R6792 gnd.n6096 gnd.n6095 33.9721
R6793 gnd.n6095 gnd.n6094 33.9721
R6794 gnd.n6094 gnd.n667 33.9721
R6795 gnd.n6088 gnd.n667 33.9721
R6796 gnd.n6088 gnd.n6087 33.9721
R6797 gnd.n6087 gnd.n6086 33.9721
R6798 gnd.n6086 gnd.n675 33.9721
R6799 gnd.n6080 gnd.n675 33.9721
R6800 gnd.n6080 gnd.n6079 33.9721
R6801 gnd.n6079 gnd.n6078 33.9721
R6802 gnd.n6078 gnd.n683 33.9721
R6803 gnd.n6072 gnd.n683 33.9721
R6804 gnd.n6072 gnd.n6071 33.9721
R6805 gnd.n6071 gnd.n6070 33.9721
R6806 gnd.n6070 gnd.n691 33.9721
R6807 gnd.n6064 gnd.n691 33.9721
R6808 gnd.n6064 gnd.n6063 33.9721
R6809 gnd.n6063 gnd.n6062 33.9721
R6810 gnd.n6062 gnd.n699 33.9721
R6811 gnd.n6056 gnd.n699 33.9721
R6812 gnd.n6056 gnd.n6055 33.9721
R6813 gnd.n6055 gnd.n6054 33.9721
R6814 gnd.n6054 gnd.n707 33.9721
R6815 gnd.n6048 gnd.n707 33.9721
R6816 gnd.n6048 gnd.n6047 33.9721
R6817 gnd.n6047 gnd.n6046 33.9721
R6818 gnd.n6046 gnd.n715 33.9721
R6819 gnd.n6040 gnd.n715 33.9721
R6820 gnd.n6040 gnd.n6039 33.9721
R6821 gnd.n6039 gnd.n6038 33.9721
R6822 gnd.n6038 gnd.n723 33.9721
R6823 gnd.n6032 gnd.n723 33.9721
R6824 gnd.n6032 gnd.n6031 33.9721
R6825 gnd.n6031 gnd.n6030 33.9721
R6826 gnd.n6030 gnd.n731 33.9721
R6827 gnd.n6024 gnd.n731 33.9721
R6828 gnd.n6024 gnd.n6023 33.9721
R6829 gnd.n6023 gnd.n6022 33.9721
R6830 gnd.n6022 gnd.n739 33.9721
R6831 gnd.n6016 gnd.n739 33.9721
R6832 gnd.n6016 gnd.n6015 33.9721
R6833 gnd.n6015 gnd.n6014 33.9721
R6834 gnd.n6014 gnd.n747 33.9721
R6835 gnd.n6008 gnd.n747 33.9721
R6836 gnd.n6008 gnd.n6007 33.9721
R6837 gnd.n6007 gnd.n6006 33.9721
R6838 gnd.n6006 gnd.n755 33.9721
R6839 gnd.n6000 gnd.n755 33.9721
R6840 gnd.n4913 gnd.n2975 32.9371
R6841 gnd.n4129 gnd.n4126 32.9371
R6842 gnd.n1473 gnd.n1367 31.8661
R6843 gnd.n1473 gnd.n1472 31.8661
R6844 gnd.n1481 gnd.n1356 31.8661
R6845 gnd.n1489 gnd.n1356 31.8661
R6846 gnd.n1489 gnd.n1350 31.8661
R6847 gnd.n1497 gnd.n1350 31.8661
R6848 gnd.n1497 gnd.n1343 31.8661
R6849 gnd.n1535 gnd.n1343 31.8661
R6850 gnd.n1545 gnd.n1276 31.8661
R6851 gnd.n5804 gnd.n2193 31.8661
R6852 gnd.n5796 gnd.n2278 31.8661
R6853 gnd.n5796 gnd.n2281 31.8661
R6854 gnd.n5790 gnd.n2281 31.8661
R6855 gnd.n5790 gnd.n2291 31.8661
R6856 gnd.n5784 gnd.n2300 31.8661
R6857 gnd.n5778 gnd.n2300 31.8661
R6858 gnd.n5772 gnd.n2316 31.8661
R6859 gnd.n5766 gnd.n2325 31.8661
R6860 gnd.n5766 gnd.n2328 31.8661
R6861 gnd.n5760 gnd.n2338 31.8661
R6862 gnd.n5754 gnd.n2338 31.8661
R6863 gnd.n5748 gnd.n2354 31.8661
R6864 gnd.n5742 gnd.n2363 31.8661
R6865 gnd.n5742 gnd.n2366 31.8661
R6866 gnd.n5736 gnd.n2376 31.8661
R6867 gnd.n5730 gnd.n2385 31.8661
R6868 gnd.n3923 gnd.n2474 31.8661
R6869 gnd.n3916 gnd.n2485 31.8661
R6870 gnd.n3916 gnd.n3398 31.8661
R6871 gnd.n3411 gnd.n3391 31.8661
R6872 gnd.n3998 gnd.n3391 31.8661
R6873 gnd.n4006 gnd.n3384 31.8661
R6874 gnd.n4006 gnd.n3376 31.8661
R6875 gnd.n4014 gnd.n3376 31.8661
R6876 gnd.n4014 gnd.n3378 31.8661
R6877 gnd.n4022 gnd.n3361 31.8661
R6878 gnd.n4042 gnd.n3361 31.8661
R6879 gnd.n4042 gnd.n3353 31.8661
R6880 gnd.n4053 gnd.n3353 31.8661
R6881 gnd.n4980 gnd.n2937 31.8661
R6882 gnd.n4988 gnd.n2931 31.8661
R6883 gnd.n4988 gnd.n2925 31.8661
R6884 gnd.n4998 gnd.n2925 31.8661
R6885 gnd.n4998 gnd.n4996 31.8661
R6886 gnd.n5006 gnd.n2914 31.8661
R6887 gnd.n5015 gnd.n2914 31.8661
R6888 gnd.n5015 gnd.n2908 31.8661
R6889 gnd.n5025 gnd.n2908 31.8661
R6890 gnd.n5051 gnd.n2901 31.8661
R6891 gnd.n5051 gnd.n2732 31.8661
R6892 gnd.n5059 gnd.n2746 31.8661
R6893 gnd.n5059 gnd.n2766 31.8661
R6894 gnd.n2886 gnd.n2804 31.8661
R6895 gnd.n6809 gnd.n195 31.8661
R6896 gnd.n6818 gnd.n189 31.8661
R6897 gnd.n6829 gnd.n172 31.8661
R6898 gnd.n6837 gnd.n172 31.8661
R6899 gnd.n7264 gnd.n74 31.8661
R6900 gnd.n7258 gnd.n86 31.8661
R6901 gnd.n7252 gnd.n86 31.8661
R6902 gnd.n7246 gnd.n104 31.8661
R6903 gnd.n7246 gnd.n107 31.8661
R6904 gnd.n7240 gnd.n116 31.8661
R6905 gnd.n7234 gnd.n126 31.8661
R6906 gnd.n7228 gnd.n126 31.8661
R6907 gnd.n7222 gnd.n143 31.8661
R6908 gnd.n7222 gnd.n146 31.8661
R6909 gnd.n7216 gnd.n146 31.8661
R6910 gnd.n7216 gnd.n155 31.8661
R6911 gnd.n7210 gnd.n165 31.8661
R6912 gnd.n2354 gnd.t45 31.5474
R6913 gnd.t121 gnd.n2376 31.5474
R6914 gnd.n6818 gnd.t62 31.5474
R6915 gnd.t79 gnd.n74 31.5474
R6916 gnd.n2316 gnd.t43 30.9101
R6917 gnd.t9 gnd.n116 30.9101
R6918 gnd.n2393 gnd.n2385 29.6355
R6919 gnd.n203 gnd.n195 29.6355
R6920 gnd.n3505 gnd.n3504 25.7944
R6921 gnd.n5401 gnd.n5400 25.7944
R6922 gnd.n6878 gnd.n6877 25.7944
R6923 gnd.n7061 gnd.n7060 25.7944
R6924 gnd.n7160 gnd.n7159 25.7944
R6925 gnd.n2827 gnd.n2826 25.7944
R6926 gnd.n2850 gnd.n2849 25.7944
R6927 gnd.n2872 gnd.n2871 25.7944
R6928 gnd.n6893 gnd.n6892 25.7944
R6929 gnd.n1336 gnd.n1335 25.7944
R6930 gnd.n785 gnd.n784 25.7944
R6931 gnd.n3510 gnd.n3509 25.7944
R6932 gnd.n3674 gnd.n3673 25.7944
R6933 gnd.n2216 gnd.n2215 25.7944
R6934 gnd.n2238 gnd.n2237 25.7944
R6935 gnd.n2260 gnd.n2259 25.7944
R6936 gnd.n2532 gnd.n2531 25.7944
R6937 gnd.n3522 gnd.n3521 25.7944
R6938 gnd.n3534 gnd.n3533 25.7944
R6939 gnd.n2751 gnd.n2750 25.7944
R6940 gnd.n1557 gnd.n1277 24.8557
R6941 gnd.n1567 gnd.n1260 24.8557
R6942 gnd.n1263 gnd.n1251 24.8557
R6943 gnd.n1588 gnd.n1252 24.8557
R6944 gnd.n1598 gnd.n1232 24.8557
R6945 gnd.n1608 gnd.n1607 24.8557
R6946 gnd.n1216 gnd.n1215 24.8557
R6947 gnd.n1645 gnd.n1208 24.8557
R6948 gnd.n1644 gnd.n1201 24.8557
R6949 gnd.n1682 gnd.n1180 24.8557
R6950 gnd.n1656 gnd.n1181 24.8557
R6951 gnd.n1675 gnd.n1045 24.8557
R6952 gnd.n1692 gnd.n1691 24.8557
R6953 gnd.n1703 gnd.n1702 24.8557
R6954 gnd.n1037 gnd.n1028 24.8557
R6955 gnd.n1723 gnd.n1011 24.8557
R6956 gnd.n1014 gnd.n1003 24.8557
R6957 gnd.n1744 gnd.n1004 24.8557
R6958 gnd.n1753 gnd.n996 24.8557
R6959 gnd.n1754 gnd.n985 24.8557
R6960 gnd.n988 gnd.n976 24.8557
R6961 gnd.n1775 gnd.n977 24.8557
R6962 gnd.n1785 gnd.n960 24.8557
R6963 gnd.n1796 gnd.n1795 24.8557
R6964 gnd.n1097 gnd.n1096 24.8557
R6965 gnd.n1806 gnd.n952 24.8557
R6966 gnd.n1816 gnd.n935 24.8557
R6967 gnd.n1827 gnd.n1826 24.8557
R6968 gnd.n1837 gnd.n927 24.8557
R6969 gnd.n1847 gnd.n909 24.8557
R6970 gnd.n1858 gnd.n1857 24.8557
R6971 gnd.n1869 gnd.n902 24.8557
R6972 gnd.n2134 gnd.n894 24.8557
R6973 gnd.n2135 gnd.n763 24.8557
R6974 gnd.n5992 gnd.n5991 24.8557
R6975 gnd.n3998 gnd.t247 24.537
R6976 gnd.t215 gnd.n2901 24.537
R6977 gnd.t270 gnd.n2579 24.2183
R6978 gnd.n3989 gnd.n3411 23.8997
R6979 gnd.n5408 gnd.n2732 23.8997
R6980 gnd.n4064 gnd.n4063 23.855
R6981 gnd.n2974 gnd.n2973 23.855
R6982 gnd.n5556 gnd.n5555 23.855
R6983 gnd.n4841 gnd.n4840 23.855
R6984 gnd.n1578 gnd.t73 23.2624
R6985 gnd.n1279 gnd.t257 22.6251
R6986 gnd.n5772 gnd.t36 21.9878
R6987 gnd.n7240 gnd.t54 21.9878
R6988 gnd.n5550 gnd.n2605 21.6691
R6989 gnd.n4140 gnd.n4137 21.6691
R6990 gnd.n4205 gnd.n3310 21.6691
R6991 gnd.n4288 gnd.n3275 21.6691
R6992 gnd.n4306 gnd.n3257 21.6691
R6993 gnd.n4344 gnd.n3236 21.6691
R6994 gnd.n4453 gnd.n3186 21.6691
R6995 gnd.n4493 gnd.n3172 21.6691
R6996 gnd.n4486 gnd.n3162 21.6691
R6997 gnd.n4525 gnd.n3154 21.6691
R6998 gnd.n4618 gnd.n3095 21.6691
R6999 gnd.n4666 gnd.n3078 21.6691
R7000 gnd.n4672 gnd.n3074 21.6691
R7001 gnd.n4772 gnd.n3009 21.6691
R7002 gnd.n4780 gnd.n4779 21.6691
R7003 gnd.n4800 gnd.n2995 21.6691
R7004 gnd.n4806 gnd.n2991 21.6691
R7005 gnd.t24 gnd.n1284 21.3504
R7006 gnd.n5748 gnd.t86 21.3504
R7007 gnd.n5736 gnd.t21 21.3504
R7008 gnd.n189 gnd.t140 21.3504
R7009 gnd.n7264 gnd.t52 21.3504
R7010 gnd.n4250 gnd.n3297 21.0318
R7011 gnd.n4260 gnd.n3290 21.0318
R7012 gnd.n4221 gnd.t85 21.0318
R7013 gnd.n4331 gnd.n3214 21.0318
R7014 gnd.n4315 gnd.n3215 21.0318
R7015 gnd.n4434 gnd.t91 21.0318
R7016 gnd.n4475 gnd.t110 21.0318
R7017 gnd.n4570 gnd.n3130 21.0318
R7018 gnd.n4577 gnd.n3124 21.0318
R7019 gnd.n4706 gnd.t51 21.0318
R7020 gnd.n4716 gnd.n4715 21.0318
R7021 gnd.n4725 gnd.n3035 21.0318
R7022 gnd.n5554 gnd.n5553 20.7615
R7023 gnd.n4908 gnd.n4907 20.7615
R7024 gnd.t39 gnd.n926 20.7131
R7025 gnd.n5760 gnd.t60 20.7131
R7026 gnd.n5724 gnd.t83 20.7131
R7027 gnd.n6796 gnd.t98 20.7131
R7028 gnd.n7252 gnd.t114 20.7131
R7029 gnd.n6000 gnd.n5999 20.3835
R7030 gnd.n1784 gnd.t23 20.0758
R7031 gnd.n5784 gnd.t19 20.0758
R7032 gnd.n2588 gnd.t202 19.8005
R7033 gnd.n2588 gnd.t227 19.8005
R7034 gnd.n2587 gnd.t305 19.8005
R7035 gnd.n2587 gnd.t205 19.8005
R7036 gnd.n4831 gnd.t262 19.8005
R7037 gnd.n4831 gnd.t199 19.8005
R7038 gnd.n4830 gnd.t241 19.8005
R7039 gnd.n4830 gnd.t220 19.8005
R7040 gnd.n5674 gnd.n2485 19.7572
R7041 gnd.n4204 gnd.n3313 19.7572
R7042 gnd.n4268 gnd.n3283 19.7572
R7043 gnd.n4382 gnd.n3222 19.7572
R7044 gnd.n4436 gnd.n3201 19.7572
R7045 gnd.n4474 gnd.n3138 19.7572
R7046 gnd.n4588 gnd.n4587 19.7572
R7047 gnd.n3058 gnd.n3056 19.7572
R7048 gnd.n4766 gnd.n4765 19.7572
R7049 gnd.n5397 gnd.n2766 19.7572
R7050 gnd.n2584 gnd.n2583 19.5087
R7051 gnd.n2597 gnd.n2584 19.5087
R7052 gnd.n2595 gnd.n2586 19.5087
R7053 gnd.n4835 gnd.n4829 19.5087
R7054 gnd.t102 gnd.n1733 19.4385
R7055 gnd.n3378 gnd.t1 19.4385
R7056 gnd.n5006 gnd.t96 19.4385
R7057 gnd.n3996 gnd.n3394 19.3944
R7058 gnd.n3996 gnd.n3382 19.3944
R7059 gnd.n4008 gnd.n3382 19.3944
R7060 gnd.n4008 gnd.n3380 19.3944
R7061 gnd.n4012 gnd.n3380 19.3944
R7062 gnd.n4012 gnd.n3368 19.3944
R7063 gnd.n4024 gnd.n3368 19.3944
R7064 gnd.n4024 gnd.n3365 19.3944
R7065 gnd.n4040 gnd.n3365 19.3944
R7066 gnd.n4040 gnd.n3366 19.3944
R7067 gnd.n4036 gnd.n3366 19.3944
R7068 gnd.n4036 gnd.n4035 19.3944
R7069 gnd.n4035 gnd.n4034 19.3944
R7070 gnd.n4034 gnd.n4031 19.3944
R7071 gnd.n4031 gnd.n2620 19.3944
R7072 gnd.n5541 gnd.n2620 19.3944
R7073 gnd.n5541 gnd.n2621 19.3944
R7074 gnd.n5537 gnd.n2621 19.3944
R7075 gnd.n5537 gnd.n5536 19.3944
R7076 gnd.n5536 gnd.n5535 19.3944
R7077 gnd.n5535 gnd.n2627 19.3944
R7078 gnd.n5531 gnd.n2627 19.3944
R7079 gnd.n5531 gnd.n5530 19.3944
R7080 gnd.n5530 gnd.n5529 19.3944
R7081 gnd.n5529 gnd.n2632 19.3944
R7082 gnd.n5525 gnd.n2632 19.3944
R7083 gnd.n5525 gnd.n5524 19.3944
R7084 gnd.n5524 gnd.n5523 19.3944
R7085 gnd.n5523 gnd.n2637 19.3944
R7086 gnd.n5519 gnd.n2637 19.3944
R7087 gnd.n5519 gnd.n5518 19.3944
R7088 gnd.n5518 gnd.n5517 19.3944
R7089 gnd.n5517 gnd.n2642 19.3944
R7090 gnd.n5513 gnd.n2642 19.3944
R7091 gnd.n5513 gnd.n5512 19.3944
R7092 gnd.n5512 gnd.n5511 19.3944
R7093 gnd.n5511 gnd.n2647 19.3944
R7094 gnd.n5507 gnd.n2647 19.3944
R7095 gnd.n5507 gnd.n5506 19.3944
R7096 gnd.n5506 gnd.n5505 19.3944
R7097 gnd.n5505 gnd.n2652 19.3944
R7098 gnd.n5501 gnd.n2652 19.3944
R7099 gnd.n5501 gnd.n5500 19.3944
R7100 gnd.n5500 gnd.n5499 19.3944
R7101 gnd.n5499 gnd.n2657 19.3944
R7102 gnd.n5495 gnd.n2657 19.3944
R7103 gnd.n5495 gnd.n5494 19.3944
R7104 gnd.n5494 gnd.n5493 19.3944
R7105 gnd.n5493 gnd.n2662 19.3944
R7106 gnd.n5489 gnd.n2662 19.3944
R7107 gnd.n5489 gnd.n5488 19.3944
R7108 gnd.n5488 gnd.n5487 19.3944
R7109 gnd.n5487 gnd.n2667 19.3944
R7110 gnd.n5483 gnd.n2667 19.3944
R7111 gnd.n5483 gnd.n5482 19.3944
R7112 gnd.n5482 gnd.n5481 19.3944
R7113 gnd.n5481 gnd.n2672 19.3944
R7114 gnd.n5477 gnd.n2672 19.3944
R7115 gnd.n5477 gnd.n5476 19.3944
R7116 gnd.n5476 gnd.n5475 19.3944
R7117 gnd.n5475 gnd.n2677 19.3944
R7118 gnd.n5471 gnd.n2677 19.3944
R7119 gnd.n5471 gnd.n5470 19.3944
R7120 gnd.n5470 gnd.n5469 19.3944
R7121 gnd.n5469 gnd.n2682 19.3944
R7122 gnd.n5465 gnd.n2682 19.3944
R7123 gnd.n5465 gnd.n5464 19.3944
R7124 gnd.n5464 gnd.n5463 19.3944
R7125 gnd.n5463 gnd.n2687 19.3944
R7126 gnd.n5459 gnd.n2687 19.3944
R7127 gnd.n5459 gnd.n5458 19.3944
R7128 gnd.n5458 gnd.n5457 19.3944
R7129 gnd.n5457 gnd.n2692 19.3944
R7130 gnd.n5453 gnd.n2692 19.3944
R7131 gnd.n5453 gnd.n5452 19.3944
R7132 gnd.n5452 gnd.n5451 19.3944
R7133 gnd.n5451 gnd.n2697 19.3944
R7134 gnd.n5447 gnd.n2697 19.3944
R7135 gnd.n5447 gnd.n5446 19.3944
R7136 gnd.n5446 gnd.n5445 19.3944
R7137 gnd.n5445 gnd.n2702 19.3944
R7138 gnd.n5441 gnd.n2702 19.3944
R7139 gnd.n5441 gnd.n5440 19.3944
R7140 gnd.n5440 gnd.n5439 19.3944
R7141 gnd.n5439 gnd.n2707 19.3944
R7142 gnd.n5435 gnd.n2707 19.3944
R7143 gnd.n5435 gnd.n5434 19.3944
R7144 gnd.n5434 gnd.n5433 19.3944
R7145 gnd.n5433 gnd.n2712 19.3944
R7146 gnd.n5429 gnd.n2712 19.3944
R7147 gnd.n5429 gnd.n5428 19.3944
R7148 gnd.n5428 gnd.n5427 19.3944
R7149 gnd.n5427 gnd.n2717 19.3944
R7150 gnd.n5423 gnd.n2717 19.3944
R7151 gnd.n5423 gnd.n5422 19.3944
R7152 gnd.n5422 gnd.n5421 19.3944
R7153 gnd.n5421 gnd.n2722 19.3944
R7154 gnd.n5417 gnd.n2722 19.3944
R7155 gnd.n5417 gnd.n5416 19.3944
R7156 gnd.n5416 gnd.n5415 19.3944
R7157 gnd.n5415 gnd.n2727 19.3944
R7158 gnd.n3516 gnd.n3514 19.3944
R7159 gnd.n3516 gnd.n3396 19.3944
R7160 gnd.n3992 gnd.n3396 19.3944
R7161 gnd.n3986 gnd.n3985 19.3944
R7162 gnd.n3985 gnd.n3440 19.3944
R7163 gnd.n3981 gnd.n3440 19.3944
R7164 gnd.n3981 gnd.n3980 19.3944
R7165 gnd.n3980 gnd.n3979 19.3944
R7166 gnd.n3979 gnd.n3445 19.3944
R7167 gnd.n3974 gnd.n3445 19.3944
R7168 gnd.n3974 gnd.n3973 19.3944
R7169 gnd.n3973 gnd.n3972 19.3944
R7170 gnd.n3972 gnd.n3452 19.3944
R7171 gnd.n3965 gnd.n3452 19.3944
R7172 gnd.n3965 gnd.n3964 19.3944
R7173 gnd.n3964 gnd.n3465 19.3944
R7174 gnd.n3957 gnd.n3465 19.3944
R7175 gnd.n3957 gnd.n3956 19.3944
R7176 gnd.n3956 gnd.n3473 19.3944
R7177 gnd.n3949 gnd.n3473 19.3944
R7178 gnd.n3949 gnd.n3948 19.3944
R7179 gnd.n3948 gnd.n3485 19.3944
R7180 gnd.n3941 gnd.n3485 19.3944
R7181 gnd.n3941 gnd.n3940 19.3944
R7182 gnd.n3940 gnd.n3493 19.3944
R7183 gnd.n3933 gnd.n3493 19.3944
R7184 gnd.n3933 gnd.n3932 19.3944
R7185 gnd.n5273 gnd.n5195 19.3944
R7186 gnd.n5273 gnd.n5272 19.3944
R7187 gnd.n5272 gnd.n5198 19.3944
R7188 gnd.n5265 gnd.n5198 19.3944
R7189 gnd.n5265 gnd.n5264 19.3944
R7190 gnd.n5264 gnd.n5208 19.3944
R7191 gnd.n5257 gnd.n5208 19.3944
R7192 gnd.n5257 gnd.n5256 19.3944
R7193 gnd.n5256 gnd.n5218 19.3944
R7194 gnd.n5249 gnd.n5218 19.3944
R7195 gnd.n5249 gnd.n5248 19.3944
R7196 gnd.n5248 gnd.n5228 19.3944
R7197 gnd.n5241 gnd.n5228 19.3944
R7198 gnd.n5241 gnd.n5240 19.3944
R7199 gnd.n5240 gnd.n2755 19.3944
R7200 gnd.n5403 gnd.n2755 19.3944
R7201 gnd.n5149 gnd.n5145 19.3944
R7202 gnd.n5149 gnd.n5148 19.3944
R7203 gnd.n5148 gnd.n5143 19.3944
R7204 gnd.n5158 gnd.n5143 19.3944
R7205 gnd.n5158 gnd.n5157 19.3944
R7206 gnd.n5157 gnd.n5100 19.3944
R7207 gnd.n5172 gnd.n5100 19.3944
R7208 gnd.n5172 gnd.n5105 19.3944
R7209 gnd.n5105 gnd.n5104 19.3944
R7210 gnd.n5104 gnd.n5101 19.3944
R7211 gnd.n5101 gnd.n220 19.3944
R7212 gnd.n6772 gnd.n220 19.3944
R7213 gnd.n6773 gnd.n6772 19.3944
R7214 gnd.n6776 gnd.n6773 19.3944
R7215 gnd.n6777 gnd.n6776 19.3944
R7216 gnd.n6777 gnd.n193 19.3944
R7217 gnd.n6811 gnd.n193 19.3944
R7218 gnd.n6814 gnd.n6811 19.3944
R7219 gnd.n6814 gnd.n6813 19.3944
R7220 gnd.n6813 gnd.n174 19.3944
R7221 gnd.n6834 gnd.n174 19.3944
R7222 gnd.n6835 gnd.n6834 19.3944
R7223 gnd.n6835 gnd.n168 19.3944
R7224 gnd.n6844 gnd.n168 19.3944
R7225 gnd.n6845 gnd.n6844 19.3944
R7226 gnd.n6847 gnd.n6845 19.3944
R7227 gnd.n6848 gnd.n6847 19.3944
R7228 gnd.n6851 gnd.n6848 19.3944
R7229 gnd.n6852 gnd.n6851 19.3944
R7230 gnd.n6854 gnd.n6852 19.3944
R7231 gnd.n6855 gnd.n6854 19.3944
R7232 gnd.n6858 gnd.n6855 19.3944
R7233 gnd.n6859 gnd.n6858 19.3944
R7234 gnd.n6861 gnd.n6859 19.3944
R7235 gnd.n6862 gnd.n6861 19.3944
R7236 gnd.n6865 gnd.n6862 19.3944
R7237 gnd.n6866 gnd.n6865 19.3944
R7238 gnd.n6868 gnd.n6866 19.3944
R7239 gnd.n6869 gnd.n6868 19.3944
R7240 gnd.n6872 gnd.n6869 19.3944
R7241 gnd.n6873 gnd.n6872 19.3944
R7242 gnd.n6874 gnd.n6873 19.3944
R7243 gnd.n7115 gnd.n7059 19.3944
R7244 gnd.n7115 gnd.n7112 19.3944
R7245 gnd.n7112 gnd.n7109 19.3944
R7246 gnd.n7109 gnd.n7108 19.3944
R7247 gnd.n7108 gnd.n7105 19.3944
R7248 gnd.n7105 gnd.n7104 19.3944
R7249 gnd.n7104 gnd.n7101 19.3944
R7250 gnd.n7101 gnd.n7100 19.3944
R7251 gnd.n7100 gnd.n7097 19.3944
R7252 gnd.n7097 gnd.n7096 19.3944
R7253 gnd.n7096 gnd.n7093 19.3944
R7254 gnd.n7093 gnd.n7092 19.3944
R7255 gnd.n7092 gnd.n7089 19.3944
R7256 gnd.n7089 gnd.n7088 19.3944
R7257 gnd.n7088 gnd.n7085 19.3944
R7258 gnd.n7085 gnd.n7084 19.3944
R7259 gnd.n7084 gnd.n7081 19.3944
R7260 gnd.n7081 gnd.n7080 19.3944
R7261 gnd.n7158 gnd.n7155 19.3944
R7262 gnd.n7155 gnd.n7154 19.3944
R7263 gnd.n7154 gnd.n7151 19.3944
R7264 gnd.n7151 gnd.n7150 19.3944
R7265 gnd.n7150 gnd.n7147 19.3944
R7266 gnd.n7147 gnd.n7146 19.3944
R7267 gnd.n7146 gnd.n7143 19.3944
R7268 gnd.n7143 gnd.n7142 19.3944
R7269 gnd.n7142 gnd.n7139 19.3944
R7270 gnd.n7139 gnd.n7138 19.3944
R7271 gnd.n7138 gnd.n7135 19.3944
R7272 gnd.n7135 gnd.n7134 19.3944
R7273 gnd.n7134 gnd.n7131 19.3944
R7274 gnd.n7131 gnd.n7130 19.3944
R7275 gnd.n7130 gnd.n7127 19.3944
R7276 gnd.n7127 gnd.n7126 19.3944
R7277 gnd.n7126 gnd.n7123 19.3944
R7278 gnd.n7123 gnd.n7122 19.3944
R7279 gnd.n7197 gnd.n7196 19.3944
R7280 gnd.n7196 gnd.n7025 19.3944
R7281 gnd.n7192 gnd.n7025 19.3944
R7282 gnd.n7192 gnd.n7189 19.3944
R7283 gnd.n7189 gnd.n7186 19.3944
R7284 gnd.n7186 gnd.n7185 19.3944
R7285 gnd.n7185 gnd.n7182 19.3944
R7286 gnd.n7182 gnd.n7181 19.3944
R7287 gnd.n7181 gnd.n7178 19.3944
R7288 gnd.n7178 gnd.n7177 19.3944
R7289 gnd.n7177 gnd.n7174 19.3944
R7290 gnd.n7174 gnd.n7173 19.3944
R7291 gnd.n7173 gnd.n7170 19.3944
R7292 gnd.n7170 gnd.n7169 19.3944
R7293 gnd.n7169 gnd.n7166 19.3944
R7294 gnd.n7166 gnd.n7165 19.3944
R7295 gnd.n7165 gnd.n7162 19.3944
R7296 gnd.n5083 gnd.n5081 19.3944
R7297 gnd.n5083 gnd.n5079 19.3944
R7298 gnd.n5182 gnd.n5079 19.3944
R7299 gnd.n5182 gnd.n5181 19.3944
R7300 gnd.n5181 gnd.n5180 19.3944
R7301 gnd.n5180 gnd.n5090 19.3944
R7302 gnd.n5090 gnd.n237 19.3944
R7303 gnd.n6753 gnd.n237 19.3944
R7304 gnd.n6753 gnd.n235 19.3944
R7305 gnd.n6759 gnd.n235 19.3944
R7306 gnd.n6759 gnd.n6758 19.3944
R7307 gnd.n6758 gnd.n209 19.3944
R7308 gnd.n6788 gnd.n209 19.3944
R7309 gnd.n6788 gnd.n207 19.3944
R7310 gnd.n6794 gnd.n207 19.3944
R7311 gnd.n6794 gnd.n6793 19.3944
R7312 gnd.n6793 gnd.n185 19.3944
R7313 gnd.n6820 gnd.n185 19.3944
R7314 gnd.n6820 gnd.n183 19.3944
R7315 gnd.n6827 gnd.n183 19.3944
R7316 gnd.n6827 gnd.n6826 19.3944
R7317 gnd.n6826 gnd.n78 19.3944
R7318 gnd.n7262 gnd.n78 19.3944
R7319 gnd.n7262 gnd.n7261 19.3944
R7320 gnd.n7261 gnd.n7260 19.3944
R7321 gnd.n7260 gnd.n82 19.3944
R7322 gnd.n7250 gnd.n82 19.3944
R7323 gnd.n7250 gnd.n7249 19.3944
R7324 gnd.n7249 gnd.n7248 19.3944
R7325 gnd.n7248 gnd.n102 19.3944
R7326 gnd.n7238 gnd.n102 19.3944
R7327 gnd.n7238 gnd.n7237 19.3944
R7328 gnd.n7237 gnd.n7236 19.3944
R7329 gnd.n7236 gnd.n122 19.3944
R7330 gnd.n7226 gnd.n122 19.3944
R7331 gnd.n7226 gnd.n7225 19.3944
R7332 gnd.n7225 gnd.n7224 19.3944
R7333 gnd.n7224 gnd.n141 19.3944
R7334 gnd.n7214 gnd.n141 19.3944
R7335 gnd.n7214 gnd.n7213 19.3944
R7336 gnd.n7213 gnd.n7212 19.3944
R7337 gnd.n7212 gnd.n161 19.3944
R7338 gnd.n5394 gnd.n5393 19.3944
R7339 gnd.n5393 gnd.n5392 19.3944
R7340 gnd.n5392 gnd.n5391 19.3944
R7341 gnd.n5391 gnd.n5389 19.3944
R7342 gnd.n5389 gnd.n5386 19.3944
R7343 gnd.n5386 gnd.n5385 19.3944
R7344 gnd.n5385 gnd.n5382 19.3944
R7345 gnd.n5382 gnd.n5381 19.3944
R7346 gnd.n5381 gnd.n5378 19.3944
R7347 gnd.n5378 gnd.n5377 19.3944
R7348 gnd.n5377 gnd.n5374 19.3944
R7349 gnd.n5374 gnd.n5373 19.3944
R7350 gnd.n5373 gnd.n5370 19.3944
R7351 gnd.n5370 gnd.n5369 19.3944
R7352 gnd.n5369 gnd.n5366 19.3944
R7353 gnd.n5366 gnd.n5365 19.3944
R7354 gnd.n5365 gnd.n5362 19.3944
R7355 gnd.n5360 gnd.n5357 19.3944
R7356 gnd.n5357 gnd.n5356 19.3944
R7357 gnd.n5356 gnd.n5353 19.3944
R7358 gnd.n5353 gnd.n5352 19.3944
R7359 gnd.n5352 gnd.n5349 19.3944
R7360 gnd.n5349 gnd.n5348 19.3944
R7361 gnd.n5348 gnd.n5345 19.3944
R7362 gnd.n5343 gnd.n5340 19.3944
R7363 gnd.n5340 gnd.n5339 19.3944
R7364 gnd.n5339 gnd.n5336 19.3944
R7365 gnd.n5336 gnd.n5335 19.3944
R7366 gnd.n5335 gnd.n5332 19.3944
R7367 gnd.n5332 gnd.n5331 19.3944
R7368 gnd.n5331 gnd.n5328 19.3944
R7369 gnd.n5328 gnd.n5327 19.3944
R7370 gnd.n5323 gnd.n5320 19.3944
R7371 gnd.n5320 gnd.n5319 19.3944
R7372 gnd.n5319 gnd.n5316 19.3944
R7373 gnd.n5316 gnd.n5315 19.3944
R7374 gnd.n5315 gnd.n5312 19.3944
R7375 gnd.n5312 gnd.n5311 19.3944
R7376 gnd.n5311 gnd.n5308 19.3944
R7377 gnd.n5308 gnd.n5307 19.3944
R7378 gnd.n5307 gnd.n5304 19.3944
R7379 gnd.n5304 gnd.n5303 19.3944
R7380 gnd.n5303 gnd.n5300 19.3944
R7381 gnd.n5300 gnd.n5299 19.3944
R7382 gnd.n5299 gnd.n5296 19.3944
R7383 gnd.n5296 gnd.n5295 19.3944
R7384 gnd.n5295 gnd.n5292 19.3944
R7385 gnd.n5292 gnd.n5291 19.3944
R7386 gnd.n5291 gnd.n5288 19.3944
R7387 gnd.n5288 gnd.n5287 19.3944
R7388 gnd.n6904 gnd.n6902 19.3944
R7389 gnd.n6907 gnd.n6904 19.3944
R7390 gnd.n6910 gnd.n6907 19.3944
R7391 gnd.n6913 gnd.n6910 19.3944
R7392 gnd.n6913 gnd.n6900 19.3944
R7393 gnd.n6917 gnd.n6900 19.3944
R7394 gnd.n6920 gnd.n6917 19.3944
R7395 gnd.n6923 gnd.n6920 19.3944
R7396 gnd.n6923 gnd.n6898 19.3944
R7397 gnd.n6927 gnd.n6898 19.3944
R7398 gnd.n6930 gnd.n6927 19.3944
R7399 gnd.n6933 gnd.n6930 19.3944
R7400 gnd.n6933 gnd.n6896 19.3944
R7401 gnd.n6937 gnd.n6896 19.3944
R7402 gnd.n6940 gnd.n6937 19.3944
R7403 gnd.n6942 gnd.n6940 19.3944
R7404 gnd.n5138 gnd.n5135 19.3944
R7405 gnd.n5138 gnd.n5133 19.3944
R7406 gnd.n5142 gnd.n5133 19.3944
R7407 gnd.n5162 gnd.n5142 19.3944
R7408 gnd.n5163 gnd.n5162 19.3944
R7409 gnd.n5163 gnd.n5130 19.3944
R7410 gnd.n5168 gnd.n5130 19.3944
R7411 gnd.n5168 gnd.n5131 19.3944
R7412 gnd.n5131 gnd.n227 19.3944
R7413 gnd.n6763 gnd.n227 19.3944
R7414 gnd.n6763 gnd.n224 19.3944
R7415 gnd.n6768 gnd.n224 19.3944
R7416 gnd.n6768 gnd.n225 19.3944
R7417 gnd.n225 gnd.n200 19.3944
R7418 gnd.n6798 gnd.n200 19.3944
R7419 gnd.n6798 gnd.n197 19.3944
R7420 gnd.n6807 gnd.n197 19.3944
R7421 gnd.n6807 gnd.n198 19.3944
R7422 gnd.n6803 gnd.n198 19.3944
R7423 gnd.n6803 gnd.n6802 19.3944
R7424 gnd.n6802 gnd.n68 19.3944
R7425 gnd.n7267 gnd.n68 19.3944
R7426 gnd.n7267 gnd.n7266 19.3944
R7427 gnd.n7266 gnd.n71 19.3944
R7428 gnd.n6955 gnd.n71 19.3944
R7429 gnd.n6957 gnd.n6955 19.3944
R7430 gnd.n6957 gnd.n6952 19.3944
R7431 gnd.n6962 gnd.n6952 19.3944
R7432 gnd.n6963 gnd.n6962 19.3944
R7433 gnd.n6965 gnd.n6963 19.3944
R7434 gnd.n6965 gnd.n6950 19.3944
R7435 gnd.n6970 gnd.n6950 19.3944
R7436 gnd.n6971 gnd.n6970 19.3944
R7437 gnd.n6973 gnd.n6971 19.3944
R7438 gnd.n6973 gnd.n6948 19.3944
R7439 gnd.n6978 gnd.n6948 19.3944
R7440 gnd.n6979 gnd.n6978 19.3944
R7441 gnd.n6981 gnd.n6979 19.3944
R7442 gnd.n6981 gnd.n6946 19.3944
R7443 gnd.n6986 gnd.n6946 19.3944
R7444 gnd.n6987 gnd.n6986 19.3944
R7445 gnd.n6988 gnd.n6987 19.3944
R7446 gnd.n5151 gnd.n2885 19.3944
R7447 gnd.n5153 gnd.n5151 19.3944
R7448 gnd.n5154 gnd.n5153 19.3944
R7449 gnd.n5154 gnd.n5098 19.3944
R7450 gnd.n5176 gnd.n5098 19.3944
R7451 gnd.n5176 gnd.n5175 19.3944
R7452 gnd.n5175 gnd.n245 19.3944
R7453 gnd.n6749 gnd.n245 19.3944
R7454 gnd.n6749 gnd.n6748 19.3944
R7455 gnd.n6748 gnd.n6747 19.3944
R7456 gnd.n6747 gnd.n6746 19.3944
R7457 gnd.n6746 gnd.n217 19.3944
R7458 gnd.n6784 gnd.n217 19.3944
R7459 gnd.n6784 gnd.n6783 19.3944
R7460 gnd.n6783 gnd.n6782 19.3944
R7461 gnd.n6782 gnd.n6781 19.3944
R7462 gnd.n6781 gnd.n191 19.3944
R7463 gnd.n6816 gnd.n191 19.3944
R7464 gnd.n6816 gnd.n176 19.3944
R7465 gnd.n6831 gnd.n176 19.3944
R7466 gnd.n6831 gnd.n170 19.3944
R7467 gnd.n6839 gnd.n170 19.3944
R7468 gnd.n6840 gnd.n6839 19.3944
R7469 gnd.n6840 gnd.n89 19.3944
R7470 gnd.n7256 gnd.n89 19.3944
R7471 gnd.n7256 gnd.n7255 19.3944
R7472 gnd.n7255 gnd.n7254 19.3944
R7473 gnd.n7254 gnd.n93 19.3944
R7474 gnd.n7244 gnd.n93 19.3944
R7475 gnd.n7244 gnd.n7243 19.3944
R7476 gnd.n7243 gnd.n7242 19.3944
R7477 gnd.n7242 gnd.n112 19.3944
R7478 gnd.n7232 gnd.n112 19.3944
R7479 gnd.n7232 gnd.n7231 19.3944
R7480 gnd.n7231 gnd.n7230 19.3944
R7481 gnd.n7230 gnd.n131 19.3944
R7482 gnd.n7220 gnd.n131 19.3944
R7483 gnd.n7220 gnd.n7219 19.3944
R7484 gnd.n7219 gnd.n7218 19.3944
R7485 gnd.n7218 gnd.n151 19.3944
R7486 gnd.n7208 gnd.n151 19.3944
R7487 gnd.n7208 gnd.n7207 19.3944
R7488 gnd.n1460 gnd.n1459 19.3944
R7489 gnd.n1459 gnd.n1458 19.3944
R7490 gnd.n1458 gnd.n1457 19.3944
R7491 gnd.n1457 gnd.n1455 19.3944
R7492 gnd.n1455 gnd.n1452 19.3944
R7493 gnd.n1452 gnd.n1451 19.3944
R7494 gnd.n1451 gnd.n1448 19.3944
R7495 gnd.n1448 gnd.n1447 19.3944
R7496 gnd.n1447 gnd.n1444 19.3944
R7497 gnd.n1444 gnd.n1443 19.3944
R7498 gnd.n1443 gnd.n1440 19.3944
R7499 gnd.n1440 gnd.n1439 19.3944
R7500 gnd.n1439 gnd.n1436 19.3944
R7501 gnd.n1436 gnd.n1435 19.3944
R7502 gnd.n1435 gnd.n1432 19.3944
R7503 gnd.n1432 gnd.n1431 19.3944
R7504 gnd.n1431 gnd.n1428 19.3944
R7505 gnd.n1428 gnd.n1427 19.3944
R7506 gnd.n1427 gnd.n1424 19.3944
R7507 gnd.n1424 gnd.n1423 19.3944
R7508 gnd.n1423 gnd.n1420 19.3944
R7509 gnd.n1420 gnd.n1419 19.3944
R7510 gnd.n1416 gnd.n1415 19.3944
R7511 gnd.n1415 gnd.n1371 19.3944
R7512 gnd.n1466 gnd.n1371 19.3944
R7513 gnd.n879 gnd.n877 19.3944
R7514 gnd.n879 gnd.n803 19.3944
R7515 gnd.n2152 gnd.n803 19.3944
R7516 gnd.n820 gnd.n819 19.3944
R7517 gnd.n824 gnd.n819 19.3944
R7518 gnd.n827 gnd.n824 19.3944
R7519 gnd.n830 gnd.n827 19.3944
R7520 gnd.n830 gnd.n816 19.3944
R7521 gnd.n834 gnd.n816 19.3944
R7522 gnd.n837 gnd.n834 19.3944
R7523 gnd.n840 gnd.n837 19.3944
R7524 gnd.n840 gnd.n814 19.3944
R7525 gnd.n844 gnd.n814 19.3944
R7526 gnd.n847 gnd.n844 19.3944
R7527 gnd.n850 gnd.n847 19.3944
R7528 gnd.n850 gnd.n812 19.3944
R7529 gnd.n854 gnd.n812 19.3944
R7530 gnd.n857 gnd.n854 19.3944
R7531 gnd.n860 gnd.n857 19.3944
R7532 gnd.n860 gnd.n810 19.3944
R7533 gnd.n864 gnd.n810 19.3944
R7534 gnd.n867 gnd.n864 19.3944
R7535 gnd.n870 gnd.n867 19.3944
R7536 gnd.n870 gnd.n808 19.3944
R7537 gnd.n874 gnd.n808 19.3944
R7538 gnd.n1559 gnd.n1268 19.3944
R7539 gnd.n1569 gnd.n1268 19.3944
R7540 gnd.n1570 gnd.n1569 19.3944
R7541 gnd.n1570 gnd.n1249 19.3944
R7542 gnd.n1590 gnd.n1249 19.3944
R7543 gnd.n1590 gnd.n1241 19.3944
R7544 gnd.n1600 gnd.n1241 19.3944
R7545 gnd.n1601 gnd.n1600 19.3944
R7546 gnd.n1602 gnd.n1601 19.3944
R7547 gnd.n1602 gnd.n1224 19.3944
R7548 gnd.n1224 gnd.n1222 19.3944
R7549 gnd.n1628 gnd.n1222 19.3944
R7550 gnd.n1628 gnd.n1204 19.3944
R7551 gnd.n1662 gnd.n1204 19.3944
R7552 gnd.n1662 gnd.n1661 19.3944
R7553 gnd.n1661 gnd.n1660 19.3944
R7554 gnd.n1660 gnd.n1655 19.3944
R7555 gnd.n1655 gnd.n1042 19.3944
R7556 gnd.n1694 gnd.n1042 19.3944
R7557 gnd.n1695 gnd.n1694 19.3944
R7558 gnd.n1695 gnd.n1026 19.3944
R7559 gnd.n1715 gnd.n1026 19.3944
R7560 gnd.n1715 gnd.n1019 19.3944
R7561 gnd.n1725 gnd.n1019 19.3944
R7562 gnd.n1726 gnd.n1725 19.3944
R7563 gnd.n1726 gnd.n1001 19.3944
R7564 gnd.n1746 gnd.n1001 19.3944
R7565 gnd.n1746 gnd.n993 19.3944
R7566 gnd.n1756 gnd.n993 19.3944
R7567 gnd.n1757 gnd.n1756 19.3944
R7568 gnd.n1757 gnd.n974 19.3944
R7569 gnd.n1777 gnd.n974 19.3944
R7570 gnd.n1777 gnd.n967 19.3944
R7571 gnd.n1787 gnd.n967 19.3944
R7572 gnd.n1788 gnd.n1787 19.3944
R7573 gnd.n1788 gnd.n950 19.3944
R7574 gnd.n1808 gnd.n950 19.3944
R7575 gnd.n1808 gnd.n943 19.3944
R7576 gnd.n1818 gnd.n943 19.3944
R7577 gnd.n1819 gnd.n1818 19.3944
R7578 gnd.n1819 gnd.n924 19.3944
R7579 gnd.n1839 gnd.n924 19.3944
R7580 gnd.n1839 gnd.n917 19.3944
R7581 gnd.n1849 gnd.n917 19.3944
R7582 gnd.n1850 gnd.n1849 19.3944
R7583 gnd.n1850 gnd.n899 19.3944
R7584 gnd.n1871 gnd.n899 19.3944
R7585 gnd.n1871 gnd.n890 19.3944
R7586 gnd.n2137 gnd.n890 19.3944
R7587 gnd.n2138 gnd.n2137 19.3944
R7588 gnd.n2140 gnd.n2138 19.3944
R7589 gnd.n2140 gnd.n782 19.3944
R7590 gnd.n5986 gnd.n782 19.3944
R7591 gnd.n1550 gnd.n1549 19.3944
R7592 gnd.n1549 gnd.n1282 19.3944
R7593 gnd.n1305 gnd.n1282 19.3944
R7594 gnd.n1308 gnd.n1305 19.3944
R7595 gnd.n1308 gnd.n1301 19.3944
R7596 gnd.n1312 gnd.n1301 19.3944
R7597 gnd.n1315 gnd.n1312 19.3944
R7598 gnd.n1318 gnd.n1315 19.3944
R7599 gnd.n1318 gnd.n1299 19.3944
R7600 gnd.n1322 gnd.n1299 19.3944
R7601 gnd.n1325 gnd.n1322 19.3944
R7602 gnd.n1328 gnd.n1325 19.3944
R7603 gnd.n1328 gnd.n1297 19.3944
R7604 gnd.n1332 gnd.n1297 19.3944
R7605 gnd.n1555 gnd.n1554 19.3944
R7606 gnd.n1554 gnd.n1258 19.3944
R7607 gnd.n1580 gnd.n1258 19.3944
R7608 gnd.n1580 gnd.n1256 19.3944
R7609 gnd.n1586 gnd.n1256 19.3944
R7610 gnd.n1586 gnd.n1585 19.3944
R7611 gnd.n1585 gnd.n1230 19.3944
R7612 gnd.n1610 gnd.n1230 19.3944
R7613 gnd.n1610 gnd.n1228 19.3944
R7614 gnd.n1622 gnd.n1228 19.3944
R7615 gnd.n1622 gnd.n1621 19.3944
R7616 gnd.n1621 gnd.n1620 19.3944
R7617 gnd.n1620 gnd.n1618 19.3944
R7618 gnd.n1618 gnd.n1200 19.3944
R7619 gnd.n1200 gnd.n1198 19.3944
R7620 gnd.n1669 gnd.n1198 19.3944
R7621 gnd.n1669 gnd.n1196 19.3944
R7622 gnd.n1673 gnd.n1196 19.3944
R7623 gnd.n1673 gnd.n1033 19.3944
R7624 gnd.n1705 gnd.n1033 19.3944
R7625 gnd.n1705 gnd.n1031 19.3944
R7626 gnd.n1711 gnd.n1031 19.3944
R7627 gnd.n1711 gnd.n1710 19.3944
R7628 gnd.n1710 gnd.n1009 19.3944
R7629 gnd.n1736 gnd.n1009 19.3944
R7630 gnd.n1736 gnd.n1007 19.3944
R7631 gnd.n1742 gnd.n1007 19.3944
R7632 gnd.n1742 gnd.n1741 19.3944
R7633 gnd.n1741 gnd.n983 19.3944
R7634 gnd.n1767 gnd.n983 19.3944
R7635 gnd.n1767 gnd.n981 19.3944
R7636 gnd.n1773 gnd.n981 19.3944
R7637 gnd.n1773 gnd.n1772 19.3944
R7638 gnd.n1772 gnd.n958 19.3944
R7639 gnd.n1798 gnd.n958 19.3944
R7640 gnd.n1798 gnd.n956 19.3944
R7641 gnd.n1804 gnd.n956 19.3944
R7642 gnd.n1804 gnd.n1803 19.3944
R7643 gnd.n1803 gnd.n933 19.3944
R7644 gnd.n1829 gnd.n933 19.3944
R7645 gnd.n1829 gnd.n931 19.3944
R7646 gnd.n1835 gnd.n931 19.3944
R7647 gnd.n1835 gnd.n1834 19.3944
R7648 gnd.n1834 gnd.n907 19.3944
R7649 gnd.n1860 gnd.n907 19.3944
R7650 gnd.n1860 gnd.n905 19.3944
R7651 gnd.n1867 gnd.n905 19.3944
R7652 gnd.n1867 gnd.n1866 19.3944
R7653 gnd.n1866 gnd.n767 19.3944
R7654 gnd.n5996 gnd.n767 19.3944
R7655 gnd.n5996 gnd.n5995 19.3944
R7656 gnd.n5995 gnd.n5994 19.3944
R7657 gnd.n5994 gnd.n771 19.3944
R7658 gnd.n5973 gnd.n5972 19.3944
R7659 gnd.n5972 gnd.n5938 19.3944
R7660 gnd.n5968 gnd.n5938 19.3944
R7661 gnd.n5968 gnd.n5965 19.3944
R7662 gnd.n5965 gnd.n5962 19.3944
R7663 gnd.n5962 gnd.n5961 19.3944
R7664 gnd.n5961 gnd.n5958 19.3944
R7665 gnd.n5958 gnd.n5957 19.3944
R7666 gnd.n5957 gnd.n5954 19.3944
R7667 gnd.n5954 gnd.n5953 19.3944
R7668 gnd.n5953 gnd.n5950 19.3944
R7669 gnd.n5950 gnd.n5949 19.3944
R7670 gnd.n5949 gnd.n788 19.3944
R7671 gnd.n5979 gnd.n788 19.3944
R7672 gnd.n1470 gnd.n1369 19.3944
R7673 gnd.n1470 gnd.n1360 19.3944
R7674 gnd.n1483 gnd.n1360 19.3944
R7675 gnd.n1483 gnd.n1358 19.3944
R7676 gnd.n1487 gnd.n1358 19.3944
R7677 gnd.n1487 gnd.n1348 19.3944
R7678 gnd.n1499 gnd.n1348 19.3944
R7679 gnd.n1499 gnd.n1346 19.3944
R7680 gnd.n1533 gnd.n1346 19.3944
R7681 gnd.n1533 gnd.n1532 19.3944
R7682 gnd.n1532 gnd.n1531 19.3944
R7683 gnd.n1531 gnd.n1530 19.3944
R7684 gnd.n1530 gnd.n1527 19.3944
R7685 gnd.n1527 gnd.n1526 19.3944
R7686 gnd.n1526 gnd.n1525 19.3944
R7687 gnd.n1525 gnd.n1523 19.3944
R7688 gnd.n1523 gnd.n1522 19.3944
R7689 gnd.n1522 gnd.n1519 19.3944
R7690 gnd.n1519 gnd.n1518 19.3944
R7691 gnd.n1518 gnd.n1517 19.3944
R7692 gnd.n1517 gnd.n1515 19.3944
R7693 gnd.n1515 gnd.n1213 19.3944
R7694 gnd.n1636 gnd.n1213 19.3944
R7695 gnd.n1636 gnd.n1211 19.3944
R7696 gnd.n1642 gnd.n1211 19.3944
R7697 gnd.n1642 gnd.n1641 19.3944
R7698 gnd.n1641 gnd.n1176 19.3944
R7699 gnd.n1684 gnd.n1176 19.3944
R7700 gnd.n1684 gnd.n1177 19.3944
R7701 gnd.n1193 gnd.n1192 19.3944
R7702 gnd.n1689 gnd.n1688 19.3944
R7703 gnd.n1124 gnd.n1048 19.3944
R7704 gnd.n1119 gnd.n1118 19.3944
R7705 gnd.n1118 gnd.n1116 19.3944
R7706 gnd.n1116 gnd.n1115 19.3944
R7707 gnd.n1115 gnd.n1112 19.3944
R7708 gnd.n1112 gnd.n1111 19.3944
R7709 gnd.n1111 gnd.n1110 19.3944
R7710 gnd.n1110 gnd.n1108 19.3944
R7711 gnd.n1108 gnd.n1107 19.3944
R7712 gnd.n1107 gnd.n1104 19.3944
R7713 gnd.n1104 gnd.n1103 19.3944
R7714 gnd.n1103 gnd.n1102 19.3944
R7715 gnd.n1102 gnd.n1100 19.3944
R7716 gnd.n1100 gnd.n1099 19.3944
R7717 gnd.n1099 gnd.n1094 19.3944
R7718 gnd.n1094 gnd.n1093 19.3944
R7719 gnd.n1093 gnd.n1092 19.3944
R7720 gnd.n1092 gnd.n1090 19.3944
R7721 gnd.n1090 gnd.n1089 19.3944
R7722 gnd.n1089 gnd.n1086 19.3944
R7723 gnd.n1086 gnd.n1085 19.3944
R7724 gnd.n1085 gnd.n1084 19.3944
R7725 gnd.n1084 gnd.n1082 19.3944
R7726 gnd.n1082 gnd.n1081 19.3944
R7727 gnd.n1081 gnd.n1078 19.3944
R7728 gnd.n1078 gnd.n1077 19.3944
R7729 gnd.n1077 gnd.n1076 19.3944
R7730 gnd.n1076 gnd.n883 19.3944
R7731 gnd.n2148 gnd.n883 19.3944
R7732 gnd.n2149 gnd.n2148 19.3944
R7733 gnd.n1475 gnd.n1365 19.3944
R7734 gnd.n1475 gnd.n1363 19.3944
R7735 gnd.n1479 gnd.n1363 19.3944
R7736 gnd.n1479 gnd.n1354 19.3944
R7737 gnd.n1491 gnd.n1354 19.3944
R7738 gnd.n1491 gnd.n1352 19.3944
R7739 gnd.n1495 gnd.n1352 19.3944
R7740 gnd.n1495 gnd.n1341 19.3944
R7741 gnd.n1537 gnd.n1341 19.3944
R7742 gnd.n1537 gnd.n1295 19.3944
R7743 gnd.n1543 gnd.n1295 19.3944
R7744 gnd.n1543 gnd.n1542 19.3944
R7745 gnd.n1542 gnd.n1273 19.3944
R7746 gnd.n1564 gnd.n1273 19.3944
R7747 gnd.n1564 gnd.n1266 19.3944
R7748 gnd.n1575 gnd.n1266 19.3944
R7749 gnd.n1575 gnd.n1574 19.3944
R7750 gnd.n1574 gnd.n1247 19.3944
R7751 gnd.n1595 gnd.n1247 19.3944
R7752 gnd.n1595 gnd.n1237 19.3944
R7753 gnd.n1605 gnd.n1237 19.3944
R7754 gnd.n1605 gnd.n1218 19.3944
R7755 gnd.n1632 gnd.n1218 19.3944
R7756 gnd.n1632 gnd.n1631 19.3944
R7757 gnd.n1631 gnd.n1206 19.3944
R7758 gnd.n1648 gnd.n1206 19.3944
R7759 gnd.n1648 gnd.n1184 19.3944
R7760 gnd.n1680 gnd.n1184 19.3944
R7761 gnd.n1680 gnd.n1679 19.3944
R7762 gnd.n1679 gnd.n1678 19.3944
R7763 gnd.n1678 gnd.n1190 19.3944
R7764 gnd.n1190 gnd.n1040 19.3944
R7765 gnd.n1700 gnd.n1040 19.3944
R7766 gnd.n1700 gnd.n1699 19.3944
R7767 gnd.n1699 gnd.n1024 19.3944
R7768 gnd.n1720 gnd.n1024 19.3944
R7769 gnd.n1720 gnd.n1017 19.3944
R7770 gnd.n1731 gnd.n1017 19.3944
R7771 gnd.n1731 gnd.n1730 19.3944
R7772 gnd.n1730 gnd.n999 19.3944
R7773 gnd.n1751 gnd.n999 19.3944
R7774 gnd.n1751 gnd.n991 19.3944
R7775 gnd.n1762 gnd.n991 19.3944
R7776 gnd.n1762 gnd.n1761 19.3944
R7777 gnd.n1761 gnd.n972 19.3944
R7778 gnd.n1782 gnd.n972 19.3944
R7779 gnd.n1782 gnd.n965 19.3944
R7780 gnd.n1793 gnd.n965 19.3944
R7781 gnd.n1793 gnd.n1792 19.3944
R7782 gnd.n1792 gnd.n948 19.3944
R7783 gnd.n1813 gnd.n948 19.3944
R7784 gnd.n1813 gnd.n941 19.3944
R7785 gnd.n1824 gnd.n941 19.3944
R7786 gnd.n1824 gnd.n1823 19.3944
R7787 gnd.n1823 gnd.n922 19.3944
R7788 gnd.n1844 gnd.n922 19.3944
R7789 gnd.n1844 gnd.n915 19.3944
R7790 gnd.n1855 gnd.n915 19.3944
R7791 gnd.n1855 gnd.n1854 19.3944
R7792 gnd.n1854 gnd.n897 19.3944
R7793 gnd.n2132 gnd.n897 19.3944
R7794 gnd.n2132 gnd.n887 19.3944
R7795 gnd.n2143 gnd.n887 19.3944
R7796 gnd.n2143 gnd.n779 19.3944
R7797 gnd.n5989 gnd.n779 19.3944
R7798 gnd.n3969 gnd.n3455 19.3944
R7799 gnd.n3969 gnd.n3968 19.3944
R7800 gnd.n3968 gnd.n3459 19.3944
R7801 gnd.n3961 gnd.n3459 19.3944
R7802 gnd.n3961 gnd.n3960 19.3944
R7803 gnd.n3960 gnd.n3469 19.3944
R7804 gnd.n3953 gnd.n3469 19.3944
R7805 gnd.n3953 gnd.n3952 19.3944
R7806 gnd.n3952 gnd.n3479 19.3944
R7807 gnd.n3945 gnd.n3479 19.3944
R7808 gnd.n3945 gnd.n3944 19.3944
R7809 gnd.n3944 gnd.n3489 19.3944
R7810 gnd.n3937 gnd.n3489 19.3944
R7811 gnd.n3937 gnd.n3936 19.3944
R7812 gnd.n3936 gnd.n3499 19.3944
R7813 gnd.n3929 gnd.n3499 19.3944
R7814 gnd.n3781 gnd.n2262 19.3944
R7815 gnd.n3784 gnd.n3781 19.3944
R7816 gnd.n3785 gnd.n3784 19.3944
R7817 gnd.n3787 gnd.n3785 19.3944
R7818 gnd.n3788 gnd.n3787 19.3944
R7819 gnd.n3791 gnd.n3788 19.3944
R7820 gnd.n3792 gnd.n3791 19.3944
R7821 gnd.n3794 gnd.n3792 19.3944
R7822 gnd.n3795 gnd.n3794 19.3944
R7823 gnd.n3798 gnd.n3795 19.3944
R7824 gnd.n3799 gnd.n3798 19.3944
R7825 gnd.n3801 gnd.n3799 19.3944
R7826 gnd.n3802 gnd.n3801 19.3944
R7827 gnd.n3805 gnd.n3802 19.3944
R7828 gnd.n3806 gnd.n3805 19.3944
R7829 gnd.n3808 gnd.n3806 19.3944
R7830 gnd.n3809 gnd.n3808 19.3944
R7831 gnd.n3812 gnd.n3809 19.3944
R7832 gnd.n3813 gnd.n3812 19.3944
R7833 gnd.n3815 gnd.n3813 19.3944
R7834 gnd.n3816 gnd.n3815 19.3944
R7835 gnd.n3819 gnd.n3816 19.3944
R7836 gnd.n3820 gnd.n3819 19.3944
R7837 gnd.n3822 gnd.n3820 19.3944
R7838 gnd.n3823 gnd.n3822 19.3944
R7839 gnd.n3826 gnd.n3823 19.3944
R7840 gnd.n3827 gnd.n3826 19.3944
R7841 gnd.n3828 gnd.n3827 19.3944
R7842 gnd.n3828 gnd.n3652 19.3944
R7843 gnd.n3840 gnd.n3652 19.3944
R7844 gnd.n3841 gnd.n3840 19.3944
R7845 gnd.n3842 gnd.n3841 19.3944
R7846 gnd.n3843 gnd.n3842 19.3944
R7847 gnd.n3847 gnd.n3843 19.3944
R7848 gnd.n3848 gnd.n3847 19.3944
R7849 gnd.n3851 gnd.n3848 19.3944
R7850 gnd.n3852 gnd.n3851 19.3944
R7851 gnd.n3856 gnd.n3852 19.3944
R7852 gnd.n3857 gnd.n3856 19.3944
R7853 gnd.n3861 gnd.n3857 19.3944
R7854 gnd.n3861 gnd.n3860 19.3944
R7855 gnd.n3860 gnd.n3859 19.3944
R7856 gnd.n3686 gnd.n3685 19.3944
R7857 gnd.n3689 gnd.n3686 19.3944
R7858 gnd.n3689 gnd.n3683 19.3944
R7859 gnd.n3695 gnd.n3683 19.3944
R7860 gnd.n3696 gnd.n3695 19.3944
R7861 gnd.n3699 gnd.n3696 19.3944
R7862 gnd.n3699 gnd.n3681 19.3944
R7863 gnd.n3705 gnd.n3681 19.3944
R7864 gnd.n3706 gnd.n3705 19.3944
R7865 gnd.n3709 gnd.n3706 19.3944
R7866 gnd.n3709 gnd.n3679 19.3944
R7867 gnd.n3715 gnd.n3679 19.3944
R7868 gnd.n3716 gnd.n3715 19.3944
R7869 gnd.n3719 gnd.n3716 19.3944
R7870 gnd.n3719 gnd.n3675 19.3944
R7871 gnd.n3723 gnd.n3675 19.3944
R7872 gnd.n3728 gnd.n3670 19.3944
R7873 gnd.n3733 gnd.n3670 19.3944
R7874 gnd.n3734 gnd.n3733 19.3944
R7875 gnd.n3736 gnd.n3734 19.3944
R7876 gnd.n3736 gnd.n3668 19.3944
R7877 gnd.n3741 gnd.n3668 19.3944
R7878 gnd.n3742 gnd.n3741 19.3944
R7879 gnd.n3744 gnd.n3742 19.3944
R7880 gnd.n3744 gnd.n3666 19.3944
R7881 gnd.n3749 gnd.n3666 19.3944
R7882 gnd.n3750 gnd.n3749 19.3944
R7883 gnd.n3752 gnd.n3750 19.3944
R7884 gnd.n3752 gnd.n3664 19.3944
R7885 gnd.n3757 gnd.n3664 19.3944
R7886 gnd.n3758 gnd.n3757 19.3944
R7887 gnd.n3760 gnd.n3758 19.3944
R7888 gnd.n3760 gnd.n3662 19.3944
R7889 gnd.n3765 gnd.n3662 19.3944
R7890 gnd.n3766 gnd.n3765 19.3944
R7891 gnd.n3768 gnd.n3766 19.3944
R7892 gnd.n3768 gnd.n3659 19.3944
R7893 gnd.n3772 gnd.n3659 19.3944
R7894 gnd.n3773 gnd.n3772 19.3944
R7895 gnd.n3775 gnd.n3773 19.3944
R7896 gnd.n3775 gnd.n3656 19.3944
R7897 gnd.n3779 gnd.n3656 19.3944
R7898 gnd.n3780 gnd.n3779 19.3944
R7899 gnd.n3832 gnd.n3780 19.3944
R7900 gnd.n3832 gnd.n3654 19.3944
R7901 gnd.n3836 gnd.n3654 19.3944
R7902 gnd.n3836 gnd.n3643 19.3944
R7903 gnd.n3881 gnd.n3643 19.3944
R7904 gnd.n3881 gnd.n3644 19.3944
R7905 gnd.n3877 gnd.n3644 19.3944
R7906 gnd.n3877 gnd.n3876 19.3944
R7907 gnd.n3876 gnd.n3875 19.3944
R7908 gnd.n3875 gnd.n3649 19.3944
R7909 gnd.n3871 gnd.n3649 19.3944
R7910 gnd.n3871 gnd.n3870 19.3944
R7911 gnd.n3870 gnd.n3869 19.3944
R7912 gnd.n3869 gnd.n3865 19.3944
R7913 gnd.n3865 gnd.n3520 19.3944
R7914 gnd.n5925 gnd.n5924 19.3944
R7915 gnd.n5924 gnd.n5923 19.3944
R7916 gnd.n5923 gnd.n5922 19.3944
R7917 gnd.n5922 gnd.n5920 19.3944
R7918 gnd.n5920 gnd.n5917 19.3944
R7919 gnd.n5917 gnd.n5916 19.3944
R7920 gnd.n5916 gnd.n5913 19.3944
R7921 gnd.n5913 gnd.n5912 19.3944
R7922 gnd.n5912 gnd.n5909 19.3944
R7923 gnd.n5909 gnd.n5908 19.3944
R7924 gnd.n5908 gnd.n5905 19.3944
R7925 gnd.n5905 gnd.n5904 19.3944
R7926 gnd.n5904 gnd.n5901 19.3944
R7927 gnd.n5901 gnd.n5900 19.3944
R7928 gnd.n5900 gnd.n5897 19.3944
R7929 gnd.n5897 gnd.n5896 19.3944
R7930 gnd.n5896 gnd.n5893 19.3944
R7931 gnd.n5891 gnd.n5888 19.3944
R7932 gnd.n5888 gnd.n5887 19.3944
R7933 gnd.n5887 gnd.n5884 19.3944
R7934 gnd.n5884 gnd.n5883 19.3944
R7935 gnd.n5883 gnd.n5880 19.3944
R7936 gnd.n5880 gnd.n5879 19.3944
R7937 gnd.n5879 gnd.n5876 19.3944
R7938 gnd.n5876 gnd.n5875 19.3944
R7939 gnd.n5875 gnd.n5872 19.3944
R7940 gnd.n5872 gnd.n5871 19.3944
R7941 gnd.n5871 gnd.n5868 19.3944
R7942 gnd.n5868 gnd.n5867 19.3944
R7943 gnd.n5867 gnd.n5864 19.3944
R7944 gnd.n5864 gnd.n5863 19.3944
R7945 gnd.n5863 gnd.n5860 19.3944
R7946 gnd.n5860 gnd.n5859 19.3944
R7947 gnd.n5859 gnd.n5856 19.3944
R7948 gnd.n5856 gnd.n5855 19.3944
R7949 gnd.n5851 gnd.n5848 19.3944
R7950 gnd.n5848 gnd.n5847 19.3944
R7951 gnd.n5847 gnd.n5844 19.3944
R7952 gnd.n5844 gnd.n5843 19.3944
R7953 gnd.n5843 gnd.n5840 19.3944
R7954 gnd.n5840 gnd.n5839 19.3944
R7955 gnd.n5839 gnd.n5836 19.3944
R7956 gnd.n5836 gnd.n5835 19.3944
R7957 gnd.n5835 gnd.n5832 19.3944
R7958 gnd.n5832 gnd.n5831 19.3944
R7959 gnd.n5831 gnd.n5828 19.3944
R7960 gnd.n5828 gnd.n5827 19.3944
R7961 gnd.n5827 gnd.n5824 19.3944
R7962 gnd.n5824 gnd.n5823 19.3944
R7963 gnd.n5823 gnd.n5820 19.3944
R7964 gnd.n5820 gnd.n5819 19.3944
R7965 gnd.n5819 gnd.n5816 19.3944
R7966 gnd.n5816 gnd.n5815 19.3944
R7967 gnd.n5676 gnd.n2472 19.3944
R7968 gnd.n5671 gnd.n2472 19.3944
R7969 gnd.n5671 gnd.n5670 19.3944
R7970 gnd.n5670 gnd.n5669 19.3944
R7971 gnd.n5669 gnd.n5666 19.3944
R7972 gnd.n5666 gnd.n5665 19.3944
R7973 gnd.n5665 gnd.n5662 19.3944
R7974 gnd.n5662 gnd.n5661 19.3944
R7975 gnd.n5661 gnd.n5658 19.3944
R7976 gnd.n5658 gnd.n5657 19.3944
R7977 gnd.n5657 gnd.n5654 19.3944
R7978 gnd.n5654 gnd.n5653 19.3944
R7979 gnd.n5653 gnd.n5650 19.3944
R7980 gnd.n5650 gnd.n5649 19.3944
R7981 gnd.n5649 gnd.n5646 19.3944
R7982 gnd.n5646 gnd.n5645 19.3944
R7983 gnd.n5645 gnd.n5642 19.3944
R7984 gnd.n3568 gnd.n3565 19.3944
R7985 gnd.n3571 gnd.n3568 19.3944
R7986 gnd.n3571 gnd.n3531 19.3944
R7987 gnd.n3575 gnd.n3531 19.3944
R7988 gnd.n3578 gnd.n3575 19.3944
R7989 gnd.n3581 gnd.n3578 19.3944
R7990 gnd.n3581 gnd.n3529 19.3944
R7991 gnd.n3585 gnd.n3529 19.3944
R7992 gnd.n3588 gnd.n3585 19.3944
R7993 gnd.n3591 gnd.n3588 19.3944
R7994 gnd.n3591 gnd.n3527 19.3944
R7995 gnd.n3595 gnd.n3527 19.3944
R7996 gnd.n3598 gnd.n3595 19.3944
R7997 gnd.n3601 gnd.n3598 19.3944
R7998 gnd.n3601 gnd.n3525 19.3944
R7999 gnd.n3605 gnd.n3525 19.3944
R8000 gnd.n3608 gnd.n3605 19.3944
R8001 gnd.n3611 gnd.n3608 19.3944
R8002 gnd.n3541 gnd.n2541 19.3944
R8003 gnd.n3545 gnd.n3541 19.3944
R8004 gnd.n3548 gnd.n3545 19.3944
R8005 gnd.n3551 gnd.n3548 19.3944
R8006 gnd.n3551 gnd.n3537 19.3944
R8007 gnd.n3555 gnd.n3537 19.3944
R8008 gnd.n3558 gnd.n3555 19.3944
R8009 gnd.n3561 gnd.n3558 19.3944
R8010 gnd.n5640 gnd.n5637 19.3944
R8011 gnd.n5637 gnd.n5636 19.3944
R8012 gnd.n5636 gnd.n5633 19.3944
R8013 gnd.n5633 gnd.n5632 19.3944
R8014 gnd.n5632 gnd.n5629 19.3944
R8015 gnd.n5629 gnd.n5628 19.3944
R8016 gnd.n5628 gnd.n5625 19.3944
R8017 gnd.n5802 gnd.n2272 19.3944
R8018 gnd.n5802 gnd.n2273 19.3944
R8019 gnd.n5798 gnd.n2273 19.3944
R8020 gnd.n5798 gnd.n2276 19.3944
R8021 gnd.n5788 gnd.n2276 19.3944
R8022 gnd.n5788 gnd.n5787 19.3944
R8023 gnd.n5787 gnd.n5786 19.3944
R8024 gnd.n5786 gnd.n2296 19.3944
R8025 gnd.n5776 gnd.n2296 19.3944
R8026 gnd.n5776 gnd.n5775 19.3944
R8027 gnd.n5775 gnd.n5774 19.3944
R8028 gnd.n5774 gnd.n2314 19.3944
R8029 gnd.n5764 gnd.n2314 19.3944
R8030 gnd.n5764 gnd.n5763 19.3944
R8031 gnd.n5763 gnd.n5762 19.3944
R8032 gnd.n5762 gnd.n2334 19.3944
R8033 gnd.n5752 gnd.n2334 19.3944
R8034 gnd.n5752 gnd.n5751 19.3944
R8035 gnd.n5751 gnd.n5750 19.3944
R8036 gnd.n5750 gnd.n2352 19.3944
R8037 gnd.n5740 gnd.n2352 19.3944
R8038 gnd.n5740 gnd.n5739 19.3944
R8039 gnd.n5739 gnd.n5738 19.3944
R8040 gnd.n5738 gnd.n2372 19.3944
R8041 gnd.n5728 gnd.n2372 19.3944
R8042 gnd.n5728 gnd.n5727 19.3944
R8043 gnd.n5727 gnd.n5726 19.3944
R8044 gnd.n5726 gnd.n2391 19.3944
R8045 gnd.n5716 gnd.n2391 19.3944
R8046 gnd.n5716 gnd.n5715 19.3944
R8047 gnd.n5715 gnd.n5714 19.3944
R8048 gnd.n5714 gnd.n2411 19.3944
R8049 gnd.n5704 gnd.n2411 19.3944
R8050 gnd.n5704 gnd.n5703 19.3944
R8051 gnd.n5703 gnd.n5702 19.3944
R8052 gnd.n5702 gnd.n2431 19.3944
R8053 gnd.n5692 gnd.n2431 19.3944
R8054 gnd.n5692 gnd.n5691 19.3944
R8055 gnd.n5691 gnd.n5690 19.3944
R8056 gnd.n5690 gnd.n2452 19.3944
R8057 gnd.n5680 gnd.n2452 19.3944
R8058 gnd.n5680 gnd.n5679 19.3944
R8059 gnd.n5807 gnd.n2264 19.3944
R8060 gnd.n2283 gnd.n2264 19.3944
R8061 gnd.n5794 gnd.n2283 19.3944
R8062 gnd.n5794 gnd.n5793 19.3944
R8063 gnd.n5793 gnd.n5792 19.3944
R8064 gnd.n5792 gnd.n2287 19.3944
R8065 gnd.n5782 gnd.n2287 19.3944
R8066 gnd.n5782 gnd.n5781 19.3944
R8067 gnd.n5781 gnd.n5780 19.3944
R8068 gnd.n5780 gnd.n2305 19.3944
R8069 gnd.n5770 gnd.n2305 19.3944
R8070 gnd.n5770 gnd.n5769 19.3944
R8071 gnd.n5769 gnd.n5768 19.3944
R8072 gnd.n5768 gnd.n2323 19.3944
R8073 gnd.n5758 gnd.n2323 19.3944
R8074 gnd.n5758 gnd.n5757 19.3944
R8075 gnd.n5757 gnd.n5756 19.3944
R8076 gnd.n5756 gnd.n2343 19.3944
R8077 gnd.n5746 gnd.n2343 19.3944
R8078 gnd.n5746 gnd.n5745 19.3944
R8079 gnd.n5745 gnd.n5744 19.3944
R8080 gnd.n5744 gnd.n2361 19.3944
R8081 gnd.n5734 gnd.n2361 19.3944
R8082 gnd.n5734 gnd.n5733 19.3944
R8083 gnd.n5733 gnd.n5732 19.3944
R8084 gnd.n5732 gnd.n2381 19.3944
R8085 gnd.n5722 gnd.n2381 19.3944
R8086 gnd.n5722 gnd.n5721 19.3944
R8087 gnd.n5721 gnd.n5720 19.3944
R8088 gnd.n5720 gnd.n2400 19.3944
R8089 gnd.n5710 gnd.n2400 19.3944
R8090 gnd.n5710 gnd.n5709 19.3944
R8091 gnd.n5709 gnd.n5708 19.3944
R8092 gnd.n5708 gnd.n2421 19.3944
R8093 gnd.n5698 gnd.n2421 19.3944
R8094 gnd.n5698 gnd.n5697 19.3944
R8095 gnd.n5697 gnd.n5696 19.3944
R8096 gnd.n5696 gnd.n2441 19.3944
R8097 gnd.n5686 gnd.n2441 19.3944
R8098 gnd.n5686 gnd.n5685 19.3944
R8099 gnd.n5685 gnd.n5684 19.3944
R8100 gnd.n5684 gnd.n2462 19.3944
R8101 gnd.n3635 gnd.n3632 19.3944
R8102 gnd.n3639 gnd.n3632 19.3944
R8103 gnd.n3639 gnd.n3630 19.3944
R8104 gnd.n3886 gnd.n3630 19.3944
R8105 gnd.n3886 gnd.n3628 19.3944
R8106 gnd.n3890 gnd.n3628 19.3944
R8107 gnd.n3890 gnd.n3626 19.3944
R8108 gnd.n3894 gnd.n3626 19.3944
R8109 gnd.n3894 gnd.n3624 19.3944
R8110 gnd.n3898 gnd.n3624 19.3944
R8111 gnd.n3898 gnd.n3622 19.3944
R8112 gnd.n3902 gnd.n3622 19.3944
R8113 gnd.n3902 gnd.n3620 19.3944
R8114 gnd.n3921 gnd.n3620 19.3944
R8115 gnd.n3921 gnd.n3920 19.3944
R8116 gnd.n3920 gnd.n3919 19.3944
R8117 gnd.n3919 gnd.n3908 19.3944
R8118 gnd.n3914 gnd.n3908 19.3944
R8119 gnd.n3914 gnd.n3913 19.3944
R8120 gnd.n3913 gnd.n3389 19.3944
R8121 gnd.n4000 gnd.n3389 19.3944
R8122 gnd.n4000 gnd.n3387 19.3944
R8123 gnd.n4004 gnd.n3387 19.3944
R8124 gnd.n4004 gnd.n3374 19.3944
R8125 gnd.n4016 gnd.n3374 19.3944
R8126 gnd.n4016 gnd.n3372 19.3944
R8127 gnd.n4020 gnd.n3372 19.3944
R8128 gnd.n4020 gnd.n3359 19.3944
R8129 gnd.n4044 gnd.n3359 19.3944
R8130 gnd.n4044 gnd.n3357 19.3944
R8131 gnd.n4051 gnd.n3357 19.3944
R8132 gnd.n4051 gnd.n4050 19.3944
R8133 gnd.n4050 gnd.n2611 19.3944
R8134 gnd.n5547 gnd.n2611 19.3944
R8135 gnd.n5547 gnd.n5546 19.3944
R8136 gnd.n5546 gnd.n5545 19.3944
R8137 gnd.n5545 gnd.n2615 19.3944
R8138 gnd.n3336 gnd.n2615 19.3944
R8139 gnd.n3336 gnd.n3318 19.3944
R8140 gnd.n4193 gnd.n3318 19.3944
R8141 gnd.n4193 gnd.n3316 19.3944
R8142 gnd.n4202 gnd.n3316 19.3944
R8143 gnd.n4202 gnd.n4201 19.3944
R8144 gnd.n4201 gnd.n4200 19.3944
R8145 gnd.n4200 gnd.n3288 19.3944
R8146 gnd.n4262 gnd.n3288 19.3944
R8147 gnd.n4262 gnd.n3286 19.3944
R8148 gnd.n4266 gnd.n3286 19.3944
R8149 gnd.n4266 gnd.n3271 19.3944
R8150 gnd.n4291 gnd.n3271 19.3944
R8151 gnd.n4291 gnd.n3269 19.3944
R8152 gnd.n4297 gnd.n3269 19.3944
R8153 gnd.n4297 gnd.n4296 19.3944
R8154 gnd.n4296 gnd.n3243 19.3944
R8155 gnd.n4365 gnd.n3243 19.3944
R8156 gnd.n4365 gnd.n3241 19.3944
R8157 gnd.n4371 gnd.n3241 19.3944
R8158 gnd.n4371 gnd.n4370 19.3944
R8159 gnd.n4370 gnd.n3220 19.3944
R8160 gnd.n4397 gnd.n3220 19.3944
R8161 gnd.n4397 gnd.n3218 19.3944
R8162 gnd.n4403 gnd.n3218 19.3944
R8163 gnd.n4403 gnd.n4402 19.3944
R8164 gnd.n4402 gnd.n3199 19.3944
R8165 gnd.n4438 gnd.n3199 19.3944
R8166 gnd.n4438 gnd.n3197 19.3944
R8167 gnd.n4444 gnd.n3197 19.3944
R8168 gnd.n4444 gnd.n4443 19.3944
R8169 gnd.n4443 gnd.n3170 19.3944
R8170 gnd.n4507 gnd.n3170 19.3944
R8171 gnd.n4507 gnd.n3168 19.3944
R8172 gnd.n4513 gnd.n3168 19.3944
R8173 gnd.n4513 gnd.n4512 19.3944
R8174 gnd.n4512 gnd.n3145 19.3944
R8175 gnd.n4539 gnd.n3145 19.3944
R8176 gnd.n4539 gnd.n3143 19.3944
R8177 gnd.n4545 gnd.n3143 19.3944
R8178 gnd.n4545 gnd.n4544 19.3944
R8179 gnd.n4544 gnd.n3122 19.3944
R8180 gnd.n4579 gnd.n3122 19.3944
R8181 gnd.n4579 gnd.n3120 19.3944
R8182 gnd.n4585 gnd.n3120 19.3944
R8183 gnd.n4585 gnd.n4584 19.3944
R8184 gnd.n4584 gnd.n3093 19.3944
R8185 gnd.n4633 gnd.n3093 19.3944
R8186 gnd.n4633 gnd.n3091 19.3944
R8187 gnd.n4639 gnd.n3091 19.3944
R8188 gnd.n4639 gnd.n4638 19.3944
R8189 gnd.n4638 gnd.n3069 19.3944
R8190 gnd.n4675 gnd.n3069 19.3944
R8191 gnd.n4675 gnd.n3067 19.3944
R8192 gnd.n4681 gnd.n3067 19.3944
R8193 gnd.n4681 gnd.n4680 19.3944
R8194 gnd.n4680 gnd.n3041 19.3944
R8195 gnd.n4718 gnd.n3041 19.3944
R8196 gnd.n4718 gnd.n3039 19.3944
R8197 gnd.n4723 gnd.n3039 19.3944
R8198 gnd.n4723 gnd.n3018 19.3944
R8199 gnd.n4763 gnd.n3018 19.3944
R8200 gnd.n4763 gnd.n4762 19.3944
R8201 gnd.n4762 gnd.n4761 19.3944
R8202 gnd.n4761 gnd.n3022 19.3944
R8203 gnd.n3025 gnd.n3022 19.3944
R8204 gnd.n3025 gnd.n2987 19.3944
R8205 gnd.n4810 gnd.n2987 19.3944
R8206 gnd.n4810 gnd.n2985 19.3944
R8207 gnd.n4814 gnd.n2985 19.3944
R8208 gnd.n4814 gnd.n2935 19.3944
R8209 gnd.n4982 gnd.n2935 19.3944
R8210 gnd.n4982 gnd.n2933 19.3944
R8211 gnd.n4986 gnd.n2933 19.3944
R8212 gnd.n4986 gnd.n2923 19.3944
R8213 gnd.n5000 gnd.n2923 19.3944
R8214 gnd.n5000 gnd.n2921 19.3944
R8215 gnd.n5004 gnd.n2921 19.3944
R8216 gnd.n5004 gnd.n2912 19.3944
R8217 gnd.n5017 gnd.n2912 19.3944
R8218 gnd.n5017 gnd.n2910 19.3944
R8219 gnd.n5023 gnd.n2910 19.3944
R8220 gnd.n5023 gnd.n5022 19.3944
R8221 gnd.n5022 gnd.n2899 19.3944
R8222 gnd.n5054 gnd.n2899 19.3944
R8223 gnd.n5054 gnd.n2897 19.3944
R8224 gnd.n5058 gnd.n2897 19.3944
R8225 gnd.n5058 gnd.n2895 19.3944
R8226 gnd.n5063 gnd.n2895 19.3944
R8227 gnd.n5063 gnd.n2893 19.3944
R8228 gnd.n5189 gnd.n2893 19.3944
R8229 gnd.n5189 gnd.n5188 19.3944
R8230 gnd.n5188 gnd.n5187 19.3944
R8231 gnd.n5187 gnd.n5069 19.3944
R8232 gnd.n5112 gnd.n5069 19.3944
R8233 gnd.n5112 gnd.n5109 19.3944
R8234 gnd.n5125 gnd.n5109 19.3944
R8235 gnd.n5125 gnd.n5124 19.3944
R8236 gnd.n5124 gnd.n5123 19.3944
R8237 gnd.n5123 gnd.n5120 19.3944
R8238 gnd.n5120 gnd.n252 19.3944
R8239 gnd.n6741 gnd.n252 19.3944
R8240 gnd.n6741 gnd.n6740 19.3944
R8241 gnd.n6740 gnd.n6739 19.3944
R8242 gnd.n6525 gnd.n379 19.3944
R8243 gnd.n6531 gnd.n379 19.3944
R8244 gnd.n6531 gnd.n377 19.3944
R8245 gnd.n6535 gnd.n377 19.3944
R8246 gnd.n6535 gnd.n373 19.3944
R8247 gnd.n6541 gnd.n373 19.3944
R8248 gnd.n6541 gnd.n371 19.3944
R8249 gnd.n6545 gnd.n371 19.3944
R8250 gnd.n6545 gnd.n367 19.3944
R8251 gnd.n6551 gnd.n367 19.3944
R8252 gnd.n6551 gnd.n365 19.3944
R8253 gnd.n6555 gnd.n365 19.3944
R8254 gnd.n6555 gnd.n361 19.3944
R8255 gnd.n6561 gnd.n361 19.3944
R8256 gnd.n6561 gnd.n359 19.3944
R8257 gnd.n6565 gnd.n359 19.3944
R8258 gnd.n6565 gnd.n355 19.3944
R8259 gnd.n6571 gnd.n355 19.3944
R8260 gnd.n6571 gnd.n353 19.3944
R8261 gnd.n6575 gnd.n353 19.3944
R8262 gnd.n6575 gnd.n349 19.3944
R8263 gnd.n6581 gnd.n349 19.3944
R8264 gnd.n6581 gnd.n347 19.3944
R8265 gnd.n6585 gnd.n347 19.3944
R8266 gnd.n6585 gnd.n343 19.3944
R8267 gnd.n6591 gnd.n343 19.3944
R8268 gnd.n6591 gnd.n341 19.3944
R8269 gnd.n6595 gnd.n341 19.3944
R8270 gnd.n6595 gnd.n337 19.3944
R8271 gnd.n6601 gnd.n337 19.3944
R8272 gnd.n6601 gnd.n335 19.3944
R8273 gnd.n6605 gnd.n335 19.3944
R8274 gnd.n6605 gnd.n331 19.3944
R8275 gnd.n6611 gnd.n331 19.3944
R8276 gnd.n6611 gnd.n329 19.3944
R8277 gnd.n6615 gnd.n329 19.3944
R8278 gnd.n6615 gnd.n325 19.3944
R8279 gnd.n6621 gnd.n325 19.3944
R8280 gnd.n6621 gnd.n323 19.3944
R8281 gnd.n6625 gnd.n323 19.3944
R8282 gnd.n6625 gnd.n319 19.3944
R8283 gnd.n6631 gnd.n319 19.3944
R8284 gnd.n6631 gnd.n317 19.3944
R8285 gnd.n6635 gnd.n317 19.3944
R8286 gnd.n6635 gnd.n313 19.3944
R8287 gnd.n6641 gnd.n313 19.3944
R8288 gnd.n6641 gnd.n311 19.3944
R8289 gnd.n6645 gnd.n311 19.3944
R8290 gnd.n6645 gnd.n307 19.3944
R8291 gnd.n6651 gnd.n307 19.3944
R8292 gnd.n6651 gnd.n305 19.3944
R8293 gnd.n6655 gnd.n305 19.3944
R8294 gnd.n6655 gnd.n301 19.3944
R8295 gnd.n6661 gnd.n301 19.3944
R8296 gnd.n6661 gnd.n299 19.3944
R8297 gnd.n6665 gnd.n299 19.3944
R8298 gnd.n6665 gnd.n295 19.3944
R8299 gnd.n6671 gnd.n295 19.3944
R8300 gnd.n6671 gnd.n293 19.3944
R8301 gnd.n6675 gnd.n293 19.3944
R8302 gnd.n6675 gnd.n289 19.3944
R8303 gnd.n6681 gnd.n289 19.3944
R8304 gnd.n6681 gnd.n287 19.3944
R8305 gnd.n6685 gnd.n287 19.3944
R8306 gnd.n6685 gnd.n283 19.3944
R8307 gnd.n6691 gnd.n283 19.3944
R8308 gnd.n6691 gnd.n281 19.3944
R8309 gnd.n6695 gnd.n281 19.3944
R8310 gnd.n6695 gnd.n277 19.3944
R8311 gnd.n6701 gnd.n277 19.3944
R8312 gnd.n6701 gnd.n275 19.3944
R8313 gnd.n6705 gnd.n275 19.3944
R8314 gnd.n6705 gnd.n271 19.3944
R8315 gnd.n6711 gnd.n271 19.3944
R8316 gnd.n6711 gnd.n269 19.3944
R8317 gnd.n6715 gnd.n269 19.3944
R8318 gnd.n6715 gnd.n265 19.3944
R8319 gnd.n6721 gnd.n265 19.3944
R8320 gnd.n6721 gnd.n263 19.3944
R8321 gnd.n6725 gnd.n263 19.3944
R8322 gnd.n6725 gnd.n259 19.3944
R8323 gnd.n6732 gnd.n259 19.3944
R8324 gnd.n6732 gnd.n257 19.3944
R8325 gnd.n6736 gnd.n257 19.3944
R8326 gnd.n6170 gnd.n592 19.3944
R8327 gnd.n6174 gnd.n592 19.3944
R8328 gnd.n6174 gnd.n588 19.3944
R8329 gnd.n6180 gnd.n588 19.3944
R8330 gnd.n6180 gnd.n586 19.3944
R8331 gnd.n6184 gnd.n586 19.3944
R8332 gnd.n6184 gnd.n582 19.3944
R8333 gnd.n6190 gnd.n582 19.3944
R8334 gnd.n6190 gnd.n580 19.3944
R8335 gnd.n6194 gnd.n580 19.3944
R8336 gnd.n6194 gnd.n576 19.3944
R8337 gnd.n6200 gnd.n576 19.3944
R8338 gnd.n6200 gnd.n574 19.3944
R8339 gnd.n6204 gnd.n574 19.3944
R8340 gnd.n6204 gnd.n570 19.3944
R8341 gnd.n6210 gnd.n570 19.3944
R8342 gnd.n6210 gnd.n568 19.3944
R8343 gnd.n6214 gnd.n568 19.3944
R8344 gnd.n6214 gnd.n564 19.3944
R8345 gnd.n6220 gnd.n564 19.3944
R8346 gnd.n6220 gnd.n562 19.3944
R8347 gnd.n6224 gnd.n562 19.3944
R8348 gnd.n6224 gnd.n558 19.3944
R8349 gnd.n6230 gnd.n558 19.3944
R8350 gnd.n6230 gnd.n556 19.3944
R8351 gnd.n6234 gnd.n556 19.3944
R8352 gnd.n6234 gnd.n552 19.3944
R8353 gnd.n6240 gnd.n552 19.3944
R8354 gnd.n6240 gnd.n550 19.3944
R8355 gnd.n6244 gnd.n550 19.3944
R8356 gnd.n6244 gnd.n546 19.3944
R8357 gnd.n6250 gnd.n546 19.3944
R8358 gnd.n6250 gnd.n544 19.3944
R8359 gnd.n6254 gnd.n544 19.3944
R8360 gnd.n6254 gnd.n540 19.3944
R8361 gnd.n6260 gnd.n540 19.3944
R8362 gnd.n6260 gnd.n538 19.3944
R8363 gnd.n6264 gnd.n538 19.3944
R8364 gnd.n6264 gnd.n534 19.3944
R8365 gnd.n6270 gnd.n534 19.3944
R8366 gnd.n6270 gnd.n532 19.3944
R8367 gnd.n6274 gnd.n532 19.3944
R8368 gnd.n6274 gnd.n528 19.3944
R8369 gnd.n6280 gnd.n528 19.3944
R8370 gnd.n6280 gnd.n526 19.3944
R8371 gnd.n6284 gnd.n526 19.3944
R8372 gnd.n6284 gnd.n522 19.3944
R8373 gnd.n6290 gnd.n522 19.3944
R8374 gnd.n6290 gnd.n520 19.3944
R8375 gnd.n6294 gnd.n520 19.3944
R8376 gnd.n6294 gnd.n516 19.3944
R8377 gnd.n6300 gnd.n516 19.3944
R8378 gnd.n6300 gnd.n514 19.3944
R8379 gnd.n6304 gnd.n514 19.3944
R8380 gnd.n6304 gnd.n510 19.3944
R8381 gnd.n6310 gnd.n510 19.3944
R8382 gnd.n6310 gnd.n508 19.3944
R8383 gnd.n6314 gnd.n508 19.3944
R8384 gnd.n6314 gnd.n504 19.3944
R8385 gnd.n6320 gnd.n504 19.3944
R8386 gnd.n6320 gnd.n502 19.3944
R8387 gnd.n6324 gnd.n502 19.3944
R8388 gnd.n6324 gnd.n498 19.3944
R8389 gnd.n6330 gnd.n498 19.3944
R8390 gnd.n6330 gnd.n496 19.3944
R8391 gnd.n6334 gnd.n496 19.3944
R8392 gnd.n6334 gnd.n492 19.3944
R8393 gnd.n6340 gnd.n492 19.3944
R8394 gnd.n6340 gnd.n490 19.3944
R8395 gnd.n6344 gnd.n490 19.3944
R8396 gnd.n6344 gnd.n486 19.3944
R8397 gnd.n6350 gnd.n486 19.3944
R8398 gnd.n6350 gnd.n484 19.3944
R8399 gnd.n6354 gnd.n484 19.3944
R8400 gnd.n6354 gnd.n480 19.3944
R8401 gnd.n6360 gnd.n480 19.3944
R8402 gnd.n6360 gnd.n478 19.3944
R8403 gnd.n6364 gnd.n478 19.3944
R8404 gnd.n6364 gnd.n474 19.3944
R8405 gnd.n6370 gnd.n474 19.3944
R8406 gnd.n6370 gnd.n472 19.3944
R8407 gnd.n6374 gnd.n472 19.3944
R8408 gnd.n6374 gnd.n468 19.3944
R8409 gnd.n6380 gnd.n468 19.3944
R8410 gnd.n6380 gnd.n466 19.3944
R8411 gnd.n6384 gnd.n466 19.3944
R8412 gnd.n6384 gnd.n462 19.3944
R8413 gnd.n6390 gnd.n462 19.3944
R8414 gnd.n6390 gnd.n460 19.3944
R8415 gnd.n6394 gnd.n460 19.3944
R8416 gnd.n6394 gnd.n456 19.3944
R8417 gnd.n6400 gnd.n456 19.3944
R8418 gnd.n6400 gnd.n454 19.3944
R8419 gnd.n6404 gnd.n454 19.3944
R8420 gnd.n6404 gnd.n450 19.3944
R8421 gnd.n6410 gnd.n450 19.3944
R8422 gnd.n6410 gnd.n448 19.3944
R8423 gnd.n6414 gnd.n448 19.3944
R8424 gnd.n6414 gnd.n444 19.3944
R8425 gnd.n6420 gnd.n444 19.3944
R8426 gnd.n6420 gnd.n442 19.3944
R8427 gnd.n6424 gnd.n442 19.3944
R8428 gnd.n6424 gnd.n438 19.3944
R8429 gnd.n6430 gnd.n438 19.3944
R8430 gnd.n6430 gnd.n436 19.3944
R8431 gnd.n6434 gnd.n436 19.3944
R8432 gnd.n6434 gnd.n432 19.3944
R8433 gnd.n6440 gnd.n432 19.3944
R8434 gnd.n6440 gnd.n430 19.3944
R8435 gnd.n6444 gnd.n430 19.3944
R8436 gnd.n6444 gnd.n426 19.3944
R8437 gnd.n6450 gnd.n426 19.3944
R8438 gnd.n6450 gnd.n424 19.3944
R8439 gnd.n6454 gnd.n424 19.3944
R8440 gnd.n6454 gnd.n420 19.3944
R8441 gnd.n6460 gnd.n420 19.3944
R8442 gnd.n6460 gnd.n418 19.3944
R8443 gnd.n6464 gnd.n418 19.3944
R8444 gnd.n6464 gnd.n414 19.3944
R8445 gnd.n6470 gnd.n414 19.3944
R8446 gnd.n6470 gnd.n412 19.3944
R8447 gnd.n6474 gnd.n412 19.3944
R8448 gnd.n6474 gnd.n408 19.3944
R8449 gnd.n6480 gnd.n408 19.3944
R8450 gnd.n6480 gnd.n406 19.3944
R8451 gnd.n6484 gnd.n406 19.3944
R8452 gnd.n6484 gnd.n402 19.3944
R8453 gnd.n6490 gnd.n402 19.3944
R8454 gnd.n6490 gnd.n400 19.3944
R8455 gnd.n6494 gnd.n400 19.3944
R8456 gnd.n6494 gnd.n396 19.3944
R8457 gnd.n6500 gnd.n396 19.3944
R8458 gnd.n6500 gnd.n394 19.3944
R8459 gnd.n6504 gnd.n394 19.3944
R8460 gnd.n6504 gnd.n390 19.3944
R8461 gnd.n6510 gnd.n390 19.3944
R8462 gnd.n6510 gnd.n388 19.3944
R8463 gnd.n6515 gnd.n388 19.3944
R8464 gnd.n6515 gnd.n384 19.3944
R8465 gnd.n6521 gnd.n384 19.3944
R8466 gnd.n6522 gnd.n6521 19.3944
R8467 gnd.n6164 gnd.n597 19.3944
R8468 gnd.n6164 gnd.n6163 19.3944
R8469 gnd.n6163 gnd.n6162 19.3944
R8470 gnd.n6162 gnd.n601 19.3944
R8471 gnd.n6156 gnd.n601 19.3944
R8472 gnd.n6156 gnd.n6155 19.3944
R8473 gnd.n6155 gnd.n6154 19.3944
R8474 gnd.n6154 gnd.n609 19.3944
R8475 gnd.n6148 gnd.n609 19.3944
R8476 gnd.n6148 gnd.n6147 19.3944
R8477 gnd.n6147 gnd.n6146 19.3944
R8478 gnd.n6146 gnd.n617 19.3944
R8479 gnd.n6140 gnd.n617 19.3944
R8480 gnd.n6140 gnd.n6139 19.3944
R8481 gnd.n6139 gnd.n6138 19.3944
R8482 gnd.n6138 gnd.n625 19.3944
R8483 gnd.n6132 gnd.n625 19.3944
R8484 gnd.n6132 gnd.n6131 19.3944
R8485 gnd.n6131 gnd.n6130 19.3944
R8486 gnd.n6130 gnd.n633 19.3944
R8487 gnd.n6124 gnd.n633 19.3944
R8488 gnd.n6124 gnd.n6123 19.3944
R8489 gnd.n6123 gnd.n6122 19.3944
R8490 gnd.n6122 gnd.n641 19.3944
R8491 gnd.n6116 gnd.n641 19.3944
R8492 gnd.n6116 gnd.n6115 19.3944
R8493 gnd.n6115 gnd.n6114 19.3944
R8494 gnd.n6114 gnd.n649 19.3944
R8495 gnd.n6108 gnd.n649 19.3944
R8496 gnd.n6108 gnd.n6107 19.3944
R8497 gnd.n6107 gnd.n6106 19.3944
R8498 gnd.n6106 gnd.n657 19.3944
R8499 gnd.n6100 gnd.n657 19.3944
R8500 gnd.n6100 gnd.n6099 19.3944
R8501 gnd.n6099 gnd.n6098 19.3944
R8502 gnd.n6098 gnd.n665 19.3944
R8503 gnd.n6092 gnd.n665 19.3944
R8504 gnd.n6092 gnd.n6091 19.3944
R8505 gnd.n6091 gnd.n6090 19.3944
R8506 gnd.n6090 gnd.n673 19.3944
R8507 gnd.n6084 gnd.n673 19.3944
R8508 gnd.n6084 gnd.n6083 19.3944
R8509 gnd.n6083 gnd.n6082 19.3944
R8510 gnd.n6082 gnd.n681 19.3944
R8511 gnd.n6076 gnd.n681 19.3944
R8512 gnd.n6076 gnd.n6075 19.3944
R8513 gnd.n6075 gnd.n6074 19.3944
R8514 gnd.n6074 gnd.n689 19.3944
R8515 gnd.n6068 gnd.n689 19.3944
R8516 gnd.n6068 gnd.n6067 19.3944
R8517 gnd.n6067 gnd.n6066 19.3944
R8518 gnd.n6066 gnd.n697 19.3944
R8519 gnd.n6060 gnd.n697 19.3944
R8520 gnd.n6060 gnd.n6059 19.3944
R8521 gnd.n6059 gnd.n6058 19.3944
R8522 gnd.n6058 gnd.n705 19.3944
R8523 gnd.n6052 gnd.n705 19.3944
R8524 gnd.n6052 gnd.n6051 19.3944
R8525 gnd.n6051 gnd.n6050 19.3944
R8526 gnd.n6050 gnd.n713 19.3944
R8527 gnd.n6044 gnd.n713 19.3944
R8528 gnd.n6044 gnd.n6043 19.3944
R8529 gnd.n6043 gnd.n6042 19.3944
R8530 gnd.n6042 gnd.n721 19.3944
R8531 gnd.n6036 gnd.n721 19.3944
R8532 gnd.n6036 gnd.n6035 19.3944
R8533 gnd.n6035 gnd.n6034 19.3944
R8534 gnd.n6034 gnd.n729 19.3944
R8535 gnd.n6028 gnd.n729 19.3944
R8536 gnd.n6028 gnd.n6027 19.3944
R8537 gnd.n6027 gnd.n6026 19.3944
R8538 gnd.n6026 gnd.n737 19.3944
R8539 gnd.n6020 gnd.n737 19.3944
R8540 gnd.n6020 gnd.n6019 19.3944
R8541 gnd.n6019 gnd.n6018 19.3944
R8542 gnd.n6018 gnd.n745 19.3944
R8543 gnd.n6012 gnd.n745 19.3944
R8544 gnd.n6012 gnd.n6011 19.3944
R8545 gnd.n6011 gnd.n6010 19.3944
R8546 gnd.n6010 gnd.n753 19.3944
R8547 gnd.n6004 gnd.n753 19.3944
R8548 gnd.n6004 gnd.n6003 19.3944
R8549 gnd.n6003 gnd.n6002 19.3944
R8550 gnd.n6002 gnd.n761 19.3944
R8551 gnd.n3437 gnd.n3436 19.3944
R8552 gnd.n3436 gnd.n3435 19.3944
R8553 gnd.n3435 gnd.n3417 19.3944
R8554 gnd.n3431 gnd.n3417 19.3944
R8555 gnd.n3431 gnd.n3430 19.3944
R8556 gnd.n3430 gnd.n3429 19.3944
R8557 gnd.n3429 gnd.n3421 19.3944
R8558 gnd.n3425 gnd.n3421 19.3944
R8559 gnd.n3425 gnd.n3424 19.3944
R8560 gnd.n3424 gnd.n3350 19.3944
R8561 gnd.n4055 gnd.n3350 19.3944
R8562 gnd.n4055 gnd.n3347 19.3944
R8563 gnd.n4059 gnd.n3347 19.3944
R8564 gnd.n4060 gnd.n4059 19.3944
R8565 gnd.n4143 gnd.n4060 19.3944
R8566 gnd.n4143 gnd.n3344 19.3944
R8567 gnd.n4161 gnd.n3344 19.3944
R8568 gnd.n4161 gnd.n3345 19.3944
R8569 gnd.n4157 gnd.n3345 19.3944
R8570 gnd.n4157 gnd.n4156 19.3944
R8571 gnd.n4156 gnd.n4155 19.3944
R8572 gnd.n4155 gnd.n4149 19.3944
R8573 gnd.n4151 gnd.n4149 19.3944
R8574 gnd.n4151 gnd.n3300 19.3944
R8575 gnd.n4246 gnd.n3300 19.3944
R8576 gnd.n4246 gnd.n3301 19.3944
R8577 gnd.n4242 gnd.n3301 19.3944
R8578 gnd.n4242 gnd.n4241 19.3944
R8579 gnd.n4241 gnd.n4240 19.3944
R8580 gnd.n4240 gnd.n4224 19.3944
R8581 gnd.n4236 gnd.n4224 19.3944
R8582 gnd.n4236 gnd.n4235 19.3944
R8583 gnd.n4235 gnd.n4234 19.3944
R8584 gnd.n4234 gnd.n4229 19.3944
R8585 gnd.n4230 gnd.n4229 19.3944
R8586 gnd.n4230 gnd.n3234 19.3944
R8587 gnd.n4375 gnd.n3234 19.3944
R8588 gnd.n4375 gnd.n3231 19.3944
R8589 gnd.n4380 gnd.n3231 19.3944
R8590 gnd.n4380 gnd.n3232 19.3944
R8591 gnd.n3232 gnd.n3212 19.3944
R8592 gnd.n4407 gnd.n3212 19.3944
R8593 gnd.n4407 gnd.n3209 19.3944
R8594 gnd.n4425 gnd.n3209 19.3944
R8595 gnd.n4425 gnd.n3210 19.3944
R8596 gnd.n4421 gnd.n3210 19.3944
R8597 gnd.n4421 gnd.n4420 19.3944
R8598 gnd.n4420 gnd.n4419 19.3944
R8599 gnd.n4419 gnd.n4414 19.3944
R8600 gnd.n4415 gnd.n4414 19.3944
R8601 gnd.n4415 gnd.n3160 19.3944
R8602 gnd.n4517 gnd.n3160 19.3944
R8603 gnd.n4517 gnd.n3157 19.3944
R8604 gnd.n4522 gnd.n3157 19.3944
R8605 gnd.n4522 gnd.n3158 19.3944
R8606 gnd.n3158 gnd.n3136 19.3944
R8607 gnd.n4549 gnd.n3136 19.3944
R8608 gnd.n4549 gnd.n3133 19.3944
R8609 gnd.n4567 gnd.n3133 19.3944
R8610 gnd.n4567 gnd.n3134 19.3944
R8611 gnd.n4563 gnd.n3134 19.3944
R8612 gnd.n4563 gnd.n4562 19.3944
R8613 gnd.n4562 gnd.n4561 19.3944
R8614 gnd.n4561 gnd.n4556 19.3944
R8615 gnd.n4557 gnd.n4556 19.3944
R8616 gnd.n4557 gnd.n3084 19.3944
R8617 gnd.n4643 gnd.n3084 19.3944
R8618 gnd.n4643 gnd.n3081 19.3944
R8619 gnd.n4662 gnd.n3081 19.3944
R8620 gnd.n4662 gnd.n3082 19.3944
R8621 gnd.n4658 gnd.n3082 19.3944
R8622 gnd.n4658 gnd.n4657 19.3944
R8623 gnd.n4657 gnd.n4656 19.3944
R8624 gnd.n4656 gnd.n4651 19.3944
R8625 gnd.n4652 gnd.n4651 19.3944
R8626 gnd.n4652 gnd.n3032 19.3944
R8627 gnd.n4727 gnd.n3032 19.3944
R8628 gnd.n4727 gnd.n3030 19.3944
R8629 gnd.n4731 gnd.n3030 19.3944
R8630 gnd.n4732 gnd.n4731 19.3944
R8631 gnd.n4737 gnd.n4732 19.3944
R8632 gnd.n4737 gnd.n3027 19.3944
R8633 gnd.n4755 gnd.n3027 19.3944
R8634 gnd.n4755 gnd.n3028 19.3944
R8635 gnd.n4751 gnd.n3028 19.3944
R8636 gnd.n4751 gnd.n4750 19.3944
R8637 gnd.n4750 gnd.n4749 19.3944
R8638 gnd.n4749 gnd.n4744 19.3944
R8639 gnd.n4745 gnd.n4744 19.3944
R8640 gnd.n4745 gnd.n2929 19.3944
R8641 gnd.n4990 gnd.n2929 19.3944
R8642 gnd.n4990 gnd.n2927 19.3944
R8643 gnd.n4994 gnd.n2927 19.3944
R8644 gnd.n4994 gnd.n2918 19.3944
R8645 gnd.n5008 gnd.n2918 19.3944
R8646 gnd.n5008 gnd.n2916 19.3944
R8647 gnd.n5012 gnd.n2916 19.3944
R8648 gnd.n5012 gnd.n2906 19.3944
R8649 gnd.n5027 gnd.n2906 19.3944
R8650 gnd.n5027 gnd.n2904 19.3944
R8651 gnd.n5049 gnd.n2904 19.3944
R8652 gnd.n5046 gnd.n5045 19.3944
R8653 gnd.n5045 gnd.n5044 19.3944
R8654 gnd.n5044 gnd.n5033 19.3944
R8655 gnd.n5040 gnd.n5033 19.3944
R8656 gnd.n5040 gnd.n5039 19.3944
R8657 gnd.n5039 gnd.n2876 19.3944
R8658 gnd.n5278 gnd.n2876 19.3944
R8659 gnd.n5278 gnd.n5277 19.3944
R8660 gnd.n5277 gnd.n5276 19.3944
R8661 gnd.n5276 gnd.n2881 19.3944
R8662 gnd.n5269 gnd.n2881 19.3944
R8663 gnd.n5269 gnd.n5268 19.3944
R8664 gnd.n5268 gnd.n5202 19.3944
R8665 gnd.n5261 gnd.n5202 19.3944
R8666 gnd.n5261 gnd.n5260 19.3944
R8667 gnd.n5260 gnd.n5214 19.3944
R8668 gnd.n5253 gnd.n5214 19.3944
R8669 gnd.n5253 gnd.n5252 19.3944
R8670 gnd.n5252 gnd.n5222 19.3944
R8671 gnd.n5245 gnd.n5222 19.3944
R8672 gnd.n5245 gnd.n5244 19.3944
R8673 gnd.n5244 gnd.n5234 19.3944
R8674 gnd.n5234 gnd.n2749 19.3944
R8675 gnd.n5406 gnd.n2749 19.3944
R8676 gnd.n2762 gnd.n2760 19.3944
R8677 gnd.n2762 gnd.n2729 19.3944
R8678 gnd.n5411 gnd.n2729 19.3944
R8679 gnd.n3830 gnd.n2402 19.1199
R8680 gnd.n5718 gnd.n2405 19.1199
R8681 gnd.n5712 gnd.n2416 19.1199
R8682 gnd.n3884 gnd.n3883 19.1199
R8683 gnd.n5706 gnd.n2425 19.1199
R8684 gnd.n3845 gnd.n2433 19.1199
R8685 gnd.n5700 gnd.n2436 19.1199
R8686 gnd.n3849 gnd.n2443 19.1199
R8687 gnd.n5694 gnd.n2446 19.1199
R8688 gnd.n3854 gnd.n2454 19.1199
R8689 gnd.n5688 gnd.n2457 19.1199
R8690 gnd.n5682 gnd.n2467 19.1199
R8691 gnd.n3924 gnd.n3923 19.1199
R8692 gnd.n4383 gnd.t50 19.1199
R8693 gnd.n3117 gnd.t314 19.1199
R8694 gnd.n5192 gnd.n2886 19.1199
R8695 gnd.n5191 gnd.n2890 19.1199
R8696 gnd.n5185 gnd.n5184 19.1199
R8697 gnd.n5160 gnd.n5075 19.1199
R8698 gnd.n5178 gnd.n5092 19.1199
R8699 gnd.n5128 gnd.n5095 19.1199
R8700 gnd.n5170 gnd.n5127 19.1199
R8701 gnd.n6751 gnd.n239 19.1199
R8702 gnd.n5102 gnd.n242 19.1199
R8703 gnd.n6761 gnd.n229 19.1199
R8704 gnd.n6744 gnd.n231 19.1199
R8705 gnd.n6786 gnd.n211 19.1199
R8706 gnd.n6774 gnd.n214 19.1199
R8707 gnd.n1676 gnd.t5 18.8012
R8708 gnd.n1121 gnd.t11 18.8012
R8709 gnd.n7228 gnd.n135 18.8012
R8710 gnd.n1546 gnd.n1545 18.4825
R8711 gnd.n4373 gnd.n3237 18.4825
R8712 gnd.n4447 gnd.n4446 18.4825
R8713 gnd.n4524 gnd.n3147 18.4825
R8714 gnd.n3108 gnd.n3103 18.4825
R8715 gnd.n5345 gnd.n5344 18.4247
R8716 gnd.n5625 gnd.n5624 18.4247
R8717 gnd.n5403 gnd.n5402 18.2308
R8718 gnd.n6942 gnd.n6894 18.2308
R8719 gnd.n3929 gnd.n3928 18.2308
R8720 gnd.n3724 gnd.n3723 18.2308
R8721 gnd.t40 gnd.n1225 18.1639
R8722 gnd.n4163 gnd.t304 17.8452
R8723 gnd.n1254 gnd.t103 17.5266
R8724 gnd.n5620 gnd.t167 17.2079
R8725 gnd.n4141 gnd.n4061 17.2079
R8726 gnd.n3338 gnd.n3333 17.2079
R8727 gnd.n4300 gnd.n4299 17.2079
R8728 gnd.n4363 gnd.n4362 17.2079
R8729 gnd.n3187 gnd.n3181 17.2079
R8730 gnd.n4515 gnd.n3163 17.2079
R8731 gnd.n4629 gnd.n3098 17.2079
R8732 gnd.n4665 gnd.n3071 17.2079
R8733 gnd.n1665 gnd.t56 16.8893
R8734 gnd.n5804 gnd.t236 16.8893
R8735 gnd.t153 gnd.n3245 16.8893
R8736 gnd.n4611 gnd.t32 16.8893
R8737 gnd.n7210 gnd.t194 16.8893
R8738 gnd.n7122 gnd.n7119 16.6793
R8739 gnd.n5327 gnd.n5324 16.6793
R8740 gnd.n5855 gnd.n5852 16.6793
R8741 gnd.n3561 gnd.n3535 16.6793
R8742 gnd.n1481 gnd.t300 16.2519
R8743 gnd.n1713 gnd.t38 16.2519
R8744 gnd.n4165 gnd.n4164 15.9333
R8745 gnd.t204 gnd.n3320 15.9333
R8746 gnd.n3258 gnd.n3252 15.9333
R8747 gnd.n4394 gnd.t77 15.9333
R8748 gnd.n4505 gnd.n4504 15.9333
R8749 gnd.n4504 gnd.n3175 15.9333
R8750 gnd.n4463 gnd.t315 15.9333
R8751 gnd.n4641 gnd.n3087 15.9333
R8752 gnd.n2983 gnd.t240 15.9333
R8753 gnd.n2108 gnd.n2106 15.6674
R8754 gnd.n2076 gnd.n2074 15.6674
R8755 gnd.n2044 gnd.n2042 15.6674
R8756 gnd.n2013 gnd.n2011 15.6674
R8757 gnd.n1981 gnd.n1979 15.6674
R8758 gnd.n1949 gnd.n1947 15.6674
R8759 gnd.n1917 gnd.n1915 15.6674
R8760 gnd.n1886 gnd.n1884 15.6674
R8761 gnd.n1472 gnd.t300 15.6146
R8762 gnd.n2145 gnd.t211 15.6146
R8763 gnd.t310 gnd.n773 15.6146
R8764 gnd.n7203 gnd.n6879 15.3217
R8765 gnd.n5284 gnd.n2870 15.3217
R8766 gnd.n5812 gnd.n2258 15.3217
R8767 gnd.n3615 gnd.n3523 15.3217
R8768 gnd.n4808 gnd.t222 15.296
R8769 gnd.n4817 gnd.t198 15.296
R8770 gnd.n4825 gnd.n4824 15.0827
R8771 gnd.n2591 gnd.n2586 15.0481
R8772 gnd.n4835 gnd.n4834 15.0481
R8773 gnd.n954 gnd.t59 14.9773
R8774 gnd.n2278 gnd.t236 14.9773
R8775 gnd.n3863 gnd.t243 14.9773
R8776 gnd.n4191 gnd.t136 14.9773
R8777 gnd.t158 gnd.n3005 14.9773
R8778 gnd.n5072 gnd.t207 14.9773
R8779 gnd.t194 gnd.n155 14.9773
R8780 gnd.n3333 gnd.n3328 14.6587
R8781 gnd.n4300 gnd.n3264 14.6587
R8782 gnd.n4673 gnd.n3071 14.6587
R8783 gnd.n4786 gnd.n3000 14.6587
R8784 gnd.n4817 gnd.n4816 14.6587
R8785 gnd.n929 gnd.t149 14.34
R8786 gnd.n912 gnd.t104 14.34
R8787 gnd.n4269 gnd.t89 14.0214
R8788 gnd.n4690 gnd.t93 14.0214
R8789 gnd.n1634 gnd.t331 13.7027
R8790 gnd.n1338 gnd.n1337 13.5763
R8791 gnd.n5983 gnd.n786 13.5763
R8792 gnd.n1546 gnd.n1284 13.384
R8793 gnd.n5549 gnd.t201 13.384
R8794 gnd.n4190 gnd.n3324 13.384
R8795 gnd.n4281 gnd.n4279 13.384
R8796 gnd.n3260 gnd.t13 13.384
R8797 gnd.n4311 gnd.n3237 13.384
R8798 gnd.n4447 gnd.n3192 13.384
R8799 gnd.n4537 gnd.n3147 13.384
R8800 gnd.n3109 gnd.n3108 13.384
R8801 gnd.n3089 gnd.t8 13.384
R8802 gnd.n4684 gnd.n4683 13.384
R8803 gnd.n4734 gnd.n4733 13.384
R8804 gnd.n2602 gnd.n2583 13.1884
R8805 gnd.n2597 gnd.n2596 13.1884
R8806 gnd.n2596 gnd.n2595 13.1884
R8807 gnd.n4828 gnd.n4823 13.1884
R8808 gnd.n4829 gnd.n4828 13.1884
R8809 gnd.n2598 gnd.n2585 13.146
R8810 gnd.n2594 gnd.n2585 13.146
R8811 gnd.n4827 gnd.n4826 13.146
R8812 gnd.n4827 gnd.n4822 13.146
R8813 gnd.n2109 gnd.n2105 12.8005
R8814 gnd.n2077 gnd.n2073 12.8005
R8815 gnd.n2045 gnd.n2041 12.8005
R8816 gnd.n2014 gnd.n2010 12.8005
R8817 gnd.n1982 gnd.n1978 12.8005
R8818 gnd.n1950 gnd.n1946 12.8005
R8819 gnd.n1918 gnd.n1914 12.8005
R8820 gnd.n1887 gnd.n1883 12.8005
R8821 gnd.n5718 gnd.n2402 12.7467
R8822 gnd.n3838 gnd.n2405 12.7467
R8823 gnd.n5712 gnd.n2413 12.7467
R8824 gnd.n3883 gnd.n2416 12.7467
R8825 gnd.n3845 gnd.n2425 12.7467
R8826 gnd.n5700 gnd.n2433 12.7467
R8827 gnd.n5694 gnd.n2443 12.7467
R8828 gnd.n3854 gnd.n2446 12.7467
R8829 gnd.n5688 gnd.n2454 12.7467
R8830 gnd.n3863 gnd.n2457 12.7467
R8831 gnd.n5682 gnd.n2464 12.7467
R8832 gnd.n3924 gnd.n2467 12.7467
R8833 gnd.t232 gnd.t226 12.7467
R8834 gnd.n4212 gnd.t164 12.7467
R8835 gnd.t41 gnd.n3036 12.7467
R8836 gnd.n4799 gnd.t261 12.7467
R8837 gnd.n5192 gnd.n5191 12.7467
R8838 gnd.n5071 gnd.n2890 12.7467
R8839 gnd.n5185 gnd.n5072 12.7467
R8840 gnd.n5184 gnd.n5075 12.7467
R8841 gnd.n5160 gnd.n5092 12.7467
R8842 gnd.n5178 gnd.n5095 12.7467
R8843 gnd.n5170 gnd.n239 12.7467
R8844 gnd.n6751 gnd.n242 12.7467
R8845 gnd.n6761 gnd.n231 12.7467
R8846 gnd.n6744 gnd.n6743 12.7467
R8847 gnd.n6770 gnd.n211 12.7467
R8848 gnd.n6786 gnd.n214 12.7467
R8849 gnd.n4022 gnd.t1 12.4281
R8850 gnd.t219 gnd.t322 12.4281
R8851 gnd.n4996 gnd.t96 12.4281
R8852 gnd.n1337 gnd.n1332 12.4126
R8853 gnd.n5979 gnd.n786 12.4126
R8854 gnd.n5617 gnd.n5554 12.1761
R8855 gnd.n4907 gnd.n4906 12.1761
R8856 gnd.n5674 gnd.n2474 12.1094
R8857 gnd.n3313 gnd.n3306 12.1094
R8858 gnd.n4222 gnd.n3283 12.1094
R8859 gnd.n4395 gnd.n3222 12.1094
R8860 gnd.n4427 gnd.n3201 12.1094
R8861 gnd.n4547 gnd.n3138 12.1094
R8862 gnd.n4588 gnd.n3114 12.1094
R8863 gnd.n3056 gnd.n3051 12.1094
R8864 gnd.n4766 gnd.n3013 12.1094
R8865 gnd.n5397 gnd.n2804 12.1094
R8866 gnd.n2113 gnd.n2112 12.0247
R8867 gnd.n2081 gnd.n2080 12.0247
R8868 gnd.n2049 gnd.n2048 12.0247
R8869 gnd.n2018 gnd.n2017 12.0247
R8870 gnd.n1986 gnd.n1985 12.0247
R8871 gnd.n1954 gnd.n1953 12.0247
R8872 gnd.n1922 gnd.n1921 12.0247
R8873 gnd.n1891 gnd.n1890 12.0247
R8874 gnd.t19 gnd.n2291 11.7908
R8875 gnd.n3884 gnd.t123 11.7908
R8876 gnd.n3849 gnd.t69 11.7908
R8877 gnd.n5128 gnd.t26 11.7908
R8878 gnd.t34 gnd.n229 11.7908
R8879 gnd.n143 gnd.t75 11.7908
R8880 gnd.n2116 gnd.n2103 11.249
R8881 gnd.n2084 gnd.n2071 11.249
R8882 gnd.n2052 gnd.n2039 11.249
R8883 gnd.n2021 gnd.n2008 11.249
R8884 gnd.n1989 gnd.n1976 11.249
R8885 gnd.n1957 gnd.n1944 11.249
R8886 gnd.n1925 gnd.n1912 11.249
R8887 gnd.n1894 gnd.n1881 11.249
R8888 gnd.n1624 gnd.t331 11.1535
R8889 gnd.t60 gnd.n2328 11.1535
R8890 gnd.n3830 gnd.t83 11.1535
R8891 gnd.n6774 gnd.t98 11.1535
R8892 gnd.n104 gnd.t114 11.1535
R8893 gnd.n4250 gnd.n4249 10.8348
R8894 gnd.n4362 gnd.t42 10.8348
R8895 gnd.n4405 gnd.n3214 10.8348
R8896 gnd.n4405 gnd.n3215 10.8348
R8897 gnd.n4570 gnd.n4569 10.8348
R8898 gnd.n4569 gnd.n3124 10.8348
R8899 gnd.t28 gnd.n4629 10.8348
R8900 gnd.n3046 gnd.n3035 10.8348
R8901 gnd.n7080 gnd.n6879 10.6672
R8902 gnd.n5287 gnd.n5284 10.6672
R8903 gnd.n5815 gnd.n5812 10.6672
R8904 gnd.n3611 gnd.n3523 10.6672
R8905 gnd.n4975 gnd.n4974 10.6151
R8906 gnd.n4974 gnd.n4971 10.6151
R8907 gnd.n4969 gnd.n4966 10.6151
R8908 gnd.n4966 gnd.n4965 10.6151
R8909 gnd.n4965 gnd.n4962 10.6151
R8910 gnd.n4962 gnd.n4961 10.6151
R8911 gnd.n4961 gnd.n4958 10.6151
R8912 gnd.n4958 gnd.n4957 10.6151
R8913 gnd.n4957 gnd.n4954 10.6151
R8914 gnd.n4954 gnd.n4953 10.6151
R8915 gnd.n4953 gnd.n4950 10.6151
R8916 gnd.n4950 gnd.n4949 10.6151
R8917 gnd.n4949 gnd.n4946 10.6151
R8918 gnd.n4946 gnd.n4945 10.6151
R8919 gnd.n4945 gnd.n4942 10.6151
R8920 gnd.n4942 gnd.n4941 10.6151
R8921 gnd.n4941 gnd.n4938 10.6151
R8922 gnd.n4938 gnd.n4937 10.6151
R8923 gnd.n4937 gnd.n4934 10.6151
R8924 gnd.n4934 gnd.n4933 10.6151
R8925 gnd.n4933 gnd.n4930 10.6151
R8926 gnd.n4930 gnd.n4929 10.6151
R8927 gnd.n4929 gnd.n4926 10.6151
R8928 gnd.n4926 gnd.n4925 10.6151
R8929 gnd.n4925 gnd.n4922 10.6151
R8930 gnd.n4922 gnd.n4921 10.6151
R8931 gnd.n4921 gnd.n4918 10.6151
R8932 gnd.n4918 gnd.n4917 10.6151
R8933 gnd.n4917 gnd.n4914 10.6151
R8934 gnd.n4914 gnd.n4913 10.6151
R8935 gnd.n4130 gnd.n4129 10.6151
R8936 gnd.n4132 gnd.n4130 10.6151
R8937 gnd.n4133 gnd.n4132 10.6151
R8938 gnd.n4135 gnd.n4133 10.6151
R8939 gnd.n4135 gnd.n4134 10.6151
R8940 gnd.n4134 gnd.n3331 10.6151
R8941 gnd.n4173 gnd.n3331 10.6151
R8942 gnd.n4174 gnd.n4173 10.6151
R8943 gnd.n4182 gnd.n4174 10.6151
R8944 gnd.n4182 gnd.n4181 10.6151
R8945 gnd.n4181 gnd.n4180 10.6151
R8946 gnd.n4180 gnd.n4179 10.6151
R8947 gnd.n4179 gnd.n4177 10.6151
R8948 gnd.n4177 gnd.n4176 10.6151
R8949 gnd.n4176 gnd.n3304 10.6151
R8950 gnd.n4214 gnd.n3304 10.6151
R8951 gnd.n4215 gnd.n4214 10.6151
R8952 gnd.n4217 gnd.n4215 10.6151
R8953 gnd.n4218 gnd.n4217 10.6151
R8954 gnd.n4219 gnd.n4218 10.6151
R8955 gnd.n4219 gnd.n3281 10.6151
R8956 gnd.n4271 gnd.n3281 10.6151
R8957 gnd.n4272 gnd.n4271 10.6151
R8958 gnd.n4277 gnd.n4272 10.6151
R8959 gnd.n4277 gnd.n4276 10.6151
R8960 gnd.n4276 gnd.n4275 10.6151
R8961 gnd.n4275 gnd.n4273 10.6151
R8962 gnd.n4273 gnd.n3255 10.6151
R8963 gnd.n4308 gnd.n3255 10.6151
R8964 gnd.n4309 gnd.n4308 10.6151
R8965 gnd.n4349 gnd.n4309 10.6151
R8966 gnd.n4349 gnd.n4348 10.6151
R8967 gnd.n4348 gnd.n4347 10.6151
R8968 gnd.n4347 gnd.n4346 10.6151
R8969 gnd.n4346 gnd.n4310 10.6151
R8970 gnd.n4340 gnd.n4310 10.6151
R8971 gnd.n4340 gnd.n4339 10.6151
R8972 gnd.n4339 gnd.n4338 10.6151
R8973 gnd.n4338 gnd.n4337 10.6151
R8974 gnd.n4337 gnd.n4335 10.6151
R8975 gnd.n4335 gnd.n4334 10.6151
R8976 gnd.n4334 gnd.n4314 10.6151
R8977 gnd.n4327 gnd.n4314 10.6151
R8978 gnd.n4327 gnd.n4326 10.6151
R8979 gnd.n4326 gnd.n4325 10.6151
R8980 gnd.n4325 gnd.n4324 10.6151
R8981 gnd.n4324 gnd.n4322 10.6151
R8982 gnd.n4322 gnd.n4321 10.6151
R8983 gnd.n4321 gnd.n4318 10.6151
R8984 gnd.n4318 gnd.n3184 10.6151
R8985 gnd.n4455 gnd.n3184 10.6151
R8986 gnd.n4456 gnd.n4455 10.6151
R8987 gnd.n4491 gnd.n4456 10.6151
R8988 gnd.n4491 gnd.n4490 10.6151
R8989 gnd.n4490 gnd.n4489 10.6151
R8990 gnd.n4489 gnd.n4488 10.6151
R8991 gnd.n4488 gnd.n4457 10.6151
R8992 gnd.n4483 gnd.n4457 10.6151
R8993 gnd.n4483 gnd.n4482 10.6151
R8994 gnd.n4482 gnd.n4481 10.6151
R8995 gnd.n4481 gnd.n4480 10.6151
R8996 gnd.n4480 gnd.n4478 10.6151
R8997 gnd.n4478 gnd.n4477 10.6151
R8998 gnd.n4477 gnd.n4459 10.6151
R8999 gnd.n4471 gnd.n4459 10.6151
R9000 gnd.n4471 gnd.n4470 10.6151
R9001 gnd.n4470 gnd.n4469 10.6151
R9002 gnd.n4469 gnd.n4468 10.6151
R9003 gnd.n4468 gnd.n4466 10.6151
R9004 gnd.n4466 gnd.n4465 10.6151
R9005 gnd.n4465 gnd.n4462 10.6151
R9006 gnd.n4462 gnd.n3106 10.6151
R9007 gnd.n4596 gnd.n3106 10.6151
R9008 gnd.n4597 gnd.n4596 10.6151
R9009 gnd.n4616 gnd.n4597 10.6151
R9010 gnd.n4616 gnd.n4615 10.6151
R9011 gnd.n4615 gnd.n4614 10.6151
R9012 gnd.n4614 gnd.n4613 10.6151
R9013 gnd.n4613 gnd.n4598 10.6151
R9014 gnd.n4608 gnd.n4598 10.6151
R9015 gnd.n4608 gnd.n4607 10.6151
R9016 gnd.n4607 gnd.n4606 10.6151
R9017 gnd.n4606 gnd.n4605 10.6151
R9018 gnd.n4605 gnd.n4603 10.6151
R9019 gnd.n4603 gnd.n4602 10.6151
R9020 gnd.n4602 gnd.n4600 10.6151
R9021 gnd.n4600 gnd.n3054 10.6151
R9022 gnd.n4692 gnd.n3054 10.6151
R9023 gnd.n4693 gnd.n4692 10.6151
R9024 gnd.n4704 gnd.n4693 10.6151
R9025 gnd.n4704 gnd.n4703 10.6151
R9026 gnd.n4703 gnd.n4702 10.6151
R9027 gnd.n4702 gnd.n4701 10.6151
R9028 gnd.n4701 gnd.n4694 10.6151
R9029 gnd.n4696 gnd.n4694 10.6151
R9030 gnd.n4696 gnd.n4695 10.6151
R9031 gnd.n4695 gnd.n3007 10.6151
R9032 gnd.n4774 gnd.n3007 10.6151
R9033 gnd.n4775 gnd.n4774 10.6151
R9034 gnd.n4777 gnd.n4775 10.6151
R9035 gnd.n4777 gnd.n4776 10.6151
R9036 gnd.n4776 gnd.n2998 10.6151
R9037 gnd.n4789 gnd.n2998 10.6151
R9038 gnd.n4790 gnd.n4789 10.6151
R9039 gnd.n4796 gnd.n4790 10.6151
R9040 gnd.n4796 gnd.n4795 10.6151
R9041 gnd.n4795 gnd.n4794 10.6151
R9042 gnd.n4794 gnd.n4792 10.6151
R9043 gnd.n4792 gnd.n4791 10.6151
R9044 gnd.n4791 gnd.n2975 10.6151
R9045 gnd.n4065 gnd.n2544 10.6151
R9046 gnd.n4068 gnd.n4065 10.6151
R9047 gnd.n4073 gnd.n4070 10.6151
R9048 gnd.n4074 gnd.n4073 10.6151
R9049 gnd.n4077 gnd.n4074 10.6151
R9050 gnd.n4078 gnd.n4077 10.6151
R9051 gnd.n4081 gnd.n4078 10.6151
R9052 gnd.n4082 gnd.n4081 10.6151
R9053 gnd.n4085 gnd.n4082 10.6151
R9054 gnd.n4086 gnd.n4085 10.6151
R9055 gnd.n4089 gnd.n4086 10.6151
R9056 gnd.n4090 gnd.n4089 10.6151
R9057 gnd.n4093 gnd.n4090 10.6151
R9058 gnd.n4094 gnd.n4093 10.6151
R9059 gnd.n4097 gnd.n4094 10.6151
R9060 gnd.n4098 gnd.n4097 10.6151
R9061 gnd.n4101 gnd.n4098 10.6151
R9062 gnd.n4102 gnd.n4101 10.6151
R9063 gnd.n4105 gnd.n4102 10.6151
R9064 gnd.n4106 gnd.n4105 10.6151
R9065 gnd.n4109 gnd.n4106 10.6151
R9066 gnd.n4110 gnd.n4109 10.6151
R9067 gnd.n4113 gnd.n4110 10.6151
R9068 gnd.n4114 gnd.n4113 10.6151
R9069 gnd.n4117 gnd.n4114 10.6151
R9070 gnd.n4118 gnd.n4117 10.6151
R9071 gnd.n4121 gnd.n4118 10.6151
R9072 gnd.n4122 gnd.n4121 10.6151
R9073 gnd.n4125 gnd.n4122 10.6151
R9074 gnd.n4126 gnd.n4125 10.6151
R9075 gnd.n5617 gnd.n5616 10.6151
R9076 gnd.n5616 gnd.n5615 10.6151
R9077 gnd.n5615 gnd.n5614 10.6151
R9078 gnd.n5614 gnd.n5612 10.6151
R9079 gnd.n5612 gnd.n5609 10.6151
R9080 gnd.n5609 gnd.n5608 10.6151
R9081 gnd.n5608 gnd.n5605 10.6151
R9082 gnd.n5605 gnd.n5604 10.6151
R9083 gnd.n5604 gnd.n5601 10.6151
R9084 gnd.n5601 gnd.n5600 10.6151
R9085 gnd.n5600 gnd.n5597 10.6151
R9086 gnd.n5597 gnd.n5596 10.6151
R9087 gnd.n5596 gnd.n5593 10.6151
R9088 gnd.n5593 gnd.n5592 10.6151
R9089 gnd.n5592 gnd.n5589 10.6151
R9090 gnd.n5589 gnd.n5588 10.6151
R9091 gnd.n5588 gnd.n5585 10.6151
R9092 gnd.n5585 gnd.n5584 10.6151
R9093 gnd.n5584 gnd.n5581 10.6151
R9094 gnd.n5581 gnd.n5580 10.6151
R9095 gnd.n5580 gnd.n5577 10.6151
R9096 gnd.n5577 gnd.n5576 10.6151
R9097 gnd.n5576 gnd.n5573 10.6151
R9098 gnd.n5573 gnd.n5572 10.6151
R9099 gnd.n5572 gnd.n5569 10.6151
R9100 gnd.n5569 gnd.n5568 10.6151
R9101 gnd.n5568 gnd.n5565 10.6151
R9102 gnd.n5565 gnd.n5564 10.6151
R9103 gnd.n5561 gnd.n5560 10.6151
R9104 gnd.n5560 gnd.n2545 10.6151
R9105 gnd.n4906 gnd.n4905 10.6151
R9106 gnd.n4905 gnd.n4902 10.6151
R9107 gnd.n4902 gnd.n4901 10.6151
R9108 gnd.n4901 gnd.n4898 10.6151
R9109 gnd.n4898 gnd.n4897 10.6151
R9110 gnd.n4897 gnd.n4894 10.6151
R9111 gnd.n4894 gnd.n4893 10.6151
R9112 gnd.n4893 gnd.n4890 10.6151
R9113 gnd.n4890 gnd.n4889 10.6151
R9114 gnd.n4889 gnd.n4886 10.6151
R9115 gnd.n4886 gnd.n4885 10.6151
R9116 gnd.n4885 gnd.n4882 10.6151
R9117 gnd.n4882 gnd.n4881 10.6151
R9118 gnd.n4881 gnd.n4878 10.6151
R9119 gnd.n4878 gnd.n4877 10.6151
R9120 gnd.n4877 gnd.n4874 10.6151
R9121 gnd.n4874 gnd.n4873 10.6151
R9122 gnd.n4873 gnd.n4870 10.6151
R9123 gnd.n4870 gnd.n4869 10.6151
R9124 gnd.n4869 gnd.n4866 10.6151
R9125 gnd.n4866 gnd.n4865 10.6151
R9126 gnd.n4865 gnd.n4862 10.6151
R9127 gnd.n4862 gnd.n4861 10.6151
R9128 gnd.n4861 gnd.n4858 10.6151
R9129 gnd.n4858 gnd.n4857 10.6151
R9130 gnd.n4857 gnd.n4854 10.6151
R9131 gnd.n4854 gnd.n4853 10.6151
R9132 gnd.n4853 gnd.n4850 10.6151
R9133 gnd.n4848 gnd.n4845 10.6151
R9134 gnd.n4845 gnd.n4844 10.6151
R9135 gnd.n5553 gnd.n5552 10.6151
R9136 gnd.n5552 gnd.n2603 10.6151
R9137 gnd.n4138 gnd.n2603 10.6151
R9138 gnd.n4138 gnd.n3340 10.6151
R9139 gnd.n4167 gnd.n3340 10.6151
R9140 gnd.n4168 gnd.n4167 10.6151
R9141 gnd.n4169 gnd.n4168 10.6151
R9142 gnd.n4169 gnd.n3326 10.6151
R9143 gnd.n4186 gnd.n3326 10.6151
R9144 gnd.n4187 gnd.n4186 10.6151
R9145 gnd.n4188 gnd.n4187 10.6151
R9146 gnd.n4188 gnd.n3308 10.6151
R9147 gnd.n4207 gnd.n3308 10.6151
R9148 gnd.n4208 gnd.n4207 10.6151
R9149 gnd.n4209 gnd.n4208 10.6151
R9150 gnd.n4209 gnd.n3295 10.6151
R9151 gnd.n4252 gnd.n3295 10.6151
R9152 gnd.n4253 gnd.n4252 10.6151
R9153 gnd.n4257 gnd.n4253 10.6151
R9154 gnd.n4257 gnd.n4256 10.6151
R9155 gnd.n4256 gnd.n4255 10.6151
R9156 gnd.n4255 gnd.n3277 10.6151
R9157 gnd.n4284 gnd.n3277 10.6151
R9158 gnd.n4285 gnd.n4284 10.6151
R9159 gnd.n4286 gnd.n4285 10.6151
R9160 gnd.n4286 gnd.n3262 10.6151
R9161 gnd.n4302 gnd.n3262 10.6151
R9162 gnd.n4303 gnd.n4302 10.6151
R9163 gnd.n4304 gnd.n4303 10.6151
R9164 gnd.n4304 gnd.n3250 10.6151
R9165 gnd.n4353 gnd.n3250 10.6151
R9166 gnd.n4354 gnd.n4353 10.6151
R9167 gnd.n4360 gnd.n4354 10.6151
R9168 gnd.n4360 gnd.n4359 10.6151
R9169 gnd.n4359 gnd.n4358 10.6151
R9170 gnd.n4358 gnd.n4355 10.6151
R9171 gnd.n4355 gnd.n3227 10.6151
R9172 gnd.n4385 gnd.n3227 10.6151
R9173 gnd.n4386 gnd.n4385 10.6151
R9174 gnd.n4392 gnd.n4386 10.6151
R9175 gnd.n4392 gnd.n4391 10.6151
R9176 gnd.n4391 gnd.n4390 10.6151
R9177 gnd.n4390 gnd.n4387 10.6151
R9178 gnd.n4387 gnd.n3205 10.6151
R9179 gnd.n4430 gnd.n3205 10.6151
R9180 gnd.n4431 gnd.n4430 10.6151
R9181 gnd.n4432 gnd.n4431 10.6151
R9182 gnd.n4432 gnd.n3190 10.6151
R9183 gnd.n4449 gnd.n3190 10.6151
R9184 gnd.n4450 gnd.n4449 10.6151
R9185 gnd.n4451 gnd.n4450 10.6151
R9186 gnd.n4451 gnd.n3178 10.6151
R9187 gnd.n4495 gnd.n3178 10.6151
R9188 gnd.n4496 gnd.n4495 10.6151
R9189 gnd.n4502 gnd.n4496 10.6151
R9190 gnd.n4502 gnd.n4501 10.6151
R9191 gnd.n4501 gnd.n4500 10.6151
R9192 gnd.n4500 gnd.n4497 10.6151
R9193 gnd.n4497 gnd.n3152 10.6151
R9194 gnd.n4527 gnd.n3152 10.6151
R9195 gnd.n4528 gnd.n4527 10.6151
R9196 gnd.n4534 gnd.n4528 10.6151
R9197 gnd.n4534 gnd.n4533 10.6151
R9198 gnd.n4533 gnd.n4532 10.6151
R9199 gnd.n4532 gnd.n4529 10.6151
R9200 gnd.n4529 gnd.n3128 10.6151
R9201 gnd.n4572 gnd.n3128 10.6151
R9202 gnd.n4573 gnd.n4572 10.6151
R9203 gnd.n4574 gnd.n4573 10.6151
R9204 gnd.n4574 gnd.n3111 10.6151
R9205 gnd.n4590 gnd.n3111 10.6151
R9206 gnd.n4591 gnd.n4590 10.6151
R9207 gnd.n4592 gnd.n4591 10.6151
R9208 gnd.n4592 gnd.n3101 10.6151
R9209 gnd.n4620 gnd.n3101 10.6151
R9210 gnd.n4621 gnd.n4620 10.6151
R9211 gnd.n4627 gnd.n4621 10.6151
R9212 gnd.n4627 gnd.n4626 10.6151
R9213 gnd.n4626 gnd.n4625 10.6151
R9214 gnd.n4625 gnd.n4622 10.6151
R9215 gnd.n4622 gnd.n3076 10.6151
R9216 gnd.n4668 gnd.n3076 10.6151
R9217 gnd.n4669 gnd.n4668 10.6151
R9218 gnd.n4670 gnd.n4669 10.6151
R9219 gnd.n4670 gnd.n3060 10.6151
R9220 gnd.n4686 gnd.n3060 10.6151
R9221 gnd.n4687 gnd.n4686 10.6151
R9222 gnd.n4688 gnd.n4687 10.6151
R9223 gnd.n4688 gnd.n3049 10.6151
R9224 gnd.n4708 gnd.n3049 10.6151
R9225 gnd.n4709 gnd.n4708 10.6151
R9226 gnd.n4713 gnd.n4709 10.6151
R9227 gnd.n4713 gnd.n4712 10.6151
R9228 gnd.n4712 gnd.n4711 10.6151
R9229 gnd.n4711 gnd.n3011 10.6151
R9230 gnd.n4768 gnd.n3011 10.6151
R9231 gnd.n4769 gnd.n4768 10.6151
R9232 gnd.n4770 gnd.n4769 10.6151
R9233 gnd.n4770 gnd.n3002 10.6151
R9234 gnd.n4782 gnd.n3002 10.6151
R9235 gnd.n4783 gnd.n4782 10.6151
R9236 gnd.n4784 gnd.n4783 10.6151
R9237 gnd.n4784 gnd.n2993 10.6151
R9238 gnd.n4802 gnd.n2993 10.6151
R9239 gnd.n4803 gnd.n4802 10.6151
R9240 gnd.n4804 gnd.n4803 10.6151
R9241 gnd.n4804 gnd.n2979 10.6151
R9242 gnd.n4819 gnd.n2979 10.6151
R9243 gnd.n4820 gnd.n4819 10.6151
R9244 gnd.n4908 gnd.n4820 10.6151
R9245 gnd.n1535 gnd.t24 10.5161
R9246 gnd.n1846 gnd.t149 10.5161
R9247 gnd.t104 gnd.n901 10.5161
R9248 gnd.n2363 gnd.t86 10.5161
R9249 gnd.t21 gnd.n2366 10.5161
R9250 gnd.n6829 gnd.t140 10.5161
R9251 gnd.n6837 gnd.t52 10.5161
R9252 gnd.n2117 gnd.n2101 10.4732
R9253 gnd.n2085 gnd.n2069 10.4732
R9254 gnd.n2053 gnd.n2037 10.4732
R9255 gnd.n2022 gnd.n2006 10.4732
R9256 gnd.n1990 gnd.n1974 10.4732
R9257 gnd.n1958 gnd.n1942 10.4732
R9258 gnd.n1926 gnd.n1910 10.4732
R9259 gnd.n1895 gnd.n1879 10.4732
R9260 gnd.n1815 gnd.t59 9.87883
R9261 gnd.n2325 gnd.t36 9.87883
R9262 gnd.n3838 gnd.t132 9.87883
R9263 gnd.t78 gnd.t116 9.87883
R9264 gnd.t16 gnd.t138 9.87883
R9265 gnd.n6770 gnd.t14 9.87883
R9266 gnd.t54 gnd.n107 9.87883
R9267 gnd.n2121 gnd.n2120 9.69747
R9268 gnd.n2089 gnd.n2088 9.69747
R9269 gnd.n2057 gnd.n2056 9.69747
R9270 gnd.n2026 gnd.n2025 9.69747
R9271 gnd.n1994 gnd.n1993 9.69747
R9272 gnd.n1962 gnd.n1961 9.69747
R9273 gnd.n1930 gnd.n1929 9.69747
R9274 gnd.n1899 gnd.n1898 9.69747
R9275 gnd.n4211 gnd.n3306 9.56018
R9276 gnd.n4222 gnd.n4221 9.56018
R9277 gnd.n4395 gnd.n4394 9.56018
R9278 gnd.n4428 gnd.n4427 9.56018
R9279 gnd.n4547 gnd.n3139 9.56018
R9280 gnd.n4463 gnd.n3114 9.56018
R9281 gnd.n4706 gnd.n3051 9.56018
R9282 gnd.n4697 gnd.n3013 9.56018
R9283 gnd.n2127 gnd.n2126 9.45567
R9284 gnd.n2095 gnd.n2094 9.45567
R9285 gnd.n2063 gnd.n2062 9.45567
R9286 gnd.n2032 gnd.n2031 9.45567
R9287 gnd.n2000 gnd.n1999 9.45567
R9288 gnd.n1968 gnd.n1967 9.45567
R9289 gnd.n1936 gnd.n1935 9.45567
R9290 gnd.n1905 gnd.n1904 9.45567
R9291 gnd.n7119 gnd.n7059 9.30959
R9292 gnd.n5324 gnd.n5323 9.30959
R9293 gnd.n5852 gnd.n5851 9.30959
R9294 gnd.n3565 gnd.n3535 9.30959
R9295 gnd.n5284 gnd.n5283 9.3005
R9296 gnd.n5287 gnd.n2869 9.3005
R9297 gnd.n5288 gnd.n2868 9.3005
R9298 gnd.n5291 gnd.n2867 9.3005
R9299 gnd.n5292 gnd.n2866 9.3005
R9300 gnd.n5295 gnd.n2865 9.3005
R9301 gnd.n5296 gnd.n2864 9.3005
R9302 gnd.n5299 gnd.n2863 9.3005
R9303 gnd.n5300 gnd.n2862 9.3005
R9304 gnd.n5303 gnd.n2861 9.3005
R9305 gnd.n5304 gnd.n2860 9.3005
R9306 gnd.n5307 gnd.n2859 9.3005
R9307 gnd.n5308 gnd.n2858 9.3005
R9308 gnd.n5311 gnd.n2857 9.3005
R9309 gnd.n5312 gnd.n2856 9.3005
R9310 gnd.n5315 gnd.n2855 9.3005
R9311 gnd.n5316 gnd.n2854 9.3005
R9312 gnd.n5319 gnd.n2853 9.3005
R9313 gnd.n5320 gnd.n2852 9.3005
R9314 gnd.n5323 gnd.n2851 9.3005
R9315 gnd.n5327 gnd.n2847 9.3005
R9316 gnd.n5328 gnd.n2846 9.3005
R9317 gnd.n5331 gnd.n2845 9.3005
R9318 gnd.n5332 gnd.n2844 9.3005
R9319 gnd.n5335 gnd.n2843 9.3005
R9320 gnd.n5336 gnd.n2842 9.3005
R9321 gnd.n5339 gnd.n2841 9.3005
R9322 gnd.n5340 gnd.n2840 9.3005
R9323 gnd.n5343 gnd.n2839 9.3005
R9324 gnd.n5345 gnd.n2835 9.3005
R9325 gnd.n5348 gnd.n2834 9.3005
R9326 gnd.n5349 gnd.n2833 9.3005
R9327 gnd.n5352 gnd.n2832 9.3005
R9328 gnd.n5353 gnd.n2831 9.3005
R9329 gnd.n5356 gnd.n2830 9.3005
R9330 gnd.n5357 gnd.n2829 9.3005
R9331 gnd.n5360 gnd.n2828 9.3005
R9332 gnd.n5362 gnd.n2825 9.3005
R9333 gnd.n5365 gnd.n2824 9.3005
R9334 gnd.n5366 gnd.n2823 9.3005
R9335 gnd.n5369 gnd.n2822 9.3005
R9336 gnd.n5370 gnd.n2821 9.3005
R9337 gnd.n5373 gnd.n2820 9.3005
R9338 gnd.n5374 gnd.n2819 9.3005
R9339 gnd.n5377 gnd.n2818 9.3005
R9340 gnd.n5378 gnd.n2817 9.3005
R9341 gnd.n5381 gnd.n2816 9.3005
R9342 gnd.n5382 gnd.n2815 9.3005
R9343 gnd.n5385 gnd.n2814 9.3005
R9344 gnd.n5386 gnd.n2813 9.3005
R9345 gnd.n5389 gnd.n2812 9.3005
R9346 gnd.n5391 gnd.n2811 9.3005
R9347 gnd.n5392 gnd.n2810 9.3005
R9348 gnd.n5393 gnd.n2809 9.3005
R9349 gnd.n5394 gnd.n2808 9.3005
R9350 gnd.n5324 gnd.n2848 9.3005
R9351 gnd.n5282 gnd.n2870 9.3005
R9352 gnd.n5084 gnd.n5083 9.3005
R9353 gnd.n5085 gnd.n5079 9.3005
R9354 gnd.n5182 gnd.n5086 9.3005
R9355 gnd.n5181 gnd.n5087 9.3005
R9356 gnd.n5180 gnd.n5088 9.3005
R9357 gnd.n5090 gnd.n5089 9.3005
R9358 gnd.n237 gnd.n236 9.3005
R9359 gnd.n6754 gnd.n6753 9.3005
R9360 gnd.n6755 gnd.n235 9.3005
R9361 gnd.n6759 gnd.n6756 9.3005
R9362 gnd.n6758 gnd.n6757 9.3005
R9363 gnd.n209 gnd.n208 9.3005
R9364 gnd.n6789 gnd.n6788 9.3005
R9365 gnd.n6790 gnd.n207 9.3005
R9366 gnd.n6794 gnd.n6791 9.3005
R9367 gnd.n6793 gnd.n6792 9.3005
R9368 gnd.n5081 gnd.n5080 9.3005
R9369 gnd.n185 gnd.n184 9.3005
R9370 gnd.n6821 gnd.n6820 9.3005
R9371 gnd.n6822 gnd.n183 9.3005
R9372 gnd.n6827 gnd.n6823 9.3005
R9373 gnd.n6826 gnd.n6825 9.3005
R9374 gnd.n6824 gnd.n78 9.3005
R9375 gnd.n7262 gnd.n79 9.3005
R9376 gnd.n7261 gnd.n80 9.3005
R9377 gnd.n7260 gnd.n81 9.3005
R9378 gnd.n98 gnd.n82 9.3005
R9379 gnd.n7250 gnd.n99 9.3005
R9380 gnd.n7249 gnd.n100 9.3005
R9381 gnd.n7248 gnd.n101 9.3005
R9382 gnd.n118 gnd.n102 9.3005
R9383 gnd.n7238 gnd.n119 9.3005
R9384 gnd.n7237 gnd.n120 9.3005
R9385 gnd.n7236 gnd.n121 9.3005
R9386 gnd.n137 gnd.n122 9.3005
R9387 gnd.n7226 gnd.n138 9.3005
R9388 gnd.n7225 gnd.n139 9.3005
R9389 gnd.n7224 gnd.n140 9.3005
R9390 gnd.n157 gnd.n141 9.3005
R9391 gnd.n7214 gnd.n158 9.3005
R9392 gnd.n7213 gnd.n159 9.3005
R9393 gnd.n7212 gnd.n160 9.3005
R9394 gnd.n7023 gnd.n161 9.3005
R9395 gnd.n7268 gnd.n7267 9.3005
R9396 gnd.n7266 gnd.n69 9.3005
R9397 gnd.n6953 gnd.n71 9.3005
R9398 gnd.n6955 gnd.n6954 9.3005
R9399 gnd.n6958 gnd.n6957 9.3005
R9400 gnd.n6959 gnd.n6952 9.3005
R9401 gnd.n6962 gnd.n6960 9.3005
R9402 gnd.n6963 gnd.n6951 9.3005
R9403 gnd.n6966 gnd.n6965 9.3005
R9404 gnd.n6967 gnd.n6950 9.3005
R9405 gnd.n6970 gnd.n6968 9.3005
R9406 gnd.n6971 gnd.n6949 9.3005
R9407 gnd.n6974 gnd.n6973 9.3005
R9408 gnd.n6975 gnd.n6948 9.3005
R9409 gnd.n6978 gnd.n6976 9.3005
R9410 gnd.n6979 gnd.n6947 9.3005
R9411 gnd.n6982 gnd.n6981 9.3005
R9412 gnd.n6983 gnd.n6946 9.3005
R9413 gnd.n6986 gnd.n6984 9.3005
R9414 gnd.n6987 gnd.n6945 9.3005
R9415 gnd.n6989 gnd.n6988 9.3005
R9416 gnd.n6905 gnd.n6904 9.3005
R9417 gnd.n6907 gnd.n6906 9.3005
R9418 gnd.n6910 gnd.n6901 9.3005
R9419 gnd.n6914 gnd.n6913 9.3005
R9420 gnd.n6915 gnd.n6900 9.3005
R9421 gnd.n6917 gnd.n6916 9.3005
R9422 gnd.n6920 gnd.n6899 9.3005
R9423 gnd.n6924 gnd.n6923 9.3005
R9424 gnd.n6925 gnd.n6898 9.3005
R9425 gnd.n6927 gnd.n6926 9.3005
R9426 gnd.n6930 gnd.n6897 9.3005
R9427 gnd.n6934 gnd.n6933 9.3005
R9428 gnd.n6935 gnd.n6896 9.3005
R9429 gnd.n6937 gnd.n6936 9.3005
R9430 gnd.n6940 gnd.n6895 9.3005
R9431 gnd.n6943 gnd.n6942 9.3005
R9432 gnd.n6944 gnd.n6894 9.3005
R9433 gnd.n6991 gnd.n6990 9.3005
R9434 gnd.n6902 gnd.n6875 9.3005
R9435 gnd.n7196 gnd.n7195 9.3005
R9436 gnd.n7194 gnd.n7025 9.3005
R9437 gnd.n7193 gnd.n7192 9.3005
R9438 gnd.n7189 gnd.n7026 9.3005
R9439 gnd.n7186 gnd.n7027 9.3005
R9440 gnd.n7185 gnd.n7028 9.3005
R9441 gnd.n7182 gnd.n7029 9.3005
R9442 gnd.n7181 gnd.n7030 9.3005
R9443 gnd.n7178 gnd.n7031 9.3005
R9444 gnd.n7177 gnd.n7032 9.3005
R9445 gnd.n7174 gnd.n7033 9.3005
R9446 gnd.n7173 gnd.n7034 9.3005
R9447 gnd.n7170 gnd.n7035 9.3005
R9448 gnd.n7169 gnd.n7036 9.3005
R9449 gnd.n7166 gnd.n7037 9.3005
R9450 gnd.n7165 gnd.n7038 9.3005
R9451 gnd.n7162 gnd.n7039 9.3005
R9452 gnd.n7158 gnd.n7040 9.3005
R9453 gnd.n7155 gnd.n7041 9.3005
R9454 gnd.n7154 gnd.n7042 9.3005
R9455 gnd.n7151 gnd.n7043 9.3005
R9456 gnd.n7150 gnd.n7044 9.3005
R9457 gnd.n7147 gnd.n7045 9.3005
R9458 gnd.n7146 gnd.n7046 9.3005
R9459 gnd.n7143 gnd.n7047 9.3005
R9460 gnd.n7142 gnd.n7048 9.3005
R9461 gnd.n7139 gnd.n7049 9.3005
R9462 gnd.n7138 gnd.n7050 9.3005
R9463 gnd.n7135 gnd.n7051 9.3005
R9464 gnd.n7134 gnd.n7052 9.3005
R9465 gnd.n7131 gnd.n7053 9.3005
R9466 gnd.n7130 gnd.n7054 9.3005
R9467 gnd.n7127 gnd.n7055 9.3005
R9468 gnd.n7126 gnd.n7056 9.3005
R9469 gnd.n7123 gnd.n7057 9.3005
R9470 gnd.n7122 gnd.n7058 9.3005
R9471 gnd.n7119 gnd.n7118 9.3005
R9472 gnd.n7117 gnd.n7059 9.3005
R9473 gnd.n7116 gnd.n7115 9.3005
R9474 gnd.n7112 gnd.n7062 9.3005
R9475 gnd.n7109 gnd.n7063 9.3005
R9476 gnd.n7108 gnd.n7064 9.3005
R9477 gnd.n7105 gnd.n7065 9.3005
R9478 gnd.n7104 gnd.n7066 9.3005
R9479 gnd.n7101 gnd.n7067 9.3005
R9480 gnd.n7100 gnd.n7068 9.3005
R9481 gnd.n7097 gnd.n7069 9.3005
R9482 gnd.n7096 gnd.n7070 9.3005
R9483 gnd.n7093 gnd.n7071 9.3005
R9484 gnd.n7092 gnd.n7072 9.3005
R9485 gnd.n7089 gnd.n7073 9.3005
R9486 gnd.n7088 gnd.n7074 9.3005
R9487 gnd.n7085 gnd.n7075 9.3005
R9488 gnd.n7084 gnd.n7076 9.3005
R9489 gnd.n7081 gnd.n7077 9.3005
R9490 gnd.n7080 gnd.n7078 9.3005
R9491 gnd.n6879 gnd.n6876 9.3005
R9492 gnd.n7204 gnd.n7203 9.3005
R9493 gnd.n7197 gnd.n7024 9.3005
R9494 gnd.n5150 gnd.n5149 9.3005
R9495 gnd.n5148 gnd.n5144 9.3005
R9496 gnd.n5155 gnd.n5143 9.3005
R9497 gnd.n5158 gnd.n5156 9.3005
R9498 gnd.n5157 gnd.n5099 9.3005
R9499 gnd.n5174 gnd.n5100 9.3005
R9500 gnd.n5173 gnd.n5172 9.3005
R9501 gnd.n5105 gnd.n246 9.3005
R9502 gnd.n5104 gnd.n247 9.3005
R9503 gnd.n5101 gnd.n248 9.3005
R9504 gnd.n249 gnd.n220 9.3005
R9505 gnd.n6772 gnd.n221 9.3005
R9506 gnd.n6773 gnd.n218 9.3005
R9507 gnd.n6776 gnd.n219 9.3005
R9508 gnd.n6778 gnd.n6777 9.3005
R9509 gnd.n6779 gnd.n193 9.3005
R9510 gnd.n6811 gnd.n192 9.3005
R9511 gnd.n6815 gnd.n6814 9.3005
R9512 gnd.n6813 gnd.n175 9.3005
R9513 gnd.n6832 gnd.n174 9.3005
R9514 gnd.n6834 gnd.n6833 9.3005
R9515 gnd.n6835 gnd.n169 9.3005
R9516 gnd.n6841 gnd.n168 9.3005
R9517 gnd.n6844 gnd.n6842 9.3005
R9518 gnd.n6845 gnd.n90 9.3005
R9519 gnd.n6847 gnd.n91 9.3005
R9520 gnd.n6848 gnd.n92 9.3005
R9521 gnd.n6851 gnd.n6849 9.3005
R9522 gnd.n6852 gnd.n109 9.3005
R9523 gnd.n6854 gnd.n110 9.3005
R9524 gnd.n6855 gnd.n111 9.3005
R9525 gnd.n6858 gnd.n6856 9.3005
R9526 gnd.n6859 gnd.n128 9.3005
R9527 gnd.n6861 gnd.n129 9.3005
R9528 gnd.n6862 gnd.n130 9.3005
R9529 gnd.n6865 gnd.n6863 9.3005
R9530 gnd.n6866 gnd.n148 9.3005
R9531 gnd.n6868 gnd.n149 9.3005
R9532 gnd.n6869 gnd.n150 9.3005
R9533 gnd.n6872 gnd.n6870 9.3005
R9534 gnd.n6873 gnd.n167 9.3005
R9535 gnd.n7206 gnd.n6874 9.3005
R9536 gnd.n5145 gnd.n2873 9.3005
R9537 gnd.n5151 gnd.n5150 9.3005
R9538 gnd.n5153 gnd.n5144 9.3005
R9539 gnd.n5155 gnd.n5154 9.3005
R9540 gnd.n5156 gnd.n5098 9.3005
R9541 gnd.n5176 gnd.n5099 9.3005
R9542 gnd.n5175 gnd.n5174 9.3005
R9543 gnd.n5173 gnd.n245 9.3005
R9544 gnd.n6749 gnd.n246 9.3005
R9545 gnd.n6748 gnd.n247 9.3005
R9546 gnd.n6747 gnd.n248 9.3005
R9547 gnd.n6746 gnd.n249 9.3005
R9548 gnd.n221 gnd.n217 9.3005
R9549 gnd.n6784 gnd.n218 9.3005
R9550 gnd.n6783 gnd.n219 9.3005
R9551 gnd.n6782 gnd.n6778 9.3005
R9552 gnd.n6781 gnd.n6779 9.3005
R9553 gnd.n192 gnd.n191 9.3005
R9554 gnd.n6816 gnd.n6815 9.3005
R9555 gnd.n176 gnd.n175 9.3005
R9556 gnd.n6832 gnd.n6831 9.3005
R9557 gnd.n6833 gnd.n170 9.3005
R9558 gnd.n6839 gnd.n169 9.3005
R9559 gnd.n6841 gnd.n6840 9.3005
R9560 gnd.n6842 gnd.n89 9.3005
R9561 gnd.n7256 gnd.n90 9.3005
R9562 gnd.n7255 gnd.n91 9.3005
R9563 gnd.n7254 gnd.n92 9.3005
R9564 gnd.n6849 gnd.n93 9.3005
R9565 gnd.n7244 gnd.n109 9.3005
R9566 gnd.n7243 gnd.n110 9.3005
R9567 gnd.n7242 gnd.n111 9.3005
R9568 gnd.n6856 gnd.n112 9.3005
R9569 gnd.n7232 gnd.n128 9.3005
R9570 gnd.n7231 gnd.n129 9.3005
R9571 gnd.n7230 gnd.n130 9.3005
R9572 gnd.n6863 gnd.n131 9.3005
R9573 gnd.n7220 gnd.n148 9.3005
R9574 gnd.n7219 gnd.n149 9.3005
R9575 gnd.n7218 gnd.n150 9.3005
R9576 gnd.n6870 gnd.n151 9.3005
R9577 gnd.n7208 gnd.n167 9.3005
R9578 gnd.n7207 gnd.n7206 9.3005
R9579 gnd.n2885 gnd.n2873 9.3005
R9580 gnd.n2126 gnd.n2125 9.3005
R9581 gnd.n2099 gnd.n2098 9.3005
R9582 gnd.n2120 gnd.n2119 9.3005
R9583 gnd.n2118 gnd.n2117 9.3005
R9584 gnd.n2103 gnd.n2102 9.3005
R9585 gnd.n2112 gnd.n2111 9.3005
R9586 gnd.n2110 gnd.n2109 9.3005
R9587 gnd.n2094 gnd.n2093 9.3005
R9588 gnd.n2067 gnd.n2066 9.3005
R9589 gnd.n2088 gnd.n2087 9.3005
R9590 gnd.n2086 gnd.n2085 9.3005
R9591 gnd.n2071 gnd.n2070 9.3005
R9592 gnd.n2080 gnd.n2079 9.3005
R9593 gnd.n2078 gnd.n2077 9.3005
R9594 gnd.n2062 gnd.n2061 9.3005
R9595 gnd.n2035 gnd.n2034 9.3005
R9596 gnd.n2056 gnd.n2055 9.3005
R9597 gnd.n2054 gnd.n2053 9.3005
R9598 gnd.n2039 gnd.n2038 9.3005
R9599 gnd.n2048 gnd.n2047 9.3005
R9600 gnd.n2046 gnd.n2045 9.3005
R9601 gnd.n2031 gnd.n2030 9.3005
R9602 gnd.n2004 gnd.n2003 9.3005
R9603 gnd.n2025 gnd.n2024 9.3005
R9604 gnd.n2023 gnd.n2022 9.3005
R9605 gnd.n2008 gnd.n2007 9.3005
R9606 gnd.n2017 gnd.n2016 9.3005
R9607 gnd.n2015 gnd.n2014 9.3005
R9608 gnd.n1999 gnd.n1998 9.3005
R9609 gnd.n1972 gnd.n1971 9.3005
R9610 gnd.n1993 gnd.n1992 9.3005
R9611 gnd.n1991 gnd.n1990 9.3005
R9612 gnd.n1976 gnd.n1975 9.3005
R9613 gnd.n1985 gnd.n1984 9.3005
R9614 gnd.n1983 gnd.n1982 9.3005
R9615 gnd.n1967 gnd.n1966 9.3005
R9616 gnd.n1940 gnd.n1939 9.3005
R9617 gnd.n1961 gnd.n1960 9.3005
R9618 gnd.n1959 gnd.n1958 9.3005
R9619 gnd.n1944 gnd.n1943 9.3005
R9620 gnd.n1953 gnd.n1952 9.3005
R9621 gnd.n1951 gnd.n1950 9.3005
R9622 gnd.n1935 gnd.n1934 9.3005
R9623 gnd.n1908 gnd.n1907 9.3005
R9624 gnd.n1929 gnd.n1928 9.3005
R9625 gnd.n1927 gnd.n1926 9.3005
R9626 gnd.n1912 gnd.n1911 9.3005
R9627 gnd.n1921 gnd.n1920 9.3005
R9628 gnd.n1919 gnd.n1918 9.3005
R9629 gnd.n1904 gnd.n1903 9.3005
R9630 gnd.n1877 gnd.n1876 9.3005
R9631 gnd.n1898 gnd.n1897 9.3005
R9632 gnd.n1896 gnd.n1895 9.3005
R9633 gnd.n1881 gnd.n1880 9.3005
R9634 gnd.n1890 gnd.n1889 9.3005
R9635 gnd.n1888 gnd.n1887 9.3005
R9636 gnd.n5972 gnd.n5971 9.3005
R9637 gnd.n5970 gnd.n5938 9.3005
R9638 gnd.n5969 gnd.n5968 9.3005
R9639 gnd.n5965 gnd.n5939 9.3005
R9640 gnd.n5962 gnd.n5940 9.3005
R9641 gnd.n5961 gnd.n5941 9.3005
R9642 gnd.n5958 gnd.n5942 9.3005
R9643 gnd.n5957 gnd.n5943 9.3005
R9644 gnd.n5954 gnd.n5944 9.3005
R9645 gnd.n5953 gnd.n5945 9.3005
R9646 gnd.n5950 gnd.n5946 9.3005
R9647 gnd.n5949 gnd.n5947 9.3005
R9648 gnd.n788 gnd.n787 9.3005
R9649 gnd.n5980 gnd.n5979 9.3005
R9650 gnd.n5981 gnd.n786 9.3005
R9651 gnd.n5983 gnd.n5982 9.3005
R9652 gnd.n5973 gnd.n5937 9.3005
R9653 gnd.n1554 gnd.n1553 9.3005
R9654 gnd.n1258 gnd.n1257 9.3005
R9655 gnd.n1581 gnd.n1580 9.3005
R9656 gnd.n1582 gnd.n1256 9.3005
R9657 gnd.n1586 gnd.n1583 9.3005
R9658 gnd.n1585 gnd.n1584 9.3005
R9659 gnd.n1230 gnd.n1229 9.3005
R9660 gnd.n1611 gnd.n1610 9.3005
R9661 gnd.n1612 gnd.n1228 9.3005
R9662 gnd.n1622 gnd.n1613 9.3005
R9663 gnd.n1621 gnd.n1614 9.3005
R9664 gnd.n1620 gnd.n1615 9.3005
R9665 gnd.n1618 gnd.n1617 9.3005
R9666 gnd.n1616 gnd.n1200 9.3005
R9667 gnd.n1198 gnd.n1197 9.3005
R9668 gnd.n1670 gnd.n1669 9.3005
R9669 gnd.n1671 gnd.n1196 9.3005
R9670 gnd.n1673 gnd.n1672 9.3005
R9671 gnd.n1033 gnd.n1032 9.3005
R9672 gnd.n1706 gnd.n1705 9.3005
R9673 gnd.n1707 gnd.n1031 9.3005
R9674 gnd.n1711 gnd.n1708 9.3005
R9675 gnd.n1710 gnd.n1709 9.3005
R9676 gnd.n1009 gnd.n1008 9.3005
R9677 gnd.n1737 gnd.n1736 9.3005
R9678 gnd.n1738 gnd.n1007 9.3005
R9679 gnd.n1742 gnd.n1739 9.3005
R9680 gnd.n1741 gnd.n1740 9.3005
R9681 gnd.n983 gnd.n982 9.3005
R9682 gnd.n1768 gnd.n1767 9.3005
R9683 gnd.n1769 gnd.n981 9.3005
R9684 gnd.n1773 gnd.n1770 9.3005
R9685 gnd.n1772 gnd.n1771 9.3005
R9686 gnd.n958 gnd.n957 9.3005
R9687 gnd.n1799 gnd.n1798 9.3005
R9688 gnd.n1800 gnd.n956 9.3005
R9689 gnd.n1804 gnd.n1801 9.3005
R9690 gnd.n1803 gnd.n1802 9.3005
R9691 gnd.n933 gnd.n932 9.3005
R9692 gnd.n1830 gnd.n1829 9.3005
R9693 gnd.n1831 gnd.n931 9.3005
R9694 gnd.n1835 gnd.n1832 9.3005
R9695 gnd.n1834 gnd.n1833 9.3005
R9696 gnd.n907 gnd.n906 9.3005
R9697 gnd.n1861 gnd.n1860 9.3005
R9698 gnd.n1862 gnd.n905 9.3005
R9699 gnd.n1867 gnd.n1863 9.3005
R9700 gnd.n1866 gnd.n1865 9.3005
R9701 gnd.n1864 gnd.n767 9.3005
R9702 gnd.n5996 gnd.n768 9.3005
R9703 gnd.n5995 gnd.n769 9.3005
R9704 gnd.n5994 gnd.n770 9.3005
R9705 gnd.n5936 gnd.n771 9.3005
R9706 gnd.n1555 gnd.n1552 9.3005
R9707 gnd.n1337 gnd.n1296 9.3005
R9708 gnd.n1332 gnd.n1331 9.3005
R9709 gnd.n1330 gnd.n1297 9.3005
R9710 gnd.n1329 gnd.n1328 9.3005
R9711 gnd.n1325 gnd.n1298 9.3005
R9712 gnd.n1322 gnd.n1321 9.3005
R9713 gnd.n1320 gnd.n1299 9.3005
R9714 gnd.n1319 gnd.n1318 9.3005
R9715 gnd.n1315 gnd.n1300 9.3005
R9716 gnd.n1312 gnd.n1311 9.3005
R9717 gnd.n1310 gnd.n1301 9.3005
R9718 gnd.n1309 gnd.n1308 9.3005
R9719 gnd.n1305 gnd.n1303 9.3005
R9720 gnd.n1302 gnd.n1282 9.3005
R9721 gnd.n1549 gnd.n1281 9.3005
R9722 gnd.n1551 gnd.n1550 9.3005
R9723 gnd.n1339 gnd.n1338 9.3005
R9724 gnd.n1562 gnd.n1268 9.3005
R9725 gnd.n1569 gnd.n1269 9.3005
R9726 gnd.n1571 gnd.n1570 9.3005
R9727 gnd.n1572 gnd.n1249 9.3005
R9728 gnd.n1591 gnd.n1590 9.3005
R9729 gnd.n1593 gnd.n1241 9.3005
R9730 gnd.n1600 gnd.n1243 9.3005
R9731 gnd.n1601 gnd.n1238 9.3005
R9732 gnd.n1603 gnd.n1602 9.3005
R9733 gnd.n1239 gnd.n1224 9.3005
R9734 gnd.n1222 gnd.n1220 9.3005
R9735 gnd.n1629 gnd.n1628 9.3005
R9736 gnd.n1205 gnd.n1204 9.3005
R9737 gnd.n1662 gnd.n1650 9.3005
R9738 gnd.n1661 gnd.n1652 9.3005
R9739 gnd.n1660 gnd.n1653 9.3005
R9740 gnd.n1655 gnd.n1654 9.3005
R9741 gnd.n1188 gnd.n1042 9.3005
R9742 gnd.n1694 gnd.n1043 9.3005
R9743 gnd.n1696 gnd.n1695 9.3005
R9744 gnd.n1697 gnd.n1026 9.3005
R9745 gnd.n1716 gnd.n1715 9.3005
R9746 gnd.n1718 gnd.n1019 9.3005
R9747 gnd.n1725 gnd.n1020 9.3005
R9748 gnd.n1727 gnd.n1726 9.3005
R9749 gnd.n1728 gnd.n1001 9.3005
R9750 gnd.n1747 gnd.n1746 9.3005
R9751 gnd.n1749 gnd.n993 9.3005
R9752 gnd.n1756 gnd.n994 9.3005
R9753 gnd.n1758 gnd.n1757 9.3005
R9754 gnd.n1759 gnd.n974 9.3005
R9755 gnd.n1778 gnd.n1777 9.3005
R9756 gnd.n1780 gnd.n967 9.3005
R9757 gnd.n1787 gnd.n968 9.3005
R9758 gnd.n1789 gnd.n1788 9.3005
R9759 gnd.n1790 gnd.n950 9.3005
R9760 gnd.n1809 gnd.n1808 9.3005
R9761 gnd.n1811 gnd.n943 9.3005
R9762 gnd.n1818 gnd.n944 9.3005
R9763 gnd.n1820 gnd.n1819 9.3005
R9764 gnd.n1821 gnd.n924 9.3005
R9765 gnd.n1840 gnd.n1839 9.3005
R9766 gnd.n1842 gnd.n917 9.3005
R9767 gnd.n1849 gnd.n918 9.3005
R9768 gnd.n1851 gnd.n1850 9.3005
R9769 gnd.n1852 gnd.n899 9.3005
R9770 gnd.n1872 gnd.n1871 9.3005
R9771 gnd.n1874 gnd.n890 9.3005
R9772 gnd.n2137 gnd.n892 9.3005
R9773 gnd.n2138 gnd.n888 9.3005
R9774 gnd.n2141 gnd.n2140 9.3005
R9775 gnd.n782 gnd.n780 9.3005
R9776 gnd.n5987 gnd.n5986 9.3005
R9777 gnd.n1560 gnd.n1559 9.3005
R9778 gnd.n822 gnd.n819 9.3005
R9779 gnd.n824 gnd.n823 9.3005
R9780 gnd.n827 gnd.n817 9.3005
R9781 gnd.n831 gnd.n830 9.3005
R9782 gnd.n832 gnd.n816 9.3005
R9783 gnd.n834 gnd.n833 9.3005
R9784 gnd.n837 gnd.n815 9.3005
R9785 gnd.n841 gnd.n840 9.3005
R9786 gnd.n842 gnd.n814 9.3005
R9787 gnd.n844 gnd.n843 9.3005
R9788 gnd.n847 gnd.n813 9.3005
R9789 gnd.n851 gnd.n850 9.3005
R9790 gnd.n852 gnd.n812 9.3005
R9791 gnd.n854 gnd.n853 9.3005
R9792 gnd.n857 gnd.n811 9.3005
R9793 gnd.n861 gnd.n860 9.3005
R9794 gnd.n862 gnd.n810 9.3005
R9795 gnd.n864 gnd.n863 9.3005
R9796 gnd.n867 gnd.n809 9.3005
R9797 gnd.n871 gnd.n870 9.3005
R9798 gnd.n872 gnd.n808 9.3005
R9799 gnd.n874 gnd.n873 9.3005
R9800 gnd.n877 gnd.n804 9.3005
R9801 gnd.n880 gnd.n879 9.3005
R9802 gnd.n881 gnd.n803 9.3005
R9803 gnd.n2152 gnd.n2151 9.3005
R9804 gnd.n821 gnd.n820 9.3005
R9805 gnd.n1118 gnd.n1049 9.3005
R9806 gnd.n1116 gnd.n1050 9.3005
R9807 gnd.n1115 gnd.n1051 9.3005
R9808 gnd.n1112 gnd.n1052 9.3005
R9809 gnd.n1111 gnd.n1053 9.3005
R9810 gnd.n1110 gnd.n1054 9.3005
R9811 gnd.n1108 gnd.n1055 9.3005
R9812 gnd.n1107 gnd.n1056 9.3005
R9813 gnd.n1104 gnd.n1057 9.3005
R9814 gnd.n1103 gnd.n1058 9.3005
R9815 gnd.n1102 gnd.n1059 9.3005
R9816 gnd.n1100 gnd.n1060 9.3005
R9817 gnd.n1099 gnd.n1061 9.3005
R9818 gnd.n1094 gnd.n1062 9.3005
R9819 gnd.n1093 gnd.n1063 9.3005
R9820 gnd.n1092 gnd.n1064 9.3005
R9821 gnd.n1090 gnd.n1065 9.3005
R9822 gnd.n1089 gnd.n1066 9.3005
R9823 gnd.n1086 gnd.n1067 9.3005
R9824 gnd.n1085 gnd.n1068 9.3005
R9825 gnd.n1084 gnd.n1069 9.3005
R9826 gnd.n1082 gnd.n1070 9.3005
R9827 gnd.n1081 gnd.n1071 9.3005
R9828 gnd.n1078 gnd.n1072 9.3005
R9829 gnd.n1077 gnd.n1073 9.3005
R9830 gnd.n1076 gnd.n1075 9.3005
R9831 gnd.n1074 gnd.n883 9.3005
R9832 gnd.n2148 gnd.n882 9.3005
R9833 gnd.n2150 gnd.n2149 9.3005
R9834 gnd.n1470 gnd.n1469 9.3005
R9835 gnd.n1360 gnd.n1359 9.3005
R9836 gnd.n1484 gnd.n1483 9.3005
R9837 gnd.n1485 gnd.n1358 9.3005
R9838 gnd.n1487 gnd.n1486 9.3005
R9839 gnd.n1348 gnd.n1347 9.3005
R9840 gnd.n1500 gnd.n1499 9.3005
R9841 gnd.n1501 gnd.n1346 9.3005
R9842 gnd.n1533 gnd.n1502 9.3005
R9843 gnd.n1532 gnd.n1503 9.3005
R9844 gnd.n1531 gnd.n1504 9.3005
R9845 gnd.n1530 gnd.n1505 9.3005
R9846 gnd.n1527 gnd.n1506 9.3005
R9847 gnd.n1526 gnd.n1507 9.3005
R9848 gnd.n1525 gnd.n1508 9.3005
R9849 gnd.n1523 gnd.n1509 9.3005
R9850 gnd.n1522 gnd.n1510 9.3005
R9851 gnd.n1519 gnd.n1511 9.3005
R9852 gnd.n1518 gnd.n1512 9.3005
R9853 gnd.n1517 gnd.n1513 9.3005
R9854 gnd.n1515 gnd.n1514 9.3005
R9855 gnd.n1213 gnd.n1212 9.3005
R9856 gnd.n1637 gnd.n1636 9.3005
R9857 gnd.n1638 gnd.n1211 9.3005
R9858 gnd.n1642 gnd.n1639 9.3005
R9859 gnd.n1641 gnd.n1640 9.3005
R9860 gnd.n1176 gnd.n1175 9.3005
R9861 gnd.n1685 gnd.n1684 9.3005
R9862 gnd.n1468 gnd.n1369 9.3005
R9863 gnd.n1371 gnd.n1370 9.3005
R9864 gnd.n1415 gnd.n1413 9.3005
R9865 gnd.n1416 gnd.n1412 9.3005
R9866 gnd.n1419 gnd.n1408 9.3005
R9867 gnd.n1420 gnd.n1407 9.3005
R9868 gnd.n1423 gnd.n1406 9.3005
R9869 gnd.n1424 gnd.n1405 9.3005
R9870 gnd.n1427 gnd.n1404 9.3005
R9871 gnd.n1428 gnd.n1403 9.3005
R9872 gnd.n1431 gnd.n1402 9.3005
R9873 gnd.n1432 gnd.n1401 9.3005
R9874 gnd.n1435 gnd.n1400 9.3005
R9875 gnd.n1436 gnd.n1399 9.3005
R9876 gnd.n1439 gnd.n1398 9.3005
R9877 gnd.n1440 gnd.n1397 9.3005
R9878 gnd.n1443 gnd.n1396 9.3005
R9879 gnd.n1444 gnd.n1395 9.3005
R9880 gnd.n1447 gnd.n1394 9.3005
R9881 gnd.n1448 gnd.n1393 9.3005
R9882 gnd.n1451 gnd.n1392 9.3005
R9883 gnd.n1452 gnd.n1391 9.3005
R9884 gnd.n1455 gnd.n1390 9.3005
R9885 gnd.n1457 gnd.n1389 9.3005
R9886 gnd.n1458 gnd.n1388 9.3005
R9887 gnd.n1459 gnd.n1387 9.3005
R9888 gnd.n1460 gnd.n1386 9.3005
R9889 gnd.n1467 gnd.n1466 9.3005
R9890 gnd.n1476 gnd.n1475 9.3005
R9891 gnd.n1477 gnd.n1363 9.3005
R9892 gnd.n1479 gnd.n1478 9.3005
R9893 gnd.n1354 gnd.n1353 9.3005
R9894 gnd.n1492 gnd.n1491 9.3005
R9895 gnd.n1493 gnd.n1352 9.3005
R9896 gnd.n1495 gnd.n1494 9.3005
R9897 gnd.n1341 gnd.n1340 9.3005
R9898 gnd.n1538 gnd.n1537 9.3005
R9899 gnd.n1539 gnd.n1295 9.3005
R9900 gnd.n1543 gnd.n1541 9.3005
R9901 gnd.n1542 gnd.n1274 9.3005
R9902 gnd.n1561 gnd.n1273 9.3005
R9903 gnd.n1564 gnd.n1563 9.3005
R9904 gnd.n1267 gnd.n1266 9.3005
R9905 gnd.n1575 gnd.n1573 9.3005
R9906 gnd.n1574 gnd.n1248 9.3005
R9907 gnd.n1592 gnd.n1247 9.3005
R9908 gnd.n1595 gnd.n1594 9.3005
R9909 gnd.n1242 gnd.n1237 9.3005
R9910 gnd.n1605 gnd.n1604 9.3005
R9911 gnd.n1240 gnd.n1218 9.3005
R9912 gnd.n1632 gnd.n1219 9.3005
R9913 gnd.n1631 gnd.n1630 9.3005
R9914 gnd.n1221 gnd.n1206 9.3005
R9915 gnd.n1649 gnd.n1648 9.3005
R9916 gnd.n1651 gnd.n1184 9.3005
R9917 gnd.n1680 gnd.n1185 9.3005
R9918 gnd.n1679 gnd.n1186 9.3005
R9919 gnd.n1678 gnd.n1187 9.3005
R9920 gnd.n1190 gnd.n1189 9.3005
R9921 gnd.n1041 gnd.n1040 9.3005
R9922 gnd.n1700 gnd.n1698 9.3005
R9923 gnd.n1699 gnd.n1025 9.3005
R9924 gnd.n1717 gnd.n1024 9.3005
R9925 gnd.n1720 gnd.n1719 9.3005
R9926 gnd.n1018 gnd.n1017 9.3005
R9927 gnd.n1731 gnd.n1729 9.3005
R9928 gnd.n1730 gnd.n1000 9.3005
R9929 gnd.n1748 gnd.n999 9.3005
R9930 gnd.n1751 gnd.n1750 9.3005
R9931 gnd.n992 gnd.n991 9.3005
R9932 gnd.n1762 gnd.n1760 9.3005
R9933 gnd.n1761 gnd.n973 9.3005
R9934 gnd.n1779 gnd.n972 9.3005
R9935 gnd.n1782 gnd.n1781 9.3005
R9936 gnd.n966 gnd.n965 9.3005
R9937 gnd.n1793 gnd.n1791 9.3005
R9938 gnd.n1792 gnd.n949 9.3005
R9939 gnd.n1810 gnd.n948 9.3005
R9940 gnd.n1813 gnd.n1812 9.3005
R9941 gnd.n942 gnd.n941 9.3005
R9942 gnd.n1824 gnd.n1822 9.3005
R9943 gnd.n1823 gnd.n923 9.3005
R9944 gnd.n1841 gnd.n922 9.3005
R9945 gnd.n1844 gnd.n1843 9.3005
R9946 gnd.n916 gnd.n915 9.3005
R9947 gnd.n1855 gnd.n1853 9.3005
R9948 gnd.n1854 gnd.n898 9.3005
R9949 gnd.n1873 gnd.n897 9.3005
R9950 gnd.n2132 gnd.n2131 9.3005
R9951 gnd.n891 gnd.n887 9.3005
R9952 gnd.n2143 gnd.n2142 9.3005
R9953 gnd.n889 gnd.n779 9.3005
R9954 gnd.n5989 gnd.n5988 9.3005
R9955 gnd.n1365 gnd.n1364 9.3005
R9956 gnd.n3770 gnd.n3659 9.3005
R9957 gnd.n3730 gnd.n3670 9.3005
R9958 gnd.n3733 gnd.n3731 9.3005
R9959 gnd.n3734 gnd.n3669 9.3005
R9960 gnd.n3737 gnd.n3736 9.3005
R9961 gnd.n3738 gnd.n3668 9.3005
R9962 gnd.n3741 gnd.n3739 9.3005
R9963 gnd.n3742 gnd.n3667 9.3005
R9964 gnd.n3745 gnd.n3744 9.3005
R9965 gnd.n3746 gnd.n3666 9.3005
R9966 gnd.n3749 gnd.n3747 9.3005
R9967 gnd.n3750 gnd.n3665 9.3005
R9968 gnd.n3753 gnd.n3752 9.3005
R9969 gnd.n3754 gnd.n3664 9.3005
R9970 gnd.n3757 gnd.n3755 9.3005
R9971 gnd.n3758 gnd.n3663 9.3005
R9972 gnd.n3761 gnd.n3760 9.3005
R9973 gnd.n3762 gnd.n3662 9.3005
R9974 gnd.n3765 gnd.n3763 9.3005
R9975 gnd.n3766 gnd.n3661 9.3005
R9976 gnd.n3769 gnd.n3768 9.3005
R9977 gnd.n3729 gnd.n3728 9.3005
R9978 gnd.n5625 gnd.n2540 9.3005
R9979 gnd.n5628 gnd.n2539 9.3005
R9980 gnd.n5629 gnd.n2538 9.3005
R9981 gnd.n5632 gnd.n2537 9.3005
R9982 gnd.n5633 gnd.n2536 9.3005
R9983 gnd.n5636 gnd.n2535 9.3005
R9984 gnd.n5637 gnd.n2534 9.3005
R9985 gnd.n5640 gnd.n2533 9.3005
R9986 gnd.n5642 gnd.n2530 9.3005
R9987 gnd.n5645 gnd.n2529 9.3005
R9988 gnd.n5646 gnd.n2528 9.3005
R9989 gnd.n5649 gnd.n2527 9.3005
R9990 gnd.n5650 gnd.n2526 9.3005
R9991 gnd.n5653 gnd.n2525 9.3005
R9992 gnd.n5654 gnd.n2524 9.3005
R9993 gnd.n5657 gnd.n2523 9.3005
R9994 gnd.n5658 gnd.n2522 9.3005
R9995 gnd.n5661 gnd.n2521 9.3005
R9996 gnd.n5662 gnd.n2520 9.3005
R9997 gnd.n5665 gnd.n2519 9.3005
R9998 gnd.n5666 gnd.n2518 9.3005
R9999 gnd.n5669 gnd.n2517 9.3005
R10000 gnd.n5670 gnd.n2516 9.3005
R10001 gnd.n5671 gnd.n2515 9.3005
R10002 gnd.n2472 gnd.n2471 9.3005
R10003 gnd.n5677 gnd.n5676 9.3005
R10004 gnd.n3543 gnd.n3541 9.3005
R10005 gnd.n3545 gnd.n3544 9.3005
R10006 gnd.n3548 gnd.n3538 9.3005
R10007 gnd.n3552 gnd.n3551 9.3005
R10008 gnd.n3553 gnd.n3537 9.3005
R10009 gnd.n3555 gnd.n3554 9.3005
R10010 gnd.n3558 gnd.n3536 9.3005
R10011 gnd.n3562 gnd.n3561 9.3005
R10012 gnd.n3563 gnd.n3535 9.3005
R10013 gnd.n3565 gnd.n3564 9.3005
R10014 gnd.n3568 gnd.n3532 9.3005
R10015 gnd.n3572 gnd.n3571 9.3005
R10016 gnd.n3573 gnd.n3531 9.3005
R10017 gnd.n3575 gnd.n3574 9.3005
R10018 gnd.n3578 gnd.n3530 9.3005
R10019 gnd.n3582 gnd.n3581 9.3005
R10020 gnd.n3583 gnd.n3529 9.3005
R10021 gnd.n3585 gnd.n3584 9.3005
R10022 gnd.n3588 gnd.n3528 9.3005
R10023 gnd.n3592 gnd.n3591 9.3005
R10024 gnd.n3593 gnd.n3527 9.3005
R10025 gnd.n3595 gnd.n3594 9.3005
R10026 gnd.n3598 gnd.n3526 9.3005
R10027 gnd.n3602 gnd.n3601 9.3005
R10028 gnd.n3603 gnd.n3525 9.3005
R10029 gnd.n3605 gnd.n3604 9.3005
R10030 gnd.n3608 gnd.n3524 9.3005
R10031 gnd.n3612 gnd.n3611 9.3005
R10032 gnd.n3613 gnd.n3523 9.3005
R10033 gnd.n3615 gnd.n3614 9.3005
R10034 gnd.n3542 gnd.n2541 9.3005
R10035 gnd.n5752 gnd.n2349 9.3005
R10036 gnd.n5751 gnd.n2350 9.3005
R10037 gnd.n5750 gnd.n2351 9.3005
R10038 gnd.n2368 gnd.n2352 9.3005
R10039 gnd.n5740 gnd.n2369 9.3005
R10040 gnd.n5739 gnd.n2370 9.3005
R10041 gnd.n5738 gnd.n2371 9.3005
R10042 gnd.n2387 gnd.n2372 9.3005
R10043 gnd.n5728 gnd.n2388 9.3005
R10044 gnd.n5727 gnd.n2389 9.3005
R10045 gnd.n5726 gnd.n2390 9.3005
R10046 gnd.n2407 gnd.n2391 9.3005
R10047 gnd.n5716 gnd.n2408 9.3005
R10048 gnd.n5715 gnd.n2409 9.3005
R10049 gnd.n5714 gnd.n2410 9.3005
R10050 gnd.n2427 gnd.n2411 9.3005
R10051 gnd.n5704 gnd.n2428 9.3005
R10052 gnd.n5703 gnd.n2429 9.3005
R10053 gnd.n5702 gnd.n2430 9.3005
R10054 gnd.n2448 gnd.n2431 9.3005
R10055 gnd.n5692 gnd.n2449 9.3005
R10056 gnd.n5691 gnd.n2450 9.3005
R10057 gnd.n5690 gnd.n2451 9.3005
R10058 gnd.n2469 gnd.n2452 9.3005
R10059 gnd.n5680 gnd.n2470 9.3005
R10060 gnd.n5679 gnd.n5678 9.3005
R10061 gnd.n5802 gnd.n5801 9.3005
R10062 gnd.n5800 gnd.n2273 9.3005
R10063 gnd.n5799 gnd.n5798 9.3005
R10064 gnd.n2276 gnd.n2275 9.3005
R10065 gnd.n5788 gnd.n2293 9.3005
R10066 gnd.n5787 gnd.n2294 9.3005
R10067 gnd.n5786 gnd.n2295 9.3005
R10068 gnd.n2310 gnd.n2296 9.3005
R10069 gnd.n5776 gnd.n2311 9.3005
R10070 gnd.n5775 gnd.n2312 9.3005
R10071 gnd.n5774 gnd.n2313 9.3005
R10072 gnd.n2330 gnd.n2314 9.3005
R10073 gnd.n5764 gnd.n2331 9.3005
R10074 gnd.n5763 gnd.n2332 9.3005
R10075 gnd.n5762 gnd.n2333 9.3005
R10076 gnd.n2348 gnd.n2334 9.3005
R10077 gnd.n2274 gnd.n2272 9.3005
R10078 gnd.n5812 gnd.n5811 9.3005
R10079 gnd.n5815 gnd.n2257 9.3005
R10080 gnd.n5816 gnd.n2256 9.3005
R10081 gnd.n5819 gnd.n2255 9.3005
R10082 gnd.n5820 gnd.n2254 9.3005
R10083 gnd.n5823 gnd.n2253 9.3005
R10084 gnd.n5824 gnd.n2252 9.3005
R10085 gnd.n5827 gnd.n2251 9.3005
R10086 gnd.n5828 gnd.n2250 9.3005
R10087 gnd.n5831 gnd.n2249 9.3005
R10088 gnd.n5832 gnd.n2248 9.3005
R10089 gnd.n5835 gnd.n2247 9.3005
R10090 gnd.n5836 gnd.n2246 9.3005
R10091 gnd.n5839 gnd.n2245 9.3005
R10092 gnd.n5840 gnd.n2244 9.3005
R10093 gnd.n5843 gnd.n2243 9.3005
R10094 gnd.n5844 gnd.n2242 9.3005
R10095 gnd.n5847 gnd.n2241 9.3005
R10096 gnd.n5848 gnd.n2240 9.3005
R10097 gnd.n5851 gnd.n2239 9.3005
R10098 gnd.n5855 gnd.n2235 9.3005
R10099 gnd.n5856 gnd.n2234 9.3005
R10100 gnd.n5859 gnd.n2233 9.3005
R10101 gnd.n5860 gnd.n2232 9.3005
R10102 gnd.n5863 gnd.n2231 9.3005
R10103 gnd.n5864 gnd.n2230 9.3005
R10104 gnd.n5867 gnd.n2229 9.3005
R10105 gnd.n5868 gnd.n2228 9.3005
R10106 gnd.n5871 gnd.n2227 9.3005
R10107 gnd.n5872 gnd.n2226 9.3005
R10108 gnd.n5875 gnd.n2225 9.3005
R10109 gnd.n5876 gnd.n2224 9.3005
R10110 gnd.n5879 gnd.n2223 9.3005
R10111 gnd.n5880 gnd.n2222 9.3005
R10112 gnd.n5883 gnd.n2221 9.3005
R10113 gnd.n5884 gnd.n2220 9.3005
R10114 gnd.n5887 gnd.n2219 9.3005
R10115 gnd.n5888 gnd.n2218 9.3005
R10116 gnd.n5891 gnd.n2217 9.3005
R10117 gnd.n5893 gnd.n2214 9.3005
R10118 gnd.n5896 gnd.n2213 9.3005
R10119 gnd.n5897 gnd.n2212 9.3005
R10120 gnd.n5900 gnd.n2211 9.3005
R10121 gnd.n5901 gnd.n2210 9.3005
R10122 gnd.n5904 gnd.n2209 9.3005
R10123 gnd.n5905 gnd.n2208 9.3005
R10124 gnd.n5908 gnd.n2207 9.3005
R10125 gnd.n5909 gnd.n2206 9.3005
R10126 gnd.n5912 gnd.n2205 9.3005
R10127 gnd.n5913 gnd.n2204 9.3005
R10128 gnd.n5916 gnd.n2203 9.3005
R10129 gnd.n5917 gnd.n2202 9.3005
R10130 gnd.n5920 gnd.n2201 9.3005
R10131 gnd.n5922 gnd.n2200 9.3005
R10132 gnd.n5923 gnd.n2199 9.3005
R10133 gnd.n5924 gnd.n2198 9.3005
R10134 gnd.n5925 gnd.n2197 9.3005
R10135 gnd.n5852 gnd.n2236 9.3005
R10136 gnd.n5810 gnd.n2258 9.3005
R10137 gnd.n3723 gnd.n3722 9.3005
R10138 gnd.n3721 gnd.n3675 9.3005
R10139 gnd.n3720 gnd.n3719 9.3005
R10140 gnd.n3716 gnd.n3678 9.3005
R10141 gnd.n3715 gnd.n3712 9.3005
R10142 gnd.n3711 gnd.n3679 9.3005
R10143 gnd.n3710 gnd.n3709 9.3005
R10144 gnd.n3706 gnd.n3680 9.3005
R10145 gnd.n3705 gnd.n3702 9.3005
R10146 gnd.n3701 gnd.n3681 9.3005
R10147 gnd.n3700 gnd.n3699 9.3005
R10148 gnd.n3696 gnd.n3682 9.3005
R10149 gnd.n3695 gnd.n3692 9.3005
R10150 gnd.n3691 gnd.n3683 9.3005
R10151 gnd.n3690 gnd.n3689 9.3005
R10152 gnd.n3686 gnd.n3684 9.3005
R10153 gnd.n3685 gnd.n2261 9.3005
R10154 gnd.n3724 gnd.n3671 9.3005
R10155 gnd.n3726 gnd.n3725 9.3005
R10156 gnd.n3781 gnd.n2263 9.3005
R10157 gnd.n3784 gnd.n3782 9.3005
R10158 gnd.n3785 gnd.n2284 9.3005
R10159 gnd.n3787 gnd.n2285 9.3005
R10160 gnd.n3788 gnd.n2286 9.3005
R10161 gnd.n3791 gnd.n3789 9.3005
R10162 gnd.n3792 gnd.n2302 9.3005
R10163 gnd.n3794 gnd.n2303 9.3005
R10164 gnd.n3795 gnd.n2304 9.3005
R10165 gnd.n3798 gnd.n3796 9.3005
R10166 gnd.n3799 gnd.n2320 9.3005
R10167 gnd.n3801 gnd.n2321 9.3005
R10168 gnd.n3802 gnd.n2322 9.3005
R10169 gnd.n3805 gnd.n3803 9.3005
R10170 gnd.n3806 gnd.n2340 9.3005
R10171 gnd.n3808 gnd.n2341 9.3005
R10172 gnd.n3809 gnd.n2342 9.3005
R10173 gnd.n3812 gnd.n3810 9.3005
R10174 gnd.n3813 gnd.n2358 9.3005
R10175 gnd.n3815 gnd.n2359 9.3005
R10176 gnd.n3816 gnd.n2360 9.3005
R10177 gnd.n3819 gnd.n3817 9.3005
R10178 gnd.n3820 gnd.n2378 9.3005
R10179 gnd.n3822 gnd.n2379 9.3005
R10180 gnd.n3823 gnd.n2380 9.3005
R10181 gnd.n3826 gnd.n3824 9.3005
R10182 gnd.n3827 gnd.n2397 9.3005
R10183 gnd.n3828 gnd.n2398 9.3005
R10184 gnd.n3652 gnd.n2399 9.3005
R10185 gnd.n3840 gnd.n3653 9.3005
R10186 gnd.n3841 gnd.n2418 9.3005
R10187 gnd.n3842 gnd.n2419 9.3005
R10188 gnd.n3843 gnd.n2420 9.3005
R10189 gnd.n3847 gnd.n3844 9.3005
R10190 gnd.n3848 gnd.n2438 9.3005
R10191 gnd.n3851 gnd.n2439 9.3005
R10192 gnd.n3852 gnd.n2440 9.3005
R10193 gnd.n3856 gnd.n3853 9.3005
R10194 gnd.n3857 gnd.n2459 9.3005
R10195 gnd.n3861 gnd.n2460 9.3005
R10196 gnd.n3860 gnd.n2461 9.3005
R10197 gnd.n3859 gnd.n3858 9.3005
R10198 gnd.n5808 gnd.n2262 9.3005
R10199 gnd.n2264 gnd.n2263 9.3005
R10200 gnd.n3782 gnd.n2283 9.3005
R10201 gnd.n5794 gnd.n2284 9.3005
R10202 gnd.n5793 gnd.n2285 9.3005
R10203 gnd.n5792 gnd.n2286 9.3005
R10204 gnd.n3789 gnd.n2287 9.3005
R10205 gnd.n5782 gnd.n2302 9.3005
R10206 gnd.n5781 gnd.n2303 9.3005
R10207 gnd.n5780 gnd.n2304 9.3005
R10208 gnd.n3796 gnd.n2305 9.3005
R10209 gnd.n5770 gnd.n2320 9.3005
R10210 gnd.n5769 gnd.n2321 9.3005
R10211 gnd.n5768 gnd.n2322 9.3005
R10212 gnd.n3803 gnd.n2323 9.3005
R10213 gnd.n5758 gnd.n2340 9.3005
R10214 gnd.n5757 gnd.n2341 9.3005
R10215 gnd.n5756 gnd.n2342 9.3005
R10216 gnd.n3810 gnd.n2343 9.3005
R10217 gnd.n5746 gnd.n2358 9.3005
R10218 gnd.n5745 gnd.n2359 9.3005
R10219 gnd.n5744 gnd.n2360 9.3005
R10220 gnd.n3817 gnd.n2361 9.3005
R10221 gnd.n5734 gnd.n2378 9.3005
R10222 gnd.n5733 gnd.n2379 9.3005
R10223 gnd.n5732 gnd.n2380 9.3005
R10224 gnd.n3824 gnd.n2381 9.3005
R10225 gnd.n5722 gnd.n2397 9.3005
R10226 gnd.n5721 gnd.n2398 9.3005
R10227 gnd.n5720 gnd.n2399 9.3005
R10228 gnd.n3653 gnd.n2400 9.3005
R10229 gnd.n5710 gnd.n2418 9.3005
R10230 gnd.n5709 gnd.n2419 9.3005
R10231 gnd.n5708 gnd.n2420 9.3005
R10232 gnd.n3844 gnd.n2421 9.3005
R10233 gnd.n5698 gnd.n2438 9.3005
R10234 gnd.n5697 gnd.n2439 9.3005
R10235 gnd.n5696 gnd.n2440 9.3005
R10236 gnd.n3853 gnd.n2441 9.3005
R10237 gnd.n5686 gnd.n2459 9.3005
R10238 gnd.n5685 gnd.n2460 9.3005
R10239 gnd.n5684 gnd.n2461 9.3005
R10240 gnd.n3858 gnd.n2462 9.3005
R10241 gnd.n5808 gnd.n5807 9.3005
R10242 gnd.n6171 gnd.n6170 9.3005
R10243 gnd.n6172 gnd.n592 9.3005
R10244 gnd.n6174 gnd.n6173 9.3005
R10245 gnd.n588 gnd.n587 9.3005
R10246 gnd.n6181 gnd.n6180 9.3005
R10247 gnd.n6182 gnd.n586 9.3005
R10248 gnd.n6184 gnd.n6183 9.3005
R10249 gnd.n582 gnd.n581 9.3005
R10250 gnd.n6191 gnd.n6190 9.3005
R10251 gnd.n6192 gnd.n580 9.3005
R10252 gnd.n6194 gnd.n6193 9.3005
R10253 gnd.n576 gnd.n575 9.3005
R10254 gnd.n6201 gnd.n6200 9.3005
R10255 gnd.n6202 gnd.n574 9.3005
R10256 gnd.n6204 gnd.n6203 9.3005
R10257 gnd.n570 gnd.n569 9.3005
R10258 gnd.n6211 gnd.n6210 9.3005
R10259 gnd.n6212 gnd.n568 9.3005
R10260 gnd.n6214 gnd.n6213 9.3005
R10261 gnd.n564 gnd.n563 9.3005
R10262 gnd.n6221 gnd.n6220 9.3005
R10263 gnd.n6222 gnd.n562 9.3005
R10264 gnd.n6224 gnd.n6223 9.3005
R10265 gnd.n558 gnd.n557 9.3005
R10266 gnd.n6231 gnd.n6230 9.3005
R10267 gnd.n6232 gnd.n556 9.3005
R10268 gnd.n6234 gnd.n6233 9.3005
R10269 gnd.n552 gnd.n551 9.3005
R10270 gnd.n6241 gnd.n6240 9.3005
R10271 gnd.n6242 gnd.n550 9.3005
R10272 gnd.n6244 gnd.n6243 9.3005
R10273 gnd.n546 gnd.n545 9.3005
R10274 gnd.n6251 gnd.n6250 9.3005
R10275 gnd.n6252 gnd.n544 9.3005
R10276 gnd.n6254 gnd.n6253 9.3005
R10277 gnd.n540 gnd.n539 9.3005
R10278 gnd.n6261 gnd.n6260 9.3005
R10279 gnd.n6262 gnd.n538 9.3005
R10280 gnd.n6264 gnd.n6263 9.3005
R10281 gnd.n534 gnd.n533 9.3005
R10282 gnd.n6271 gnd.n6270 9.3005
R10283 gnd.n6272 gnd.n532 9.3005
R10284 gnd.n6274 gnd.n6273 9.3005
R10285 gnd.n528 gnd.n527 9.3005
R10286 gnd.n6281 gnd.n6280 9.3005
R10287 gnd.n6282 gnd.n526 9.3005
R10288 gnd.n6284 gnd.n6283 9.3005
R10289 gnd.n522 gnd.n521 9.3005
R10290 gnd.n6291 gnd.n6290 9.3005
R10291 gnd.n6292 gnd.n520 9.3005
R10292 gnd.n6294 gnd.n6293 9.3005
R10293 gnd.n516 gnd.n515 9.3005
R10294 gnd.n6301 gnd.n6300 9.3005
R10295 gnd.n6302 gnd.n514 9.3005
R10296 gnd.n6304 gnd.n6303 9.3005
R10297 gnd.n510 gnd.n509 9.3005
R10298 gnd.n6311 gnd.n6310 9.3005
R10299 gnd.n6312 gnd.n508 9.3005
R10300 gnd.n6314 gnd.n6313 9.3005
R10301 gnd.n504 gnd.n503 9.3005
R10302 gnd.n6321 gnd.n6320 9.3005
R10303 gnd.n6322 gnd.n502 9.3005
R10304 gnd.n6324 gnd.n6323 9.3005
R10305 gnd.n498 gnd.n497 9.3005
R10306 gnd.n6331 gnd.n6330 9.3005
R10307 gnd.n6332 gnd.n496 9.3005
R10308 gnd.n6334 gnd.n6333 9.3005
R10309 gnd.n492 gnd.n491 9.3005
R10310 gnd.n6341 gnd.n6340 9.3005
R10311 gnd.n6342 gnd.n490 9.3005
R10312 gnd.n6344 gnd.n6343 9.3005
R10313 gnd.n486 gnd.n485 9.3005
R10314 gnd.n6351 gnd.n6350 9.3005
R10315 gnd.n6352 gnd.n484 9.3005
R10316 gnd.n6354 gnd.n6353 9.3005
R10317 gnd.n480 gnd.n479 9.3005
R10318 gnd.n6361 gnd.n6360 9.3005
R10319 gnd.n6362 gnd.n478 9.3005
R10320 gnd.n6364 gnd.n6363 9.3005
R10321 gnd.n474 gnd.n473 9.3005
R10322 gnd.n6371 gnd.n6370 9.3005
R10323 gnd.n6372 gnd.n472 9.3005
R10324 gnd.n6374 gnd.n6373 9.3005
R10325 gnd.n468 gnd.n467 9.3005
R10326 gnd.n6381 gnd.n6380 9.3005
R10327 gnd.n6382 gnd.n466 9.3005
R10328 gnd.n6384 gnd.n6383 9.3005
R10329 gnd.n462 gnd.n461 9.3005
R10330 gnd.n6391 gnd.n6390 9.3005
R10331 gnd.n6392 gnd.n460 9.3005
R10332 gnd.n6394 gnd.n6393 9.3005
R10333 gnd.n456 gnd.n455 9.3005
R10334 gnd.n6401 gnd.n6400 9.3005
R10335 gnd.n6402 gnd.n454 9.3005
R10336 gnd.n6404 gnd.n6403 9.3005
R10337 gnd.n450 gnd.n449 9.3005
R10338 gnd.n6411 gnd.n6410 9.3005
R10339 gnd.n6412 gnd.n448 9.3005
R10340 gnd.n6414 gnd.n6413 9.3005
R10341 gnd.n444 gnd.n443 9.3005
R10342 gnd.n6421 gnd.n6420 9.3005
R10343 gnd.n6422 gnd.n442 9.3005
R10344 gnd.n6424 gnd.n6423 9.3005
R10345 gnd.n438 gnd.n437 9.3005
R10346 gnd.n6431 gnd.n6430 9.3005
R10347 gnd.n6432 gnd.n436 9.3005
R10348 gnd.n6434 gnd.n6433 9.3005
R10349 gnd.n432 gnd.n431 9.3005
R10350 gnd.n6441 gnd.n6440 9.3005
R10351 gnd.n6442 gnd.n430 9.3005
R10352 gnd.n6444 gnd.n6443 9.3005
R10353 gnd.n426 gnd.n425 9.3005
R10354 gnd.n6451 gnd.n6450 9.3005
R10355 gnd.n6452 gnd.n424 9.3005
R10356 gnd.n6454 gnd.n6453 9.3005
R10357 gnd.n420 gnd.n419 9.3005
R10358 gnd.n6461 gnd.n6460 9.3005
R10359 gnd.n6462 gnd.n418 9.3005
R10360 gnd.n6464 gnd.n6463 9.3005
R10361 gnd.n414 gnd.n413 9.3005
R10362 gnd.n6471 gnd.n6470 9.3005
R10363 gnd.n6472 gnd.n412 9.3005
R10364 gnd.n6474 gnd.n6473 9.3005
R10365 gnd.n408 gnd.n407 9.3005
R10366 gnd.n6481 gnd.n6480 9.3005
R10367 gnd.n6482 gnd.n406 9.3005
R10368 gnd.n6484 gnd.n6483 9.3005
R10369 gnd.n402 gnd.n401 9.3005
R10370 gnd.n6491 gnd.n6490 9.3005
R10371 gnd.n6492 gnd.n400 9.3005
R10372 gnd.n6494 gnd.n6493 9.3005
R10373 gnd.n396 gnd.n395 9.3005
R10374 gnd.n6501 gnd.n6500 9.3005
R10375 gnd.n6502 gnd.n394 9.3005
R10376 gnd.n6504 gnd.n6503 9.3005
R10377 gnd.n390 gnd.n389 9.3005
R10378 gnd.n6511 gnd.n6510 9.3005
R10379 gnd.n6512 gnd.n388 9.3005
R10380 gnd.n6515 gnd.n6514 9.3005
R10381 gnd.n6513 gnd.n384 9.3005
R10382 gnd.n6521 gnd.n383 9.3005
R10383 gnd.n6523 gnd.n6522 9.3005
R10384 gnd.n379 gnd.n378 9.3005
R10385 gnd.n6532 gnd.n6531 9.3005
R10386 gnd.n6533 gnd.n377 9.3005
R10387 gnd.n6535 gnd.n6534 9.3005
R10388 gnd.n373 gnd.n372 9.3005
R10389 gnd.n6542 gnd.n6541 9.3005
R10390 gnd.n6543 gnd.n371 9.3005
R10391 gnd.n6545 gnd.n6544 9.3005
R10392 gnd.n367 gnd.n366 9.3005
R10393 gnd.n6552 gnd.n6551 9.3005
R10394 gnd.n6553 gnd.n365 9.3005
R10395 gnd.n6555 gnd.n6554 9.3005
R10396 gnd.n361 gnd.n360 9.3005
R10397 gnd.n6562 gnd.n6561 9.3005
R10398 gnd.n6563 gnd.n359 9.3005
R10399 gnd.n6565 gnd.n6564 9.3005
R10400 gnd.n355 gnd.n354 9.3005
R10401 gnd.n6572 gnd.n6571 9.3005
R10402 gnd.n6573 gnd.n353 9.3005
R10403 gnd.n6575 gnd.n6574 9.3005
R10404 gnd.n349 gnd.n348 9.3005
R10405 gnd.n6582 gnd.n6581 9.3005
R10406 gnd.n6583 gnd.n347 9.3005
R10407 gnd.n6585 gnd.n6584 9.3005
R10408 gnd.n343 gnd.n342 9.3005
R10409 gnd.n6592 gnd.n6591 9.3005
R10410 gnd.n6593 gnd.n341 9.3005
R10411 gnd.n6595 gnd.n6594 9.3005
R10412 gnd.n337 gnd.n336 9.3005
R10413 gnd.n6602 gnd.n6601 9.3005
R10414 gnd.n6603 gnd.n335 9.3005
R10415 gnd.n6605 gnd.n6604 9.3005
R10416 gnd.n331 gnd.n330 9.3005
R10417 gnd.n6612 gnd.n6611 9.3005
R10418 gnd.n6613 gnd.n329 9.3005
R10419 gnd.n6615 gnd.n6614 9.3005
R10420 gnd.n325 gnd.n324 9.3005
R10421 gnd.n6622 gnd.n6621 9.3005
R10422 gnd.n6623 gnd.n323 9.3005
R10423 gnd.n6625 gnd.n6624 9.3005
R10424 gnd.n319 gnd.n318 9.3005
R10425 gnd.n6632 gnd.n6631 9.3005
R10426 gnd.n6633 gnd.n317 9.3005
R10427 gnd.n6635 gnd.n6634 9.3005
R10428 gnd.n313 gnd.n312 9.3005
R10429 gnd.n6642 gnd.n6641 9.3005
R10430 gnd.n6643 gnd.n311 9.3005
R10431 gnd.n6645 gnd.n6644 9.3005
R10432 gnd.n307 gnd.n306 9.3005
R10433 gnd.n6652 gnd.n6651 9.3005
R10434 gnd.n6653 gnd.n305 9.3005
R10435 gnd.n6655 gnd.n6654 9.3005
R10436 gnd.n301 gnd.n300 9.3005
R10437 gnd.n6662 gnd.n6661 9.3005
R10438 gnd.n6663 gnd.n299 9.3005
R10439 gnd.n6665 gnd.n6664 9.3005
R10440 gnd.n295 gnd.n294 9.3005
R10441 gnd.n6672 gnd.n6671 9.3005
R10442 gnd.n6673 gnd.n293 9.3005
R10443 gnd.n6675 gnd.n6674 9.3005
R10444 gnd.n289 gnd.n288 9.3005
R10445 gnd.n6682 gnd.n6681 9.3005
R10446 gnd.n6683 gnd.n287 9.3005
R10447 gnd.n6685 gnd.n6684 9.3005
R10448 gnd.n283 gnd.n282 9.3005
R10449 gnd.n6692 gnd.n6691 9.3005
R10450 gnd.n6693 gnd.n281 9.3005
R10451 gnd.n6695 gnd.n6694 9.3005
R10452 gnd.n277 gnd.n276 9.3005
R10453 gnd.n6702 gnd.n6701 9.3005
R10454 gnd.n6703 gnd.n275 9.3005
R10455 gnd.n6705 gnd.n6704 9.3005
R10456 gnd.n271 gnd.n270 9.3005
R10457 gnd.n6712 gnd.n6711 9.3005
R10458 gnd.n6713 gnd.n269 9.3005
R10459 gnd.n6715 gnd.n6714 9.3005
R10460 gnd.n265 gnd.n264 9.3005
R10461 gnd.n6722 gnd.n6721 9.3005
R10462 gnd.n6723 gnd.n263 9.3005
R10463 gnd.n6725 gnd.n6724 9.3005
R10464 gnd.n259 gnd.n258 9.3005
R10465 gnd.n6733 gnd.n6732 9.3005
R10466 gnd.n6734 gnd.n257 9.3005
R10467 gnd.n6736 gnd.n6735 9.3005
R10468 gnd.n6525 gnd.n6524 9.3005
R10469 gnd.n3637 gnd.n3632 9.3005
R10470 gnd.n3639 gnd.n3638 9.3005
R10471 gnd.n3630 gnd.n3629 9.3005
R10472 gnd.n3887 gnd.n3886 9.3005
R10473 gnd.n3888 gnd.n3628 9.3005
R10474 gnd.n3890 gnd.n3889 9.3005
R10475 gnd.n3626 gnd.n3625 9.3005
R10476 gnd.n3895 gnd.n3894 9.3005
R10477 gnd.n3896 gnd.n3624 9.3005
R10478 gnd.n3898 gnd.n3897 9.3005
R10479 gnd.n3622 gnd.n3621 9.3005
R10480 gnd.n3903 gnd.n3902 9.3005
R10481 gnd.n3904 gnd.n3620 9.3005
R10482 gnd.n3921 gnd.n3905 9.3005
R10483 gnd.n3920 gnd.n3906 9.3005
R10484 gnd.n3919 gnd.n3907 9.3005
R10485 gnd.n3910 gnd.n3908 9.3005
R10486 gnd.n3914 gnd.n3911 9.3005
R10487 gnd.n3913 gnd.n3912 9.3005
R10488 gnd.n3389 gnd.n3388 9.3005
R10489 gnd.n4001 gnd.n4000 9.3005
R10490 gnd.n4002 gnd.n3387 9.3005
R10491 gnd.n4004 gnd.n4003 9.3005
R10492 gnd.n3374 gnd.n3373 9.3005
R10493 gnd.n4017 gnd.n4016 9.3005
R10494 gnd.n4018 gnd.n3372 9.3005
R10495 gnd.n4020 gnd.n4019 9.3005
R10496 gnd.n3359 gnd.n3358 9.3005
R10497 gnd.n4045 gnd.n4044 9.3005
R10498 gnd.n4046 gnd.n3357 9.3005
R10499 gnd.n4051 gnd.n4047 9.3005
R10500 gnd.n4050 gnd.n4049 9.3005
R10501 gnd.n4048 gnd.n2611 9.3005
R10502 gnd.n5547 gnd.n2612 9.3005
R10503 gnd.n5546 gnd.n2613 9.3005
R10504 gnd.n5545 gnd.n2614 9.3005
R10505 gnd.n3334 gnd.n2615 9.3005
R10506 gnd.n3336 gnd.n3335 9.3005
R10507 gnd.n3318 gnd.n3317 9.3005
R10508 gnd.n4194 gnd.n4193 9.3005
R10509 gnd.n4195 gnd.n3316 9.3005
R10510 gnd.n4202 gnd.n4196 9.3005
R10511 gnd.n4201 gnd.n4197 9.3005
R10512 gnd.n4200 gnd.n4198 9.3005
R10513 gnd.n3288 gnd.n3287 9.3005
R10514 gnd.n4263 gnd.n4262 9.3005
R10515 gnd.n4264 gnd.n3286 9.3005
R10516 gnd.n4266 gnd.n4265 9.3005
R10517 gnd.n3271 gnd.n3270 9.3005
R10518 gnd.n4292 gnd.n4291 9.3005
R10519 gnd.n4293 gnd.n3269 9.3005
R10520 gnd.n4297 gnd.n4294 9.3005
R10521 gnd.n4296 gnd.n4295 9.3005
R10522 gnd.n3243 gnd.n3242 9.3005
R10523 gnd.n4366 gnd.n4365 9.3005
R10524 gnd.n4367 gnd.n3241 9.3005
R10525 gnd.n4371 gnd.n4368 9.3005
R10526 gnd.n4370 gnd.n4369 9.3005
R10527 gnd.n3220 gnd.n3219 9.3005
R10528 gnd.n4398 gnd.n4397 9.3005
R10529 gnd.n4399 gnd.n3218 9.3005
R10530 gnd.n4403 gnd.n4400 9.3005
R10531 gnd.n4402 gnd.n4401 9.3005
R10532 gnd.n3199 gnd.n3198 9.3005
R10533 gnd.n4439 gnd.n4438 9.3005
R10534 gnd.n4440 gnd.n3197 9.3005
R10535 gnd.n4444 gnd.n4441 9.3005
R10536 gnd.n4443 gnd.n4442 9.3005
R10537 gnd.n3170 gnd.n3169 9.3005
R10538 gnd.n4508 gnd.n4507 9.3005
R10539 gnd.n4509 gnd.n3168 9.3005
R10540 gnd.n4513 gnd.n4510 9.3005
R10541 gnd.n4512 gnd.n4511 9.3005
R10542 gnd.n3145 gnd.n3144 9.3005
R10543 gnd.n4540 gnd.n4539 9.3005
R10544 gnd.n4541 gnd.n3143 9.3005
R10545 gnd.n4545 gnd.n4542 9.3005
R10546 gnd.n4544 gnd.n4543 9.3005
R10547 gnd.n3122 gnd.n3121 9.3005
R10548 gnd.n4580 gnd.n4579 9.3005
R10549 gnd.n4581 gnd.n3120 9.3005
R10550 gnd.n4585 gnd.n4582 9.3005
R10551 gnd.n4584 gnd.n4583 9.3005
R10552 gnd.n3093 gnd.n3092 9.3005
R10553 gnd.n4634 gnd.n4633 9.3005
R10554 gnd.n4635 gnd.n3091 9.3005
R10555 gnd.n4639 gnd.n4636 9.3005
R10556 gnd.n4638 gnd.n4637 9.3005
R10557 gnd.n3069 gnd.n3068 9.3005
R10558 gnd.n4676 gnd.n4675 9.3005
R10559 gnd.n4677 gnd.n3067 9.3005
R10560 gnd.n4681 gnd.n4678 9.3005
R10561 gnd.n4680 gnd.n4679 9.3005
R10562 gnd.n3041 gnd.n3040 9.3005
R10563 gnd.n4719 gnd.n4718 9.3005
R10564 gnd.n4720 gnd.n3039 9.3005
R10565 gnd.n4723 gnd.n4722 9.3005
R10566 gnd.n4721 gnd.n3018 9.3005
R10567 gnd.n4763 gnd.n3019 9.3005
R10568 gnd.n4762 gnd.n3020 9.3005
R10569 gnd.n4761 gnd.n3021 9.3005
R10570 gnd.n3023 gnd.n3022 9.3005
R10571 gnd.n3025 gnd.n3024 9.3005
R10572 gnd.n2987 gnd.n2986 9.3005
R10573 gnd.n4811 gnd.n4810 9.3005
R10574 gnd.n4812 gnd.n2985 9.3005
R10575 gnd.n4814 gnd.n4813 9.3005
R10576 gnd.n2935 gnd.n2934 9.3005
R10577 gnd.n4983 gnd.n4982 9.3005
R10578 gnd.n4984 gnd.n2933 9.3005
R10579 gnd.n4986 gnd.n4985 9.3005
R10580 gnd.n2923 gnd.n2922 9.3005
R10581 gnd.n5001 gnd.n5000 9.3005
R10582 gnd.n5002 gnd.n2921 9.3005
R10583 gnd.n5004 gnd.n5003 9.3005
R10584 gnd.n2912 gnd.n2911 9.3005
R10585 gnd.n5018 gnd.n5017 9.3005
R10586 gnd.n5019 gnd.n2910 9.3005
R10587 gnd.n5023 gnd.n5020 9.3005
R10588 gnd.n5022 gnd.n5021 9.3005
R10589 gnd.n2899 gnd.n2898 9.3005
R10590 gnd.n5055 gnd.n5054 9.3005
R10591 gnd.n5056 gnd.n2897 9.3005
R10592 gnd.n5058 gnd.n5057 9.3005
R10593 gnd.n2895 gnd.n2894 9.3005
R10594 gnd.n5064 gnd.n5063 9.3005
R10595 gnd.n5065 gnd.n2893 9.3005
R10596 gnd.n5189 gnd.n5066 9.3005
R10597 gnd.n5188 gnd.n5067 9.3005
R10598 gnd.n5187 gnd.n5068 9.3005
R10599 gnd.n5110 gnd.n5069 9.3005
R10600 gnd.n5113 gnd.n5112 9.3005
R10601 gnd.n5114 gnd.n5109 9.3005
R10602 gnd.n5125 gnd.n5115 9.3005
R10603 gnd.n5124 gnd.n5116 9.3005
R10604 gnd.n5123 gnd.n5117 9.3005
R10605 gnd.n5120 gnd.n5119 9.3005
R10606 gnd.n5118 gnd.n252 9.3005
R10607 gnd.n6741 gnd.n253 9.3005
R10608 gnd.n6740 gnd.n254 9.3005
R10609 gnd.n6739 gnd.n255 9.3005
R10610 gnd.n3636 gnd.n3635 9.3005
R10611 gnd.n6002 gnd.n760 9.3005
R10612 gnd.n6003 gnd.n759 9.3005
R10613 gnd.n6004 gnd.n758 9.3005
R10614 gnd.n757 gnd.n753 9.3005
R10615 gnd.n6010 gnd.n752 9.3005
R10616 gnd.n6011 gnd.n751 9.3005
R10617 gnd.n6012 gnd.n750 9.3005
R10618 gnd.n749 gnd.n745 9.3005
R10619 gnd.n6018 gnd.n744 9.3005
R10620 gnd.n6019 gnd.n743 9.3005
R10621 gnd.n6020 gnd.n742 9.3005
R10622 gnd.n741 gnd.n737 9.3005
R10623 gnd.n6026 gnd.n736 9.3005
R10624 gnd.n6027 gnd.n735 9.3005
R10625 gnd.n6028 gnd.n734 9.3005
R10626 gnd.n733 gnd.n729 9.3005
R10627 gnd.n6034 gnd.n728 9.3005
R10628 gnd.n6035 gnd.n727 9.3005
R10629 gnd.n6036 gnd.n726 9.3005
R10630 gnd.n725 gnd.n721 9.3005
R10631 gnd.n6042 gnd.n720 9.3005
R10632 gnd.n6043 gnd.n719 9.3005
R10633 gnd.n6044 gnd.n718 9.3005
R10634 gnd.n717 gnd.n713 9.3005
R10635 gnd.n6050 gnd.n712 9.3005
R10636 gnd.n6051 gnd.n711 9.3005
R10637 gnd.n6052 gnd.n710 9.3005
R10638 gnd.n709 gnd.n705 9.3005
R10639 gnd.n6058 gnd.n704 9.3005
R10640 gnd.n6059 gnd.n703 9.3005
R10641 gnd.n6060 gnd.n702 9.3005
R10642 gnd.n701 gnd.n697 9.3005
R10643 gnd.n6066 gnd.n696 9.3005
R10644 gnd.n6067 gnd.n695 9.3005
R10645 gnd.n6068 gnd.n694 9.3005
R10646 gnd.n693 gnd.n689 9.3005
R10647 gnd.n6074 gnd.n688 9.3005
R10648 gnd.n6075 gnd.n687 9.3005
R10649 gnd.n6076 gnd.n686 9.3005
R10650 gnd.n685 gnd.n681 9.3005
R10651 gnd.n6082 gnd.n680 9.3005
R10652 gnd.n6083 gnd.n679 9.3005
R10653 gnd.n6084 gnd.n678 9.3005
R10654 gnd.n677 gnd.n673 9.3005
R10655 gnd.n6090 gnd.n672 9.3005
R10656 gnd.n6091 gnd.n671 9.3005
R10657 gnd.n6092 gnd.n670 9.3005
R10658 gnd.n669 gnd.n665 9.3005
R10659 gnd.n6098 gnd.n664 9.3005
R10660 gnd.n6099 gnd.n663 9.3005
R10661 gnd.n6100 gnd.n662 9.3005
R10662 gnd.n661 gnd.n657 9.3005
R10663 gnd.n6106 gnd.n656 9.3005
R10664 gnd.n6107 gnd.n655 9.3005
R10665 gnd.n6108 gnd.n654 9.3005
R10666 gnd.n653 gnd.n649 9.3005
R10667 gnd.n6114 gnd.n648 9.3005
R10668 gnd.n6115 gnd.n647 9.3005
R10669 gnd.n6116 gnd.n646 9.3005
R10670 gnd.n645 gnd.n641 9.3005
R10671 gnd.n6122 gnd.n640 9.3005
R10672 gnd.n6123 gnd.n639 9.3005
R10673 gnd.n6124 gnd.n638 9.3005
R10674 gnd.n637 gnd.n633 9.3005
R10675 gnd.n6130 gnd.n632 9.3005
R10676 gnd.n6131 gnd.n631 9.3005
R10677 gnd.n6132 gnd.n630 9.3005
R10678 gnd.n629 gnd.n625 9.3005
R10679 gnd.n6138 gnd.n624 9.3005
R10680 gnd.n6139 gnd.n623 9.3005
R10681 gnd.n6140 gnd.n622 9.3005
R10682 gnd.n621 gnd.n617 9.3005
R10683 gnd.n6146 gnd.n616 9.3005
R10684 gnd.n6147 gnd.n615 9.3005
R10685 gnd.n6148 gnd.n614 9.3005
R10686 gnd.n613 gnd.n609 9.3005
R10687 gnd.n6154 gnd.n608 9.3005
R10688 gnd.n6155 gnd.n607 9.3005
R10689 gnd.n6156 gnd.n606 9.3005
R10690 gnd.n605 gnd.n601 9.3005
R10691 gnd.n6162 gnd.n600 9.3005
R10692 gnd.n6163 gnd.n599 9.3005
R10693 gnd.n6164 gnd.n598 9.3005
R10694 gnd.n597 gnd.n593 9.3005
R10695 gnd.n3633 gnd.n761 9.3005
R10696 gnd.n5412 gnd.n5411 9.3005
R10697 gnd.n3996 gnd.n3995 9.3005
R10698 gnd.n3382 gnd.n3381 9.3005
R10699 gnd.n4009 gnd.n4008 9.3005
R10700 gnd.n4010 gnd.n3380 9.3005
R10701 gnd.n4012 gnd.n4011 9.3005
R10702 gnd.n3368 gnd.n3367 9.3005
R10703 gnd.n4025 gnd.n4024 9.3005
R10704 gnd.n4026 gnd.n3365 9.3005
R10705 gnd.n4040 gnd.n4039 9.3005
R10706 gnd.n4038 gnd.n3366 9.3005
R10707 gnd.n4037 gnd.n4036 9.3005
R10708 gnd.n4035 gnd.n4027 9.3005
R10709 gnd.n4034 gnd.n4033 9.3005
R10710 gnd.n4032 gnd.n4031 9.3005
R10711 gnd.n2622 gnd.n2620 9.3005
R10712 gnd.n5541 gnd.n5540 9.3005
R10713 gnd.n5539 gnd.n2621 9.3005
R10714 gnd.n5538 gnd.n5537 9.3005
R10715 gnd.n5536 gnd.n2623 9.3005
R10716 gnd.n5535 gnd.n5534 9.3005
R10717 gnd.n5533 gnd.n2627 9.3005
R10718 gnd.n5532 gnd.n5531 9.3005
R10719 gnd.n5530 gnd.n2628 9.3005
R10720 gnd.n5529 gnd.n5528 9.3005
R10721 gnd.n5527 gnd.n2632 9.3005
R10722 gnd.n5526 gnd.n5525 9.3005
R10723 gnd.n5524 gnd.n2633 9.3005
R10724 gnd.n5523 gnd.n5522 9.3005
R10725 gnd.n5521 gnd.n2637 9.3005
R10726 gnd.n5520 gnd.n5519 9.3005
R10727 gnd.n5518 gnd.n2638 9.3005
R10728 gnd.n5517 gnd.n5516 9.3005
R10729 gnd.n5515 gnd.n2642 9.3005
R10730 gnd.n5514 gnd.n5513 9.3005
R10731 gnd.n5512 gnd.n2643 9.3005
R10732 gnd.n5511 gnd.n5510 9.3005
R10733 gnd.n5509 gnd.n2647 9.3005
R10734 gnd.n5508 gnd.n5507 9.3005
R10735 gnd.n5506 gnd.n2648 9.3005
R10736 gnd.n5505 gnd.n5504 9.3005
R10737 gnd.n5503 gnd.n2652 9.3005
R10738 gnd.n5502 gnd.n5501 9.3005
R10739 gnd.n5500 gnd.n2653 9.3005
R10740 gnd.n5499 gnd.n5498 9.3005
R10741 gnd.n5497 gnd.n2657 9.3005
R10742 gnd.n5496 gnd.n5495 9.3005
R10743 gnd.n5494 gnd.n2658 9.3005
R10744 gnd.n5493 gnd.n5492 9.3005
R10745 gnd.n5491 gnd.n2662 9.3005
R10746 gnd.n5490 gnd.n5489 9.3005
R10747 gnd.n5488 gnd.n2663 9.3005
R10748 gnd.n5487 gnd.n5486 9.3005
R10749 gnd.n5485 gnd.n2667 9.3005
R10750 gnd.n5484 gnd.n5483 9.3005
R10751 gnd.n5482 gnd.n2668 9.3005
R10752 gnd.n5481 gnd.n5480 9.3005
R10753 gnd.n5479 gnd.n2672 9.3005
R10754 gnd.n5478 gnd.n5477 9.3005
R10755 gnd.n5476 gnd.n2673 9.3005
R10756 gnd.n5475 gnd.n5474 9.3005
R10757 gnd.n5473 gnd.n2677 9.3005
R10758 gnd.n5472 gnd.n5471 9.3005
R10759 gnd.n5470 gnd.n2678 9.3005
R10760 gnd.n5469 gnd.n5468 9.3005
R10761 gnd.n5467 gnd.n2682 9.3005
R10762 gnd.n5466 gnd.n5465 9.3005
R10763 gnd.n5464 gnd.n2683 9.3005
R10764 gnd.n5463 gnd.n5462 9.3005
R10765 gnd.n5461 gnd.n2687 9.3005
R10766 gnd.n5460 gnd.n5459 9.3005
R10767 gnd.n5458 gnd.n2688 9.3005
R10768 gnd.n5457 gnd.n5456 9.3005
R10769 gnd.n5455 gnd.n2692 9.3005
R10770 gnd.n5454 gnd.n5453 9.3005
R10771 gnd.n5452 gnd.n2693 9.3005
R10772 gnd.n5451 gnd.n5450 9.3005
R10773 gnd.n5449 gnd.n2697 9.3005
R10774 gnd.n5448 gnd.n5447 9.3005
R10775 gnd.n5446 gnd.n2698 9.3005
R10776 gnd.n5445 gnd.n5444 9.3005
R10777 gnd.n5443 gnd.n2702 9.3005
R10778 gnd.n5442 gnd.n5441 9.3005
R10779 gnd.n5440 gnd.n2703 9.3005
R10780 gnd.n5439 gnd.n5438 9.3005
R10781 gnd.n5437 gnd.n2707 9.3005
R10782 gnd.n5436 gnd.n5435 9.3005
R10783 gnd.n5434 gnd.n2708 9.3005
R10784 gnd.n5433 gnd.n5432 9.3005
R10785 gnd.n5431 gnd.n2712 9.3005
R10786 gnd.n5430 gnd.n5429 9.3005
R10787 gnd.n5428 gnd.n2713 9.3005
R10788 gnd.n5427 gnd.n5426 9.3005
R10789 gnd.n5425 gnd.n2717 9.3005
R10790 gnd.n5424 gnd.n5423 9.3005
R10791 gnd.n5422 gnd.n2718 9.3005
R10792 gnd.n5421 gnd.n5420 9.3005
R10793 gnd.n5419 gnd.n2722 9.3005
R10794 gnd.n5418 gnd.n5417 9.3005
R10795 gnd.n5416 gnd.n2723 9.3005
R10796 gnd.n5415 gnd.n5414 9.3005
R10797 gnd.n5413 gnd.n2727 9.3005
R10798 gnd.n3994 gnd.n3394 9.3005
R10799 gnd.n3993 gnd.n3992 9.3005
R10800 gnd.n3772 gnd.n3771 9.3005
R10801 gnd.n3773 gnd.n3658 9.3005
R10802 gnd.n3776 gnd.n3775 9.3005
R10803 gnd.n3777 gnd.n3656 9.3005
R10804 gnd.n3779 gnd.n3778 9.3005
R10805 gnd.n3780 gnd.n3655 9.3005
R10806 gnd.n3833 gnd.n3832 9.3005
R10807 gnd.n3834 gnd.n3654 9.3005
R10808 gnd.n3836 gnd.n3835 9.3005
R10809 gnd.n3645 gnd.n3643 9.3005
R10810 gnd.n3881 gnd.n3880 9.3005
R10811 gnd.n3879 gnd.n3644 9.3005
R10812 gnd.n3878 gnd.n3877 9.3005
R10813 gnd.n3876 gnd.n3646 9.3005
R10814 gnd.n3875 gnd.n3874 9.3005
R10815 gnd.n3873 gnd.n3649 9.3005
R10816 gnd.n3872 gnd.n3871 9.3005
R10817 gnd.n3870 gnd.n3650 9.3005
R10818 gnd.n3869 gnd.n3868 9.3005
R10819 gnd.n3867 gnd.n3865 9.3005
R10820 gnd.n3866 gnd.n3520 9.3005
R10821 gnd.n3970 gnd.n3969 9.3005
R10822 gnd.n3968 gnd.n3967 9.3005
R10823 gnd.n3460 gnd.n3459 9.3005
R10824 gnd.n3962 gnd.n3961 9.3005
R10825 gnd.n3960 gnd.n3959 9.3005
R10826 gnd.n3470 gnd.n3469 9.3005
R10827 gnd.n3954 gnd.n3953 9.3005
R10828 gnd.n3952 gnd.n3951 9.3005
R10829 gnd.n3480 gnd.n3479 9.3005
R10830 gnd.n3946 gnd.n3945 9.3005
R10831 gnd.n3944 gnd.n3943 9.3005
R10832 gnd.n3490 gnd.n3489 9.3005
R10833 gnd.n3938 gnd.n3937 9.3005
R10834 gnd.n3936 gnd.n3935 9.3005
R10835 gnd.n3500 gnd.n3499 9.3005
R10836 gnd.n3930 gnd.n3929 9.3005
R10837 gnd.n3928 gnd.n3511 9.3005
R10838 gnd.n3927 gnd.n3519 9.3005
R10839 gnd.n3455 gnd.n3453 9.3005
R10840 gnd.n3518 gnd.n3396 9.3005
R10841 gnd.n3517 gnd.n3516 9.3005
R10842 gnd.n3514 gnd.n3507 9.3005
R10843 gnd.n3932 gnd.n3931 9.3005
R10844 gnd.n3934 gnd.n3933 9.3005
R10845 gnd.n3494 gnd.n3493 9.3005
R10846 gnd.n3940 gnd.n3939 9.3005
R10847 gnd.n3942 gnd.n3941 9.3005
R10848 gnd.n3486 gnd.n3485 9.3005
R10849 gnd.n3948 gnd.n3947 9.3005
R10850 gnd.n3950 gnd.n3949 9.3005
R10851 gnd.n3474 gnd.n3473 9.3005
R10852 gnd.n3956 gnd.n3955 9.3005
R10853 gnd.n3958 gnd.n3957 9.3005
R10854 gnd.n3466 gnd.n3465 9.3005
R10855 gnd.n3964 gnd.n3963 9.3005
R10856 gnd.n3966 gnd.n3965 9.3005
R10857 gnd.n3454 gnd.n3452 9.3005
R10858 gnd.n3972 gnd.n3971 9.3005
R10859 gnd.n3973 gnd.n3447 9.3005
R10860 gnd.n3975 gnd.n3974 9.3005
R10861 gnd.n3977 gnd.n3445 9.3005
R10862 gnd.n3979 gnd.n3978 9.3005
R10863 gnd.n3980 gnd.n3441 9.3005
R10864 gnd.n3982 gnd.n3981 9.3005
R10865 gnd.n3983 gnd.n3440 9.3005
R10866 gnd.n3985 gnd.n3984 9.3005
R10867 gnd.n3986 gnd.n3439 9.3005
R10868 gnd.n3436 gnd.n3415 9.3005
R10869 gnd.n3435 gnd.n3434 9.3005
R10870 gnd.n3433 gnd.n3417 9.3005
R10871 gnd.n3432 gnd.n3431 9.3005
R10872 gnd.n3430 gnd.n3418 9.3005
R10873 gnd.n3429 gnd.n3428 9.3005
R10874 gnd.n3427 gnd.n3421 9.3005
R10875 gnd.n3426 gnd.n3425 9.3005
R10876 gnd.n3424 gnd.n3422 9.3005
R10877 gnd.n3350 gnd.n3349 9.3005
R10878 gnd.n4056 gnd.n4055 9.3005
R10879 gnd.n4057 gnd.n3347 9.3005
R10880 gnd.n4059 gnd.n4058 9.3005
R10881 gnd.n4060 gnd.n3346 9.3005
R10882 gnd.n4144 gnd.n4143 9.3005
R10883 gnd.n4145 gnd.n3344 9.3005
R10884 gnd.n4161 gnd.n4160 9.3005
R10885 gnd.n4159 gnd.n3345 9.3005
R10886 gnd.n4158 gnd.n4157 9.3005
R10887 gnd.n4156 gnd.n4146 9.3005
R10888 gnd.n4155 gnd.n4154 9.3005
R10889 gnd.n4153 gnd.n4149 9.3005
R10890 gnd.n4152 gnd.n4151 9.3005
R10891 gnd.n3302 gnd.n3300 9.3005
R10892 gnd.n4246 gnd.n4245 9.3005
R10893 gnd.n4244 gnd.n3301 9.3005
R10894 gnd.n4243 gnd.n4242 9.3005
R10895 gnd.n4241 gnd.n3303 9.3005
R10896 gnd.n4240 gnd.n4239 9.3005
R10897 gnd.n4238 gnd.n4224 9.3005
R10898 gnd.n4237 gnd.n4236 9.3005
R10899 gnd.n4235 gnd.n4225 9.3005
R10900 gnd.n4234 gnd.n4233 9.3005
R10901 gnd.n4232 gnd.n4229 9.3005
R10902 gnd.n4231 gnd.n4230 9.3005
R10903 gnd.n3234 gnd.n3233 9.3005
R10904 gnd.n4376 gnd.n4375 9.3005
R10905 gnd.n4377 gnd.n3231 9.3005
R10906 gnd.n4380 gnd.n4379 9.3005
R10907 gnd.n4378 gnd.n3232 9.3005
R10908 gnd.n3212 gnd.n3211 9.3005
R10909 gnd.n4408 gnd.n4407 9.3005
R10910 gnd.n4409 gnd.n3209 9.3005
R10911 gnd.n4425 gnd.n4424 9.3005
R10912 gnd.n4423 gnd.n3210 9.3005
R10913 gnd.n4422 gnd.n4421 9.3005
R10914 gnd.n4420 gnd.n4410 9.3005
R10915 gnd.n4419 gnd.n4418 9.3005
R10916 gnd.n4417 gnd.n4414 9.3005
R10917 gnd.n4416 gnd.n4415 9.3005
R10918 gnd.n3160 gnd.n3159 9.3005
R10919 gnd.n4518 gnd.n4517 9.3005
R10920 gnd.n4519 gnd.n3157 9.3005
R10921 gnd.n4522 gnd.n4521 9.3005
R10922 gnd.n4520 gnd.n3158 9.3005
R10923 gnd.n3136 gnd.n3135 9.3005
R10924 gnd.n4550 gnd.n4549 9.3005
R10925 gnd.n4551 gnd.n3133 9.3005
R10926 gnd.n4567 gnd.n4566 9.3005
R10927 gnd.n4565 gnd.n3134 9.3005
R10928 gnd.n4564 gnd.n4563 9.3005
R10929 gnd.n4562 gnd.n4552 9.3005
R10930 gnd.n4561 gnd.n4560 9.3005
R10931 gnd.n4559 gnd.n4556 9.3005
R10932 gnd.n4558 gnd.n4557 9.3005
R10933 gnd.n3084 gnd.n3083 9.3005
R10934 gnd.n4644 gnd.n4643 9.3005
R10935 gnd.n4645 gnd.n3081 9.3005
R10936 gnd.n4662 gnd.n4661 9.3005
R10937 gnd.n4660 gnd.n3082 9.3005
R10938 gnd.n4659 gnd.n4658 9.3005
R10939 gnd.n4657 gnd.n4646 9.3005
R10940 gnd.n4656 gnd.n4655 9.3005
R10941 gnd.n4654 gnd.n4651 9.3005
R10942 gnd.n4653 gnd.n4652 9.3005
R10943 gnd.n3032 gnd.n3031 9.3005
R10944 gnd.n4728 gnd.n4727 9.3005
R10945 gnd.n4729 gnd.n3030 9.3005
R10946 gnd.n4731 gnd.n4730 9.3005
R10947 gnd.n4732 gnd.n3029 9.3005
R10948 gnd.n4738 gnd.n4737 9.3005
R10949 gnd.n4739 gnd.n3027 9.3005
R10950 gnd.n4755 gnd.n4754 9.3005
R10951 gnd.n4753 gnd.n3028 9.3005
R10952 gnd.n4752 gnd.n4751 9.3005
R10953 gnd.n4750 gnd.n4740 9.3005
R10954 gnd.n4749 gnd.n4748 9.3005
R10955 gnd.n4747 gnd.n4744 9.3005
R10956 gnd.n4746 gnd.n4745 9.3005
R10957 gnd.n2929 gnd.n2928 9.3005
R10958 gnd.n4991 gnd.n4990 9.3005
R10959 gnd.n4992 gnd.n2927 9.3005
R10960 gnd.n4994 gnd.n4993 9.3005
R10961 gnd.n2918 gnd.n2917 9.3005
R10962 gnd.n5009 gnd.n5008 9.3005
R10963 gnd.n5010 gnd.n2916 9.3005
R10964 gnd.n5012 gnd.n5011 9.3005
R10965 gnd.n2906 gnd.n2905 9.3005
R10966 gnd.n5028 gnd.n5027 9.3005
R10967 gnd.n5029 gnd.n2904 9.3005
R10968 gnd.n5049 gnd.n5048 9.3005
R10969 gnd.n3438 gnd.n3437 9.3005
R10970 gnd.n5045 gnd.n5030 9.3005
R10971 gnd.n5044 gnd.n5043 9.3005
R10972 gnd.n5042 gnd.n5033 9.3005
R10973 gnd.n5041 gnd.n5040 9.3005
R10974 gnd.n5039 gnd.n5034 9.3005
R10975 gnd.n2876 gnd.n2874 9.3005
R10976 gnd.n5047 gnd.n5046 9.3005
R10977 gnd.n5404 gnd.n5403 9.3005
R10978 gnd.n2755 gnd.n2753 9.3005
R10979 gnd.n5240 gnd.n5239 9.3005
R10980 gnd.n5242 gnd.n5241 9.3005
R10981 gnd.n5229 gnd.n5228 9.3005
R10982 gnd.n5248 gnd.n5247 9.3005
R10983 gnd.n5250 gnd.n5249 9.3005
R10984 gnd.n5219 gnd.n5218 9.3005
R10985 gnd.n5256 gnd.n5255 9.3005
R10986 gnd.n5258 gnd.n5257 9.3005
R10987 gnd.n5209 gnd.n5208 9.3005
R10988 gnd.n5264 gnd.n5263 9.3005
R10989 gnd.n5266 gnd.n5265 9.3005
R10990 gnd.n5199 gnd.n5198 9.3005
R10991 gnd.n5272 gnd.n5271 9.3005
R10992 gnd.n5274 gnd.n5273 9.3005
R10993 gnd.n5195 gnd.n2882 9.3005
R10994 gnd.n5402 gnd.n2764 9.3005
R10995 gnd.n2759 gnd.n2757 9.3005
R10996 gnd.n5279 gnd.n5278 9.3005
R10997 gnd.n5277 gnd.n2875 9.3005
R10998 gnd.n5276 gnd.n5275 9.3005
R10999 gnd.n2883 gnd.n2881 9.3005
R11000 gnd.n5270 gnd.n5269 9.3005
R11001 gnd.n5268 gnd.n5267 9.3005
R11002 gnd.n5203 gnd.n5202 9.3005
R11003 gnd.n5262 gnd.n5261 9.3005
R11004 gnd.n5260 gnd.n5259 9.3005
R11005 gnd.n5215 gnd.n5214 9.3005
R11006 gnd.n5254 gnd.n5253 9.3005
R11007 gnd.n5252 gnd.n5251 9.3005
R11008 gnd.n5223 gnd.n5222 9.3005
R11009 gnd.n5246 gnd.n5245 9.3005
R11010 gnd.n5244 gnd.n5243 9.3005
R11011 gnd.n5235 gnd.n5234 9.3005
R11012 gnd.n5238 gnd.n2749 9.3005
R11013 gnd.n5406 gnd.n5405 9.3005
R11014 gnd.n2760 gnd.n2754 9.3005
R11015 gnd.n2763 gnd.n2762 9.3005
R11016 gnd.n2758 gnd.n2729 9.3005
R11017 gnd.n5139 gnd.n5138 9.3005
R11018 gnd.n5140 gnd.n5133 9.3005
R11019 gnd.n5142 gnd.n5141 9.3005
R11020 gnd.n5162 gnd.n5132 9.3005
R11021 gnd.n5164 gnd.n5163 9.3005
R11022 gnd.n5165 gnd.n5130 9.3005
R11023 gnd.n5168 gnd.n5167 9.3005
R11024 gnd.n5166 gnd.n5131 9.3005
R11025 gnd.n227 gnd.n226 9.3005
R11026 gnd.n6764 gnd.n6763 9.3005
R11027 gnd.n6765 gnd.n224 9.3005
R11028 gnd.n6768 gnd.n6767 9.3005
R11029 gnd.n6766 gnd.n225 9.3005
R11030 gnd.n200 gnd.n199 9.3005
R11031 gnd.n6799 gnd.n6798 9.3005
R11032 gnd.n6800 gnd.n197 9.3005
R11033 gnd.n6807 gnd.n6806 9.3005
R11034 gnd.n6805 gnd.n198 9.3005
R11035 gnd.n6804 gnd.n6803 9.3005
R11036 gnd.n6802 gnd.n67 9.3005
R11037 gnd.n5135 gnd.n5134 9.3005
R11038 gnd.n7269 gnd.n68 9.3005
R11039 gnd.t3 gnd.n1764 9.24152
R11040 gnd.n5998 gnd.t211 9.24152
R11041 gnd.n885 gnd.t310 9.24152
R11042 gnd.t132 gnd.n2413 9.24152
R11043 gnd.n4279 gnd.t67 9.24152
R11044 gnd.n4289 gnd.t67 9.24152
R11045 gnd.n4647 gnd.t105 9.24152
R11046 gnd.n4684 gnd.t105 9.24152
R11047 gnd.n6743 gnd.t14 9.24152
R11048 gnd.t48 gnd.t3 8.92286
R11049 gnd.t164 gnd.n4211 8.92286
R11050 gnd.n4697 gnd.t41 8.92286
R11051 gnd.n4786 gnd.t282 8.92286
R11052 gnd.n2124 gnd.n2099 8.92171
R11053 gnd.n2092 gnd.n2067 8.92171
R11054 gnd.n2060 gnd.n2035 8.92171
R11055 gnd.n2029 gnd.n2004 8.92171
R11056 gnd.n1997 gnd.n1972 8.92171
R11057 gnd.n1965 gnd.n1940 8.92171
R11058 gnd.n1933 gnd.n1908 8.92171
R11059 gnd.n1902 gnd.n1877 8.92171
R11060 gnd.n4839 gnd.n4821 8.72777
R11061 gnd.n1122 gnd.t38 8.60421
R11062 gnd.t17 gnd.n3187 8.60421
R11063 gnd.t112 gnd.n3163 8.60421
R11064 gnd.n1148 gnd.n1136 8.43656
R11065 gnd.n42 gnd.n30 8.43656
R11066 gnd.n4282 gnd.n4281 8.28555
R11067 gnd.n4312 gnd.n4311 8.28555
R11068 gnd.n4319 gnd.n3192 8.28555
R11069 gnd.n4537 gnd.n4536 8.28555
R11070 gnd.n4594 gnd.n3109 8.28555
R11071 gnd.n4683 gnd.n3064 8.28555
R11072 gnd.n4757 gnd.t282 8.28555
R11073 gnd.n2125 gnd.n2097 8.14595
R11074 gnd.n2093 gnd.n2065 8.14595
R11075 gnd.n2061 gnd.n2033 8.14595
R11076 gnd.n2030 gnd.n2002 8.14595
R11077 gnd.n1998 gnd.n1970 8.14595
R11078 gnd.n1966 gnd.n1938 8.14595
R11079 gnd.n1934 gnd.n1906 8.14595
R11080 gnd.n1903 gnd.n1875 8.14595
R11081 gnd.n3770 gnd.n0 8.10675
R11082 gnd.n7270 gnd.n7269 8.10675
R11083 gnd.n2130 gnd.n2129 7.97301
R11084 gnd.t56 gnd.n1664 7.9669
R11085 gnd.n3989 gnd.n3398 7.9669
R11086 gnd.t94 gnd.n3290 7.9669
R11087 gnd.n4715 gnd.t165 7.9669
R11088 gnd.n5408 gnd.n2746 7.9669
R11089 gnd.n7270 gnd.n66 7.78567
R11090 gnd.n5402 gnd.n2757 7.75808
R11091 gnd.n6991 gnd.n6894 7.75808
R11092 gnd.n3928 gnd.n3927 7.75808
R11093 gnd.n3725 gnd.n3724 7.75808
R11094 gnd.n4029 gnd.t270 7.64824
R11095 gnd.n4282 gnd.t89 7.64824
R11096 gnd.n4316 gnd.t78 7.64824
R11097 gnd.n4460 gnd.t16 7.64824
R11098 gnd.n3064 gnd.t93 7.64824
R11099 gnd.n1173 gnd.n1172 7.53171
R11100 gnd.n1597 gnd.t103 7.32958
R11101 gnd.t247 gnd.n3384 7.32958
R11102 gnd.n4053 gnd.t167 7.32958
R11103 gnd.n5620 gnd.n2579 7.32958
R11104 gnd.n4980 gnd.n4978 7.32958
R11105 gnd.t322 gnd.n2931 7.32958
R11106 gnd.n5025 gnd.t215 7.32958
R11107 gnd.n2601 gnd.n2600 7.30353
R11108 gnd.n4838 gnd.n4837 7.30353
R11109 gnd.n1557 gnd.n1276 7.01093
R11110 gnd.n1279 gnd.n1277 7.01093
R11111 gnd.n1567 gnd.n1566 7.01093
R11112 gnd.n1578 gnd.n1260 7.01093
R11113 gnd.n1577 gnd.n1263 7.01093
R11114 gnd.n1588 gnd.n1251 7.01093
R11115 gnd.n1254 gnd.n1252 7.01093
R11116 gnd.n1598 gnd.n1597 7.01093
R11117 gnd.n1608 gnd.n1232 7.01093
R11118 gnd.n1607 gnd.n1235 7.01093
R11119 gnd.n1624 gnd.n1225 7.01093
R11120 gnd.n1634 gnd.n1216 7.01093
R11121 gnd.n1645 gnd.n1644 7.01093
R11122 gnd.n1665 gnd.n1201 7.01093
R11123 gnd.n1664 gnd.n1180 7.01093
R11124 gnd.n1682 gnd.n1181 7.01093
R11125 gnd.n1676 gnd.n1675 7.01093
R11126 gnd.n1692 gnd.n1045 7.01093
R11127 gnd.n1702 gnd.n1037 7.01093
R11128 gnd.n1713 gnd.n1028 7.01093
R11129 gnd.n1122 gnd.n1121 7.01093
R11130 gnd.n1723 gnd.n1722 7.01093
R11131 gnd.n1734 gnd.n1011 7.01093
R11132 gnd.n1733 gnd.n1014 7.01093
R11133 gnd.n1744 gnd.n1003 7.01093
R11134 gnd.n1754 gnd.n1753 7.01093
R11135 gnd.n1765 gnd.n985 7.01093
R11136 gnd.n1764 gnd.n988 7.01093
R11137 gnd.n1775 gnd.n976 7.01093
R11138 gnd.n979 gnd.n977 7.01093
R11139 gnd.n1785 gnd.n1784 7.01093
R11140 gnd.n1796 gnd.n960 7.01093
R11141 gnd.n954 gnd.n952 7.01093
R11142 gnd.n1816 gnd.n1815 7.01093
R11143 gnd.n1827 gnd.n935 7.01093
R11144 gnd.n1826 gnd.n938 7.01093
R11145 gnd.n1837 gnd.n926 7.01093
R11146 gnd.n929 gnd.n927 7.01093
R11147 gnd.n1858 gnd.n909 7.01093
R11148 gnd.n1857 gnd.n912 7.01093
R11149 gnd.n1869 gnd.n901 7.01093
R11150 gnd.n902 gnd.n894 7.01093
R11151 gnd.n2135 gnd.n2134 7.01093
R11152 gnd.n2145 gnd.n885 7.01093
R11153 gnd.n5992 gnd.n773 7.01093
R11154 gnd.n5991 gnd.n776 7.01093
R11155 gnd.n5550 gnd.n5549 7.01093
R11156 gnd.n4184 gnd.n3328 7.01093
R11157 gnd.n4344 gnd.n4343 7.01093
R11158 gnd.n4453 gnd.n3188 7.01093
R11159 gnd.n3166 gnd.n3154 7.01093
R11160 gnd.n4631 gnd.n3095 7.01093
R11161 gnd.n4779 gnd.n3000 7.01093
R11162 gnd.n4816 gnd.n2983 7.01093
R11163 gnd.n1235 gnd.t40 6.69227
R11164 gnd.n1765 gnd.t48 6.69227
R11165 gnd.n1847 gnd.t147 6.69227
R11166 gnd.n4971 gnd.n4970 6.5566
R11167 gnd.n4069 gnd.n4068 6.5566
R11168 gnd.n5561 gnd.n5557 6.5566
R11169 gnd.n4849 gnd.n4848 6.5566
R11170 gnd.n3514 gnd.n3506 6.20656
R11171 gnd.n2760 gnd.n2752 6.20656
R11172 gnd.t6 gnd.n1656 6.05496
R11173 gnd.n1657 gnd.t5 6.05496
R11174 gnd.n1722 gnd.t11 6.05496
R11175 gnd.n1096 gnd.t58 6.05496
R11176 gnd.n2127 gnd.n2097 5.81868
R11177 gnd.n2095 gnd.n2065 5.81868
R11178 gnd.n2063 gnd.n2033 5.81868
R11179 gnd.n2032 gnd.n2002 5.81868
R11180 gnd.n2000 gnd.n1970 5.81868
R11181 gnd.n1968 gnd.n1938 5.81868
R11182 gnd.n1936 gnd.n1906 5.81868
R11183 gnd.n1905 gnd.n1875 5.81868
R11184 gnd.n4164 gnd.n4163 5.73631
R11185 gnd.n4184 gnd.t204 5.73631
R11186 gnd.n3275 gnd.t92 5.73631
R11187 gnd.n4306 gnd.n3260 5.73631
R11188 gnd.n4351 gnd.n3252 5.73631
R11189 gnd.n4332 gnd.t77 5.73631
R11190 gnd.n3188 gnd.t145 5.73631
R11191 gnd.n4505 gnd.n3172 5.73631
R11192 gnd.n4486 gnd.n3175 5.73631
R11193 gnd.n3166 gnd.t29 5.73631
R11194 gnd.n4576 gnd.t315 5.73631
R11195 gnd.n4641 gnd.n3086 5.73631
R11196 gnd.n3089 gnd.n3078 5.73631
R11197 gnd.t90 gnd.n4672 5.73631
R11198 gnd.n4800 gnd.n4799 5.73631
R11199 gnd.n4910 gnd.t240 5.73631
R11200 gnd.n4975 gnd.n2836 5.62001
R11201 gnd.n5623 gnd.n2544 5.62001
R11202 gnd.n5623 gnd.n2545 5.62001
R11203 gnd.n4844 gnd.n2836 5.62001
R11204 gnd.n1416 gnd.n1411 5.4308
R11205 gnd.n877 gnd.n807 5.4308
R11206 gnd.n1734 gnd.t102 5.41765
R11207 gnd.t57 gnd.n996 5.41765
R11208 gnd.n1806 gnd.t108 5.41765
R11209 gnd.n2125 gnd.n2124 5.04292
R11210 gnd.n2093 gnd.n2092 5.04292
R11211 gnd.n2061 gnd.n2060 5.04292
R11212 gnd.n2030 gnd.n2029 5.04292
R11213 gnd.n1998 gnd.n1997 5.04292
R11214 gnd.n1966 gnd.n1965 5.04292
R11215 gnd.n1934 gnd.n1933 5.04292
R11216 gnd.n1903 gnd.n1902 5.04292
R11217 gnd.n1703 gnd.t71 4.78034
R11218 gnd.n979 gnd.t23 4.78034
R11219 gnd.n5999 gnd.n5998 4.78034
R11220 gnd.n5543 gnd.t30 4.78034
R11221 gnd.n4351 gnd.t153 4.78034
R11222 gnd.t32 gnd.n3086 4.78034
R11223 gnd.n4808 gnd.t118 4.78034
R11224 gnd.n4978 gnd.t219 4.78034
R11225 gnd.n1177 gnd.n1174 4.74817
R11226 gnd.n1689 gnd.n1047 4.74817
R11227 gnd.n1687 gnd.n1048 4.74817
R11228 gnd.n1125 gnd.n1119 4.74817
R11229 gnd.n1193 gnd.n1174 4.74817
R11230 gnd.n1192 gnd.n1047 4.74817
R11231 gnd.n1688 gnd.n1687 4.74817
R11232 gnd.n1125 gnd.n1124 4.74817
R11233 gnd.n1172 gnd.n1171 4.74296
R11234 gnd.n66 gnd.n65 4.74296
R11235 gnd.n1148 gnd.n1147 4.7074
R11236 gnd.n1160 gnd.n1159 4.7074
R11237 gnd.n42 gnd.n41 4.7074
R11238 gnd.n54 gnd.n53 4.7074
R11239 gnd.n1172 gnd.n1160 4.65959
R11240 gnd.n66 gnd.n54 4.65959
R11241 gnd.n5344 gnd.n2838 4.6132
R11242 gnd.n5624 gnd.n2543 4.6132
R11243 gnd.n4141 gnd.n4140 4.46168
R11244 gnd.n4171 gnd.n3338 4.46168
R11245 gnd.t111 gnd.n3310 4.46168
R11246 gnd.n4299 gnd.n3257 4.46168
R11247 gnd.n4363 gnd.n3245 4.46168
R11248 gnd.n4493 gnd.n3181 4.46168
R11249 gnd.n4515 gnd.n3162 4.46168
R11250 gnd.n4611 gnd.n3098 4.46168
R11251 gnd.n4666 gnd.n4665 4.46168
R11252 gnd.n4772 gnd.t0 4.46168
R11253 gnd.n4757 gnd.n2995 4.46168
R11254 gnd.n4741 gnd.n2991 4.46168
R11255 gnd.n4834 gnd.n4821 4.46111
R11256 gnd.n2110 gnd.n2106 4.38594
R11257 gnd.n2078 gnd.n2074 4.38594
R11258 gnd.n2046 gnd.n2042 4.38594
R11259 gnd.n2015 gnd.n2011 4.38594
R11260 gnd.n1983 gnd.n1979 4.38594
R11261 gnd.n1951 gnd.n1947 4.38594
R11262 gnd.n1919 gnd.n1915 4.38594
R11263 gnd.n1888 gnd.n1884 4.38594
R11264 gnd.n2121 gnd.n2099 4.26717
R11265 gnd.n2089 gnd.n2067 4.26717
R11266 gnd.n2057 gnd.n2035 4.26717
R11267 gnd.n2026 gnd.n2004 4.26717
R11268 gnd.n1994 gnd.n1972 4.26717
R11269 gnd.n1962 gnd.n1940 4.26717
R11270 gnd.n1930 gnd.n1908 4.26717
R11271 gnd.n1899 gnd.n1877 4.26717
R11272 gnd.t4 gnd.n1208 4.14303
R11273 gnd.n938 gnd.t39 4.14303
R11274 gnd.t243 gnd.n2464 4.14303
R11275 gnd.n4428 gnd.t116 4.14303
R11276 gnd.t138 gnd.n3139 4.14303
R11277 gnd.t207 gnd.n5071 4.14303
R11278 gnd.n2129 gnd.n2128 4.08274
R11279 gnd.n4970 gnd.n4969 4.05904
R11280 gnd.n4070 gnd.n4069 4.05904
R11281 gnd.n5564 gnd.n5557 4.05904
R11282 gnd.n4850 gnd.n4849 4.05904
R11283 gnd.n19 gnd.n9 3.99943
R11284 gnd.n4171 gnd.t304 3.82437
R11285 gnd.n3324 gnd.t111 3.82437
R11286 gnd.n4343 gnd.t42 3.82437
R11287 gnd.n4631 gnd.t28 3.82437
R11288 gnd.n4734 gnd.t0 3.82437
R11289 gnd.n1686 gnd.n1173 3.81325
R11290 gnd.n1160 gnd.n1148 3.72967
R11291 gnd.n54 gnd.n42 3.72967
R11292 gnd.n2129 gnd.n2001 3.70378
R11293 gnd.n19 gnd.n18 3.60163
R11294 gnd.t136 gnd.n4190 3.50571
R11295 gnd.n4733 gnd.t158 3.50571
R11296 gnd.n2120 gnd.n2101 3.49141
R11297 gnd.n2088 gnd.n2069 3.49141
R11298 gnd.n2056 gnd.n2037 3.49141
R11299 gnd.n2025 gnd.n2006 3.49141
R11300 gnd.n1993 gnd.n1974 3.49141
R11301 gnd.n1961 gnd.n1942 3.49141
R11302 gnd.n1929 gnd.n1910 3.49141
R11303 gnd.n1898 gnd.n1879 3.49141
R11304 gnd.n7161 gnd.n7158 3.29747
R11305 gnd.n7162 gnd.n7161 3.29747
R11306 gnd.n5362 gnd.n5361 3.29747
R11307 gnd.n5361 gnd.n5360 3.29747
R11308 gnd.n5893 gnd.n5892 3.29747
R11309 gnd.n5892 gnd.n5891 3.29747
R11310 gnd.n5642 gnd.n5641 3.29747
R11311 gnd.n5641 gnd.n5640 3.29747
R11312 gnd.n4029 gnd.n2605 3.18706
R11313 gnd.n4191 gnd.n3320 3.18706
R11314 gnd.n4289 gnd.n4288 3.18706
R11315 gnd.n4373 gnd.n3236 3.18706
R11316 gnd.n4446 gnd.n3186 3.18706
R11317 gnd.n4525 gnd.n4524 3.18706
R11318 gnd.n4618 gnd.n3103 3.18706
R11319 gnd.n4647 gnd.n3074 3.18706
R11320 gnd.n4780 gnd.n3005 3.18706
R11321 gnd.t261 gnd.n4798 3.18706
R11322 gnd.n4910 gnd.n2937 3.18706
R11323 gnd.n1215 gnd.t4 2.8684
R11324 gnd.n4249 gnd.t94 2.8684
R11325 gnd.t165 gnd.n3046 2.8684
R11326 gnd.n1161 gnd.t176 2.82907
R11327 gnd.n1161 gnd.t324 2.82907
R11328 gnd.n1163 gnd.t175 2.82907
R11329 gnd.n1163 gnd.t101 2.82907
R11330 gnd.n1165 gnd.t87 2.82907
R11331 gnd.n1165 gnd.t88 2.82907
R11332 gnd.n1167 gnd.t187 2.82907
R11333 gnd.n1167 gnd.t46 2.82907
R11334 gnd.n1169 gnd.t44 2.82907
R11335 gnd.n1169 gnd.t127 2.82907
R11336 gnd.n1126 gnd.t133 2.82907
R11337 gnd.n1126 gnd.t183 2.82907
R11338 gnd.n1128 gnd.t170 2.82907
R11339 gnd.n1128 gnd.t84 2.82907
R11340 gnd.n1130 gnd.t163 2.82907
R11341 gnd.n1130 gnd.t321 2.82907
R11342 gnd.n1132 gnd.t129 2.82907
R11343 gnd.n1132 gnd.t148 2.82907
R11344 gnd.n1134 gnd.t160 2.82907
R11345 gnd.n1134 gnd.t186 2.82907
R11346 gnd.n1137 gnd.t157 2.82907
R11347 gnd.n1137 gnd.t134 2.82907
R11348 gnd.n1139 gnd.t190 2.82907
R11349 gnd.n1139 gnd.t151 2.82907
R11350 gnd.n1141 gnd.t192 2.82907
R11351 gnd.n1141 gnd.t329 2.82907
R11352 gnd.n1143 gnd.t61 2.82907
R11353 gnd.n1143 gnd.t326 2.82907
R11354 gnd.n1145 gnd.t189 2.82907
R11355 gnd.n1145 gnd.t177 2.82907
R11356 gnd.n1149 gnd.t142 2.82907
R11357 gnd.n1149 gnd.t124 2.82907
R11358 gnd.n1151 gnd.t122 2.82907
R11359 gnd.n1151 gnd.t161 2.82907
R11360 gnd.n1153 gnd.t181 2.82907
R11361 gnd.n1153 gnd.t22 2.82907
R11362 gnd.n1155 gnd.t144 2.82907
R11363 gnd.n1155 gnd.t146 2.82907
R11364 gnd.n1157 gnd.t174 2.82907
R11365 gnd.n1157 gnd.t37 2.82907
R11366 gnd.n63 gnd.t135 2.82907
R11367 gnd.n63 gnd.t47 2.82907
R11368 gnd.n61 gnd.t120 2.82907
R11369 gnd.n61 gnd.t335 2.82907
R11370 gnd.n59 gnd.t313 2.82907
R11371 gnd.n59 gnd.t100 2.82907
R11372 gnd.n57 gnd.t156 2.82907
R11373 gnd.n57 gnd.t63 2.82907
R11374 gnd.n55 gnd.t35 2.82907
R11375 gnd.n55 gnd.t82 2.82907
R11376 gnd.n28 gnd.t191 2.82907
R11377 gnd.n28 gnd.t178 2.82907
R11378 gnd.n26 gnd.t80 2.82907
R11379 gnd.n26 gnd.t319 2.82907
R11380 gnd.n24 gnd.t179 2.82907
R11381 gnd.n24 gnd.t188 2.82907
R11382 gnd.n22 gnd.t333 2.82907
R11383 gnd.n22 gnd.t328 2.82907
R11384 gnd.n20 gnd.t325 2.82907
R11385 gnd.n20 gnd.t72 2.82907
R11386 gnd.n39 gnd.t55 2.82907
R11387 gnd.n39 gnd.t130 2.82907
R11388 gnd.n37 gnd.t107 2.82907
R11389 gnd.n37 gnd.t115 2.82907
R11390 gnd.n35 gnd.t141 2.82907
R11391 gnd.n35 gnd.t53 2.82907
R11392 gnd.n33 gnd.t184 2.82907
R11393 gnd.n33 gnd.t128 2.82907
R11394 gnd.n31 gnd.t182 2.82907
R11395 gnd.n31 gnd.t15 2.82907
R11396 gnd.n51 gnd.t171 2.82907
R11397 gnd.n51 gnd.t10 2.82907
R11398 gnd.n49 gnd.t318 2.82907
R11399 gnd.n49 gnd.t185 2.82907
R11400 gnd.n47 gnd.t327 2.82907
R11401 gnd.n47 gnd.t162 2.82907
R11402 gnd.n45 gnd.t99 2.82907
R11403 gnd.n45 gnd.t152 2.82907
R11404 gnd.n43 gnd.t64 2.82907
R11405 gnd.n43 gnd.t330 2.82907
R11406 gnd.n2117 gnd.n2116 2.71565
R11407 gnd.n2085 gnd.n2084 2.71565
R11408 gnd.n2053 gnd.n2052 2.71565
R11409 gnd.n2022 gnd.n2021 2.71565
R11410 gnd.n1990 gnd.n1989 2.71565
R11411 gnd.n1958 gnd.n1957 2.71565
R11412 gnd.n1926 gnd.n1925 2.71565
R11413 gnd.n1895 gnd.n1894 2.71565
R11414 gnd.n5543 gnd.t226 2.54975
R11415 gnd.t13 gnd.n3258 2.54975
R11416 gnd.n4312 gnd.t50 2.54975
R11417 gnd.n4594 gnd.t314 2.54975
R11418 gnd.t8 gnd.n3087 2.54975
R11419 gnd.n1686 gnd.n1174 2.27742
R11420 gnd.n1686 gnd.n1047 2.27742
R11421 gnd.n1687 gnd.n1686 2.27742
R11422 gnd.n1686 gnd.n1125 2.27742
R11423 gnd.n1566 gnd.t257 2.23109
R11424 gnd.n1691 gnd.t71 2.23109
R11425 gnd.n5999 gnd.n763 2.23109
R11426 gnd.n5724 gnd.n2393 2.23109
R11427 gnd.n6796 gnd.n203 2.23109
R11428 gnd.n2113 gnd.n2103 1.93989
R11429 gnd.n2081 gnd.n2071 1.93989
R11430 gnd.n2049 gnd.n2039 1.93989
R11431 gnd.n2018 gnd.n2008 1.93989
R11432 gnd.n1986 gnd.n1976 1.93989
R11433 gnd.n1954 gnd.n1944 1.93989
R11434 gnd.n1922 gnd.n1912 1.93989
R11435 gnd.n1891 gnd.n1881 1.93989
R11436 gnd.n4205 gnd.n4204 1.91244
R11437 gnd.n4269 gnd.n4268 1.91244
R11438 gnd.n4436 gnd.n4434 1.91244
R11439 gnd.n4475 gnd.n4474 1.91244
R11440 gnd.n4690 gnd.n3058 1.91244
R11441 gnd.n4765 gnd.n3009 1.91244
R11442 gnd.n4741 gnd.t198 1.91244
R11443 gnd.t73 gnd.n1577 1.59378
R11444 gnd.n1004 gnd.t57 1.59378
R11445 gnd.n1097 gnd.t108 1.59378
R11446 gnd.t316 gnd.n4382 1.59378
R11447 gnd.n4587 gnd.t65 1.59378
R11448 gnd.n4061 gnd.t201 1.27512
R11449 gnd.t92 gnd.n3264 1.27512
R11450 gnd.n4673 gnd.t90 1.27512
R11451 gnd.t75 gnd.n135 1.27512
R11452 gnd.n1419 gnd.n1411 1.16414
R11453 gnd.n874 gnd.n807 1.16414
R11454 gnd.n2112 gnd.n2105 1.16414
R11455 gnd.n2080 gnd.n2073 1.16414
R11456 gnd.n2048 gnd.n2041 1.16414
R11457 gnd.n2017 gnd.n2010 1.16414
R11458 gnd.n1985 gnd.n1978 1.16414
R11459 gnd.n1953 gnd.n1946 1.16414
R11460 gnd.n1921 gnd.n1914 1.16414
R11461 gnd.n1890 gnd.n1883 1.16414
R11462 gnd.n5344 gnd.n5343 0.970197
R11463 gnd.n5624 gnd.n2541 0.970197
R11464 gnd.n2096 gnd.n2064 0.962709
R11465 gnd.n2128 gnd.n2096 0.962709
R11466 gnd.n1969 gnd.n1937 0.962709
R11467 gnd.n2001 gnd.n1969 0.962709
R11468 gnd.n1657 gnd.t6 0.956468
R11469 gnd.n1795 gnd.t58 0.956468
R11470 gnd.n5778 gnd.t43 0.956468
R11471 gnd.n5706 gnd.t123 0.956468
R11472 gnd.t69 gnd.n2436 0.956468
R11473 gnd.n4137 gnd.t30 0.956468
R11474 gnd.t118 gnd.n4806 0.956468
R11475 gnd.t26 gnd.n5127 0.956468
R11476 gnd.n5102 gnd.t34 0.956468
R11477 gnd.n7234 gnd.t9 0.956468
R11478 gnd.n2 gnd.n1 0.672012
R11479 gnd.n3 gnd.n2 0.672012
R11480 gnd.n4 gnd.n3 0.672012
R11481 gnd.n5 gnd.n4 0.672012
R11482 gnd.n6 gnd.n5 0.672012
R11483 gnd.n7 gnd.n6 0.672012
R11484 gnd.n8 gnd.n7 0.672012
R11485 gnd.n9 gnd.n8 0.672012
R11486 gnd.n11 gnd.n10 0.672012
R11487 gnd.n12 gnd.n11 0.672012
R11488 gnd.n13 gnd.n12 0.672012
R11489 gnd.n14 gnd.n13 0.672012
R11490 gnd.n15 gnd.n14 0.672012
R11491 gnd.n16 gnd.n15 0.672012
R11492 gnd.n17 gnd.n16 0.672012
R11493 gnd.n18 gnd.n17 0.672012
R11494 gnd.n4165 gnd.t232 0.637812
R11495 gnd.n4212 gnd.n3297 0.637812
R11496 gnd.n4260 gnd.n4259 0.637812
R11497 gnd.n4259 gnd.t85 0.637812
R11498 gnd.n4332 gnd.n4331 0.637812
R11499 gnd.n4316 gnd.n4315 0.637812
R11500 gnd.n4319 gnd.t91 0.637812
R11501 gnd.n4536 gnd.t110 0.637812
R11502 gnd.n4460 gnd.n3130 0.637812
R11503 gnd.n4577 gnd.n4576 0.637812
R11504 gnd.t51 gnd.n3043 0.637812
R11505 gnd.n4716 gnd.n3043 0.637812
R11506 gnd.n4725 gnd.n3036 0.637812
R11507 gnd.n4798 gnd.t222 0.637812
R11508 gnd gnd.n0 0.624033
R11509 gnd.n1171 gnd.n1170 0.573776
R11510 gnd.n1170 gnd.n1168 0.573776
R11511 gnd.n1168 gnd.n1166 0.573776
R11512 gnd.n1166 gnd.n1164 0.573776
R11513 gnd.n1164 gnd.n1162 0.573776
R11514 gnd.n1136 gnd.n1135 0.573776
R11515 gnd.n1135 gnd.n1133 0.573776
R11516 gnd.n1133 gnd.n1131 0.573776
R11517 gnd.n1131 gnd.n1129 0.573776
R11518 gnd.n1129 gnd.n1127 0.573776
R11519 gnd.n1147 gnd.n1146 0.573776
R11520 gnd.n1146 gnd.n1144 0.573776
R11521 gnd.n1144 gnd.n1142 0.573776
R11522 gnd.n1142 gnd.n1140 0.573776
R11523 gnd.n1140 gnd.n1138 0.573776
R11524 gnd.n1159 gnd.n1158 0.573776
R11525 gnd.n1158 gnd.n1156 0.573776
R11526 gnd.n1156 gnd.n1154 0.573776
R11527 gnd.n1154 gnd.n1152 0.573776
R11528 gnd.n1152 gnd.n1150 0.573776
R11529 gnd.n58 gnd.n56 0.573776
R11530 gnd.n60 gnd.n58 0.573776
R11531 gnd.n62 gnd.n60 0.573776
R11532 gnd.n64 gnd.n62 0.573776
R11533 gnd.n65 gnd.n64 0.573776
R11534 gnd.n23 gnd.n21 0.573776
R11535 gnd.n25 gnd.n23 0.573776
R11536 gnd.n27 gnd.n25 0.573776
R11537 gnd.n29 gnd.n27 0.573776
R11538 gnd.n30 gnd.n29 0.573776
R11539 gnd.n34 gnd.n32 0.573776
R11540 gnd.n36 gnd.n34 0.573776
R11541 gnd.n38 gnd.n36 0.573776
R11542 gnd.n40 gnd.n38 0.573776
R11543 gnd.n41 gnd.n40 0.573776
R11544 gnd.n46 gnd.n44 0.573776
R11545 gnd.n48 gnd.n46 0.573776
R11546 gnd.n50 gnd.n48 0.573776
R11547 gnd.n52 gnd.n50 0.573776
R11548 gnd.n53 gnd.n52 0.573776
R11549 gnd.n6990 gnd.n6989 0.532512
R11550 gnd.n3729 gnd.n3726 0.532512
R11551 gnd.n7024 gnd.n7023 0.497451
R11552 gnd.n5678 gnd.n5677 0.497451
R11553 gnd.n5080 gnd.n2808 0.497451
R11554 gnd.n2274 gnd.n2197 0.497451
R11555 gnd.n2151 gnd.n2150 0.486781
R11556 gnd.n1468 gnd.n1467 0.48678
R11557 gnd.n5937 gnd.n5936 0.480683
R11558 gnd.n1552 gnd.n1551 0.480683
R11559 gnd.n7271 gnd.n7270 0.4705
R11560 gnd.n5413 gnd.n5412 0.451719
R11561 gnd.n3994 gnd.n3993 0.451719
R11562 gnd.n3439 gnd.n3438 0.451719
R11563 gnd.n5048 gnd.n5047 0.451719
R11564 gnd.n6171 gnd.n593 0.438
R11565 gnd.n6524 gnd.n6523 0.438
R11566 gnd.n6735 gnd.n255 0.438
R11567 gnd.n3636 gnd.n3633 0.438
R11568 gnd.n3932 gnd.n3506 0.388379
R11569 gnd.n2109 gnd.n2108 0.388379
R11570 gnd.n2077 gnd.n2076 0.388379
R11571 gnd.n2045 gnd.n2044 0.388379
R11572 gnd.n2014 gnd.n2013 0.388379
R11573 gnd.n1982 gnd.n1981 0.388379
R11574 gnd.n1950 gnd.n1949 0.388379
R11575 gnd.n1918 gnd.n1917 0.388379
R11576 gnd.n1887 gnd.n1886 0.388379
R11577 gnd.n5406 gnd.n2752 0.388379
R11578 gnd.n7271 gnd.n19 0.374463
R11579 gnd gnd.n7271 0.367492
R11580 gnd.t147 gnd.n1846 0.319156
R11581 gnd.n5754 gnd.t45 0.319156
R11582 gnd.n5730 gnd.t121 0.319156
R11583 gnd.n4383 gnd.t316 0.319156
R11584 gnd.t145 gnd.t17 0.319156
R11585 gnd.t29 gnd.t112 0.319156
R11586 gnd.t65 gnd.n3117 0.319156
R11587 gnd.n6809 gnd.t62 0.319156
R11588 gnd.n7258 gnd.t79 0.319156
R11589 gnd.n1386 gnd.n1364 0.311721
R11590 gnd.n3866 gnd.n3395 0.302329
R11591 gnd.n5134 gnd.n2728 0.302329
R11592 gnd.n7205 gnd.n6875 0.293183
R11593 gnd.n5809 gnd.n2261 0.293183
R11594 gnd.n5982 gnd.n781 0.268793
R11595 gnd.n5282 gnd.n5281 0.258122
R11596 gnd.n7205 gnd.n7204 0.258122
R11597 gnd.n3614 gnd.n3446 0.258122
R11598 gnd.n5810 gnd.n5809 0.258122
R11599 gnd.n821 gnd.n781 0.241354
R11600 gnd.n2838 gnd.n2835 0.229039
R11601 gnd.n2839 gnd.n2838 0.229039
R11602 gnd.n2543 gnd.n2540 0.229039
R11603 gnd.n3542 gnd.n2543 0.229039
R11604 gnd.n1540 gnd.n1339 0.206293
R11605 gnd.n2126 gnd.n2098 0.155672
R11606 gnd.n2119 gnd.n2098 0.155672
R11607 gnd.n2119 gnd.n2118 0.155672
R11608 gnd.n2118 gnd.n2102 0.155672
R11609 gnd.n2111 gnd.n2102 0.155672
R11610 gnd.n2111 gnd.n2110 0.155672
R11611 gnd.n2094 gnd.n2066 0.155672
R11612 gnd.n2087 gnd.n2066 0.155672
R11613 gnd.n2087 gnd.n2086 0.155672
R11614 gnd.n2086 gnd.n2070 0.155672
R11615 gnd.n2079 gnd.n2070 0.155672
R11616 gnd.n2079 gnd.n2078 0.155672
R11617 gnd.n2062 gnd.n2034 0.155672
R11618 gnd.n2055 gnd.n2034 0.155672
R11619 gnd.n2055 gnd.n2054 0.155672
R11620 gnd.n2054 gnd.n2038 0.155672
R11621 gnd.n2047 gnd.n2038 0.155672
R11622 gnd.n2047 gnd.n2046 0.155672
R11623 gnd.n2031 gnd.n2003 0.155672
R11624 gnd.n2024 gnd.n2003 0.155672
R11625 gnd.n2024 gnd.n2023 0.155672
R11626 gnd.n2023 gnd.n2007 0.155672
R11627 gnd.n2016 gnd.n2007 0.155672
R11628 gnd.n2016 gnd.n2015 0.155672
R11629 gnd.n1999 gnd.n1971 0.155672
R11630 gnd.n1992 gnd.n1971 0.155672
R11631 gnd.n1992 gnd.n1991 0.155672
R11632 gnd.n1991 gnd.n1975 0.155672
R11633 gnd.n1984 gnd.n1975 0.155672
R11634 gnd.n1984 gnd.n1983 0.155672
R11635 gnd.n1967 gnd.n1939 0.155672
R11636 gnd.n1960 gnd.n1939 0.155672
R11637 gnd.n1960 gnd.n1959 0.155672
R11638 gnd.n1959 gnd.n1943 0.155672
R11639 gnd.n1952 gnd.n1943 0.155672
R11640 gnd.n1952 gnd.n1951 0.155672
R11641 gnd.n1935 gnd.n1907 0.155672
R11642 gnd.n1928 gnd.n1907 0.155672
R11643 gnd.n1928 gnd.n1927 0.155672
R11644 gnd.n1927 gnd.n1911 0.155672
R11645 gnd.n1920 gnd.n1911 0.155672
R11646 gnd.n1920 gnd.n1919 0.155672
R11647 gnd.n1904 gnd.n1876 0.155672
R11648 gnd.n1897 gnd.n1876 0.155672
R11649 gnd.n1897 gnd.n1896 0.155672
R11650 gnd.n1896 gnd.n1880 0.155672
R11651 gnd.n1889 gnd.n1880 0.155672
R11652 gnd.n1889 gnd.n1888 0.155672
R11653 gnd.n2809 gnd.n2808 0.152939
R11654 gnd.n2810 gnd.n2809 0.152939
R11655 gnd.n2811 gnd.n2810 0.152939
R11656 gnd.n2812 gnd.n2811 0.152939
R11657 gnd.n2813 gnd.n2812 0.152939
R11658 gnd.n2814 gnd.n2813 0.152939
R11659 gnd.n2815 gnd.n2814 0.152939
R11660 gnd.n2816 gnd.n2815 0.152939
R11661 gnd.n2817 gnd.n2816 0.152939
R11662 gnd.n2818 gnd.n2817 0.152939
R11663 gnd.n2819 gnd.n2818 0.152939
R11664 gnd.n2820 gnd.n2819 0.152939
R11665 gnd.n2821 gnd.n2820 0.152939
R11666 gnd.n2822 gnd.n2821 0.152939
R11667 gnd.n2823 gnd.n2822 0.152939
R11668 gnd.n2824 gnd.n2823 0.152939
R11669 gnd.n2825 gnd.n2824 0.152939
R11670 gnd.n2828 gnd.n2825 0.152939
R11671 gnd.n2829 gnd.n2828 0.152939
R11672 gnd.n2830 gnd.n2829 0.152939
R11673 gnd.n2831 gnd.n2830 0.152939
R11674 gnd.n2832 gnd.n2831 0.152939
R11675 gnd.n2833 gnd.n2832 0.152939
R11676 gnd.n2834 gnd.n2833 0.152939
R11677 gnd.n2835 gnd.n2834 0.152939
R11678 gnd.n2840 gnd.n2839 0.152939
R11679 gnd.n2841 gnd.n2840 0.152939
R11680 gnd.n2842 gnd.n2841 0.152939
R11681 gnd.n2843 gnd.n2842 0.152939
R11682 gnd.n2844 gnd.n2843 0.152939
R11683 gnd.n2845 gnd.n2844 0.152939
R11684 gnd.n2846 gnd.n2845 0.152939
R11685 gnd.n2847 gnd.n2846 0.152939
R11686 gnd.n2848 gnd.n2847 0.152939
R11687 gnd.n2851 gnd.n2848 0.152939
R11688 gnd.n2852 gnd.n2851 0.152939
R11689 gnd.n2853 gnd.n2852 0.152939
R11690 gnd.n2854 gnd.n2853 0.152939
R11691 gnd.n2855 gnd.n2854 0.152939
R11692 gnd.n2856 gnd.n2855 0.152939
R11693 gnd.n2857 gnd.n2856 0.152939
R11694 gnd.n2858 gnd.n2857 0.152939
R11695 gnd.n2859 gnd.n2858 0.152939
R11696 gnd.n2860 gnd.n2859 0.152939
R11697 gnd.n2861 gnd.n2860 0.152939
R11698 gnd.n2862 gnd.n2861 0.152939
R11699 gnd.n2863 gnd.n2862 0.152939
R11700 gnd.n2864 gnd.n2863 0.152939
R11701 gnd.n2865 gnd.n2864 0.152939
R11702 gnd.n2866 gnd.n2865 0.152939
R11703 gnd.n2867 gnd.n2866 0.152939
R11704 gnd.n2868 gnd.n2867 0.152939
R11705 gnd.n2869 gnd.n2868 0.152939
R11706 gnd.n5283 gnd.n2869 0.152939
R11707 gnd.n5283 gnd.n5282 0.152939
R11708 gnd.n5084 gnd.n5080 0.152939
R11709 gnd.n5085 gnd.n5084 0.152939
R11710 gnd.n5086 gnd.n5085 0.152939
R11711 gnd.n5087 gnd.n5086 0.152939
R11712 gnd.n5088 gnd.n5087 0.152939
R11713 gnd.n5089 gnd.n5088 0.152939
R11714 gnd.n5089 gnd.n236 0.152939
R11715 gnd.n6754 gnd.n236 0.152939
R11716 gnd.n6755 gnd.n6754 0.152939
R11717 gnd.n6756 gnd.n6755 0.152939
R11718 gnd.n6757 gnd.n6756 0.152939
R11719 gnd.n6757 gnd.n208 0.152939
R11720 gnd.n6789 gnd.n208 0.152939
R11721 gnd.n6790 gnd.n6789 0.152939
R11722 gnd.n6791 gnd.n6790 0.152939
R11723 gnd.n6792 gnd.n6791 0.152939
R11724 gnd.n99 gnd.n98 0.152939
R11725 gnd.n100 gnd.n99 0.152939
R11726 gnd.n101 gnd.n100 0.152939
R11727 gnd.n118 gnd.n101 0.152939
R11728 gnd.n119 gnd.n118 0.152939
R11729 gnd.n120 gnd.n119 0.152939
R11730 gnd.n121 gnd.n120 0.152939
R11731 gnd.n137 gnd.n121 0.152939
R11732 gnd.n138 gnd.n137 0.152939
R11733 gnd.n139 gnd.n138 0.152939
R11734 gnd.n140 gnd.n139 0.152939
R11735 gnd.n157 gnd.n140 0.152939
R11736 gnd.n158 gnd.n157 0.152939
R11737 gnd.n159 gnd.n158 0.152939
R11738 gnd.n160 gnd.n159 0.152939
R11739 gnd.n7023 gnd.n160 0.152939
R11740 gnd.n7268 gnd.n69 0.152939
R11741 gnd.n6953 gnd.n69 0.152939
R11742 gnd.n6954 gnd.n6953 0.152939
R11743 gnd.n6958 gnd.n6954 0.152939
R11744 gnd.n6959 gnd.n6958 0.152939
R11745 gnd.n6960 gnd.n6959 0.152939
R11746 gnd.n6960 gnd.n6951 0.152939
R11747 gnd.n6966 gnd.n6951 0.152939
R11748 gnd.n6967 gnd.n6966 0.152939
R11749 gnd.n6968 gnd.n6967 0.152939
R11750 gnd.n6968 gnd.n6949 0.152939
R11751 gnd.n6974 gnd.n6949 0.152939
R11752 gnd.n6975 gnd.n6974 0.152939
R11753 gnd.n6976 gnd.n6975 0.152939
R11754 gnd.n6976 gnd.n6947 0.152939
R11755 gnd.n6982 gnd.n6947 0.152939
R11756 gnd.n6983 gnd.n6982 0.152939
R11757 gnd.n6984 gnd.n6983 0.152939
R11758 gnd.n6984 gnd.n6945 0.152939
R11759 gnd.n6989 gnd.n6945 0.152939
R11760 gnd.n6905 gnd.n6875 0.152939
R11761 gnd.n6906 gnd.n6905 0.152939
R11762 gnd.n6906 gnd.n6901 0.152939
R11763 gnd.n6914 gnd.n6901 0.152939
R11764 gnd.n6915 gnd.n6914 0.152939
R11765 gnd.n6916 gnd.n6915 0.152939
R11766 gnd.n6916 gnd.n6899 0.152939
R11767 gnd.n6924 gnd.n6899 0.152939
R11768 gnd.n6925 gnd.n6924 0.152939
R11769 gnd.n6926 gnd.n6925 0.152939
R11770 gnd.n6926 gnd.n6897 0.152939
R11771 gnd.n6934 gnd.n6897 0.152939
R11772 gnd.n6935 gnd.n6934 0.152939
R11773 gnd.n6936 gnd.n6935 0.152939
R11774 gnd.n6936 gnd.n6895 0.152939
R11775 gnd.n6943 gnd.n6895 0.152939
R11776 gnd.n6944 gnd.n6943 0.152939
R11777 gnd.n6990 gnd.n6944 0.152939
R11778 gnd.n7195 gnd.n7024 0.152939
R11779 gnd.n7195 gnd.n7194 0.152939
R11780 gnd.n7194 gnd.n7193 0.152939
R11781 gnd.n7193 gnd.n7026 0.152939
R11782 gnd.n7027 gnd.n7026 0.152939
R11783 gnd.n7028 gnd.n7027 0.152939
R11784 gnd.n7029 gnd.n7028 0.152939
R11785 gnd.n7030 gnd.n7029 0.152939
R11786 gnd.n7031 gnd.n7030 0.152939
R11787 gnd.n7032 gnd.n7031 0.152939
R11788 gnd.n7033 gnd.n7032 0.152939
R11789 gnd.n7034 gnd.n7033 0.152939
R11790 gnd.n7035 gnd.n7034 0.152939
R11791 gnd.n7036 gnd.n7035 0.152939
R11792 gnd.n7037 gnd.n7036 0.152939
R11793 gnd.n7038 gnd.n7037 0.152939
R11794 gnd.n7039 gnd.n7038 0.152939
R11795 gnd.n7040 gnd.n7039 0.152939
R11796 gnd.n7041 gnd.n7040 0.152939
R11797 gnd.n7042 gnd.n7041 0.152939
R11798 gnd.n7043 gnd.n7042 0.152939
R11799 gnd.n7044 gnd.n7043 0.152939
R11800 gnd.n7045 gnd.n7044 0.152939
R11801 gnd.n7046 gnd.n7045 0.152939
R11802 gnd.n7047 gnd.n7046 0.152939
R11803 gnd.n7048 gnd.n7047 0.152939
R11804 gnd.n7049 gnd.n7048 0.152939
R11805 gnd.n7050 gnd.n7049 0.152939
R11806 gnd.n7051 gnd.n7050 0.152939
R11807 gnd.n7052 gnd.n7051 0.152939
R11808 gnd.n7053 gnd.n7052 0.152939
R11809 gnd.n7054 gnd.n7053 0.152939
R11810 gnd.n7055 gnd.n7054 0.152939
R11811 gnd.n7056 gnd.n7055 0.152939
R11812 gnd.n7057 gnd.n7056 0.152939
R11813 gnd.n7058 gnd.n7057 0.152939
R11814 gnd.n7118 gnd.n7058 0.152939
R11815 gnd.n7118 gnd.n7117 0.152939
R11816 gnd.n7117 gnd.n7116 0.152939
R11817 gnd.n7116 gnd.n7062 0.152939
R11818 gnd.n7063 gnd.n7062 0.152939
R11819 gnd.n7064 gnd.n7063 0.152939
R11820 gnd.n7065 gnd.n7064 0.152939
R11821 gnd.n7066 gnd.n7065 0.152939
R11822 gnd.n7067 gnd.n7066 0.152939
R11823 gnd.n7068 gnd.n7067 0.152939
R11824 gnd.n7069 gnd.n7068 0.152939
R11825 gnd.n7070 gnd.n7069 0.152939
R11826 gnd.n7071 gnd.n7070 0.152939
R11827 gnd.n7072 gnd.n7071 0.152939
R11828 gnd.n7073 gnd.n7072 0.152939
R11829 gnd.n7074 gnd.n7073 0.152939
R11830 gnd.n7075 gnd.n7074 0.152939
R11831 gnd.n7076 gnd.n7075 0.152939
R11832 gnd.n7077 gnd.n7076 0.152939
R11833 gnd.n7078 gnd.n7077 0.152939
R11834 gnd.n7078 gnd.n6876 0.152939
R11835 gnd.n7204 gnd.n6876 0.152939
R11836 gnd.n5971 gnd.n5937 0.152939
R11837 gnd.n5971 gnd.n5970 0.152939
R11838 gnd.n5970 gnd.n5969 0.152939
R11839 gnd.n5969 gnd.n5939 0.152939
R11840 gnd.n5940 gnd.n5939 0.152939
R11841 gnd.n5941 gnd.n5940 0.152939
R11842 gnd.n5942 gnd.n5941 0.152939
R11843 gnd.n5943 gnd.n5942 0.152939
R11844 gnd.n5944 gnd.n5943 0.152939
R11845 gnd.n5945 gnd.n5944 0.152939
R11846 gnd.n5946 gnd.n5945 0.152939
R11847 gnd.n5947 gnd.n5946 0.152939
R11848 gnd.n5947 gnd.n787 0.152939
R11849 gnd.n5980 gnd.n787 0.152939
R11850 gnd.n5981 gnd.n5980 0.152939
R11851 gnd.n5982 gnd.n5981 0.152939
R11852 gnd.n1553 gnd.n1552 0.152939
R11853 gnd.n1553 gnd.n1257 0.152939
R11854 gnd.n1581 gnd.n1257 0.152939
R11855 gnd.n1582 gnd.n1581 0.152939
R11856 gnd.n1583 gnd.n1582 0.152939
R11857 gnd.n1584 gnd.n1583 0.152939
R11858 gnd.n1584 gnd.n1229 0.152939
R11859 gnd.n1611 gnd.n1229 0.152939
R11860 gnd.n1612 gnd.n1611 0.152939
R11861 gnd.n1613 gnd.n1612 0.152939
R11862 gnd.n1614 gnd.n1613 0.152939
R11863 gnd.n1615 gnd.n1614 0.152939
R11864 gnd.n1617 gnd.n1615 0.152939
R11865 gnd.n1617 gnd.n1616 0.152939
R11866 gnd.n1616 gnd.n1197 0.152939
R11867 gnd.n1670 gnd.n1197 0.152939
R11868 gnd.n1671 gnd.n1670 0.152939
R11869 gnd.n1672 gnd.n1671 0.152939
R11870 gnd.n1672 gnd.n1032 0.152939
R11871 gnd.n1706 gnd.n1032 0.152939
R11872 gnd.n1707 gnd.n1706 0.152939
R11873 gnd.n1708 gnd.n1707 0.152939
R11874 gnd.n1709 gnd.n1708 0.152939
R11875 gnd.n1709 gnd.n1008 0.152939
R11876 gnd.n1737 gnd.n1008 0.152939
R11877 gnd.n1738 gnd.n1737 0.152939
R11878 gnd.n1739 gnd.n1738 0.152939
R11879 gnd.n1740 gnd.n1739 0.152939
R11880 gnd.n1740 gnd.n982 0.152939
R11881 gnd.n1768 gnd.n982 0.152939
R11882 gnd.n1769 gnd.n1768 0.152939
R11883 gnd.n1770 gnd.n1769 0.152939
R11884 gnd.n1771 gnd.n1770 0.152939
R11885 gnd.n1771 gnd.n957 0.152939
R11886 gnd.n1799 gnd.n957 0.152939
R11887 gnd.n1800 gnd.n1799 0.152939
R11888 gnd.n1801 gnd.n1800 0.152939
R11889 gnd.n1802 gnd.n1801 0.152939
R11890 gnd.n1802 gnd.n932 0.152939
R11891 gnd.n1830 gnd.n932 0.152939
R11892 gnd.n1831 gnd.n1830 0.152939
R11893 gnd.n1832 gnd.n1831 0.152939
R11894 gnd.n1833 gnd.n1832 0.152939
R11895 gnd.n1833 gnd.n906 0.152939
R11896 gnd.n1861 gnd.n906 0.152939
R11897 gnd.n1862 gnd.n1861 0.152939
R11898 gnd.n1863 gnd.n1862 0.152939
R11899 gnd.n1865 gnd.n1863 0.152939
R11900 gnd.n1865 gnd.n1864 0.152939
R11901 gnd.n1864 gnd.n768 0.152939
R11902 gnd.n769 gnd.n768 0.152939
R11903 gnd.n770 gnd.n769 0.152939
R11904 gnd.n5936 gnd.n770 0.152939
R11905 gnd.n1551 gnd.n1281 0.152939
R11906 gnd.n1302 gnd.n1281 0.152939
R11907 gnd.n1303 gnd.n1302 0.152939
R11908 gnd.n1309 gnd.n1303 0.152939
R11909 gnd.n1310 gnd.n1309 0.152939
R11910 gnd.n1311 gnd.n1310 0.152939
R11911 gnd.n1311 gnd.n1300 0.152939
R11912 gnd.n1319 gnd.n1300 0.152939
R11913 gnd.n1320 gnd.n1319 0.152939
R11914 gnd.n1321 gnd.n1320 0.152939
R11915 gnd.n1321 gnd.n1298 0.152939
R11916 gnd.n1329 gnd.n1298 0.152939
R11917 gnd.n1330 gnd.n1329 0.152939
R11918 gnd.n1331 gnd.n1330 0.152939
R11919 gnd.n1331 gnd.n1296 0.152939
R11920 gnd.n1339 gnd.n1296 0.152939
R11921 gnd.n822 gnd.n821 0.152939
R11922 gnd.n823 gnd.n822 0.152939
R11923 gnd.n823 gnd.n817 0.152939
R11924 gnd.n831 gnd.n817 0.152939
R11925 gnd.n832 gnd.n831 0.152939
R11926 gnd.n833 gnd.n832 0.152939
R11927 gnd.n833 gnd.n815 0.152939
R11928 gnd.n841 gnd.n815 0.152939
R11929 gnd.n842 gnd.n841 0.152939
R11930 gnd.n843 gnd.n842 0.152939
R11931 gnd.n843 gnd.n813 0.152939
R11932 gnd.n851 gnd.n813 0.152939
R11933 gnd.n852 gnd.n851 0.152939
R11934 gnd.n853 gnd.n852 0.152939
R11935 gnd.n853 gnd.n811 0.152939
R11936 gnd.n861 gnd.n811 0.152939
R11937 gnd.n862 gnd.n861 0.152939
R11938 gnd.n863 gnd.n862 0.152939
R11939 gnd.n863 gnd.n809 0.152939
R11940 gnd.n871 gnd.n809 0.152939
R11941 gnd.n872 gnd.n871 0.152939
R11942 gnd.n873 gnd.n872 0.152939
R11943 gnd.n873 gnd.n804 0.152939
R11944 gnd.n880 gnd.n804 0.152939
R11945 gnd.n881 gnd.n880 0.152939
R11946 gnd.n2151 gnd.n881 0.152939
R11947 gnd.n1050 gnd.n1049 0.152939
R11948 gnd.n1051 gnd.n1050 0.152939
R11949 gnd.n1052 gnd.n1051 0.152939
R11950 gnd.n1053 gnd.n1052 0.152939
R11951 gnd.n1054 gnd.n1053 0.152939
R11952 gnd.n1055 gnd.n1054 0.152939
R11953 gnd.n1056 gnd.n1055 0.152939
R11954 gnd.n1057 gnd.n1056 0.152939
R11955 gnd.n1058 gnd.n1057 0.152939
R11956 gnd.n1059 gnd.n1058 0.152939
R11957 gnd.n1060 gnd.n1059 0.152939
R11958 gnd.n1061 gnd.n1060 0.152939
R11959 gnd.n1062 gnd.n1061 0.152939
R11960 gnd.n1063 gnd.n1062 0.152939
R11961 gnd.n1064 gnd.n1063 0.152939
R11962 gnd.n1065 gnd.n1064 0.152939
R11963 gnd.n1066 gnd.n1065 0.152939
R11964 gnd.n1067 gnd.n1066 0.152939
R11965 gnd.n1068 gnd.n1067 0.152939
R11966 gnd.n1069 gnd.n1068 0.152939
R11967 gnd.n1070 gnd.n1069 0.152939
R11968 gnd.n1071 gnd.n1070 0.152939
R11969 gnd.n1072 gnd.n1071 0.152939
R11970 gnd.n1073 gnd.n1072 0.152939
R11971 gnd.n1075 gnd.n1073 0.152939
R11972 gnd.n1075 gnd.n1074 0.152939
R11973 gnd.n1074 gnd.n882 0.152939
R11974 gnd.n2150 gnd.n882 0.152939
R11975 gnd.n1469 gnd.n1468 0.152939
R11976 gnd.n1469 gnd.n1359 0.152939
R11977 gnd.n1484 gnd.n1359 0.152939
R11978 gnd.n1485 gnd.n1484 0.152939
R11979 gnd.n1486 gnd.n1485 0.152939
R11980 gnd.n1486 gnd.n1347 0.152939
R11981 gnd.n1500 gnd.n1347 0.152939
R11982 gnd.n1501 gnd.n1500 0.152939
R11983 gnd.n1502 gnd.n1501 0.152939
R11984 gnd.n1503 gnd.n1502 0.152939
R11985 gnd.n1504 gnd.n1503 0.152939
R11986 gnd.n1505 gnd.n1504 0.152939
R11987 gnd.n1506 gnd.n1505 0.152939
R11988 gnd.n1507 gnd.n1506 0.152939
R11989 gnd.n1508 gnd.n1507 0.152939
R11990 gnd.n1509 gnd.n1508 0.152939
R11991 gnd.n1510 gnd.n1509 0.152939
R11992 gnd.n1511 gnd.n1510 0.152939
R11993 gnd.n1512 gnd.n1511 0.152939
R11994 gnd.n1513 gnd.n1512 0.152939
R11995 gnd.n1514 gnd.n1513 0.152939
R11996 gnd.n1514 gnd.n1212 0.152939
R11997 gnd.n1637 gnd.n1212 0.152939
R11998 gnd.n1638 gnd.n1637 0.152939
R11999 gnd.n1639 gnd.n1638 0.152939
R12000 gnd.n1640 gnd.n1639 0.152939
R12001 gnd.n1640 gnd.n1175 0.152939
R12002 gnd.n1685 gnd.n1175 0.152939
R12003 gnd.n1387 gnd.n1386 0.152939
R12004 gnd.n1388 gnd.n1387 0.152939
R12005 gnd.n1389 gnd.n1388 0.152939
R12006 gnd.n1390 gnd.n1389 0.152939
R12007 gnd.n1391 gnd.n1390 0.152939
R12008 gnd.n1392 gnd.n1391 0.152939
R12009 gnd.n1393 gnd.n1392 0.152939
R12010 gnd.n1394 gnd.n1393 0.152939
R12011 gnd.n1395 gnd.n1394 0.152939
R12012 gnd.n1396 gnd.n1395 0.152939
R12013 gnd.n1397 gnd.n1396 0.152939
R12014 gnd.n1398 gnd.n1397 0.152939
R12015 gnd.n1399 gnd.n1398 0.152939
R12016 gnd.n1400 gnd.n1399 0.152939
R12017 gnd.n1401 gnd.n1400 0.152939
R12018 gnd.n1402 gnd.n1401 0.152939
R12019 gnd.n1403 gnd.n1402 0.152939
R12020 gnd.n1404 gnd.n1403 0.152939
R12021 gnd.n1405 gnd.n1404 0.152939
R12022 gnd.n1406 gnd.n1405 0.152939
R12023 gnd.n1407 gnd.n1406 0.152939
R12024 gnd.n1408 gnd.n1407 0.152939
R12025 gnd.n1412 gnd.n1408 0.152939
R12026 gnd.n1413 gnd.n1412 0.152939
R12027 gnd.n1413 gnd.n1370 0.152939
R12028 gnd.n1467 gnd.n1370 0.152939
R12029 gnd.n3730 gnd.n3729 0.152939
R12030 gnd.n3731 gnd.n3730 0.152939
R12031 gnd.n3731 gnd.n3669 0.152939
R12032 gnd.n3737 gnd.n3669 0.152939
R12033 gnd.n3738 gnd.n3737 0.152939
R12034 gnd.n3739 gnd.n3738 0.152939
R12035 gnd.n3739 gnd.n3667 0.152939
R12036 gnd.n3745 gnd.n3667 0.152939
R12037 gnd.n3746 gnd.n3745 0.152939
R12038 gnd.n3747 gnd.n3746 0.152939
R12039 gnd.n3747 gnd.n3665 0.152939
R12040 gnd.n3753 gnd.n3665 0.152939
R12041 gnd.n3754 gnd.n3753 0.152939
R12042 gnd.n3755 gnd.n3754 0.152939
R12043 gnd.n3755 gnd.n3663 0.152939
R12044 gnd.n3761 gnd.n3663 0.152939
R12045 gnd.n3762 gnd.n3761 0.152939
R12046 gnd.n3763 gnd.n3762 0.152939
R12047 gnd.n3763 gnd.n3661 0.152939
R12048 gnd.n3769 gnd.n3661 0.152939
R12049 gnd.n5677 gnd.n2471 0.152939
R12050 gnd.n2515 gnd.n2471 0.152939
R12051 gnd.n2516 gnd.n2515 0.152939
R12052 gnd.n2517 gnd.n2516 0.152939
R12053 gnd.n2518 gnd.n2517 0.152939
R12054 gnd.n2519 gnd.n2518 0.152939
R12055 gnd.n2520 gnd.n2519 0.152939
R12056 gnd.n2521 gnd.n2520 0.152939
R12057 gnd.n2522 gnd.n2521 0.152939
R12058 gnd.n2523 gnd.n2522 0.152939
R12059 gnd.n2524 gnd.n2523 0.152939
R12060 gnd.n2525 gnd.n2524 0.152939
R12061 gnd.n2526 gnd.n2525 0.152939
R12062 gnd.n2527 gnd.n2526 0.152939
R12063 gnd.n2528 gnd.n2527 0.152939
R12064 gnd.n2529 gnd.n2528 0.152939
R12065 gnd.n2530 gnd.n2529 0.152939
R12066 gnd.n2533 gnd.n2530 0.152939
R12067 gnd.n2534 gnd.n2533 0.152939
R12068 gnd.n2535 gnd.n2534 0.152939
R12069 gnd.n2536 gnd.n2535 0.152939
R12070 gnd.n2537 gnd.n2536 0.152939
R12071 gnd.n2538 gnd.n2537 0.152939
R12072 gnd.n2539 gnd.n2538 0.152939
R12073 gnd.n2540 gnd.n2539 0.152939
R12074 gnd.n3543 gnd.n3542 0.152939
R12075 gnd.n3544 gnd.n3543 0.152939
R12076 gnd.n3544 gnd.n3538 0.152939
R12077 gnd.n3552 gnd.n3538 0.152939
R12078 gnd.n3553 gnd.n3552 0.152939
R12079 gnd.n3554 gnd.n3553 0.152939
R12080 gnd.n3554 gnd.n3536 0.152939
R12081 gnd.n3562 gnd.n3536 0.152939
R12082 gnd.n3563 gnd.n3562 0.152939
R12083 gnd.n3564 gnd.n3563 0.152939
R12084 gnd.n3564 gnd.n3532 0.152939
R12085 gnd.n3572 gnd.n3532 0.152939
R12086 gnd.n3573 gnd.n3572 0.152939
R12087 gnd.n3574 gnd.n3573 0.152939
R12088 gnd.n3574 gnd.n3530 0.152939
R12089 gnd.n3582 gnd.n3530 0.152939
R12090 gnd.n3583 gnd.n3582 0.152939
R12091 gnd.n3584 gnd.n3583 0.152939
R12092 gnd.n3584 gnd.n3528 0.152939
R12093 gnd.n3592 gnd.n3528 0.152939
R12094 gnd.n3593 gnd.n3592 0.152939
R12095 gnd.n3594 gnd.n3593 0.152939
R12096 gnd.n3594 gnd.n3526 0.152939
R12097 gnd.n3602 gnd.n3526 0.152939
R12098 gnd.n3603 gnd.n3602 0.152939
R12099 gnd.n3604 gnd.n3603 0.152939
R12100 gnd.n3604 gnd.n3524 0.152939
R12101 gnd.n3612 gnd.n3524 0.152939
R12102 gnd.n3613 gnd.n3612 0.152939
R12103 gnd.n3614 gnd.n3613 0.152939
R12104 gnd.n2390 gnd.n2389 0.152939
R12105 gnd.n2407 gnd.n2390 0.152939
R12106 gnd.n2408 gnd.n2407 0.152939
R12107 gnd.n2409 gnd.n2408 0.152939
R12108 gnd.n2410 gnd.n2409 0.152939
R12109 gnd.n2427 gnd.n2410 0.152939
R12110 gnd.n2428 gnd.n2427 0.152939
R12111 gnd.n2429 gnd.n2428 0.152939
R12112 gnd.n2430 gnd.n2429 0.152939
R12113 gnd.n2448 gnd.n2430 0.152939
R12114 gnd.n2449 gnd.n2448 0.152939
R12115 gnd.n2450 gnd.n2449 0.152939
R12116 gnd.n2451 gnd.n2450 0.152939
R12117 gnd.n2469 gnd.n2451 0.152939
R12118 gnd.n2470 gnd.n2469 0.152939
R12119 gnd.n5678 gnd.n2470 0.152939
R12120 gnd.n5801 gnd.n2274 0.152939
R12121 gnd.n5801 gnd.n5800 0.152939
R12122 gnd.n5800 gnd.n5799 0.152939
R12123 gnd.n5799 gnd.n2275 0.152939
R12124 gnd.n2293 gnd.n2275 0.152939
R12125 gnd.n2294 gnd.n2293 0.152939
R12126 gnd.n2295 gnd.n2294 0.152939
R12127 gnd.n2310 gnd.n2295 0.152939
R12128 gnd.n2311 gnd.n2310 0.152939
R12129 gnd.n2312 gnd.n2311 0.152939
R12130 gnd.n2313 gnd.n2312 0.152939
R12131 gnd.n2330 gnd.n2313 0.152939
R12132 gnd.n2331 gnd.n2330 0.152939
R12133 gnd.n2332 gnd.n2331 0.152939
R12134 gnd.n2333 gnd.n2332 0.152939
R12135 gnd.n2348 gnd.n2333 0.152939
R12136 gnd.n2198 gnd.n2197 0.152939
R12137 gnd.n2199 gnd.n2198 0.152939
R12138 gnd.n2200 gnd.n2199 0.152939
R12139 gnd.n2201 gnd.n2200 0.152939
R12140 gnd.n2202 gnd.n2201 0.152939
R12141 gnd.n2203 gnd.n2202 0.152939
R12142 gnd.n2204 gnd.n2203 0.152939
R12143 gnd.n2205 gnd.n2204 0.152939
R12144 gnd.n2206 gnd.n2205 0.152939
R12145 gnd.n2207 gnd.n2206 0.152939
R12146 gnd.n2208 gnd.n2207 0.152939
R12147 gnd.n2209 gnd.n2208 0.152939
R12148 gnd.n2210 gnd.n2209 0.152939
R12149 gnd.n2211 gnd.n2210 0.152939
R12150 gnd.n2212 gnd.n2211 0.152939
R12151 gnd.n2213 gnd.n2212 0.152939
R12152 gnd.n2214 gnd.n2213 0.152939
R12153 gnd.n2217 gnd.n2214 0.152939
R12154 gnd.n2218 gnd.n2217 0.152939
R12155 gnd.n2219 gnd.n2218 0.152939
R12156 gnd.n2220 gnd.n2219 0.152939
R12157 gnd.n2221 gnd.n2220 0.152939
R12158 gnd.n2222 gnd.n2221 0.152939
R12159 gnd.n2223 gnd.n2222 0.152939
R12160 gnd.n2224 gnd.n2223 0.152939
R12161 gnd.n2225 gnd.n2224 0.152939
R12162 gnd.n2226 gnd.n2225 0.152939
R12163 gnd.n2227 gnd.n2226 0.152939
R12164 gnd.n2228 gnd.n2227 0.152939
R12165 gnd.n2229 gnd.n2228 0.152939
R12166 gnd.n2230 gnd.n2229 0.152939
R12167 gnd.n2231 gnd.n2230 0.152939
R12168 gnd.n2232 gnd.n2231 0.152939
R12169 gnd.n2233 gnd.n2232 0.152939
R12170 gnd.n2234 gnd.n2233 0.152939
R12171 gnd.n2235 gnd.n2234 0.152939
R12172 gnd.n2236 gnd.n2235 0.152939
R12173 gnd.n2239 gnd.n2236 0.152939
R12174 gnd.n2240 gnd.n2239 0.152939
R12175 gnd.n2241 gnd.n2240 0.152939
R12176 gnd.n2242 gnd.n2241 0.152939
R12177 gnd.n2243 gnd.n2242 0.152939
R12178 gnd.n2244 gnd.n2243 0.152939
R12179 gnd.n2245 gnd.n2244 0.152939
R12180 gnd.n2246 gnd.n2245 0.152939
R12181 gnd.n2247 gnd.n2246 0.152939
R12182 gnd.n2248 gnd.n2247 0.152939
R12183 gnd.n2249 gnd.n2248 0.152939
R12184 gnd.n2250 gnd.n2249 0.152939
R12185 gnd.n2251 gnd.n2250 0.152939
R12186 gnd.n2252 gnd.n2251 0.152939
R12187 gnd.n2253 gnd.n2252 0.152939
R12188 gnd.n2254 gnd.n2253 0.152939
R12189 gnd.n2255 gnd.n2254 0.152939
R12190 gnd.n2256 gnd.n2255 0.152939
R12191 gnd.n2257 gnd.n2256 0.152939
R12192 gnd.n5811 gnd.n2257 0.152939
R12193 gnd.n5811 gnd.n5810 0.152939
R12194 gnd.n3684 gnd.n2261 0.152939
R12195 gnd.n3690 gnd.n3684 0.152939
R12196 gnd.n3691 gnd.n3690 0.152939
R12197 gnd.n3692 gnd.n3691 0.152939
R12198 gnd.n3692 gnd.n3682 0.152939
R12199 gnd.n3700 gnd.n3682 0.152939
R12200 gnd.n3701 gnd.n3700 0.152939
R12201 gnd.n3702 gnd.n3701 0.152939
R12202 gnd.n3702 gnd.n3680 0.152939
R12203 gnd.n3710 gnd.n3680 0.152939
R12204 gnd.n3711 gnd.n3710 0.152939
R12205 gnd.n3712 gnd.n3711 0.152939
R12206 gnd.n3712 gnd.n3678 0.152939
R12207 gnd.n3720 gnd.n3678 0.152939
R12208 gnd.n3721 gnd.n3720 0.152939
R12209 gnd.n3722 gnd.n3721 0.152939
R12210 gnd.n3722 gnd.n3671 0.152939
R12211 gnd.n3726 gnd.n3671 0.152939
R12212 gnd.n6172 gnd.n6171 0.152939
R12213 gnd.n6173 gnd.n6172 0.152939
R12214 gnd.n6173 gnd.n587 0.152939
R12215 gnd.n6181 gnd.n587 0.152939
R12216 gnd.n6182 gnd.n6181 0.152939
R12217 gnd.n6183 gnd.n6182 0.152939
R12218 gnd.n6183 gnd.n581 0.152939
R12219 gnd.n6191 gnd.n581 0.152939
R12220 gnd.n6192 gnd.n6191 0.152939
R12221 gnd.n6193 gnd.n6192 0.152939
R12222 gnd.n6193 gnd.n575 0.152939
R12223 gnd.n6201 gnd.n575 0.152939
R12224 gnd.n6202 gnd.n6201 0.152939
R12225 gnd.n6203 gnd.n6202 0.152939
R12226 gnd.n6203 gnd.n569 0.152939
R12227 gnd.n6211 gnd.n569 0.152939
R12228 gnd.n6212 gnd.n6211 0.152939
R12229 gnd.n6213 gnd.n6212 0.152939
R12230 gnd.n6213 gnd.n563 0.152939
R12231 gnd.n6221 gnd.n563 0.152939
R12232 gnd.n6222 gnd.n6221 0.152939
R12233 gnd.n6223 gnd.n6222 0.152939
R12234 gnd.n6223 gnd.n557 0.152939
R12235 gnd.n6231 gnd.n557 0.152939
R12236 gnd.n6232 gnd.n6231 0.152939
R12237 gnd.n6233 gnd.n6232 0.152939
R12238 gnd.n6233 gnd.n551 0.152939
R12239 gnd.n6241 gnd.n551 0.152939
R12240 gnd.n6242 gnd.n6241 0.152939
R12241 gnd.n6243 gnd.n6242 0.152939
R12242 gnd.n6243 gnd.n545 0.152939
R12243 gnd.n6251 gnd.n545 0.152939
R12244 gnd.n6252 gnd.n6251 0.152939
R12245 gnd.n6253 gnd.n6252 0.152939
R12246 gnd.n6253 gnd.n539 0.152939
R12247 gnd.n6261 gnd.n539 0.152939
R12248 gnd.n6262 gnd.n6261 0.152939
R12249 gnd.n6263 gnd.n6262 0.152939
R12250 gnd.n6263 gnd.n533 0.152939
R12251 gnd.n6271 gnd.n533 0.152939
R12252 gnd.n6272 gnd.n6271 0.152939
R12253 gnd.n6273 gnd.n6272 0.152939
R12254 gnd.n6273 gnd.n527 0.152939
R12255 gnd.n6281 gnd.n527 0.152939
R12256 gnd.n6282 gnd.n6281 0.152939
R12257 gnd.n6283 gnd.n6282 0.152939
R12258 gnd.n6283 gnd.n521 0.152939
R12259 gnd.n6291 gnd.n521 0.152939
R12260 gnd.n6292 gnd.n6291 0.152939
R12261 gnd.n6293 gnd.n6292 0.152939
R12262 gnd.n6293 gnd.n515 0.152939
R12263 gnd.n6301 gnd.n515 0.152939
R12264 gnd.n6302 gnd.n6301 0.152939
R12265 gnd.n6303 gnd.n6302 0.152939
R12266 gnd.n6303 gnd.n509 0.152939
R12267 gnd.n6311 gnd.n509 0.152939
R12268 gnd.n6312 gnd.n6311 0.152939
R12269 gnd.n6313 gnd.n6312 0.152939
R12270 gnd.n6313 gnd.n503 0.152939
R12271 gnd.n6321 gnd.n503 0.152939
R12272 gnd.n6322 gnd.n6321 0.152939
R12273 gnd.n6323 gnd.n6322 0.152939
R12274 gnd.n6323 gnd.n497 0.152939
R12275 gnd.n6331 gnd.n497 0.152939
R12276 gnd.n6332 gnd.n6331 0.152939
R12277 gnd.n6333 gnd.n6332 0.152939
R12278 gnd.n6333 gnd.n491 0.152939
R12279 gnd.n6341 gnd.n491 0.152939
R12280 gnd.n6342 gnd.n6341 0.152939
R12281 gnd.n6343 gnd.n6342 0.152939
R12282 gnd.n6343 gnd.n485 0.152939
R12283 gnd.n6351 gnd.n485 0.152939
R12284 gnd.n6352 gnd.n6351 0.152939
R12285 gnd.n6353 gnd.n6352 0.152939
R12286 gnd.n6353 gnd.n479 0.152939
R12287 gnd.n6361 gnd.n479 0.152939
R12288 gnd.n6362 gnd.n6361 0.152939
R12289 gnd.n6363 gnd.n6362 0.152939
R12290 gnd.n6363 gnd.n473 0.152939
R12291 gnd.n6371 gnd.n473 0.152939
R12292 gnd.n6372 gnd.n6371 0.152939
R12293 gnd.n6373 gnd.n6372 0.152939
R12294 gnd.n6373 gnd.n467 0.152939
R12295 gnd.n6381 gnd.n467 0.152939
R12296 gnd.n6382 gnd.n6381 0.152939
R12297 gnd.n6383 gnd.n6382 0.152939
R12298 gnd.n6383 gnd.n461 0.152939
R12299 gnd.n6391 gnd.n461 0.152939
R12300 gnd.n6392 gnd.n6391 0.152939
R12301 gnd.n6393 gnd.n6392 0.152939
R12302 gnd.n6393 gnd.n455 0.152939
R12303 gnd.n6401 gnd.n455 0.152939
R12304 gnd.n6402 gnd.n6401 0.152939
R12305 gnd.n6403 gnd.n6402 0.152939
R12306 gnd.n6403 gnd.n449 0.152939
R12307 gnd.n6411 gnd.n449 0.152939
R12308 gnd.n6412 gnd.n6411 0.152939
R12309 gnd.n6413 gnd.n6412 0.152939
R12310 gnd.n6413 gnd.n443 0.152939
R12311 gnd.n6421 gnd.n443 0.152939
R12312 gnd.n6422 gnd.n6421 0.152939
R12313 gnd.n6423 gnd.n6422 0.152939
R12314 gnd.n6423 gnd.n437 0.152939
R12315 gnd.n6431 gnd.n437 0.152939
R12316 gnd.n6432 gnd.n6431 0.152939
R12317 gnd.n6433 gnd.n6432 0.152939
R12318 gnd.n6433 gnd.n431 0.152939
R12319 gnd.n6441 gnd.n431 0.152939
R12320 gnd.n6442 gnd.n6441 0.152939
R12321 gnd.n6443 gnd.n6442 0.152939
R12322 gnd.n6443 gnd.n425 0.152939
R12323 gnd.n6451 gnd.n425 0.152939
R12324 gnd.n6452 gnd.n6451 0.152939
R12325 gnd.n6453 gnd.n6452 0.152939
R12326 gnd.n6453 gnd.n419 0.152939
R12327 gnd.n6461 gnd.n419 0.152939
R12328 gnd.n6462 gnd.n6461 0.152939
R12329 gnd.n6463 gnd.n6462 0.152939
R12330 gnd.n6463 gnd.n413 0.152939
R12331 gnd.n6471 gnd.n413 0.152939
R12332 gnd.n6472 gnd.n6471 0.152939
R12333 gnd.n6473 gnd.n6472 0.152939
R12334 gnd.n6473 gnd.n407 0.152939
R12335 gnd.n6481 gnd.n407 0.152939
R12336 gnd.n6482 gnd.n6481 0.152939
R12337 gnd.n6483 gnd.n6482 0.152939
R12338 gnd.n6483 gnd.n401 0.152939
R12339 gnd.n6491 gnd.n401 0.152939
R12340 gnd.n6492 gnd.n6491 0.152939
R12341 gnd.n6493 gnd.n6492 0.152939
R12342 gnd.n6493 gnd.n395 0.152939
R12343 gnd.n6501 gnd.n395 0.152939
R12344 gnd.n6502 gnd.n6501 0.152939
R12345 gnd.n6503 gnd.n6502 0.152939
R12346 gnd.n6503 gnd.n389 0.152939
R12347 gnd.n6511 gnd.n389 0.152939
R12348 gnd.n6512 gnd.n6511 0.152939
R12349 gnd.n6514 gnd.n6512 0.152939
R12350 gnd.n6514 gnd.n6513 0.152939
R12351 gnd.n6513 gnd.n383 0.152939
R12352 gnd.n6523 gnd.n383 0.152939
R12353 gnd.n6524 gnd.n378 0.152939
R12354 gnd.n6532 gnd.n378 0.152939
R12355 gnd.n6533 gnd.n6532 0.152939
R12356 gnd.n6534 gnd.n6533 0.152939
R12357 gnd.n6534 gnd.n372 0.152939
R12358 gnd.n6542 gnd.n372 0.152939
R12359 gnd.n6543 gnd.n6542 0.152939
R12360 gnd.n6544 gnd.n6543 0.152939
R12361 gnd.n6544 gnd.n366 0.152939
R12362 gnd.n6552 gnd.n366 0.152939
R12363 gnd.n6553 gnd.n6552 0.152939
R12364 gnd.n6554 gnd.n6553 0.152939
R12365 gnd.n6554 gnd.n360 0.152939
R12366 gnd.n6562 gnd.n360 0.152939
R12367 gnd.n6563 gnd.n6562 0.152939
R12368 gnd.n6564 gnd.n6563 0.152939
R12369 gnd.n6564 gnd.n354 0.152939
R12370 gnd.n6572 gnd.n354 0.152939
R12371 gnd.n6573 gnd.n6572 0.152939
R12372 gnd.n6574 gnd.n6573 0.152939
R12373 gnd.n6574 gnd.n348 0.152939
R12374 gnd.n6582 gnd.n348 0.152939
R12375 gnd.n6583 gnd.n6582 0.152939
R12376 gnd.n6584 gnd.n6583 0.152939
R12377 gnd.n6584 gnd.n342 0.152939
R12378 gnd.n6592 gnd.n342 0.152939
R12379 gnd.n6593 gnd.n6592 0.152939
R12380 gnd.n6594 gnd.n6593 0.152939
R12381 gnd.n6594 gnd.n336 0.152939
R12382 gnd.n6602 gnd.n336 0.152939
R12383 gnd.n6603 gnd.n6602 0.152939
R12384 gnd.n6604 gnd.n6603 0.152939
R12385 gnd.n6604 gnd.n330 0.152939
R12386 gnd.n6612 gnd.n330 0.152939
R12387 gnd.n6613 gnd.n6612 0.152939
R12388 gnd.n6614 gnd.n6613 0.152939
R12389 gnd.n6614 gnd.n324 0.152939
R12390 gnd.n6622 gnd.n324 0.152939
R12391 gnd.n6623 gnd.n6622 0.152939
R12392 gnd.n6624 gnd.n6623 0.152939
R12393 gnd.n6624 gnd.n318 0.152939
R12394 gnd.n6632 gnd.n318 0.152939
R12395 gnd.n6633 gnd.n6632 0.152939
R12396 gnd.n6634 gnd.n6633 0.152939
R12397 gnd.n6634 gnd.n312 0.152939
R12398 gnd.n6642 gnd.n312 0.152939
R12399 gnd.n6643 gnd.n6642 0.152939
R12400 gnd.n6644 gnd.n6643 0.152939
R12401 gnd.n6644 gnd.n306 0.152939
R12402 gnd.n6652 gnd.n306 0.152939
R12403 gnd.n6653 gnd.n6652 0.152939
R12404 gnd.n6654 gnd.n6653 0.152939
R12405 gnd.n6654 gnd.n300 0.152939
R12406 gnd.n6662 gnd.n300 0.152939
R12407 gnd.n6663 gnd.n6662 0.152939
R12408 gnd.n6664 gnd.n6663 0.152939
R12409 gnd.n6664 gnd.n294 0.152939
R12410 gnd.n6672 gnd.n294 0.152939
R12411 gnd.n6673 gnd.n6672 0.152939
R12412 gnd.n6674 gnd.n6673 0.152939
R12413 gnd.n6674 gnd.n288 0.152939
R12414 gnd.n6682 gnd.n288 0.152939
R12415 gnd.n6683 gnd.n6682 0.152939
R12416 gnd.n6684 gnd.n6683 0.152939
R12417 gnd.n6684 gnd.n282 0.152939
R12418 gnd.n6692 gnd.n282 0.152939
R12419 gnd.n6693 gnd.n6692 0.152939
R12420 gnd.n6694 gnd.n6693 0.152939
R12421 gnd.n6694 gnd.n276 0.152939
R12422 gnd.n6702 gnd.n276 0.152939
R12423 gnd.n6703 gnd.n6702 0.152939
R12424 gnd.n6704 gnd.n6703 0.152939
R12425 gnd.n6704 gnd.n270 0.152939
R12426 gnd.n6712 gnd.n270 0.152939
R12427 gnd.n6713 gnd.n6712 0.152939
R12428 gnd.n6714 gnd.n6713 0.152939
R12429 gnd.n6714 gnd.n264 0.152939
R12430 gnd.n6722 gnd.n264 0.152939
R12431 gnd.n6723 gnd.n6722 0.152939
R12432 gnd.n6724 gnd.n6723 0.152939
R12433 gnd.n6724 gnd.n258 0.152939
R12434 gnd.n6733 gnd.n258 0.152939
R12435 gnd.n6734 gnd.n6733 0.152939
R12436 gnd.n6735 gnd.n6734 0.152939
R12437 gnd.n3637 gnd.n3636 0.152939
R12438 gnd.n3638 gnd.n3637 0.152939
R12439 gnd.n3638 gnd.n3629 0.152939
R12440 gnd.n3887 gnd.n3629 0.152939
R12441 gnd.n3888 gnd.n3887 0.152939
R12442 gnd.n3889 gnd.n3888 0.152939
R12443 gnd.n3889 gnd.n3625 0.152939
R12444 gnd.n3895 gnd.n3625 0.152939
R12445 gnd.n3896 gnd.n3895 0.152939
R12446 gnd.n3897 gnd.n3896 0.152939
R12447 gnd.n3897 gnd.n3621 0.152939
R12448 gnd.n3903 gnd.n3621 0.152939
R12449 gnd.n3904 gnd.n3903 0.152939
R12450 gnd.n3905 gnd.n3904 0.152939
R12451 gnd.n3906 gnd.n3905 0.152939
R12452 gnd.n3907 gnd.n3906 0.152939
R12453 gnd.n3910 gnd.n3907 0.152939
R12454 gnd.n3911 gnd.n3910 0.152939
R12455 gnd.n3912 gnd.n3911 0.152939
R12456 gnd.n3912 gnd.n3388 0.152939
R12457 gnd.n4001 gnd.n3388 0.152939
R12458 gnd.n4002 gnd.n4001 0.152939
R12459 gnd.n4003 gnd.n4002 0.152939
R12460 gnd.n4003 gnd.n3373 0.152939
R12461 gnd.n4017 gnd.n3373 0.152939
R12462 gnd.n4018 gnd.n4017 0.152939
R12463 gnd.n4019 gnd.n4018 0.152939
R12464 gnd.n4019 gnd.n3358 0.152939
R12465 gnd.n4045 gnd.n3358 0.152939
R12466 gnd.n4046 gnd.n4045 0.152939
R12467 gnd.n4047 gnd.n4046 0.152939
R12468 gnd.n4049 gnd.n4047 0.152939
R12469 gnd.n4049 gnd.n4048 0.152939
R12470 gnd.n4048 gnd.n2612 0.152939
R12471 gnd.n2613 gnd.n2612 0.152939
R12472 gnd.n2614 gnd.n2613 0.152939
R12473 gnd.n3334 gnd.n2614 0.152939
R12474 gnd.n3335 gnd.n3334 0.152939
R12475 gnd.n3335 gnd.n3317 0.152939
R12476 gnd.n4194 gnd.n3317 0.152939
R12477 gnd.n4195 gnd.n4194 0.152939
R12478 gnd.n4196 gnd.n4195 0.152939
R12479 gnd.n4197 gnd.n4196 0.152939
R12480 gnd.n4198 gnd.n4197 0.152939
R12481 gnd.n4198 gnd.n3287 0.152939
R12482 gnd.n4263 gnd.n3287 0.152939
R12483 gnd.n4264 gnd.n4263 0.152939
R12484 gnd.n4265 gnd.n4264 0.152939
R12485 gnd.n4265 gnd.n3270 0.152939
R12486 gnd.n4292 gnd.n3270 0.152939
R12487 gnd.n4293 gnd.n4292 0.152939
R12488 gnd.n4294 gnd.n4293 0.152939
R12489 gnd.n4295 gnd.n4294 0.152939
R12490 gnd.n4295 gnd.n3242 0.152939
R12491 gnd.n4366 gnd.n3242 0.152939
R12492 gnd.n4367 gnd.n4366 0.152939
R12493 gnd.n4368 gnd.n4367 0.152939
R12494 gnd.n4369 gnd.n4368 0.152939
R12495 gnd.n4369 gnd.n3219 0.152939
R12496 gnd.n4398 gnd.n3219 0.152939
R12497 gnd.n4399 gnd.n4398 0.152939
R12498 gnd.n4400 gnd.n4399 0.152939
R12499 gnd.n4401 gnd.n4400 0.152939
R12500 gnd.n4401 gnd.n3198 0.152939
R12501 gnd.n4439 gnd.n3198 0.152939
R12502 gnd.n4440 gnd.n4439 0.152939
R12503 gnd.n4441 gnd.n4440 0.152939
R12504 gnd.n4442 gnd.n4441 0.152939
R12505 gnd.n4442 gnd.n3169 0.152939
R12506 gnd.n4508 gnd.n3169 0.152939
R12507 gnd.n4509 gnd.n4508 0.152939
R12508 gnd.n4510 gnd.n4509 0.152939
R12509 gnd.n4511 gnd.n4510 0.152939
R12510 gnd.n4511 gnd.n3144 0.152939
R12511 gnd.n4540 gnd.n3144 0.152939
R12512 gnd.n4541 gnd.n4540 0.152939
R12513 gnd.n4542 gnd.n4541 0.152939
R12514 gnd.n4543 gnd.n4542 0.152939
R12515 gnd.n4543 gnd.n3121 0.152939
R12516 gnd.n4580 gnd.n3121 0.152939
R12517 gnd.n4581 gnd.n4580 0.152939
R12518 gnd.n4582 gnd.n4581 0.152939
R12519 gnd.n4583 gnd.n4582 0.152939
R12520 gnd.n4583 gnd.n3092 0.152939
R12521 gnd.n4634 gnd.n3092 0.152939
R12522 gnd.n4635 gnd.n4634 0.152939
R12523 gnd.n4636 gnd.n4635 0.152939
R12524 gnd.n4637 gnd.n4636 0.152939
R12525 gnd.n4637 gnd.n3068 0.152939
R12526 gnd.n4676 gnd.n3068 0.152939
R12527 gnd.n4677 gnd.n4676 0.152939
R12528 gnd.n4678 gnd.n4677 0.152939
R12529 gnd.n4679 gnd.n4678 0.152939
R12530 gnd.n4679 gnd.n3040 0.152939
R12531 gnd.n4719 gnd.n3040 0.152939
R12532 gnd.n4720 gnd.n4719 0.152939
R12533 gnd.n4722 gnd.n4720 0.152939
R12534 gnd.n4722 gnd.n4721 0.152939
R12535 gnd.n4721 gnd.n3019 0.152939
R12536 gnd.n3020 gnd.n3019 0.152939
R12537 gnd.n3021 gnd.n3020 0.152939
R12538 gnd.n3023 gnd.n3021 0.152939
R12539 gnd.n3024 gnd.n3023 0.152939
R12540 gnd.n3024 gnd.n2986 0.152939
R12541 gnd.n4811 gnd.n2986 0.152939
R12542 gnd.n4812 gnd.n4811 0.152939
R12543 gnd.n4813 gnd.n4812 0.152939
R12544 gnd.n4813 gnd.n2934 0.152939
R12545 gnd.n4983 gnd.n2934 0.152939
R12546 gnd.n4984 gnd.n4983 0.152939
R12547 gnd.n4985 gnd.n4984 0.152939
R12548 gnd.n4985 gnd.n2922 0.152939
R12549 gnd.n5001 gnd.n2922 0.152939
R12550 gnd.n5002 gnd.n5001 0.152939
R12551 gnd.n5003 gnd.n5002 0.152939
R12552 gnd.n5003 gnd.n2911 0.152939
R12553 gnd.n5018 gnd.n2911 0.152939
R12554 gnd.n5019 gnd.n5018 0.152939
R12555 gnd.n5020 gnd.n5019 0.152939
R12556 gnd.n5021 gnd.n5020 0.152939
R12557 gnd.n5021 gnd.n2898 0.152939
R12558 gnd.n5055 gnd.n2898 0.152939
R12559 gnd.n5056 gnd.n5055 0.152939
R12560 gnd.n5057 gnd.n5056 0.152939
R12561 gnd.n5057 gnd.n2894 0.152939
R12562 gnd.n5064 gnd.n2894 0.152939
R12563 gnd.n5065 gnd.n5064 0.152939
R12564 gnd.n5066 gnd.n5065 0.152939
R12565 gnd.n5067 gnd.n5066 0.152939
R12566 gnd.n5068 gnd.n5067 0.152939
R12567 gnd.n5110 gnd.n5068 0.152939
R12568 gnd.n5113 gnd.n5110 0.152939
R12569 gnd.n5114 gnd.n5113 0.152939
R12570 gnd.n5115 gnd.n5114 0.152939
R12571 gnd.n5116 gnd.n5115 0.152939
R12572 gnd.n5117 gnd.n5116 0.152939
R12573 gnd.n5119 gnd.n5117 0.152939
R12574 gnd.n5119 gnd.n5118 0.152939
R12575 gnd.n5118 gnd.n253 0.152939
R12576 gnd.n254 gnd.n253 0.152939
R12577 gnd.n255 gnd.n254 0.152939
R12578 gnd.n598 gnd.n593 0.152939
R12579 gnd.n599 gnd.n598 0.152939
R12580 gnd.n600 gnd.n599 0.152939
R12581 gnd.n605 gnd.n600 0.152939
R12582 gnd.n606 gnd.n605 0.152939
R12583 gnd.n607 gnd.n606 0.152939
R12584 gnd.n608 gnd.n607 0.152939
R12585 gnd.n613 gnd.n608 0.152939
R12586 gnd.n614 gnd.n613 0.152939
R12587 gnd.n615 gnd.n614 0.152939
R12588 gnd.n616 gnd.n615 0.152939
R12589 gnd.n621 gnd.n616 0.152939
R12590 gnd.n622 gnd.n621 0.152939
R12591 gnd.n623 gnd.n622 0.152939
R12592 gnd.n624 gnd.n623 0.152939
R12593 gnd.n629 gnd.n624 0.152939
R12594 gnd.n630 gnd.n629 0.152939
R12595 gnd.n631 gnd.n630 0.152939
R12596 gnd.n632 gnd.n631 0.152939
R12597 gnd.n637 gnd.n632 0.152939
R12598 gnd.n638 gnd.n637 0.152939
R12599 gnd.n639 gnd.n638 0.152939
R12600 gnd.n640 gnd.n639 0.152939
R12601 gnd.n645 gnd.n640 0.152939
R12602 gnd.n646 gnd.n645 0.152939
R12603 gnd.n647 gnd.n646 0.152939
R12604 gnd.n648 gnd.n647 0.152939
R12605 gnd.n653 gnd.n648 0.152939
R12606 gnd.n654 gnd.n653 0.152939
R12607 gnd.n655 gnd.n654 0.152939
R12608 gnd.n656 gnd.n655 0.152939
R12609 gnd.n661 gnd.n656 0.152939
R12610 gnd.n662 gnd.n661 0.152939
R12611 gnd.n663 gnd.n662 0.152939
R12612 gnd.n664 gnd.n663 0.152939
R12613 gnd.n669 gnd.n664 0.152939
R12614 gnd.n670 gnd.n669 0.152939
R12615 gnd.n671 gnd.n670 0.152939
R12616 gnd.n672 gnd.n671 0.152939
R12617 gnd.n677 gnd.n672 0.152939
R12618 gnd.n678 gnd.n677 0.152939
R12619 gnd.n679 gnd.n678 0.152939
R12620 gnd.n680 gnd.n679 0.152939
R12621 gnd.n685 gnd.n680 0.152939
R12622 gnd.n686 gnd.n685 0.152939
R12623 gnd.n687 gnd.n686 0.152939
R12624 gnd.n688 gnd.n687 0.152939
R12625 gnd.n693 gnd.n688 0.152939
R12626 gnd.n694 gnd.n693 0.152939
R12627 gnd.n695 gnd.n694 0.152939
R12628 gnd.n696 gnd.n695 0.152939
R12629 gnd.n701 gnd.n696 0.152939
R12630 gnd.n702 gnd.n701 0.152939
R12631 gnd.n703 gnd.n702 0.152939
R12632 gnd.n704 gnd.n703 0.152939
R12633 gnd.n709 gnd.n704 0.152939
R12634 gnd.n710 gnd.n709 0.152939
R12635 gnd.n711 gnd.n710 0.152939
R12636 gnd.n712 gnd.n711 0.152939
R12637 gnd.n717 gnd.n712 0.152939
R12638 gnd.n718 gnd.n717 0.152939
R12639 gnd.n719 gnd.n718 0.152939
R12640 gnd.n720 gnd.n719 0.152939
R12641 gnd.n725 gnd.n720 0.152939
R12642 gnd.n726 gnd.n725 0.152939
R12643 gnd.n727 gnd.n726 0.152939
R12644 gnd.n728 gnd.n727 0.152939
R12645 gnd.n733 gnd.n728 0.152939
R12646 gnd.n734 gnd.n733 0.152939
R12647 gnd.n735 gnd.n734 0.152939
R12648 gnd.n736 gnd.n735 0.152939
R12649 gnd.n741 gnd.n736 0.152939
R12650 gnd.n742 gnd.n741 0.152939
R12651 gnd.n743 gnd.n742 0.152939
R12652 gnd.n744 gnd.n743 0.152939
R12653 gnd.n749 gnd.n744 0.152939
R12654 gnd.n750 gnd.n749 0.152939
R12655 gnd.n751 gnd.n750 0.152939
R12656 gnd.n752 gnd.n751 0.152939
R12657 gnd.n757 gnd.n752 0.152939
R12658 gnd.n758 gnd.n757 0.152939
R12659 gnd.n759 gnd.n758 0.152939
R12660 gnd.n760 gnd.n759 0.152939
R12661 gnd.n3633 gnd.n760 0.152939
R12662 gnd.n3995 gnd.n3994 0.152939
R12663 gnd.n3995 gnd.n3381 0.152939
R12664 gnd.n4009 gnd.n3381 0.152939
R12665 gnd.n4010 gnd.n4009 0.152939
R12666 gnd.n4011 gnd.n4010 0.152939
R12667 gnd.n4011 gnd.n3367 0.152939
R12668 gnd.n4025 gnd.n3367 0.152939
R12669 gnd.n4026 gnd.n4025 0.152939
R12670 gnd.n4039 gnd.n4026 0.152939
R12671 gnd.n4039 gnd.n4038 0.152939
R12672 gnd.n4038 gnd.n4037 0.152939
R12673 gnd.n4037 gnd.n4027 0.152939
R12674 gnd.n4033 gnd.n4027 0.152939
R12675 gnd.n4033 gnd.n4032 0.152939
R12676 gnd.n4032 gnd.n2622 0.152939
R12677 gnd.n5540 gnd.n2622 0.152939
R12678 gnd.n5540 gnd.n5539 0.152939
R12679 gnd.n5539 gnd.n5538 0.152939
R12680 gnd.n5538 gnd.n2623 0.152939
R12681 gnd.n5534 gnd.n2623 0.152939
R12682 gnd.n5534 gnd.n5533 0.152939
R12683 gnd.n5533 gnd.n5532 0.152939
R12684 gnd.n5532 gnd.n2628 0.152939
R12685 gnd.n5528 gnd.n2628 0.152939
R12686 gnd.n5528 gnd.n5527 0.152939
R12687 gnd.n5527 gnd.n5526 0.152939
R12688 gnd.n5526 gnd.n2633 0.152939
R12689 gnd.n5522 gnd.n2633 0.152939
R12690 gnd.n5522 gnd.n5521 0.152939
R12691 gnd.n5521 gnd.n5520 0.152939
R12692 gnd.n5520 gnd.n2638 0.152939
R12693 gnd.n5516 gnd.n2638 0.152939
R12694 gnd.n5516 gnd.n5515 0.152939
R12695 gnd.n5515 gnd.n5514 0.152939
R12696 gnd.n5514 gnd.n2643 0.152939
R12697 gnd.n5510 gnd.n2643 0.152939
R12698 gnd.n5510 gnd.n5509 0.152939
R12699 gnd.n5509 gnd.n5508 0.152939
R12700 gnd.n5508 gnd.n2648 0.152939
R12701 gnd.n5504 gnd.n2648 0.152939
R12702 gnd.n5504 gnd.n5503 0.152939
R12703 gnd.n5503 gnd.n5502 0.152939
R12704 gnd.n5502 gnd.n2653 0.152939
R12705 gnd.n5498 gnd.n2653 0.152939
R12706 gnd.n5498 gnd.n5497 0.152939
R12707 gnd.n5497 gnd.n5496 0.152939
R12708 gnd.n5496 gnd.n2658 0.152939
R12709 gnd.n5492 gnd.n2658 0.152939
R12710 gnd.n5492 gnd.n5491 0.152939
R12711 gnd.n5491 gnd.n5490 0.152939
R12712 gnd.n5490 gnd.n2663 0.152939
R12713 gnd.n5486 gnd.n2663 0.152939
R12714 gnd.n5486 gnd.n5485 0.152939
R12715 gnd.n5485 gnd.n5484 0.152939
R12716 gnd.n5484 gnd.n2668 0.152939
R12717 gnd.n5480 gnd.n2668 0.152939
R12718 gnd.n5480 gnd.n5479 0.152939
R12719 gnd.n5479 gnd.n5478 0.152939
R12720 gnd.n5478 gnd.n2673 0.152939
R12721 gnd.n5474 gnd.n2673 0.152939
R12722 gnd.n5474 gnd.n5473 0.152939
R12723 gnd.n5473 gnd.n5472 0.152939
R12724 gnd.n5472 gnd.n2678 0.152939
R12725 gnd.n5468 gnd.n2678 0.152939
R12726 gnd.n5468 gnd.n5467 0.152939
R12727 gnd.n5467 gnd.n5466 0.152939
R12728 gnd.n5466 gnd.n2683 0.152939
R12729 gnd.n5462 gnd.n2683 0.152939
R12730 gnd.n5462 gnd.n5461 0.152939
R12731 gnd.n5461 gnd.n5460 0.152939
R12732 gnd.n5460 gnd.n2688 0.152939
R12733 gnd.n5456 gnd.n2688 0.152939
R12734 gnd.n5456 gnd.n5455 0.152939
R12735 gnd.n5455 gnd.n5454 0.152939
R12736 gnd.n5454 gnd.n2693 0.152939
R12737 gnd.n5450 gnd.n2693 0.152939
R12738 gnd.n5450 gnd.n5449 0.152939
R12739 gnd.n5449 gnd.n5448 0.152939
R12740 gnd.n5448 gnd.n2698 0.152939
R12741 gnd.n5444 gnd.n2698 0.152939
R12742 gnd.n5444 gnd.n5443 0.152939
R12743 gnd.n5443 gnd.n5442 0.152939
R12744 gnd.n5442 gnd.n2703 0.152939
R12745 gnd.n5438 gnd.n2703 0.152939
R12746 gnd.n5438 gnd.n5437 0.152939
R12747 gnd.n5437 gnd.n5436 0.152939
R12748 gnd.n5436 gnd.n2708 0.152939
R12749 gnd.n5432 gnd.n2708 0.152939
R12750 gnd.n5432 gnd.n5431 0.152939
R12751 gnd.n5431 gnd.n5430 0.152939
R12752 gnd.n5430 gnd.n2713 0.152939
R12753 gnd.n5426 gnd.n2713 0.152939
R12754 gnd.n5426 gnd.n5425 0.152939
R12755 gnd.n5425 gnd.n5424 0.152939
R12756 gnd.n5424 gnd.n2718 0.152939
R12757 gnd.n5420 gnd.n2718 0.152939
R12758 gnd.n5420 gnd.n5419 0.152939
R12759 gnd.n5419 gnd.n5418 0.152939
R12760 gnd.n5418 gnd.n2723 0.152939
R12761 gnd.n5414 gnd.n2723 0.152939
R12762 gnd.n5414 gnd.n5413 0.152939
R12763 gnd.n3771 gnd.n3658 0.152939
R12764 gnd.n3776 gnd.n3658 0.152939
R12765 gnd.n3777 gnd.n3776 0.152939
R12766 gnd.n3778 gnd.n3777 0.152939
R12767 gnd.n3778 gnd.n3655 0.152939
R12768 gnd.n3833 gnd.n3655 0.152939
R12769 gnd.n3834 gnd.n3833 0.152939
R12770 gnd.n3835 gnd.n3834 0.152939
R12771 gnd.n3835 gnd.n3645 0.152939
R12772 gnd.n3880 gnd.n3645 0.152939
R12773 gnd.n3880 gnd.n3879 0.152939
R12774 gnd.n3879 gnd.n3878 0.152939
R12775 gnd.n3878 gnd.n3646 0.152939
R12776 gnd.n3874 gnd.n3646 0.152939
R12777 gnd.n3874 gnd.n3873 0.152939
R12778 gnd.n3873 gnd.n3872 0.152939
R12779 gnd.n3872 gnd.n3650 0.152939
R12780 gnd.n3868 gnd.n3650 0.152939
R12781 gnd.n3868 gnd.n3867 0.152939
R12782 gnd.n3867 gnd.n3866 0.152939
R12783 gnd.n3984 gnd.n3439 0.152939
R12784 gnd.n3984 gnd.n3983 0.152939
R12785 gnd.n3983 gnd.n3982 0.152939
R12786 gnd.n3982 gnd.n3441 0.152939
R12787 gnd.n3978 gnd.n3441 0.152939
R12788 gnd.n3978 gnd.n3977 0.152939
R12789 gnd.n3438 gnd.n3415 0.152939
R12790 gnd.n3434 gnd.n3415 0.152939
R12791 gnd.n3434 gnd.n3433 0.152939
R12792 gnd.n3433 gnd.n3432 0.152939
R12793 gnd.n3432 gnd.n3418 0.152939
R12794 gnd.n3428 gnd.n3418 0.152939
R12795 gnd.n3428 gnd.n3427 0.152939
R12796 gnd.n3427 gnd.n3426 0.152939
R12797 gnd.n3426 gnd.n3422 0.152939
R12798 gnd.n3422 gnd.n3349 0.152939
R12799 gnd.n4056 gnd.n3349 0.152939
R12800 gnd.n4057 gnd.n4056 0.152939
R12801 gnd.n4058 gnd.n4057 0.152939
R12802 gnd.n4058 gnd.n3346 0.152939
R12803 gnd.n4144 gnd.n3346 0.152939
R12804 gnd.n4145 gnd.n4144 0.152939
R12805 gnd.n4160 gnd.n4145 0.152939
R12806 gnd.n4160 gnd.n4159 0.152939
R12807 gnd.n4159 gnd.n4158 0.152939
R12808 gnd.n4158 gnd.n4146 0.152939
R12809 gnd.n4154 gnd.n4146 0.152939
R12810 gnd.n4154 gnd.n4153 0.152939
R12811 gnd.n4153 gnd.n4152 0.152939
R12812 gnd.n4152 gnd.n3302 0.152939
R12813 gnd.n4245 gnd.n3302 0.152939
R12814 gnd.n4245 gnd.n4244 0.152939
R12815 gnd.n4244 gnd.n4243 0.152939
R12816 gnd.n4243 gnd.n3303 0.152939
R12817 gnd.n4239 gnd.n3303 0.152939
R12818 gnd.n4239 gnd.n4238 0.152939
R12819 gnd.n4238 gnd.n4237 0.152939
R12820 gnd.n4237 gnd.n4225 0.152939
R12821 gnd.n4233 gnd.n4225 0.152939
R12822 gnd.n4233 gnd.n4232 0.152939
R12823 gnd.n4232 gnd.n4231 0.152939
R12824 gnd.n4231 gnd.n3233 0.152939
R12825 gnd.n4376 gnd.n3233 0.152939
R12826 gnd.n4377 gnd.n4376 0.152939
R12827 gnd.n4379 gnd.n4377 0.152939
R12828 gnd.n4379 gnd.n4378 0.152939
R12829 gnd.n4378 gnd.n3211 0.152939
R12830 gnd.n4408 gnd.n3211 0.152939
R12831 gnd.n4409 gnd.n4408 0.152939
R12832 gnd.n4424 gnd.n4409 0.152939
R12833 gnd.n4424 gnd.n4423 0.152939
R12834 gnd.n4423 gnd.n4422 0.152939
R12835 gnd.n4422 gnd.n4410 0.152939
R12836 gnd.n4418 gnd.n4410 0.152939
R12837 gnd.n4418 gnd.n4417 0.152939
R12838 gnd.n4417 gnd.n4416 0.152939
R12839 gnd.n4416 gnd.n3159 0.152939
R12840 gnd.n4518 gnd.n3159 0.152939
R12841 gnd.n4519 gnd.n4518 0.152939
R12842 gnd.n4521 gnd.n4519 0.152939
R12843 gnd.n4521 gnd.n4520 0.152939
R12844 gnd.n4520 gnd.n3135 0.152939
R12845 gnd.n4550 gnd.n3135 0.152939
R12846 gnd.n4551 gnd.n4550 0.152939
R12847 gnd.n4566 gnd.n4551 0.152939
R12848 gnd.n4566 gnd.n4565 0.152939
R12849 gnd.n4565 gnd.n4564 0.152939
R12850 gnd.n4564 gnd.n4552 0.152939
R12851 gnd.n4560 gnd.n4552 0.152939
R12852 gnd.n4560 gnd.n4559 0.152939
R12853 gnd.n4559 gnd.n4558 0.152939
R12854 gnd.n4558 gnd.n3083 0.152939
R12855 gnd.n4644 gnd.n3083 0.152939
R12856 gnd.n4645 gnd.n4644 0.152939
R12857 gnd.n4661 gnd.n4645 0.152939
R12858 gnd.n4661 gnd.n4660 0.152939
R12859 gnd.n4660 gnd.n4659 0.152939
R12860 gnd.n4659 gnd.n4646 0.152939
R12861 gnd.n4655 gnd.n4646 0.152939
R12862 gnd.n4655 gnd.n4654 0.152939
R12863 gnd.n4654 gnd.n4653 0.152939
R12864 gnd.n4653 gnd.n3031 0.152939
R12865 gnd.n4728 gnd.n3031 0.152939
R12866 gnd.n4729 gnd.n4728 0.152939
R12867 gnd.n4730 gnd.n4729 0.152939
R12868 gnd.n4730 gnd.n3029 0.152939
R12869 gnd.n4738 gnd.n3029 0.152939
R12870 gnd.n4739 gnd.n4738 0.152939
R12871 gnd.n4754 gnd.n4739 0.152939
R12872 gnd.n4754 gnd.n4753 0.152939
R12873 gnd.n4753 gnd.n4752 0.152939
R12874 gnd.n4752 gnd.n4740 0.152939
R12875 gnd.n4748 gnd.n4740 0.152939
R12876 gnd.n4748 gnd.n4747 0.152939
R12877 gnd.n4747 gnd.n4746 0.152939
R12878 gnd.n4746 gnd.n2928 0.152939
R12879 gnd.n4991 gnd.n2928 0.152939
R12880 gnd.n4992 gnd.n4991 0.152939
R12881 gnd.n4993 gnd.n4992 0.152939
R12882 gnd.n4993 gnd.n2917 0.152939
R12883 gnd.n5009 gnd.n2917 0.152939
R12884 gnd.n5010 gnd.n5009 0.152939
R12885 gnd.n5011 gnd.n5010 0.152939
R12886 gnd.n5011 gnd.n2905 0.152939
R12887 gnd.n5028 gnd.n2905 0.152939
R12888 gnd.n5029 gnd.n5028 0.152939
R12889 gnd.n5048 gnd.n5029 0.152939
R12890 gnd.n5047 gnd.n5030 0.152939
R12891 gnd.n5043 gnd.n5030 0.152939
R12892 gnd.n5043 gnd.n5042 0.152939
R12893 gnd.n5042 gnd.n5041 0.152939
R12894 gnd.n5041 gnd.n5034 0.152939
R12895 gnd.n5034 gnd.n2874 0.152939
R12896 gnd.n5139 gnd.n5134 0.152939
R12897 gnd.n5140 gnd.n5139 0.152939
R12898 gnd.n5141 gnd.n5140 0.152939
R12899 gnd.n5141 gnd.n5132 0.152939
R12900 gnd.n5164 gnd.n5132 0.152939
R12901 gnd.n5165 gnd.n5164 0.152939
R12902 gnd.n5167 gnd.n5165 0.152939
R12903 gnd.n5167 gnd.n5166 0.152939
R12904 gnd.n5166 gnd.n226 0.152939
R12905 gnd.n6764 gnd.n226 0.152939
R12906 gnd.n6765 gnd.n6764 0.152939
R12907 gnd.n6767 gnd.n6765 0.152939
R12908 gnd.n6767 gnd.n6766 0.152939
R12909 gnd.n6766 gnd.n199 0.152939
R12910 gnd.n6799 gnd.n199 0.152939
R12911 gnd.n6800 gnd.n6799 0.152939
R12912 gnd.n6806 gnd.n6800 0.152939
R12913 gnd.n6806 gnd.n6805 0.152939
R12914 gnd.n6805 gnd.n6804 0.152939
R12915 gnd.n6804 gnd.n67 0.152939
R12916 gnd.n7269 gnd.n7268 0.145814
R12917 gnd.n3770 gnd.n3769 0.145814
R12918 gnd.n3771 gnd.n3770 0.145814
R12919 gnd.n7269 gnd.n67 0.145814
R12920 gnd.n3977 gnd.n3976 0.128549
R12921 gnd.n5280 gnd.n2874 0.128549
R12922 gnd.n1173 gnd.n0 0.127478
R12923 gnd.n1686 gnd.n1049 0.0767195
R12924 gnd.n1686 gnd.n1685 0.0767195
R12925 gnd.n3976 gnd.n3446 0.063
R12926 gnd.n5281 gnd.n5280 0.063
R12927 gnd.n5281 gnd.n2873 0.0538288
R12928 gnd.n7206 gnd.n7205 0.0538288
R12929 gnd.n5809 gnd.n5808 0.0538288
R12930 gnd.n3858 gnd.n3446 0.0538288
R12931 gnd.n5987 gnd.n781 0.0477147
R12932 gnd.n1476 gnd.n1364 0.0442063
R12933 gnd.n1477 gnd.n1476 0.0442063
R12934 gnd.n1478 gnd.n1477 0.0442063
R12935 gnd.n1478 gnd.n1353 0.0442063
R12936 gnd.n1492 gnd.n1353 0.0442063
R12937 gnd.n1493 gnd.n1492 0.0442063
R12938 gnd.n1494 gnd.n1493 0.0442063
R12939 gnd.n1494 gnd.n1340 0.0442063
R12940 gnd.n1538 gnd.n1340 0.0442063
R12941 gnd.n1539 gnd.n1538 0.0442063
R12942 gnd.n5150 gnd.n2873 0.0344674
R12943 gnd.n5150 gnd.n5144 0.0344674
R12944 gnd.n5155 gnd.n5144 0.0344674
R12945 gnd.n5156 gnd.n5155 0.0344674
R12946 gnd.n5156 gnd.n5099 0.0344674
R12947 gnd.n5174 gnd.n5099 0.0344674
R12948 gnd.n5174 gnd.n5173 0.0344674
R12949 gnd.n5173 gnd.n246 0.0344674
R12950 gnd.n247 gnd.n246 0.0344674
R12951 gnd.n248 gnd.n247 0.0344674
R12952 gnd.n249 gnd.n248 0.0344674
R12953 gnd.n249 gnd.n221 0.0344674
R12954 gnd.n221 gnd.n218 0.0344674
R12955 gnd.n219 gnd.n218 0.0344674
R12956 gnd.n6778 gnd.n219 0.0344674
R12957 gnd.n6779 gnd.n6778 0.0344674
R12958 gnd.n6779 gnd.n192 0.0344674
R12959 gnd.n6815 gnd.n192 0.0344674
R12960 gnd.n6815 gnd.n175 0.0344674
R12961 gnd.n6832 gnd.n175 0.0344674
R12962 gnd.n6833 gnd.n6832 0.0344674
R12963 gnd.n6833 gnd.n169 0.0344674
R12964 gnd.n6841 gnd.n169 0.0344674
R12965 gnd.n6842 gnd.n6841 0.0344674
R12966 gnd.n6842 gnd.n90 0.0344674
R12967 gnd.n91 gnd.n90 0.0344674
R12968 gnd.n92 gnd.n91 0.0344674
R12969 gnd.n6849 gnd.n92 0.0344674
R12970 gnd.n6849 gnd.n109 0.0344674
R12971 gnd.n110 gnd.n109 0.0344674
R12972 gnd.n111 gnd.n110 0.0344674
R12973 gnd.n6856 gnd.n111 0.0344674
R12974 gnd.n6856 gnd.n128 0.0344674
R12975 gnd.n129 gnd.n128 0.0344674
R12976 gnd.n130 gnd.n129 0.0344674
R12977 gnd.n6863 gnd.n130 0.0344674
R12978 gnd.n6863 gnd.n148 0.0344674
R12979 gnd.n149 gnd.n148 0.0344674
R12980 gnd.n150 gnd.n149 0.0344674
R12981 gnd.n6870 gnd.n150 0.0344674
R12982 gnd.n6870 gnd.n167 0.0344674
R12983 gnd.n7206 gnd.n167 0.0344674
R12984 gnd.n1541 gnd.n1274 0.0344674
R12985 gnd.n5808 gnd.n2263 0.0344674
R12986 gnd.n3782 gnd.n2263 0.0344674
R12987 gnd.n3782 gnd.n2284 0.0344674
R12988 gnd.n2285 gnd.n2284 0.0344674
R12989 gnd.n2286 gnd.n2285 0.0344674
R12990 gnd.n3789 gnd.n2286 0.0344674
R12991 gnd.n3789 gnd.n2302 0.0344674
R12992 gnd.n2303 gnd.n2302 0.0344674
R12993 gnd.n2304 gnd.n2303 0.0344674
R12994 gnd.n3796 gnd.n2304 0.0344674
R12995 gnd.n3796 gnd.n2320 0.0344674
R12996 gnd.n2321 gnd.n2320 0.0344674
R12997 gnd.n2322 gnd.n2321 0.0344674
R12998 gnd.n3803 gnd.n2322 0.0344674
R12999 gnd.n3803 gnd.n2340 0.0344674
R13000 gnd.n2341 gnd.n2340 0.0344674
R13001 gnd.n2342 gnd.n2341 0.0344674
R13002 gnd.n3810 gnd.n2342 0.0344674
R13003 gnd.n3810 gnd.n2358 0.0344674
R13004 gnd.n2359 gnd.n2358 0.0344674
R13005 gnd.n2360 gnd.n2359 0.0344674
R13006 gnd.n3817 gnd.n2360 0.0344674
R13007 gnd.n3817 gnd.n2378 0.0344674
R13008 gnd.n2379 gnd.n2378 0.0344674
R13009 gnd.n2380 gnd.n2379 0.0344674
R13010 gnd.n3824 gnd.n2380 0.0344674
R13011 gnd.n3824 gnd.n2397 0.0344674
R13012 gnd.n2398 gnd.n2397 0.0344674
R13013 gnd.n2399 gnd.n2398 0.0344674
R13014 gnd.n3653 gnd.n2399 0.0344674
R13015 gnd.n3653 gnd.n2418 0.0344674
R13016 gnd.n2419 gnd.n2418 0.0344674
R13017 gnd.n2420 gnd.n2419 0.0344674
R13018 gnd.n3844 gnd.n2420 0.0344674
R13019 gnd.n3844 gnd.n2438 0.0344674
R13020 gnd.n2439 gnd.n2438 0.0344674
R13021 gnd.n2440 gnd.n2439 0.0344674
R13022 gnd.n3853 gnd.n2440 0.0344674
R13023 gnd.n3853 gnd.n2459 0.0344674
R13024 gnd.n2460 gnd.n2459 0.0344674
R13025 gnd.n2461 gnd.n2460 0.0344674
R13026 gnd.n3858 gnd.n2461 0.0344674
R13027 gnd.n3975 gnd.n3447 0.0343753
R13028 gnd.n5279 gnd.n2875 0.0343753
R13029 gnd.n3518 gnd.n3395 0.0296328
R13030 gnd.n2758 gnd.n2728 0.0296328
R13031 gnd.n1561 gnd.n1560 0.0269946
R13032 gnd.n1563 gnd.n1562 0.0269946
R13033 gnd.n1269 gnd.n1267 0.0269946
R13034 gnd.n1573 gnd.n1571 0.0269946
R13035 gnd.n1572 gnd.n1248 0.0269946
R13036 gnd.n1592 gnd.n1591 0.0269946
R13037 gnd.n1594 gnd.n1593 0.0269946
R13038 gnd.n1243 gnd.n1242 0.0269946
R13039 gnd.n1604 gnd.n1238 0.0269946
R13040 gnd.n1603 gnd.n1240 0.0269946
R13041 gnd.n1239 gnd.n1219 0.0269946
R13042 gnd.n1630 gnd.n1220 0.0269946
R13043 gnd.n1629 gnd.n1221 0.0269946
R13044 gnd.n1649 gnd.n1205 0.0269946
R13045 gnd.n1651 gnd.n1650 0.0269946
R13046 gnd.n1652 gnd.n1185 0.0269946
R13047 gnd.n1653 gnd.n1186 0.0269946
R13048 gnd.n1654 gnd.n1187 0.0269946
R13049 gnd.n1189 gnd.n1188 0.0269946
R13050 gnd.n1043 gnd.n1041 0.0269946
R13051 gnd.n1698 gnd.n1696 0.0269946
R13052 gnd.n1697 gnd.n1025 0.0269946
R13053 gnd.n1717 gnd.n1716 0.0269946
R13054 gnd.n1719 gnd.n1718 0.0269946
R13055 gnd.n1020 gnd.n1018 0.0269946
R13056 gnd.n1729 gnd.n1727 0.0269946
R13057 gnd.n1728 gnd.n1000 0.0269946
R13058 gnd.n1748 gnd.n1747 0.0269946
R13059 gnd.n1750 gnd.n1749 0.0269946
R13060 gnd.n994 gnd.n992 0.0269946
R13061 gnd.n1760 gnd.n1758 0.0269946
R13062 gnd.n1759 gnd.n973 0.0269946
R13063 gnd.n1779 gnd.n1778 0.0269946
R13064 gnd.n1781 gnd.n1780 0.0269946
R13065 gnd.n968 gnd.n966 0.0269946
R13066 gnd.n1791 gnd.n1789 0.0269946
R13067 gnd.n1790 gnd.n949 0.0269946
R13068 gnd.n1810 gnd.n1809 0.0269946
R13069 gnd.n1812 gnd.n1811 0.0269946
R13070 gnd.n944 gnd.n942 0.0269946
R13071 gnd.n1822 gnd.n1820 0.0269946
R13072 gnd.n1821 gnd.n923 0.0269946
R13073 gnd.n1841 gnd.n1840 0.0269946
R13074 gnd.n1843 gnd.n1842 0.0269946
R13075 gnd.n918 gnd.n916 0.0269946
R13076 gnd.n1853 gnd.n1851 0.0269946
R13077 gnd.n1852 gnd.n898 0.0269946
R13078 gnd.n1873 gnd.n1872 0.0269946
R13079 gnd.n892 gnd.n891 0.0269946
R13080 gnd.n2142 gnd.n888 0.0269946
R13081 gnd.n2141 gnd.n889 0.0269946
R13082 gnd.n5988 gnd.n780 0.0269946
R13083 gnd.n3971 gnd.n3453 0.022519
R13084 gnd.n3970 gnd.n3454 0.022519
R13085 gnd.n3967 gnd.n3966 0.022519
R13086 gnd.n3963 gnd.n3460 0.022519
R13087 gnd.n3962 gnd.n3466 0.022519
R13088 gnd.n3959 gnd.n3958 0.022519
R13089 gnd.n3955 gnd.n3470 0.022519
R13090 gnd.n3954 gnd.n3474 0.022519
R13091 gnd.n3951 gnd.n3950 0.022519
R13092 gnd.n3947 gnd.n3480 0.022519
R13093 gnd.n3946 gnd.n3486 0.022519
R13094 gnd.n3943 gnd.n3942 0.022519
R13095 gnd.n3939 gnd.n3490 0.022519
R13096 gnd.n3938 gnd.n3494 0.022519
R13097 gnd.n3935 gnd.n3934 0.022519
R13098 gnd.n3931 gnd.n3500 0.022519
R13099 gnd.n3930 gnd.n3507 0.022519
R13100 gnd.n3517 gnd.n3511 0.022519
R13101 gnd.n3519 gnd.n3518 0.022519
R13102 gnd.n5275 gnd.n2882 0.022519
R13103 gnd.n5274 gnd.n2883 0.022519
R13104 gnd.n5271 gnd.n5270 0.022519
R13105 gnd.n5267 gnd.n5199 0.022519
R13106 gnd.n5266 gnd.n5203 0.022519
R13107 gnd.n5263 gnd.n5262 0.022519
R13108 gnd.n5259 gnd.n5209 0.022519
R13109 gnd.n5258 gnd.n5215 0.022519
R13110 gnd.n5255 gnd.n5254 0.022519
R13111 gnd.n5251 gnd.n5219 0.022519
R13112 gnd.n5250 gnd.n5223 0.022519
R13113 gnd.n5247 gnd.n5246 0.022519
R13114 gnd.n5243 gnd.n5229 0.022519
R13115 gnd.n5242 gnd.n5235 0.022519
R13116 gnd.n5239 gnd.n5238 0.022519
R13117 gnd.n5405 gnd.n2753 0.022519
R13118 gnd.n5404 gnd.n2754 0.022519
R13119 gnd.n2764 gnd.n2763 0.022519
R13120 gnd.n2759 gnd.n2758 0.022519
R13121 gnd.n5412 gnd.n2728 0.0218415
R13122 gnd.n3993 gnd.n3395 0.0218415
R13123 gnd.n1541 gnd.n1540 0.0202011
R13124 gnd.n1540 gnd.n1539 0.0148637
R13125 gnd.n2130 gnd.n1874 0.0144266
R13126 gnd.n2131 gnd.n2130 0.0130679
R13127 gnd.n3453 gnd.n3447 0.0123564
R13128 gnd.n3971 gnd.n3970 0.0123564
R13129 gnd.n3967 gnd.n3454 0.0123564
R13130 gnd.n3966 gnd.n3460 0.0123564
R13131 gnd.n3963 gnd.n3962 0.0123564
R13132 gnd.n3959 gnd.n3466 0.0123564
R13133 gnd.n3958 gnd.n3470 0.0123564
R13134 gnd.n3955 gnd.n3954 0.0123564
R13135 gnd.n3951 gnd.n3474 0.0123564
R13136 gnd.n3950 gnd.n3480 0.0123564
R13137 gnd.n3947 gnd.n3946 0.0123564
R13138 gnd.n3943 gnd.n3486 0.0123564
R13139 gnd.n3942 gnd.n3490 0.0123564
R13140 gnd.n3939 gnd.n3938 0.0123564
R13141 gnd.n3935 gnd.n3494 0.0123564
R13142 gnd.n3934 gnd.n3500 0.0123564
R13143 gnd.n3931 gnd.n3930 0.0123564
R13144 gnd.n3511 gnd.n3507 0.0123564
R13145 gnd.n3519 gnd.n3517 0.0123564
R13146 gnd.n2882 gnd.n2875 0.0123564
R13147 gnd.n5275 gnd.n5274 0.0123564
R13148 gnd.n5271 gnd.n2883 0.0123564
R13149 gnd.n5270 gnd.n5199 0.0123564
R13150 gnd.n5267 gnd.n5266 0.0123564
R13151 gnd.n5263 gnd.n5203 0.0123564
R13152 gnd.n5262 gnd.n5209 0.0123564
R13153 gnd.n5259 gnd.n5258 0.0123564
R13154 gnd.n5255 gnd.n5215 0.0123564
R13155 gnd.n5254 gnd.n5219 0.0123564
R13156 gnd.n5251 gnd.n5250 0.0123564
R13157 gnd.n5247 gnd.n5223 0.0123564
R13158 gnd.n5246 gnd.n5229 0.0123564
R13159 gnd.n5243 gnd.n5242 0.0123564
R13160 gnd.n5239 gnd.n5235 0.0123564
R13161 gnd.n5238 gnd.n2753 0.0123564
R13162 gnd.n5405 gnd.n5404 0.0123564
R13163 gnd.n2764 gnd.n2754 0.0123564
R13164 gnd.n2763 gnd.n2759 0.0123564
R13165 gnd.n1560 gnd.n1274 0.00797283
R13166 gnd.n1562 gnd.n1561 0.00797283
R13167 gnd.n1563 gnd.n1269 0.00797283
R13168 gnd.n1571 gnd.n1267 0.00797283
R13169 gnd.n1573 gnd.n1572 0.00797283
R13170 gnd.n1591 gnd.n1248 0.00797283
R13171 gnd.n1593 gnd.n1592 0.00797283
R13172 gnd.n1594 gnd.n1243 0.00797283
R13173 gnd.n1242 gnd.n1238 0.00797283
R13174 gnd.n1604 gnd.n1603 0.00797283
R13175 gnd.n1240 gnd.n1239 0.00797283
R13176 gnd.n1220 gnd.n1219 0.00797283
R13177 gnd.n1630 gnd.n1629 0.00797283
R13178 gnd.n1221 gnd.n1205 0.00797283
R13179 gnd.n1650 gnd.n1649 0.00797283
R13180 gnd.n1652 gnd.n1651 0.00797283
R13181 gnd.n1653 gnd.n1185 0.00797283
R13182 gnd.n1654 gnd.n1186 0.00797283
R13183 gnd.n1188 gnd.n1187 0.00797283
R13184 gnd.n1189 gnd.n1043 0.00797283
R13185 gnd.n1696 gnd.n1041 0.00797283
R13186 gnd.n1698 gnd.n1697 0.00797283
R13187 gnd.n1716 gnd.n1025 0.00797283
R13188 gnd.n1718 gnd.n1717 0.00797283
R13189 gnd.n1719 gnd.n1020 0.00797283
R13190 gnd.n1727 gnd.n1018 0.00797283
R13191 gnd.n1729 gnd.n1728 0.00797283
R13192 gnd.n1747 gnd.n1000 0.00797283
R13193 gnd.n1749 gnd.n1748 0.00797283
R13194 gnd.n1750 gnd.n994 0.00797283
R13195 gnd.n1758 gnd.n992 0.00797283
R13196 gnd.n1760 gnd.n1759 0.00797283
R13197 gnd.n1778 gnd.n973 0.00797283
R13198 gnd.n1780 gnd.n1779 0.00797283
R13199 gnd.n1781 gnd.n968 0.00797283
R13200 gnd.n1789 gnd.n966 0.00797283
R13201 gnd.n1791 gnd.n1790 0.00797283
R13202 gnd.n1809 gnd.n949 0.00797283
R13203 gnd.n1811 gnd.n1810 0.00797283
R13204 gnd.n1812 gnd.n944 0.00797283
R13205 gnd.n1820 gnd.n942 0.00797283
R13206 gnd.n1822 gnd.n1821 0.00797283
R13207 gnd.n1840 gnd.n923 0.00797283
R13208 gnd.n1842 gnd.n1841 0.00797283
R13209 gnd.n1843 gnd.n918 0.00797283
R13210 gnd.n1851 gnd.n916 0.00797283
R13211 gnd.n1853 gnd.n1852 0.00797283
R13212 gnd.n1872 gnd.n898 0.00797283
R13213 gnd.n1874 gnd.n1873 0.00797283
R13214 gnd.n2131 gnd.n892 0.00797283
R13215 gnd.n891 gnd.n888 0.00797283
R13216 gnd.n2142 gnd.n2141 0.00797283
R13217 gnd.n889 gnd.n780 0.00797283
R13218 gnd.n5988 gnd.n5987 0.00797283
R13219 gnd.n3976 gnd.n3975 0.00592005
R13220 gnd.n5280 gnd.n5279 0.00592005
R13221 gnd.n6792 gnd.n184 0.00417647
R13222 gnd.n6821 gnd.n184 0.00417647
R13223 gnd.n6822 gnd.n6821 0.00417647
R13224 gnd.n6823 gnd.n6822 0.00417647
R13225 gnd.n6825 gnd.n6823 0.00417647
R13226 gnd.n6825 gnd.n6824 0.00417647
R13227 gnd.n6824 gnd.n79 0.00417647
R13228 gnd.n80 gnd.n79 0.00417647
R13229 gnd.n81 gnd.n80 0.00417647
R13230 gnd.n98 gnd.n81 0.00417647
R13231 gnd.n2349 gnd.n2348 0.00417647
R13232 gnd.n2350 gnd.n2349 0.00417647
R13233 gnd.n2351 gnd.n2350 0.00417647
R13234 gnd.n2368 gnd.n2351 0.00417647
R13235 gnd.n2369 gnd.n2368 0.00417647
R13236 gnd.n2370 gnd.n2369 0.00417647
R13237 gnd.n2371 gnd.n2370 0.00417647
R13238 gnd.n2387 gnd.n2371 0.00417647
R13239 gnd.n2388 gnd.n2387 0.00417647
R13240 gnd.n2389 gnd.n2388 0.00417647
R13241 commonsourceibias.n25 commonsourceibias.t34 230.006
R13242 commonsourceibias.n91 commonsourceibias.t95 230.006
R13243 commonsourceibias.n218 commonsourceibias.t117 230.006
R13244 commonsourceibias.n154 commonsourceibias.t97 230.006
R13245 commonsourceibias.n322 commonsourceibias.t4 230.006
R13246 commonsourceibias.n281 commonsourceibias.t70 230.006
R13247 commonsourceibias.n483 commonsourceibias.t55 230.006
R13248 commonsourceibias.n419 commonsourceibias.t80 230.006
R13249 commonsourceibias.n70 commonsourceibias.t16 207.983
R13250 commonsourceibias.n136 commonsourceibias.t56 207.983
R13251 commonsourceibias.n263 commonsourceibias.t111 207.983
R13252 commonsourceibias.n199 commonsourceibias.t89 207.983
R13253 commonsourceibias.n368 commonsourceibias.t26 207.983
R13254 commonsourceibias.n402 commonsourceibias.t114 207.983
R13255 commonsourceibias.n529 commonsourceibias.t51 207.983
R13256 commonsourceibias.n465 commonsourceibias.t74 207.983
R13257 commonsourceibias.n10 commonsourceibias.t30 168.701
R13258 commonsourceibias.n63 commonsourceibias.t2 168.701
R13259 commonsourceibias.n57 commonsourceibias.t22 168.701
R13260 commonsourceibias.n16 commonsourceibias.t42 168.701
R13261 commonsourceibias.n49 commonsourceibias.t18 168.701
R13262 commonsourceibias.n43 commonsourceibias.t32 168.701
R13263 commonsourceibias.n19 commonsourceibias.t40 168.701
R13264 commonsourceibias.n21 commonsourceibias.t24 168.701
R13265 commonsourceibias.n23 commonsourceibias.t44 168.701
R13266 commonsourceibias.n26 commonsourceibias.t6 168.701
R13267 commonsourceibias.n1 commonsourceibias.t109 168.701
R13268 commonsourceibias.n129 commonsourceibias.t69 168.701
R13269 commonsourceibias.n123 commonsourceibias.t119 168.701
R13270 commonsourceibias.n7 commonsourceibias.t85 168.701
R13271 commonsourceibias.n115 commonsourceibias.t54 168.701
R13272 commonsourceibias.n109 commonsourceibias.t100 168.701
R13273 commonsourceibias.n85 commonsourceibias.t87 168.701
R13274 commonsourceibias.n87 commonsourceibias.t115 168.701
R13275 commonsourceibias.n89 commonsourceibias.t79 168.701
R13276 commonsourceibias.n92 commonsourceibias.t66 168.701
R13277 commonsourceibias.n219 commonsourceibias.t75 168.701
R13278 commonsourceibias.n216 commonsourceibias.t59 168.701
R13279 commonsourceibias.n214 commonsourceibias.t49 168.701
R13280 commonsourceibias.n212 commonsourceibias.t84 168.701
R13281 commonsourceibias.n236 commonsourceibias.t93 168.701
R13282 commonsourceibias.n242 commonsourceibias.t52 168.701
R13283 commonsourceibias.n209 commonsourceibias.t118 168.701
R13284 commonsourceibias.n250 commonsourceibias.t104 168.701
R13285 commonsourceibias.n256 commonsourceibias.t60 168.701
R13286 commonsourceibias.n203 commonsourceibias.t50 168.701
R13287 commonsourceibias.n139 commonsourceibias.t106 168.701
R13288 commonsourceibias.n192 commonsourceibias.t101 168.701
R13289 commonsourceibias.n186 commonsourceibias.t88 168.701
R13290 commonsourceibias.n145 commonsourceibias.t105 168.701
R13291 commonsourceibias.n178 commonsourceibias.t99 168.701
R13292 commonsourceibias.n172 commonsourceibias.t86 168.701
R13293 commonsourceibias.n148 commonsourceibias.t108 168.701
R13294 commonsourceibias.n150 commonsourceibias.t98 168.701
R13295 commonsourceibias.n152 commonsourceibias.t112 168.701
R13296 commonsourceibias.n155 commonsourceibias.t107 168.701
R13297 commonsourceibias.n323 commonsourceibias.t14 168.701
R13298 commonsourceibias.n320 commonsourceibias.t12 168.701
R13299 commonsourceibias.n318 commonsourceibias.t38 168.701
R13300 commonsourceibias.n316 commonsourceibias.t8 168.701
R13301 commonsourceibias.n340 commonsourceibias.t0 168.701
R13302 commonsourceibias.n346 commonsourceibias.t28 168.701
R13303 commonsourceibias.n348 commonsourceibias.t10 168.701
R13304 commonsourceibias.n355 commonsourceibias.t36 168.701
R13305 commonsourceibias.n361 commonsourceibias.t20 168.701
R13306 commonsourceibias.n308 commonsourceibias.t46 168.701
R13307 commonsourceibias.n267 commonsourceibias.t78 168.701
R13308 commonsourceibias.n395 commonsourceibias.t53 168.701
R13309 commonsourceibias.n389 commonsourceibias.t94 168.701
R13310 commonsourceibias.n382 commonsourceibias.t64 168.701
R13311 commonsourceibias.n380 commonsourceibias.t113 168.701
R13312 commonsourceibias.n282 commonsourceibias.t58 168.701
R13313 commonsourceibias.n279 commonsourceibias.t63 168.701
R13314 commonsourceibias.n277 commonsourceibias.t92 168.701
R13315 commonsourceibias.n275 commonsourceibias.t65 168.701
R13316 commonsourceibias.n299 commonsourceibias.t76 168.701
R13317 commonsourceibias.n484 commonsourceibias.t68 168.701
R13318 commonsourceibias.n481 commonsourceibias.t72 168.701
R13319 commonsourceibias.n479 commonsourceibias.t61 168.701
R13320 commonsourceibias.n477 commonsourceibias.t110 168.701
R13321 commonsourceibias.n501 commonsourceibias.t77 168.701
R13322 commonsourceibias.n507 commonsourceibias.t67 168.701
R13323 commonsourceibias.n509 commonsourceibias.t57 168.701
R13324 commonsourceibias.n516 commonsourceibias.t48 168.701
R13325 commonsourceibias.n522 commonsourceibias.t71 168.701
R13326 commonsourceibias.n469 commonsourceibias.t62 168.701
R13327 commonsourceibias.n420 commonsourceibias.t116 168.701
R13328 commonsourceibias.n417 commonsourceibias.t102 168.701
R13329 commonsourceibias.n415 commonsourceibias.t81 168.701
R13330 commonsourceibias.n413 commonsourceibias.t96 168.701
R13331 commonsourceibias.n437 commonsourceibias.t103 168.701
R13332 commonsourceibias.n443 commonsourceibias.t82 168.701
R13333 commonsourceibias.n445 commonsourceibias.t90 168.701
R13334 commonsourceibias.n452 commonsourceibias.t73 168.701
R13335 commonsourceibias.n458 commonsourceibias.t83 168.701
R13336 commonsourceibias.n405 commonsourceibias.t91 168.701
R13337 commonsourceibias.n27 commonsourceibias.n24 161.3
R13338 commonsourceibias.n29 commonsourceibias.n28 161.3
R13339 commonsourceibias.n31 commonsourceibias.n30 161.3
R13340 commonsourceibias.n32 commonsourceibias.n22 161.3
R13341 commonsourceibias.n34 commonsourceibias.n33 161.3
R13342 commonsourceibias.n36 commonsourceibias.n35 161.3
R13343 commonsourceibias.n37 commonsourceibias.n20 161.3
R13344 commonsourceibias.n39 commonsourceibias.n38 161.3
R13345 commonsourceibias.n41 commonsourceibias.n40 161.3
R13346 commonsourceibias.n42 commonsourceibias.n18 161.3
R13347 commonsourceibias.n45 commonsourceibias.n44 161.3
R13348 commonsourceibias.n46 commonsourceibias.n17 161.3
R13349 commonsourceibias.n48 commonsourceibias.n47 161.3
R13350 commonsourceibias.n50 commonsourceibias.n15 161.3
R13351 commonsourceibias.n52 commonsourceibias.n51 161.3
R13352 commonsourceibias.n53 commonsourceibias.n14 161.3
R13353 commonsourceibias.n55 commonsourceibias.n54 161.3
R13354 commonsourceibias.n56 commonsourceibias.n13 161.3
R13355 commonsourceibias.n59 commonsourceibias.n58 161.3
R13356 commonsourceibias.n60 commonsourceibias.n12 161.3
R13357 commonsourceibias.n62 commonsourceibias.n61 161.3
R13358 commonsourceibias.n64 commonsourceibias.n11 161.3
R13359 commonsourceibias.n66 commonsourceibias.n65 161.3
R13360 commonsourceibias.n68 commonsourceibias.n67 161.3
R13361 commonsourceibias.n69 commonsourceibias.n9 161.3
R13362 commonsourceibias.n93 commonsourceibias.n90 161.3
R13363 commonsourceibias.n95 commonsourceibias.n94 161.3
R13364 commonsourceibias.n97 commonsourceibias.n96 161.3
R13365 commonsourceibias.n98 commonsourceibias.n88 161.3
R13366 commonsourceibias.n100 commonsourceibias.n99 161.3
R13367 commonsourceibias.n102 commonsourceibias.n101 161.3
R13368 commonsourceibias.n103 commonsourceibias.n86 161.3
R13369 commonsourceibias.n105 commonsourceibias.n104 161.3
R13370 commonsourceibias.n107 commonsourceibias.n106 161.3
R13371 commonsourceibias.n108 commonsourceibias.n84 161.3
R13372 commonsourceibias.n111 commonsourceibias.n110 161.3
R13373 commonsourceibias.n112 commonsourceibias.n8 161.3
R13374 commonsourceibias.n114 commonsourceibias.n113 161.3
R13375 commonsourceibias.n116 commonsourceibias.n6 161.3
R13376 commonsourceibias.n118 commonsourceibias.n117 161.3
R13377 commonsourceibias.n119 commonsourceibias.n5 161.3
R13378 commonsourceibias.n121 commonsourceibias.n120 161.3
R13379 commonsourceibias.n122 commonsourceibias.n4 161.3
R13380 commonsourceibias.n125 commonsourceibias.n124 161.3
R13381 commonsourceibias.n126 commonsourceibias.n3 161.3
R13382 commonsourceibias.n128 commonsourceibias.n127 161.3
R13383 commonsourceibias.n130 commonsourceibias.n2 161.3
R13384 commonsourceibias.n132 commonsourceibias.n131 161.3
R13385 commonsourceibias.n134 commonsourceibias.n133 161.3
R13386 commonsourceibias.n135 commonsourceibias.n0 161.3
R13387 commonsourceibias.n262 commonsourceibias.n202 161.3
R13388 commonsourceibias.n261 commonsourceibias.n260 161.3
R13389 commonsourceibias.n259 commonsourceibias.n258 161.3
R13390 commonsourceibias.n257 commonsourceibias.n204 161.3
R13391 commonsourceibias.n255 commonsourceibias.n254 161.3
R13392 commonsourceibias.n253 commonsourceibias.n205 161.3
R13393 commonsourceibias.n252 commonsourceibias.n251 161.3
R13394 commonsourceibias.n249 commonsourceibias.n206 161.3
R13395 commonsourceibias.n248 commonsourceibias.n247 161.3
R13396 commonsourceibias.n246 commonsourceibias.n207 161.3
R13397 commonsourceibias.n245 commonsourceibias.n244 161.3
R13398 commonsourceibias.n243 commonsourceibias.n208 161.3
R13399 commonsourceibias.n241 commonsourceibias.n240 161.3
R13400 commonsourceibias.n239 commonsourceibias.n210 161.3
R13401 commonsourceibias.n238 commonsourceibias.n237 161.3
R13402 commonsourceibias.n235 commonsourceibias.n211 161.3
R13403 commonsourceibias.n234 commonsourceibias.n233 161.3
R13404 commonsourceibias.n232 commonsourceibias.n231 161.3
R13405 commonsourceibias.n230 commonsourceibias.n213 161.3
R13406 commonsourceibias.n229 commonsourceibias.n228 161.3
R13407 commonsourceibias.n227 commonsourceibias.n226 161.3
R13408 commonsourceibias.n225 commonsourceibias.n215 161.3
R13409 commonsourceibias.n224 commonsourceibias.n223 161.3
R13410 commonsourceibias.n222 commonsourceibias.n221 161.3
R13411 commonsourceibias.n220 commonsourceibias.n217 161.3
R13412 commonsourceibias.n156 commonsourceibias.n153 161.3
R13413 commonsourceibias.n158 commonsourceibias.n157 161.3
R13414 commonsourceibias.n160 commonsourceibias.n159 161.3
R13415 commonsourceibias.n161 commonsourceibias.n151 161.3
R13416 commonsourceibias.n163 commonsourceibias.n162 161.3
R13417 commonsourceibias.n165 commonsourceibias.n164 161.3
R13418 commonsourceibias.n166 commonsourceibias.n149 161.3
R13419 commonsourceibias.n168 commonsourceibias.n167 161.3
R13420 commonsourceibias.n170 commonsourceibias.n169 161.3
R13421 commonsourceibias.n171 commonsourceibias.n147 161.3
R13422 commonsourceibias.n174 commonsourceibias.n173 161.3
R13423 commonsourceibias.n175 commonsourceibias.n146 161.3
R13424 commonsourceibias.n177 commonsourceibias.n176 161.3
R13425 commonsourceibias.n179 commonsourceibias.n144 161.3
R13426 commonsourceibias.n181 commonsourceibias.n180 161.3
R13427 commonsourceibias.n182 commonsourceibias.n143 161.3
R13428 commonsourceibias.n184 commonsourceibias.n183 161.3
R13429 commonsourceibias.n185 commonsourceibias.n142 161.3
R13430 commonsourceibias.n188 commonsourceibias.n187 161.3
R13431 commonsourceibias.n189 commonsourceibias.n141 161.3
R13432 commonsourceibias.n191 commonsourceibias.n190 161.3
R13433 commonsourceibias.n193 commonsourceibias.n140 161.3
R13434 commonsourceibias.n195 commonsourceibias.n194 161.3
R13435 commonsourceibias.n197 commonsourceibias.n196 161.3
R13436 commonsourceibias.n198 commonsourceibias.n138 161.3
R13437 commonsourceibias.n367 commonsourceibias.n307 161.3
R13438 commonsourceibias.n366 commonsourceibias.n365 161.3
R13439 commonsourceibias.n364 commonsourceibias.n363 161.3
R13440 commonsourceibias.n362 commonsourceibias.n309 161.3
R13441 commonsourceibias.n360 commonsourceibias.n359 161.3
R13442 commonsourceibias.n358 commonsourceibias.n310 161.3
R13443 commonsourceibias.n357 commonsourceibias.n356 161.3
R13444 commonsourceibias.n354 commonsourceibias.n311 161.3
R13445 commonsourceibias.n353 commonsourceibias.n352 161.3
R13446 commonsourceibias.n351 commonsourceibias.n312 161.3
R13447 commonsourceibias.n350 commonsourceibias.n349 161.3
R13448 commonsourceibias.n347 commonsourceibias.n313 161.3
R13449 commonsourceibias.n345 commonsourceibias.n344 161.3
R13450 commonsourceibias.n343 commonsourceibias.n314 161.3
R13451 commonsourceibias.n342 commonsourceibias.n341 161.3
R13452 commonsourceibias.n339 commonsourceibias.n315 161.3
R13453 commonsourceibias.n338 commonsourceibias.n337 161.3
R13454 commonsourceibias.n336 commonsourceibias.n335 161.3
R13455 commonsourceibias.n334 commonsourceibias.n317 161.3
R13456 commonsourceibias.n333 commonsourceibias.n332 161.3
R13457 commonsourceibias.n331 commonsourceibias.n330 161.3
R13458 commonsourceibias.n329 commonsourceibias.n319 161.3
R13459 commonsourceibias.n328 commonsourceibias.n327 161.3
R13460 commonsourceibias.n326 commonsourceibias.n325 161.3
R13461 commonsourceibias.n324 commonsourceibias.n321 161.3
R13462 commonsourceibias.n301 commonsourceibias.n300 161.3
R13463 commonsourceibias.n298 commonsourceibias.n274 161.3
R13464 commonsourceibias.n297 commonsourceibias.n296 161.3
R13465 commonsourceibias.n295 commonsourceibias.n294 161.3
R13466 commonsourceibias.n293 commonsourceibias.n276 161.3
R13467 commonsourceibias.n292 commonsourceibias.n291 161.3
R13468 commonsourceibias.n290 commonsourceibias.n289 161.3
R13469 commonsourceibias.n288 commonsourceibias.n278 161.3
R13470 commonsourceibias.n287 commonsourceibias.n286 161.3
R13471 commonsourceibias.n285 commonsourceibias.n284 161.3
R13472 commonsourceibias.n283 commonsourceibias.n280 161.3
R13473 commonsourceibias.n377 commonsourceibias.n273 161.3
R13474 commonsourceibias.n401 commonsourceibias.n266 161.3
R13475 commonsourceibias.n400 commonsourceibias.n399 161.3
R13476 commonsourceibias.n398 commonsourceibias.n397 161.3
R13477 commonsourceibias.n396 commonsourceibias.n268 161.3
R13478 commonsourceibias.n394 commonsourceibias.n393 161.3
R13479 commonsourceibias.n392 commonsourceibias.n269 161.3
R13480 commonsourceibias.n391 commonsourceibias.n390 161.3
R13481 commonsourceibias.n388 commonsourceibias.n270 161.3
R13482 commonsourceibias.n387 commonsourceibias.n386 161.3
R13483 commonsourceibias.n385 commonsourceibias.n271 161.3
R13484 commonsourceibias.n384 commonsourceibias.n383 161.3
R13485 commonsourceibias.n381 commonsourceibias.n272 161.3
R13486 commonsourceibias.n379 commonsourceibias.n378 161.3
R13487 commonsourceibias.n528 commonsourceibias.n468 161.3
R13488 commonsourceibias.n527 commonsourceibias.n526 161.3
R13489 commonsourceibias.n525 commonsourceibias.n524 161.3
R13490 commonsourceibias.n523 commonsourceibias.n470 161.3
R13491 commonsourceibias.n521 commonsourceibias.n520 161.3
R13492 commonsourceibias.n519 commonsourceibias.n471 161.3
R13493 commonsourceibias.n518 commonsourceibias.n517 161.3
R13494 commonsourceibias.n515 commonsourceibias.n472 161.3
R13495 commonsourceibias.n514 commonsourceibias.n513 161.3
R13496 commonsourceibias.n512 commonsourceibias.n473 161.3
R13497 commonsourceibias.n511 commonsourceibias.n510 161.3
R13498 commonsourceibias.n508 commonsourceibias.n474 161.3
R13499 commonsourceibias.n506 commonsourceibias.n505 161.3
R13500 commonsourceibias.n504 commonsourceibias.n475 161.3
R13501 commonsourceibias.n503 commonsourceibias.n502 161.3
R13502 commonsourceibias.n500 commonsourceibias.n476 161.3
R13503 commonsourceibias.n499 commonsourceibias.n498 161.3
R13504 commonsourceibias.n497 commonsourceibias.n496 161.3
R13505 commonsourceibias.n495 commonsourceibias.n478 161.3
R13506 commonsourceibias.n494 commonsourceibias.n493 161.3
R13507 commonsourceibias.n492 commonsourceibias.n491 161.3
R13508 commonsourceibias.n490 commonsourceibias.n480 161.3
R13509 commonsourceibias.n489 commonsourceibias.n488 161.3
R13510 commonsourceibias.n487 commonsourceibias.n486 161.3
R13511 commonsourceibias.n485 commonsourceibias.n482 161.3
R13512 commonsourceibias.n464 commonsourceibias.n404 161.3
R13513 commonsourceibias.n463 commonsourceibias.n462 161.3
R13514 commonsourceibias.n461 commonsourceibias.n460 161.3
R13515 commonsourceibias.n459 commonsourceibias.n406 161.3
R13516 commonsourceibias.n457 commonsourceibias.n456 161.3
R13517 commonsourceibias.n455 commonsourceibias.n407 161.3
R13518 commonsourceibias.n454 commonsourceibias.n453 161.3
R13519 commonsourceibias.n451 commonsourceibias.n408 161.3
R13520 commonsourceibias.n450 commonsourceibias.n449 161.3
R13521 commonsourceibias.n448 commonsourceibias.n409 161.3
R13522 commonsourceibias.n447 commonsourceibias.n446 161.3
R13523 commonsourceibias.n444 commonsourceibias.n410 161.3
R13524 commonsourceibias.n442 commonsourceibias.n441 161.3
R13525 commonsourceibias.n440 commonsourceibias.n411 161.3
R13526 commonsourceibias.n439 commonsourceibias.n438 161.3
R13527 commonsourceibias.n436 commonsourceibias.n412 161.3
R13528 commonsourceibias.n435 commonsourceibias.n434 161.3
R13529 commonsourceibias.n433 commonsourceibias.n432 161.3
R13530 commonsourceibias.n431 commonsourceibias.n414 161.3
R13531 commonsourceibias.n430 commonsourceibias.n429 161.3
R13532 commonsourceibias.n428 commonsourceibias.n427 161.3
R13533 commonsourceibias.n426 commonsourceibias.n416 161.3
R13534 commonsourceibias.n425 commonsourceibias.n424 161.3
R13535 commonsourceibias.n423 commonsourceibias.n422 161.3
R13536 commonsourceibias.n421 commonsourceibias.n418 161.3
R13537 commonsourceibias.n80 commonsourceibias.n78 81.5057
R13538 commonsourceibias.n304 commonsourceibias.n302 81.5057
R13539 commonsourceibias.n80 commonsourceibias.n79 80.9324
R13540 commonsourceibias.n82 commonsourceibias.n81 80.9324
R13541 commonsourceibias.n77 commonsourceibias.n76 80.9324
R13542 commonsourceibias.n75 commonsourceibias.n74 80.9324
R13543 commonsourceibias.n73 commonsourceibias.n72 80.9324
R13544 commonsourceibias.n371 commonsourceibias.n370 80.9324
R13545 commonsourceibias.n373 commonsourceibias.n372 80.9324
R13546 commonsourceibias.n375 commonsourceibias.n374 80.9324
R13547 commonsourceibias.n306 commonsourceibias.n305 80.9324
R13548 commonsourceibias.n304 commonsourceibias.n303 80.9324
R13549 commonsourceibias.n71 commonsourceibias.n70 80.6037
R13550 commonsourceibias.n137 commonsourceibias.n136 80.6037
R13551 commonsourceibias.n264 commonsourceibias.n263 80.6037
R13552 commonsourceibias.n200 commonsourceibias.n199 80.6037
R13553 commonsourceibias.n369 commonsourceibias.n368 80.6037
R13554 commonsourceibias.n403 commonsourceibias.n402 80.6037
R13555 commonsourceibias.n530 commonsourceibias.n529 80.6037
R13556 commonsourceibias.n466 commonsourceibias.n465 80.6037
R13557 commonsourceibias.n65 commonsourceibias.n64 56.5617
R13558 commonsourceibias.n51 commonsourceibias.n50 56.5617
R13559 commonsourceibias.n42 commonsourceibias.n41 56.5617
R13560 commonsourceibias.n28 commonsourceibias.n27 56.5617
R13561 commonsourceibias.n131 commonsourceibias.n130 56.5617
R13562 commonsourceibias.n117 commonsourceibias.n116 56.5617
R13563 commonsourceibias.n108 commonsourceibias.n107 56.5617
R13564 commonsourceibias.n94 commonsourceibias.n93 56.5617
R13565 commonsourceibias.n221 commonsourceibias.n220 56.5617
R13566 commonsourceibias.n235 commonsourceibias.n234 56.5617
R13567 commonsourceibias.n244 commonsourceibias.n243 56.5617
R13568 commonsourceibias.n258 commonsourceibias.n257 56.5617
R13569 commonsourceibias.n194 commonsourceibias.n193 56.5617
R13570 commonsourceibias.n180 commonsourceibias.n179 56.5617
R13571 commonsourceibias.n171 commonsourceibias.n170 56.5617
R13572 commonsourceibias.n157 commonsourceibias.n156 56.5617
R13573 commonsourceibias.n325 commonsourceibias.n324 56.5617
R13574 commonsourceibias.n339 commonsourceibias.n338 56.5617
R13575 commonsourceibias.n349 commonsourceibias.n347 56.5617
R13576 commonsourceibias.n363 commonsourceibias.n362 56.5617
R13577 commonsourceibias.n397 commonsourceibias.n396 56.5617
R13578 commonsourceibias.n383 commonsourceibias.n381 56.5617
R13579 commonsourceibias.n284 commonsourceibias.n283 56.5617
R13580 commonsourceibias.n298 commonsourceibias.n297 56.5617
R13581 commonsourceibias.n486 commonsourceibias.n485 56.5617
R13582 commonsourceibias.n500 commonsourceibias.n499 56.5617
R13583 commonsourceibias.n510 commonsourceibias.n508 56.5617
R13584 commonsourceibias.n524 commonsourceibias.n523 56.5617
R13585 commonsourceibias.n422 commonsourceibias.n421 56.5617
R13586 commonsourceibias.n436 commonsourceibias.n435 56.5617
R13587 commonsourceibias.n446 commonsourceibias.n444 56.5617
R13588 commonsourceibias.n460 commonsourceibias.n459 56.5617
R13589 commonsourceibias.n56 commonsourceibias.n55 56.0773
R13590 commonsourceibias.n37 commonsourceibias.n36 56.0773
R13591 commonsourceibias.n122 commonsourceibias.n121 56.0773
R13592 commonsourceibias.n103 commonsourceibias.n102 56.0773
R13593 commonsourceibias.n230 commonsourceibias.n229 56.0773
R13594 commonsourceibias.n249 commonsourceibias.n248 56.0773
R13595 commonsourceibias.n185 commonsourceibias.n184 56.0773
R13596 commonsourceibias.n166 commonsourceibias.n165 56.0773
R13597 commonsourceibias.n334 commonsourceibias.n333 56.0773
R13598 commonsourceibias.n354 commonsourceibias.n353 56.0773
R13599 commonsourceibias.n388 commonsourceibias.n387 56.0773
R13600 commonsourceibias.n293 commonsourceibias.n292 56.0773
R13601 commonsourceibias.n495 commonsourceibias.n494 56.0773
R13602 commonsourceibias.n515 commonsourceibias.n514 56.0773
R13603 commonsourceibias.n431 commonsourceibias.n430 56.0773
R13604 commonsourceibias.n451 commonsourceibias.n450 56.0773
R13605 commonsourceibias.n70 commonsourceibias.n69 46.0096
R13606 commonsourceibias.n136 commonsourceibias.n135 46.0096
R13607 commonsourceibias.n263 commonsourceibias.n262 46.0096
R13608 commonsourceibias.n199 commonsourceibias.n198 46.0096
R13609 commonsourceibias.n368 commonsourceibias.n367 46.0096
R13610 commonsourceibias.n402 commonsourceibias.n401 46.0096
R13611 commonsourceibias.n529 commonsourceibias.n528 46.0096
R13612 commonsourceibias.n465 commonsourceibias.n464 46.0096
R13613 commonsourceibias.n58 commonsourceibias.n12 41.5458
R13614 commonsourceibias.n33 commonsourceibias.n32 41.5458
R13615 commonsourceibias.n124 commonsourceibias.n3 41.5458
R13616 commonsourceibias.n99 commonsourceibias.n98 41.5458
R13617 commonsourceibias.n226 commonsourceibias.n225 41.5458
R13618 commonsourceibias.n251 commonsourceibias.n205 41.5458
R13619 commonsourceibias.n187 commonsourceibias.n141 41.5458
R13620 commonsourceibias.n162 commonsourceibias.n161 41.5458
R13621 commonsourceibias.n330 commonsourceibias.n329 41.5458
R13622 commonsourceibias.n356 commonsourceibias.n310 41.5458
R13623 commonsourceibias.n390 commonsourceibias.n269 41.5458
R13624 commonsourceibias.n289 commonsourceibias.n288 41.5458
R13625 commonsourceibias.n491 commonsourceibias.n490 41.5458
R13626 commonsourceibias.n517 commonsourceibias.n471 41.5458
R13627 commonsourceibias.n427 commonsourceibias.n426 41.5458
R13628 commonsourceibias.n453 commonsourceibias.n407 41.5458
R13629 commonsourceibias.n48 commonsourceibias.n17 40.577
R13630 commonsourceibias.n44 commonsourceibias.n17 40.577
R13631 commonsourceibias.n114 commonsourceibias.n8 40.577
R13632 commonsourceibias.n110 commonsourceibias.n8 40.577
R13633 commonsourceibias.n237 commonsourceibias.n210 40.577
R13634 commonsourceibias.n241 commonsourceibias.n210 40.577
R13635 commonsourceibias.n177 commonsourceibias.n146 40.577
R13636 commonsourceibias.n173 commonsourceibias.n146 40.577
R13637 commonsourceibias.n341 commonsourceibias.n314 40.577
R13638 commonsourceibias.n345 commonsourceibias.n314 40.577
R13639 commonsourceibias.n379 commonsourceibias.n273 40.577
R13640 commonsourceibias.n300 commonsourceibias.n273 40.577
R13641 commonsourceibias.n502 commonsourceibias.n475 40.577
R13642 commonsourceibias.n506 commonsourceibias.n475 40.577
R13643 commonsourceibias.n438 commonsourceibias.n411 40.577
R13644 commonsourceibias.n442 commonsourceibias.n411 40.577
R13645 commonsourceibias.n62 commonsourceibias.n12 39.6083
R13646 commonsourceibias.n32 commonsourceibias.n31 39.6083
R13647 commonsourceibias.n128 commonsourceibias.n3 39.6083
R13648 commonsourceibias.n98 commonsourceibias.n97 39.6083
R13649 commonsourceibias.n225 commonsourceibias.n224 39.6083
R13650 commonsourceibias.n255 commonsourceibias.n205 39.6083
R13651 commonsourceibias.n191 commonsourceibias.n141 39.6083
R13652 commonsourceibias.n161 commonsourceibias.n160 39.6083
R13653 commonsourceibias.n329 commonsourceibias.n328 39.6083
R13654 commonsourceibias.n360 commonsourceibias.n310 39.6083
R13655 commonsourceibias.n394 commonsourceibias.n269 39.6083
R13656 commonsourceibias.n288 commonsourceibias.n287 39.6083
R13657 commonsourceibias.n490 commonsourceibias.n489 39.6083
R13658 commonsourceibias.n521 commonsourceibias.n471 39.6083
R13659 commonsourceibias.n426 commonsourceibias.n425 39.6083
R13660 commonsourceibias.n457 commonsourceibias.n407 39.6083
R13661 commonsourceibias.n26 commonsourceibias.n25 33.0515
R13662 commonsourceibias.n92 commonsourceibias.n91 33.0515
R13663 commonsourceibias.n155 commonsourceibias.n154 33.0515
R13664 commonsourceibias.n219 commonsourceibias.n218 33.0515
R13665 commonsourceibias.n323 commonsourceibias.n322 33.0515
R13666 commonsourceibias.n282 commonsourceibias.n281 33.0515
R13667 commonsourceibias.n484 commonsourceibias.n483 33.0515
R13668 commonsourceibias.n420 commonsourceibias.n419 33.0515
R13669 commonsourceibias.n25 commonsourceibias.n24 28.5514
R13670 commonsourceibias.n91 commonsourceibias.n90 28.5514
R13671 commonsourceibias.n218 commonsourceibias.n217 28.5514
R13672 commonsourceibias.n154 commonsourceibias.n153 28.5514
R13673 commonsourceibias.n322 commonsourceibias.n321 28.5514
R13674 commonsourceibias.n281 commonsourceibias.n280 28.5514
R13675 commonsourceibias.n483 commonsourceibias.n482 28.5514
R13676 commonsourceibias.n419 commonsourceibias.n418 28.5514
R13677 commonsourceibias.n69 commonsourceibias.n68 26.0455
R13678 commonsourceibias.n135 commonsourceibias.n134 26.0455
R13679 commonsourceibias.n262 commonsourceibias.n261 26.0455
R13680 commonsourceibias.n198 commonsourceibias.n197 26.0455
R13681 commonsourceibias.n367 commonsourceibias.n366 26.0455
R13682 commonsourceibias.n401 commonsourceibias.n400 26.0455
R13683 commonsourceibias.n528 commonsourceibias.n527 26.0455
R13684 commonsourceibias.n464 commonsourceibias.n463 26.0455
R13685 commonsourceibias.n55 commonsourceibias.n14 25.0767
R13686 commonsourceibias.n38 commonsourceibias.n37 25.0767
R13687 commonsourceibias.n121 commonsourceibias.n5 25.0767
R13688 commonsourceibias.n104 commonsourceibias.n103 25.0767
R13689 commonsourceibias.n231 commonsourceibias.n230 25.0767
R13690 commonsourceibias.n248 commonsourceibias.n207 25.0767
R13691 commonsourceibias.n184 commonsourceibias.n143 25.0767
R13692 commonsourceibias.n167 commonsourceibias.n166 25.0767
R13693 commonsourceibias.n335 commonsourceibias.n334 25.0767
R13694 commonsourceibias.n353 commonsourceibias.n312 25.0767
R13695 commonsourceibias.n387 commonsourceibias.n271 25.0767
R13696 commonsourceibias.n294 commonsourceibias.n293 25.0767
R13697 commonsourceibias.n496 commonsourceibias.n495 25.0767
R13698 commonsourceibias.n514 commonsourceibias.n473 25.0767
R13699 commonsourceibias.n432 commonsourceibias.n431 25.0767
R13700 commonsourceibias.n450 commonsourceibias.n409 25.0767
R13701 commonsourceibias.n51 commonsourceibias.n16 24.3464
R13702 commonsourceibias.n41 commonsourceibias.n19 24.3464
R13703 commonsourceibias.n117 commonsourceibias.n7 24.3464
R13704 commonsourceibias.n107 commonsourceibias.n85 24.3464
R13705 commonsourceibias.n234 commonsourceibias.n212 24.3464
R13706 commonsourceibias.n244 commonsourceibias.n209 24.3464
R13707 commonsourceibias.n180 commonsourceibias.n145 24.3464
R13708 commonsourceibias.n170 commonsourceibias.n148 24.3464
R13709 commonsourceibias.n338 commonsourceibias.n316 24.3464
R13710 commonsourceibias.n349 commonsourceibias.n348 24.3464
R13711 commonsourceibias.n383 commonsourceibias.n382 24.3464
R13712 commonsourceibias.n297 commonsourceibias.n275 24.3464
R13713 commonsourceibias.n499 commonsourceibias.n477 24.3464
R13714 commonsourceibias.n510 commonsourceibias.n509 24.3464
R13715 commonsourceibias.n435 commonsourceibias.n413 24.3464
R13716 commonsourceibias.n446 commonsourceibias.n445 24.3464
R13717 commonsourceibias.n65 commonsourceibias.n10 23.8546
R13718 commonsourceibias.n27 commonsourceibias.n26 23.8546
R13719 commonsourceibias.n131 commonsourceibias.n1 23.8546
R13720 commonsourceibias.n93 commonsourceibias.n92 23.8546
R13721 commonsourceibias.n220 commonsourceibias.n219 23.8546
R13722 commonsourceibias.n258 commonsourceibias.n203 23.8546
R13723 commonsourceibias.n194 commonsourceibias.n139 23.8546
R13724 commonsourceibias.n156 commonsourceibias.n155 23.8546
R13725 commonsourceibias.n324 commonsourceibias.n323 23.8546
R13726 commonsourceibias.n363 commonsourceibias.n308 23.8546
R13727 commonsourceibias.n397 commonsourceibias.n267 23.8546
R13728 commonsourceibias.n283 commonsourceibias.n282 23.8546
R13729 commonsourceibias.n485 commonsourceibias.n484 23.8546
R13730 commonsourceibias.n524 commonsourceibias.n469 23.8546
R13731 commonsourceibias.n421 commonsourceibias.n420 23.8546
R13732 commonsourceibias.n460 commonsourceibias.n405 23.8546
R13733 commonsourceibias.n64 commonsourceibias.n63 16.9689
R13734 commonsourceibias.n28 commonsourceibias.n23 16.9689
R13735 commonsourceibias.n130 commonsourceibias.n129 16.9689
R13736 commonsourceibias.n94 commonsourceibias.n89 16.9689
R13737 commonsourceibias.n221 commonsourceibias.n216 16.9689
R13738 commonsourceibias.n257 commonsourceibias.n256 16.9689
R13739 commonsourceibias.n193 commonsourceibias.n192 16.9689
R13740 commonsourceibias.n157 commonsourceibias.n152 16.9689
R13741 commonsourceibias.n325 commonsourceibias.n320 16.9689
R13742 commonsourceibias.n362 commonsourceibias.n361 16.9689
R13743 commonsourceibias.n396 commonsourceibias.n395 16.9689
R13744 commonsourceibias.n284 commonsourceibias.n279 16.9689
R13745 commonsourceibias.n486 commonsourceibias.n481 16.9689
R13746 commonsourceibias.n523 commonsourceibias.n522 16.9689
R13747 commonsourceibias.n422 commonsourceibias.n417 16.9689
R13748 commonsourceibias.n459 commonsourceibias.n458 16.9689
R13749 commonsourceibias.n50 commonsourceibias.n49 16.477
R13750 commonsourceibias.n43 commonsourceibias.n42 16.477
R13751 commonsourceibias.n116 commonsourceibias.n115 16.477
R13752 commonsourceibias.n109 commonsourceibias.n108 16.477
R13753 commonsourceibias.n236 commonsourceibias.n235 16.477
R13754 commonsourceibias.n243 commonsourceibias.n242 16.477
R13755 commonsourceibias.n179 commonsourceibias.n178 16.477
R13756 commonsourceibias.n172 commonsourceibias.n171 16.477
R13757 commonsourceibias.n340 commonsourceibias.n339 16.477
R13758 commonsourceibias.n347 commonsourceibias.n346 16.477
R13759 commonsourceibias.n381 commonsourceibias.n380 16.477
R13760 commonsourceibias.n299 commonsourceibias.n298 16.477
R13761 commonsourceibias.n501 commonsourceibias.n500 16.477
R13762 commonsourceibias.n508 commonsourceibias.n507 16.477
R13763 commonsourceibias.n437 commonsourceibias.n436 16.477
R13764 commonsourceibias.n444 commonsourceibias.n443 16.477
R13765 commonsourceibias.n57 commonsourceibias.n56 15.9852
R13766 commonsourceibias.n36 commonsourceibias.n21 15.9852
R13767 commonsourceibias.n123 commonsourceibias.n122 15.9852
R13768 commonsourceibias.n102 commonsourceibias.n87 15.9852
R13769 commonsourceibias.n229 commonsourceibias.n214 15.9852
R13770 commonsourceibias.n250 commonsourceibias.n249 15.9852
R13771 commonsourceibias.n186 commonsourceibias.n185 15.9852
R13772 commonsourceibias.n165 commonsourceibias.n150 15.9852
R13773 commonsourceibias.n333 commonsourceibias.n318 15.9852
R13774 commonsourceibias.n355 commonsourceibias.n354 15.9852
R13775 commonsourceibias.n389 commonsourceibias.n388 15.9852
R13776 commonsourceibias.n292 commonsourceibias.n277 15.9852
R13777 commonsourceibias.n494 commonsourceibias.n479 15.9852
R13778 commonsourceibias.n516 commonsourceibias.n515 15.9852
R13779 commonsourceibias.n430 commonsourceibias.n415 15.9852
R13780 commonsourceibias.n452 commonsourceibias.n451 15.9852
R13781 commonsourceibias.n73 commonsourceibias.n71 13.2057
R13782 commonsourceibias.n371 commonsourceibias.n369 13.2057
R13783 commonsourceibias.n532 commonsourceibias.n265 10.4122
R13784 commonsourceibias.n112 commonsourceibias.n83 9.50363
R13785 commonsourceibias.n377 commonsourceibias.n376 9.50363
R13786 commonsourceibias.n201 commonsourceibias.n137 8.7339
R13787 commonsourceibias.n467 commonsourceibias.n403 8.7339
R13788 commonsourceibias.n58 commonsourceibias.n57 8.60764
R13789 commonsourceibias.n33 commonsourceibias.n21 8.60764
R13790 commonsourceibias.n124 commonsourceibias.n123 8.60764
R13791 commonsourceibias.n99 commonsourceibias.n87 8.60764
R13792 commonsourceibias.n226 commonsourceibias.n214 8.60764
R13793 commonsourceibias.n251 commonsourceibias.n250 8.60764
R13794 commonsourceibias.n187 commonsourceibias.n186 8.60764
R13795 commonsourceibias.n162 commonsourceibias.n150 8.60764
R13796 commonsourceibias.n330 commonsourceibias.n318 8.60764
R13797 commonsourceibias.n356 commonsourceibias.n355 8.60764
R13798 commonsourceibias.n390 commonsourceibias.n389 8.60764
R13799 commonsourceibias.n289 commonsourceibias.n277 8.60764
R13800 commonsourceibias.n491 commonsourceibias.n479 8.60764
R13801 commonsourceibias.n517 commonsourceibias.n516 8.60764
R13802 commonsourceibias.n427 commonsourceibias.n415 8.60764
R13803 commonsourceibias.n453 commonsourceibias.n452 8.60764
R13804 commonsourceibias.n532 commonsourceibias.n531 8.46921
R13805 commonsourceibias.n49 commonsourceibias.n48 8.11581
R13806 commonsourceibias.n44 commonsourceibias.n43 8.11581
R13807 commonsourceibias.n115 commonsourceibias.n114 8.11581
R13808 commonsourceibias.n110 commonsourceibias.n109 8.11581
R13809 commonsourceibias.n237 commonsourceibias.n236 8.11581
R13810 commonsourceibias.n242 commonsourceibias.n241 8.11581
R13811 commonsourceibias.n178 commonsourceibias.n177 8.11581
R13812 commonsourceibias.n173 commonsourceibias.n172 8.11581
R13813 commonsourceibias.n341 commonsourceibias.n340 8.11581
R13814 commonsourceibias.n346 commonsourceibias.n345 8.11581
R13815 commonsourceibias.n380 commonsourceibias.n379 8.11581
R13816 commonsourceibias.n300 commonsourceibias.n299 8.11581
R13817 commonsourceibias.n502 commonsourceibias.n501 8.11581
R13818 commonsourceibias.n507 commonsourceibias.n506 8.11581
R13819 commonsourceibias.n438 commonsourceibias.n437 8.11581
R13820 commonsourceibias.n443 commonsourceibias.n442 8.11581
R13821 commonsourceibias.n63 commonsourceibias.n62 7.62397
R13822 commonsourceibias.n31 commonsourceibias.n23 7.62397
R13823 commonsourceibias.n129 commonsourceibias.n128 7.62397
R13824 commonsourceibias.n97 commonsourceibias.n89 7.62397
R13825 commonsourceibias.n224 commonsourceibias.n216 7.62397
R13826 commonsourceibias.n256 commonsourceibias.n255 7.62397
R13827 commonsourceibias.n192 commonsourceibias.n191 7.62397
R13828 commonsourceibias.n160 commonsourceibias.n152 7.62397
R13829 commonsourceibias.n328 commonsourceibias.n320 7.62397
R13830 commonsourceibias.n361 commonsourceibias.n360 7.62397
R13831 commonsourceibias.n395 commonsourceibias.n394 7.62397
R13832 commonsourceibias.n287 commonsourceibias.n279 7.62397
R13833 commonsourceibias.n489 commonsourceibias.n481 7.62397
R13834 commonsourceibias.n522 commonsourceibias.n521 7.62397
R13835 commonsourceibias.n425 commonsourceibias.n417 7.62397
R13836 commonsourceibias.n458 commonsourceibias.n457 7.62397
R13837 commonsourceibias.n265 commonsourceibias.n264 5.00473
R13838 commonsourceibias.n201 commonsourceibias.n200 5.00473
R13839 commonsourceibias.n531 commonsourceibias.n530 5.00473
R13840 commonsourceibias.n467 commonsourceibias.n466 5.00473
R13841 commonsourceibias commonsourceibias.n532 3.87639
R13842 commonsourceibias.n265 commonsourceibias.n201 3.72967
R13843 commonsourceibias.n531 commonsourceibias.n467 3.72967
R13844 commonsourceibias.n78 commonsourceibias.t7 2.82907
R13845 commonsourceibias.n78 commonsourceibias.t35 2.82907
R13846 commonsourceibias.n79 commonsourceibias.t25 2.82907
R13847 commonsourceibias.n79 commonsourceibias.t45 2.82907
R13848 commonsourceibias.n81 commonsourceibias.t33 2.82907
R13849 commonsourceibias.n81 commonsourceibias.t41 2.82907
R13850 commonsourceibias.n76 commonsourceibias.t43 2.82907
R13851 commonsourceibias.n76 commonsourceibias.t19 2.82907
R13852 commonsourceibias.n74 commonsourceibias.t3 2.82907
R13853 commonsourceibias.n74 commonsourceibias.t23 2.82907
R13854 commonsourceibias.n72 commonsourceibias.t17 2.82907
R13855 commonsourceibias.n72 commonsourceibias.t31 2.82907
R13856 commonsourceibias.n370 commonsourceibias.t47 2.82907
R13857 commonsourceibias.n370 commonsourceibias.t27 2.82907
R13858 commonsourceibias.n372 commonsourceibias.t37 2.82907
R13859 commonsourceibias.n372 commonsourceibias.t21 2.82907
R13860 commonsourceibias.n374 commonsourceibias.t29 2.82907
R13861 commonsourceibias.n374 commonsourceibias.t11 2.82907
R13862 commonsourceibias.n305 commonsourceibias.t9 2.82907
R13863 commonsourceibias.n305 commonsourceibias.t1 2.82907
R13864 commonsourceibias.n303 commonsourceibias.t13 2.82907
R13865 commonsourceibias.n303 commonsourceibias.t39 2.82907
R13866 commonsourceibias.n302 commonsourceibias.t5 2.82907
R13867 commonsourceibias.n302 commonsourceibias.t15 2.82907
R13868 commonsourceibias.n68 commonsourceibias.n10 0.738255
R13869 commonsourceibias.n134 commonsourceibias.n1 0.738255
R13870 commonsourceibias.n261 commonsourceibias.n203 0.738255
R13871 commonsourceibias.n197 commonsourceibias.n139 0.738255
R13872 commonsourceibias.n366 commonsourceibias.n308 0.738255
R13873 commonsourceibias.n400 commonsourceibias.n267 0.738255
R13874 commonsourceibias.n527 commonsourceibias.n469 0.738255
R13875 commonsourceibias.n463 commonsourceibias.n405 0.738255
R13876 commonsourceibias.n75 commonsourceibias.n73 0.573776
R13877 commonsourceibias.n77 commonsourceibias.n75 0.573776
R13878 commonsourceibias.n82 commonsourceibias.n80 0.573776
R13879 commonsourceibias.n306 commonsourceibias.n304 0.573776
R13880 commonsourceibias.n375 commonsourceibias.n373 0.573776
R13881 commonsourceibias.n373 commonsourceibias.n371 0.573776
R13882 commonsourceibias.n83 commonsourceibias.n77 0.287138
R13883 commonsourceibias.n83 commonsourceibias.n82 0.287138
R13884 commonsourceibias.n376 commonsourceibias.n306 0.287138
R13885 commonsourceibias.n376 commonsourceibias.n375 0.287138
R13886 commonsourceibias.n71 commonsourceibias.n9 0.285035
R13887 commonsourceibias.n137 commonsourceibias.n0 0.285035
R13888 commonsourceibias.n264 commonsourceibias.n202 0.285035
R13889 commonsourceibias.n200 commonsourceibias.n138 0.285035
R13890 commonsourceibias.n369 commonsourceibias.n307 0.285035
R13891 commonsourceibias.n403 commonsourceibias.n266 0.285035
R13892 commonsourceibias.n530 commonsourceibias.n468 0.285035
R13893 commonsourceibias.n466 commonsourceibias.n404 0.285035
R13894 commonsourceibias.n16 commonsourceibias.n14 0.246418
R13895 commonsourceibias.n38 commonsourceibias.n19 0.246418
R13896 commonsourceibias.n7 commonsourceibias.n5 0.246418
R13897 commonsourceibias.n104 commonsourceibias.n85 0.246418
R13898 commonsourceibias.n231 commonsourceibias.n212 0.246418
R13899 commonsourceibias.n209 commonsourceibias.n207 0.246418
R13900 commonsourceibias.n145 commonsourceibias.n143 0.246418
R13901 commonsourceibias.n167 commonsourceibias.n148 0.246418
R13902 commonsourceibias.n335 commonsourceibias.n316 0.246418
R13903 commonsourceibias.n348 commonsourceibias.n312 0.246418
R13904 commonsourceibias.n382 commonsourceibias.n271 0.246418
R13905 commonsourceibias.n294 commonsourceibias.n275 0.246418
R13906 commonsourceibias.n496 commonsourceibias.n477 0.246418
R13907 commonsourceibias.n509 commonsourceibias.n473 0.246418
R13908 commonsourceibias.n432 commonsourceibias.n413 0.246418
R13909 commonsourceibias.n445 commonsourceibias.n409 0.246418
R13910 commonsourceibias.n67 commonsourceibias.n9 0.189894
R13911 commonsourceibias.n67 commonsourceibias.n66 0.189894
R13912 commonsourceibias.n66 commonsourceibias.n11 0.189894
R13913 commonsourceibias.n61 commonsourceibias.n11 0.189894
R13914 commonsourceibias.n61 commonsourceibias.n60 0.189894
R13915 commonsourceibias.n60 commonsourceibias.n59 0.189894
R13916 commonsourceibias.n59 commonsourceibias.n13 0.189894
R13917 commonsourceibias.n54 commonsourceibias.n13 0.189894
R13918 commonsourceibias.n54 commonsourceibias.n53 0.189894
R13919 commonsourceibias.n53 commonsourceibias.n52 0.189894
R13920 commonsourceibias.n52 commonsourceibias.n15 0.189894
R13921 commonsourceibias.n47 commonsourceibias.n15 0.189894
R13922 commonsourceibias.n47 commonsourceibias.n46 0.189894
R13923 commonsourceibias.n46 commonsourceibias.n45 0.189894
R13924 commonsourceibias.n45 commonsourceibias.n18 0.189894
R13925 commonsourceibias.n40 commonsourceibias.n18 0.189894
R13926 commonsourceibias.n40 commonsourceibias.n39 0.189894
R13927 commonsourceibias.n39 commonsourceibias.n20 0.189894
R13928 commonsourceibias.n35 commonsourceibias.n20 0.189894
R13929 commonsourceibias.n35 commonsourceibias.n34 0.189894
R13930 commonsourceibias.n34 commonsourceibias.n22 0.189894
R13931 commonsourceibias.n30 commonsourceibias.n22 0.189894
R13932 commonsourceibias.n30 commonsourceibias.n29 0.189894
R13933 commonsourceibias.n29 commonsourceibias.n24 0.189894
R13934 commonsourceibias.n111 commonsourceibias.n84 0.189894
R13935 commonsourceibias.n106 commonsourceibias.n84 0.189894
R13936 commonsourceibias.n106 commonsourceibias.n105 0.189894
R13937 commonsourceibias.n105 commonsourceibias.n86 0.189894
R13938 commonsourceibias.n101 commonsourceibias.n86 0.189894
R13939 commonsourceibias.n101 commonsourceibias.n100 0.189894
R13940 commonsourceibias.n100 commonsourceibias.n88 0.189894
R13941 commonsourceibias.n96 commonsourceibias.n88 0.189894
R13942 commonsourceibias.n96 commonsourceibias.n95 0.189894
R13943 commonsourceibias.n95 commonsourceibias.n90 0.189894
R13944 commonsourceibias.n133 commonsourceibias.n0 0.189894
R13945 commonsourceibias.n133 commonsourceibias.n132 0.189894
R13946 commonsourceibias.n132 commonsourceibias.n2 0.189894
R13947 commonsourceibias.n127 commonsourceibias.n2 0.189894
R13948 commonsourceibias.n127 commonsourceibias.n126 0.189894
R13949 commonsourceibias.n126 commonsourceibias.n125 0.189894
R13950 commonsourceibias.n125 commonsourceibias.n4 0.189894
R13951 commonsourceibias.n120 commonsourceibias.n4 0.189894
R13952 commonsourceibias.n120 commonsourceibias.n119 0.189894
R13953 commonsourceibias.n119 commonsourceibias.n118 0.189894
R13954 commonsourceibias.n118 commonsourceibias.n6 0.189894
R13955 commonsourceibias.n113 commonsourceibias.n6 0.189894
R13956 commonsourceibias.n260 commonsourceibias.n202 0.189894
R13957 commonsourceibias.n260 commonsourceibias.n259 0.189894
R13958 commonsourceibias.n259 commonsourceibias.n204 0.189894
R13959 commonsourceibias.n254 commonsourceibias.n204 0.189894
R13960 commonsourceibias.n254 commonsourceibias.n253 0.189894
R13961 commonsourceibias.n253 commonsourceibias.n252 0.189894
R13962 commonsourceibias.n252 commonsourceibias.n206 0.189894
R13963 commonsourceibias.n247 commonsourceibias.n206 0.189894
R13964 commonsourceibias.n247 commonsourceibias.n246 0.189894
R13965 commonsourceibias.n246 commonsourceibias.n245 0.189894
R13966 commonsourceibias.n245 commonsourceibias.n208 0.189894
R13967 commonsourceibias.n240 commonsourceibias.n208 0.189894
R13968 commonsourceibias.n240 commonsourceibias.n239 0.189894
R13969 commonsourceibias.n239 commonsourceibias.n238 0.189894
R13970 commonsourceibias.n238 commonsourceibias.n211 0.189894
R13971 commonsourceibias.n233 commonsourceibias.n211 0.189894
R13972 commonsourceibias.n233 commonsourceibias.n232 0.189894
R13973 commonsourceibias.n232 commonsourceibias.n213 0.189894
R13974 commonsourceibias.n228 commonsourceibias.n213 0.189894
R13975 commonsourceibias.n228 commonsourceibias.n227 0.189894
R13976 commonsourceibias.n227 commonsourceibias.n215 0.189894
R13977 commonsourceibias.n223 commonsourceibias.n215 0.189894
R13978 commonsourceibias.n223 commonsourceibias.n222 0.189894
R13979 commonsourceibias.n222 commonsourceibias.n217 0.189894
R13980 commonsourceibias.n196 commonsourceibias.n138 0.189894
R13981 commonsourceibias.n196 commonsourceibias.n195 0.189894
R13982 commonsourceibias.n195 commonsourceibias.n140 0.189894
R13983 commonsourceibias.n190 commonsourceibias.n140 0.189894
R13984 commonsourceibias.n190 commonsourceibias.n189 0.189894
R13985 commonsourceibias.n189 commonsourceibias.n188 0.189894
R13986 commonsourceibias.n188 commonsourceibias.n142 0.189894
R13987 commonsourceibias.n183 commonsourceibias.n142 0.189894
R13988 commonsourceibias.n183 commonsourceibias.n182 0.189894
R13989 commonsourceibias.n182 commonsourceibias.n181 0.189894
R13990 commonsourceibias.n181 commonsourceibias.n144 0.189894
R13991 commonsourceibias.n176 commonsourceibias.n144 0.189894
R13992 commonsourceibias.n176 commonsourceibias.n175 0.189894
R13993 commonsourceibias.n175 commonsourceibias.n174 0.189894
R13994 commonsourceibias.n174 commonsourceibias.n147 0.189894
R13995 commonsourceibias.n169 commonsourceibias.n147 0.189894
R13996 commonsourceibias.n169 commonsourceibias.n168 0.189894
R13997 commonsourceibias.n168 commonsourceibias.n149 0.189894
R13998 commonsourceibias.n164 commonsourceibias.n149 0.189894
R13999 commonsourceibias.n164 commonsourceibias.n163 0.189894
R14000 commonsourceibias.n163 commonsourceibias.n151 0.189894
R14001 commonsourceibias.n159 commonsourceibias.n151 0.189894
R14002 commonsourceibias.n159 commonsourceibias.n158 0.189894
R14003 commonsourceibias.n158 commonsourceibias.n153 0.189894
R14004 commonsourceibias.n326 commonsourceibias.n321 0.189894
R14005 commonsourceibias.n327 commonsourceibias.n326 0.189894
R14006 commonsourceibias.n327 commonsourceibias.n319 0.189894
R14007 commonsourceibias.n331 commonsourceibias.n319 0.189894
R14008 commonsourceibias.n332 commonsourceibias.n331 0.189894
R14009 commonsourceibias.n332 commonsourceibias.n317 0.189894
R14010 commonsourceibias.n336 commonsourceibias.n317 0.189894
R14011 commonsourceibias.n337 commonsourceibias.n336 0.189894
R14012 commonsourceibias.n337 commonsourceibias.n315 0.189894
R14013 commonsourceibias.n342 commonsourceibias.n315 0.189894
R14014 commonsourceibias.n343 commonsourceibias.n342 0.189894
R14015 commonsourceibias.n344 commonsourceibias.n343 0.189894
R14016 commonsourceibias.n344 commonsourceibias.n313 0.189894
R14017 commonsourceibias.n350 commonsourceibias.n313 0.189894
R14018 commonsourceibias.n351 commonsourceibias.n350 0.189894
R14019 commonsourceibias.n352 commonsourceibias.n351 0.189894
R14020 commonsourceibias.n352 commonsourceibias.n311 0.189894
R14021 commonsourceibias.n357 commonsourceibias.n311 0.189894
R14022 commonsourceibias.n358 commonsourceibias.n357 0.189894
R14023 commonsourceibias.n359 commonsourceibias.n358 0.189894
R14024 commonsourceibias.n359 commonsourceibias.n309 0.189894
R14025 commonsourceibias.n364 commonsourceibias.n309 0.189894
R14026 commonsourceibias.n365 commonsourceibias.n364 0.189894
R14027 commonsourceibias.n365 commonsourceibias.n307 0.189894
R14028 commonsourceibias.n285 commonsourceibias.n280 0.189894
R14029 commonsourceibias.n286 commonsourceibias.n285 0.189894
R14030 commonsourceibias.n286 commonsourceibias.n278 0.189894
R14031 commonsourceibias.n290 commonsourceibias.n278 0.189894
R14032 commonsourceibias.n291 commonsourceibias.n290 0.189894
R14033 commonsourceibias.n291 commonsourceibias.n276 0.189894
R14034 commonsourceibias.n295 commonsourceibias.n276 0.189894
R14035 commonsourceibias.n296 commonsourceibias.n295 0.189894
R14036 commonsourceibias.n296 commonsourceibias.n274 0.189894
R14037 commonsourceibias.n301 commonsourceibias.n274 0.189894
R14038 commonsourceibias.n378 commonsourceibias.n272 0.189894
R14039 commonsourceibias.n384 commonsourceibias.n272 0.189894
R14040 commonsourceibias.n385 commonsourceibias.n384 0.189894
R14041 commonsourceibias.n386 commonsourceibias.n385 0.189894
R14042 commonsourceibias.n386 commonsourceibias.n270 0.189894
R14043 commonsourceibias.n391 commonsourceibias.n270 0.189894
R14044 commonsourceibias.n392 commonsourceibias.n391 0.189894
R14045 commonsourceibias.n393 commonsourceibias.n392 0.189894
R14046 commonsourceibias.n393 commonsourceibias.n268 0.189894
R14047 commonsourceibias.n398 commonsourceibias.n268 0.189894
R14048 commonsourceibias.n399 commonsourceibias.n398 0.189894
R14049 commonsourceibias.n399 commonsourceibias.n266 0.189894
R14050 commonsourceibias.n487 commonsourceibias.n482 0.189894
R14051 commonsourceibias.n488 commonsourceibias.n487 0.189894
R14052 commonsourceibias.n488 commonsourceibias.n480 0.189894
R14053 commonsourceibias.n492 commonsourceibias.n480 0.189894
R14054 commonsourceibias.n493 commonsourceibias.n492 0.189894
R14055 commonsourceibias.n493 commonsourceibias.n478 0.189894
R14056 commonsourceibias.n497 commonsourceibias.n478 0.189894
R14057 commonsourceibias.n498 commonsourceibias.n497 0.189894
R14058 commonsourceibias.n498 commonsourceibias.n476 0.189894
R14059 commonsourceibias.n503 commonsourceibias.n476 0.189894
R14060 commonsourceibias.n504 commonsourceibias.n503 0.189894
R14061 commonsourceibias.n505 commonsourceibias.n504 0.189894
R14062 commonsourceibias.n505 commonsourceibias.n474 0.189894
R14063 commonsourceibias.n511 commonsourceibias.n474 0.189894
R14064 commonsourceibias.n512 commonsourceibias.n511 0.189894
R14065 commonsourceibias.n513 commonsourceibias.n512 0.189894
R14066 commonsourceibias.n513 commonsourceibias.n472 0.189894
R14067 commonsourceibias.n518 commonsourceibias.n472 0.189894
R14068 commonsourceibias.n519 commonsourceibias.n518 0.189894
R14069 commonsourceibias.n520 commonsourceibias.n519 0.189894
R14070 commonsourceibias.n520 commonsourceibias.n470 0.189894
R14071 commonsourceibias.n525 commonsourceibias.n470 0.189894
R14072 commonsourceibias.n526 commonsourceibias.n525 0.189894
R14073 commonsourceibias.n526 commonsourceibias.n468 0.189894
R14074 commonsourceibias.n423 commonsourceibias.n418 0.189894
R14075 commonsourceibias.n424 commonsourceibias.n423 0.189894
R14076 commonsourceibias.n424 commonsourceibias.n416 0.189894
R14077 commonsourceibias.n428 commonsourceibias.n416 0.189894
R14078 commonsourceibias.n429 commonsourceibias.n428 0.189894
R14079 commonsourceibias.n429 commonsourceibias.n414 0.189894
R14080 commonsourceibias.n433 commonsourceibias.n414 0.189894
R14081 commonsourceibias.n434 commonsourceibias.n433 0.189894
R14082 commonsourceibias.n434 commonsourceibias.n412 0.189894
R14083 commonsourceibias.n439 commonsourceibias.n412 0.189894
R14084 commonsourceibias.n440 commonsourceibias.n439 0.189894
R14085 commonsourceibias.n441 commonsourceibias.n440 0.189894
R14086 commonsourceibias.n441 commonsourceibias.n410 0.189894
R14087 commonsourceibias.n447 commonsourceibias.n410 0.189894
R14088 commonsourceibias.n448 commonsourceibias.n447 0.189894
R14089 commonsourceibias.n449 commonsourceibias.n448 0.189894
R14090 commonsourceibias.n449 commonsourceibias.n408 0.189894
R14091 commonsourceibias.n454 commonsourceibias.n408 0.189894
R14092 commonsourceibias.n455 commonsourceibias.n454 0.189894
R14093 commonsourceibias.n456 commonsourceibias.n455 0.189894
R14094 commonsourceibias.n456 commonsourceibias.n406 0.189894
R14095 commonsourceibias.n461 commonsourceibias.n406 0.189894
R14096 commonsourceibias.n462 commonsourceibias.n461 0.189894
R14097 commonsourceibias.n462 commonsourceibias.n404 0.189894
R14098 commonsourceibias.n112 commonsourceibias.n111 0.170955
R14099 commonsourceibias.n113 commonsourceibias.n112 0.170955
R14100 commonsourceibias.n377 commonsourceibias.n301 0.170955
R14101 commonsourceibias.n378 commonsourceibias.n377 0.170955
R14102 vdd.n303 vdd.n267 756.745
R14103 vdd.n252 vdd.n216 756.745
R14104 vdd.n209 vdd.n173 756.745
R14105 vdd.n158 vdd.n122 756.745
R14106 vdd.n116 vdd.n80 756.745
R14107 vdd.n65 vdd.n29 756.745
R14108 vdd.n1498 vdd.n1462 756.745
R14109 vdd.n1549 vdd.n1513 756.745
R14110 vdd.n1404 vdd.n1368 756.745
R14111 vdd.n1455 vdd.n1419 756.745
R14112 vdd.n1311 vdd.n1275 756.745
R14113 vdd.n1362 vdd.n1326 756.745
R14114 vdd.n1889 vdd.t97 640.208
R14115 vdd.n793 vdd.t82 640.208
R14116 vdd.n1863 vdd.t124 640.208
R14117 vdd.n785 vdd.t108 640.208
R14118 vdd.n2634 vdd.t69 640.208
R14119 vdd.n2354 vdd.t105 640.208
R14120 vdd.n661 vdd.t86 640.208
R14121 vdd.n2351 vdd.t90 640.208
R14122 vdd.n625 vdd.t94 640.208
R14123 vdd.n855 vdd.t101 640.208
R14124 vdd.n1110 vdd.t118 592.009
R14125 vdd.n1147 vdd.t65 592.009
R14126 vdd.n1021 vdd.t76 592.009
R14127 vdd.n2045 vdd.t61 592.009
R14128 vdd.n1682 vdd.t73 592.009
R14129 vdd.n1642 vdd.t79 592.009
R14130 vdd.n3021 vdd.t121 592.009
R14131 vdd.n427 vdd.t114 592.009
R14132 vdd.n387 vdd.t127 592.009
R14133 vdd.n580 vdd.t54 592.009
R14134 vdd.n543 vdd.t58 592.009
R14135 vdd.n2808 vdd.t111 592.009
R14136 vdd.n304 vdd.n303 585
R14137 vdd.n302 vdd.n269 585
R14138 vdd.n301 vdd.n300 585
R14139 vdd.n272 vdd.n270 585
R14140 vdd.n295 vdd.n294 585
R14141 vdd.n293 vdd.n292 585
R14142 vdd.n276 vdd.n275 585
R14143 vdd.n287 vdd.n286 585
R14144 vdd.n285 vdd.n284 585
R14145 vdd.n280 vdd.n279 585
R14146 vdd.n253 vdd.n252 585
R14147 vdd.n251 vdd.n218 585
R14148 vdd.n250 vdd.n249 585
R14149 vdd.n221 vdd.n219 585
R14150 vdd.n244 vdd.n243 585
R14151 vdd.n242 vdd.n241 585
R14152 vdd.n225 vdd.n224 585
R14153 vdd.n236 vdd.n235 585
R14154 vdd.n234 vdd.n233 585
R14155 vdd.n229 vdd.n228 585
R14156 vdd.n210 vdd.n209 585
R14157 vdd.n208 vdd.n175 585
R14158 vdd.n207 vdd.n206 585
R14159 vdd.n178 vdd.n176 585
R14160 vdd.n201 vdd.n200 585
R14161 vdd.n199 vdd.n198 585
R14162 vdd.n182 vdd.n181 585
R14163 vdd.n193 vdd.n192 585
R14164 vdd.n191 vdd.n190 585
R14165 vdd.n186 vdd.n185 585
R14166 vdd.n159 vdd.n158 585
R14167 vdd.n157 vdd.n124 585
R14168 vdd.n156 vdd.n155 585
R14169 vdd.n127 vdd.n125 585
R14170 vdd.n150 vdd.n149 585
R14171 vdd.n148 vdd.n147 585
R14172 vdd.n131 vdd.n130 585
R14173 vdd.n142 vdd.n141 585
R14174 vdd.n140 vdd.n139 585
R14175 vdd.n135 vdd.n134 585
R14176 vdd.n117 vdd.n116 585
R14177 vdd.n115 vdd.n82 585
R14178 vdd.n114 vdd.n113 585
R14179 vdd.n85 vdd.n83 585
R14180 vdd.n108 vdd.n107 585
R14181 vdd.n106 vdd.n105 585
R14182 vdd.n89 vdd.n88 585
R14183 vdd.n100 vdd.n99 585
R14184 vdd.n98 vdd.n97 585
R14185 vdd.n93 vdd.n92 585
R14186 vdd.n66 vdd.n65 585
R14187 vdd.n64 vdd.n31 585
R14188 vdd.n63 vdd.n62 585
R14189 vdd.n34 vdd.n32 585
R14190 vdd.n57 vdd.n56 585
R14191 vdd.n55 vdd.n54 585
R14192 vdd.n38 vdd.n37 585
R14193 vdd.n49 vdd.n48 585
R14194 vdd.n47 vdd.n46 585
R14195 vdd.n42 vdd.n41 585
R14196 vdd.n1499 vdd.n1498 585
R14197 vdd.n1497 vdd.n1464 585
R14198 vdd.n1496 vdd.n1495 585
R14199 vdd.n1467 vdd.n1465 585
R14200 vdd.n1490 vdd.n1489 585
R14201 vdd.n1488 vdd.n1487 585
R14202 vdd.n1471 vdd.n1470 585
R14203 vdd.n1482 vdd.n1481 585
R14204 vdd.n1480 vdd.n1479 585
R14205 vdd.n1475 vdd.n1474 585
R14206 vdd.n1550 vdd.n1549 585
R14207 vdd.n1548 vdd.n1515 585
R14208 vdd.n1547 vdd.n1546 585
R14209 vdd.n1518 vdd.n1516 585
R14210 vdd.n1541 vdd.n1540 585
R14211 vdd.n1539 vdd.n1538 585
R14212 vdd.n1522 vdd.n1521 585
R14213 vdd.n1533 vdd.n1532 585
R14214 vdd.n1531 vdd.n1530 585
R14215 vdd.n1526 vdd.n1525 585
R14216 vdd.n1405 vdd.n1404 585
R14217 vdd.n1403 vdd.n1370 585
R14218 vdd.n1402 vdd.n1401 585
R14219 vdd.n1373 vdd.n1371 585
R14220 vdd.n1396 vdd.n1395 585
R14221 vdd.n1394 vdd.n1393 585
R14222 vdd.n1377 vdd.n1376 585
R14223 vdd.n1388 vdd.n1387 585
R14224 vdd.n1386 vdd.n1385 585
R14225 vdd.n1381 vdd.n1380 585
R14226 vdd.n1456 vdd.n1455 585
R14227 vdd.n1454 vdd.n1421 585
R14228 vdd.n1453 vdd.n1452 585
R14229 vdd.n1424 vdd.n1422 585
R14230 vdd.n1447 vdd.n1446 585
R14231 vdd.n1445 vdd.n1444 585
R14232 vdd.n1428 vdd.n1427 585
R14233 vdd.n1439 vdd.n1438 585
R14234 vdd.n1437 vdd.n1436 585
R14235 vdd.n1432 vdd.n1431 585
R14236 vdd.n1312 vdd.n1311 585
R14237 vdd.n1310 vdd.n1277 585
R14238 vdd.n1309 vdd.n1308 585
R14239 vdd.n1280 vdd.n1278 585
R14240 vdd.n1303 vdd.n1302 585
R14241 vdd.n1301 vdd.n1300 585
R14242 vdd.n1284 vdd.n1283 585
R14243 vdd.n1295 vdd.n1294 585
R14244 vdd.n1293 vdd.n1292 585
R14245 vdd.n1288 vdd.n1287 585
R14246 vdd.n1363 vdd.n1362 585
R14247 vdd.n1361 vdd.n1328 585
R14248 vdd.n1360 vdd.n1359 585
R14249 vdd.n1331 vdd.n1329 585
R14250 vdd.n1354 vdd.n1353 585
R14251 vdd.n1352 vdd.n1351 585
R14252 vdd.n1335 vdd.n1334 585
R14253 vdd.n1346 vdd.n1345 585
R14254 vdd.n1344 vdd.n1343 585
R14255 vdd.n1339 vdd.n1338 585
R14256 vdd.n3137 vdd.n352 488.781
R14257 vdd.n3019 vdd.n350 488.781
R14258 vdd.n2941 vdd.n515 488.781
R14259 vdd.n2939 vdd.n517 488.781
R14260 vdd.n2040 vdd.n903 488.781
R14261 vdd.n2043 vdd.n2042 488.781
R14262 vdd.n1216 vdd.n981 488.781
R14263 vdd.n1214 vdd.n984 488.781
R14264 vdd.n281 vdd.t223 329.043
R14265 vdd.n230 vdd.t22 329.043
R14266 vdd.n187 vdd.t153 329.043
R14267 vdd.n136 vdd.t27 329.043
R14268 vdd.n94 vdd.t230 329.043
R14269 vdd.n43 vdd.t175 329.043
R14270 vdd.n1476 vdd.t43 329.043
R14271 vdd.n1527 vdd.t202 329.043
R14272 vdd.n1382 vdd.t195 329.043
R14273 vdd.n1433 vdd.t47 329.043
R14274 vdd.n1289 vdd.t176 329.043
R14275 vdd.n1340 vdd.t214 329.043
R14276 vdd.n1110 vdd.t120 319.788
R14277 vdd.n1147 vdd.t68 319.788
R14278 vdd.n1021 vdd.t78 319.788
R14279 vdd.n2045 vdd.t63 319.788
R14280 vdd.n1682 vdd.t74 319.788
R14281 vdd.n1642 vdd.t80 319.788
R14282 vdd.n3021 vdd.t122 319.788
R14283 vdd.n427 vdd.t116 319.788
R14284 vdd.n387 vdd.t128 319.788
R14285 vdd.n580 vdd.t57 319.788
R14286 vdd.n543 vdd.t60 319.788
R14287 vdd.n2808 vdd.t113 319.788
R14288 vdd.n1111 vdd.t119 303.69
R14289 vdd.n1148 vdd.t67 303.69
R14290 vdd.n1022 vdd.t77 303.69
R14291 vdd.n2046 vdd.t64 303.69
R14292 vdd.n1683 vdd.t75 303.69
R14293 vdd.n1643 vdd.t81 303.69
R14294 vdd.n3022 vdd.t123 303.69
R14295 vdd.n428 vdd.t117 303.69
R14296 vdd.n388 vdd.t129 303.69
R14297 vdd.n581 vdd.t56 303.69
R14298 vdd.n544 vdd.t59 303.69
R14299 vdd.n2809 vdd.t112 303.69
R14300 vdd.n2577 vdd.n741 297.074
R14301 vdd.n2770 vdd.n635 297.074
R14302 vdd.n2707 vdd.n632 297.074
R14303 vdd.n2500 vdd.n742 297.074
R14304 vdd.n2315 vdd.n782 297.074
R14305 vdd.n2246 vdd.n2245 297.074
R14306 vdd.n1992 vdd.n878 297.074
R14307 vdd.n2088 vdd.n876 297.074
R14308 vdd.n2686 vdd.n633 297.074
R14309 vdd.n2773 vdd.n2772 297.074
R14310 vdd.n2349 vdd.n743 297.074
R14311 vdd.n2575 vdd.n744 297.074
R14312 vdd.n2243 vdd.n791 297.074
R14313 vdd.n789 vdd.n764 297.074
R14314 vdd.n1929 vdd.n879 297.074
R14315 vdd.n2086 vdd.n880 297.074
R14316 vdd.n2688 vdd.n633 185
R14317 vdd.n2771 vdd.n633 185
R14318 vdd.n2690 vdd.n2689 185
R14319 vdd.n2689 vdd.n631 185
R14320 vdd.n2691 vdd.n667 185
R14321 vdd.n2701 vdd.n667 185
R14322 vdd.n2692 vdd.n676 185
R14323 vdd.n676 vdd.n674 185
R14324 vdd.n2694 vdd.n2693 185
R14325 vdd.n2695 vdd.n2694 185
R14326 vdd.n2647 vdd.n675 185
R14327 vdd.n675 vdd.n671 185
R14328 vdd.n2646 vdd.n2645 185
R14329 vdd.n2645 vdd.n2644 185
R14330 vdd.n678 vdd.n677 185
R14331 vdd.n679 vdd.n678 185
R14332 vdd.n2637 vdd.n2636 185
R14333 vdd.n2638 vdd.n2637 185
R14334 vdd.n2633 vdd.n688 185
R14335 vdd.n688 vdd.n685 185
R14336 vdd.n2632 vdd.n2631 185
R14337 vdd.n2631 vdd.n2630 185
R14338 vdd.n690 vdd.n689 185
R14339 vdd.n698 vdd.n690 185
R14340 vdd.n2623 vdd.n2622 185
R14341 vdd.n2624 vdd.n2623 185
R14342 vdd.n2621 vdd.n699 185
R14343 vdd.n2472 vdd.n699 185
R14344 vdd.n2620 vdd.n2619 185
R14345 vdd.n2619 vdd.n2618 185
R14346 vdd.n701 vdd.n700 185
R14347 vdd.n702 vdd.n701 185
R14348 vdd.n2611 vdd.n2610 185
R14349 vdd.n2612 vdd.n2611 185
R14350 vdd.n2609 vdd.n711 185
R14351 vdd.n711 vdd.n708 185
R14352 vdd.n2608 vdd.n2607 185
R14353 vdd.n2607 vdd.n2606 185
R14354 vdd.n713 vdd.n712 185
R14355 vdd.n721 vdd.n713 185
R14356 vdd.n2599 vdd.n2598 185
R14357 vdd.n2600 vdd.n2599 185
R14358 vdd.n2597 vdd.n722 185
R14359 vdd.n728 vdd.n722 185
R14360 vdd.n2596 vdd.n2595 185
R14361 vdd.n2595 vdd.n2594 185
R14362 vdd.n724 vdd.n723 185
R14363 vdd.n725 vdd.n724 185
R14364 vdd.n2587 vdd.n2586 185
R14365 vdd.n2588 vdd.n2587 185
R14366 vdd.n2585 vdd.n734 185
R14367 vdd.n2493 vdd.n734 185
R14368 vdd.n2584 vdd.n2583 185
R14369 vdd.n2583 vdd.n2582 185
R14370 vdd.n736 vdd.n735 185
R14371 vdd.t170 vdd.n736 185
R14372 vdd.n2575 vdd.n2574 185
R14373 vdd.n2576 vdd.n2575 185
R14374 vdd.n2573 vdd.n744 185
R14375 vdd.n2572 vdd.n2571 185
R14376 vdd.n746 vdd.n745 185
R14377 vdd.n2358 vdd.n2357 185
R14378 vdd.n2360 vdd.n2359 185
R14379 vdd.n2362 vdd.n2361 185
R14380 vdd.n2364 vdd.n2363 185
R14381 vdd.n2366 vdd.n2365 185
R14382 vdd.n2368 vdd.n2367 185
R14383 vdd.n2370 vdd.n2369 185
R14384 vdd.n2372 vdd.n2371 185
R14385 vdd.n2374 vdd.n2373 185
R14386 vdd.n2376 vdd.n2375 185
R14387 vdd.n2378 vdd.n2377 185
R14388 vdd.n2380 vdd.n2379 185
R14389 vdd.n2382 vdd.n2381 185
R14390 vdd.n2384 vdd.n2383 185
R14391 vdd.n2386 vdd.n2385 185
R14392 vdd.n2388 vdd.n2387 185
R14393 vdd.n2390 vdd.n2389 185
R14394 vdd.n2392 vdd.n2391 185
R14395 vdd.n2394 vdd.n2393 185
R14396 vdd.n2396 vdd.n2395 185
R14397 vdd.n2398 vdd.n2397 185
R14398 vdd.n2400 vdd.n2399 185
R14399 vdd.n2402 vdd.n2401 185
R14400 vdd.n2404 vdd.n2403 185
R14401 vdd.n2406 vdd.n2405 185
R14402 vdd.n2408 vdd.n2407 185
R14403 vdd.n2410 vdd.n2409 185
R14404 vdd.n2412 vdd.n2411 185
R14405 vdd.n2414 vdd.n2413 185
R14406 vdd.n2416 vdd.n2415 185
R14407 vdd.n2418 vdd.n2417 185
R14408 vdd.n2419 vdd.n2349 185
R14409 vdd.n2569 vdd.n2349 185
R14410 vdd.n2774 vdd.n2773 185
R14411 vdd.n2775 vdd.n624 185
R14412 vdd.n2777 vdd.n2776 185
R14413 vdd.n2779 vdd.n622 185
R14414 vdd.n2781 vdd.n2780 185
R14415 vdd.n2782 vdd.n621 185
R14416 vdd.n2784 vdd.n2783 185
R14417 vdd.n2786 vdd.n619 185
R14418 vdd.n2788 vdd.n2787 185
R14419 vdd.n2789 vdd.n618 185
R14420 vdd.n2791 vdd.n2790 185
R14421 vdd.n2793 vdd.n616 185
R14422 vdd.n2795 vdd.n2794 185
R14423 vdd.n2796 vdd.n615 185
R14424 vdd.n2798 vdd.n2797 185
R14425 vdd.n2800 vdd.n614 185
R14426 vdd.n2801 vdd.n611 185
R14427 vdd.n2804 vdd.n2803 185
R14428 vdd.n612 vdd.n610 185
R14429 vdd.n2660 vdd.n2659 185
R14430 vdd.n2662 vdd.n2661 185
R14431 vdd.n2664 vdd.n2656 185
R14432 vdd.n2666 vdd.n2665 185
R14433 vdd.n2667 vdd.n2655 185
R14434 vdd.n2669 vdd.n2668 185
R14435 vdd.n2671 vdd.n2653 185
R14436 vdd.n2673 vdd.n2672 185
R14437 vdd.n2674 vdd.n2652 185
R14438 vdd.n2676 vdd.n2675 185
R14439 vdd.n2678 vdd.n2650 185
R14440 vdd.n2680 vdd.n2679 185
R14441 vdd.n2681 vdd.n2649 185
R14442 vdd.n2683 vdd.n2682 185
R14443 vdd.n2685 vdd.n2648 185
R14444 vdd.n2687 vdd.n2686 185
R14445 vdd.n2686 vdd.n613 185
R14446 vdd.n2772 vdd.n628 185
R14447 vdd.n2772 vdd.n2771 185
R14448 vdd.n2424 vdd.n630 185
R14449 vdd.n631 vdd.n630 185
R14450 vdd.n2425 vdd.n666 185
R14451 vdd.n2701 vdd.n666 185
R14452 vdd.n2427 vdd.n2426 185
R14453 vdd.n2426 vdd.n674 185
R14454 vdd.n2428 vdd.n673 185
R14455 vdd.n2695 vdd.n673 185
R14456 vdd.n2430 vdd.n2429 185
R14457 vdd.n2429 vdd.n671 185
R14458 vdd.n2431 vdd.n681 185
R14459 vdd.n2644 vdd.n681 185
R14460 vdd.n2433 vdd.n2432 185
R14461 vdd.n2432 vdd.n679 185
R14462 vdd.n2434 vdd.n687 185
R14463 vdd.n2638 vdd.n687 185
R14464 vdd.n2436 vdd.n2435 185
R14465 vdd.n2435 vdd.n685 185
R14466 vdd.n2437 vdd.n692 185
R14467 vdd.n2630 vdd.n692 185
R14468 vdd.n2439 vdd.n2438 185
R14469 vdd.n2438 vdd.n698 185
R14470 vdd.n2440 vdd.n697 185
R14471 vdd.n2624 vdd.n697 185
R14472 vdd.n2474 vdd.n2473 185
R14473 vdd.n2473 vdd.n2472 185
R14474 vdd.n2475 vdd.n704 185
R14475 vdd.n2618 vdd.n704 185
R14476 vdd.n2477 vdd.n2476 185
R14477 vdd.n2476 vdd.n702 185
R14478 vdd.n2478 vdd.n710 185
R14479 vdd.n2612 vdd.n710 185
R14480 vdd.n2480 vdd.n2479 185
R14481 vdd.n2479 vdd.n708 185
R14482 vdd.n2481 vdd.n715 185
R14483 vdd.n2606 vdd.n715 185
R14484 vdd.n2483 vdd.n2482 185
R14485 vdd.n2482 vdd.n721 185
R14486 vdd.n2484 vdd.n720 185
R14487 vdd.n2600 vdd.n720 185
R14488 vdd.n2486 vdd.n2485 185
R14489 vdd.n2485 vdd.n728 185
R14490 vdd.n2487 vdd.n727 185
R14491 vdd.n2594 vdd.n727 185
R14492 vdd.n2489 vdd.n2488 185
R14493 vdd.n2488 vdd.n725 185
R14494 vdd.n2490 vdd.n733 185
R14495 vdd.n2588 vdd.n733 185
R14496 vdd.n2492 vdd.n2491 185
R14497 vdd.n2493 vdd.n2492 185
R14498 vdd.n2423 vdd.n738 185
R14499 vdd.n2582 vdd.n738 185
R14500 vdd.n2422 vdd.n2421 185
R14501 vdd.n2421 vdd.t170 185
R14502 vdd.n2420 vdd.n743 185
R14503 vdd.n2576 vdd.n743 185
R14504 vdd.n2040 vdd.n2039 185
R14505 vdd.n2041 vdd.n2040 185
R14506 vdd.n904 vdd.n902 185
R14507 vdd.n1606 vdd.n902 185
R14508 vdd.n1609 vdd.n1608 185
R14509 vdd.n1608 vdd.n1607 185
R14510 vdd.n907 vdd.n906 185
R14511 vdd.n908 vdd.n907 185
R14512 vdd.n1595 vdd.n1594 185
R14513 vdd.n1596 vdd.n1595 185
R14514 vdd.n916 vdd.n915 185
R14515 vdd.n1587 vdd.n915 185
R14516 vdd.n1590 vdd.n1589 185
R14517 vdd.n1589 vdd.n1588 185
R14518 vdd.n919 vdd.n918 185
R14519 vdd.n925 vdd.n919 185
R14520 vdd.n1578 vdd.n1577 185
R14521 vdd.n1579 vdd.n1578 185
R14522 vdd.n927 vdd.n926 185
R14523 vdd.n1570 vdd.n926 185
R14524 vdd.n1573 vdd.n1572 185
R14525 vdd.n1572 vdd.n1571 185
R14526 vdd.n930 vdd.n929 185
R14527 vdd.n931 vdd.n930 185
R14528 vdd.n1561 vdd.n1560 185
R14529 vdd.n1562 vdd.n1561 185
R14530 vdd.n939 vdd.n938 185
R14531 vdd.n938 vdd.n937 185
R14532 vdd.n1274 vdd.n1273 185
R14533 vdd.n1273 vdd.n1272 185
R14534 vdd.n942 vdd.n941 185
R14535 vdd.n948 vdd.n942 185
R14536 vdd.n1263 vdd.n1262 185
R14537 vdd.n1264 vdd.n1263 185
R14538 vdd.n950 vdd.n949 185
R14539 vdd.n1255 vdd.n949 185
R14540 vdd.n1258 vdd.n1257 185
R14541 vdd.n1257 vdd.n1256 185
R14542 vdd.n953 vdd.n952 185
R14543 vdd.n960 vdd.n953 185
R14544 vdd.n1246 vdd.n1245 185
R14545 vdd.n1247 vdd.n1246 185
R14546 vdd.n962 vdd.n961 185
R14547 vdd.n961 vdd.n959 185
R14548 vdd.n1241 vdd.n1240 185
R14549 vdd.n1240 vdd.n1239 185
R14550 vdd.n965 vdd.n964 185
R14551 vdd.n966 vdd.n965 185
R14552 vdd.n1230 vdd.n1229 185
R14553 vdd.n1231 vdd.n1230 185
R14554 vdd.n974 vdd.n973 185
R14555 vdd.n973 vdd.n972 185
R14556 vdd.n1225 vdd.n1224 185
R14557 vdd.n1224 vdd.n1223 185
R14558 vdd.n977 vdd.n976 185
R14559 vdd.n983 vdd.n977 185
R14560 vdd.n1214 vdd.n1213 185
R14561 vdd.n1215 vdd.n1214 185
R14562 vdd.n1210 vdd.n984 185
R14563 vdd.n1209 vdd.n987 185
R14564 vdd.n1208 vdd.n988 185
R14565 vdd.n988 vdd.n982 185
R14566 vdd.n991 vdd.n989 185
R14567 vdd.n1204 vdd.n993 185
R14568 vdd.n1203 vdd.n994 185
R14569 vdd.n1202 vdd.n996 185
R14570 vdd.n999 vdd.n997 185
R14571 vdd.n1198 vdd.n1001 185
R14572 vdd.n1197 vdd.n1002 185
R14573 vdd.n1196 vdd.n1004 185
R14574 vdd.n1007 vdd.n1005 185
R14575 vdd.n1192 vdd.n1009 185
R14576 vdd.n1191 vdd.n1010 185
R14577 vdd.n1190 vdd.n1012 185
R14578 vdd.n1015 vdd.n1013 185
R14579 vdd.n1186 vdd.n1017 185
R14580 vdd.n1185 vdd.n1018 185
R14581 vdd.n1184 vdd.n1020 185
R14582 vdd.n1025 vdd.n1023 185
R14583 vdd.n1180 vdd.n1027 185
R14584 vdd.n1179 vdd.n1028 185
R14585 vdd.n1178 vdd.n1030 185
R14586 vdd.n1033 vdd.n1031 185
R14587 vdd.n1174 vdd.n1035 185
R14588 vdd.n1173 vdd.n1036 185
R14589 vdd.n1172 vdd.n1038 185
R14590 vdd.n1041 vdd.n1039 185
R14591 vdd.n1168 vdd.n1043 185
R14592 vdd.n1167 vdd.n1044 185
R14593 vdd.n1166 vdd.n1046 185
R14594 vdd.n1049 vdd.n1047 185
R14595 vdd.n1162 vdd.n1051 185
R14596 vdd.n1161 vdd.n1052 185
R14597 vdd.n1160 vdd.n1054 185
R14598 vdd.n1057 vdd.n1055 185
R14599 vdd.n1156 vdd.n1059 185
R14600 vdd.n1155 vdd.n1060 185
R14601 vdd.n1154 vdd.n1062 185
R14602 vdd.n1065 vdd.n1063 185
R14603 vdd.n1150 vdd.n1067 185
R14604 vdd.n1149 vdd.n1146 185
R14605 vdd.n1144 vdd.n1068 185
R14606 vdd.n1143 vdd.n1142 185
R14607 vdd.n1073 vdd.n1070 185
R14608 vdd.n1138 vdd.n1074 185
R14609 vdd.n1137 vdd.n1076 185
R14610 vdd.n1136 vdd.n1077 185
R14611 vdd.n1081 vdd.n1078 185
R14612 vdd.n1132 vdd.n1082 185
R14613 vdd.n1131 vdd.n1084 185
R14614 vdd.n1130 vdd.n1085 185
R14615 vdd.n1089 vdd.n1086 185
R14616 vdd.n1126 vdd.n1090 185
R14617 vdd.n1125 vdd.n1092 185
R14618 vdd.n1124 vdd.n1093 185
R14619 vdd.n1097 vdd.n1094 185
R14620 vdd.n1120 vdd.n1098 185
R14621 vdd.n1119 vdd.n1100 185
R14622 vdd.n1118 vdd.n1101 185
R14623 vdd.n1105 vdd.n1102 185
R14624 vdd.n1114 vdd.n1106 185
R14625 vdd.n1113 vdd.n1108 185
R14626 vdd.n1109 vdd.n981 185
R14627 vdd.n982 vdd.n981 185
R14628 vdd.n2044 vdd.n2043 185
R14629 vdd.n2048 vdd.n897 185
R14630 vdd.n1711 vdd.n896 185
R14631 vdd.n1714 vdd.n1713 185
R14632 vdd.n1716 vdd.n1715 185
R14633 vdd.n1719 vdd.n1718 185
R14634 vdd.n1721 vdd.n1720 185
R14635 vdd.n1723 vdd.n1709 185
R14636 vdd.n1725 vdd.n1724 185
R14637 vdd.n1726 vdd.n1703 185
R14638 vdd.n1728 vdd.n1727 185
R14639 vdd.n1730 vdd.n1701 185
R14640 vdd.n1732 vdd.n1731 185
R14641 vdd.n1733 vdd.n1696 185
R14642 vdd.n1735 vdd.n1734 185
R14643 vdd.n1737 vdd.n1694 185
R14644 vdd.n1739 vdd.n1738 185
R14645 vdd.n1740 vdd.n1690 185
R14646 vdd.n1742 vdd.n1741 185
R14647 vdd.n1744 vdd.n1687 185
R14648 vdd.n1746 vdd.n1745 185
R14649 vdd.n1688 vdd.n1681 185
R14650 vdd.n1750 vdd.n1685 185
R14651 vdd.n1751 vdd.n1677 185
R14652 vdd.n1753 vdd.n1752 185
R14653 vdd.n1755 vdd.n1675 185
R14654 vdd.n1757 vdd.n1756 185
R14655 vdd.n1758 vdd.n1670 185
R14656 vdd.n1760 vdd.n1759 185
R14657 vdd.n1762 vdd.n1668 185
R14658 vdd.n1764 vdd.n1763 185
R14659 vdd.n1765 vdd.n1663 185
R14660 vdd.n1767 vdd.n1766 185
R14661 vdd.n1769 vdd.n1661 185
R14662 vdd.n1771 vdd.n1770 185
R14663 vdd.n1772 vdd.n1656 185
R14664 vdd.n1774 vdd.n1773 185
R14665 vdd.n1776 vdd.n1654 185
R14666 vdd.n1778 vdd.n1777 185
R14667 vdd.n1779 vdd.n1650 185
R14668 vdd.n1781 vdd.n1780 185
R14669 vdd.n1783 vdd.n1647 185
R14670 vdd.n1785 vdd.n1784 185
R14671 vdd.n1648 vdd.n1641 185
R14672 vdd.n1789 vdd.n1645 185
R14673 vdd.n1790 vdd.n1637 185
R14674 vdd.n1792 vdd.n1791 185
R14675 vdd.n1794 vdd.n1635 185
R14676 vdd.n1796 vdd.n1795 185
R14677 vdd.n1797 vdd.n1630 185
R14678 vdd.n1799 vdd.n1798 185
R14679 vdd.n1801 vdd.n1628 185
R14680 vdd.n1803 vdd.n1802 185
R14681 vdd.n1804 vdd.n1623 185
R14682 vdd.n1806 vdd.n1805 185
R14683 vdd.n1808 vdd.n1622 185
R14684 vdd.n1809 vdd.n1619 185
R14685 vdd.n1812 vdd.n1811 185
R14686 vdd.n1621 vdd.n1617 185
R14687 vdd.n2029 vdd.n1615 185
R14688 vdd.n2031 vdd.n2030 185
R14689 vdd.n2033 vdd.n1613 185
R14690 vdd.n2035 vdd.n2034 185
R14691 vdd.n2036 vdd.n903 185
R14692 vdd.n2042 vdd.n900 185
R14693 vdd.n2042 vdd.n2041 185
R14694 vdd.n911 vdd.n899 185
R14695 vdd.n1606 vdd.n899 185
R14696 vdd.n1605 vdd.n1604 185
R14697 vdd.n1607 vdd.n1605 185
R14698 vdd.n910 vdd.n909 185
R14699 vdd.n909 vdd.n908 185
R14700 vdd.n1598 vdd.n1597 185
R14701 vdd.n1597 vdd.n1596 185
R14702 vdd.n914 vdd.n913 185
R14703 vdd.n1587 vdd.n914 185
R14704 vdd.n1586 vdd.n1585 185
R14705 vdd.n1588 vdd.n1586 185
R14706 vdd.n921 vdd.n920 185
R14707 vdd.n925 vdd.n920 185
R14708 vdd.n1581 vdd.n1580 185
R14709 vdd.n1580 vdd.n1579 185
R14710 vdd.n924 vdd.n923 185
R14711 vdd.n1570 vdd.n924 185
R14712 vdd.n1569 vdd.n1568 185
R14713 vdd.n1571 vdd.n1569 185
R14714 vdd.n933 vdd.n932 185
R14715 vdd.n932 vdd.n931 185
R14716 vdd.n1564 vdd.n1563 185
R14717 vdd.n1563 vdd.n1562 185
R14718 vdd.n936 vdd.n935 185
R14719 vdd.n937 vdd.n936 185
R14720 vdd.n1271 vdd.n1270 185
R14721 vdd.n1272 vdd.n1271 185
R14722 vdd.n944 vdd.n943 185
R14723 vdd.n948 vdd.n943 185
R14724 vdd.n1266 vdd.n1265 185
R14725 vdd.n1265 vdd.n1264 185
R14726 vdd.n947 vdd.n946 185
R14727 vdd.n1255 vdd.n947 185
R14728 vdd.n1254 vdd.n1253 185
R14729 vdd.n1256 vdd.n1254 185
R14730 vdd.n955 vdd.n954 185
R14731 vdd.n960 vdd.n954 185
R14732 vdd.n1249 vdd.n1248 185
R14733 vdd.n1248 vdd.n1247 185
R14734 vdd.n958 vdd.n957 185
R14735 vdd.n959 vdd.n958 185
R14736 vdd.n1238 vdd.n1237 185
R14737 vdd.n1239 vdd.n1238 185
R14738 vdd.n968 vdd.n967 185
R14739 vdd.n967 vdd.n966 185
R14740 vdd.n1233 vdd.n1232 185
R14741 vdd.n1232 vdd.n1231 185
R14742 vdd.n971 vdd.n970 185
R14743 vdd.n972 vdd.n971 185
R14744 vdd.n1222 vdd.n1221 185
R14745 vdd.n1223 vdd.n1222 185
R14746 vdd.n979 vdd.n978 185
R14747 vdd.n983 vdd.n978 185
R14748 vdd.n1217 vdd.n1216 185
R14749 vdd.n1216 vdd.n1215 185
R14750 vdd.n784 vdd.n782 185
R14751 vdd.n2244 vdd.n782 185
R14752 vdd.n2166 vdd.n801 185
R14753 vdd.n801 vdd.t144 185
R14754 vdd.n2168 vdd.n2167 185
R14755 vdd.n2169 vdd.n2168 185
R14756 vdd.n2165 vdd.n800 185
R14757 vdd.n1868 vdd.n800 185
R14758 vdd.n2164 vdd.n2163 185
R14759 vdd.n2163 vdd.n2162 185
R14760 vdd.n803 vdd.n802 185
R14761 vdd.n804 vdd.n803 185
R14762 vdd.n2153 vdd.n2152 185
R14763 vdd.n2154 vdd.n2153 185
R14764 vdd.n2151 vdd.n814 185
R14765 vdd.n814 vdd.n811 185
R14766 vdd.n2150 vdd.n2149 185
R14767 vdd.n2149 vdd.n2148 185
R14768 vdd.n816 vdd.n815 185
R14769 vdd.n817 vdd.n816 185
R14770 vdd.n2141 vdd.n2140 185
R14771 vdd.n2142 vdd.n2141 185
R14772 vdd.n2139 vdd.n825 185
R14773 vdd.n830 vdd.n825 185
R14774 vdd.n2138 vdd.n2137 185
R14775 vdd.n2137 vdd.n2136 185
R14776 vdd.n827 vdd.n826 185
R14777 vdd.n836 vdd.n827 185
R14778 vdd.n2129 vdd.n2128 185
R14779 vdd.n2130 vdd.n2129 185
R14780 vdd.n2127 vdd.n837 185
R14781 vdd.n1969 vdd.n837 185
R14782 vdd.n2126 vdd.n2125 185
R14783 vdd.n2125 vdd.n2124 185
R14784 vdd.n839 vdd.n838 185
R14785 vdd.n840 vdd.n839 185
R14786 vdd.n2117 vdd.n2116 185
R14787 vdd.n2118 vdd.n2117 185
R14788 vdd.n2115 vdd.n849 185
R14789 vdd.n849 vdd.n846 185
R14790 vdd.n2114 vdd.n2113 185
R14791 vdd.n2113 vdd.n2112 185
R14792 vdd.n851 vdd.n850 185
R14793 vdd.n861 vdd.n851 185
R14794 vdd.n2104 vdd.n2103 185
R14795 vdd.n2105 vdd.n2104 185
R14796 vdd.n2102 vdd.n862 185
R14797 vdd.n862 vdd.n858 185
R14798 vdd.n2101 vdd.n2100 185
R14799 vdd.n2100 vdd.n2099 185
R14800 vdd.n864 vdd.n863 185
R14801 vdd.n865 vdd.n864 185
R14802 vdd.n2092 vdd.n2091 185
R14803 vdd.n2093 vdd.n2092 185
R14804 vdd.n2090 vdd.n874 185
R14805 vdd.n874 vdd.n871 185
R14806 vdd.n2089 vdd.n2088 185
R14807 vdd.n2088 vdd.n2087 185
R14808 vdd.n876 vdd.n875 185
R14809 vdd.n1824 vdd.n1823 185
R14810 vdd.n1825 vdd.n1821 185
R14811 vdd.n1821 vdd.n877 185
R14812 vdd.n1827 vdd.n1826 185
R14813 vdd.n1829 vdd.n1820 185
R14814 vdd.n1832 vdd.n1831 185
R14815 vdd.n1833 vdd.n1819 185
R14816 vdd.n1835 vdd.n1834 185
R14817 vdd.n1837 vdd.n1818 185
R14818 vdd.n1840 vdd.n1839 185
R14819 vdd.n1841 vdd.n1817 185
R14820 vdd.n1843 vdd.n1842 185
R14821 vdd.n1845 vdd.n1816 185
R14822 vdd.n1848 vdd.n1847 185
R14823 vdd.n1849 vdd.n1815 185
R14824 vdd.n1851 vdd.n1850 185
R14825 vdd.n1853 vdd.n1814 185
R14826 vdd.n2026 vdd.n1854 185
R14827 vdd.n2025 vdd.n2024 185
R14828 vdd.n2022 vdd.n1855 185
R14829 vdd.n2020 vdd.n2019 185
R14830 vdd.n2018 vdd.n1856 185
R14831 vdd.n2017 vdd.n2016 185
R14832 vdd.n2014 vdd.n1857 185
R14833 vdd.n2012 vdd.n2011 185
R14834 vdd.n2010 vdd.n1858 185
R14835 vdd.n2009 vdd.n2008 185
R14836 vdd.n2006 vdd.n1859 185
R14837 vdd.n2004 vdd.n2003 185
R14838 vdd.n2002 vdd.n1860 185
R14839 vdd.n2001 vdd.n2000 185
R14840 vdd.n1998 vdd.n1861 185
R14841 vdd.n1996 vdd.n1995 185
R14842 vdd.n1994 vdd.n1862 185
R14843 vdd.n1993 vdd.n1992 185
R14844 vdd.n2247 vdd.n2246 185
R14845 vdd.n2249 vdd.n2248 185
R14846 vdd.n2251 vdd.n2250 185
R14847 vdd.n2254 vdd.n2253 185
R14848 vdd.n2256 vdd.n2255 185
R14849 vdd.n2258 vdd.n2257 185
R14850 vdd.n2260 vdd.n2259 185
R14851 vdd.n2262 vdd.n2261 185
R14852 vdd.n2264 vdd.n2263 185
R14853 vdd.n2266 vdd.n2265 185
R14854 vdd.n2268 vdd.n2267 185
R14855 vdd.n2270 vdd.n2269 185
R14856 vdd.n2272 vdd.n2271 185
R14857 vdd.n2274 vdd.n2273 185
R14858 vdd.n2276 vdd.n2275 185
R14859 vdd.n2278 vdd.n2277 185
R14860 vdd.n2280 vdd.n2279 185
R14861 vdd.n2282 vdd.n2281 185
R14862 vdd.n2284 vdd.n2283 185
R14863 vdd.n2286 vdd.n2285 185
R14864 vdd.n2288 vdd.n2287 185
R14865 vdd.n2290 vdd.n2289 185
R14866 vdd.n2292 vdd.n2291 185
R14867 vdd.n2294 vdd.n2293 185
R14868 vdd.n2296 vdd.n2295 185
R14869 vdd.n2298 vdd.n2297 185
R14870 vdd.n2300 vdd.n2299 185
R14871 vdd.n2302 vdd.n2301 185
R14872 vdd.n2304 vdd.n2303 185
R14873 vdd.n2306 vdd.n2305 185
R14874 vdd.n2308 vdd.n2307 185
R14875 vdd.n2310 vdd.n2309 185
R14876 vdd.n2312 vdd.n2311 185
R14877 vdd.n2313 vdd.n783 185
R14878 vdd.n2315 vdd.n2314 185
R14879 vdd.n2316 vdd.n2315 185
R14880 vdd.n2245 vdd.n787 185
R14881 vdd.n2245 vdd.n2244 185
R14882 vdd.n1866 vdd.n788 185
R14883 vdd.t144 vdd.n788 185
R14884 vdd.n1867 vdd.n798 185
R14885 vdd.n2169 vdd.n798 185
R14886 vdd.n1870 vdd.n1869 185
R14887 vdd.n1869 vdd.n1868 185
R14888 vdd.n1871 vdd.n805 185
R14889 vdd.n2162 vdd.n805 185
R14890 vdd.n1873 vdd.n1872 185
R14891 vdd.n1872 vdd.n804 185
R14892 vdd.n1874 vdd.n812 185
R14893 vdd.n2154 vdd.n812 185
R14894 vdd.n1876 vdd.n1875 185
R14895 vdd.n1875 vdd.n811 185
R14896 vdd.n1877 vdd.n818 185
R14897 vdd.n2148 vdd.n818 185
R14898 vdd.n1879 vdd.n1878 185
R14899 vdd.n1878 vdd.n817 185
R14900 vdd.n1880 vdd.n823 185
R14901 vdd.n2142 vdd.n823 185
R14902 vdd.n1882 vdd.n1881 185
R14903 vdd.n1881 vdd.n830 185
R14904 vdd.n1883 vdd.n828 185
R14905 vdd.n2136 vdd.n828 185
R14906 vdd.n1885 vdd.n1884 185
R14907 vdd.n1884 vdd.n836 185
R14908 vdd.n1886 vdd.n834 185
R14909 vdd.n2130 vdd.n834 185
R14910 vdd.n1971 vdd.n1970 185
R14911 vdd.n1970 vdd.n1969 185
R14912 vdd.n1972 vdd.n841 185
R14913 vdd.n2124 vdd.n841 185
R14914 vdd.n1974 vdd.n1973 185
R14915 vdd.n1973 vdd.n840 185
R14916 vdd.n1975 vdd.n847 185
R14917 vdd.n2118 vdd.n847 185
R14918 vdd.n1977 vdd.n1976 185
R14919 vdd.n1976 vdd.n846 185
R14920 vdd.n1978 vdd.n852 185
R14921 vdd.n2112 vdd.n852 185
R14922 vdd.n1980 vdd.n1979 185
R14923 vdd.n1979 vdd.n861 185
R14924 vdd.n1981 vdd.n859 185
R14925 vdd.n2105 vdd.n859 185
R14926 vdd.n1983 vdd.n1982 185
R14927 vdd.n1982 vdd.n858 185
R14928 vdd.n1984 vdd.n866 185
R14929 vdd.n2099 vdd.n866 185
R14930 vdd.n1986 vdd.n1985 185
R14931 vdd.n1985 vdd.n865 185
R14932 vdd.n1987 vdd.n872 185
R14933 vdd.n2093 vdd.n872 185
R14934 vdd.n1989 vdd.n1988 185
R14935 vdd.n1988 vdd.n871 185
R14936 vdd.n1990 vdd.n878 185
R14937 vdd.n2087 vdd.n878 185
R14938 vdd.n3137 vdd.n3136 185
R14939 vdd.n3138 vdd.n3137 185
R14940 vdd.n347 vdd.n346 185
R14941 vdd.n3139 vdd.n347 185
R14942 vdd.n3142 vdd.n3141 185
R14943 vdd.n3141 vdd.n3140 185
R14944 vdd.n3143 vdd.n341 185
R14945 vdd.n341 vdd.n340 185
R14946 vdd.n3145 vdd.n3144 185
R14947 vdd.n3146 vdd.n3145 185
R14948 vdd.n336 vdd.n335 185
R14949 vdd.n3147 vdd.n336 185
R14950 vdd.n3150 vdd.n3149 185
R14951 vdd.n3149 vdd.n3148 185
R14952 vdd.n3151 vdd.n330 185
R14953 vdd.n330 vdd.n329 185
R14954 vdd.n3153 vdd.n3152 185
R14955 vdd.n3154 vdd.n3153 185
R14956 vdd.n324 vdd.n323 185
R14957 vdd.n3155 vdd.n324 185
R14958 vdd.n3158 vdd.n3157 185
R14959 vdd.n3157 vdd.n3156 185
R14960 vdd.n3159 vdd.n319 185
R14961 vdd.n325 vdd.n319 185
R14962 vdd.n3161 vdd.n3160 185
R14963 vdd.n3162 vdd.n3161 185
R14964 vdd.n315 vdd.n313 185
R14965 vdd.n3163 vdd.n315 185
R14966 vdd.n3166 vdd.n3165 185
R14967 vdd.n3165 vdd.n3164 185
R14968 vdd.n314 vdd.n312 185
R14969 vdd.n481 vdd.n314 185
R14970 vdd.n2988 vdd.n2987 185
R14971 vdd.n2989 vdd.n2988 185
R14972 vdd.n483 vdd.n482 185
R14973 vdd.n2980 vdd.n482 185
R14974 vdd.n2983 vdd.n2982 185
R14975 vdd.n2982 vdd.n2981 185
R14976 vdd.n486 vdd.n485 185
R14977 vdd.n493 vdd.n486 185
R14978 vdd.n2971 vdd.n2970 185
R14979 vdd.n2972 vdd.n2971 185
R14980 vdd.n495 vdd.n494 185
R14981 vdd.n494 vdd.n492 185
R14982 vdd.n2966 vdd.n2965 185
R14983 vdd.n2965 vdd.n2964 185
R14984 vdd.n498 vdd.n497 185
R14985 vdd.n499 vdd.n498 185
R14986 vdd.n2955 vdd.n2954 185
R14987 vdd.n2956 vdd.n2955 185
R14988 vdd.n507 vdd.n506 185
R14989 vdd.n506 vdd.n505 185
R14990 vdd.n2950 vdd.n2949 185
R14991 vdd.n2949 vdd.n2948 185
R14992 vdd.n510 vdd.n509 185
R14993 vdd.n511 vdd.n510 185
R14994 vdd.n2939 vdd.n2938 185
R14995 vdd.n2940 vdd.n2939 185
R14996 vdd.n2935 vdd.n517 185
R14997 vdd.n2934 vdd.n2933 185
R14998 vdd.n2931 vdd.n519 185
R14999 vdd.n2931 vdd.n516 185
R15000 vdd.n2930 vdd.n2929 185
R15001 vdd.n2928 vdd.n2927 185
R15002 vdd.n2926 vdd.n2925 185
R15003 vdd.n2924 vdd.n2923 185
R15004 vdd.n2922 vdd.n525 185
R15005 vdd.n2920 vdd.n2919 185
R15006 vdd.n2918 vdd.n526 185
R15007 vdd.n2917 vdd.n2916 185
R15008 vdd.n2914 vdd.n531 185
R15009 vdd.n2912 vdd.n2911 185
R15010 vdd.n2910 vdd.n532 185
R15011 vdd.n2909 vdd.n2908 185
R15012 vdd.n2906 vdd.n537 185
R15013 vdd.n2904 vdd.n2903 185
R15014 vdd.n2902 vdd.n538 185
R15015 vdd.n2901 vdd.n2900 185
R15016 vdd.n2898 vdd.n545 185
R15017 vdd.n2896 vdd.n2895 185
R15018 vdd.n2894 vdd.n546 185
R15019 vdd.n2893 vdd.n2892 185
R15020 vdd.n2890 vdd.n551 185
R15021 vdd.n2888 vdd.n2887 185
R15022 vdd.n2886 vdd.n552 185
R15023 vdd.n2885 vdd.n2884 185
R15024 vdd.n2882 vdd.n557 185
R15025 vdd.n2880 vdd.n2879 185
R15026 vdd.n2878 vdd.n558 185
R15027 vdd.n2877 vdd.n2876 185
R15028 vdd.n2874 vdd.n563 185
R15029 vdd.n2872 vdd.n2871 185
R15030 vdd.n2870 vdd.n564 185
R15031 vdd.n2869 vdd.n2868 185
R15032 vdd.n2866 vdd.n569 185
R15033 vdd.n2864 vdd.n2863 185
R15034 vdd.n2862 vdd.n570 185
R15035 vdd.n2861 vdd.n2860 185
R15036 vdd.n2858 vdd.n575 185
R15037 vdd.n2856 vdd.n2855 185
R15038 vdd.n2854 vdd.n576 185
R15039 vdd.n585 vdd.n579 185
R15040 vdd.n2850 vdd.n2849 185
R15041 vdd.n2847 vdd.n583 185
R15042 vdd.n2846 vdd.n2845 185
R15043 vdd.n2844 vdd.n2843 185
R15044 vdd.n2842 vdd.n589 185
R15045 vdd.n2840 vdd.n2839 185
R15046 vdd.n2838 vdd.n590 185
R15047 vdd.n2837 vdd.n2836 185
R15048 vdd.n2834 vdd.n595 185
R15049 vdd.n2832 vdd.n2831 185
R15050 vdd.n2830 vdd.n596 185
R15051 vdd.n2829 vdd.n2828 185
R15052 vdd.n2826 vdd.n601 185
R15053 vdd.n2824 vdd.n2823 185
R15054 vdd.n2822 vdd.n602 185
R15055 vdd.n2821 vdd.n2820 185
R15056 vdd.n2818 vdd.n2817 185
R15057 vdd.n2816 vdd.n2815 185
R15058 vdd.n2814 vdd.n2813 185
R15059 vdd.n2812 vdd.n2811 185
R15060 vdd.n2807 vdd.n515 185
R15061 vdd.n516 vdd.n515 185
R15062 vdd.n3020 vdd.n3019 185
R15063 vdd.n3024 vdd.n462 185
R15064 vdd.n3026 vdd.n3025 185
R15065 vdd.n3028 vdd.n460 185
R15066 vdd.n3030 vdd.n3029 185
R15067 vdd.n3031 vdd.n455 185
R15068 vdd.n3033 vdd.n3032 185
R15069 vdd.n3035 vdd.n453 185
R15070 vdd.n3037 vdd.n3036 185
R15071 vdd.n3038 vdd.n448 185
R15072 vdd.n3040 vdd.n3039 185
R15073 vdd.n3042 vdd.n446 185
R15074 vdd.n3044 vdd.n3043 185
R15075 vdd.n3045 vdd.n441 185
R15076 vdd.n3047 vdd.n3046 185
R15077 vdd.n3049 vdd.n439 185
R15078 vdd.n3051 vdd.n3050 185
R15079 vdd.n3052 vdd.n435 185
R15080 vdd.n3054 vdd.n3053 185
R15081 vdd.n3056 vdd.n432 185
R15082 vdd.n3058 vdd.n3057 185
R15083 vdd.n433 vdd.n426 185
R15084 vdd.n3062 vdd.n430 185
R15085 vdd.n3063 vdd.n422 185
R15086 vdd.n3065 vdd.n3064 185
R15087 vdd.n3067 vdd.n420 185
R15088 vdd.n3069 vdd.n3068 185
R15089 vdd.n3070 vdd.n415 185
R15090 vdd.n3072 vdd.n3071 185
R15091 vdd.n3074 vdd.n413 185
R15092 vdd.n3076 vdd.n3075 185
R15093 vdd.n3077 vdd.n408 185
R15094 vdd.n3079 vdd.n3078 185
R15095 vdd.n3081 vdd.n406 185
R15096 vdd.n3083 vdd.n3082 185
R15097 vdd.n3084 vdd.n401 185
R15098 vdd.n3086 vdd.n3085 185
R15099 vdd.n3088 vdd.n399 185
R15100 vdd.n3090 vdd.n3089 185
R15101 vdd.n3091 vdd.n395 185
R15102 vdd.n3093 vdd.n3092 185
R15103 vdd.n3095 vdd.n392 185
R15104 vdd.n3097 vdd.n3096 185
R15105 vdd.n393 vdd.n386 185
R15106 vdd.n3101 vdd.n390 185
R15107 vdd.n3102 vdd.n382 185
R15108 vdd.n3104 vdd.n3103 185
R15109 vdd.n3106 vdd.n380 185
R15110 vdd.n3108 vdd.n3107 185
R15111 vdd.n3109 vdd.n375 185
R15112 vdd.n3111 vdd.n3110 185
R15113 vdd.n3113 vdd.n373 185
R15114 vdd.n3115 vdd.n3114 185
R15115 vdd.n3116 vdd.n368 185
R15116 vdd.n3118 vdd.n3117 185
R15117 vdd.n3120 vdd.n366 185
R15118 vdd.n3122 vdd.n3121 185
R15119 vdd.n3123 vdd.n360 185
R15120 vdd.n3125 vdd.n3124 185
R15121 vdd.n3127 vdd.n359 185
R15122 vdd.n3128 vdd.n358 185
R15123 vdd.n3131 vdd.n3130 185
R15124 vdd.n3132 vdd.n356 185
R15125 vdd.n3133 vdd.n352 185
R15126 vdd.n3015 vdd.n350 185
R15127 vdd.n3138 vdd.n350 185
R15128 vdd.n3014 vdd.n349 185
R15129 vdd.n3139 vdd.n349 185
R15130 vdd.n3013 vdd.n348 185
R15131 vdd.n3140 vdd.n348 185
R15132 vdd.n468 vdd.n467 185
R15133 vdd.n467 vdd.n340 185
R15134 vdd.n3009 vdd.n339 185
R15135 vdd.n3146 vdd.n339 185
R15136 vdd.n3008 vdd.n338 185
R15137 vdd.n3147 vdd.n338 185
R15138 vdd.n3007 vdd.n337 185
R15139 vdd.n3148 vdd.n337 185
R15140 vdd.n471 vdd.n470 185
R15141 vdd.n470 vdd.n329 185
R15142 vdd.n3003 vdd.n328 185
R15143 vdd.n3154 vdd.n328 185
R15144 vdd.n3002 vdd.n327 185
R15145 vdd.n3155 vdd.n327 185
R15146 vdd.n3001 vdd.n326 185
R15147 vdd.n3156 vdd.n326 185
R15148 vdd.n474 vdd.n473 185
R15149 vdd.n473 vdd.n325 185
R15150 vdd.n2997 vdd.n318 185
R15151 vdd.n3162 vdd.n318 185
R15152 vdd.n2996 vdd.n317 185
R15153 vdd.n3163 vdd.n317 185
R15154 vdd.n2995 vdd.n316 185
R15155 vdd.n3164 vdd.n316 185
R15156 vdd.n480 vdd.n476 185
R15157 vdd.n481 vdd.n480 185
R15158 vdd.n2991 vdd.n2990 185
R15159 vdd.n2990 vdd.n2989 185
R15160 vdd.n479 vdd.n478 185
R15161 vdd.n2980 vdd.n479 185
R15162 vdd.n2979 vdd.n2978 185
R15163 vdd.n2981 vdd.n2979 185
R15164 vdd.n488 vdd.n487 185
R15165 vdd.n493 vdd.n487 185
R15166 vdd.n2974 vdd.n2973 185
R15167 vdd.n2973 vdd.n2972 185
R15168 vdd.n491 vdd.n490 185
R15169 vdd.n492 vdd.n491 185
R15170 vdd.n2963 vdd.n2962 185
R15171 vdd.n2964 vdd.n2963 185
R15172 vdd.n501 vdd.n500 185
R15173 vdd.n500 vdd.n499 185
R15174 vdd.n2958 vdd.n2957 185
R15175 vdd.n2957 vdd.n2956 185
R15176 vdd.n504 vdd.n503 185
R15177 vdd.n505 vdd.n504 185
R15178 vdd.n2947 vdd.n2946 185
R15179 vdd.n2948 vdd.n2947 185
R15180 vdd.n513 vdd.n512 185
R15181 vdd.n512 vdd.n511 185
R15182 vdd.n2942 vdd.n2941 185
R15183 vdd.n2941 vdd.n2940 185
R15184 vdd.n741 vdd.n740 185
R15185 vdd.n2567 vdd.n2566 185
R15186 vdd.n2565 vdd.n2350 185
R15187 vdd.n2569 vdd.n2350 185
R15188 vdd.n2564 vdd.n2563 185
R15189 vdd.n2562 vdd.n2561 185
R15190 vdd.n2560 vdd.n2559 185
R15191 vdd.n2558 vdd.n2557 185
R15192 vdd.n2556 vdd.n2555 185
R15193 vdd.n2554 vdd.n2553 185
R15194 vdd.n2552 vdd.n2551 185
R15195 vdd.n2550 vdd.n2549 185
R15196 vdd.n2548 vdd.n2547 185
R15197 vdd.n2546 vdd.n2545 185
R15198 vdd.n2544 vdd.n2543 185
R15199 vdd.n2542 vdd.n2541 185
R15200 vdd.n2540 vdd.n2539 185
R15201 vdd.n2538 vdd.n2537 185
R15202 vdd.n2536 vdd.n2535 185
R15203 vdd.n2534 vdd.n2533 185
R15204 vdd.n2532 vdd.n2531 185
R15205 vdd.n2530 vdd.n2529 185
R15206 vdd.n2528 vdd.n2527 185
R15207 vdd.n2526 vdd.n2525 185
R15208 vdd.n2524 vdd.n2523 185
R15209 vdd.n2522 vdd.n2521 185
R15210 vdd.n2520 vdd.n2519 185
R15211 vdd.n2518 vdd.n2517 185
R15212 vdd.n2516 vdd.n2515 185
R15213 vdd.n2514 vdd.n2513 185
R15214 vdd.n2512 vdd.n2511 185
R15215 vdd.n2510 vdd.n2509 185
R15216 vdd.n2508 vdd.n2507 185
R15217 vdd.n2505 vdd.n2504 185
R15218 vdd.n2503 vdd.n2502 185
R15219 vdd.n2501 vdd.n2500 185
R15220 vdd.n2708 vdd.n2707 185
R15221 vdd.n2709 vdd.n660 185
R15222 vdd.n2711 vdd.n2710 185
R15223 vdd.n2713 vdd.n658 185
R15224 vdd.n2715 vdd.n2714 185
R15225 vdd.n2716 vdd.n657 185
R15226 vdd.n2718 vdd.n2717 185
R15227 vdd.n2720 vdd.n655 185
R15228 vdd.n2722 vdd.n2721 185
R15229 vdd.n2723 vdd.n654 185
R15230 vdd.n2725 vdd.n2724 185
R15231 vdd.n2727 vdd.n652 185
R15232 vdd.n2729 vdd.n2728 185
R15233 vdd.n2730 vdd.n651 185
R15234 vdd.n2732 vdd.n2731 185
R15235 vdd.n2734 vdd.n649 185
R15236 vdd.n2736 vdd.n2735 185
R15237 vdd.n2738 vdd.n648 185
R15238 vdd.n2740 vdd.n2739 185
R15239 vdd.n2742 vdd.n646 185
R15240 vdd.n2744 vdd.n2743 185
R15241 vdd.n2745 vdd.n645 185
R15242 vdd.n2747 vdd.n2746 185
R15243 vdd.n2749 vdd.n643 185
R15244 vdd.n2751 vdd.n2750 185
R15245 vdd.n2752 vdd.n642 185
R15246 vdd.n2754 vdd.n2753 185
R15247 vdd.n2756 vdd.n640 185
R15248 vdd.n2758 vdd.n2757 185
R15249 vdd.n2759 vdd.n639 185
R15250 vdd.n2761 vdd.n2760 185
R15251 vdd.n2763 vdd.n638 185
R15252 vdd.n2764 vdd.n637 185
R15253 vdd.n2767 vdd.n2766 185
R15254 vdd.n2768 vdd.n635 185
R15255 vdd.n635 vdd.n613 185
R15256 vdd.n2705 vdd.n632 185
R15257 vdd.n2771 vdd.n632 185
R15258 vdd.n2704 vdd.n2703 185
R15259 vdd.n2703 vdd.n631 185
R15260 vdd.n2702 vdd.n664 185
R15261 vdd.n2702 vdd.n2701 185
R15262 vdd.n2456 vdd.n665 185
R15263 vdd.n674 vdd.n665 185
R15264 vdd.n2457 vdd.n672 185
R15265 vdd.n2695 vdd.n672 185
R15266 vdd.n2459 vdd.n2458 185
R15267 vdd.n2458 vdd.n671 185
R15268 vdd.n2460 vdd.n680 185
R15269 vdd.n2644 vdd.n680 185
R15270 vdd.n2462 vdd.n2461 185
R15271 vdd.n2461 vdd.n679 185
R15272 vdd.n2463 vdd.n686 185
R15273 vdd.n2638 vdd.n686 185
R15274 vdd.n2465 vdd.n2464 185
R15275 vdd.n2464 vdd.n685 185
R15276 vdd.n2466 vdd.n691 185
R15277 vdd.n2630 vdd.n691 185
R15278 vdd.n2468 vdd.n2467 185
R15279 vdd.n2467 vdd.n698 185
R15280 vdd.n2469 vdd.n696 185
R15281 vdd.n2624 vdd.n696 185
R15282 vdd.n2471 vdd.n2470 185
R15283 vdd.n2472 vdd.n2471 185
R15284 vdd.n2455 vdd.n703 185
R15285 vdd.n2618 vdd.n703 185
R15286 vdd.n2454 vdd.n2453 185
R15287 vdd.n2453 vdd.n702 185
R15288 vdd.n2452 vdd.n709 185
R15289 vdd.n2612 vdd.n709 185
R15290 vdd.n2451 vdd.n2450 185
R15291 vdd.n2450 vdd.n708 185
R15292 vdd.n2449 vdd.n714 185
R15293 vdd.n2606 vdd.n714 185
R15294 vdd.n2448 vdd.n2447 185
R15295 vdd.n2447 vdd.n721 185
R15296 vdd.n2446 vdd.n719 185
R15297 vdd.n2600 vdd.n719 185
R15298 vdd.n2445 vdd.n2444 185
R15299 vdd.n2444 vdd.n728 185
R15300 vdd.n2443 vdd.n726 185
R15301 vdd.n2594 vdd.n726 185
R15302 vdd.n2442 vdd.n2441 185
R15303 vdd.n2441 vdd.n725 185
R15304 vdd.n2353 vdd.n732 185
R15305 vdd.n2588 vdd.n732 185
R15306 vdd.n2495 vdd.n2494 185
R15307 vdd.n2494 vdd.n2493 185
R15308 vdd.n2496 vdd.n737 185
R15309 vdd.n2582 vdd.n737 185
R15310 vdd.n2498 vdd.n2497 185
R15311 vdd.n2497 vdd.t170 185
R15312 vdd.n2499 vdd.n742 185
R15313 vdd.n2576 vdd.n742 185
R15314 vdd.n2578 vdd.n2577 185
R15315 vdd.n2577 vdd.n2576 185
R15316 vdd.n2579 vdd.n739 185
R15317 vdd.n739 vdd.t170 185
R15318 vdd.n2581 vdd.n2580 185
R15319 vdd.n2582 vdd.n2581 185
R15320 vdd.n731 vdd.n730 185
R15321 vdd.n2493 vdd.n731 185
R15322 vdd.n2590 vdd.n2589 185
R15323 vdd.n2589 vdd.n2588 185
R15324 vdd.n2591 vdd.n729 185
R15325 vdd.n729 vdd.n725 185
R15326 vdd.n2593 vdd.n2592 185
R15327 vdd.n2594 vdd.n2593 185
R15328 vdd.n718 vdd.n717 185
R15329 vdd.n728 vdd.n718 185
R15330 vdd.n2602 vdd.n2601 185
R15331 vdd.n2601 vdd.n2600 185
R15332 vdd.n2603 vdd.n716 185
R15333 vdd.n721 vdd.n716 185
R15334 vdd.n2605 vdd.n2604 185
R15335 vdd.n2606 vdd.n2605 185
R15336 vdd.n707 vdd.n706 185
R15337 vdd.n708 vdd.n707 185
R15338 vdd.n2614 vdd.n2613 185
R15339 vdd.n2613 vdd.n2612 185
R15340 vdd.n2615 vdd.n705 185
R15341 vdd.n705 vdd.n702 185
R15342 vdd.n2617 vdd.n2616 185
R15343 vdd.n2618 vdd.n2617 185
R15344 vdd.n695 vdd.n694 185
R15345 vdd.n2472 vdd.n695 185
R15346 vdd.n2626 vdd.n2625 185
R15347 vdd.n2625 vdd.n2624 185
R15348 vdd.n2627 vdd.n693 185
R15349 vdd.n698 vdd.n693 185
R15350 vdd.n2629 vdd.n2628 185
R15351 vdd.n2630 vdd.n2629 185
R15352 vdd.n684 vdd.n683 185
R15353 vdd.n685 vdd.n684 185
R15354 vdd.n2640 vdd.n2639 185
R15355 vdd.n2639 vdd.n2638 185
R15356 vdd.n2641 vdd.n682 185
R15357 vdd.n682 vdd.n679 185
R15358 vdd.n2643 vdd.n2642 185
R15359 vdd.n2644 vdd.n2643 185
R15360 vdd.n670 vdd.n669 185
R15361 vdd.n671 vdd.n670 185
R15362 vdd.n2697 vdd.n2696 185
R15363 vdd.n2696 vdd.n2695 185
R15364 vdd.n2698 vdd.n668 185
R15365 vdd.n674 vdd.n668 185
R15366 vdd.n2700 vdd.n2699 185
R15367 vdd.n2701 vdd.n2700 185
R15368 vdd.n636 vdd.n634 185
R15369 vdd.n634 vdd.n631 185
R15370 vdd.n2770 vdd.n2769 185
R15371 vdd.n2771 vdd.n2770 185
R15372 vdd.n2243 vdd.n2242 185
R15373 vdd.n2244 vdd.n2243 185
R15374 vdd.n792 vdd.n790 185
R15375 vdd.n790 vdd.t144 185
R15376 vdd.n2158 vdd.n799 185
R15377 vdd.n2169 vdd.n799 185
R15378 vdd.n2159 vdd.n808 185
R15379 vdd.n1868 vdd.n808 185
R15380 vdd.n2161 vdd.n2160 185
R15381 vdd.n2162 vdd.n2161 185
R15382 vdd.n2157 vdd.n807 185
R15383 vdd.n807 vdd.n804 185
R15384 vdd.n2156 vdd.n2155 185
R15385 vdd.n2155 vdd.n2154 185
R15386 vdd.n810 vdd.n809 185
R15387 vdd.n811 vdd.n810 185
R15388 vdd.n2147 vdd.n2146 185
R15389 vdd.n2148 vdd.n2147 185
R15390 vdd.n2145 vdd.n820 185
R15391 vdd.n820 vdd.n817 185
R15392 vdd.n2144 vdd.n2143 185
R15393 vdd.n2143 vdd.n2142 185
R15394 vdd.n822 vdd.n821 185
R15395 vdd.n830 vdd.n822 185
R15396 vdd.n2135 vdd.n2134 185
R15397 vdd.n2136 vdd.n2135 185
R15398 vdd.n2133 vdd.n831 185
R15399 vdd.n836 vdd.n831 185
R15400 vdd.n2132 vdd.n2131 185
R15401 vdd.n2131 vdd.n2130 185
R15402 vdd.n833 vdd.n832 185
R15403 vdd.n1969 vdd.n833 185
R15404 vdd.n2123 vdd.n2122 185
R15405 vdd.n2124 vdd.n2123 185
R15406 vdd.n2121 vdd.n843 185
R15407 vdd.n843 vdd.n840 185
R15408 vdd.n2120 vdd.n2119 185
R15409 vdd.n2119 vdd.n2118 185
R15410 vdd.n845 vdd.n844 185
R15411 vdd.n846 vdd.n845 185
R15412 vdd.n2111 vdd.n2110 185
R15413 vdd.n2112 vdd.n2111 185
R15414 vdd.n2108 vdd.n854 185
R15415 vdd.n861 vdd.n854 185
R15416 vdd.n2107 vdd.n2106 185
R15417 vdd.n2106 vdd.n2105 185
R15418 vdd.n857 vdd.n856 185
R15419 vdd.n858 vdd.n857 185
R15420 vdd.n2098 vdd.n2097 185
R15421 vdd.n2099 vdd.n2098 185
R15422 vdd.n2096 vdd.n868 185
R15423 vdd.n868 vdd.n865 185
R15424 vdd.n2095 vdd.n2094 185
R15425 vdd.n2094 vdd.n2093 185
R15426 vdd.n870 vdd.n869 185
R15427 vdd.n871 vdd.n870 185
R15428 vdd.n2086 vdd.n2085 185
R15429 vdd.n2087 vdd.n2086 185
R15430 vdd.n2174 vdd.n764 185
R15431 vdd.n2316 vdd.n764 185
R15432 vdd.n2176 vdd.n2175 185
R15433 vdd.n2178 vdd.n2177 185
R15434 vdd.n2180 vdd.n2179 185
R15435 vdd.n2182 vdd.n2181 185
R15436 vdd.n2184 vdd.n2183 185
R15437 vdd.n2186 vdd.n2185 185
R15438 vdd.n2188 vdd.n2187 185
R15439 vdd.n2190 vdd.n2189 185
R15440 vdd.n2192 vdd.n2191 185
R15441 vdd.n2194 vdd.n2193 185
R15442 vdd.n2196 vdd.n2195 185
R15443 vdd.n2198 vdd.n2197 185
R15444 vdd.n2200 vdd.n2199 185
R15445 vdd.n2202 vdd.n2201 185
R15446 vdd.n2204 vdd.n2203 185
R15447 vdd.n2206 vdd.n2205 185
R15448 vdd.n2208 vdd.n2207 185
R15449 vdd.n2210 vdd.n2209 185
R15450 vdd.n2212 vdd.n2211 185
R15451 vdd.n2214 vdd.n2213 185
R15452 vdd.n2216 vdd.n2215 185
R15453 vdd.n2218 vdd.n2217 185
R15454 vdd.n2220 vdd.n2219 185
R15455 vdd.n2222 vdd.n2221 185
R15456 vdd.n2224 vdd.n2223 185
R15457 vdd.n2226 vdd.n2225 185
R15458 vdd.n2228 vdd.n2227 185
R15459 vdd.n2230 vdd.n2229 185
R15460 vdd.n2232 vdd.n2231 185
R15461 vdd.n2234 vdd.n2233 185
R15462 vdd.n2236 vdd.n2235 185
R15463 vdd.n2238 vdd.n2237 185
R15464 vdd.n2240 vdd.n2239 185
R15465 vdd.n2241 vdd.n791 185
R15466 vdd.n2173 vdd.n789 185
R15467 vdd.n2244 vdd.n789 185
R15468 vdd.n2172 vdd.n2171 185
R15469 vdd.n2171 vdd.t144 185
R15470 vdd.n2170 vdd.n796 185
R15471 vdd.n2170 vdd.n2169 185
R15472 vdd.n1950 vdd.n797 185
R15473 vdd.n1868 vdd.n797 185
R15474 vdd.n1951 vdd.n806 185
R15475 vdd.n2162 vdd.n806 185
R15476 vdd.n1953 vdd.n1952 185
R15477 vdd.n1952 vdd.n804 185
R15478 vdd.n1954 vdd.n813 185
R15479 vdd.n2154 vdd.n813 185
R15480 vdd.n1956 vdd.n1955 185
R15481 vdd.n1955 vdd.n811 185
R15482 vdd.n1957 vdd.n819 185
R15483 vdd.n2148 vdd.n819 185
R15484 vdd.n1959 vdd.n1958 185
R15485 vdd.n1958 vdd.n817 185
R15486 vdd.n1960 vdd.n824 185
R15487 vdd.n2142 vdd.n824 185
R15488 vdd.n1962 vdd.n1961 185
R15489 vdd.n1961 vdd.n830 185
R15490 vdd.n1963 vdd.n829 185
R15491 vdd.n2136 vdd.n829 185
R15492 vdd.n1965 vdd.n1964 185
R15493 vdd.n1964 vdd.n836 185
R15494 vdd.n1966 vdd.n835 185
R15495 vdd.n2130 vdd.n835 185
R15496 vdd.n1968 vdd.n1967 185
R15497 vdd.n1969 vdd.n1968 185
R15498 vdd.n1949 vdd.n842 185
R15499 vdd.n2124 vdd.n842 185
R15500 vdd.n1948 vdd.n1947 185
R15501 vdd.n1947 vdd.n840 185
R15502 vdd.n1946 vdd.n848 185
R15503 vdd.n2118 vdd.n848 185
R15504 vdd.n1945 vdd.n1944 185
R15505 vdd.n1944 vdd.n846 185
R15506 vdd.n1943 vdd.n853 185
R15507 vdd.n2112 vdd.n853 185
R15508 vdd.n1942 vdd.n1941 185
R15509 vdd.n1941 vdd.n861 185
R15510 vdd.n1940 vdd.n860 185
R15511 vdd.n2105 vdd.n860 185
R15512 vdd.n1939 vdd.n1938 185
R15513 vdd.n1938 vdd.n858 185
R15514 vdd.n1937 vdd.n867 185
R15515 vdd.n2099 vdd.n867 185
R15516 vdd.n1936 vdd.n1935 185
R15517 vdd.n1935 vdd.n865 185
R15518 vdd.n1934 vdd.n873 185
R15519 vdd.n2093 vdd.n873 185
R15520 vdd.n1933 vdd.n1932 185
R15521 vdd.n1932 vdd.n871 185
R15522 vdd.n1931 vdd.n879 185
R15523 vdd.n2087 vdd.n879 185
R15524 vdd.n2084 vdd.n880 185
R15525 vdd.n2083 vdd.n2082 185
R15526 vdd.n2080 vdd.n881 185
R15527 vdd.n2078 vdd.n2077 185
R15528 vdd.n2076 vdd.n882 185
R15529 vdd.n2075 vdd.n2074 185
R15530 vdd.n2072 vdd.n883 185
R15531 vdd.n2070 vdd.n2069 185
R15532 vdd.n2068 vdd.n884 185
R15533 vdd.n2067 vdd.n2066 185
R15534 vdd.n2064 vdd.n885 185
R15535 vdd.n2062 vdd.n2061 185
R15536 vdd.n2060 vdd.n886 185
R15537 vdd.n2059 vdd.n2058 185
R15538 vdd.n2056 vdd.n887 185
R15539 vdd.n2054 vdd.n2053 185
R15540 vdd.n2052 vdd.n888 185
R15541 vdd.n2051 vdd.n890 185
R15542 vdd.n1896 vdd.n891 185
R15543 vdd.n1899 vdd.n1898 185
R15544 vdd.n1901 vdd.n1900 185
R15545 vdd.n1903 vdd.n1895 185
R15546 vdd.n1906 vdd.n1905 185
R15547 vdd.n1907 vdd.n1894 185
R15548 vdd.n1909 vdd.n1908 185
R15549 vdd.n1911 vdd.n1893 185
R15550 vdd.n1914 vdd.n1913 185
R15551 vdd.n1915 vdd.n1892 185
R15552 vdd.n1917 vdd.n1916 185
R15553 vdd.n1919 vdd.n1891 185
R15554 vdd.n1922 vdd.n1921 185
R15555 vdd.n1923 vdd.n1888 185
R15556 vdd.n1926 vdd.n1925 185
R15557 vdd.n1928 vdd.n1887 185
R15558 vdd.n1930 vdd.n1929 185
R15559 vdd.n1929 vdd.n877 185
R15560 vdd.n303 vdd.n302 171.744
R15561 vdd.n302 vdd.n301 171.744
R15562 vdd.n301 vdd.n270 171.744
R15563 vdd.n294 vdd.n270 171.744
R15564 vdd.n294 vdd.n293 171.744
R15565 vdd.n293 vdd.n275 171.744
R15566 vdd.n286 vdd.n275 171.744
R15567 vdd.n286 vdd.n285 171.744
R15568 vdd.n285 vdd.n279 171.744
R15569 vdd.n252 vdd.n251 171.744
R15570 vdd.n251 vdd.n250 171.744
R15571 vdd.n250 vdd.n219 171.744
R15572 vdd.n243 vdd.n219 171.744
R15573 vdd.n243 vdd.n242 171.744
R15574 vdd.n242 vdd.n224 171.744
R15575 vdd.n235 vdd.n224 171.744
R15576 vdd.n235 vdd.n234 171.744
R15577 vdd.n234 vdd.n228 171.744
R15578 vdd.n209 vdd.n208 171.744
R15579 vdd.n208 vdd.n207 171.744
R15580 vdd.n207 vdd.n176 171.744
R15581 vdd.n200 vdd.n176 171.744
R15582 vdd.n200 vdd.n199 171.744
R15583 vdd.n199 vdd.n181 171.744
R15584 vdd.n192 vdd.n181 171.744
R15585 vdd.n192 vdd.n191 171.744
R15586 vdd.n191 vdd.n185 171.744
R15587 vdd.n158 vdd.n157 171.744
R15588 vdd.n157 vdd.n156 171.744
R15589 vdd.n156 vdd.n125 171.744
R15590 vdd.n149 vdd.n125 171.744
R15591 vdd.n149 vdd.n148 171.744
R15592 vdd.n148 vdd.n130 171.744
R15593 vdd.n141 vdd.n130 171.744
R15594 vdd.n141 vdd.n140 171.744
R15595 vdd.n140 vdd.n134 171.744
R15596 vdd.n116 vdd.n115 171.744
R15597 vdd.n115 vdd.n114 171.744
R15598 vdd.n114 vdd.n83 171.744
R15599 vdd.n107 vdd.n83 171.744
R15600 vdd.n107 vdd.n106 171.744
R15601 vdd.n106 vdd.n88 171.744
R15602 vdd.n99 vdd.n88 171.744
R15603 vdd.n99 vdd.n98 171.744
R15604 vdd.n98 vdd.n92 171.744
R15605 vdd.n65 vdd.n64 171.744
R15606 vdd.n64 vdd.n63 171.744
R15607 vdd.n63 vdd.n32 171.744
R15608 vdd.n56 vdd.n32 171.744
R15609 vdd.n56 vdd.n55 171.744
R15610 vdd.n55 vdd.n37 171.744
R15611 vdd.n48 vdd.n37 171.744
R15612 vdd.n48 vdd.n47 171.744
R15613 vdd.n47 vdd.n41 171.744
R15614 vdd.n1498 vdd.n1497 171.744
R15615 vdd.n1497 vdd.n1496 171.744
R15616 vdd.n1496 vdd.n1465 171.744
R15617 vdd.n1489 vdd.n1465 171.744
R15618 vdd.n1489 vdd.n1488 171.744
R15619 vdd.n1488 vdd.n1470 171.744
R15620 vdd.n1481 vdd.n1470 171.744
R15621 vdd.n1481 vdd.n1480 171.744
R15622 vdd.n1480 vdd.n1474 171.744
R15623 vdd.n1549 vdd.n1548 171.744
R15624 vdd.n1548 vdd.n1547 171.744
R15625 vdd.n1547 vdd.n1516 171.744
R15626 vdd.n1540 vdd.n1516 171.744
R15627 vdd.n1540 vdd.n1539 171.744
R15628 vdd.n1539 vdd.n1521 171.744
R15629 vdd.n1532 vdd.n1521 171.744
R15630 vdd.n1532 vdd.n1531 171.744
R15631 vdd.n1531 vdd.n1525 171.744
R15632 vdd.n1404 vdd.n1403 171.744
R15633 vdd.n1403 vdd.n1402 171.744
R15634 vdd.n1402 vdd.n1371 171.744
R15635 vdd.n1395 vdd.n1371 171.744
R15636 vdd.n1395 vdd.n1394 171.744
R15637 vdd.n1394 vdd.n1376 171.744
R15638 vdd.n1387 vdd.n1376 171.744
R15639 vdd.n1387 vdd.n1386 171.744
R15640 vdd.n1386 vdd.n1380 171.744
R15641 vdd.n1455 vdd.n1454 171.744
R15642 vdd.n1454 vdd.n1453 171.744
R15643 vdd.n1453 vdd.n1422 171.744
R15644 vdd.n1446 vdd.n1422 171.744
R15645 vdd.n1446 vdd.n1445 171.744
R15646 vdd.n1445 vdd.n1427 171.744
R15647 vdd.n1438 vdd.n1427 171.744
R15648 vdd.n1438 vdd.n1437 171.744
R15649 vdd.n1437 vdd.n1431 171.744
R15650 vdd.n1311 vdd.n1310 171.744
R15651 vdd.n1310 vdd.n1309 171.744
R15652 vdd.n1309 vdd.n1278 171.744
R15653 vdd.n1302 vdd.n1278 171.744
R15654 vdd.n1302 vdd.n1301 171.744
R15655 vdd.n1301 vdd.n1283 171.744
R15656 vdd.n1294 vdd.n1283 171.744
R15657 vdd.n1294 vdd.n1293 171.744
R15658 vdd.n1293 vdd.n1287 171.744
R15659 vdd.n1362 vdd.n1361 171.744
R15660 vdd.n1361 vdd.n1360 171.744
R15661 vdd.n1360 vdd.n1329 171.744
R15662 vdd.n1353 vdd.n1329 171.744
R15663 vdd.n1353 vdd.n1352 171.744
R15664 vdd.n1352 vdd.n1334 171.744
R15665 vdd.n1345 vdd.n1334 171.744
R15666 vdd.n1345 vdd.n1344 171.744
R15667 vdd.n1344 vdd.n1338 171.744
R15668 vdd.n3130 vdd.n356 146.341
R15669 vdd.n3128 vdd.n3127 146.341
R15670 vdd.n3125 vdd.n360 146.341
R15671 vdd.n3121 vdd.n3120 146.341
R15672 vdd.n3118 vdd.n368 146.341
R15673 vdd.n3114 vdd.n3113 146.341
R15674 vdd.n3111 vdd.n375 146.341
R15675 vdd.n3107 vdd.n3106 146.341
R15676 vdd.n3104 vdd.n382 146.341
R15677 vdd.n393 vdd.n390 146.341
R15678 vdd.n3096 vdd.n3095 146.341
R15679 vdd.n3093 vdd.n395 146.341
R15680 vdd.n3089 vdd.n3088 146.341
R15681 vdd.n3086 vdd.n401 146.341
R15682 vdd.n3082 vdd.n3081 146.341
R15683 vdd.n3079 vdd.n408 146.341
R15684 vdd.n3075 vdd.n3074 146.341
R15685 vdd.n3072 vdd.n415 146.341
R15686 vdd.n3068 vdd.n3067 146.341
R15687 vdd.n3065 vdd.n422 146.341
R15688 vdd.n433 vdd.n430 146.341
R15689 vdd.n3057 vdd.n3056 146.341
R15690 vdd.n3054 vdd.n435 146.341
R15691 vdd.n3050 vdd.n3049 146.341
R15692 vdd.n3047 vdd.n441 146.341
R15693 vdd.n3043 vdd.n3042 146.341
R15694 vdd.n3040 vdd.n448 146.341
R15695 vdd.n3036 vdd.n3035 146.341
R15696 vdd.n3033 vdd.n455 146.341
R15697 vdd.n3029 vdd.n3028 146.341
R15698 vdd.n3026 vdd.n462 146.341
R15699 vdd.n2941 vdd.n512 146.341
R15700 vdd.n2947 vdd.n512 146.341
R15701 vdd.n2947 vdd.n504 146.341
R15702 vdd.n2957 vdd.n504 146.341
R15703 vdd.n2957 vdd.n500 146.341
R15704 vdd.n2963 vdd.n500 146.341
R15705 vdd.n2963 vdd.n491 146.341
R15706 vdd.n2973 vdd.n491 146.341
R15707 vdd.n2973 vdd.n487 146.341
R15708 vdd.n2979 vdd.n487 146.341
R15709 vdd.n2979 vdd.n479 146.341
R15710 vdd.n2990 vdd.n479 146.341
R15711 vdd.n2990 vdd.n480 146.341
R15712 vdd.n480 vdd.n316 146.341
R15713 vdd.n317 vdd.n316 146.341
R15714 vdd.n318 vdd.n317 146.341
R15715 vdd.n473 vdd.n318 146.341
R15716 vdd.n473 vdd.n326 146.341
R15717 vdd.n327 vdd.n326 146.341
R15718 vdd.n328 vdd.n327 146.341
R15719 vdd.n470 vdd.n328 146.341
R15720 vdd.n470 vdd.n337 146.341
R15721 vdd.n338 vdd.n337 146.341
R15722 vdd.n339 vdd.n338 146.341
R15723 vdd.n467 vdd.n339 146.341
R15724 vdd.n467 vdd.n348 146.341
R15725 vdd.n349 vdd.n348 146.341
R15726 vdd.n350 vdd.n349 146.341
R15727 vdd.n2933 vdd.n2931 146.341
R15728 vdd.n2931 vdd.n2930 146.341
R15729 vdd.n2927 vdd.n2926 146.341
R15730 vdd.n2923 vdd.n2922 146.341
R15731 vdd.n2920 vdd.n526 146.341
R15732 vdd.n2916 vdd.n2914 146.341
R15733 vdd.n2912 vdd.n532 146.341
R15734 vdd.n2908 vdd.n2906 146.341
R15735 vdd.n2904 vdd.n538 146.341
R15736 vdd.n2900 vdd.n2898 146.341
R15737 vdd.n2896 vdd.n546 146.341
R15738 vdd.n2892 vdd.n2890 146.341
R15739 vdd.n2888 vdd.n552 146.341
R15740 vdd.n2884 vdd.n2882 146.341
R15741 vdd.n2880 vdd.n558 146.341
R15742 vdd.n2876 vdd.n2874 146.341
R15743 vdd.n2872 vdd.n564 146.341
R15744 vdd.n2868 vdd.n2866 146.341
R15745 vdd.n2864 vdd.n570 146.341
R15746 vdd.n2860 vdd.n2858 146.341
R15747 vdd.n2856 vdd.n576 146.341
R15748 vdd.n2849 vdd.n585 146.341
R15749 vdd.n2847 vdd.n2846 146.341
R15750 vdd.n2843 vdd.n2842 146.341
R15751 vdd.n2840 vdd.n590 146.341
R15752 vdd.n2836 vdd.n2834 146.341
R15753 vdd.n2832 vdd.n596 146.341
R15754 vdd.n2828 vdd.n2826 146.341
R15755 vdd.n2824 vdd.n602 146.341
R15756 vdd.n2820 vdd.n2818 146.341
R15757 vdd.n2815 vdd.n2814 146.341
R15758 vdd.n2811 vdd.n515 146.341
R15759 vdd.n2939 vdd.n510 146.341
R15760 vdd.n2949 vdd.n510 146.341
R15761 vdd.n2949 vdd.n506 146.341
R15762 vdd.n2955 vdd.n506 146.341
R15763 vdd.n2955 vdd.n498 146.341
R15764 vdd.n2965 vdd.n498 146.341
R15765 vdd.n2965 vdd.n494 146.341
R15766 vdd.n2971 vdd.n494 146.341
R15767 vdd.n2971 vdd.n486 146.341
R15768 vdd.n2982 vdd.n486 146.341
R15769 vdd.n2982 vdd.n482 146.341
R15770 vdd.n2988 vdd.n482 146.341
R15771 vdd.n2988 vdd.n314 146.341
R15772 vdd.n3165 vdd.n314 146.341
R15773 vdd.n3165 vdd.n315 146.341
R15774 vdd.n3161 vdd.n315 146.341
R15775 vdd.n3161 vdd.n319 146.341
R15776 vdd.n3157 vdd.n319 146.341
R15777 vdd.n3157 vdd.n324 146.341
R15778 vdd.n3153 vdd.n324 146.341
R15779 vdd.n3153 vdd.n330 146.341
R15780 vdd.n3149 vdd.n330 146.341
R15781 vdd.n3149 vdd.n336 146.341
R15782 vdd.n3145 vdd.n336 146.341
R15783 vdd.n3145 vdd.n341 146.341
R15784 vdd.n3141 vdd.n341 146.341
R15785 vdd.n3141 vdd.n347 146.341
R15786 vdd.n3137 vdd.n347 146.341
R15787 vdd.n2034 vdd.n2033 146.341
R15788 vdd.n2031 vdd.n1615 146.341
R15789 vdd.n1811 vdd.n1621 146.341
R15790 vdd.n1809 vdd.n1808 146.341
R15791 vdd.n1806 vdd.n1623 146.341
R15792 vdd.n1802 vdd.n1801 146.341
R15793 vdd.n1799 vdd.n1630 146.341
R15794 vdd.n1795 vdd.n1794 146.341
R15795 vdd.n1792 vdd.n1637 146.341
R15796 vdd.n1648 vdd.n1645 146.341
R15797 vdd.n1784 vdd.n1783 146.341
R15798 vdd.n1781 vdd.n1650 146.341
R15799 vdd.n1777 vdd.n1776 146.341
R15800 vdd.n1774 vdd.n1656 146.341
R15801 vdd.n1770 vdd.n1769 146.341
R15802 vdd.n1767 vdd.n1663 146.341
R15803 vdd.n1763 vdd.n1762 146.341
R15804 vdd.n1760 vdd.n1670 146.341
R15805 vdd.n1756 vdd.n1755 146.341
R15806 vdd.n1753 vdd.n1677 146.341
R15807 vdd.n1688 vdd.n1685 146.341
R15808 vdd.n1745 vdd.n1744 146.341
R15809 vdd.n1742 vdd.n1690 146.341
R15810 vdd.n1738 vdd.n1737 146.341
R15811 vdd.n1735 vdd.n1696 146.341
R15812 vdd.n1731 vdd.n1730 146.341
R15813 vdd.n1728 vdd.n1703 146.341
R15814 vdd.n1724 vdd.n1723 146.341
R15815 vdd.n1721 vdd.n1718 146.341
R15816 vdd.n1716 vdd.n1713 146.341
R15817 vdd.n1711 vdd.n897 146.341
R15818 vdd.n1216 vdd.n978 146.341
R15819 vdd.n1222 vdd.n978 146.341
R15820 vdd.n1222 vdd.n971 146.341
R15821 vdd.n1232 vdd.n971 146.341
R15822 vdd.n1232 vdd.n967 146.341
R15823 vdd.n1238 vdd.n967 146.341
R15824 vdd.n1238 vdd.n958 146.341
R15825 vdd.n1248 vdd.n958 146.341
R15826 vdd.n1248 vdd.n954 146.341
R15827 vdd.n1254 vdd.n954 146.341
R15828 vdd.n1254 vdd.n947 146.341
R15829 vdd.n1265 vdd.n947 146.341
R15830 vdd.n1265 vdd.n943 146.341
R15831 vdd.n1271 vdd.n943 146.341
R15832 vdd.n1271 vdd.n936 146.341
R15833 vdd.n1563 vdd.n936 146.341
R15834 vdd.n1563 vdd.n932 146.341
R15835 vdd.n1569 vdd.n932 146.341
R15836 vdd.n1569 vdd.n924 146.341
R15837 vdd.n1580 vdd.n924 146.341
R15838 vdd.n1580 vdd.n920 146.341
R15839 vdd.n1586 vdd.n920 146.341
R15840 vdd.n1586 vdd.n914 146.341
R15841 vdd.n1597 vdd.n914 146.341
R15842 vdd.n1597 vdd.n909 146.341
R15843 vdd.n1605 vdd.n909 146.341
R15844 vdd.n1605 vdd.n899 146.341
R15845 vdd.n2042 vdd.n899 146.341
R15846 vdd.n988 vdd.n987 146.341
R15847 vdd.n991 vdd.n988 146.341
R15848 vdd.n994 vdd.n993 146.341
R15849 vdd.n999 vdd.n996 146.341
R15850 vdd.n1002 vdd.n1001 146.341
R15851 vdd.n1007 vdd.n1004 146.341
R15852 vdd.n1010 vdd.n1009 146.341
R15853 vdd.n1015 vdd.n1012 146.341
R15854 vdd.n1018 vdd.n1017 146.341
R15855 vdd.n1025 vdd.n1020 146.341
R15856 vdd.n1028 vdd.n1027 146.341
R15857 vdd.n1033 vdd.n1030 146.341
R15858 vdd.n1036 vdd.n1035 146.341
R15859 vdd.n1041 vdd.n1038 146.341
R15860 vdd.n1044 vdd.n1043 146.341
R15861 vdd.n1049 vdd.n1046 146.341
R15862 vdd.n1052 vdd.n1051 146.341
R15863 vdd.n1057 vdd.n1054 146.341
R15864 vdd.n1060 vdd.n1059 146.341
R15865 vdd.n1065 vdd.n1062 146.341
R15866 vdd.n1146 vdd.n1067 146.341
R15867 vdd.n1144 vdd.n1143 146.341
R15868 vdd.n1074 vdd.n1073 146.341
R15869 vdd.n1077 vdd.n1076 146.341
R15870 vdd.n1082 vdd.n1081 146.341
R15871 vdd.n1085 vdd.n1084 146.341
R15872 vdd.n1090 vdd.n1089 146.341
R15873 vdd.n1093 vdd.n1092 146.341
R15874 vdd.n1098 vdd.n1097 146.341
R15875 vdd.n1101 vdd.n1100 146.341
R15876 vdd.n1106 vdd.n1105 146.341
R15877 vdd.n1108 vdd.n981 146.341
R15878 vdd.n1214 vdd.n977 146.341
R15879 vdd.n1224 vdd.n977 146.341
R15880 vdd.n1224 vdd.n973 146.341
R15881 vdd.n1230 vdd.n973 146.341
R15882 vdd.n1230 vdd.n965 146.341
R15883 vdd.n1240 vdd.n965 146.341
R15884 vdd.n1240 vdd.n961 146.341
R15885 vdd.n1246 vdd.n961 146.341
R15886 vdd.n1246 vdd.n953 146.341
R15887 vdd.n1257 vdd.n953 146.341
R15888 vdd.n1257 vdd.n949 146.341
R15889 vdd.n1263 vdd.n949 146.341
R15890 vdd.n1263 vdd.n942 146.341
R15891 vdd.n1273 vdd.n942 146.341
R15892 vdd.n1273 vdd.n938 146.341
R15893 vdd.n1561 vdd.n938 146.341
R15894 vdd.n1561 vdd.n930 146.341
R15895 vdd.n1572 vdd.n930 146.341
R15896 vdd.n1572 vdd.n926 146.341
R15897 vdd.n1578 vdd.n926 146.341
R15898 vdd.n1578 vdd.n919 146.341
R15899 vdd.n1589 vdd.n919 146.341
R15900 vdd.n1589 vdd.n915 146.341
R15901 vdd.n1595 vdd.n915 146.341
R15902 vdd.n1595 vdd.n907 146.341
R15903 vdd.n1608 vdd.n907 146.341
R15904 vdd.n1608 vdd.n902 146.341
R15905 vdd.n2040 vdd.n902 146.341
R15906 vdd.n901 vdd.n877 141.707
R15907 vdd.n613 vdd.n516 141.707
R15908 vdd.n1889 vdd.t100 127.284
R15909 vdd.n793 vdd.t84 127.284
R15910 vdd.n1863 vdd.t126 127.284
R15911 vdd.n785 vdd.t109 127.284
R15912 vdd.n2634 vdd.t71 127.284
R15913 vdd.n2634 vdd.t72 127.284
R15914 vdd.n2354 vdd.t107 127.284
R15915 vdd.n661 vdd.t88 127.284
R15916 vdd.n2351 vdd.t93 127.284
R15917 vdd.n625 vdd.t95 127.284
R15918 vdd.n855 vdd.t103 127.284
R15919 vdd.n855 vdd.t104 127.284
R15920 vdd.n22 vdd.n20 117.314
R15921 vdd.n17 vdd.n15 117.314
R15922 vdd.n27 vdd.n26 116.927
R15923 vdd.n24 vdd.n23 116.927
R15924 vdd.n22 vdd.n21 116.927
R15925 vdd.n17 vdd.n16 116.927
R15926 vdd.n19 vdd.n18 116.927
R15927 vdd.n27 vdd.n25 116.927
R15928 vdd.n1890 vdd.t99 111.188
R15929 vdd.n794 vdd.t85 111.188
R15930 vdd.n1864 vdd.t125 111.188
R15931 vdd.n786 vdd.t110 111.188
R15932 vdd.n2355 vdd.t106 111.188
R15933 vdd.n662 vdd.t89 111.188
R15934 vdd.n2352 vdd.t92 111.188
R15935 vdd.n626 vdd.t96 111.188
R15936 vdd.n2577 vdd.n739 99.5127
R15937 vdd.n2581 vdd.n739 99.5127
R15938 vdd.n2581 vdd.n731 99.5127
R15939 vdd.n2589 vdd.n731 99.5127
R15940 vdd.n2589 vdd.n729 99.5127
R15941 vdd.n2593 vdd.n729 99.5127
R15942 vdd.n2593 vdd.n718 99.5127
R15943 vdd.n2601 vdd.n718 99.5127
R15944 vdd.n2601 vdd.n716 99.5127
R15945 vdd.n2605 vdd.n716 99.5127
R15946 vdd.n2605 vdd.n707 99.5127
R15947 vdd.n2613 vdd.n707 99.5127
R15948 vdd.n2613 vdd.n705 99.5127
R15949 vdd.n2617 vdd.n705 99.5127
R15950 vdd.n2617 vdd.n695 99.5127
R15951 vdd.n2625 vdd.n695 99.5127
R15952 vdd.n2625 vdd.n693 99.5127
R15953 vdd.n2629 vdd.n693 99.5127
R15954 vdd.n2629 vdd.n684 99.5127
R15955 vdd.n2639 vdd.n684 99.5127
R15956 vdd.n2639 vdd.n682 99.5127
R15957 vdd.n2643 vdd.n682 99.5127
R15958 vdd.n2643 vdd.n670 99.5127
R15959 vdd.n2696 vdd.n670 99.5127
R15960 vdd.n2696 vdd.n668 99.5127
R15961 vdd.n2700 vdd.n668 99.5127
R15962 vdd.n2700 vdd.n634 99.5127
R15963 vdd.n2770 vdd.n634 99.5127
R15964 vdd.n2766 vdd.n635 99.5127
R15965 vdd.n2764 vdd.n2763 99.5127
R15966 vdd.n2761 vdd.n639 99.5127
R15967 vdd.n2757 vdd.n2756 99.5127
R15968 vdd.n2754 vdd.n642 99.5127
R15969 vdd.n2750 vdd.n2749 99.5127
R15970 vdd.n2747 vdd.n645 99.5127
R15971 vdd.n2743 vdd.n2742 99.5127
R15972 vdd.n2740 vdd.n648 99.5127
R15973 vdd.n2735 vdd.n2734 99.5127
R15974 vdd.n2732 vdd.n651 99.5127
R15975 vdd.n2728 vdd.n2727 99.5127
R15976 vdd.n2725 vdd.n654 99.5127
R15977 vdd.n2721 vdd.n2720 99.5127
R15978 vdd.n2718 vdd.n657 99.5127
R15979 vdd.n2714 vdd.n2713 99.5127
R15980 vdd.n2711 vdd.n660 99.5127
R15981 vdd.n2497 vdd.n742 99.5127
R15982 vdd.n2497 vdd.n737 99.5127
R15983 vdd.n2494 vdd.n737 99.5127
R15984 vdd.n2494 vdd.n732 99.5127
R15985 vdd.n2441 vdd.n732 99.5127
R15986 vdd.n2441 vdd.n726 99.5127
R15987 vdd.n2444 vdd.n726 99.5127
R15988 vdd.n2444 vdd.n719 99.5127
R15989 vdd.n2447 vdd.n719 99.5127
R15990 vdd.n2447 vdd.n714 99.5127
R15991 vdd.n2450 vdd.n714 99.5127
R15992 vdd.n2450 vdd.n709 99.5127
R15993 vdd.n2453 vdd.n709 99.5127
R15994 vdd.n2453 vdd.n703 99.5127
R15995 vdd.n2471 vdd.n703 99.5127
R15996 vdd.n2471 vdd.n696 99.5127
R15997 vdd.n2467 vdd.n696 99.5127
R15998 vdd.n2467 vdd.n691 99.5127
R15999 vdd.n2464 vdd.n691 99.5127
R16000 vdd.n2464 vdd.n686 99.5127
R16001 vdd.n2461 vdd.n686 99.5127
R16002 vdd.n2461 vdd.n680 99.5127
R16003 vdd.n2458 vdd.n680 99.5127
R16004 vdd.n2458 vdd.n672 99.5127
R16005 vdd.n672 vdd.n665 99.5127
R16006 vdd.n2702 vdd.n665 99.5127
R16007 vdd.n2703 vdd.n2702 99.5127
R16008 vdd.n2703 vdd.n632 99.5127
R16009 vdd.n2567 vdd.n2350 99.5127
R16010 vdd.n2563 vdd.n2350 99.5127
R16011 vdd.n2561 vdd.n2560 99.5127
R16012 vdd.n2557 vdd.n2556 99.5127
R16013 vdd.n2553 vdd.n2552 99.5127
R16014 vdd.n2549 vdd.n2548 99.5127
R16015 vdd.n2545 vdd.n2544 99.5127
R16016 vdd.n2541 vdd.n2540 99.5127
R16017 vdd.n2537 vdd.n2536 99.5127
R16018 vdd.n2533 vdd.n2532 99.5127
R16019 vdd.n2529 vdd.n2528 99.5127
R16020 vdd.n2525 vdd.n2524 99.5127
R16021 vdd.n2521 vdd.n2520 99.5127
R16022 vdd.n2517 vdd.n2516 99.5127
R16023 vdd.n2513 vdd.n2512 99.5127
R16024 vdd.n2509 vdd.n2508 99.5127
R16025 vdd.n2504 vdd.n2503 99.5127
R16026 vdd.n2315 vdd.n783 99.5127
R16027 vdd.n2311 vdd.n2310 99.5127
R16028 vdd.n2307 vdd.n2306 99.5127
R16029 vdd.n2303 vdd.n2302 99.5127
R16030 vdd.n2299 vdd.n2298 99.5127
R16031 vdd.n2295 vdd.n2294 99.5127
R16032 vdd.n2291 vdd.n2290 99.5127
R16033 vdd.n2287 vdd.n2286 99.5127
R16034 vdd.n2283 vdd.n2282 99.5127
R16035 vdd.n2279 vdd.n2278 99.5127
R16036 vdd.n2275 vdd.n2274 99.5127
R16037 vdd.n2271 vdd.n2270 99.5127
R16038 vdd.n2267 vdd.n2266 99.5127
R16039 vdd.n2263 vdd.n2262 99.5127
R16040 vdd.n2259 vdd.n2258 99.5127
R16041 vdd.n2255 vdd.n2254 99.5127
R16042 vdd.n2250 vdd.n2249 99.5127
R16043 vdd.n1988 vdd.n878 99.5127
R16044 vdd.n1988 vdd.n872 99.5127
R16045 vdd.n1985 vdd.n872 99.5127
R16046 vdd.n1985 vdd.n866 99.5127
R16047 vdd.n1982 vdd.n866 99.5127
R16048 vdd.n1982 vdd.n859 99.5127
R16049 vdd.n1979 vdd.n859 99.5127
R16050 vdd.n1979 vdd.n852 99.5127
R16051 vdd.n1976 vdd.n852 99.5127
R16052 vdd.n1976 vdd.n847 99.5127
R16053 vdd.n1973 vdd.n847 99.5127
R16054 vdd.n1973 vdd.n841 99.5127
R16055 vdd.n1970 vdd.n841 99.5127
R16056 vdd.n1970 vdd.n834 99.5127
R16057 vdd.n1884 vdd.n834 99.5127
R16058 vdd.n1884 vdd.n828 99.5127
R16059 vdd.n1881 vdd.n828 99.5127
R16060 vdd.n1881 vdd.n823 99.5127
R16061 vdd.n1878 vdd.n823 99.5127
R16062 vdd.n1878 vdd.n818 99.5127
R16063 vdd.n1875 vdd.n818 99.5127
R16064 vdd.n1875 vdd.n812 99.5127
R16065 vdd.n1872 vdd.n812 99.5127
R16066 vdd.n1872 vdd.n805 99.5127
R16067 vdd.n1869 vdd.n805 99.5127
R16068 vdd.n1869 vdd.n798 99.5127
R16069 vdd.n798 vdd.n788 99.5127
R16070 vdd.n2245 vdd.n788 99.5127
R16071 vdd.n1823 vdd.n1821 99.5127
R16072 vdd.n1827 vdd.n1821 99.5127
R16073 vdd.n1831 vdd.n1829 99.5127
R16074 vdd.n1835 vdd.n1819 99.5127
R16075 vdd.n1839 vdd.n1837 99.5127
R16076 vdd.n1843 vdd.n1817 99.5127
R16077 vdd.n1847 vdd.n1845 99.5127
R16078 vdd.n1851 vdd.n1815 99.5127
R16079 vdd.n1854 vdd.n1853 99.5127
R16080 vdd.n2024 vdd.n2022 99.5127
R16081 vdd.n2020 vdd.n1856 99.5127
R16082 vdd.n2016 vdd.n2014 99.5127
R16083 vdd.n2012 vdd.n1858 99.5127
R16084 vdd.n2008 vdd.n2006 99.5127
R16085 vdd.n2004 vdd.n1860 99.5127
R16086 vdd.n2000 vdd.n1998 99.5127
R16087 vdd.n1996 vdd.n1862 99.5127
R16088 vdd.n2088 vdd.n874 99.5127
R16089 vdd.n2092 vdd.n874 99.5127
R16090 vdd.n2092 vdd.n864 99.5127
R16091 vdd.n2100 vdd.n864 99.5127
R16092 vdd.n2100 vdd.n862 99.5127
R16093 vdd.n2104 vdd.n862 99.5127
R16094 vdd.n2104 vdd.n851 99.5127
R16095 vdd.n2113 vdd.n851 99.5127
R16096 vdd.n2113 vdd.n849 99.5127
R16097 vdd.n2117 vdd.n849 99.5127
R16098 vdd.n2117 vdd.n839 99.5127
R16099 vdd.n2125 vdd.n839 99.5127
R16100 vdd.n2125 vdd.n837 99.5127
R16101 vdd.n2129 vdd.n837 99.5127
R16102 vdd.n2129 vdd.n827 99.5127
R16103 vdd.n2137 vdd.n827 99.5127
R16104 vdd.n2137 vdd.n825 99.5127
R16105 vdd.n2141 vdd.n825 99.5127
R16106 vdd.n2141 vdd.n816 99.5127
R16107 vdd.n2149 vdd.n816 99.5127
R16108 vdd.n2149 vdd.n814 99.5127
R16109 vdd.n2153 vdd.n814 99.5127
R16110 vdd.n2153 vdd.n803 99.5127
R16111 vdd.n2163 vdd.n803 99.5127
R16112 vdd.n2163 vdd.n800 99.5127
R16113 vdd.n2168 vdd.n800 99.5127
R16114 vdd.n2168 vdd.n801 99.5127
R16115 vdd.n801 vdd.n782 99.5127
R16116 vdd.n2686 vdd.n2685 99.5127
R16117 vdd.n2683 vdd.n2649 99.5127
R16118 vdd.n2679 vdd.n2678 99.5127
R16119 vdd.n2676 vdd.n2652 99.5127
R16120 vdd.n2672 vdd.n2671 99.5127
R16121 vdd.n2669 vdd.n2655 99.5127
R16122 vdd.n2665 vdd.n2664 99.5127
R16123 vdd.n2662 vdd.n2659 99.5127
R16124 vdd.n2803 vdd.n612 99.5127
R16125 vdd.n2801 vdd.n2800 99.5127
R16126 vdd.n2798 vdd.n615 99.5127
R16127 vdd.n2794 vdd.n2793 99.5127
R16128 vdd.n2791 vdd.n618 99.5127
R16129 vdd.n2787 vdd.n2786 99.5127
R16130 vdd.n2784 vdd.n621 99.5127
R16131 vdd.n2780 vdd.n2779 99.5127
R16132 vdd.n2777 vdd.n624 99.5127
R16133 vdd.n2421 vdd.n743 99.5127
R16134 vdd.n2421 vdd.n738 99.5127
R16135 vdd.n2492 vdd.n738 99.5127
R16136 vdd.n2492 vdd.n733 99.5127
R16137 vdd.n2488 vdd.n733 99.5127
R16138 vdd.n2488 vdd.n727 99.5127
R16139 vdd.n2485 vdd.n727 99.5127
R16140 vdd.n2485 vdd.n720 99.5127
R16141 vdd.n2482 vdd.n720 99.5127
R16142 vdd.n2482 vdd.n715 99.5127
R16143 vdd.n2479 vdd.n715 99.5127
R16144 vdd.n2479 vdd.n710 99.5127
R16145 vdd.n2476 vdd.n710 99.5127
R16146 vdd.n2476 vdd.n704 99.5127
R16147 vdd.n2473 vdd.n704 99.5127
R16148 vdd.n2473 vdd.n697 99.5127
R16149 vdd.n2438 vdd.n697 99.5127
R16150 vdd.n2438 vdd.n692 99.5127
R16151 vdd.n2435 vdd.n692 99.5127
R16152 vdd.n2435 vdd.n687 99.5127
R16153 vdd.n2432 vdd.n687 99.5127
R16154 vdd.n2432 vdd.n681 99.5127
R16155 vdd.n2429 vdd.n681 99.5127
R16156 vdd.n2429 vdd.n673 99.5127
R16157 vdd.n2426 vdd.n673 99.5127
R16158 vdd.n2426 vdd.n666 99.5127
R16159 vdd.n666 vdd.n630 99.5127
R16160 vdd.n2772 vdd.n630 99.5127
R16161 vdd.n2571 vdd.n746 99.5127
R16162 vdd.n2359 vdd.n2358 99.5127
R16163 vdd.n2363 vdd.n2362 99.5127
R16164 vdd.n2367 vdd.n2366 99.5127
R16165 vdd.n2371 vdd.n2370 99.5127
R16166 vdd.n2375 vdd.n2374 99.5127
R16167 vdd.n2379 vdd.n2378 99.5127
R16168 vdd.n2383 vdd.n2382 99.5127
R16169 vdd.n2387 vdd.n2386 99.5127
R16170 vdd.n2391 vdd.n2390 99.5127
R16171 vdd.n2395 vdd.n2394 99.5127
R16172 vdd.n2399 vdd.n2398 99.5127
R16173 vdd.n2403 vdd.n2402 99.5127
R16174 vdd.n2407 vdd.n2406 99.5127
R16175 vdd.n2411 vdd.n2410 99.5127
R16176 vdd.n2415 vdd.n2414 99.5127
R16177 vdd.n2417 vdd.n2349 99.5127
R16178 vdd.n2575 vdd.n736 99.5127
R16179 vdd.n2583 vdd.n736 99.5127
R16180 vdd.n2583 vdd.n734 99.5127
R16181 vdd.n2587 vdd.n734 99.5127
R16182 vdd.n2587 vdd.n724 99.5127
R16183 vdd.n2595 vdd.n724 99.5127
R16184 vdd.n2595 vdd.n722 99.5127
R16185 vdd.n2599 vdd.n722 99.5127
R16186 vdd.n2599 vdd.n713 99.5127
R16187 vdd.n2607 vdd.n713 99.5127
R16188 vdd.n2607 vdd.n711 99.5127
R16189 vdd.n2611 vdd.n711 99.5127
R16190 vdd.n2611 vdd.n701 99.5127
R16191 vdd.n2619 vdd.n701 99.5127
R16192 vdd.n2619 vdd.n699 99.5127
R16193 vdd.n2623 vdd.n699 99.5127
R16194 vdd.n2623 vdd.n690 99.5127
R16195 vdd.n2631 vdd.n690 99.5127
R16196 vdd.n2631 vdd.n688 99.5127
R16197 vdd.n2637 vdd.n688 99.5127
R16198 vdd.n2637 vdd.n678 99.5127
R16199 vdd.n2645 vdd.n678 99.5127
R16200 vdd.n2645 vdd.n675 99.5127
R16201 vdd.n2694 vdd.n675 99.5127
R16202 vdd.n2694 vdd.n676 99.5127
R16203 vdd.n676 vdd.n667 99.5127
R16204 vdd.n2689 vdd.n667 99.5127
R16205 vdd.n2689 vdd.n633 99.5127
R16206 vdd.n2239 vdd.n2238 99.5127
R16207 vdd.n2235 vdd.n2234 99.5127
R16208 vdd.n2231 vdd.n2230 99.5127
R16209 vdd.n2227 vdd.n2226 99.5127
R16210 vdd.n2223 vdd.n2222 99.5127
R16211 vdd.n2219 vdd.n2218 99.5127
R16212 vdd.n2215 vdd.n2214 99.5127
R16213 vdd.n2211 vdd.n2210 99.5127
R16214 vdd.n2207 vdd.n2206 99.5127
R16215 vdd.n2203 vdd.n2202 99.5127
R16216 vdd.n2199 vdd.n2198 99.5127
R16217 vdd.n2195 vdd.n2194 99.5127
R16218 vdd.n2191 vdd.n2190 99.5127
R16219 vdd.n2187 vdd.n2186 99.5127
R16220 vdd.n2183 vdd.n2182 99.5127
R16221 vdd.n2179 vdd.n2178 99.5127
R16222 vdd.n2175 vdd.n764 99.5127
R16223 vdd.n1932 vdd.n879 99.5127
R16224 vdd.n1932 vdd.n873 99.5127
R16225 vdd.n1935 vdd.n873 99.5127
R16226 vdd.n1935 vdd.n867 99.5127
R16227 vdd.n1938 vdd.n867 99.5127
R16228 vdd.n1938 vdd.n860 99.5127
R16229 vdd.n1941 vdd.n860 99.5127
R16230 vdd.n1941 vdd.n853 99.5127
R16231 vdd.n1944 vdd.n853 99.5127
R16232 vdd.n1944 vdd.n848 99.5127
R16233 vdd.n1947 vdd.n848 99.5127
R16234 vdd.n1947 vdd.n842 99.5127
R16235 vdd.n1968 vdd.n842 99.5127
R16236 vdd.n1968 vdd.n835 99.5127
R16237 vdd.n1964 vdd.n835 99.5127
R16238 vdd.n1964 vdd.n829 99.5127
R16239 vdd.n1961 vdd.n829 99.5127
R16240 vdd.n1961 vdd.n824 99.5127
R16241 vdd.n1958 vdd.n824 99.5127
R16242 vdd.n1958 vdd.n819 99.5127
R16243 vdd.n1955 vdd.n819 99.5127
R16244 vdd.n1955 vdd.n813 99.5127
R16245 vdd.n1952 vdd.n813 99.5127
R16246 vdd.n1952 vdd.n806 99.5127
R16247 vdd.n806 vdd.n797 99.5127
R16248 vdd.n2170 vdd.n797 99.5127
R16249 vdd.n2171 vdd.n2170 99.5127
R16250 vdd.n2171 vdd.n789 99.5127
R16251 vdd.n2082 vdd.n2080 99.5127
R16252 vdd.n2078 vdd.n882 99.5127
R16253 vdd.n2074 vdd.n2072 99.5127
R16254 vdd.n2070 vdd.n884 99.5127
R16255 vdd.n2066 vdd.n2064 99.5127
R16256 vdd.n2062 vdd.n886 99.5127
R16257 vdd.n2058 vdd.n2056 99.5127
R16258 vdd.n2054 vdd.n888 99.5127
R16259 vdd.n1896 vdd.n890 99.5127
R16260 vdd.n1901 vdd.n1898 99.5127
R16261 vdd.n1905 vdd.n1903 99.5127
R16262 vdd.n1909 vdd.n1894 99.5127
R16263 vdd.n1913 vdd.n1911 99.5127
R16264 vdd.n1917 vdd.n1892 99.5127
R16265 vdd.n1921 vdd.n1919 99.5127
R16266 vdd.n1926 vdd.n1888 99.5127
R16267 vdd.n1929 vdd.n1928 99.5127
R16268 vdd.n2086 vdd.n870 99.5127
R16269 vdd.n2094 vdd.n870 99.5127
R16270 vdd.n2094 vdd.n868 99.5127
R16271 vdd.n2098 vdd.n868 99.5127
R16272 vdd.n2098 vdd.n857 99.5127
R16273 vdd.n2106 vdd.n857 99.5127
R16274 vdd.n2106 vdd.n854 99.5127
R16275 vdd.n2111 vdd.n854 99.5127
R16276 vdd.n2111 vdd.n845 99.5127
R16277 vdd.n2119 vdd.n845 99.5127
R16278 vdd.n2119 vdd.n843 99.5127
R16279 vdd.n2123 vdd.n843 99.5127
R16280 vdd.n2123 vdd.n833 99.5127
R16281 vdd.n2131 vdd.n833 99.5127
R16282 vdd.n2131 vdd.n831 99.5127
R16283 vdd.n2135 vdd.n831 99.5127
R16284 vdd.n2135 vdd.n822 99.5127
R16285 vdd.n2143 vdd.n822 99.5127
R16286 vdd.n2143 vdd.n820 99.5127
R16287 vdd.n2147 vdd.n820 99.5127
R16288 vdd.n2147 vdd.n810 99.5127
R16289 vdd.n2155 vdd.n810 99.5127
R16290 vdd.n2155 vdd.n807 99.5127
R16291 vdd.n2161 vdd.n807 99.5127
R16292 vdd.n2161 vdd.n808 99.5127
R16293 vdd.n808 vdd.n799 99.5127
R16294 vdd.n799 vdd.n790 99.5127
R16295 vdd.n2243 vdd.n790 99.5127
R16296 vdd.n9 vdd.n7 98.9633
R16297 vdd.n2 vdd.n0 98.9633
R16298 vdd.n9 vdd.n8 98.6055
R16299 vdd.n11 vdd.n10 98.6055
R16300 vdd.n13 vdd.n12 98.6055
R16301 vdd.n6 vdd.n5 98.6055
R16302 vdd.n4 vdd.n3 98.6055
R16303 vdd.n2 vdd.n1 98.6055
R16304 vdd.t223 vdd.n279 85.8723
R16305 vdd.t22 vdd.n228 85.8723
R16306 vdd.t153 vdd.n185 85.8723
R16307 vdd.t27 vdd.n134 85.8723
R16308 vdd.t230 vdd.n92 85.8723
R16309 vdd.t175 vdd.n41 85.8723
R16310 vdd.t43 vdd.n1474 85.8723
R16311 vdd.t202 vdd.n1525 85.8723
R16312 vdd.t195 vdd.n1380 85.8723
R16313 vdd.t47 vdd.n1431 85.8723
R16314 vdd.t176 vdd.n1287 85.8723
R16315 vdd.t214 vdd.n1338 85.8723
R16316 vdd.n2635 vdd.n2634 78.546
R16317 vdd.n2109 vdd.n855 78.546
R16318 vdd.n266 vdd.n265 75.1835
R16319 vdd.n264 vdd.n263 75.1835
R16320 vdd.n262 vdd.n261 75.1835
R16321 vdd.n260 vdd.n259 75.1835
R16322 vdd.n258 vdd.n257 75.1835
R16323 vdd.n172 vdd.n171 75.1835
R16324 vdd.n170 vdd.n169 75.1835
R16325 vdd.n168 vdd.n167 75.1835
R16326 vdd.n166 vdd.n165 75.1835
R16327 vdd.n164 vdd.n163 75.1835
R16328 vdd.n79 vdd.n78 75.1835
R16329 vdd.n77 vdd.n76 75.1835
R16330 vdd.n75 vdd.n74 75.1835
R16331 vdd.n73 vdd.n72 75.1835
R16332 vdd.n71 vdd.n70 75.1835
R16333 vdd.n1504 vdd.n1503 75.1835
R16334 vdd.n1506 vdd.n1505 75.1835
R16335 vdd.n1508 vdd.n1507 75.1835
R16336 vdd.n1510 vdd.n1509 75.1835
R16337 vdd.n1512 vdd.n1511 75.1835
R16338 vdd.n1410 vdd.n1409 75.1835
R16339 vdd.n1412 vdd.n1411 75.1835
R16340 vdd.n1414 vdd.n1413 75.1835
R16341 vdd.n1416 vdd.n1415 75.1835
R16342 vdd.n1418 vdd.n1417 75.1835
R16343 vdd.n1317 vdd.n1316 75.1835
R16344 vdd.n1319 vdd.n1318 75.1835
R16345 vdd.n1321 vdd.n1320 75.1835
R16346 vdd.n1323 vdd.n1322 75.1835
R16347 vdd.n1325 vdd.n1324 75.1835
R16348 vdd.n2570 vdd.n2569 72.8958
R16349 vdd.n2569 vdd.n2333 72.8958
R16350 vdd.n2569 vdd.n2334 72.8958
R16351 vdd.n2569 vdd.n2335 72.8958
R16352 vdd.n2569 vdd.n2336 72.8958
R16353 vdd.n2569 vdd.n2337 72.8958
R16354 vdd.n2569 vdd.n2338 72.8958
R16355 vdd.n2569 vdd.n2339 72.8958
R16356 vdd.n2569 vdd.n2340 72.8958
R16357 vdd.n2569 vdd.n2341 72.8958
R16358 vdd.n2569 vdd.n2342 72.8958
R16359 vdd.n2569 vdd.n2343 72.8958
R16360 vdd.n2569 vdd.n2344 72.8958
R16361 vdd.n2569 vdd.n2345 72.8958
R16362 vdd.n2569 vdd.n2346 72.8958
R16363 vdd.n2569 vdd.n2347 72.8958
R16364 vdd.n2569 vdd.n2348 72.8958
R16365 vdd.n629 vdd.n613 72.8958
R16366 vdd.n2778 vdd.n613 72.8958
R16367 vdd.n623 vdd.n613 72.8958
R16368 vdd.n2785 vdd.n613 72.8958
R16369 vdd.n620 vdd.n613 72.8958
R16370 vdd.n2792 vdd.n613 72.8958
R16371 vdd.n617 vdd.n613 72.8958
R16372 vdd.n2799 vdd.n613 72.8958
R16373 vdd.n2802 vdd.n613 72.8958
R16374 vdd.n2658 vdd.n613 72.8958
R16375 vdd.n2663 vdd.n613 72.8958
R16376 vdd.n2657 vdd.n613 72.8958
R16377 vdd.n2670 vdd.n613 72.8958
R16378 vdd.n2654 vdd.n613 72.8958
R16379 vdd.n2677 vdd.n613 72.8958
R16380 vdd.n2651 vdd.n613 72.8958
R16381 vdd.n2684 vdd.n613 72.8958
R16382 vdd.n1822 vdd.n877 72.8958
R16383 vdd.n1828 vdd.n877 72.8958
R16384 vdd.n1830 vdd.n877 72.8958
R16385 vdd.n1836 vdd.n877 72.8958
R16386 vdd.n1838 vdd.n877 72.8958
R16387 vdd.n1844 vdd.n877 72.8958
R16388 vdd.n1846 vdd.n877 72.8958
R16389 vdd.n1852 vdd.n877 72.8958
R16390 vdd.n2023 vdd.n877 72.8958
R16391 vdd.n2021 vdd.n877 72.8958
R16392 vdd.n2015 vdd.n877 72.8958
R16393 vdd.n2013 vdd.n877 72.8958
R16394 vdd.n2007 vdd.n877 72.8958
R16395 vdd.n2005 vdd.n877 72.8958
R16396 vdd.n1999 vdd.n877 72.8958
R16397 vdd.n1997 vdd.n877 72.8958
R16398 vdd.n1991 vdd.n877 72.8958
R16399 vdd.n2316 vdd.n765 72.8958
R16400 vdd.n2316 vdd.n766 72.8958
R16401 vdd.n2316 vdd.n767 72.8958
R16402 vdd.n2316 vdd.n768 72.8958
R16403 vdd.n2316 vdd.n769 72.8958
R16404 vdd.n2316 vdd.n770 72.8958
R16405 vdd.n2316 vdd.n771 72.8958
R16406 vdd.n2316 vdd.n772 72.8958
R16407 vdd.n2316 vdd.n773 72.8958
R16408 vdd.n2316 vdd.n774 72.8958
R16409 vdd.n2316 vdd.n775 72.8958
R16410 vdd.n2316 vdd.n776 72.8958
R16411 vdd.n2316 vdd.n777 72.8958
R16412 vdd.n2316 vdd.n778 72.8958
R16413 vdd.n2316 vdd.n779 72.8958
R16414 vdd.n2316 vdd.n780 72.8958
R16415 vdd.n2316 vdd.n781 72.8958
R16416 vdd.n2569 vdd.n2568 72.8958
R16417 vdd.n2569 vdd.n2317 72.8958
R16418 vdd.n2569 vdd.n2318 72.8958
R16419 vdd.n2569 vdd.n2319 72.8958
R16420 vdd.n2569 vdd.n2320 72.8958
R16421 vdd.n2569 vdd.n2321 72.8958
R16422 vdd.n2569 vdd.n2322 72.8958
R16423 vdd.n2569 vdd.n2323 72.8958
R16424 vdd.n2569 vdd.n2324 72.8958
R16425 vdd.n2569 vdd.n2325 72.8958
R16426 vdd.n2569 vdd.n2326 72.8958
R16427 vdd.n2569 vdd.n2327 72.8958
R16428 vdd.n2569 vdd.n2328 72.8958
R16429 vdd.n2569 vdd.n2329 72.8958
R16430 vdd.n2569 vdd.n2330 72.8958
R16431 vdd.n2569 vdd.n2331 72.8958
R16432 vdd.n2569 vdd.n2332 72.8958
R16433 vdd.n2706 vdd.n613 72.8958
R16434 vdd.n2712 vdd.n613 72.8958
R16435 vdd.n659 vdd.n613 72.8958
R16436 vdd.n2719 vdd.n613 72.8958
R16437 vdd.n656 vdd.n613 72.8958
R16438 vdd.n2726 vdd.n613 72.8958
R16439 vdd.n653 vdd.n613 72.8958
R16440 vdd.n2733 vdd.n613 72.8958
R16441 vdd.n650 vdd.n613 72.8958
R16442 vdd.n2741 vdd.n613 72.8958
R16443 vdd.n647 vdd.n613 72.8958
R16444 vdd.n2748 vdd.n613 72.8958
R16445 vdd.n644 vdd.n613 72.8958
R16446 vdd.n2755 vdd.n613 72.8958
R16447 vdd.n641 vdd.n613 72.8958
R16448 vdd.n2762 vdd.n613 72.8958
R16449 vdd.n2765 vdd.n613 72.8958
R16450 vdd.n2316 vdd.n763 72.8958
R16451 vdd.n2316 vdd.n762 72.8958
R16452 vdd.n2316 vdd.n761 72.8958
R16453 vdd.n2316 vdd.n760 72.8958
R16454 vdd.n2316 vdd.n759 72.8958
R16455 vdd.n2316 vdd.n758 72.8958
R16456 vdd.n2316 vdd.n757 72.8958
R16457 vdd.n2316 vdd.n756 72.8958
R16458 vdd.n2316 vdd.n755 72.8958
R16459 vdd.n2316 vdd.n754 72.8958
R16460 vdd.n2316 vdd.n753 72.8958
R16461 vdd.n2316 vdd.n752 72.8958
R16462 vdd.n2316 vdd.n751 72.8958
R16463 vdd.n2316 vdd.n750 72.8958
R16464 vdd.n2316 vdd.n749 72.8958
R16465 vdd.n2316 vdd.n748 72.8958
R16466 vdd.n2316 vdd.n747 72.8958
R16467 vdd.n2081 vdd.n877 72.8958
R16468 vdd.n2079 vdd.n877 72.8958
R16469 vdd.n2073 vdd.n877 72.8958
R16470 vdd.n2071 vdd.n877 72.8958
R16471 vdd.n2065 vdd.n877 72.8958
R16472 vdd.n2063 vdd.n877 72.8958
R16473 vdd.n2057 vdd.n877 72.8958
R16474 vdd.n2055 vdd.n877 72.8958
R16475 vdd.n889 vdd.n877 72.8958
R16476 vdd.n1897 vdd.n877 72.8958
R16477 vdd.n1902 vdd.n877 72.8958
R16478 vdd.n1904 vdd.n877 72.8958
R16479 vdd.n1910 vdd.n877 72.8958
R16480 vdd.n1912 vdd.n877 72.8958
R16481 vdd.n1918 vdd.n877 72.8958
R16482 vdd.n1920 vdd.n877 72.8958
R16483 vdd.n1927 vdd.n877 72.8958
R16484 vdd.n986 vdd.n982 66.2847
R16485 vdd.n992 vdd.n982 66.2847
R16486 vdd.n995 vdd.n982 66.2847
R16487 vdd.n1000 vdd.n982 66.2847
R16488 vdd.n1003 vdd.n982 66.2847
R16489 vdd.n1008 vdd.n982 66.2847
R16490 vdd.n1011 vdd.n982 66.2847
R16491 vdd.n1016 vdd.n982 66.2847
R16492 vdd.n1019 vdd.n982 66.2847
R16493 vdd.n1026 vdd.n982 66.2847
R16494 vdd.n1029 vdd.n982 66.2847
R16495 vdd.n1034 vdd.n982 66.2847
R16496 vdd.n1037 vdd.n982 66.2847
R16497 vdd.n1042 vdd.n982 66.2847
R16498 vdd.n1045 vdd.n982 66.2847
R16499 vdd.n1050 vdd.n982 66.2847
R16500 vdd.n1053 vdd.n982 66.2847
R16501 vdd.n1058 vdd.n982 66.2847
R16502 vdd.n1061 vdd.n982 66.2847
R16503 vdd.n1066 vdd.n982 66.2847
R16504 vdd.n1145 vdd.n982 66.2847
R16505 vdd.n1069 vdd.n982 66.2847
R16506 vdd.n1075 vdd.n982 66.2847
R16507 vdd.n1080 vdd.n982 66.2847
R16508 vdd.n1083 vdd.n982 66.2847
R16509 vdd.n1088 vdd.n982 66.2847
R16510 vdd.n1091 vdd.n982 66.2847
R16511 vdd.n1096 vdd.n982 66.2847
R16512 vdd.n1099 vdd.n982 66.2847
R16513 vdd.n1104 vdd.n982 66.2847
R16514 vdd.n1107 vdd.n982 66.2847
R16515 vdd.n901 vdd.n898 66.2847
R16516 vdd.n1712 vdd.n901 66.2847
R16517 vdd.n1717 vdd.n901 66.2847
R16518 vdd.n1722 vdd.n901 66.2847
R16519 vdd.n1710 vdd.n901 66.2847
R16520 vdd.n1729 vdd.n901 66.2847
R16521 vdd.n1702 vdd.n901 66.2847
R16522 vdd.n1736 vdd.n901 66.2847
R16523 vdd.n1695 vdd.n901 66.2847
R16524 vdd.n1743 vdd.n901 66.2847
R16525 vdd.n1689 vdd.n901 66.2847
R16526 vdd.n1684 vdd.n901 66.2847
R16527 vdd.n1754 vdd.n901 66.2847
R16528 vdd.n1676 vdd.n901 66.2847
R16529 vdd.n1761 vdd.n901 66.2847
R16530 vdd.n1669 vdd.n901 66.2847
R16531 vdd.n1768 vdd.n901 66.2847
R16532 vdd.n1662 vdd.n901 66.2847
R16533 vdd.n1775 vdd.n901 66.2847
R16534 vdd.n1655 vdd.n901 66.2847
R16535 vdd.n1782 vdd.n901 66.2847
R16536 vdd.n1649 vdd.n901 66.2847
R16537 vdd.n1644 vdd.n901 66.2847
R16538 vdd.n1793 vdd.n901 66.2847
R16539 vdd.n1636 vdd.n901 66.2847
R16540 vdd.n1800 vdd.n901 66.2847
R16541 vdd.n1629 vdd.n901 66.2847
R16542 vdd.n1807 vdd.n901 66.2847
R16543 vdd.n1810 vdd.n901 66.2847
R16544 vdd.n1620 vdd.n901 66.2847
R16545 vdd.n2032 vdd.n901 66.2847
R16546 vdd.n1614 vdd.n901 66.2847
R16547 vdd.n2932 vdd.n516 66.2847
R16548 vdd.n520 vdd.n516 66.2847
R16549 vdd.n523 vdd.n516 66.2847
R16550 vdd.n2921 vdd.n516 66.2847
R16551 vdd.n2915 vdd.n516 66.2847
R16552 vdd.n2913 vdd.n516 66.2847
R16553 vdd.n2907 vdd.n516 66.2847
R16554 vdd.n2905 vdd.n516 66.2847
R16555 vdd.n2899 vdd.n516 66.2847
R16556 vdd.n2897 vdd.n516 66.2847
R16557 vdd.n2891 vdd.n516 66.2847
R16558 vdd.n2889 vdd.n516 66.2847
R16559 vdd.n2883 vdd.n516 66.2847
R16560 vdd.n2881 vdd.n516 66.2847
R16561 vdd.n2875 vdd.n516 66.2847
R16562 vdd.n2873 vdd.n516 66.2847
R16563 vdd.n2867 vdd.n516 66.2847
R16564 vdd.n2865 vdd.n516 66.2847
R16565 vdd.n2859 vdd.n516 66.2847
R16566 vdd.n2857 vdd.n516 66.2847
R16567 vdd.n584 vdd.n516 66.2847
R16568 vdd.n2848 vdd.n516 66.2847
R16569 vdd.n586 vdd.n516 66.2847
R16570 vdd.n2841 vdd.n516 66.2847
R16571 vdd.n2835 vdd.n516 66.2847
R16572 vdd.n2833 vdd.n516 66.2847
R16573 vdd.n2827 vdd.n516 66.2847
R16574 vdd.n2825 vdd.n516 66.2847
R16575 vdd.n2819 vdd.n516 66.2847
R16576 vdd.n607 vdd.n516 66.2847
R16577 vdd.n609 vdd.n516 66.2847
R16578 vdd.n3018 vdd.n351 66.2847
R16579 vdd.n3027 vdd.n351 66.2847
R16580 vdd.n461 vdd.n351 66.2847
R16581 vdd.n3034 vdd.n351 66.2847
R16582 vdd.n454 vdd.n351 66.2847
R16583 vdd.n3041 vdd.n351 66.2847
R16584 vdd.n447 vdd.n351 66.2847
R16585 vdd.n3048 vdd.n351 66.2847
R16586 vdd.n440 vdd.n351 66.2847
R16587 vdd.n3055 vdd.n351 66.2847
R16588 vdd.n434 vdd.n351 66.2847
R16589 vdd.n429 vdd.n351 66.2847
R16590 vdd.n3066 vdd.n351 66.2847
R16591 vdd.n421 vdd.n351 66.2847
R16592 vdd.n3073 vdd.n351 66.2847
R16593 vdd.n414 vdd.n351 66.2847
R16594 vdd.n3080 vdd.n351 66.2847
R16595 vdd.n407 vdd.n351 66.2847
R16596 vdd.n3087 vdd.n351 66.2847
R16597 vdd.n400 vdd.n351 66.2847
R16598 vdd.n3094 vdd.n351 66.2847
R16599 vdd.n394 vdd.n351 66.2847
R16600 vdd.n389 vdd.n351 66.2847
R16601 vdd.n3105 vdd.n351 66.2847
R16602 vdd.n381 vdd.n351 66.2847
R16603 vdd.n3112 vdd.n351 66.2847
R16604 vdd.n374 vdd.n351 66.2847
R16605 vdd.n3119 vdd.n351 66.2847
R16606 vdd.n367 vdd.n351 66.2847
R16607 vdd.n3126 vdd.n351 66.2847
R16608 vdd.n3129 vdd.n351 66.2847
R16609 vdd.n355 vdd.n351 66.2847
R16610 vdd.n356 vdd.n355 52.4337
R16611 vdd.n3129 vdd.n3128 52.4337
R16612 vdd.n3126 vdd.n3125 52.4337
R16613 vdd.n3121 vdd.n367 52.4337
R16614 vdd.n3119 vdd.n3118 52.4337
R16615 vdd.n3114 vdd.n374 52.4337
R16616 vdd.n3112 vdd.n3111 52.4337
R16617 vdd.n3107 vdd.n381 52.4337
R16618 vdd.n3105 vdd.n3104 52.4337
R16619 vdd.n390 vdd.n389 52.4337
R16620 vdd.n3096 vdd.n394 52.4337
R16621 vdd.n3094 vdd.n3093 52.4337
R16622 vdd.n3089 vdd.n400 52.4337
R16623 vdd.n3087 vdd.n3086 52.4337
R16624 vdd.n3082 vdd.n407 52.4337
R16625 vdd.n3080 vdd.n3079 52.4337
R16626 vdd.n3075 vdd.n414 52.4337
R16627 vdd.n3073 vdd.n3072 52.4337
R16628 vdd.n3068 vdd.n421 52.4337
R16629 vdd.n3066 vdd.n3065 52.4337
R16630 vdd.n430 vdd.n429 52.4337
R16631 vdd.n3057 vdd.n434 52.4337
R16632 vdd.n3055 vdd.n3054 52.4337
R16633 vdd.n3050 vdd.n440 52.4337
R16634 vdd.n3048 vdd.n3047 52.4337
R16635 vdd.n3043 vdd.n447 52.4337
R16636 vdd.n3041 vdd.n3040 52.4337
R16637 vdd.n3036 vdd.n454 52.4337
R16638 vdd.n3034 vdd.n3033 52.4337
R16639 vdd.n3029 vdd.n461 52.4337
R16640 vdd.n3027 vdd.n3026 52.4337
R16641 vdd.n3019 vdd.n3018 52.4337
R16642 vdd.n2932 vdd.n517 52.4337
R16643 vdd.n2930 vdd.n520 52.4337
R16644 vdd.n2926 vdd.n523 52.4337
R16645 vdd.n2922 vdd.n2921 52.4337
R16646 vdd.n2915 vdd.n526 52.4337
R16647 vdd.n2914 vdd.n2913 52.4337
R16648 vdd.n2907 vdd.n532 52.4337
R16649 vdd.n2906 vdd.n2905 52.4337
R16650 vdd.n2899 vdd.n538 52.4337
R16651 vdd.n2898 vdd.n2897 52.4337
R16652 vdd.n2891 vdd.n546 52.4337
R16653 vdd.n2890 vdd.n2889 52.4337
R16654 vdd.n2883 vdd.n552 52.4337
R16655 vdd.n2882 vdd.n2881 52.4337
R16656 vdd.n2875 vdd.n558 52.4337
R16657 vdd.n2874 vdd.n2873 52.4337
R16658 vdd.n2867 vdd.n564 52.4337
R16659 vdd.n2866 vdd.n2865 52.4337
R16660 vdd.n2859 vdd.n570 52.4337
R16661 vdd.n2858 vdd.n2857 52.4337
R16662 vdd.n584 vdd.n576 52.4337
R16663 vdd.n2849 vdd.n2848 52.4337
R16664 vdd.n2846 vdd.n586 52.4337
R16665 vdd.n2842 vdd.n2841 52.4337
R16666 vdd.n2835 vdd.n590 52.4337
R16667 vdd.n2834 vdd.n2833 52.4337
R16668 vdd.n2827 vdd.n596 52.4337
R16669 vdd.n2826 vdd.n2825 52.4337
R16670 vdd.n2819 vdd.n602 52.4337
R16671 vdd.n2818 vdd.n607 52.4337
R16672 vdd.n2814 vdd.n609 52.4337
R16673 vdd.n2034 vdd.n1614 52.4337
R16674 vdd.n2032 vdd.n2031 52.4337
R16675 vdd.n1621 vdd.n1620 52.4337
R16676 vdd.n1810 vdd.n1809 52.4337
R16677 vdd.n1807 vdd.n1806 52.4337
R16678 vdd.n1802 vdd.n1629 52.4337
R16679 vdd.n1800 vdd.n1799 52.4337
R16680 vdd.n1795 vdd.n1636 52.4337
R16681 vdd.n1793 vdd.n1792 52.4337
R16682 vdd.n1645 vdd.n1644 52.4337
R16683 vdd.n1784 vdd.n1649 52.4337
R16684 vdd.n1782 vdd.n1781 52.4337
R16685 vdd.n1777 vdd.n1655 52.4337
R16686 vdd.n1775 vdd.n1774 52.4337
R16687 vdd.n1770 vdd.n1662 52.4337
R16688 vdd.n1768 vdd.n1767 52.4337
R16689 vdd.n1763 vdd.n1669 52.4337
R16690 vdd.n1761 vdd.n1760 52.4337
R16691 vdd.n1756 vdd.n1676 52.4337
R16692 vdd.n1754 vdd.n1753 52.4337
R16693 vdd.n1685 vdd.n1684 52.4337
R16694 vdd.n1745 vdd.n1689 52.4337
R16695 vdd.n1743 vdd.n1742 52.4337
R16696 vdd.n1738 vdd.n1695 52.4337
R16697 vdd.n1736 vdd.n1735 52.4337
R16698 vdd.n1731 vdd.n1702 52.4337
R16699 vdd.n1729 vdd.n1728 52.4337
R16700 vdd.n1724 vdd.n1710 52.4337
R16701 vdd.n1722 vdd.n1721 52.4337
R16702 vdd.n1717 vdd.n1716 52.4337
R16703 vdd.n1712 vdd.n1711 52.4337
R16704 vdd.n2043 vdd.n898 52.4337
R16705 vdd.n986 vdd.n984 52.4337
R16706 vdd.n992 vdd.n991 52.4337
R16707 vdd.n995 vdd.n994 52.4337
R16708 vdd.n1000 vdd.n999 52.4337
R16709 vdd.n1003 vdd.n1002 52.4337
R16710 vdd.n1008 vdd.n1007 52.4337
R16711 vdd.n1011 vdd.n1010 52.4337
R16712 vdd.n1016 vdd.n1015 52.4337
R16713 vdd.n1019 vdd.n1018 52.4337
R16714 vdd.n1026 vdd.n1025 52.4337
R16715 vdd.n1029 vdd.n1028 52.4337
R16716 vdd.n1034 vdd.n1033 52.4337
R16717 vdd.n1037 vdd.n1036 52.4337
R16718 vdd.n1042 vdd.n1041 52.4337
R16719 vdd.n1045 vdd.n1044 52.4337
R16720 vdd.n1050 vdd.n1049 52.4337
R16721 vdd.n1053 vdd.n1052 52.4337
R16722 vdd.n1058 vdd.n1057 52.4337
R16723 vdd.n1061 vdd.n1060 52.4337
R16724 vdd.n1066 vdd.n1065 52.4337
R16725 vdd.n1146 vdd.n1145 52.4337
R16726 vdd.n1143 vdd.n1069 52.4337
R16727 vdd.n1075 vdd.n1074 52.4337
R16728 vdd.n1080 vdd.n1077 52.4337
R16729 vdd.n1083 vdd.n1082 52.4337
R16730 vdd.n1088 vdd.n1085 52.4337
R16731 vdd.n1091 vdd.n1090 52.4337
R16732 vdd.n1096 vdd.n1093 52.4337
R16733 vdd.n1099 vdd.n1098 52.4337
R16734 vdd.n1104 vdd.n1101 52.4337
R16735 vdd.n1107 vdd.n1106 52.4337
R16736 vdd.n987 vdd.n986 52.4337
R16737 vdd.n993 vdd.n992 52.4337
R16738 vdd.n996 vdd.n995 52.4337
R16739 vdd.n1001 vdd.n1000 52.4337
R16740 vdd.n1004 vdd.n1003 52.4337
R16741 vdd.n1009 vdd.n1008 52.4337
R16742 vdd.n1012 vdd.n1011 52.4337
R16743 vdd.n1017 vdd.n1016 52.4337
R16744 vdd.n1020 vdd.n1019 52.4337
R16745 vdd.n1027 vdd.n1026 52.4337
R16746 vdd.n1030 vdd.n1029 52.4337
R16747 vdd.n1035 vdd.n1034 52.4337
R16748 vdd.n1038 vdd.n1037 52.4337
R16749 vdd.n1043 vdd.n1042 52.4337
R16750 vdd.n1046 vdd.n1045 52.4337
R16751 vdd.n1051 vdd.n1050 52.4337
R16752 vdd.n1054 vdd.n1053 52.4337
R16753 vdd.n1059 vdd.n1058 52.4337
R16754 vdd.n1062 vdd.n1061 52.4337
R16755 vdd.n1067 vdd.n1066 52.4337
R16756 vdd.n1145 vdd.n1144 52.4337
R16757 vdd.n1073 vdd.n1069 52.4337
R16758 vdd.n1076 vdd.n1075 52.4337
R16759 vdd.n1081 vdd.n1080 52.4337
R16760 vdd.n1084 vdd.n1083 52.4337
R16761 vdd.n1089 vdd.n1088 52.4337
R16762 vdd.n1092 vdd.n1091 52.4337
R16763 vdd.n1097 vdd.n1096 52.4337
R16764 vdd.n1100 vdd.n1099 52.4337
R16765 vdd.n1105 vdd.n1104 52.4337
R16766 vdd.n1108 vdd.n1107 52.4337
R16767 vdd.n898 vdd.n897 52.4337
R16768 vdd.n1713 vdd.n1712 52.4337
R16769 vdd.n1718 vdd.n1717 52.4337
R16770 vdd.n1723 vdd.n1722 52.4337
R16771 vdd.n1710 vdd.n1703 52.4337
R16772 vdd.n1730 vdd.n1729 52.4337
R16773 vdd.n1702 vdd.n1696 52.4337
R16774 vdd.n1737 vdd.n1736 52.4337
R16775 vdd.n1695 vdd.n1690 52.4337
R16776 vdd.n1744 vdd.n1743 52.4337
R16777 vdd.n1689 vdd.n1688 52.4337
R16778 vdd.n1684 vdd.n1677 52.4337
R16779 vdd.n1755 vdd.n1754 52.4337
R16780 vdd.n1676 vdd.n1670 52.4337
R16781 vdd.n1762 vdd.n1761 52.4337
R16782 vdd.n1669 vdd.n1663 52.4337
R16783 vdd.n1769 vdd.n1768 52.4337
R16784 vdd.n1662 vdd.n1656 52.4337
R16785 vdd.n1776 vdd.n1775 52.4337
R16786 vdd.n1655 vdd.n1650 52.4337
R16787 vdd.n1783 vdd.n1782 52.4337
R16788 vdd.n1649 vdd.n1648 52.4337
R16789 vdd.n1644 vdd.n1637 52.4337
R16790 vdd.n1794 vdd.n1793 52.4337
R16791 vdd.n1636 vdd.n1630 52.4337
R16792 vdd.n1801 vdd.n1800 52.4337
R16793 vdd.n1629 vdd.n1623 52.4337
R16794 vdd.n1808 vdd.n1807 52.4337
R16795 vdd.n1811 vdd.n1810 52.4337
R16796 vdd.n1620 vdd.n1615 52.4337
R16797 vdd.n2033 vdd.n2032 52.4337
R16798 vdd.n1614 vdd.n903 52.4337
R16799 vdd.n2933 vdd.n2932 52.4337
R16800 vdd.n2927 vdd.n520 52.4337
R16801 vdd.n2923 vdd.n523 52.4337
R16802 vdd.n2921 vdd.n2920 52.4337
R16803 vdd.n2916 vdd.n2915 52.4337
R16804 vdd.n2913 vdd.n2912 52.4337
R16805 vdd.n2908 vdd.n2907 52.4337
R16806 vdd.n2905 vdd.n2904 52.4337
R16807 vdd.n2900 vdd.n2899 52.4337
R16808 vdd.n2897 vdd.n2896 52.4337
R16809 vdd.n2892 vdd.n2891 52.4337
R16810 vdd.n2889 vdd.n2888 52.4337
R16811 vdd.n2884 vdd.n2883 52.4337
R16812 vdd.n2881 vdd.n2880 52.4337
R16813 vdd.n2876 vdd.n2875 52.4337
R16814 vdd.n2873 vdd.n2872 52.4337
R16815 vdd.n2868 vdd.n2867 52.4337
R16816 vdd.n2865 vdd.n2864 52.4337
R16817 vdd.n2860 vdd.n2859 52.4337
R16818 vdd.n2857 vdd.n2856 52.4337
R16819 vdd.n585 vdd.n584 52.4337
R16820 vdd.n2848 vdd.n2847 52.4337
R16821 vdd.n2843 vdd.n586 52.4337
R16822 vdd.n2841 vdd.n2840 52.4337
R16823 vdd.n2836 vdd.n2835 52.4337
R16824 vdd.n2833 vdd.n2832 52.4337
R16825 vdd.n2828 vdd.n2827 52.4337
R16826 vdd.n2825 vdd.n2824 52.4337
R16827 vdd.n2820 vdd.n2819 52.4337
R16828 vdd.n2815 vdd.n607 52.4337
R16829 vdd.n2811 vdd.n609 52.4337
R16830 vdd.n3018 vdd.n462 52.4337
R16831 vdd.n3028 vdd.n3027 52.4337
R16832 vdd.n461 vdd.n455 52.4337
R16833 vdd.n3035 vdd.n3034 52.4337
R16834 vdd.n454 vdd.n448 52.4337
R16835 vdd.n3042 vdd.n3041 52.4337
R16836 vdd.n447 vdd.n441 52.4337
R16837 vdd.n3049 vdd.n3048 52.4337
R16838 vdd.n440 vdd.n435 52.4337
R16839 vdd.n3056 vdd.n3055 52.4337
R16840 vdd.n434 vdd.n433 52.4337
R16841 vdd.n429 vdd.n422 52.4337
R16842 vdd.n3067 vdd.n3066 52.4337
R16843 vdd.n421 vdd.n415 52.4337
R16844 vdd.n3074 vdd.n3073 52.4337
R16845 vdd.n414 vdd.n408 52.4337
R16846 vdd.n3081 vdd.n3080 52.4337
R16847 vdd.n407 vdd.n401 52.4337
R16848 vdd.n3088 vdd.n3087 52.4337
R16849 vdd.n400 vdd.n395 52.4337
R16850 vdd.n3095 vdd.n3094 52.4337
R16851 vdd.n394 vdd.n393 52.4337
R16852 vdd.n389 vdd.n382 52.4337
R16853 vdd.n3106 vdd.n3105 52.4337
R16854 vdd.n381 vdd.n375 52.4337
R16855 vdd.n3113 vdd.n3112 52.4337
R16856 vdd.n374 vdd.n368 52.4337
R16857 vdd.n3120 vdd.n3119 52.4337
R16858 vdd.n367 vdd.n360 52.4337
R16859 vdd.n3127 vdd.n3126 52.4337
R16860 vdd.n3130 vdd.n3129 52.4337
R16861 vdd.n355 vdd.n352 52.4337
R16862 vdd.t200 vdd.t17 51.4683
R16863 vdd.n258 vdd.n256 42.0461
R16864 vdd.n164 vdd.n162 42.0461
R16865 vdd.n71 vdd.n69 42.0461
R16866 vdd.n1504 vdd.n1502 42.0461
R16867 vdd.n1410 vdd.n1408 42.0461
R16868 vdd.n1317 vdd.n1315 42.0461
R16869 vdd.n308 vdd.n307 41.6884
R16870 vdd.n214 vdd.n213 41.6884
R16871 vdd.n121 vdd.n120 41.6884
R16872 vdd.n1554 vdd.n1553 41.6884
R16873 vdd.n1460 vdd.n1459 41.6884
R16874 vdd.n1367 vdd.n1366 41.6884
R16875 vdd.n1112 vdd.n1111 41.1157
R16876 vdd.n1149 vdd.n1148 41.1157
R16877 vdd.n1023 vdd.n1022 41.1157
R16878 vdd.n3023 vdd.n3022 41.1157
R16879 vdd.n3062 vdd.n428 41.1157
R16880 vdd.n3101 vdd.n388 41.1157
R16881 vdd.n2765 vdd.n2764 39.2114
R16882 vdd.n2762 vdd.n2761 39.2114
R16883 vdd.n2757 vdd.n641 39.2114
R16884 vdd.n2755 vdd.n2754 39.2114
R16885 vdd.n2750 vdd.n644 39.2114
R16886 vdd.n2748 vdd.n2747 39.2114
R16887 vdd.n2743 vdd.n647 39.2114
R16888 vdd.n2741 vdd.n2740 39.2114
R16889 vdd.n2735 vdd.n650 39.2114
R16890 vdd.n2733 vdd.n2732 39.2114
R16891 vdd.n2728 vdd.n653 39.2114
R16892 vdd.n2726 vdd.n2725 39.2114
R16893 vdd.n2721 vdd.n656 39.2114
R16894 vdd.n2719 vdd.n2718 39.2114
R16895 vdd.n2714 vdd.n659 39.2114
R16896 vdd.n2712 vdd.n2711 39.2114
R16897 vdd.n2707 vdd.n2706 39.2114
R16898 vdd.n2568 vdd.n741 39.2114
R16899 vdd.n2563 vdd.n2317 39.2114
R16900 vdd.n2560 vdd.n2318 39.2114
R16901 vdd.n2556 vdd.n2319 39.2114
R16902 vdd.n2552 vdd.n2320 39.2114
R16903 vdd.n2548 vdd.n2321 39.2114
R16904 vdd.n2544 vdd.n2322 39.2114
R16905 vdd.n2540 vdd.n2323 39.2114
R16906 vdd.n2536 vdd.n2324 39.2114
R16907 vdd.n2532 vdd.n2325 39.2114
R16908 vdd.n2528 vdd.n2326 39.2114
R16909 vdd.n2524 vdd.n2327 39.2114
R16910 vdd.n2520 vdd.n2328 39.2114
R16911 vdd.n2516 vdd.n2329 39.2114
R16912 vdd.n2512 vdd.n2330 39.2114
R16913 vdd.n2508 vdd.n2331 39.2114
R16914 vdd.n2503 vdd.n2332 39.2114
R16915 vdd.n2311 vdd.n781 39.2114
R16916 vdd.n2307 vdd.n780 39.2114
R16917 vdd.n2303 vdd.n779 39.2114
R16918 vdd.n2299 vdd.n778 39.2114
R16919 vdd.n2295 vdd.n777 39.2114
R16920 vdd.n2291 vdd.n776 39.2114
R16921 vdd.n2287 vdd.n775 39.2114
R16922 vdd.n2283 vdd.n774 39.2114
R16923 vdd.n2279 vdd.n773 39.2114
R16924 vdd.n2275 vdd.n772 39.2114
R16925 vdd.n2271 vdd.n771 39.2114
R16926 vdd.n2267 vdd.n770 39.2114
R16927 vdd.n2263 vdd.n769 39.2114
R16928 vdd.n2259 vdd.n768 39.2114
R16929 vdd.n2255 vdd.n767 39.2114
R16930 vdd.n2250 vdd.n766 39.2114
R16931 vdd.n2246 vdd.n765 39.2114
R16932 vdd.n1822 vdd.n876 39.2114
R16933 vdd.n1828 vdd.n1827 39.2114
R16934 vdd.n1831 vdd.n1830 39.2114
R16935 vdd.n1836 vdd.n1835 39.2114
R16936 vdd.n1839 vdd.n1838 39.2114
R16937 vdd.n1844 vdd.n1843 39.2114
R16938 vdd.n1847 vdd.n1846 39.2114
R16939 vdd.n1852 vdd.n1851 39.2114
R16940 vdd.n2023 vdd.n1854 39.2114
R16941 vdd.n2022 vdd.n2021 39.2114
R16942 vdd.n2015 vdd.n1856 39.2114
R16943 vdd.n2014 vdd.n2013 39.2114
R16944 vdd.n2007 vdd.n1858 39.2114
R16945 vdd.n2006 vdd.n2005 39.2114
R16946 vdd.n1999 vdd.n1860 39.2114
R16947 vdd.n1998 vdd.n1997 39.2114
R16948 vdd.n1991 vdd.n1862 39.2114
R16949 vdd.n2684 vdd.n2683 39.2114
R16950 vdd.n2679 vdd.n2651 39.2114
R16951 vdd.n2677 vdd.n2676 39.2114
R16952 vdd.n2672 vdd.n2654 39.2114
R16953 vdd.n2670 vdd.n2669 39.2114
R16954 vdd.n2665 vdd.n2657 39.2114
R16955 vdd.n2663 vdd.n2662 39.2114
R16956 vdd.n2658 vdd.n612 39.2114
R16957 vdd.n2802 vdd.n2801 39.2114
R16958 vdd.n2799 vdd.n2798 39.2114
R16959 vdd.n2794 vdd.n617 39.2114
R16960 vdd.n2792 vdd.n2791 39.2114
R16961 vdd.n2787 vdd.n620 39.2114
R16962 vdd.n2785 vdd.n2784 39.2114
R16963 vdd.n2780 vdd.n623 39.2114
R16964 vdd.n2778 vdd.n2777 39.2114
R16965 vdd.n2773 vdd.n629 39.2114
R16966 vdd.n2570 vdd.n744 39.2114
R16967 vdd.n2333 vdd.n746 39.2114
R16968 vdd.n2359 vdd.n2334 39.2114
R16969 vdd.n2363 vdd.n2335 39.2114
R16970 vdd.n2367 vdd.n2336 39.2114
R16971 vdd.n2371 vdd.n2337 39.2114
R16972 vdd.n2375 vdd.n2338 39.2114
R16973 vdd.n2379 vdd.n2339 39.2114
R16974 vdd.n2383 vdd.n2340 39.2114
R16975 vdd.n2387 vdd.n2341 39.2114
R16976 vdd.n2391 vdd.n2342 39.2114
R16977 vdd.n2395 vdd.n2343 39.2114
R16978 vdd.n2399 vdd.n2344 39.2114
R16979 vdd.n2403 vdd.n2345 39.2114
R16980 vdd.n2407 vdd.n2346 39.2114
R16981 vdd.n2411 vdd.n2347 39.2114
R16982 vdd.n2415 vdd.n2348 39.2114
R16983 vdd.n2571 vdd.n2570 39.2114
R16984 vdd.n2358 vdd.n2333 39.2114
R16985 vdd.n2362 vdd.n2334 39.2114
R16986 vdd.n2366 vdd.n2335 39.2114
R16987 vdd.n2370 vdd.n2336 39.2114
R16988 vdd.n2374 vdd.n2337 39.2114
R16989 vdd.n2378 vdd.n2338 39.2114
R16990 vdd.n2382 vdd.n2339 39.2114
R16991 vdd.n2386 vdd.n2340 39.2114
R16992 vdd.n2390 vdd.n2341 39.2114
R16993 vdd.n2394 vdd.n2342 39.2114
R16994 vdd.n2398 vdd.n2343 39.2114
R16995 vdd.n2402 vdd.n2344 39.2114
R16996 vdd.n2406 vdd.n2345 39.2114
R16997 vdd.n2410 vdd.n2346 39.2114
R16998 vdd.n2414 vdd.n2347 39.2114
R16999 vdd.n2417 vdd.n2348 39.2114
R17000 vdd.n629 vdd.n624 39.2114
R17001 vdd.n2779 vdd.n2778 39.2114
R17002 vdd.n623 vdd.n621 39.2114
R17003 vdd.n2786 vdd.n2785 39.2114
R17004 vdd.n620 vdd.n618 39.2114
R17005 vdd.n2793 vdd.n2792 39.2114
R17006 vdd.n617 vdd.n615 39.2114
R17007 vdd.n2800 vdd.n2799 39.2114
R17008 vdd.n2803 vdd.n2802 39.2114
R17009 vdd.n2659 vdd.n2658 39.2114
R17010 vdd.n2664 vdd.n2663 39.2114
R17011 vdd.n2657 vdd.n2655 39.2114
R17012 vdd.n2671 vdd.n2670 39.2114
R17013 vdd.n2654 vdd.n2652 39.2114
R17014 vdd.n2678 vdd.n2677 39.2114
R17015 vdd.n2651 vdd.n2649 39.2114
R17016 vdd.n2685 vdd.n2684 39.2114
R17017 vdd.n1823 vdd.n1822 39.2114
R17018 vdd.n1829 vdd.n1828 39.2114
R17019 vdd.n1830 vdd.n1819 39.2114
R17020 vdd.n1837 vdd.n1836 39.2114
R17021 vdd.n1838 vdd.n1817 39.2114
R17022 vdd.n1845 vdd.n1844 39.2114
R17023 vdd.n1846 vdd.n1815 39.2114
R17024 vdd.n1853 vdd.n1852 39.2114
R17025 vdd.n2024 vdd.n2023 39.2114
R17026 vdd.n2021 vdd.n2020 39.2114
R17027 vdd.n2016 vdd.n2015 39.2114
R17028 vdd.n2013 vdd.n2012 39.2114
R17029 vdd.n2008 vdd.n2007 39.2114
R17030 vdd.n2005 vdd.n2004 39.2114
R17031 vdd.n2000 vdd.n1999 39.2114
R17032 vdd.n1997 vdd.n1996 39.2114
R17033 vdd.n1992 vdd.n1991 39.2114
R17034 vdd.n2249 vdd.n765 39.2114
R17035 vdd.n2254 vdd.n766 39.2114
R17036 vdd.n2258 vdd.n767 39.2114
R17037 vdd.n2262 vdd.n768 39.2114
R17038 vdd.n2266 vdd.n769 39.2114
R17039 vdd.n2270 vdd.n770 39.2114
R17040 vdd.n2274 vdd.n771 39.2114
R17041 vdd.n2278 vdd.n772 39.2114
R17042 vdd.n2282 vdd.n773 39.2114
R17043 vdd.n2286 vdd.n774 39.2114
R17044 vdd.n2290 vdd.n775 39.2114
R17045 vdd.n2294 vdd.n776 39.2114
R17046 vdd.n2298 vdd.n777 39.2114
R17047 vdd.n2302 vdd.n778 39.2114
R17048 vdd.n2306 vdd.n779 39.2114
R17049 vdd.n2310 vdd.n780 39.2114
R17050 vdd.n783 vdd.n781 39.2114
R17051 vdd.n2568 vdd.n2567 39.2114
R17052 vdd.n2561 vdd.n2317 39.2114
R17053 vdd.n2557 vdd.n2318 39.2114
R17054 vdd.n2553 vdd.n2319 39.2114
R17055 vdd.n2549 vdd.n2320 39.2114
R17056 vdd.n2545 vdd.n2321 39.2114
R17057 vdd.n2541 vdd.n2322 39.2114
R17058 vdd.n2537 vdd.n2323 39.2114
R17059 vdd.n2533 vdd.n2324 39.2114
R17060 vdd.n2529 vdd.n2325 39.2114
R17061 vdd.n2525 vdd.n2326 39.2114
R17062 vdd.n2521 vdd.n2327 39.2114
R17063 vdd.n2517 vdd.n2328 39.2114
R17064 vdd.n2513 vdd.n2329 39.2114
R17065 vdd.n2509 vdd.n2330 39.2114
R17066 vdd.n2504 vdd.n2331 39.2114
R17067 vdd.n2500 vdd.n2332 39.2114
R17068 vdd.n2706 vdd.n660 39.2114
R17069 vdd.n2713 vdd.n2712 39.2114
R17070 vdd.n659 vdd.n657 39.2114
R17071 vdd.n2720 vdd.n2719 39.2114
R17072 vdd.n656 vdd.n654 39.2114
R17073 vdd.n2727 vdd.n2726 39.2114
R17074 vdd.n653 vdd.n651 39.2114
R17075 vdd.n2734 vdd.n2733 39.2114
R17076 vdd.n650 vdd.n648 39.2114
R17077 vdd.n2742 vdd.n2741 39.2114
R17078 vdd.n647 vdd.n645 39.2114
R17079 vdd.n2749 vdd.n2748 39.2114
R17080 vdd.n644 vdd.n642 39.2114
R17081 vdd.n2756 vdd.n2755 39.2114
R17082 vdd.n641 vdd.n639 39.2114
R17083 vdd.n2763 vdd.n2762 39.2114
R17084 vdd.n2766 vdd.n2765 39.2114
R17085 vdd.n791 vdd.n747 39.2114
R17086 vdd.n2238 vdd.n748 39.2114
R17087 vdd.n2234 vdd.n749 39.2114
R17088 vdd.n2230 vdd.n750 39.2114
R17089 vdd.n2226 vdd.n751 39.2114
R17090 vdd.n2222 vdd.n752 39.2114
R17091 vdd.n2218 vdd.n753 39.2114
R17092 vdd.n2214 vdd.n754 39.2114
R17093 vdd.n2210 vdd.n755 39.2114
R17094 vdd.n2206 vdd.n756 39.2114
R17095 vdd.n2202 vdd.n757 39.2114
R17096 vdd.n2198 vdd.n758 39.2114
R17097 vdd.n2194 vdd.n759 39.2114
R17098 vdd.n2190 vdd.n760 39.2114
R17099 vdd.n2186 vdd.n761 39.2114
R17100 vdd.n2182 vdd.n762 39.2114
R17101 vdd.n2178 vdd.n763 39.2114
R17102 vdd.n2081 vdd.n880 39.2114
R17103 vdd.n2080 vdd.n2079 39.2114
R17104 vdd.n2073 vdd.n882 39.2114
R17105 vdd.n2072 vdd.n2071 39.2114
R17106 vdd.n2065 vdd.n884 39.2114
R17107 vdd.n2064 vdd.n2063 39.2114
R17108 vdd.n2057 vdd.n886 39.2114
R17109 vdd.n2056 vdd.n2055 39.2114
R17110 vdd.n889 vdd.n888 39.2114
R17111 vdd.n1897 vdd.n1896 39.2114
R17112 vdd.n1902 vdd.n1901 39.2114
R17113 vdd.n1905 vdd.n1904 39.2114
R17114 vdd.n1910 vdd.n1909 39.2114
R17115 vdd.n1913 vdd.n1912 39.2114
R17116 vdd.n1918 vdd.n1917 39.2114
R17117 vdd.n1921 vdd.n1920 39.2114
R17118 vdd.n1927 vdd.n1926 39.2114
R17119 vdd.n2175 vdd.n763 39.2114
R17120 vdd.n2179 vdd.n762 39.2114
R17121 vdd.n2183 vdd.n761 39.2114
R17122 vdd.n2187 vdd.n760 39.2114
R17123 vdd.n2191 vdd.n759 39.2114
R17124 vdd.n2195 vdd.n758 39.2114
R17125 vdd.n2199 vdd.n757 39.2114
R17126 vdd.n2203 vdd.n756 39.2114
R17127 vdd.n2207 vdd.n755 39.2114
R17128 vdd.n2211 vdd.n754 39.2114
R17129 vdd.n2215 vdd.n753 39.2114
R17130 vdd.n2219 vdd.n752 39.2114
R17131 vdd.n2223 vdd.n751 39.2114
R17132 vdd.n2227 vdd.n750 39.2114
R17133 vdd.n2231 vdd.n749 39.2114
R17134 vdd.n2235 vdd.n748 39.2114
R17135 vdd.n2239 vdd.n747 39.2114
R17136 vdd.n2082 vdd.n2081 39.2114
R17137 vdd.n2079 vdd.n2078 39.2114
R17138 vdd.n2074 vdd.n2073 39.2114
R17139 vdd.n2071 vdd.n2070 39.2114
R17140 vdd.n2066 vdd.n2065 39.2114
R17141 vdd.n2063 vdd.n2062 39.2114
R17142 vdd.n2058 vdd.n2057 39.2114
R17143 vdd.n2055 vdd.n2054 39.2114
R17144 vdd.n890 vdd.n889 39.2114
R17145 vdd.n1898 vdd.n1897 39.2114
R17146 vdd.n1903 vdd.n1902 39.2114
R17147 vdd.n1904 vdd.n1894 39.2114
R17148 vdd.n1911 vdd.n1910 39.2114
R17149 vdd.n1912 vdd.n1892 39.2114
R17150 vdd.n1919 vdd.n1918 39.2114
R17151 vdd.n1920 vdd.n1888 39.2114
R17152 vdd.n1928 vdd.n1927 39.2114
R17153 vdd.n2047 vdd.n2046 37.2369
R17154 vdd.n1750 vdd.n1683 37.2369
R17155 vdd.n1789 vdd.n1643 37.2369
R17156 vdd.n2854 vdd.n581 37.2369
R17157 vdd.n545 vdd.n544 37.2369
R17158 vdd.n2810 vdd.n2809 37.2369
R17159 vdd.n2089 vdd.n875 31.6883
R17160 vdd.n2314 vdd.n784 31.6883
R17161 vdd.n2247 vdd.n787 31.6883
R17162 vdd.n1993 vdd.n1990 31.6883
R17163 vdd.n2501 vdd.n2499 31.6883
R17164 vdd.n2708 vdd.n2705 31.6883
R17165 vdd.n2578 vdd.n740 31.6883
R17166 vdd.n2769 vdd.n2768 31.6883
R17167 vdd.n2688 vdd.n2687 31.6883
R17168 vdd.n2774 vdd.n628 31.6883
R17169 vdd.n2420 vdd.n2419 31.6883
R17170 vdd.n2574 vdd.n2573 31.6883
R17171 vdd.n2085 vdd.n2084 31.6883
R17172 vdd.n2242 vdd.n2241 31.6883
R17173 vdd.n2174 vdd.n2173 31.6883
R17174 vdd.n1931 vdd.n1930 31.6883
R17175 vdd.n1924 vdd.n1890 30.449
R17176 vdd.n795 vdd.n794 30.449
R17177 vdd.n1865 vdd.n1864 30.449
R17178 vdd.n2252 vdd.n786 30.449
R17179 vdd.n2356 vdd.n2355 30.449
R17180 vdd.n663 vdd.n662 30.449
R17181 vdd.n2506 vdd.n2352 30.449
R17182 vdd.n627 vdd.n626 30.449
R17183 vdd.n1215 vdd.n982 20.633
R17184 vdd.n2041 vdd.n901 20.633
R17185 vdd.n2940 vdd.n516 20.633
R17186 vdd.n3138 vdd.n351 20.633
R17187 vdd.n1217 vdd.n979 19.3944
R17188 vdd.n1221 vdd.n979 19.3944
R17189 vdd.n1221 vdd.n970 19.3944
R17190 vdd.n1233 vdd.n970 19.3944
R17191 vdd.n1233 vdd.n968 19.3944
R17192 vdd.n1237 vdd.n968 19.3944
R17193 vdd.n1237 vdd.n957 19.3944
R17194 vdd.n1249 vdd.n957 19.3944
R17195 vdd.n1249 vdd.n955 19.3944
R17196 vdd.n1253 vdd.n955 19.3944
R17197 vdd.n1253 vdd.n946 19.3944
R17198 vdd.n1266 vdd.n946 19.3944
R17199 vdd.n1266 vdd.n944 19.3944
R17200 vdd.n1270 vdd.n944 19.3944
R17201 vdd.n1270 vdd.n935 19.3944
R17202 vdd.n1564 vdd.n935 19.3944
R17203 vdd.n1564 vdd.n933 19.3944
R17204 vdd.n1568 vdd.n933 19.3944
R17205 vdd.n1568 vdd.n923 19.3944
R17206 vdd.n1581 vdd.n923 19.3944
R17207 vdd.n1581 vdd.n921 19.3944
R17208 vdd.n1585 vdd.n921 19.3944
R17209 vdd.n1585 vdd.n913 19.3944
R17210 vdd.n1598 vdd.n913 19.3944
R17211 vdd.n1598 vdd.n910 19.3944
R17212 vdd.n1604 vdd.n910 19.3944
R17213 vdd.n1604 vdd.n911 19.3944
R17214 vdd.n911 vdd.n900 19.3944
R17215 vdd.n1142 vdd.n1068 19.3944
R17216 vdd.n1142 vdd.n1070 19.3944
R17217 vdd.n1138 vdd.n1070 19.3944
R17218 vdd.n1138 vdd.n1137 19.3944
R17219 vdd.n1137 vdd.n1136 19.3944
R17220 vdd.n1136 vdd.n1078 19.3944
R17221 vdd.n1132 vdd.n1078 19.3944
R17222 vdd.n1132 vdd.n1131 19.3944
R17223 vdd.n1131 vdd.n1130 19.3944
R17224 vdd.n1130 vdd.n1086 19.3944
R17225 vdd.n1126 vdd.n1086 19.3944
R17226 vdd.n1126 vdd.n1125 19.3944
R17227 vdd.n1125 vdd.n1124 19.3944
R17228 vdd.n1124 vdd.n1094 19.3944
R17229 vdd.n1120 vdd.n1094 19.3944
R17230 vdd.n1120 vdd.n1119 19.3944
R17231 vdd.n1119 vdd.n1118 19.3944
R17232 vdd.n1118 vdd.n1102 19.3944
R17233 vdd.n1114 vdd.n1102 19.3944
R17234 vdd.n1114 vdd.n1113 19.3944
R17235 vdd.n1180 vdd.n1179 19.3944
R17236 vdd.n1179 vdd.n1178 19.3944
R17237 vdd.n1178 vdd.n1031 19.3944
R17238 vdd.n1174 vdd.n1031 19.3944
R17239 vdd.n1174 vdd.n1173 19.3944
R17240 vdd.n1173 vdd.n1172 19.3944
R17241 vdd.n1172 vdd.n1039 19.3944
R17242 vdd.n1168 vdd.n1039 19.3944
R17243 vdd.n1168 vdd.n1167 19.3944
R17244 vdd.n1167 vdd.n1166 19.3944
R17245 vdd.n1166 vdd.n1047 19.3944
R17246 vdd.n1162 vdd.n1047 19.3944
R17247 vdd.n1162 vdd.n1161 19.3944
R17248 vdd.n1161 vdd.n1160 19.3944
R17249 vdd.n1160 vdd.n1055 19.3944
R17250 vdd.n1156 vdd.n1055 19.3944
R17251 vdd.n1156 vdd.n1155 19.3944
R17252 vdd.n1155 vdd.n1154 19.3944
R17253 vdd.n1154 vdd.n1063 19.3944
R17254 vdd.n1150 vdd.n1063 19.3944
R17255 vdd.n1210 vdd.n1209 19.3944
R17256 vdd.n1209 vdd.n1208 19.3944
R17257 vdd.n1208 vdd.n989 19.3944
R17258 vdd.n1204 vdd.n989 19.3944
R17259 vdd.n1204 vdd.n1203 19.3944
R17260 vdd.n1203 vdd.n1202 19.3944
R17261 vdd.n1202 vdd.n997 19.3944
R17262 vdd.n1198 vdd.n997 19.3944
R17263 vdd.n1198 vdd.n1197 19.3944
R17264 vdd.n1197 vdd.n1196 19.3944
R17265 vdd.n1196 vdd.n1005 19.3944
R17266 vdd.n1192 vdd.n1005 19.3944
R17267 vdd.n1192 vdd.n1191 19.3944
R17268 vdd.n1191 vdd.n1190 19.3944
R17269 vdd.n1190 vdd.n1013 19.3944
R17270 vdd.n1186 vdd.n1013 19.3944
R17271 vdd.n1186 vdd.n1185 19.3944
R17272 vdd.n1185 vdd.n1184 19.3944
R17273 vdd.n1746 vdd.n1681 19.3944
R17274 vdd.n1746 vdd.n1687 19.3944
R17275 vdd.n1741 vdd.n1687 19.3944
R17276 vdd.n1741 vdd.n1740 19.3944
R17277 vdd.n1740 vdd.n1739 19.3944
R17278 vdd.n1739 vdd.n1694 19.3944
R17279 vdd.n1734 vdd.n1694 19.3944
R17280 vdd.n1734 vdd.n1733 19.3944
R17281 vdd.n1733 vdd.n1732 19.3944
R17282 vdd.n1732 vdd.n1701 19.3944
R17283 vdd.n1727 vdd.n1701 19.3944
R17284 vdd.n1727 vdd.n1726 19.3944
R17285 vdd.n1726 vdd.n1725 19.3944
R17286 vdd.n1725 vdd.n1709 19.3944
R17287 vdd.n1720 vdd.n1709 19.3944
R17288 vdd.n1720 vdd.n1719 19.3944
R17289 vdd.n1715 vdd.n1714 19.3944
R17290 vdd.n2048 vdd.n896 19.3944
R17291 vdd.n1785 vdd.n1641 19.3944
R17292 vdd.n1785 vdd.n1647 19.3944
R17293 vdd.n1780 vdd.n1647 19.3944
R17294 vdd.n1780 vdd.n1779 19.3944
R17295 vdd.n1779 vdd.n1778 19.3944
R17296 vdd.n1778 vdd.n1654 19.3944
R17297 vdd.n1773 vdd.n1654 19.3944
R17298 vdd.n1773 vdd.n1772 19.3944
R17299 vdd.n1772 vdd.n1771 19.3944
R17300 vdd.n1771 vdd.n1661 19.3944
R17301 vdd.n1766 vdd.n1661 19.3944
R17302 vdd.n1766 vdd.n1765 19.3944
R17303 vdd.n1765 vdd.n1764 19.3944
R17304 vdd.n1764 vdd.n1668 19.3944
R17305 vdd.n1759 vdd.n1668 19.3944
R17306 vdd.n1759 vdd.n1758 19.3944
R17307 vdd.n1758 vdd.n1757 19.3944
R17308 vdd.n1757 vdd.n1675 19.3944
R17309 vdd.n1752 vdd.n1675 19.3944
R17310 vdd.n1752 vdd.n1751 19.3944
R17311 vdd.n2036 vdd.n2035 19.3944
R17312 vdd.n2035 vdd.n1613 19.3944
R17313 vdd.n2030 vdd.n2029 19.3944
R17314 vdd.n1812 vdd.n1617 19.3944
R17315 vdd.n1812 vdd.n1619 19.3944
R17316 vdd.n1622 vdd.n1619 19.3944
R17317 vdd.n1805 vdd.n1622 19.3944
R17318 vdd.n1805 vdd.n1804 19.3944
R17319 vdd.n1804 vdd.n1803 19.3944
R17320 vdd.n1803 vdd.n1628 19.3944
R17321 vdd.n1798 vdd.n1628 19.3944
R17322 vdd.n1798 vdd.n1797 19.3944
R17323 vdd.n1797 vdd.n1796 19.3944
R17324 vdd.n1796 vdd.n1635 19.3944
R17325 vdd.n1791 vdd.n1635 19.3944
R17326 vdd.n1791 vdd.n1790 19.3944
R17327 vdd.n1213 vdd.n976 19.3944
R17328 vdd.n1225 vdd.n976 19.3944
R17329 vdd.n1225 vdd.n974 19.3944
R17330 vdd.n1229 vdd.n974 19.3944
R17331 vdd.n1229 vdd.n964 19.3944
R17332 vdd.n1241 vdd.n964 19.3944
R17333 vdd.n1241 vdd.n962 19.3944
R17334 vdd.n1245 vdd.n962 19.3944
R17335 vdd.n1245 vdd.n952 19.3944
R17336 vdd.n1258 vdd.n952 19.3944
R17337 vdd.n1258 vdd.n950 19.3944
R17338 vdd.n1262 vdd.n950 19.3944
R17339 vdd.n1262 vdd.n941 19.3944
R17340 vdd.n1274 vdd.n941 19.3944
R17341 vdd.n1274 vdd.n939 19.3944
R17342 vdd.n1560 vdd.n939 19.3944
R17343 vdd.n1560 vdd.n929 19.3944
R17344 vdd.n1573 vdd.n929 19.3944
R17345 vdd.n1573 vdd.n927 19.3944
R17346 vdd.n1577 vdd.n927 19.3944
R17347 vdd.n1577 vdd.n918 19.3944
R17348 vdd.n1590 vdd.n918 19.3944
R17349 vdd.n1590 vdd.n916 19.3944
R17350 vdd.n1594 vdd.n916 19.3944
R17351 vdd.n1594 vdd.n906 19.3944
R17352 vdd.n1609 vdd.n906 19.3944
R17353 vdd.n1609 vdd.n904 19.3944
R17354 vdd.n2039 vdd.n904 19.3944
R17355 vdd.n2942 vdd.n513 19.3944
R17356 vdd.n2946 vdd.n513 19.3944
R17357 vdd.n2946 vdd.n503 19.3944
R17358 vdd.n2958 vdd.n503 19.3944
R17359 vdd.n2958 vdd.n501 19.3944
R17360 vdd.n2962 vdd.n501 19.3944
R17361 vdd.n2962 vdd.n490 19.3944
R17362 vdd.n2974 vdd.n490 19.3944
R17363 vdd.n2974 vdd.n488 19.3944
R17364 vdd.n2978 vdd.n488 19.3944
R17365 vdd.n2978 vdd.n478 19.3944
R17366 vdd.n2991 vdd.n478 19.3944
R17367 vdd.n2991 vdd.n476 19.3944
R17368 vdd.n2995 vdd.n476 19.3944
R17369 vdd.n2996 vdd.n2995 19.3944
R17370 vdd.n2997 vdd.n2996 19.3944
R17371 vdd.n2997 vdd.n474 19.3944
R17372 vdd.n3001 vdd.n474 19.3944
R17373 vdd.n3002 vdd.n3001 19.3944
R17374 vdd.n3003 vdd.n3002 19.3944
R17375 vdd.n3003 vdd.n471 19.3944
R17376 vdd.n3007 vdd.n471 19.3944
R17377 vdd.n3008 vdd.n3007 19.3944
R17378 vdd.n3009 vdd.n3008 19.3944
R17379 vdd.n3009 vdd.n468 19.3944
R17380 vdd.n3013 vdd.n468 19.3944
R17381 vdd.n3014 vdd.n3013 19.3944
R17382 vdd.n3015 vdd.n3014 19.3944
R17383 vdd.n3058 vdd.n426 19.3944
R17384 vdd.n3058 vdd.n432 19.3944
R17385 vdd.n3053 vdd.n432 19.3944
R17386 vdd.n3053 vdd.n3052 19.3944
R17387 vdd.n3052 vdd.n3051 19.3944
R17388 vdd.n3051 vdd.n439 19.3944
R17389 vdd.n3046 vdd.n439 19.3944
R17390 vdd.n3046 vdd.n3045 19.3944
R17391 vdd.n3045 vdd.n3044 19.3944
R17392 vdd.n3044 vdd.n446 19.3944
R17393 vdd.n3039 vdd.n446 19.3944
R17394 vdd.n3039 vdd.n3038 19.3944
R17395 vdd.n3038 vdd.n3037 19.3944
R17396 vdd.n3037 vdd.n453 19.3944
R17397 vdd.n3032 vdd.n453 19.3944
R17398 vdd.n3032 vdd.n3031 19.3944
R17399 vdd.n3031 vdd.n3030 19.3944
R17400 vdd.n3030 vdd.n460 19.3944
R17401 vdd.n3025 vdd.n460 19.3944
R17402 vdd.n3025 vdd.n3024 19.3944
R17403 vdd.n3097 vdd.n386 19.3944
R17404 vdd.n3097 vdd.n392 19.3944
R17405 vdd.n3092 vdd.n392 19.3944
R17406 vdd.n3092 vdd.n3091 19.3944
R17407 vdd.n3091 vdd.n3090 19.3944
R17408 vdd.n3090 vdd.n399 19.3944
R17409 vdd.n3085 vdd.n399 19.3944
R17410 vdd.n3085 vdd.n3084 19.3944
R17411 vdd.n3084 vdd.n3083 19.3944
R17412 vdd.n3083 vdd.n406 19.3944
R17413 vdd.n3078 vdd.n406 19.3944
R17414 vdd.n3078 vdd.n3077 19.3944
R17415 vdd.n3077 vdd.n3076 19.3944
R17416 vdd.n3076 vdd.n413 19.3944
R17417 vdd.n3071 vdd.n413 19.3944
R17418 vdd.n3071 vdd.n3070 19.3944
R17419 vdd.n3070 vdd.n3069 19.3944
R17420 vdd.n3069 vdd.n420 19.3944
R17421 vdd.n3064 vdd.n420 19.3944
R17422 vdd.n3064 vdd.n3063 19.3944
R17423 vdd.n3133 vdd.n3132 19.3944
R17424 vdd.n3132 vdd.n3131 19.3944
R17425 vdd.n3131 vdd.n358 19.3944
R17426 vdd.n359 vdd.n358 19.3944
R17427 vdd.n3124 vdd.n359 19.3944
R17428 vdd.n3124 vdd.n3123 19.3944
R17429 vdd.n3123 vdd.n3122 19.3944
R17430 vdd.n3122 vdd.n366 19.3944
R17431 vdd.n3117 vdd.n366 19.3944
R17432 vdd.n3117 vdd.n3116 19.3944
R17433 vdd.n3116 vdd.n3115 19.3944
R17434 vdd.n3115 vdd.n373 19.3944
R17435 vdd.n3110 vdd.n373 19.3944
R17436 vdd.n3110 vdd.n3109 19.3944
R17437 vdd.n3109 vdd.n3108 19.3944
R17438 vdd.n3108 vdd.n380 19.3944
R17439 vdd.n3103 vdd.n380 19.3944
R17440 vdd.n3103 vdd.n3102 19.3944
R17441 vdd.n2938 vdd.n509 19.3944
R17442 vdd.n2950 vdd.n509 19.3944
R17443 vdd.n2950 vdd.n507 19.3944
R17444 vdd.n2954 vdd.n507 19.3944
R17445 vdd.n2954 vdd.n497 19.3944
R17446 vdd.n2966 vdd.n497 19.3944
R17447 vdd.n2966 vdd.n495 19.3944
R17448 vdd.n2970 vdd.n495 19.3944
R17449 vdd.n2970 vdd.n485 19.3944
R17450 vdd.n2983 vdd.n485 19.3944
R17451 vdd.n2983 vdd.n483 19.3944
R17452 vdd.n2987 vdd.n483 19.3944
R17453 vdd.n2987 vdd.n312 19.3944
R17454 vdd.n3166 vdd.n312 19.3944
R17455 vdd.n3166 vdd.n313 19.3944
R17456 vdd.n3160 vdd.n313 19.3944
R17457 vdd.n3160 vdd.n3159 19.3944
R17458 vdd.n3159 vdd.n3158 19.3944
R17459 vdd.n3158 vdd.n323 19.3944
R17460 vdd.n3152 vdd.n323 19.3944
R17461 vdd.n3152 vdd.n3151 19.3944
R17462 vdd.n3151 vdd.n3150 19.3944
R17463 vdd.n3150 vdd.n335 19.3944
R17464 vdd.n3144 vdd.n335 19.3944
R17465 vdd.n3144 vdd.n3143 19.3944
R17466 vdd.n3143 vdd.n3142 19.3944
R17467 vdd.n3142 vdd.n346 19.3944
R17468 vdd.n3136 vdd.n346 19.3944
R17469 vdd.n2895 vdd.n2894 19.3944
R17470 vdd.n2894 vdd.n2893 19.3944
R17471 vdd.n2893 vdd.n551 19.3944
R17472 vdd.n2887 vdd.n551 19.3944
R17473 vdd.n2887 vdd.n2886 19.3944
R17474 vdd.n2886 vdd.n2885 19.3944
R17475 vdd.n2885 vdd.n557 19.3944
R17476 vdd.n2879 vdd.n557 19.3944
R17477 vdd.n2879 vdd.n2878 19.3944
R17478 vdd.n2878 vdd.n2877 19.3944
R17479 vdd.n2877 vdd.n563 19.3944
R17480 vdd.n2871 vdd.n563 19.3944
R17481 vdd.n2871 vdd.n2870 19.3944
R17482 vdd.n2870 vdd.n2869 19.3944
R17483 vdd.n2869 vdd.n569 19.3944
R17484 vdd.n2863 vdd.n569 19.3944
R17485 vdd.n2863 vdd.n2862 19.3944
R17486 vdd.n2862 vdd.n2861 19.3944
R17487 vdd.n2861 vdd.n575 19.3944
R17488 vdd.n2855 vdd.n575 19.3944
R17489 vdd.n2935 vdd.n2934 19.3944
R17490 vdd.n2934 vdd.n519 19.3944
R17491 vdd.n2929 vdd.n2928 19.3944
R17492 vdd.n2925 vdd.n2924 19.3944
R17493 vdd.n2924 vdd.n525 19.3944
R17494 vdd.n2919 vdd.n525 19.3944
R17495 vdd.n2919 vdd.n2918 19.3944
R17496 vdd.n2918 vdd.n2917 19.3944
R17497 vdd.n2917 vdd.n531 19.3944
R17498 vdd.n2911 vdd.n531 19.3944
R17499 vdd.n2911 vdd.n2910 19.3944
R17500 vdd.n2910 vdd.n2909 19.3944
R17501 vdd.n2909 vdd.n537 19.3944
R17502 vdd.n2903 vdd.n537 19.3944
R17503 vdd.n2903 vdd.n2902 19.3944
R17504 vdd.n2902 vdd.n2901 19.3944
R17505 vdd.n2850 vdd.n579 19.3944
R17506 vdd.n2850 vdd.n583 19.3944
R17507 vdd.n2845 vdd.n583 19.3944
R17508 vdd.n2845 vdd.n2844 19.3944
R17509 vdd.n2844 vdd.n589 19.3944
R17510 vdd.n2839 vdd.n589 19.3944
R17511 vdd.n2839 vdd.n2838 19.3944
R17512 vdd.n2838 vdd.n2837 19.3944
R17513 vdd.n2837 vdd.n595 19.3944
R17514 vdd.n2831 vdd.n595 19.3944
R17515 vdd.n2831 vdd.n2830 19.3944
R17516 vdd.n2830 vdd.n2829 19.3944
R17517 vdd.n2829 vdd.n601 19.3944
R17518 vdd.n2823 vdd.n601 19.3944
R17519 vdd.n2823 vdd.n2822 19.3944
R17520 vdd.n2822 vdd.n2821 19.3944
R17521 vdd.n2817 vdd.n2816 19.3944
R17522 vdd.n2813 vdd.n2812 19.3944
R17523 vdd.n1149 vdd.n1068 19.0066
R17524 vdd.n1750 vdd.n1681 19.0066
R17525 vdd.n3062 vdd.n426 19.0066
R17526 vdd.n2854 vdd.n579 19.0066
R17527 vdd.n1890 vdd.n1889 16.0975
R17528 vdd.n794 vdd.n793 16.0975
R17529 vdd.n1111 vdd.n1110 16.0975
R17530 vdd.n1148 vdd.n1147 16.0975
R17531 vdd.n1022 vdd.n1021 16.0975
R17532 vdd.n2046 vdd.n2045 16.0975
R17533 vdd.n1683 vdd.n1682 16.0975
R17534 vdd.n1643 vdd.n1642 16.0975
R17535 vdd.n1864 vdd.n1863 16.0975
R17536 vdd.n786 vdd.n785 16.0975
R17537 vdd.n2355 vdd.n2354 16.0975
R17538 vdd.n3022 vdd.n3021 16.0975
R17539 vdd.n428 vdd.n427 16.0975
R17540 vdd.n388 vdd.n387 16.0975
R17541 vdd.n581 vdd.n580 16.0975
R17542 vdd.n544 vdd.n543 16.0975
R17543 vdd.n662 vdd.n661 16.0975
R17544 vdd.n2352 vdd.n2351 16.0975
R17545 vdd.n2809 vdd.n2808 16.0975
R17546 vdd.n626 vdd.n625 16.0975
R17547 vdd.t17 vdd.n2316 15.4182
R17548 vdd.n2569 vdd.t200 15.4182
R17549 vdd.n28 vdd.n27 14.5458
R17550 vdd.n2087 vdd.n877 14.5112
R17551 vdd.n2771 vdd.n613 14.5112
R17552 vdd.n304 vdd.n269 13.1884
R17553 vdd.n253 vdd.n218 13.1884
R17554 vdd.n210 vdd.n175 13.1884
R17555 vdd.n159 vdd.n124 13.1884
R17556 vdd.n117 vdd.n82 13.1884
R17557 vdd.n66 vdd.n31 13.1884
R17558 vdd.n1499 vdd.n1464 13.1884
R17559 vdd.n1550 vdd.n1515 13.1884
R17560 vdd.n1405 vdd.n1370 13.1884
R17561 vdd.n1456 vdd.n1421 13.1884
R17562 vdd.n1312 vdd.n1277 13.1884
R17563 vdd.n1363 vdd.n1328 13.1884
R17564 vdd.n1180 vdd.n1023 12.9944
R17565 vdd.n1184 vdd.n1023 12.9944
R17566 vdd.n1789 vdd.n1641 12.9944
R17567 vdd.n1790 vdd.n1789 12.9944
R17568 vdd.n3101 vdd.n386 12.9944
R17569 vdd.n3102 vdd.n3101 12.9944
R17570 vdd.n2895 vdd.n545 12.9944
R17571 vdd.n2901 vdd.n545 12.9944
R17572 vdd.n305 vdd.n267 12.8005
R17573 vdd.n300 vdd.n271 12.8005
R17574 vdd.n254 vdd.n216 12.8005
R17575 vdd.n249 vdd.n220 12.8005
R17576 vdd.n211 vdd.n173 12.8005
R17577 vdd.n206 vdd.n177 12.8005
R17578 vdd.n160 vdd.n122 12.8005
R17579 vdd.n155 vdd.n126 12.8005
R17580 vdd.n118 vdd.n80 12.8005
R17581 vdd.n113 vdd.n84 12.8005
R17582 vdd.n67 vdd.n29 12.8005
R17583 vdd.n62 vdd.n33 12.8005
R17584 vdd.n1500 vdd.n1462 12.8005
R17585 vdd.n1495 vdd.n1466 12.8005
R17586 vdd.n1551 vdd.n1513 12.8005
R17587 vdd.n1546 vdd.n1517 12.8005
R17588 vdd.n1406 vdd.n1368 12.8005
R17589 vdd.n1401 vdd.n1372 12.8005
R17590 vdd.n1457 vdd.n1419 12.8005
R17591 vdd.n1452 vdd.n1423 12.8005
R17592 vdd.n1313 vdd.n1275 12.8005
R17593 vdd.n1308 vdd.n1279 12.8005
R17594 vdd.n1364 vdd.n1326 12.8005
R17595 vdd.n1359 vdd.n1330 12.8005
R17596 vdd.n299 vdd.n272 12.0247
R17597 vdd.n248 vdd.n221 12.0247
R17598 vdd.n205 vdd.n178 12.0247
R17599 vdd.n154 vdd.n127 12.0247
R17600 vdd.n112 vdd.n85 12.0247
R17601 vdd.n61 vdd.n34 12.0247
R17602 vdd.n1494 vdd.n1467 12.0247
R17603 vdd.n1545 vdd.n1518 12.0247
R17604 vdd.n1400 vdd.n1373 12.0247
R17605 vdd.n1451 vdd.n1424 12.0247
R17606 vdd.n1307 vdd.n1280 12.0247
R17607 vdd.n1358 vdd.n1331 12.0247
R17608 vdd.n1215 vdd.n983 11.337
R17609 vdd.n1223 vdd.n972 11.337
R17610 vdd.n1231 vdd.n972 11.337
R17611 vdd.n1239 vdd.n966 11.337
R17612 vdd.n1247 vdd.n959 11.337
R17613 vdd.n1256 vdd.n1255 11.337
R17614 vdd.n1264 vdd.n948 11.337
R17615 vdd.n1562 vdd.n937 11.337
R17616 vdd.n1571 vdd.n931 11.337
R17617 vdd.n1579 vdd.n925 11.337
R17618 vdd.n1588 vdd.n1587 11.337
R17619 vdd.n1596 vdd.n908 11.337
R17620 vdd.n1607 vdd.n908 11.337
R17621 vdd.n1607 vdd.n1606 11.337
R17622 vdd.n2948 vdd.n511 11.337
R17623 vdd.n2948 vdd.n505 11.337
R17624 vdd.n2956 vdd.n505 11.337
R17625 vdd.n2964 vdd.n499 11.337
R17626 vdd.n2972 vdd.n492 11.337
R17627 vdd.n2981 vdd.n2980 11.337
R17628 vdd.n2989 vdd.n481 11.337
R17629 vdd.n3163 vdd.n3162 11.337
R17630 vdd.n3156 vdd.n325 11.337
R17631 vdd.n3154 vdd.n329 11.337
R17632 vdd.n3148 vdd.n3147 11.337
R17633 vdd.n3146 vdd.n340 11.337
R17634 vdd.n3140 vdd.n340 11.337
R17635 vdd.n3139 vdd.n3138 11.337
R17636 vdd.n296 vdd.n295 11.249
R17637 vdd.n245 vdd.n244 11.249
R17638 vdd.n202 vdd.n201 11.249
R17639 vdd.n151 vdd.n150 11.249
R17640 vdd.n109 vdd.n108 11.249
R17641 vdd.n58 vdd.n57 11.249
R17642 vdd.n1491 vdd.n1490 11.249
R17643 vdd.n1542 vdd.n1541 11.249
R17644 vdd.n1397 vdd.n1396 11.249
R17645 vdd.n1448 vdd.n1447 11.249
R17646 vdd.n1304 vdd.n1303 11.249
R17647 vdd.n1355 vdd.n1354 11.249
R17648 vdd.n2244 vdd.t163 11.1103
R17649 vdd.n2576 vdd.t172 11.1103
R17650 vdd.n1231 vdd.t46 10.9969
R17651 vdd.t152 vdd.n3146 10.9969
R17652 vdd.n960 vdd.t32 10.7702
R17653 vdd.t138 vdd.n3155 10.7702
R17654 vdd.n281 vdd.n280 10.7238
R17655 vdd.n230 vdd.n229 10.7238
R17656 vdd.n187 vdd.n186 10.7238
R17657 vdd.n136 vdd.n135 10.7238
R17658 vdd.n94 vdd.n93 10.7238
R17659 vdd.n43 vdd.n42 10.7238
R17660 vdd.n1476 vdd.n1475 10.7238
R17661 vdd.n1527 vdd.n1526 10.7238
R17662 vdd.n1382 vdd.n1381 10.7238
R17663 vdd.n1433 vdd.n1432 10.7238
R17664 vdd.n1289 vdd.n1288 10.7238
R17665 vdd.n1340 vdd.n1339 10.7238
R17666 vdd.n2090 vdd.n2089 10.6151
R17667 vdd.n2091 vdd.n2090 10.6151
R17668 vdd.n2091 vdd.n863 10.6151
R17669 vdd.n2101 vdd.n863 10.6151
R17670 vdd.n2102 vdd.n2101 10.6151
R17671 vdd.n2103 vdd.n2102 10.6151
R17672 vdd.n2103 vdd.n850 10.6151
R17673 vdd.n2114 vdd.n850 10.6151
R17674 vdd.n2115 vdd.n2114 10.6151
R17675 vdd.n2116 vdd.n2115 10.6151
R17676 vdd.n2116 vdd.n838 10.6151
R17677 vdd.n2126 vdd.n838 10.6151
R17678 vdd.n2127 vdd.n2126 10.6151
R17679 vdd.n2128 vdd.n2127 10.6151
R17680 vdd.n2128 vdd.n826 10.6151
R17681 vdd.n2138 vdd.n826 10.6151
R17682 vdd.n2139 vdd.n2138 10.6151
R17683 vdd.n2140 vdd.n2139 10.6151
R17684 vdd.n2140 vdd.n815 10.6151
R17685 vdd.n2150 vdd.n815 10.6151
R17686 vdd.n2151 vdd.n2150 10.6151
R17687 vdd.n2152 vdd.n2151 10.6151
R17688 vdd.n2152 vdd.n802 10.6151
R17689 vdd.n2164 vdd.n802 10.6151
R17690 vdd.n2165 vdd.n2164 10.6151
R17691 vdd.n2167 vdd.n2165 10.6151
R17692 vdd.n2167 vdd.n2166 10.6151
R17693 vdd.n2166 vdd.n784 10.6151
R17694 vdd.n2314 vdd.n2313 10.6151
R17695 vdd.n2313 vdd.n2312 10.6151
R17696 vdd.n2312 vdd.n2309 10.6151
R17697 vdd.n2309 vdd.n2308 10.6151
R17698 vdd.n2308 vdd.n2305 10.6151
R17699 vdd.n2305 vdd.n2304 10.6151
R17700 vdd.n2304 vdd.n2301 10.6151
R17701 vdd.n2301 vdd.n2300 10.6151
R17702 vdd.n2300 vdd.n2297 10.6151
R17703 vdd.n2297 vdd.n2296 10.6151
R17704 vdd.n2296 vdd.n2293 10.6151
R17705 vdd.n2293 vdd.n2292 10.6151
R17706 vdd.n2292 vdd.n2289 10.6151
R17707 vdd.n2289 vdd.n2288 10.6151
R17708 vdd.n2288 vdd.n2285 10.6151
R17709 vdd.n2285 vdd.n2284 10.6151
R17710 vdd.n2284 vdd.n2281 10.6151
R17711 vdd.n2281 vdd.n2280 10.6151
R17712 vdd.n2280 vdd.n2277 10.6151
R17713 vdd.n2277 vdd.n2276 10.6151
R17714 vdd.n2276 vdd.n2273 10.6151
R17715 vdd.n2273 vdd.n2272 10.6151
R17716 vdd.n2272 vdd.n2269 10.6151
R17717 vdd.n2269 vdd.n2268 10.6151
R17718 vdd.n2268 vdd.n2265 10.6151
R17719 vdd.n2265 vdd.n2264 10.6151
R17720 vdd.n2264 vdd.n2261 10.6151
R17721 vdd.n2261 vdd.n2260 10.6151
R17722 vdd.n2260 vdd.n2257 10.6151
R17723 vdd.n2257 vdd.n2256 10.6151
R17724 vdd.n2256 vdd.n2253 10.6151
R17725 vdd.n2251 vdd.n2248 10.6151
R17726 vdd.n2248 vdd.n2247 10.6151
R17727 vdd.n1990 vdd.n1989 10.6151
R17728 vdd.n1989 vdd.n1987 10.6151
R17729 vdd.n1987 vdd.n1986 10.6151
R17730 vdd.n1986 vdd.n1984 10.6151
R17731 vdd.n1984 vdd.n1983 10.6151
R17732 vdd.n1983 vdd.n1981 10.6151
R17733 vdd.n1981 vdd.n1980 10.6151
R17734 vdd.n1980 vdd.n1978 10.6151
R17735 vdd.n1978 vdd.n1977 10.6151
R17736 vdd.n1977 vdd.n1975 10.6151
R17737 vdd.n1975 vdd.n1974 10.6151
R17738 vdd.n1974 vdd.n1972 10.6151
R17739 vdd.n1972 vdd.n1971 10.6151
R17740 vdd.n1971 vdd.n1886 10.6151
R17741 vdd.n1886 vdd.n1885 10.6151
R17742 vdd.n1885 vdd.n1883 10.6151
R17743 vdd.n1883 vdd.n1882 10.6151
R17744 vdd.n1882 vdd.n1880 10.6151
R17745 vdd.n1880 vdd.n1879 10.6151
R17746 vdd.n1879 vdd.n1877 10.6151
R17747 vdd.n1877 vdd.n1876 10.6151
R17748 vdd.n1876 vdd.n1874 10.6151
R17749 vdd.n1874 vdd.n1873 10.6151
R17750 vdd.n1873 vdd.n1871 10.6151
R17751 vdd.n1871 vdd.n1870 10.6151
R17752 vdd.n1870 vdd.n1867 10.6151
R17753 vdd.n1867 vdd.n1866 10.6151
R17754 vdd.n1866 vdd.n787 10.6151
R17755 vdd.n1824 vdd.n875 10.6151
R17756 vdd.n1825 vdd.n1824 10.6151
R17757 vdd.n1826 vdd.n1825 10.6151
R17758 vdd.n1826 vdd.n1820 10.6151
R17759 vdd.n1832 vdd.n1820 10.6151
R17760 vdd.n1833 vdd.n1832 10.6151
R17761 vdd.n1834 vdd.n1833 10.6151
R17762 vdd.n1834 vdd.n1818 10.6151
R17763 vdd.n1840 vdd.n1818 10.6151
R17764 vdd.n1841 vdd.n1840 10.6151
R17765 vdd.n1842 vdd.n1841 10.6151
R17766 vdd.n1842 vdd.n1816 10.6151
R17767 vdd.n1848 vdd.n1816 10.6151
R17768 vdd.n1849 vdd.n1848 10.6151
R17769 vdd.n1850 vdd.n1849 10.6151
R17770 vdd.n1850 vdd.n1814 10.6151
R17771 vdd.n2026 vdd.n1814 10.6151
R17772 vdd.n2026 vdd.n2025 10.6151
R17773 vdd.n2025 vdd.n1855 10.6151
R17774 vdd.n2019 vdd.n1855 10.6151
R17775 vdd.n2019 vdd.n2018 10.6151
R17776 vdd.n2018 vdd.n2017 10.6151
R17777 vdd.n2017 vdd.n1857 10.6151
R17778 vdd.n2011 vdd.n1857 10.6151
R17779 vdd.n2011 vdd.n2010 10.6151
R17780 vdd.n2010 vdd.n2009 10.6151
R17781 vdd.n2009 vdd.n1859 10.6151
R17782 vdd.n2003 vdd.n1859 10.6151
R17783 vdd.n2003 vdd.n2002 10.6151
R17784 vdd.n2002 vdd.n2001 10.6151
R17785 vdd.n2001 vdd.n1861 10.6151
R17786 vdd.n1995 vdd.n1994 10.6151
R17787 vdd.n1994 vdd.n1993 10.6151
R17788 vdd.n2499 vdd.n2498 10.6151
R17789 vdd.n2498 vdd.n2496 10.6151
R17790 vdd.n2496 vdd.n2495 10.6151
R17791 vdd.n2495 vdd.n2353 10.6151
R17792 vdd.n2442 vdd.n2353 10.6151
R17793 vdd.n2443 vdd.n2442 10.6151
R17794 vdd.n2445 vdd.n2443 10.6151
R17795 vdd.n2446 vdd.n2445 10.6151
R17796 vdd.n2448 vdd.n2446 10.6151
R17797 vdd.n2449 vdd.n2448 10.6151
R17798 vdd.n2451 vdd.n2449 10.6151
R17799 vdd.n2452 vdd.n2451 10.6151
R17800 vdd.n2454 vdd.n2452 10.6151
R17801 vdd.n2455 vdd.n2454 10.6151
R17802 vdd.n2470 vdd.n2455 10.6151
R17803 vdd.n2470 vdd.n2469 10.6151
R17804 vdd.n2469 vdd.n2468 10.6151
R17805 vdd.n2468 vdd.n2466 10.6151
R17806 vdd.n2466 vdd.n2465 10.6151
R17807 vdd.n2465 vdd.n2463 10.6151
R17808 vdd.n2463 vdd.n2462 10.6151
R17809 vdd.n2462 vdd.n2460 10.6151
R17810 vdd.n2460 vdd.n2459 10.6151
R17811 vdd.n2459 vdd.n2457 10.6151
R17812 vdd.n2457 vdd.n2456 10.6151
R17813 vdd.n2456 vdd.n664 10.6151
R17814 vdd.n2704 vdd.n664 10.6151
R17815 vdd.n2705 vdd.n2704 10.6151
R17816 vdd.n2566 vdd.n740 10.6151
R17817 vdd.n2566 vdd.n2565 10.6151
R17818 vdd.n2565 vdd.n2564 10.6151
R17819 vdd.n2564 vdd.n2562 10.6151
R17820 vdd.n2562 vdd.n2559 10.6151
R17821 vdd.n2559 vdd.n2558 10.6151
R17822 vdd.n2558 vdd.n2555 10.6151
R17823 vdd.n2555 vdd.n2554 10.6151
R17824 vdd.n2554 vdd.n2551 10.6151
R17825 vdd.n2551 vdd.n2550 10.6151
R17826 vdd.n2550 vdd.n2547 10.6151
R17827 vdd.n2547 vdd.n2546 10.6151
R17828 vdd.n2546 vdd.n2543 10.6151
R17829 vdd.n2543 vdd.n2542 10.6151
R17830 vdd.n2542 vdd.n2539 10.6151
R17831 vdd.n2539 vdd.n2538 10.6151
R17832 vdd.n2538 vdd.n2535 10.6151
R17833 vdd.n2535 vdd.n2534 10.6151
R17834 vdd.n2534 vdd.n2531 10.6151
R17835 vdd.n2531 vdd.n2530 10.6151
R17836 vdd.n2530 vdd.n2527 10.6151
R17837 vdd.n2527 vdd.n2526 10.6151
R17838 vdd.n2526 vdd.n2523 10.6151
R17839 vdd.n2523 vdd.n2522 10.6151
R17840 vdd.n2522 vdd.n2519 10.6151
R17841 vdd.n2519 vdd.n2518 10.6151
R17842 vdd.n2518 vdd.n2515 10.6151
R17843 vdd.n2515 vdd.n2514 10.6151
R17844 vdd.n2514 vdd.n2511 10.6151
R17845 vdd.n2511 vdd.n2510 10.6151
R17846 vdd.n2510 vdd.n2507 10.6151
R17847 vdd.n2505 vdd.n2502 10.6151
R17848 vdd.n2502 vdd.n2501 10.6151
R17849 vdd.n2579 vdd.n2578 10.6151
R17850 vdd.n2580 vdd.n2579 10.6151
R17851 vdd.n2580 vdd.n730 10.6151
R17852 vdd.n2590 vdd.n730 10.6151
R17853 vdd.n2591 vdd.n2590 10.6151
R17854 vdd.n2592 vdd.n2591 10.6151
R17855 vdd.n2592 vdd.n717 10.6151
R17856 vdd.n2602 vdd.n717 10.6151
R17857 vdd.n2603 vdd.n2602 10.6151
R17858 vdd.n2604 vdd.n2603 10.6151
R17859 vdd.n2604 vdd.n706 10.6151
R17860 vdd.n2614 vdd.n706 10.6151
R17861 vdd.n2615 vdd.n2614 10.6151
R17862 vdd.n2616 vdd.n2615 10.6151
R17863 vdd.n2616 vdd.n694 10.6151
R17864 vdd.n2626 vdd.n694 10.6151
R17865 vdd.n2627 vdd.n2626 10.6151
R17866 vdd.n2628 vdd.n2627 10.6151
R17867 vdd.n2628 vdd.n683 10.6151
R17868 vdd.n2640 vdd.n683 10.6151
R17869 vdd.n2641 vdd.n2640 10.6151
R17870 vdd.n2642 vdd.n2641 10.6151
R17871 vdd.n2642 vdd.n669 10.6151
R17872 vdd.n2697 vdd.n669 10.6151
R17873 vdd.n2698 vdd.n2697 10.6151
R17874 vdd.n2699 vdd.n2698 10.6151
R17875 vdd.n2699 vdd.n636 10.6151
R17876 vdd.n2769 vdd.n636 10.6151
R17877 vdd.n2768 vdd.n2767 10.6151
R17878 vdd.n2767 vdd.n637 10.6151
R17879 vdd.n638 vdd.n637 10.6151
R17880 vdd.n2760 vdd.n638 10.6151
R17881 vdd.n2760 vdd.n2759 10.6151
R17882 vdd.n2759 vdd.n2758 10.6151
R17883 vdd.n2758 vdd.n640 10.6151
R17884 vdd.n2753 vdd.n640 10.6151
R17885 vdd.n2753 vdd.n2752 10.6151
R17886 vdd.n2752 vdd.n2751 10.6151
R17887 vdd.n2751 vdd.n643 10.6151
R17888 vdd.n2746 vdd.n643 10.6151
R17889 vdd.n2746 vdd.n2745 10.6151
R17890 vdd.n2745 vdd.n2744 10.6151
R17891 vdd.n2744 vdd.n646 10.6151
R17892 vdd.n2739 vdd.n646 10.6151
R17893 vdd.n2739 vdd.n2738 10.6151
R17894 vdd.n2738 vdd.n2736 10.6151
R17895 vdd.n2736 vdd.n649 10.6151
R17896 vdd.n2731 vdd.n649 10.6151
R17897 vdd.n2731 vdd.n2730 10.6151
R17898 vdd.n2730 vdd.n2729 10.6151
R17899 vdd.n2729 vdd.n652 10.6151
R17900 vdd.n2724 vdd.n652 10.6151
R17901 vdd.n2724 vdd.n2723 10.6151
R17902 vdd.n2723 vdd.n2722 10.6151
R17903 vdd.n2722 vdd.n655 10.6151
R17904 vdd.n2717 vdd.n655 10.6151
R17905 vdd.n2717 vdd.n2716 10.6151
R17906 vdd.n2716 vdd.n2715 10.6151
R17907 vdd.n2715 vdd.n658 10.6151
R17908 vdd.n2710 vdd.n2709 10.6151
R17909 vdd.n2709 vdd.n2708 10.6151
R17910 vdd.n2687 vdd.n2648 10.6151
R17911 vdd.n2682 vdd.n2648 10.6151
R17912 vdd.n2682 vdd.n2681 10.6151
R17913 vdd.n2681 vdd.n2680 10.6151
R17914 vdd.n2680 vdd.n2650 10.6151
R17915 vdd.n2675 vdd.n2650 10.6151
R17916 vdd.n2675 vdd.n2674 10.6151
R17917 vdd.n2674 vdd.n2673 10.6151
R17918 vdd.n2673 vdd.n2653 10.6151
R17919 vdd.n2668 vdd.n2653 10.6151
R17920 vdd.n2668 vdd.n2667 10.6151
R17921 vdd.n2667 vdd.n2666 10.6151
R17922 vdd.n2666 vdd.n2656 10.6151
R17923 vdd.n2661 vdd.n2656 10.6151
R17924 vdd.n2661 vdd.n2660 10.6151
R17925 vdd.n2660 vdd.n610 10.6151
R17926 vdd.n2804 vdd.n610 10.6151
R17927 vdd.n2804 vdd.n611 10.6151
R17928 vdd.n614 vdd.n611 10.6151
R17929 vdd.n2797 vdd.n614 10.6151
R17930 vdd.n2797 vdd.n2796 10.6151
R17931 vdd.n2796 vdd.n2795 10.6151
R17932 vdd.n2795 vdd.n616 10.6151
R17933 vdd.n2790 vdd.n616 10.6151
R17934 vdd.n2790 vdd.n2789 10.6151
R17935 vdd.n2789 vdd.n2788 10.6151
R17936 vdd.n2788 vdd.n619 10.6151
R17937 vdd.n2783 vdd.n619 10.6151
R17938 vdd.n2783 vdd.n2782 10.6151
R17939 vdd.n2782 vdd.n2781 10.6151
R17940 vdd.n2781 vdd.n622 10.6151
R17941 vdd.n2776 vdd.n2775 10.6151
R17942 vdd.n2775 vdd.n2774 10.6151
R17943 vdd.n2422 vdd.n2420 10.6151
R17944 vdd.n2423 vdd.n2422 10.6151
R17945 vdd.n2491 vdd.n2423 10.6151
R17946 vdd.n2491 vdd.n2490 10.6151
R17947 vdd.n2490 vdd.n2489 10.6151
R17948 vdd.n2489 vdd.n2487 10.6151
R17949 vdd.n2487 vdd.n2486 10.6151
R17950 vdd.n2486 vdd.n2484 10.6151
R17951 vdd.n2484 vdd.n2483 10.6151
R17952 vdd.n2483 vdd.n2481 10.6151
R17953 vdd.n2481 vdd.n2480 10.6151
R17954 vdd.n2480 vdd.n2478 10.6151
R17955 vdd.n2478 vdd.n2477 10.6151
R17956 vdd.n2477 vdd.n2475 10.6151
R17957 vdd.n2475 vdd.n2474 10.6151
R17958 vdd.n2474 vdd.n2440 10.6151
R17959 vdd.n2440 vdd.n2439 10.6151
R17960 vdd.n2439 vdd.n2437 10.6151
R17961 vdd.n2437 vdd.n2436 10.6151
R17962 vdd.n2436 vdd.n2434 10.6151
R17963 vdd.n2434 vdd.n2433 10.6151
R17964 vdd.n2433 vdd.n2431 10.6151
R17965 vdd.n2431 vdd.n2430 10.6151
R17966 vdd.n2430 vdd.n2428 10.6151
R17967 vdd.n2428 vdd.n2427 10.6151
R17968 vdd.n2427 vdd.n2425 10.6151
R17969 vdd.n2425 vdd.n2424 10.6151
R17970 vdd.n2424 vdd.n628 10.6151
R17971 vdd.n2573 vdd.n2572 10.6151
R17972 vdd.n2572 vdd.n745 10.6151
R17973 vdd.n2357 vdd.n745 10.6151
R17974 vdd.n2360 vdd.n2357 10.6151
R17975 vdd.n2361 vdd.n2360 10.6151
R17976 vdd.n2364 vdd.n2361 10.6151
R17977 vdd.n2365 vdd.n2364 10.6151
R17978 vdd.n2368 vdd.n2365 10.6151
R17979 vdd.n2369 vdd.n2368 10.6151
R17980 vdd.n2372 vdd.n2369 10.6151
R17981 vdd.n2373 vdd.n2372 10.6151
R17982 vdd.n2376 vdd.n2373 10.6151
R17983 vdd.n2377 vdd.n2376 10.6151
R17984 vdd.n2380 vdd.n2377 10.6151
R17985 vdd.n2381 vdd.n2380 10.6151
R17986 vdd.n2384 vdd.n2381 10.6151
R17987 vdd.n2385 vdd.n2384 10.6151
R17988 vdd.n2388 vdd.n2385 10.6151
R17989 vdd.n2389 vdd.n2388 10.6151
R17990 vdd.n2392 vdd.n2389 10.6151
R17991 vdd.n2393 vdd.n2392 10.6151
R17992 vdd.n2396 vdd.n2393 10.6151
R17993 vdd.n2397 vdd.n2396 10.6151
R17994 vdd.n2400 vdd.n2397 10.6151
R17995 vdd.n2401 vdd.n2400 10.6151
R17996 vdd.n2404 vdd.n2401 10.6151
R17997 vdd.n2405 vdd.n2404 10.6151
R17998 vdd.n2408 vdd.n2405 10.6151
R17999 vdd.n2409 vdd.n2408 10.6151
R18000 vdd.n2412 vdd.n2409 10.6151
R18001 vdd.n2413 vdd.n2412 10.6151
R18002 vdd.n2418 vdd.n2416 10.6151
R18003 vdd.n2419 vdd.n2418 10.6151
R18004 vdd.n2574 vdd.n735 10.6151
R18005 vdd.n2584 vdd.n735 10.6151
R18006 vdd.n2585 vdd.n2584 10.6151
R18007 vdd.n2586 vdd.n2585 10.6151
R18008 vdd.n2586 vdd.n723 10.6151
R18009 vdd.n2596 vdd.n723 10.6151
R18010 vdd.n2597 vdd.n2596 10.6151
R18011 vdd.n2598 vdd.n2597 10.6151
R18012 vdd.n2598 vdd.n712 10.6151
R18013 vdd.n2608 vdd.n712 10.6151
R18014 vdd.n2609 vdd.n2608 10.6151
R18015 vdd.n2610 vdd.n2609 10.6151
R18016 vdd.n2610 vdd.n700 10.6151
R18017 vdd.n2620 vdd.n700 10.6151
R18018 vdd.n2621 vdd.n2620 10.6151
R18019 vdd.n2622 vdd.n2621 10.6151
R18020 vdd.n2622 vdd.n689 10.6151
R18021 vdd.n2632 vdd.n689 10.6151
R18022 vdd.n2633 vdd.n2632 10.6151
R18023 vdd.n2636 vdd.n2633 10.6151
R18024 vdd.n2646 vdd.n677 10.6151
R18025 vdd.n2647 vdd.n2646 10.6151
R18026 vdd.n2693 vdd.n2647 10.6151
R18027 vdd.n2693 vdd.n2692 10.6151
R18028 vdd.n2692 vdd.n2691 10.6151
R18029 vdd.n2691 vdd.n2690 10.6151
R18030 vdd.n2690 vdd.n2688 10.6151
R18031 vdd.n2085 vdd.n869 10.6151
R18032 vdd.n2095 vdd.n869 10.6151
R18033 vdd.n2096 vdd.n2095 10.6151
R18034 vdd.n2097 vdd.n2096 10.6151
R18035 vdd.n2097 vdd.n856 10.6151
R18036 vdd.n2107 vdd.n856 10.6151
R18037 vdd.n2108 vdd.n2107 10.6151
R18038 vdd.n2110 vdd.n844 10.6151
R18039 vdd.n2120 vdd.n844 10.6151
R18040 vdd.n2121 vdd.n2120 10.6151
R18041 vdd.n2122 vdd.n2121 10.6151
R18042 vdd.n2122 vdd.n832 10.6151
R18043 vdd.n2132 vdd.n832 10.6151
R18044 vdd.n2133 vdd.n2132 10.6151
R18045 vdd.n2134 vdd.n2133 10.6151
R18046 vdd.n2134 vdd.n821 10.6151
R18047 vdd.n2144 vdd.n821 10.6151
R18048 vdd.n2145 vdd.n2144 10.6151
R18049 vdd.n2146 vdd.n2145 10.6151
R18050 vdd.n2146 vdd.n809 10.6151
R18051 vdd.n2156 vdd.n809 10.6151
R18052 vdd.n2157 vdd.n2156 10.6151
R18053 vdd.n2160 vdd.n2157 10.6151
R18054 vdd.n2160 vdd.n2159 10.6151
R18055 vdd.n2159 vdd.n2158 10.6151
R18056 vdd.n2158 vdd.n792 10.6151
R18057 vdd.n2242 vdd.n792 10.6151
R18058 vdd.n2241 vdd.n2240 10.6151
R18059 vdd.n2240 vdd.n2237 10.6151
R18060 vdd.n2237 vdd.n2236 10.6151
R18061 vdd.n2236 vdd.n2233 10.6151
R18062 vdd.n2233 vdd.n2232 10.6151
R18063 vdd.n2232 vdd.n2229 10.6151
R18064 vdd.n2229 vdd.n2228 10.6151
R18065 vdd.n2228 vdd.n2225 10.6151
R18066 vdd.n2225 vdd.n2224 10.6151
R18067 vdd.n2224 vdd.n2221 10.6151
R18068 vdd.n2221 vdd.n2220 10.6151
R18069 vdd.n2220 vdd.n2217 10.6151
R18070 vdd.n2217 vdd.n2216 10.6151
R18071 vdd.n2216 vdd.n2213 10.6151
R18072 vdd.n2213 vdd.n2212 10.6151
R18073 vdd.n2212 vdd.n2209 10.6151
R18074 vdd.n2209 vdd.n2208 10.6151
R18075 vdd.n2208 vdd.n2205 10.6151
R18076 vdd.n2205 vdd.n2204 10.6151
R18077 vdd.n2204 vdd.n2201 10.6151
R18078 vdd.n2201 vdd.n2200 10.6151
R18079 vdd.n2200 vdd.n2197 10.6151
R18080 vdd.n2197 vdd.n2196 10.6151
R18081 vdd.n2196 vdd.n2193 10.6151
R18082 vdd.n2193 vdd.n2192 10.6151
R18083 vdd.n2192 vdd.n2189 10.6151
R18084 vdd.n2189 vdd.n2188 10.6151
R18085 vdd.n2188 vdd.n2185 10.6151
R18086 vdd.n2185 vdd.n2184 10.6151
R18087 vdd.n2184 vdd.n2181 10.6151
R18088 vdd.n2181 vdd.n2180 10.6151
R18089 vdd.n2177 vdd.n2176 10.6151
R18090 vdd.n2176 vdd.n2174 10.6151
R18091 vdd.n1933 vdd.n1931 10.6151
R18092 vdd.n1934 vdd.n1933 10.6151
R18093 vdd.n1936 vdd.n1934 10.6151
R18094 vdd.n1937 vdd.n1936 10.6151
R18095 vdd.n1939 vdd.n1937 10.6151
R18096 vdd.n1940 vdd.n1939 10.6151
R18097 vdd.n1942 vdd.n1940 10.6151
R18098 vdd.n1943 vdd.n1942 10.6151
R18099 vdd.n1945 vdd.n1943 10.6151
R18100 vdd.n1946 vdd.n1945 10.6151
R18101 vdd.n1948 vdd.n1946 10.6151
R18102 vdd.n1949 vdd.n1948 10.6151
R18103 vdd.n1967 vdd.n1949 10.6151
R18104 vdd.n1967 vdd.n1966 10.6151
R18105 vdd.n1966 vdd.n1965 10.6151
R18106 vdd.n1965 vdd.n1963 10.6151
R18107 vdd.n1963 vdd.n1962 10.6151
R18108 vdd.n1962 vdd.n1960 10.6151
R18109 vdd.n1960 vdd.n1959 10.6151
R18110 vdd.n1959 vdd.n1957 10.6151
R18111 vdd.n1957 vdd.n1956 10.6151
R18112 vdd.n1956 vdd.n1954 10.6151
R18113 vdd.n1954 vdd.n1953 10.6151
R18114 vdd.n1953 vdd.n1951 10.6151
R18115 vdd.n1951 vdd.n1950 10.6151
R18116 vdd.n1950 vdd.n796 10.6151
R18117 vdd.n2172 vdd.n796 10.6151
R18118 vdd.n2173 vdd.n2172 10.6151
R18119 vdd.n2084 vdd.n2083 10.6151
R18120 vdd.n2083 vdd.n881 10.6151
R18121 vdd.n2077 vdd.n881 10.6151
R18122 vdd.n2077 vdd.n2076 10.6151
R18123 vdd.n2076 vdd.n2075 10.6151
R18124 vdd.n2075 vdd.n883 10.6151
R18125 vdd.n2069 vdd.n883 10.6151
R18126 vdd.n2069 vdd.n2068 10.6151
R18127 vdd.n2068 vdd.n2067 10.6151
R18128 vdd.n2067 vdd.n885 10.6151
R18129 vdd.n2061 vdd.n885 10.6151
R18130 vdd.n2061 vdd.n2060 10.6151
R18131 vdd.n2060 vdd.n2059 10.6151
R18132 vdd.n2059 vdd.n887 10.6151
R18133 vdd.n2053 vdd.n887 10.6151
R18134 vdd.n2053 vdd.n2052 10.6151
R18135 vdd.n2052 vdd.n2051 10.6151
R18136 vdd.n2051 vdd.n891 10.6151
R18137 vdd.n1899 vdd.n891 10.6151
R18138 vdd.n1900 vdd.n1899 10.6151
R18139 vdd.n1900 vdd.n1895 10.6151
R18140 vdd.n1906 vdd.n1895 10.6151
R18141 vdd.n1907 vdd.n1906 10.6151
R18142 vdd.n1908 vdd.n1907 10.6151
R18143 vdd.n1908 vdd.n1893 10.6151
R18144 vdd.n1914 vdd.n1893 10.6151
R18145 vdd.n1915 vdd.n1914 10.6151
R18146 vdd.n1916 vdd.n1915 10.6151
R18147 vdd.n1916 vdd.n1891 10.6151
R18148 vdd.n1922 vdd.n1891 10.6151
R18149 vdd.n1923 vdd.n1922 10.6151
R18150 vdd.n1925 vdd.n1887 10.6151
R18151 vdd.n1930 vdd.n1887 10.6151
R18152 vdd.n1272 vdd.t178 10.5435
R18153 vdd.n2041 vdd.t62 10.5435
R18154 vdd.n2940 vdd.t55 10.5435
R18155 vdd.n3164 vdd.t35 10.5435
R18156 vdd.n292 vdd.n274 10.4732
R18157 vdd.n241 vdd.n223 10.4732
R18158 vdd.n198 vdd.n180 10.4732
R18159 vdd.n147 vdd.n129 10.4732
R18160 vdd.n105 vdd.n87 10.4732
R18161 vdd.n54 vdd.n36 10.4732
R18162 vdd.n1487 vdd.n1469 10.4732
R18163 vdd.n1538 vdd.n1520 10.4732
R18164 vdd.n1393 vdd.n1375 10.4732
R18165 vdd.n1444 vdd.n1426 10.4732
R18166 vdd.n1300 vdd.n1282 10.4732
R18167 vdd.n1351 vdd.n1333 10.4732
R18168 vdd.n1570 vdd.t4 10.3167
R18169 vdd.t28 vdd.n493 10.3167
R18170 vdd.n1223 vdd.t66 9.86327
R18171 vdd.n3140 vdd.t115 9.86327
R18172 vdd.n291 vdd.n276 9.69747
R18173 vdd.n240 vdd.n225 9.69747
R18174 vdd.n197 vdd.n182 9.69747
R18175 vdd.n146 vdd.n131 9.69747
R18176 vdd.n104 vdd.n89 9.69747
R18177 vdd.n53 vdd.n38 9.69747
R18178 vdd.n1486 vdd.n1471 9.69747
R18179 vdd.n1537 vdd.n1522 9.69747
R18180 vdd.n1392 vdd.n1377 9.69747
R18181 vdd.n1443 vdd.n1428 9.69747
R18182 vdd.n1299 vdd.n1284 9.69747
R18183 vdd.n1350 vdd.n1335 9.69747
R18184 vdd.n2027 vdd.n2026 9.67831
R18185 vdd.n2738 vdd.n2737 9.67831
R18186 vdd.n2805 vdd.n2804 9.67831
R18187 vdd.n2051 vdd.n2050 9.67831
R18188 vdd.n307 vdd.n306 9.45567
R18189 vdd.n256 vdd.n255 9.45567
R18190 vdd.n213 vdd.n212 9.45567
R18191 vdd.n162 vdd.n161 9.45567
R18192 vdd.n120 vdd.n119 9.45567
R18193 vdd.n69 vdd.n68 9.45567
R18194 vdd.n1502 vdd.n1501 9.45567
R18195 vdd.n1553 vdd.n1552 9.45567
R18196 vdd.n1408 vdd.n1407 9.45567
R18197 vdd.n1459 vdd.n1458 9.45567
R18198 vdd.n1315 vdd.n1314 9.45567
R18199 vdd.n1366 vdd.n1365 9.45567
R18200 vdd.n1787 vdd.n1641 9.3005
R18201 vdd.n1786 vdd.n1785 9.3005
R18202 vdd.n1647 vdd.n1646 9.3005
R18203 vdd.n1780 vdd.n1651 9.3005
R18204 vdd.n1779 vdd.n1652 9.3005
R18205 vdd.n1778 vdd.n1653 9.3005
R18206 vdd.n1657 vdd.n1654 9.3005
R18207 vdd.n1773 vdd.n1658 9.3005
R18208 vdd.n1772 vdd.n1659 9.3005
R18209 vdd.n1771 vdd.n1660 9.3005
R18210 vdd.n1664 vdd.n1661 9.3005
R18211 vdd.n1766 vdd.n1665 9.3005
R18212 vdd.n1765 vdd.n1666 9.3005
R18213 vdd.n1764 vdd.n1667 9.3005
R18214 vdd.n1671 vdd.n1668 9.3005
R18215 vdd.n1759 vdd.n1672 9.3005
R18216 vdd.n1758 vdd.n1673 9.3005
R18217 vdd.n1757 vdd.n1674 9.3005
R18218 vdd.n1678 vdd.n1675 9.3005
R18219 vdd.n1752 vdd.n1679 9.3005
R18220 vdd.n1751 vdd.n1680 9.3005
R18221 vdd.n1750 vdd.n1749 9.3005
R18222 vdd.n1748 vdd.n1681 9.3005
R18223 vdd.n1747 vdd.n1746 9.3005
R18224 vdd.n1687 vdd.n1686 9.3005
R18225 vdd.n1741 vdd.n1691 9.3005
R18226 vdd.n1740 vdd.n1692 9.3005
R18227 vdd.n1739 vdd.n1693 9.3005
R18228 vdd.n1697 vdd.n1694 9.3005
R18229 vdd.n1734 vdd.n1698 9.3005
R18230 vdd.n1733 vdd.n1699 9.3005
R18231 vdd.n1732 vdd.n1700 9.3005
R18232 vdd.n1704 vdd.n1701 9.3005
R18233 vdd.n1727 vdd.n1705 9.3005
R18234 vdd.n1726 vdd.n1706 9.3005
R18235 vdd.n1725 vdd.n1707 9.3005
R18236 vdd.n1709 vdd.n1708 9.3005
R18237 vdd.n1720 vdd.n892 9.3005
R18238 vdd.n1789 vdd.n1788 9.3005
R18239 vdd.n1813 vdd.n1812 9.3005
R18240 vdd.n1619 vdd.n1618 9.3005
R18241 vdd.n1624 vdd.n1622 9.3005
R18242 vdd.n1805 vdd.n1625 9.3005
R18243 vdd.n1804 vdd.n1626 9.3005
R18244 vdd.n1803 vdd.n1627 9.3005
R18245 vdd.n1631 vdd.n1628 9.3005
R18246 vdd.n1798 vdd.n1632 9.3005
R18247 vdd.n1797 vdd.n1633 9.3005
R18248 vdd.n1796 vdd.n1634 9.3005
R18249 vdd.n1638 vdd.n1635 9.3005
R18250 vdd.n1791 vdd.n1639 9.3005
R18251 vdd.n1790 vdd.n1640 9.3005
R18252 vdd.n2035 vdd.n1612 9.3005
R18253 vdd.n2037 vdd.n2036 9.3005
R18254 vdd.n1558 vdd.n939 9.3005
R18255 vdd.n1560 vdd.n1559 9.3005
R18256 vdd.n929 vdd.n928 9.3005
R18257 vdd.n1574 vdd.n1573 9.3005
R18258 vdd.n1575 vdd.n927 9.3005
R18259 vdd.n1577 vdd.n1576 9.3005
R18260 vdd.n918 vdd.n917 9.3005
R18261 vdd.n1591 vdd.n1590 9.3005
R18262 vdd.n1592 vdd.n916 9.3005
R18263 vdd.n1594 vdd.n1593 9.3005
R18264 vdd.n906 vdd.n905 9.3005
R18265 vdd.n1610 vdd.n1609 9.3005
R18266 vdd.n1611 vdd.n904 9.3005
R18267 vdd.n2039 vdd.n2038 9.3005
R18268 vdd.n283 vdd.n282 9.3005
R18269 vdd.n278 vdd.n277 9.3005
R18270 vdd.n289 vdd.n288 9.3005
R18271 vdd.n291 vdd.n290 9.3005
R18272 vdd.n274 vdd.n273 9.3005
R18273 vdd.n297 vdd.n296 9.3005
R18274 vdd.n299 vdd.n298 9.3005
R18275 vdd.n271 vdd.n268 9.3005
R18276 vdd.n306 vdd.n305 9.3005
R18277 vdd.n232 vdd.n231 9.3005
R18278 vdd.n227 vdd.n226 9.3005
R18279 vdd.n238 vdd.n237 9.3005
R18280 vdd.n240 vdd.n239 9.3005
R18281 vdd.n223 vdd.n222 9.3005
R18282 vdd.n246 vdd.n245 9.3005
R18283 vdd.n248 vdd.n247 9.3005
R18284 vdd.n220 vdd.n217 9.3005
R18285 vdd.n255 vdd.n254 9.3005
R18286 vdd.n189 vdd.n188 9.3005
R18287 vdd.n184 vdd.n183 9.3005
R18288 vdd.n195 vdd.n194 9.3005
R18289 vdd.n197 vdd.n196 9.3005
R18290 vdd.n180 vdd.n179 9.3005
R18291 vdd.n203 vdd.n202 9.3005
R18292 vdd.n205 vdd.n204 9.3005
R18293 vdd.n177 vdd.n174 9.3005
R18294 vdd.n212 vdd.n211 9.3005
R18295 vdd.n138 vdd.n137 9.3005
R18296 vdd.n133 vdd.n132 9.3005
R18297 vdd.n144 vdd.n143 9.3005
R18298 vdd.n146 vdd.n145 9.3005
R18299 vdd.n129 vdd.n128 9.3005
R18300 vdd.n152 vdd.n151 9.3005
R18301 vdd.n154 vdd.n153 9.3005
R18302 vdd.n126 vdd.n123 9.3005
R18303 vdd.n161 vdd.n160 9.3005
R18304 vdd.n96 vdd.n95 9.3005
R18305 vdd.n91 vdd.n90 9.3005
R18306 vdd.n102 vdd.n101 9.3005
R18307 vdd.n104 vdd.n103 9.3005
R18308 vdd.n87 vdd.n86 9.3005
R18309 vdd.n110 vdd.n109 9.3005
R18310 vdd.n112 vdd.n111 9.3005
R18311 vdd.n84 vdd.n81 9.3005
R18312 vdd.n119 vdd.n118 9.3005
R18313 vdd.n45 vdd.n44 9.3005
R18314 vdd.n40 vdd.n39 9.3005
R18315 vdd.n51 vdd.n50 9.3005
R18316 vdd.n53 vdd.n52 9.3005
R18317 vdd.n36 vdd.n35 9.3005
R18318 vdd.n59 vdd.n58 9.3005
R18319 vdd.n61 vdd.n60 9.3005
R18320 vdd.n33 vdd.n30 9.3005
R18321 vdd.n68 vdd.n67 9.3005
R18322 vdd.n2854 vdd.n2853 9.3005
R18323 vdd.n2855 vdd.n578 9.3005
R18324 vdd.n577 vdd.n575 9.3005
R18325 vdd.n2861 vdd.n574 9.3005
R18326 vdd.n2862 vdd.n573 9.3005
R18327 vdd.n2863 vdd.n572 9.3005
R18328 vdd.n571 vdd.n569 9.3005
R18329 vdd.n2869 vdd.n568 9.3005
R18330 vdd.n2870 vdd.n567 9.3005
R18331 vdd.n2871 vdd.n566 9.3005
R18332 vdd.n565 vdd.n563 9.3005
R18333 vdd.n2877 vdd.n562 9.3005
R18334 vdd.n2878 vdd.n561 9.3005
R18335 vdd.n2879 vdd.n560 9.3005
R18336 vdd.n559 vdd.n557 9.3005
R18337 vdd.n2885 vdd.n556 9.3005
R18338 vdd.n2886 vdd.n555 9.3005
R18339 vdd.n2887 vdd.n554 9.3005
R18340 vdd.n553 vdd.n551 9.3005
R18341 vdd.n2893 vdd.n550 9.3005
R18342 vdd.n2894 vdd.n549 9.3005
R18343 vdd.n2895 vdd.n548 9.3005
R18344 vdd.n547 vdd.n545 9.3005
R18345 vdd.n2901 vdd.n542 9.3005
R18346 vdd.n2902 vdd.n541 9.3005
R18347 vdd.n2903 vdd.n540 9.3005
R18348 vdd.n539 vdd.n537 9.3005
R18349 vdd.n2909 vdd.n536 9.3005
R18350 vdd.n2910 vdd.n535 9.3005
R18351 vdd.n2911 vdd.n534 9.3005
R18352 vdd.n533 vdd.n531 9.3005
R18353 vdd.n2917 vdd.n530 9.3005
R18354 vdd.n2918 vdd.n529 9.3005
R18355 vdd.n2919 vdd.n528 9.3005
R18356 vdd.n527 vdd.n525 9.3005
R18357 vdd.n2924 vdd.n524 9.3005
R18358 vdd.n2934 vdd.n518 9.3005
R18359 vdd.n2936 vdd.n2935 9.3005
R18360 vdd.n509 vdd.n508 9.3005
R18361 vdd.n2951 vdd.n2950 9.3005
R18362 vdd.n2952 vdd.n507 9.3005
R18363 vdd.n2954 vdd.n2953 9.3005
R18364 vdd.n497 vdd.n496 9.3005
R18365 vdd.n2967 vdd.n2966 9.3005
R18366 vdd.n2968 vdd.n495 9.3005
R18367 vdd.n2970 vdd.n2969 9.3005
R18368 vdd.n485 vdd.n484 9.3005
R18369 vdd.n2984 vdd.n2983 9.3005
R18370 vdd.n2985 vdd.n483 9.3005
R18371 vdd.n2987 vdd.n2986 9.3005
R18372 vdd.n312 vdd.n310 9.3005
R18373 vdd.n2938 vdd.n2937 9.3005
R18374 vdd.n3167 vdd.n3166 9.3005
R18375 vdd.n313 vdd.n311 9.3005
R18376 vdd.n3160 vdd.n320 9.3005
R18377 vdd.n3159 vdd.n321 9.3005
R18378 vdd.n3158 vdd.n322 9.3005
R18379 vdd.n331 vdd.n323 9.3005
R18380 vdd.n3152 vdd.n332 9.3005
R18381 vdd.n3151 vdd.n333 9.3005
R18382 vdd.n3150 vdd.n334 9.3005
R18383 vdd.n342 vdd.n335 9.3005
R18384 vdd.n3144 vdd.n343 9.3005
R18385 vdd.n3143 vdd.n344 9.3005
R18386 vdd.n3142 vdd.n345 9.3005
R18387 vdd.n353 vdd.n346 9.3005
R18388 vdd.n3136 vdd.n3135 9.3005
R18389 vdd.n3132 vdd.n354 9.3005
R18390 vdd.n3131 vdd.n357 9.3005
R18391 vdd.n361 vdd.n358 9.3005
R18392 vdd.n362 vdd.n359 9.3005
R18393 vdd.n3124 vdd.n363 9.3005
R18394 vdd.n3123 vdd.n364 9.3005
R18395 vdd.n3122 vdd.n365 9.3005
R18396 vdd.n369 vdd.n366 9.3005
R18397 vdd.n3117 vdd.n370 9.3005
R18398 vdd.n3116 vdd.n371 9.3005
R18399 vdd.n3115 vdd.n372 9.3005
R18400 vdd.n376 vdd.n373 9.3005
R18401 vdd.n3110 vdd.n377 9.3005
R18402 vdd.n3109 vdd.n378 9.3005
R18403 vdd.n3108 vdd.n379 9.3005
R18404 vdd.n383 vdd.n380 9.3005
R18405 vdd.n3103 vdd.n384 9.3005
R18406 vdd.n3102 vdd.n385 9.3005
R18407 vdd.n3101 vdd.n3100 9.3005
R18408 vdd.n3099 vdd.n386 9.3005
R18409 vdd.n3098 vdd.n3097 9.3005
R18410 vdd.n392 vdd.n391 9.3005
R18411 vdd.n3092 vdd.n396 9.3005
R18412 vdd.n3091 vdd.n397 9.3005
R18413 vdd.n3090 vdd.n398 9.3005
R18414 vdd.n402 vdd.n399 9.3005
R18415 vdd.n3085 vdd.n403 9.3005
R18416 vdd.n3084 vdd.n404 9.3005
R18417 vdd.n3083 vdd.n405 9.3005
R18418 vdd.n409 vdd.n406 9.3005
R18419 vdd.n3078 vdd.n410 9.3005
R18420 vdd.n3077 vdd.n411 9.3005
R18421 vdd.n3076 vdd.n412 9.3005
R18422 vdd.n416 vdd.n413 9.3005
R18423 vdd.n3071 vdd.n417 9.3005
R18424 vdd.n3070 vdd.n418 9.3005
R18425 vdd.n3069 vdd.n419 9.3005
R18426 vdd.n423 vdd.n420 9.3005
R18427 vdd.n3064 vdd.n424 9.3005
R18428 vdd.n3063 vdd.n425 9.3005
R18429 vdd.n3062 vdd.n3061 9.3005
R18430 vdd.n3060 vdd.n426 9.3005
R18431 vdd.n3059 vdd.n3058 9.3005
R18432 vdd.n432 vdd.n431 9.3005
R18433 vdd.n3053 vdd.n436 9.3005
R18434 vdd.n3052 vdd.n437 9.3005
R18435 vdd.n3051 vdd.n438 9.3005
R18436 vdd.n442 vdd.n439 9.3005
R18437 vdd.n3046 vdd.n443 9.3005
R18438 vdd.n3045 vdd.n444 9.3005
R18439 vdd.n3044 vdd.n445 9.3005
R18440 vdd.n449 vdd.n446 9.3005
R18441 vdd.n3039 vdd.n450 9.3005
R18442 vdd.n3038 vdd.n451 9.3005
R18443 vdd.n3037 vdd.n452 9.3005
R18444 vdd.n456 vdd.n453 9.3005
R18445 vdd.n3032 vdd.n457 9.3005
R18446 vdd.n3031 vdd.n458 9.3005
R18447 vdd.n3030 vdd.n459 9.3005
R18448 vdd.n463 vdd.n460 9.3005
R18449 vdd.n3025 vdd.n464 9.3005
R18450 vdd.n3024 vdd.n465 9.3005
R18451 vdd.n3020 vdd.n3017 9.3005
R18452 vdd.n3134 vdd.n3133 9.3005
R18453 vdd.n2944 vdd.n513 9.3005
R18454 vdd.n2946 vdd.n2945 9.3005
R18455 vdd.n503 vdd.n502 9.3005
R18456 vdd.n2959 vdd.n2958 9.3005
R18457 vdd.n2960 vdd.n501 9.3005
R18458 vdd.n2962 vdd.n2961 9.3005
R18459 vdd.n490 vdd.n489 9.3005
R18460 vdd.n2975 vdd.n2974 9.3005
R18461 vdd.n2976 vdd.n488 9.3005
R18462 vdd.n2978 vdd.n2977 9.3005
R18463 vdd.n478 vdd.n477 9.3005
R18464 vdd.n2992 vdd.n2991 9.3005
R18465 vdd.n2993 vdd.n476 9.3005
R18466 vdd.n2995 vdd.n2994 9.3005
R18467 vdd.n2996 vdd.n475 9.3005
R18468 vdd.n2998 vdd.n2997 9.3005
R18469 vdd.n2999 vdd.n474 9.3005
R18470 vdd.n3001 vdd.n3000 9.3005
R18471 vdd.n3002 vdd.n472 9.3005
R18472 vdd.n3004 vdd.n3003 9.3005
R18473 vdd.n3005 vdd.n471 9.3005
R18474 vdd.n3007 vdd.n3006 9.3005
R18475 vdd.n3008 vdd.n469 9.3005
R18476 vdd.n3010 vdd.n3009 9.3005
R18477 vdd.n3011 vdd.n468 9.3005
R18478 vdd.n3013 vdd.n3012 9.3005
R18479 vdd.n3014 vdd.n466 9.3005
R18480 vdd.n3016 vdd.n3015 9.3005
R18481 vdd.n2943 vdd.n2942 9.3005
R18482 vdd.n2807 vdd.n514 9.3005
R18483 vdd.n2812 vdd.n2806 9.3005
R18484 vdd.n2822 vdd.n605 9.3005
R18485 vdd.n2823 vdd.n604 9.3005
R18486 vdd.n603 vdd.n601 9.3005
R18487 vdd.n2829 vdd.n600 9.3005
R18488 vdd.n2830 vdd.n599 9.3005
R18489 vdd.n2831 vdd.n598 9.3005
R18490 vdd.n597 vdd.n595 9.3005
R18491 vdd.n2837 vdd.n594 9.3005
R18492 vdd.n2838 vdd.n593 9.3005
R18493 vdd.n2839 vdd.n592 9.3005
R18494 vdd.n591 vdd.n589 9.3005
R18495 vdd.n2844 vdd.n588 9.3005
R18496 vdd.n2845 vdd.n587 9.3005
R18497 vdd.n583 vdd.n582 9.3005
R18498 vdd.n2851 vdd.n2850 9.3005
R18499 vdd.n2852 vdd.n579 9.3005
R18500 vdd.n2049 vdd.n2048 9.3005
R18501 vdd.n2044 vdd.n895 9.3005
R18502 vdd.n1219 vdd.n979 9.3005
R18503 vdd.n1221 vdd.n1220 9.3005
R18504 vdd.n970 vdd.n969 9.3005
R18505 vdd.n1234 vdd.n1233 9.3005
R18506 vdd.n1235 vdd.n968 9.3005
R18507 vdd.n1237 vdd.n1236 9.3005
R18508 vdd.n957 vdd.n956 9.3005
R18509 vdd.n1250 vdd.n1249 9.3005
R18510 vdd.n1251 vdd.n955 9.3005
R18511 vdd.n1253 vdd.n1252 9.3005
R18512 vdd.n946 vdd.n945 9.3005
R18513 vdd.n1267 vdd.n1266 9.3005
R18514 vdd.n1268 vdd.n944 9.3005
R18515 vdd.n1270 vdd.n1269 9.3005
R18516 vdd.n935 vdd.n934 9.3005
R18517 vdd.n1565 vdd.n1564 9.3005
R18518 vdd.n1566 vdd.n933 9.3005
R18519 vdd.n1568 vdd.n1567 9.3005
R18520 vdd.n923 vdd.n922 9.3005
R18521 vdd.n1582 vdd.n1581 9.3005
R18522 vdd.n1583 vdd.n921 9.3005
R18523 vdd.n1585 vdd.n1584 9.3005
R18524 vdd.n913 vdd.n912 9.3005
R18525 vdd.n1599 vdd.n1598 9.3005
R18526 vdd.n1600 vdd.n910 9.3005
R18527 vdd.n1604 vdd.n1603 9.3005
R18528 vdd.n1602 vdd.n911 9.3005
R18529 vdd.n1601 vdd.n900 9.3005
R18530 vdd.n1218 vdd.n1217 9.3005
R18531 vdd.n1113 vdd.n1103 9.3005
R18532 vdd.n1115 vdd.n1114 9.3005
R18533 vdd.n1116 vdd.n1102 9.3005
R18534 vdd.n1118 vdd.n1117 9.3005
R18535 vdd.n1119 vdd.n1095 9.3005
R18536 vdd.n1121 vdd.n1120 9.3005
R18537 vdd.n1122 vdd.n1094 9.3005
R18538 vdd.n1124 vdd.n1123 9.3005
R18539 vdd.n1125 vdd.n1087 9.3005
R18540 vdd.n1127 vdd.n1126 9.3005
R18541 vdd.n1128 vdd.n1086 9.3005
R18542 vdd.n1130 vdd.n1129 9.3005
R18543 vdd.n1131 vdd.n1079 9.3005
R18544 vdd.n1133 vdd.n1132 9.3005
R18545 vdd.n1134 vdd.n1078 9.3005
R18546 vdd.n1136 vdd.n1135 9.3005
R18547 vdd.n1137 vdd.n1072 9.3005
R18548 vdd.n1139 vdd.n1138 9.3005
R18549 vdd.n1140 vdd.n1070 9.3005
R18550 vdd.n1142 vdd.n1141 9.3005
R18551 vdd.n1071 vdd.n1068 9.3005
R18552 vdd.n1149 vdd.n1064 9.3005
R18553 vdd.n1151 vdd.n1150 9.3005
R18554 vdd.n1152 vdd.n1063 9.3005
R18555 vdd.n1154 vdd.n1153 9.3005
R18556 vdd.n1155 vdd.n1056 9.3005
R18557 vdd.n1157 vdd.n1156 9.3005
R18558 vdd.n1158 vdd.n1055 9.3005
R18559 vdd.n1160 vdd.n1159 9.3005
R18560 vdd.n1161 vdd.n1048 9.3005
R18561 vdd.n1163 vdd.n1162 9.3005
R18562 vdd.n1164 vdd.n1047 9.3005
R18563 vdd.n1166 vdd.n1165 9.3005
R18564 vdd.n1167 vdd.n1040 9.3005
R18565 vdd.n1169 vdd.n1168 9.3005
R18566 vdd.n1170 vdd.n1039 9.3005
R18567 vdd.n1172 vdd.n1171 9.3005
R18568 vdd.n1173 vdd.n1032 9.3005
R18569 vdd.n1175 vdd.n1174 9.3005
R18570 vdd.n1176 vdd.n1031 9.3005
R18571 vdd.n1178 vdd.n1177 9.3005
R18572 vdd.n1179 vdd.n1024 9.3005
R18573 vdd.n1181 vdd.n1180 9.3005
R18574 vdd.n1182 vdd.n1023 9.3005
R18575 vdd.n1184 vdd.n1183 9.3005
R18576 vdd.n1185 vdd.n1014 9.3005
R18577 vdd.n1187 vdd.n1186 9.3005
R18578 vdd.n1188 vdd.n1013 9.3005
R18579 vdd.n1190 vdd.n1189 9.3005
R18580 vdd.n1191 vdd.n1006 9.3005
R18581 vdd.n1193 vdd.n1192 9.3005
R18582 vdd.n1194 vdd.n1005 9.3005
R18583 vdd.n1196 vdd.n1195 9.3005
R18584 vdd.n1197 vdd.n998 9.3005
R18585 vdd.n1199 vdd.n1198 9.3005
R18586 vdd.n1200 vdd.n997 9.3005
R18587 vdd.n1202 vdd.n1201 9.3005
R18588 vdd.n1203 vdd.n990 9.3005
R18589 vdd.n1205 vdd.n1204 9.3005
R18590 vdd.n1206 vdd.n989 9.3005
R18591 vdd.n1208 vdd.n1207 9.3005
R18592 vdd.n1209 vdd.n985 9.3005
R18593 vdd.n1211 vdd.n1210 9.3005
R18594 vdd.n1109 vdd.n980 9.3005
R18595 vdd.n976 vdd.n975 9.3005
R18596 vdd.n1226 vdd.n1225 9.3005
R18597 vdd.n1227 vdd.n974 9.3005
R18598 vdd.n1229 vdd.n1228 9.3005
R18599 vdd.n964 vdd.n963 9.3005
R18600 vdd.n1242 vdd.n1241 9.3005
R18601 vdd.n1243 vdd.n962 9.3005
R18602 vdd.n1245 vdd.n1244 9.3005
R18603 vdd.n952 vdd.n951 9.3005
R18604 vdd.n1259 vdd.n1258 9.3005
R18605 vdd.n1260 vdd.n950 9.3005
R18606 vdd.n1262 vdd.n1261 9.3005
R18607 vdd.n941 vdd.n940 9.3005
R18608 vdd.n1213 vdd.n1212 9.3005
R18609 vdd.n1557 vdd.n1274 9.3005
R18610 vdd.n1478 vdd.n1477 9.3005
R18611 vdd.n1473 vdd.n1472 9.3005
R18612 vdd.n1484 vdd.n1483 9.3005
R18613 vdd.n1486 vdd.n1485 9.3005
R18614 vdd.n1469 vdd.n1468 9.3005
R18615 vdd.n1492 vdd.n1491 9.3005
R18616 vdd.n1494 vdd.n1493 9.3005
R18617 vdd.n1466 vdd.n1463 9.3005
R18618 vdd.n1501 vdd.n1500 9.3005
R18619 vdd.n1529 vdd.n1528 9.3005
R18620 vdd.n1524 vdd.n1523 9.3005
R18621 vdd.n1535 vdd.n1534 9.3005
R18622 vdd.n1537 vdd.n1536 9.3005
R18623 vdd.n1520 vdd.n1519 9.3005
R18624 vdd.n1543 vdd.n1542 9.3005
R18625 vdd.n1545 vdd.n1544 9.3005
R18626 vdd.n1517 vdd.n1514 9.3005
R18627 vdd.n1552 vdd.n1551 9.3005
R18628 vdd.n1384 vdd.n1383 9.3005
R18629 vdd.n1379 vdd.n1378 9.3005
R18630 vdd.n1390 vdd.n1389 9.3005
R18631 vdd.n1392 vdd.n1391 9.3005
R18632 vdd.n1375 vdd.n1374 9.3005
R18633 vdd.n1398 vdd.n1397 9.3005
R18634 vdd.n1400 vdd.n1399 9.3005
R18635 vdd.n1372 vdd.n1369 9.3005
R18636 vdd.n1407 vdd.n1406 9.3005
R18637 vdd.n1435 vdd.n1434 9.3005
R18638 vdd.n1430 vdd.n1429 9.3005
R18639 vdd.n1441 vdd.n1440 9.3005
R18640 vdd.n1443 vdd.n1442 9.3005
R18641 vdd.n1426 vdd.n1425 9.3005
R18642 vdd.n1449 vdd.n1448 9.3005
R18643 vdd.n1451 vdd.n1450 9.3005
R18644 vdd.n1423 vdd.n1420 9.3005
R18645 vdd.n1458 vdd.n1457 9.3005
R18646 vdd.n1291 vdd.n1290 9.3005
R18647 vdd.n1286 vdd.n1285 9.3005
R18648 vdd.n1297 vdd.n1296 9.3005
R18649 vdd.n1299 vdd.n1298 9.3005
R18650 vdd.n1282 vdd.n1281 9.3005
R18651 vdd.n1305 vdd.n1304 9.3005
R18652 vdd.n1307 vdd.n1306 9.3005
R18653 vdd.n1279 vdd.n1276 9.3005
R18654 vdd.n1314 vdd.n1313 9.3005
R18655 vdd.n1342 vdd.n1341 9.3005
R18656 vdd.n1337 vdd.n1336 9.3005
R18657 vdd.n1348 vdd.n1347 9.3005
R18658 vdd.n1350 vdd.n1349 9.3005
R18659 vdd.n1333 vdd.n1332 9.3005
R18660 vdd.n1356 vdd.n1355 9.3005
R18661 vdd.n1358 vdd.n1357 9.3005
R18662 vdd.n1330 vdd.n1327 9.3005
R18663 vdd.n1365 vdd.n1364 9.3005
R18664 vdd.n288 vdd.n287 8.92171
R18665 vdd.n237 vdd.n236 8.92171
R18666 vdd.n194 vdd.n193 8.92171
R18667 vdd.n143 vdd.n142 8.92171
R18668 vdd.n101 vdd.n100 8.92171
R18669 vdd.n50 vdd.n49 8.92171
R18670 vdd.n1483 vdd.n1482 8.92171
R18671 vdd.n1534 vdd.n1533 8.92171
R18672 vdd.n1389 vdd.n1388 8.92171
R18673 vdd.n1440 vdd.n1439 8.92171
R18674 vdd.n1296 vdd.n1295 8.92171
R18675 vdd.n1347 vdd.n1346 8.92171
R18676 vdd.n215 vdd.n121 8.81535
R18677 vdd.n1461 vdd.n1367 8.81535
R18678 vdd.n1596 vdd.t42 8.72962
R18679 vdd.n2956 vdd.t21 8.72962
R18680 vdd.t39 vdd.n1570 8.50289
R18681 vdd.n493 vdd.t147 8.50289
R18682 vdd.n28 vdd.n14 8.42249
R18683 vdd.n1272 vdd.t208 8.27616
R18684 vdd.n3164 vdd.t187 8.27616
R18685 vdd.n3168 vdd.n3167 8.16225
R18686 vdd.n1557 vdd.n1556 8.16225
R18687 vdd.n284 vdd.n278 8.14595
R18688 vdd.n233 vdd.n227 8.14595
R18689 vdd.n190 vdd.n184 8.14595
R18690 vdd.n139 vdd.n133 8.14595
R18691 vdd.n97 vdd.n91 8.14595
R18692 vdd.n46 vdd.n40 8.14595
R18693 vdd.n1479 vdd.n1473 8.14595
R18694 vdd.n1530 vdd.n1524 8.14595
R18695 vdd.n1385 vdd.n1379 8.14595
R18696 vdd.n1436 vdd.n1430 8.14595
R18697 vdd.n1292 vdd.n1286 8.14595
R18698 vdd.n1343 vdd.n1337 8.14595
R18699 vdd.n2635 vdd.n677 8.11757
R18700 vdd.n2109 vdd.n2108 8.11757
R18701 vdd.t168 vdd.n960 8.04943
R18702 vdd.n3155 vdd.t149 8.04943
R18703 vdd.n2087 vdd.n871 7.70933
R18704 vdd.n2093 vdd.n871 7.70933
R18705 vdd.n2099 vdd.n865 7.70933
R18706 vdd.n2099 vdd.n858 7.70933
R18707 vdd.n2105 vdd.n858 7.70933
R18708 vdd.n2105 vdd.n861 7.70933
R18709 vdd.n2112 vdd.n846 7.70933
R18710 vdd.n2118 vdd.n846 7.70933
R18711 vdd.n2124 vdd.n840 7.70933
R18712 vdd.n2130 vdd.n836 7.70933
R18713 vdd.n2136 vdd.n830 7.70933
R18714 vdd.n2148 vdd.n817 7.70933
R18715 vdd.n2154 vdd.n811 7.70933
R18716 vdd.n2154 vdd.n804 7.70933
R18717 vdd.n2162 vdd.n804 7.70933
R18718 vdd.n2169 vdd.t144 7.70933
R18719 vdd.n2244 vdd.t144 7.70933
R18720 vdd.n2576 vdd.t170 7.70933
R18721 vdd.n2582 vdd.t170 7.70933
R18722 vdd.n2588 vdd.n725 7.70933
R18723 vdd.n2594 vdd.n725 7.70933
R18724 vdd.n2594 vdd.n728 7.70933
R18725 vdd.n2600 vdd.n721 7.70933
R18726 vdd.n2612 vdd.n708 7.70933
R18727 vdd.n2618 vdd.n702 7.70933
R18728 vdd.n2624 vdd.n698 7.70933
R18729 vdd.n2630 vdd.n685 7.70933
R18730 vdd.n2638 vdd.n685 7.70933
R18731 vdd.n2644 vdd.n679 7.70933
R18732 vdd.n2644 vdd.n671 7.70933
R18733 vdd.n2695 vdd.n671 7.70933
R18734 vdd.n2695 vdd.n674 7.70933
R18735 vdd.n2701 vdd.n631 7.70933
R18736 vdd.n2771 vdd.n631 7.70933
R18737 vdd.n283 vdd.n280 7.3702
R18738 vdd.n232 vdd.n229 7.3702
R18739 vdd.n189 vdd.n186 7.3702
R18740 vdd.n138 vdd.n135 7.3702
R18741 vdd.n96 vdd.n93 7.3702
R18742 vdd.n45 vdd.n42 7.3702
R18743 vdd.n1478 vdd.n1475 7.3702
R18744 vdd.n1529 vdd.n1526 7.3702
R18745 vdd.n1384 vdd.n1381 7.3702
R18746 vdd.n1435 vdd.n1432 7.3702
R18747 vdd.n1291 vdd.n1288 7.3702
R18748 vdd.n1342 vdd.n1339 7.3702
R18749 vdd.n1239 vdd.t48 7.1425
R18750 vdd.n3148 vdd.t154 7.1425
R18751 vdd.n1150 vdd.n1149 6.98232
R18752 vdd.n1751 vdd.n1750 6.98232
R18753 vdd.n3063 vdd.n3062 6.98232
R18754 vdd.n2855 vdd.n2854 6.98232
R18755 vdd.n1255 vdd.t25 6.91577
R18756 vdd.n325 vdd.t23 6.91577
R18757 vdd.n1562 vdd.t30 6.68904
R18758 vdd.n2989 vdd.t6 6.68904
R18759 vdd.n925 vdd.t44 6.46231
R18760 vdd.t19 vdd.n492 6.46231
R18761 vdd.n3168 vdd.n309 6.27748
R18762 vdd.n1556 vdd.n1555 6.27748
R18763 vdd.n2124 vdd.t151 6.00885
R18764 vdd.n2624 vdd.t143 6.00885
R18765 vdd.n861 vdd.t102 5.89549
R18766 vdd.t70 vdd.n679 5.89549
R18767 vdd.n284 vdd.n283 5.81868
R18768 vdd.n233 vdd.n232 5.81868
R18769 vdd.n190 vdd.n189 5.81868
R18770 vdd.n139 vdd.n138 5.81868
R18771 vdd.n97 vdd.n96 5.81868
R18772 vdd.n46 vdd.n45 5.81868
R18773 vdd.n1479 vdd.n1478 5.81868
R18774 vdd.n1530 vdd.n1529 5.81868
R18775 vdd.n1385 vdd.n1384 5.81868
R18776 vdd.n1436 vdd.n1435 5.81868
R18777 vdd.n1292 vdd.n1291 5.81868
R18778 vdd.n1343 vdd.n1342 5.81868
R18779 vdd.t98 vdd.n865 5.78212
R18780 vdd.n1868 vdd.t83 5.78212
R18781 vdd.n2493 vdd.t91 5.78212
R18782 vdd.n674 vdd.t87 5.78212
R18783 vdd.n2252 vdd.n2251 5.77611
R18784 vdd.n1995 vdd.n1865 5.77611
R18785 vdd.n2506 vdd.n2505 5.77611
R18786 vdd.n2710 vdd.n663 5.77611
R18787 vdd.n2776 vdd.n627 5.77611
R18788 vdd.n2416 vdd.n2356 5.77611
R18789 vdd.n2177 vdd.n795 5.77611
R18790 vdd.n1925 vdd.n1924 5.77611
R18791 vdd.n1112 vdd.n1109 5.62474
R18792 vdd.n2047 vdd.n2044 5.62474
R18793 vdd.n3023 vdd.n3020 5.62474
R18794 vdd.n2810 vdd.n2807 5.62474
R18795 vdd.t159 vdd.n817 5.44203
R18796 vdd.n721 vdd.t165 5.44203
R18797 vdd.t174 vdd.n840 5.10193
R18798 vdd.n830 vdd.t132 5.10193
R18799 vdd.t34 vdd.n708 5.10193
R18800 vdd.n698 vdd.t146 5.10193
R18801 vdd.n287 vdd.n278 5.04292
R18802 vdd.n236 vdd.n227 5.04292
R18803 vdd.n193 vdd.n184 5.04292
R18804 vdd.n142 vdd.n133 5.04292
R18805 vdd.n100 vdd.n91 5.04292
R18806 vdd.n49 vdd.n40 5.04292
R18807 vdd.n1482 vdd.n1473 5.04292
R18808 vdd.n1533 vdd.n1524 5.04292
R18809 vdd.n1388 vdd.n1379 5.04292
R18810 vdd.n1439 vdd.n1430 5.04292
R18811 vdd.n1295 vdd.n1286 5.04292
R18812 vdd.n1346 vdd.n1337 5.04292
R18813 vdd.n1588 vdd.t44 4.8752
R18814 vdd.t219 vdd.t184 4.8752
R18815 vdd.t9 vdd.t226 4.8752
R18816 vdd.t130 vdd.t15 4.8752
R18817 vdd.t161 vdd.t16 4.8752
R18818 vdd.n2964 vdd.t19 4.8752
R18819 vdd.n2253 vdd.n2252 4.83952
R18820 vdd.n1865 vdd.n1861 4.83952
R18821 vdd.n2507 vdd.n2506 4.83952
R18822 vdd.n663 vdd.n658 4.83952
R18823 vdd.n627 vdd.n622 4.83952
R18824 vdd.n2413 vdd.n2356 4.83952
R18825 vdd.n2180 vdd.n795 4.83952
R18826 vdd.n1924 vdd.n1923 4.83952
R18827 vdd.n1719 vdd.n893 4.74817
R18828 vdd.n1714 vdd.n894 4.74817
R18829 vdd.n1616 vdd.n1613 4.74817
R18830 vdd.n2028 vdd.n1617 4.74817
R18831 vdd.n2030 vdd.n1616 4.74817
R18832 vdd.n2029 vdd.n2028 4.74817
R18833 vdd.n521 vdd.n519 4.74817
R18834 vdd.n2925 vdd.n522 4.74817
R18835 vdd.n2928 vdd.n522 4.74817
R18836 vdd.n2929 vdd.n521 4.74817
R18837 vdd.n2817 vdd.n606 4.74817
R18838 vdd.n2813 vdd.n608 4.74817
R18839 vdd.n2816 vdd.n608 4.74817
R18840 vdd.n2821 vdd.n606 4.74817
R18841 vdd.n1715 vdd.n893 4.74817
R18842 vdd.n896 vdd.n894 4.74817
R18843 vdd.n309 vdd.n308 4.7074
R18844 vdd.n215 vdd.n214 4.7074
R18845 vdd.n1555 vdd.n1554 4.7074
R18846 vdd.n1461 vdd.n1460 4.7074
R18847 vdd.t30 vdd.n931 4.64847
R18848 vdd.n2980 vdd.t6 4.64847
R18849 vdd.n2130 vdd.t220 4.53511
R18850 vdd.n2618 vdd.t198 4.53511
R18851 vdd.n1264 vdd.t25 4.42174
R18852 vdd.n3162 vdd.t23 4.42174
R18853 vdd.n2162 vdd.t196 4.30838
R18854 vdd.n2588 vdd.t13 4.30838
R18855 vdd.n288 vdd.n276 4.26717
R18856 vdd.n237 vdd.n225 4.26717
R18857 vdd.n194 vdd.n182 4.26717
R18858 vdd.n143 vdd.n131 4.26717
R18859 vdd.n101 vdd.n89 4.26717
R18860 vdd.n50 vdd.n38 4.26717
R18861 vdd.n1483 vdd.n1471 4.26717
R18862 vdd.n1534 vdd.n1522 4.26717
R18863 vdd.n1389 vdd.n1377 4.26717
R18864 vdd.n1440 vdd.n1428 4.26717
R18865 vdd.n1296 vdd.n1284 4.26717
R18866 vdd.n1347 vdd.n1335 4.26717
R18867 vdd.t48 vdd.n959 4.19501
R18868 vdd.t154 vdd.n329 4.19501
R18869 vdd.n309 vdd.n215 4.10845
R18870 vdd.n1555 vdd.n1461 4.10845
R18871 vdd.n265 vdd.t150 4.06363
R18872 vdd.n265 vdd.t167 4.06363
R18873 vdd.n263 vdd.t186 4.06363
R18874 vdd.n263 vdd.t211 4.06363
R18875 vdd.n261 vdd.t37 4.06363
R18876 vdd.n261 vdd.t213 4.06363
R18877 vdd.n259 vdd.t228 4.06363
R18878 vdd.n259 vdd.t224 4.06363
R18879 vdd.n257 vdd.t20 4.06363
R18880 vdd.n257 vdd.t194 4.06363
R18881 vdd.n171 vdd.t204 4.06363
R18882 vdd.n171 vdd.t155 4.06363
R18883 vdd.n169 vdd.t193 4.06363
R18884 vdd.n169 vdd.t192 4.06363
R18885 vdd.n167 vdd.t142 4.06363
R18886 vdd.n167 vdd.t190 4.06363
R18887 vdd.n165 vdd.t177 4.06363
R18888 vdd.n165 vdd.t7 4.06363
R18889 vdd.n163 vdd.t210 4.06363
R18890 vdd.n163 vdd.t141 4.06363
R18891 vdd.n78 vdd.t180 4.06363
R18892 vdd.n78 vdd.t217 4.06363
R18893 vdd.n76 vdd.t24 4.06363
R18894 vdd.n76 vdd.t139 4.06363
R18895 vdd.n74 vdd.t36 4.06363
R18896 vdd.n74 vdd.t188 4.06363
R18897 vdd.n72 vdd.t148 4.06363
R18898 vdd.n72 vdd.t183 4.06363
R18899 vdd.n70 vdd.t133 4.06363
R18900 vdd.n70 vdd.t29 4.06363
R18901 vdd.n1503 vdd.t216 4.06363
R18902 vdd.n1503 vdd.t45 4.06363
R18903 vdd.n1505 vdd.t31 4.06363
R18904 vdd.n1505 vdd.t136 4.06363
R18905 vdd.n1507 vdd.t209 4.06363
R18906 vdd.n1507 vdd.t229 4.06363
R18907 vdd.n1509 vdd.t191 4.06363
R18908 vdd.n1509 vdd.t137 4.06363
R18909 vdd.n1511 vdd.t203 4.06363
R18910 vdd.n1511 vdd.t169 4.06363
R18911 vdd.n1409 vdd.t231 4.06363
R18912 vdd.n1409 vdd.t134 4.06363
R18913 vdd.n1411 vdd.t207 4.06363
R18914 vdd.n1411 vdd.t40 4.06363
R18915 vdd.n1413 vdd.t212 4.06363
R18916 vdd.n1413 vdd.t179 4.06363
R18917 vdd.n1415 vdd.t33 4.06363
R18918 vdd.n1415 vdd.t41 4.06363
R18919 vdd.n1417 vdd.t49 4.06363
R18920 vdd.n1417 vdd.t182 4.06363
R18921 vdd.n1316 vdd.t5 4.06363
R18922 vdd.n1316 vdd.t205 4.06363
R18923 vdd.n1318 vdd.t215 4.06363
R18924 vdd.n1318 vdd.t140 4.06363
R18925 vdd.n1320 vdd.t222 4.06363
R18926 vdd.n1320 vdd.t206 4.06363
R18927 vdd.n1322 vdd.t225 4.06363
R18928 vdd.n1322 vdd.t26 4.06363
R18929 vdd.n1324 vdd.t218 4.06363
R18930 vdd.n1324 vdd.t181 4.06363
R18931 vdd.n26 vdd.t51 3.9605
R18932 vdd.n26 vdd.t0 3.9605
R18933 vdd.n23 vdd.t2 3.9605
R18934 vdd.n23 vdd.t135 3.9605
R18935 vdd.n21 vdd.t1 3.9605
R18936 vdd.n21 vdd.t50 3.9605
R18937 vdd.n20 vdd.t157 3.9605
R18938 vdd.n20 vdd.t12 3.9605
R18939 vdd.n15 vdd.t189 3.9605
R18940 vdd.n15 vdd.t158 3.9605
R18941 vdd.n16 vdd.t53 3.9605
R18942 vdd.n16 vdd.t11 3.9605
R18943 vdd.n18 vdd.t8 3.9605
R18944 vdd.n18 vdd.t52 3.9605
R18945 vdd.n25 vdd.t10 3.9605
R18946 vdd.n25 vdd.t156 3.9605
R18947 vdd.n7 vdd.t162 3.61217
R18948 vdd.n7 vdd.t199 3.61217
R18949 vdd.n8 vdd.t131 3.61217
R18950 vdd.n8 vdd.t166 3.61217
R18951 vdd.n10 vdd.t171 3.61217
R18952 vdd.n10 vdd.t14 3.61217
R18953 vdd.n12 vdd.t201 3.61217
R18954 vdd.n12 vdd.t173 3.61217
R18955 vdd.n5 vdd.t164 3.61217
R18956 vdd.n5 vdd.t18 3.61217
R18957 vdd.n3 vdd.t197 3.61217
R18958 vdd.n3 vdd.t145 3.61217
R18959 vdd.n1 vdd.t160 3.61217
R18960 vdd.n1 vdd.t227 3.61217
R18961 vdd.n0 vdd.t221 3.61217
R18962 vdd.n0 vdd.t185 3.61217
R18963 vdd.n292 vdd.n291 3.49141
R18964 vdd.n241 vdd.n240 3.49141
R18965 vdd.n198 vdd.n197 3.49141
R18966 vdd.n147 vdd.n146 3.49141
R18967 vdd.n105 vdd.n104 3.49141
R18968 vdd.n54 vdd.n53 3.49141
R18969 vdd.n1487 vdd.n1486 3.49141
R18970 vdd.n1538 vdd.n1537 3.49141
R18971 vdd.n1393 vdd.n1392 3.49141
R18972 vdd.n1444 vdd.n1443 3.49141
R18973 vdd.n1300 vdd.n1299 3.49141
R18974 vdd.n1351 vdd.n1350 3.49141
R18975 vdd.n1868 vdd.t196 3.40145
R18976 vdd.n2316 vdd.t163 3.40145
R18977 vdd.n2569 vdd.t172 3.40145
R18978 vdd.n2493 vdd.t13 3.40145
R18979 vdd.n1247 vdd.t168 3.28809
R18980 vdd.t149 vdd.n3154 3.28809
R18981 vdd.n1969 vdd.t220 3.17472
R18982 vdd.n2472 vdd.t198 3.17472
R18983 vdd.n948 vdd.t208 3.06136
R18984 vdd.t187 vdd.n3163 3.06136
R18985 vdd.n1571 vdd.t39 2.83463
R18986 vdd.n2981 vdd.t147 2.83463
R18987 vdd.n295 vdd.n274 2.71565
R18988 vdd.n244 vdd.n223 2.71565
R18989 vdd.n201 vdd.n180 2.71565
R18990 vdd.n150 vdd.n129 2.71565
R18991 vdd.n108 vdd.n87 2.71565
R18992 vdd.n57 vdd.n36 2.71565
R18993 vdd.n1490 vdd.n1469 2.71565
R18994 vdd.n1541 vdd.n1520 2.71565
R18995 vdd.n1396 vdd.n1375 2.71565
R18996 vdd.n1447 vdd.n1426 2.71565
R18997 vdd.n1303 vdd.n1282 2.71565
R18998 vdd.n1354 vdd.n1333 2.71565
R18999 vdd.n1587 vdd.t42 2.6079
R19000 vdd.n2118 vdd.t174 2.6079
R19001 vdd.n2142 vdd.t132 2.6079
R19002 vdd.n2606 vdd.t34 2.6079
R19003 vdd.n2630 vdd.t146 2.6079
R19004 vdd.t21 vdd.n499 2.6079
R19005 vdd.n2636 vdd.n2635 2.49806
R19006 vdd.n2110 vdd.n2109 2.49806
R19007 vdd.n282 vdd.n281 2.4129
R19008 vdd.n231 vdd.n230 2.4129
R19009 vdd.n188 vdd.n187 2.4129
R19010 vdd.n137 vdd.n136 2.4129
R19011 vdd.n95 vdd.n94 2.4129
R19012 vdd.n44 vdd.n43 2.4129
R19013 vdd.n1477 vdd.n1476 2.4129
R19014 vdd.n1528 vdd.n1527 2.4129
R19015 vdd.n1383 vdd.n1382 2.4129
R19016 vdd.n1434 vdd.n1433 2.4129
R19017 vdd.n1290 vdd.n1289 2.4129
R19018 vdd.n1341 vdd.n1340 2.4129
R19019 vdd.n2027 vdd.n1616 2.27742
R19020 vdd.n2028 vdd.n2027 2.27742
R19021 vdd.n2737 vdd.n522 2.27742
R19022 vdd.n2737 vdd.n521 2.27742
R19023 vdd.n2805 vdd.n608 2.27742
R19024 vdd.n2805 vdd.n606 2.27742
R19025 vdd.n2050 vdd.n893 2.27742
R19026 vdd.n2050 vdd.n894 2.27742
R19027 vdd.n2142 vdd.t159 2.2678
R19028 vdd.n2606 vdd.t165 2.2678
R19029 vdd.t226 vdd.n811 2.04107
R19030 vdd.n728 vdd.t130 2.04107
R19031 vdd.n296 vdd.n272 1.93989
R19032 vdd.n245 vdd.n221 1.93989
R19033 vdd.n202 vdd.n178 1.93989
R19034 vdd.n151 vdd.n127 1.93989
R19035 vdd.n109 vdd.n85 1.93989
R19036 vdd.n58 vdd.n34 1.93989
R19037 vdd.n1491 vdd.n1467 1.93989
R19038 vdd.n1542 vdd.n1518 1.93989
R19039 vdd.n1397 vdd.n1373 1.93989
R19040 vdd.n1448 vdd.n1424 1.93989
R19041 vdd.n1304 vdd.n1280 1.93989
R19042 vdd.n1355 vdd.n1331 1.93989
R19043 vdd.n2093 vdd.t98 1.92771
R19044 vdd.n2169 vdd.t83 1.92771
R19045 vdd.n2582 vdd.t91 1.92771
R19046 vdd.n2701 vdd.t87 1.92771
R19047 vdd.n1969 vdd.t151 1.70098
R19048 vdd.n836 vdd.t219 1.70098
R19049 vdd.t16 vdd.n702 1.70098
R19050 vdd.n2472 vdd.t143 1.70098
R19051 vdd.n983 vdd.t66 1.47425
R19052 vdd.t115 vdd.n3139 1.47425
R19053 vdd.n307 vdd.n267 1.16414
R19054 vdd.n300 vdd.n299 1.16414
R19055 vdd.n256 vdd.n216 1.16414
R19056 vdd.n249 vdd.n248 1.16414
R19057 vdd.n213 vdd.n173 1.16414
R19058 vdd.n206 vdd.n205 1.16414
R19059 vdd.n162 vdd.n122 1.16414
R19060 vdd.n155 vdd.n154 1.16414
R19061 vdd.n120 vdd.n80 1.16414
R19062 vdd.n113 vdd.n112 1.16414
R19063 vdd.n69 vdd.n29 1.16414
R19064 vdd.n62 vdd.n61 1.16414
R19065 vdd.n1502 vdd.n1462 1.16414
R19066 vdd.n1495 vdd.n1494 1.16414
R19067 vdd.n1553 vdd.n1513 1.16414
R19068 vdd.n1546 vdd.n1545 1.16414
R19069 vdd.n1408 vdd.n1368 1.16414
R19070 vdd.n1401 vdd.n1400 1.16414
R19071 vdd.n1459 vdd.n1419 1.16414
R19072 vdd.n1452 vdd.n1451 1.16414
R19073 vdd.n1315 vdd.n1275 1.16414
R19074 vdd.n1308 vdd.n1307 1.16414
R19075 vdd.n1366 vdd.n1326 1.16414
R19076 vdd.n1359 vdd.n1358 1.16414
R19077 vdd.n2136 vdd.t184 1.13415
R19078 vdd.n2612 vdd.t161 1.13415
R19079 vdd.n1579 vdd.t4 1.02079
R19080 vdd.t102 vdd.t3 1.02079
R19081 vdd.t38 vdd.t70 1.02079
R19082 vdd.n2972 vdd.t28 1.02079
R19083 vdd.n1113 vdd.n1112 0.970197
R19084 vdd.n2048 vdd.n2047 0.970197
R19085 vdd.n3024 vdd.n3023 0.970197
R19086 vdd.n2812 vdd.n2810 0.970197
R19087 vdd.n1556 vdd.n28 0.800283
R19088 vdd.t178 vdd.n937 0.794056
R19089 vdd.n1606 vdd.t62 0.794056
R19090 vdd.n2112 vdd.t3 0.794056
R19091 vdd.n2148 vdd.t9 0.794056
R19092 vdd.n2600 vdd.t15 0.794056
R19093 vdd.n2638 vdd.t38 0.794056
R19094 vdd.t55 vdd.n511 0.794056
R19095 vdd.n481 vdd.t35 0.794056
R19096 vdd vdd.n3168 0.79245
R19097 vdd.n1256 vdd.t32 0.567326
R19098 vdd.n3156 vdd.t138 0.567326
R19099 vdd.n2038 vdd.n2037 0.509646
R19100 vdd.n2937 vdd.n2936 0.509646
R19101 vdd.n3135 vdd.n3134 0.509646
R19102 vdd.n3017 vdd.n3016 0.509646
R19103 vdd.n2943 vdd.n514 0.509646
R19104 vdd.n1601 vdd.n895 0.509646
R19105 vdd.n1218 vdd.n980 0.509646
R19106 vdd.n1212 vdd.n1211 0.509646
R19107 vdd.n4 vdd.n2 0.459552
R19108 vdd.n11 vdd.n9 0.459552
R19109 vdd.n305 vdd.n304 0.388379
R19110 vdd.n271 vdd.n269 0.388379
R19111 vdd.n254 vdd.n253 0.388379
R19112 vdd.n220 vdd.n218 0.388379
R19113 vdd.n211 vdd.n210 0.388379
R19114 vdd.n177 vdd.n175 0.388379
R19115 vdd.n160 vdd.n159 0.388379
R19116 vdd.n126 vdd.n124 0.388379
R19117 vdd.n118 vdd.n117 0.388379
R19118 vdd.n84 vdd.n82 0.388379
R19119 vdd.n67 vdd.n66 0.388379
R19120 vdd.n33 vdd.n31 0.388379
R19121 vdd.n1500 vdd.n1499 0.388379
R19122 vdd.n1466 vdd.n1464 0.388379
R19123 vdd.n1551 vdd.n1550 0.388379
R19124 vdd.n1517 vdd.n1515 0.388379
R19125 vdd.n1406 vdd.n1405 0.388379
R19126 vdd.n1372 vdd.n1370 0.388379
R19127 vdd.n1457 vdd.n1456 0.388379
R19128 vdd.n1423 vdd.n1421 0.388379
R19129 vdd.n1313 vdd.n1312 0.388379
R19130 vdd.n1279 vdd.n1277 0.388379
R19131 vdd.n1364 vdd.n1363 0.388379
R19132 vdd.n1330 vdd.n1328 0.388379
R19133 vdd.n19 vdd.n17 0.387128
R19134 vdd.n24 vdd.n22 0.387128
R19135 vdd.n6 vdd.n4 0.358259
R19136 vdd.n13 vdd.n11 0.358259
R19137 vdd.n260 vdd.n258 0.358259
R19138 vdd.n262 vdd.n260 0.358259
R19139 vdd.n264 vdd.n262 0.358259
R19140 vdd.n266 vdd.n264 0.358259
R19141 vdd.n308 vdd.n266 0.358259
R19142 vdd.n166 vdd.n164 0.358259
R19143 vdd.n168 vdd.n166 0.358259
R19144 vdd.n170 vdd.n168 0.358259
R19145 vdd.n172 vdd.n170 0.358259
R19146 vdd.n214 vdd.n172 0.358259
R19147 vdd.n73 vdd.n71 0.358259
R19148 vdd.n75 vdd.n73 0.358259
R19149 vdd.n77 vdd.n75 0.358259
R19150 vdd.n79 vdd.n77 0.358259
R19151 vdd.n121 vdd.n79 0.358259
R19152 vdd.n1554 vdd.n1512 0.358259
R19153 vdd.n1512 vdd.n1510 0.358259
R19154 vdd.n1510 vdd.n1508 0.358259
R19155 vdd.n1508 vdd.n1506 0.358259
R19156 vdd.n1506 vdd.n1504 0.358259
R19157 vdd.n1460 vdd.n1418 0.358259
R19158 vdd.n1418 vdd.n1416 0.358259
R19159 vdd.n1416 vdd.n1414 0.358259
R19160 vdd.n1414 vdd.n1412 0.358259
R19161 vdd.n1412 vdd.n1410 0.358259
R19162 vdd.n1367 vdd.n1325 0.358259
R19163 vdd.n1325 vdd.n1323 0.358259
R19164 vdd.n1323 vdd.n1321 0.358259
R19165 vdd.n1321 vdd.n1319 0.358259
R19166 vdd.n1319 vdd.n1317 0.358259
R19167 vdd.t46 vdd.n966 0.340595
R19168 vdd.n3147 vdd.t152 0.340595
R19169 vdd.n14 vdd.n6 0.334552
R19170 vdd.n14 vdd.n13 0.334552
R19171 vdd.n27 vdd.n19 0.21707
R19172 vdd.n27 vdd.n24 0.21707
R19173 vdd.n306 vdd.n268 0.155672
R19174 vdd.n298 vdd.n268 0.155672
R19175 vdd.n298 vdd.n297 0.155672
R19176 vdd.n297 vdd.n273 0.155672
R19177 vdd.n290 vdd.n273 0.155672
R19178 vdd.n290 vdd.n289 0.155672
R19179 vdd.n289 vdd.n277 0.155672
R19180 vdd.n282 vdd.n277 0.155672
R19181 vdd.n255 vdd.n217 0.155672
R19182 vdd.n247 vdd.n217 0.155672
R19183 vdd.n247 vdd.n246 0.155672
R19184 vdd.n246 vdd.n222 0.155672
R19185 vdd.n239 vdd.n222 0.155672
R19186 vdd.n239 vdd.n238 0.155672
R19187 vdd.n238 vdd.n226 0.155672
R19188 vdd.n231 vdd.n226 0.155672
R19189 vdd.n212 vdd.n174 0.155672
R19190 vdd.n204 vdd.n174 0.155672
R19191 vdd.n204 vdd.n203 0.155672
R19192 vdd.n203 vdd.n179 0.155672
R19193 vdd.n196 vdd.n179 0.155672
R19194 vdd.n196 vdd.n195 0.155672
R19195 vdd.n195 vdd.n183 0.155672
R19196 vdd.n188 vdd.n183 0.155672
R19197 vdd.n161 vdd.n123 0.155672
R19198 vdd.n153 vdd.n123 0.155672
R19199 vdd.n153 vdd.n152 0.155672
R19200 vdd.n152 vdd.n128 0.155672
R19201 vdd.n145 vdd.n128 0.155672
R19202 vdd.n145 vdd.n144 0.155672
R19203 vdd.n144 vdd.n132 0.155672
R19204 vdd.n137 vdd.n132 0.155672
R19205 vdd.n119 vdd.n81 0.155672
R19206 vdd.n111 vdd.n81 0.155672
R19207 vdd.n111 vdd.n110 0.155672
R19208 vdd.n110 vdd.n86 0.155672
R19209 vdd.n103 vdd.n86 0.155672
R19210 vdd.n103 vdd.n102 0.155672
R19211 vdd.n102 vdd.n90 0.155672
R19212 vdd.n95 vdd.n90 0.155672
R19213 vdd.n68 vdd.n30 0.155672
R19214 vdd.n60 vdd.n30 0.155672
R19215 vdd.n60 vdd.n59 0.155672
R19216 vdd.n59 vdd.n35 0.155672
R19217 vdd.n52 vdd.n35 0.155672
R19218 vdd.n52 vdd.n51 0.155672
R19219 vdd.n51 vdd.n39 0.155672
R19220 vdd.n44 vdd.n39 0.155672
R19221 vdd.n1501 vdd.n1463 0.155672
R19222 vdd.n1493 vdd.n1463 0.155672
R19223 vdd.n1493 vdd.n1492 0.155672
R19224 vdd.n1492 vdd.n1468 0.155672
R19225 vdd.n1485 vdd.n1468 0.155672
R19226 vdd.n1485 vdd.n1484 0.155672
R19227 vdd.n1484 vdd.n1472 0.155672
R19228 vdd.n1477 vdd.n1472 0.155672
R19229 vdd.n1552 vdd.n1514 0.155672
R19230 vdd.n1544 vdd.n1514 0.155672
R19231 vdd.n1544 vdd.n1543 0.155672
R19232 vdd.n1543 vdd.n1519 0.155672
R19233 vdd.n1536 vdd.n1519 0.155672
R19234 vdd.n1536 vdd.n1535 0.155672
R19235 vdd.n1535 vdd.n1523 0.155672
R19236 vdd.n1528 vdd.n1523 0.155672
R19237 vdd.n1407 vdd.n1369 0.155672
R19238 vdd.n1399 vdd.n1369 0.155672
R19239 vdd.n1399 vdd.n1398 0.155672
R19240 vdd.n1398 vdd.n1374 0.155672
R19241 vdd.n1391 vdd.n1374 0.155672
R19242 vdd.n1391 vdd.n1390 0.155672
R19243 vdd.n1390 vdd.n1378 0.155672
R19244 vdd.n1383 vdd.n1378 0.155672
R19245 vdd.n1458 vdd.n1420 0.155672
R19246 vdd.n1450 vdd.n1420 0.155672
R19247 vdd.n1450 vdd.n1449 0.155672
R19248 vdd.n1449 vdd.n1425 0.155672
R19249 vdd.n1442 vdd.n1425 0.155672
R19250 vdd.n1442 vdd.n1441 0.155672
R19251 vdd.n1441 vdd.n1429 0.155672
R19252 vdd.n1434 vdd.n1429 0.155672
R19253 vdd.n1314 vdd.n1276 0.155672
R19254 vdd.n1306 vdd.n1276 0.155672
R19255 vdd.n1306 vdd.n1305 0.155672
R19256 vdd.n1305 vdd.n1281 0.155672
R19257 vdd.n1298 vdd.n1281 0.155672
R19258 vdd.n1298 vdd.n1297 0.155672
R19259 vdd.n1297 vdd.n1285 0.155672
R19260 vdd.n1290 vdd.n1285 0.155672
R19261 vdd.n1365 vdd.n1327 0.155672
R19262 vdd.n1357 vdd.n1327 0.155672
R19263 vdd.n1357 vdd.n1356 0.155672
R19264 vdd.n1356 vdd.n1332 0.155672
R19265 vdd.n1349 vdd.n1332 0.155672
R19266 vdd.n1349 vdd.n1348 0.155672
R19267 vdd.n1348 vdd.n1336 0.155672
R19268 vdd.n1341 vdd.n1336 0.155672
R19269 vdd.n1813 vdd.n1618 0.152939
R19270 vdd.n1624 vdd.n1618 0.152939
R19271 vdd.n1625 vdd.n1624 0.152939
R19272 vdd.n1626 vdd.n1625 0.152939
R19273 vdd.n1627 vdd.n1626 0.152939
R19274 vdd.n1631 vdd.n1627 0.152939
R19275 vdd.n1632 vdd.n1631 0.152939
R19276 vdd.n1633 vdd.n1632 0.152939
R19277 vdd.n1634 vdd.n1633 0.152939
R19278 vdd.n1638 vdd.n1634 0.152939
R19279 vdd.n1639 vdd.n1638 0.152939
R19280 vdd.n1640 vdd.n1639 0.152939
R19281 vdd.n1788 vdd.n1640 0.152939
R19282 vdd.n1788 vdd.n1787 0.152939
R19283 vdd.n1787 vdd.n1786 0.152939
R19284 vdd.n1786 vdd.n1646 0.152939
R19285 vdd.n1651 vdd.n1646 0.152939
R19286 vdd.n1652 vdd.n1651 0.152939
R19287 vdd.n1653 vdd.n1652 0.152939
R19288 vdd.n1657 vdd.n1653 0.152939
R19289 vdd.n1658 vdd.n1657 0.152939
R19290 vdd.n1659 vdd.n1658 0.152939
R19291 vdd.n1660 vdd.n1659 0.152939
R19292 vdd.n1664 vdd.n1660 0.152939
R19293 vdd.n1665 vdd.n1664 0.152939
R19294 vdd.n1666 vdd.n1665 0.152939
R19295 vdd.n1667 vdd.n1666 0.152939
R19296 vdd.n1671 vdd.n1667 0.152939
R19297 vdd.n1672 vdd.n1671 0.152939
R19298 vdd.n1673 vdd.n1672 0.152939
R19299 vdd.n1674 vdd.n1673 0.152939
R19300 vdd.n1678 vdd.n1674 0.152939
R19301 vdd.n1679 vdd.n1678 0.152939
R19302 vdd.n1680 vdd.n1679 0.152939
R19303 vdd.n1749 vdd.n1680 0.152939
R19304 vdd.n1749 vdd.n1748 0.152939
R19305 vdd.n1748 vdd.n1747 0.152939
R19306 vdd.n1747 vdd.n1686 0.152939
R19307 vdd.n1691 vdd.n1686 0.152939
R19308 vdd.n1692 vdd.n1691 0.152939
R19309 vdd.n1693 vdd.n1692 0.152939
R19310 vdd.n1697 vdd.n1693 0.152939
R19311 vdd.n1698 vdd.n1697 0.152939
R19312 vdd.n1699 vdd.n1698 0.152939
R19313 vdd.n1700 vdd.n1699 0.152939
R19314 vdd.n1704 vdd.n1700 0.152939
R19315 vdd.n1705 vdd.n1704 0.152939
R19316 vdd.n1706 vdd.n1705 0.152939
R19317 vdd.n1707 vdd.n1706 0.152939
R19318 vdd.n1708 vdd.n1707 0.152939
R19319 vdd.n1708 vdd.n892 0.152939
R19320 vdd.n2037 vdd.n1612 0.152939
R19321 vdd.n1559 vdd.n1558 0.152939
R19322 vdd.n1559 vdd.n928 0.152939
R19323 vdd.n1574 vdd.n928 0.152939
R19324 vdd.n1575 vdd.n1574 0.152939
R19325 vdd.n1576 vdd.n1575 0.152939
R19326 vdd.n1576 vdd.n917 0.152939
R19327 vdd.n1591 vdd.n917 0.152939
R19328 vdd.n1592 vdd.n1591 0.152939
R19329 vdd.n1593 vdd.n1592 0.152939
R19330 vdd.n1593 vdd.n905 0.152939
R19331 vdd.n1610 vdd.n905 0.152939
R19332 vdd.n1611 vdd.n1610 0.152939
R19333 vdd.n2038 vdd.n1611 0.152939
R19334 vdd.n527 vdd.n524 0.152939
R19335 vdd.n528 vdd.n527 0.152939
R19336 vdd.n529 vdd.n528 0.152939
R19337 vdd.n530 vdd.n529 0.152939
R19338 vdd.n533 vdd.n530 0.152939
R19339 vdd.n534 vdd.n533 0.152939
R19340 vdd.n535 vdd.n534 0.152939
R19341 vdd.n536 vdd.n535 0.152939
R19342 vdd.n539 vdd.n536 0.152939
R19343 vdd.n540 vdd.n539 0.152939
R19344 vdd.n541 vdd.n540 0.152939
R19345 vdd.n542 vdd.n541 0.152939
R19346 vdd.n547 vdd.n542 0.152939
R19347 vdd.n548 vdd.n547 0.152939
R19348 vdd.n549 vdd.n548 0.152939
R19349 vdd.n550 vdd.n549 0.152939
R19350 vdd.n553 vdd.n550 0.152939
R19351 vdd.n554 vdd.n553 0.152939
R19352 vdd.n555 vdd.n554 0.152939
R19353 vdd.n556 vdd.n555 0.152939
R19354 vdd.n559 vdd.n556 0.152939
R19355 vdd.n560 vdd.n559 0.152939
R19356 vdd.n561 vdd.n560 0.152939
R19357 vdd.n562 vdd.n561 0.152939
R19358 vdd.n565 vdd.n562 0.152939
R19359 vdd.n566 vdd.n565 0.152939
R19360 vdd.n567 vdd.n566 0.152939
R19361 vdd.n568 vdd.n567 0.152939
R19362 vdd.n571 vdd.n568 0.152939
R19363 vdd.n572 vdd.n571 0.152939
R19364 vdd.n573 vdd.n572 0.152939
R19365 vdd.n574 vdd.n573 0.152939
R19366 vdd.n577 vdd.n574 0.152939
R19367 vdd.n578 vdd.n577 0.152939
R19368 vdd.n2853 vdd.n578 0.152939
R19369 vdd.n2853 vdd.n2852 0.152939
R19370 vdd.n2852 vdd.n2851 0.152939
R19371 vdd.n2851 vdd.n582 0.152939
R19372 vdd.n587 vdd.n582 0.152939
R19373 vdd.n588 vdd.n587 0.152939
R19374 vdd.n591 vdd.n588 0.152939
R19375 vdd.n592 vdd.n591 0.152939
R19376 vdd.n593 vdd.n592 0.152939
R19377 vdd.n594 vdd.n593 0.152939
R19378 vdd.n597 vdd.n594 0.152939
R19379 vdd.n598 vdd.n597 0.152939
R19380 vdd.n599 vdd.n598 0.152939
R19381 vdd.n600 vdd.n599 0.152939
R19382 vdd.n603 vdd.n600 0.152939
R19383 vdd.n604 vdd.n603 0.152939
R19384 vdd.n605 vdd.n604 0.152939
R19385 vdd.n2936 vdd.n518 0.152939
R19386 vdd.n2937 vdd.n508 0.152939
R19387 vdd.n2951 vdd.n508 0.152939
R19388 vdd.n2952 vdd.n2951 0.152939
R19389 vdd.n2953 vdd.n2952 0.152939
R19390 vdd.n2953 vdd.n496 0.152939
R19391 vdd.n2967 vdd.n496 0.152939
R19392 vdd.n2968 vdd.n2967 0.152939
R19393 vdd.n2969 vdd.n2968 0.152939
R19394 vdd.n2969 vdd.n484 0.152939
R19395 vdd.n2984 vdd.n484 0.152939
R19396 vdd.n2985 vdd.n2984 0.152939
R19397 vdd.n2986 vdd.n2985 0.152939
R19398 vdd.n2986 vdd.n310 0.152939
R19399 vdd.n320 vdd.n311 0.152939
R19400 vdd.n321 vdd.n320 0.152939
R19401 vdd.n322 vdd.n321 0.152939
R19402 vdd.n331 vdd.n322 0.152939
R19403 vdd.n332 vdd.n331 0.152939
R19404 vdd.n333 vdd.n332 0.152939
R19405 vdd.n334 vdd.n333 0.152939
R19406 vdd.n342 vdd.n334 0.152939
R19407 vdd.n343 vdd.n342 0.152939
R19408 vdd.n344 vdd.n343 0.152939
R19409 vdd.n345 vdd.n344 0.152939
R19410 vdd.n353 vdd.n345 0.152939
R19411 vdd.n3135 vdd.n353 0.152939
R19412 vdd.n3134 vdd.n354 0.152939
R19413 vdd.n357 vdd.n354 0.152939
R19414 vdd.n361 vdd.n357 0.152939
R19415 vdd.n362 vdd.n361 0.152939
R19416 vdd.n363 vdd.n362 0.152939
R19417 vdd.n364 vdd.n363 0.152939
R19418 vdd.n365 vdd.n364 0.152939
R19419 vdd.n369 vdd.n365 0.152939
R19420 vdd.n370 vdd.n369 0.152939
R19421 vdd.n371 vdd.n370 0.152939
R19422 vdd.n372 vdd.n371 0.152939
R19423 vdd.n376 vdd.n372 0.152939
R19424 vdd.n377 vdd.n376 0.152939
R19425 vdd.n378 vdd.n377 0.152939
R19426 vdd.n379 vdd.n378 0.152939
R19427 vdd.n383 vdd.n379 0.152939
R19428 vdd.n384 vdd.n383 0.152939
R19429 vdd.n385 vdd.n384 0.152939
R19430 vdd.n3100 vdd.n385 0.152939
R19431 vdd.n3100 vdd.n3099 0.152939
R19432 vdd.n3099 vdd.n3098 0.152939
R19433 vdd.n3098 vdd.n391 0.152939
R19434 vdd.n396 vdd.n391 0.152939
R19435 vdd.n397 vdd.n396 0.152939
R19436 vdd.n398 vdd.n397 0.152939
R19437 vdd.n402 vdd.n398 0.152939
R19438 vdd.n403 vdd.n402 0.152939
R19439 vdd.n404 vdd.n403 0.152939
R19440 vdd.n405 vdd.n404 0.152939
R19441 vdd.n409 vdd.n405 0.152939
R19442 vdd.n410 vdd.n409 0.152939
R19443 vdd.n411 vdd.n410 0.152939
R19444 vdd.n412 vdd.n411 0.152939
R19445 vdd.n416 vdd.n412 0.152939
R19446 vdd.n417 vdd.n416 0.152939
R19447 vdd.n418 vdd.n417 0.152939
R19448 vdd.n419 vdd.n418 0.152939
R19449 vdd.n423 vdd.n419 0.152939
R19450 vdd.n424 vdd.n423 0.152939
R19451 vdd.n425 vdd.n424 0.152939
R19452 vdd.n3061 vdd.n425 0.152939
R19453 vdd.n3061 vdd.n3060 0.152939
R19454 vdd.n3060 vdd.n3059 0.152939
R19455 vdd.n3059 vdd.n431 0.152939
R19456 vdd.n436 vdd.n431 0.152939
R19457 vdd.n437 vdd.n436 0.152939
R19458 vdd.n438 vdd.n437 0.152939
R19459 vdd.n442 vdd.n438 0.152939
R19460 vdd.n443 vdd.n442 0.152939
R19461 vdd.n444 vdd.n443 0.152939
R19462 vdd.n445 vdd.n444 0.152939
R19463 vdd.n449 vdd.n445 0.152939
R19464 vdd.n450 vdd.n449 0.152939
R19465 vdd.n451 vdd.n450 0.152939
R19466 vdd.n452 vdd.n451 0.152939
R19467 vdd.n456 vdd.n452 0.152939
R19468 vdd.n457 vdd.n456 0.152939
R19469 vdd.n458 vdd.n457 0.152939
R19470 vdd.n459 vdd.n458 0.152939
R19471 vdd.n463 vdd.n459 0.152939
R19472 vdd.n464 vdd.n463 0.152939
R19473 vdd.n465 vdd.n464 0.152939
R19474 vdd.n3017 vdd.n465 0.152939
R19475 vdd.n2944 vdd.n2943 0.152939
R19476 vdd.n2945 vdd.n2944 0.152939
R19477 vdd.n2945 vdd.n502 0.152939
R19478 vdd.n2959 vdd.n502 0.152939
R19479 vdd.n2960 vdd.n2959 0.152939
R19480 vdd.n2961 vdd.n2960 0.152939
R19481 vdd.n2961 vdd.n489 0.152939
R19482 vdd.n2975 vdd.n489 0.152939
R19483 vdd.n2976 vdd.n2975 0.152939
R19484 vdd.n2977 vdd.n2976 0.152939
R19485 vdd.n2977 vdd.n477 0.152939
R19486 vdd.n2992 vdd.n477 0.152939
R19487 vdd.n2993 vdd.n2992 0.152939
R19488 vdd.n2994 vdd.n2993 0.152939
R19489 vdd.n2994 vdd.n475 0.152939
R19490 vdd.n2998 vdd.n475 0.152939
R19491 vdd.n2999 vdd.n2998 0.152939
R19492 vdd.n3000 vdd.n2999 0.152939
R19493 vdd.n3000 vdd.n472 0.152939
R19494 vdd.n3004 vdd.n472 0.152939
R19495 vdd.n3005 vdd.n3004 0.152939
R19496 vdd.n3006 vdd.n3005 0.152939
R19497 vdd.n3006 vdd.n469 0.152939
R19498 vdd.n3010 vdd.n469 0.152939
R19499 vdd.n3011 vdd.n3010 0.152939
R19500 vdd.n3012 vdd.n3011 0.152939
R19501 vdd.n3012 vdd.n466 0.152939
R19502 vdd.n3016 vdd.n466 0.152939
R19503 vdd.n2806 vdd.n514 0.152939
R19504 vdd.n2049 vdd.n895 0.152939
R19505 vdd.n1219 vdd.n1218 0.152939
R19506 vdd.n1220 vdd.n1219 0.152939
R19507 vdd.n1220 vdd.n969 0.152939
R19508 vdd.n1234 vdd.n969 0.152939
R19509 vdd.n1235 vdd.n1234 0.152939
R19510 vdd.n1236 vdd.n1235 0.152939
R19511 vdd.n1236 vdd.n956 0.152939
R19512 vdd.n1250 vdd.n956 0.152939
R19513 vdd.n1251 vdd.n1250 0.152939
R19514 vdd.n1252 vdd.n1251 0.152939
R19515 vdd.n1252 vdd.n945 0.152939
R19516 vdd.n1267 vdd.n945 0.152939
R19517 vdd.n1268 vdd.n1267 0.152939
R19518 vdd.n1269 vdd.n1268 0.152939
R19519 vdd.n1269 vdd.n934 0.152939
R19520 vdd.n1565 vdd.n934 0.152939
R19521 vdd.n1566 vdd.n1565 0.152939
R19522 vdd.n1567 vdd.n1566 0.152939
R19523 vdd.n1567 vdd.n922 0.152939
R19524 vdd.n1582 vdd.n922 0.152939
R19525 vdd.n1583 vdd.n1582 0.152939
R19526 vdd.n1584 vdd.n1583 0.152939
R19527 vdd.n1584 vdd.n912 0.152939
R19528 vdd.n1599 vdd.n912 0.152939
R19529 vdd.n1600 vdd.n1599 0.152939
R19530 vdd.n1603 vdd.n1600 0.152939
R19531 vdd.n1603 vdd.n1602 0.152939
R19532 vdd.n1602 vdd.n1601 0.152939
R19533 vdd.n1211 vdd.n985 0.152939
R19534 vdd.n1207 vdd.n985 0.152939
R19535 vdd.n1207 vdd.n1206 0.152939
R19536 vdd.n1206 vdd.n1205 0.152939
R19537 vdd.n1205 vdd.n990 0.152939
R19538 vdd.n1201 vdd.n990 0.152939
R19539 vdd.n1201 vdd.n1200 0.152939
R19540 vdd.n1200 vdd.n1199 0.152939
R19541 vdd.n1199 vdd.n998 0.152939
R19542 vdd.n1195 vdd.n998 0.152939
R19543 vdd.n1195 vdd.n1194 0.152939
R19544 vdd.n1194 vdd.n1193 0.152939
R19545 vdd.n1193 vdd.n1006 0.152939
R19546 vdd.n1189 vdd.n1006 0.152939
R19547 vdd.n1189 vdd.n1188 0.152939
R19548 vdd.n1188 vdd.n1187 0.152939
R19549 vdd.n1187 vdd.n1014 0.152939
R19550 vdd.n1183 vdd.n1014 0.152939
R19551 vdd.n1183 vdd.n1182 0.152939
R19552 vdd.n1182 vdd.n1181 0.152939
R19553 vdd.n1181 vdd.n1024 0.152939
R19554 vdd.n1177 vdd.n1024 0.152939
R19555 vdd.n1177 vdd.n1176 0.152939
R19556 vdd.n1176 vdd.n1175 0.152939
R19557 vdd.n1175 vdd.n1032 0.152939
R19558 vdd.n1171 vdd.n1032 0.152939
R19559 vdd.n1171 vdd.n1170 0.152939
R19560 vdd.n1170 vdd.n1169 0.152939
R19561 vdd.n1169 vdd.n1040 0.152939
R19562 vdd.n1165 vdd.n1040 0.152939
R19563 vdd.n1165 vdd.n1164 0.152939
R19564 vdd.n1164 vdd.n1163 0.152939
R19565 vdd.n1163 vdd.n1048 0.152939
R19566 vdd.n1159 vdd.n1048 0.152939
R19567 vdd.n1159 vdd.n1158 0.152939
R19568 vdd.n1158 vdd.n1157 0.152939
R19569 vdd.n1157 vdd.n1056 0.152939
R19570 vdd.n1153 vdd.n1056 0.152939
R19571 vdd.n1153 vdd.n1152 0.152939
R19572 vdd.n1152 vdd.n1151 0.152939
R19573 vdd.n1151 vdd.n1064 0.152939
R19574 vdd.n1071 vdd.n1064 0.152939
R19575 vdd.n1141 vdd.n1071 0.152939
R19576 vdd.n1141 vdd.n1140 0.152939
R19577 vdd.n1140 vdd.n1139 0.152939
R19578 vdd.n1139 vdd.n1072 0.152939
R19579 vdd.n1135 vdd.n1072 0.152939
R19580 vdd.n1135 vdd.n1134 0.152939
R19581 vdd.n1134 vdd.n1133 0.152939
R19582 vdd.n1133 vdd.n1079 0.152939
R19583 vdd.n1129 vdd.n1079 0.152939
R19584 vdd.n1129 vdd.n1128 0.152939
R19585 vdd.n1128 vdd.n1127 0.152939
R19586 vdd.n1127 vdd.n1087 0.152939
R19587 vdd.n1123 vdd.n1087 0.152939
R19588 vdd.n1123 vdd.n1122 0.152939
R19589 vdd.n1122 vdd.n1121 0.152939
R19590 vdd.n1121 vdd.n1095 0.152939
R19591 vdd.n1117 vdd.n1095 0.152939
R19592 vdd.n1117 vdd.n1116 0.152939
R19593 vdd.n1116 vdd.n1115 0.152939
R19594 vdd.n1115 vdd.n1103 0.152939
R19595 vdd.n1103 vdd.n980 0.152939
R19596 vdd.n1212 vdd.n975 0.152939
R19597 vdd.n1226 vdd.n975 0.152939
R19598 vdd.n1227 vdd.n1226 0.152939
R19599 vdd.n1228 vdd.n1227 0.152939
R19600 vdd.n1228 vdd.n963 0.152939
R19601 vdd.n1242 vdd.n963 0.152939
R19602 vdd.n1243 vdd.n1242 0.152939
R19603 vdd.n1244 vdd.n1243 0.152939
R19604 vdd.n1244 vdd.n951 0.152939
R19605 vdd.n1259 vdd.n951 0.152939
R19606 vdd.n1260 vdd.n1259 0.152939
R19607 vdd.n1261 vdd.n1260 0.152939
R19608 vdd.n1261 vdd.n940 0.152939
R19609 vdd.n1558 vdd.n1557 0.145814
R19610 vdd.n3167 vdd.n310 0.145814
R19611 vdd.n3167 vdd.n311 0.145814
R19612 vdd.n1557 vdd.n940 0.145814
R19613 vdd.n2027 vdd.n1612 0.110256
R19614 vdd.n2737 vdd.n518 0.110256
R19615 vdd.n2806 vdd.n2805 0.110256
R19616 vdd.n2050 vdd.n2049 0.110256
R19617 vdd.n2027 vdd.n1813 0.0431829
R19618 vdd.n2050 vdd.n892 0.0431829
R19619 vdd.n2737 vdd.n524 0.0431829
R19620 vdd.n2805 vdd.n605 0.0431829
R19621 vdd vdd.n28 0.00833333
R19622 a_n6308_8799.n143 a_n6308_8799.t83 490.524
R19623 a_n6308_8799.n154 a_n6308_8799.t90 490.524
R19624 a_n6308_8799.n166 a_n6308_8799.t100 490.524
R19625 a_n6308_8799.n109 a_n6308_8799.t60 490.524
R19626 a_n6308_8799.n120 a_n6308_8799.t66 490.524
R19627 a_n6308_8799.n132 a_n6308_8799.t99 490.524
R19628 a_n6308_8799.n30 a_n6308_8799.t69 484.3
R19629 a_n6308_8799.n149 a_n6308_8799.t68 464.166
R19630 a_n6308_8799.n148 a_n6308_8799.t50 464.166
R19631 a_n6308_8799.n139 a_n6308_8799.t96 464.166
R19632 a_n6308_8799.n147 a_n6308_8799.t70 464.166
R19633 a_n6308_8799.n146 a_n6308_8799.t55 464.166
R19634 a_n6308_8799.n140 a_n6308_8799.t98 464.166
R19635 a_n6308_8799.n145 a_n6308_8799.t80 464.166
R19636 a_n6308_8799.n144 a_n6308_8799.t78 464.166
R19637 a_n6308_8799.n141 a_n6308_8799.t39 464.166
R19638 a_n6308_8799.n142 a_n6308_8799.t84 464.166
R19639 a_n6308_8799.n39 a_n6308_8799.t74 484.3
R19640 a_n6308_8799.n160 a_n6308_8799.t73 464.166
R19641 a_n6308_8799.n159 a_n6308_8799.t62 464.166
R19642 a_n6308_8799.n150 a_n6308_8799.t104 464.166
R19643 a_n6308_8799.n158 a_n6308_8799.t77 464.166
R19644 a_n6308_8799.n157 a_n6308_8799.t63 464.166
R19645 a_n6308_8799.n151 a_n6308_8799.t36 464.166
R19646 a_n6308_8799.n156 a_n6308_8799.t89 464.166
R19647 a_n6308_8799.n155 a_n6308_8799.t88 464.166
R19648 a_n6308_8799.n152 a_n6308_8799.t46 464.166
R19649 a_n6308_8799.n153 a_n6308_8799.t91 464.166
R19650 a_n6308_8799.n48 a_n6308_8799.t106 484.3
R19651 a_n6308_8799.n172 a_n6308_8799.t48 464.166
R19652 a_n6308_8799.n171 a_n6308_8799.t75 464.166
R19653 a_n6308_8799.n162 a_n6308_8799.t38 464.166
R19654 a_n6308_8799.n170 a_n6308_8799.t93 464.166
R19655 a_n6308_8799.n169 a_n6308_8799.t54 464.166
R19656 a_n6308_8799.n163 a_n6308_8799.t81 464.166
R19657 a_n6308_8799.n168 a_n6308_8799.t40 464.166
R19658 a_n6308_8799.n167 a_n6308_8799.t58 464.166
R19659 a_n6308_8799.n164 a_n6308_8799.t102 464.166
R19660 a_n6308_8799.n165 a_n6308_8799.t86 464.166
R19661 a_n6308_8799.n108 a_n6308_8799.t61 464.166
R19662 a_n6308_8799.n107 a_n6308_8799.t85 464.166
R19663 a_n6308_8799.n110 a_n6308_8799.t37 464.166
R19664 a_n6308_8799.n106 a_n6308_8799.t57 464.166
R19665 a_n6308_8799.n111 a_n6308_8799.t72 464.166
R19666 a_n6308_8799.n112 a_n6308_8799.t97 464.166
R19667 a_n6308_8799.n105 a_n6308_8799.t44 464.166
R19668 a_n6308_8799.n113 a_n6308_8799.t56 464.166
R19669 a_n6308_8799.n104 a_n6308_8799.t95 464.166
R19670 a_n6308_8799.n114 a_n6308_8799.t43 464.166
R19671 a_n6308_8799.n119 a_n6308_8799.t67 464.166
R19672 a_n6308_8799.n118 a_n6308_8799.t92 464.166
R19673 a_n6308_8799.n121 a_n6308_8799.t45 464.166
R19674 a_n6308_8799.n117 a_n6308_8799.t65 464.166
R19675 a_n6308_8799.n122 a_n6308_8799.t79 464.166
R19676 a_n6308_8799.n123 a_n6308_8799.t105 464.166
R19677 a_n6308_8799.n116 a_n6308_8799.t53 464.166
R19678 a_n6308_8799.n124 a_n6308_8799.t64 464.166
R19679 a_n6308_8799.n115 a_n6308_8799.t101 464.166
R19680 a_n6308_8799.n125 a_n6308_8799.t49 464.166
R19681 a_n6308_8799.n131 a_n6308_8799.t87 464.166
R19682 a_n6308_8799.n130 a_n6308_8799.t103 464.166
R19683 a_n6308_8799.n133 a_n6308_8799.t71 464.166
R19684 a_n6308_8799.n129 a_n6308_8799.t41 464.166
R19685 a_n6308_8799.n134 a_n6308_8799.t82 464.166
R19686 a_n6308_8799.n135 a_n6308_8799.t52 464.166
R19687 a_n6308_8799.n128 a_n6308_8799.t94 464.166
R19688 a_n6308_8799.n136 a_n6308_8799.t59 464.166
R19689 a_n6308_8799.n127 a_n6308_8799.t76 464.166
R19690 a_n6308_8799.n137 a_n6308_8799.t47 464.166
R19691 a_n6308_8799.n38 a_n6308_8799.n37 75.3623
R19692 a_n6308_8799.n36 a_n6308_8799.n20 70.3058
R19693 a_n6308_8799.n20 a_n6308_8799.n35 70.1674
R19694 a_n6308_8799.n35 a_n6308_8799.n140 20.9683
R19695 a_n6308_8799.n34 a_n6308_8799.n21 75.0448
R19696 a_n6308_8799.n146 a_n6308_8799.n34 11.2134
R19697 a_n6308_8799.n33 a_n6308_8799.n21 80.4688
R19698 a_n6308_8799.n23 a_n6308_8799.n32 74.73
R19699 a_n6308_8799.n31 a_n6308_8799.n23 70.1674
R19700 a_n6308_8799.n149 a_n6308_8799.n31 20.9683
R19701 a_n6308_8799.n22 a_n6308_8799.n30 70.5844
R19702 a_n6308_8799.n47 a_n6308_8799.n46 75.3623
R19703 a_n6308_8799.n45 a_n6308_8799.n16 70.3058
R19704 a_n6308_8799.n16 a_n6308_8799.n44 70.1674
R19705 a_n6308_8799.n44 a_n6308_8799.n151 20.9683
R19706 a_n6308_8799.n43 a_n6308_8799.n17 75.0448
R19707 a_n6308_8799.n157 a_n6308_8799.n43 11.2134
R19708 a_n6308_8799.n42 a_n6308_8799.n17 80.4688
R19709 a_n6308_8799.n19 a_n6308_8799.n41 74.73
R19710 a_n6308_8799.n40 a_n6308_8799.n19 70.1674
R19711 a_n6308_8799.n160 a_n6308_8799.n40 20.9683
R19712 a_n6308_8799.n18 a_n6308_8799.n39 70.5844
R19713 a_n6308_8799.n56 a_n6308_8799.n55 75.3623
R19714 a_n6308_8799.n54 a_n6308_8799.n12 70.3058
R19715 a_n6308_8799.n12 a_n6308_8799.n53 70.1674
R19716 a_n6308_8799.n53 a_n6308_8799.n163 20.9683
R19717 a_n6308_8799.n52 a_n6308_8799.n13 75.0448
R19718 a_n6308_8799.n169 a_n6308_8799.n52 11.2134
R19719 a_n6308_8799.n51 a_n6308_8799.n13 80.4688
R19720 a_n6308_8799.n15 a_n6308_8799.n50 74.73
R19721 a_n6308_8799.n49 a_n6308_8799.n15 70.1674
R19722 a_n6308_8799.n172 a_n6308_8799.n49 20.9683
R19723 a_n6308_8799.n14 a_n6308_8799.n48 70.5844
R19724 a_n6308_8799.n8 a_n6308_8799.n65 70.5844
R19725 a_n6308_8799.n64 a_n6308_8799.n9 70.1674
R19726 a_n6308_8799.n64 a_n6308_8799.n104 20.9683
R19727 a_n6308_8799.n9 a_n6308_8799.n63 74.73
R19728 a_n6308_8799.n113 a_n6308_8799.n63 11.843
R19729 a_n6308_8799.n62 a_n6308_8799.n10 80.4688
R19730 a_n6308_8799.n62 a_n6308_8799.n105 0.365327
R19731 a_n6308_8799.n10 a_n6308_8799.n61 75.0448
R19732 a_n6308_8799.n60 a_n6308_8799.n11 70.1674
R19733 a_n6308_8799.n60 a_n6308_8799.n106 20.9683
R19734 a_n6308_8799.n11 a_n6308_8799.n59 70.3058
R19735 a_n6308_8799.n110 a_n6308_8799.n59 20.6913
R19736 a_n6308_8799.n58 a_n6308_8799.n57 75.3623
R19737 a_n6308_8799.n4 a_n6308_8799.n74 70.5844
R19738 a_n6308_8799.n73 a_n6308_8799.n5 70.1674
R19739 a_n6308_8799.n73 a_n6308_8799.n115 20.9683
R19740 a_n6308_8799.n5 a_n6308_8799.n72 74.73
R19741 a_n6308_8799.n124 a_n6308_8799.n72 11.843
R19742 a_n6308_8799.n71 a_n6308_8799.n6 80.4688
R19743 a_n6308_8799.n71 a_n6308_8799.n116 0.365327
R19744 a_n6308_8799.n6 a_n6308_8799.n70 75.0448
R19745 a_n6308_8799.n69 a_n6308_8799.n7 70.1674
R19746 a_n6308_8799.n69 a_n6308_8799.n117 20.9683
R19747 a_n6308_8799.n7 a_n6308_8799.n68 70.3058
R19748 a_n6308_8799.n121 a_n6308_8799.n68 20.6913
R19749 a_n6308_8799.n67 a_n6308_8799.n66 75.3623
R19750 a_n6308_8799.n0 a_n6308_8799.n83 70.5844
R19751 a_n6308_8799.n82 a_n6308_8799.n1 70.1674
R19752 a_n6308_8799.n82 a_n6308_8799.n127 20.9683
R19753 a_n6308_8799.n1 a_n6308_8799.n81 74.73
R19754 a_n6308_8799.n136 a_n6308_8799.n81 11.843
R19755 a_n6308_8799.n80 a_n6308_8799.n2 80.4688
R19756 a_n6308_8799.n80 a_n6308_8799.n128 0.365327
R19757 a_n6308_8799.n2 a_n6308_8799.n79 75.0448
R19758 a_n6308_8799.n78 a_n6308_8799.n3 70.1674
R19759 a_n6308_8799.n78 a_n6308_8799.n129 20.9683
R19760 a_n6308_8799.n3 a_n6308_8799.n77 70.3058
R19761 a_n6308_8799.n133 a_n6308_8799.n77 20.6913
R19762 a_n6308_8799.n76 a_n6308_8799.n75 75.3623
R19763 a_n6308_8799.n179 a_n6308_8799.n25 98.9632
R19764 a_n6308_8799.n24 a_n6308_8799.n84 98.9631
R19765 a_n6308_8799.n25 a_n6308_8799.n177 98.6055
R19766 a_n6308_8799.n25 a_n6308_8799.n178 98.6055
R19767 a_n6308_8799.n24 a_n6308_8799.n85 98.6055
R19768 a_n6308_8799.n24 a_n6308_8799.n86 98.6055
R19769 a_n6308_8799.n89 a_n6308_8799.n87 81.4626
R19770 a_n6308_8799.n97 a_n6308_8799.n95 81.4626
R19771 a_n6308_8799.n93 a_n6308_8799.n91 81.4626
R19772 a_n6308_8799.n100 a_n6308_8799.n99 80.9324
R19773 a_n6308_8799.n102 a_n6308_8799.n101 80.9324
R19774 a_n6308_8799.n29 a_n6308_8799.n103 80.9324
R19775 a_n6308_8799.n28 a_n6308_8799.n90 80.9324
R19776 a_n6308_8799.n89 a_n6308_8799.n88 80.9324
R19777 a_n6308_8799.n97 a_n6308_8799.n96 80.9324
R19778 a_n6308_8799.n27 a_n6308_8799.n98 80.9324
R19779 a_n6308_8799.n26 a_n6308_8799.n94 80.9324
R19780 a_n6308_8799.n93 a_n6308_8799.n92 80.9324
R19781 a_n6308_8799.n31 a_n6308_8799.n148 20.9683
R19782 a_n6308_8799.n147 a_n6308_8799.n146 48.2005
R19783 a_n6308_8799.n145 a_n6308_8799.n35 20.9683
R19784 a_n6308_8799.n142 a_n6308_8799.n141 48.2005
R19785 a_n6308_8799.n40 a_n6308_8799.n159 20.9683
R19786 a_n6308_8799.n158 a_n6308_8799.n157 48.2005
R19787 a_n6308_8799.n156 a_n6308_8799.n44 20.9683
R19788 a_n6308_8799.n153 a_n6308_8799.n152 48.2005
R19789 a_n6308_8799.n49 a_n6308_8799.n171 20.9683
R19790 a_n6308_8799.n170 a_n6308_8799.n169 48.2005
R19791 a_n6308_8799.n168 a_n6308_8799.n53 20.9683
R19792 a_n6308_8799.n165 a_n6308_8799.n164 48.2005
R19793 a_n6308_8799.n108 a_n6308_8799.n107 48.2005
R19794 a_n6308_8799.n111 a_n6308_8799.n60 20.9683
R19795 a_n6308_8799.n112 a_n6308_8799.n105 48.2005
R19796 a_n6308_8799.n114 a_n6308_8799.n64 20.9683
R19797 a_n6308_8799.n119 a_n6308_8799.n118 48.2005
R19798 a_n6308_8799.n122 a_n6308_8799.n69 20.9683
R19799 a_n6308_8799.n123 a_n6308_8799.n116 48.2005
R19800 a_n6308_8799.n125 a_n6308_8799.n73 20.9683
R19801 a_n6308_8799.n131 a_n6308_8799.n130 48.2005
R19802 a_n6308_8799.n134 a_n6308_8799.n78 20.9683
R19803 a_n6308_8799.n135 a_n6308_8799.n128 48.2005
R19804 a_n6308_8799.n137 a_n6308_8799.n82 20.9683
R19805 a_n6308_8799.n33 a_n6308_8799.n139 47.835
R19806 a_n6308_8799.n36 a_n6308_8799.n144 20.6913
R19807 a_n6308_8799.n42 a_n6308_8799.n150 47.835
R19808 a_n6308_8799.n45 a_n6308_8799.n155 20.6913
R19809 a_n6308_8799.n51 a_n6308_8799.n162 47.835
R19810 a_n6308_8799.n54 a_n6308_8799.n167 20.6913
R19811 a_n6308_8799.n106 a_n6308_8799.n59 21.4216
R19812 a_n6308_8799.n117 a_n6308_8799.n68 21.4216
R19813 a_n6308_8799.n129 a_n6308_8799.n77 21.4216
R19814 a_n6308_8799.t42 a_n6308_8799.n65 484.3
R19815 a_n6308_8799.t51 a_n6308_8799.n74 484.3
R19816 a_n6308_8799.t107 a_n6308_8799.n83 484.3
R19817 a_n6308_8799.n58 a_n6308_8799.n109 45.0871
R19818 a_n6308_8799.n67 a_n6308_8799.n120 45.0871
R19819 a_n6308_8799.n76 a_n6308_8799.n132 45.0871
R19820 a_n6308_8799.n38 a_n6308_8799.n143 45.0871
R19821 a_n6308_8799.n47 a_n6308_8799.n154 45.0871
R19822 a_n6308_8799.n56 a_n6308_8799.n166 45.0871
R19823 a_n6308_8799.n100 a_n6308_8799.n27 34.3237
R19824 a_n6308_8799.n32 a_n6308_8799.n139 11.843
R19825 a_n6308_8799.n144 a_n6308_8799.n37 36.139
R19826 a_n6308_8799.n41 a_n6308_8799.n150 11.843
R19827 a_n6308_8799.n155 a_n6308_8799.n46 36.139
R19828 a_n6308_8799.n50 a_n6308_8799.n162 11.843
R19829 a_n6308_8799.n167 a_n6308_8799.n55 36.139
R19830 a_n6308_8799.n110 a_n6308_8799.n57 36.139
R19831 a_n6308_8799.n104 a_n6308_8799.n63 34.4824
R19832 a_n6308_8799.n121 a_n6308_8799.n66 36.139
R19833 a_n6308_8799.n115 a_n6308_8799.n72 34.4824
R19834 a_n6308_8799.n133 a_n6308_8799.n75 36.139
R19835 a_n6308_8799.n127 a_n6308_8799.n81 34.4824
R19836 a_n6308_8799.n34 a_n6308_8799.n140 35.3134
R19837 a_n6308_8799.n43 a_n6308_8799.n151 35.3134
R19838 a_n6308_8799.n52 a_n6308_8799.n163 35.3134
R19839 a_n6308_8799.n61 a_n6308_8799.n111 35.3134
R19840 a_n6308_8799.n112 a_n6308_8799.n61 11.2134
R19841 a_n6308_8799.n70 a_n6308_8799.n122 35.3134
R19842 a_n6308_8799.n123 a_n6308_8799.n70 11.2134
R19843 a_n6308_8799.n79 a_n6308_8799.n134 35.3134
R19844 a_n6308_8799.n135 a_n6308_8799.n79 11.2134
R19845 a_n6308_8799.n148 a_n6308_8799.n32 34.4824
R19846 a_n6308_8799.n37 a_n6308_8799.n141 10.5784
R19847 a_n6308_8799.n159 a_n6308_8799.n41 34.4824
R19848 a_n6308_8799.n46 a_n6308_8799.n152 10.5784
R19849 a_n6308_8799.n171 a_n6308_8799.n50 34.4824
R19850 a_n6308_8799.n55 a_n6308_8799.n164 10.5784
R19851 a_n6308_8799.n57 a_n6308_8799.n107 10.5784
R19852 a_n6308_8799.n66 a_n6308_8799.n118 10.5784
R19853 a_n6308_8799.n75 a_n6308_8799.n130 10.5784
R19854 a_n6308_8799.n143 a_n6308_8799.n142 14.1472
R19855 a_n6308_8799.n154 a_n6308_8799.n153 14.1472
R19856 a_n6308_8799.n166 a_n6308_8799.n165 14.1472
R19857 a_n6308_8799.n109 a_n6308_8799.n108 14.1472
R19858 a_n6308_8799.n120 a_n6308_8799.n119 14.1472
R19859 a_n6308_8799.n132 a_n6308_8799.n131 14.1472
R19860 a_n6308_8799.n175 a_n6308_8799.n29 12.3339
R19861 a_n6308_8799.n176 a_n6308_8799.n175 11.4887
R19862 a_n6308_8799.n161 a_n6308_8799.n22 9.01755
R19863 a_n6308_8799.n126 a_n6308_8799.n8 9.01755
R19864 a_n6308_8799.n174 a_n6308_8799.n138 6.93972
R19865 a_n6308_8799.n174 a_n6308_8799.n173 6.44309
R19866 a_n6308_8799.n161 a_n6308_8799.n18 4.90959
R19867 a_n6308_8799.n173 a_n6308_8799.n14 4.90959
R19868 a_n6308_8799.n126 a_n6308_8799.n4 4.90959
R19869 a_n6308_8799.n138 a_n6308_8799.n0 4.90959
R19870 a_n6308_8799.n173 a_n6308_8799.n161 4.10845
R19871 a_n6308_8799.n138 a_n6308_8799.n126 4.10845
R19872 a_n6308_8799.n177 a_n6308_8799.t16 3.61217
R19873 a_n6308_8799.n177 a_n6308_8799.t20 3.61217
R19874 a_n6308_8799.n178 a_n6308_8799.t2 3.61217
R19875 a_n6308_8799.n178 a_n6308_8799.t6 3.61217
R19876 a_n6308_8799.n84 a_n6308_8799.t5 3.61217
R19877 a_n6308_8799.n84 a_n6308_8799.t8 3.61217
R19878 a_n6308_8799.n85 a_n6308_8799.t7 3.61217
R19879 a_n6308_8799.n85 a_n6308_8799.t29 3.61217
R19880 a_n6308_8799.n86 a_n6308_8799.t21 3.61217
R19881 a_n6308_8799.n86 a_n6308_8799.t22 3.61217
R19882 a_n6308_8799.t1 a_n6308_8799.n179 3.61217
R19883 a_n6308_8799.n179 a_n6308_8799.t32 3.61217
R19884 a_n6308_8799.n175 a_n6308_8799.n174 3.4105
R19885 a_n6308_8799.n99 a_n6308_8799.t18 2.82907
R19886 a_n6308_8799.n99 a_n6308_8799.t0 2.82907
R19887 a_n6308_8799.n101 a_n6308_8799.t19 2.82907
R19888 a_n6308_8799.n101 a_n6308_8799.t25 2.82907
R19889 a_n6308_8799.n103 a_n6308_8799.t10 2.82907
R19890 a_n6308_8799.n103 a_n6308_8799.t13 2.82907
R19891 a_n6308_8799.n90 a_n6308_8799.t26 2.82907
R19892 a_n6308_8799.n90 a_n6308_8799.t3 2.82907
R19893 a_n6308_8799.n88 a_n6308_8799.t15 2.82907
R19894 a_n6308_8799.n88 a_n6308_8799.t34 2.82907
R19895 a_n6308_8799.n87 a_n6308_8799.t9 2.82907
R19896 a_n6308_8799.n87 a_n6308_8799.t11 2.82907
R19897 a_n6308_8799.n95 a_n6308_8799.t12 2.82907
R19898 a_n6308_8799.n95 a_n6308_8799.t31 2.82907
R19899 a_n6308_8799.n96 a_n6308_8799.t24 2.82907
R19900 a_n6308_8799.n96 a_n6308_8799.t17 2.82907
R19901 a_n6308_8799.n98 a_n6308_8799.t23 2.82907
R19902 a_n6308_8799.n98 a_n6308_8799.t4 2.82907
R19903 a_n6308_8799.n94 a_n6308_8799.t33 2.82907
R19904 a_n6308_8799.n94 a_n6308_8799.t30 2.82907
R19905 a_n6308_8799.n92 a_n6308_8799.t28 2.82907
R19906 a_n6308_8799.n92 a_n6308_8799.t14 2.82907
R19907 a_n6308_8799.n91 a_n6308_8799.t27 2.82907
R19908 a_n6308_8799.n91 a_n6308_8799.t35 2.82907
R19909 a_n6308_8799.n30 a_n6308_8799.n149 22.3251
R19910 a_n6308_8799.n39 a_n6308_8799.n160 22.3251
R19911 a_n6308_8799.n48 a_n6308_8799.n172 22.3251
R19912 a_n6308_8799.n65 a_n6308_8799.n114 22.3251
R19913 a_n6308_8799.n74 a_n6308_8799.n125 22.3251
R19914 a_n6308_8799.n83 a_n6308_8799.n137 22.3251
R19915 a_n6308_8799.n33 a_n6308_8799.n147 0.365327
R19916 a_n6308_8799.n145 a_n6308_8799.n36 21.4216
R19917 a_n6308_8799.n42 a_n6308_8799.n158 0.365327
R19918 a_n6308_8799.n156 a_n6308_8799.n45 21.4216
R19919 a_n6308_8799.n51 a_n6308_8799.n170 0.365327
R19920 a_n6308_8799.n168 a_n6308_8799.n54 21.4216
R19921 a_n6308_8799.n113 a_n6308_8799.n62 47.835
R19922 a_n6308_8799.n124 a_n6308_8799.n71 47.835
R19923 a_n6308_8799.n136 a_n6308_8799.n80 47.835
R19924 a_n6308_8799.n176 a_n6308_8799.n24 31.5519
R19925 a_n6308_8799.n25 a_n6308_8799.n176 17.6132
R19926 a_n6308_8799.n23 a_n6308_8799.n21 0.758076
R19927 a_n6308_8799.n21 a_n6308_8799.n20 0.758076
R19928 a_n6308_8799.n38 a_n6308_8799.n20 0.758076
R19929 a_n6308_8799.n19 a_n6308_8799.n17 0.758076
R19930 a_n6308_8799.n17 a_n6308_8799.n16 0.758076
R19931 a_n6308_8799.n47 a_n6308_8799.n16 0.758076
R19932 a_n6308_8799.n15 a_n6308_8799.n13 0.758076
R19933 a_n6308_8799.n13 a_n6308_8799.n12 0.758076
R19934 a_n6308_8799.n56 a_n6308_8799.n12 0.758076
R19935 a_n6308_8799.n11 a_n6308_8799.n10 0.758076
R19936 a_n6308_8799.n10 a_n6308_8799.n9 0.758076
R19937 a_n6308_8799.n9 a_n6308_8799.n8 0.758076
R19938 a_n6308_8799.n7 a_n6308_8799.n6 0.758076
R19939 a_n6308_8799.n6 a_n6308_8799.n5 0.758076
R19940 a_n6308_8799.n5 a_n6308_8799.n4 0.758076
R19941 a_n6308_8799.n3 a_n6308_8799.n2 0.758076
R19942 a_n6308_8799.n2 a_n6308_8799.n1 0.758076
R19943 a_n6308_8799.n1 a_n6308_8799.n0 0.758076
R19944 a_n6308_8799.n76 a_n6308_8799.n3 0.568682
R19945 a_n6308_8799.n67 a_n6308_8799.n7 0.568682
R19946 a_n6308_8799.n58 a_n6308_8799.n11 0.568682
R19947 a_n6308_8799.n15 a_n6308_8799.n14 0.568682
R19948 a_n6308_8799.n19 a_n6308_8799.n18 0.568682
R19949 a_n6308_8799.n23 a_n6308_8799.n22 0.568682
R19950 a_n6308_8799.n26 a_n6308_8799.n93 0.530672
R19951 a_n6308_8799.n27 a_n6308_8799.n97 0.530672
R19952 a_n6308_8799.n28 a_n6308_8799.n89 0.530672
R19953 a_n6308_8799.n29 a_n6308_8799.n102 0.530672
R19954 a_n6308_8799.n102 a_n6308_8799.n100 0.530672
R19955 a_n6308_8799.n29 a_n6308_8799.n28 0.530672
R19956 a_n6308_8799.n27 a_n6308_8799.n26 0.530672
R19957 CSoutput.n19 CSoutput.t161 184.661
R19958 CSoutput.n78 CSoutput.n77 165.8
R19959 CSoutput.n76 CSoutput.n0 165.8
R19960 CSoutput.n75 CSoutput.n74 165.8
R19961 CSoutput.n73 CSoutput.n72 165.8
R19962 CSoutput.n71 CSoutput.n2 165.8
R19963 CSoutput.n69 CSoutput.n68 165.8
R19964 CSoutput.n67 CSoutput.n3 165.8
R19965 CSoutput.n66 CSoutput.n65 165.8
R19966 CSoutput.n63 CSoutput.n4 165.8
R19967 CSoutput.n61 CSoutput.n60 165.8
R19968 CSoutput.n59 CSoutput.n5 165.8
R19969 CSoutput.n58 CSoutput.n57 165.8
R19970 CSoutput.n55 CSoutput.n6 165.8
R19971 CSoutput.n54 CSoutput.n53 165.8
R19972 CSoutput.n52 CSoutput.n51 165.8
R19973 CSoutput.n50 CSoutput.n8 165.8
R19974 CSoutput.n48 CSoutput.n47 165.8
R19975 CSoutput.n46 CSoutput.n9 165.8
R19976 CSoutput.n45 CSoutput.n44 165.8
R19977 CSoutput.n42 CSoutput.n10 165.8
R19978 CSoutput.n41 CSoutput.n40 165.8
R19979 CSoutput.n39 CSoutput.n38 165.8
R19980 CSoutput.n37 CSoutput.n12 165.8
R19981 CSoutput.n35 CSoutput.n34 165.8
R19982 CSoutput.n33 CSoutput.n13 165.8
R19983 CSoutput.n32 CSoutput.n31 165.8
R19984 CSoutput.n29 CSoutput.n14 165.8
R19985 CSoutput.n28 CSoutput.n27 165.8
R19986 CSoutput.n26 CSoutput.n25 165.8
R19987 CSoutput.n24 CSoutput.n16 165.8
R19988 CSoutput.n22 CSoutput.n21 165.8
R19989 CSoutput.n20 CSoutput.n17 165.8
R19990 CSoutput.n77 CSoutput.t162 162.194
R19991 CSoutput.n18 CSoutput.t150 120.501
R19992 CSoutput.n23 CSoutput.t152 120.501
R19993 CSoutput.n15 CSoutput.t163 120.501
R19994 CSoutput.n30 CSoutput.t153 120.501
R19995 CSoutput.n36 CSoutput.t154 120.501
R19996 CSoutput.n11 CSoutput.t148 120.501
R19997 CSoutput.n43 CSoutput.t160 120.501
R19998 CSoutput.n49 CSoutput.t157 120.501
R19999 CSoutput.n7 CSoutput.t151 120.501
R20000 CSoutput.n56 CSoutput.t147 120.501
R20001 CSoutput.n62 CSoutput.t158 120.501
R20002 CSoutput.n64 CSoutput.t159 120.501
R20003 CSoutput.n70 CSoutput.t149 120.501
R20004 CSoutput.n1 CSoutput.t144 120.501
R20005 CSoutput.n290 CSoutput.n288 103.469
R20006 CSoutput.n278 CSoutput.n276 103.469
R20007 CSoutput.n267 CSoutput.n265 103.469
R20008 CSoutput.n104 CSoutput.n102 103.469
R20009 CSoutput.n92 CSoutput.n90 103.469
R20010 CSoutput.n81 CSoutput.n79 103.469
R20011 CSoutput.n296 CSoutput.n295 103.111
R20012 CSoutput.n294 CSoutput.n293 103.111
R20013 CSoutput.n292 CSoutput.n291 103.111
R20014 CSoutput.n290 CSoutput.n289 103.111
R20015 CSoutput.n286 CSoutput.n285 103.111
R20016 CSoutput.n284 CSoutput.n283 103.111
R20017 CSoutput.n282 CSoutput.n281 103.111
R20018 CSoutput.n280 CSoutput.n279 103.111
R20019 CSoutput.n278 CSoutput.n277 103.111
R20020 CSoutput.n275 CSoutput.n274 103.111
R20021 CSoutput.n273 CSoutput.n272 103.111
R20022 CSoutput.n271 CSoutput.n270 103.111
R20023 CSoutput.n269 CSoutput.n268 103.111
R20024 CSoutput.n267 CSoutput.n266 103.111
R20025 CSoutput.n104 CSoutput.n103 103.111
R20026 CSoutput.n106 CSoutput.n105 103.111
R20027 CSoutput.n108 CSoutput.n107 103.111
R20028 CSoutput.n110 CSoutput.n109 103.111
R20029 CSoutput.n112 CSoutput.n111 103.111
R20030 CSoutput.n92 CSoutput.n91 103.111
R20031 CSoutput.n94 CSoutput.n93 103.111
R20032 CSoutput.n96 CSoutput.n95 103.111
R20033 CSoutput.n98 CSoutput.n97 103.111
R20034 CSoutput.n100 CSoutput.n99 103.111
R20035 CSoutput.n81 CSoutput.n80 103.111
R20036 CSoutput.n83 CSoutput.n82 103.111
R20037 CSoutput.n85 CSoutput.n84 103.111
R20038 CSoutput.n87 CSoutput.n86 103.111
R20039 CSoutput.n89 CSoutput.n88 103.111
R20040 CSoutput.n298 CSoutput.n297 103.111
R20041 CSoutput.n326 CSoutput.n324 81.5057
R20042 CSoutput.n314 CSoutput.n312 81.5057
R20043 CSoutput.n303 CSoutput.n301 81.5057
R20044 CSoutput.n362 CSoutput.n360 81.5057
R20045 CSoutput.n350 CSoutput.n348 81.5057
R20046 CSoutput.n339 CSoutput.n337 81.5057
R20047 CSoutput.n334 CSoutput.n333 80.9324
R20048 CSoutput.n332 CSoutput.n331 80.9324
R20049 CSoutput.n330 CSoutput.n329 80.9324
R20050 CSoutput.n328 CSoutput.n327 80.9324
R20051 CSoutput.n326 CSoutput.n325 80.9324
R20052 CSoutput.n322 CSoutput.n321 80.9324
R20053 CSoutput.n320 CSoutput.n319 80.9324
R20054 CSoutput.n318 CSoutput.n317 80.9324
R20055 CSoutput.n316 CSoutput.n315 80.9324
R20056 CSoutput.n314 CSoutput.n313 80.9324
R20057 CSoutput.n311 CSoutput.n310 80.9324
R20058 CSoutput.n309 CSoutput.n308 80.9324
R20059 CSoutput.n307 CSoutput.n306 80.9324
R20060 CSoutput.n305 CSoutput.n304 80.9324
R20061 CSoutput.n303 CSoutput.n302 80.9324
R20062 CSoutput.n362 CSoutput.n361 80.9324
R20063 CSoutput.n364 CSoutput.n363 80.9324
R20064 CSoutput.n366 CSoutput.n365 80.9324
R20065 CSoutput.n368 CSoutput.n367 80.9324
R20066 CSoutput.n370 CSoutput.n369 80.9324
R20067 CSoutput.n350 CSoutput.n349 80.9324
R20068 CSoutput.n352 CSoutput.n351 80.9324
R20069 CSoutput.n354 CSoutput.n353 80.9324
R20070 CSoutput.n356 CSoutput.n355 80.9324
R20071 CSoutput.n358 CSoutput.n357 80.9324
R20072 CSoutput.n339 CSoutput.n338 80.9324
R20073 CSoutput.n341 CSoutput.n340 80.9324
R20074 CSoutput.n343 CSoutput.n342 80.9324
R20075 CSoutput.n345 CSoutput.n344 80.9324
R20076 CSoutput.n347 CSoutput.n346 80.9324
R20077 CSoutput.n25 CSoutput.n24 48.1486
R20078 CSoutput.n69 CSoutput.n3 48.1486
R20079 CSoutput.n38 CSoutput.n37 48.1486
R20080 CSoutput.n42 CSoutput.n41 48.1486
R20081 CSoutput.n51 CSoutput.n50 48.1486
R20082 CSoutput.n55 CSoutput.n54 48.1486
R20083 CSoutput.n22 CSoutput.n17 46.462
R20084 CSoutput.n72 CSoutput.n71 46.462
R20085 CSoutput.n20 CSoutput.n19 44.9055
R20086 CSoutput.n29 CSoutput.n28 43.7635
R20087 CSoutput.n65 CSoutput.n63 43.7635
R20088 CSoutput.n35 CSoutput.n13 41.7396
R20089 CSoutput.n57 CSoutput.n5 41.7396
R20090 CSoutput.n44 CSoutput.n9 37.0171
R20091 CSoutput.n48 CSoutput.n9 37.0171
R20092 CSoutput.n76 CSoutput.n75 34.9932
R20093 CSoutput.n31 CSoutput.n13 32.2947
R20094 CSoutput.n61 CSoutput.n5 32.2947
R20095 CSoutput.n30 CSoutput.n29 29.6014
R20096 CSoutput.n63 CSoutput.n62 29.6014
R20097 CSoutput.n19 CSoutput.n18 28.4085
R20098 CSoutput.n18 CSoutput.n17 25.1176
R20099 CSoutput.n72 CSoutput.n1 25.1176
R20100 CSoutput.n43 CSoutput.n42 22.0922
R20101 CSoutput.n50 CSoutput.n49 22.0922
R20102 CSoutput.n77 CSoutput.n76 21.8586
R20103 CSoutput.n37 CSoutput.n36 18.9681
R20104 CSoutput.n56 CSoutput.n55 18.9681
R20105 CSoutput.n25 CSoutput.n15 17.6292
R20106 CSoutput.n64 CSoutput.n3 17.6292
R20107 CSoutput.n24 CSoutput.n23 15.844
R20108 CSoutput.n70 CSoutput.n69 15.844
R20109 CSoutput.n38 CSoutput.n11 14.5051
R20110 CSoutput.n54 CSoutput.n7 14.5051
R20111 CSoutput.n373 CSoutput.n78 11.4982
R20112 CSoutput.n41 CSoutput.n11 11.3811
R20113 CSoutput.n51 CSoutput.n7 11.3811
R20114 CSoutput.n23 CSoutput.n22 10.0422
R20115 CSoutput.n71 CSoutput.n70 10.0422
R20116 CSoutput.n287 CSoutput.n275 9.25285
R20117 CSoutput.n101 CSoutput.n89 9.25285
R20118 CSoutput.n323 CSoutput.n311 8.98182
R20119 CSoutput.n359 CSoutput.n347 8.98182
R20120 CSoutput.n336 CSoutput.n300 8.96934
R20121 CSoutput.n28 CSoutput.n15 8.25698
R20122 CSoutput.n65 CSoutput.n64 8.25698
R20123 CSoutput.n300 CSoutput.n299 7.12641
R20124 CSoutput.n114 CSoutput.n113 7.12641
R20125 CSoutput.n36 CSoutput.n35 6.91809
R20126 CSoutput.n57 CSoutput.n56 6.91809
R20127 CSoutput.n336 CSoutput.n335 6.02792
R20128 CSoutput.n372 CSoutput.n371 6.02792
R20129 CSoutput.n373 CSoutput.n114 5.3769
R20130 CSoutput.n335 CSoutput.n334 5.25266
R20131 CSoutput.n323 CSoutput.n322 5.25266
R20132 CSoutput.n371 CSoutput.n370 5.25266
R20133 CSoutput.n359 CSoutput.n358 5.25266
R20134 CSoutput.n299 CSoutput.n298 5.1449
R20135 CSoutput.n287 CSoutput.n286 5.1449
R20136 CSoutput.n113 CSoutput.n112 5.1449
R20137 CSoutput.n101 CSoutput.n100 5.1449
R20138 CSoutput.n205 CSoutput.n158 4.5005
R20139 CSoutput.n174 CSoutput.n158 4.5005
R20140 CSoutput.n169 CSoutput.n153 4.5005
R20141 CSoutput.n169 CSoutput.n155 4.5005
R20142 CSoutput.n169 CSoutput.n152 4.5005
R20143 CSoutput.n169 CSoutput.n156 4.5005
R20144 CSoutput.n169 CSoutput.n151 4.5005
R20145 CSoutput.n169 CSoutput.t164 4.5005
R20146 CSoutput.n169 CSoutput.n150 4.5005
R20147 CSoutput.n169 CSoutput.n157 4.5005
R20148 CSoutput.n169 CSoutput.n158 4.5005
R20149 CSoutput.n167 CSoutput.n153 4.5005
R20150 CSoutput.n167 CSoutput.n155 4.5005
R20151 CSoutput.n167 CSoutput.n152 4.5005
R20152 CSoutput.n167 CSoutput.n156 4.5005
R20153 CSoutput.n167 CSoutput.n151 4.5005
R20154 CSoutput.n167 CSoutput.t164 4.5005
R20155 CSoutput.n167 CSoutput.n150 4.5005
R20156 CSoutput.n167 CSoutput.n157 4.5005
R20157 CSoutput.n167 CSoutput.n158 4.5005
R20158 CSoutput.n166 CSoutput.n153 4.5005
R20159 CSoutput.n166 CSoutput.n155 4.5005
R20160 CSoutput.n166 CSoutput.n152 4.5005
R20161 CSoutput.n166 CSoutput.n156 4.5005
R20162 CSoutput.n166 CSoutput.n151 4.5005
R20163 CSoutput.n166 CSoutput.t164 4.5005
R20164 CSoutput.n166 CSoutput.n150 4.5005
R20165 CSoutput.n166 CSoutput.n157 4.5005
R20166 CSoutput.n166 CSoutput.n158 4.5005
R20167 CSoutput.n251 CSoutput.n153 4.5005
R20168 CSoutput.n251 CSoutput.n155 4.5005
R20169 CSoutput.n251 CSoutput.n152 4.5005
R20170 CSoutput.n251 CSoutput.n156 4.5005
R20171 CSoutput.n251 CSoutput.n151 4.5005
R20172 CSoutput.n251 CSoutput.t164 4.5005
R20173 CSoutput.n251 CSoutput.n150 4.5005
R20174 CSoutput.n251 CSoutput.n157 4.5005
R20175 CSoutput.n251 CSoutput.n158 4.5005
R20176 CSoutput.n249 CSoutput.n153 4.5005
R20177 CSoutput.n249 CSoutput.n155 4.5005
R20178 CSoutput.n249 CSoutput.n152 4.5005
R20179 CSoutput.n249 CSoutput.n156 4.5005
R20180 CSoutput.n249 CSoutput.n151 4.5005
R20181 CSoutput.n249 CSoutput.t164 4.5005
R20182 CSoutput.n249 CSoutput.n150 4.5005
R20183 CSoutput.n249 CSoutput.n157 4.5005
R20184 CSoutput.n247 CSoutput.n153 4.5005
R20185 CSoutput.n247 CSoutput.n155 4.5005
R20186 CSoutput.n247 CSoutput.n152 4.5005
R20187 CSoutput.n247 CSoutput.n156 4.5005
R20188 CSoutput.n247 CSoutput.n151 4.5005
R20189 CSoutput.n247 CSoutput.t164 4.5005
R20190 CSoutput.n247 CSoutput.n150 4.5005
R20191 CSoutput.n247 CSoutput.n157 4.5005
R20192 CSoutput.n177 CSoutput.n153 4.5005
R20193 CSoutput.n177 CSoutput.n155 4.5005
R20194 CSoutput.n177 CSoutput.n152 4.5005
R20195 CSoutput.n177 CSoutput.n156 4.5005
R20196 CSoutput.n177 CSoutput.n151 4.5005
R20197 CSoutput.n177 CSoutput.t164 4.5005
R20198 CSoutput.n177 CSoutput.n150 4.5005
R20199 CSoutput.n177 CSoutput.n157 4.5005
R20200 CSoutput.n177 CSoutput.n158 4.5005
R20201 CSoutput.n176 CSoutput.n153 4.5005
R20202 CSoutput.n176 CSoutput.n155 4.5005
R20203 CSoutput.n176 CSoutput.n152 4.5005
R20204 CSoutput.n176 CSoutput.n156 4.5005
R20205 CSoutput.n176 CSoutput.n151 4.5005
R20206 CSoutput.n176 CSoutput.t164 4.5005
R20207 CSoutput.n176 CSoutput.n150 4.5005
R20208 CSoutput.n176 CSoutput.n157 4.5005
R20209 CSoutput.n176 CSoutput.n158 4.5005
R20210 CSoutput.n180 CSoutput.n153 4.5005
R20211 CSoutput.n180 CSoutput.n155 4.5005
R20212 CSoutput.n180 CSoutput.n152 4.5005
R20213 CSoutput.n180 CSoutput.n156 4.5005
R20214 CSoutput.n180 CSoutput.n151 4.5005
R20215 CSoutput.n180 CSoutput.t164 4.5005
R20216 CSoutput.n180 CSoutput.n150 4.5005
R20217 CSoutput.n180 CSoutput.n157 4.5005
R20218 CSoutput.n180 CSoutput.n158 4.5005
R20219 CSoutput.n179 CSoutput.n153 4.5005
R20220 CSoutput.n179 CSoutput.n155 4.5005
R20221 CSoutput.n179 CSoutput.n152 4.5005
R20222 CSoutput.n179 CSoutput.n156 4.5005
R20223 CSoutput.n179 CSoutput.n151 4.5005
R20224 CSoutput.n179 CSoutput.t164 4.5005
R20225 CSoutput.n179 CSoutput.n150 4.5005
R20226 CSoutput.n179 CSoutput.n157 4.5005
R20227 CSoutput.n179 CSoutput.n158 4.5005
R20228 CSoutput.n162 CSoutput.n153 4.5005
R20229 CSoutput.n162 CSoutput.n155 4.5005
R20230 CSoutput.n162 CSoutput.n152 4.5005
R20231 CSoutput.n162 CSoutput.n156 4.5005
R20232 CSoutput.n162 CSoutput.n151 4.5005
R20233 CSoutput.n162 CSoutput.t164 4.5005
R20234 CSoutput.n162 CSoutput.n150 4.5005
R20235 CSoutput.n162 CSoutput.n157 4.5005
R20236 CSoutput.n162 CSoutput.n158 4.5005
R20237 CSoutput.n254 CSoutput.n153 4.5005
R20238 CSoutput.n254 CSoutput.n155 4.5005
R20239 CSoutput.n254 CSoutput.n152 4.5005
R20240 CSoutput.n254 CSoutput.n156 4.5005
R20241 CSoutput.n254 CSoutput.n151 4.5005
R20242 CSoutput.n254 CSoutput.t164 4.5005
R20243 CSoutput.n254 CSoutput.n150 4.5005
R20244 CSoutput.n254 CSoutput.n157 4.5005
R20245 CSoutput.n254 CSoutput.n158 4.5005
R20246 CSoutput.n241 CSoutput.n212 4.5005
R20247 CSoutput.n241 CSoutput.n218 4.5005
R20248 CSoutput.n199 CSoutput.n188 4.5005
R20249 CSoutput.n199 CSoutput.n190 4.5005
R20250 CSoutput.n199 CSoutput.n187 4.5005
R20251 CSoutput.n199 CSoutput.n191 4.5005
R20252 CSoutput.n199 CSoutput.n186 4.5005
R20253 CSoutput.n199 CSoutput.t156 4.5005
R20254 CSoutput.n199 CSoutput.n185 4.5005
R20255 CSoutput.n199 CSoutput.n192 4.5005
R20256 CSoutput.n241 CSoutput.n199 4.5005
R20257 CSoutput.n220 CSoutput.n188 4.5005
R20258 CSoutput.n220 CSoutput.n190 4.5005
R20259 CSoutput.n220 CSoutput.n187 4.5005
R20260 CSoutput.n220 CSoutput.n191 4.5005
R20261 CSoutput.n220 CSoutput.n186 4.5005
R20262 CSoutput.n220 CSoutput.t156 4.5005
R20263 CSoutput.n220 CSoutput.n185 4.5005
R20264 CSoutput.n220 CSoutput.n192 4.5005
R20265 CSoutput.n241 CSoutput.n220 4.5005
R20266 CSoutput.n198 CSoutput.n188 4.5005
R20267 CSoutput.n198 CSoutput.n190 4.5005
R20268 CSoutput.n198 CSoutput.n187 4.5005
R20269 CSoutput.n198 CSoutput.n191 4.5005
R20270 CSoutput.n198 CSoutput.n186 4.5005
R20271 CSoutput.n198 CSoutput.t156 4.5005
R20272 CSoutput.n198 CSoutput.n185 4.5005
R20273 CSoutput.n198 CSoutput.n192 4.5005
R20274 CSoutput.n241 CSoutput.n198 4.5005
R20275 CSoutput.n222 CSoutput.n188 4.5005
R20276 CSoutput.n222 CSoutput.n190 4.5005
R20277 CSoutput.n222 CSoutput.n187 4.5005
R20278 CSoutput.n222 CSoutput.n191 4.5005
R20279 CSoutput.n222 CSoutput.n186 4.5005
R20280 CSoutput.n222 CSoutput.t156 4.5005
R20281 CSoutput.n222 CSoutput.n185 4.5005
R20282 CSoutput.n222 CSoutput.n192 4.5005
R20283 CSoutput.n241 CSoutput.n222 4.5005
R20284 CSoutput.n188 CSoutput.n183 4.5005
R20285 CSoutput.n190 CSoutput.n183 4.5005
R20286 CSoutput.n187 CSoutput.n183 4.5005
R20287 CSoutput.n191 CSoutput.n183 4.5005
R20288 CSoutput.n186 CSoutput.n183 4.5005
R20289 CSoutput.t156 CSoutput.n183 4.5005
R20290 CSoutput.n185 CSoutput.n183 4.5005
R20291 CSoutput.n192 CSoutput.n183 4.5005
R20292 CSoutput.n244 CSoutput.n188 4.5005
R20293 CSoutput.n244 CSoutput.n190 4.5005
R20294 CSoutput.n244 CSoutput.n187 4.5005
R20295 CSoutput.n244 CSoutput.n191 4.5005
R20296 CSoutput.n244 CSoutput.n186 4.5005
R20297 CSoutput.n244 CSoutput.t156 4.5005
R20298 CSoutput.n244 CSoutput.n185 4.5005
R20299 CSoutput.n244 CSoutput.n192 4.5005
R20300 CSoutput.n242 CSoutput.n188 4.5005
R20301 CSoutput.n242 CSoutput.n190 4.5005
R20302 CSoutput.n242 CSoutput.n187 4.5005
R20303 CSoutput.n242 CSoutput.n191 4.5005
R20304 CSoutput.n242 CSoutput.n186 4.5005
R20305 CSoutput.n242 CSoutput.t156 4.5005
R20306 CSoutput.n242 CSoutput.n185 4.5005
R20307 CSoutput.n242 CSoutput.n192 4.5005
R20308 CSoutput.n242 CSoutput.n241 4.5005
R20309 CSoutput.n224 CSoutput.n188 4.5005
R20310 CSoutput.n224 CSoutput.n190 4.5005
R20311 CSoutput.n224 CSoutput.n187 4.5005
R20312 CSoutput.n224 CSoutput.n191 4.5005
R20313 CSoutput.n224 CSoutput.n186 4.5005
R20314 CSoutput.n224 CSoutput.t156 4.5005
R20315 CSoutput.n224 CSoutput.n185 4.5005
R20316 CSoutput.n224 CSoutput.n192 4.5005
R20317 CSoutput.n241 CSoutput.n224 4.5005
R20318 CSoutput.n196 CSoutput.n188 4.5005
R20319 CSoutput.n196 CSoutput.n190 4.5005
R20320 CSoutput.n196 CSoutput.n187 4.5005
R20321 CSoutput.n196 CSoutput.n191 4.5005
R20322 CSoutput.n196 CSoutput.n186 4.5005
R20323 CSoutput.n196 CSoutput.t156 4.5005
R20324 CSoutput.n196 CSoutput.n185 4.5005
R20325 CSoutput.n196 CSoutput.n192 4.5005
R20326 CSoutput.n241 CSoutput.n196 4.5005
R20327 CSoutput.n226 CSoutput.n188 4.5005
R20328 CSoutput.n226 CSoutput.n190 4.5005
R20329 CSoutput.n226 CSoutput.n187 4.5005
R20330 CSoutput.n226 CSoutput.n191 4.5005
R20331 CSoutput.n226 CSoutput.n186 4.5005
R20332 CSoutput.n226 CSoutput.t156 4.5005
R20333 CSoutput.n226 CSoutput.n185 4.5005
R20334 CSoutput.n226 CSoutput.n192 4.5005
R20335 CSoutput.n241 CSoutput.n226 4.5005
R20336 CSoutput.n195 CSoutput.n188 4.5005
R20337 CSoutput.n195 CSoutput.n190 4.5005
R20338 CSoutput.n195 CSoutput.n187 4.5005
R20339 CSoutput.n195 CSoutput.n191 4.5005
R20340 CSoutput.n195 CSoutput.n186 4.5005
R20341 CSoutput.n195 CSoutput.t156 4.5005
R20342 CSoutput.n195 CSoutput.n185 4.5005
R20343 CSoutput.n195 CSoutput.n192 4.5005
R20344 CSoutput.n241 CSoutput.n195 4.5005
R20345 CSoutput.n240 CSoutput.n188 4.5005
R20346 CSoutput.n240 CSoutput.n190 4.5005
R20347 CSoutput.n240 CSoutput.n187 4.5005
R20348 CSoutput.n240 CSoutput.n191 4.5005
R20349 CSoutput.n240 CSoutput.n186 4.5005
R20350 CSoutput.n240 CSoutput.t156 4.5005
R20351 CSoutput.n240 CSoutput.n185 4.5005
R20352 CSoutput.n240 CSoutput.n192 4.5005
R20353 CSoutput.n241 CSoutput.n240 4.5005
R20354 CSoutput.n239 CSoutput.n124 4.5005
R20355 CSoutput.n140 CSoutput.n124 4.5005
R20356 CSoutput.n135 CSoutput.n119 4.5005
R20357 CSoutput.n135 CSoutput.n121 4.5005
R20358 CSoutput.n135 CSoutput.n118 4.5005
R20359 CSoutput.n135 CSoutput.n122 4.5005
R20360 CSoutput.n135 CSoutput.n117 4.5005
R20361 CSoutput.n135 CSoutput.t155 4.5005
R20362 CSoutput.n135 CSoutput.n116 4.5005
R20363 CSoutput.n135 CSoutput.n123 4.5005
R20364 CSoutput.n135 CSoutput.n124 4.5005
R20365 CSoutput.n133 CSoutput.n119 4.5005
R20366 CSoutput.n133 CSoutput.n121 4.5005
R20367 CSoutput.n133 CSoutput.n118 4.5005
R20368 CSoutput.n133 CSoutput.n122 4.5005
R20369 CSoutput.n133 CSoutput.n117 4.5005
R20370 CSoutput.n133 CSoutput.t155 4.5005
R20371 CSoutput.n133 CSoutput.n116 4.5005
R20372 CSoutput.n133 CSoutput.n123 4.5005
R20373 CSoutput.n133 CSoutput.n124 4.5005
R20374 CSoutput.n132 CSoutput.n119 4.5005
R20375 CSoutput.n132 CSoutput.n121 4.5005
R20376 CSoutput.n132 CSoutput.n118 4.5005
R20377 CSoutput.n132 CSoutput.n122 4.5005
R20378 CSoutput.n132 CSoutput.n117 4.5005
R20379 CSoutput.n132 CSoutput.t155 4.5005
R20380 CSoutput.n132 CSoutput.n116 4.5005
R20381 CSoutput.n132 CSoutput.n123 4.5005
R20382 CSoutput.n132 CSoutput.n124 4.5005
R20383 CSoutput.n261 CSoutput.n119 4.5005
R20384 CSoutput.n261 CSoutput.n121 4.5005
R20385 CSoutput.n261 CSoutput.n118 4.5005
R20386 CSoutput.n261 CSoutput.n122 4.5005
R20387 CSoutput.n261 CSoutput.n117 4.5005
R20388 CSoutput.n261 CSoutput.t155 4.5005
R20389 CSoutput.n261 CSoutput.n116 4.5005
R20390 CSoutput.n261 CSoutput.n123 4.5005
R20391 CSoutput.n261 CSoutput.n124 4.5005
R20392 CSoutput.n259 CSoutput.n119 4.5005
R20393 CSoutput.n259 CSoutput.n121 4.5005
R20394 CSoutput.n259 CSoutput.n118 4.5005
R20395 CSoutput.n259 CSoutput.n122 4.5005
R20396 CSoutput.n259 CSoutput.n117 4.5005
R20397 CSoutput.n259 CSoutput.t155 4.5005
R20398 CSoutput.n259 CSoutput.n116 4.5005
R20399 CSoutput.n259 CSoutput.n123 4.5005
R20400 CSoutput.n257 CSoutput.n119 4.5005
R20401 CSoutput.n257 CSoutput.n121 4.5005
R20402 CSoutput.n257 CSoutput.n118 4.5005
R20403 CSoutput.n257 CSoutput.n122 4.5005
R20404 CSoutput.n257 CSoutput.n117 4.5005
R20405 CSoutput.n257 CSoutput.t155 4.5005
R20406 CSoutput.n257 CSoutput.n116 4.5005
R20407 CSoutput.n257 CSoutput.n123 4.5005
R20408 CSoutput.n143 CSoutput.n119 4.5005
R20409 CSoutput.n143 CSoutput.n121 4.5005
R20410 CSoutput.n143 CSoutput.n118 4.5005
R20411 CSoutput.n143 CSoutput.n122 4.5005
R20412 CSoutput.n143 CSoutput.n117 4.5005
R20413 CSoutput.n143 CSoutput.t155 4.5005
R20414 CSoutput.n143 CSoutput.n116 4.5005
R20415 CSoutput.n143 CSoutput.n123 4.5005
R20416 CSoutput.n143 CSoutput.n124 4.5005
R20417 CSoutput.n142 CSoutput.n119 4.5005
R20418 CSoutput.n142 CSoutput.n121 4.5005
R20419 CSoutput.n142 CSoutput.n118 4.5005
R20420 CSoutput.n142 CSoutput.n122 4.5005
R20421 CSoutput.n142 CSoutput.n117 4.5005
R20422 CSoutput.n142 CSoutput.t155 4.5005
R20423 CSoutput.n142 CSoutput.n116 4.5005
R20424 CSoutput.n142 CSoutput.n123 4.5005
R20425 CSoutput.n142 CSoutput.n124 4.5005
R20426 CSoutput.n146 CSoutput.n119 4.5005
R20427 CSoutput.n146 CSoutput.n121 4.5005
R20428 CSoutput.n146 CSoutput.n118 4.5005
R20429 CSoutput.n146 CSoutput.n122 4.5005
R20430 CSoutput.n146 CSoutput.n117 4.5005
R20431 CSoutput.n146 CSoutput.t155 4.5005
R20432 CSoutput.n146 CSoutput.n116 4.5005
R20433 CSoutput.n146 CSoutput.n123 4.5005
R20434 CSoutput.n146 CSoutput.n124 4.5005
R20435 CSoutput.n145 CSoutput.n119 4.5005
R20436 CSoutput.n145 CSoutput.n121 4.5005
R20437 CSoutput.n145 CSoutput.n118 4.5005
R20438 CSoutput.n145 CSoutput.n122 4.5005
R20439 CSoutput.n145 CSoutput.n117 4.5005
R20440 CSoutput.n145 CSoutput.t155 4.5005
R20441 CSoutput.n145 CSoutput.n116 4.5005
R20442 CSoutput.n145 CSoutput.n123 4.5005
R20443 CSoutput.n145 CSoutput.n124 4.5005
R20444 CSoutput.n128 CSoutput.n119 4.5005
R20445 CSoutput.n128 CSoutput.n121 4.5005
R20446 CSoutput.n128 CSoutput.n118 4.5005
R20447 CSoutput.n128 CSoutput.n122 4.5005
R20448 CSoutput.n128 CSoutput.n117 4.5005
R20449 CSoutput.n128 CSoutput.t155 4.5005
R20450 CSoutput.n128 CSoutput.n116 4.5005
R20451 CSoutput.n128 CSoutput.n123 4.5005
R20452 CSoutput.n128 CSoutput.n124 4.5005
R20453 CSoutput.n264 CSoutput.n119 4.5005
R20454 CSoutput.n264 CSoutput.n121 4.5005
R20455 CSoutput.n264 CSoutput.n118 4.5005
R20456 CSoutput.n264 CSoutput.n122 4.5005
R20457 CSoutput.n264 CSoutput.n117 4.5005
R20458 CSoutput.n264 CSoutput.t155 4.5005
R20459 CSoutput.n264 CSoutput.n116 4.5005
R20460 CSoutput.n264 CSoutput.n123 4.5005
R20461 CSoutput.n264 CSoutput.n124 4.5005
R20462 CSoutput.n299 CSoutput.n287 4.10845
R20463 CSoutput.n113 CSoutput.n101 4.10845
R20464 CSoutput.n297 CSoutput.t95 4.06363
R20465 CSoutput.n297 CSoutput.t96 4.06363
R20466 CSoutput.n295 CSoutput.t101 4.06363
R20467 CSoutput.n295 CSoutput.t140 4.06363
R20468 CSoutput.n293 CSoutput.t81 4.06363
R20469 CSoutput.n293 CSoutput.t99 4.06363
R20470 CSoutput.n291 CSoutput.t109 4.06363
R20471 CSoutput.n291 CSoutput.t124 4.06363
R20472 CSoutput.n289 CSoutput.t129 4.06363
R20473 CSoutput.n289 CSoutput.t83 4.06363
R20474 CSoutput.n288 CSoutput.t110 4.06363
R20475 CSoutput.n288 CSoutput.t111 4.06363
R20476 CSoutput.n285 CSoutput.t88 4.06363
R20477 CSoutput.n285 CSoutput.t89 4.06363
R20478 CSoutput.n283 CSoutput.t91 4.06363
R20479 CSoutput.n283 CSoutput.t133 4.06363
R20480 CSoutput.n281 CSoutput.t143 4.06363
R20481 CSoutput.n281 CSoutput.t90 4.06363
R20482 CSoutput.n279 CSoutput.t102 4.06363
R20483 CSoutput.n279 CSoutput.t116 4.06363
R20484 CSoutput.n277 CSoutput.t117 4.06363
R20485 CSoutput.n277 CSoutput.t75 4.06363
R20486 CSoutput.n276 CSoutput.t105 4.06363
R20487 CSoutput.n276 CSoutput.t106 4.06363
R20488 CSoutput.n274 CSoutput.t93 4.06363
R20489 CSoutput.n274 CSoutput.t79 4.06363
R20490 CSoutput.n272 CSoutput.t121 4.06363
R20491 CSoutput.n272 CSoutput.t77 4.06363
R20492 CSoutput.n270 CSoutput.t98 4.06363
R20493 CSoutput.n270 CSoutput.t139 4.06363
R20494 CSoutput.n268 CSoutput.t86 4.06363
R20495 CSoutput.n268 CSoutput.t125 4.06363
R20496 CSoutput.n266 CSoutput.t104 4.06363
R20497 CSoutput.n266 CSoutput.t141 4.06363
R20498 CSoutput.n265 CSoutput.t73 4.06363
R20499 CSoutput.n265 CSoutput.t131 4.06363
R20500 CSoutput.n102 CSoutput.t136 4.06363
R20501 CSoutput.n102 CSoutput.t137 4.06363
R20502 CSoutput.n103 CSoutput.t123 4.06363
R20503 CSoutput.n103 CSoutput.t84 4.06363
R20504 CSoutput.n105 CSoutput.t82 4.06363
R20505 CSoutput.n105 CSoutput.t135 4.06363
R20506 CSoutput.n107 CSoutput.t122 4.06363
R20507 CSoutput.n107 CSoutput.t107 4.06363
R20508 CSoutput.n109 CSoutput.t94 4.06363
R20509 CSoutput.n109 CSoutput.t142 4.06363
R20510 CSoutput.n111 CSoutput.t119 4.06363
R20511 CSoutput.n111 CSoutput.t118 4.06363
R20512 CSoutput.n90 CSoutput.t130 4.06363
R20513 CSoutput.n90 CSoutput.t128 4.06363
R20514 CSoutput.n91 CSoutput.t115 4.06363
R20515 CSoutput.n91 CSoutput.t78 4.06363
R20516 CSoutput.n93 CSoutput.t74 4.06363
R20517 CSoutput.n93 CSoutput.t126 4.06363
R20518 CSoutput.n95 CSoutput.t114 4.06363
R20519 CSoutput.n95 CSoutput.t100 4.06363
R20520 CSoutput.n97 CSoutput.t87 4.06363
R20521 CSoutput.n97 CSoutput.t134 4.06363
R20522 CSoutput.n99 CSoutput.t113 4.06363
R20523 CSoutput.n99 CSoutput.t112 4.06363
R20524 CSoutput.n79 CSoutput.t132 4.06363
R20525 CSoutput.n79 CSoutput.t72 4.06363
R20526 CSoutput.n80 CSoutput.t120 4.06363
R20527 CSoutput.n80 CSoutput.t103 4.06363
R20528 CSoutput.n82 CSoutput.t127 4.06363
R20529 CSoutput.n82 CSoutput.t85 4.06363
R20530 CSoutput.n84 CSoutput.t138 4.06363
R20531 CSoutput.n84 CSoutput.t97 4.06363
R20532 CSoutput.n86 CSoutput.t76 4.06363
R20533 CSoutput.n86 CSoutput.t108 4.06363
R20534 CSoutput.n88 CSoutput.t80 4.06363
R20535 CSoutput.n88 CSoutput.t92 4.06363
R20536 CSoutput.n44 CSoutput.n43 3.79402
R20537 CSoutput.n49 CSoutput.n48 3.79402
R20538 CSoutput.n335 CSoutput.n323 3.72967
R20539 CSoutput.n371 CSoutput.n359 3.72967
R20540 CSoutput.n373 CSoutput.n372 3.57343
R20541 CSoutput.n372 CSoutput.n336 3.04641
R20542 CSoutput.n333 CSoutput.t44 2.82907
R20543 CSoutput.n333 CSoutput.t2 2.82907
R20544 CSoutput.n331 CSoutput.t70 2.82907
R20545 CSoutput.n331 CSoutput.t60 2.82907
R20546 CSoutput.n329 CSoutput.t26 2.82907
R20547 CSoutput.n329 CSoutput.t35 2.82907
R20548 CSoutput.n327 CSoutput.t1 2.82907
R20549 CSoutput.n327 CSoutput.t67 2.82907
R20550 CSoutput.n325 CSoutput.t59 2.82907
R20551 CSoutput.n325 CSoutput.t15 2.82907
R20552 CSoutput.n324 CSoutput.t8 2.82907
R20553 CSoutput.n324 CSoutput.t69 2.82907
R20554 CSoutput.n321 CSoutput.t12 2.82907
R20555 CSoutput.n321 CSoutput.t22 2.82907
R20556 CSoutput.n319 CSoutput.t21 2.82907
R20557 CSoutput.n319 CSoutput.t7 2.82907
R20558 CSoutput.n317 CSoutput.t33 2.82907
R20559 CSoutput.n317 CSoutput.t11 2.82907
R20560 CSoutput.n315 CSoutput.t14 2.82907
R20561 CSoutput.n315 CSoutput.t20 2.82907
R20562 CSoutput.n313 CSoutput.t18 2.82907
R20563 CSoutput.n313 CSoutput.t31 2.82907
R20564 CSoutput.n312 CSoutput.t30 2.82907
R20565 CSoutput.n312 CSoutput.t13 2.82907
R20566 CSoutput.n310 CSoutput.t53 2.82907
R20567 CSoutput.n310 CSoutput.t24 2.82907
R20568 CSoutput.n308 CSoutput.t4 2.82907
R20569 CSoutput.n308 CSoutput.t40 2.82907
R20570 CSoutput.n306 CSoutput.t19 2.82907
R20571 CSoutput.n306 CSoutput.t32 2.82907
R20572 CSoutput.n304 CSoutput.t34 2.82907
R20573 CSoutput.n304 CSoutput.t65 2.82907
R20574 CSoutput.n302 CSoutput.t50 2.82907
R20575 CSoutput.n302 CSoutput.t0 2.82907
R20576 CSoutput.n301 CSoutput.t63 2.82907
R20577 CSoutput.n301 CSoutput.t10 2.82907
R20578 CSoutput.n360 CSoutput.t57 2.82907
R20579 CSoutput.n360 CSoutput.t68 2.82907
R20580 CSoutput.n361 CSoutput.t71 2.82907
R20581 CSoutput.n361 CSoutput.t48 2.82907
R20582 CSoutput.n363 CSoutput.t52 2.82907
R20583 CSoutput.n363 CSoutput.t62 2.82907
R20584 CSoutput.n365 CSoutput.t9 2.82907
R20585 CSoutput.n365 CSoutput.t42 2.82907
R20586 CSoutput.n367 CSoutput.t47 2.82907
R20587 CSoutput.n367 CSoutput.t58 2.82907
R20588 CSoutput.n369 CSoutput.t64 2.82907
R20589 CSoutput.n369 CSoutput.t51 2.82907
R20590 CSoutput.n348 CSoutput.t28 2.82907
R20591 CSoutput.n348 CSoutput.t45 2.82907
R20592 CSoutput.n349 CSoutput.t46 2.82907
R20593 CSoutput.n349 CSoutput.t36 2.82907
R20594 CSoutput.n351 CSoutput.t37 2.82907
R20595 CSoutput.n351 CSoutput.t29 2.82907
R20596 CSoutput.n353 CSoutput.t23 2.82907
R20597 CSoutput.n353 CSoutput.t16 2.82907
R20598 CSoutput.n355 CSoutput.t17 2.82907
R20599 CSoutput.n355 CSoutput.t38 2.82907
R20600 CSoutput.n357 CSoutput.t39 2.82907
R20601 CSoutput.n357 CSoutput.t3 2.82907
R20602 CSoutput.n337 CSoutput.t41 2.82907
R20603 CSoutput.n337 CSoutput.t5 2.82907
R20604 CSoutput.n338 CSoutput.t25 2.82907
R20605 CSoutput.n338 CSoutput.t66 2.82907
R20606 CSoutput.n340 CSoutput.t6 2.82907
R20607 CSoutput.n340 CSoutput.t55 2.82907
R20608 CSoutput.n342 CSoutput.t54 2.82907
R20609 CSoutput.n342 CSoutput.t43 2.82907
R20610 CSoutput.n344 CSoutput.t56 2.82907
R20611 CSoutput.n344 CSoutput.t27 2.82907
R20612 CSoutput.n346 CSoutput.t49 2.82907
R20613 CSoutput.n346 CSoutput.t61 2.82907
R20614 CSoutput.n75 CSoutput.n1 2.45513
R20615 CSoutput.n205 CSoutput.n203 2.251
R20616 CSoutput.n205 CSoutput.n202 2.251
R20617 CSoutput.n205 CSoutput.n201 2.251
R20618 CSoutput.n205 CSoutput.n200 2.251
R20619 CSoutput.n174 CSoutput.n173 2.251
R20620 CSoutput.n174 CSoutput.n172 2.251
R20621 CSoutput.n174 CSoutput.n171 2.251
R20622 CSoutput.n174 CSoutput.n170 2.251
R20623 CSoutput.n247 CSoutput.n246 2.251
R20624 CSoutput.n212 CSoutput.n210 2.251
R20625 CSoutput.n212 CSoutput.n209 2.251
R20626 CSoutput.n212 CSoutput.n208 2.251
R20627 CSoutput.n230 CSoutput.n212 2.251
R20628 CSoutput.n218 CSoutput.n217 2.251
R20629 CSoutput.n218 CSoutput.n216 2.251
R20630 CSoutput.n218 CSoutput.n215 2.251
R20631 CSoutput.n218 CSoutput.n214 2.251
R20632 CSoutput.n244 CSoutput.n184 2.251
R20633 CSoutput.n239 CSoutput.n237 2.251
R20634 CSoutput.n239 CSoutput.n236 2.251
R20635 CSoutput.n239 CSoutput.n235 2.251
R20636 CSoutput.n239 CSoutput.n234 2.251
R20637 CSoutput.n140 CSoutput.n139 2.251
R20638 CSoutput.n140 CSoutput.n138 2.251
R20639 CSoutput.n140 CSoutput.n137 2.251
R20640 CSoutput.n140 CSoutput.n136 2.251
R20641 CSoutput.n257 CSoutput.n256 2.251
R20642 CSoutput.n174 CSoutput.n154 2.2505
R20643 CSoutput.n169 CSoutput.n154 2.2505
R20644 CSoutput.n167 CSoutput.n154 2.2505
R20645 CSoutput.n166 CSoutput.n154 2.2505
R20646 CSoutput.n251 CSoutput.n154 2.2505
R20647 CSoutput.n249 CSoutput.n154 2.2505
R20648 CSoutput.n247 CSoutput.n154 2.2505
R20649 CSoutput.n177 CSoutput.n154 2.2505
R20650 CSoutput.n176 CSoutput.n154 2.2505
R20651 CSoutput.n180 CSoutput.n154 2.2505
R20652 CSoutput.n179 CSoutput.n154 2.2505
R20653 CSoutput.n162 CSoutput.n154 2.2505
R20654 CSoutput.n254 CSoutput.n154 2.2505
R20655 CSoutput.n254 CSoutput.n253 2.2505
R20656 CSoutput.n218 CSoutput.n189 2.2505
R20657 CSoutput.n199 CSoutput.n189 2.2505
R20658 CSoutput.n220 CSoutput.n189 2.2505
R20659 CSoutput.n198 CSoutput.n189 2.2505
R20660 CSoutput.n222 CSoutput.n189 2.2505
R20661 CSoutput.n189 CSoutput.n183 2.2505
R20662 CSoutput.n244 CSoutput.n189 2.2505
R20663 CSoutput.n242 CSoutput.n189 2.2505
R20664 CSoutput.n224 CSoutput.n189 2.2505
R20665 CSoutput.n196 CSoutput.n189 2.2505
R20666 CSoutput.n226 CSoutput.n189 2.2505
R20667 CSoutput.n195 CSoutput.n189 2.2505
R20668 CSoutput.n240 CSoutput.n189 2.2505
R20669 CSoutput.n240 CSoutput.n193 2.2505
R20670 CSoutput.n140 CSoutput.n120 2.2505
R20671 CSoutput.n135 CSoutput.n120 2.2505
R20672 CSoutput.n133 CSoutput.n120 2.2505
R20673 CSoutput.n132 CSoutput.n120 2.2505
R20674 CSoutput.n261 CSoutput.n120 2.2505
R20675 CSoutput.n259 CSoutput.n120 2.2505
R20676 CSoutput.n257 CSoutput.n120 2.2505
R20677 CSoutput.n143 CSoutput.n120 2.2505
R20678 CSoutput.n142 CSoutput.n120 2.2505
R20679 CSoutput.n146 CSoutput.n120 2.2505
R20680 CSoutput.n145 CSoutput.n120 2.2505
R20681 CSoutput.n128 CSoutput.n120 2.2505
R20682 CSoutput.n264 CSoutput.n120 2.2505
R20683 CSoutput.n264 CSoutput.n263 2.2505
R20684 CSoutput.n182 CSoutput.n175 2.25024
R20685 CSoutput.n182 CSoutput.n168 2.25024
R20686 CSoutput.n250 CSoutput.n182 2.25024
R20687 CSoutput.n182 CSoutput.n178 2.25024
R20688 CSoutput.n182 CSoutput.n181 2.25024
R20689 CSoutput.n182 CSoutput.n149 2.25024
R20690 CSoutput.n232 CSoutput.n229 2.25024
R20691 CSoutput.n232 CSoutput.n228 2.25024
R20692 CSoutput.n232 CSoutput.n227 2.25024
R20693 CSoutput.n232 CSoutput.n194 2.25024
R20694 CSoutput.n232 CSoutput.n231 2.25024
R20695 CSoutput.n233 CSoutput.n232 2.25024
R20696 CSoutput.n148 CSoutput.n141 2.25024
R20697 CSoutput.n148 CSoutput.n134 2.25024
R20698 CSoutput.n260 CSoutput.n148 2.25024
R20699 CSoutput.n148 CSoutput.n144 2.25024
R20700 CSoutput.n148 CSoutput.n147 2.25024
R20701 CSoutput.n148 CSoutput.n115 2.25024
R20702 CSoutput.n300 CSoutput.n114 2.15937
R20703 CSoutput.n249 CSoutput.n159 1.50111
R20704 CSoutput.n197 CSoutput.n183 1.50111
R20705 CSoutput.n259 CSoutput.n125 1.50111
R20706 CSoutput.n205 CSoutput.n204 1.501
R20707 CSoutput.n212 CSoutput.n211 1.501
R20708 CSoutput.n239 CSoutput.n238 1.501
R20709 CSoutput.n253 CSoutput.n164 1.12536
R20710 CSoutput.n253 CSoutput.n165 1.12536
R20711 CSoutput.n253 CSoutput.n252 1.12536
R20712 CSoutput.n213 CSoutput.n193 1.12536
R20713 CSoutput.n219 CSoutput.n193 1.12536
R20714 CSoutput.n221 CSoutput.n193 1.12536
R20715 CSoutput.n263 CSoutput.n130 1.12536
R20716 CSoutput.n263 CSoutput.n131 1.12536
R20717 CSoutput.n263 CSoutput.n262 1.12536
R20718 CSoutput.n253 CSoutput.n160 1.12536
R20719 CSoutput.n253 CSoutput.n161 1.12536
R20720 CSoutput.n253 CSoutput.n163 1.12536
R20721 CSoutput.n243 CSoutput.n193 1.12536
R20722 CSoutput.n223 CSoutput.n193 1.12536
R20723 CSoutput.n225 CSoutput.n193 1.12536
R20724 CSoutput.n263 CSoutput.n126 1.12536
R20725 CSoutput.n263 CSoutput.n127 1.12536
R20726 CSoutput.n263 CSoutput.n129 1.12536
R20727 CSoutput.n31 CSoutput.n30 0.669944
R20728 CSoutput.n62 CSoutput.n61 0.669944
R20729 CSoutput.n328 CSoutput.n326 0.573776
R20730 CSoutput.n330 CSoutput.n328 0.573776
R20731 CSoutput.n332 CSoutput.n330 0.573776
R20732 CSoutput.n334 CSoutput.n332 0.573776
R20733 CSoutput.n316 CSoutput.n314 0.573776
R20734 CSoutput.n318 CSoutput.n316 0.573776
R20735 CSoutput.n320 CSoutput.n318 0.573776
R20736 CSoutput.n322 CSoutput.n320 0.573776
R20737 CSoutput.n305 CSoutput.n303 0.573776
R20738 CSoutput.n307 CSoutput.n305 0.573776
R20739 CSoutput.n309 CSoutput.n307 0.573776
R20740 CSoutput.n311 CSoutput.n309 0.573776
R20741 CSoutput.n370 CSoutput.n368 0.573776
R20742 CSoutput.n368 CSoutput.n366 0.573776
R20743 CSoutput.n366 CSoutput.n364 0.573776
R20744 CSoutput.n364 CSoutput.n362 0.573776
R20745 CSoutput.n358 CSoutput.n356 0.573776
R20746 CSoutput.n356 CSoutput.n354 0.573776
R20747 CSoutput.n354 CSoutput.n352 0.573776
R20748 CSoutput.n352 CSoutput.n350 0.573776
R20749 CSoutput.n347 CSoutput.n345 0.573776
R20750 CSoutput.n345 CSoutput.n343 0.573776
R20751 CSoutput.n343 CSoutput.n341 0.573776
R20752 CSoutput.n341 CSoutput.n339 0.573776
R20753 CSoutput.n373 CSoutput.n264 0.53442
R20754 CSoutput.n292 CSoutput.n290 0.358259
R20755 CSoutput.n294 CSoutput.n292 0.358259
R20756 CSoutput.n296 CSoutput.n294 0.358259
R20757 CSoutput.n298 CSoutput.n296 0.358259
R20758 CSoutput.n280 CSoutput.n278 0.358259
R20759 CSoutput.n282 CSoutput.n280 0.358259
R20760 CSoutput.n284 CSoutput.n282 0.358259
R20761 CSoutput.n286 CSoutput.n284 0.358259
R20762 CSoutput.n269 CSoutput.n267 0.358259
R20763 CSoutput.n271 CSoutput.n269 0.358259
R20764 CSoutput.n273 CSoutput.n271 0.358259
R20765 CSoutput.n275 CSoutput.n273 0.358259
R20766 CSoutput.n112 CSoutput.n110 0.358259
R20767 CSoutput.n110 CSoutput.n108 0.358259
R20768 CSoutput.n108 CSoutput.n106 0.358259
R20769 CSoutput.n106 CSoutput.n104 0.358259
R20770 CSoutput.n100 CSoutput.n98 0.358259
R20771 CSoutput.n98 CSoutput.n96 0.358259
R20772 CSoutput.n96 CSoutput.n94 0.358259
R20773 CSoutput.n94 CSoutput.n92 0.358259
R20774 CSoutput.n89 CSoutput.n87 0.358259
R20775 CSoutput.n87 CSoutput.n85 0.358259
R20776 CSoutput.n85 CSoutput.n83 0.358259
R20777 CSoutput.n83 CSoutput.n81 0.358259
R20778 CSoutput.n21 CSoutput.n20 0.169105
R20779 CSoutput.n21 CSoutput.n16 0.169105
R20780 CSoutput.n26 CSoutput.n16 0.169105
R20781 CSoutput.n27 CSoutput.n26 0.169105
R20782 CSoutput.n27 CSoutput.n14 0.169105
R20783 CSoutput.n32 CSoutput.n14 0.169105
R20784 CSoutput.n33 CSoutput.n32 0.169105
R20785 CSoutput.n34 CSoutput.n33 0.169105
R20786 CSoutput.n34 CSoutput.n12 0.169105
R20787 CSoutput.n39 CSoutput.n12 0.169105
R20788 CSoutput.n40 CSoutput.n39 0.169105
R20789 CSoutput.n40 CSoutput.n10 0.169105
R20790 CSoutput.n45 CSoutput.n10 0.169105
R20791 CSoutput.n46 CSoutput.n45 0.169105
R20792 CSoutput.n47 CSoutput.n46 0.169105
R20793 CSoutput.n47 CSoutput.n8 0.169105
R20794 CSoutput.n52 CSoutput.n8 0.169105
R20795 CSoutput.n53 CSoutput.n52 0.169105
R20796 CSoutput.n53 CSoutput.n6 0.169105
R20797 CSoutput.n58 CSoutput.n6 0.169105
R20798 CSoutput.n59 CSoutput.n58 0.169105
R20799 CSoutput.n60 CSoutput.n59 0.169105
R20800 CSoutput.n60 CSoutput.n4 0.169105
R20801 CSoutput.n66 CSoutput.n4 0.169105
R20802 CSoutput.n67 CSoutput.n66 0.169105
R20803 CSoutput.n68 CSoutput.n67 0.169105
R20804 CSoutput.n68 CSoutput.n2 0.169105
R20805 CSoutput.n73 CSoutput.n2 0.169105
R20806 CSoutput.n74 CSoutput.n73 0.169105
R20807 CSoutput.n74 CSoutput.n0 0.169105
R20808 CSoutput.n78 CSoutput.n0 0.169105
R20809 CSoutput.n207 CSoutput.n206 0.0910737
R20810 CSoutput.n258 CSoutput.n255 0.0723685
R20811 CSoutput.n212 CSoutput.n207 0.0522944
R20812 CSoutput.n255 CSoutput.n254 0.0499135
R20813 CSoutput.n206 CSoutput.n205 0.0499135
R20814 CSoutput.n240 CSoutput.n239 0.0464294
R20815 CSoutput.n248 CSoutput.n245 0.0391444
R20816 CSoutput.n207 CSoutput.t165 0.023435
R20817 CSoutput.n255 CSoutput.t145 0.02262
R20818 CSoutput.n206 CSoutput.t146 0.02262
R20819 CSoutput CSoutput.n373 0.0052
R20820 CSoutput.n177 CSoutput.n160 0.00365111
R20821 CSoutput.n180 CSoutput.n161 0.00365111
R20822 CSoutput.n163 CSoutput.n162 0.00365111
R20823 CSoutput.n205 CSoutput.n164 0.00365111
R20824 CSoutput.n169 CSoutput.n165 0.00365111
R20825 CSoutput.n252 CSoutput.n166 0.00365111
R20826 CSoutput.n243 CSoutput.n242 0.00365111
R20827 CSoutput.n223 CSoutput.n196 0.00365111
R20828 CSoutput.n225 CSoutput.n195 0.00365111
R20829 CSoutput.n213 CSoutput.n212 0.00365111
R20830 CSoutput.n219 CSoutput.n199 0.00365111
R20831 CSoutput.n221 CSoutput.n198 0.00365111
R20832 CSoutput.n143 CSoutput.n126 0.00365111
R20833 CSoutput.n146 CSoutput.n127 0.00365111
R20834 CSoutput.n129 CSoutput.n128 0.00365111
R20835 CSoutput.n239 CSoutput.n130 0.00365111
R20836 CSoutput.n135 CSoutput.n131 0.00365111
R20837 CSoutput.n262 CSoutput.n132 0.00365111
R20838 CSoutput.n174 CSoutput.n164 0.00340054
R20839 CSoutput.n167 CSoutput.n165 0.00340054
R20840 CSoutput.n252 CSoutput.n251 0.00340054
R20841 CSoutput.n247 CSoutput.n160 0.00340054
R20842 CSoutput.n176 CSoutput.n161 0.00340054
R20843 CSoutput.n179 CSoutput.n163 0.00340054
R20844 CSoutput.n218 CSoutput.n213 0.00340054
R20845 CSoutput.n220 CSoutput.n219 0.00340054
R20846 CSoutput.n222 CSoutput.n221 0.00340054
R20847 CSoutput.n244 CSoutput.n243 0.00340054
R20848 CSoutput.n224 CSoutput.n223 0.00340054
R20849 CSoutput.n226 CSoutput.n225 0.00340054
R20850 CSoutput.n140 CSoutput.n130 0.00340054
R20851 CSoutput.n133 CSoutput.n131 0.00340054
R20852 CSoutput.n262 CSoutput.n261 0.00340054
R20853 CSoutput.n257 CSoutput.n126 0.00340054
R20854 CSoutput.n142 CSoutput.n127 0.00340054
R20855 CSoutput.n145 CSoutput.n129 0.00340054
R20856 CSoutput.n175 CSoutput.n169 0.00252698
R20857 CSoutput.n168 CSoutput.n166 0.00252698
R20858 CSoutput.n250 CSoutput.n249 0.00252698
R20859 CSoutput.n178 CSoutput.n176 0.00252698
R20860 CSoutput.n181 CSoutput.n179 0.00252698
R20861 CSoutput.n254 CSoutput.n149 0.00252698
R20862 CSoutput.n175 CSoutput.n174 0.00252698
R20863 CSoutput.n168 CSoutput.n167 0.00252698
R20864 CSoutput.n251 CSoutput.n250 0.00252698
R20865 CSoutput.n178 CSoutput.n177 0.00252698
R20866 CSoutput.n181 CSoutput.n180 0.00252698
R20867 CSoutput.n162 CSoutput.n149 0.00252698
R20868 CSoutput.n229 CSoutput.n199 0.00252698
R20869 CSoutput.n228 CSoutput.n198 0.00252698
R20870 CSoutput.n227 CSoutput.n183 0.00252698
R20871 CSoutput.n224 CSoutput.n194 0.00252698
R20872 CSoutput.n231 CSoutput.n226 0.00252698
R20873 CSoutput.n240 CSoutput.n233 0.00252698
R20874 CSoutput.n229 CSoutput.n218 0.00252698
R20875 CSoutput.n228 CSoutput.n220 0.00252698
R20876 CSoutput.n227 CSoutput.n222 0.00252698
R20877 CSoutput.n242 CSoutput.n194 0.00252698
R20878 CSoutput.n231 CSoutput.n196 0.00252698
R20879 CSoutput.n233 CSoutput.n195 0.00252698
R20880 CSoutput.n141 CSoutput.n135 0.00252698
R20881 CSoutput.n134 CSoutput.n132 0.00252698
R20882 CSoutput.n260 CSoutput.n259 0.00252698
R20883 CSoutput.n144 CSoutput.n142 0.00252698
R20884 CSoutput.n147 CSoutput.n145 0.00252698
R20885 CSoutput.n264 CSoutput.n115 0.00252698
R20886 CSoutput.n141 CSoutput.n140 0.00252698
R20887 CSoutput.n134 CSoutput.n133 0.00252698
R20888 CSoutput.n261 CSoutput.n260 0.00252698
R20889 CSoutput.n144 CSoutput.n143 0.00252698
R20890 CSoutput.n147 CSoutput.n146 0.00252698
R20891 CSoutput.n128 CSoutput.n115 0.00252698
R20892 CSoutput.n249 CSoutput.n248 0.0020275
R20893 CSoutput.n248 CSoutput.n247 0.0020275
R20894 CSoutput.n245 CSoutput.n183 0.0020275
R20895 CSoutput.n245 CSoutput.n244 0.0020275
R20896 CSoutput.n259 CSoutput.n258 0.0020275
R20897 CSoutput.n258 CSoutput.n257 0.0020275
R20898 CSoutput.n159 CSoutput.n158 0.00166668
R20899 CSoutput.n241 CSoutput.n197 0.00166668
R20900 CSoutput.n125 CSoutput.n124 0.00166668
R20901 CSoutput.n263 CSoutput.n125 0.00133328
R20902 CSoutput.n197 CSoutput.n193 0.00133328
R20903 CSoutput.n253 CSoutput.n159 0.00133328
R20904 CSoutput.n256 CSoutput.n148 0.001
R20905 CSoutput.n234 CSoutput.n148 0.001
R20906 CSoutput.n136 CSoutput.n116 0.001
R20907 CSoutput.n235 CSoutput.n116 0.001
R20908 CSoutput.n137 CSoutput.n117 0.001
R20909 CSoutput.n236 CSoutput.n117 0.001
R20910 CSoutput.n138 CSoutput.n118 0.001
R20911 CSoutput.n237 CSoutput.n118 0.001
R20912 CSoutput.n139 CSoutput.n119 0.001
R20913 CSoutput.n238 CSoutput.n119 0.001
R20914 CSoutput.n232 CSoutput.n184 0.001
R20915 CSoutput.n232 CSoutput.n230 0.001
R20916 CSoutput.n214 CSoutput.n185 0.001
R20917 CSoutput.n208 CSoutput.n185 0.001
R20918 CSoutput.n215 CSoutput.n186 0.001
R20919 CSoutput.n209 CSoutput.n186 0.001
R20920 CSoutput.n216 CSoutput.n187 0.001
R20921 CSoutput.n210 CSoutput.n187 0.001
R20922 CSoutput.n217 CSoutput.n188 0.001
R20923 CSoutput.n211 CSoutput.n188 0.001
R20924 CSoutput.n246 CSoutput.n182 0.001
R20925 CSoutput.n200 CSoutput.n182 0.001
R20926 CSoutput.n170 CSoutput.n150 0.001
R20927 CSoutput.n201 CSoutput.n150 0.001
R20928 CSoutput.n171 CSoutput.n151 0.001
R20929 CSoutput.n202 CSoutput.n151 0.001
R20930 CSoutput.n172 CSoutput.n152 0.001
R20931 CSoutput.n203 CSoutput.n152 0.001
R20932 CSoutput.n173 CSoutput.n153 0.001
R20933 CSoutput.n204 CSoutput.n153 0.001
R20934 CSoutput.n204 CSoutput.n154 0.001
R20935 CSoutput.n203 CSoutput.n155 0.001
R20936 CSoutput.n202 CSoutput.n156 0.001
R20937 CSoutput.n201 CSoutput.t164 0.001
R20938 CSoutput.n200 CSoutput.n157 0.001
R20939 CSoutput.n173 CSoutput.n155 0.001
R20940 CSoutput.n172 CSoutput.n156 0.001
R20941 CSoutput.n171 CSoutput.t164 0.001
R20942 CSoutput.n170 CSoutput.n157 0.001
R20943 CSoutput.n246 CSoutput.n158 0.001
R20944 CSoutput.n211 CSoutput.n189 0.001
R20945 CSoutput.n210 CSoutput.n190 0.001
R20946 CSoutput.n209 CSoutput.n191 0.001
R20947 CSoutput.n208 CSoutput.t156 0.001
R20948 CSoutput.n230 CSoutput.n192 0.001
R20949 CSoutput.n217 CSoutput.n190 0.001
R20950 CSoutput.n216 CSoutput.n191 0.001
R20951 CSoutput.n215 CSoutput.t156 0.001
R20952 CSoutput.n214 CSoutput.n192 0.001
R20953 CSoutput.n241 CSoutput.n184 0.001
R20954 CSoutput.n238 CSoutput.n120 0.001
R20955 CSoutput.n237 CSoutput.n121 0.001
R20956 CSoutput.n236 CSoutput.n122 0.001
R20957 CSoutput.n235 CSoutput.t155 0.001
R20958 CSoutput.n234 CSoutput.n123 0.001
R20959 CSoutput.n139 CSoutput.n121 0.001
R20960 CSoutput.n138 CSoutput.n122 0.001
R20961 CSoutput.n137 CSoutput.t155 0.001
R20962 CSoutput.n136 CSoutput.n123 0.001
R20963 CSoutput.n256 CSoutput.n124 0.001
R20964 a_n2848_n452.n3 a_n2848_n452.t75 539.01
R20965 a_n2848_n452.n55 a_n2848_n452.t58 512.366
R20966 a_n2848_n452.n54 a_n2848_n452.t62 512.366
R20967 a_n2848_n452.n52 a_n2848_n452.t52 512.366
R20968 a_n2848_n452.n53 a_n2848_n452.t67 512.366
R20969 a_n2848_n452.n44 a_n2848_n452.t24 533.058
R20970 a_n2848_n452.n56 a_n2848_n452.t14 512.366
R20971 a_n2848_n452.n57 a_n2848_n452.t20 512.366
R20972 a_n2848_n452.n49 a_n2848_n452.t22 512.366
R20973 a_n2848_n452.n78 a_n2848_n452.t12 512.366
R20974 a_n2848_n452.n76 a_n2848_n452.t16 512.366
R20975 a_n2848_n452.n17 a_n2848_n452.t10 539.01
R20976 a_n2848_n452.n100 a_n2848_n452.t30 512.366
R20977 a_n2848_n452.n101 a_n2848_n452.t32 512.366
R20978 a_n2848_n452.n50 a_n2848_n452.t26 512.366
R20979 a_n2848_n452.n102 a_n2848_n452.t28 512.366
R20980 a_n2848_n452.n21 a_n2848_n452.t70 539.01
R20981 a_n2848_n452.n97 a_n2848_n452.t71 512.366
R20982 a_n2848_n452.n98 a_n2848_n452.t50 512.366
R20983 a_n2848_n452.n51 a_n2848_n452.t56 512.366
R20984 a_n2848_n452.n99 a_n2848_n452.t65 512.366
R20985 a_n2848_n452.n89 a_n2848_n452.t64 512.366
R20986 a_n2848_n452.n88 a_n2848_n452.t55 512.366
R20987 a_n2848_n452.n87 a_n2848_n452.t49 512.366
R20988 a_n2848_n452.n91 a_n2848_n452.t72 512.366
R20989 a_n2848_n452.n90 a_n2848_n452.t61 512.366
R20990 a_n2848_n452.n86 a_n2848_n452.t60 512.366
R20991 a_n2848_n452.n93 a_n2848_n452.t68 512.366
R20992 a_n2848_n452.n92 a_n2848_n452.t53 512.366
R20993 a_n2848_n452.n85 a_n2848_n452.t54 512.366
R20994 a_n2848_n452.n95 a_n2848_n452.t57 512.366
R20995 a_n2848_n452.n94 a_n2848_n452.t66 512.366
R20996 a_n2848_n452.n84 a_n2848_n452.t48 512.366
R20997 a_n2848_n452.n47 a_n2848_n452.n1 70.3058
R20998 a_n2848_n452.n48 a_n2848_n452.n5 70.1674
R20999 a_n2848_n452.n14 a_n2848_n452.n33 70.3058
R21000 a_n2848_n452.n18 a_n2848_n452.n30 70.3058
R21001 a_n2848_n452.n29 a_n2848_n452.n19 70.1674
R21002 a_n2848_n452.n29 a_n2848_n452.n51 20.9683
R21003 a_n2848_n452.n19 a_n2848_n452.n28 75.0448
R21004 a_n2848_n452.n98 a_n2848_n452.n28 11.2134
R21005 a_n2848_n452.n20 a_n2848_n452.n21 44.8194
R21006 a_n2848_n452.n32 a_n2848_n452.n15 70.1674
R21007 a_n2848_n452.n32 a_n2848_n452.n50 20.9683
R21008 a_n2848_n452.n15 a_n2848_n452.n31 75.0448
R21009 a_n2848_n452.n101 a_n2848_n452.n31 11.2134
R21010 a_n2848_n452.n16 a_n2848_n452.n17 44.8194
R21011 a_n2848_n452.n6 a_n2848_n452.n42 70.1674
R21012 a_n2848_n452.n8 a_n2848_n452.n39 70.1674
R21013 a_n2848_n452.n10 a_n2848_n452.n37 70.1674
R21014 a_n2848_n452.n12 a_n2848_n452.n35 70.1674
R21015 a_n2848_n452.n35 a_n2848_n452.n84 20.9683
R21016 a_n2848_n452.n34 a_n2848_n452.n13 75.0448
R21017 a_n2848_n452.n94 a_n2848_n452.n34 11.2134
R21018 a_n2848_n452.n13 a_n2848_n452.n95 161.3
R21019 a_n2848_n452.n37 a_n2848_n452.n85 20.9683
R21020 a_n2848_n452.n36 a_n2848_n452.n11 75.0448
R21021 a_n2848_n452.n92 a_n2848_n452.n36 11.2134
R21022 a_n2848_n452.n11 a_n2848_n452.n93 161.3
R21023 a_n2848_n452.n39 a_n2848_n452.n86 20.9683
R21024 a_n2848_n452.n38 a_n2848_n452.n9 75.0448
R21025 a_n2848_n452.n90 a_n2848_n452.n38 11.2134
R21026 a_n2848_n452.n9 a_n2848_n452.n91 161.3
R21027 a_n2848_n452.n42 a_n2848_n452.n87 20.9683
R21028 a_n2848_n452.n40 a_n2848_n452.n7 75.0448
R21029 a_n2848_n452.n88 a_n2848_n452.n40 11.2134
R21030 a_n2848_n452.n7 a_n2848_n452.n89 161.3
R21031 a_n2848_n452.n77 a_n2848_n452.n5 161.3
R21032 a_n2848_n452.n79 a_n2848_n452.n78 161.3
R21033 a_n2848_n452.n48 a_n2848_n452.n49 20.9683
R21034 a_n2848_n452.n4 a_n2848_n452.n44 70.3058
R21035 a_n2848_n452.n43 a_n2848_n452.n5 70.1674
R21036 a_n2848_n452.n57 a_n2848_n452.n43 20.9683
R21037 a_n2848_n452.n5 a_n2848_n452.n58 161.3
R21038 a_n2848_n452.n2 a_n2848_n452.n46 70.1674
R21039 a_n2848_n452.n46 a_n2848_n452.n52 20.9683
R21040 a_n2848_n452.n45 a_n2848_n452.n2 75.0448
R21041 a_n2848_n452.n54 a_n2848_n452.n45 11.2134
R21042 a_n2848_n452.n0 a_n2848_n452.n3 44.8194
R21043 a_n2848_n452.n74 a_n2848_n452.n72 81.4626
R21044 a_n2848_n452.n65 a_n2848_n452.n63 81.4626
R21045 a_n2848_n452.n61 a_n2848_n452.n59 81.4626
R21046 a_n2848_n452.n74 a_n2848_n452.n73 80.9324
R21047 a_n2848_n452.n27 a_n2848_n452.n75 80.9324
R21048 a_n2848_n452.n26 a_n2848_n452.n71 80.9324
R21049 a_n2848_n452.n70 a_n2848_n452.n69 80.9324
R21050 a_n2848_n452.n68 a_n2848_n452.n67 80.9324
R21051 a_n2848_n452.n65 a_n2848_n452.n64 80.9324
R21052 a_n2848_n452.n25 a_n2848_n452.n66 80.9324
R21053 a_n2848_n452.n24 a_n2848_n452.n62 80.9324
R21054 a_n2848_n452.n61 a_n2848_n452.n60 80.9324
R21055 a_n2848_n452.n22 a_n2848_n452.t25 74.6477
R21056 a_n2848_n452.t11 a_n2848_n452.n106 74.6477
R21057 a_n2848_n452.n82 a_n2848_n452.t13 74.2899
R21058 a_n2848_n452.n23 a_n2848_n452.t19 74.2897
R21059 a_n2848_n452.n23 a_n2848_n452.n104 70.6783
R21060 a_n2848_n452.n106 a_n2848_n452.n105 70.6783
R21061 a_n2848_n452.n22 a_n2848_n452.n80 70.6783
R21062 a_n2848_n452.n22 a_n2848_n452.n81 70.6783
R21063 a_n2848_n452.n55 a_n2848_n452.n54 48.2005
R21064 a_n2848_n452.n53 a_n2848_n452.n46 20.9683
R21065 a_n2848_n452.n43 a_n2848_n452.n56 20.9683
R21066 a_n2848_n452.n76 a_n2848_n452.n48 20.9683
R21067 a_n2848_n452.n101 a_n2848_n452.n100 48.2005
R21068 a_n2848_n452.n102 a_n2848_n452.n32 20.9683
R21069 a_n2848_n452.n98 a_n2848_n452.n97 48.2005
R21070 a_n2848_n452.n99 a_n2848_n452.n29 20.9683
R21071 a_n2848_n452.n89 a_n2848_n452.n88 48.2005
R21072 a_n2848_n452.t69 a_n2848_n452.n42 533.335
R21073 a_n2848_n452.n91 a_n2848_n452.n90 48.2005
R21074 a_n2848_n452.t74 a_n2848_n452.n39 533.335
R21075 a_n2848_n452.n93 a_n2848_n452.n92 48.2005
R21076 a_n2848_n452.t63 a_n2848_n452.n37 533.335
R21077 a_n2848_n452.n95 a_n2848_n452.n94 48.2005
R21078 a_n2848_n452.t59 a_n2848_n452.n35 533.335
R21079 a_n2848_n452.n47 a_n2848_n452.t73 533.058
R21080 a_n2848_n452.n78 a_n2848_n452.n77 47.4702
R21081 a_n2848_n452.t18 a_n2848_n452.n33 533.058
R21082 a_n2848_n452.t51 a_n2848_n452.n30 533.058
R21083 a_n2848_n452.n68 a_n2848_n452.n25 33.585
R21084 a_n2848_n452.n45 a_n2848_n452.n52 35.3134
R21085 a_n2848_n452.n58 a_n2848_n452.n49 24.1005
R21086 a_n2848_n452.n58 a_n2848_n452.n57 24.1005
R21087 a_n2848_n452.n50 a_n2848_n452.n31 35.3134
R21088 a_n2848_n452.n51 a_n2848_n452.n28 35.3134
R21089 a_n2848_n452.n40 a_n2848_n452.n87 35.3134
R21090 a_n2848_n452.n38 a_n2848_n452.n86 35.3134
R21091 a_n2848_n452.n36 a_n2848_n452.n85 35.3134
R21092 a_n2848_n452.n34 a_n2848_n452.n84 35.3134
R21093 a_n2848_n452.n5 a_n2848_n452.n27 23.891
R21094 a_n2848_n452.n20 a_n2848_n452.n96 12.046
R21095 a_n2848_n452.n1 a_n2848_n452.n41 11.8414
R21096 a_n2848_n452.n83 a_n2848_n452.n79 10.5365
R21097 a_n2848_n452.n23 a_n2848_n452.n103 9.50122
R21098 a_n2848_n452.n6 a_n2848_n452.n41 7.47588
R21099 a_n2848_n452.n96 a_n2848_n452.n13 7.47588
R21100 a_n2848_n452.n103 a_n2848_n452.n14 6.70126
R21101 a_n2848_n452.n83 a_n2848_n452.n82 5.65783
R21102 a_n2848_n452.n103 a_n2848_n452.n41 5.3452
R21103 a_n2848_n452.n16 a_n2848_n452.n18 3.95126
R21104 a_n2848_n452.n4 a_n2848_n452.n0 3.95126
R21105 a_n2848_n452.n104 a_n2848_n452.t27 3.61217
R21106 a_n2848_n452.n104 a_n2848_n452.t29 3.61217
R21107 a_n2848_n452.n105 a_n2848_n452.t31 3.61217
R21108 a_n2848_n452.n105 a_n2848_n452.t33 3.61217
R21109 a_n2848_n452.n80 a_n2848_n452.t21 3.61217
R21110 a_n2848_n452.n80 a_n2848_n452.t15 3.61217
R21111 a_n2848_n452.n81 a_n2848_n452.t17 3.61217
R21112 a_n2848_n452.n81 a_n2848_n452.t23 3.61217
R21113 a_n2848_n452.n72 a_n2848_n452.t39 2.82907
R21114 a_n2848_n452.n72 a_n2848_n452.t43 2.82907
R21115 a_n2848_n452.n73 a_n2848_n452.t34 2.82907
R21116 a_n2848_n452.n73 a_n2848_n452.t35 2.82907
R21117 a_n2848_n452.n75 a_n2848_n452.t7 2.82907
R21118 a_n2848_n452.n75 a_n2848_n452.t8 2.82907
R21119 a_n2848_n452.n71 a_n2848_n452.t40 2.82907
R21120 a_n2848_n452.n71 a_n2848_n452.t1 2.82907
R21121 a_n2848_n452.n69 a_n2848_n452.t36 2.82907
R21122 a_n2848_n452.n69 a_n2848_n452.t37 2.82907
R21123 a_n2848_n452.n67 a_n2848_n452.t42 2.82907
R21124 a_n2848_n452.n67 a_n2848_n452.t45 2.82907
R21125 a_n2848_n452.n63 a_n2848_n452.t5 2.82907
R21126 a_n2848_n452.n63 a_n2848_n452.t6 2.82907
R21127 a_n2848_n452.n64 a_n2848_n452.t41 2.82907
R21128 a_n2848_n452.n64 a_n2848_n452.t9 2.82907
R21129 a_n2848_n452.n66 a_n2848_n452.t0 2.82907
R21130 a_n2848_n452.n66 a_n2848_n452.t38 2.82907
R21131 a_n2848_n452.n62 a_n2848_n452.t47 2.82907
R21132 a_n2848_n452.n62 a_n2848_n452.t3 2.82907
R21133 a_n2848_n452.n60 a_n2848_n452.t2 2.82907
R21134 a_n2848_n452.n60 a_n2848_n452.t46 2.82907
R21135 a_n2848_n452.n59 a_n2848_n452.t4 2.82907
R21136 a_n2848_n452.n59 a_n2848_n452.t44 2.82907
R21137 a_n2848_n452.n96 a_n2848_n452.n83 1.30542
R21138 a_n2848_n452.n10 a_n2848_n452.n9 1.04595
R21139 a_n2848_n452.n3 a_n2848_n452.n55 13.657
R21140 a_n2848_n452.n53 a_n2848_n452.n47 21.4216
R21141 a_n2848_n452.n56 a_n2848_n452.n44 21.4216
R21142 a_n2848_n452.n77 a_n2848_n452.n76 0.730803
R21143 a_n2848_n452.n100 a_n2848_n452.n17 13.657
R21144 a_n2848_n452.n33 a_n2848_n452.n102 21.4216
R21145 a_n2848_n452.n97 a_n2848_n452.n21 13.657
R21146 a_n2848_n452.n30 a_n2848_n452.n99 21.4216
R21147 a_n2848_n452.n20 a_n2848_n452.n19 0.758076
R21148 a_n2848_n452.n19 a_n2848_n452.n18 0.758076
R21149 a_n2848_n452.n16 a_n2848_n452.n15 0.758076
R21150 a_n2848_n452.n15 a_n2848_n452.n14 0.758076
R21151 a_n2848_n452.n13 a_n2848_n452.n12 0.758076
R21152 a_n2848_n452.n11 a_n2848_n452.n10 0.758076
R21153 a_n2848_n452.n9 a_n2848_n452.n8 0.758076
R21154 a_n2848_n452.n7 a_n2848_n452.n6 0.758076
R21155 a_n2848_n452.n5 a_n2848_n452.n4 0.758076
R21156 a_n2848_n452.n2 a_n2848_n452.n0 0.758076
R21157 a_n2848_n452.n2 a_n2848_n452.n1 0.758076
R21158 a_n2848_n452.n79 a_n2848_n452.n5 0.720197
R21159 a_n2848_n452.n106 a_n2848_n452.n23 0.716017
R21160 a_n2848_n452.n82 a_n2848_n452.n22 0.716017
R21161 a_n2848_n452.n12 a_n2848_n452.n11 0.67853
R21162 a_n2848_n452.n8 a_n2848_n452.n7 0.67853
R21163 a_n2848_n452.n24 a_n2848_n452.n61 0.530672
R21164 a_n2848_n452.n25 a_n2848_n452.n65 0.530672
R21165 a_n2848_n452.n70 a_n2848_n452.n68 0.530672
R21166 a_n2848_n452.n26 a_n2848_n452.n70 0.530672
R21167 a_n2848_n452.n27 a_n2848_n452.n74 0.530672
R21168 a_n2848_n452.n27 a_n2848_n452.n26 0.530672
R21169 a_n2848_n452.n25 a_n2848_n452.n24 0.530672
R21170 a_n1986_8322.n6 a_n1986_8322.t18 74.6477
R21171 a_n1986_8322.n1 a_n1986_8322.t5 74.6477
R21172 a_n1986_8322.n16 a_n1986_8322.t14 74.6474
R21173 a_n1986_8322.n14 a_n1986_8322.t7 74.2899
R21174 a_n1986_8322.n7 a_n1986_8322.t16 74.2899
R21175 a_n1986_8322.n8 a_n1986_8322.t19 74.2899
R21176 a_n1986_8322.n11 a_n1986_8322.t20 74.2899
R21177 a_n1986_8322.n4 a_n1986_8322.t4 74.2899
R21178 a_n1986_8322.n16 a_n1986_8322.n15 70.6783
R21179 a_n1986_8322.n6 a_n1986_8322.n5 70.6783
R21180 a_n1986_8322.n10 a_n1986_8322.n9 70.6783
R21181 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R21182 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R21183 a_n1986_8322.n18 a_n1986_8322.n17 70.6782
R21184 a_n1986_8322.n12 a_n1986_8322.n4 22.7556
R21185 a_n1986_8322.n13 a_n1986_8322.t0 9.94227
R21186 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R21187 a_n1986_8322.n14 a_n1986_8322.n13 5.83671
R21188 a_n1986_8322.n13 a_n1986_8322.n12 5.3452
R21189 a_n1986_8322.n15 a_n1986_8322.t12 3.61217
R21190 a_n1986_8322.n15 a_n1986_8322.t9 3.61217
R21191 a_n1986_8322.n5 a_n1986_8322.t22 3.61217
R21192 a_n1986_8322.n5 a_n1986_8322.t21 3.61217
R21193 a_n1986_8322.n9 a_n1986_8322.t17 3.61217
R21194 a_n1986_8322.n9 a_n1986_8322.t23 3.61217
R21195 a_n1986_8322.n0 a_n1986_8322.t13 3.61217
R21196 a_n1986_8322.n0 a_n1986_8322.t8 3.61217
R21197 a_n1986_8322.n2 a_n1986_8322.t11 3.61217
R21198 a_n1986_8322.n2 a_n1986_8322.t10 3.61217
R21199 a_n1986_8322.n18 a_n1986_8322.t6 3.61217
R21200 a_n1986_8322.t15 a_n1986_8322.n18 3.61217
R21201 a_n1986_8322.n11 a_n1986_8322.n10 0.358259
R21202 a_n1986_8322.n10 a_n1986_8322.n8 0.358259
R21203 a_n1986_8322.n7 a_n1986_8322.n6 0.358259
R21204 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R21205 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R21206 a_n1986_8322.n17 a_n1986_8322.n14 0.358259
R21207 a_n1986_8322.n17 a_n1986_8322.n16 0.358259
R21208 a_n1986_8322.n8 a_n1986_8322.n7 0.101793
R21209 a_n1986_8322.t3 a_n1986_8322.t2 0.0788333
R21210 a_n1986_8322.t1 a_n1986_8322.t3 0.0631667
R21211 a_n1986_8322.t0 a_n1986_8322.t1 0.0471944
R21212 a_n1986_8322.t0 a_n1986_8322.t2 0.0453889
R21213 a_n1808_13878.n5 a_n1808_13878.n3 98.9633
R21214 a_n1808_13878.n2 a_n1808_13878.n0 98.7517
R21215 a_n1808_13878.n2 a_n1808_13878.n1 98.6055
R21216 a_n1808_13878.n5 a_n1808_13878.n4 98.6055
R21217 a_n1808_13878.n17 a_n1808_13878.n16 98.6054
R21218 a_n1808_13878.n7 a_n1808_13878.n6 98.6054
R21219 a_n1808_13878.n9 a_n1808_13878.t13 74.6477
R21220 a_n1808_13878.n14 a_n1808_13878.t14 74.2899
R21221 a_n1808_13878.n11 a_n1808_13878.t15 74.2899
R21222 a_n1808_13878.n10 a_n1808_13878.t12 74.2899
R21223 a_n1808_13878.n13 a_n1808_13878.n12 70.6783
R21224 a_n1808_13878.n9 a_n1808_13878.n8 70.6783
R21225 a_n1808_13878.n16 a_n1808_13878.n15 13.5694
R21226 a_n1808_13878.n15 a_n1808_13878.n7 11.5762
R21227 a_n1808_13878.n15 a_n1808_13878.n14 6.2408
R21228 a_n1808_13878.n1 a_n1808_13878.t6 3.61217
R21229 a_n1808_13878.n1 a_n1808_13878.t1 3.61217
R21230 a_n1808_13878.n0 a_n1808_13878.t0 3.61217
R21231 a_n1808_13878.n0 a_n1808_13878.t2 3.61217
R21232 a_n1808_13878.n6 a_n1808_13878.t7 3.61217
R21233 a_n1808_13878.n6 a_n1808_13878.t8 3.61217
R21234 a_n1808_13878.n4 a_n1808_13878.t10 3.61217
R21235 a_n1808_13878.n4 a_n1808_13878.t3 3.61217
R21236 a_n1808_13878.n3 a_n1808_13878.t5 3.61217
R21237 a_n1808_13878.n3 a_n1808_13878.t9 3.61217
R21238 a_n1808_13878.n12 a_n1808_13878.t18 3.61217
R21239 a_n1808_13878.n12 a_n1808_13878.t19 3.61217
R21240 a_n1808_13878.n8 a_n1808_13878.t16 3.61217
R21241 a_n1808_13878.n8 a_n1808_13878.t17 3.61217
R21242 a_n1808_13878.n17 a_n1808_13878.t4 3.61217
R21243 a_n1808_13878.t11 a_n1808_13878.n17 3.61217
R21244 a_n1808_13878.n7 a_n1808_13878.n5 0.358259
R21245 a_n1808_13878.n10 a_n1808_13878.n9 0.358259
R21246 a_n1808_13878.n13 a_n1808_13878.n11 0.358259
R21247 a_n1808_13878.n14 a_n1808_13878.n13 0.358259
R21248 a_n1808_13878.n16 a_n1808_13878.n2 0.146627
R21249 a_n1808_13878.n11 a_n1808_13878.n10 0.101793
R21250 plus.n76 plus.t11 250.337
R21251 plus.n15 plus.t14 250.337
R21252 plus.n124 plus.t1 243.97
R21253 plus.n120 plus.t24 231.093
R21254 plus.n59 plus.t20 231.093
R21255 plus.n124 plus.n123 223.454
R21256 plus.n126 plus.n125 223.454
R21257 plus.n77 plus.t5 187.445
R21258 plus.n74 plus.t22 187.445
R21259 plus.n72 plus.t21 187.445
R21260 plus.n89 plus.t16 187.445
R21261 plus.n95 plus.t17 187.445
R21262 plus.n68 plus.t13 187.445
R21263 plus.n66 plus.t15 187.445
R21264 plus.n107 plus.t10 187.445
R21265 plus.n113 plus.t26 187.445
R21266 plus.n62 plus.t28 187.445
R21267 plus.n1 plus.t23 187.445
R21268 plus.n52 plus.t6 187.445
R21269 plus.n46 plus.t12 187.445
R21270 plus.n5 plus.t8 187.445
R21271 plus.n7 plus.t7 187.445
R21272 plus.n34 plus.t19 187.445
R21273 plus.n28 plus.t18 187.445
R21274 plus.n11 plus.t27 187.445
R21275 plus.n13 plus.t25 187.445
R21276 plus.n16 plus.t9 187.445
R21277 plus.n121 plus.n120 161.3
R21278 plus.n119 plus.n61 161.3
R21279 plus.n118 plus.n117 161.3
R21280 plus.n116 plus.n115 161.3
R21281 plus.n114 plus.n63 161.3
R21282 plus.n112 plus.n111 161.3
R21283 plus.n110 plus.n64 161.3
R21284 plus.n109 plus.n108 161.3
R21285 plus.n106 plus.n65 161.3
R21286 plus.n105 plus.n104 161.3
R21287 plus.n103 plus.n102 161.3
R21288 plus.n101 plus.n67 161.3
R21289 plus.n100 plus.n99 161.3
R21290 plus.n98 plus.n97 161.3
R21291 plus.n96 plus.n69 161.3
R21292 plus.n94 plus.n93 161.3
R21293 plus.n92 plus.n70 161.3
R21294 plus.n91 plus.n90 161.3
R21295 plus.n88 plus.n71 161.3
R21296 plus.n87 plus.n86 161.3
R21297 plus.n85 plus.n84 161.3
R21298 plus.n83 plus.n73 161.3
R21299 plus.n82 plus.n81 161.3
R21300 plus.n80 plus.n79 161.3
R21301 plus.n78 plus.n75 161.3
R21302 plus.n17 plus.n14 161.3
R21303 plus.n19 plus.n18 161.3
R21304 plus.n21 plus.n20 161.3
R21305 plus.n22 plus.n12 161.3
R21306 plus.n24 plus.n23 161.3
R21307 plus.n26 plus.n25 161.3
R21308 plus.n27 plus.n10 161.3
R21309 plus.n30 plus.n29 161.3
R21310 plus.n31 plus.n9 161.3
R21311 plus.n33 plus.n32 161.3
R21312 plus.n35 plus.n8 161.3
R21313 plus.n37 plus.n36 161.3
R21314 plus.n39 plus.n38 161.3
R21315 plus.n40 plus.n6 161.3
R21316 plus.n42 plus.n41 161.3
R21317 plus.n44 plus.n43 161.3
R21318 plus.n45 plus.n4 161.3
R21319 plus.n48 plus.n47 161.3
R21320 plus.n49 plus.n3 161.3
R21321 plus.n51 plus.n50 161.3
R21322 plus.n53 plus.n2 161.3
R21323 plus.n55 plus.n54 161.3
R21324 plus.n57 plus.n56 161.3
R21325 plus.n58 plus.n0 161.3
R21326 plus.n60 plus.n59 161.3
R21327 plus.n88 plus.n87 56.5617
R21328 plus.n97 plus.n96 56.5617
R21329 plus.n106 plus.n105 56.5617
R21330 plus.n45 plus.n44 56.5617
R21331 plus.n36 plus.n35 56.5617
R21332 plus.n27 plus.n26 56.5617
R21333 plus.n79 plus.n78 56.5617
R21334 plus.n115 plus.n114 56.5617
R21335 plus.n54 plus.n53 56.5617
R21336 plus.n18 plus.n17 56.5617
R21337 plus.n119 plus.n118 50.2647
R21338 plus.n58 plus.n57 50.2647
R21339 plus.n84 plus.n83 46.3896
R21340 plus.n108 plus.n64 46.3896
R21341 plus.n47 plus.n3 46.3896
R21342 plus.n23 plus.n22 46.3896
R21343 plus.n76 plus.n75 43.1929
R21344 plus.n15 plus.n14 43.1929
R21345 plus.n94 plus.n70 42.5146
R21346 plus.n101 plus.n100 42.5146
R21347 plus.n40 plus.n39 42.5146
R21348 plus.n33 plus.n9 42.5146
R21349 plus.n77 plus.n76 40.6041
R21350 plus.n16 plus.n15 40.6041
R21351 plus.n90 plus.n70 38.6395
R21352 plus.n102 plus.n101 38.6395
R21353 plus.n41 plus.n40 38.6395
R21354 plus.n29 plus.n9 38.6395
R21355 plus.n122 plus.n121 35.2031
R21356 plus.n83 plus.n82 34.7644
R21357 plus.n112 plus.n64 34.7644
R21358 plus.n51 plus.n3 34.7644
R21359 plus.n22 plus.n21 34.7644
R21360 plus.n79 plus.n74 21.8872
R21361 plus.n114 plus.n113 21.8872
R21362 plus.n53 plus.n52 21.8872
R21363 plus.n18 plus.n13 21.8872
R21364 plus.n89 plus.n88 19.9199
R21365 plus.n105 plus.n66 19.9199
R21366 plus.n44 plus.n5 19.9199
R21367 plus.n28 plus.n27 19.9199
R21368 plus.n123 plus.t2 19.8005
R21369 plus.n123 plus.t4 19.8005
R21370 plus.n125 plus.t3 19.8005
R21371 plus.n125 plus.t0 19.8005
R21372 plus.n96 plus.n95 17.9525
R21373 plus.n97 plus.n68 17.9525
R21374 plus.n36 plus.n7 17.9525
R21375 plus.n35 plus.n34 17.9525
R21376 plus.n87 plus.n72 15.9852
R21377 plus.n107 plus.n106 15.9852
R21378 plus.n46 plus.n45 15.9852
R21379 plus.n26 plus.n11 15.9852
R21380 plus plus.n127 14.6928
R21381 plus.n78 plus.n77 14.0178
R21382 plus.n115 plus.n62 14.0178
R21383 plus.n54 plus.n1 14.0178
R21384 plus.n17 plus.n16 14.0178
R21385 plus.n122 plus.n60 11.9342
R21386 plus.n118 plus.n62 10.575
R21387 plus.n57 plus.n1 10.575
R21388 plus.n120 plus.n119 9.49444
R21389 plus.n59 plus.n58 9.49444
R21390 plus.n84 plus.n72 8.60764
R21391 plus.n108 plus.n107 8.60764
R21392 plus.n47 plus.n46 8.60764
R21393 plus.n23 plus.n11 8.60764
R21394 plus.n95 plus.n94 6.6403
R21395 plus.n100 plus.n68 6.6403
R21396 plus.n39 plus.n7 6.6403
R21397 plus.n34 plus.n33 6.6403
R21398 plus.n127 plus.n126 5.40567
R21399 plus.n90 plus.n89 4.67295
R21400 plus.n102 plus.n66 4.67295
R21401 plus.n41 plus.n5 4.67295
R21402 plus.n29 plus.n28 4.67295
R21403 plus.n82 plus.n74 2.7056
R21404 plus.n113 plus.n112 2.7056
R21405 plus.n52 plus.n51 2.7056
R21406 plus.n21 plus.n13 2.7056
R21407 plus.n127 plus.n122 1.188
R21408 plus.n126 plus.n124 0.716017
R21409 plus.n80 plus.n75 0.189894
R21410 plus.n81 plus.n80 0.189894
R21411 plus.n81 plus.n73 0.189894
R21412 plus.n85 plus.n73 0.189894
R21413 plus.n86 plus.n85 0.189894
R21414 plus.n86 plus.n71 0.189894
R21415 plus.n91 plus.n71 0.189894
R21416 plus.n92 plus.n91 0.189894
R21417 plus.n93 plus.n92 0.189894
R21418 plus.n93 plus.n69 0.189894
R21419 plus.n98 plus.n69 0.189894
R21420 plus.n99 plus.n98 0.189894
R21421 plus.n99 plus.n67 0.189894
R21422 plus.n103 plus.n67 0.189894
R21423 plus.n104 plus.n103 0.189894
R21424 plus.n104 plus.n65 0.189894
R21425 plus.n109 plus.n65 0.189894
R21426 plus.n110 plus.n109 0.189894
R21427 plus.n111 plus.n110 0.189894
R21428 plus.n111 plus.n63 0.189894
R21429 plus.n116 plus.n63 0.189894
R21430 plus.n117 plus.n116 0.189894
R21431 plus.n117 plus.n61 0.189894
R21432 plus.n121 plus.n61 0.189894
R21433 plus.n60 plus.n0 0.189894
R21434 plus.n56 plus.n0 0.189894
R21435 plus.n56 plus.n55 0.189894
R21436 plus.n55 plus.n2 0.189894
R21437 plus.n50 plus.n2 0.189894
R21438 plus.n50 plus.n49 0.189894
R21439 plus.n49 plus.n48 0.189894
R21440 plus.n48 plus.n4 0.189894
R21441 plus.n43 plus.n4 0.189894
R21442 plus.n43 plus.n42 0.189894
R21443 plus.n42 plus.n6 0.189894
R21444 plus.n38 plus.n6 0.189894
R21445 plus.n38 plus.n37 0.189894
R21446 plus.n37 plus.n8 0.189894
R21447 plus.n32 plus.n8 0.189894
R21448 plus.n32 plus.n31 0.189894
R21449 plus.n31 plus.n30 0.189894
R21450 plus.n30 plus.n10 0.189894
R21451 plus.n25 plus.n10 0.189894
R21452 plus.n25 plus.n24 0.189894
R21453 plus.n24 plus.n12 0.189894
R21454 plus.n20 plus.n12 0.189894
R21455 plus.n20 plus.n19 0.189894
R21456 plus.n19 plus.n14 0.189894
R21457 a_n3827_n3924.n22 a_n3827_n3924.t0 214.938
R21458 a_n3827_n3924.n1 a_n3827_n3924.t57 214.409
R21459 a_n3827_n3924.n14 a_n3827_n3924.t52 214.321
R21460 a_n3827_n3924.n15 a_n3827_n3924.t46 214.321
R21461 a_n3827_n3924.n16 a_n3827_n3924.t12 214.321
R21462 a_n3827_n3924.n17 a_n3827_n3924.t48 214.321
R21463 a_n3827_n3924.n18 a_n3827_n3924.t49 214.321
R21464 a_n3827_n3924.n19 a_n3827_n3924.t51 214.321
R21465 a_n3827_n3924.n20 a_n3827_n3924.t45 214.321
R21466 a_n3827_n3924.n21 a_n3827_n3924.t6 214.321
R21467 a_n3827_n3924.n0 a_n3827_n3924.t32 55.8337
R21468 a_n3827_n3924.n2 a_n3827_n3924.t50 55.8337
R21469 a_n3827_n3924.n13 a_n3827_n3924.t47 55.8337
R21470 a_n3827_n3924.n49 a_n3827_n3924.t19 55.8335
R21471 a_n3827_n3924.n47 a_n3827_n3924.t8 55.8335
R21472 a_n3827_n3924.n36 a_n3827_n3924.t5 55.8335
R21473 a_n3827_n3924.n35 a_n3827_n3924.t29 55.8335
R21474 a_n3827_n3924.n24 a_n3827_n3924.t23 55.8335
R21475 a_n3827_n3924.n51 a_n3827_n3924.n50 53.0052
R21476 a_n3827_n3924.n53 a_n3827_n3924.n52 53.0052
R21477 a_n3827_n3924.n55 a_n3827_n3924.n54 53.0052
R21478 a_n3827_n3924.n57 a_n3827_n3924.n56 53.0052
R21479 a_n3827_n3924.n4 a_n3827_n3924.n3 53.0052
R21480 a_n3827_n3924.n6 a_n3827_n3924.n5 53.0052
R21481 a_n3827_n3924.n8 a_n3827_n3924.n7 53.0052
R21482 a_n3827_n3924.n10 a_n3827_n3924.n9 53.0052
R21483 a_n3827_n3924.n12 a_n3827_n3924.n11 53.0052
R21484 a_n3827_n3924.n46 a_n3827_n3924.n45 53.0051
R21485 a_n3827_n3924.n44 a_n3827_n3924.n43 53.0051
R21486 a_n3827_n3924.n42 a_n3827_n3924.n41 53.0051
R21487 a_n3827_n3924.n40 a_n3827_n3924.n39 53.0051
R21488 a_n3827_n3924.n38 a_n3827_n3924.n37 53.0051
R21489 a_n3827_n3924.n34 a_n3827_n3924.n33 53.0051
R21490 a_n3827_n3924.n32 a_n3827_n3924.n31 53.0051
R21491 a_n3827_n3924.n30 a_n3827_n3924.n29 53.0051
R21492 a_n3827_n3924.n28 a_n3827_n3924.n27 53.0051
R21493 a_n3827_n3924.n26 a_n3827_n3924.n25 53.0051
R21494 a_n3827_n3924.n59 a_n3827_n3924.n58 53.0051
R21495 a_n3827_n3924.n23 a_n3827_n3924.n13 12.2417
R21496 a_n3827_n3924.n49 a_n3827_n3924.n48 12.2417
R21497 a_n3827_n3924.n24 a_n3827_n3924.n23 5.16214
R21498 a_n3827_n3924.n48 a_n3827_n3924.n47 5.16214
R21499 a_n3827_n3924.n50 a_n3827_n3924.t17 2.82907
R21500 a_n3827_n3924.n50 a_n3827_n3924.t15 2.82907
R21501 a_n3827_n3924.n52 a_n3827_n3924.t28 2.82907
R21502 a_n3827_n3924.n52 a_n3827_n3924.t33 2.82907
R21503 a_n3827_n3924.n54 a_n3827_n3924.t26 2.82907
R21504 a_n3827_n3924.n54 a_n3827_n3924.t30 2.82907
R21505 a_n3827_n3924.n56 a_n3827_n3924.t22 2.82907
R21506 a_n3827_n3924.n56 a_n3827_n3924.t27 2.82907
R21507 a_n3827_n3924.n3 a_n3827_n3924.t14 2.82907
R21508 a_n3827_n3924.n3 a_n3827_n3924.t42 2.82907
R21509 a_n3827_n3924.n5 a_n3827_n3924.t10 2.82907
R21510 a_n3827_n3924.n5 a_n3827_n3924.t13 2.82907
R21511 a_n3827_n3924.n7 a_n3827_n3924.t2 2.82907
R21512 a_n3827_n3924.n7 a_n3827_n3924.t9 2.82907
R21513 a_n3827_n3924.n9 a_n3827_n3924.t40 2.82907
R21514 a_n3827_n3924.n9 a_n3827_n3924.t43 2.82907
R21515 a_n3827_n3924.n11 a_n3827_n3924.t54 2.82907
R21516 a_n3827_n3924.n11 a_n3827_n3924.t39 2.82907
R21517 a_n3827_n3924.n45 a_n3827_n3924.t11 2.82907
R21518 a_n3827_n3924.n45 a_n3827_n3924.t7 2.82907
R21519 a_n3827_n3924.n43 a_n3827_n3924.t41 2.82907
R21520 a_n3827_n3924.n43 a_n3827_n3924.t44 2.82907
R21521 a_n3827_n3924.n41 a_n3827_n3924.t4 2.82907
R21522 a_n3827_n3924.n41 a_n3827_n3924.t1 2.82907
R21523 a_n3827_n3924.n39 a_n3827_n3924.t55 2.82907
R21524 a_n3827_n3924.n39 a_n3827_n3924.t56 2.82907
R21525 a_n3827_n3924.n37 a_n3827_n3924.t53 2.82907
R21526 a_n3827_n3924.n37 a_n3827_n3924.t3 2.82907
R21527 a_n3827_n3924.n33 a_n3827_n3924.t18 2.82907
R21528 a_n3827_n3924.n33 a_n3827_n3924.t34 2.82907
R21529 a_n3827_n3924.n31 a_n3827_n3924.t25 2.82907
R21530 a_n3827_n3924.n31 a_n3827_n3924.t16 2.82907
R21531 a_n3827_n3924.n29 a_n3827_n3924.t36 2.82907
R21532 a_n3827_n3924.n29 a_n3827_n3924.t24 2.82907
R21533 a_n3827_n3924.n27 a_n3827_n3924.t31 2.82907
R21534 a_n3827_n3924.n27 a_n3827_n3924.t35 2.82907
R21535 a_n3827_n3924.n25 a_n3827_n3924.t20 2.82907
R21536 a_n3827_n3924.n25 a_n3827_n3924.t37 2.82907
R21537 a_n3827_n3924.t38 a_n3827_n3924.n59 2.82907
R21538 a_n3827_n3924.n59 a_n3827_n3924.t21 2.82907
R21539 a_n3827_n3924.n48 a_n3827_n3924.n1 1.95694
R21540 a_n3827_n3924.n23 a_n3827_n3924.n22 1.95694
R21541 a_n3827_n3924.n21 a_n3827_n3924.n20 0.672012
R21542 a_n3827_n3924.n20 a_n3827_n3924.n19 0.672012
R21543 a_n3827_n3924.n19 a_n3827_n3924.n18 0.672012
R21544 a_n3827_n3924.n18 a_n3827_n3924.n17 0.672012
R21545 a_n3827_n3924.n17 a_n3827_n3924.n16 0.672012
R21546 a_n3827_n3924.n16 a_n3827_n3924.n15 0.672012
R21547 a_n3827_n3924.n15 a_n3827_n3924.n14 0.672012
R21548 a_n3827_n3924.n14 a_n3827_n3924.n1 0.585529
R21549 a_n3827_n3924.n26 a_n3827_n3924.n24 0.530672
R21550 a_n3827_n3924.n28 a_n3827_n3924.n26 0.530672
R21551 a_n3827_n3924.n30 a_n3827_n3924.n28 0.530672
R21552 a_n3827_n3924.n32 a_n3827_n3924.n30 0.530672
R21553 a_n3827_n3924.n34 a_n3827_n3924.n32 0.530672
R21554 a_n3827_n3924.n35 a_n3827_n3924.n34 0.530672
R21555 a_n3827_n3924.n38 a_n3827_n3924.n36 0.530672
R21556 a_n3827_n3924.n40 a_n3827_n3924.n38 0.530672
R21557 a_n3827_n3924.n42 a_n3827_n3924.n40 0.530672
R21558 a_n3827_n3924.n44 a_n3827_n3924.n42 0.530672
R21559 a_n3827_n3924.n46 a_n3827_n3924.n44 0.530672
R21560 a_n3827_n3924.n47 a_n3827_n3924.n46 0.530672
R21561 a_n3827_n3924.n13 a_n3827_n3924.n12 0.530672
R21562 a_n3827_n3924.n12 a_n3827_n3924.n10 0.530672
R21563 a_n3827_n3924.n10 a_n3827_n3924.n8 0.530672
R21564 a_n3827_n3924.n8 a_n3827_n3924.n6 0.530672
R21565 a_n3827_n3924.n6 a_n3827_n3924.n4 0.530672
R21566 a_n3827_n3924.n4 a_n3827_n3924.n2 0.530672
R21567 a_n3827_n3924.n58 a_n3827_n3924.n0 0.530672
R21568 a_n3827_n3924.n58 a_n3827_n3924.n57 0.530672
R21569 a_n3827_n3924.n57 a_n3827_n3924.n55 0.530672
R21570 a_n3827_n3924.n55 a_n3827_n3924.n53 0.530672
R21571 a_n3827_n3924.n53 a_n3827_n3924.n51 0.530672
R21572 a_n3827_n3924.n51 a_n3827_n3924.n49 0.530672
R21573 a_n3827_n3924.n36 a_n3827_n3924.n35 0.235414
R21574 a_n3827_n3924.n2 a_n3827_n3924.n0 0.235414
R21575 a_n3827_n3924.n22 a_n3827_n3924.n21 0.0564593
R21576 diffpairibias.n0 diffpairibias.t27 436.822
R21577 diffpairibias.n27 diffpairibias.t24 435.479
R21578 diffpairibias.n26 diffpairibias.t21 435.479
R21579 diffpairibias.n25 diffpairibias.t22 435.479
R21580 diffpairibias.n24 diffpairibias.t26 435.479
R21581 diffpairibias.n23 diffpairibias.t20 435.479
R21582 diffpairibias.n0 diffpairibias.t23 435.479
R21583 diffpairibias.n1 diffpairibias.t28 435.479
R21584 diffpairibias.n2 diffpairibias.t25 435.479
R21585 diffpairibias.n3 diffpairibias.t29 435.479
R21586 diffpairibias.n13 diffpairibias.t14 377.536
R21587 diffpairibias.n13 diffpairibias.t0 376.193
R21588 diffpairibias.n14 diffpairibias.t10 376.193
R21589 diffpairibias.n15 diffpairibias.t12 376.193
R21590 diffpairibias.n16 diffpairibias.t6 376.193
R21591 diffpairibias.n17 diffpairibias.t2 376.193
R21592 diffpairibias.n18 diffpairibias.t16 376.193
R21593 diffpairibias.n19 diffpairibias.t4 376.193
R21594 diffpairibias.n20 diffpairibias.t18 376.193
R21595 diffpairibias.n21 diffpairibias.t8 376.193
R21596 diffpairibias.n4 diffpairibias.t15 113.368
R21597 diffpairibias.n4 diffpairibias.t1 112.698
R21598 diffpairibias.n5 diffpairibias.t11 112.698
R21599 diffpairibias.n6 diffpairibias.t13 112.698
R21600 diffpairibias.n7 diffpairibias.t7 112.698
R21601 diffpairibias.n8 diffpairibias.t3 112.698
R21602 diffpairibias.n9 diffpairibias.t17 112.698
R21603 diffpairibias.n10 diffpairibias.t5 112.698
R21604 diffpairibias.n11 diffpairibias.t19 112.698
R21605 diffpairibias.n12 diffpairibias.t9 112.698
R21606 diffpairibias.n22 diffpairibias.n21 4.77242
R21607 diffpairibias.n22 diffpairibias.n12 4.30807
R21608 diffpairibias.n23 diffpairibias.n22 4.13945
R21609 diffpairibias.n21 diffpairibias.n20 1.34352
R21610 diffpairibias.n20 diffpairibias.n19 1.34352
R21611 diffpairibias.n19 diffpairibias.n18 1.34352
R21612 diffpairibias.n18 diffpairibias.n17 1.34352
R21613 diffpairibias.n17 diffpairibias.n16 1.34352
R21614 diffpairibias.n16 diffpairibias.n15 1.34352
R21615 diffpairibias.n15 diffpairibias.n14 1.34352
R21616 diffpairibias.n14 diffpairibias.n13 1.34352
R21617 diffpairibias.n3 diffpairibias.n2 1.34352
R21618 diffpairibias.n2 diffpairibias.n1 1.34352
R21619 diffpairibias.n1 diffpairibias.n0 1.34352
R21620 diffpairibias.n24 diffpairibias.n23 1.34352
R21621 diffpairibias.n25 diffpairibias.n24 1.34352
R21622 diffpairibias.n26 diffpairibias.n25 1.34352
R21623 diffpairibias.n27 diffpairibias.n26 1.34352
R21624 diffpairibias.n28 diffpairibias.n27 0.862419
R21625 diffpairibias diffpairibias.n28 0.684875
R21626 diffpairibias.n12 diffpairibias.n11 0.672012
R21627 diffpairibias.n11 diffpairibias.n10 0.672012
R21628 diffpairibias.n10 diffpairibias.n9 0.672012
R21629 diffpairibias.n9 diffpairibias.n8 0.672012
R21630 diffpairibias.n8 diffpairibias.n7 0.672012
R21631 diffpairibias.n7 diffpairibias.n6 0.672012
R21632 diffpairibias.n6 diffpairibias.n5 0.672012
R21633 diffpairibias.n5 diffpairibias.n4 0.672012
R21634 diffpairibias.n28 diffpairibias.n3 0.190907
R21635 outputibias.n27 outputibias.n1 289.615
R21636 outputibias.n58 outputibias.n32 289.615
R21637 outputibias.n90 outputibias.n64 289.615
R21638 outputibias.n122 outputibias.n96 289.615
R21639 outputibias.n28 outputibias.n27 185
R21640 outputibias.n26 outputibias.n25 185
R21641 outputibias.n5 outputibias.n4 185
R21642 outputibias.n20 outputibias.n19 185
R21643 outputibias.n18 outputibias.n17 185
R21644 outputibias.n9 outputibias.n8 185
R21645 outputibias.n12 outputibias.n11 185
R21646 outputibias.n59 outputibias.n58 185
R21647 outputibias.n57 outputibias.n56 185
R21648 outputibias.n36 outputibias.n35 185
R21649 outputibias.n51 outputibias.n50 185
R21650 outputibias.n49 outputibias.n48 185
R21651 outputibias.n40 outputibias.n39 185
R21652 outputibias.n43 outputibias.n42 185
R21653 outputibias.n91 outputibias.n90 185
R21654 outputibias.n89 outputibias.n88 185
R21655 outputibias.n68 outputibias.n67 185
R21656 outputibias.n83 outputibias.n82 185
R21657 outputibias.n81 outputibias.n80 185
R21658 outputibias.n72 outputibias.n71 185
R21659 outputibias.n75 outputibias.n74 185
R21660 outputibias.n123 outputibias.n122 185
R21661 outputibias.n121 outputibias.n120 185
R21662 outputibias.n100 outputibias.n99 185
R21663 outputibias.n115 outputibias.n114 185
R21664 outputibias.n113 outputibias.n112 185
R21665 outputibias.n104 outputibias.n103 185
R21666 outputibias.n107 outputibias.n106 185
R21667 outputibias.n0 outputibias.t10 178.945
R21668 outputibias.n133 outputibias.t8 177.018
R21669 outputibias.n132 outputibias.t11 177.018
R21670 outputibias.n0 outputibias.t9 177.018
R21671 outputibias.t7 outputibias.n10 147.661
R21672 outputibias.t1 outputibias.n41 147.661
R21673 outputibias.t3 outputibias.n73 147.661
R21674 outputibias.t5 outputibias.n105 147.661
R21675 outputibias.n128 outputibias.t6 132.363
R21676 outputibias.n128 outputibias.t0 130.436
R21677 outputibias.n129 outputibias.t2 130.436
R21678 outputibias.n130 outputibias.t4 130.436
R21679 outputibias.n27 outputibias.n26 104.615
R21680 outputibias.n26 outputibias.n4 104.615
R21681 outputibias.n19 outputibias.n4 104.615
R21682 outputibias.n19 outputibias.n18 104.615
R21683 outputibias.n18 outputibias.n8 104.615
R21684 outputibias.n11 outputibias.n8 104.615
R21685 outputibias.n58 outputibias.n57 104.615
R21686 outputibias.n57 outputibias.n35 104.615
R21687 outputibias.n50 outputibias.n35 104.615
R21688 outputibias.n50 outputibias.n49 104.615
R21689 outputibias.n49 outputibias.n39 104.615
R21690 outputibias.n42 outputibias.n39 104.615
R21691 outputibias.n90 outputibias.n89 104.615
R21692 outputibias.n89 outputibias.n67 104.615
R21693 outputibias.n82 outputibias.n67 104.615
R21694 outputibias.n82 outputibias.n81 104.615
R21695 outputibias.n81 outputibias.n71 104.615
R21696 outputibias.n74 outputibias.n71 104.615
R21697 outputibias.n122 outputibias.n121 104.615
R21698 outputibias.n121 outputibias.n99 104.615
R21699 outputibias.n114 outputibias.n99 104.615
R21700 outputibias.n114 outputibias.n113 104.615
R21701 outputibias.n113 outputibias.n103 104.615
R21702 outputibias.n106 outputibias.n103 104.615
R21703 outputibias.n63 outputibias.n31 95.6354
R21704 outputibias.n63 outputibias.n62 94.6732
R21705 outputibias.n95 outputibias.n94 94.6732
R21706 outputibias.n127 outputibias.n126 94.6732
R21707 outputibias.n11 outputibias.t7 52.3082
R21708 outputibias.n42 outputibias.t1 52.3082
R21709 outputibias.n74 outputibias.t3 52.3082
R21710 outputibias.n106 outputibias.t5 52.3082
R21711 outputibias.n12 outputibias.n10 15.6674
R21712 outputibias.n43 outputibias.n41 15.6674
R21713 outputibias.n75 outputibias.n73 15.6674
R21714 outputibias.n107 outputibias.n105 15.6674
R21715 outputibias.n13 outputibias.n9 12.8005
R21716 outputibias.n44 outputibias.n40 12.8005
R21717 outputibias.n76 outputibias.n72 12.8005
R21718 outputibias.n108 outputibias.n104 12.8005
R21719 outputibias.n17 outputibias.n16 12.0247
R21720 outputibias.n48 outputibias.n47 12.0247
R21721 outputibias.n80 outputibias.n79 12.0247
R21722 outputibias.n112 outputibias.n111 12.0247
R21723 outputibias.n20 outputibias.n7 11.249
R21724 outputibias.n51 outputibias.n38 11.249
R21725 outputibias.n83 outputibias.n70 11.249
R21726 outputibias.n115 outputibias.n102 11.249
R21727 outputibias.n21 outputibias.n5 10.4732
R21728 outputibias.n52 outputibias.n36 10.4732
R21729 outputibias.n84 outputibias.n68 10.4732
R21730 outputibias.n116 outputibias.n100 10.4732
R21731 outputibias.n25 outputibias.n24 9.69747
R21732 outputibias.n56 outputibias.n55 9.69747
R21733 outputibias.n88 outputibias.n87 9.69747
R21734 outputibias.n120 outputibias.n119 9.69747
R21735 outputibias.n31 outputibias.n30 9.45567
R21736 outputibias.n62 outputibias.n61 9.45567
R21737 outputibias.n94 outputibias.n93 9.45567
R21738 outputibias.n126 outputibias.n125 9.45567
R21739 outputibias.n30 outputibias.n29 9.3005
R21740 outputibias.n3 outputibias.n2 9.3005
R21741 outputibias.n24 outputibias.n23 9.3005
R21742 outputibias.n22 outputibias.n21 9.3005
R21743 outputibias.n7 outputibias.n6 9.3005
R21744 outputibias.n16 outputibias.n15 9.3005
R21745 outputibias.n14 outputibias.n13 9.3005
R21746 outputibias.n61 outputibias.n60 9.3005
R21747 outputibias.n34 outputibias.n33 9.3005
R21748 outputibias.n55 outputibias.n54 9.3005
R21749 outputibias.n53 outputibias.n52 9.3005
R21750 outputibias.n38 outputibias.n37 9.3005
R21751 outputibias.n47 outputibias.n46 9.3005
R21752 outputibias.n45 outputibias.n44 9.3005
R21753 outputibias.n93 outputibias.n92 9.3005
R21754 outputibias.n66 outputibias.n65 9.3005
R21755 outputibias.n87 outputibias.n86 9.3005
R21756 outputibias.n85 outputibias.n84 9.3005
R21757 outputibias.n70 outputibias.n69 9.3005
R21758 outputibias.n79 outputibias.n78 9.3005
R21759 outputibias.n77 outputibias.n76 9.3005
R21760 outputibias.n125 outputibias.n124 9.3005
R21761 outputibias.n98 outputibias.n97 9.3005
R21762 outputibias.n119 outputibias.n118 9.3005
R21763 outputibias.n117 outputibias.n116 9.3005
R21764 outputibias.n102 outputibias.n101 9.3005
R21765 outputibias.n111 outputibias.n110 9.3005
R21766 outputibias.n109 outputibias.n108 9.3005
R21767 outputibias.n28 outputibias.n3 8.92171
R21768 outputibias.n59 outputibias.n34 8.92171
R21769 outputibias.n91 outputibias.n66 8.92171
R21770 outputibias.n123 outputibias.n98 8.92171
R21771 outputibias.n29 outputibias.n1 8.14595
R21772 outputibias.n60 outputibias.n32 8.14595
R21773 outputibias.n92 outputibias.n64 8.14595
R21774 outputibias.n124 outputibias.n96 8.14595
R21775 outputibias.n31 outputibias.n1 5.81868
R21776 outputibias.n62 outputibias.n32 5.81868
R21777 outputibias.n94 outputibias.n64 5.81868
R21778 outputibias.n126 outputibias.n96 5.81868
R21779 outputibias.n131 outputibias.n130 5.20947
R21780 outputibias.n29 outputibias.n28 5.04292
R21781 outputibias.n60 outputibias.n59 5.04292
R21782 outputibias.n92 outputibias.n91 5.04292
R21783 outputibias.n124 outputibias.n123 5.04292
R21784 outputibias.n131 outputibias.n127 4.42209
R21785 outputibias.n14 outputibias.n10 4.38594
R21786 outputibias.n45 outputibias.n41 4.38594
R21787 outputibias.n77 outputibias.n73 4.38594
R21788 outputibias.n109 outputibias.n105 4.38594
R21789 outputibias.n132 outputibias.n131 4.28454
R21790 outputibias.n25 outputibias.n3 4.26717
R21791 outputibias.n56 outputibias.n34 4.26717
R21792 outputibias.n88 outputibias.n66 4.26717
R21793 outputibias.n120 outputibias.n98 4.26717
R21794 outputibias.n24 outputibias.n5 3.49141
R21795 outputibias.n55 outputibias.n36 3.49141
R21796 outputibias.n87 outputibias.n68 3.49141
R21797 outputibias.n119 outputibias.n100 3.49141
R21798 outputibias.n21 outputibias.n20 2.71565
R21799 outputibias.n52 outputibias.n51 2.71565
R21800 outputibias.n84 outputibias.n83 2.71565
R21801 outputibias.n116 outputibias.n115 2.71565
R21802 outputibias.n17 outputibias.n7 1.93989
R21803 outputibias.n48 outputibias.n38 1.93989
R21804 outputibias.n80 outputibias.n70 1.93989
R21805 outputibias.n112 outputibias.n102 1.93989
R21806 outputibias.n130 outputibias.n129 1.9266
R21807 outputibias.n129 outputibias.n128 1.9266
R21808 outputibias.n133 outputibias.n132 1.92658
R21809 outputibias.n134 outputibias.n133 1.29913
R21810 outputibias.n16 outputibias.n9 1.16414
R21811 outputibias.n47 outputibias.n40 1.16414
R21812 outputibias.n79 outputibias.n72 1.16414
R21813 outputibias.n111 outputibias.n104 1.16414
R21814 outputibias.n127 outputibias.n95 0.962709
R21815 outputibias.n95 outputibias.n63 0.962709
R21816 outputibias.n13 outputibias.n12 0.388379
R21817 outputibias.n44 outputibias.n43 0.388379
R21818 outputibias.n76 outputibias.n75 0.388379
R21819 outputibias.n108 outputibias.n107 0.388379
R21820 outputibias.n134 outputibias.n0 0.337251
R21821 outputibias outputibias.n134 0.302375
R21822 outputibias.n30 outputibias.n2 0.155672
R21823 outputibias.n23 outputibias.n2 0.155672
R21824 outputibias.n23 outputibias.n22 0.155672
R21825 outputibias.n22 outputibias.n6 0.155672
R21826 outputibias.n15 outputibias.n6 0.155672
R21827 outputibias.n15 outputibias.n14 0.155672
R21828 outputibias.n61 outputibias.n33 0.155672
R21829 outputibias.n54 outputibias.n33 0.155672
R21830 outputibias.n54 outputibias.n53 0.155672
R21831 outputibias.n53 outputibias.n37 0.155672
R21832 outputibias.n46 outputibias.n37 0.155672
R21833 outputibias.n46 outputibias.n45 0.155672
R21834 outputibias.n93 outputibias.n65 0.155672
R21835 outputibias.n86 outputibias.n65 0.155672
R21836 outputibias.n86 outputibias.n85 0.155672
R21837 outputibias.n85 outputibias.n69 0.155672
R21838 outputibias.n78 outputibias.n69 0.155672
R21839 outputibias.n78 outputibias.n77 0.155672
R21840 outputibias.n125 outputibias.n97 0.155672
R21841 outputibias.n118 outputibias.n97 0.155672
R21842 outputibias.n118 outputibias.n117 0.155672
R21843 outputibias.n117 outputibias.n101 0.155672
R21844 outputibias.n110 outputibias.n101 0.155672
R21845 outputibias.n110 outputibias.n109 0.155672
R21846 output.n41 output.n15 289.615
R21847 output.n72 output.n46 289.615
R21848 output.n104 output.n78 289.615
R21849 output.n136 output.n110 289.615
R21850 output.n77 output.n45 197.26
R21851 output.n77 output.n76 196.298
R21852 output.n109 output.n108 196.298
R21853 output.n141 output.n140 196.298
R21854 output.n42 output.n41 185
R21855 output.n40 output.n39 185
R21856 output.n19 output.n18 185
R21857 output.n34 output.n33 185
R21858 output.n32 output.n31 185
R21859 output.n23 output.n22 185
R21860 output.n26 output.n25 185
R21861 output.n73 output.n72 185
R21862 output.n71 output.n70 185
R21863 output.n50 output.n49 185
R21864 output.n65 output.n64 185
R21865 output.n63 output.n62 185
R21866 output.n54 output.n53 185
R21867 output.n57 output.n56 185
R21868 output.n105 output.n104 185
R21869 output.n103 output.n102 185
R21870 output.n82 output.n81 185
R21871 output.n97 output.n96 185
R21872 output.n95 output.n94 185
R21873 output.n86 output.n85 185
R21874 output.n89 output.n88 185
R21875 output.n137 output.n136 185
R21876 output.n135 output.n134 185
R21877 output.n114 output.n113 185
R21878 output.n129 output.n128 185
R21879 output.n127 output.n126 185
R21880 output.n118 output.n117 185
R21881 output.n121 output.n120 185
R21882 output.t1 output.n24 147.661
R21883 output.t2 output.n55 147.661
R21884 output.t3 output.n87 147.661
R21885 output.t0 output.n119 147.661
R21886 output.n41 output.n40 104.615
R21887 output.n40 output.n18 104.615
R21888 output.n33 output.n18 104.615
R21889 output.n33 output.n32 104.615
R21890 output.n32 output.n22 104.615
R21891 output.n25 output.n22 104.615
R21892 output.n72 output.n71 104.615
R21893 output.n71 output.n49 104.615
R21894 output.n64 output.n49 104.615
R21895 output.n64 output.n63 104.615
R21896 output.n63 output.n53 104.615
R21897 output.n56 output.n53 104.615
R21898 output.n104 output.n103 104.615
R21899 output.n103 output.n81 104.615
R21900 output.n96 output.n81 104.615
R21901 output.n96 output.n95 104.615
R21902 output.n95 output.n85 104.615
R21903 output.n88 output.n85 104.615
R21904 output.n136 output.n135 104.615
R21905 output.n135 output.n113 104.615
R21906 output.n128 output.n113 104.615
R21907 output.n128 output.n127 104.615
R21908 output.n127 output.n117 104.615
R21909 output.n120 output.n117 104.615
R21910 output.n1 output.t5 77.056
R21911 output.n14 output.t6 76.6694
R21912 output.n1 output.n0 72.7095
R21913 output.n3 output.n2 72.7095
R21914 output.n5 output.n4 72.7095
R21915 output.n7 output.n6 72.7095
R21916 output.n9 output.n8 72.7095
R21917 output.n11 output.n10 72.7095
R21918 output.n13 output.n12 72.7095
R21919 output.n25 output.t1 52.3082
R21920 output.n56 output.t2 52.3082
R21921 output.n88 output.t3 52.3082
R21922 output.n120 output.t0 52.3082
R21923 output.n26 output.n24 15.6674
R21924 output.n57 output.n55 15.6674
R21925 output.n89 output.n87 15.6674
R21926 output.n121 output.n119 15.6674
R21927 output.n27 output.n23 12.8005
R21928 output.n58 output.n54 12.8005
R21929 output.n90 output.n86 12.8005
R21930 output.n122 output.n118 12.8005
R21931 output.n31 output.n30 12.0247
R21932 output.n62 output.n61 12.0247
R21933 output.n94 output.n93 12.0247
R21934 output.n126 output.n125 12.0247
R21935 output.n34 output.n21 11.249
R21936 output.n65 output.n52 11.249
R21937 output.n97 output.n84 11.249
R21938 output.n129 output.n116 11.249
R21939 output.n35 output.n19 10.4732
R21940 output.n66 output.n50 10.4732
R21941 output.n98 output.n82 10.4732
R21942 output.n130 output.n114 10.4732
R21943 output.n39 output.n38 9.69747
R21944 output.n70 output.n69 9.69747
R21945 output.n102 output.n101 9.69747
R21946 output.n134 output.n133 9.69747
R21947 output.n45 output.n44 9.45567
R21948 output.n76 output.n75 9.45567
R21949 output.n108 output.n107 9.45567
R21950 output.n140 output.n139 9.45567
R21951 output.n44 output.n43 9.3005
R21952 output.n17 output.n16 9.3005
R21953 output.n38 output.n37 9.3005
R21954 output.n36 output.n35 9.3005
R21955 output.n21 output.n20 9.3005
R21956 output.n30 output.n29 9.3005
R21957 output.n28 output.n27 9.3005
R21958 output.n75 output.n74 9.3005
R21959 output.n48 output.n47 9.3005
R21960 output.n69 output.n68 9.3005
R21961 output.n67 output.n66 9.3005
R21962 output.n52 output.n51 9.3005
R21963 output.n61 output.n60 9.3005
R21964 output.n59 output.n58 9.3005
R21965 output.n107 output.n106 9.3005
R21966 output.n80 output.n79 9.3005
R21967 output.n101 output.n100 9.3005
R21968 output.n99 output.n98 9.3005
R21969 output.n84 output.n83 9.3005
R21970 output.n93 output.n92 9.3005
R21971 output.n91 output.n90 9.3005
R21972 output.n139 output.n138 9.3005
R21973 output.n112 output.n111 9.3005
R21974 output.n133 output.n132 9.3005
R21975 output.n131 output.n130 9.3005
R21976 output.n116 output.n115 9.3005
R21977 output.n125 output.n124 9.3005
R21978 output.n123 output.n122 9.3005
R21979 output.n42 output.n17 8.92171
R21980 output.n73 output.n48 8.92171
R21981 output.n105 output.n80 8.92171
R21982 output.n137 output.n112 8.92171
R21983 output output.n141 8.15037
R21984 output.n43 output.n15 8.14595
R21985 output.n74 output.n46 8.14595
R21986 output.n106 output.n78 8.14595
R21987 output.n138 output.n110 8.14595
R21988 output.n45 output.n15 5.81868
R21989 output.n76 output.n46 5.81868
R21990 output.n108 output.n78 5.81868
R21991 output.n140 output.n110 5.81868
R21992 output.n43 output.n42 5.04292
R21993 output.n74 output.n73 5.04292
R21994 output.n106 output.n105 5.04292
R21995 output.n138 output.n137 5.04292
R21996 output.n28 output.n24 4.38594
R21997 output.n59 output.n55 4.38594
R21998 output.n91 output.n87 4.38594
R21999 output.n123 output.n119 4.38594
R22000 output.n39 output.n17 4.26717
R22001 output.n70 output.n48 4.26717
R22002 output.n102 output.n80 4.26717
R22003 output.n134 output.n112 4.26717
R22004 output.n0 output.t16 3.9605
R22005 output.n0 output.t19 3.9605
R22006 output.n2 output.t9 3.9605
R22007 output.n2 output.t8 3.9605
R22008 output.n4 output.t14 3.9605
R22009 output.n4 output.t18 3.9605
R22010 output.n6 output.t7 3.9605
R22011 output.n6 output.t10 3.9605
R22012 output.n8 output.t11 3.9605
R22013 output.n8 output.t17 3.9605
R22014 output.n10 output.t4 3.9605
R22015 output.n10 output.t12 3.9605
R22016 output.n12 output.t15 3.9605
R22017 output.n12 output.t13 3.9605
R22018 output.n38 output.n19 3.49141
R22019 output.n69 output.n50 3.49141
R22020 output.n101 output.n82 3.49141
R22021 output.n133 output.n114 3.49141
R22022 output.n35 output.n34 2.71565
R22023 output.n66 output.n65 2.71565
R22024 output.n98 output.n97 2.71565
R22025 output.n130 output.n129 2.71565
R22026 output.n31 output.n21 1.93989
R22027 output.n62 output.n52 1.93989
R22028 output.n94 output.n84 1.93989
R22029 output.n126 output.n116 1.93989
R22030 output.n30 output.n23 1.16414
R22031 output.n61 output.n54 1.16414
R22032 output.n93 output.n86 1.16414
R22033 output.n125 output.n118 1.16414
R22034 output.n141 output.n109 0.962709
R22035 output.n109 output.n77 0.962709
R22036 output.n27 output.n26 0.388379
R22037 output.n58 output.n57 0.388379
R22038 output.n90 output.n89 0.388379
R22039 output.n122 output.n121 0.388379
R22040 output.n14 output.n13 0.387128
R22041 output.n13 output.n11 0.387128
R22042 output.n11 output.n9 0.387128
R22043 output.n9 output.n7 0.387128
R22044 output.n7 output.n5 0.387128
R22045 output.n5 output.n3 0.387128
R22046 output.n3 output.n1 0.387128
R22047 output.n44 output.n16 0.155672
R22048 output.n37 output.n16 0.155672
R22049 output.n37 output.n36 0.155672
R22050 output.n36 output.n20 0.155672
R22051 output.n29 output.n20 0.155672
R22052 output.n29 output.n28 0.155672
R22053 output.n75 output.n47 0.155672
R22054 output.n68 output.n47 0.155672
R22055 output.n68 output.n67 0.155672
R22056 output.n67 output.n51 0.155672
R22057 output.n60 output.n51 0.155672
R22058 output.n60 output.n59 0.155672
R22059 output.n107 output.n79 0.155672
R22060 output.n100 output.n79 0.155672
R22061 output.n100 output.n99 0.155672
R22062 output.n99 output.n83 0.155672
R22063 output.n92 output.n83 0.155672
R22064 output.n92 output.n91 0.155672
R22065 output.n139 output.n111 0.155672
R22066 output.n132 output.n111 0.155672
R22067 output.n132 output.n131 0.155672
R22068 output.n131 output.n115 0.155672
R22069 output.n124 output.n115 0.155672
R22070 output.n124 output.n123 0.155672
R22071 output output.n14 0.126227
R22072 minus.n76 minus.t28 250.337
R22073 minus.n15 minus.t20 250.337
R22074 minus.n126 minus.t1 243.255
R22075 minus.n120 minus.t8 231.093
R22076 minus.n59 minus.t10 231.093
R22077 minus.n125 minus.n123 224.169
R22078 minus.n125 minus.n124 223.454
R22079 minus.n62 minus.t12 187.445
R22080 minus.n113 minus.t18 187.445
R22081 minus.n107 minus.t25 187.445
R22082 minus.n66 minus.t22 187.445
R22083 minus.n68 minus.t19 187.445
R22084 minus.n95 minus.t7 187.445
R22085 minus.n89 minus.t6 187.445
R22086 minus.n72 minus.t16 187.445
R22087 minus.n74 minus.t15 187.445
R22088 minus.n77 minus.t23 187.445
R22089 minus.n16 minus.t14 187.445
R22090 minus.n13 minus.t9 187.445
R22091 minus.n11 minus.t5 187.445
R22092 minus.n28 minus.t26 187.445
R22093 minus.n34 minus.t27 187.445
R22094 minus.n7 minus.t21 187.445
R22095 minus.n5 minus.t24 187.445
R22096 minus.n46 minus.t17 187.445
R22097 minus.n52 minus.t11 187.445
R22098 minus.n1 minus.t13 187.445
R22099 minus.n78 minus.n75 161.3
R22100 minus.n80 minus.n79 161.3
R22101 minus.n82 minus.n81 161.3
R22102 minus.n83 minus.n73 161.3
R22103 minus.n85 minus.n84 161.3
R22104 minus.n87 minus.n86 161.3
R22105 minus.n88 minus.n71 161.3
R22106 minus.n91 minus.n90 161.3
R22107 minus.n92 minus.n70 161.3
R22108 minus.n94 minus.n93 161.3
R22109 minus.n96 minus.n69 161.3
R22110 minus.n98 minus.n97 161.3
R22111 minus.n100 minus.n99 161.3
R22112 minus.n101 minus.n67 161.3
R22113 minus.n103 minus.n102 161.3
R22114 minus.n105 minus.n104 161.3
R22115 minus.n106 minus.n65 161.3
R22116 minus.n109 minus.n108 161.3
R22117 minus.n110 minus.n64 161.3
R22118 minus.n112 minus.n111 161.3
R22119 minus.n114 minus.n63 161.3
R22120 minus.n116 minus.n115 161.3
R22121 minus.n118 minus.n117 161.3
R22122 minus.n119 minus.n61 161.3
R22123 minus.n121 minus.n120 161.3
R22124 minus.n60 minus.n59 161.3
R22125 minus.n58 minus.n0 161.3
R22126 minus.n57 minus.n56 161.3
R22127 minus.n55 minus.n54 161.3
R22128 minus.n53 minus.n2 161.3
R22129 minus.n51 minus.n50 161.3
R22130 minus.n49 minus.n3 161.3
R22131 minus.n48 minus.n47 161.3
R22132 minus.n45 minus.n4 161.3
R22133 minus.n44 minus.n43 161.3
R22134 minus.n42 minus.n41 161.3
R22135 minus.n40 minus.n6 161.3
R22136 minus.n39 minus.n38 161.3
R22137 minus.n37 minus.n36 161.3
R22138 minus.n35 minus.n8 161.3
R22139 minus.n33 minus.n32 161.3
R22140 minus.n31 minus.n9 161.3
R22141 minus.n30 minus.n29 161.3
R22142 minus.n27 minus.n10 161.3
R22143 minus.n26 minus.n25 161.3
R22144 minus.n24 minus.n23 161.3
R22145 minus.n22 minus.n12 161.3
R22146 minus.n21 minus.n20 161.3
R22147 minus.n19 minus.n18 161.3
R22148 minus.n17 minus.n14 161.3
R22149 minus.n106 minus.n105 56.5617
R22150 minus.n97 minus.n96 56.5617
R22151 minus.n88 minus.n87 56.5617
R22152 minus.n27 minus.n26 56.5617
R22153 minus.n36 minus.n35 56.5617
R22154 minus.n45 minus.n44 56.5617
R22155 minus.n115 minus.n114 56.5617
R22156 minus.n79 minus.n78 56.5617
R22157 minus.n18 minus.n17 56.5617
R22158 minus.n54 minus.n53 56.5617
R22159 minus.n119 minus.n118 50.2647
R22160 minus.n58 minus.n57 50.2647
R22161 minus.n108 minus.n64 46.3896
R22162 minus.n84 minus.n83 46.3896
R22163 minus.n23 minus.n22 46.3896
R22164 minus.n47 minus.n3 46.3896
R22165 minus.n76 minus.n75 43.1929
R22166 minus.n15 minus.n14 43.1929
R22167 minus.n101 minus.n100 42.5146
R22168 minus.n94 minus.n70 42.5146
R22169 minus.n33 minus.n9 42.5146
R22170 minus.n40 minus.n39 42.5146
R22171 minus.n77 minus.n76 40.6041
R22172 minus.n16 minus.n15 40.6041
R22173 minus.n102 minus.n101 38.6395
R22174 minus.n90 minus.n70 38.6395
R22175 minus.n29 minus.n9 38.6395
R22176 minus.n41 minus.n40 38.6395
R22177 minus.n122 minus.n121 35.4191
R22178 minus.n112 minus.n64 34.7644
R22179 minus.n83 minus.n82 34.7644
R22180 minus.n22 minus.n21 34.7644
R22181 minus.n51 minus.n3 34.7644
R22182 minus.n114 minus.n113 21.8872
R22183 minus.n79 minus.n74 21.8872
R22184 minus.n18 minus.n13 21.8872
R22185 minus.n53 minus.n52 21.8872
R22186 minus.n105 minus.n66 19.9199
R22187 minus.n89 minus.n88 19.9199
R22188 minus.n28 minus.n27 19.9199
R22189 minus.n44 minus.n5 19.9199
R22190 minus.n124 minus.t0 19.8005
R22191 minus.n124 minus.t2 19.8005
R22192 minus.n123 minus.t4 19.8005
R22193 minus.n123 minus.t3 19.8005
R22194 minus.n97 minus.n68 17.9525
R22195 minus.n96 minus.n95 17.9525
R22196 minus.n35 minus.n34 17.9525
R22197 minus.n36 minus.n7 17.9525
R22198 minus.n107 minus.n106 15.9852
R22199 minus.n87 minus.n72 15.9852
R22200 minus.n26 minus.n11 15.9852
R22201 minus.n46 minus.n45 15.9852
R22202 minus.n115 minus.n62 14.0178
R22203 minus.n78 minus.n77 14.0178
R22204 minus.n17 minus.n16 14.0178
R22205 minus.n54 minus.n1 14.0178
R22206 minus.n122 minus.n60 12.1501
R22207 minus minus.n127 11.2056
R22208 minus.n118 minus.n62 10.575
R22209 minus.n57 minus.n1 10.575
R22210 minus.n120 minus.n119 9.49444
R22211 minus.n59 minus.n58 9.49444
R22212 minus.n108 minus.n107 8.60764
R22213 minus.n84 minus.n72 8.60764
R22214 minus.n23 minus.n11 8.60764
R22215 minus.n47 minus.n46 8.60764
R22216 minus.n100 minus.n68 6.6403
R22217 minus.n95 minus.n94 6.6403
R22218 minus.n34 minus.n33 6.6403
R22219 minus.n39 minus.n7 6.6403
R22220 minus.n127 minus.n126 4.80222
R22221 minus.n102 minus.n66 4.67295
R22222 minus.n90 minus.n89 4.67295
R22223 minus.n29 minus.n28 4.67295
R22224 minus.n41 minus.n5 4.67295
R22225 minus.n113 minus.n112 2.7056
R22226 minus.n82 minus.n74 2.7056
R22227 minus.n21 minus.n13 2.7056
R22228 minus.n52 minus.n51 2.7056
R22229 minus.n127 minus.n122 0.972091
R22230 minus.n126 minus.n125 0.716017
R22231 minus.n121 minus.n61 0.189894
R22232 minus.n117 minus.n61 0.189894
R22233 minus.n117 minus.n116 0.189894
R22234 minus.n116 minus.n63 0.189894
R22235 minus.n111 minus.n63 0.189894
R22236 minus.n111 minus.n110 0.189894
R22237 minus.n110 minus.n109 0.189894
R22238 minus.n109 minus.n65 0.189894
R22239 minus.n104 minus.n65 0.189894
R22240 minus.n104 minus.n103 0.189894
R22241 minus.n103 minus.n67 0.189894
R22242 minus.n99 minus.n67 0.189894
R22243 minus.n99 minus.n98 0.189894
R22244 minus.n98 minus.n69 0.189894
R22245 minus.n93 minus.n69 0.189894
R22246 minus.n93 minus.n92 0.189894
R22247 minus.n92 minus.n91 0.189894
R22248 minus.n91 minus.n71 0.189894
R22249 minus.n86 minus.n71 0.189894
R22250 minus.n86 minus.n85 0.189894
R22251 minus.n85 minus.n73 0.189894
R22252 minus.n81 minus.n73 0.189894
R22253 minus.n81 minus.n80 0.189894
R22254 minus.n80 minus.n75 0.189894
R22255 minus.n19 minus.n14 0.189894
R22256 minus.n20 minus.n19 0.189894
R22257 minus.n20 minus.n12 0.189894
R22258 minus.n24 minus.n12 0.189894
R22259 minus.n25 minus.n24 0.189894
R22260 minus.n25 minus.n10 0.189894
R22261 minus.n30 minus.n10 0.189894
R22262 minus.n31 minus.n30 0.189894
R22263 minus.n32 minus.n31 0.189894
R22264 minus.n32 minus.n8 0.189894
R22265 minus.n37 minus.n8 0.189894
R22266 minus.n38 minus.n37 0.189894
R22267 minus.n38 minus.n6 0.189894
R22268 minus.n42 minus.n6 0.189894
R22269 minus.n43 minus.n42 0.189894
R22270 minus.n43 minus.n4 0.189894
R22271 minus.n48 minus.n4 0.189894
R22272 minus.n49 minus.n48 0.189894
R22273 minus.n50 minus.n49 0.189894
R22274 minus.n50 minus.n2 0.189894
R22275 minus.n55 minus.n2 0.189894
R22276 minus.n56 minus.n55 0.189894
R22277 minus.n56 minus.n0 0.189894
R22278 minus.n60 minus.n0 0.189894
C0 minus commonsourceibias 0.343793f
C1 plus commonsourceibias 0.290384f
C2 output outputibias 2.34152f
C3 vdd output 7.23429f
C4 CSoutput output 6.13881f
C5 CSoutput outputibias 0.032386f
C6 vdd CSoutput 91.9904f
C7 minus diffpairibias 5.39e-19
C8 commonsourceibias output 0.006808f
C9 vdd plus 0.080622f
C10 CSoutput minus 2.49197f
C11 plus diffpairibias 4.4e-19
C12 commonsourceibias outputibias 0.003832f
C13 vdd commonsourceibias 0.004218f
C14 CSoutput plus 0.892246f
C15 commonsourceibias diffpairibias 0.064336f
C16 minus plus 10.004901f
C17 CSoutput commonsourceibias 42.3358f
C18 diffpairibias gnd 60.003128f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.145005p
C22 plus gnd 38.5963f
C23 minus gnd 30.044651f
C24 CSoutput gnd 0.10808p
C25 vdd gnd 0.376447p
C26 minus.n0 gnd 0.031282f
C27 minus.t13 gnd 0.525996f
C28 minus.n1 gnd 0.212736f
C29 minus.n2 gnd 0.031282f
C30 minus.t11 gnd 0.525996f
C31 minus.n3 gnd 0.026731f
C32 minus.n4 gnd 0.031282f
C33 minus.t17 gnd 0.525996f
C34 minus.t24 gnd 0.525996f
C35 minus.n5 gnd 0.212736f
C36 minus.n6 gnd 0.031282f
C37 minus.t21 gnd 0.525996f
C38 minus.n7 gnd 0.212736f
C39 minus.n8 gnd 0.031282f
C40 minus.t27 gnd 0.525996f
C41 minus.n9 gnd 0.025425f
C42 minus.n10 gnd 0.031282f
C43 minus.t26 gnd 0.525996f
C44 minus.t5 gnd 0.525996f
C45 minus.n11 gnd 0.212736f
C46 minus.n12 gnd 0.031282f
C47 minus.t9 gnd 0.525996f
C48 minus.n13 gnd 0.212736f
C49 minus.n14 gnd 0.132756f
C50 minus.t14 gnd 0.525996f
C51 minus.t20 gnd 0.588422f
C52 minus.n15 gnd 0.24871f
C53 minus.n16 gnd 0.243623f
C54 minus.n17 gnd 0.040082f
C55 minus.n18 gnd 0.035399f
C56 minus.n19 gnd 0.031282f
C57 minus.n20 gnd 0.031282f
C58 minus.n21 gnd 0.037382f
C59 minus.n22 gnd 0.026731f
C60 minus.n23 gnd 0.04074f
C61 minus.n24 gnd 0.031282f
C62 minus.n25 gnd 0.031282f
C63 minus.n26 gnd 0.038912f
C64 minus.n27 gnd 0.03657f
C65 minus.n28 gnd 0.212736f
C66 minus.n29 gnd 0.039185f
C67 minus.n30 gnd 0.031282f
C68 minus.n31 gnd 0.031282f
C69 minus.n32 gnd 0.031282f
C70 minus.n33 gnd 0.040243f
C71 minus.n34 gnd 0.212736f
C72 minus.n35 gnd 0.037741f
C73 minus.n36 gnd 0.037741f
C74 minus.n37 gnd 0.031282f
C75 minus.n38 gnd 0.031282f
C76 minus.n39 gnd 0.040243f
C77 minus.n40 gnd 0.025425f
C78 minus.n41 gnd 0.039185f
C79 minus.n42 gnd 0.031282f
C80 minus.n43 gnd 0.031282f
C81 minus.n44 gnd 0.03657f
C82 minus.n45 gnd 0.038912f
C83 minus.n46 gnd 0.212736f
C84 minus.n47 gnd 0.04074f
C85 minus.n48 gnd 0.031282f
C86 minus.n49 gnd 0.031282f
C87 minus.n50 gnd 0.031282f
C88 minus.n51 gnd 0.037382f
C89 minus.n52 gnd 0.212736f
C90 minus.n53 gnd 0.035399f
C91 minus.n54 gnd 0.040082f
C92 minus.n55 gnd 0.031282f
C93 minus.n56 gnd 0.031282f
C94 minus.n57 gnd 0.040808f
C95 minus.n58 gnd 0.011369f
C96 minus.t10 gnd 0.568865f
C97 minus.n59 gnd 0.246313f
C98 minus.n60 gnd 0.366453f
C99 minus.n61 gnd 0.031282f
C100 minus.t8 gnd 0.568865f
C101 minus.t12 gnd 0.525996f
C102 minus.n62 gnd 0.212736f
C103 minus.n63 gnd 0.031282f
C104 minus.t18 gnd 0.525996f
C105 minus.n64 gnd 0.026731f
C106 minus.n65 gnd 0.031282f
C107 minus.t25 gnd 0.525996f
C108 minus.t22 gnd 0.525996f
C109 minus.n66 gnd 0.212736f
C110 minus.n67 gnd 0.031282f
C111 minus.t19 gnd 0.525996f
C112 minus.n68 gnd 0.212736f
C113 minus.n69 gnd 0.031282f
C114 minus.t7 gnd 0.525996f
C115 minus.n70 gnd 0.025425f
C116 minus.n71 gnd 0.031282f
C117 minus.t6 gnd 0.525996f
C118 minus.t16 gnd 0.525996f
C119 minus.n72 gnd 0.212736f
C120 minus.n73 gnd 0.031282f
C121 minus.t15 gnd 0.525996f
C122 minus.n74 gnd 0.212736f
C123 minus.n75 gnd 0.132756f
C124 minus.t23 gnd 0.525996f
C125 minus.t28 gnd 0.588422f
C126 minus.n76 gnd 0.24871f
C127 minus.n77 gnd 0.243623f
C128 minus.n78 gnd 0.040082f
C129 minus.n79 gnd 0.035399f
C130 minus.n80 gnd 0.031282f
C131 minus.n81 gnd 0.031282f
C132 minus.n82 gnd 0.037382f
C133 minus.n83 gnd 0.026731f
C134 minus.n84 gnd 0.04074f
C135 minus.n85 gnd 0.031282f
C136 minus.n86 gnd 0.031282f
C137 minus.n87 gnd 0.038912f
C138 minus.n88 gnd 0.03657f
C139 minus.n89 gnd 0.212736f
C140 minus.n90 gnd 0.039185f
C141 minus.n91 gnd 0.031282f
C142 minus.n92 gnd 0.031282f
C143 minus.n93 gnd 0.031282f
C144 minus.n94 gnd 0.040243f
C145 minus.n95 gnd 0.212736f
C146 minus.n96 gnd 0.037741f
C147 minus.n97 gnd 0.037741f
C148 minus.n98 gnd 0.031282f
C149 minus.n99 gnd 0.031282f
C150 minus.n100 gnd 0.040243f
C151 minus.n101 gnd 0.025425f
C152 minus.n102 gnd 0.039185f
C153 minus.n103 gnd 0.031282f
C154 minus.n104 gnd 0.031282f
C155 minus.n105 gnd 0.03657f
C156 minus.n106 gnd 0.038912f
C157 minus.n107 gnd 0.212736f
C158 minus.n108 gnd 0.04074f
C159 minus.n109 gnd 0.031282f
C160 minus.n110 gnd 0.031282f
C161 minus.n111 gnd 0.031282f
C162 minus.n112 gnd 0.037382f
C163 minus.n113 gnd 0.212736f
C164 minus.n114 gnd 0.035399f
C165 minus.n115 gnd 0.040082f
C166 minus.n116 gnd 0.031282f
C167 minus.n117 gnd 0.031282f
C168 minus.n118 gnd 0.040808f
C169 minus.n119 gnd 0.011369f
C170 minus.n120 gnd 0.246313f
C171 minus.n121 gnd 1.14114f
C172 minus.n122 gnd 1.67625f
C173 minus.t4 gnd 0.009643f
C174 minus.t3 gnd 0.009643f
C175 minus.n123 gnd 0.031709f
C176 minus.t0 gnd 0.009643f
C177 minus.t2 gnd 0.009643f
C178 minus.n124 gnd 0.031275f
C179 minus.n125 gnd 0.266915f
C180 minus.t1 gnd 0.053673f
C181 minus.n126 gnd 0.145653f
C182 minus.n127 gnd 1.75318f
C183 output.t5 gnd 0.464308f
C184 output.t16 gnd 0.044422f
C185 output.t19 gnd 0.044422f
C186 output.n0 gnd 0.364624f
C187 output.n1 gnd 0.614102f
C188 output.t9 gnd 0.044422f
C189 output.t8 gnd 0.044422f
C190 output.n2 gnd 0.364624f
C191 output.n3 gnd 0.350265f
C192 output.t14 gnd 0.044422f
C193 output.t18 gnd 0.044422f
C194 output.n4 gnd 0.364624f
C195 output.n5 gnd 0.350265f
C196 output.t7 gnd 0.044422f
C197 output.t10 gnd 0.044422f
C198 output.n6 gnd 0.364624f
C199 output.n7 gnd 0.350265f
C200 output.t11 gnd 0.044422f
C201 output.t17 gnd 0.044422f
C202 output.n8 gnd 0.364624f
C203 output.n9 gnd 0.350265f
C204 output.t4 gnd 0.044422f
C205 output.t12 gnd 0.044422f
C206 output.n10 gnd 0.364624f
C207 output.n11 gnd 0.350265f
C208 output.t15 gnd 0.044422f
C209 output.t13 gnd 0.044422f
C210 output.n12 gnd 0.364624f
C211 output.n13 gnd 0.350265f
C212 output.t6 gnd 0.462979f
C213 output.n14 gnd 0.28994f
C214 output.n15 gnd 0.015803f
C215 output.n16 gnd 0.011243f
C216 output.n17 gnd 0.006041f
C217 output.n18 gnd 0.01428f
C218 output.n19 gnd 0.006397f
C219 output.n20 gnd 0.011243f
C220 output.n21 gnd 0.006041f
C221 output.n22 gnd 0.01428f
C222 output.n23 gnd 0.006397f
C223 output.n24 gnd 0.048111f
C224 output.t1 gnd 0.023274f
C225 output.n25 gnd 0.01071f
C226 output.n26 gnd 0.008435f
C227 output.n27 gnd 0.006041f
C228 output.n28 gnd 0.267512f
C229 output.n29 gnd 0.011243f
C230 output.n30 gnd 0.006041f
C231 output.n31 gnd 0.006397f
C232 output.n32 gnd 0.01428f
C233 output.n33 gnd 0.01428f
C234 output.n34 gnd 0.006397f
C235 output.n35 gnd 0.006041f
C236 output.n36 gnd 0.011243f
C237 output.n37 gnd 0.011243f
C238 output.n38 gnd 0.006041f
C239 output.n39 gnd 0.006397f
C240 output.n40 gnd 0.01428f
C241 output.n41 gnd 0.030913f
C242 output.n42 gnd 0.006397f
C243 output.n43 gnd 0.006041f
C244 output.n44 gnd 0.025987f
C245 output.n45 gnd 0.097665f
C246 output.n46 gnd 0.015803f
C247 output.n47 gnd 0.011243f
C248 output.n48 gnd 0.006041f
C249 output.n49 gnd 0.01428f
C250 output.n50 gnd 0.006397f
C251 output.n51 gnd 0.011243f
C252 output.n52 gnd 0.006041f
C253 output.n53 gnd 0.01428f
C254 output.n54 gnd 0.006397f
C255 output.n55 gnd 0.048111f
C256 output.t2 gnd 0.023274f
C257 output.n56 gnd 0.01071f
C258 output.n57 gnd 0.008435f
C259 output.n58 gnd 0.006041f
C260 output.n59 gnd 0.267512f
C261 output.n60 gnd 0.011243f
C262 output.n61 gnd 0.006041f
C263 output.n62 gnd 0.006397f
C264 output.n63 gnd 0.01428f
C265 output.n64 gnd 0.01428f
C266 output.n65 gnd 0.006397f
C267 output.n66 gnd 0.006041f
C268 output.n67 gnd 0.011243f
C269 output.n68 gnd 0.011243f
C270 output.n69 gnd 0.006041f
C271 output.n70 gnd 0.006397f
C272 output.n71 gnd 0.01428f
C273 output.n72 gnd 0.030913f
C274 output.n73 gnd 0.006397f
C275 output.n74 gnd 0.006041f
C276 output.n75 gnd 0.025987f
C277 output.n76 gnd 0.09306f
C278 output.n77 gnd 1.65264f
C279 output.n78 gnd 0.015803f
C280 output.n79 gnd 0.011243f
C281 output.n80 gnd 0.006041f
C282 output.n81 gnd 0.01428f
C283 output.n82 gnd 0.006397f
C284 output.n83 gnd 0.011243f
C285 output.n84 gnd 0.006041f
C286 output.n85 gnd 0.01428f
C287 output.n86 gnd 0.006397f
C288 output.n87 gnd 0.048111f
C289 output.t3 gnd 0.023274f
C290 output.n88 gnd 0.01071f
C291 output.n89 gnd 0.008435f
C292 output.n90 gnd 0.006041f
C293 output.n91 gnd 0.267512f
C294 output.n92 gnd 0.011243f
C295 output.n93 gnd 0.006041f
C296 output.n94 gnd 0.006397f
C297 output.n95 gnd 0.01428f
C298 output.n96 gnd 0.01428f
C299 output.n97 gnd 0.006397f
C300 output.n98 gnd 0.006041f
C301 output.n99 gnd 0.011243f
C302 output.n100 gnd 0.011243f
C303 output.n101 gnd 0.006041f
C304 output.n102 gnd 0.006397f
C305 output.n103 gnd 0.01428f
C306 output.n104 gnd 0.030913f
C307 output.n105 gnd 0.006397f
C308 output.n106 gnd 0.006041f
C309 output.n107 gnd 0.025987f
C310 output.n108 gnd 0.09306f
C311 output.n109 gnd 0.713089f
C312 output.n110 gnd 0.015803f
C313 output.n111 gnd 0.011243f
C314 output.n112 gnd 0.006041f
C315 output.n113 gnd 0.01428f
C316 output.n114 gnd 0.006397f
C317 output.n115 gnd 0.011243f
C318 output.n116 gnd 0.006041f
C319 output.n117 gnd 0.01428f
C320 output.n118 gnd 0.006397f
C321 output.n119 gnd 0.048111f
C322 output.t0 gnd 0.023274f
C323 output.n120 gnd 0.01071f
C324 output.n121 gnd 0.008435f
C325 output.n122 gnd 0.006041f
C326 output.n123 gnd 0.267512f
C327 output.n124 gnd 0.011243f
C328 output.n125 gnd 0.006041f
C329 output.n126 gnd 0.006397f
C330 output.n127 gnd 0.01428f
C331 output.n128 gnd 0.01428f
C332 output.n129 gnd 0.006397f
C333 output.n130 gnd 0.006041f
C334 output.n131 gnd 0.011243f
C335 output.n132 gnd 0.011243f
C336 output.n133 gnd 0.006041f
C337 output.n134 gnd 0.006397f
C338 output.n135 gnd 0.01428f
C339 output.n136 gnd 0.030913f
C340 output.n137 gnd 0.006397f
C341 output.n138 gnd 0.006041f
C342 output.n139 gnd 0.025987f
C343 output.n140 gnd 0.09306f
C344 output.n141 gnd 1.67353f
C345 outputibias.t9 gnd 0.11477f
C346 outputibias.t10 gnd 0.115567f
C347 outputibias.n0 gnd 0.130108f
C348 outputibias.n1 gnd 0.001372f
C349 outputibias.n2 gnd 9.76e-19
C350 outputibias.n3 gnd 5.24e-19
C351 outputibias.n4 gnd 0.001239f
C352 outputibias.n5 gnd 5.55e-19
C353 outputibias.n6 gnd 9.76e-19
C354 outputibias.n7 gnd 5.24e-19
C355 outputibias.n8 gnd 0.001239f
C356 outputibias.n9 gnd 5.55e-19
C357 outputibias.n10 gnd 0.004176f
C358 outputibias.t7 gnd 0.00202f
C359 outputibias.n11 gnd 9.3e-19
C360 outputibias.n12 gnd 7.32e-19
C361 outputibias.n13 gnd 5.24e-19
C362 outputibias.n14 gnd 0.02322f
C363 outputibias.n15 gnd 9.76e-19
C364 outputibias.n16 gnd 5.24e-19
C365 outputibias.n17 gnd 5.55e-19
C366 outputibias.n18 gnd 0.001239f
C367 outputibias.n19 gnd 0.001239f
C368 outputibias.n20 gnd 5.55e-19
C369 outputibias.n21 gnd 5.24e-19
C370 outputibias.n22 gnd 9.76e-19
C371 outputibias.n23 gnd 9.76e-19
C372 outputibias.n24 gnd 5.24e-19
C373 outputibias.n25 gnd 5.55e-19
C374 outputibias.n26 gnd 0.001239f
C375 outputibias.n27 gnd 0.002683f
C376 outputibias.n28 gnd 5.55e-19
C377 outputibias.n29 gnd 5.24e-19
C378 outputibias.n30 gnd 0.002256f
C379 outputibias.n31 gnd 0.005781f
C380 outputibias.n32 gnd 0.001372f
C381 outputibias.n33 gnd 9.76e-19
C382 outputibias.n34 gnd 5.24e-19
C383 outputibias.n35 gnd 0.001239f
C384 outputibias.n36 gnd 5.55e-19
C385 outputibias.n37 gnd 9.76e-19
C386 outputibias.n38 gnd 5.24e-19
C387 outputibias.n39 gnd 0.001239f
C388 outputibias.n40 gnd 5.55e-19
C389 outputibias.n41 gnd 0.004176f
C390 outputibias.t1 gnd 0.00202f
C391 outputibias.n42 gnd 9.3e-19
C392 outputibias.n43 gnd 7.32e-19
C393 outputibias.n44 gnd 5.24e-19
C394 outputibias.n45 gnd 0.02322f
C395 outputibias.n46 gnd 9.76e-19
C396 outputibias.n47 gnd 5.24e-19
C397 outputibias.n48 gnd 5.55e-19
C398 outputibias.n49 gnd 0.001239f
C399 outputibias.n50 gnd 0.001239f
C400 outputibias.n51 gnd 5.55e-19
C401 outputibias.n52 gnd 5.24e-19
C402 outputibias.n53 gnd 9.76e-19
C403 outputibias.n54 gnd 9.76e-19
C404 outputibias.n55 gnd 5.24e-19
C405 outputibias.n56 gnd 5.55e-19
C406 outputibias.n57 gnd 0.001239f
C407 outputibias.n58 gnd 0.002683f
C408 outputibias.n59 gnd 5.55e-19
C409 outputibias.n60 gnd 5.24e-19
C410 outputibias.n61 gnd 0.002256f
C411 outputibias.n62 gnd 0.005197f
C412 outputibias.n63 gnd 0.121892f
C413 outputibias.n64 gnd 0.001372f
C414 outputibias.n65 gnd 9.76e-19
C415 outputibias.n66 gnd 5.24e-19
C416 outputibias.n67 gnd 0.001239f
C417 outputibias.n68 gnd 5.55e-19
C418 outputibias.n69 gnd 9.76e-19
C419 outputibias.n70 gnd 5.24e-19
C420 outputibias.n71 gnd 0.001239f
C421 outputibias.n72 gnd 5.55e-19
C422 outputibias.n73 gnd 0.004176f
C423 outputibias.t3 gnd 0.00202f
C424 outputibias.n74 gnd 9.3e-19
C425 outputibias.n75 gnd 7.32e-19
C426 outputibias.n76 gnd 5.24e-19
C427 outputibias.n77 gnd 0.02322f
C428 outputibias.n78 gnd 9.76e-19
C429 outputibias.n79 gnd 5.24e-19
C430 outputibias.n80 gnd 5.55e-19
C431 outputibias.n81 gnd 0.001239f
C432 outputibias.n82 gnd 0.001239f
C433 outputibias.n83 gnd 5.55e-19
C434 outputibias.n84 gnd 5.24e-19
C435 outputibias.n85 gnd 9.76e-19
C436 outputibias.n86 gnd 9.76e-19
C437 outputibias.n87 gnd 5.24e-19
C438 outputibias.n88 gnd 5.55e-19
C439 outputibias.n89 gnd 0.001239f
C440 outputibias.n90 gnd 0.002683f
C441 outputibias.n91 gnd 5.55e-19
C442 outputibias.n92 gnd 5.24e-19
C443 outputibias.n93 gnd 0.002256f
C444 outputibias.n94 gnd 0.005197f
C445 outputibias.n95 gnd 0.064513f
C446 outputibias.n96 gnd 0.001372f
C447 outputibias.n97 gnd 9.76e-19
C448 outputibias.n98 gnd 5.24e-19
C449 outputibias.n99 gnd 0.001239f
C450 outputibias.n100 gnd 5.55e-19
C451 outputibias.n101 gnd 9.76e-19
C452 outputibias.n102 gnd 5.24e-19
C453 outputibias.n103 gnd 0.001239f
C454 outputibias.n104 gnd 5.55e-19
C455 outputibias.n105 gnd 0.004176f
C456 outputibias.t5 gnd 0.00202f
C457 outputibias.n106 gnd 9.3e-19
C458 outputibias.n107 gnd 7.32e-19
C459 outputibias.n108 gnd 5.24e-19
C460 outputibias.n109 gnd 0.02322f
C461 outputibias.n110 gnd 9.76e-19
C462 outputibias.n111 gnd 5.24e-19
C463 outputibias.n112 gnd 5.55e-19
C464 outputibias.n113 gnd 0.001239f
C465 outputibias.n114 gnd 0.001239f
C466 outputibias.n115 gnd 5.55e-19
C467 outputibias.n116 gnd 5.24e-19
C468 outputibias.n117 gnd 9.76e-19
C469 outputibias.n118 gnd 9.76e-19
C470 outputibias.n119 gnd 5.24e-19
C471 outputibias.n120 gnd 5.55e-19
C472 outputibias.n121 gnd 0.001239f
C473 outputibias.n122 gnd 0.002683f
C474 outputibias.n123 gnd 5.55e-19
C475 outputibias.n124 gnd 5.24e-19
C476 outputibias.n125 gnd 0.002256f
C477 outputibias.n126 gnd 0.005197f
C478 outputibias.n127 gnd 0.084814f
C479 outputibias.t4 gnd 0.108319f
C480 outputibias.t2 gnd 0.108319f
C481 outputibias.t0 gnd 0.108319f
C482 outputibias.t6 gnd 0.109238f
C483 outputibias.n128 gnd 0.134674f
C484 outputibias.n129 gnd 0.07244f
C485 outputibias.n130 gnd 0.079818f
C486 outputibias.n131 gnd 0.164901f
C487 outputibias.t11 gnd 0.11477f
C488 outputibias.n132 gnd 0.067481f
C489 outputibias.t8 gnd 0.11477f
C490 outputibias.n133 gnd 0.065115f
C491 outputibias.n134 gnd 0.029159f
C492 diffpairibias.t27 gnd 0.090128f
C493 diffpairibias.t23 gnd 0.08996f
C494 diffpairibias.n0 gnd 0.105991f
C495 diffpairibias.t28 gnd 0.08996f
C496 diffpairibias.n1 gnd 0.051736f
C497 diffpairibias.t25 gnd 0.08996f
C498 diffpairibias.n2 gnd 0.051736f
C499 diffpairibias.t29 gnd 0.08996f
C500 diffpairibias.n3 gnd 0.041084f
C501 diffpairibias.t15 gnd 0.086371f
C502 diffpairibias.t1 gnd 0.085993f
C503 diffpairibias.n4 gnd 0.13579f
C504 diffpairibias.t11 gnd 0.085993f
C505 diffpairibias.n5 gnd 0.072463f
C506 diffpairibias.t13 gnd 0.085993f
C507 diffpairibias.n6 gnd 0.072463f
C508 diffpairibias.t7 gnd 0.085993f
C509 diffpairibias.n7 gnd 0.072463f
C510 diffpairibias.t3 gnd 0.085993f
C511 diffpairibias.n8 gnd 0.072463f
C512 diffpairibias.t17 gnd 0.085993f
C513 diffpairibias.n9 gnd 0.072463f
C514 diffpairibias.t5 gnd 0.085993f
C515 diffpairibias.n10 gnd 0.072463f
C516 diffpairibias.t19 gnd 0.085993f
C517 diffpairibias.n11 gnd 0.072463f
C518 diffpairibias.t9 gnd 0.085993f
C519 diffpairibias.n12 gnd 0.102883f
C520 diffpairibias.t14 gnd 0.086899f
C521 diffpairibias.t0 gnd 0.086748f
C522 diffpairibias.n13 gnd 0.094648f
C523 diffpairibias.t10 gnd 0.086748f
C524 diffpairibias.n14 gnd 0.052262f
C525 diffpairibias.t12 gnd 0.086748f
C526 diffpairibias.n15 gnd 0.052262f
C527 diffpairibias.t6 gnd 0.086748f
C528 diffpairibias.n16 gnd 0.052262f
C529 diffpairibias.t2 gnd 0.086748f
C530 diffpairibias.n17 gnd 0.052262f
C531 diffpairibias.t16 gnd 0.086748f
C532 diffpairibias.n18 gnd 0.052262f
C533 diffpairibias.t4 gnd 0.086748f
C534 diffpairibias.n19 gnd 0.052262f
C535 diffpairibias.t18 gnd 0.086748f
C536 diffpairibias.n20 gnd 0.052262f
C537 diffpairibias.t8 gnd 0.086748f
C538 diffpairibias.n21 gnd 0.061849f
C539 diffpairibias.n22 gnd 0.233513f
C540 diffpairibias.t20 gnd 0.08996f
C541 diffpairibias.n23 gnd 0.051747f
C542 diffpairibias.t26 gnd 0.08996f
C543 diffpairibias.n24 gnd 0.051736f
C544 diffpairibias.t22 gnd 0.08996f
C545 diffpairibias.n25 gnd 0.051736f
C546 diffpairibias.t21 gnd 0.08996f
C547 diffpairibias.n26 gnd 0.051736f
C548 diffpairibias.t24 gnd 0.08996f
C549 diffpairibias.n27 gnd 0.04729f
C550 diffpairibias.n28 gnd 0.047711f
C551 a_n3827_n3924.t21 gnd 0.095164f
C552 a_n3827_n3924.t32 gnd 0.989057f
C553 a_n3827_n3924.n0 gnd 0.373908f
C554 a_n3827_n3924.t57 gnd 1.2292f
C555 a_n3827_n3924.n1 gnd 1.25966f
C556 a_n3827_n3924.t50 gnd 0.989057f
C557 a_n3827_n3924.n2 gnd 0.373908f
C558 a_n3827_n3924.t14 gnd 0.095164f
C559 a_n3827_n3924.t42 gnd 0.095164f
C560 a_n3827_n3924.n3 gnd 0.777221f
C561 a_n3827_n3924.n4 gnd 0.391675f
C562 a_n3827_n3924.t10 gnd 0.095164f
C563 a_n3827_n3924.t13 gnd 0.095164f
C564 a_n3827_n3924.n5 gnd 0.777221f
C565 a_n3827_n3924.n6 gnd 0.391675f
C566 a_n3827_n3924.t2 gnd 0.095164f
C567 a_n3827_n3924.t9 gnd 0.095164f
C568 a_n3827_n3924.n7 gnd 0.777221f
C569 a_n3827_n3924.n8 gnd 0.391675f
C570 a_n3827_n3924.t40 gnd 0.095164f
C571 a_n3827_n3924.t43 gnd 0.095164f
C572 a_n3827_n3924.n9 gnd 0.777221f
C573 a_n3827_n3924.n10 gnd 0.391675f
C574 a_n3827_n3924.t54 gnd 0.095164f
C575 a_n3827_n3924.t39 gnd 0.095164f
C576 a_n3827_n3924.n11 gnd 0.777221f
C577 a_n3827_n3924.n12 gnd 0.391675f
C578 a_n3827_n3924.t47 gnd 0.989057f
C579 a_n3827_n3924.n13 gnd 0.925833f
C580 a_n3827_n3924.t0 gnd 1.23041f
C581 a_n3827_n3924.t52 gnd 1.22888f
C582 a_n3827_n3924.n14 gnd 0.823361f
C583 a_n3827_n3924.t46 gnd 1.22888f
C584 a_n3827_n3924.n15 gnd 0.865521f
C585 a_n3827_n3924.t12 gnd 1.22888f
C586 a_n3827_n3924.n16 gnd 0.865521f
C587 a_n3827_n3924.t48 gnd 1.22888f
C588 a_n3827_n3924.n17 gnd 0.865521f
C589 a_n3827_n3924.t49 gnd 1.22888f
C590 a_n3827_n3924.n18 gnd 0.865521f
C591 a_n3827_n3924.t51 gnd 1.22888f
C592 a_n3827_n3924.n19 gnd 0.865521f
C593 a_n3827_n3924.t45 gnd 1.22888f
C594 a_n3827_n3924.n20 gnd 0.865521f
C595 a_n3827_n3924.t6 gnd 1.22888f
C596 a_n3827_n3924.n21 gnd 0.565437f
C597 a_n3827_n3924.n22 gnd 1.00053f
C598 a_n3827_n3924.n23 gnd 0.897154f
C599 a_n3827_n3924.t23 gnd 0.989054f
C600 a_n3827_n3924.n24 gnd 0.61435f
C601 a_n3827_n3924.t20 gnd 0.095164f
C602 a_n3827_n3924.t37 gnd 0.095164f
C603 a_n3827_n3924.n25 gnd 0.777219f
C604 a_n3827_n3924.n26 gnd 0.391677f
C605 a_n3827_n3924.t31 gnd 0.095164f
C606 a_n3827_n3924.t35 gnd 0.095164f
C607 a_n3827_n3924.n27 gnd 0.777219f
C608 a_n3827_n3924.n28 gnd 0.391677f
C609 a_n3827_n3924.t36 gnd 0.095164f
C610 a_n3827_n3924.t24 gnd 0.095164f
C611 a_n3827_n3924.n29 gnd 0.777219f
C612 a_n3827_n3924.n30 gnd 0.391677f
C613 a_n3827_n3924.t25 gnd 0.095164f
C614 a_n3827_n3924.t16 gnd 0.095164f
C615 a_n3827_n3924.n31 gnd 0.777219f
C616 a_n3827_n3924.n32 gnd 0.391677f
C617 a_n3827_n3924.t18 gnd 0.095164f
C618 a_n3827_n3924.t34 gnd 0.095164f
C619 a_n3827_n3924.n33 gnd 0.777219f
C620 a_n3827_n3924.n34 gnd 0.391677f
C621 a_n3827_n3924.t29 gnd 0.989054f
C622 a_n3827_n3924.n35 gnd 0.373911f
C623 a_n3827_n3924.t5 gnd 0.989054f
C624 a_n3827_n3924.n36 gnd 0.373911f
C625 a_n3827_n3924.t53 gnd 0.095164f
C626 a_n3827_n3924.t3 gnd 0.095164f
C627 a_n3827_n3924.n37 gnd 0.777219f
C628 a_n3827_n3924.n38 gnd 0.391677f
C629 a_n3827_n3924.t55 gnd 0.095164f
C630 a_n3827_n3924.t56 gnd 0.095164f
C631 a_n3827_n3924.n39 gnd 0.777219f
C632 a_n3827_n3924.n40 gnd 0.391677f
C633 a_n3827_n3924.t4 gnd 0.095164f
C634 a_n3827_n3924.t1 gnd 0.095164f
C635 a_n3827_n3924.n41 gnd 0.777219f
C636 a_n3827_n3924.n42 gnd 0.391677f
C637 a_n3827_n3924.t41 gnd 0.095164f
C638 a_n3827_n3924.t44 gnd 0.095164f
C639 a_n3827_n3924.n43 gnd 0.777219f
C640 a_n3827_n3924.n44 gnd 0.391677f
C641 a_n3827_n3924.t11 gnd 0.095164f
C642 a_n3827_n3924.t7 gnd 0.095164f
C643 a_n3827_n3924.n45 gnd 0.777219f
C644 a_n3827_n3924.n46 gnd 0.391677f
C645 a_n3827_n3924.t8 gnd 0.989054f
C646 a_n3827_n3924.n47 gnd 0.61435f
C647 a_n3827_n3924.n48 gnd 0.897154f
C648 a_n3827_n3924.t19 gnd 0.989053f
C649 a_n3827_n3924.n49 gnd 0.925837f
C650 a_n3827_n3924.t17 gnd 0.095164f
C651 a_n3827_n3924.t15 gnd 0.095164f
C652 a_n3827_n3924.n50 gnd 0.777221f
C653 a_n3827_n3924.n51 gnd 0.391675f
C654 a_n3827_n3924.t28 gnd 0.095164f
C655 a_n3827_n3924.t33 gnd 0.095164f
C656 a_n3827_n3924.n52 gnd 0.777221f
C657 a_n3827_n3924.n53 gnd 0.391675f
C658 a_n3827_n3924.t26 gnd 0.095164f
C659 a_n3827_n3924.t30 gnd 0.095164f
C660 a_n3827_n3924.n54 gnd 0.777221f
C661 a_n3827_n3924.n55 gnd 0.391675f
C662 a_n3827_n3924.t22 gnd 0.095164f
C663 a_n3827_n3924.t27 gnd 0.095164f
C664 a_n3827_n3924.n56 gnd 0.777221f
C665 a_n3827_n3924.n57 gnd 0.391675f
C666 a_n3827_n3924.n58 gnd 0.391674f
C667 a_n3827_n3924.n59 gnd 0.777222f
C668 a_n3827_n3924.t38 gnd 0.095164f
C669 plus.n0 gnd 0.023283f
C670 plus.t20 gnd 0.423413f
C671 plus.t23 gnd 0.391505f
C672 plus.n1 gnd 0.158342f
C673 plus.n2 gnd 0.023283f
C674 plus.t6 gnd 0.391505f
C675 plus.n3 gnd 0.019896f
C676 plus.n4 gnd 0.023283f
C677 plus.t12 gnd 0.391505f
C678 plus.t8 gnd 0.391505f
C679 plus.n5 gnd 0.158342f
C680 plus.n6 gnd 0.023283f
C681 plus.t7 gnd 0.391505f
C682 plus.n7 gnd 0.158342f
C683 plus.n8 gnd 0.023283f
C684 plus.t19 gnd 0.391505f
C685 plus.n9 gnd 0.018924f
C686 plus.n10 gnd 0.023283f
C687 plus.t18 gnd 0.391505f
C688 plus.t27 gnd 0.391505f
C689 plus.n11 gnd 0.158342f
C690 plus.n12 gnd 0.023283f
C691 plus.t25 gnd 0.391505f
C692 plus.n13 gnd 0.158342f
C693 plus.n14 gnd 0.098812f
C694 plus.t9 gnd 0.391505f
C695 plus.t14 gnd 0.43797f
C696 plus.n15 gnd 0.185118f
C697 plus.n16 gnd 0.181331f
C698 plus.n17 gnd 0.029834f
C699 plus.n18 gnd 0.026348f
C700 plus.n19 gnd 0.023283f
C701 plus.n20 gnd 0.023283f
C702 plus.n21 gnd 0.027824f
C703 plus.n22 gnd 0.019896f
C704 plus.n23 gnd 0.030323f
C705 plus.n24 gnd 0.023283f
C706 plus.n25 gnd 0.023283f
C707 plus.n26 gnd 0.028962f
C708 plus.n27 gnd 0.027219f
C709 plus.n28 gnd 0.158342f
C710 plus.n29 gnd 0.029166f
C711 plus.n30 gnd 0.023283f
C712 plus.n31 gnd 0.023283f
C713 plus.n32 gnd 0.023283f
C714 plus.n33 gnd 0.029953f
C715 plus.n34 gnd 0.158342f
C716 plus.n35 gnd 0.028091f
C717 plus.n36 gnd 0.028091f
C718 plus.n37 gnd 0.023283f
C719 plus.n38 gnd 0.023283f
C720 plus.n39 gnd 0.029953f
C721 plus.n40 gnd 0.018924f
C722 plus.n41 gnd 0.029166f
C723 plus.n42 gnd 0.023283f
C724 plus.n43 gnd 0.023283f
C725 plus.n44 gnd 0.027219f
C726 plus.n45 gnd 0.028962f
C727 plus.n46 gnd 0.158342f
C728 plus.n47 gnd 0.030323f
C729 plus.n48 gnd 0.023283f
C730 plus.n49 gnd 0.023283f
C731 plus.n50 gnd 0.023283f
C732 plus.n51 gnd 0.027824f
C733 plus.n52 gnd 0.158342f
C734 plus.n53 gnd 0.026348f
C735 plus.n54 gnd 0.029834f
C736 plus.n55 gnd 0.023283f
C737 plus.n56 gnd 0.023283f
C738 plus.n57 gnd 0.030374f
C739 plus.n58 gnd 0.008462f
C740 plus.n59 gnd 0.183334f
C741 plus.n60 gnd 0.266765f
C742 plus.n61 gnd 0.023283f
C743 plus.t28 gnd 0.391505f
C744 plus.n62 gnd 0.158342f
C745 plus.n63 gnd 0.023283f
C746 plus.t26 gnd 0.391505f
C747 plus.n64 gnd 0.019896f
C748 plus.n65 gnd 0.023283f
C749 plus.t10 gnd 0.391505f
C750 plus.t15 gnd 0.391505f
C751 plus.n66 gnd 0.158342f
C752 plus.n67 gnd 0.023283f
C753 plus.t13 gnd 0.391505f
C754 plus.n68 gnd 0.158342f
C755 plus.n69 gnd 0.023283f
C756 plus.t17 gnd 0.391505f
C757 plus.n70 gnd 0.018924f
C758 plus.n71 gnd 0.023283f
C759 plus.t16 gnd 0.391505f
C760 plus.t21 gnd 0.391505f
C761 plus.n72 gnd 0.158342f
C762 plus.n73 gnd 0.023283f
C763 plus.t22 gnd 0.391505f
C764 plus.n74 gnd 0.158342f
C765 plus.n75 gnd 0.098812f
C766 plus.t5 gnd 0.391505f
C767 plus.t11 gnd 0.43797f
C768 plus.n76 gnd 0.185118f
C769 plus.n77 gnd 0.181331f
C770 plus.n78 gnd 0.029834f
C771 plus.n79 gnd 0.026348f
C772 plus.n80 gnd 0.023283f
C773 plus.n81 gnd 0.023283f
C774 plus.n82 gnd 0.027824f
C775 plus.n83 gnd 0.019896f
C776 plus.n84 gnd 0.030323f
C777 plus.n85 gnd 0.023283f
C778 plus.n86 gnd 0.023283f
C779 plus.n87 gnd 0.028962f
C780 plus.n88 gnd 0.027219f
C781 plus.n89 gnd 0.158342f
C782 plus.n90 gnd 0.029166f
C783 plus.n91 gnd 0.023283f
C784 plus.n92 gnd 0.023283f
C785 plus.n93 gnd 0.023283f
C786 plus.n94 gnd 0.029953f
C787 plus.n95 gnd 0.158342f
C788 plus.n96 gnd 0.028091f
C789 plus.n97 gnd 0.028091f
C790 plus.n98 gnd 0.023283f
C791 plus.n99 gnd 0.023283f
C792 plus.n100 gnd 0.029953f
C793 plus.n101 gnd 0.018924f
C794 plus.n102 gnd 0.029166f
C795 plus.n103 gnd 0.023283f
C796 plus.n104 gnd 0.023283f
C797 plus.n105 gnd 0.027219f
C798 plus.n106 gnd 0.028962f
C799 plus.n107 gnd 0.158342f
C800 plus.n108 gnd 0.030323f
C801 plus.n109 gnd 0.023283f
C802 plus.n110 gnd 0.023283f
C803 plus.n111 gnd 0.023283f
C804 plus.n112 gnd 0.027824f
C805 plus.n113 gnd 0.158342f
C806 plus.n114 gnd 0.026348f
C807 plus.n115 gnd 0.029834f
C808 plus.n116 gnd 0.023283f
C809 plus.n117 gnd 0.023283f
C810 plus.n118 gnd 0.030374f
C811 plus.n119 gnd 0.008462f
C812 plus.t24 gnd 0.423413f
C813 plus.n120 gnd 0.183334f
C814 plus.n121 gnd 0.840053f
C815 plus.n122 gnd 1.23841f
C816 plus.t1 gnd 0.040194f
C817 plus.t2 gnd 0.007178f
C818 plus.t4 gnd 0.007178f
C819 plus.n123 gnd 0.023278f
C820 plus.n124 gnd 0.18071f
C821 plus.t3 gnd 0.007178f
C822 plus.t0 gnd 0.007178f
C823 plus.n125 gnd 0.023278f
C824 plus.n126 gnd 0.135645f
C825 plus.n127 gnd 2.80941f
C826 a_n1808_13878.t4 gnd 0.185195f
C827 a_n1808_13878.t0 gnd 0.185195f
C828 a_n1808_13878.t2 gnd 0.185195f
C829 a_n1808_13878.n0 gnd 1.4598f
C830 a_n1808_13878.t6 gnd 0.185195f
C831 a_n1808_13878.t1 gnd 0.185195f
C832 a_n1808_13878.n1 gnd 1.45825f
C833 a_n1808_13878.n2 gnd 2.03762f
C834 a_n1808_13878.t5 gnd 0.185195f
C835 a_n1808_13878.t9 gnd 0.185195f
C836 a_n1808_13878.n3 gnd 1.46067f
C837 a_n1808_13878.t10 gnd 0.185195f
C838 a_n1808_13878.t3 gnd 0.185195f
C839 a_n1808_13878.n4 gnd 1.45825f
C840 a_n1808_13878.n5 gnd 1.31079f
C841 a_n1808_13878.t7 gnd 0.185195f
C842 a_n1808_13878.t8 gnd 0.185195f
C843 a_n1808_13878.n6 gnd 1.45825f
C844 a_n1808_13878.n7 gnd 1.80025f
C845 a_n1808_13878.t13 gnd 1.73408f
C846 a_n1808_13878.t16 gnd 0.185195f
C847 a_n1808_13878.t17 gnd 0.185195f
C848 a_n1808_13878.n8 gnd 1.30452f
C849 a_n1808_13878.n9 gnd 1.4576f
C850 a_n1808_13878.t12 gnd 1.73062f
C851 a_n1808_13878.n10 gnd 0.733487f
C852 a_n1808_13878.t15 gnd 1.73062f
C853 a_n1808_13878.n11 gnd 0.733487f
C854 a_n1808_13878.t18 gnd 0.185195f
C855 a_n1808_13878.t19 gnd 0.185195f
C856 a_n1808_13878.n12 gnd 1.30452f
C857 a_n1808_13878.n13 gnd 0.74059f
C858 a_n1808_13878.t14 gnd 1.73062f
C859 a_n1808_13878.n14 gnd 1.7272f
C860 a_n1808_13878.n15 gnd 2.51438f
C861 a_n1808_13878.n16 gnd 3.69301f
C862 a_n1808_13878.n17 gnd 1.45826f
C863 a_n1808_13878.t11 gnd 0.185195f
C864 a_n1986_8322.t2 gnd 38.652897f
C865 a_n1986_8322.t0 gnd 28.1251f
C866 a_n1986_8322.t3 gnd 19.258501f
C867 a_n1986_8322.t1 gnd 38.652897f
C868 a_n1986_8322.t6 gnd 0.093486f
C869 a_n1986_8322.t5 gnd 0.875352f
C870 a_n1986_8322.t13 gnd 0.093486f
C871 a_n1986_8322.t8 gnd 0.093486f
C872 a_n1986_8322.n0 gnd 0.658513f
C873 a_n1986_8322.n1 gnd 0.735791f
C874 a_n1986_8322.t11 gnd 0.093486f
C875 a_n1986_8322.t10 gnd 0.093486f
C876 a_n1986_8322.n2 gnd 0.658513f
C877 a_n1986_8322.n3 gnd 0.373846f
C878 a_n1986_8322.t4 gnd 0.873609f
C879 a_n1986_8322.n4 gnd 1.39826f
C880 a_n1986_8322.t18 gnd 0.875352f
C881 a_n1986_8322.t22 gnd 0.093486f
C882 a_n1986_8322.t21 gnd 0.093486f
C883 a_n1986_8322.n5 gnd 0.658513f
C884 a_n1986_8322.n6 gnd 0.735791f
C885 a_n1986_8322.t16 gnd 0.873609f
C886 a_n1986_8322.n7 gnd 0.37026f
C887 a_n1986_8322.t19 gnd 0.873609f
C888 a_n1986_8322.n8 gnd 0.37026f
C889 a_n1986_8322.t17 gnd 0.093486f
C890 a_n1986_8322.t23 gnd 0.093486f
C891 a_n1986_8322.n9 gnd 0.658513f
C892 a_n1986_8322.n10 gnd 0.373846f
C893 a_n1986_8322.t20 gnd 0.873609f
C894 a_n1986_8322.n11 gnd 0.871879f
C895 a_n1986_8322.n12 gnd 1.58991f
C896 a_n1986_8322.n13 gnd 3.44798f
C897 a_n1986_8322.t7 gnd 0.873609f
C898 a_n1986_8322.n14 gnd 0.766135f
C899 a_n1986_8322.t14 gnd 0.875349f
C900 a_n1986_8322.t12 gnd 0.093486f
C901 a_n1986_8322.t9 gnd 0.093486f
C902 a_n1986_8322.n15 gnd 0.658513f
C903 a_n1986_8322.n16 gnd 0.735793f
C904 a_n1986_8322.n17 gnd 0.373844f
C905 a_n1986_8322.n18 gnd 0.658514f
C906 a_n1986_8322.t15 gnd 0.093486f
C907 a_n2848_n452.n0 gnd 0.492472f
C908 a_n2848_n452.n1 gnd 0.664435f
C909 a_n2848_n452.n2 gnd 0.215942f
C910 a_n2848_n452.n3 gnd 0.282512f
C911 a_n2848_n452.n4 gnd 0.438486f
C912 a_n2848_n452.n5 gnd 2.99175f
C913 a_n2848_n452.n6 gnd 0.526038f
C914 a_n2848_n452.n7 gnd 0.204894f
C915 a_n2848_n452.n8 gnd 0.150908f
C916 a_n2848_n452.n9 gnd 0.23718f
C917 a_n2848_n452.n10 gnd 0.183194f
C918 a_n2848_n452.n11 gnd 0.204894f
C919 a_n2848_n452.n12 gnd 0.150908f
C920 a_n2848_n452.n13 gnd 0.580023f
C921 a_n2848_n452.n14 gnd 0.432289f
C922 a_n2848_n452.n15 gnd 0.215942f
C923 a_n2848_n452.n16 gnd 0.492472f
C924 a_n2848_n452.n17 gnd 0.282512f
C925 a_n2848_n452.n18 gnd 0.438486f
C926 a_n2848_n452.n19 gnd 0.215942f
C927 a_n2848_n452.n20 gnd 0.731535f
C928 a_n2848_n452.n21 gnd 0.282512f
C929 a_n2848_n452.n22 gnd 1.77783f
C930 a_n2848_n452.n23 gnd 1.91568f
C931 a_n2848_n452.n24 gnd 0.377489f
C932 a_n2848_n452.n25 gnd 3.11576f
C933 a_n2848_n452.n26 gnd 0.377488f
C934 a_n2848_n452.n27 gnd 3.20158f
C935 a_n2848_n452.n28 gnd 0.008361f
C936 a_n2848_n452.n30 gnd 0.285666f
C937 a_n2848_n452.n31 gnd 0.008361f
C938 a_n2848_n452.n33 gnd 0.285666f
C939 a_n2848_n452.n34 gnd 0.008361f
C940 a_n2848_n452.n35 gnd 0.28526f
C941 a_n2848_n452.n36 gnd 0.008361f
C942 a_n2848_n452.n37 gnd 0.28526f
C943 a_n2848_n452.n38 gnd 0.008361f
C944 a_n2848_n452.n39 gnd 0.28526f
C945 a_n2848_n452.n40 gnd 0.008361f
C946 a_n2848_n452.n41 gnd 1.33845f
C947 a_n2848_n452.n42 gnd 0.28526f
C948 a_n2848_n452.n44 gnd 0.285666f
C949 a_n2848_n452.n45 gnd 0.008361f
C950 a_n2848_n452.n47 gnd 0.285666f
C951 a_n2848_n452.n49 gnd 0.302425f
C952 a_n2848_n452.t26 gnd 0.696704f
C953 a_n2848_n452.n50 gnd 0.306315f
C954 a_n2848_n452.t28 gnd 0.696704f
C955 a_n2848_n452.t30 gnd 0.696704f
C956 a_n2848_n452.t56 gnd 0.696704f
C957 a_n2848_n452.n51 gnd 0.306315f
C958 a_n2848_n452.t65 gnd 0.696704f
C959 a_n2848_n452.t71 gnd 0.696704f
C960 a_n2848_n452.t12 gnd 0.696704f
C961 a_n2848_n452.t22 gnd 0.696704f
C962 a_n2848_n452.t16 gnd 0.696704f
C963 a_n2848_n452.t14 gnd 0.696704f
C964 a_n2848_n452.t75 gnd 0.711378f
C965 a_n2848_n452.t58 gnd 0.696704f
C966 a_n2848_n452.t62 gnd 0.696704f
C967 a_n2848_n452.t52 gnd 0.696704f
C968 a_n2848_n452.n52 gnd 0.306315f
C969 a_n2848_n452.t67 gnd 0.696704f
C970 a_n2848_n452.t73 gnd 0.708223f
C971 a_n2848_n452.n53 gnd 0.308933f
C972 a_n2848_n452.n54 gnd 0.302425f
C973 a_n2848_n452.n55 gnd 0.308932f
C974 a_n2848_n452.t24 gnd 0.708223f
C975 a_n2848_n452.n56 gnd 0.308933f
C976 a_n2848_n452.t20 gnd 0.696704f
C977 a_n2848_n452.n57 gnd 0.302425f
C978 a_n2848_n452.n58 gnd 0.01225f
C979 a_n2848_n452.t4 gnd 0.116496f
C980 a_n2848_n452.t44 gnd 0.116496f
C981 a_n2848_n452.n59 gnd 1.03243f
C982 a_n2848_n452.t2 gnd 0.116496f
C983 a_n2848_n452.t46 gnd 0.116496f
C984 a_n2848_n452.n60 gnd 1.0294f
C985 a_n2848_n452.n61 gnd 0.912817f
C986 a_n2848_n452.t47 gnd 0.116496f
C987 a_n2848_n452.t3 gnd 0.116496f
C988 a_n2848_n452.n62 gnd 1.0294f
C989 a_n2848_n452.t5 gnd 0.116496f
C990 a_n2848_n452.t6 gnd 0.116496f
C991 a_n2848_n452.n63 gnd 1.03243f
C992 a_n2848_n452.t41 gnd 0.116496f
C993 a_n2848_n452.t9 gnd 0.116496f
C994 a_n2848_n452.n64 gnd 1.0294f
C995 a_n2848_n452.n65 gnd 0.912817f
C996 a_n2848_n452.t0 gnd 0.116496f
C997 a_n2848_n452.t38 gnd 0.116496f
C998 a_n2848_n452.n66 gnd 1.0294f
C999 a_n2848_n452.t42 gnd 0.116496f
C1000 a_n2848_n452.t45 gnd 0.116496f
C1001 a_n2848_n452.n67 gnd 1.0294f
C1002 a_n2848_n452.n68 gnd 3.15028f
C1003 a_n2848_n452.t36 gnd 0.116496f
C1004 a_n2848_n452.t37 gnd 0.116496f
C1005 a_n2848_n452.n69 gnd 1.0294f
C1006 a_n2848_n452.n70 gnd 0.449443f
C1007 a_n2848_n452.t40 gnd 0.116496f
C1008 a_n2848_n452.t1 gnd 0.116496f
C1009 a_n2848_n452.n71 gnd 1.0294f
C1010 a_n2848_n452.t39 gnd 0.116496f
C1011 a_n2848_n452.t43 gnd 0.116496f
C1012 a_n2848_n452.n72 gnd 1.03243f
C1013 a_n2848_n452.t34 gnd 0.116496f
C1014 a_n2848_n452.t35 gnd 0.116496f
C1015 a_n2848_n452.n73 gnd 1.0294f
C1016 a_n2848_n452.n74 gnd 0.912815f
C1017 a_n2848_n452.t7 gnd 0.116496f
C1018 a_n2848_n452.t8 gnd 0.116496f
C1019 a_n2848_n452.n75 gnd 1.0294f
C1020 a_n2848_n452.n76 gnd 0.2971f
C1021 a_n2848_n452.n77 gnd 0.01225f
C1022 a_n2848_n452.n78 gnd 0.296767f
C1023 a_n2848_n452.n79 gnd 0.531228f
C1024 a_n2848_n452.t25 gnd 1.40246f
C1025 a_n2848_n452.t21 gnd 0.14978f
C1026 a_n2848_n452.t15 gnd 0.14978f
C1027 a_n2848_n452.n80 gnd 1.05505f
C1028 a_n2848_n452.t17 gnd 0.14978f
C1029 a_n2848_n452.t23 gnd 0.14978f
C1030 a_n2848_n452.n81 gnd 1.05505f
C1031 a_n2848_n452.t13 gnd 1.39967f
C1032 a_n2848_n452.n82 gnd 1.14458f
C1033 a_n2848_n452.n83 gnd 0.786935f
C1034 a_n2848_n452.t57 gnd 0.696704f
C1035 a_n2848_n452.t66 gnd 0.696704f
C1036 a_n2848_n452.t48 gnd 0.696704f
C1037 a_n2848_n452.n84 gnd 0.306315f
C1038 a_n2848_n452.t68 gnd 0.696704f
C1039 a_n2848_n452.t53 gnd 0.696704f
C1040 a_n2848_n452.t54 gnd 0.696704f
C1041 a_n2848_n452.n85 gnd 0.306315f
C1042 a_n2848_n452.t72 gnd 0.696704f
C1043 a_n2848_n452.t61 gnd 0.696704f
C1044 a_n2848_n452.t60 gnd 0.696704f
C1045 a_n2848_n452.n86 gnd 0.306315f
C1046 a_n2848_n452.t64 gnd 0.696704f
C1047 a_n2848_n452.t55 gnd 0.696704f
C1048 a_n2848_n452.t49 gnd 0.696704f
C1049 a_n2848_n452.n87 gnd 0.306315f
C1050 a_n2848_n452.t69 gnd 0.708378f
C1051 a_n2848_n452.n88 gnd 0.302425f
C1052 a_n2848_n452.n89 gnd 0.296933f
C1053 a_n2848_n452.t74 gnd 0.708378f
C1054 a_n2848_n452.n90 gnd 0.302425f
C1055 a_n2848_n452.n91 gnd 0.296933f
C1056 a_n2848_n452.t63 gnd 0.708378f
C1057 a_n2848_n452.n92 gnd 0.302425f
C1058 a_n2848_n452.n93 gnd 0.296933f
C1059 a_n2848_n452.t59 gnd 0.708378f
C1060 a_n2848_n452.n94 gnd 0.302425f
C1061 a_n2848_n452.n95 gnd 0.296933f
C1062 a_n2848_n452.n96 gnd 1.0063f
C1063 a_n2848_n452.t70 gnd 0.711378f
C1064 a_n2848_n452.n97 gnd 0.308932f
C1065 a_n2848_n452.t50 gnd 0.696704f
C1066 a_n2848_n452.n98 gnd 0.302425f
C1067 a_n2848_n452.n99 gnd 0.308933f
C1068 a_n2848_n452.t51 gnd 0.708223f
C1069 a_n2848_n452.t10 gnd 0.711378f
C1070 a_n2848_n452.n100 gnd 0.308932f
C1071 a_n2848_n452.t32 gnd 0.696704f
C1072 a_n2848_n452.n101 gnd 0.302425f
C1073 a_n2848_n452.n102 gnd 0.308933f
C1074 a_n2848_n452.t18 gnd 0.708223f
C1075 a_n2848_n452.n103 gnd 1.13204f
C1076 a_n2848_n452.t19 gnd 1.39967f
C1077 a_n2848_n452.t27 gnd 0.14978f
C1078 a_n2848_n452.t29 gnd 0.14978f
C1079 a_n2848_n452.n104 gnd 1.05505f
C1080 a_n2848_n452.t31 gnd 0.14978f
C1081 a_n2848_n452.t33 gnd 0.14978f
C1082 a_n2848_n452.n105 gnd 1.05505f
C1083 a_n2848_n452.n106 gnd 1.17886f
C1084 a_n2848_n452.t11 gnd 1.40246f
C1085 CSoutput.n0 gnd 0.041285f
C1086 CSoutput.t144 gnd 0.273089f
C1087 CSoutput.n1 gnd 0.123313f
C1088 CSoutput.n2 gnd 0.041285f
C1089 CSoutput.t149 gnd 0.273089f
C1090 CSoutput.n3 gnd 0.032721f
C1091 CSoutput.n4 gnd 0.041285f
C1092 CSoutput.t158 gnd 0.273089f
C1093 CSoutput.n5 gnd 0.028216f
C1094 CSoutput.n6 gnd 0.041285f
C1095 CSoutput.t147 gnd 0.273089f
C1096 CSoutput.t151 gnd 0.273089f
C1097 CSoutput.n7 gnd 0.121969f
C1098 CSoutput.n8 gnd 0.041285f
C1099 CSoutput.t157 gnd 0.273089f
C1100 CSoutput.n9 gnd 0.026902f
C1101 CSoutput.n10 gnd 0.041285f
C1102 CSoutput.t160 gnd 0.273089f
C1103 CSoutput.t148 gnd 0.273089f
C1104 CSoutput.n11 gnd 0.121969f
C1105 CSoutput.n12 gnd 0.041285f
C1106 CSoutput.t154 gnd 0.273089f
C1107 CSoutput.n13 gnd 0.028216f
C1108 CSoutput.n14 gnd 0.041285f
C1109 CSoutput.t153 gnd 0.273089f
C1110 CSoutput.t163 gnd 0.273089f
C1111 CSoutput.n15 gnd 0.121969f
C1112 CSoutput.n16 gnd 0.041285f
C1113 CSoutput.t152 gnd 0.273089f
C1114 CSoutput.n17 gnd 0.030136f
C1115 CSoutput.t161 gnd 0.326348f
C1116 CSoutput.t150 gnd 0.273089f
C1117 CSoutput.n18 gnd 0.155707f
C1118 CSoutput.n19 gnd 0.15109f
C1119 CSoutput.n20 gnd 0.175282f
C1120 CSoutput.n21 gnd 0.041285f
C1121 CSoutput.n22 gnd 0.034457f
C1122 CSoutput.n23 gnd 0.121969f
C1123 CSoutput.n24 gnd 0.033215f
C1124 CSoutput.n25 gnd 0.032721f
C1125 CSoutput.n26 gnd 0.041285f
C1126 CSoutput.n27 gnd 0.041285f
C1127 CSoutput.n28 gnd 0.034192f
C1128 CSoutput.n29 gnd 0.02903f
C1129 CSoutput.n30 gnd 0.124684f
C1130 CSoutput.n31 gnd 0.029429f
C1131 CSoutput.n32 gnd 0.041285f
C1132 CSoutput.n33 gnd 0.041285f
C1133 CSoutput.n34 gnd 0.041285f
C1134 CSoutput.n35 gnd 0.033827f
C1135 CSoutput.n36 gnd 0.121969f
C1136 CSoutput.n37 gnd 0.032351f
C1137 CSoutput.n38 gnd 0.033585f
C1138 CSoutput.n39 gnd 0.041285f
C1139 CSoutput.n40 gnd 0.041285f
C1140 CSoutput.n41 gnd 0.03445f
C1141 CSoutput.n42 gnd 0.031487f
C1142 CSoutput.n43 gnd 0.121969f
C1143 CSoutput.n44 gnd 0.032285f
C1144 CSoutput.n45 gnd 0.041285f
C1145 CSoutput.n46 gnd 0.041285f
C1146 CSoutput.n47 gnd 0.041285f
C1147 CSoutput.n48 gnd 0.032285f
C1148 CSoutput.n49 gnd 0.121969f
C1149 CSoutput.n50 gnd 0.031487f
C1150 CSoutput.n51 gnd 0.03445f
C1151 CSoutput.n52 gnd 0.041285f
C1152 CSoutput.n53 gnd 0.041285f
C1153 CSoutput.n54 gnd 0.033585f
C1154 CSoutput.n55 gnd 0.032351f
C1155 CSoutput.n56 gnd 0.121969f
C1156 CSoutput.n57 gnd 0.033827f
C1157 CSoutput.n58 gnd 0.041285f
C1158 CSoutput.n59 gnd 0.041285f
C1159 CSoutput.n60 gnd 0.041285f
C1160 CSoutput.n61 gnd 0.029429f
C1161 CSoutput.n62 gnd 0.124684f
C1162 CSoutput.n63 gnd 0.02903f
C1163 CSoutput.t159 gnd 0.273089f
C1164 CSoutput.n64 gnd 0.121969f
C1165 CSoutput.n65 gnd 0.034192f
C1166 CSoutput.n66 gnd 0.041285f
C1167 CSoutput.n67 gnd 0.041285f
C1168 CSoutput.n68 gnd 0.041285f
C1169 CSoutput.n69 gnd 0.033215f
C1170 CSoutput.n70 gnd 0.121969f
C1171 CSoutput.n71 gnd 0.034457f
C1172 CSoutput.n72 gnd 0.030136f
C1173 CSoutput.n73 gnd 0.041285f
C1174 CSoutput.n74 gnd 0.041285f
C1175 CSoutput.n75 gnd 0.031253f
C1176 CSoutput.n76 gnd 0.018561f
C1177 CSoutput.t162 gnd 0.306835f
C1178 CSoutput.n77 gnd 0.152423f
C1179 CSoutput.n78 gnd 0.623555f
C1180 CSoutput.t132 gnd 0.051497f
C1181 CSoutput.t72 gnd 0.051497f
C1182 CSoutput.n79 gnd 0.398705f
C1183 CSoutput.t120 gnd 0.051497f
C1184 CSoutput.t103 gnd 0.051497f
C1185 CSoutput.n80 gnd 0.397994f
C1186 CSoutput.n81 gnd 0.403963f
C1187 CSoutput.t127 gnd 0.051497f
C1188 CSoutput.t85 gnd 0.051497f
C1189 CSoutput.n82 gnd 0.397994f
C1190 CSoutput.n83 gnd 0.199056f
C1191 CSoutput.t138 gnd 0.051497f
C1192 CSoutput.t97 gnd 0.051497f
C1193 CSoutput.n84 gnd 0.397994f
C1194 CSoutput.n85 gnd 0.199056f
C1195 CSoutput.t76 gnd 0.051497f
C1196 CSoutput.t108 gnd 0.051497f
C1197 CSoutput.n86 gnd 0.397994f
C1198 CSoutput.n87 gnd 0.199056f
C1199 CSoutput.t80 gnd 0.051497f
C1200 CSoutput.t92 gnd 0.051497f
C1201 CSoutput.n88 gnd 0.397994f
C1202 CSoutput.n89 gnd 0.365023f
C1203 CSoutput.t130 gnd 0.051497f
C1204 CSoutput.t128 gnd 0.051497f
C1205 CSoutput.n90 gnd 0.398705f
C1206 CSoutput.t115 gnd 0.051497f
C1207 CSoutput.t78 gnd 0.051497f
C1208 CSoutput.n91 gnd 0.397994f
C1209 CSoutput.n92 gnd 0.403963f
C1210 CSoutput.t74 gnd 0.051497f
C1211 CSoutput.t126 gnd 0.051497f
C1212 CSoutput.n93 gnd 0.397994f
C1213 CSoutput.n94 gnd 0.199056f
C1214 CSoutput.t114 gnd 0.051497f
C1215 CSoutput.t100 gnd 0.051497f
C1216 CSoutput.n95 gnd 0.397994f
C1217 CSoutput.n96 gnd 0.199056f
C1218 CSoutput.t87 gnd 0.051497f
C1219 CSoutput.t134 gnd 0.051497f
C1220 CSoutput.n97 gnd 0.397994f
C1221 CSoutput.n98 gnd 0.199056f
C1222 CSoutput.t113 gnd 0.051497f
C1223 CSoutput.t112 gnd 0.051497f
C1224 CSoutput.n99 gnd 0.397994f
C1225 CSoutput.n100 gnd 0.296842f
C1226 CSoutput.n101 gnd 0.374317f
C1227 CSoutput.t136 gnd 0.051497f
C1228 CSoutput.t137 gnd 0.051497f
C1229 CSoutput.n102 gnd 0.398705f
C1230 CSoutput.t123 gnd 0.051497f
C1231 CSoutput.t84 gnd 0.051497f
C1232 CSoutput.n103 gnd 0.397994f
C1233 CSoutput.n104 gnd 0.403963f
C1234 CSoutput.t82 gnd 0.051497f
C1235 CSoutput.t135 gnd 0.051497f
C1236 CSoutput.n105 gnd 0.397994f
C1237 CSoutput.n106 gnd 0.199056f
C1238 CSoutput.t122 gnd 0.051497f
C1239 CSoutput.t107 gnd 0.051497f
C1240 CSoutput.n107 gnd 0.397994f
C1241 CSoutput.n108 gnd 0.199056f
C1242 CSoutput.t94 gnd 0.051497f
C1243 CSoutput.t142 gnd 0.051497f
C1244 CSoutput.n109 gnd 0.397994f
C1245 CSoutput.n110 gnd 0.199056f
C1246 CSoutput.t119 gnd 0.051497f
C1247 CSoutput.t118 gnd 0.051497f
C1248 CSoutput.n111 gnd 0.397994f
C1249 CSoutput.n112 gnd 0.296842f
C1250 CSoutput.n113 gnd 0.41839f
C1251 CSoutput.n114 gnd 7.55102f
C1252 CSoutput.n116 gnd 0.730317f
C1253 CSoutput.n117 gnd 0.547738f
C1254 CSoutput.n118 gnd 0.730317f
C1255 CSoutput.n119 gnd 0.730317f
C1256 CSoutput.n120 gnd 1.96624f
C1257 CSoutput.n121 gnd 0.730317f
C1258 CSoutput.n122 gnd 0.730317f
C1259 CSoutput.t155 gnd 0.912896f
C1260 CSoutput.n123 gnd 0.730317f
C1261 CSoutput.n124 gnd 0.730317f
C1262 CSoutput.n128 gnd 0.730317f
C1263 CSoutput.n132 gnd 0.730317f
C1264 CSoutput.n133 gnd 0.730317f
C1265 CSoutput.n135 gnd 0.730317f
C1266 CSoutput.n140 gnd 0.730317f
C1267 CSoutput.n142 gnd 0.730317f
C1268 CSoutput.n143 gnd 0.730317f
C1269 CSoutput.n145 gnd 0.730317f
C1270 CSoutput.n146 gnd 0.730317f
C1271 CSoutput.n148 gnd 0.730317f
C1272 CSoutput.t145 gnd 12.2035f
C1273 CSoutput.n150 gnd 0.730317f
C1274 CSoutput.n151 gnd 0.547738f
C1275 CSoutput.n152 gnd 0.730317f
C1276 CSoutput.n153 gnd 0.730317f
C1277 CSoutput.n154 gnd 1.96624f
C1278 CSoutput.n155 gnd 0.730317f
C1279 CSoutput.n156 gnd 0.730317f
C1280 CSoutput.t164 gnd 0.912896f
C1281 CSoutput.n157 gnd 0.730317f
C1282 CSoutput.n158 gnd 0.730317f
C1283 CSoutput.n162 gnd 0.730317f
C1284 CSoutput.n166 gnd 0.730317f
C1285 CSoutput.n167 gnd 0.730317f
C1286 CSoutput.n169 gnd 0.730317f
C1287 CSoutput.n174 gnd 0.730317f
C1288 CSoutput.n176 gnd 0.730317f
C1289 CSoutput.n177 gnd 0.730317f
C1290 CSoutput.n179 gnd 0.730317f
C1291 CSoutput.n180 gnd 0.730317f
C1292 CSoutput.n182 gnd 0.730317f
C1293 CSoutput.n183 gnd 0.547738f
C1294 CSoutput.n185 gnd 0.730317f
C1295 CSoutput.n186 gnd 0.547738f
C1296 CSoutput.n187 gnd 0.730317f
C1297 CSoutput.n188 gnd 0.730317f
C1298 CSoutput.n189 gnd 1.96624f
C1299 CSoutput.n190 gnd 0.730317f
C1300 CSoutput.n191 gnd 0.730317f
C1301 CSoutput.t156 gnd 0.912896f
C1302 CSoutput.n192 gnd 0.730317f
C1303 CSoutput.n193 gnd 1.96624f
C1304 CSoutput.n195 gnd 0.730317f
C1305 CSoutput.n196 gnd 0.730317f
C1306 CSoutput.n198 gnd 0.730317f
C1307 CSoutput.n199 gnd 0.730317f
C1308 CSoutput.t165 gnd 12.0046f
C1309 CSoutput.t146 gnd 12.2035f
C1310 CSoutput.n205 gnd 2.29111f
C1311 CSoutput.n206 gnd 9.33316f
C1312 CSoutput.n207 gnd 9.72369f
C1313 CSoutput.n212 gnd 2.48189f
C1314 CSoutput.n218 gnd 0.730317f
C1315 CSoutput.n220 gnd 0.730317f
C1316 CSoutput.n222 gnd 0.730317f
C1317 CSoutput.n224 gnd 0.730317f
C1318 CSoutput.n226 gnd 0.730317f
C1319 CSoutput.n232 gnd 0.730317f
C1320 CSoutput.n239 gnd 1.33985f
C1321 CSoutput.n240 gnd 1.33985f
C1322 CSoutput.n241 gnd 0.730317f
C1323 CSoutput.n242 gnd 0.730317f
C1324 CSoutput.n244 gnd 0.547738f
C1325 CSoutput.n245 gnd 0.469088f
C1326 CSoutput.n247 gnd 0.547738f
C1327 CSoutput.n248 gnd 0.469088f
C1328 CSoutput.n249 gnd 0.547738f
C1329 CSoutput.n251 gnd 0.730317f
C1330 CSoutput.n253 gnd 1.96624f
C1331 CSoutput.n254 gnd 2.29111f
C1332 CSoutput.n255 gnd 8.5841f
C1333 CSoutput.n257 gnd 0.547738f
C1334 CSoutput.n258 gnd 1.40936f
C1335 CSoutput.n259 gnd 0.547738f
C1336 CSoutput.n261 gnd 0.730317f
C1337 CSoutput.n263 gnd 1.96624f
C1338 CSoutput.n264 gnd 4.28278f
C1339 CSoutput.t73 gnd 0.051497f
C1340 CSoutput.t131 gnd 0.051497f
C1341 CSoutput.n265 gnd 0.398705f
C1342 CSoutput.t104 gnd 0.051497f
C1343 CSoutput.t141 gnd 0.051497f
C1344 CSoutput.n266 gnd 0.397994f
C1345 CSoutput.n267 gnd 0.403963f
C1346 CSoutput.t86 gnd 0.051497f
C1347 CSoutput.t125 gnd 0.051497f
C1348 CSoutput.n268 gnd 0.397994f
C1349 CSoutput.n269 gnd 0.199056f
C1350 CSoutput.t98 gnd 0.051497f
C1351 CSoutput.t139 gnd 0.051497f
C1352 CSoutput.n270 gnd 0.397994f
C1353 CSoutput.n271 gnd 0.199056f
C1354 CSoutput.t121 gnd 0.051497f
C1355 CSoutput.t77 gnd 0.051497f
C1356 CSoutput.n272 gnd 0.397994f
C1357 CSoutput.n273 gnd 0.199056f
C1358 CSoutput.t93 gnd 0.051497f
C1359 CSoutput.t79 gnd 0.051497f
C1360 CSoutput.n274 gnd 0.397994f
C1361 CSoutput.n275 gnd 0.365023f
C1362 CSoutput.t105 gnd 0.051497f
C1363 CSoutput.t106 gnd 0.051497f
C1364 CSoutput.n276 gnd 0.398705f
C1365 CSoutput.t117 gnd 0.051497f
C1366 CSoutput.t75 gnd 0.051497f
C1367 CSoutput.n277 gnd 0.397994f
C1368 CSoutput.n278 gnd 0.403963f
C1369 CSoutput.t102 gnd 0.051497f
C1370 CSoutput.t116 gnd 0.051497f
C1371 CSoutput.n279 gnd 0.397994f
C1372 CSoutput.n280 gnd 0.199056f
C1373 CSoutput.t143 gnd 0.051497f
C1374 CSoutput.t90 gnd 0.051497f
C1375 CSoutput.n281 gnd 0.397994f
C1376 CSoutput.n282 gnd 0.199056f
C1377 CSoutput.t91 gnd 0.051497f
C1378 CSoutput.t133 gnd 0.051497f
C1379 CSoutput.n283 gnd 0.397994f
C1380 CSoutput.n284 gnd 0.199056f
C1381 CSoutput.t88 gnd 0.051497f
C1382 CSoutput.t89 gnd 0.051497f
C1383 CSoutput.n285 gnd 0.397994f
C1384 CSoutput.n286 gnd 0.296842f
C1385 CSoutput.n287 gnd 0.374317f
C1386 CSoutput.t110 gnd 0.051497f
C1387 CSoutput.t111 gnd 0.051497f
C1388 CSoutput.n288 gnd 0.398705f
C1389 CSoutput.t129 gnd 0.051497f
C1390 CSoutput.t83 gnd 0.051497f
C1391 CSoutput.n289 gnd 0.397994f
C1392 CSoutput.n290 gnd 0.403963f
C1393 CSoutput.t109 gnd 0.051497f
C1394 CSoutput.t124 gnd 0.051497f
C1395 CSoutput.n291 gnd 0.397994f
C1396 CSoutput.n292 gnd 0.199056f
C1397 CSoutput.t81 gnd 0.051497f
C1398 CSoutput.t99 gnd 0.051497f
C1399 CSoutput.n293 gnd 0.397994f
C1400 CSoutput.n294 gnd 0.199056f
C1401 CSoutput.t101 gnd 0.051497f
C1402 CSoutput.t140 gnd 0.051497f
C1403 CSoutput.n295 gnd 0.397994f
C1404 CSoutput.n296 gnd 0.199056f
C1405 CSoutput.t95 gnd 0.051497f
C1406 CSoutput.t96 gnd 0.051497f
C1407 CSoutput.n297 gnd 0.397992f
C1408 CSoutput.n298 gnd 0.296844f
C1409 CSoutput.n299 gnd 0.41839f
C1410 CSoutput.n300 gnd 10.8432f
C1411 CSoutput.t63 gnd 0.04506f
C1412 CSoutput.t10 gnd 0.04506f
C1413 CSoutput.n301 gnd 0.399495f
C1414 CSoutput.t50 gnd 0.04506f
C1415 CSoutput.t0 gnd 0.04506f
C1416 CSoutput.n302 gnd 0.398163f
C1417 CSoutput.n303 gnd 0.371013f
C1418 CSoutput.t34 gnd 0.04506f
C1419 CSoutput.t65 gnd 0.04506f
C1420 CSoutput.n304 gnd 0.398163f
C1421 CSoutput.n305 gnd 0.182892f
C1422 CSoutput.t19 gnd 0.04506f
C1423 CSoutput.t32 gnd 0.04506f
C1424 CSoutput.n306 gnd 0.398163f
C1425 CSoutput.n307 gnd 0.182892f
C1426 CSoutput.t4 gnd 0.04506f
C1427 CSoutput.t40 gnd 0.04506f
C1428 CSoutput.n308 gnd 0.398163f
C1429 CSoutput.n309 gnd 0.182892f
C1430 CSoutput.t53 gnd 0.04506f
C1431 CSoutput.t24 gnd 0.04506f
C1432 CSoutput.n310 gnd 0.398163f
C1433 CSoutput.n311 gnd 0.337334f
C1434 CSoutput.t30 gnd 0.04506f
C1435 CSoutput.t13 gnd 0.04506f
C1436 CSoutput.n312 gnd 0.399495f
C1437 CSoutput.t18 gnd 0.04506f
C1438 CSoutput.t31 gnd 0.04506f
C1439 CSoutput.n313 gnd 0.398163f
C1440 CSoutput.n314 gnd 0.371013f
C1441 CSoutput.t14 gnd 0.04506f
C1442 CSoutput.t20 gnd 0.04506f
C1443 CSoutput.n315 gnd 0.398163f
C1444 CSoutput.n316 gnd 0.182892f
C1445 CSoutput.t33 gnd 0.04506f
C1446 CSoutput.t11 gnd 0.04506f
C1447 CSoutput.n317 gnd 0.398163f
C1448 CSoutput.n318 gnd 0.182892f
C1449 CSoutput.t21 gnd 0.04506f
C1450 CSoutput.t7 gnd 0.04506f
C1451 CSoutput.n319 gnd 0.398163f
C1452 CSoutput.n320 gnd 0.182892f
C1453 CSoutput.t12 gnd 0.04506f
C1454 CSoutput.t22 gnd 0.04506f
C1455 CSoutput.n321 gnd 0.398163f
C1456 CSoutput.n322 gnd 0.277669f
C1457 CSoutput.n323 gnd 0.350227f
C1458 CSoutput.t8 gnd 0.04506f
C1459 CSoutput.t69 gnd 0.04506f
C1460 CSoutput.n324 gnd 0.399495f
C1461 CSoutput.t59 gnd 0.04506f
C1462 CSoutput.t15 gnd 0.04506f
C1463 CSoutput.n325 gnd 0.398163f
C1464 CSoutput.n326 gnd 0.371013f
C1465 CSoutput.t1 gnd 0.04506f
C1466 CSoutput.t67 gnd 0.04506f
C1467 CSoutput.n327 gnd 0.398163f
C1468 CSoutput.n328 gnd 0.182892f
C1469 CSoutput.t26 gnd 0.04506f
C1470 CSoutput.t35 gnd 0.04506f
C1471 CSoutput.n329 gnd 0.398163f
C1472 CSoutput.n330 gnd 0.182892f
C1473 CSoutput.t70 gnd 0.04506f
C1474 CSoutput.t60 gnd 0.04506f
C1475 CSoutput.n331 gnd 0.398163f
C1476 CSoutput.n332 gnd 0.182892f
C1477 CSoutput.t44 gnd 0.04506f
C1478 CSoutput.t2 gnd 0.04506f
C1479 CSoutput.n333 gnd 0.398163f
C1480 CSoutput.n334 gnd 0.277669f
C1481 CSoutput.n335 gnd 0.376089f
C1482 CSoutput.n336 gnd 11.4074f
C1483 CSoutput.t41 gnd 0.04506f
C1484 CSoutput.t5 gnd 0.04506f
C1485 CSoutput.n337 gnd 0.399495f
C1486 CSoutput.t25 gnd 0.04506f
C1487 CSoutput.t66 gnd 0.04506f
C1488 CSoutput.n338 gnd 0.398163f
C1489 CSoutput.n339 gnd 0.371013f
C1490 CSoutput.t6 gnd 0.04506f
C1491 CSoutput.t55 gnd 0.04506f
C1492 CSoutput.n340 gnd 0.398163f
C1493 CSoutput.n341 gnd 0.182892f
C1494 CSoutput.t54 gnd 0.04506f
C1495 CSoutput.t43 gnd 0.04506f
C1496 CSoutput.n342 gnd 0.398163f
C1497 CSoutput.n343 gnd 0.182892f
C1498 CSoutput.t56 gnd 0.04506f
C1499 CSoutput.t27 gnd 0.04506f
C1500 CSoutput.n344 gnd 0.398163f
C1501 CSoutput.n345 gnd 0.182892f
C1502 CSoutput.t49 gnd 0.04506f
C1503 CSoutput.t61 gnd 0.04506f
C1504 CSoutput.n346 gnd 0.398163f
C1505 CSoutput.n347 gnd 0.337334f
C1506 CSoutput.t28 gnd 0.04506f
C1507 CSoutput.t45 gnd 0.04506f
C1508 CSoutput.n348 gnd 0.399495f
C1509 CSoutput.t46 gnd 0.04506f
C1510 CSoutput.t36 gnd 0.04506f
C1511 CSoutput.n349 gnd 0.398163f
C1512 CSoutput.n350 gnd 0.371013f
C1513 CSoutput.t37 gnd 0.04506f
C1514 CSoutput.t29 gnd 0.04506f
C1515 CSoutput.n351 gnd 0.398163f
C1516 CSoutput.n352 gnd 0.182892f
C1517 CSoutput.t23 gnd 0.04506f
C1518 CSoutput.t16 gnd 0.04506f
C1519 CSoutput.n353 gnd 0.398163f
C1520 CSoutput.n354 gnd 0.182892f
C1521 CSoutput.t17 gnd 0.04506f
C1522 CSoutput.t38 gnd 0.04506f
C1523 CSoutput.n355 gnd 0.398163f
C1524 CSoutput.n356 gnd 0.182892f
C1525 CSoutput.t39 gnd 0.04506f
C1526 CSoutput.t3 gnd 0.04506f
C1527 CSoutput.n357 gnd 0.398163f
C1528 CSoutput.n358 gnd 0.277669f
C1529 CSoutput.n359 gnd 0.350227f
C1530 CSoutput.t57 gnd 0.04506f
C1531 CSoutput.t68 gnd 0.04506f
C1532 CSoutput.n360 gnd 0.399495f
C1533 CSoutput.t71 gnd 0.04506f
C1534 CSoutput.t48 gnd 0.04506f
C1535 CSoutput.n361 gnd 0.398163f
C1536 CSoutput.n362 gnd 0.371013f
C1537 CSoutput.t52 gnd 0.04506f
C1538 CSoutput.t62 gnd 0.04506f
C1539 CSoutput.n363 gnd 0.398163f
C1540 CSoutput.n364 gnd 0.182892f
C1541 CSoutput.t9 gnd 0.04506f
C1542 CSoutput.t42 gnd 0.04506f
C1543 CSoutput.n365 gnd 0.398163f
C1544 CSoutput.n366 gnd 0.182892f
C1545 CSoutput.t47 gnd 0.04506f
C1546 CSoutput.t58 gnd 0.04506f
C1547 CSoutput.n367 gnd 0.398163f
C1548 CSoutput.n368 gnd 0.182892f
C1549 CSoutput.t64 gnd 0.04506f
C1550 CSoutput.t51 gnd 0.04506f
C1551 CSoutput.n369 gnd 0.398163f
C1552 CSoutput.n370 gnd 0.277669f
C1553 CSoutput.n371 gnd 0.376089f
C1554 CSoutput.n372 gnd 6.47972f
C1555 CSoutput.n373 gnd 12.6361f
C1556 a_n6308_8799.n0 gnd 0.177227f
C1557 a_n6308_8799.n1 gnd 0.207544f
C1558 a_n6308_8799.n2 gnd 0.207544f
C1559 a_n6308_8799.n3 gnd 0.207544f
C1560 a_n6308_8799.n4 gnd 0.177227f
C1561 a_n6308_8799.n5 gnd 0.207544f
C1562 a_n6308_8799.n6 gnd 0.207544f
C1563 a_n6308_8799.n7 gnd 0.207544f
C1564 a_n6308_8799.n8 gnd 0.342341f
C1565 a_n6308_8799.n9 gnd 0.207544f
C1566 a_n6308_8799.n10 gnd 0.207544f
C1567 a_n6308_8799.n11 gnd 0.207544f
C1568 a_n6308_8799.n12 gnd 0.207544f
C1569 a_n6308_8799.n13 gnd 0.207544f
C1570 a_n6308_8799.n14 gnd 0.177227f
C1571 a_n6308_8799.n15 gnd 0.207544f
C1572 a_n6308_8799.n16 gnd 0.207544f
C1573 a_n6308_8799.n17 gnd 0.207544f
C1574 a_n6308_8799.n18 gnd 0.177227f
C1575 a_n6308_8799.n19 gnd 0.207544f
C1576 a_n6308_8799.n20 gnd 0.207544f
C1577 a_n6308_8799.n21 gnd 0.207544f
C1578 a_n6308_8799.n22 gnd 0.342341f
C1579 a_n6308_8799.n23 gnd 0.207544f
C1580 a_n6308_8799.n24 gnd 4.02437f
C1581 a_n6308_8799.n25 gnd 2.7877f
C1582 a_n6308_8799.n26 gnd 0.362808f
C1583 a_n6308_8799.n27 gnd 3.04066f
C1584 a_n6308_8799.n28 gnd 0.362807f
C1585 a_n6308_8799.n29 gnd 0.855106f
C1586 a_n6308_8799.n30 gnd 0.250989f
C1587 a_n6308_8799.n32 gnd 0.00773f
C1588 a_n6308_8799.n33 gnd 0.011684f
C1589 a_n6308_8799.n34 gnd 0.008035f
C1590 a_n6308_8799.n36 gnd 4.01e-19
C1591 a_n6308_8799.n37 gnd 0.008328f
C1592 a_n6308_8799.n38 gnd 0.262565f
C1593 a_n6308_8799.n39 gnd 0.250989f
C1594 a_n6308_8799.n41 gnd 0.00773f
C1595 a_n6308_8799.n42 gnd 0.011684f
C1596 a_n6308_8799.n43 gnd 0.008035f
C1597 a_n6308_8799.n45 gnd 4.01e-19
C1598 a_n6308_8799.n46 gnd 0.008328f
C1599 a_n6308_8799.n47 gnd 0.262565f
C1600 a_n6308_8799.n48 gnd 0.250989f
C1601 a_n6308_8799.n50 gnd 0.00773f
C1602 a_n6308_8799.n51 gnd 0.011684f
C1603 a_n6308_8799.n52 gnd 0.008035f
C1604 a_n6308_8799.n54 gnd 4.01e-19
C1605 a_n6308_8799.n55 gnd 0.008328f
C1606 a_n6308_8799.n56 gnd 0.262565f
C1607 a_n6308_8799.n57 gnd 0.008328f
C1608 a_n6308_8799.n58 gnd 0.262565f
C1609 a_n6308_8799.n59 gnd 4.01e-19
C1610 a_n6308_8799.n61 gnd 0.008035f
C1611 a_n6308_8799.n62 gnd 0.011684f
C1612 a_n6308_8799.n63 gnd 0.00773f
C1613 a_n6308_8799.n65 gnd 0.250989f
C1614 a_n6308_8799.n66 gnd 0.008328f
C1615 a_n6308_8799.n67 gnd 0.262565f
C1616 a_n6308_8799.n68 gnd 4.01e-19
C1617 a_n6308_8799.n70 gnd 0.008035f
C1618 a_n6308_8799.n71 gnd 0.011684f
C1619 a_n6308_8799.n72 gnd 0.00773f
C1620 a_n6308_8799.n74 gnd 0.250989f
C1621 a_n6308_8799.n75 gnd 0.008328f
C1622 a_n6308_8799.n76 gnd 0.262565f
C1623 a_n6308_8799.n77 gnd 4.01e-19
C1624 a_n6308_8799.n79 gnd 0.008035f
C1625 a_n6308_8799.n80 gnd 0.011684f
C1626 a_n6308_8799.n81 gnd 0.00773f
C1627 a_n6308_8799.n83 gnd 0.250989f
C1628 a_n6308_8799.t32 gnd 0.143955f
C1629 a_n6308_8799.t5 gnd 0.143955f
C1630 a_n6308_8799.t8 gnd 0.143955f
C1631 a_n6308_8799.n84 gnd 1.13539f
C1632 a_n6308_8799.t7 gnd 0.143955f
C1633 a_n6308_8799.t29 gnd 0.143955f
C1634 a_n6308_8799.n85 gnd 1.13352f
C1635 a_n6308_8799.t21 gnd 0.143955f
C1636 a_n6308_8799.t22 gnd 0.143955f
C1637 a_n6308_8799.n86 gnd 1.13352f
C1638 a_n6308_8799.t9 gnd 0.111965f
C1639 a_n6308_8799.t11 gnd 0.111965f
C1640 a_n6308_8799.n87 gnd 0.992279f
C1641 a_n6308_8799.t15 gnd 0.111965f
C1642 a_n6308_8799.t34 gnd 0.111965f
C1643 a_n6308_8799.n88 gnd 0.989362f
C1644 a_n6308_8799.n89 gnd 0.877314f
C1645 a_n6308_8799.t26 gnd 0.111965f
C1646 a_n6308_8799.t3 gnd 0.111965f
C1647 a_n6308_8799.n90 gnd 0.989362f
C1648 a_n6308_8799.t27 gnd 0.111965f
C1649 a_n6308_8799.t35 gnd 0.111965f
C1650 a_n6308_8799.n91 gnd 0.992278f
C1651 a_n6308_8799.t28 gnd 0.111965f
C1652 a_n6308_8799.t14 gnd 0.111965f
C1653 a_n6308_8799.n92 gnd 0.989361f
C1654 a_n6308_8799.n93 gnd 0.877316f
C1655 a_n6308_8799.t33 gnd 0.111965f
C1656 a_n6308_8799.t30 gnd 0.111965f
C1657 a_n6308_8799.n94 gnd 0.989361f
C1658 a_n6308_8799.t12 gnd 0.111965f
C1659 a_n6308_8799.t31 gnd 0.111965f
C1660 a_n6308_8799.n95 gnd 0.992278f
C1661 a_n6308_8799.t24 gnd 0.111965f
C1662 a_n6308_8799.t17 gnd 0.111965f
C1663 a_n6308_8799.n96 gnd 0.989361f
C1664 a_n6308_8799.n97 gnd 0.877316f
C1665 a_n6308_8799.t23 gnd 0.111965f
C1666 a_n6308_8799.t4 gnd 0.111965f
C1667 a_n6308_8799.n98 gnd 0.989361f
C1668 a_n6308_8799.t18 gnd 0.111965f
C1669 a_n6308_8799.t0 gnd 0.111965f
C1670 a_n6308_8799.n99 gnd 0.989362f
C1671 a_n6308_8799.n100 gnd 3.0863f
C1672 a_n6308_8799.t19 gnd 0.111965f
C1673 a_n6308_8799.t25 gnd 0.111965f
C1674 a_n6308_8799.n101 gnd 0.989362f
C1675 a_n6308_8799.n102 gnd 0.431963f
C1676 a_n6308_8799.t10 gnd 0.111965f
C1677 a_n6308_8799.t13 gnd 0.111965f
C1678 a_n6308_8799.n103 gnd 0.989362f
C1679 a_n6308_8799.t95 gnd 0.596904f
C1680 a_n6308_8799.n104 gnd 0.270153f
C1681 a_n6308_8799.t43 gnd 0.596904f
C1682 a_n6308_8799.t44 gnd 0.596904f
C1683 a_n6308_8799.n105 gnd 0.26131f
C1684 a_n6308_8799.t57 gnd 0.596904f
C1685 a_n6308_8799.n106 gnd 0.272683f
C1686 a_n6308_8799.t72 gnd 0.596904f
C1687 a_n6308_8799.t85 gnd 0.596904f
C1688 a_n6308_8799.n107 gnd 0.266109f
C1689 a_n6308_8799.t60 gnd 0.610933f
C1690 a_n6308_8799.t61 gnd 0.596904f
C1691 a_n6308_8799.n108 gnd 0.272248f
C1692 a_n6308_8799.n109 gnd 0.248822f
C1693 a_n6308_8799.t37 gnd 0.596904f
C1694 a_n6308_8799.n110 gnd 0.270035f
C1695 a_n6308_8799.n111 gnd 0.270167f
C1696 a_n6308_8799.t97 gnd 0.596904f
C1697 a_n6308_8799.n112 gnd 0.266429f
C1698 a_n6308_8799.t56 gnd 0.596904f
C1699 a_n6308_8799.n113 gnd 0.266679f
C1700 a_n6308_8799.n114 gnd 0.272249f
C1701 a_n6308_8799.t42 gnd 0.607741f
C1702 a_n6308_8799.t101 gnd 0.596904f
C1703 a_n6308_8799.n115 gnd 0.270153f
C1704 a_n6308_8799.t49 gnd 0.596904f
C1705 a_n6308_8799.t53 gnd 0.596904f
C1706 a_n6308_8799.n116 gnd 0.26131f
C1707 a_n6308_8799.t65 gnd 0.596904f
C1708 a_n6308_8799.n117 gnd 0.272683f
C1709 a_n6308_8799.t79 gnd 0.596904f
C1710 a_n6308_8799.t92 gnd 0.596904f
C1711 a_n6308_8799.n118 gnd 0.266109f
C1712 a_n6308_8799.t66 gnd 0.610933f
C1713 a_n6308_8799.t67 gnd 0.596904f
C1714 a_n6308_8799.n119 gnd 0.272248f
C1715 a_n6308_8799.n120 gnd 0.248822f
C1716 a_n6308_8799.t45 gnd 0.596904f
C1717 a_n6308_8799.n121 gnd 0.270035f
C1718 a_n6308_8799.n122 gnd 0.270167f
C1719 a_n6308_8799.t105 gnd 0.596904f
C1720 a_n6308_8799.n123 gnd 0.266429f
C1721 a_n6308_8799.t64 gnd 0.596904f
C1722 a_n6308_8799.n124 gnd 0.266679f
C1723 a_n6308_8799.n125 gnd 0.272249f
C1724 a_n6308_8799.t51 gnd 0.607741f
C1725 a_n6308_8799.n126 gnd 0.896117f
C1726 a_n6308_8799.t76 gnd 0.596904f
C1727 a_n6308_8799.n127 gnd 0.270153f
C1728 a_n6308_8799.t47 gnd 0.596904f
C1729 a_n6308_8799.t94 gnd 0.596904f
C1730 a_n6308_8799.n128 gnd 0.26131f
C1731 a_n6308_8799.t41 gnd 0.596904f
C1732 a_n6308_8799.n129 gnd 0.272683f
C1733 a_n6308_8799.t82 gnd 0.596904f
C1734 a_n6308_8799.t103 gnd 0.596904f
C1735 a_n6308_8799.n130 gnd 0.266109f
C1736 a_n6308_8799.t99 gnd 0.610933f
C1737 a_n6308_8799.t87 gnd 0.596904f
C1738 a_n6308_8799.n131 gnd 0.272248f
C1739 a_n6308_8799.n132 gnd 0.248822f
C1740 a_n6308_8799.t71 gnd 0.596904f
C1741 a_n6308_8799.n133 gnd 0.270035f
C1742 a_n6308_8799.n134 gnd 0.270167f
C1743 a_n6308_8799.t52 gnd 0.596904f
C1744 a_n6308_8799.n135 gnd 0.266429f
C1745 a_n6308_8799.t59 gnd 0.596904f
C1746 a_n6308_8799.n136 gnd 0.266679f
C1747 a_n6308_8799.n137 gnd 0.272249f
C1748 a_n6308_8799.t107 gnd 0.607741f
C1749 a_n6308_8799.n138 gnd 1.53643f
C1750 a_n6308_8799.t69 gnd 0.607741f
C1751 a_n6308_8799.t68 gnd 0.596904f
C1752 a_n6308_8799.t50 gnd 0.596904f
C1753 a_n6308_8799.t96 gnd 0.596904f
C1754 a_n6308_8799.n139 gnd 0.266679f
C1755 a_n6308_8799.t70 gnd 0.596904f
C1756 a_n6308_8799.t55 gnd 0.596904f
C1757 a_n6308_8799.t98 gnd 0.596904f
C1758 a_n6308_8799.n140 gnd 0.270167f
C1759 a_n6308_8799.t80 gnd 0.596904f
C1760 a_n6308_8799.t78 gnd 0.596904f
C1761 a_n6308_8799.t39 gnd 0.596904f
C1762 a_n6308_8799.n141 gnd 0.266109f
C1763 a_n6308_8799.t83 gnd 0.610933f
C1764 a_n6308_8799.t84 gnd 0.596904f
C1765 a_n6308_8799.n142 gnd 0.272248f
C1766 a_n6308_8799.n143 gnd 0.248822f
C1767 a_n6308_8799.n144 gnd 0.270035f
C1768 a_n6308_8799.n145 gnd 0.272683f
C1769 a_n6308_8799.n146 gnd 0.266429f
C1770 a_n6308_8799.n147 gnd 0.26131f
C1771 a_n6308_8799.n148 gnd 0.270153f
C1772 a_n6308_8799.n149 gnd 0.272249f
C1773 a_n6308_8799.t74 gnd 0.607741f
C1774 a_n6308_8799.t73 gnd 0.596904f
C1775 a_n6308_8799.t62 gnd 0.596904f
C1776 a_n6308_8799.t104 gnd 0.596904f
C1777 a_n6308_8799.n150 gnd 0.266679f
C1778 a_n6308_8799.t77 gnd 0.596904f
C1779 a_n6308_8799.t63 gnd 0.596904f
C1780 a_n6308_8799.t36 gnd 0.596904f
C1781 a_n6308_8799.n151 gnd 0.270167f
C1782 a_n6308_8799.t89 gnd 0.596904f
C1783 a_n6308_8799.t88 gnd 0.596904f
C1784 a_n6308_8799.t46 gnd 0.596904f
C1785 a_n6308_8799.n152 gnd 0.266109f
C1786 a_n6308_8799.t90 gnd 0.610933f
C1787 a_n6308_8799.t91 gnd 0.596904f
C1788 a_n6308_8799.n153 gnd 0.272248f
C1789 a_n6308_8799.n154 gnd 0.248822f
C1790 a_n6308_8799.n155 gnd 0.270035f
C1791 a_n6308_8799.n156 gnd 0.272683f
C1792 a_n6308_8799.n157 gnd 0.266429f
C1793 a_n6308_8799.n158 gnd 0.26131f
C1794 a_n6308_8799.n159 gnd 0.270153f
C1795 a_n6308_8799.n160 gnd 0.272249f
C1796 a_n6308_8799.n161 gnd 0.896117f
C1797 a_n6308_8799.t106 gnd 0.607741f
C1798 a_n6308_8799.t48 gnd 0.596904f
C1799 a_n6308_8799.t75 gnd 0.596904f
C1800 a_n6308_8799.t38 gnd 0.596904f
C1801 a_n6308_8799.n162 gnd 0.266679f
C1802 a_n6308_8799.t93 gnd 0.596904f
C1803 a_n6308_8799.t54 gnd 0.596904f
C1804 a_n6308_8799.t81 gnd 0.596904f
C1805 a_n6308_8799.n163 gnd 0.270167f
C1806 a_n6308_8799.t40 gnd 0.596904f
C1807 a_n6308_8799.t58 gnd 0.596904f
C1808 a_n6308_8799.t102 gnd 0.596904f
C1809 a_n6308_8799.n164 gnd 0.266109f
C1810 a_n6308_8799.t100 gnd 0.610933f
C1811 a_n6308_8799.t86 gnd 0.596904f
C1812 a_n6308_8799.n165 gnd 0.272248f
C1813 a_n6308_8799.n166 gnd 0.248822f
C1814 a_n6308_8799.n167 gnd 0.270035f
C1815 a_n6308_8799.n168 gnd 0.272683f
C1816 a_n6308_8799.n169 gnd 0.266429f
C1817 a_n6308_8799.n170 gnd 0.26131f
C1818 a_n6308_8799.n171 gnd 0.270153f
C1819 a_n6308_8799.n172 gnd 0.272249f
C1820 a_n6308_8799.n173 gnd 1.08397f
C1821 a_n6308_8799.n174 gnd 12.191501f
C1822 a_n6308_8799.n175 gnd 4.36847f
C1823 a_n6308_8799.n176 gnd 5.66783f
C1824 a_n6308_8799.t16 gnd 0.143955f
C1825 a_n6308_8799.t20 gnd 0.143955f
C1826 a_n6308_8799.n177 gnd 1.13352f
C1827 a_n6308_8799.t2 gnd 0.143955f
C1828 a_n6308_8799.t6 gnd 0.143955f
C1829 a_n6308_8799.n178 gnd 1.13352f
C1830 a_n6308_8799.n179 gnd 1.1354f
C1831 a_n6308_8799.t1 gnd 0.143955f
C1832 vdd.t221 gnd 0.035939f
C1833 vdd.t185 gnd 0.035939f
C1834 vdd.n0 gnd 0.283454f
C1835 vdd.t160 gnd 0.035939f
C1836 vdd.t227 gnd 0.035939f
C1837 vdd.n1 gnd 0.282986f
C1838 vdd.n2 gnd 0.260967f
C1839 vdd.t197 gnd 0.035939f
C1840 vdd.t145 gnd 0.035939f
C1841 vdd.n3 gnd 0.282986f
C1842 vdd.n4 gnd 0.131981f
C1843 vdd.t164 gnd 0.035939f
C1844 vdd.t18 gnd 0.035939f
C1845 vdd.n5 gnd 0.282986f
C1846 vdd.n6 gnd 0.12384f
C1847 vdd.t162 gnd 0.035939f
C1848 vdd.t199 gnd 0.035939f
C1849 vdd.n7 gnd 0.283454f
C1850 vdd.t131 gnd 0.035939f
C1851 vdd.t166 gnd 0.035939f
C1852 vdd.n8 gnd 0.282986f
C1853 vdd.n9 gnd 0.260967f
C1854 vdd.t171 gnd 0.035939f
C1855 vdd.t14 gnd 0.035939f
C1856 vdd.n10 gnd 0.282986f
C1857 vdd.n11 gnd 0.131981f
C1858 vdd.t201 gnd 0.035939f
C1859 vdd.t173 gnd 0.035939f
C1860 vdd.n12 gnd 0.282986f
C1861 vdd.n13 gnd 0.12384f
C1862 vdd.n14 gnd 0.087552f
C1863 vdd.t189 gnd 0.019966f
C1864 vdd.t158 gnd 0.019966f
C1865 vdd.n15 gnd 0.183778f
C1866 vdd.t53 gnd 0.019966f
C1867 vdd.t11 gnd 0.019966f
C1868 vdd.n16 gnd 0.18324f
C1869 vdd.n17 gnd 0.318895f
C1870 vdd.t8 gnd 0.019966f
C1871 vdd.t52 gnd 0.019966f
C1872 vdd.n18 gnd 0.18324f
C1873 vdd.n19 gnd 0.131931f
C1874 vdd.t157 gnd 0.019966f
C1875 vdd.t12 gnd 0.019966f
C1876 vdd.n20 gnd 0.183778f
C1877 vdd.t1 gnd 0.019966f
C1878 vdd.t50 gnd 0.019966f
C1879 vdd.n21 gnd 0.18324f
C1880 vdd.n22 gnd 0.318895f
C1881 vdd.t2 gnd 0.019966f
C1882 vdd.t135 gnd 0.019966f
C1883 vdd.n23 gnd 0.18324f
C1884 vdd.n24 gnd 0.131931f
C1885 vdd.t10 gnd 0.019966f
C1886 vdd.t156 gnd 0.019966f
C1887 vdd.n25 gnd 0.18324f
C1888 vdd.t51 gnd 0.019966f
C1889 vdd.t0 gnd 0.019966f
C1890 vdd.n26 gnd 0.18324f
C1891 vdd.n27 gnd 20.061699f
C1892 vdd.n28 gnd 7.54208f
C1893 vdd.n29 gnd 0.005446f
C1894 vdd.n30 gnd 0.005053f
C1895 vdd.n31 gnd 0.002795f
C1896 vdd.n32 gnd 0.006418f
C1897 vdd.n33 gnd 0.002715f
C1898 vdd.n34 gnd 0.002875f
C1899 vdd.n35 gnd 0.005053f
C1900 vdd.n36 gnd 0.002715f
C1901 vdd.n37 gnd 0.006418f
C1902 vdd.n38 gnd 0.002875f
C1903 vdd.n39 gnd 0.005053f
C1904 vdd.n40 gnd 0.002715f
C1905 vdd.n41 gnd 0.004814f
C1906 vdd.n42 gnd 0.004828f
C1907 vdd.t175 gnd 0.013789f
C1908 vdd.n43 gnd 0.03068f
C1909 vdd.n44 gnd 0.159666f
C1910 vdd.n45 gnd 0.002715f
C1911 vdd.n46 gnd 0.002875f
C1912 vdd.n47 gnd 0.006418f
C1913 vdd.n48 gnd 0.006418f
C1914 vdd.n49 gnd 0.002875f
C1915 vdd.n50 gnd 0.002715f
C1916 vdd.n51 gnd 0.005053f
C1917 vdd.n52 gnd 0.005053f
C1918 vdd.n53 gnd 0.002715f
C1919 vdd.n54 gnd 0.002875f
C1920 vdd.n55 gnd 0.006418f
C1921 vdd.n56 gnd 0.006418f
C1922 vdd.n57 gnd 0.002875f
C1923 vdd.n58 gnd 0.002715f
C1924 vdd.n59 gnd 0.005053f
C1925 vdd.n60 gnd 0.005053f
C1926 vdd.n61 gnd 0.002715f
C1927 vdd.n62 gnd 0.002875f
C1928 vdd.n63 gnd 0.006418f
C1929 vdd.n64 gnd 0.006418f
C1930 vdd.n65 gnd 0.015174f
C1931 vdd.n66 gnd 0.002795f
C1932 vdd.n67 gnd 0.002715f
C1933 vdd.n68 gnd 0.013061f
C1934 vdd.n69 gnd 0.009118f
C1935 vdd.t133 gnd 0.031946f
C1936 vdd.t29 gnd 0.031946f
C1937 vdd.n70 gnd 0.219551f
C1938 vdd.n71 gnd 0.172644f
C1939 vdd.t148 gnd 0.031946f
C1940 vdd.t183 gnd 0.031946f
C1941 vdd.n72 gnd 0.219551f
C1942 vdd.n73 gnd 0.139322f
C1943 vdd.t36 gnd 0.031946f
C1944 vdd.t188 gnd 0.031946f
C1945 vdd.n74 gnd 0.219551f
C1946 vdd.n75 gnd 0.139322f
C1947 vdd.t24 gnd 0.031946f
C1948 vdd.t139 gnd 0.031946f
C1949 vdd.n76 gnd 0.219551f
C1950 vdd.n77 gnd 0.139322f
C1951 vdd.t180 gnd 0.031946f
C1952 vdd.t217 gnd 0.031946f
C1953 vdd.n78 gnd 0.219551f
C1954 vdd.n79 gnd 0.139322f
C1955 vdd.n80 gnd 0.005446f
C1956 vdd.n81 gnd 0.005053f
C1957 vdd.n82 gnd 0.002795f
C1958 vdd.n83 gnd 0.006418f
C1959 vdd.n84 gnd 0.002715f
C1960 vdd.n85 gnd 0.002875f
C1961 vdd.n86 gnd 0.005053f
C1962 vdd.n87 gnd 0.002715f
C1963 vdd.n88 gnd 0.006418f
C1964 vdd.n89 gnd 0.002875f
C1965 vdd.n90 gnd 0.005053f
C1966 vdd.n91 gnd 0.002715f
C1967 vdd.n92 gnd 0.004814f
C1968 vdd.n93 gnd 0.004828f
C1969 vdd.t230 gnd 0.013789f
C1970 vdd.n94 gnd 0.03068f
C1971 vdd.n95 gnd 0.159666f
C1972 vdd.n96 gnd 0.002715f
C1973 vdd.n97 gnd 0.002875f
C1974 vdd.n98 gnd 0.006418f
C1975 vdd.n99 gnd 0.006418f
C1976 vdd.n100 gnd 0.002875f
C1977 vdd.n101 gnd 0.002715f
C1978 vdd.n102 gnd 0.005053f
C1979 vdd.n103 gnd 0.005053f
C1980 vdd.n104 gnd 0.002715f
C1981 vdd.n105 gnd 0.002875f
C1982 vdd.n106 gnd 0.006418f
C1983 vdd.n107 gnd 0.006418f
C1984 vdd.n108 gnd 0.002875f
C1985 vdd.n109 gnd 0.002715f
C1986 vdd.n110 gnd 0.005053f
C1987 vdd.n111 gnd 0.005053f
C1988 vdd.n112 gnd 0.002715f
C1989 vdd.n113 gnd 0.002875f
C1990 vdd.n114 gnd 0.006418f
C1991 vdd.n115 gnd 0.006418f
C1992 vdd.n116 gnd 0.015174f
C1993 vdd.n117 gnd 0.002795f
C1994 vdd.n118 gnd 0.002715f
C1995 vdd.n119 gnd 0.013061f
C1996 vdd.n120 gnd 0.008832f
C1997 vdd.n121 gnd 0.103657f
C1998 vdd.n122 gnd 0.005446f
C1999 vdd.n123 gnd 0.005053f
C2000 vdd.n124 gnd 0.002795f
C2001 vdd.n125 gnd 0.006418f
C2002 vdd.n126 gnd 0.002715f
C2003 vdd.n127 gnd 0.002875f
C2004 vdd.n128 gnd 0.005053f
C2005 vdd.n129 gnd 0.002715f
C2006 vdd.n130 gnd 0.006418f
C2007 vdd.n131 gnd 0.002875f
C2008 vdd.n132 gnd 0.005053f
C2009 vdd.n133 gnd 0.002715f
C2010 vdd.n134 gnd 0.004814f
C2011 vdd.n135 gnd 0.004828f
C2012 vdd.t27 gnd 0.013789f
C2013 vdd.n136 gnd 0.03068f
C2014 vdd.n137 gnd 0.159666f
C2015 vdd.n138 gnd 0.002715f
C2016 vdd.n139 gnd 0.002875f
C2017 vdd.n140 gnd 0.006418f
C2018 vdd.n141 gnd 0.006418f
C2019 vdd.n142 gnd 0.002875f
C2020 vdd.n143 gnd 0.002715f
C2021 vdd.n144 gnd 0.005053f
C2022 vdd.n145 gnd 0.005053f
C2023 vdd.n146 gnd 0.002715f
C2024 vdd.n147 gnd 0.002875f
C2025 vdd.n148 gnd 0.006418f
C2026 vdd.n149 gnd 0.006418f
C2027 vdd.n150 gnd 0.002875f
C2028 vdd.n151 gnd 0.002715f
C2029 vdd.n152 gnd 0.005053f
C2030 vdd.n153 gnd 0.005053f
C2031 vdd.n154 gnd 0.002715f
C2032 vdd.n155 gnd 0.002875f
C2033 vdd.n156 gnd 0.006418f
C2034 vdd.n157 gnd 0.006418f
C2035 vdd.n158 gnd 0.015174f
C2036 vdd.n159 gnd 0.002795f
C2037 vdd.n160 gnd 0.002715f
C2038 vdd.n161 gnd 0.013061f
C2039 vdd.n162 gnd 0.009118f
C2040 vdd.t210 gnd 0.031946f
C2041 vdd.t141 gnd 0.031946f
C2042 vdd.n163 gnd 0.219551f
C2043 vdd.n164 gnd 0.172644f
C2044 vdd.t177 gnd 0.031946f
C2045 vdd.t7 gnd 0.031946f
C2046 vdd.n165 gnd 0.219551f
C2047 vdd.n166 gnd 0.139322f
C2048 vdd.t142 gnd 0.031946f
C2049 vdd.t190 gnd 0.031946f
C2050 vdd.n167 gnd 0.219551f
C2051 vdd.n168 gnd 0.139322f
C2052 vdd.t193 gnd 0.031946f
C2053 vdd.t192 gnd 0.031946f
C2054 vdd.n169 gnd 0.219551f
C2055 vdd.n170 gnd 0.139322f
C2056 vdd.t204 gnd 0.031946f
C2057 vdd.t155 gnd 0.031946f
C2058 vdd.n171 gnd 0.219551f
C2059 vdd.n172 gnd 0.139322f
C2060 vdd.n173 gnd 0.005446f
C2061 vdd.n174 gnd 0.005053f
C2062 vdd.n175 gnd 0.002795f
C2063 vdd.n176 gnd 0.006418f
C2064 vdd.n177 gnd 0.002715f
C2065 vdd.n178 gnd 0.002875f
C2066 vdd.n179 gnd 0.005053f
C2067 vdd.n180 gnd 0.002715f
C2068 vdd.n181 gnd 0.006418f
C2069 vdd.n182 gnd 0.002875f
C2070 vdd.n183 gnd 0.005053f
C2071 vdd.n184 gnd 0.002715f
C2072 vdd.n185 gnd 0.004814f
C2073 vdd.n186 gnd 0.004828f
C2074 vdd.t153 gnd 0.013789f
C2075 vdd.n187 gnd 0.03068f
C2076 vdd.n188 gnd 0.159666f
C2077 vdd.n189 gnd 0.002715f
C2078 vdd.n190 gnd 0.002875f
C2079 vdd.n191 gnd 0.006418f
C2080 vdd.n192 gnd 0.006418f
C2081 vdd.n193 gnd 0.002875f
C2082 vdd.n194 gnd 0.002715f
C2083 vdd.n195 gnd 0.005053f
C2084 vdd.n196 gnd 0.005053f
C2085 vdd.n197 gnd 0.002715f
C2086 vdd.n198 gnd 0.002875f
C2087 vdd.n199 gnd 0.006418f
C2088 vdd.n200 gnd 0.006418f
C2089 vdd.n201 gnd 0.002875f
C2090 vdd.n202 gnd 0.002715f
C2091 vdd.n203 gnd 0.005053f
C2092 vdd.n204 gnd 0.005053f
C2093 vdd.n205 gnd 0.002715f
C2094 vdd.n206 gnd 0.002875f
C2095 vdd.n207 gnd 0.006418f
C2096 vdd.n208 gnd 0.006418f
C2097 vdd.n209 gnd 0.015174f
C2098 vdd.n210 gnd 0.002795f
C2099 vdd.n211 gnd 0.002715f
C2100 vdd.n212 gnd 0.013061f
C2101 vdd.n213 gnd 0.008832f
C2102 vdd.n214 gnd 0.061665f
C2103 vdd.n215 gnd 0.222196f
C2104 vdd.n216 gnd 0.005446f
C2105 vdd.n217 gnd 0.005053f
C2106 vdd.n218 gnd 0.002795f
C2107 vdd.n219 gnd 0.006418f
C2108 vdd.n220 gnd 0.002715f
C2109 vdd.n221 gnd 0.002875f
C2110 vdd.n222 gnd 0.005053f
C2111 vdd.n223 gnd 0.002715f
C2112 vdd.n224 gnd 0.006418f
C2113 vdd.n225 gnd 0.002875f
C2114 vdd.n226 gnd 0.005053f
C2115 vdd.n227 gnd 0.002715f
C2116 vdd.n228 gnd 0.004814f
C2117 vdd.n229 gnd 0.004828f
C2118 vdd.t22 gnd 0.013789f
C2119 vdd.n230 gnd 0.03068f
C2120 vdd.n231 gnd 0.159666f
C2121 vdd.n232 gnd 0.002715f
C2122 vdd.n233 gnd 0.002875f
C2123 vdd.n234 gnd 0.006418f
C2124 vdd.n235 gnd 0.006418f
C2125 vdd.n236 gnd 0.002875f
C2126 vdd.n237 gnd 0.002715f
C2127 vdd.n238 gnd 0.005053f
C2128 vdd.n239 gnd 0.005053f
C2129 vdd.n240 gnd 0.002715f
C2130 vdd.n241 gnd 0.002875f
C2131 vdd.n242 gnd 0.006418f
C2132 vdd.n243 gnd 0.006418f
C2133 vdd.n244 gnd 0.002875f
C2134 vdd.n245 gnd 0.002715f
C2135 vdd.n246 gnd 0.005053f
C2136 vdd.n247 gnd 0.005053f
C2137 vdd.n248 gnd 0.002715f
C2138 vdd.n249 gnd 0.002875f
C2139 vdd.n250 gnd 0.006418f
C2140 vdd.n251 gnd 0.006418f
C2141 vdd.n252 gnd 0.015174f
C2142 vdd.n253 gnd 0.002795f
C2143 vdd.n254 gnd 0.002715f
C2144 vdd.n255 gnd 0.013061f
C2145 vdd.n256 gnd 0.009118f
C2146 vdd.t20 gnd 0.031946f
C2147 vdd.t194 gnd 0.031946f
C2148 vdd.n257 gnd 0.219551f
C2149 vdd.n258 gnd 0.172644f
C2150 vdd.t228 gnd 0.031946f
C2151 vdd.t224 gnd 0.031946f
C2152 vdd.n259 gnd 0.219551f
C2153 vdd.n260 gnd 0.139322f
C2154 vdd.t37 gnd 0.031946f
C2155 vdd.t213 gnd 0.031946f
C2156 vdd.n261 gnd 0.219551f
C2157 vdd.n262 gnd 0.139322f
C2158 vdd.t186 gnd 0.031946f
C2159 vdd.t211 gnd 0.031946f
C2160 vdd.n263 gnd 0.219551f
C2161 vdd.n264 gnd 0.139322f
C2162 vdd.t150 gnd 0.031946f
C2163 vdd.t167 gnd 0.031946f
C2164 vdd.n265 gnd 0.219551f
C2165 vdd.n266 gnd 0.139322f
C2166 vdd.n267 gnd 0.005446f
C2167 vdd.n268 gnd 0.005053f
C2168 vdd.n269 gnd 0.002795f
C2169 vdd.n270 gnd 0.006418f
C2170 vdd.n271 gnd 0.002715f
C2171 vdd.n272 gnd 0.002875f
C2172 vdd.n273 gnd 0.005053f
C2173 vdd.n274 gnd 0.002715f
C2174 vdd.n275 gnd 0.006418f
C2175 vdd.n276 gnd 0.002875f
C2176 vdd.n277 gnd 0.005053f
C2177 vdd.n278 gnd 0.002715f
C2178 vdd.n279 gnd 0.004814f
C2179 vdd.n280 gnd 0.004828f
C2180 vdd.t223 gnd 0.013789f
C2181 vdd.n281 gnd 0.03068f
C2182 vdd.n282 gnd 0.159666f
C2183 vdd.n283 gnd 0.002715f
C2184 vdd.n284 gnd 0.002875f
C2185 vdd.n285 gnd 0.006418f
C2186 vdd.n286 gnd 0.006418f
C2187 vdd.n287 gnd 0.002875f
C2188 vdd.n288 gnd 0.002715f
C2189 vdd.n289 gnd 0.005053f
C2190 vdd.n290 gnd 0.005053f
C2191 vdd.n291 gnd 0.002715f
C2192 vdd.n292 gnd 0.002875f
C2193 vdd.n293 gnd 0.006418f
C2194 vdd.n294 gnd 0.006418f
C2195 vdd.n295 gnd 0.002875f
C2196 vdd.n296 gnd 0.002715f
C2197 vdd.n297 gnd 0.005053f
C2198 vdd.n298 gnd 0.005053f
C2199 vdd.n299 gnd 0.002715f
C2200 vdd.n300 gnd 0.002875f
C2201 vdd.n301 gnd 0.006418f
C2202 vdd.n302 gnd 0.006418f
C2203 vdd.n303 gnd 0.015174f
C2204 vdd.n304 gnd 0.002795f
C2205 vdd.n305 gnd 0.002715f
C2206 vdd.n306 gnd 0.013061f
C2207 vdd.n307 gnd 0.008832f
C2208 vdd.n308 gnd 0.061665f
C2209 vdd.n309 gnd 0.244201f
C2210 vdd.n310 gnd 0.009888f
C2211 vdd.n311 gnd 0.009888f
C2212 vdd.n312 gnd 0.007986f
C2213 vdd.n313 gnd 0.007986f
C2214 vdd.n314 gnd 0.009922f
C2215 vdd.n315 gnd 0.009922f
C2216 vdd.t35 gnd 0.507014f
C2217 vdd.n316 gnd 0.009922f
C2218 vdd.n317 gnd 0.009922f
C2219 vdd.n318 gnd 0.009922f
C2220 vdd.t23 gnd 0.507014f
C2221 vdd.n319 gnd 0.009922f
C2222 vdd.n320 gnd 0.009922f
C2223 vdd.n321 gnd 0.009922f
C2224 vdd.n322 gnd 0.009922f
C2225 vdd.n323 gnd 0.007986f
C2226 vdd.n324 gnd 0.009922f
C2227 vdd.n325 gnd 0.816292f
C2228 vdd.n326 gnd 0.009922f
C2229 vdd.n327 gnd 0.009922f
C2230 vdd.n328 gnd 0.009922f
C2231 vdd.n329 gnd 0.694609f
C2232 vdd.n330 gnd 0.009922f
C2233 vdd.n331 gnd 0.009922f
C2234 vdd.n332 gnd 0.009922f
C2235 vdd.n333 gnd 0.009922f
C2236 vdd.n334 gnd 0.009922f
C2237 vdd.n335 gnd 0.007986f
C2238 vdd.n336 gnd 0.009922f
C2239 vdd.t154 gnd 0.507014f
C2240 vdd.n337 gnd 0.009922f
C2241 vdd.n338 gnd 0.009922f
C2242 vdd.n339 gnd 0.009922f
C2243 vdd.n340 gnd 1.01403f
C2244 vdd.n341 gnd 0.009922f
C2245 vdd.n342 gnd 0.009922f
C2246 vdd.n343 gnd 0.009922f
C2247 vdd.n344 gnd 0.009922f
C2248 vdd.n345 gnd 0.009922f
C2249 vdd.n346 gnd 0.007986f
C2250 vdd.n347 gnd 0.009922f
C2251 vdd.n348 gnd 0.009922f
C2252 vdd.n349 gnd 0.009922f
C2253 vdd.n350 gnd 0.023383f
C2254 vdd.n351 gnd 2.33226f
C2255 vdd.n352 gnd 0.023749f
C2256 vdd.n353 gnd 0.009922f
C2257 vdd.n354 gnd 0.009922f
C2258 vdd.n356 gnd 0.009922f
C2259 vdd.n357 gnd 0.009922f
C2260 vdd.n358 gnd 0.007986f
C2261 vdd.n359 gnd 0.007986f
C2262 vdd.n360 gnd 0.009922f
C2263 vdd.n361 gnd 0.009922f
C2264 vdd.n362 gnd 0.009922f
C2265 vdd.n363 gnd 0.009922f
C2266 vdd.n364 gnd 0.009922f
C2267 vdd.n365 gnd 0.009922f
C2268 vdd.n366 gnd 0.007986f
C2269 vdd.n368 gnd 0.009922f
C2270 vdd.n369 gnd 0.009922f
C2271 vdd.n370 gnd 0.009922f
C2272 vdd.n371 gnd 0.009922f
C2273 vdd.n372 gnd 0.009922f
C2274 vdd.n373 gnd 0.007986f
C2275 vdd.n375 gnd 0.009922f
C2276 vdd.n376 gnd 0.009922f
C2277 vdd.n377 gnd 0.009922f
C2278 vdd.n378 gnd 0.009922f
C2279 vdd.n379 gnd 0.009922f
C2280 vdd.n380 gnd 0.007986f
C2281 vdd.n382 gnd 0.009922f
C2282 vdd.n383 gnd 0.009922f
C2283 vdd.n384 gnd 0.009922f
C2284 vdd.n385 gnd 0.009922f
C2285 vdd.n386 gnd 0.006669f
C2286 vdd.t129 gnd 0.122072f
C2287 vdd.t128 gnd 0.130462f
C2288 vdd.t127 gnd 0.159425f
C2289 vdd.n387 gnd 0.20436f
C2290 vdd.n388 gnd 0.172498f
C2291 vdd.n390 gnd 0.009922f
C2292 vdd.n391 gnd 0.009922f
C2293 vdd.n392 gnd 0.007986f
C2294 vdd.n393 gnd 0.009922f
C2295 vdd.n395 gnd 0.009922f
C2296 vdd.n396 gnd 0.009922f
C2297 vdd.n397 gnd 0.009922f
C2298 vdd.n398 gnd 0.009922f
C2299 vdd.n399 gnd 0.007986f
C2300 vdd.n401 gnd 0.009922f
C2301 vdd.n402 gnd 0.009922f
C2302 vdd.n403 gnd 0.009922f
C2303 vdd.n404 gnd 0.009922f
C2304 vdd.n405 gnd 0.009922f
C2305 vdd.n406 gnd 0.007986f
C2306 vdd.n408 gnd 0.009922f
C2307 vdd.n409 gnd 0.009922f
C2308 vdd.n410 gnd 0.009922f
C2309 vdd.n411 gnd 0.009922f
C2310 vdd.n412 gnd 0.009922f
C2311 vdd.n413 gnd 0.007986f
C2312 vdd.n415 gnd 0.009922f
C2313 vdd.n416 gnd 0.009922f
C2314 vdd.n417 gnd 0.009922f
C2315 vdd.n418 gnd 0.009922f
C2316 vdd.n419 gnd 0.009922f
C2317 vdd.n420 gnd 0.007986f
C2318 vdd.n422 gnd 0.009922f
C2319 vdd.n423 gnd 0.009922f
C2320 vdd.n424 gnd 0.009922f
C2321 vdd.n425 gnd 0.009922f
C2322 vdd.n426 gnd 0.007907f
C2323 vdd.t117 gnd 0.122072f
C2324 vdd.t116 gnd 0.130462f
C2325 vdd.t114 gnd 0.159425f
C2326 vdd.n427 gnd 0.20436f
C2327 vdd.n428 gnd 0.172498f
C2328 vdd.n430 gnd 0.009922f
C2329 vdd.n431 gnd 0.009922f
C2330 vdd.n432 gnd 0.007986f
C2331 vdd.n433 gnd 0.009922f
C2332 vdd.n435 gnd 0.009922f
C2333 vdd.n436 gnd 0.009922f
C2334 vdd.n437 gnd 0.009922f
C2335 vdd.n438 gnd 0.009922f
C2336 vdd.n439 gnd 0.007986f
C2337 vdd.n441 gnd 0.009922f
C2338 vdd.n442 gnd 0.009922f
C2339 vdd.n443 gnd 0.009922f
C2340 vdd.n444 gnd 0.009922f
C2341 vdd.n445 gnd 0.009922f
C2342 vdd.n446 gnd 0.007986f
C2343 vdd.n448 gnd 0.009922f
C2344 vdd.n449 gnd 0.009922f
C2345 vdd.n450 gnd 0.009922f
C2346 vdd.n451 gnd 0.009922f
C2347 vdd.n452 gnd 0.009922f
C2348 vdd.n453 gnd 0.007986f
C2349 vdd.n455 gnd 0.009922f
C2350 vdd.n456 gnd 0.009922f
C2351 vdd.n457 gnd 0.009922f
C2352 vdd.n458 gnd 0.009922f
C2353 vdd.n459 gnd 0.009922f
C2354 vdd.n460 gnd 0.007986f
C2355 vdd.n462 gnd 0.009922f
C2356 vdd.n463 gnd 0.009922f
C2357 vdd.n464 gnd 0.009922f
C2358 vdd.n465 gnd 0.009922f
C2359 vdd.n466 gnd 0.009922f
C2360 vdd.n467 gnd 0.009922f
C2361 vdd.n468 gnd 0.007986f
C2362 vdd.n469 gnd 0.009922f
C2363 vdd.n470 gnd 0.009922f
C2364 vdd.n471 gnd 0.007986f
C2365 vdd.n472 gnd 0.009922f
C2366 vdd.n473 gnd 0.009922f
C2367 vdd.n474 gnd 0.007986f
C2368 vdd.n475 gnd 0.009922f
C2369 vdd.n476 gnd 0.007986f
C2370 vdd.n477 gnd 0.009922f
C2371 vdd.n478 gnd 0.007986f
C2372 vdd.n479 gnd 0.009922f
C2373 vdd.n480 gnd 0.009922f
C2374 vdd.t6 gnd 0.507014f
C2375 vdd.n481 gnd 0.542505f
C2376 vdd.n482 gnd 0.009922f
C2377 vdd.n483 gnd 0.007986f
C2378 vdd.n484 gnd 0.009922f
C2379 vdd.n485 gnd 0.007986f
C2380 vdd.n486 gnd 0.009922f
C2381 vdd.t147 gnd 0.507014f
C2382 vdd.n487 gnd 0.009922f
C2383 vdd.n488 gnd 0.007986f
C2384 vdd.n489 gnd 0.009922f
C2385 vdd.n490 gnd 0.007986f
C2386 vdd.n491 gnd 0.009922f
C2387 vdd.n492 gnd 0.796012f
C2388 vdd.n493 gnd 0.841643f
C2389 vdd.t28 gnd 0.507014f
C2390 vdd.n494 gnd 0.009922f
C2391 vdd.n495 gnd 0.007986f
C2392 vdd.n496 gnd 0.009922f
C2393 vdd.n497 gnd 0.007986f
C2394 vdd.n498 gnd 0.009922f
C2395 vdd.n499 gnd 0.623627f
C2396 vdd.n500 gnd 0.009922f
C2397 vdd.n501 gnd 0.007986f
C2398 vdd.n502 gnd 0.009922f
C2399 vdd.n503 gnd 0.007986f
C2400 vdd.n504 gnd 0.009922f
C2401 vdd.n505 gnd 1.01403f
C2402 vdd.t21 gnd 0.507014f
C2403 vdd.n506 gnd 0.009922f
C2404 vdd.n507 gnd 0.007986f
C2405 vdd.n508 gnd 0.009922f
C2406 vdd.n509 gnd 0.007986f
C2407 vdd.n510 gnd 0.009922f
C2408 vdd.n511 gnd 0.542505f
C2409 vdd.n512 gnd 0.009922f
C2410 vdd.n513 gnd 0.007986f
C2411 vdd.n514 gnd 0.023749f
C2412 vdd.n515 gnd 0.023749f
C2413 vdd.n516 gnd 7.26044f
C2414 vdd.t55 gnd 0.507014f
C2415 vdd.n517 gnd 0.023749f
C2416 vdd.n518 gnd 0.008533f
C2417 vdd.n519 gnd 0.007986f
C2418 vdd.n524 gnd 0.00635f
C2419 vdd.n525 gnd 0.007986f
C2420 vdd.n526 gnd 0.009922f
C2421 vdd.n527 gnd 0.009922f
C2422 vdd.n528 gnd 0.009922f
C2423 vdd.n529 gnd 0.009922f
C2424 vdd.n530 gnd 0.009922f
C2425 vdd.n531 gnd 0.007986f
C2426 vdd.n532 gnd 0.009922f
C2427 vdd.n533 gnd 0.009922f
C2428 vdd.n534 gnd 0.009922f
C2429 vdd.n535 gnd 0.009922f
C2430 vdd.n536 gnd 0.009922f
C2431 vdd.n537 gnd 0.007986f
C2432 vdd.n538 gnd 0.009922f
C2433 vdd.n539 gnd 0.009922f
C2434 vdd.n540 gnd 0.009922f
C2435 vdd.n541 gnd 0.009922f
C2436 vdd.n542 gnd 0.009922f
C2437 vdd.t59 gnd 0.122072f
C2438 vdd.t60 gnd 0.130462f
C2439 vdd.t58 gnd 0.159425f
C2440 vdd.n543 gnd 0.20436f
C2441 vdd.n544 gnd 0.171699f
C2442 vdd.n545 gnd 0.016292f
C2443 vdd.n546 gnd 0.009922f
C2444 vdd.n547 gnd 0.009922f
C2445 vdd.n548 gnd 0.009922f
C2446 vdd.n549 gnd 0.009922f
C2447 vdd.n550 gnd 0.009922f
C2448 vdd.n551 gnd 0.007986f
C2449 vdd.n552 gnd 0.009922f
C2450 vdd.n553 gnd 0.009922f
C2451 vdd.n554 gnd 0.009922f
C2452 vdd.n555 gnd 0.009922f
C2453 vdd.n556 gnd 0.009922f
C2454 vdd.n557 gnd 0.007986f
C2455 vdd.n558 gnd 0.009922f
C2456 vdd.n559 gnd 0.009922f
C2457 vdd.n560 gnd 0.009922f
C2458 vdd.n561 gnd 0.009922f
C2459 vdd.n562 gnd 0.009922f
C2460 vdd.n563 gnd 0.007986f
C2461 vdd.n564 gnd 0.009922f
C2462 vdd.n565 gnd 0.009922f
C2463 vdd.n566 gnd 0.009922f
C2464 vdd.n567 gnd 0.009922f
C2465 vdd.n568 gnd 0.009922f
C2466 vdd.n569 gnd 0.007986f
C2467 vdd.n570 gnd 0.009922f
C2468 vdd.n571 gnd 0.009922f
C2469 vdd.n572 gnd 0.009922f
C2470 vdd.n573 gnd 0.009922f
C2471 vdd.n574 gnd 0.009922f
C2472 vdd.n575 gnd 0.007986f
C2473 vdd.n576 gnd 0.009922f
C2474 vdd.n577 gnd 0.009922f
C2475 vdd.n578 gnd 0.009922f
C2476 vdd.n579 gnd 0.007907f
C2477 vdd.t56 gnd 0.122072f
C2478 vdd.t57 gnd 0.130462f
C2479 vdd.t54 gnd 0.159425f
C2480 vdd.n580 gnd 0.20436f
C2481 vdd.n581 gnd 0.171699f
C2482 vdd.n582 gnd 0.009922f
C2483 vdd.n583 gnd 0.007986f
C2484 vdd.n585 gnd 0.009922f
C2485 vdd.n587 gnd 0.009922f
C2486 vdd.n588 gnd 0.009922f
C2487 vdd.n589 gnd 0.007986f
C2488 vdd.n590 gnd 0.009922f
C2489 vdd.n591 gnd 0.009922f
C2490 vdd.n592 gnd 0.009922f
C2491 vdd.n593 gnd 0.009922f
C2492 vdd.n594 gnd 0.009922f
C2493 vdd.n595 gnd 0.007986f
C2494 vdd.n596 gnd 0.009922f
C2495 vdd.n597 gnd 0.009922f
C2496 vdd.n598 gnd 0.009922f
C2497 vdd.n599 gnd 0.009922f
C2498 vdd.n600 gnd 0.009922f
C2499 vdd.n601 gnd 0.007986f
C2500 vdd.n602 gnd 0.009922f
C2501 vdd.n603 gnd 0.009922f
C2502 vdd.n604 gnd 0.009922f
C2503 vdd.n605 gnd 0.00635f
C2504 vdd.n610 gnd 0.006747f
C2505 vdd.n611 gnd 0.006747f
C2506 vdd.n612 gnd 0.006747f
C2507 vdd.n613 gnd 6.98665f
C2508 vdd.n614 gnd 0.006747f
C2509 vdd.n615 gnd 0.006747f
C2510 vdd.n616 gnd 0.006747f
C2511 vdd.n618 gnd 0.006747f
C2512 vdd.n619 gnd 0.006747f
C2513 vdd.n621 gnd 0.006747f
C2514 vdd.n622 gnd 0.004912f
C2515 vdd.n624 gnd 0.006747f
C2516 vdd.t96 gnd 0.272656f
C2517 vdd.t95 gnd 0.279098f
C2518 vdd.t94 gnd 0.178f
C2519 vdd.n625 gnd 0.096199f
C2520 vdd.n626 gnd 0.054567f
C2521 vdd.n627 gnd 0.009643f
C2522 vdd.n628 gnd 0.01577f
C2523 vdd.n630 gnd 0.006747f
C2524 vdd.n631 gnd 0.689539f
C2525 vdd.n632 gnd 0.014948f
C2526 vdd.n633 gnd 0.014948f
C2527 vdd.n634 gnd 0.006747f
C2528 vdd.n635 gnd 0.01601f
C2529 vdd.n636 gnd 0.006747f
C2530 vdd.n637 gnd 0.006747f
C2531 vdd.n638 gnd 0.006747f
C2532 vdd.n639 gnd 0.006747f
C2533 vdd.n640 gnd 0.006747f
C2534 vdd.n642 gnd 0.006747f
C2535 vdd.n643 gnd 0.006747f
C2536 vdd.n645 gnd 0.006747f
C2537 vdd.n646 gnd 0.006747f
C2538 vdd.n648 gnd 0.006747f
C2539 vdd.n649 gnd 0.006747f
C2540 vdd.n651 gnd 0.006747f
C2541 vdd.n652 gnd 0.006747f
C2542 vdd.n654 gnd 0.006747f
C2543 vdd.n655 gnd 0.006747f
C2544 vdd.n657 gnd 0.006747f
C2545 vdd.n658 gnd 0.004912f
C2546 vdd.n660 gnd 0.006747f
C2547 vdd.t89 gnd 0.272656f
C2548 vdd.t88 gnd 0.279098f
C2549 vdd.t86 gnd 0.178f
C2550 vdd.n661 gnd 0.096199f
C2551 vdd.n662 gnd 0.054567f
C2552 vdd.n663 gnd 0.009643f
C2553 vdd.n664 gnd 0.006747f
C2554 vdd.n665 gnd 0.006747f
C2555 vdd.t87 gnd 0.344769f
C2556 vdd.n666 gnd 0.006747f
C2557 vdd.n667 gnd 0.006747f
C2558 vdd.n668 gnd 0.006747f
C2559 vdd.n669 gnd 0.006747f
C2560 vdd.n670 gnd 0.006747f
C2561 vdd.n671 gnd 0.689539f
C2562 vdd.n672 gnd 0.006747f
C2563 vdd.n673 gnd 0.006747f
C2564 vdd.n674 gnd 0.603347f
C2565 vdd.n675 gnd 0.006747f
C2566 vdd.n676 gnd 0.006747f
C2567 vdd.n677 gnd 0.005953f
C2568 vdd.n678 gnd 0.006747f
C2569 vdd.n679 gnd 0.608417f
C2570 vdd.n680 gnd 0.006747f
C2571 vdd.n681 gnd 0.006747f
C2572 vdd.n682 gnd 0.006747f
C2573 vdd.n683 gnd 0.006747f
C2574 vdd.n684 gnd 0.006747f
C2575 vdd.n685 gnd 0.689539f
C2576 vdd.n686 gnd 0.006747f
C2577 vdd.n687 gnd 0.006747f
C2578 vdd.t70 gnd 0.309278f
C2579 vdd.t38 gnd 0.081122f
C2580 vdd.n688 gnd 0.006747f
C2581 vdd.n689 gnd 0.006747f
C2582 vdd.n690 gnd 0.006747f
C2583 vdd.t146 gnd 0.344769f
C2584 vdd.n691 gnd 0.006747f
C2585 vdd.n692 gnd 0.006747f
C2586 vdd.n693 gnd 0.006747f
C2587 vdd.n694 gnd 0.006747f
C2588 vdd.n695 gnd 0.006747f
C2589 vdd.t143 gnd 0.344769f
C2590 vdd.n696 gnd 0.006747f
C2591 vdd.n697 gnd 0.006747f
C2592 vdd.n698 gnd 0.572926f
C2593 vdd.n699 gnd 0.006747f
C2594 vdd.n700 gnd 0.006747f
C2595 vdd.n701 gnd 0.006747f
C2596 vdd.n702 gnd 0.420822f
C2597 vdd.n703 gnd 0.006747f
C2598 vdd.n704 gnd 0.006747f
C2599 vdd.t198 gnd 0.344769f
C2600 vdd.n705 gnd 0.006747f
C2601 vdd.n706 gnd 0.006747f
C2602 vdd.n707 gnd 0.006747f
C2603 vdd.n708 gnd 0.572926f
C2604 vdd.n709 gnd 0.006747f
C2605 vdd.n710 gnd 0.006747f
C2606 vdd.t16 gnd 0.294068f
C2607 vdd.t161 gnd 0.268717f
C2608 vdd.n711 gnd 0.006747f
C2609 vdd.n712 gnd 0.006747f
C2610 vdd.n713 gnd 0.006747f
C2611 vdd.t165 gnd 0.344769f
C2612 vdd.n714 gnd 0.006747f
C2613 vdd.n715 gnd 0.006747f
C2614 vdd.t34 gnd 0.344769f
C2615 vdd.n716 gnd 0.006747f
C2616 vdd.n717 gnd 0.006747f
C2617 vdd.n718 gnd 0.006747f
C2618 vdd.t15 gnd 0.253507f
C2619 vdd.n719 gnd 0.006747f
C2620 vdd.n720 gnd 0.006747f
C2621 vdd.n721 gnd 0.588136f
C2622 vdd.n722 gnd 0.006747f
C2623 vdd.n723 gnd 0.006747f
C2624 vdd.n724 gnd 0.006747f
C2625 vdd.n725 gnd 0.689539f
C2626 vdd.n726 gnd 0.006747f
C2627 vdd.n727 gnd 0.006747f
C2628 vdd.t130 gnd 0.309278f
C2629 vdd.n728 gnd 0.436032f
C2630 vdd.n729 gnd 0.006747f
C2631 vdd.n730 gnd 0.006747f
C2632 vdd.n731 gnd 0.006747f
C2633 vdd.t13 gnd 0.344769f
C2634 vdd.n732 gnd 0.006747f
C2635 vdd.n733 gnd 0.006747f
C2636 vdd.n734 gnd 0.006747f
C2637 vdd.n735 gnd 0.006747f
C2638 vdd.n736 gnd 0.006747f
C2639 vdd.t170 gnd 0.689539f
C2640 vdd.n737 gnd 0.006747f
C2641 vdd.n738 gnd 0.006747f
C2642 vdd.t91 gnd 0.344769f
C2643 vdd.n739 gnd 0.006747f
C2644 vdd.n740 gnd 0.01601f
C2645 vdd.n741 gnd 0.01601f
C2646 vdd.t172 gnd 0.648978f
C2647 vdd.n742 gnd 0.014948f
C2648 vdd.n743 gnd 0.014948f
C2649 vdd.n744 gnd 0.01601f
C2650 vdd.n745 gnd 0.006747f
C2651 vdd.n746 gnd 0.006747f
C2652 vdd.t163 gnd 0.648978f
C2653 vdd.n764 gnd 0.01601f
C2654 vdd.n782 gnd 0.014948f
C2655 vdd.n783 gnd 0.006747f
C2656 vdd.n784 gnd 0.014948f
C2657 vdd.t110 gnd 0.272656f
C2658 vdd.t109 gnd 0.279098f
C2659 vdd.t108 gnd 0.178f
C2660 vdd.n785 gnd 0.096199f
C2661 vdd.n786 gnd 0.054567f
C2662 vdd.n787 gnd 0.01577f
C2663 vdd.n788 gnd 0.006747f
C2664 vdd.t144 gnd 0.689539f
C2665 vdd.n789 gnd 0.014948f
C2666 vdd.n790 gnd 0.006747f
C2667 vdd.n791 gnd 0.01601f
C2668 vdd.n792 gnd 0.006747f
C2669 vdd.t85 gnd 0.272656f
C2670 vdd.t84 gnd 0.279098f
C2671 vdd.t82 gnd 0.178f
C2672 vdd.n793 gnd 0.096199f
C2673 vdd.n794 gnd 0.054567f
C2674 vdd.n795 gnd 0.009643f
C2675 vdd.n796 gnd 0.006747f
C2676 vdd.n797 gnd 0.006747f
C2677 vdd.t83 gnd 0.344769f
C2678 vdd.n798 gnd 0.006747f
C2679 vdd.n799 gnd 0.006747f
C2680 vdd.n800 gnd 0.006747f
C2681 vdd.n801 gnd 0.006747f
C2682 vdd.n802 gnd 0.006747f
C2683 vdd.n803 gnd 0.006747f
C2684 vdd.n804 gnd 0.689539f
C2685 vdd.n805 gnd 0.006747f
C2686 vdd.n806 gnd 0.006747f
C2687 vdd.t196 gnd 0.344769f
C2688 vdd.n807 gnd 0.006747f
C2689 vdd.n808 gnd 0.006747f
C2690 vdd.n809 gnd 0.006747f
C2691 vdd.n810 gnd 0.006747f
C2692 vdd.n811 gnd 0.436032f
C2693 vdd.n812 gnd 0.006747f
C2694 vdd.n813 gnd 0.006747f
C2695 vdd.n814 gnd 0.006747f
C2696 vdd.n815 gnd 0.006747f
C2697 vdd.n816 gnd 0.006747f
C2698 vdd.n817 gnd 0.588136f
C2699 vdd.n818 gnd 0.006747f
C2700 vdd.n819 gnd 0.006747f
C2701 vdd.t226 gnd 0.309278f
C2702 vdd.t9 gnd 0.253507f
C2703 vdd.n820 gnd 0.006747f
C2704 vdd.n821 gnd 0.006747f
C2705 vdd.n822 gnd 0.006747f
C2706 vdd.t132 gnd 0.344769f
C2707 vdd.n823 gnd 0.006747f
C2708 vdd.n824 gnd 0.006747f
C2709 vdd.t159 gnd 0.344769f
C2710 vdd.n825 gnd 0.006747f
C2711 vdd.n826 gnd 0.006747f
C2712 vdd.n827 gnd 0.006747f
C2713 vdd.t184 gnd 0.268717f
C2714 vdd.n828 gnd 0.006747f
C2715 vdd.n829 gnd 0.006747f
C2716 vdd.n830 gnd 0.572926f
C2717 vdd.n831 gnd 0.006747f
C2718 vdd.n832 gnd 0.006747f
C2719 vdd.n833 gnd 0.006747f
C2720 vdd.t220 gnd 0.344769f
C2721 vdd.n834 gnd 0.006747f
C2722 vdd.n835 gnd 0.006747f
C2723 vdd.t219 gnd 0.294068f
C2724 vdd.n836 gnd 0.420822f
C2725 vdd.n837 gnd 0.006747f
C2726 vdd.n838 gnd 0.006747f
C2727 vdd.n839 gnd 0.006747f
C2728 vdd.n840 gnd 0.572926f
C2729 vdd.n841 gnd 0.006747f
C2730 vdd.n842 gnd 0.006747f
C2731 vdd.t151 gnd 0.344769f
C2732 vdd.n843 gnd 0.006747f
C2733 vdd.n844 gnd 0.006747f
C2734 vdd.n845 gnd 0.006747f
C2735 vdd.n846 gnd 0.689539f
C2736 vdd.n847 gnd 0.006747f
C2737 vdd.n848 gnd 0.006747f
C2738 vdd.t174 gnd 0.344769f
C2739 vdd.n849 gnd 0.006747f
C2740 vdd.n850 gnd 0.006747f
C2741 vdd.n851 gnd 0.006747f
C2742 vdd.t3 gnd 0.081122f
C2743 vdd.n852 gnd 0.006747f
C2744 vdd.n853 gnd 0.006747f
C2745 vdd.n854 gnd 0.006747f
C2746 vdd.t103 gnd 0.279098f
C2747 vdd.t101 gnd 0.178f
C2748 vdd.t104 gnd 0.279098f
C2749 vdd.n855 gnd 0.156864f
C2750 vdd.n856 gnd 0.006747f
C2751 vdd.n857 gnd 0.006747f
C2752 vdd.n858 gnd 0.689539f
C2753 vdd.n859 gnd 0.006747f
C2754 vdd.n860 gnd 0.006747f
C2755 vdd.t102 gnd 0.309278f
C2756 vdd.n861 gnd 0.608417f
C2757 vdd.n862 gnd 0.006747f
C2758 vdd.n863 gnd 0.006747f
C2759 vdd.n864 gnd 0.006747f
C2760 vdd.n865 gnd 0.603347f
C2761 vdd.n866 gnd 0.006747f
C2762 vdd.n867 gnd 0.006747f
C2763 vdd.n868 gnd 0.006747f
C2764 vdd.n869 gnd 0.006747f
C2765 vdd.n870 gnd 0.006747f
C2766 vdd.n871 gnd 0.689539f
C2767 vdd.n872 gnd 0.006747f
C2768 vdd.n873 gnd 0.006747f
C2769 vdd.t98 gnd 0.344769f
C2770 vdd.n874 gnd 0.006747f
C2771 vdd.n875 gnd 0.01601f
C2772 vdd.n876 gnd 0.01601f
C2773 vdd.n877 gnd 6.98665f
C2774 vdd.n878 gnd 0.014948f
C2775 vdd.n879 gnd 0.014948f
C2776 vdd.n880 gnd 0.01601f
C2777 vdd.n881 gnd 0.006747f
C2778 vdd.n882 gnd 0.006747f
C2779 vdd.n883 gnd 0.006747f
C2780 vdd.n884 gnd 0.006747f
C2781 vdd.n885 gnd 0.006747f
C2782 vdd.n886 gnd 0.006747f
C2783 vdd.n887 gnd 0.006747f
C2784 vdd.n888 gnd 0.006747f
C2785 vdd.n890 gnd 0.006747f
C2786 vdd.n891 gnd 0.006747f
C2787 vdd.n892 gnd 0.00635f
C2788 vdd.n895 gnd 0.023749f
C2789 vdd.n896 gnd 0.007986f
C2790 vdd.n897 gnd 0.009922f
C2791 vdd.n899 gnd 0.009922f
C2792 vdd.n900 gnd 0.006629f
C2793 vdd.t62 gnd 0.507014f
C2794 vdd.n901 gnd 7.26044f
C2795 vdd.n902 gnd 0.009922f
C2796 vdd.n903 gnd 0.023749f
C2797 vdd.n904 gnd 0.007986f
C2798 vdd.n905 gnd 0.009922f
C2799 vdd.n906 gnd 0.007986f
C2800 vdd.n907 gnd 0.009922f
C2801 vdd.n908 gnd 1.01403f
C2802 vdd.n909 gnd 0.009922f
C2803 vdd.n910 gnd 0.007986f
C2804 vdd.n911 gnd 0.007986f
C2805 vdd.n912 gnd 0.009922f
C2806 vdd.n913 gnd 0.007986f
C2807 vdd.n914 gnd 0.009922f
C2808 vdd.t42 gnd 0.507014f
C2809 vdd.n915 gnd 0.009922f
C2810 vdd.n916 gnd 0.007986f
C2811 vdd.n917 gnd 0.009922f
C2812 vdd.n918 gnd 0.007986f
C2813 vdd.n919 gnd 0.009922f
C2814 vdd.t44 gnd 0.507014f
C2815 vdd.n920 gnd 0.009922f
C2816 vdd.n921 gnd 0.007986f
C2817 vdd.n922 gnd 0.009922f
C2818 vdd.n923 gnd 0.007986f
C2819 vdd.n924 gnd 0.009922f
C2820 vdd.t4 gnd 0.507014f
C2821 vdd.n925 gnd 0.796012f
C2822 vdd.n926 gnd 0.009922f
C2823 vdd.n927 gnd 0.007986f
C2824 vdd.n928 gnd 0.009922f
C2825 vdd.n929 gnd 0.007986f
C2826 vdd.n930 gnd 0.009922f
C2827 vdd.n931 gnd 0.71489f
C2828 vdd.n932 gnd 0.009922f
C2829 vdd.n933 gnd 0.007986f
C2830 vdd.n934 gnd 0.009922f
C2831 vdd.n935 gnd 0.007986f
C2832 vdd.n936 gnd 0.009922f
C2833 vdd.n937 gnd 0.542505f
C2834 vdd.t30 gnd 0.507014f
C2835 vdd.n938 gnd 0.009922f
C2836 vdd.n939 gnd 0.007986f
C2837 vdd.n940 gnd 0.009888f
C2838 vdd.n941 gnd 0.007986f
C2839 vdd.n942 gnd 0.009922f
C2840 vdd.t208 gnd 0.507014f
C2841 vdd.n943 gnd 0.009922f
C2842 vdd.n944 gnd 0.007986f
C2843 vdd.n945 gnd 0.009922f
C2844 vdd.n946 gnd 0.007986f
C2845 vdd.n947 gnd 0.009922f
C2846 vdd.t25 gnd 0.507014f
C2847 vdd.n948 gnd 0.643908f
C2848 vdd.n949 gnd 0.009922f
C2849 vdd.n950 gnd 0.007986f
C2850 vdd.n951 gnd 0.009922f
C2851 vdd.n952 gnd 0.007986f
C2852 vdd.n953 gnd 0.009922f
C2853 vdd.t32 gnd 0.507014f
C2854 vdd.n954 gnd 0.009922f
C2855 vdd.n955 gnd 0.007986f
C2856 vdd.n956 gnd 0.009922f
C2857 vdd.n957 gnd 0.007986f
C2858 vdd.n958 gnd 0.009922f
C2859 vdd.n959 gnd 0.694609f
C2860 vdd.n960 gnd 0.841643f
C2861 vdd.t168 gnd 0.507014f
C2862 vdd.n961 gnd 0.009922f
C2863 vdd.n962 gnd 0.007986f
C2864 vdd.n963 gnd 0.009922f
C2865 vdd.n964 gnd 0.007986f
C2866 vdd.n965 gnd 0.009922f
C2867 vdd.n966 gnd 0.522224f
C2868 vdd.n967 gnd 0.009922f
C2869 vdd.n968 gnd 0.007986f
C2870 vdd.n969 gnd 0.009922f
C2871 vdd.n970 gnd 0.007986f
C2872 vdd.n971 gnd 0.009922f
C2873 vdd.n972 gnd 1.01403f
C2874 vdd.t46 gnd 0.507014f
C2875 vdd.n973 gnd 0.009922f
C2876 vdd.n974 gnd 0.007986f
C2877 vdd.n975 gnd 0.009922f
C2878 vdd.n976 gnd 0.007986f
C2879 vdd.n977 gnd 0.009922f
C2880 vdd.t66 gnd 0.507014f
C2881 vdd.n978 gnd 0.009922f
C2882 vdd.n979 gnd 0.007986f
C2883 vdd.n980 gnd 0.023749f
C2884 vdd.n981 gnd 0.023749f
C2885 vdd.n982 gnd 2.33226f
C2886 vdd.n983 gnd 0.572926f
C2887 vdd.n984 gnd 0.023749f
C2888 vdd.n985 gnd 0.009922f
C2889 vdd.n987 gnd 0.009922f
C2890 vdd.n988 gnd 0.009922f
C2891 vdd.n989 gnd 0.007986f
C2892 vdd.n990 gnd 0.009922f
C2893 vdd.n991 gnd 0.009922f
C2894 vdd.n993 gnd 0.009922f
C2895 vdd.n994 gnd 0.009922f
C2896 vdd.n996 gnd 0.009922f
C2897 vdd.n997 gnd 0.007986f
C2898 vdd.n998 gnd 0.009922f
C2899 vdd.n999 gnd 0.009922f
C2900 vdd.n1001 gnd 0.009922f
C2901 vdd.n1002 gnd 0.009922f
C2902 vdd.n1004 gnd 0.009922f
C2903 vdd.n1005 gnd 0.007986f
C2904 vdd.n1006 gnd 0.009922f
C2905 vdd.n1007 gnd 0.009922f
C2906 vdd.n1009 gnd 0.009922f
C2907 vdd.n1010 gnd 0.009922f
C2908 vdd.n1012 gnd 0.009922f
C2909 vdd.n1013 gnd 0.007986f
C2910 vdd.n1014 gnd 0.009922f
C2911 vdd.n1015 gnd 0.009922f
C2912 vdd.n1017 gnd 0.009922f
C2913 vdd.n1018 gnd 0.009922f
C2914 vdd.n1020 gnd 0.009922f
C2915 vdd.t77 gnd 0.122072f
C2916 vdd.t78 gnd 0.130462f
C2917 vdd.t76 gnd 0.159425f
C2918 vdd.n1021 gnd 0.20436f
C2919 vdd.n1022 gnd 0.172498f
C2920 vdd.n1023 gnd 0.017091f
C2921 vdd.n1024 gnd 0.009922f
C2922 vdd.n1025 gnd 0.009922f
C2923 vdd.n1027 gnd 0.009922f
C2924 vdd.n1028 gnd 0.009922f
C2925 vdd.n1030 gnd 0.009922f
C2926 vdd.n1031 gnd 0.007986f
C2927 vdd.n1032 gnd 0.009922f
C2928 vdd.n1033 gnd 0.009922f
C2929 vdd.n1035 gnd 0.009922f
C2930 vdd.n1036 gnd 0.009922f
C2931 vdd.n1038 gnd 0.009922f
C2932 vdd.n1039 gnd 0.007986f
C2933 vdd.n1040 gnd 0.009922f
C2934 vdd.n1041 gnd 0.009922f
C2935 vdd.n1043 gnd 0.009922f
C2936 vdd.n1044 gnd 0.009922f
C2937 vdd.n1046 gnd 0.009922f
C2938 vdd.n1047 gnd 0.007986f
C2939 vdd.n1048 gnd 0.009922f
C2940 vdd.n1049 gnd 0.009922f
C2941 vdd.n1051 gnd 0.009922f
C2942 vdd.n1052 gnd 0.009922f
C2943 vdd.n1054 gnd 0.009922f
C2944 vdd.n1055 gnd 0.007986f
C2945 vdd.n1056 gnd 0.009922f
C2946 vdd.n1057 gnd 0.009922f
C2947 vdd.n1059 gnd 0.009922f
C2948 vdd.n1060 gnd 0.009922f
C2949 vdd.n1062 gnd 0.009922f
C2950 vdd.n1063 gnd 0.007986f
C2951 vdd.n1064 gnd 0.009922f
C2952 vdd.n1065 gnd 0.009922f
C2953 vdd.n1067 gnd 0.009922f
C2954 vdd.n1068 gnd 0.007907f
C2955 vdd.n1070 gnd 0.007986f
C2956 vdd.n1071 gnd 0.009922f
C2957 vdd.n1072 gnd 0.009922f
C2958 vdd.n1073 gnd 0.009922f
C2959 vdd.n1074 gnd 0.009922f
C2960 vdd.n1076 gnd 0.009922f
C2961 vdd.n1077 gnd 0.009922f
C2962 vdd.n1078 gnd 0.007986f
C2963 vdd.n1079 gnd 0.009922f
C2964 vdd.n1081 gnd 0.009922f
C2965 vdd.n1082 gnd 0.009922f
C2966 vdd.n1084 gnd 0.009922f
C2967 vdd.n1085 gnd 0.009922f
C2968 vdd.n1086 gnd 0.007986f
C2969 vdd.n1087 gnd 0.009922f
C2970 vdd.n1089 gnd 0.009922f
C2971 vdd.n1090 gnd 0.009922f
C2972 vdd.n1092 gnd 0.009922f
C2973 vdd.n1093 gnd 0.009922f
C2974 vdd.n1094 gnd 0.007986f
C2975 vdd.n1095 gnd 0.009922f
C2976 vdd.n1097 gnd 0.009922f
C2977 vdd.n1098 gnd 0.009922f
C2978 vdd.n1100 gnd 0.009922f
C2979 vdd.n1101 gnd 0.009922f
C2980 vdd.n1102 gnd 0.007986f
C2981 vdd.n1103 gnd 0.009922f
C2982 vdd.n1105 gnd 0.009922f
C2983 vdd.n1106 gnd 0.009922f
C2984 vdd.n1108 gnd 0.009922f
C2985 vdd.n1109 gnd 0.003794f
C2986 vdd.t119 gnd 0.122072f
C2987 vdd.t120 gnd 0.130462f
C2988 vdd.t118 gnd 0.159425f
C2989 vdd.n1110 gnd 0.20436f
C2990 vdd.n1111 gnd 0.172498f
C2991 vdd.n1112 gnd 0.013098f
C2992 vdd.n1113 gnd 0.004193f
C2993 vdd.n1114 gnd 0.007986f
C2994 vdd.n1115 gnd 0.009922f
C2995 vdd.n1116 gnd 0.009922f
C2996 vdd.n1117 gnd 0.009922f
C2997 vdd.n1118 gnd 0.007986f
C2998 vdd.n1119 gnd 0.007986f
C2999 vdd.n1120 gnd 0.007986f
C3000 vdd.n1121 gnd 0.009922f
C3001 vdd.n1122 gnd 0.009922f
C3002 vdd.n1123 gnd 0.009922f
C3003 vdd.n1124 gnd 0.007986f
C3004 vdd.n1125 gnd 0.007986f
C3005 vdd.n1126 gnd 0.007986f
C3006 vdd.n1127 gnd 0.009922f
C3007 vdd.n1128 gnd 0.009922f
C3008 vdd.n1129 gnd 0.009922f
C3009 vdd.n1130 gnd 0.007986f
C3010 vdd.n1131 gnd 0.007986f
C3011 vdd.n1132 gnd 0.007986f
C3012 vdd.n1133 gnd 0.009922f
C3013 vdd.n1134 gnd 0.009922f
C3014 vdd.n1135 gnd 0.009922f
C3015 vdd.n1136 gnd 0.007986f
C3016 vdd.n1137 gnd 0.007986f
C3017 vdd.n1138 gnd 0.007986f
C3018 vdd.n1139 gnd 0.009922f
C3019 vdd.n1140 gnd 0.009922f
C3020 vdd.n1141 gnd 0.009922f
C3021 vdd.n1142 gnd 0.007986f
C3022 vdd.n1143 gnd 0.009922f
C3023 vdd.n1144 gnd 0.009922f
C3024 vdd.n1146 gnd 0.009922f
C3025 vdd.t67 gnd 0.122072f
C3026 vdd.t68 gnd 0.130462f
C3027 vdd.t65 gnd 0.159425f
C3028 vdd.n1147 gnd 0.20436f
C3029 vdd.n1148 gnd 0.172498f
C3030 vdd.n1149 gnd 0.017091f
C3031 vdd.n1150 gnd 0.005431f
C3032 vdd.n1151 gnd 0.009922f
C3033 vdd.n1152 gnd 0.009922f
C3034 vdd.n1153 gnd 0.009922f
C3035 vdd.n1154 gnd 0.007986f
C3036 vdd.n1155 gnd 0.007986f
C3037 vdd.n1156 gnd 0.007986f
C3038 vdd.n1157 gnd 0.009922f
C3039 vdd.n1158 gnd 0.009922f
C3040 vdd.n1159 gnd 0.009922f
C3041 vdd.n1160 gnd 0.007986f
C3042 vdd.n1161 gnd 0.007986f
C3043 vdd.n1162 gnd 0.007986f
C3044 vdd.n1163 gnd 0.009922f
C3045 vdd.n1164 gnd 0.009922f
C3046 vdd.n1165 gnd 0.009922f
C3047 vdd.n1166 gnd 0.007986f
C3048 vdd.n1167 gnd 0.007986f
C3049 vdd.n1168 gnd 0.007986f
C3050 vdd.n1169 gnd 0.009922f
C3051 vdd.n1170 gnd 0.009922f
C3052 vdd.n1171 gnd 0.009922f
C3053 vdd.n1172 gnd 0.007986f
C3054 vdd.n1173 gnd 0.007986f
C3055 vdd.n1174 gnd 0.007986f
C3056 vdd.n1175 gnd 0.009922f
C3057 vdd.n1176 gnd 0.009922f
C3058 vdd.n1177 gnd 0.009922f
C3059 vdd.n1178 gnd 0.007986f
C3060 vdd.n1179 gnd 0.007986f
C3061 vdd.n1180 gnd 0.006669f
C3062 vdd.n1181 gnd 0.009922f
C3063 vdd.n1182 gnd 0.009922f
C3064 vdd.n1183 gnd 0.009922f
C3065 vdd.n1184 gnd 0.006669f
C3066 vdd.n1185 gnd 0.007986f
C3067 vdd.n1186 gnd 0.007986f
C3068 vdd.n1187 gnd 0.009922f
C3069 vdd.n1188 gnd 0.009922f
C3070 vdd.n1189 gnd 0.009922f
C3071 vdd.n1190 gnd 0.007986f
C3072 vdd.n1191 gnd 0.007986f
C3073 vdd.n1192 gnd 0.007986f
C3074 vdd.n1193 gnd 0.009922f
C3075 vdd.n1194 gnd 0.009922f
C3076 vdd.n1195 gnd 0.009922f
C3077 vdd.n1196 gnd 0.007986f
C3078 vdd.n1197 gnd 0.007986f
C3079 vdd.n1198 gnd 0.007986f
C3080 vdd.n1199 gnd 0.009922f
C3081 vdd.n1200 gnd 0.009922f
C3082 vdd.n1201 gnd 0.009922f
C3083 vdd.n1202 gnd 0.007986f
C3084 vdd.n1203 gnd 0.007986f
C3085 vdd.n1204 gnd 0.007986f
C3086 vdd.n1205 gnd 0.009922f
C3087 vdd.n1206 gnd 0.009922f
C3088 vdd.n1207 gnd 0.009922f
C3089 vdd.n1208 gnd 0.007986f
C3090 vdd.n1209 gnd 0.007986f
C3091 vdd.n1210 gnd 0.006629f
C3092 vdd.n1211 gnd 0.023749f
C3093 vdd.n1212 gnd 0.023383f
C3094 vdd.n1213 gnd 0.006629f
C3095 vdd.n1214 gnd 0.023383f
C3096 vdd.n1215 gnd 1.42978f
C3097 vdd.n1216 gnd 0.023383f
C3098 vdd.n1217 gnd 0.006629f
C3099 vdd.n1218 gnd 0.023383f
C3100 vdd.n1219 gnd 0.009922f
C3101 vdd.n1220 gnd 0.009922f
C3102 vdd.n1221 gnd 0.007986f
C3103 vdd.n1222 gnd 0.009922f
C3104 vdd.n1223 gnd 0.948116f
C3105 vdd.n1224 gnd 0.009922f
C3106 vdd.n1225 gnd 0.007986f
C3107 vdd.n1226 gnd 0.009922f
C3108 vdd.n1227 gnd 0.009922f
C3109 vdd.n1228 gnd 0.009922f
C3110 vdd.n1229 gnd 0.007986f
C3111 vdd.n1230 gnd 0.009922f
C3112 vdd.n1231 gnd 0.998817f
C3113 vdd.n1232 gnd 0.009922f
C3114 vdd.n1233 gnd 0.007986f
C3115 vdd.n1234 gnd 0.009922f
C3116 vdd.n1235 gnd 0.009922f
C3117 vdd.n1236 gnd 0.009922f
C3118 vdd.n1237 gnd 0.007986f
C3119 vdd.n1238 gnd 0.009922f
C3120 vdd.t48 gnd 0.507014f
C3121 vdd.n1239 gnd 0.826433f
C3122 vdd.n1240 gnd 0.009922f
C3123 vdd.n1241 gnd 0.007986f
C3124 vdd.n1242 gnd 0.009922f
C3125 vdd.n1243 gnd 0.009922f
C3126 vdd.n1244 gnd 0.009922f
C3127 vdd.n1245 gnd 0.007986f
C3128 vdd.n1246 gnd 0.009922f
C3129 vdd.n1247 gnd 0.654048f
C3130 vdd.n1248 gnd 0.009922f
C3131 vdd.n1249 gnd 0.007986f
C3132 vdd.n1250 gnd 0.009922f
C3133 vdd.n1251 gnd 0.009922f
C3134 vdd.n1252 gnd 0.009922f
C3135 vdd.n1253 gnd 0.007986f
C3136 vdd.n1254 gnd 0.009922f
C3137 vdd.n1255 gnd 0.816292f
C3138 vdd.n1256 gnd 0.532365f
C3139 vdd.n1257 gnd 0.009922f
C3140 vdd.n1258 gnd 0.007986f
C3141 vdd.n1259 gnd 0.009922f
C3142 vdd.n1260 gnd 0.009922f
C3143 vdd.n1261 gnd 0.009922f
C3144 vdd.n1262 gnd 0.007986f
C3145 vdd.n1263 gnd 0.009922f
C3146 vdd.n1264 gnd 0.704749f
C3147 vdd.n1265 gnd 0.009922f
C3148 vdd.n1266 gnd 0.007986f
C3149 vdd.n1267 gnd 0.009922f
C3150 vdd.n1268 gnd 0.009922f
C3151 vdd.n1269 gnd 0.009922f
C3152 vdd.n1270 gnd 0.007986f
C3153 vdd.n1271 gnd 0.009922f
C3154 vdd.t178 gnd 0.507014f
C3155 vdd.n1272 gnd 0.841643f
C3156 vdd.n1273 gnd 0.009922f
C3157 vdd.n1274 gnd 0.007986f
C3158 vdd.n1275 gnd 0.005446f
C3159 vdd.n1276 gnd 0.005053f
C3160 vdd.n1277 gnd 0.002795f
C3161 vdd.n1278 gnd 0.006418f
C3162 vdd.n1279 gnd 0.002715f
C3163 vdd.n1280 gnd 0.002875f
C3164 vdd.n1281 gnd 0.005053f
C3165 vdd.n1282 gnd 0.002715f
C3166 vdd.n1283 gnd 0.006418f
C3167 vdd.n1284 gnd 0.002875f
C3168 vdd.n1285 gnd 0.005053f
C3169 vdd.n1286 gnd 0.002715f
C3170 vdd.n1287 gnd 0.004814f
C3171 vdd.n1288 gnd 0.004828f
C3172 vdd.t176 gnd 0.013789f
C3173 vdd.n1289 gnd 0.03068f
C3174 vdd.n1290 gnd 0.159666f
C3175 vdd.n1291 gnd 0.002715f
C3176 vdd.n1292 gnd 0.002875f
C3177 vdd.n1293 gnd 0.006418f
C3178 vdd.n1294 gnd 0.006418f
C3179 vdd.n1295 gnd 0.002875f
C3180 vdd.n1296 gnd 0.002715f
C3181 vdd.n1297 gnd 0.005053f
C3182 vdd.n1298 gnd 0.005053f
C3183 vdd.n1299 gnd 0.002715f
C3184 vdd.n1300 gnd 0.002875f
C3185 vdd.n1301 gnd 0.006418f
C3186 vdd.n1302 gnd 0.006418f
C3187 vdd.n1303 gnd 0.002875f
C3188 vdd.n1304 gnd 0.002715f
C3189 vdd.n1305 gnd 0.005053f
C3190 vdd.n1306 gnd 0.005053f
C3191 vdd.n1307 gnd 0.002715f
C3192 vdd.n1308 gnd 0.002875f
C3193 vdd.n1309 gnd 0.006418f
C3194 vdd.n1310 gnd 0.006418f
C3195 vdd.n1311 gnd 0.015174f
C3196 vdd.n1312 gnd 0.002795f
C3197 vdd.n1313 gnd 0.002715f
C3198 vdd.n1314 gnd 0.013061f
C3199 vdd.n1315 gnd 0.009118f
C3200 vdd.t5 gnd 0.031946f
C3201 vdd.t205 gnd 0.031946f
C3202 vdd.n1316 gnd 0.219551f
C3203 vdd.n1317 gnd 0.172644f
C3204 vdd.t215 gnd 0.031946f
C3205 vdd.t140 gnd 0.031946f
C3206 vdd.n1318 gnd 0.219551f
C3207 vdd.n1319 gnd 0.139322f
C3208 vdd.t222 gnd 0.031946f
C3209 vdd.t206 gnd 0.031946f
C3210 vdd.n1320 gnd 0.219551f
C3211 vdd.n1321 gnd 0.139322f
C3212 vdd.t225 gnd 0.031946f
C3213 vdd.t26 gnd 0.031946f
C3214 vdd.n1322 gnd 0.219551f
C3215 vdd.n1323 gnd 0.139322f
C3216 vdd.t218 gnd 0.031946f
C3217 vdd.t181 gnd 0.031946f
C3218 vdd.n1324 gnd 0.219551f
C3219 vdd.n1325 gnd 0.139322f
C3220 vdd.n1326 gnd 0.005446f
C3221 vdd.n1327 gnd 0.005053f
C3222 vdd.n1328 gnd 0.002795f
C3223 vdd.n1329 gnd 0.006418f
C3224 vdd.n1330 gnd 0.002715f
C3225 vdd.n1331 gnd 0.002875f
C3226 vdd.n1332 gnd 0.005053f
C3227 vdd.n1333 gnd 0.002715f
C3228 vdd.n1334 gnd 0.006418f
C3229 vdd.n1335 gnd 0.002875f
C3230 vdd.n1336 gnd 0.005053f
C3231 vdd.n1337 gnd 0.002715f
C3232 vdd.n1338 gnd 0.004814f
C3233 vdd.n1339 gnd 0.004828f
C3234 vdd.t214 gnd 0.013789f
C3235 vdd.n1340 gnd 0.03068f
C3236 vdd.n1341 gnd 0.159666f
C3237 vdd.n1342 gnd 0.002715f
C3238 vdd.n1343 gnd 0.002875f
C3239 vdd.n1344 gnd 0.006418f
C3240 vdd.n1345 gnd 0.006418f
C3241 vdd.n1346 gnd 0.002875f
C3242 vdd.n1347 gnd 0.002715f
C3243 vdd.n1348 gnd 0.005053f
C3244 vdd.n1349 gnd 0.005053f
C3245 vdd.n1350 gnd 0.002715f
C3246 vdd.n1351 gnd 0.002875f
C3247 vdd.n1352 gnd 0.006418f
C3248 vdd.n1353 gnd 0.006418f
C3249 vdd.n1354 gnd 0.002875f
C3250 vdd.n1355 gnd 0.002715f
C3251 vdd.n1356 gnd 0.005053f
C3252 vdd.n1357 gnd 0.005053f
C3253 vdd.n1358 gnd 0.002715f
C3254 vdd.n1359 gnd 0.002875f
C3255 vdd.n1360 gnd 0.006418f
C3256 vdd.n1361 gnd 0.006418f
C3257 vdd.n1362 gnd 0.015174f
C3258 vdd.n1363 gnd 0.002795f
C3259 vdd.n1364 gnd 0.002715f
C3260 vdd.n1365 gnd 0.013061f
C3261 vdd.n1366 gnd 0.008832f
C3262 vdd.n1367 gnd 0.103657f
C3263 vdd.n1368 gnd 0.005446f
C3264 vdd.n1369 gnd 0.005053f
C3265 vdd.n1370 gnd 0.002795f
C3266 vdd.n1371 gnd 0.006418f
C3267 vdd.n1372 gnd 0.002715f
C3268 vdd.n1373 gnd 0.002875f
C3269 vdd.n1374 gnd 0.005053f
C3270 vdd.n1375 gnd 0.002715f
C3271 vdd.n1376 gnd 0.006418f
C3272 vdd.n1377 gnd 0.002875f
C3273 vdd.n1378 gnd 0.005053f
C3274 vdd.n1379 gnd 0.002715f
C3275 vdd.n1380 gnd 0.004814f
C3276 vdd.n1381 gnd 0.004828f
C3277 vdd.t195 gnd 0.013789f
C3278 vdd.n1382 gnd 0.03068f
C3279 vdd.n1383 gnd 0.159666f
C3280 vdd.n1384 gnd 0.002715f
C3281 vdd.n1385 gnd 0.002875f
C3282 vdd.n1386 gnd 0.006418f
C3283 vdd.n1387 gnd 0.006418f
C3284 vdd.n1388 gnd 0.002875f
C3285 vdd.n1389 gnd 0.002715f
C3286 vdd.n1390 gnd 0.005053f
C3287 vdd.n1391 gnd 0.005053f
C3288 vdd.n1392 gnd 0.002715f
C3289 vdd.n1393 gnd 0.002875f
C3290 vdd.n1394 gnd 0.006418f
C3291 vdd.n1395 gnd 0.006418f
C3292 vdd.n1396 gnd 0.002875f
C3293 vdd.n1397 gnd 0.002715f
C3294 vdd.n1398 gnd 0.005053f
C3295 vdd.n1399 gnd 0.005053f
C3296 vdd.n1400 gnd 0.002715f
C3297 vdd.n1401 gnd 0.002875f
C3298 vdd.n1402 gnd 0.006418f
C3299 vdd.n1403 gnd 0.006418f
C3300 vdd.n1404 gnd 0.015174f
C3301 vdd.n1405 gnd 0.002795f
C3302 vdd.n1406 gnd 0.002715f
C3303 vdd.n1407 gnd 0.013061f
C3304 vdd.n1408 gnd 0.009118f
C3305 vdd.t231 gnd 0.031946f
C3306 vdd.t134 gnd 0.031946f
C3307 vdd.n1409 gnd 0.219551f
C3308 vdd.n1410 gnd 0.172644f
C3309 vdd.t207 gnd 0.031946f
C3310 vdd.t40 gnd 0.031946f
C3311 vdd.n1411 gnd 0.219551f
C3312 vdd.n1412 gnd 0.139322f
C3313 vdd.t212 gnd 0.031946f
C3314 vdd.t179 gnd 0.031946f
C3315 vdd.n1413 gnd 0.219551f
C3316 vdd.n1414 gnd 0.139322f
C3317 vdd.t33 gnd 0.031946f
C3318 vdd.t41 gnd 0.031946f
C3319 vdd.n1415 gnd 0.219551f
C3320 vdd.n1416 gnd 0.139322f
C3321 vdd.t49 gnd 0.031946f
C3322 vdd.t182 gnd 0.031946f
C3323 vdd.n1417 gnd 0.219551f
C3324 vdd.n1418 gnd 0.139322f
C3325 vdd.n1419 gnd 0.005446f
C3326 vdd.n1420 gnd 0.005053f
C3327 vdd.n1421 gnd 0.002795f
C3328 vdd.n1422 gnd 0.006418f
C3329 vdd.n1423 gnd 0.002715f
C3330 vdd.n1424 gnd 0.002875f
C3331 vdd.n1425 gnd 0.005053f
C3332 vdd.n1426 gnd 0.002715f
C3333 vdd.n1427 gnd 0.006418f
C3334 vdd.n1428 gnd 0.002875f
C3335 vdd.n1429 gnd 0.005053f
C3336 vdd.n1430 gnd 0.002715f
C3337 vdd.n1431 gnd 0.004814f
C3338 vdd.n1432 gnd 0.004828f
C3339 vdd.t47 gnd 0.013789f
C3340 vdd.n1433 gnd 0.03068f
C3341 vdd.n1434 gnd 0.159666f
C3342 vdd.n1435 gnd 0.002715f
C3343 vdd.n1436 gnd 0.002875f
C3344 vdd.n1437 gnd 0.006418f
C3345 vdd.n1438 gnd 0.006418f
C3346 vdd.n1439 gnd 0.002875f
C3347 vdd.n1440 gnd 0.002715f
C3348 vdd.n1441 gnd 0.005053f
C3349 vdd.n1442 gnd 0.005053f
C3350 vdd.n1443 gnd 0.002715f
C3351 vdd.n1444 gnd 0.002875f
C3352 vdd.n1445 gnd 0.006418f
C3353 vdd.n1446 gnd 0.006418f
C3354 vdd.n1447 gnd 0.002875f
C3355 vdd.n1448 gnd 0.002715f
C3356 vdd.n1449 gnd 0.005053f
C3357 vdd.n1450 gnd 0.005053f
C3358 vdd.n1451 gnd 0.002715f
C3359 vdd.n1452 gnd 0.002875f
C3360 vdd.n1453 gnd 0.006418f
C3361 vdd.n1454 gnd 0.006418f
C3362 vdd.n1455 gnd 0.015174f
C3363 vdd.n1456 gnd 0.002795f
C3364 vdd.n1457 gnd 0.002715f
C3365 vdd.n1458 gnd 0.013061f
C3366 vdd.n1459 gnd 0.008832f
C3367 vdd.n1460 gnd 0.061665f
C3368 vdd.n1461 gnd 0.222196f
C3369 vdd.n1462 gnd 0.005446f
C3370 vdd.n1463 gnd 0.005053f
C3371 vdd.n1464 gnd 0.002795f
C3372 vdd.n1465 gnd 0.006418f
C3373 vdd.n1466 gnd 0.002715f
C3374 vdd.n1467 gnd 0.002875f
C3375 vdd.n1468 gnd 0.005053f
C3376 vdd.n1469 gnd 0.002715f
C3377 vdd.n1470 gnd 0.006418f
C3378 vdd.n1471 gnd 0.002875f
C3379 vdd.n1472 gnd 0.005053f
C3380 vdd.n1473 gnd 0.002715f
C3381 vdd.n1474 gnd 0.004814f
C3382 vdd.n1475 gnd 0.004828f
C3383 vdd.t43 gnd 0.013789f
C3384 vdd.n1476 gnd 0.03068f
C3385 vdd.n1477 gnd 0.159666f
C3386 vdd.n1478 gnd 0.002715f
C3387 vdd.n1479 gnd 0.002875f
C3388 vdd.n1480 gnd 0.006418f
C3389 vdd.n1481 gnd 0.006418f
C3390 vdd.n1482 gnd 0.002875f
C3391 vdd.n1483 gnd 0.002715f
C3392 vdd.n1484 gnd 0.005053f
C3393 vdd.n1485 gnd 0.005053f
C3394 vdd.n1486 gnd 0.002715f
C3395 vdd.n1487 gnd 0.002875f
C3396 vdd.n1488 gnd 0.006418f
C3397 vdd.n1489 gnd 0.006418f
C3398 vdd.n1490 gnd 0.002875f
C3399 vdd.n1491 gnd 0.002715f
C3400 vdd.n1492 gnd 0.005053f
C3401 vdd.n1493 gnd 0.005053f
C3402 vdd.n1494 gnd 0.002715f
C3403 vdd.n1495 gnd 0.002875f
C3404 vdd.n1496 gnd 0.006418f
C3405 vdd.n1497 gnd 0.006418f
C3406 vdd.n1498 gnd 0.015174f
C3407 vdd.n1499 gnd 0.002795f
C3408 vdd.n1500 gnd 0.002715f
C3409 vdd.n1501 gnd 0.013061f
C3410 vdd.n1502 gnd 0.009118f
C3411 vdd.t216 gnd 0.031946f
C3412 vdd.t45 gnd 0.031946f
C3413 vdd.n1503 gnd 0.219551f
C3414 vdd.n1504 gnd 0.172644f
C3415 vdd.t31 gnd 0.031946f
C3416 vdd.t136 gnd 0.031946f
C3417 vdd.n1505 gnd 0.219551f
C3418 vdd.n1506 gnd 0.139322f
C3419 vdd.t209 gnd 0.031946f
C3420 vdd.t229 gnd 0.031946f
C3421 vdd.n1507 gnd 0.219551f
C3422 vdd.n1508 gnd 0.139322f
C3423 vdd.t191 gnd 0.031946f
C3424 vdd.t137 gnd 0.031946f
C3425 vdd.n1509 gnd 0.219551f
C3426 vdd.n1510 gnd 0.139322f
C3427 vdd.t203 gnd 0.031946f
C3428 vdd.t169 gnd 0.031946f
C3429 vdd.n1511 gnd 0.219551f
C3430 vdd.n1512 gnd 0.139322f
C3431 vdd.n1513 gnd 0.005446f
C3432 vdd.n1514 gnd 0.005053f
C3433 vdd.n1515 gnd 0.002795f
C3434 vdd.n1516 gnd 0.006418f
C3435 vdd.n1517 gnd 0.002715f
C3436 vdd.n1518 gnd 0.002875f
C3437 vdd.n1519 gnd 0.005053f
C3438 vdd.n1520 gnd 0.002715f
C3439 vdd.n1521 gnd 0.006418f
C3440 vdd.n1522 gnd 0.002875f
C3441 vdd.n1523 gnd 0.005053f
C3442 vdd.n1524 gnd 0.002715f
C3443 vdd.n1525 gnd 0.004814f
C3444 vdd.n1526 gnd 0.004828f
C3445 vdd.t202 gnd 0.013789f
C3446 vdd.n1527 gnd 0.03068f
C3447 vdd.n1528 gnd 0.159666f
C3448 vdd.n1529 gnd 0.002715f
C3449 vdd.n1530 gnd 0.002875f
C3450 vdd.n1531 gnd 0.006418f
C3451 vdd.n1532 gnd 0.006418f
C3452 vdd.n1533 gnd 0.002875f
C3453 vdd.n1534 gnd 0.002715f
C3454 vdd.n1535 gnd 0.005053f
C3455 vdd.n1536 gnd 0.005053f
C3456 vdd.n1537 gnd 0.002715f
C3457 vdd.n1538 gnd 0.002875f
C3458 vdd.n1539 gnd 0.006418f
C3459 vdd.n1540 gnd 0.006418f
C3460 vdd.n1541 gnd 0.002875f
C3461 vdd.n1542 gnd 0.002715f
C3462 vdd.n1543 gnd 0.005053f
C3463 vdd.n1544 gnd 0.005053f
C3464 vdd.n1545 gnd 0.002715f
C3465 vdd.n1546 gnd 0.002875f
C3466 vdd.n1547 gnd 0.006418f
C3467 vdd.n1548 gnd 0.006418f
C3468 vdd.n1549 gnd 0.015174f
C3469 vdd.n1550 gnd 0.002795f
C3470 vdd.n1551 gnd 0.002715f
C3471 vdd.n1552 gnd 0.013061f
C3472 vdd.n1553 gnd 0.008832f
C3473 vdd.n1554 gnd 0.061665f
C3474 vdd.n1555 gnd 0.244201f
C3475 vdd.n1556 gnd 2.19785f
C3476 vdd.n1557 gnd 0.590662f
C3477 vdd.n1558 gnd 0.009888f
C3478 vdd.n1559 gnd 0.009922f
C3479 vdd.n1560 gnd 0.007986f
C3480 vdd.n1561 gnd 0.009922f
C3481 vdd.n1562 gnd 0.806152f
C3482 vdd.n1563 gnd 0.009922f
C3483 vdd.n1564 gnd 0.007986f
C3484 vdd.n1565 gnd 0.009922f
C3485 vdd.n1566 gnd 0.009922f
C3486 vdd.n1567 gnd 0.009922f
C3487 vdd.n1568 gnd 0.007986f
C3488 vdd.n1569 gnd 0.009922f
C3489 vdd.n1570 gnd 0.841643f
C3490 vdd.t39 gnd 0.507014f
C3491 vdd.n1571 gnd 0.633767f
C3492 vdd.n1572 gnd 0.009922f
C3493 vdd.n1573 gnd 0.007986f
C3494 vdd.n1574 gnd 0.009922f
C3495 vdd.n1575 gnd 0.009922f
C3496 vdd.n1576 gnd 0.009922f
C3497 vdd.n1577 gnd 0.007986f
C3498 vdd.n1578 gnd 0.009922f
C3499 vdd.n1579 gnd 0.552645f
C3500 vdd.n1580 gnd 0.009922f
C3501 vdd.n1581 gnd 0.007986f
C3502 vdd.n1582 gnd 0.009922f
C3503 vdd.n1583 gnd 0.009922f
C3504 vdd.n1584 gnd 0.009922f
C3505 vdd.n1585 gnd 0.007986f
C3506 vdd.n1586 gnd 0.009922f
C3507 vdd.n1587 gnd 0.623627f
C3508 vdd.n1588 gnd 0.72503f
C3509 vdd.n1589 gnd 0.009922f
C3510 vdd.n1590 gnd 0.007986f
C3511 vdd.n1591 gnd 0.009922f
C3512 vdd.n1592 gnd 0.009922f
C3513 vdd.n1593 gnd 0.009922f
C3514 vdd.n1594 gnd 0.007986f
C3515 vdd.n1595 gnd 0.009922f
C3516 vdd.n1596 gnd 0.897415f
C3517 vdd.n1597 gnd 0.009922f
C3518 vdd.n1598 gnd 0.007986f
C3519 vdd.n1599 gnd 0.009922f
C3520 vdd.n1600 gnd 0.009922f
C3521 vdd.n1601 gnd 0.023383f
C3522 vdd.n1602 gnd 0.009922f
C3523 vdd.n1603 gnd 0.009922f
C3524 vdd.n1604 gnd 0.007986f
C3525 vdd.n1605 gnd 0.009922f
C3526 vdd.n1606 gnd 0.542505f
C3527 vdd.n1607 gnd 1.01403f
C3528 vdd.n1608 gnd 0.009922f
C3529 vdd.n1609 gnd 0.007986f
C3530 vdd.n1610 gnd 0.009922f
C3531 vdd.n1611 gnd 0.009922f
C3532 vdd.n1612 gnd 0.008533f
C3533 vdd.n1613 gnd 0.007986f
C3534 vdd.n1615 gnd 0.009922f
C3535 vdd.n1617 gnd 0.007986f
C3536 vdd.n1618 gnd 0.009922f
C3537 vdd.n1619 gnd 0.007986f
C3538 vdd.n1621 gnd 0.009922f
C3539 vdd.n1622 gnd 0.007986f
C3540 vdd.n1623 gnd 0.009922f
C3541 vdd.n1624 gnd 0.009922f
C3542 vdd.n1625 gnd 0.009922f
C3543 vdd.n1626 gnd 0.009922f
C3544 vdd.n1627 gnd 0.009922f
C3545 vdd.n1628 gnd 0.007986f
C3546 vdd.n1630 gnd 0.009922f
C3547 vdd.n1631 gnd 0.009922f
C3548 vdd.n1632 gnd 0.009922f
C3549 vdd.n1633 gnd 0.009922f
C3550 vdd.n1634 gnd 0.009922f
C3551 vdd.n1635 gnd 0.007986f
C3552 vdd.n1637 gnd 0.009922f
C3553 vdd.n1638 gnd 0.009922f
C3554 vdd.n1639 gnd 0.009922f
C3555 vdd.n1640 gnd 0.009922f
C3556 vdd.n1641 gnd 0.006669f
C3557 vdd.t81 gnd 0.122072f
C3558 vdd.t80 gnd 0.130462f
C3559 vdd.t79 gnd 0.159425f
C3560 vdd.n1642 gnd 0.20436f
C3561 vdd.n1643 gnd 0.171699f
C3562 vdd.n1645 gnd 0.009922f
C3563 vdd.n1646 gnd 0.009922f
C3564 vdd.n1647 gnd 0.007986f
C3565 vdd.n1648 gnd 0.009922f
C3566 vdd.n1650 gnd 0.009922f
C3567 vdd.n1651 gnd 0.009922f
C3568 vdd.n1652 gnd 0.009922f
C3569 vdd.n1653 gnd 0.009922f
C3570 vdd.n1654 gnd 0.007986f
C3571 vdd.n1656 gnd 0.009922f
C3572 vdd.n1657 gnd 0.009922f
C3573 vdd.n1658 gnd 0.009922f
C3574 vdd.n1659 gnd 0.009922f
C3575 vdd.n1660 gnd 0.009922f
C3576 vdd.n1661 gnd 0.007986f
C3577 vdd.n1663 gnd 0.009922f
C3578 vdd.n1664 gnd 0.009922f
C3579 vdd.n1665 gnd 0.009922f
C3580 vdd.n1666 gnd 0.009922f
C3581 vdd.n1667 gnd 0.009922f
C3582 vdd.n1668 gnd 0.007986f
C3583 vdd.n1670 gnd 0.009922f
C3584 vdd.n1671 gnd 0.009922f
C3585 vdd.n1672 gnd 0.009922f
C3586 vdd.n1673 gnd 0.009922f
C3587 vdd.n1674 gnd 0.009922f
C3588 vdd.n1675 gnd 0.007986f
C3589 vdd.n1677 gnd 0.009922f
C3590 vdd.n1678 gnd 0.009922f
C3591 vdd.n1679 gnd 0.009922f
C3592 vdd.n1680 gnd 0.009922f
C3593 vdd.n1681 gnd 0.007907f
C3594 vdd.t75 gnd 0.122072f
C3595 vdd.t74 gnd 0.130462f
C3596 vdd.t73 gnd 0.159425f
C3597 vdd.n1682 gnd 0.20436f
C3598 vdd.n1683 gnd 0.171699f
C3599 vdd.n1685 gnd 0.009922f
C3600 vdd.n1686 gnd 0.009922f
C3601 vdd.n1687 gnd 0.007986f
C3602 vdd.n1688 gnd 0.009922f
C3603 vdd.n1690 gnd 0.009922f
C3604 vdd.n1691 gnd 0.009922f
C3605 vdd.n1692 gnd 0.009922f
C3606 vdd.n1693 gnd 0.009922f
C3607 vdd.n1694 gnd 0.007986f
C3608 vdd.n1696 gnd 0.009922f
C3609 vdd.n1697 gnd 0.009922f
C3610 vdd.n1698 gnd 0.009922f
C3611 vdd.n1699 gnd 0.009922f
C3612 vdd.n1700 gnd 0.009922f
C3613 vdd.n1701 gnd 0.007986f
C3614 vdd.n1703 gnd 0.009922f
C3615 vdd.n1704 gnd 0.009922f
C3616 vdd.n1705 gnd 0.009922f
C3617 vdd.n1706 gnd 0.009922f
C3618 vdd.n1707 gnd 0.009922f
C3619 vdd.n1708 gnd 0.009922f
C3620 vdd.n1709 gnd 0.007986f
C3621 vdd.n1711 gnd 0.009922f
C3622 vdd.n1713 gnd 0.009922f
C3623 vdd.n1714 gnd 0.007986f
C3624 vdd.n1715 gnd 0.007986f
C3625 vdd.n1716 gnd 0.009922f
C3626 vdd.n1718 gnd 0.009922f
C3627 vdd.n1719 gnd 0.007986f
C3628 vdd.n1720 gnd 0.007986f
C3629 vdd.n1721 gnd 0.009922f
C3630 vdd.n1723 gnd 0.009922f
C3631 vdd.n1724 gnd 0.009922f
C3632 vdd.n1725 gnd 0.007986f
C3633 vdd.n1726 gnd 0.007986f
C3634 vdd.n1727 gnd 0.007986f
C3635 vdd.n1728 gnd 0.009922f
C3636 vdd.n1730 gnd 0.009922f
C3637 vdd.n1731 gnd 0.009922f
C3638 vdd.n1732 gnd 0.007986f
C3639 vdd.n1733 gnd 0.007986f
C3640 vdd.n1734 gnd 0.007986f
C3641 vdd.n1735 gnd 0.009922f
C3642 vdd.n1737 gnd 0.009922f
C3643 vdd.n1738 gnd 0.009922f
C3644 vdd.n1739 gnd 0.007986f
C3645 vdd.n1740 gnd 0.007986f
C3646 vdd.n1741 gnd 0.007986f
C3647 vdd.n1742 gnd 0.009922f
C3648 vdd.n1744 gnd 0.009922f
C3649 vdd.n1745 gnd 0.009922f
C3650 vdd.n1746 gnd 0.007986f
C3651 vdd.n1747 gnd 0.009922f
C3652 vdd.n1748 gnd 0.009922f
C3653 vdd.n1749 gnd 0.009922f
C3654 vdd.n1750 gnd 0.016292f
C3655 vdd.n1751 gnd 0.005431f
C3656 vdd.n1752 gnd 0.007986f
C3657 vdd.n1753 gnd 0.009922f
C3658 vdd.n1755 gnd 0.009922f
C3659 vdd.n1756 gnd 0.009922f
C3660 vdd.n1757 gnd 0.007986f
C3661 vdd.n1758 gnd 0.007986f
C3662 vdd.n1759 gnd 0.007986f
C3663 vdd.n1760 gnd 0.009922f
C3664 vdd.n1762 gnd 0.009922f
C3665 vdd.n1763 gnd 0.009922f
C3666 vdd.n1764 gnd 0.007986f
C3667 vdd.n1765 gnd 0.007986f
C3668 vdd.n1766 gnd 0.007986f
C3669 vdd.n1767 gnd 0.009922f
C3670 vdd.n1769 gnd 0.009922f
C3671 vdd.n1770 gnd 0.009922f
C3672 vdd.n1771 gnd 0.007986f
C3673 vdd.n1772 gnd 0.007986f
C3674 vdd.n1773 gnd 0.007986f
C3675 vdd.n1774 gnd 0.009922f
C3676 vdd.n1776 gnd 0.009922f
C3677 vdd.n1777 gnd 0.009922f
C3678 vdd.n1778 gnd 0.007986f
C3679 vdd.n1779 gnd 0.007986f
C3680 vdd.n1780 gnd 0.007986f
C3681 vdd.n1781 gnd 0.009922f
C3682 vdd.n1783 gnd 0.009922f
C3683 vdd.n1784 gnd 0.009922f
C3684 vdd.n1785 gnd 0.007986f
C3685 vdd.n1786 gnd 0.009922f
C3686 vdd.n1787 gnd 0.009922f
C3687 vdd.n1788 gnd 0.009922f
C3688 vdd.n1789 gnd 0.016292f
C3689 vdd.n1790 gnd 0.006669f
C3690 vdd.n1791 gnd 0.007986f
C3691 vdd.n1792 gnd 0.009922f
C3692 vdd.n1794 gnd 0.009922f
C3693 vdd.n1795 gnd 0.009922f
C3694 vdd.n1796 gnd 0.007986f
C3695 vdd.n1797 gnd 0.007986f
C3696 vdd.n1798 gnd 0.007986f
C3697 vdd.n1799 gnd 0.009922f
C3698 vdd.n1801 gnd 0.009922f
C3699 vdd.n1802 gnd 0.009922f
C3700 vdd.n1803 gnd 0.007986f
C3701 vdd.n1804 gnd 0.007986f
C3702 vdd.n1805 gnd 0.007986f
C3703 vdd.n1806 gnd 0.009922f
C3704 vdd.n1808 gnd 0.009922f
C3705 vdd.n1809 gnd 0.009922f
C3706 vdd.n1811 gnd 0.009922f
C3707 vdd.n1812 gnd 0.007986f
C3708 vdd.n1813 gnd 0.00635f
C3709 vdd.n1814 gnd 0.006747f
C3710 vdd.n1815 gnd 0.006747f
C3711 vdd.n1816 gnd 0.006747f
C3712 vdd.n1817 gnd 0.006747f
C3713 vdd.n1818 gnd 0.006747f
C3714 vdd.n1819 gnd 0.006747f
C3715 vdd.n1820 gnd 0.006747f
C3716 vdd.n1821 gnd 0.006747f
C3717 vdd.n1823 gnd 0.006747f
C3718 vdd.n1824 gnd 0.006747f
C3719 vdd.n1825 gnd 0.006747f
C3720 vdd.n1826 gnd 0.006747f
C3721 vdd.n1827 gnd 0.006747f
C3722 vdd.n1829 gnd 0.006747f
C3723 vdd.n1831 gnd 0.006747f
C3724 vdd.n1832 gnd 0.006747f
C3725 vdd.n1833 gnd 0.006747f
C3726 vdd.n1834 gnd 0.006747f
C3727 vdd.n1835 gnd 0.006747f
C3728 vdd.n1837 gnd 0.006747f
C3729 vdd.n1839 gnd 0.006747f
C3730 vdd.n1840 gnd 0.006747f
C3731 vdd.n1841 gnd 0.006747f
C3732 vdd.n1842 gnd 0.006747f
C3733 vdd.n1843 gnd 0.006747f
C3734 vdd.n1845 gnd 0.006747f
C3735 vdd.n1847 gnd 0.006747f
C3736 vdd.n1848 gnd 0.006747f
C3737 vdd.n1849 gnd 0.006747f
C3738 vdd.n1850 gnd 0.006747f
C3739 vdd.n1851 gnd 0.006747f
C3740 vdd.n1853 gnd 0.006747f
C3741 vdd.n1854 gnd 0.006747f
C3742 vdd.n1855 gnd 0.006747f
C3743 vdd.n1856 gnd 0.006747f
C3744 vdd.n1857 gnd 0.006747f
C3745 vdd.n1858 gnd 0.006747f
C3746 vdd.n1859 gnd 0.006747f
C3747 vdd.n1860 gnd 0.006747f
C3748 vdd.n1861 gnd 0.004912f
C3749 vdd.n1862 gnd 0.006747f
C3750 vdd.t125 gnd 0.272656f
C3751 vdd.t126 gnd 0.279098f
C3752 vdd.t124 gnd 0.178f
C3753 vdd.n1863 gnd 0.096199f
C3754 vdd.n1864 gnd 0.054567f
C3755 vdd.n1865 gnd 0.009643f
C3756 vdd.n1866 gnd 0.006747f
C3757 vdd.n1867 gnd 0.006747f
C3758 vdd.n1868 gnd 0.410681f
C3759 vdd.n1869 gnd 0.006747f
C3760 vdd.n1870 gnd 0.006747f
C3761 vdd.n1871 gnd 0.006747f
C3762 vdd.n1872 gnd 0.006747f
C3763 vdd.n1873 gnd 0.006747f
C3764 vdd.n1874 gnd 0.006747f
C3765 vdd.n1875 gnd 0.006747f
C3766 vdd.n1876 gnd 0.006747f
C3767 vdd.n1877 gnd 0.006747f
C3768 vdd.n1878 gnd 0.006747f
C3769 vdd.n1879 gnd 0.006747f
C3770 vdd.n1880 gnd 0.006747f
C3771 vdd.n1881 gnd 0.006747f
C3772 vdd.n1882 gnd 0.006747f
C3773 vdd.n1883 gnd 0.006747f
C3774 vdd.n1884 gnd 0.006747f
C3775 vdd.n1885 gnd 0.006747f
C3776 vdd.n1886 gnd 0.006747f
C3777 vdd.n1887 gnd 0.006747f
C3778 vdd.n1888 gnd 0.006747f
C3779 vdd.t99 gnd 0.272656f
C3780 vdd.t100 gnd 0.279098f
C3781 vdd.t97 gnd 0.178f
C3782 vdd.n1889 gnd 0.096199f
C3783 vdd.n1890 gnd 0.054567f
C3784 vdd.n1891 gnd 0.006747f
C3785 vdd.n1892 gnd 0.006747f
C3786 vdd.n1893 gnd 0.006747f
C3787 vdd.n1894 gnd 0.006747f
C3788 vdd.n1895 gnd 0.006747f
C3789 vdd.n1896 gnd 0.006747f
C3790 vdd.n1898 gnd 0.006747f
C3791 vdd.n1899 gnd 0.006747f
C3792 vdd.n1900 gnd 0.006747f
C3793 vdd.n1901 gnd 0.006747f
C3794 vdd.n1903 gnd 0.006747f
C3795 vdd.n1905 gnd 0.006747f
C3796 vdd.n1906 gnd 0.006747f
C3797 vdd.n1907 gnd 0.006747f
C3798 vdd.n1908 gnd 0.006747f
C3799 vdd.n1909 gnd 0.006747f
C3800 vdd.n1911 gnd 0.006747f
C3801 vdd.n1913 gnd 0.006747f
C3802 vdd.n1914 gnd 0.006747f
C3803 vdd.n1915 gnd 0.006747f
C3804 vdd.n1916 gnd 0.006747f
C3805 vdd.n1917 gnd 0.006747f
C3806 vdd.n1919 gnd 0.006747f
C3807 vdd.n1921 gnd 0.006747f
C3808 vdd.n1922 gnd 0.006747f
C3809 vdd.n1923 gnd 0.004912f
C3810 vdd.n1924 gnd 0.009643f
C3811 vdd.n1925 gnd 0.005209f
C3812 vdd.n1926 gnd 0.006747f
C3813 vdd.n1928 gnd 0.006747f
C3814 vdd.n1929 gnd 0.01601f
C3815 vdd.n1930 gnd 0.01601f
C3816 vdd.n1931 gnd 0.014948f
C3817 vdd.n1932 gnd 0.006747f
C3818 vdd.n1933 gnd 0.006747f
C3819 vdd.n1934 gnd 0.006747f
C3820 vdd.n1935 gnd 0.006747f
C3821 vdd.n1936 gnd 0.006747f
C3822 vdd.n1937 gnd 0.006747f
C3823 vdd.n1938 gnd 0.006747f
C3824 vdd.n1939 gnd 0.006747f
C3825 vdd.n1940 gnd 0.006747f
C3826 vdd.n1941 gnd 0.006747f
C3827 vdd.n1942 gnd 0.006747f
C3828 vdd.n1943 gnd 0.006747f
C3829 vdd.n1944 gnd 0.006747f
C3830 vdd.n1945 gnd 0.006747f
C3831 vdd.n1946 gnd 0.006747f
C3832 vdd.n1947 gnd 0.006747f
C3833 vdd.n1948 gnd 0.006747f
C3834 vdd.n1949 gnd 0.006747f
C3835 vdd.n1950 gnd 0.006747f
C3836 vdd.n1951 gnd 0.006747f
C3837 vdd.n1952 gnd 0.006747f
C3838 vdd.n1953 gnd 0.006747f
C3839 vdd.n1954 gnd 0.006747f
C3840 vdd.n1955 gnd 0.006747f
C3841 vdd.n1956 gnd 0.006747f
C3842 vdd.n1957 gnd 0.006747f
C3843 vdd.n1958 gnd 0.006747f
C3844 vdd.n1959 gnd 0.006747f
C3845 vdd.n1960 gnd 0.006747f
C3846 vdd.n1961 gnd 0.006747f
C3847 vdd.n1962 gnd 0.006747f
C3848 vdd.n1963 gnd 0.006747f
C3849 vdd.n1964 gnd 0.006747f
C3850 vdd.n1965 gnd 0.006747f
C3851 vdd.n1966 gnd 0.006747f
C3852 vdd.n1967 gnd 0.006747f
C3853 vdd.n1968 gnd 0.006747f
C3854 vdd.n1969 gnd 0.218016f
C3855 vdd.n1970 gnd 0.006747f
C3856 vdd.n1971 gnd 0.006747f
C3857 vdd.n1972 gnd 0.006747f
C3858 vdd.n1973 gnd 0.006747f
C3859 vdd.n1974 gnd 0.006747f
C3860 vdd.n1975 gnd 0.006747f
C3861 vdd.n1976 gnd 0.006747f
C3862 vdd.n1977 gnd 0.006747f
C3863 vdd.n1978 gnd 0.006747f
C3864 vdd.n1979 gnd 0.006747f
C3865 vdd.n1980 gnd 0.006747f
C3866 vdd.n1981 gnd 0.006747f
C3867 vdd.n1982 gnd 0.006747f
C3868 vdd.n1983 gnd 0.006747f
C3869 vdd.n1984 gnd 0.006747f
C3870 vdd.n1985 gnd 0.006747f
C3871 vdd.n1986 gnd 0.006747f
C3872 vdd.n1987 gnd 0.006747f
C3873 vdd.n1988 gnd 0.006747f
C3874 vdd.n1989 gnd 0.006747f
C3875 vdd.n1990 gnd 0.014948f
C3876 vdd.n1992 gnd 0.01601f
C3877 vdd.n1993 gnd 0.01601f
C3878 vdd.n1994 gnd 0.006747f
C3879 vdd.n1995 gnd 0.005209f
C3880 vdd.n1996 gnd 0.006747f
C3881 vdd.n1998 gnd 0.006747f
C3882 vdd.n2000 gnd 0.006747f
C3883 vdd.n2001 gnd 0.006747f
C3884 vdd.n2002 gnd 0.006747f
C3885 vdd.n2003 gnd 0.006747f
C3886 vdd.n2004 gnd 0.006747f
C3887 vdd.n2006 gnd 0.006747f
C3888 vdd.n2008 gnd 0.006747f
C3889 vdd.n2009 gnd 0.006747f
C3890 vdd.n2010 gnd 0.006747f
C3891 vdd.n2011 gnd 0.006747f
C3892 vdd.n2012 gnd 0.006747f
C3893 vdd.n2014 gnd 0.006747f
C3894 vdd.n2016 gnd 0.006747f
C3895 vdd.n2017 gnd 0.006747f
C3896 vdd.n2018 gnd 0.006747f
C3897 vdd.n2019 gnd 0.006747f
C3898 vdd.n2020 gnd 0.006747f
C3899 vdd.n2022 gnd 0.006747f
C3900 vdd.n2024 gnd 0.006747f
C3901 vdd.n2025 gnd 0.006747f
C3902 vdd.n2026 gnd 0.020126f
C3903 vdd.n2027 gnd 0.596611f
C3904 vdd.n2029 gnd 0.007986f
C3905 vdd.n2030 gnd 0.007986f
C3906 vdd.n2031 gnd 0.009922f
C3907 vdd.n2033 gnd 0.009922f
C3908 vdd.n2034 gnd 0.009922f
C3909 vdd.n2035 gnd 0.007986f
C3910 vdd.n2036 gnd 0.006629f
C3911 vdd.n2037 gnd 0.023749f
C3912 vdd.n2038 gnd 0.023383f
C3913 vdd.n2039 gnd 0.006629f
C3914 vdd.n2040 gnd 0.023383f
C3915 vdd.n2041 gnd 1.39429f
C3916 vdd.n2042 gnd 0.023383f
C3917 vdd.n2043 gnd 0.023749f
C3918 vdd.n2044 gnd 0.003794f
C3919 vdd.t64 gnd 0.122072f
C3920 vdd.t63 gnd 0.130462f
C3921 vdd.t61 gnd 0.159425f
C3922 vdd.n2045 gnd 0.20436f
C3923 vdd.n2046 gnd 0.171699f
C3924 vdd.n2047 gnd 0.012299f
C3925 vdd.n2048 gnd 0.004193f
C3926 vdd.n2049 gnd 0.008533f
C3927 vdd.n2050 gnd 0.596611f
C3928 vdd.n2051 gnd 0.020126f
C3929 vdd.n2052 gnd 0.006747f
C3930 vdd.n2053 gnd 0.006747f
C3931 vdd.n2054 gnd 0.006747f
C3932 vdd.n2056 gnd 0.006747f
C3933 vdd.n2058 gnd 0.006747f
C3934 vdd.n2059 gnd 0.006747f
C3935 vdd.n2060 gnd 0.006747f
C3936 vdd.n2061 gnd 0.006747f
C3937 vdd.n2062 gnd 0.006747f
C3938 vdd.n2064 gnd 0.006747f
C3939 vdd.n2066 gnd 0.006747f
C3940 vdd.n2067 gnd 0.006747f
C3941 vdd.n2068 gnd 0.006747f
C3942 vdd.n2069 gnd 0.006747f
C3943 vdd.n2070 gnd 0.006747f
C3944 vdd.n2072 gnd 0.006747f
C3945 vdd.n2074 gnd 0.006747f
C3946 vdd.n2075 gnd 0.006747f
C3947 vdd.n2076 gnd 0.006747f
C3948 vdd.n2077 gnd 0.006747f
C3949 vdd.n2078 gnd 0.006747f
C3950 vdd.n2080 gnd 0.006747f
C3951 vdd.n2082 gnd 0.006747f
C3952 vdd.n2083 gnd 0.006747f
C3953 vdd.n2084 gnd 0.01601f
C3954 vdd.n2085 gnd 0.014948f
C3955 vdd.n2086 gnd 0.014948f
C3956 vdd.n2087 gnd 0.993747f
C3957 vdd.n2088 gnd 0.014948f
C3958 vdd.n2089 gnd 0.014948f
C3959 vdd.n2090 gnd 0.006747f
C3960 vdd.n2091 gnd 0.006747f
C3961 vdd.n2092 gnd 0.006747f
C3962 vdd.n2093 gnd 0.430962f
C3963 vdd.n2094 gnd 0.006747f
C3964 vdd.n2095 gnd 0.006747f
C3965 vdd.n2096 gnd 0.006747f
C3966 vdd.n2097 gnd 0.006747f
C3967 vdd.n2098 gnd 0.006747f
C3968 vdd.n2099 gnd 0.689539f
C3969 vdd.n2100 gnd 0.006747f
C3970 vdd.n2101 gnd 0.006747f
C3971 vdd.n2102 gnd 0.006747f
C3972 vdd.n2103 gnd 0.006747f
C3973 vdd.n2104 gnd 0.006747f
C3974 vdd.n2105 gnd 0.689539f
C3975 vdd.n2106 gnd 0.006747f
C3976 vdd.n2107 gnd 0.006747f
C3977 vdd.n2108 gnd 0.005953f
C3978 vdd.n2109 gnd 0.019546f
C3979 vdd.n2110 gnd 0.004167f
C3980 vdd.n2111 gnd 0.006747f
C3981 vdd.n2112 gnd 0.38026f
C3982 vdd.n2113 gnd 0.006747f
C3983 vdd.n2114 gnd 0.006747f
C3984 vdd.n2115 gnd 0.006747f
C3985 vdd.n2116 gnd 0.006747f
C3986 vdd.n2117 gnd 0.006747f
C3987 vdd.n2118 gnd 0.461383f
C3988 vdd.n2119 gnd 0.006747f
C3989 vdd.n2120 gnd 0.006747f
C3990 vdd.n2121 gnd 0.006747f
C3991 vdd.n2122 gnd 0.006747f
C3992 vdd.n2123 gnd 0.006747f
C3993 vdd.n2124 gnd 0.613487f
C3994 vdd.n2125 gnd 0.006747f
C3995 vdd.n2126 gnd 0.006747f
C3996 vdd.n2127 gnd 0.006747f
C3997 vdd.n2128 gnd 0.006747f
C3998 vdd.n2129 gnd 0.006747f
C3999 vdd.n2130 gnd 0.547575f
C4000 vdd.n2131 gnd 0.006747f
C4001 vdd.n2132 gnd 0.006747f
C4002 vdd.n2133 gnd 0.006747f
C4003 vdd.n2134 gnd 0.006747f
C4004 vdd.n2135 gnd 0.006747f
C4005 vdd.n2136 gnd 0.395471f
C4006 vdd.n2137 gnd 0.006747f
C4007 vdd.n2138 gnd 0.006747f
C4008 vdd.n2139 gnd 0.006747f
C4009 vdd.n2140 gnd 0.006747f
C4010 vdd.n2141 gnd 0.006747f
C4011 vdd.n2142 gnd 0.218016f
C4012 vdd.n2143 gnd 0.006747f
C4013 vdd.n2144 gnd 0.006747f
C4014 vdd.n2145 gnd 0.006747f
C4015 vdd.n2146 gnd 0.006747f
C4016 vdd.n2147 gnd 0.006747f
C4017 vdd.n2148 gnd 0.38026f
C4018 vdd.n2149 gnd 0.006747f
C4019 vdd.n2150 gnd 0.006747f
C4020 vdd.n2151 gnd 0.006747f
C4021 vdd.n2152 gnd 0.006747f
C4022 vdd.n2153 gnd 0.006747f
C4023 vdd.n2154 gnd 0.689539f
C4024 vdd.n2155 gnd 0.006747f
C4025 vdd.n2156 gnd 0.006747f
C4026 vdd.n2157 gnd 0.006747f
C4027 vdd.n2158 gnd 0.006747f
C4028 vdd.n2159 gnd 0.006747f
C4029 vdd.n2160 gnd 0.006747f
C4030 vdd.n2161 gnd 0.006747f
C4031 vdd.n2162 gnd 0.537435f
C4032 vdd.n2163 gnd 0.006747f
C4033 vdd.n2164 gnd 0.006747f
C4034 vdd.n2165 gnd 0.006747f
C4035 vdd.n2166 gnd 0.006747f
C4036 vdd.n2167 gnd 0.006747f
C4037 vdd.n2168 gnd 0.006747f
C4038 vdd.n2169 gnd 0.430962f
C4039 vdd.n2170 gnd 0.006747f
C4040 vdd.n2171 gnd 0.006747f
C4041 vdd.n2172 gnd 0.006747f
C4042 vdd.n2173 gnd 0.01577f
C4043 vdd.n2174 gnd 0.015189f
C4044 vdd.n2175 gnd 0.006747f
C4045 vdd.n2176 gnd 0.006747f
C4046 vdd.n2177 gnd 0.005209f
C4047 vdd.n2178 gnd 0.006747f
C4048 vdd.n2179 gnd 0.006747f
C4049 vdd.n2180 gnd 0.004912f
C4050 vdd.n2181 gnd 0.006747f
C4051 vdd.n2182 gnd 0.006747f
C4052 vdd.n2183 gnd 0.006747f
C4053 vdd.n2184 gnd 0.006747f
C4054 vdd.n2185 gnd 0.006747f
C4055 vdd.n2186 gnd 0.006747f
C4056 vdd.n2187 gnd 0.006747f
C4057 vdd.n2188 gnd 0.006747f
C4058 vdd.n2189 gnd 0.006747f
C4059 vdd.n2190 gnd 0.006747f
C4060 vdd.n2191 gnd 0.006747f
C4061 vdd.n2192 gnd 0.006747f
C4062 vdd.n2193 gnd 0.006747f
C4063 vdd.n2194 gnd 0.006747f
C4064 vdd.n2195 gnd 0.006747f
C4065 vdd.n2196 gnd 0.006747f
C4066 vdd.n2197 gnd 0.006747f
C4067 vdd.n2198 gnd 0.006747f
C4068 vdd.n2199 gnd 0.006747f
C4069 vdd.n2200 gnd 0.006747f
C4070 vdd.n2201 gnd 0.006747f
C4071 vdd.n2202 gnd 0.006747f
C4072 vdd.n2203 gnd 0.006747f
C4073 vdd.n2204 gnd 0.006747f
C4074 vdd.n2205 gnd 0.006747f
C4075 vdd.n2206 gnd 0.006747f
C4076 vdd.n2207 gnd 0.006747f
C4077 vdd.n2208 gnd 0.006747f
C4078 vdd.n2209 gnd 0.006747f
C4079 vdd.n2210 gnd 0.006747f
C4080 vdd.n2211 gnd 0.006747f
C4081 vdd.n2212 gnd 0.006747f
C4082 vdd.n2213 gnd 0.006747f
C4083 vdd.n2214 gnd 0.006747f
C4084 vdd.n2215 gnd 0.006747f
C4085 vdd.n2216 gnd 0.006747f
C4086 vdd.n2217 gnd 0.006747f
C4087 vdd.n2218 gnd 0.006747f
C4088 vdd.n2219 gnd 0.006747f
C4089 vdd.n2220 gnd 0.006747f
C4090 vdd.n2221 gnd 0.006747f
C4091 vdd.n2222 gnd 0.006747f
C4092 vdd.n2223 gnd 0.006747f
C4093 vdd.n2224 gnd 0.006747f
C4094 vdd.n2225 gnd 0.006747f
C4095 vdd.n2226 gnd 0.006747f
C4096 vdd.n2227 gnd 0.006747f
C4097 vdd.n2228 gnd 0.006747f
C4098 vdd.n2229 gnd 0.006747f
C4099 vdd.n2230 gnd 0.006747f
C4100 vdd.n2231 gnd 0.006747f
C4101 vdd.n2232 gnd 0.006747f
C4102 vdd.n2233 gnd 0.006747f
C4103 vdd.n2234 gnd 0.006747f
C4104 vdd.n2235 gnd 0.006747f
C4105 vdd.n2236 gnd 0.006747f
C4106 vdd.n2237 gnd 0.006747f
C4107 vdd.n2238 gnd 0.006747f
C4108 vdd.n2239 gnd 0.006747f
C4109 vdd.n2240 gnd 0.006747f
C4110 vdd.n2241 gnd 0.01601f
C4111 vdd.n2242 gnd 0.014948f
C4112 vdd.n2243 gnd 0.014948f
C4113 vdd.n2244 gnd 0.841643f
C4114 vdd.n2245 gnd 0.014948f
C4115 vdd.n2246 gnd 0.01601f
C4116 vdd.n2247 gnd 0.015189f
C4117 vdd.n2248 gnd 0.006747f
C4118 vdd.n2249 gnd 0.006747f
C4119 vdd.n2250 gnd 0.006747f
C4120 vdd.n2251 gnd 0.005209f
C4121 vdd.n2252 gnd 0.009643f
C4122 vdd.n2253 gnd 0.004912f
C4123 vdd.n2254 gnd 0.006747f
C4124 vdd.n2255 gnd 0.006747f
C4125 vdd.n2256 gnd 0.006747f
C4126 vdd.n2257 gnd 0.006747f
C4127 vdd.n2258 gnd 0.006747f
C4128 vdd.n2259 gnd 0.006747f
C4129 vdd.n2260 gnd 0.006747f
C4130 vdd.n2261 gnd 0.006747f
C4131 vdd.n2262 gnd 0.006747f
C4132 vdd.n2263 gnd 0.006747f
C4133 vdd.n2264 gnd 0.006747f
C4134 vdd.n2265 gnd 0.006747f
C4135 vdd.n2266 gnd 0.006747f
C4136 vdd.n2267 gnd 0.006747f
C4137 vdd.n2268 gnd 0.006747f
C4138 vdd.n2269 gnd 0.006747f
C4139 vdd.n2270 gnd 0.006747f
C4140 vdd.n2271 gnd 0.006747f
C4141 vdd.n2272 gnd 0.006747f
C4142 vdd.n2273 gnd 0.006747f
C4143 vdd.n2274 gnd 0.006747f
C4144 vdd.n2275 gnd 0.006747f
C4145 vdd.n2276 gnd 0.006747f
C4146 vdd.n2277 gnd 0.006747f
C4147 vdd.n2278 gnd 0.006747f
C4148 vdd.n2279 gnd 0.006747f
C4149 vdd.n2280 gnd 0.006747f
C4150 vdd.n2281 gnd 0.006747f
C4151 vdd.n2282 gnd 0.006747f
C4152 vdd.n2283 gnd 0.006747f
C4153 vdd.n2284 gnd 0.006747f
C4154 vdd.n2285 gnd 0.006747f
C4155 vdd.n2286 gnd 0.006747f
C4156 vdd.n2287 gnd 0.006747f
C4157 vdd.n2288 gnd 0.006747f
C4158 vdd.n2289 gnd 0.006747f
C4159 vdd.n2290 gnd 0.006747f
C4160 vdd.n2291 gnd 0.006747f
C4161 vdd.n2292 gnd 0.006747f
C4162 vdd.n2293 gnd 0.006747f
C4163 vdd.n2294 gnd 0.006747f
C4164 vdd.n2295 gnd 0.006747f
C4165 vdd.n2296 gnd 0.006747f
C4166 vdd.n2297 gnd 0.006747f
C4167 vdd.n2298 gnd 0.006747f
C4168 vdd.n2299 gnd 0.006747f
C4169 vdd.n2300 gnd 0.006747f
C4170 vdd.n2301 gnd 0.006747f
C4171 vdd.n2302 gnd 0.006747f
C4172 vdd.n2303 gnd 0.006747f
C4173 vdd.n2304 gnd 0.006747f
C4174 vdd.n2305 gnd 0.006747f
C4175 vdd.n2306 gnd 0.006747f
C4176 vdd.n2307 gnd 0.006747f
C4177 vdd.n2308 gnd 0.006747f
C4178 vdd.n2309 gnd 0.006747f
C4179 vdd.n2310 gnd 0.006747f
C4180 vdd.n2311 gnd 0.006747f
C4181 vdd.n2312 gnd 0.006747f
C4182 vdd.n2313 gnd 0.006747f
C4183 vdd.n2314 gnd 0.01601f
C4184 vdd.n2315 gnd 0.01601f
C4185 vdd.n2316 gnd 0.841643f
C4186 vdd.t17 gnd 2.99138f
C4187 vdd.t200 gnd 2.99138f
C4188 vdd.n2349 gnd 0.01601f
C4189 vdd.n2350 gnd 0.006747f
C4190 vdd.t92 gnd 0.272656f
C4191 vdd.t93 gnd 0.279098f
C4192 vdd.t90 gnd 0.178f
C4193 vdd.n2351 gnd 0.096199f
C4194 vdd.n2352 gnd 0.054567f
C4195 vdd.n2353 gnd 0.006747f
C4196 vdd.t106 gnd 0.272656f
C4197 vdd.t107 gnd 0.279098f
C4198 vdd.t105 gnd 0.178f
C4199 vdd.n2354 gnd 0.096199f
C4200 vdd.n2355 gnd 0.054567f
C4201 vdd.n2356 gnd 0.009643f
C4202 vdd.n2357 gnd 0.006747f
C4203 vdd.n2358 gnd 0.006747f
C4204 vdd.n2359 gnd 0.006747f
C4205 vdd.n2360 gnd 0.006747f
C4206 vdd.n2361 gnd 0.006747f
C4207 vdd.n2362 gnd 0.006747f
C4208 vdd.n2363 gnd 0.006747f
C4209 vdd.n2364 gnd 0.006747f
C4210 vdd.n2365 gnd 0.006747f
C4211 vdd.n2366 gnd 0.006747f
C4212 vdd.n2367 gnd 0.006747f
C4213 vdd.n2368 gnd 0.006747f
C4214 vdd.n2369 gnd 0.006747f
C4215 vdd.n2370 gnd 0.006747f
C4216 vdd.n2371 gnd 0.006747f
C4217 vdd.n2372 gnd 0.006747f
C4218 vdd.n2373 gnd 0.006747f
C4219 vdd.n2374 gnd 0.006747f
C4220 vdd.n2375 gnd 0.006747f
C4221 vdd.n2376 gnd 0.006747f
C4222 vdd.n2377 gnd 0.006747f
C4223 vdd.n2378 gnd 0.006747f
C4224 vdd.n2379 gnd 0.006747f
C4225 vdd.n2380 gnd 0.006747f
C4226 vdd.n2381 gnd 0.006747f
C4227 vdd.n2382 gnd 0.006747f
C4228 vdd.n2383 gnd 0.006747f
C4229 vdd.n2384 gnd 0.006747f
C4230 vdd.n2385 gnd 0.006747f
C4231 vdd.n2386 gnd 0.006747f
C4232 vdd.n2387 gnd 0.006747f
C4233 vdd.n2388 gnd 0.006747f
C4234 vdd.n2389 gnd 0.006747f
C4235 vdd.n2390 gnd 0.006747f
C4236 vdd.n2391 gnd 0.006747f
C4237 vdd.n2392 gnd 0.006747f
C4238 vdd.n2393 gnd 0.006747f
C4239 vdd.n2394 gnd 0.006747f
C4240 vdd.n2395 gnd 0.006747f
C4241 vdd.n2396 gnd 0.006747f
C4242 vdd.n2397 gnd 0.006747f
C4243 vdd.n2398 gnd 0.006747f
C4244 vdd.n2399 gnd 0.006747f
C4245 vdd.n2400 gnd 0.006747f
C4246 vdd.n2401 gnd 0.006747f
C4247 vdd.n2402 gnd 0.006747f
C4248 vdd.n2403 gnd 0.006747f
C4249 vdd.n2404 gnd 0.006747f
C4250 vdd.n2405 gnd 0.006747f
C4251 vdd.n2406 gnd 0.006747f
C4252 vdd.n2407 gnd 0.006747f
C4253 vdd.n2408 gnd 0.006747f
C4254 vdd.n2409 gnd 0.006747f
C4255 vdd.n2410 gnd 0.006747f
C4256 vdd.n2411 gnd 0.006747f
C4257 vdd.n2412 gnd 0.006747f
C4258 vdd.n2413 gnd 0.004912f
C4259 vdd.n2414 gnd 0.006747f
C4260 vdd.n2415 gnd 0.006747f
C4261 vdd.n2416 gnd 0.005209f
C4262 vdd.n2417 gnd 0.006747f
C4263 vdd.n2418 gnd 0.006747f
C4264 vdd.n2419 gnd 0.01601f
C4265 vdd.n2420 gnd 0.014948f
C4266 vdd.n2421 gnd 0.006747f
C4267 vdd.n2422 gnd 0.006747f
C4268 vdd.n2423 gnd 0.006747f
C4269 vdd.n2424 gnd 0.006747f
C4270 vdd.n2425 gnd 0.006747f
C4271 vdd.n2426 gnd 0.006747f
C4272 vdd.n2427 gnd 0.006747f
C4273 vdd.n2428 gnd 0.006747f
C4274 vdd.n2429 gnd 0.006747f
C4275 vdd.n2430 gnd 0.006747f
C4276 vdd.n2431 gnd 0.006747f
C4277 vdd.n2432 gnd 0.006747f
C4278 vdd.n2433 gnd 0.006747f
C4279 vdd.n2434 gnd 0.006747f
C4280 vdd.n2435 gnd 0.006747f
C4281 vdd.n2436 gnd 0.006747f
C4282 vdd.n2437 gnd 0.006747f
C4283 vdd.n2438 gnd 0.006747f
C4284 vdd.n2439 gnd 0.006747f
C4285 vdd.n2440 gnd 0.006747f
C4286 vdd.n2441 gnd 0.006747f
C4287 vdd.n2442 gnd 0.006747f
C4288 vdd.n2443 gnd 0.006747f
C4289 vdd.n2444 gnd 0.006747f
C4290 vdd.n2445 gnd 0.006747f
C4291 vdd.n2446 gnd 0.006747f
C4292 vdd.n2447 gnd 0.006747f
C4293 vdd.n2448 gnd 0.006747f
C4294 vdd.n2449 gnd 0.006747f
C4295 vdd.n2450 gnd 0.006747f
C4296 vdd.n2451 gnd 0.006747f
C4297 vdd.n2452 gnd 0.006747f
C4298 vdd.n2453 gnd 0.006747f
C4299 vdd.n2454 gnd 0.006747f
C4300 vdd.n2455 gnd 0.006747f
C4301 vdd.n2456 gnd 0.006747f
C4302 vdd.n2457 gnd 0.006747f
C4303 vdd.n2458 gnd 0.006747f
C4304 vdd.n2459 gnd 0.006747f
C4305 vdd.n2460 gnd 0.006747f
C4306 vdd.n2461 gnd 0.006747f
C4307 vdd.n2462 gnd 0.006747f
C4308 vdd.n2463 gnd 0.006747f
C4309 vdd.n2464 gnd 0.006747f
C4310 vdd.n2465 gnd 0.006747f
C4311 vdd.n2466 gnd 0.006747f
C4312 vdd.n2467 gnd 0.006747f
C4313 vdd.n2468 gnd 0.006747f
C4314 vdd.n2469 gnd 0.006747f
C4315 vdd.n2470 gnd 0.006747f
C4316 vdd.n2471 gnd 0.006747f
C4317 vdd.n2472 gnd 0.218016f
C4318 vdd.n2473 gnd 0.006747f
C4319 vdd.n2474 gnd 0.006747f
C4320 vdd.n2475 gnd 0.006747f
C4321 vdd.n2476 gnd 0.006747f
C4322 vdd.n2477 gnd 0.006747f
C4323 vdd.n2478 gnd 0.006747f
C4324 vdd.n2479 gnd 0.006747f
C4325 vdd.n2480 gnd 0.006747f
C4326 vdd.n2481 gnd 0.006747f
C4327 vdd.n2482 gnd 0.006747f
C4328 vdd.n2483 gnd 0.006747f
C4329 vdd.n2484 gnd 0.006747f
C4330 vdd.n2485 gnd 0.006747f
C4331 vdd.n2486 gnd 0.006747f
C4332 vdd.n2487 gnd 0.006747f
C4333 vdd.n2488 gnd 0.006747f
C4334 vdd.n2489 gnd 0.006747f
C4335 vdd.n2490 gnd 0.006747f
C4336 vdd.n2491 gnd 0.006747f
C4337 vdd.n2492 gnd 0.006747f
C4338 vdd.n2493 gnd 0.410681f
C4339 vdd.n2494 gnd 0.006747f
C4340 vdd.n2495 gnd 0.006747f
C4341 vdd.n2496 gnd 0.006747f
C4342 vdd.n2497 gnd 0.006747f
C4343 vdd.n2498 gnd 0.006747f
C4344 vdd.n2499 gnd 0.014948f
C4345 vdd.n2500 gnd 0.01601f
C4346 vdd.n2501 gnd 0.01601f
C4347 vdd.n2502 gnd 0.006747f
C4348 vdd.n2503 gnd 0.006747f
C4349 vdd.n2504 gnd 0.006747f
C4350 vdd.n2505 gnd 0.005209f
C4351 vdd.n2506 gnd 0.009643f
C4352 vdd.n2507 gnd 0.004912f
C4353 vdd.n2508 gnd 0.006747f
C4354 vdd.n2509 gnd 0.006747f
C4355 vdd.n2510 gnd 0.006747f
C4356 vdd.n2511 gnd 0.006747f
C4357 vdd.n2512 gnd 0.006747f
C4358 vdd.n2513 gnd 0.006747f
C4359 vdd.n2514 gnd 0.006747f
C4360 vdd.n2515 gnd 0.006747f
C4361 vdd.n2516 gnd 0.006747f
C4362 vdd.n2517 gnd 0.006747f
C4363 vdd.n2518 gnd 0.006747f
C4364 vdd.n2519 gnd 0.006747f
C4365 vdd.n2520 gnd 0.006747f
C4366 vdd.n2521 gnd 0.006747f
C4367 vdd.n2522 gnd 0.006747f
C4368 vdd.n2523 gnd 0.006747f
C4369 vdd.n2524 gnd 0.006747f
C4370 vdd.n2525 gnd 0.006747f
C4371 vdd.n2526 gnd 0.006747f
C4372 vdd.n2527 gnd 0.006747f
C4373 vdd.n2528 gnd 0.006747f
C4374 vdd.n2529 gnd 0.006747f
C4375 vdd.n2530 gnd 0.006747f
C4376 vdd.n2531 gnd 0.006747f
C4377 vdd.n2532 gnd 0.006747f
C4378 vdd.n2533 gnd 0.006747f
C4379 vdd.n2534 gnd 0.006747f
C4380 vdd.n2535 gnd 0.006747f
C4381 vdd.n2536 gnd 0.006747f
C4382 vdd.n2537 gnd 0.006747f
C4383 vdd.n2538 gnd 0.006747f
C4384 vdd.n2539 gnd 0.006747f
C4385 vdd.n2540 gnd 0.006747f
C4386 vdd.n2541 gnd 0.006747f
C4387 vdd.n2542 gnd 0.006747f
C4388 vdd.n2543 gnd 0.006747f
C4389 vdd.n2544 gnd 0.006747f
C4390 vdd.n2545 gnd 0.006747f
C4391 vdd.n2546 gnd 0.006747f
C4392 vdd.n2547 gnd 0.006747f
C4393 vdd.n2548 gnd 0.006747f
C4394 vdd.n2549 gnd 0.006747f
C4395 vdd.n2550 gnd 0.006747f
C4396 vdd.n2551 gnd 0.006747f
C4397 vdd.n2552 gnd 0.006747f
C4398 vdd.n2553 gnd 0.006747f
C4399 vdd.n2554 gnd 0.006747f
C4400 vdd.n2555 gnd 0.006747f
C4401 vdd.n2556 gnd 0.006747f
C4402 vdd.n2557 gnd 0.006747f
C4403 vdd.n2558 gnd 0.006747f
C4404 vdd.n2559 gnd 0.006747f
C4405 vdd.n2560 gnd 0.006747f
C4406 vdd.n2561 gnd 0.006747f
C4407 vdd.n2562 gnd 0.006747f
C4408 vdd.n2563 gnd 0.006747f
C4409 vdd.n2564 gnd 0.006747f
C4410 vdd.n2565 gnd 0.006747f
C4411 vdd.n2566 gnd 0.006747f
C4412 vdd.n2567 gnd 0.006747f
C4413 vdd.n2569 gnd 0.841643f
C4414 vdd.n2571 gnd 0.006747f
C4415 vdd.n2572 gnd 0.006747f
C4416 vdd.n2573 gnd 0.01601f
C4417 vdd.n2574 gnd 0.014948f
C4418 vdd.n2575 gnd 0.014948f
C4419 vdd.n2576 gnd 0.841643f
C4420 vdd.n2577 gnd 0.014948f
C4421 vdd.n2578 gnd 0.014948f
C4422 vdd.n2579 gnd 0.006747f
C4423 vdd.n2580 gnd 0.006747f
C4424 vdd.n2581 gnd 0.006747f
C4425 vdd.n2582 gnd 0.430962f
C4426 vdd.n2583 gnd 0.006747f
C4427 vdd.n2584 gnd 0.006747f
C4428 vdd.n2585 gnd 0.006747f
C4429 vdd.n2586 gnd 0.006747f
C4430 vdd.n2587 gnd 0.006747f
C4431 vdd.n2588 gnd 0.537435f
C4432 vdd.n2589 gnd 0.006747f
C4433 vdd.n2590 gnd 0.006747f
C4434 vdd.n2591 gnd 0.006747f
C4435 vdd.n2592 gnd 0.006747f
C4436 vdd.n2593 gnd 0.006747f
C4437 vdd.n2594 gnd 0.689539f
C4438 vdd.n2595 gnd 0.006747f
C4439 vdd.n2596 gnd 0.006747f
C4440 vdd.n2597 gnd 0.006747f
C4441 vdd.n2598 gnd 0.006747f
C4442 vdd.n2599 gnd 0.006747f
C4443 vdd.n2600 gnd 0.38026f
C4444 vdd.n2601 gnd 0.006747f
C4445 vdd.n2602 gnd 0.006747f
C4446 vdd.n2603 gnd 0.006747f
C4447 vdd.n2604 gnd 0.006747f
C4448 vdd.n2605 gnd 0.006747f
C4449 vdd.n2606 gnd 0.218016f
C4450 vdd.n2607 gnd 0.006747f
C4451 vdd.n2608 gnd 0.006747f
C4452 vdd.n2609 gnd 0.006747f
C4453 vdd.n2610 gnd 0.006747f
C4454 vdd.n2611 gnd 0.006747f
C4455 vdd.n2612 gnd 0.395471f
C4456 vdd.n2613 gnd 0.006747f
C4457 vdd.n2614 gnd 0.006747f
C4458 vdd.n2615 gnd 0.006747f
C4459 vdd.n2616 gnd 0.006747f
C4460 vdd.n2617 gnd 0.006747f
C4461 vdd.n2618 gnd 0.547575f
C4462 vdd.n2619 gnd 0.006747f
C4463 vdd.n2620 gnd 0.006747f
C4464 vdd.n2621 gnd 0.006747f
C4465 vdd.n2622 gnd 0.006747f
C4466 vdd.n2623 gnd 0.006747f
C4467 vdd.n2624 gnd 0.613487f
C4468 vdd.n2625 gnd 0.006747f
C4469 vdd.n2626 gnd 0.006747f
C4470 vdd.n2627 gnd 0.006747f
C4471 vdd.n2628 gnd 0.006747f
C4472 vdd.n2629 gnd 0.006747f
C4473 vdd.n2630 gnd 0.461383f
C4474 vdd.n2631 gnd 0.006747f
C4475 vdd.n2632 gnd 0.006747f
C4476 vdd.n2633 gnd 0.006747f
C4477 vdd.t71 gnd 0.279098f
C4478 vdd.t69 gnd 0.178f
C4479 vdd.t72 gnd 0.279098f
C4480 vdd.n2634 gnd 0.156864f
C4481 vdd.n2635 gnd 0.019546f
C4482 vdd.n2636 gnd 0.004167f
C4483 vdd.n2637 gnd 0.006747f
C4484 vdd.n2638 gnd 0.38026f
C4485 vdd.n2639 gnd 0.006747f
C4486 vdd.n2640 gnd 0.006747f
C4487 vdd.n2641 gnd 0.006747f
C4488 vdd.n2642 gnd 0.006747f
C4489 vdd.n2643 gnd 0.006747f
C4490 vdd.n2644 gnd 0.689539f
C4491 vdd.n2645 gnd 0.006747f
C4492 vdd.n2646 gnd 0.006747f
C4493 vdd.n2647 gnd 0.006747f
C4494 vdd.n2648 gnd 0.006747f
C4495 vdd.n2649 gnd 0.006747f
C4496 vdd.n2650 gnd 0.006747f
C4497 vdd.n2652 gnd 0.006747f
C4498 vdd.n2653 gnd 0.006747f
C4499 vdd.n2655 gnd 0.006747f
C4500 vdd.n2656 gnd 0.006747f
C4501 vdd.n2659 gnd 0.006747f
C4502 vdd.n2660 gnd 0.006747f
C4503 vdd.n2661 gnd 0.006747f
C4504 vdd.n2662 gnd 0.006747f
C4505 vdd.n2664 gnd 0.006747f
C4506 vdd.n2665 gnd 0.006747f
C4507 vdd.n2666 gnd 0.006747f
C4508 vdd.n2667 gnd 0.006747f
C4509 vdd.n2668 gnd 0.006747f
C4510 vdd.n2669 gnd 0.006747f
C4511 vdd.n2671 gnd 0.006747f
C4512 vdd.n2672 gnd 0.006747f
C4513 vdd.n2673 gnd 0.006747f
C4514 vdd.n2674 gnd 0.006747f
C4515 vdd.n2675 gnd 0.006747f
C4516 vdd.n2676 gnd 0.006747f
C4517 vdd.n2678 gnd 0.006747f
C4518 vdd.n2679 gnd 0.006747f
C4519 vdd.n2680 gnd 0.006747f
C4520 vdd.n2681 gnd 0.006747f
C4521 vdd.n2682 gnd 0.006747f
C4522 vdd.n2683 gnd 0.006747f
C4523 vdd.n2685 gnd 0.006747f
C4524 vdd.n2686 gnd 0.01601f
C4525 vdd.n2687 gnd 0.01601f
C4526 vdd.n2688 gnd 0.014948f
C4527 vdd.n2689 gnd 0.006747f
C4528 vdd.n2690 gnd 0.006747f
C4529 vdd.n2691 gnd 0.006747f
C4530 vdd.n2692 gnd 0.006747f
C4531 vdd.n2693 gnd 0.006747f
C4532 vdd.n2694 gnd 0.006747f
C4533 vdd.n2695 gnd 0.689539f
C4534 vdd.n2696 gnd 0.006747f
C4535 vdd.n2697 gnd 0.006747f
C4536 vdd.n2698 gnd 0.006747f
C4537 vdd.n2699 gnd 0.006747f
C4538 vdd.n2700 gnd 0.006747f
C4539 vdd.n2701 gnd 0.430962f
C4540 vdd.n2702 gnd 0.006747f
C4541 vdd.n2703 gnd 0.006747f
C4542 vdd.n2704 gnd 0.006747f
C4543 vdd.n2705 gnd 0.01577f
C4544 vdd.n2707 gnd 0.01601f
C4545 vdd.n2708 gnd 0.015189f
C4546 vdd.n2709 gnd 0.006747f
C4547 vdd.n2710 gnd 0.005209f
C4548 vdd.n2711 gnd 0.006747f
C4549 vdd.n2713 gnd 0.006747f
C4550 vdd.n2714 gnd 0.006747f
C4551 vdd.n2715 gnd 0.006747f
C4552 vdd.n2716 gnd 0.006747f
C4553 vdd.n2717 gnd 0.006747f
C4554 vdd.n2718 gnd 0.006747f
C4555 vdd.n2720 gnd 0.006747f
C4556 vdd.n2721 gnd 0.006747f
C4557 vdd.n2722 gnd 0.006747f
C4558 vdd.n2723 gnd 0.006747f
C4559 vdd.n2724 gnd 0.006747f
C4560 vdd.n2725 gnd 0.006747f
C4561 vdd.n2727 gnd 0.006747f
C4562 vdd.n2728 gnd 0.006747f
C4563 vdd.n2729 gnd 0.006747f
C4564 vdd.n2730 gnd 0.006747f
C4565 vdd.n2731 gnd 0.006747f
C4566 vdd.n2732 gnd 0.006747f
C4567 vdd.n2734 gnd 0.006747f
C4568 vdd.n2735 gnd 0.006747f
C4569 vdd.n2736 gnd 0.006747f
C4570 vdd.n2737 gnd 0.600523f
C4571 vdd.n2738 gnd 0.016214f
C4572 vdd.n2739 gnd 0.006747f
C4573 vdd.n2740 gnd 0.006747f
C4574 vdd.n2742 gnd 0.006747f
C4575 vdd.n2743 gnd 0.006747f
C4576 vdd.n2744 gnd 0.006747f
C4577 vdd.n2745 gnd 0.006747f
C4578 vdd.n2746 gnd 0.006747f
C4579 vdd.n2747 gnd 0.006747f
C4580 vdd.n2749 gnd 0.006747f
C4581 vdd.n2750 gnd 0.006747f
C4582 vdd.n2751 gnd 0.006747f
C4583 vdd.n2752 gnd 0.006747f
C4584 vdd.n2753 gnd 0.006747f
C4585 vdd.n2754 gnd 0.006747f
C4586 vdd.n2756 gnd 0.006747f
C4587 vdd.n2757 gnd 0.006747f
C4588 vdd.n2758 gnd 0.006747f
C4589 vdd.n2759 gnd 0.006747f
C4590 vdd.n2760 gnd 0.006747f
C4591 vdd.n2761 gnd 0.006747f
C4592 vdd.n2763 gnd 0.006747f
C4593 vdd.n2764 gnd 0.006747f
C4594 vdd.n2766 gnd 0.006747f
C4595 vdd.n2767 gnd 0.006747f
C4596 vdd.n2768 gnd 0.01601f
C4597 vdd.n2769 gnd 0.014948f
C4598 vdd.n2770 gnd 0.014948f
C4599 vdd.n2771 gnd 0.993747f
C4600 vdd.n2772 gnd 0.014948f
C4601 vdd.n2773 gnd 0.01601f
C4602 vdd.n2774 gnd 0.015189f
C4603 vdd.n2775 gnd 0.006747f
C4604 vdd.n2776 gnd 0.005209f
C4605 vdd.n2777 gnd 0.006747f
C4606 vdd.n2779 gnd 0.006747f
C4607 vdd.n2780 gnd 0.006747f
C4608 vdd.n2781 gnd 0.006747f
C4609 vdd.n2782 gnd 0.006747f
C4610 vdd.n2783 gnd 0.006747f
C4611 vdd.n2784 gnd 0.006747f
C4612 vdd.n2786 gnd 0.006747f
C4613 vdd.n2787 gnd 0.006747f
C4614 vdd.n2788 gnd 0.006747f
C4615 vdd.n2789 gnd 0.006747f
C4616 vdd.n2790 gnd 0.006747f
C4617 vdd.n2791 gnd 0.006747f
C4618 vdd.n2793 gnd 0.006747f
C4619 vdd.n2794 gnd 0.006747f
C4620 vdd.n2795 gnd 0.006747f
C4621 vdd.n2796 gnd 0.006747f
C4622 vdd.n2797 gnd 0.006747f
C4623 vdd.n2798 gnd 0.006747f
C4624 vdd.n2800 gnd 0.006747f
C4625 vdd.n2801 gnd 0.006747f
C4626 vdd.n2803 gnd 0.006747f
C4627 vdd.n2804 gnd 0.016214f
C4628 vdd.n2805 gnd 0.600523f
C4629 vdd.n2806 gnd 0.008533f
C4630 vdd.n2807 gnd 0.003794f
C4631 vdd.t112 gnd 0.122072f
C4632 vdd.t113 gnd 0.130462f
C4633 vdd.t111 gnd 0.159425f
C4634 vdd.n2808 gnd 0.20436f
C4635 vdd.n2809 gnd 0.171699f
C4636 vdd.n2810 gnd 0.012299f
C4637 vdd.n2811 gnd 0.009922f
C4638 vdd.n2812 gnd 0.004193f
C4639 vdd.n2813 gnd 0.007986f
C4640 vdd.n2814 gnd 0.009922f
C4641 vdd.n2815 gnd 0.009922f
C4642 vdd.n2816 gnd 0.007986f
C4643 vdd.n2817 gnd 0.007986f
C4644 vdd.n2818 gnd 0.009922f
C4645 vdd.n2820 gnd 0.009922f
C4646 vdd.n2821 gnd 0.007986f
C4647 vdd.n2822 gnd 0.007986f
C4648 vdd.n2823 gnd 0.007986f
C4649 vdd.n2824 gnd 0.009922f
C4650 vdd.n2826 gnd 0.009922f
C4651 vdd.n2828 gnd 0.009922f
C4652 vdd.n2829 gnd 0.007986f
C4653 vdd.n2830 gnd 0.007986f
C4654 vdd.n2831 gnd 0.007986f
C4655 vdd.n2832 gnd 0.009922f
C4656 vdd.n2834 gnd 0.009922f
C4657 vdd.n2836 gnd 0.009922f
C4658 vdd.n2837 gnd 0.007986f
C4659 vdd.n2838 gnd 0.007986f
C4660 vdd.n2839 gnd 0.007986f
C4661 vdd.n2840 gnd 0.009922f
C4662 vdd.n2842 gnd 0.009922f
C4663 vdd.n2843 gnd 0.009922f
C4664 vdd.n2844 gnd 0.007986f
C4665 vdd.n2845 gnd 0.007986f
C4666 vdd.n2846 gnd 0.009922f
C4667 vdd.n2847 gnd 0.009922f
C4668 vdd.n2849 gnd 0.009922f
C4669 vdd.n2850 gnd 0.007986f
C4670 vdd.n2851 gnd 0.009922f
C4671 vdd.n2852 gnd 0.009922f
C4672 vdd.n2853 gnd 0.009922f
C4673 vdd.n2854 gnd 0.016292f
C4674 vdd.n2855 gnd 0.005431f
C4675 vdd.n2856 gnd 0.009922f
C4676 vdd.n2858 gnd 0.009922f
C4677 vdd.n2860 gnd 0.009922f
C4678 vdd.n2861 gnd 0.007986f
C4679 vdd.n2862 gnd 0.007986f
C4680 vdd.n2863 gnd 0.007986f
C4681 vdd.n2864 gnd 0.009922f
C4682 vdd.n2866 gnd 0.009922f
C4683 vdd.n2868 gnd 0.009922f
C4684 vdd.n2869 gnd 0.007986f
C4685 vdd.n2870 gnd 0.007986f
C4686 vdd.n2871 gnd 0.007986f
C4687 vdd.n2872 gnd 0.009922f
C4688 vdd.n2874 gnd 0.009922f
C4689 vdd.n2876 gnd 0.009922f
C4690 vdd.n2877 gnd 0.007986f
C4691 vdd.n2878 gnd 0.007986f
C4692 vdd.n2879 gnd 0.007986f
C4693 vdd.n2880 gnd 0.009922f
C4694 vdd.n2882 gnd 0.009922f
C4695 vdd.n2884 gnd 0.009922f
C4696 vdd.n2885 gnd 0.007986f
C4697 vdd.n2886 gnd 0.007986f
C4698 vdd.n2887 gnd 0.007986f
C4699 vdd.n2888 gnd 0.009922f
C4700 vdd.n2890 gnd 0.009922f
C4701 vdd.n2892 gnd 0.009922f
C4702 vdd.n2893 gnd 0.007986f
C4703 vdd.n2894 gnd 0.007986f
C4704 vdd.n2895 gnd 0.006669f
C4705 vdd.n2896 gnd 0.009922f
C4706 vdd.n2898 gnd 0.009922f
C4707 vdd.n2900 gnd 0.009922f
C4708 vdd.n2901 gnd 0.006669f
C4709 vdd.n2902 gnd 0.007986f
C4710 vdd.n2903 gnd 0.007986f
C4711 vdd.n2904 gnd 0.009922f
C4712 vdd.n2906 gnd 0.009922f
C4713 vdd.n2908 gnd 0.009922f
C4714 vdd.n2909 gnd 0.007986f
C4715 vdd.n2910 gnd 0.007986f
C4716 vdd.n2911 gnd 0.007986f
C4717 vdd.n2912 gnd 0.009922f
C4718 vdd.n2914 gnd 0.009922f
C4719 vdd.n2916 gnd 0.009922f
C4720 vdd.n2917 gnd 0.007986f
C4721 vdd.n2918 gnd 0.007986f
C4722 vdd.n2919 gnd 0.007986f
C4723 vdd.n2920 gnd 0.009922f
C4724 vdd.n2922 gnd 0.009922f
C4725 vdd.n2923 gnd 0.009922f
C4726 vdd.n2924 gnd 0.007986f
C4727 vdd.n2925 gnd 0.007986f
C4728 vdd.n2926 gnd 0.009922f
C4729 vdd.n2927 gnd 0.009922f
C4730 vdd.n2928 gnd 0.007986f
C4731 vdd.n2929 gnd 0.007986f
C4732 vdd.n2930 gnd 0.009922f
C4733 vdd.n2931 gnd 0.009922f
C4734 vdd.n2933 gnd 0.009922f
C4735 vdd.n2934 gnd 0.007986f
C4736 vdd.n2935 gnd 0.006629f
C4737 vdd.n2936 gnd 0.023749f
C4738 vdd.n2937 gnd 0.023383f
C4739 vdd.n2938 gnd 0.006629f
C4740 vdd.n2939 gnd 0.023383f
C4741 vdd.n2940 gnd 1.39429f
C4742 vdd.n2941 gnd 0.023383f
C4743 vdd.n2942 gnd 0.006629f
C4744 vdd.n2943 gnd 0.023383f
C4745 vdd.n2944 gnd 0.009922f
C4746 vdd.n2945 gnd 0.009922f
C4747 vdd.n2946 gnd 0.007986f
C4748 vdd.n2947 gnd 0.009922f
C4749 vdd.n2948 gnd 1.01403f
C4750 vdd.n2949 gnd 0.009922f
C4751 vdd.n2950 gnd 0.007986f
C4752 vdd.n2951 gnd 0.009922f
C4753 vdd.n2952 gnd 0.009922f
C4754 vdd.n2953 gnd 0.009922f
C4755 vdd.n2954 gnd 0.007986f
C4756 vdd.n2955 gnd 0.009922f
C4757 vdd.n2956 gnd 0.897415f
C4758 vdd.n2957 gnd 0.009922f
C4759 vdd.n2958 gnd 0.007986f
C4760 vdd.n2959 gnd 0.009922f
C4761 vdd.n2960 gnd 0.009922f
C4762 vdd.n2961 gnd 0.009922f
C4763 vdd.n2962 gnd 0.007986f
C4764 vdd.n2963 gnd 0.009922f
C4765 vdd.t19 gnd 0.507014f
C4766 vdd.n2964 gnd 0.72503f
C4767 vdd.n2965 gnd 0.009922f
C4768 vdd.n2966 gnd 0.007986f
C4769 vdd.n2967 gnd 0.009922f
C4770 vdd.n2968 gnd 0.009922f
C4771 vdd.n2969 gnd 0.009922f
C4772 vdd.n2970 gnd 0.007986f
C4773 vdd.n2971 gnd 0.009922f
C4774 vdd.n2972 gnd 0.552645f
C4775 vdd.n2973 gnd 0.009922f
C4776 vdd.n2974 gnd 0.007986f
C4777 vdd.n2975 gnd 0.009922f
C4778 vdd.n2976 gnd 0.009922f
C4779 vdd.n2977 gnd 0.009922f
C4780 vdd.n2978 gnd 0.007986f
C4781 vdd.n2979 gnd 0.009922f
C4782 vdd.n2980 gnd 0.71489f
C4783 vdd.n2981 gnd 0.633767f
C4784 vdd.n2982 gnd 0.009922f
C4785 vdd.n2983 gnd 0.007986f
C4786 vdd.n2984 gnd 0.009922f
C4787 vdd.n2985 gnd 0.009922f
C4788 vdd.n2986 gnd 0.009922f
C4789 vdd.n2987 gnd 0.007986f
C4790 vdd.n2988 gnd 0.009922f
C4791 vdd.n2989 gnd 0.806152f
C4792 vdd.n2990 gnd 0.009922f
C4793 vdd.n2991 gnd 0.007986f
C4794 vdd.n2992 gnd 0.009922f
C4795 vdd.n2993 gnd 0.009922f
C4796 vdd.n2994 gnd 0.009922f
C4797 vdd.n2995 gnd 0.007986f
C4798 vdd.n2996 gnd 0.007986f
C4799 vdd.n2997 gnd 0.007986f
C4800 vdd.n2998 gnd 0.009922f
C4801 vdd.n2999 gnd 0.009922f
C4802 vdd.n3000 gnd 0.009922f
C4803 vdd.n3001 gnd 0.007986f
C4804 vdd.n3002 gnd 0.007986f
C4805 vdd.n3003 gnd 0.007986f
C4806 vdd.n3004 gnd 0.009922f
C4807 vdd.n3005 gnd 0.009922f
C4808 vdd.n3006 gnd 0.009922f
C4809 vdd.n3007 gnd 0.007986f
C4810 vdd.n3008 gnd 0.007986f
C4811 vdd.n3009 gnd 0.007986f
C4812 vdd.n3010 gnd 0.009922f
C4813 vdd.n3011 gnd 0.009922f
C4814 vdd.n3012 gnd 0.009922f
C4815 vdd.n3013 gnd 0.007986f
C4816 vdd.n3014 gnd 0.007986f
C4817 vdd.n3015 gnd 0.006629f
C4818 vdd.n3016 gnd 0.023383f
C4819 vdd.n3017 gnd 0.023749f
C4820 vdd.n3019 gnd 0.023749f
C4821 vdd.n3020 gnd 0.003794f
C4822 vdd.t123 gnd 0.122072f
C4823 vdd.t122 gnd 0.130462f
C4824 vdd.t121 gnd 0.159425f
C4825 vdd.n3021 gnd 0.20436f
C4826 vdd.n3022 gnd 0.172498f
C4827 vdd.n3023 gnd 0.013098f
C4828 vdd.n3024 gnd 0.004193f
C4829 vdd.n3025 gnd 0.007986f
C4830 vdd.n3026 gnd 0.009922f
C4831 vdd.n3028 gnd 0.009922f
C4832 vdd.n3029 gnd 0.009922f
C4833 vdd.n3030 gnd 0.007986f
C4834 vdd.n3031 gnd 0.007986f
C4835 vdd.n3032 gnd 0.007986f
C4836 vdd.n3033 gnd 0.009922f
C4837 vdd.n3035 gnd 0.009922f
C4838 vdd.n3036 gnd 0.009922f
C4839 vdd.n3037 gnd 0.007986f
C4840 vdd.n3038 gnd 0.007986f
C4841 vdd.n3039 gnd 0.007986f
C4842 vdd.n3040 gnd 0.009922f
C4843 vdd.n3042 gnd 0.009922f
C4844 vdd.n3043 gnd 0.009922f
C4845 vdd.n3044 gnd 0.007986f
C4846 vdd.n3045 gnd 0.007986f
C4847 vdd.n3046 gnd 0.007986f
C4848 vdd.n3047 gnd 0.009922f
C4849 vdd.n3049 gnd 0.009922f
C4850 vdd.n3050 gnd 0.009922f
C4851 vdd.n3051 gnd 0.007986f
C4852 vdd.n3052 gnd 0.007986f
C4853 vdd.n3053 gnd 0.007986f
C4854 vdd.n3054 gnd 0.009922f
C4855 vdd.n3056 gnd 0.009922f
C4856 vdd.n3057 gnd 0.009922f
C4857 vdd.n3058 gnd 0.007986f
C4858 vdd.n3059 gnd 0.009922f
C4859 vdd.n3060 gnd 0.009922f
C4860 vdd.n3061 gnd 0.009922f
C4861 vdd.n3062 gnd 0.017091f
C4862 vdd.n3063 gnd 0.005431f
C4863 vdd.n3064 gnd 0.007986f
C4864 vdd.n3065 gnd 0.009922f
C4865 vdd.n3067 gnd 0.009922f
C4866 vdd.n3068 gnd 0.009922f
C4867 vdd.n3069 gnd 0.007986f
C4868 vdd.n3070 gnd 0.007986f
C4869 vdd.n3071 gnd 0.007986f
C4870 vdd.n3072 gnd 0.009922f
C4871 vdd.n3074 gnd 0.009922f
C4872 vdd.n3075 gnd 0.009922f
C4873 vdd.n3076 gnd 0.007986f
C4874 vdd.n3077 gnd 0.007986f
C4875 vdd.n3078 gnd 0.007986f
C4876 vdd.n3079 gnd 0.009922f
C4877 vdd.n3081 gnd 0.009922f
C4878 vdd.n3082 gnd 0.009922f
C4879 vdd.n3083 gnd 0.007986f
C4880 vdd.n3084 gnd 0.007986f
C4881 vdd.n3085 gnd 0.007986f
C4882 vdd.n3086 gnd 0.009922f
C4883 vdd.n3088 gnd 0.009922f
C4884 vdd.n3089 gnd 0.009922f
C4885 vdd.n3090 gnd 0.007986f
C4886 vdd.n3091 gnd 0.007986f
C4887 vdd.n3092 gnd 0.007986f
C4888 vdd.n3093 gnd 0.009922f
C4889 vdd.n3095 gnd 0.009922f
C4890 vdd.n3096 gnd 0.009922f
C4891 vdd.n3097 gnd 0.007986f
C4892 vdd.n3098 gnd 0.009922f
C4893 vdd.n3099 gnd 0.009922f
C4894 vdd.n3100 gnd 0.009922f
C4895 vdd.n3101 gnd 0.017091f
C4896 vdd.n3102 gnd 0.006669f
C4897 vdd.n3103 gnd 0.007986f
C4898 vdd.n3104 gnd 0.009922f
C4899 vdd.n3106 gnd 0.009922f
C4900 vdd.n3107 gnd 0.009922f
C4901 vdd.n3108 gnd 0.007986f
C4902 vdd.n3109 gnd 0.007986f
C4903 vdd.n3110 gnd 0.007986f
C4904 vdd.n3111 gnd 0.009922f
C4905 vdd.n3113 gnd 0.009922f
C4906 vdd.n3114 gnd 0.009922f
C4907 vdd.n3115 gnd 0.007986f
C4908 vdd.n3116 gnd 0.007986f
C4909 vdd.n3117 gnd 0.007986f
C4910 vdd.n3118 gnd 0.009922f
C4911 vdd.n3120 gnd 0.009922f
C4912 vdd.n3121 gnd 0.009922f
C4913 vdd.n3122 gnd 0.007986f
C4914 vdd.n3123 gnd 0.007986f
C4915 vdd.n3124 gnd 0.007986f
C4916 vdd.n3125 gnd 0.009922f
C4917 vdd.n3127 gnd 0.009922f
C4918 vdd.n3128 gnd 0.009922f
C4919 vdd.n3130 gnd 0.009922f
C4920 vdd.n3131 gnd 0.007986f
C4921 vdd.n3132 gnd 0.007986f
C4922 vdd.n3133 gnd 0.006629f
C4923 vdd.n3134 gnd 0.023749f
C4924 vdd.n3135 gnd 0.023383f
C4925 vdd.n3136 gnd 0.006629f
C4926 vdd.n3137 gnd 0.023383f
C4927 vdd.n3138 gnd 1.42978f
C4928 vdd.n3139 gnd 0.572926f
C4929 vdd.t115 gnd 0.507014f
C4930 vdd.n3140 gnd 0.948116f
C4931 vdd.n3141 gnd 0.009922f
C4932 vdd.n3142 gnd 0.007986f
C4933 vdd.n3143 gnd 0.007986f
C4934 vdd.n3144 gnd 0.007986f
C4935 vdd.n3145 gnd 0.009922f
C4936 vdd.n3146 gnd 0.998817f
C4937 vdd.t152 gnd 0.507014f
C4938 vdd.n3147 gnd 0.522224f
C4939 vdd.n3148 gnd 0.826433f
C4940 vdd.n3149 gnd 0.009922f
C4941 vdd.n3150 gnd 0.007986f
C4942 vdd.n3151 gnd 0.007986f
C4943 vdd.n3152 gnd 0.007986f
C4944 vdd.n3153 gnd 0.009922f
C4945 vdd.n3154 gnd 0.654048f
C4946 vdd.t149 gnd 0.507014f
C4947 vdd.n3155 gnd 0.841643f
C4948 vdd.t138 gnd 0.507014f
C4949 vdd.n3156 gnd 0.532365f
C4950 vdd.n3157 gnd 0.009922f
C4951 vdd.n3158 gnd 0.007986f
C4952 vdd.n3159 gnd 0.007986f
C4953 vdd.n3160 gnd 0.007986f
C4954 vdd.n3161 gnd 0.009922f
C4955 vdd.n3162 gnd 0.704749f
C4956 vdd.n3163 gnd 0.643908f
C4957 vdd.t187 gnd 0.507014f
C4958 vdd.n3164 gnd 0.841643f
C4959 vdd.n3165 gnd 0.009922f
C4960 vdd.n3166 gnd 0.007986f
C4961 vdd.n3167 gnd 0.590662f
C4962 vdd.n3168 gnd 2.18642f
C4963 commonsourceibias.n0 gnd 0.012299f
C4964 commonsourceibias.t56 gnd 0.18623f
C4965 commonsourceibias.t109 gnd 0.172196f
C4966 commonsourceibias.n1 gnd 0.068706f
C4967 commonsourceibias.n2 gnd 0.009217f
C4968 commonsourceibias.t69 gnd 0.172196f
C4969 commonsourceibias.n3 gnd 0.007456f
C4970 commonsourceibias.n4 gnd 0.009217f
C4971 commonsourceibias.t119 gnd 0.172196f
C4972 commonsourceibias.n5 gnd 0.008898f
C4973 commonsourceibias.n6 gnd 0.009217f
C4974 commonsourceibias.t85 gnd 0.172196f
C4975 commonsourceibias.n7 gnd 0.068706f
C4976 commonsourceibias.t54 gnd 0.172196f
C4977 commonsourceibias.n8 gnd 0.007444f
C4978 commonsourceibias.n9 gnd 0.012299f
C4979 commonsourceibias.t16 gnd 0.18623f
C4980 commonsourceibias.t30 gnd 0.172196f
C4981 commonsourceibias.n10 gnd 0.068706f
C4982 commonsourceibias.n11 gnd 0.009217f
C4983 commonsourceibias.t2 gnd 0.172196f
C4984 commonsourceibias.n12 gnd 0.007456f
C4985 commonsourceibias.n13 gnd 0.009217f
C4986 commonsourceibias.t22 gnd 0.172196f
C4987 commonsourceibias.n14 gnd 0.008898f
C4988 commonsourceibias.n15 gnd 0.009217f
C4989 commonsourceibias.t42 gnd 0.172196f
C4990 commonsourceibias.n16 gnd 0.068706f
C4991 commonsourceibias.t18 gnd 0.172196f
C4992 commonsourceibias.n17 gnd 0.007444f
C4993 commonsourceibias.n18 gnd 0.009217f
C4994 commonsourceibias.t32 gnd 0.172196f
C4995 commonsourceibias.t40 gnd 0.172196f
C4996 commonsourceibias.n19 gnd 0.068706f
C4997 commonsourceibias.n20 gnd 0.009217f
C4998 commonsourceibias.t24 gnd 0.172196f
C4999 commonsourceibias.n21 gnd 0.068706f
C5000 commonsourceibias.n22 gnd 0.009217f
C5001 commonsourceibias.t44 gnd 0.172196f
C5002 commonsourceibias.n23 gnd 0.068706f
C5003 commonsourceibias.n24 gnd 0.046399f
C5004 commonsourceibias.t6 gnd 0.172196f
C5005 commonsourceibias.t34 gnd 0.194303f
C5006 commonsourceibias.n25 gnd 0.079733f
C5007 commonsourceibias.n26 gnd 0.082545f
C5008 commonsourceibias.n27 gnd 0.01136f
C5009 commonsourceibias.n28 gnd 0.012567f
C5010 commonsourceibias.n29 gnd 0.009217f
C5011 commonsourceibias.n30 gnd 0.009217f
C5012 commonsourceibias.n31 gnd 0.012485f
C5013 commonsourceibias.n32 gnd 0.007456f
C5014 commonsourceibias.n33 gnd 0.01264f
C5015 commonsourceibias.n34 gnd 0.009217f
C5016 commonsourceibias.n35 gnd 0.009217f
C5017 commonsourceibias.n36 gnd 0.012717f
C5018 commonsourceibias.n37 gnd 0.010966f
C5019 commonsourceibias.n38 gnd 0.008898f
C5020 commonsourceibias.n39 gnd 0.009217f
C5021 commonsourceibias.n40 gnd 0.009217f
C5022 commonsourceibias.n41 gnd 0.011274f
C5023 commonsourceibias.n42 gnd 0.012653f
C5024 commonsourceibias.n43 gnd 0.068706f
C5025 commonsourceibias.n44 gnd 0.012568f
C5026 commonsourceibias.n45 gnd 0.009217f
C5027 commonsourceibias.n46 gnd 0.009217f
C5028 commonsourceibias.n47 gnd 0.009217f
C5029 commonsourceibias.n48 gnd 0.012568f
C5030 commonsourceibias.n49 gnd 0.068706f
C5031 commonsourceibias.n50 gnd 0.012653f
C5032 commonsourceibias.n51 gnd 0.011274f
C5033 commonsourceibias.n52 gnd 0.009217f
C5034 commonsourceibias.n53 gnd 0.009217f
C5035 commonsourceibias.n54 gnd 0.009217f
C5036 commonsourceibias.n55 gnd 0.010966f
C5037 commonsourceibias.n56 gnd 0.012717f
C5038 commonsourceibias.n57 gnd 0.068706f
C5039 commonsourceibias.n58 gnd 0.01264f
C5040 commonsourceibias.n59 gnd 0.009217f
C5041 commonsourceibias.n60 gnd 0.009217f
C5042 commonsourceibias.n61 gnd 0.009217f
C5043 commonsourceibias.n62 gnd 0.012485f
C5044 commonsourceibias.n63 gnd 0.068706f
C5045 commonsourceibias.n64 gnd 0.012567f
C5046 commonsourceibias.n65 gnd 0.01136f
C5047 commonsourceibias.n66 gnd 0.009217f
C5048 commonsourceibias.n67 gnd 0.009217f
C5049 commonsourceibias.n68 gnd 0.009349f
C5050 commonsourceibias.n69 gnd 0.009666f
C5051 commonsourceibias.n70 gnd 0.082208f
C5052 commonsourceibias.n71 gnd 0.091197f
C5053 commonsourceibias.t17 gnd 0.019889f
C5054 commonsourceibias.t31 gnd 0.019889f
C5055 commonsourceibias.n72 gnd 0.175743f
C5056 commonsourceibias.n73 gnd 0.151855f
C5057 commonsourceibias.t3 gnd 0.019889f
C5058 commonsourceibias.t23 gnd 0.019889f
C5059 commonsourceibias.n74 gnd 0.175743f
C5060 commonsourceibias.n75 gnd 0.080726f
C5061 commonsourceibias.t43 gnd 0.019889f
C5062 commonsourceibias.t19 gnd 0.019889f
C5063 commonsourceibias.n76 gnd 0.175743f
C5064 commonsourceibias.n77 gnd 0.067443f
C5065 commonsourceibias.t7 gnd 0.019889f
C5066 commonsourceibias.t35 gnd 0.019889f
C5067 commonsourceibias.n78 gnd 0.176331f
C5068 commonsourceibias.t25 gnd 0.019889f
C5069 commonsourceibias.t45 gnd 0.019889f
C5070 commonsourceibias.n79 gnd 0.175743f
C5071 commonsourceibias.n80 gnd 0.16376f
C5072 commonsourceibias.t33 gnd 0.019889f
C5073 commonsourceibias.t41 gnd 0.019889f
C5074 commonsourceibias.n81 gnd 0.175743f
C5075 commonsourceibias.n82 gnd 0.067443f
C5076 commonsourceibias.n83 gnd 0.081666f
C5077 commonsourceibias.n84 gnd 0.009217f
C5078 commonsourceibias.t100 gnd 0.172196f
C5079 commonsourceibias.t87 gnd 0.172196f
C5080 commonsourceibias.n85 gnd 0.068706f
C5081 commonsourceibias.n86 gnd 0.009217f
C5082 commonsourceibias.t115 gnd 0.172196f
C5083 commonsourceibias.n87 gnd 0.068706f
C5084 commonsourceibias.n88 gnd 0.009217f
C5085 commonsourceibias.t79 gnd 0.172196f
C5086 commonsourceibias.n89 gnd 0.068706f
C5087 commonsourceibias.n90 gnd 0.046399f
C5088 commonsourceibias.t66 gnd 0.172196f
C5089 commonsourceibias.t95 gnd 0.194303f
C5090 commonsourceibias.n91 gnd 0.079733f
C5091 commonsourceibias.n92 gnd 0.082545f
C5092 commonsourceibias.n93 gnd 0.01136f
C5093 commonsourceibias.n94 gnd 0.012567f
C5094 commonsourceibias.n95 gnd 0.009217f
C5095 commonsourceibias.n96 gnd 0.009217f
C5096 commonsourceibias.n97 gnd 0.012485f
C5097 commonsourceibias.n98 gnd 0.007456f
C5098 commonsourceibias.n99 gnd 0.01264f
C5099 commonsourceibias.n100 gnd 0.009217f
C5100 commonsourceibias.n101 gnd 0.009217f
C5101 commonsourceibias.n102 gnd 0.012717f
C5102 commonsourceibias.n103 gnd 0.010966f
C5103 commonsourceibias.n104 gnd 0.008898f
C5104 commonsourceibias.n105 gnd 0.009217f
C5105 commonsourceibias.n106 gnd 0.009217f
C5106 commonsourceibias.n107 gnd 0.011274f
C5107 commonsourceibias.n108 gnd 0.012653f
C5108 commonsourceibias.n109 gnd 0.068706f
C5109 commonsourceibias.n110 gnd 0.012568f
C5110 commonsourceibias.n111 gnd 0.009172f
C5111 commonsourceibias.n112 gnd 0.066626f
C5112 commonsourceibias.n113 gnd 0.009172f
C5113 commonsourceibias.n114 gnd 0.012568f
C5114 commonsourceibias.n115 gnd 0.068706f
C5115 commonsourceibias.n116 gnd 0.012653f
C5116 commonsourceibias.n117 gnd 0.011274f
C5117 commonsourceibias.n118 gnd 0.009217f
C5118 commonsourceibias.n119 gnd 0.009217f
C5119 commonsourceibias.n120 gnd 0.009217f
C5120 commonsourceibias.n121 gnd 0.010966f
C5121 commonsourceibias.n122 gnd 0.012717f
C5122 commonsourceibias.n123 gnd 0.068706f
C5123 commonsourceibias.n124 gnd 0.01264f
C5124 commonsourceibias.n125 gnd 0.009217f
C5125 commonsourceibias.n126 gnd 0.009217f
C5126 commonsourceibias.n127 gnd 0.009217f
C5127 commonsourceibias.n128 gnd 0.012485f
C5128 commonsourceibias.n129 gnd 0.068706f
C5129 commonsourceibias.n130 gnd 0.012567f
C5130 commonsourceibias.n131 gnd 0.01136f
C5131 commonsourceibias.n132 gnd 0.009217f
C5132 commonsourceibias.n133 gnd 0.009217f
C5133 commonsourceibias.n134 gnd 0.009349f
C5134 commonsourceibias.n135 gnd 0.009666f
C5135 commonsourceibias.n136 gnd 0.082208f
C5136 commonsourceibias.n137 gnd 0.05322f
C5137 commonsourceibias.n138 gnd 0.012299f
C5138 commonsourceibias.t89 gnd 0.18623f
C5139 commonsourceibias.t106 gnd 0.172196f
C5140 commonsourceibias.n139 gnd 0.068706f
C5141 commonsourceibias.n140 gnd 0.009217f
C5142 commonsourceibias.t101 gnd 0.172196f
C5143 commonsourceibias.n141 gnd 0.007456f
C5144 commonsourceibias.n142 gnd 0.009217f
C5145 commonsourceibias.t88 gnd 0.172196f
C5146 commonsourceibias.n143 gnd 0.008898f
C5147 commonsourceibias.n144 gnd 0.009217f
C5148 commonsourceibias.t105 gnd 0.172196f
C5149 commonsourceibias.n145 gnd 0.068706f
C5150 commonsourceibias.t99 gnd 0.172196f
C5151 commonsourceibias.n146 gnd 0.007444f
C5152 commonsourceibias.n147 gnd 0.009217f
C5153 commonsourceibias.t86 gnd 0.172196f
C5154 commonsourceibias.t108 gnd 0.172196f
C5155 commonsourceibias.n148 gnd 0.068706f
C5156 commonsourceibias.n149 gnd 0.009217f
C5157 commonsourceibias.t98 gnd 0.172196f
C5158 commonsourceibias.n150 gnd 0.068706f
C5159 commonsourceibias.n151 gnd 0.009217f
C5160 commonsourceibias.t112 gnd 0.172196f
C5161 commonsourceibias.n152 gnd 0.068706f
C5162 commonsourceibias.n153 gnd 0.046399f
C5163 commonsourceibias.t107 gnd 0.172196f
C5164 commonsourceibias.t97 gnd 0.194303f
C5165 commonsourceibias.n154 gnd 0.079733f
C5166 commonsourceibias.n155 gnd 0.082545f
C5167 commonsourceibias.n156 gnd 0.01136f
C5168 commonsourceibias.n157 gnd 0.012567f
C5169 commonsourceibias.n158 gnd 0.009217f
C5170 commonsourceibias.n159 gnd 0.009217f
C5171 commonsourceibias.n160 gnd 0.012485f
C5172 commonsourceibias.n161 gnd 0.007456f
C5173 commonsourceibias.n162 gnd 0.01264f
C5174 commonsourceibias.n163 gnd 0.009217f
C5175 commonsourceibias.n164 gnd 0.009217f
C5176 commonsourceibias.n165 gnd 0.012717f
C5177 commonsourceibias.n166 gnd 0.010966f
C5178 commonsourceibias.n167 gnd 0.008898f
C5179 commonsourceibias.n168 gnd 0.009217f
C5180 commonsourceibias.n169 gnd 0.009217f
C5181 commonsourceibias.n170 gnd 0.011274f
C5182 commonsourceibias.n171 gnd 0.012653f
C5183 commonsourceibias.n172 gnd 0.068706f
C5184 commonsourceibias.n173 gnd 0.012568f
C5185 commonsourceibias.n174 gnd 0.009217f
C5186 commonsourceibias.n175 gnd 0.009217f
C5187 commonsourceibias.n176 gnd 0.009217f
C5188 commonsourceibias.n177 gnd 0.012568f
C5189 commonsourceibias.n178 gnd 0.068706f
C5190 commonsourceibias.n179 gnd 0.012653f
C5191 commonsourceibias.n180 gnd 0.011274f
C5192 commonsourceibias.n181 gnd 0.009217f
C5193 commonsourceibias.n182 gnd 0.009217f
C5194 commonsourceibias.n183 gnd 0.009217f
C5195 commonsourceibias.n184 gnd 0.010966f
C5196 commonsourceibias.n185 gnd 0.012717f
C5197 commonsourceibias.n186 gnd 0.068706f
C5198 commonsourceibias.n187 gnd 0.01264f
C5199 commonsourceibias.n188 gnd 0.009217f
C5200 commonsourceibias.n189 gnd 0.009217f
C5201 commonsourceibias.n190 gnd 0.009217f
C5202 commonsourceibias.n191 gnd 0.012485f
C5203 commonsourceibias.n192 gnd 0.068706f
C5204 commonsourceibias.n193 gnd 0.012567f
C5205 commonsourceibias.n194 gnd 0.01136f
C5206 commonsourceibias.n195 gnd 0.009217f
C5207 commonsourceibias.n196 gnd 0.009217f
C5208 commonsourceibias.n197 gnd 0.009349f
C5209 commonsourceibias.n198 gnd 0.009666f
C5210 commonsourceibias.n199 gnd 0.082208f
C5211 commonsourceibias.n200 gnd 0.027976f
C5212 commonsourceibias.n201 gnd 0.147064f
C5213 commonsourceibias.n202 gnd 0.012299f
C5214 commonsourceibias.t50 gnd 0.172196f
C5215 commonsourceibias.n203 gnd 0.068706f
C5216 commonsourceibias.n204 gnd 0.009217f
C5217 commonsourceibias.t60 gnd 0.172196f
C5218 commonsourceibias.n205 gnd 0.007456f
C5219 commonsourceibias.n206 gnd 0.009217f
C5220 commonsourceibias.t104 gnd 0.172196f
C5221 commonsourceibias.n207 gnd 0.008898f
C5222 commonsourceibias.n208 gnd 0.009217f
C5223 commonsourceibias.t118 gnd 0.172196f
C5224 commonsourceibias.n209 gnd 0.068706f
C5225 commonsourceibias.t52 gnd 0.172196f
C5226 commonsourceibias.n210 gnd 0.007444f
C5227 commonsourceibias.n211 gnd 0.009217f
C5228 commonsourceibias.t93 gnd 0.172196f
C5229 commonsourceibias.t84 gnd 0.172196f
C5230 commonsourceibias.n212 gnd 0.068706f
C5231 commonsourceibias.n213 gnd 0.009217f
C5232 commonsourceibias.t49 gnd 0.172196f
C5233 commonsourceibias.n214 gnd 0.068706f
C5234 commonsourceibias.n215 gnd 0.009217f
C5235 commonsourceibias.t59 gnd 0.172196f
C5236 commonsourceibias.n216 gnd 0.068706f
C5237 commonsourceibias.n217 gnd 0.046399f
C5238 commonsourceibias.t75 gnd 0.172196f
C5239 commonsourceibias.t117 gnd 0.194303f
C5240 commonsourceibias.n218 gnd 0.079733f
C5241 commonsourceibias.n219 gnd 0.082545f
C5242 commonsourceibias.n220 gnd 0.01136f
C5243 commonsourceibias.n221 gnd 0.012567f
C5244 commonsourceibias.n222 gnd 0.009217f
C5245 commonsourceibias.n223 gnd 0.009217f
C5246 commonsourceibias.n224 gnd 0.012485f
C5247 commonsourceibias.n225 gnd 0.007456f
C5248 commonsourceibias.n226 gnd 0.01264f
C5249 commonsourceibias.n227 gnd 0.009217f
C5250 commonsourceibias.n228 gnd 0.009217f
C5251 commonsourceibias.n229 gnd 0.012717f
C5252 commonsourceibias.n230 gnd 0.010966f
C5253 commonsourceibias.n231 gnd 0.008898f
C5254 commonsourceibias.n232 gnd 0.009217f
C5255 commonsourceibias.n233 gnd 0.009217f
C5256 commonsourceibias.n234 gnd 0.011274f
C5257 commonsourceibias.n235 gnd 0.012653f
C5258 commonsourceibias.n236 gnd 0.068706f
C5259 commonsourceibias.n237 gnd 0.012568f
C5260 commonsourceibias.n238 gnd 0.009217f
C5261 commonsourceibias.n239 gnd 0.009217f
C5262 commonsourceibias.n240 gnd 0.009217f
C5263 commonsourceibias.n241 gnd 0.012568f
C5264 commonsourceibias.n242 gnd 0.068706f
C5265 commonsourceibias.n243 gnd 0.012653f
C5266 commonsourceibias.n244 gnd 0.011274f
C5267 commonsourceibias.n245 gnd 0.009217f
C5268 commonsourceibias.n246 gnd 0.009217f
C5269 commonsourceibias.n247 gnd 0.009217f
C5270 commonsourceibias.n248 gnd 0.010966f
C5271 commonsourceibias.n249 gnd 0.012717f
C5272 commonsourceibias.n250 gnd 0.068706f
C5273 commonsourceibias.n251 gnd 0.01264f
C5274 commonsourceibias.n252 gnd 0.009217f
C5275 commonsourceibias.n253 gnd 0.009217f
C5276 commonsourceibias.n254 gnd 0.009217f
C5277 commonsourceibias.n255 gnd 0.012485f
C5278 commonsourceibias.n256 gnd 0.068706f
C5279 commonsourceibias.n257 gnd 0.012567f
C5280 commonsourceibias.n258 gnd 0.01136f
C5281 commonsourceibias.n259 gnd 0.009217f
C5282 commonsourceibias.n260 gnd 0.009217f
C5283 commonsourceibias.n261 gnd 0.009349f
C5284 commonsourceibias.n262 gnd 0.009666f
C5285 commonsourceibias.t111 gnd 0.18623f
C5286 commonsourceibias.n263 gnd 0.082208f
C5287 commonsourceibias.n264 gnd 0.027976f
C5288 commonsourceibias.n265 gnd 0.517265f
C5289 commonsourceibias.n266 gnd 0.012299f
C5290 commonsourceibias.t114 gnd 0.18623f
C5291 commonsourceibias.t78 gnd 0.172196f
C5292 commonsourceibias.n267 gnd 0.068706f
C5293 commonsourceibias.n268 gnd 0.009217f
C5294 commonsourceibias.t53 gnd 0.172196f
C5295 commonsourceibias.n269 gnd 0.007456f
C5296 commonsourceibias.n270 gnd 0.009217f
C5297 commonsourceibias.t94 gnd 0.172196f
C5298 commonsourceibias.n271 gnd 0.008898f
C5299 commonsourceibias.n272 gnd 0.009217f
C5300 commonsourceibias.t113 gnd 0.172196f
C5301 commonsourceibias.n273 gnd 0.007444f
C5302 commonsourceibias.n274 gnd 0.009217f
C5303 commonsourceibias.t76 gnd 0.172196f
C5304 commonsourceibias.t65 gnd 0.172196f
C5305 commonsourceibias.n275 gnd 0.068706f
C5306 commonsourceibias.n276 gnd 0.009217f
C5307 commonsourceibias.t92 gnd 0.172196f
C5308 commonsourceibias.n277 gnd 0.068706f
C5309 commonsourceibias.n278 gnd 0.009217f
C5310 commonsourceibias.t63 gnd 0.172196f
C5311 commonsourceibias.n279 gnd 0.068706f
C5312 commonsourceibias.n280 gnd 0.046399f
C5313 commonsourceibias.t58 gnd 0.172196f
C5314 commonsourceibias.t70 gnd 0.194303f
C5315 commonsourceibias.n281 gnd 0.079733f
C5316 commonsourceibias.n282 gnd 0.082545f
C5317 commonsourceibias.n283 gnd 0.01136f
C5318 commonsourceibias.n284 gnd 0.012567f
C5319 commonsourceibias.n285 gnd 0.009217f
C5320 commonsourceibias.n286 gnd 0.009217f
C5321 commonsourceibias.n287 gnd 0.012485f
C5322 commonsourceibias.n288 gnd 0.007456f
C5323 commonsourceibias.n289 gnd 0.01264f
C5324 commonsourceibias.n290 gnd 0.009217f
C5325 commonsourceibias.n291 gnd 0.009217f
C5326 commonsourceibias.n292 gnd 0.012717f
C5327 commonsourceibias.n293 gnd 0.010966f
C5328 commonsourceibias.n294 gnd 0.008898f
C5329 commonsourceibias.n295 gnd 0.009217f
C5330 commonsourceibias.n296 gnd 0.009217f
C5331 commonsourceibias.n297 gnd 0.011274f
C5332 commonsourceibias.n298 gnd 0.012653f
C5333 commonsourceibias.n299 gnd 0.068706f
C5334 commonsourceibias.n300 gnd 0.012568f
C5335 commonsourceibias.n301 gnd 0.009172f
C5336 commonsourceibias.t5 gnd 0.019889f
C5337 commonsourceibias.t15 gnd 0.019889f
C5338 commonsourceibias.n302 gnd 0.176331f
C5339 commonsourceibias.t13 gnd 0.019889f
C5340 commonsourceibias.t39 gnd 0.019889f
C5341 commonsourceibias.n303 gnd 0.175743f
C5342 commonsourceibias.n304 gnd 0.16376f
C5343 commonsourceibias.t9 gnd 0.019889f
C5344 commonsourceibias.t1 gnd 0.019889f
C5345 commonsourceibias.n305 gnd 0.175743f
C5346 commonsourceibias.n306 gnd 0.067443f
C5347 commonsourceibias.n307 gnd 0.012299f
C5348 commonsourceibias.t46 gnd 0.172196f
C5349 commonsourceibias.n308 gnd 0.068706f
C5350 commonsourceibias.n309 gnd 0.009217f
C5351 commonsourceibias.t20 gnd 0.172196f
C5352 commonsourceibias.n310 gnd 0.007456f
C5353 commonsourceibias.n311 gnd 0.009217f
C5354 commonsourceibias.t36 gnd 0.172196f
C5355 commonsourceibias.n312 gnd 0.008898f
C5356 commonsourceibias.n313 gnd 0.009217f
C5357 commonsourceibias.t28 gnd 0.172196f
C5358 commonsourceibias.n314 gnd 0.007444f
C5359 commonsourceibias.n315 gnd 0.009217f
C5360 commonsourceibias.t0 gnd 0.172196f
C5361 commonsourceibias.t8 gnd 0.172196f
C5362 commonsourceibias.n316 gnd 0.068706f
C5363 commonsourceibias.n317 gnd 0.009217f
C5364 commonsourceibias.t38 gnd 0.172196f
C5365 commonsourceibias.n318 gnd 0.068706f
C5366 commonsourceibias.n319 gnd 0.009217f
C5367 commonsourceibias.t12 gnd 0.172196f
C5368 commonsourceibias.n320 gnd 0.068706f
C5369 commonsourceibias.n321 gnd 0.046399f
C5370 commonsourceibias.t14 gnd 0.172196f
C5371 commonsourceibias.t4 gnd 0.194303f
C5372 commonsourceibias.n322 gnd 0.079733f
C5373 commonsourceibias.n323 gnd 0.082545f
C5374 commonsourceibias.n324 gnd 0.01136f
C5375 commonsourceibias.n325 gnd 0.012567f
C5376 commonsourceibias.n326 gnd 0.009217f
C5377 commonsourceibias.n327 gnd 0.009217f
C5378 commonsourceibias.n328 gnd 0.012485f
C5379 commonsourceibias.n329 gnd 0.007456f
C5380 commonsourceibias.n330 gnd 0.01264f
C5381 commonsourceibias.n331 gnd 0.009217f
C5382 commonsourceibias.n332 gnd 0.009217f
C5383 commonsourceibias.n333 gnd 0.012717f
C5384 commonsourceibias.n334 gnd 0.010966f
C5385 commonsourceibias.n335 gnd 0.008898f
C5386 commonsourceibias.n336 gnd 0.009217f
C5387 commonsourceibias.n337 gnd 0.009217f
C5388 commonsourceibias.n338 gnd 0.011274f
C5389 commonsourceibias.n339 gnd 0.012653f
C5390 commonsourceibias.n340 gnd 0.068706f
C5391 commonsourceibias.n341 gnd 0.012568f
C5392 commonsourceibias.n342 gnd 0.009217f
C5393 commonsourceibias.n343 gnd 0.009217f
C5394 commonsourceibias.n344 gnd 0.009217f
C5395 commonsourceibias.n345 gnd 0.012568f
C5396 commonsourceibias.n346 gnd 0.068706f
C5397 commonsourceibias.n347 gnd 0.012653f
C5398 commonsourceibias.t10 gnd 0.172196f
C5399 commonsourceibias.n348 gnd 0.068706f
C5400 commonsourceibias.n349 gnd 0.011274f
C5401 commonsourceibias.n350 gnd 0.009217f
C5402 commonsourceibias.n351 gnd 0.009217f
C5403 commonsourceibias.n352 gnd 0.009217f
C5404 commonsourceibias.n353 gnd 0.010966f
C5405 commonsourceibias.n354 gnd 0.012717f
C5406 commonsourceibias.n355 gnd 0.068706f
C5407 commonsourceibias.n356 gnd 0.01264f
C5408 commonsourceibias.n357 gnd 0.009217f
C5409 commonsourceibias.n358 gnd 0.009217f
C5410 commonsourceibias.n359 gnd 0.009217f
C5411 commonsourceibias.n360 gnd 0.012485f
C5412 commonsourceibias.n361 gnd 0.068706f
C5413 commonsourceibias.n362 gnd 0.012567f
C5414 commonsourceibias.n363 gnd 0.01136f
C5415 commonsourceibias.n364 gnd 0.009217f
C5416 commonsourceibias.n365 gnd 0.009217f
C5417 commonsourceibias.n366 gnd 0.009349f
C5418 commonsourceibias.n367 gnd 0.009666f
C5419 commonsourceibias.t26 gnd 0.18623f
C5420 commonsourceibias.n368 gnd 0.082208f
C5421 commonsourceibias.n369 gnd 0.091197f
C5422 commonsourceibias.t47 gnd 0.019889f
C5423 commonsourceibias.t27 gnd 0.019889f
C5424 commonsourceibias.n370 gnd 0.175743f
C5425 commonsourceibias.n371 gnd 0.151855f
C5426 commonsourceibias.t37 gnd 0.019889f
C5427 commonsourceibias.t21 gnd 0.019889f
C5428 commonsourceibias.n372 gnd 0.175743f
C5429 commonsourceibias.n373 gnd 0.080726f
C5430 commonsourceibias.t29 gnd 0.019889f
C5431 commonsourceibias.t11 gnd 0.019889f
C5432 commonsourceibias.n374 gnd 0.175743f
C5433 commonsourceibias.n375 gnd 0.067443f
C5434 commonsourceibias.n376 gnd 0.081666f
C5435 commonsourceibias.n377 gnd 0.066626f
C5436 commonsourceibias.n378 gnd 0.009172f
C5437 commonsourceibias.n379 gnd 0.012568f
C5438 commonsourceibias.n380 gnd 0.068706f
C5439 commonsourceibias.n381 gnd 0.012653f
C5440 commonsourceibias.t64 gnd 0.172196f
C5441 commonsourceibias.n382 gnd 0.068706f
C5442 commonsourceibias.n383 gnd 0.011274f
C5443 commonsourceibias.n384 gnd 0.009217f
C5444 commonsourceibias.n385 gnd 0.009217f
C5445 commonsourceibias.n386 gnd 0.009217f
C5446 commonsourceibias.n387 gnd 0.010966f
C5447 commonsourceibias.n388 gnd 0.012717f
C5448 commonsourceibias.n389 gnd 0.068706f
C5449 commonsourceibias.n390 gnd 0.01264f
C5450 commonsourceibias.n391 gnd 0.009217f
C5451 commonsourceibias.n392 gnd 0.009217f
C5452 commonsourceibias.n393 gnd 0.009217f
C5453 commonsourceibias.n394 gnd 0.012485f
C5454 commonsourceibias.n395 gnd 0.068706f
C5455 commonsourceibias.n396 gnd 0.012567f
C5456 commonsourceibias.n397 gnd 0.01136f
C5457 commonsourceibias.n398 gnd 0.009217f
C5458 commonsourceibias.n399 gnd 0.009217f
C5459 commonsourceibias.n400 gnd 0.009349f
C5460 commonsourceibias.n401 gnd 0.009666f
C5461 commonsourceibias.n402 gnd 0.082208f
C5462 commonsourceibias.n403 gnd 0.05322f
C5463 commonsourceibias.n404 gnd 0.012299f
C5464 commonsourceibias.t91 gnd 0.172196f
C5465 commonsourceibias.n405 gnd 0.068706f
C5466 commonsourceibias.n406 gnd 0.009217f
C5467 commonsourceibias.t83 gnd 0.172196f
C5468 commonsourceibias.n407 gnd 0.007456f
C5469 commonsourceibias.n408 gnd 0.009217f
C5470 commonsourceibias.t73 gnd 0.172196f
C5471 commonsourceibias.n409 gnd 0.008898f
C5472 commonsourceibias.n410 gnd 0.009217f
C5473 commonsourceibias.t82 gnd 0.172196f
C5474 commonsourceibias.n411 gnd 0.007444f
C5475 commonsourceibias.n412 gnd 0.009217f
C5476 commonsourceibias.t103 gnd 0.172196f
C5477 commonsourceibias.t96 gnd 0.172196f
C5478 commonsourceibias.n413 gnd 0.068706f
C5479 commonsourceibias.n414 gnd 0.009217f
C5480 commonsourceibias.t81 gnd 0.172196f
C5481 commonsourceibias.n415 gnd 0.068706f
C5482 commonsourceibias.n416 gnd 0.009217f
C5483 commonsourceibias.t102 gnd 0.172196f
C5484 commonsourceibias.n417 gnd 0.068706f
C5485 commonsourceibias.n418 gnd 0.046399f
C5486 commonsourceibias.t116 gnd 0.172196f
C5487 commonsourceibias.t80 gnd 0.194303f
C5488 commonsourceibias.n419 gnd 0.079733f
C5489 commonsourceibias.n420 gnd 0.082545f
C5490 commonsourceibias.n421 gnd 0.01136f
C5491 commonsourceibias.n422 gnd 0.012567f
C5492 commonsourceibias.n423 gnd 0.009217f
C5493 commonsourceibias.n424 gnd 0.009217f
C5494 commonsourceibias.n425 gnd 0.012485f
C5495 commonsourceibias.n426 gnd 0.007456f
C5496 commonsourceibias.n427 gnd 0.01264f
C5497 commonsourceibias.n428 gnd 0.009217f
C5498 commonsourceibias.n429 gnd 0.009217f
C5499 commonsourceibias.n430 gnd 0.012717f
C5500 commonsourceibias.n431 gnd 0.010966f
C5501 commonsourceibias.n432 gnd 0.008898f
C5502 commonsourceibias.n433 gnd 0.009217f
C5503 commonsourceibias.n434 gnd 0.009217f
C5504 commonsourceibias.n435 gnd 0.011274f
C5505 commonsourceibias.n436 gnd 0.012653f
C5506 commonsourceibias.n437 gnd 0.068706f
C5507 commonsourceibias.n438 gnd 0.012568f
C5508 commonsourceibias.n439 gnd 0.009217f
C5509 commonsourceibias.n440 gnd 0.009217f
C5510 commonsourceibias.n441 gnd 0.009217f
C5511 commonsourceibias.n442 gnd 0.012568f
C5512 commonsourceibias.n443 gnd 0.068706f
C5513 commonsourceibias.n444 gnd 0.012653f
C5514 commonsourceibias.t90 gnd 0.172196f
C5515 commonsourceibias.n445 gnd 0.068706f
C5516 commonsourceibias.n446 gnd 0.011274f
C5517 commonsourceibias.n447 gnd 0.009217f
C5518 commonsourceibias.n448 gnd 0.009217f
C5519 commonsourceibias.n449 gnd 0.009217f
C5520 commonsourceibias.n450 gnd 0.010966f
C5521 commonsourceibias.n451 gnd 0.012717f
C5522 commonsourceibias.n452 gnd 0.068706f
C5523 commonsourceibias.n453 gnd 0.01264f
C5524 commonsourceibias.n454 gnd 0.009217f
C5525 commonsourceibias.n455 gnd 0.009217f
C5526 commonsourceibias.n456 gnd 0.009217f
C5527 commonsourceibias.n457 gnd 0.012485f
C5528 commonsourceibias.n458 gnd 0.068706f
C5529 commonsourceibias.n459 gnd 0.012567f
C5530 commonsourceibias.n460 gnd 0.01136f
C5531 commonsourceibias.n461 gnd 0.009217f
C5532 commonsourceibias.n462 gnd 0.009217f
C5533 commonsourceibias.n463 gnd 0.009349f
C5534 commonsourceibias.n464 gnd 0.009666f
C5535 commonsourceibias.t74 gnd 0.18623f
C5536 commonsourceibias.n465 gnd 0.082208f
C5537 commonsourceibias.n466 gnd 0.027976f
C5538 commonsourceibias.n467 gnd 0.147064f
C5539 commonsourceibias.n468 gnd 0.012299f
C5540 commonsourceibias.t62 gnd 0.172196f
C5541 commonsourceibias.n469 gnd 0.068706f
C5542 commonsourceibias.n470 gnd 0.009217f
C5543 commonsourceibias.t71 gnd 0.172196f
C5544 commonsourceibias.n471 gnd 0.007456f
C5545 commonsourceibias.n472 gnd 0.009217f
C5546 commonsourceibias.t48 gnd 0.172196f
C5547 commonsourceibias.n473 gnd 0.008898f
C5548 commonsourceibias.n474 gnd 0.009217f
C5549 commonsourceibias.t67 gnd 0.172196f
C5550 commonsourceibias.n475 gnd 0.007444f
C5551 commonsourceibias.n476 gnd 0.009217f
C5552 commonsourceibias.t77 gnd 0.172196f
C5553 commonsourceibias.t110 gnd 0.172196f
C5554 commonsourceibias.n477 gnd 0.068706f
C5555 commonsourceibias.n478 gnd 0.009217f
C5556 commonsourceibias.t61 gnd 0.172196f
C5557 commonsourceibias.n479 gnd 0.068706f
C5558 commonsourceibias.n480 gnd 0.009217f
C5559 commonsourceibias.t72 gnd 0.172196f
C5560 commonsourceibias.n481 gnd 0.068706f
C5561 commonsourceibias.n482 gnd 0.046399f
C5562 commonsourceibias.t68 gnd 0.172196f
C5563 commonsourceibias.t55 gnd 0.194303f
C5564 commonsourceibias.n483 gnd 0.079733f
C5565 commonsourceibias.n484 gnd 0.082545f
C5566 commonsourceibias.n485 gnd 0.01136f
C5567 commonsourceibias.n486 gnd 0.012567f
C5568 commonsourceibias.n487 gnd 0.009217f
C5569 commonsourceibias.n488 gnd 0.009217f
C5570 commonsourceibias.n489 gnd 0.012485f
C5571 commonsourceibias.n490 gnd 0.007456f
C5572 commonsourceibias.n491 gnd 0.01264f
C5573 commonsourceibias.n492 gnd 0.009217f
C5574 commonsourceibias.n493 gnd 0.009217f
C5575 commonsourceibias.n494 gnd 0.012717f
C5576 commonsourceibias.n495 gnd 0.010966f
C5577 commonsourceibias.n496 gnd 0.008898f
C5578 commonsourceibias.n497 gnd 0.009217f
C5579 commonsourceibias.n498 gnd 0.009217f
C5580 commonsourceibias.n499 gnd 0.011274f
C5581 commonsourceibias.n500 gnd 0.012653f
C5582 commonsourceibias.n501 gnd 0.068706f
C5583 commonsourceibias.n502 gnd 0.012568f
C5584 commonsourceibias.n503 gnd 0.009217f
C5585 commonsourceibias.n504 gnd 0.009217f
C5586 commonsourceibias.n505 gnd 0.009217f
C5587 commonsourceibias.n506 gnd 0.012568f
C5588 commonsourceibias.n507 gnd 0.068706f
C5589 commonsourceibias.n508 gnd 0.012653f
C5590 commonsourceibias.t57 gnd 0.172196f
C5591 commonsourceibias.n509 gnd 0.068706f
C5592 commonsourceibias.n510 gnd 0.011274f
C5593 commonsourceibias.n511 gnd 0.009217f
C5594 commonsourceibias.n512 gnd 0.009217f
C5595 commonsourceibias.n513 gnd 0.009217f
C5596 commonsourceibias.n514 gnd 0.010966f
C5597 commonsourceibias.n515 gnd 0.012717f
C5598 commonsourceibias.n516 gnd 0.068706f
C5599 commonsourceibias.n517 gnd 0.01264f
C5600 commonsourceibias.n518 gnd 0.009217f
C5601 commonsourceibias.n519 gnd 0.009217f
C5602 commonsourceibias.n520 gnd 0.009217f
C5603 commonsourceibias.n521 gnd 0.012485f
C5604 commonsourceibias.n522 gnd 0.068706f
C5605 commonsourceibias.n523 gnd 0.012567f
C5606 commonsourceibias.n524 gnd 0.01136f
C5607 commonsourceibias.n525 gnd 0.009217f
C5608 commonsourceibias.n526 gnd 0.009217f
C5609 commonsourceibias.n527 gnd 0.009349f
C5610 commonsourceibias.n528 gnd 0.009666f
C5611 commonsourceibias.t51 gnd 0.18623f
C5612 commonsourceibias.n529 gnd 0.082208f
C5613 commonsourceibias.n530 gnd 0.027976f
C5614 commonsourceibias.n531 gnd 0.194274f
C5615 commonsourceibias.n532 gnd 5.09694f
.ends

