* NGSPICE file created from opamp125.ext - technology: sky130A

.subckt opamp125 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 gnd.t406 commonsourceibias.t4 commonsourceibias.t5 gnd.t309 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X1 a_n7636_8799.t29 plus.t5 a_n3827_n3924.t8 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X2 a_n2804_13878.t26 a_n2982_13878.t26 a_n2982_13878.t27 vdd.t49 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 a_n2804_13878.t1 a_n2982_13878.t72 vdd.t60 vdd.t59 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 gnd.t206 gnd.t204 gnd.t205 gnd.t157 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X5 gnd.t405 commonsourceibias.t80 CSoutput.t119 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X6 gnd.t404 commonsourceibias.t81 CSoutput.t118 gnd.t263 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 CSoutput.t117 commonsourceibias.t82 gnd.t402 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 vdd.t211 a_n7636_8799.t48 CSoutput.t167 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X9 commonsourceibias.t3 commonsourceibias.t2 gnd.t403 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X10 gnd.t401 commonsourceibias.t83 CSoutput.t116 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X11 gnd.t203 gnd.t201 minus.t4 gnd.t202 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X12 gnd.t400 commonsourceibias.t0 commonsourceibias.t1 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X13 a_n3827_n3924.t45 diffpairibias.t20 gnd.t64 gnd.t63 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X14 CSoutput.t115 commonsourceibias.t84 gnd.t399 gnd.t347 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X15 a_n3827_n3924.t14 plus.t6 a_n7636_8799.t28 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X16 gnd.t398 commonsourceibias.t48 commonsourceibias.t49 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X17 vdd.t142 vdd.t140 vdd.t141 vdd.t101 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X18 a_n3827_n3924.t2 minus.t5 a_n2982_13878.t2 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X19 a_n2982_8322.t31 a_n2982_13878.t73 a_n7636_8799.t4 vdd.t57 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X20 commonsourceibias.t47 commonsourceibias.t46 gnd.t397 gnd.t259 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X21 gnd.t396 commonsourceibias.t85 CSoutput.t114 gnd.t301 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X22 CSoutput.t166 a_n7636_8799.t49 vdd.t210 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X23 vdd.t209 a_n7636_8799.t50 CSoutput.t165 vdd.t182 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X24 a_n2982_13878.t71 minus.t6 a_n3827_n3924.t56 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X25 gnd.t200 gnd.t198 gnd.t199 gnd.t124 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X26 a_n7636_8799.t45 a_n2982_13878.t74 a_n2982_8322.t30 vdd.t45 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X27 CSoutput.t113 commonsourceibias.t86 gnd.t395 gnd.t278 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X28 gnd.t197 gnd.t194 gnd.t196 gnd.t195 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X29 CSoutput.t112 commonsourceibias.t87 gnd.t394 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X30 a_n2982_13878.t67 minus.t7 a_n3827_n3924.t47 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X31 vdd.t208 a_n7636_8799.t51 CSoutput.t164 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X32 commonsourceibias.t45 commonsourceibias.t44 gnd.t393 gnd.t307 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X33 a_n7636_8799.t3 a_n2982_13878.t75 a_n2982_8322.t29 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X34 gnd.t392 commonsourceibias.t88 CSoutput.t111 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 gnd.t193 gnd.t191 gnd.t192 gnd.t113 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X36 CSoutput.t110 commonsourceibias.t89 gnd.t391 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X37 a_n3827_n3924.t3 minus.t8 a_n2982_13878.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X38 CSoutput.t109 commonsourceibias.t90 gnd.t390 gnd.t347 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X39 gnd.t389 commonsourceibias.t42 commonsourceibias.t43 gnd.t301 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X40 outputibias.t7 outputibias.t6 gnd.t408 gnd.t407 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X41 gnd.t388 commonsourceibias.t40 commonsourceibias.t41 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X42 CSoutput.t108 commonsourceibias.t91 gnd.t373 gnd.t311 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X43 a_n3827_n3924.t48 diffpairibias.t21 gnd.t72 gnd.t71 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X44 commonsourceibias.t39 commonsourceibias.t38 gnd.t387 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X45 CSoutput.t107 commonsourceibias.t92 gnd.t386 gnd.t311 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X46 a_n3827_n3924.t16 plus.t7 a_n7636_8799.t27 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X47 gnd.t385 commonsourceibias.t36 commonsourceibias.t37 gnd.t294 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X48 CSoutput.t106 commonsourceibias.t93 gnd.t384 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X49 a_n2804_13878.t25 a_n2982_13878.t20 a_n2982_13878.t21 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X50 vdd.t139 vdd.t137 vdd.t138 vdd.t101 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X51 a_n7636_8799.t26 plus.t8 a_n3827_n3924.t11 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X52 a_n2982_13878.t23 a_n2982_13878.t22 a_n2804_13878.t24 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X53 a_n7636_8799.t25 plus.t9 a_n3827_n3924.t23 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X54 CSoutput.t163 a_n7636_8799.t52 vdd.t207 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X55 vdd.t136 vdd.t134 vdd.t135 vdd.t117 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X56 vdd.t206 a_n7636_8799.t53 CSoutput.t162 vdd.t182 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X57 CSoutput.t105 commonsourceibias.t94 gnd.t383 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X58 vdd.t61 CSoutput.t168 output.t19 gnd.t30 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X59 gnd.t382 commonsourceibias.t95 CSoutput.t104 gnd.t263 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X60 diffpairibias.t19 diffpairibias.t18 gnd.t7 gnd.t6 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X61 CSoutput.t103 commonsourceibias.t96 gnd.t379 gnd.t269 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X62 a_n3827_n3924.t20 plus.t10 a_n7636_8799.t24 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X63 a_n2982_13878.t65 minus.t9 a_n3827_n3924.t44 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X64 a_n2982_13878.t31 a_n2982_13878.t30 a_n2804_13878.t23 vdd.t44 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X65 a_n7636_8799.t2 a_n2982_13878.t76 a_n2982_8322.t28 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X66 CSoutput.t102 commonsourceibias.t97 gnd.t381 gnd.t322 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X67 CSoutput.t101 commonsourceibias.t98 gnd.t380 gnd.t291 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X68 CSoutput.t161 a_n7636_8799.t54 vdd.t205 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X69 commonsourceibias.t57 commonsourceibias.t56 gnd.t378 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X70 gnd.t190 gnd.t188 plus.t4 gnd.t189 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X71 a_n2982_13878.t11 a_n2982_13878.t10 a_n2804_13878.t22 vdd.t58 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X72 gnd.t187 gnd.t185 gnd.t186 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X73 vdd.t204 a_n7636_8799.t55 CSoutput.t160 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X74 vdd.t203 a_n7636_8799.t56 CSoutput.t159 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X75 CSoutput.t100 commonsourceibias.t99 gnd.t377 gnd.t347 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X76 a_n7636_8799.t36 a_n2982_13878.t77 a_n2982_8322.t27 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X77 diffpairibias.t17 diffpairibias.t16 gnd.t24 gnd.t23 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X78 CSoutput.t158 a_n7636_8799.t57 vdd.t202 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X79 gnd.t184 gnd.t182 gnd.t183 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X80 a_n7636_8799.t40 a_n2982_13878.t78 a_n2982_8322.t26 vdd.t52 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X81 a_n2982_8322.t25 a_n2982_13878.t79 a_n7636_8799.t42 vdd.t58 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X82 CSoutput.t99 commonsourceibias.t100 gnd.t375 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X83 CSoutput.t98 commonsourceibias.t101 gnd.t376 gnd.t291 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X84 gnd.t181 gnd.t179 gnd.t180 gnd.t131 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X85 CSoutput.t157 a_n7636_8799.t58 vdd.t201 vdd.t177 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X86 gnd.t374 commonsourceibias.t102 CSoutput.t97 gnd.t265 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X87 gnd.t178 gnd.t176 gnd.t177 gnd.t106 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X88 gnd.t175 gnd.t173 plus.t3 gnd.t174 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X89 CSoutput.t96 commonsourceibias.t103 gnd.t372 gnd.t287 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 gnd.t371 commonsourceibias.t104 CSoutput.t95 gnd.t244 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X91 a_n3827_n3924.t17 plus.t11 a_n7636_8799.t23 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X92 gnd.t172 gnd.t170 gnd.t171 gnd.t124 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X93 output.t3 outputibias.t8 gnd.t80 gnd.t79 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X94 a_n3827_n3924.t42 diffpairibias.t22 gnd.t58 gnd.t57 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X95 vdd.t200 a_n7636_8799.t59 CSoutput.t156 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X96 CSoutput.t94 commonsourceibias.t105 gnd.t370 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X97 a_n2982_13878.t13 a_n2982_13878.t12 a_n2804_13878.t21 vdd.t57 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X98 a_n7636_8799.t35 a_n2982_13878.t80 a_n2982_8322.t24 vdd.t48 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X99 a_n2982_13878.t9 a_n2982_13878.t8 a_n2804_13878.t20 vdd.t9 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X100 gnd.t369 commonsourceibias.t106 CSoutput.t93 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X101 vdd.t62 CSoutput.t169 output.t18 gnd.t31 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X102 commonsourceibias.t55 commonsourceibias.t54 gnd.t368 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X103 gnd.t367 commonsourceibias.t107 CSoutput.t92 gnd.t261 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X104 gnd.t169 gnd.t166 gnd.t168 gnd.t167 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X105 CSoutput.t91 commonsourceibias.t108 gnd.t366 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X106 CSoutput.t170 a_n2982_8322.t37 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X107 gnd.t365 commonsourceibias.t52 commonsourceibias.t53 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 CSoutput.t90 commonsourceibias.t109 gnd.t364 gnd.t311 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X109 diffpairibias.t15 diffpairibias.t14 gnd.t21 gnd.t20 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X110 a_n2982_13878.t69 minus.t10 a_n3827_n3924.t51 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X111 vdd.t133 vdd.t131 vdd.t132 vdd.t124 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X112 CSoutput.t155 a_n7636_8799.t60 vdd.t199 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X113 vdd.t130 vdd.t127 vdd.t129 vdd.t128 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X114 gnd.t363 commonsourceibias.t110 CSoutput.t89 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X115 a_n2804_13878.t19 a_n2982_13878.t28 a_n2982_13878.t29 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X116 a_n3827_n3924.t50 minus.t11 a_n2982_13878.t68 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X117 vdd.t56 a_n2982_13878.t81 a_n2982_8322.t7 vdd.t55 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X118 gnd.t362 commonsourceibias.t50 commonsourceibias.t51 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X119 a_n2982_13878.t25 a_n2982_13878.t24 a_n2804_13878.t18 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X120 CSoutput.t88 commonsourceibias.t111 gnd.t361 gnd.t256 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X121 CSoutput.t87 commonsourceibias.t112 gnd.t360 gnd.t307 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X122 a_n2982_8322.t6 a_n2982_13878.t82 vdd.t41 vdd.t40 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X123 a_n3827_n3924.t57 diffpairibias.t23 gnd.t415 gnd.t414 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X124 CSoutput.t154 a_n7636_8799.t61 vdd.t198 vdd.t177 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X125 gnd.t359 commonsourceibias.t113 CSoutput.t86 gnd.t309 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X126 a_n3827_n3924.t40 minus.t12 a_n2982_13878.t63 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X127 a_n3827_n3924.t34 minus.t13 a_n2982_13878.t57 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X128 commonsourceibias.t71 commonsourceibias.t70 gnd.t358 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X129 vdd.t54 a_n2982_13878.t83 a_n2804_13878.t27 vdd.t53 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X130 gnd.t357 commonsourceibias.t114 CSoutput.t85 gnd.t283 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X131 commonsourceibias.t69 commonsourceibias.t68 gnd.t356 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X132 a_n2982_13878.t4 minus.t14 a_n3827_n3924.t29 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X133 a_n3827_n3924.t10 plus.t12 a_n7636_8799.t22 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X134 a_n3827_n3924.t28 plus.t13 a_n7636_8799.t21 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X135 vdd.t126 vdd.t123 vdd.t125 vdd.t124 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X136 gnd.t355 commonsourceibias.t66 commonsourceibias.t67 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X137 output.t17 CSoutput.t171 vdd.t65 gnd.t42 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X138 CSoutput.t84 commonsourceibias.t115 gnd.t354 gnd.t269 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X139 gnd.t353 commonsourceibias.t116 CSoutput.t83 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X140 a_n2982_13878.t59 minus.t15 a_n3827_n3924.t36 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X141 a_n2804_13878.t17 a_n2982_13878.t6 a_n2982_13878.t7 vdd.t52 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X142 a_n2982_8322.t23 a_n2982_13878.t84 a_n7636_8799.t43 vdd.t36 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X143 gnd.t165 gnd.t163 plus.t2 gnd.t164 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X144 CSoutput.t82 commonsourceibias.t117 gnd.t352 gnd.t287 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X145 a_n7636_8799.t20 plus.t14 a_n3827_n3924.t25 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X146 a_n7636_8799.t19 plus.t15 a_n3827_n3924.t15 gnd.t413 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X147 vdd.t122 vdd.t120 vdd.t121 vdd.t86 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X148 commonsourceibias.t65 commonsourceibias.t64 gnd.t351 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X149 vdd.t119 vdd.t116 vdd.t118 vdd.t117 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X150 a_n2982_8322.t5 a_n2982_13878.t85 vdd.t51 vdd.t50 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X151 a_n7636_8799.t32 a_n2982_13878.t86 a_n2982_8322.t22 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X152 gnd.t350 commonsourceibias.t118 CSoutput.t81 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X153 CSoutput.t153 a_n7636_8799.t62 vdd.t197 vdd.t166 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X154 diffpairibias.t13 diffpairibias.t12 gnd.t33 gnd.t32 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X155 CSoutput.t172 a_n2982_8322.t36 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X156 vdd.t196 a_n7636_8799.t63 CSoutput.t152 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X157 a_n2982_13878.t0 minus.t16 a_n3827_n3924.t0 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X158 a_n2982_13878.t33 a_n2982_13878.t32 a_n2804_13878.t16 vdd.t30 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X159 a_n7636_8799.t44 a_n2982_13878.t87 a_n2982_8322.t21 vdd.t49 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X160 gnd.t349 commonsourceibias.t62 commonsourceibias.t63 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X161 a_n2804_13878.t15 a_n2982_13878.t14 a_n2982_13878.t15 vdd.t48 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X162 commonsourceibias.t61 commonsourceibias.t60 gnd.t348 gnd.t347 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X163 a_n3827_n3924.t32 minus.t17 a_n2982_13878.t55 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X164 gnd.t346 commonsourceibias.t119 CSoutput.t80 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 gnd.t162 gnd.t160 gnd.t161 gnd.t131 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X166 output.t16 CSoutput.t173 vdd.t66 gnd.t43 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X167 gnd.t345 commonsourceibias.t120 CSoutput.t79 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X168 vdd.t115 vdd.t113 vdd.t114 vdd.t72 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X169 CSoutput.t151 a_n7636_8799.t64 vdd.t194 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X170 gnd.t159 gnd.t156 gnd.t158 gnd.t157 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X171 vdd.t47 a_n2982_13878.t88 a_n2982_8322.t4 vdd.t46 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X172 a_n2804_13878.t14 a_n2982_13878.t40 a_n2982_13878.t41 vdd.t45 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X173 output.t2 outputibias.t9 gnd.t60 gnd.t59 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X174 vdd.t193 a_n7636_8799.t65 CSoutput.t150 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X175 a_n2982_13878.t39 a_n2982_13878.t38 a_n2804_13878.t13 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X176 gnd.t155 gnd.t153 gnd.t154 gnd.t124 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X177 output.t15 CSoutput.t174 vdd.t3 gnd.t17 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X178 minus.t3 gnd.t150 gnd.t152 gnd.t151 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X179 vdd.t4 CSoutput.t175 output.t14 gnd.t18 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X180 CSoutput.t78 commonsourceibias.t121 gnd.t344 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X181 gnd.t343 commonsourceibias.t122 CSoutput.t77 gnd.t265 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X182 commonsourceibias.t59 commonsourceibias.t58 gnd.t342 gnd.t278 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X183 gnd.t341 commonsourceibias.t123 CSoutput.t76 gnd.t263 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X184 a_n3827_n3924.t27 plus.t16 a_n7636_8799.t18 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X185 gnd.t340 commonsourceibias.t124 CSoutput.t75 gnd.t261 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X186 vdd.t192 a_n7636_8799.t66 CSoutput.t149 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X187 a_n3827_n3924.t49 diffpairibias.t24 gnd.t74 gnd.t73 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X188 a_n3827_n3924.t53 diffpairibias.t25 gnd.t84 gnd.t83 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X189 vdd.t191 a_n7636_8799.t67 CSoutput.t148 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X190 a_n7636_8799.t17 plus.t17 a_n3827_n3924.t18 gnd.t37 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X191 vdd.t112 vdd.t110 vdd.t111 vdd.t86 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X192 a_n2804_13878.t12 a_n2982_13878.t46 a_n2982_13878.t47 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X193 CSoutput.t176 a_n2982_8322.t35 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X194 a_n2982_8322.t20 a_n2982_13878.t89 a_n7636_8799.t0 vdd.t44 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X195 CSoutput.t147 a_n7636_8799.t68 vdd.t190 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X196 CSoutput.t177 a_n2982_8322.t34 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X197 CSoutput.t74 commonsourceibias.t125 gnd.t339 gnd.t322 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X198 output.t13 CSoutput.t178 vdd.t146 gnd.t69 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X199 gnd.t149 gnd.t147 gnd.t148 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X200 gnd.t338 commonsourceibias.t126 CSoutput.t73 gnd.t283 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X201 diffpairibias.t11 diffpairibias.t10 gnd.t62 gnd.t61 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X202 gnd.t146 gnd.t144 gnd.t145 gnd.t113 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X203 a_n2804_13878.t29 a_n2982_13878.t90 vdd.t43 vdd.t42 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X204 vdd.t39 a_n2982_13878.t91 a_n2804_13878.t0 vdd.t38 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X205 gnd.t337 commonsourceibias.t127 CSoutput.t72 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X206 vdd.t109 vdd.t107 vdd.t108 vdd.t94 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X207 CSoutput.t146 a_n7636_8799.t69 vdd.t189 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X208 gnd.t336 commonsourceibias.t128 CSoutput.t71 gnd.t301 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X209 CSoutput.t70 commonsourceibias.t129 gnd.t335 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X210 vdd.t187 a_n7636_8799.t70 CSoutput.t145 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X211 output.t12 CSoutput.t179 vdd.t147 gnd.t70 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X212 vdd.t106 vdd.t104 vdd.t105 vdd.t94 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X213 outputibias.t5 outputibias.t4 gnd.t410 gnd.t409 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X214 plus.t1 gnd.t141 gnd.t143 gnd.t142 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X215 a_n2804_13878.t11 a_n2982_13878.t48 a_n2982_13878.t49 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X216 diffpairibias.t9 diffpairibias.t8 gnd.t11 gnd.t10 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X217 gnd.t210 commonsourceibias.t130 CSoutput.t69 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X218 a_n3827_n3924.t30 minus.t18 a_n2982_13878.t5 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X219 gnd.t334 commonsourceibias.t131 CSoutput.t68 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X220 vdd.t185 a_n7636_8799.t71 CSoutput.t144 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X221 commonsourceibias.t79 commonsourceibias.t78 gnd.t333 gnd.t322 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X222 a_n2982_13878.t66 minus.t19 a_n3827_n3924.t46 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X223 a_n2982_8322.t19 a_n2982_13878.t92 a_n7636_8799.t41 vdd.t5 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X224 a_n2982_13878.t43 a_n2982_13878.t42 a_n2804_13878.t10 vdd.t36 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X225 CSoutput.t143 a_n7636_8799.t72 vdd.t184 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X226 diffpairibias.t7 diffpairibias.t6 gnd.t56 gnd.t55 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X227 vdd.t183 a_n7636_8799.t73 CSoutput.t142 vdd.t182 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X228 a_n2804_13878.t9 a_n2982_13878.t34 a_n2982_13878.t35 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X229 a_n2982_13878.t58 minus.t20 a_n3827_n3924.t35 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X230 a_n2982_13878.t54 minus.t21 a_n3827_n3924.t31 gnd.t27 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X231 vdd.t34 a_n2982_13878.t93 a_n2982_8322.t3 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X232 vdd.t181 a_n7636_8799.t74 CSoutput.t141 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X233 a_n3827_n3924.t37 minus.t22 a_n2982_13878.t60 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X234 CSoutput.t67 commonsourceibias.t132 gnd.t332 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 a_n7636_8799.t16 plus.t18 a_n3827_n3924.t26 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X236 gnd.t140 gnd.t138 gnd.t139 gnd.t131 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X237 commonsourceibias.t77 commonsourceibias.t76 gnd.t331 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X238 commonsourceibias.t75 commonsourceibias.t74 gnd.t330 gnd.t291 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X239 a_n3827_n3924.t43 minus.t23 a_n2982_13878.t64 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X240 gnd.t137 gnd.t134 gnd.t136 gnd.t135 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X241 gnd.t133 gnd.t130 gnd.t132 gnd.t131 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X242 a_n2804_13878.t28 a_n2982_13878.t94 vdd.t32 vdd.t31 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X243 vdd.t63 CSoutput.t180 output.t11 gnd.t40 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X244 CSoutput.t66 commonsourceibias.t133 gnd.t329 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X245 gnd.t318 commonsourceibias.t134 CSoutput.t65 gnd.t309 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X246 gnd.t328 commonsourceibias.t72 commonsourceibias.t73 gnd.t244 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X247 gnd.t129 gnd.t127 minus.t2 gnd.t128 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X248 gnd.t327 commonsourceibias.t135 CSoutput.t64 gnd.t265 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X249 CSoutput.t63 commonsourceibias.t136 gnd.t325 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X250 gnd.t126 gnd.t123 gnd.t125 gnd.t124 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X251 CSoutput.t62 commonsourceibias.t137 gnd.t326 gnd.t307 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X252 vdd.t103 vdd.t100 vdd.t102 vdd.t101 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X253 gnd.t324 commonsourceibias.t138 CSoutput.t61 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X254 CSoutput.t60 commonsourceibias.t139 gnd.t323 gnd.t322 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X255 vdd.t99 vdd.t97 vdd.t98 vdd.t76 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X256 gnd.t122 gnd.t120 gnd.t121 gnd.t113 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X257 a_n3827_n3924.t54 diffpairibias.t26 gnd.t86 gnd.t85 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X258 gnd.t321 commonsourceibias.t140 CSoutput.t59 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X259 a_n2982_8322.t18 a_n2982_13878.t95 a_n7636_8799.t47 vdd.t30 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X260 commonsourceibias.t13 commonsourceibias.t12 gnd.t320 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X261 vdd.t64 CSoutput.t181 output.t10 gnd.t41 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X262 vdd.t96 vdd.t93 vdd.t95 vdd.t94 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X263 vdd.t29 a_n2982_13878.t96 a_n2982_8322.t2 vdd.t28 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X264 CSoutput.t58 commonsourceibias.t141 gnd.t319 gnd.t259 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X265 gnd.t317 commonsourceibias.t142 CSoutput.t57 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X266 a_n7636_8799.t15 plus.t19 a_n3827_n3924.t7 gnd.t66 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X267 CSoutput.t56 commonsourceibias.t143 gnd.t316 gnd.t259 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X268 outputibias.t3 outputibias.t2 gnd.t45 gnd.t44 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X269 gnd.t315 commonsourceibias.t144 CSoutput.t55 gnd.t294 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X270 gnd.t314 commonsourceibias.t145 CSoutput.t54 gnd.t244 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X271 CSoutput.t53 commonsourceibias.t146 gnd.t313 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X272 gnd.t119 gnd.t116 gnd.t118 gnd.t117 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X273 commonsourceibias.t11 commonsourceibias.t10 gnd.t312 gnd.t311 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X274 vdd.t92 vdd.t89 vdd.t91 vdd.t90 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X275 a_n3827_n3924.t21 plus.t20 a_n7636_8799.t14 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X276 vdd.t179 a_n7636_8799.t75 CSoutput.t140 vdd.t150 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X277 CSoutput.t139 a_n7636_8799.t76 vdd.t178 vdd.t177 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X278 CSoutput.t138 a_n7636_8799.t77 vdd.t176 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X279 a_n2804_13878.t8 a_n2982_13878.t16 a_n2982_13878.t17 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X280 CSoutput.t52 commonsourceibias.t147 gnd.t290 gnd.t287 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X281 a_n2982_8322.t17 a_n2982_13878.t97 a_n7636_8799.t38 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X282 output.t1 outputibias.t10 gnd.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X283 diffpairibias.t5 diffpairibias.t4 gnd.t35 gnd.t34 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X284 gnd.t310 commonsourceibias.t148 CSoutput.t51 gnd.t309 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X285 CSoutput.t50 commonsourceibias.t149 gnd.t308 gnd.t307 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X286 gnd.t306 commonsourceibias.t8 commonsourceibias.t9 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X287 gnd.t115 gnd.t112 gnd.t114 gnd.t113 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X288 outputibias.t1 outputibias.t0 gnd.t412 gnd.t411 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X289 commonsourceibias.t7 commonsourceibias.t6 gnd.t305 gnd.t256 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X290 CSoutput.t137 a_n7636_8799.t78 vdd.t175 vdd.t166 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X291 gnd.t304 commonsourceibias.t150 CSoutput.t49 gnd.t294 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X292 a_n3827_n3924.t52 diffpairibias.t27 gnd.t82 gnd.t81 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X293 vdd.t88 vdd.t85 vdd.t87 vdd.t86 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X294 gnd.t303 commonsourceibias.t151 CSoutput.t48 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X295 gnd.t302 commonsourceibias.t152 CSoutput.t47 gnd.t301 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X296 gnd.t300 commonsourceibias.t153 CSoutput.t46 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X297 CSoutput.t182 a_n2982_8322.t33 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X298 a_n2982_8322.t1 a_n2982_13878.t98 vdd.t26 vdd.t25 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X299 gnd.t299 commonsourceibias.t154 CSoutput.t45 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X300 CSoutput.t44 commonsourceibias.t155 gnd.t298 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X301 output.t9 CSoutput.t183 vdd.t0 gnd.t14 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X302 gnd.t297 commonsourceibias.t32 commonsourceibias.t33 gnd.t283 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X303 commonsourceibias.t31 commonsourceibias.t30 gnd.t296 gnd.t269 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X304 vdd.t24 a_n2982_13878.t99 a_n2804_13878.t31 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X305 plus.t0 gnd.t109 gnd.t111 gnd.t110 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X306 CSoutput.t136 a_n7636_8799.t79 vdd.t174 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X307 gnd.t295 commonsourceibias.t156 CSoutput.t43 gnd.t294 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X308 CSoutput.t42 commonsourceibias.t157 gnd.t293 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X309 CSoutput.t41 commonsourceibias.t158 gnd.t292 gnd.t291 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X310 gnd.t289 commonsourceibias.t159 CSoutput.t40 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X311 commonsourceibias.t29 commonsourceibias.t28 gnd.t288 gnd.t287 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X312 gnd.t286 commonsourceibias.t160 CSoutput.t39 gnd.t261 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X313 a_n3827_n3924.t12 plus.t21 a_n7636_8799.t13 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X314 gnd.t285 commonsourceibias.t26 commonsourceibias.t27 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X315 a_n3827_n3924.t39 minus.t24 a_n2982_13878.t62 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X316 a_n2982_8322.t16 a_n2982_13878.t100 a_n7636_8799.t31 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X317 a_n7636_8799.t46 a_n2982_13878.t101 a_n2982_8322.t15 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X318 output.t0 outputibias.t11 gnd.t78 gnd.t77 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X319 gnd.t284 commonsourceibias.t161 CSoutput.t38 gnd.t283 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X320 a_n7636_8799.t12 plus.t22 a_n3827_n3924.t24 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X321 a_n2804_13878.t30 a_n2982_13878.t102 vdd.t21 vdd.t20 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X322 CSoutput.t37 commonsourceibias.t162 gnd.t280 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X323 vdd.t84 vdd.t82 vdd.t83 vdd.t68 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X324 CSoutput.t36 commonsourceibias.t163 gnd.t282 gnd.t278 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X325 vdd.t172 a_n7636_8799.t80 CSoutput.t135 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X326 gnd.t281 commonsourceibias.t164 CSoutput.t35 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X327 CSoutput.t34 commonsourceibias.t165 gnd.t279 gnd.t278 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X328 a_n2982_13878.t56 minus.t25 a_n3827_n3924.t33 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X329 CSoutput.t134 a_n7636_8799.t81 vdd.t171 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X330 a_n2982_13878.t45 a_n2982_13878.t44 a_n2804_13878.t7 vdd.t10 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X331 vdd.t1 CSoutput.t184 output.t8 gnd.t15 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X332 gnd.t277 commonsourceibias.t20 commonsourceibias.t21 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X333 CSoutput.t33 commonsourceibias.t166 gnd.t276 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X334 a_n7636_8799.t33 a_n2982_13878.t103 a_n2982_8322.t14 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X335 CSoutput.t32 commonsourceibias.t167 gnd.t275 gnd.t256 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X336 a_n7636_8799.t30 a_n2982_13878.t104 a_n2982_8322.t13 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X337 CSoutput.t31 commonsourceibias.t168 gnd.t274 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X338 gnd.t273 commonsourceibias.t169 CSoutput.t30 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X339 a_n2982_8322.t12 a_n2982_13878.t105 a_n7636_8799.t39 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X340 a_n7636_8799.t11 plus.t23 a_n3827_n3924.t22 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X341 gnd.t108 gnd.t105 gnd.t107 gnd.t106 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X342 CSoutput.t29 commonsourceibias.t170 gnd.t272 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X343 gnd.t104 gnd.t102 minus.t1 gnd.t103 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X344 a_n3827_n3924.t38 minus.t26 a_n2982_13878.t61 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X345 vdd.t169 a_n7636_8799.t82 CSoutput.t133 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X346 CSoutput.t132 a_n7636_8799.t83 vdd.t167 vdd.t166 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X347 CSoutput.t131 a_n7636_8799.t84 vdd.t165 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X348 CSoutput.t28 commonsourceibias.t171 gnd.t270 gnd.t269 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X349 CSoutput.t27 commonsourceibias.t172 gnd.t268 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X350 gnd.t267 commonsourceibias.t173 CSoutput.t26 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X351 CSoutput.t130 a_n7636_8799.t85 vdd.t164 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X352 a_n2804_13878.t6 a_n2982_13878.t50 a_n2982_13878.t51 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X353 vdd.t163 a_n7636_8799.t86 CSoutput.t129 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X354 output.t7 CSoutput.t185 vdd.t2 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X355 a_n3827_n3924.t19 plus.t24 a_n7636_8799.t10 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X356 gnd.t266 commonsourceibias.t18 commonsourceibias.t19 gnd.t265 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X357 CSoutput.t186 a_n2982_8322.t32 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X358 gnd.t264 commonsourceibias.t16 commonsourceibias.t17 gnd.t263 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X359 gnd.t262 commonsourceibias.t14 commonsourceibias.t15 gnd.t261 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X360 a_n3827_n3924.t4 diffpairibias.t28 gnd.t13 gnd.t12 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X361 vdd.t162 a_n7636_8799.t87 CSoutput.t128 vdd.t150 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X362 CSoutput.t25 commonsourceibias.t174 gnd.t260 gnd.t259 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X363 gnd.t258 commonsourceibias.t175 CSoutput.t24 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X364 CSoutput.t127 a_n7636_8799.t88 vdd.t161 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X365 a_n2982_13878.t53 a_n2982_13878.t52 a_n2804_13878.t5 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X366 a_n7636_8799.t1 a_n2982_13878.t106 a_n2982_8322.t11 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X367 vdd.t160 a_n7636_8799.t89 CSoutput.t126 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X368 CSoutput.t125 a_n7636_8799.t90 vdd.t159 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X369 vdd.t81 vdd.t79 vdd.t80 vdd.t76 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X370 CSoutput.t23 commonsourceibias.t176 gnd.t257 gnd.t256 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X371 a_n7636_8799.t9 plus.t25 a_n3827_n3924.t9 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X372 gnd.t101 gnd.t98 gnd.t100 gnd.t99 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X373 gnd.t255 commonsourceibias.t177 CSoutput.t22 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X374 gnd.t254 commonsourceibias.t178 CSoutput.t21 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X375 gnd.t252 commonsourceibias.t179 CSoutput.t20 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X376 diffpairibias.t3 diffpairibias.t2 gnd.t49 gnd.t48 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X377 gnd.t250 commonsourceibias.t180 CSoutput.t19 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X378 CSoutput.t18 commonsourceibias.t181 gnd.t249 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X379 output.t6 CSoutput.t187 vdd.t144 gnd.t67 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X380 a_n2982_8322.t10 a_n2982_13878.t107 a_n7636_8799.t37 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X381 vdd.t145 CSoutput.t188 output.t5 gnd.t68 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X382 a_n3827_n3924.t5 plus.t26 a_n7636_8799.t8 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X383 gnd.t247 commonsourceibias.t182 CSoutput.t17 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X384 gnd.t245 commonsourceibias.t183 CSoutput.t16 gnd.t244 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X385 vdd.t157 a_n7636_8799.t91 CSoutput.t124 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X386 gnd.t97 gnd.t94 gnd.t96 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X387 gnd.t93 gnd.t90 gnd.t92 gnd.t91 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X388 diffpairibias.t1 diffpairibias.t0 gnd.t76 gnd.t75 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X389 CSoutput.t15 commonsourceibias.t184 gnd.t243 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X390 CSoutput.t14 commonsourceibias.t185 gnd.t241 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X391 gnd.t239 commonsourceibias.t34 commonsourceibias.t35 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X392 a_n3827_n3924.t13 plus.t27 a_n7636_8799.t7 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X393 gnd.t237 commonsourceibias.t186 CSoutput.t13 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X394 vdd.t12 a_n2982_13878.t108 a_n2804_13878.t2 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X395 a_n7636_8799.t6 plus.t28 a_n3827_n3924.t6 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X396 CSoutput.t123 a_n7636_8799.t92 vdd.t155 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X397 a_n3827_n3924.t1 minus.t27 a_n2982_13878.t1 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X398 gnd.t236 commonsourceibias.t187 CSoutput.t12 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X399 vdd.t153 a_n7636_8799.t93 CSoutput.t122 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X400 gnd.t234 commonsourceibias.t24 commonsourceibias.t25 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X401 gnd.t232 commonsourceibias.t188 CSoutput.t11 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X402 CSoutput.t10 commonsourceibias.t189 gnd.t231 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X403 a_n2982_8322.t9 a_n2982_13878.t109 a_n7636_8799.t34 vdd.t10 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X404 gnd.t230 commonsourceibias.t190 CSoutput.t9 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X405 a_n2982_13878.t70 minus.t28 a_n3827_n3924.t55 gnd.t413 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X406 a_n2982_8322.t8 a_n2982_13878.t110 a_n7636_8799.t5 vdd.t9 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X407 CSoutput.t8 commonsourceibias.t191 gnd.t228 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X408 CSoutput.t7 commonsourceibias.t192 gnd.t226 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X409 vdd.t151 a_n7636_8799.t94 CSoutput.t121 vdd.t150 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X410 CSoutput.t120 a_n7636_8799.t95 vdd.t149 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X411 gnd.t224 commonsourceibias.t193 CSoutput.t6 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X412 commonsourceibias.t23 commonsourceibias.t22 gnd.t222 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X413 gnd.t212 commonsourceibias.t194 CSoutput.t5 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X414 CSoutput.t4 commonsourceibias.t195 gnd.t220 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X415 vdd.t78 vdd.t75 vdd.t77 vdd.t76 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X416 a_n2982_8322.t0 a_n2982_13878.t111 vdd.t8 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X417 gnd.t218 commonsourceibias.t196 CSoutput.t3 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X418 a_n2804_13878.t4 a_n2982_13878.t18 a_n2982_13878.t19 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X419 vdd.t143 CSoutput.t189 output.t4 gnd.t54 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X420 minus.t0 gnd.t87 gnd.t89 gnd.t88 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X421 vdd.t74 vdd.t71 vdd.t73 vdd.t72 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X422 a_n3827_n3924.t41 diffpairibias.t29 gnd.t53 gnd.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X423 vdd.t70 vdd.t67 vdd.t69 vdd.t68 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X424 CSoutput.t2 commonsourceibias.t197 gnd.t216 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X425 CSoutput.t1 commonsourceibias.t198 gnd.t214 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X426 a_n2982_13878.t37 a_n2982_13878.t36 a_n2804_13878.t3 vdd.t5 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X427 gnd.t208 commonsourceibias.t199 CSoutput.t0 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
R0 commonsourceibias.n397 commonsourceibias.t184 222.032
R1 commonsourceibias.n281 commonsourceibias.t94 222.032
R2 commonsourceibias.n44 commonsourceibias.t76 222.032
R3 commonsourceibias.n166 commonsourceibias.t100 222.032
R4 commonsourceibias.n875 commonsourceibias.t196 222.032
R5 commonsourceibias.n759 commonsourceibias.t188 222.032
R6 commonsourceibias.n529 commonsourceibias.t40 222.032
R7 commonsourceibias.n645 commonsourceibias.t153 222.032
R8 commonsourceibias.n480 commonsourceibias.t183 207.983
R9 commonsourceibias.n364 commonsourceibias.t145 207.983
R10 commonsourceibias.n127 commonsourceibias.t72 207.983
R11 commonsourceibias.n249 commonsourceibias.t104 207.983
R12 commonsourceibias.n963 commonsourceibias.t93 207.983
R13 commonsourceibias.n847 commonsourceibias.t129 207.983
R14 commonsourceibias.n617 commonsourceibias.t70 207.983
R15 commonsourceibias.n732 commonsourceibias.t191 207.983
R16 commonsourceibias.n396 commonsourceibias.t151 168.701
R17 commonsourceibias.n402 commonsourceibias.t99 168.701
R18 commonsourceibias.n408 commonsourceibias.t81 168.701
R19 commonsourceibias.n392 commonsourceibias.t170 168.701
R20 commonsourceibias.n416 commonsourceibias.t177 168.701
R21 commonsourceibias.n422 commonsourceibias.t92 168.701
R22 commonsourceibias.n387 commonsourceibias.t186 168.701
R23 commonsourceibias.n430 commonsourceibias.t198 168.701
R24 commonsourceibias.n436 commonsourceibias.t130 168.701
R25 commonsourceibias.n382 commonsourceibias.t108 168.701
R26 commonsourceibias.n444 commonsourceibias.t88 168.701
R27 commonsourceibias.n450 commonsourceibias.t141 168.701
R28 commonsourceibias.n377 commonsourceibias.t150 168.701
R29 commonsourceibias.n458 commonsourceibias.t98 168.701
R30 commonsourceibias.n464 commonsourceibias.t199 168.701
R31 commonsourceibias.n372 commonsourceibias.t168 168.701
R32 commonsourceibias.n472 commonsourceibias.t107 168.701
R33 commonsourceibias.n478 commonsourceibias.t89 168.701
R34 commonsourceibias.n362 commonsourceibias.t172 168.701
R35 commonsourceibias.n356 commonsourceibias.t160 168.701
R36 commonsourceibias.n256 commonsourceibias.t146 168.701
R37 commonsourceibias.n348 commonsourceibias.t173 168.701
R38 commonsourceibias.n342 commonsourceibias.t158 168.701
R39 commonsourceibias.n261 commonsourceibias.t144 168.701
R40 commonsourceibias.n334 commonsourceibias.t174 168.701
R41 commonsourceibias.n328 commonsourceibias.t159 168.701
R42 commonsourceibias.n266 commonsourceibias.t185 168.701
R43 commonsourceibias.n320 commonsourceibias.t175 168.701
R44 commonsourceibias.n314 commonsourceibias.t157 168.701
R45 commonsourceibias.n271 commonsourceibias.t190 168.701
R46 commonsourceibias.n306 commonsourceibias.t91 168.701
R47 commonsourceibias.n300 commonsourceibias.t169 168.701
R48 commonsourceibias.n276 commonsourceibias.t82 168.701
R49 commonsourceibias.n292 commonsourceibias.t95 168.701
R50 commonsourceibias.n286 commonsourceibias.t90 168.701
R51 commonsourceibias.n280 commonsourceibias.t80 168.701
R52 commonsourceibias.n125 commonsourceibias.t54 168.701
R53 commonsourceibias.n119 commonsourceibias.t14 168.701
R54 commonsourceibias.n19 commonsourceibias.t64 168.701
R55 commonsourceibias.n111 commonsourceibias.t48 168.701
R56 commonsourceibias.n105 commonsourceibias.t74 168.701
R57 commonsourceibias.n24 commonsourceibias.t36 168.701
R58 commonsourceibias.n97 commonsourceibias.t46 168.701
R59 commonsourceibias.n91 commonsourceibias.t66 168.701
R60 commonsourceibias.n29 commonsourceibias.t2 168.701
R61 commonsourceibias.n83 commonsourceibias.t20 168.701
R62 commonsourceibias.n77 commonsourceibias.t38 168.701
R63 commonsourceibias.n34 commonsourceibias.t0 168.701
R64 commonsourceibias.n69 commonsourceibias.t10 168.701
R65 commonsourceibias.n63 commonsourceibias.t52 168.701
R66 commonsourceibias.n39 commonsourceibias.t56 168.701
R67 commonsourceibias.n55 commonsourceibias.t16 168.701
R68 commonsourceibias.n49 commonsourceibias.t60 168.701
R69 commonsourceibias.n43 commonsourceibias.t24 168.701
R70 commonsourceibias.n247 commonsourceibias.t181 168.701
R71 commonsourceibias.n241 commonsourceibias.t124 168.701
R72 commonsourceibias.n5 commonsourceibias.t197 168.701
R73 commonsourceibias.n233 commonsourceibias.t142 168.701
R74 commonsourceibias.n227 commonsourceibias.t101 168.701
R75 commonsourceibias.n10 commonsourceibias.t156 168.701
R76 commonsourceibias.n219 commonsourceibias.t143 168.701
R77 commonsourceibias.n213 commonsourceibias.t193 168.701
R78 commonsourceibias.n150 commonsourceibias.t136 168.701
R79 commonsourceibias.n151 commonsourceibias.t119 168.701
R80 commonsourceibias.n153 commonsourceibias.t155 168.701
R81 commonsourceibias.n155 commonsourceibias.t140 168.701
R82 commonsourceibias.n191 commonsourceibias.t109 168.701
R83 commonsourceibias.n185 commonsourceibias.t182 168.701
R84 commonsourceibias.n161 commonsourceibias.t166 168.701
R85 commonsourceibias.n177 commonsourceibias.t123 168.701
R86 commonsourceibias.n171 commonsourceibias.t84 168.701
R87 commonsourceibias.n165 commonsourceibias.t131 168.701
R88 commonsourceibias.n874 commonsourceibias.t165 168.701
R89 commonsourceibias.n880 commonsourceibias.t106 168.701
R90 commonsourceibias.n886 commonsourceibias.t87 168.701
R91 commonsourceibias.n888 commonsourceibias.t178 168.701
R92 commonsourceibias.n895 commonsourceibias.t167 168.701
R93 commonsourceibias.n901 commonsourceibias.t116 168.701
R94 commonsourceibias.n903 commonsourceibias.t96 168.701
R95 commonsourceibias.n910 commonsourceibias.t102 168.701
R96 commonsourceibias.n916 commonsourceibias.t121 168.701
R97 commonsourceibias.n918 commonsourceibias.t126 168.701
R98 commonsourceibias.n925 commonsourceibias.t112 168.701
R99 commonsourceibias.n931 commonsourceibias.t179 168.701
R100 commonsourceibias.n933 commonsourceibias.t133 168.701
R101 commonsourceibias.n940 commonsourceibias.t120 168.701
R102 commonsourceibias.n946 commonsourceibias.t103 168.701
R103 commonsourceibias.n948 commonsourceibias.t85 168.701
R104 commonsourceibias.n955 commonsourceibias.t125 168.701
R105 commonsourceibias.n961 commonsourceibias.t113 168.701
R106 commonsourceibias.n758 commonsourceibias.t163 168.701
R107 commonsourceibias.n764 commonsourceibias.t180 168.701
R108 commonsourceibias.n770 commonsourceibias.t189 168.701
R109 commonsourceibias.n772 commonsourceibias.t164 168.701
R110 commonsourceibias.n779 commonsourceibias.t176 168.701
R111 commonsourceibias.n785 commonsourceibias.t194 168.701
R112 commonsourceibias.n787 commonsourceibias.t171 168.701
R113 commonsourceibias.n794 commonsourceibias.t135 168.701
R114 commonsourceibias.n800 commonsourceibias.t195 168.701
R115 commonsourceibias.n802 commonsourceibias.t161 168.701
R116 commonsourceibias.n809 commonsourceibias.t137 168.701
R117 commonsourceibias.n815 commonsourceibias.t154 168.701
R118 commonsourceibias.n817 commonsourceibias.t162 168.701
R119 commonsourceibias.n824 commonsourceibias.t138 168.701
R120 commonsourceibias.n830 commonsourceibias.t147 168.701
R121 commonsourceibias.n832 commonsourceibias.t128 168.701
R122 commonsourceibias.n839 commonsourceibias.t139 168.701
R123 commonsourceibias.n845 commonsourceibias.t148 168.701
R124 commonsourceibias.n528 commonsourceibias.t58 168.701
R125 commonsourceibias.n534 commonsourceibias.t34 168.701
R126 commonsourceibias.n540 commonsourceibias.t68 168.701
R127 commonsourceibias.n542 commonsourceibias.t8 168.701
R128 commonsourceibias.n549 commonsourceibias.t6 168.701
R129 commonsourceibias.n555 commonsourceibias.t62 168.701
R130 commonsourceibias.n557 commonsourceibias.t30 168.701
R131 commonsourceibias.n564 commonsourceibias.t18 168.701
R132 commonsourceibias.n570 commonsourceibias.t12 168.701
R133 commonsourceibias.n572 commonsourceibias.t32 168.701
R134 commonsourceibias.n579 commonsourceibias.t44 168.701
R135 commonsourceibias.n585 commonsourceibias.t26 168.701
R136 commonsourceibias.n587 commonsourceibias.t22 168.701
R137 commonsourceibias.n594 commonsourceibias.t50 168.701
R138 commonsourceibias.n600 commonsourceibias.t28 168.701
R139 commonsourceibias.n602 commonsourceibias.t42 168.701
R140 commonsourceibias.n609 commonsourceibias.t78 168.701
R141 commonsourceibias.n615 commonsourceibias.t4 168.701
R142 commonsourceibias.n730 commonsourceibias.t134 168.701
R143 commonsourceibias.n724 commonsourceibias.t97 168.701
R144 commonsourceibias.n717 commonsourceibias.t152 168.701
R145 commonsourceibias.n715 commonsourceibias.t117 168.701
R146 commonsourceibias.n709 commonsourceibias.t187 168.701
R147 commonsourceibias.n702 commonsourceibias.t132 168.701
R148 commonsourceibias.n700 commonsourceibias.t118 168.701
R149 commonsourceibias.n694 commonsourceibias.t149 168.701
R150 commonsourceibias.n687 commonsourceibias.t114 168.701
R151 commonsourceibias.n644 commonsourceibias.t86 168.701
R152 commonsourceibias.n650 commonsourceibias.t127 168.701
R153 commonsourceibias.n656 commonsourceibias.t192 168.701
R154 commonsourceibias.n658 commonsourceibias.t110 168.701
R155 commonsourceibias.n665 commonsourceibias.t111 168.701
R156 commonsourceibias.n671 commonsourceibias.t83 168.701
R157 commonsourceibias.n635 commonsourceibias.t115 168.701
R158 commonsourceibias.n633 commonsourceibias.t122 168.701
R159 commonsourceibias.n631 commonsourceibias.t105 168.701
R160 commonsourceibias.n479 commonsourceibias.n367 161.3
R161 commonsourceibias.n477 commonsourceibias.n476 161.3
R162 commonsourceibias.n475 commonsourceibias.n368 161.3
R163 commonsourceibias.n474 commonsourceibias.n473 161.3
R164 commonsourceibias.n471 commonsourceibias.n369 161.3
R165 commonsourceibias.n470 commonsourceibias.n469 161.3
R166 commonsourceibias.n468 commonsourceibias.n370 161.3
R167 commonsourceibias.n467 commonsourceibias.n466 161.3
R168 commonsourceibias.n465 commonsourceibias.n371 161.3
R169 commonsourceibias.n463 commonsourceibias.n462 161.3
R170 commonsourceibias.n461 commonsourceibias.n373 161.3
R171 commonsourceibias.n460 commonsourceibias.n459 161.3
R172 commonsourceibias.n457 commonsourceibias.n374 161.3
R173 commonsourceibias.n456 commonsourceibias.n455 161.3
R174 commonsourceibias.n454 commonsourceibias.n375 161.3
R175 commonsourceibias.n453 commonsourceibias.n452 161.3
R176 commonsourceibias.n451 commonsourceibias.n376 161.3
R177 commonsourceibias.n449 commonsourceibias.n448 161.3
R178 commonsourceibias.n447 commonsourceibias.n378 161.3
R179 commonsourceibias.n446 commonsourceibias.n445 161.3
R180 commonsourceibias.n443 commonsourceibias.n379 161.3
R181 commonsourceibias.n442 commonsourceibias.n441 161.3
R182 commonsourceibias.n440 commonsourceibias.n380 161.3
R183 commonsourceibias.n439 commonsourceibias.n438 161.3
R184 commonsourceibias.n437 commonsourceibias.n381 161.3
R185 commonsourceibias.n435 commonsourceibias.n434 161.3
R186 commonsourceibias.n433 commonsourceibias.n383 161.3
R187 commonsourceibias.n432 commonsourceibias.n431 161.3
R188 commonsourceibias.n429 commonsourceibias.n384 161.3
R189 commonsourceibias.n428 commonsourceibias.n427 161.3
R190 commonsourceibias.n426 commonsourceibias.n385 161.3
R191 commonsourceibias.n425 commonsourceibias.n424 161.3
R192 commonsourceibias.n423 commonsourceibias.n386 161.3
R193 commonsourceibias.n421 commonsourceibias.n420 161.3
R194 commonsourceibias.n419 commonsourceibias.n388 161.3
R195 commonsourceibias.n418 commonsourceibias.n417 161.3
R196 commonsourceibias.n415 commonsourceibias.n389 161.3
R197 commonsourceibias.n414 commonsourceibias.n413 161.3
R198 commonsourceibias.n412 commonsourceibias.n390 161.3
R199 commonsourceibias.n411 commonsourceibias.n410 161.3
R200 commonsourceibias.n409 commonsourceibias.n391 161.3
R201 commonsourceibias.n407 commonsourceibias.n406 161.3
R202 commonsourceibias.n405 commonsourceibias.n393 161.3
R203 commonsourceibias.n404 commonsourceibias.n403 161.3
R204 commonsourceibias.n401 commonsourceibias.n394 161.3
R205 commonsourceibias.n400 commonsourceibias.n399 161.3
R206 commonsourceibias.n398 commonsourceibias.n395 161.3
R207 commonsourceibias.n282 commonsourceibias.n279 161.3
R208 commonsourceibias.n284 commonsourceibias.n283 161.3
R209 commonsourceibias.n285 commonsourceibias.n278 161.3
R210 commonsourceibias.n288 commonsourceibias.n287 161.3
R211 commonsourceibias.n289 commonsourceibias.n277 161.3
R212 commonsourceibias.n291 commonsourceibias.n290 161.3
R213 commonsourceibias.n293 commonsourceibias.n275 161.3
R214 commonsourceibias.n295 commonsourceibias.n294 161.3
R215 commonsourceibias.n296 commonsourceibias.n274 161.3
R216 commonsourceibias.n298 commonsourceibias.n297 161.3
R217 commonsourceibias.n299 commonsourceibias.n273 161.3
R218 commonsourceibias.n302 commonsourceibias.n301 161.3
R219 commonsourceibias.n303 commonsourceibias.n272 161.3
R220 commonsourceibias.n305 commonsourceibias.n304 161.3
R221 commonsourceibias.n307 commonsourceibias.n270 161.3
R222 commonsourceibias.n309 commonsourceibias.n308 161.3
R223 commonsourceibias.n310 commonsourceibias.n269 161.3
R224 commonsourceibias.n312 commonsourceibias.n311 161.3
R225 commonsourceibias.n313 commonsourceibias.n268 161.3
R226 commonsourceibias.n316 commonsourceibias.n315 161.3
R227 commonsourceibias.n317 commonsourceibias.n267 161.3
R228 commonsourceibias.n319 commonsourceibias.n318 161.3
R229 commonsourceibias.n321 commonsourceibias.n265 161.3
R230 commonsourceibias.n323 commonsourceibias.n322 161.3
R231 commonsourceibias.n324 commonsourceibias.n264 161.3
R232 commonsourceibias.n326 commonsourceibias.n325 161.3
R233 commonsourceibias.n327 commonsourceibias.n263 161.3
R234 commonsourceibias.n330 commonsourceibias.n329 161.3
R235 commonsourceibias.n331 commonsourceibias.n262 161.3
R236 commonsourceibias.n333 commonsourceibias.n332 161.3
R237 commonsourceibias.n335 commonsourceibias.n260 161.3
R238 commonsourceibias.n337 commonsourceibias.n336 161.3
R239 commonsourceibias.n338 commonsourceibias.n259 161.3
R240 commonsourceibias.n340 commonsourceibias.n339 161.3
R241 commonsourceibias.n341 commonsourceibias.n258 161.3
R242 commonsourceibias.n344 commonsourceibias.n343 161.3
R243 commonsourceibias.n345 commonsourceibias.n257 161.3
R244 commonsourceibias.n347 commonsourceibias.n346 161.3
R245 commonsourceibias.n349 commonsourceibias.n255 161.3
R246 commonsourceibias.n351 commonsourceibias.n350 161.3
R247 commonsourceibias.n352 commonsourceibias.n254 161.3
R248 commonsourceibias.n354 commonsourceibias.n353 161.3
R249 commonsourceibias.n355 commonsourceibias.n253 161.3
R250 commonsourceibias.n358 commonsourceibias.n357 161.3
R251 commonsourceibias.n359 commonsourceibias.n252 161.3
R252 commonsourceibias.n361 commonsourceibias.n360 161.3
R253 commonsourceibias.n363 commonsourceibias.n251 161.3
R254 commonsourceibias.n45 commonsourceibias.n42 161.3
R255 commonsourceibias.n47 commonsourceibias.n46 161.3
R256 commonsourceibias.n48 commonsourceibias.n41 161.3
R257 commonsourceibias.n51 commonsourceibias.n50 161.3
R258 commonsourceibias.n52 commonsourceibias.n40 161.3
R259 commonsourceibias.n54 commonsourceibias.n53 161.3
R260 commonsourceibias.n56 commonsourceibias.n38 161.3
R261 commonsourceibias.n58 commonsourceibias.n57 161.3
R262 commonsourceibias.n59 commonsourceibias.n37 161.3
R263 commonsourceibias.n61 commonsourceibias.n60 161.3
R264 commonsourceibias.n62 commonsourceibias.n36 161.3
R265 commonsourceibias.n65 commonsourceibias.n64 161.3
R266 commonsourceibias.n66 commonsourceibias.n35 161.3
R267 commonsourceibias.n68 commonsourceibias.n67 161.3
R268 commonsourceibias.n70 commonsourceibias.n33 161.3
R269 commonsourceibias.n72 commonsourceibias.n71 161.3
R270 commonsourceibias.n73 commonsourceibias.n32 161.3
R271 commonsourceibias.n75 commonsourceibias.n74 161.3
R272 commonsourceibias.n76 commonsourceibias.n31 161.3
R273 commonsourceibias.n79 commonsourceibias.n78 161.3
R274 commonsourceibias.n80 commonsourceibias.n30 161.3
R275 commonsourceibias.n82 commonsourceibias.n81 161.3
R276 commonsourceibias.n84 commonsourceibias.n28 161.3
R277 commonsourceibias.n86 commonsourceibias.n85 161.3
R278 commonsourceibias.n87 commonsourceibias.n27 161.3
R279 commonsourceibias.n89 commonsourceibias.n88 161.3
R280 commonsourceibias.n90 commonsourceibias.n26 161.3
R281 commonsourceibias.n93 commonsourceibias.n92 161.3
R282 commonsourceibias.n94 commonsourceibias.n25 161.3
R283 commonsourceibias.n96 commonsourceibias.n95 161.3
R284 commonsourceibias.n98 commonsourceibias.n23 161.3
R285 commonsourceibias.n100 commonsourceibias.n99 161.3
R286 commonsourceibias.n101 commonsourceibias.n22 161.3
R287 commonsourceibias.n103 commonsourceibias.n102 161.3
R288 commonsourceibias.n104 commonsourceibias.n21 161.3
R289 commonsourceibias.n107 commonsourceibias.n106 161.3
R290 commonsourceibias.n108 commonsourceibias.n20 161.3
R291 commonsourceibias.n110 commonsourceibias.n109 161.3
R292 commonsourceibias.n112 commonsourceibias.n18 161.3
R293 commonsourceibias.n114 commonsourceibias.n113 161.3
R294 commonsourceibias.n115 commonsourceibias.n17 161.3
R295 commonsourceibias.n117 commonsourceibias.n116 161.3
R296 commonsourceibias.n118 commonsourceibias.n16 161.3
R297 commonsourceibias.n121 commonsourceibias.n120 161.3
R298 commonsourceibias.n122 commonsourceibias.n15 161.3
R299 commonsourceibias.n124 commonsourceibias.n123 161.3
R300 commonsourceibias.n126 commonsourceibias.n14 161.3
R301 commonsourceibias.n167 commonsourceibias.n164 161.3
R302 commonsourceibias.n169 commonsourceibias.n168 161.3
R303 commonsourceibias.n170 commonsourceibias.n163 161.3
R304 commonsourceibias.n173 commonsourceibias.n172 161.3
R305 commonsourceibias.n174 commonsourceibias.n162 161.3
R306 commonsourceibias.n176 commonsourceibias.n175 161.3
R307 commonsourceibias.n178 commonsourceibias.n160 161.3
R308 commonsourceibias.n180 commonsourceibias.n179 161.3
R309 commonsourceibias.n181 commonsourceibias.n159 161.3
R310 commonsourceibias.n183 commonsourceibias.n182 161.3
R311 commonsourceibias.n184 commonsourceibias.n158 161.3
R312 commonsourceibias.n187 commonsourceibias.n186 161.3
R313 commonsourceibias.n188 commonsourceibias.n157 161.3
R314 commonsourceibias.n190 commonsourceibias.n189 161.3
R315 commonsourceibias.n192 commonsourceibias.n156 161.3
R316 commonsourceibias.n194 commonsourceibias.n193 161.3
R317 commonsourceibias.n196 commonsourceibias.n195 161.3
R318 commonsourceibias.n197 commonsourceibias.n154 161.3
R319 commonsourceibias.n199 commonsourceibias.n198 161.3
R320 commonsourceibias.n201 commonsourceibias.n200 161.3
R321 commonsourceibias.n202 commonsourceibias.n152 161.3
R322 commonsourceibias.n204 commonsourceibias.n203 161.3
R323 commonsourceibias.n206 commonsourceibias.n205 161.3
R324 commonsourceibias.n208 commonsourceibias.n207 161.3
R325 commonsourceibias.n209 commonsourceibias.n13 161.3
R326 commonsourceibias.n211 commonsourceibias.n210 161.3
R327 commonsourceibias.n212 commonsourceibias.n12 161.3
R328 commonsourceibias.n215 commonsourceibias.n214 161.3
R329 commonsourceibias.n216 commonsourceibias.n11 161.3
R330 commonsourceibias.n218 commonsourceibias.n217 161.3
R331 commonsourceibias.n220 commonsourceibias.n9 161.3
R332 commonsourceibias.n222 commonsourceibias.n221 161.3
R333 commonsourceibias.n223 commonsourceibias.n8 161.3
R334 commonsourceibias.n225 commonsourceibias.n224 161.3
R335 commonsourceibias.n226 commonsourceibias.n7 161.3
R336 commonsourceibias.n229 commonsourceibias.n228 161.3
R337 commonsourceibias.n230 commonsourceibias.n6 161.3
R338 commonsourceibias.n232 commonsourceibias.n231 161.3
R339 commonsourceibias.n234 commonsourceibias.n4 161.3
R340 commonsourceibias.n236 commonsourceibias.n235 161.3
R341 commonsourceibias.n237 commonsourceibias.n3 161.3
R342 commonsourceibias.n239 commonsourceibias.n238 161.3
R343 commonsourceibias.n240 commonsourceibias.n2 161.3
R344 commonsourceibias.n243 commonsourceibias.n242 161.3
R345 commonsourceibias.n244 commonsourceibias.n1 161.3
R346 commonsourceibias.n246 commonsourceibias.n245 161.3
R347 commonsourceibias.n248 commonsourceibias.n0 161.3
R348 commonsourceibias.n962 commonsourceibias.n850 161.3
R349 commonsourceibias.n960 commonsourceibias.n959 161.3
R350 commonsourceibias.n958 commonsourceibias.n851 161.3
R351 commonsourceibias.n957 commonsourceibias.n956 161.3
R352 commonsourceibias.n954 commonsourceibias.n852 161.3
R353 commonsourceibias.n953 commonsourceibias.n952 161.3
R354 commonsourceibias.n951 commonsourceibias.n853 161.3
R355 commonsourceibias.n950 commonsourceibias.n949 161.3
R356 commonsourceibias.n947 commonsourceibias.n854 161.3
R357 commonsourceibias.n945 commonsourceibias.n944 161.3
R358 commonsourceibias.n943 commonsourceibias.n855 161.3
R359 commonsourceibias.n942 commonsourceibias.n941 161.3
R360 commonsourceibias.n939 commonsourceibias.n856 161.3
R361 commonsourceibias.n938 commonsourceibias.n937 161.3
R362 commonsourceibias.n936 commonsourceibias.n857 161.3
R363 commonsourceibias.n935 commonsourceibias.n934 161.3
R364 commonsourceibias.n932 commonsourceibias.n858 161.3
R365 commonsourceibias.n930 commonsourceibias.n929 161.3
R366 commonsourceibias.n928 commonsourceibias.n859 161.3
R367 commonsourceibias.n927 commonsourceibias.n926 161.3
R368 commonsourceibias.n924 commonsourceibias.n860 161.3
R369 commonsourceibias.n923 commonsourceibias.n922 161.3
R370 commonsourceibias.n921 commonsourceibias.n861 161.3
R371 commonsourceibias.n920 commonsourceibias.n919 161.3
R372 commonsourceibias.n917 commonsourceibias.n862 161.3
R373 commonsourceibias.n915 commonsourceibias.n914 161.3
R374 commonsourceibias.n913 commonsourceibias.n863 161.3
R375 commonsourceibias.n912 commonsourceibias.n911 161.3
R376 commonsourceibias.n909 commonsourceibias.n864 161.3
R377 commonsourceibias.n908 commonsourceibias.n907 161.3
R378 commonsourceibias.n906 commonsourceibias.n865 161.3
R379 commonsourceibias.n905 commonsourceibias.n904 161.3
R380 commonsourceibias.n902 commonsourceibias.n866 161.3
R381 commonsourceibias.n900 commonsourceibias.n899 161.3
R382 commonsourceibias.n898 commonsourceibias.n867 161.3
R383 commonsourceibias.n897 commonsourceibias.n896 161.3
R384 commonsourceibias.n894 commonsourceibias.n868 161.3
R385 commonsourceibias.n893 commonsourceibias.n892 161.3
R386 commonsourceibias.n891 commonsourceibias.n869 161.3
R387 commonsourceibias.n890 commonsourceibias.n889 161.3
R388 commonsourceibias.n887 commonsourceibias.n870 161.3
R389 commonsourceibias.n885 commonsourceibias.n884 161.3
R390 commonsourceibias.n883 commonsourceibias.n871 161.3
R391 commonsourceibias.n882 commonsourceibias.n881 161.3
R392 commonsourceibias.n879 commonsourceibias.n872 161.3
R393 commonsourceibias.n878 commonsourceibias.n877 161.3
R394 commonsourceibias.n876 commonsourceibias.n873 161.3
R395 commonsourceibias.n846 commonsourceibias.n734 161.3
R396 commonsourceibias.n844 commonsourceibias.n843 161.3
R397 commonsourceibias.n842 commonsourceibias.n735 161.3
R398 commonsourceibias.n841 commonsourceibias.n840 161.3
R399 commonsourceibias.n838 commonsourceibias.n736 161.3
R400 commonsourceibias.n837 commonsourceibias.n836 161.3
R401 commonsourceibias.n835 commonsourceibias.n737 161.3
R402 commonsourceibias.n834 commonsourceibias.n833 161.3
R403 commonsourceibias.n831 commonsourceibias.n738 161.3
R404 commonsourceibias.n829 commonsourceibias.n828 161.3
R405 commonsourceibias.n827 commonsourceibias.n739 161.3
R406 commonsourceibias.n826 commonsourceibias.n825 161.3
R407 commonsourceibias.n823 commonsourceibias.n740 161.3
R408 commonsourceibias.n822 commonsourceibias.n821 161.3
R409 commonsourceibias.n820 commonsourceibias.n741 161.3
R410 commonsourceibias.n819 commonsourceibias.n818 161.3
R411 commonsourceibias.n816 commonsourceibias.n742 161.3
R412 commonsourceibias.n814 commonsourceibias.n813 161.3
R413 commonsourceibias.n812 commonsourceibias.n743 161.3
R414 commonsourceibias.n811 commonsourceibias.n810 161.3
R415 commonsourceibias.n808 commonsourceibias.n744 161.3
R416 commonsourceibias.n807 commonsourceibias.n806 161.3
R417 commonsourceibias.n805 commonsourceibias.n745 161.3
R418 commonsourceibias.n804 commonsourceibias.n803 161.3
R419 commonsourceibias.n801 commonsourceibias.n746 161.3
R420 commonsourceibias.n799 commonsourceibias.n798 161.3
R421 commonsourceibias.n797 commonsourceibias.n747 161.3
R422 commonsourceibias.n796 commonsourceibias.n795 161.3
R423 commonsourceibias.n793 commonsourceibias.n748 161.3
R424 commonsourceibias.n792 commonsourceibias.n791 161.3
R425 commonsourceibias.n790 commonsourceibias.n749 161.3
R426 commonsourceibias.n789 commonsourceibias.n788 161.3
R427 commonsourceibias.n786 commonsourceibias.n750 161.3
R428 commonsourceibias.n784 commonsourceibias.n783 161.3
R429 commonsourceibias.n782 commonsourceibias.n751 161.3
R430 commonsourceibias.n781 commonsourceibias.n780 161.3
R431 commonsourceibias.n778 commonsourceibias.n752 161.3
R432 commonsourceibias.n777 commonsourceibias.n776 161.3
R433 commonsourceibias.n775 commonsourceibias.n753 161.3
R434 commonsourceibias.n774 commonsourceibias.n773 161.3
R435 commonsourceibias.n771 commonsourceibias.n754 161.3
R436 commonsourceibias.n769 commonsourceibias.n768 161.3
R437 commonsourceibias.n767 commonsourceibias.n755 161.3
R438 commonsourceibias.n766 commonsourceibias.n765 161.3
R439 commonsourceibias.n763 commonsourceibias.n756 161.3
R440 commonsourceibias.n762 commonsourceibias.n761 161.3
R441 commonsourceibias.n760 commonsourceibias.n757 161.3
R442 commonsourceibias.n616 commonsourceibias.n504 161.3
R443 commonsourceibias.n614 commonsourceibias.n613 161.3
R444 commonsourceibias.n612 commonsourceibias.n505 161.3
R445 commonsourceibias.n611 commonsourceibias.n610 161.3
R446 commonsourceibias.n608 commonsourceibias.n506 161.3
R447 commonsourceibias.n607 commonsourceibias.n606 161.3
R448 commonsourceibias.n605 commonsourceibias.n507 161.3
R449 commonsourceibias.n604 commonsourceibias.n603 161.3
R450 commonsourceibias.n601 commonsourceibias.n508 161.3
R451 commonsourceibias.n599 commonsourceibias.n598 161.3
R452 commonsourceibias.n597 commonsourceibias.n509 161.3
R453 commonsourceibias.n596 commonsourceibias.n595 161.3
R454 commonsourceibias.n593 commonsourceibias.n510 161.3
R455 commonsourceibias.n592 commonsourceibias.n591 161.3
R456 commonsourceibias.n590 commonsourceibias.n511 161.3
R457 commonsourceibias.n589 commonsourceibias.n588 161.3
R458 commonsourceibias.n586 commonsourceibias.n512 161.3
R459 commonsourceibias.n584 commonsourceibias.n583 161.3
R460 commonsourceibias.n582 commonsourceibias.n513 161.3
R461 commonsourceibias.n581 commonsourceibias.n580 161.3
R462 commonsourceibias.n578 commonsourceibias.n514 161.3
R463 commonsourceibias.n577 commonsourceibias.n576 161.3
R464 commonsourceibias.n575 commonsourceibias.n515 161.3
R465 commonsourceibias.n574 commonsourceibias.n573 161.3
R466 commonsourceibias.n571 commonsourceibias.n516 161.3
R467 commonsourceibias.n569 commonsourceibias.n568 161.3
R468 commonsourceibias.n567 commonsourceibias.n517 161.3
R469 commonsourceibias.n566 commonsourceibias.n565 161.3
R470 commonsourceibias.n563 commonsourceibias.n518 161.3
R471 commonsourceibias.n562 commonsourceibias.n561 161.3
R472 commonsourceibias.n560 commonsourceibias.n519 161.3
R473 commonsourceibias.n559 commonsourceibias.n558 161.3
R474 commonsourceibias.n556 commonsourceibias.n520 161.3
R475 commonsourceibias.n554 commonsourceibias.n553 161.3
R476 commonsourceibias.n552 commonsourceibias.n521 161.3
R477 commonsourceibias.n551 commonsourceibias.n550 161.3
R478 commonsourceibias.n548 commonsourceibias.n522 161.3
R479 commonsourceibias.n547 commonsourceibias.n546 161.3
R480 commonsourceibias.n545 commonsourceibias.n523 161.3
R481 commonsourceibias.n544 commonsourceibias.n543 161.3
R482 commonsourceibias.n541 commonsourceibias.n524 161.3
R483 commonsourceibias.n539 commonsourceibias.n538 161.3
R484 commonsourceibias.n537 commonsourceibias.n525 161.3
R485 commonsourceibias.n536 commonsourceibias.n535 161.3
R486 commonsourceibias.n533 commonsourceibias.n526 161.3
R487 commonsourceibias.n532 commonsourceibias.n531 161.3
R488 commonsourceibias.n530 commonsourceibias.n527 161.3
R489 commonsourceibias.n686 commonsourceibias.n685 161.3
R490 commonsourceibias.n684 commonsourceibias.n683 161.3
R491 commonsourceibias.n682 commonsourceibias.n632 161.3
R492 commonsourceibias.n681 commonsourceibias.n680 161.3
R493 commonsourceibias.n679 commonsourceibias.n678 161.3
R494 commonsourceibias.n677 commonsourceibias.n634 161.3
R495 commonsourceibias.n676 commonsourceibias.n675 161.3
R496 commonsourceibias.n674 commonsourceibias.n673 161.3
R497 commonsourceibias.n672 commonsourceibias.n636 161.3
R498 commonsourceibias.n670 commonsourceibias.n669 161.3
R499 commonsourceibias.n668 commonsourceibias.n637 161.3
R500 commonsourceibias.n667 commonsourceibias.n666 161.3
R501 commonsourceibias.n664 commonsourceibias.n638 161.3
R502 commonsourceibias.n663 commonsourceibias.n662 161.3
R503 commonsourceibias.n661 commonsourceibias.n639 161.3
R504 commonsourceibias.n660 commonsourceibias.n659 161.3
R505 commonsourceibias.n657 commonsourceibias.n640 161.3
R506 commonsourceibias.n655 commonsourceibias.n654 161.3
R507 commonsourceibias.n653 commonsourceibias.n641 161.3
R508 commonsourceibias.n652 commonsourceibias.n651 161.3
R509 commonsourceibias.n649 commonsourceibias.n642 161.3
R510 commonsourceibias.n648 commonsourceibias.n647 161.3
R511 commonsourceibias.n646 commonsourceibias.n643 161.3
R512 commonsourceibias.n731 commonsourceibias.n483 161.3
R513 commonsourceibias.n729 commonsourceibias.n728 161.3
R514 commonsourceibias.n727 commonsourceibias.n484 161.3
R515 commonsourceibias.n726 commonsourceibias.n725 161.3
R516 commonsourceibias.n723 commonsourceibias.n485 161.3
R517 commonsourceibias.n722 commonsourceibias.n721 161.3
R518 commonsourceibias.n720 commonsourceibias.n486 161.3
R519 commonsourceibias.n719 commonsourceibias.n718 161.3
R520 commonsourceibias.n716 commonsourceibias.n487 161.3
R521 commonsourceibias.n714 commonsourceibias.n713 161.3
R522 commonsourceibias.n712 commonsourceibias.n488 161.3
R523 commonsourceibias.n711 commonsourceibias.n710 161.3
R524 commonsourceibias.n708 commonsourceibias.n489 161.3
R525 commonsourceibias.n707 commonsourceibias.n706 161.3
R526 commonsourceibias.n705 commonsourceibias.n490 161.3
R527 commonsourceibias.n704 commonsourceibias.n703 161.3
R528 commonsourceibias.n701 commonsourceibias.n491 161.3
R529 commonsourceibias.n699 commonsourceibias.n698 161.3
R530 commonsourceibias.n697 commonsourceibias.n492 161.3
R531 commonsourceibias.n696 commonsourceibias.n695 161.3
R532 commonsourceibias.n693 commonsourceibias.n493 161.3
R533 commonsourceibias.n692 commonsourceibias.n691 161.3
R534 commonsourceibias.n690 commonsourceibias.n494 161.3
R535 commonsourceibias.n689 commonsourceibias.n688 161.3
R536 commonsourceibias.n141 commonsourceibias.n139 81.5057
R537 commonsourceibias.n497 commonsourceibias.n495 81.5057
R538 commonsourceibias.n141 commonsourceibias.n140 80.9324
R539 commonsourceibias.n143 commonsourceibias.n142 80.9324
R540 commonsourceibias.n145 commonsourceibias.n144 80.9324
R541 commonsourceibias.n147 commonsourceibias.n146 80.9324
R542 commonsourceibias.n138 commonsourceibias.n137 80.9324
R543 commonsourceibias.n136 commonsourceibias.n135 80.9324
R544 commonsourceibias.n134 commonsourceibias.n133 80.9324
R545 commonsourceibias.n132 commonsourceibias.n131 80.9324
R546 commonsourceibias.n130 commonsourceibias.n129 80.9324
R547 commonsourceibias.n620 commonsourceibias.n619 80.9324
R548 commonsourceibias.n622 commonsourceibias.n621 80.9324
R549 commonsourceibias.n624 commonsourceibias.n623 80.9324
R550 commonsourceibias.n626 commonsourceibias.n625 80.9324
R551 commonsourceibias.n628 commonsourceibias.n627 80.9324
R552 commonsourceibias.n503 commonsourceibias.n502 80.9324
R553 commonsourceibias.n501 commonsourceibias.n500 80.9324
R554 commonsourceibias.n499 commonsourceibias.n498 80.9324
R555 commonsourceibias.n497 commonsourceibias.n496 80.9324
R556 commonsourceibias.n481 commonsourceibias.n480 80.6037
R557 commonsourceibias.n365 commonsourceibias.n364 80.6037
R558 commonsourceibias.n128 commonsourceibias.n127 80.6037
R559 commonsourceibias.n250 commonsourceibias.n249 80.6037
R560 commonsourceibias.n964 commonsourceibias.n963 80.6037
R561 commonsourceibias.n848 commonsourceibias.n847 80.6037
R562 commonsourceibias.n618 commonsourceibias.n617 80.6037
R563 commonsourceibias.n733 commonsourceibias.n732 80.6037
R564 commonsourceibias.n438 commonsourceibias.n437 56.5617
R565 commonsourceibias.n452 commonsourceibias.n451 56.5617
R566 commonsourceibias.n322 commonsourceibias.n321 56.5617
R567 commonsourceibias.n308 commonsourceibias.n307 56.5617
R568 commonsourceibias.n85 commonsourceibias.n84 56.5617
R569 commonsourceibias.n71 commonsourceibias.n70 56.5617
R570 commonsourceibias.n207 commonsourceibias.n206 56.5617
R571 commonsourceibias.n193 commonsourceibias.n192 56.5617
R572 commonsourceibias.n919 commonsourceibias.n917 56.5617
R573 commonsourceibias.n934 commonsourceibias.n932 56.5617
R574 commonsourceibias.n803 commonsourceibias.n801 56.5617
R575 commonsourceibias.n818 commonsourceibias.n816 56.5617
R576 commonsourceibias.n573 commonsourceibias.n571 56.5617
R577 commonsourceibias.n588 commonsourceibias.n586 56.5617
R578 commonsourceibias.n688 commonsourceibias.n686 56.5617
R579 commonsourceibias.n410 commonsourceibias.n409 56.5617
R580 commonsourceibias.n424 commonsourceibias.n423 56.5617
R581 commonsourceibias.n466 commonsourceibias.n465 56.5617
R582 commonsourceibias.n350 commonsourceibias.n349 56.5617
R583 commonsourceibias.n336 commonsourceibias.n335 56.5617
R584 commonsourceibias.n294 commonsourceibias.n293 56.5617
R585 commonsourceibias.n113 commonsourceibias.n112 56.5617
R586 commonsourceibias.n99 commonsourceibias.n98 56.5617
R587 commonsourceibias.n57 commonsourceibias.n56 56.5617
R588 commonsourceibias.n235 commonsourceibias.n234 56.5617
R589 commonsourceibias.n221 commonsourceibias.n220 56.5617
R590 commonsourceibias.n179 commonsourceibias.n178 56.5617
R591 commonsourceibias.n889 commonsourceibias.n887 56.5617
R592 commonsourceibias.n904 commonsourceibias.n902 56.5617
R593 commonsourceibias.n949 commonsourceibias.n947 56.5617
R594 commonsourceibias.n773 commonsourceibias.n771 56.5617
R595 commonsourceibias.n788 commonsourceibias.n786 56.5617
R596 commonsourceibias.n833 commonsourceibias.n831 56.5617
R597 commonsourceibias.n543 commonsourceibias.n541 56.5617
R598 commonsourceibias.n558 commonsourceibias.n556 56.5617
R599 commonsourceibias.n603 commonsourceibias.n601 56.5617
R600 commonsourceibias.n718 commonsourceibias.n716 56.5617
R601 commonsourceibias.n703 commonsourceibias.n701 56.5617
R602 commonsourceibias.n659 commonsourceibias.n657 56.5617
R603 commonsourceibias.n673 commonsourceibias.n672 56.5617
R604 commonsourceibias.n401 commonsourceibias.n400 51.2335
R605 commonsourceibias.n473 commonsourceibias.n368 51.2335
R606 commonsourceibias.n357 commonsourceibias.n252 51.2335
R607 commonsourceibias.n285 commonsourceibias.n284 51.2335
R608 commonsourceibias.n120 commonsourceibias.n15 51.2335
R609 commonsourceibias.n48 commonsourceibias.n47 51.2335
R610 commonsourceibias.n242 commonsourceibias.n1 51.2335
R611 commonsourceibias.n170 commonsourceibias.n169 51.2335
R612 commonsourceibias.n879 commonsourceibias.n878 51.2335
R613 commonsourceibias.n956 commonsourceibias.n851 51.2335
R614 commonsourceibias.n763 commonsourceibias.n762 51.2335
R615 commonsourceibias.n840 commonsourceibias.n735 51.2335
R616 commonsourceibias.n533 commonsourceibias.n532 51.2335
R617 commonsourceibias.n610 commonsourceibias.n505 51.2335
R618 commonsourceibias.n725 commonsourceibias.n484 51.2335
R619 commonsourceibias.n649 commonsourceibias.n648 51.2335
R620 commonsourceibias.n480 commonsourceibias.n479 50.9056
R621 commonsourceibias.n364 commonsourceibias.n363 50.9056
R622 commonsourceibias.n127 commonsourceibias.n126 50.9056
R623 commonsourceibias.n249 commonsourceibias.n248 50.9056
R624 commonsourceibias.n963 commonsourceibias.n962 50.9056
R625 commonsourceibias.n847 commonsourceibias.n846 50.9056
R626 commonsourceibias.n617 commonsourceibias.n616 50.9056
R627 commonsourceibias.n732 commonsourceibias.n731 50.9056
R628 commonsourceibias.n415 commonsourceibias.n414 50.2647
R629 commonsourceibias.n459 commonsourceibias.n373 50.2647
R630 commonsourceibias.n343 commonsourceibias.n257 50.2647
R631 commonsourceibias.n299 commonsourceibias.n298 50.2647
R632 commonsourceibias.n106 commonsourceibias.n20 50.2647
R633 commonsourceibias.n62 commonsourceibias.n61 50.2647
R634 commonsourceibias.n228 commonsourceibias.n6 50.2647
R635 commonsourceibias.n184 commonsourceibias.n183 50.2647
R636 commonsourceibias.n894 commonsourceibias.n893 50.2647
R637 commonsourceibias.n941 commonsourceibias.n855 50.2647
R638 commonsourceibias.n778 commonsourceibias.n777 50.2647
R639 commonsourceibias.n825 commonsourceibias.n739 50.2647
R640 commonsourceibias.n548 commonsourceibias.n547 50.2647
R641 commonsourceibias.n595 commonsourceibias.n509 50.2647
R642 commonsourceibias.n710 commonsourceibias.n488 50.2647
R643 commonsourceibias.n664 commonsourceibias.n663 50.2647
R644 commonsourceibias.n397 commonsourceibias.n396 49.9027
R645 commonsourceibias.n281 commonsourceibias.n280 49.9027
R646 commonsourceibias.n44 commonsourceibias.n43 49.9027
R647 commonsourceibias.n166 commonsourceibias.n165 49.9027
R648 commonsourceibias.n875 commonsourceibias.n874 49.9027
R649 commonsourceibias.n759 commonsourceibias.n758 49.9027
R650 commonsourceibias.n529 commonsourceibias.n528 49.9027
R651 commonsourceibias.n645 commonsourceibias.n644 49.9027
R652 commonsourceibias.n429 commonsourceibias.n428 49.296
R653 commonsourceibias.n445 commonsourceibias.n378 49.296
R654 commonsourceibias.n329 commonsourceibias.n262 49.296
R655 commonsourceibias.n313 commonsourceibias.n312 49.296
R656 commonsourceibias.n92 commonsourceibias.n25 49.296
R657 commonsourceibias.n76 commonsourceibias.n75 49.296
R658 commonsourceibias.n214 commonsourceibias.n11 49.296
R659 commonsourceibias.n198 commonsourceibias.n197 49.296
R660 commonsourceibias.n909 commonsourceibias.n908 49.296
R661 commonsourceibias.n926 commonsourceibias.n859 49.296
R662 commonsourceibias.n793 commonsourceibias.n792 49.296
R663 commonsourceibias.n810 commonsourceibias.n743 49.296
R664 commonsourceibias.n563 commonsourceibias.n562 49.296
R665 commonsourceibias.n580 commonsourceibias.n513 49.296
R666 commonsourceibias.n695 commonsourceibias.n492 49.296
R667 commonsourceibias.n678 commonsourceibias.n677 49.296
R668 commonsourceibias.n431 commonsourceibias.n383 48.3272
R669 commonsourceibias.n443 commonsourceibias.n442 48.3272
R670 commonsourceibias.n327 commonsourceibias.n326 48.3272
R671 commonsourceibias.n315 commonsourceibias.n267 48.3272
R672 commonsourceibias.n90 commonsourceibias.n89 48.3272
R673 commonsourceibias.n78 commonsourceibias.n30 48.3272
R674 commonsourceibias.n212 commonsourceibias.n211 48.3272
R675 commonsourceibias.n202 commonsourceibias.n201 48.3272
R676 commonsourceibias.n911 commonsourceibias.n863 48.3272
R677 commonsourceibias.n924 commonsourceibias.n923 48.3272
R678 commonsourceibias.n795 commonsourceibias.n747 48.3272
R679 commonsourceibias.n808 commonsourceibias.n807 48.3272
R680 commonsourceibias.n565 commonsourceibias.n517 48.3272
R681 commonsourceibias.n578 commonsourceibias.n577 48.3272
R682 commonsourceibias.n693 commonsourceibias.n692 48.3272
R683 commonsourceibias.n682 commonsourceibias.n681 48.3272
R684 commonsourceibias.n417 commonsourceibias.n388 47.3584
R685 commonsourceibias.n457 commonsourceibias.n456 47.3584
R686 commonsourceibias.n341 commonsourceibias.n340 47.3584
R687 commonsourceibias.n301 commonsourceibias.n272 47.3584
R688 commonsourceibias.n104 commonsourceibias.n103 47.3584
R689 commonsourceibias.n64 commonsourceibias.n35 47.3584
R690 commonsourceibias.n226 commonsourceibias.n225 47.3584
R691 commonsourceibias.n186 commonsourceibias.n157 47.3584
R692 commonsourceibias.n896 commonsourceibias.n867 47.3584
R693 commonsourceibias.n939 commonsourceibias.n938 47.3584
R694 commonsourceibias.n780 commonsourceibias.n751 47.3584
R695 commonsourceibias.n823 commonsourceibias.n822 47.3584
R696 commonsourceibias.n550 commonsourceibias.n521 47.3584
R697 commonsourceibias.n593 commonsourceibias.n592 47.3584
R698 commonsourceibias.n708 commonsourceibias.n707 47.3584
R699 commonsourceibias.n666 commonsourceibias.n637 47.3584
R700 commonsourceibias.n403 commonsourceibias.n393 46.3896
R701 commonsourceibias.n471 commonsourceibias.n470 46.3896
R702 commonsourceibias.n355 commonsourceibias.n354 46.3896
R703 commonsourceibias.n287 commonsourceibias.n277 46.3896
R704 commonsourceibias.n118 commonsourceibias.n117 46.3896
R705 commonsourceibias.n50 commonsourceibias.n40 46.3896
R706 commonsourceibias.n240 commonsourceibias.n239 46.3896
R707 commonsourceibias.n172 commonsourceibias.n162 46.3896
R708 commonsourceibias.n881 commonsourceibias.n871 46.3896
R709 commonsourceibias.n954 commonsourceibias.n953 46.3896
R710 commonsourceibias.n765 commonsourceibias.n755 46.3896
R711 commonsourceibias.n838 commonsourceibias.n837 46.3896
R712 commonsourceibias.n535 commonsourceibias.n525 46.3896
R713 commonsourceibias.n608 commonsourceibias.n607 46.3896
R714 commonsourceibias.n723 commonsourceibias.n722 46.3896
R715 commonsourceibias.n651 commonsourceibias.n641 46.3896
R716 commonsourceibias.n398 commonsourceibias.n397 44.7059
R717 commonsourceibias.n876 commonsourceibias.n875 44.7059
R718 commonsourceibias.n760 commonsourceibias.n759 44.7059
R719 commonsourceibias.n530 commonsourceibias.n529 44.7059
R720 commonsourceibias.n646 commonsourceibias.n645 44.7059
R721 commonsourceibias.n282 commonsourceibias.n281 44.7059
R722 commonsourceibias.n45 commonsourceibias.n44 44.7059
R723 commonsourceibias.n167 commonsourceibias.n166 44.7059
R724 commonsourceibias.n407 commonsourceibias.n393 34.7644
R725 commonsourceibias.n470 commonsourceibias.n370 34.7644
R726 commonsourceibias.n354 commonsourceibias.n254 34.7644
R727 commonsourceibias.n291 commonsourceibias.n277 34.7644
R728 commonsourceibias.n117 commonsourceibias.n17 34.7644
R729 commonsourceibias.n54 commonsourceibias.n40 34.7644
R730 commonsourceibias.n239 commonsourceibias.n3 34.7644
R731 commonsourceibias.n176 commonsourceibias.n162 34.7644
R732 commonsourceibias.n885 commonsourceibias.n871 34.7644
R733 commonsourceibias.n953 commonsourceibias.n853 34.7644
R734 commonsourceibias.n769 commonsourceibias.n755 34.7644
R735 commonsourceibias.n837 commonsourceibias.n737 34.7644
R736 commonsourceibias.n539 commonsourceibias.n525 34.7644
R737 commonsourceibias.n607 commonsourceibias.n507 34.7644
R738 commonsourceibias.n722 commonsourceibias.n486 34.7644
R739 commonsourceibias.n655 commonsourceibias.n641 34.7644
R740 commonsourceibias.n421 commonsourceibias.n388 33.7956
R741 commonsourceibias.n456 commonsourceibias.n375 33.7956
R742 commonsourceibias.n340 commonsourceibias.n259 33.7956
R743 commonsourceibias.n305 commonsourceibias.n272 33.7956
R744 commonsourceibias.n103 commonsourceibias.n22 33.7956
R745 commonsourceibias.n68 commonsourceibias.n35 33.7956
R746 commonsourceibias.n225 commonsourceibias.n8 33.7956
R747 commonsourceibias.n190 commonsourceibias.n157 33.7956
R748 commonsourceibias.n900 commonsourceibias.n867 33.7956
R749 commonsourceibias.n938 commonsourceibias.n857 33.7956
R750 commonsourceibias.n784 commonsourceibias.n751 33.7956
R751 commonsourceibias.n822 commonsourceibias.n741 33.7956
R752 commonsourceibias.n554 commonsourceibias.n521 33.7956
R753 commonsourceibias.n592 commonsourceibias.n511 33.7956
R754 commonsourceibias.n707 commonsourceibias.n490 33.7956
R755 commonsourceibias.n670 commonsourceibias.n637 33.7956
R756 commonsourceibias.n435 commonsourceibias.n383 32.8269
R757 commonsourceibias.n442 commonsourceibias.n380 32.8269
R758 commonsourceibias.n326 commonsourceibias.n264 32.8269
R759 commonsourceibias.n319 commonsourceibias.n267 32.8269
R760 commonsourceibias.n89 commonsourceibias.n27 32.8269
R761 commonsourceibias.n82 commonsourceibias.n30 32.8269
R762 commonsourceibias.n211 commonsourceibias.n13 32.8269
R763 commonsourceibias.n203 commonsourceibias.n202 32.8269
R764 commonsourceibias.n915 commonsourceibias.n863 32.8269
R765 commonsourceibias.n923 commonsourceibias.n861 32.8269
R766 commonsourceibias.n799 commonsourceibias.n747 32.8269
R767 commonsourceibias.n807 commonsourceibias.n745 32.8269
R768 commonsourceibias.n569 commonsourceibias.n517 32.8269
R769 commonsourceibias.n577 commonsourceibias.n515 32.8269
R770 commonsourceibias.n692 commonsourceibias.n494 32.8269
R771 commonsourceibias.n683 commonsourceibias.n682 32.8269
R772 commonsourceibias.n428 commonsourceibias.n385 31.8581
R773 commonsourceibias.n449 commonsourceibias.n378 31.8581
R774 commonsourceibias.n333 commonsourceibias.n262 31.8581
R775 commonsourceibias.n312 commonsourceibias.n269 31.8581
R776 commonsourceibias.n96 commonsourceibias.n25 31.8581
R777 commonsourceibias.n75 commonsourceibias.n32 31.8581
R778 commonsourceibias.n218 commonsourceibias.n11 31.8581
R779 commonsourceibias.n197 commonsourceibias.n196 31.8581
R780 commonsourceibias.n908 commonsourceibias.n865 31.8581
R781 commonsourceibias.n930 commonsourceibias.n859 31.8581
R782 commonsourceibias.n792 commonsourceibias.n749 31.8581
R783 commonsourceibias.n814 commonsourceibias.n743 31.8581
R784 commonsourceibias.n562 commonsourceibias.n519 31.8581
R785 commonsourceibias.n584 commonsourceibias.n513 31.8581
R786 commonsourceibias.n699 commonsourceibias.n492 31.8581
R787 commonsourceibias.n677 commonsourceibias.n676 31.8581
R788 commonsourceibias.n414 commonsourceibias.n390 30.8893
R789 commonsourceibias.n463 commonsourceibias.n373 30.8893
R790 commonsourceibias.n347 commonsourceibias.n257 30.8893
R791 commonsourceibias.n298 commonsourceibias.n274 30.8893
R792 commonsourceibias.n110 commonsourceibias.n20 30.8893
R793 commonsourceibias.n61 commonsourceibias.n37 30.8893
R794 commonsourceibias.n232 commonsourceibias.n6 30.8893
R795 commonsourceibias.n183 commonsourceibias.n159 30.8893
R796 commonsourceibias.n893 commonsourceibias.n869 30.8893
R797 commonsourceibias.n945 commonsourceibias.n855 30.8893
R798 commonsourceibias.n777 commonsourceibias.n753 30.8893
R799 commonsourceibias.n829 commonsourceibias.n739 30.8893
R800 commonsourceibias.n547 commonsourceibias.n523 30.8893
R801 commonsourceibias.n599 commonsourceibias.n509 30.8893
R802 commonsourceibias.n714 commonsourceibias.n488 30.8893
R803 commonsourceibias.n663 commonsourceibias.n639 30.8893
R804 commonsourceibias.n400 commonsourceibias.n395 29.9206
R805 commonsourceibias.n477 commonsourceibias.n368 29.9206
R806 commonsourceibias.n361 commonsourceibias.n252 29.9206
R807 commonsourceibias.n284 commonsourceibias.n279 29.9206
R808 commonsourceibias.n124 commonsourceibias.n15 29.9206
R809 commonsourceibias.n47 commonsourceibias.n42 29.9206
R810 commonsourceibias.n246 commonsourceibias.n1 29.9206
R811 commonsourceibias.n169 commonsourceibias.n164 29.9206
R812 commonsourceibias.n878 commonsourceibias.n873 29.9206
R813 commonsourceibias.n960 commonsourceibias.n851 29.9206
R814 commonsourceibias.n762 commonsourceibias.n757 29.9206
R815 commonsourceibias.n844 commonsourceibias.n735 29.9206
R816 commonsourceibias.n532 commonsourceibias.n527 29.9206
R817 commonsourceibias.n614 commonsourceibias.n505 29.9206
R818 commonsourceibias.n729 commonsourceibias.n484 29.9206
R819 commonsourceibias.n648 commonsourceibias.n643 29.9206
R820 commonsourceibias.n479 commonsourceibias.n478 21.8872
R821 commonsourceibias.n363 commonsourceibias.n362 21.8872
R822 commonsourceibias.n126 commonsourceibias.n125 21.8872
R823 commonsourceibias.n248 commonsourceibias.n247 21.8872
R824 commonsourceibias.n962 commonsourceibias.n961 21.8872
R825 commonsourceibias.n846 commonsourceibias.n845 21.8872
R826 commonsourceibias.n616 commonsourceibias.n615 21.8872
R827 commonsourceibias.n731 commonsourceibias.n730 21.8872
R828 commonsourceibias.n410 commonsourceibias.n392 21.3954
R829 commonsourceibias.n465 commonsourceibias.n464 21.3954
R830 commonsourceibias.n349 commonsourceibias.n348 21.3954
R831 commonsourceibias.n294 commonsourceibias.n276 21.3954
R832 commonsourceibias.n112 commonsourceibias.n111 21.3954
R833 commonsourceibias.n57 commonsourceibias.n39 21.3954
R834 commonsourceibias.n234 commonsourceibias.n233 21.3954
R835 commonsourceibias.n179 commonsourceibias.n161 21.3954
R836 commonsourceibias.n889 commonsourceibias.n888 21.3954
R837 commonsourceibias.n947 commonsourceibias.n946 21.3954
R838 commonsourceibias.n773 commonsourceibias.n772 21.3954
R839 commonsourceibias.n831 commonsourceibias.n830 21.3954
R840 commonsourceibias.n543 commonsourceibias.n542 21.3954
R841 commonsourceibias.n601 commonsourceibias.n600 21.3954
R842 commonsourceibias.n716 commonsourceibias.n715 21.3954
R843 commonsourceibias.n659 commonsourceibias.n658 21.3954
R844 commonsourceibias.n424 commonsourceibias.n387 20.9036
R845 commonsourceibias.n451 commonsourceibias.n450 20.9036
R846 commonsourceibias.n335 commonsourceibias.n334 20.9036
R847 commonsourceibias.n308 commonsourceibias.n271 20.9036
R848 commonsourceibias.n98 commonsourceibias.n97 20.9036
R849 commonsourceibias.n71 commonsourceibias.n34 20.9036
R850 commonsourceibias.n220 commonsourceibias.n219 20.9036
R851 commonsourceibias.n193 commonsourceibias.n155 20.9036
R852 commonsourceibias.n904 commonsourceibias.n903 20.9036
R853 commonsourceibias.n932 commonsourceibias.n931 20.9036
R854 commonsourceibias.n788 commonsourceibias.n787 20.9036
R855 commonsourceibias.n816 commonsourceibias.n815 20.9036
R856 commonsourceibias.n558 commonsourceibias.n557 20.9036
R857 commonsourceibias.n586 commonsourceibias.n585 20.9036
R858 commonsourceibias.n701 commonsourceibias.n700 20.9036
R859 commonsourceibias.n673 commonsourceibias.n635 20.9036
R860 commonsourceibias.n437 commonsourceibias.n436 20.4117
R861 commonsourceibias.n438 commonsourceibias.n382 20.4117
R862 commonsourceibias.n322 commonsourceibias.n266 20.4117
R863 commonsourceibias.n321 commonsourceibias.n320 20.4117
R864 commonsourceibias.n85 commonsourceibias.n29 20.4117
R865 commonsourceibias.n84 commonsourceibias.n83 20.4117
R866 commonsourceibias.n207 commonsourceibias.n150 20.4117
R867 commonsourceibias.n206 commonsourceibias.n151 20.4117
R868 commonsourceibias.n917 commonsourceibias.n916 20.4117
R869 commonsourceibias.n919 commonsourceibias.n918 20.4117
R870 commonsourceibias.n801 commonsourceibias.n800 20.4117
R871 commonsourceibias.n803 commonsourceibias.n802 20.4117
R872 commonsourceibias.n571 commonsourceibias.n570 20.4117
R873 commonsourceibias.n573 commonsourceibias.n572 20.4117
R874 commonsourceibias.n688 commonsourceibias.n687 20.4117
R875 commonsourceibias.n686 commonsourceibias.n631 20.4117
R876 commonsourceibias.n423 commonsourceibias.n422 19.9199
R877 commonsourceibias.n452 commonsourceibias.n377 19.9199
R878 commonsourceibias.n336 commonsourceibias.n261 19.9199
R879 commonsourceibias.n307 commonsourceibias.n306 19.9199
R880 commonsourceibias.n99 commonsourceibias.n24 19.9199
R881 commonsourceibias.n70 commonsourceibias.n69 19.9199
R882 commonsourceibias.n221 commonsourceibias.n10 19.9199
R883 commonsourceibias.n192 commonsourceibias.n191 19.9199
R884 commonsourceibias.n902 commonsourceibias.n901 19.9199
R885 commonsourceibias.n934 commonsourceibias.n933 19.9199
R886 commonsourceibias.n786 commonsourceibias.n785 19.9199
R887 commonsourceibias.n818 commonsourceibias.n817 19.9199
R888 commonsourceibias.n556 commonsourceibias.n555 19.9199
R889 commonsourceibias.n588 commonsourceibias.n587 19.9199
R890 commonsourceibias.n703 commonsourceibias.n702 19.9199
R891 commonsourceibias.n672 commonsourceibias.n671 19.9199
R892 commonsourceibias.n409 commonsourceibias.n408 19.4281
R893 commonsourceibias.n466 commonsourceibias.n372 19.4281
R894 commonsourceibias.n350 commonsourceibias.n256 19.4281
R895 commonsourceibias.n293 commonsourceibias.n292 19.4281
R896 commonsourceibias.n113 commonsourceibias.n19 19.4281
R897 commonsourceibias.n56 commonsourceibias.n55 19.4281
R898 commonsourceibias.n235 commonsourceibias.n5 19.4281
R899 commonsourceibias.n178 commonsourceibias.n177 19.4281
R900 commonsourceibias.n887 commonsourceibias.n886 19.4281
R901 commonsourceibias.n949 commonsourceibias.n948 19.4281
R902 commonsourceibias.n771 commonsourceibias.n770 19.4281
R903 commonsourceibias.n833 commonsourceibias.n832 19.4281
R904 commonsourceibias.n541 commonsourceibias.n540 19.4281
R905 commonsourceibias.n603 commonsourceibias.n602 19.4281
R906 commonsourceibias.n718 commonsourceibias.n717 19.4281
R907 commonsourceibias.n657 commonsourceibias.n656 19.4281
R908 commonsourceibias.n402 commonsourceibias.n401 13.526
R909 commonsourceibias.n473 commonsourceibias.n472 13.526
R910 commonsourceibias.n357 commonsourceibias.n356 13.526
R911 commonsourceibias.n286 commonsourceibias.n285 13.526
R912 commonsourceibias.n120 commonsourceibias.n119 13.526
R913 commonsourceibias.n49 commonsourceibias.n48 13.526
R914 commonsourceibias.n242 commonsourceibias.n241 13.526
R915 commonsourceibias.n171 commonsourceibias.n170 13.526
R916 commonsourceibias.n880 commonsourceibias.n879 13.526
R917 commonsourceibias.n956 commonsourceibias.n955 13.526
R918 commonsourceibias.n764 commonsourceibias.n763 13.526
R919 commonsourceibias.n840 commonsourceibias.n839 13.526
R920 commonsourceibias.n534 commonsourceibias.n533 13.526
R921 commonsourceibias.n610 commonsourceibias.n609 13.526
R922 commonsourceibias.n725 commonsourceibias.n724 13.526
R923 commonsourceibias.n650 commonsourceibias.n649 13.526
R924 commonsourceibias.n130 commonsourceibias.n128 13.2322
R925 commonsourceibias.n620 commonsourceibias.n618 13.2322
R926 commonsourceibias.n416 commonsourceibias.n415 13.0342
R927 commonsourceibias.n459 commonsourceibias.n458 13.0342
R928 commonsourceibias.n343 commonsourceibias.n342 13.0342
R929 commonsourceibias.n300 commonsourceibias.n299 13.0342
R930 commonsourceibias.n106 commonsourceibias.n105 13.0342
R931 commonsourceibias.n63 commonsourceibias.n62 13.0342
R932 commonsourceibias.n228 commonsourceibias.n227 13.0342
R933 commonsourceibias.n185 commonsourceibias.n184 13.0342
R934 commonsourceibias.n895 commonsourceibias.n894 13.0342
R935 commonsourceibias.n941 commonsourceibias.n940 13.0342
R936 commonsourceibias.n779 commonsourceibias.n778 13.0342
R937 commonsourceibias.n825 commonsourceibias.n824 13.0342
R938 commonsourceibias.n549 commonsourceibias.n548 13.0342
R939 commonsourceibias.n595 commonsourceibias.n594 13.0342
R940 commonsourceibias.n710 commonsourceibias.n709 13.0342
R941 commonsourceibias.n665 commonsourceibias.n664 13.0342
R942 commonsourceibias.n430 commonsourceibias.n429 12.5423
R943 commonsourceibias.n445 commonsourceibias.n444 12.5423
R944 commonsourceibias.n329 commonsourceibias.n328 12.5423
R945 commonsourceibias.n314 commonsourceibias.n313 12.5423
R946 commonsourceibias.n92 commonsourceibias.n91 12.5423
R947 commonsourceibias.n77 commonsourceibias.n76 12.5423
R948 commonsourceibias.n214 commonsourceibias.n213 12.5423
R949 commonsourceibias.n198 commonsourceibias.n153 12.5423
R950 commonsourceibias.n910 commonsourceibias.n909 12.5423
R951 commonsourceibias.n926 commonsourceibias.n925 12.5423
R952 commonsourceibias.n794 commonsourceibias.n793 12.5423
R953 commonsourceibias.n810 commonsourceibias.n809 12.5423
R954 commonsourceibias.n564 commonsourceibias.n563 12.5423
R955 commonsourceibias.n580 commonsourceibias.n579 12.5423
R956 commonsourceibias.n695 commonsourceibias.n694 12.5423
R957 commonsourceibias.n678 commonsourceibias.n633 12.5423
R958 commonsourceibias.n431 commonsourceibias.n430 12.0505
R959 commonsourceibias.n444 commonsourceibias.n443 12.0505
R960 commonsourceibias.n328 commonsourceibias.n327 12.0505
R961 commonsourceibias.n315 commonsourceibias.n314 12.0505
R962 commonsourceibias.n91 commonsourceibias.n90 12.0505
R963 commonsourceibias.n78 commonsourceibias.n77 12.0505
R964 commonsourceibias.n213 commonsourceibias.n212 12.0505
R965 commonsourceibias.n201 commonsourceibias.n153 12.0505
R966 commonsourceibias.n911 commonsourceibias.n910 12.0505
R967 commonsourceibias.n925 commonsourceibias.n924 12.0505
R968 commonsourceibias.n795 commonsourceibias.n794 12.0505
R969 commonsourceibias.n809 commonsourceibias.n808 12.0505
R970 commonsourceibias.n565 commonsourceibias.n564 12.0505
R971 commonsourceibias.n579 commonsourceibias.n578 12.0505
R972 commonsourceibias.n694 commonsourceibias.n693 12.0505
R973 commonsourceibias.n681 commonsourceibias.n633 12.0505
R974 commonsourceibias.n417 commonsourceibias.n416 11.5587
R975 commonsourceibias.n458 commonsourceibias.n457 11.5587
R976 commonsourceibias.n342 commonsourceibias.n341 11.5587
R977 commonsourceibias.n301 commonsourceibias.n300 11.5587
R978 commonsourceibias.n105 commonsourceibias.n104 11.5587
R979 commonsourceibias.n64 commonsourceibias.n63 11.5587
R980 commonsourceibias.n227 commonsourceibias.n226 11.5587
R981 commonsourceibias.n186 commonsourceibias.n185 11.5587
R982 commonsourceibias.n896 commonsourceibias.n895 11.5587
R983 commonsourceibias.n940 commonsourceibias.n939 11.5587
R984 commonsourceibias.n780 commonsourceibias.n779 11.5587
R985 commonsourceibias.n824 commonsourceibias.n823 11.5587
R986 commonsourceibias.n550 commonsourceibias.n549 11.5587
R987 commonsourceibias.n594 commonsourceibias.n593 11.5587
R988 commonsourceibias.n709 commonsourceibias.n708 11.5587
R989 commonsourceibias.n666 commonsourceibias.n665 11.5587
R990 commonsourceibias.n403 commonsourceibias.n402 11.0668
R991 commonsourceibias.n472 commonsourceibias.n471 11.0668
R992 commonsourceibias.n356 commonsourceibias.n355 11.0668
R993 commonsourceibias.n287 commonsourceibias.n286 11.0668
R994 commonsourceibias.n119 commonsourceibias.n118 11.0668
R995 commonsourceibias.n50 commonsourceibias.n49 11.0668
R996 commonsourceibias.n241 commonsourceibias.n240 11.0668
R997 commonsourceibias.n172 commonsourceibias.n171 11.0668
R998 commonsourceibias.n881 commonsourceibias.n880 11.0668
R999 commonsourceibias.n955 commonsourceibias.n954 11.0668
R1000 commonsourceibias.n765 commonsourceibias.n764 11.0668
R1001 commonsourceibias.n839 commonsourceibias.n838 11.0668
R1002 commonsourceibias.n535 commonsourceibias.n534 11.0668
R1003 commonsourceibias.n609 commonsourceibias.n608 11.0668
R1004 commonsourceibias.n724 commonsourceibias.n723 11.0668
R1005 commonsourceibias.n651 commonsourceibias.n650 11.0668
R1006 commonsourceibias.n966 commonsourceibias.n482 10.4122
R1007 commonsourceibias.n149 commonsourceibias.n148 9.50363
R1008 commonsourceibias.n630 commonsourceibias.n629 9.50363
R1009 commonsourceibias.n366 commonsourceibias.n250 8.76042
R1010 commonsourceibias.n849 commonsourceibias.n733 8.76042
R1011 commonsourceibias.n966 commonsourceibias.n965 8.46921
R1012 commonsourceibias.n408 commonsourceibias.n407 5.16479
R1013 commonsourceibias.n372 commonsourceibias.n370 5.16479
R1014 commonsourceibias.n256 commonsourceibias.n254 5.16479
R1015 commonsourceibias.n292 commonsourceibias.n291 5.16479
R1016 commonsourceibias.n19 commonsourceibias.n17 5.16479
R1017 commonsourceibias.n55 commonsourceibias.n54 5.16479
R1018 commonsourceibias.n5 commonsourceibias.n3 5.16479
R1019 commonsourceibias.n177 commonsourceibias.n176 5.16479
R1020 commonsourceibias.n886 commonsourceibias.n885 5.16479
R1021 commonsourceibias.n948 commonsourceibias.n853 5.16479
R1022 commonsourceibias.n770 commonsourceibias.n769 5.16479
R1023 commonsourceibias.n832 commonsourceibias.n737 5.16479
R1024 commonsourceibias.n540 commonsourceibias.n539 5.16479
R1025 commonsourceibias.n602 commonsourceibias.n507 5.16479
R1026 commonsourceibias.n717 commonsourceibias.n486 5.16479
R1027 commonsourceibias.n656 commonsourceibias.n655 5.16479
R1028 commonsourceibias.n482 commonsourceibias.n481 5.03125
R1029 commonsourceibias.n366 commonsourceibias.n365 5.03125
R1030 commonsourceibias.n965 commonsourceibias.n964 5.03125
R1031 commonsourceibias.n849 commonsourceibias.n848 5.03125
R1032 commonsourceibias.n422 commonsourceibias.n421 4.67295
R1033 commonsourceibias.n377 commonsourceibias.n375 4.67295
R1034 commonsourceibias.n261 commonsourceibias.n259 4.67295
R1035 commonsourceibias.n306 commonsourceibias.n305 4.67295
R1036 commonsourceibias.n24 commonsourceibias.n22 4.67295
R1037 commonsourceibias.n69 commonsourceibias.n68 4.67295
R1038 commonsourceibias.n10 commonsourceibias.n8 4.67295
R1039 commonsourceibias.n191 commonsourceibias.n190 4.67295
R1040 commonsourceibias.n901 commonsourceibias.n900 4.67295
R1041 commonsourceibias.n933 commonsourceibias.n857 4.67295
R1042 commonsourceibias.n785 commonsourceibias.n784 4.67295
R1043 commonsourceibias.n817 commonsourceibias.n741 4.67295
R1044 commonsourceibias.n555 commonsourceibias.n554 4.67295
R1045 commonsourceibias.n587 commonsourceibias.n511 4.67295
R1046 commonsourceibias.n702 commonsourceibias.n490 4.67295
R1047 commonsourceibias.n671 commonsourceibias.n670 4.67295
R1048 commonsourceibias commonsourceibias.n966 4.20978
R1049 commonsourceibias.n436 commonsourceibias.n435 4.18111
R1050 commonsourceibias.n382 commonsourceibias.n380 4.18111
R1051 commonsourceibias.n266 commonsourceibias.n264 4.18111
R1052 commonsourceibias.n320 commonsourceibias.n319 4.18111
R1053 commonsourceibias.n29 commonsourceibias.n27 4.18111
R1054 commonsourceibias.n83 commonsourceibias.n82 4.18111
R1055 commonsourceibias.n150 commonsourceibias.n13 4.18111
R1056 commonsourceibias.n203 commonsourceibias.n151 4.18111
R1057 commonsourceibias.n916 commonsourceibias.n915 4.18111
R1058 commonsourceibias.n918 commonsourceibias.n861 4.18111
R1059 commonsourceibias.n800 commonsourceibias.n799 4.18111
R1060 commonsourceibias.n802 commonsourceibias.n745 4.18111
R1061 commonsourceibias.n570 commonsourceibias.n569 4.18111
R1062 commonsourceibias.n572 commonsourceibias.n515 4.18111
R1063 commonsourceibias.n687 commonsourceibias.n494 4.18111
R1064 commonsourceibias.n683 commonsourceibias.n631 4.18111
R1065 commonsourceibias.n482 commonsourceibias.n366 3.72967
R1066 commonsourceibias.n965 commonsourceibias.n849 3.72967
R1067 commonsourceibias.n387 commonsourceibias.n385 3.68928
R1068 commonsourceibias.n450 commonsourceibias.n449 3.68928
R1069 commonsourceibias.n334 commonsourceibias.n333 3.68928
R1070 commonsourceibias.n271 commonsourceibias.n269 3.68928
R1071 commonsourceibias.n97 commonsourceibias.n96 3.68928
R1072 commonsourceibias.n34 commonsourceibias.n32 3.68928
R1073 commonsourceibias.n219 commonsourceibias.n218 3.68928
R1074 commonsourceibias.n196 commonsourceibias.n155 3.68928
R1075 commonsourceibias.n903 commonsourceibias.n865 3.68928
R1076 commonsourceibias.n931 commonsourceibias.n930 3.68928
R1077 commonsourceibias.n787 commonsourceibias.n749 3.68928
R1078 commonsourceibias.n815 commonsourceibias.n814 3.68928
R1079 commonsourceibias.n557 commonsourceibias.n519 3.68928
R1080 commonsourceibias.n585 commonsourceibias.n584 3.68928
R1081 commonsourceibias.n700 commonsourceibias.n699 3.68928
R1082 commonsourceibias.n676 commonsourceibias.n635 3.68928
R1083 commonsourceibias.n392 commonsourceibias.n390 3.19744
R1084 commonsourceibias.n464 commonsourceibias.n463 3.19744
R1085 commonsourceibias.n348 commonsourceibias.n347 3.19744
R1086 commonsourceibias.n276 commonsourceibias.n274 3.19744
R1087 commonsourceibias.n111 commonsourceibias.n110 3.19744
R1088 commonsourceibias.n39 commonsourceibias.n37 3.19744
R1089 commonsourceibias.n233 commonsourceibias.n232 3.19744
R1090 commonsourceibias.n161 commonsourceibias.n159 3.19744
R1091 commonsourceibias.n888 commonsourceibias.n869 3.19744
R1092 commonsourceibias.n946 commonsourceibias.n945 3.19744
R1093 commonsourceibias.n772 commonsourceibias.n753 3.19744
R1094 commonsourceibias.n830 commonsourceibias.n829 3.19744
R1095 commonsourceibias.n542 commonsourceibias.n523 3.19744
R1096 commonsourceibias.n600 commonsourceibias.n599 3.19744
R1097 commonsourceibias.n715 commonsourceibias.n714 3.19744
R1098 commonsourceibias.n658 commonsourceibias.n639 3.19744
R1099 commonsourceibias.n139 commonsourceibias.t25 2.82907
R1100 commonsourceibias.n139 commonsourceibias.t77 2.82907
R1101 commonsourceibias.n140 commonsourceibias.t17 2.82907
R1102 commonsourceibias.n140 commonsourceibias.t61 2.82907
R1103 commonsourceibias.n142 commonsourceibias.t53 2.82907
R1104 commonsourceibias.n142 commonsourceibias.t57 2.82907
R1105 commonsourceibias.n144 commonsourceibias.t1 2.82907
R1106 commonsourceibias.n144 commonsourceibias.t11 2.82907
R1107 commonsourceibias.n146 commonsourceibias.t21 2.82907
R1108 commonsourceibias.n146 commonsourceibias.t39 2.82907
R1109 commonsourceibias.n137 commonsourceibias.t67 2.82907
R1110 commonsourceibias.n137 commonsourceibias.t3 2.82907
R1111 commonsourceibias.n135 commonsourceibias.t37 2.82907
R1112 commonsourceibias.n135 commonsourceibias.t47 2.82907
R1113 commonsourceibias.n133 commonsourceibias.t49 2.82907
R1114 commonsourceibias.n133 commonsourceibias.t75 2.82907
R1115 commonsourceibias.n131 commonsourceibias.t15 2.82907
R1116 commonsourceibias.n131 commonsourceibias.t65 2.82907
R1117 commonsourceibias.n129 commonsourceibias.t73 2.82907
R1118 commonsourceibias.n129 commonsourceibias.t55 2.82907
R1119 commonsourceibias.n619 commonsourceibias.t5 2.82907
R1120 commonsourceibias.n619 commonsourceibias.t71 2.82907
R1121 commonsourceibias.n621 commonsourceibias.t43 2.82907
R1122 commonsourceibias.n621 commonsourceibias.t79 2.82907
R1123 commonsourceibias.n623 commonsourceibias.t51 2.82907
R1124 commonsourceibias.n623 commonsourceibias.t29 2.82907
R1125 commonsourceibias.n625 commonsourceibias.t27 2.82907
R1126 commonsourceibias.n625 commonsourceibias.t23 2.82907
R1127 commonsourceibias.n627 commonsourceibias.t33 2.82907
R1128 commonsourceibias.n627 commonsourceibias.t45 2.82907
R1129 commonsourceibias.n502 commonsourceibias.t19 2.82907
R1130 commonsourceibias.n502 commonsourceibias.t13 2.82907
R1131 commonsourceibias.n500 commonsourceibias.t63 2.82907
R1132 commonsourceibias.n500 commonsourceibias.t31 2.82907
R1133 commonsourceibias.n498 commonsourceibias.t9 2.82907
R1134 commonsourceibias.n498 commonsourceibias.t7 2.82907
R1135 commonsourceibias.n496 commonsourceibias.t35 2.82907
R1136 commonsourceibias.n496 commonsourceibias.t69 2.82907
R1137 commonsourceibias.n495 commonsourceibias.t41 2.82907
R1138 commonsourceibias.n495 commonsourceibias.t59 2.82907
R1139 commonsourceibias.n396 commonsourceibias.n395 2.7056
R1140 commonsourceibias.n478 commonsourceibias.n477 2.7056
R1141 commonsourceibias.n362 commonsourceibias.n361 2.7056
R1142 commonsourceibias.n280 commonsourceibias.n279 2.7056
R1143 commonsourceibias.n125 commonsourceibias.n124 2.7056
R1144 commonsourceibias.n43 commonsourceibias.n42 2.7056
R1145 commonsourceibias.n247 commonsourceibias.n246 2.7056
R1146 commonsourceibias.n165 commonsourceibias.n164 2.7056
R1147 commonsourceibias.n874 commonsourceibias.n873 2.7056
R1148 commonsourceibias.n961 commonsourceibias.n960 2.7056
R1149 commonsourceibias.n758 commonsourceibias.n757 2.7056
R1150 commonsourceibias.n845 commonsourceibias.n844 2.7056
R1151 commonsourceibias.n528 commonsourceibias.n527 2.7056
R1152 commonsourceibias.n615 commonsourceibias.n614 2.7056
R1153 commonsourceibias.n730 commonsourceibias.n729 2.7056
R1154 commonsourceibias.n644 commonsourceibias.n643 2.7056
R1155 commonsourceibias.n132 commonsourceibias.n130 0.573776
R1156 commonsourceibias.n134 commonsourceibias.n132 0.573776
R1157 commonsourceibias.n136 commonsourceibias.n134 0.573776
R1158 commonsourceibias.n138 commonsourceibias.n136 0.573776
R1159 commonsourceibias.n147 commonsourceibias.n145 0.573776
R1160 commonsourceibias.n145 commonsourceibias.n143 0.573776
R1161 commonsourceibias.n143 commonsourceibias.n141 0.573776
R1162 commonsourceibias.n499 commonsourceibias.n497 0.573776
R1163 commonsourceibias.n501 commonsourceibias.n499 0.573776
R1164 commonsourceibias.n503 commonsourceibias.n501 0.573776
R1165 commonsourceibias.n628 commonsourceibias.n626 0.573776
R1166 commonsourceibias.n626 commonsourceibias.n624 0.573776
R1167 commonsourceibias.n624 commonsourceibias.n622 0.573776
R1168 commonsourceibias.n622 commonsourceibias.n620 0.573776
R1169 commonsourceibias.n148 commonsourceibias.n138 0.287138
R1170 commonsourceibias.n148 commonsourceibias.n147 0.287138
R1171 commonsourceibias.n629 commonsourceibias.n503 0.287138
R1172 commonsourceibias.n629 commonsourceibias.n628 0.287138
R1173 commonsourceibias.n481 commonsourceibias.n367 0.285035
R1174 commonsourceibias.n365 commonsourceibias.n251 0.285035
R1175 commonsourceibias.n128 commonsourceibias.n14 0.285035
R1176 commonsourceibias.n250 commonsourceibias.n0 0.285035
R1177 commonsourceibias.n964 commonsourceibias.n850 0.285035
R1178 commonsourceibias.n848 commonsourceibias.n734 0.285035
R1179 commonsourceibias.n618 commonsourceibias.n504 0.285035
R1180 commonsourceibias.n733 commonsourceibias.n483 0.285035
R1181 commonsourceibias.n476 commonsourceibias.n367 0.189894
R1182 commonsourceibias.n476 commonsourceibias.n475 0.189894
R1183 commonsourceibias.n475 commonsourceibias.n474 0.189894
R1184 commonsourceibias.n474 commonsourceibias.n369 0.189894
R1185 commonsourceibias.n469 commonsourceibias.n369 0.189894
R1186 commonsourceibias.n469 commonsourceibias.n468 0.189894
R1187 commonsourceibias.n468 commonsourceibias.n467 0.189894
R1188 commonsourceibias.n467 commonsourceibias.n371 0.189894
R1189 commonsourceibias.n462 commonsourceibias.n371 0.189894
R1190 commonsourceibias.n462 commonsourceibias.n461 0.189894
R1191 commonsourceibias.n461 commonsourceibias.n460 0.189894
R1192 commonsourceibias.n460 commonsourceibias.n374 0.189894
R1193 commonsourceibias.n455 commonsourceibias.n374 0.189894
R1194 commonsourceibias.n455 commonsourceibias.n454 0.189894
R1195 commonsourceibias.n454 commonsourceibias.n453 0.189894
R1196 commonsourceibias.n453 commonsourceibias.n376 0.189894
R1197 commonsourceibias.n448 commonsourceibias.n376 0.189894
R1198 commonsourceibias.n448 commonsourceibias.n447 0.189894
R1199 commonsourceibias.n447 commonsourceibias.n446 0.189894
R1200 commonsourceibias.n446 commonsourceibias.n379 0.189894
R1201 commonsourceibias.n441 commonsourceibias.n379 0.189894
R1202 commonsourceibias.n441 commonsourceibias.n440 0.189894
R1203 commonsourceibias.n440 commonsourceibias.n439 0.189894
R1204 commonsourceibias.n439 commonsourceibias.n381 0.189894
R1205 commonsourceibias.n434 commonsourceibias.n381 0.189894
R1206 commonsourceibias.n434 commonsourceibias.n433 0.189894
R1207 commonsourceibias.n433 commonsourceibias.n432 0.189894
R1208 commonsourceibias.n432 commonsourceibias.n384 0.189894
R1209 commonsourceibias.n427 commonsourceibias.n384 0.189894
R1210 commonsourceibias.n427 commonsourceibias.n426 0.189894
R1211 commonsourceibias.n426 commonsourceibias.n425 0.189894
R1212 commonsourceibias.n425 commonsourceibias.n386 0.189894
R1213 commonsourceibias.n420 commonsourceibias.n386 0.189894
R1214 commonsourceibias.n420 commonsourceibias.n419 0.189894
R1215 commonsourceibias.n419 commonsourceibias.n418 0.189894
R1216 commonsourceibias.n418 commonsourceibias.n389 0.189894
R1217 commonsourceibias.n413 commonsourceibias.n389 0.189894
R1218 commonsourceibias.n413 commonsourceibias.n412 0.189894
R1219 commonsourceibias.n412 commonsourceibias.n411 0.189894
R1220 commonsourceibias.n411 commonsourceibias.n391 0.189894
R1221 commonsourceibias.n406 commonsourceibias.n391 0.189894
R1222 commonsourceibias.n406 commonsourceibias.n405 0.189894
R1223 commonsourceibias.n405 commonsourceibias.n404 0.189894
R1224 commonsourceibias.n404 commonsourceibias.n394 0.189894
R1225 commonsourceibias.n399 commonsourceibias.n394 0.189894
R1226 commonsourceibias.n399 commonsourceibias.n398 0.189894
R1227 commonsourceibias.n360 commonsourceibias.n251 0.189894
R1228 commonsourceibias.n360 commonsourceibias.n359 0.189894
R1229 commonsourceibias.n359 commonsourceibias.n358 0.189894
R1230 commonsourceibias.n358 commonsourceibias.n253 0.189894
R1231 commonsourceibias.n353 commonsourceibias.n253 0.189894
R1232 commonsourceibias.n353 commonsourceibias.n352 0.189894
R1233 commonsourceibias.n352 commonsourceibias.n351 0.189894
R1234 commonsourceibias.n351 commonsourceibias.n255 0.189894
R1235 commonsourceibias.n346 commonsourceibias.n255 0.189894
R1236 commonsourceibias.n346 commonsourceibias.n345 0.189894
R1237 commonsourceibias.n345 commonsourceibias.n344 0.189894
R1238 commonsourceibias.n344 commonsourceibias.n258 0.189894
R1239 commonsourceibias.n339 commonsourceibias.n258 0.189894
R1240 commonsourceibias.n339 commonsourceibias.n338 0.189894
R1241 commonsourceibias.n338 commonsourceibias.n337 0.189894
R1242 commonsourceibias.n337 commonsourceibias.n260 0.189894
R1243 commonsourceibias.n332 commonsourceibias.n260 0.189894
R1244 commonsourceibias.n332 commonsourceibias.n331 0.189894
R1245 commonsourceibias.n331 commonsourceibias.n330 0.189894
R1246 commonsourceibias.n330 commonsourceibias.n263 0.189894
R1247 commonsourceibias.n325 commonsourceibias.n263 0.189894
R1248 commonsourceibias.n325 commonsourceibias.n324 0.189894
R1249 commonsourceibias.n324 commonsourceibias.n323 0.189894
R1250 commonsourceibias.n323 commonsourceibias.n265 0.189894
R1251 commonsourceibias.n318 commonsourceibias.n265 0.189894
R1252 commonsourceibias.n318 commonsourceibias.n317 0.189894
R1253 commonsourceibias.n317 commonsourceibias.n316 0.189894
R1254 commonsourceibias.n316 commonsourceibias.n268 0.189894
R1255 commonsourceibias.n311 commonsourceibias.n268 0.189894
R1256 commonsourceibias.n311 commonsourceibias.n310 0.189894
R1257 commonsourceibias.n310 commonsourceibias.n309 0.189894
R1258 commonsourceibias.n309 commonsourceibias.n270 0.189894
R1259 commonsourceibias.n304 commonsourceibias.n270 0.189894
R1260 commonsourceibias.n304 commonsourceibias.n303 0.189894
R1261 commonsourceibias.n303 commonsourceibias.n302 0.189894
R1262 commonsourceibias.n302 commonsourceibias.n273 0.189894
R1263 commonsourceibias.n297 commonsourceibias.n273 0.189894
R1264 commonsourceibias.n297 commonsourceibias.n296 0.189894
R1265 commonsourceibias.n296 commonsourceibias.n295 0.189894
R1266 commonsourceibias.n295 commonsourceibias.n275 0.189894
R1267 commonsourceibias.n290 commonsourceibias.n275 0.189894
R1268 commonsourceibias.n290 commonsourceibias.n289 0.189894
R1269 commonsourceibias.n289 commonsourceibias.n288 0.189894
R1270 commonsourceibias.n288 commonsourceibias.n278 0.189894
R1271 commonsourceibias.n283 commonsourceibias.n278 0.189894
R1272 commonsourceibias.n283 commonsourceibias.n282 0.189894
R1273 commonsourceibias.n123 commonsourceibias.n14 0.189894
R1274 commonsourceibias.n123 commonsourceibias.n122 0.189894
R1275 commonsourceibias.n122 commonsourceibias.n121 0.189894
R1276 commonsourceibias.n121 commonsourceibias.n16 0.189894
R1277 commonsourceibias.n116 commonsourceibias.n16 0.189894
R1278 commonsourceibias.n116 commonsourceibias.n115 0.189894
R1279 commonsourceibias.n115 commonsourceibias.n114 0.189894
R1280 commonsourceibias.n114 commonsourceibias.n18 0.189894
R1281 commonsourceibias.n109 commonsourceibias.n18 0.189894
R1282 commonsourceibias.n109 commonsourceibias.n108 0.189894
R1283 commonsourceibias.n108 commonsourceibias.n107 0.189894
R1284 commonsourceibias.n107 commonsourceibias.n21 0.189894
R1285 commonsourceibias.n102 commonsourceibias.n21 0.189894
R1286 commonsourceibias.n102 commonsourceibias.n101 0.189894
R1287 commonsourceibias.n101 commonsourceibias.n100 0.189894
R1288 commonsourceibias.n100 commonsourceibias.n23 0.189894
R1289 commonsourceibias.n95 commonsourceibias.n23 0.189894
R1290 commonsourceibias.n95 commonsourceibias.n94 0.189894
R1291 commonsourceibias.n94 commonsourceibias.n93 0.189894
R1292 commonsourceibias.n93 commonsourceibias.n26 0.189894
R1293 commonsourceibias.n88 commonsourceibias.n26 0.189894
R1294 commonsourceibias.n88 commonsourceibias.n87 0.189894
R1295 commonsourceibias.n87 commonsourceibias.n86 0.189894
R1296 commonsourceibias.n86 commonsourceibias.n28 0.189894
R1297 commonsourceibias.n81 commonsourceibias.n28 0.189894
R1298 commonsourceibias.n81 commonsourceibias.n80 0.189894
R1299 commonsourceibias.n80 commonsourceibias.n79 0.189894
R1300 commonsourceibias.n79 commonsourceibias.n31 0.189894
R1301 commonsourceibias.n74 commonsourceibias.n31 0.189894
R1302 commonsourceibias.n74 commonsourceibias.n73 0.189894
R1303 commonsourceibias.n73 commonsourceibias.n72 0.189894
R1304 commonsourceibias.n72 commonsourceibias.n33 0.189894
R1305 commonsourceibias.n67 commonsourceibias.n33 0.189894
R1306 commonsourceibias.n67 commonsourceibias.n66 0.189894
R1307 commonsourceibias.n66 commonsourceibias.n65 0.189894
R1308 commonsourceibias.n65 commonsourceibias.n36 0.189894
R1309 commonsourceibias.n60 commonsourceibias.n36 0.189894
R1310 commonsourceibias.n60 commonsourceibias.n59 0.189894
R1311 commonsourceibias.n59 commonsourceibias.n58 0.189894
R1312 commonsourceibias.n58 commonsourceibias.n38 0.189894
R1313 commonsourceibias.n53 commonsourceibias.n38 0.189894
R1314 commonsourceibias.n53 commonsourceibias.n52 0.189894
R1315 commonsourceibias.n52 commonsourceibias.n51 0.189894
R1316 commonsourceibias.n51 commonsourceibias.n41 0.189894
R1317 commonsourceibias.n46 commonsourceibias.n41 0.189894
R1318 commonsourceibias.n46 commonsourceibias.n45 0.189894
R1319 commonsourceibias.n205 commonsourceibias.n204 0.189894
R1320 commonsourceibias.n204 commonsourceibias.n152 0.189894
R1321 commonsourceibias.n200 commonsourceibias.n152 0.189894
R1322 commonsourceibias.n200 commonsourceibias.n199 0.189894
R1323 commonsourceibias.n199 commonsourceibias.n154 0.189894
R1324 commonsourceibias.n195 commonsourceibias.n154 0.189894
R1325 commonsourceibias.n195 commonsourceibias.n194 0.189894
R1326 commonsourceibias.n194 commonsourceibias.n156 0.189894
R1327 commonsourceibias.n189 commonsourceibias.n156 0.189894
R1328 commonsourceibias.n189 commonsourceibias.n188 0.189894
R1329 commonsourceibias.n188 commonsourceibias.n187 0.189894
R1330 commonsourceibias.n187 commonsourceibias.n158 0.189894
R1331 commonsourceibias.n182 commonsourceibias.n158 0.189894
R1332 commonsourceibias.n182 commonsourceibias.n181 0.189894
R1333 commonsourceibias.n181 commonsourceibias.n180 0.189894
R1334 commonsourceibias.n180 commonsourceibias.n160 0.189894
R1335 commonsourceibias.n175 commonsourceibias.n160 0.189894
R1336 commonsourceibias.n175 commonsourceibias.n174 0.189894
R1337 commonsourceibias.n174 commonsourceibias.n173 0.189894
R1338 commonsourceibias.n173 commonsourceibias.n163 0.189894
R1339 commonsourceibias.n168 commonsourceibias.n163 0.189894
R1340 commonsourceibias.n168 commonsourceibias.n167 0.189894
R1341 commonsourceibias.n245 commonsourceibias.n0 0.189894
R1342 commonsourceibias.n245 commonsourceibias.n244 0.189894
R1343 commonsourceibias.n244 commonsourceibias.n243 0.189894
R1344 commonsourceibias.n243 commonsourceibias.n2 0.189894
R1345 commonsourceibias.n238 commonsourceibias.n2 0.189894
R1346 commonsourceibias.n238 commonsourceibias.n237 0.189894
R1347 commonsourceibias.n237 commonsourceibias.n236 0.189894
R1348 commonsourceibias.n236 commonsourceibias.n4 0.189894
R1349 commonsourceibias.n231 commonsourceibias.n4 0.189894
R1350 commonsourceibias.n231 commonsourceibias.n230 0.189894
R1351 commonsourceibias.n230 commonsourceibias.n229 0.189894
R1352 commonsourceibias.n229 commonsourceibias.n7 0.189894
R1353 commonsourceibias.n224 commonsourceibias.n7 0.189894
R1354 commonsourceibias.n224 commonsourceibias.n223 0.189894
R1355 commonsourceibias.n223 commonsourceibias.n222 0.189894
R1356 commonsourceibias.n222 commonsourceibias.n9 0.189894
R1357 commonsourceibias.n217 commonsourceibias.n9 0.189894
R1358 commonsourceibias.n217 commonsourceibias.n216 0.189894
R1359 commonsourceibias.n216 commonsourceibias.n215 0.189894
R1360 commonsourceibias.n215 commonsourceibias.n12 0.189894
R1361 commonsourceibias.n210 commonsourceibias.n12 0.189894
R1362 commonsourceibias.n210 commonsourceibias.n209 0.189894
R1363 commonsourceibias.n209 commonsourceibias.n208 0.189894
R1364 commonsourceibias.n877 commonsourceibias.n876 0.189894
R1365 commonsourceibias.n877 commonsourceibias.n872 0.189894
R1366 commonsourceibias.n882 commonsourceibias.n872 0.189894
R1367 commonsourceibias.n883 commonsourceibias.n882 0.189894
R1368 commonsourceibias.n884 commonsourceibias.n883 0.189894
R1369 commonsourceibias.n884 commonsourceibias.n870 0.189894
R1370 commonsourceibias.n890 commonsourceibias.n870 0.189894
R1371 commonsourceibias.n891 commonsourceibias.n890 0.189894
R1372 commonsourceibias.n892 commonsourceibias.n891 0.189894
R1373 commonsourceibias.n892 commonsourceibias.n868 0.189894
R1374 commonsourceibias.n897 commonsourceibias.n868 0.189894
R1375 commonsourceibias.n898 commonsourceibias.n897 0.189894
R1376 commonsourceibias.n899 commonsourceibias.n898 0.189894
R1377 commonsourceibias.n899 commonsourceibias.n866 0.189894
R1378 commonsourceibias.n905 commonsourceibias.n866 0.189894
R1379 commonsourceibias.n906 commonsourceibias.n905 0.189894
R1380 commonsourceibias.n907 commonsourceibias.n906 0.189894
R1381 commonsourceibias.n907 commonsourceibias.n864 0.189894
R1382 commonsourceibias.n912 commonsourceibias.n864 0.189894
R1383 commonsourceibias.n913 commonsourceibias.n912 0.189894
R1384 commonsourceibias.n914 commonsourceibias.n913 0.189894
R1385 commonsourceibias.n914 commonsourceibias.n862 0.189894
R1386 commonsourceibias.n920 commonsourceibias.n862 0.189894
R1387 commonsourceibias.n921 commonsourceibias.n920 0.189894
R1388 commonsourceibias.n922 commonsourceibias.n921 0.189894
R1389 commonsourceibias.n922 commonsourceibias.n860 0.189894
R1390 commonsourceibias.n927 commonsourceibias.n860 0.189894
R1391 commonsourceibias.n928 commonsourceibias.n927 0.189894
R1392 commonsourceibias.n929 commonsourceibias.n928 0.189894
R1393 commonsourceibias.n929 commonsourceibias.n858 0.189894
R1394 commonsourceibias.n935 commonsourceibias.n858 0.189894
R1395 commonsourceibias.n936 commonsourceibias.n935 0.189894
R1396 commonsourceibias.n937 commonsourceibias.n936 0.189894
R1397 commonsourceibias.n937 commonsourceibias.n856 0.189894
R1398 commonsourceibias.n942 commonsourceibias.n856 0.189894
R1399 commonsourceibias.n943 commonsourceibias.n942 0.189894
R1400 commonsourceibias.n944 commonsourceibias.n943 0.189894
R1401 commonsourceibias.n944 commonsourceibias.n854 0.189894
R1402 commonsourceibias.n950 commonsourceibias.n854 0.189894
R1403 commonsourceibias.n951 commonsourceibias.n950 0.189894
R1404 commonsourceibias.n952 commonsourceibias.n951 0.189894
R1405 commonsourceibias.n952 commonsourceibias.n852 0.189894
R1406 commonsourceibias.n957 commonsourceibias.n852 0.189894
R1407 commonsourceibias.n958 commonsourceibias.n957 0.189894
R1408 commonsourceibias.n959 commonsourceibias.n958 0.189894
R1409 commonsourceibias.n959 commonsourceibias.n850 0.189894
R1410 commonsourceibias.n761 commonsourceibias.n760 0.189894
R1411 commonsourceibias.n761 commonsourceibias.n756 0.189894
R1412 commonsourceibias.n766 commonsourceibias.n756 0.189894
R1413 commonsourceibias.n767 commonsourceibias.n766 0.189894
R1414 commonsourceibias.n768 commonsourceibias.n767 0.189894
R1415 commonsourceibias.n768 commonsourceibias.n754 0.189894
R1416 commonsourceibias.n774 commonsourceibias.n754 0.189894
R1417 commonsourceibias.n775 commonsourceibias.n774 0.189894
R1418 commonsourceibias.n776 commonsourceibias.n775 0.189894
R1419 commonsourceibias.n776 commonsourceibias.n752 0.189894
R1420 commonsourceibias.n781 commonsourceibias.n752 0.189894
R1421 commonsourceibias.n782 commonsourceibias.n781 0.189894
R1422 commonsourceibias.n783 commonsourceibias.n782 0.189894
R1423 commonsourceibias.n783 commonsourceibias.n750 0.189894
R1424 commonsourceibias.n789 commonsourceibias.n750 0.189894
R1425 commonsourceibias.n790 commonsourceibias.n789 0.189894
R1426 commonsourceibias.n791 commonsourceibias.n790 0.189894
R1427 commonsourceibias.n791 commonsourceibias.n748 0.189894
R1428 commonsourceibias.n796 commonsourceibias.n748 0.189894
R1429 commonsourceibias.n797 commonsourceibias.n796 0.189894
R1430 commonsourceibias.n798 commonsourceibias.n797 0.189894
R1431 commonsourceibias.n798 commonsourceibias.n746 0.189894
R1432 commonsourceibias.n804 commonsourceibias.n746 0.189894
R1433 commonsourceibias.n805 commonsourceibias.n804 0.189894
R1434 commonsourceibias.n806 commonsourceibias.n805 0.189894
R1435 commonsourceibias.n806 commonsourceibias.n744 0.189894
R1436 commonsourceibias.n811 commonsourceibias.n744 0.189894
R1437 commonsourceibias.n812 commonsourceibias.n811 0.189894
R1438 commonsourceibias.n813 commonsourceibias.n812 0.189894
R1439 commonsourceibias.n813 commonsourceibias.n742 0.189894
R1440 commonsourceibias.n819 commonsourceibias.n742 0.189894
R1441 commonsourceibias.n820 commonsourceibias.n819 0.189894
R1442 commonsourceibias.n821 commonsourceibias.n820 0.189894
R1443 commonsourceibias.n821 commonsourceibias.n740 0.189894
R1444 commonsourceibias.n826 commonsourceibias.n740 0.189894
R1445 commonsourceibias.n827 commonsourceibias.n826 0.189894
R1446 commonsourceibias.n828 commonsourceibias.n827 0.189894
R1447 commonsourceibias.n828 commonsourceibias.n738 0.189894
R1448 commonsourceibias.n834 commonsourceibias.n738 0.189894
R1449 commonsourceibias.n835 commonsourceibias.n834 0.189894
R1450 commonsourceibias.n836 commonsourceibias.n835 0.189894
R1451 commonsourceibias.n836 commonsourceibias.n736 0.189894
R1452 commonsourceibias.n841 commonsourceibias.n736 0.189894
R1453 commonsourceibias.n842 commonsourceibias.n841 0.189894
R1454 commonsourceibias.n843 commonsourceibias.n842 0.189894
R1455 commonsourceibias.n843 commonsourceibias.n734 0.189894
R1456 commonsourceibias.n531 commonsourceibias.n530 0.189894
R1457 commonsourceibias.n531 commonsourceibias.n526 0.189894
R1458 commonsourceibias.n536 commonsourceibias.n526 0.189894
R1459 commonsourceibias.n537 commonsourceibias.n536 0.189894
R1460 commonsourceibias.n538 commonsourceibias.n537 0.189894
R1461 commonsourceibias.n538 commonsourceibias.n524 0.189894
R1462 commonsourceibias.n544 commonsourceibias.n524 0.189894
R1463 commonsourceibias.n545 commonsourceibias.n544 0.189894
R1464 commonsourceibias.n546 commonsourceibias.n545 0.189894
R1465 commonsourceibias.n546 commonsourceibias.n522 0.189894
R1466 commonsourceibias.n551 commonsourceibias.n522 0.189894
R1467 commonsourceibias.n552 commonsourceibias.n551 0.189894
R1468 commonsourceibias.n553 commonsourceibias.n552 0.189894
R1469 commonsourceibias.n553 commonsourceibias.n520 0.189894
R1470 commonsourceibias.n559 commonsourceibias.n520 0.189894
R1471 commonsourceibias.n560 commonsourceibias.n559 0.189894
R1472 commonsourceibias.n561 commonsourceibias.n560 0.189894
R1473 commonsourceibias.n561 commonsourceibias.n518 0.189894
R1474 commonsourceibias.n566 commonsourceibias.n518 0.189894
R1475 commonsourceibias.n567 commonsourceibias.n566 0.189894
R1476 commonsourceibias.n568 commonsourceibias.n567 0.189894
R1477 commonsourceibias.n568 commonsourceibias.n516 0.189894
R1478 commonsourceibias.n574 commonsourceibias.n516 0.189894
R1479 commonsourceibias.n575 commonsourceibias.n574 0.189894
R1480 commonsourceibias.n576 commonsourceibias.n575 0.189894
R1481 commonsourceibias.n576 commonsourceibias.n514 0.189894
R1482 commonsourceibias.n581 commonsourceibias.n514 0.189894
R1483 commonsourceibias.n582 commonsourceibias.n581 0.189894
R1484 commonsourceibias.n583 commonsourceibias.n582 0.189894
R1485 commonsourceibias.n583 commonsourceibias.n512 0.189894
R1486 commonsourceibias.n589 commonsourceibias.n512 0.189894
R1487 commonsourceibias.n590 commonsourceibias.n589 0.189894
R1488 commonsourceibias.n591 commonsourceibias.n590 0.189894
R1489 commonsourceibias.n591 commonsourceibias.n510 0.189894
R1490 commonsourceibias.n596 commonsourceibias.n510 0.189894
R1491 commonsourceibias.n597 commonsourceibias.n596 0.189894
R1492 commonsourceibias.n598 commonsourceibias.n597 0.189894
R1493 commonsourceibias.n598 commonsourceibias.n508 0.189894
R1494 commonsourceibias.n604 commonsourceibias.n508 0.189894
R1495 commonsourceibias.n605 commonsourceibias.n604 0.189894
R1496 commonsourceibias.n606 commonsourceibias.n605 0.189894
R1497 commonsourceibias.n606 commonsourceibias.n506 0.189894
R1498 commonsourceibias.n611 commonsourceibias.n506 0.189894
R1499 commonsourceibias.n612 commonsourceibias.n611 0.189894
R1500 commonsourceibias.n613 commonsourceibias.n612 0.189894
R1501 commonsourceibias.n613 commonsourceibias.n504 0.189894
R1502 commonsourceibias.n647 commonsourceibias.n646 0.189894
R1503 commonsourceibias.n647 commonsourceibias.n642 0.189894
R1504 commonsourceibias.n652 commonsourceibias.n642 0.189894
R1505 commonsourceibias.n653 commonsourceibias.n652 0.189894
R1506 commonsourceibias.n654 commonsourceibias.n653 0.189894
R1507 commonsourceibias.n654 commonsourceibias.n640 0.189894
R1508 commonsourceibias.n660 commonsourceibias.n640 0.189894
R1509 commonsourceibias.n661 commonsourceibias.n660 0.189894
R1510 commonsourceibias.n662 commonsourceibias.n661 0.189894
R1511 commonsourceibias.n662 commonsourceibias.n638 0.189894
R1512 commonsourceibias.n667 commonsourceibias.n638 0.189894
R1513 commonsourceibias.n668 commonsourceibias.n667 0.189894
R1514 commonsourceibias.n669 commonsourceibias.n668 0.189894
R1515 commonsourceibias.n669 commonsourceibias.n636 0.189894
R1516 commonsourceibias.n674 commonsourceibias.n636 0.189894
R1517 commonsourceibias.n675 commonsourceibias.n674 0.189894
R1518 commonsourceibias.n675 commonsourceibias.n634 0.189894
R1519 commonsourceibias.n679 commonsourceibias.n634 0.189894
R1520 commonsourceibias.n680 commonsourceibias.n679 0.189894
R1521 commonsourceibias.n680 commonsourceibias.n632 0.189894
R1522 commonsourceibias.n684 commonsourceibias.n632 0.189894
R1523 commonsourceibias.n685 commonsourceibias.n684 0.189894
R1524 commonsourceibias.n690 commonsourceibias.n689 0.189894
R1525 commonsourceibias.n691 commonsourceibias.n690 0.189894
R1526 commonsourceibias.n691 commonsourceibias.n493 0.189894
R1527 commonsourceibias.n696 commonsourceibias.n493 0.189894
R1528 commonsourceibias.n697 commonsourceibias.n696 0.189894
R1529 commonsourceibias.n698 commonsourceibias.n697 0.189894
R1530 commonsourceibias.n698 commonsourceibias.n491 0.189894
R1531 commonsourceibias.n704 commonsourceibias.n491 0.189894
R1532 commonsourceibias.n705 commonsourceibias.n704 0.189894
R1533 commonsourceibias.n706 commonsourceibias.n705 0.189894
R1534 commonsourceibias.n706 commonsourceibias.n489 0.189894
R1535 commonsourceibias.n711 commonsourceibias.n489 0.189894
R1536 commonsourceibias.n712 commonsourceibias.n711 0.189894
R1537 commonsourceibias.n713 commonsourceibias.n712 0.189894
R1538 commonsourceibias.n713 commonsourceibias.n487 0.189894
R1539 commonsourceibias.n719 commonsourceibias.n487 0.189894
R1540 commonsourceibias.n720 commonsourceibias.n719 0.189894
R1541 commonsourceibias.n721 commonsourceibias.n720 0.189894
R1542 commonsourceibias.n721 commonsourceibias.n485 0.189894
R1543 commonsourceibias.n726 commonsourceibias.n485 0.189894
R1544 commonsourceibias.n727 commonsourceibias.n726 0.189894
R1545 commonsourceibias.n728 commonsourceibias.n727 0.189894
R1546 commonsourceibias.n728 commonsourceibias.n483 0.189894
R1547 commonsourceibias.n205 commonsourceibias.n149 0.0762576
R1548 commonsourceibias.n208 commonsourceibias.n149 0.0762576
R1549 commonsourceibias.n685 commonsourceibias.n630 0.0762576
R1550 commonsourceibias.n689 commonsourceibias.n630 0.0762576
R1551 gnd.n2609 gnd.n2267 965.481
R1552 gnd.n5312 gnd.n3833 939.716
R1553 gnd.n5220 gnd.n3150 766.379
R1554 gnd.n5223 gnd.n5222 766.379
R1555 gnd.n4462 gnd.n4365 766.379
R1556 gnd.n4458 gnd.n4363 766.379
R1557 gnd.n5311 gnd.n3842 756.769
R1558 gnd.n5214 gnd.n5213 756.769
R1559 gnd.n4555 gnd.n4272 756.769
R1560 gnd.n4553 gnd.n4275 756.769
R1561 gnd.n2946 gnd.n1935 756.769
R1562 gnd.n2608 gnd.n2268 756.769
R1563 gnd.n7517 gnd.n398 756.769
R1564 gnd.n5322 gnd.n1809 756.769
R1565 gnd.n255 gnd.n245 751.963
R1566 gnd.n7724 gnd.n7723 751.963
R1567 gnd.n609 gnd.n553 751.963
R1568 gnd.n7309 gnd.n555 751.963
R1569 gnd.n5615 gnd.n1246 751.963
R1570 gnd.n6154 gnd.n6153 751.963
R1571 gnd.n3474 gnd.n3201 751.963
R1572 gnd.n3430 gnd.n3429 751.963
R1573 gnd.n5740 gnd.n1230 711.122
R1574 gnd.n7093 gnd.n749 711.122
R1575 gnd.n6163 gnd.n1232 711.122
R1576 gnd.n7095 gnd.n744 711.122
R1577 gnd.n7884 gnd.n249 696.707
R1578 gnd.n7760 gnd.n7759 696.707
R1579 gnd.n673 gnd.n552 696.707
R1580 gnd.n7311 gnd.n550 696.707
R1581 gnd.n6151 gnd.n1248 696.707
R1582 gnd.n1588 gnd.n1244 696.707
R1583 gnd.n3711 gnd.n3274 696.707
R1584 gnd.n3831 gnd.n3205 696.707
R1585 gnd.n2946 gnd.n2945 585
R1586 gnd.n2947 gnd.n2946 585
R1587 gnd.n1933 gnd.n1932 585
R1588 gnd.n2948 gnd.n1933 585
R1589 gnd.n2951 gnd.n2950 585
R1590 gnd.n2950 gnd.n2949 585
R1591 gnd.n1930 gnd.n1929 585
R1592 gnd.n1929 gnd.n1928 585
R1593 gnd.n2956 gnd.n2955 585
R1594 gnd.n2957 gnd.n2956 585
R1595 gnd.n1927 gnd.n1926 585
R1596 gnd.n2958 gnd.n1927 585
R1597 gnd.n2961 gnd.n2960 585
R1598 gnd.n2960 gnd.n2959 585
R1599 gnd.n1924 gnd.n1923 585
R1600 gnd.n1923 gnd.n1922 585
R1601 gnd.n2966 gnd.n2965 585
R1602 gnd.n2967 gnd.n2966 585
R1603 gnd.n1921 gnd.n1920 585
R1604 gnd.n2968 gnd.n1921 585
R1605 gnd.n2971 gnd.n2970 585
R1606 gnd.n2970 gnd.n2969 585
R1607 gnd.n1918 gnd.n1917 585
R1608 gnd.n1917 gnd.n1916 585
R1609 gnd.n2976 gnd.n2975 585
R1610 gnd.n2977 gnd.n2976 585
R1611 gnd.n1915 gnd.n1914 585
R1612 gnd.n2978 gnd.n1915 585
R1613 gnd.n2981 gnd.n2980 585
R1614 gnd.n2980 gnd.n2979 585
R1615 gnd.n1912 gnd.n1911 585
R1616 gnd.n1911 gnd.n1910 585
R1617 gnd.n2986 gnd.n2985 585
R1618 gnd.n2987 gnd.n2986 585
R1619 gnd.n1909 gnd.n1908 585
R1620 gnd.n2988 gnd.n1909 585
R1621 gnd.n2991 gnd.n2990 585
R1622 gnd.n2990 gnd.n2989 585
R1623 gnd.n1906 gnd.n1905 585
R1624 gnd.n1905 gnd.n1904 585
R1625 gnd.n2996 gnd.n2995 585
R1626 gnd.n2997 gnd.n2996 585
R1627 gnd.n1903 gnd.n1902 585
R1628 gnd.n2998 gnd.n1903 585
R1629 gnd.n3001 gnd.n3000 585
R1630 gnd.n3000 gnd.n2999 585
R1631 gnd.n1900 gnd.n1899 585
R1632 gnd.n1899 gnd.n1898 585
R1633 gnd.n3006 gnd.n3005 585
R1634 gnd.n3007 gnd.n3006 585
R1635 gnd.n1897 gnd.n1896 585
R1636 gnd.n3008 gnd.n1897 585
R1637 gnd.n3011 gnd.n3010 585
R1638 gnd.n3010 gnd.n3009 585
R1639 gnd.n1894 gnd.n1893 585
R1640 gnd.n1893 gnd.n1892 585
R1641 gnd.n3016 gnd.n3015 585
R1642 gnd.n3017 gnd.n3016 585
R1643 gnd.n1891 gnd.n1890 585
R1644 gnd.n3018 gnd.n1891 585
R1645 gnd.n3021 gnd.n3020 585
R1646 gnd.n3020 gnd.n3019 585
R1647 gnd.n1888 gnd.n1887 585
R1648 gnd.n1887 gnd.n1886 585
R1649 gnd.n3026 gnd.n3025 585
R1650 gnd.n3027 gnd.n3026 585
R1651 gnd.n1885 gnd.n1884 585
R1652 gnd.n3028 gnd.n1885 585
R1653 gnd.n3031 gnd.n3030 585
R1654 gnd.n3030 gnd.n3029 585
R1655 gnd.n1882 gnd.n1881 585
R1656 gnd.n1881 gnd.n1880 585
R1657 gnd.n3036 gnd.n3035 585
R1658 gnd.n3037 gnd.n3036 585
R1659 gnd.n1879 gnd.n1878 585
R1660 gnd.n3038 gnd.n1879 585
R1661 gnd.n3041 gnd.n3040 585
R1662 gnd.n3040 gnd.n3039 585
R1663 gnd.n1876 gnd.n1875 585
R1664 gnd.n1875 gnd.n1874 585
R1665 gnd.n3046 gnd.n3045 585
R1666 gnd.n3047 gnd.n3046 585
R1667 gnd.n1873 gnd.n1872 585
R1668 gnd.n3048 gnd.n1873 585
R1669 gnd.n3051 gnd.n3050 585
R1670 gnd.n3050 gnd.n3049 585
R1671 gnd.n1870 gnd.n1869 585
R1672 gnd.n1869 gnd.n1868 585
R1673 gnd.n3056 gnd.n3055 585
R1674 gnd.n3057 gnd.n3056 585
R1675 gnd.n1867 gnd.n1866 585
R1676 gnd.n3058 gnd.n1867 585
R1677 gnd.n3061 gnd.n3060 585
R1678 gnd.n3060 gnd.n3059 585
R1679 gnd.n1864 gnd.n1863 585
R1680 gnd.n1863 gnd.n1862 585
R1681 gnd.n3066 gnd.n3065 585
R1682 gnd.n3067 gnd.n3066 585
R1683 gnd.n1861 gnd.n1860 585
R1684 gnd.n3068 gnd.n1861 585
R1685 gnd.n3071 gnd.n3070 585
R1686 gnd.n3070 gnd.n3069 585
R1687 gnd.n1858 gnd.n1857 585
R1688 gnd.n1857 gnd.n1856 585
R1689 gnd.n3076 gnd.n3075 585
R1690 gnd.n3077 gnd.n3076 585
R1691 gnd.n1855 gnd.n1854 585
R1692 gnd.n3078 gnd.n1855 585
R1693 gnd.n3081 gnd.n3080 585
R1694 gnd.n3080 gnd.n3079 585
R1695 gnd.n1852 gnd.n1851 585
R1696 gnd.n1851 gnd.n1850 585
R1697 gnd.n3086 gnd.n3085 585
R1698 gnd.n3087 gnd.n3086 585
R1699 gnd.n1849 gnd.n1848 585
R1700 gnd.n3088 gnd.n1849 585
R1701 gnd.n3091 gnd.n3090 585
R1702 gnd.n3090 gnd.n3089 585
R1703 gnd.n1846 gnd.n1845 585
R1704 gnd.n1845 gnd.n1844 585
R1705 gnd.n3096 gnd.n3095 585
R1706 gnd.n3097 gnd.n3096 585
R1707 gnd.n1843 gnd.n1842 585
R1708 gnd.n3098 gnd.n1843 585
R1709 gnd.n3101 gnd.n3100 585
R1710 gnd.n3100 gnd.n3099 585
R1711 gnd.n1840 gnd.n1839 585
R1712 gnd.n1839 gnd.n1838 585
R1713 gnd.n3106 gnd.n3105 585
R1714 gnd.n3107 gnd.n3106 585
R1715 gnd.n1837 gnd.n1836 585
R1716 gnd.n3108 gnd.n1837 585
R1717 gnd.n3111 gnd.n3110 585
R1718 gnd.n3110 gnd.n3109 585
R1719 gnd.n1834 gnd.n1833 585
R1720 gnd.n1833 gnd.n1832 585
R1721 gnd.n3116 gnd.n3115 585
R1722 gnd.n3117 gnd.n3116 585
R1723 gnd.n1831 gnd.n1830 585
R1724 gnd.n3118 gnd.n1831 585
R1725 gnd.n3121 gnd.n3120 585
R1726 gnd.n3120 gnd.n3119 585
R1727 gnd.n1828 gnd.n1827 585
R1728 gnd.n1827 gnd.n1826 585
R1729 gnd.n3126 gnd.n3125 585
R1730 gnd.n3127 gnd.n3126 585
R1731 gnd.n1825 gnd.n1824 585
R1732 gnd.n3128 gnd.n1825 585
R1733 gnd.n3131 gnd.n3130 585
R1734 gnd.n3130 gnd.n3129 585
R1735 gnd.n1822 gnd.n1821 585
R1736 gnd.n1821 gnd.n1820 585
R1737 gnd.n3136 gnd.n3135 585
R1738 gnd.n3137 gnd.n3136 585
R1739 gnd.n1819 gnd.n1818 585
R1740 gnd.n3138 gnd.n1819 585
R1741 gnd.n3141 gnd.n3140 585
R1742 gnd.n3140 gnd.n3139 585
R1743 gnd.n1816 gnd.n1815 585
R1744 gnd.n1815 gnd.n1814 585
R1745 gnd.n3146 gnd.n3145 585
R1746 gnd.n3147 gnd.n3146 585
R1747 gnd.n1813 gnd.n1812 585
R1748 gnd.n3148 gnd.n1813 585
R1749 gnd.n5317 gnd.n5316 585
R1750 gnd.n5316 gnd.n5315 585
R1751 gnd.n1810 gnd.n1808 585
R1752 gnd.n5314 gnd.n1808 585
R1753 gnd.n2942 gnd.n1935 585
R1754 gnd.n1935 gnd.n1934 585
R1755 gnd.n2941 gnd.n2940 585
R1756 gnd.n2940 gnd.n2939 585
R1757 gnd.n1938 gnd.n1937 585
R1758 gnd.n2938 gnd.n1938 585
R1759 gnd.n2936 gnd.n2935 585
R1760 gnd.n2937 gnd.n2936 585
R1761 gnd.n2934 gnd.n1940 585
R1762 gnd.n1940 gnd.n1939 585
R1763 gnd.n2933 gnd.n2932 585
R1764 gnd.n2932 gnd.n2931 585
R1765 gnd.n1946 gnd.n1945 585
R1766 gnd.n2930 gnd.n1946 585
R1767 gnd.n2928 gnd.n2927 585
R1768 gnd.n2929 gnd.n2928 585
R1769 gnd.n2926 gnd.n1948 585
R1770 gnd.n1948 gnd.n1947 585
R1771 gnd.n2925 gnd.n2924 585
R1772 gnd.n2924 gnd.n2923 585
R1773 gnd.n1954 gnd.n1953 585
R1774 gnd.n2922 gnd.n1954 585
R1775 gnd.n2920 gnd.n2919 585
R1776 gnd.n2921 gnd.n2920 585
R1777 gnd.n2918 gnd.n1956 585
R1778 gnd.n1956 gnd.n1955 585
R1779 gnd.n2917 gnd.n2916 585
R1780 gnd.n2916 gnd.n2915 585
R1781 gnd.n1962 gnd.n1961 585
R1782 gnd.n2914 gnd.n1962 585
R1783 gnd.n2912 gnd.n2911 585
R1784 gnd.n2913 gnd.n2912 585
R1785 gnd.n2910 gnd.n1964 585
R1786 gnd.n1964 gnd.n1963 585
R1787 gnd.n2909 gnd.n2908 585
R1788 gnd.n2908 gnd.n2907 585
R1789 gnd.n1970 gnd.n1969 585
R1790 gnd.n2906 gnd.n1970 585
R1791 gnd.n2904 gnd.n2903 585
R1792 gnd.n2905 gnd.n2904 585
R1793 gnd.n2902 gnd.n1972 585
R1794 gnd.n1972 gnd.n1971 585
R1795 gnd.n2901 gnd.n2900 585
R1796 gnd.n2900 gnd.n2899 585
R1797 gnd.n1978 gnd.n1977 585
R1798 gnd.n2898 gnd.n1978 585
R1799 gnd.n2896 gnd.n2895 585
R1800 gnd.n2897 gnd.n2896 585
R1801 gnd.n2894 gnd.n1980 585
R1802 gnd.n1980 gnd.n1979 585
R1803 gnd.n2893 gnd.n2892 585
R1804 gnd.n2892 gnd.n2891 585
R1805 gnd.n1986 gnd.n1985 585
R1806 gnd.n2890 gnd.n1986 585
R1807 gnd.n2888 gnd.n2887 585
R1808 gnd.n2889 gnd.n2888 585
R1809 gnd.n2886 gnd.n1988 585
R1810 gnd.n1988 gnd.n1987 585
R1811 gnd.n2885 gnd.n2884 585
R1812 gnd.n2884 gnd.n2883 585
R1813 gnd.n1994 gnd.n1993 585
R1814 gnd.n2882 gnd.n1994 585
R1815 gnd.n2880 gnd.n2879 585
R1816 gnd.n2881 gnd.n2880 585
R1817 gnd.n2878 gnd.n1996 585
R1818 gnd.n1996 gnd.n1995 585
R1819 gnd.n2877 gnd.n2876 585
R1820 gnd.n2876 gnd.n2875 585
R1821 gnd.n2002 gnd.n2001 585
R1822 gnd.n2874 gnd.n2002 585
R1823 gnd.n2872 gnd.n2871 585
R1824 gnd.n2873 gnd.n2872 585
R1825 gnd.n2870 gnd.n2004 585
R1826 gnd.n2004 gnd.n2003 585
R1827 gnd.n2869 gnd.n2868 585
R1828 gnd.n2868 gnd.n2867 585
R1829 gnd.n2010 gnd.n2009 585
R1830 gnd.n2866 gnd.n2010 585
R1831 gnd.n2864 gnd.n2863 585
R1832 gnd.n2865 gnd.n2864 585
R1833 gnd.n2862 gnd.n2012 585
R1834 gnd.n2012 gnd.n2011 585
R1835 gnd.n2861 gnd.n2860 585
R1836 gnd.n2860 gnd.n2859 585
R1837 gnd.n2018 gnd.n2017 585
R1838 gnd.n2858 gnd.n2018 585
R1839 gnd.n2856 gnd.n2855 585
R1840 gnd.n2857 gnd.n2856 585
R1841 gnd.n2854 gnd.n2020 585
R1842 gnd.n2020 gnd.n2019 585
R1843 gnd.n2853 gnd.n2852 585
R1844 gnd.n2852 gnd.n2851 585
R1845 gnd.n2026 gnd.n2025 585
R1846 gnd.n2850 gnd.n2026 585
R1847 gnd.n2848 gnd.n2847 585
R1848 gnd.n2849 gnd.n2848 585
R1849 gnd.n2846 gnd.n2028 585
R1850 gnd.n2028 gnd.n2027 585
R1851 gnd.n2845 gnd.n2844 585
R1852 gnd.n2844 gnd.n2843 585
R1853 gnd.n2034 gnd.n2033 585
R1854 gnd.n2842 gnd.n2034 585
R1855 gnd.n2840 gnd.n2839 585
R1856 gnd.n2841 gnd.n2840 585
R1857 gnd.n2838 gnd.n2036 585
R1858 gnd.n2036 gnd.n2035 585
R1859 gnd.n2837 gnd.n2836 585
R1860 gnd.n2836 gnd.n2835 585
R1861 gnd.n2042 gnd.n2041 585
R1862 gnd.n2834 gnd.n2042 585
R1863 gnd.n2832 gnd.n2831 585
R1864 gnd.n2833 gnd.n2832 585
R1865 gnd.n2830 gnd.n2044 585
R1866 gnd.n2044 gnd.n2043 585
R1867 gnd.n2829 gnd.n2828 585
R1868 gnd.n2828 gnd.n2827 585
R1869 gnd.n2050 gnd.n2049 585
R1870 gnd.n2826 gnd.n2050 585
R1871 gnd.n2824 gnd.n2823 585
R1872 gnd.n2825 gnd.n2824 585
R1873 gnd.n2822 gnd.n2052 585
R1874 gnd.n2052 gnd.n2051 585
R1875 gnd.n2821 gnd.n2820 585
R1876 gnd.n2820 gnd.n2819 585
R1877 gnd.n2058 gnd.n2057 585
R1878 gnd.n2818 gnd.n2058 585
R1879 gnd.n2816 gnd.n2815 585
R1880 gnd.n2817 gnd.n2816 585
R1881 gnd.n2814 gnd.n2060 585
R1882 gnd.n2060 gnd.n2059 585
R1883 gnd.n2813 gnd.n2812 585
R1884 gnd.n2812 gnd.n2811 585
R1885 gnd.n2066 gnd.n2065 585
R1886 gnd.n2810 gnd.n2066 585
R1887 gnd.n2808 gnd.n2807 585
R1888 gnd.n2809 gnd.n2808 585
R1889 gnd.n2806 gnd.n2068 585
R1890 gnd.n2068 gnd.n2067 585
R1891 gnd.n2805 gnd.n2804 585
R1892 gnd.n2804 gnd.n2803 585
R1893 gnd.n2074 gnd.n2073 585
R1894 gnd.n2802 gnd.n2074 585
R1895 gnd.n2800 gnd.n2799 585
R1896 gnd.n2801 gnd.n2800 585
R1897 gnd.n2798 gnd.n2076 585
R1898 gnd.n2076 gnd.n2075 585
R1899 gnd.n2797 gnd.n2796 585
R1900 gnd.n2796 gnd.n2795 585
R1901 gnd.n2082 gnd.n2081 585
R1902 gnd.n2794 gnd.n2082 585
R1903 gnd.n2792 gnd.n2791 585
R1904 gnd.n2793 gnd.n2792 585
R1905 gnd.n2790 gnd.n2084 585
R1906 gnd.n2084 gnd.n2083 585
R1907 gnd.n2789 gnd.n2788 585
R1908 gnd.n2788 gnd.n2787 585
R1909 gnd.n2090 gnd.n2089 585
R1910 gnd.n2786 gnd.n2090 585
R1911 gnd.n2784 gnd.n2783 585
R1912 gnd.n2785 gnd.n2784 585
R1913 gnd.n2782 gnd.n2092 585
R1914 gnd.n2092 gnd.n2091 585
R1915 gnd.n2781 gnd.n2780 585
R1916 gnd.n2780 gnd.n2779 585
R1917 gnd.n2098 gnd.n2097 585
R1918 gnd.n2778 gnd.n2098 585
R1919 gnd.n2776 gnd.n2775 585
R1920 gnd.n2777 gnd.n2776 585
R1921 gnd.n2774 gnd.n2100 585
R1922 gnd.n2100 gnd.n2099 585
R1923 gnd.n2773 gnd.n2772 585
R1924 gnd.n2772 gnd.n2771 585
R1925 gnd.n2106 gnd.n2105 585
R1926 gnd.n2770 gnd.n2106 585
R1927 gnd.n2768 gnd.n2767 585
R1928 gnd.n2769 gnd.n2768 585
R1929 gnd.n2766 gnd.n2108 585
R1930 gnd.n2108 gnd.n2107 585
R1931 gnd.n2765 gnd.n2764 585
R1932 gnd.n2764 gnd.n2763 585
R1933 gnd.n2114 gnd.n2113 585
R1934 gnd.n2762 gnd.n2114 585
R1935 gnd.n2760 gnd.n2759 585
R1936 gnd.n2761 gnd.n2760 585
R1937 gnd.n2758 gnd.n2116 585
R1938 gnd.n2116 gnd.n2115 585
R1939 gnd.n2757 gnd.n2756 585
R1940 gnd.n2756 gnd.n2755 585
R1941 gnd.n2122 gnd.n2121 585
R1942 gnd.n2754 gnd.n2122 585
R1943 gnd.n2752 gnd.n2751 585
R1944 gnd.n2753 gnd.n2752 585
R1945 gnd.n2750 gnd.n2124 585
R1946 gnd.n2124 gnd.n2123 585
R1947 gnd.n2749 gnd.n2748 585
R1948 gnd.n2748 gnd.n2747 585
R1949 gnd.n2130 gnd.n2129 585
R1950 gnd.n2746 gnd.n2130 585
R1951 gnd.n2744 gnd.n2743 585
R1952 gnd.n2745 gnd.n2744 585
R1953 gnd.n2742 gnd.n2132 585
R1954 gnd.n2132 gnd.n2131 585
R1955 gnd.n2741 gnd.n2740 585
R1956 gnd.n2740 gnd.n2739 585
R1957 gnd.n2138 gnd.n2137 585
R1958 gnd.n2738 gnd.n2138 585
R1959 gnd.n2736 gnd.n2735 585
R1960 gnd.n2737 gnd.n2736 585
R1961 gnd.n2734 gnd.n2140 585
R1962 gnd.n2140 gnd.n2139 585
R1963 gnd.n2733 gnd.n2732 585
R1964 gnd.n2732 gnd.n2731 585
R1965 gnd.n2146 gnd.n2145 585
R1966 gnd.n2730 gnd.n2146 585
R1967 gnd.n2728 gnd.n2727 585
R1968 gnd.n2729 gnd.n2728 585
R1969 gnd.n2726 gnd.n2148 585
R1970 gnd.n2148 gnd.n2147 585
R1971 gnd.n2725 gnd.n2724 585
R1972 gnd.n2724 gnd.n2723 585
R1973 gnd.n2154 gnd.n2153 585
R1974 gnd.n2722 gnd.n2154 585
R1975 gnd.n2720 gnd.n2719 585
R1976 gnd.n2721 gnd.n2720 585
R1977 gnd.n2718 gnd.n2156 585
R1978 gnd.n2156 gnd.n2155 585
R1979 gnd.n2717 gnd.n2716 585
R1980 gnd.n2716 gnd.n2715 585
R1981 gnd.n2162 gnd.n2161 585
R1982 gnd.n2714 gnd.n2162 585
R1983 gnd.n2712 gnd.n2711 585
R1984 gnd.n2713 gnd.n2712 585
R1985 gnd.n2710 gnd.n2164 585
R1986 gnd.n2164 gnd.n2163 585
R1987 gnd.n2709 gnd.n2708 585
R1988 gnd.n2708 gnd.n2707 585
R1989 gnd.n2170 gnd.n2169 585
R1990 gnd.n2706 gnd.n2170 585
R1991 gnd.n2704 gnd.n2703 585
R1992 gnd.n2705 gnd.n2704 585
R1993 gnd.n2702 gnd.n2172 585
R1994 gnd.n2172 gnd.n2171 585
R1995 gnd.n2701 gnd.n2700 585
R1996 gnd.n2700 gnd.n2699 585
R1997 gnd.n2178 gnd.n2177 585
R1998 gnd.n2698 gnd.n2178 585
R1999 gnd.n2696 gnd.n2695 585
R2000 gnd.n2697 gnd.n2696 585
R2001 gnd.n2694 gnd.n2180 585
R2002 gnd.n2180 gnd.n2179 585
R2003 gnd.n2693 gnd.n2692 585
R2004 gnd.n2692 gnd.n2691 585
R2005 gnd.n2186 gnd.n2185 585
R2006 gnd.n2690 gnd.n2186 585
R2007 gnd.n2688 gnd.n2687 585
R2008 gnd.n2689 gnd.n2688 585
R2009 gnd.n2686 gnd.n2188 585
R2010 gnd.n2188 gnd.n2187 585
R2011 gnd.n2685 gnd.n2684 585
R2012 gnd.n2684 gnd.n2683 585
R2013 gnd.n2194 gnd.n2193 585
R2014 gnd.n2682 gnd.n2194 585
R2015 gnd.n2680 gnd.n2679 585
R2016 gnd.n2681 gnd.n2680 585
R2017 gnd.n2678 gnd.n2196 585
R2018 gnd.n2196 gnd.n2195 585
R2019 gnd.n2677 gnd.n2676 585
R2020 gnd.n2676 gnd.n2675 585
R2021 gnd.n2202 gnd.n2201 585
R2022 gnd.n2674 gnd.n2202 585
R2023 gnd.n2672 gnd.n2671 585
R2024 gnd.n2673 gnd.n2672 585
R2025 gnd.n2670 gnd.n2204 585
R2026 gnd.n2204 gnd.n2203 585
R2027 gnd.n2669 gnd.n2668 585
R2028 gnd.n2668 gnd.n2667 585
R2029 gnd.n2210 gnd.n2209 585
R2030 gnd.n2666 gnd.n2210 585
R2031 gnd.n2664 gnd.n2663 585
R2032 gnd.n2665 gnd.n2664 585
R2033 gnd.n2662 gnd.n2212 585
R2034 gnd.n2212 gnd.n2211 585
R2035 gnd.n2661 gnd.n2660 585
R2036 gnd.n2660 gnd.n2659 585
R2037 gnd.n2218 gnd.n2217 585
R2038 gnd.n2658 gnd.n2218 585
R2039 gnd.n2656 gnd.n2655 585
R2040 gnd.n2657 gnd.n2656 585
R2041 gnd.n2654 gnd.n2220 585
R2042 gnd.n2220 gnd.n2219 585
R2043 gnd.n2653 gnd.n2652 585
R2044 gnd.n2652 gnd.n2651 585
R2045 gnd.n2226 gnd.n2225 585
R2046 gnd.n2650 gnd.n2226 585
R2047 gnd.n2648 gnd.n2647 585
R2048 gnd.n2649 gnd.n2648 585
R2049 gnd.n2646 gnd.n2228 585
R2050 gnd.n2228 gnd.n2227 585
R2051 gnd.n2645 gnd.n2644 585
R2052 gnd.n2644 gnd.n2643 585
R2053 gnd.n2234 gnd.n2233 585
R2054 gnd.n2642 gnd.n2234 585
R2055 gnd.n2640 gnd.n2639 585
R2056 gnd.n2641 gnd.n2640 585
R2057 gnd.n2638 gnd.n2236 585
R2058 gnd.n2236 gnd.n2235 585
R2059 gnd.n2637 gnd.n2636 585
R2060 gnd.n2636 gnd.n2635 585
R2061 gnd.n2242 gnd.n2241 585
R2062 gnd.n2634 gnd.n2242 585
R2063 gnd.n2632 gnd.n2631 585
R2064 gnd.n2633 gnd.n2632 585
R2065 gnd.n2630 gnd.n2244 585
R2066 gnd.n2244 gnd.n2243 585
R2067 gnd.n2629 gnd.n2628 585
R2068 gnd.n2628 gnd.n2627 585
R2069 gnd.n2250 gnd.n2249 585
R2070 gnd.n2626 gnd.n2250 585
R2071 gnd.n2624 gnd.n2623 585
R2072 gnd.n2625 gnd.n2624 585
R2073 gnd.n2622 gnd.n2252 585
R2074 gnd.n2252 gnd.n2251 585
R2075 gnd.n2621 gnd.n2620 585
R2076 gnd.n2620 gnd.n2619 585
R2077 gnd.n2258 gnd.n2257 585
R2078 gnd.n2618 gnd.n2258 585
R2079 gnd.n2616 gnd.n2615 585
R2080 gnd.n2617 gnd.n2616 585
R2081 gnd.n2614 gnd.n2260 585
R2082 gnd.n2260 gnd.n2259 585
R2083 gnd.n2613 gnd.n2612 585
R2084 gnd.n2612 gnd.n2611 585
R2085 gnd.n2266 gnd.n2265 585
R2086 gnd.n2610 gnd.n2266 585
R2087 gnd.n2608 gnd.n2607 585
R2088 gnd.n2609 gnd.n2608 585
R2089 gnd.n2438 gnd.n2437 585
R2090 gnd.n2439 gnd.n2438 585
R2091 gnd.n2442 gnd.n2441 585
R2092 gnd.n2441 gnd.n2440 585
R2093 gnd.n2443 gnd.n2429 585
R2094 gnd.n2429 gnd.n2428 585
R2095 gnd.n2445 gnd.n2444 585
R2096 gnd.n2446 gnd.n2445 585
R2097 gnd.n2427 gnd.n2426 585
R2098 gnd.n2447 gnd.n2427 585
R2099 gnd.n2450 gnd.n2449 585
R2100 gnd.n2449 gnd.n2448 585
R2101 gnd.n2451 gnd.n2421 585
R2102 gnd.n2421 gnd.n2420 585
R2103 gnd.n2453 gnd.n2452 585
R2104 gnd.n2454 gnd.n2453 585
R2105 gnd.n2419 gnd.n2418 585
R2106 gnd.n2455 gnd.n2419 585
R2107 gnd.n2458 gnd.n2457 585
R2108 gnd.n2457 gnd.n2456 585
R2109 gnd.n2459 gnd.n2413 585
R2110 gnd.n2413 gnd.n2412 585
R2111 gnd.n2461 gnd.n2460 585
R2112 gnd.n2462 gnd.n2461 585
R2113 gnd.n2411 gnd.n2410 585
R2114 gnd.n2463 gnd.n2411 585
R2115 gnd.n2466 gnd.n2465 585
R2116 gnd.n2465 gnd.n2464 585
R2117 gnd.n2467 gnd.n2405 585
R2118 gnd.n2405 gnd.n2404 585
R2119 gnd.n2469 gnd.n2468 585
R2120 gnd.n2470 gnd.n2469 585
R2121 gnd.n2403 gnd.n2402 585
R2122 gnd.n2471 gnd.n2403 585
R2123 gnd.n2474 gnd.n2473 585
R2124 gnd.n2473 gnd.n2472 585
R2125 gnd.n2475 gnd.n2397 585
R2126 gnd.n2397 gnd.n2396 585
R2127 gnd.n2477 gnd.n2476 585
R2128 gnd.n2478 gnd.n2477 585
R2129 gnd.n2395 gnd.n2394 585
R2130 gnd.n2479 gnd.n2395 585
R2131 gnd.n2482 gnd.n2481 585
R2132 gnd.n2481 gnd.n2480 585
R2133 gnd.n2483 gnd.n2389 585
R2134 gnd.n2389 gnd.n2388 585
R2135 gnd.n2485 gnd.n2484 585
R2136 gnd.n2486 gnd.n2485 585
R2137 gnd.n2387 gnd.n2386 585
R2138 gnd.n2487 gnd.n2387 585
R2139 gnd.n2490 gnd.n2489 585
R2140 gnd.n2489 gnd.n2488 585
R2141 gnd.n2491 gnd.n2381 585
R2142 gnd.n2381 gnd.n2380 585
R2143 gnd.n2493 gnd.n2492 585
R2144 gnd.n2494 gnd.n2493 585
R2145 gnd.n2379 gnd.n2378 585
R2146 gnd.n2495 gnd.n2379 585
R2147 gnd.n2498 gnd.n2497 585
R2148 gnd.n2497 gnd.n2496 585
R2149 gnd.n2499 gnd.n2373 585
R2150 gnd.n2373 gnd.n2372 585
R2151 gnd.n2501 gnd.n2500 585
R2152 gnd.n2502 gnd.n2501 585
R2153 gnd.n2371 gnd.n2370 585
R2154 gnd.n2503 gnd.n2371 585
R2155 gnd.n2506 gnd.n2505 585
R2156 gnd.n2505 gnd.n2504 585
R2157 gnd.n2507 gnd.n2365 585
R2158 gnd.n2365 gnd.n2364 585
R2159 gnd.n2509 gnd.n2508 585
R2160 gnd.n2510 gnd.n2509 585
R2161 gnd.n2363 gnd.n2362 585
R2162 gnd.n2511 gnd.n2363 585
R2163 gnd.n2514 gnd.n2513 585
R2164 gnd.n2513 gnd.n2512 585
R2165 gnd.n2515 gnd.n2357 585
R2166 gnd.n2357 gnd.n2356 585
R2167 gnd.n2517 gnd.n2516 585
R2168 gnd.n2518 gnd.n2517 585
R2169 gnd.n2355 gnd.n2354 585
R2170 gnd.n2519 gnd.n2355 585
R2171 gnd.n2522 gnd.n2521 585
R2172 gnd.n2521 gnd.n2520 585
R2173 gnd.n2523 gnd.n2349 585
R2174 gnd.n2349 gnd.n2348 585
R2175 gnd.n2525 gnd.n2524 585
R2176 gnd.n2526 gnd.n2525 585
R2177 gnd.n2347 gnd.n2346 585
R2178 gnd.n2527 gnd.n2347 585
R2179 gnd.n2530 gnd.n2529 585
R2180 gnd.n2529 gnd.n2528 585
R2181 gnd.n2531 gnd.n2341 585
R2182 gnd.n2341 gnd.n2340 585
R2183 gnd.n2533 gnd.n2532 585
R2184 gnd.n2534 gnd.n2533 585
R2185 gnd.n2339 gnd.n2338 585
R2186 gnd.n2535 gnd.n2339 585
R2187 gnd.n2538 gnd.n2537 585
R2188 gnd.n2537 gnd.n2536 585
R2189 gnd.n2539 gnd.n2333 585
R2190 gnd.n2333 gnd.n2332 585
R2191 gnd.n2541 gnd.n2540 585
R2192 gnd.n2542 gnd.n2541 585
R2193 gnd.n2331 gnd.n2330 585
R2194 gnd.n2543 gnd.n2331 585
R2195 gnd.n2546 gnd.n2545 585
R2196 gnd.n2545 gnd.n2544 585
R2197 gnd.n2547 gnd.n2325 585
R2198 gnd.n2325 gnd.n2324 585
R2199 gnd.n2549 gnd.n2548 585
R2200 gnd.n2550 gnd.n2549 585
R2201 gnd.n2323 gnd.n2322 585
R2202 gnd.n2551 gnd.n2323 585
R2203 gnd.n2554 gnd.n2553 585
R2204 gnd.n2553 gnd.n2552 585
R2205 gnd.n2555 gnd.n2317 585
R2206 gnd.n2317 gnd.n2316 585
R2207 gnd.n2557 gnd.n2556 585
R2208 gnd.n2558 gnd.n2557 585
R2209 gnd.n2315 gnd.n2314 585
R2210 gnd.n2559 gnd.n2315 585
R2211 gnd.n2562 gnd.n2561 585
R2212 gnd.n2561 gnd.n2560 585
R2213 gnd.n2563 gnd.n2309 585
R2214 gnd.n2309 gnd.n2308 585
R2215 gnd.n2565 gnd.n2564 585
R2216 gnd.n2566 gnd.n2565 585
R2217 gnd.n2307 gnd.n2306 585
R2218 gnd.n2567 gnd.n2307 585
R2219 gnd.n2570 gnd.n2569 585
R2220 gnd.n2569 gnd.n2568 585
R2221 gnd.n2571 gnd.n2301 585
R2222 gnd.n2301 gnd.n2300 585
R2223 gnd.n2573 gnd.n2572 585
R2224 gnd.n2574 gnd.n2573 585
R2225 gnd.n2299 gnd.n2298 585
R2226 gnd.n2575 gnd.n2299 585
R2227 gnd.n2578 gnd.n2577 585
R2228 gnd.n2577 gnd.n2576 585
R2229 gnd.n2579 gnd.n2293 585
R2230 gnd.n2293 gnd.n2292 585
R2231 gnd.n2581 gnd.n2580 585
R2232 gnd.n2582 gnd.n2581 585
R2233 gnd.n2291 gnd.n2290 585
R2234 gnd.n2583 gnd.n2291 585
R2235 gnd.n2586 gnd.n2585 585
R2236 gnd.n2585 gnd.n2584 585
R2237 gnd.n2587 gnd.n2285 585
R2238 gnd.n2285 gnd.n2284 585
R2239 gnd.n2589 gnd.n2588 585
R2240 gnd.n2590 gnd.n2589 585
R2241 gnd.n2283 gnd.n2282 585
R2242 gnd.n2591 gnd.n2283 585
R2243 gnd.n2594 gnd.n2593 585
R2244 gnd.n2593 gnd.n2592 585
R2245 gnd.n2595 gnd.n2277 585
R2246 gnd.n2277 gnd.n2276 585
R2247 gnd.n2597 gnd.n2596 585
R2248 gnd.n2598 gnd.n2597 585
R2249 gnd.n2274 gnd.n2273 585
R2250 gnd.n2599 gnd.n2274 585
R2251 gnd.n2602 gnd.n2601 585
R2252 gnd.n2601 gnd.n2600 585
R2253 gnd.n2603 gnd.n2271 585
R2254 gnd.n2275 gnd.n2271 585
R2255 gnd.n2604 gnd.n2268 585
R2256 gnd.n2268 gnd.n2267 585
R2257 gnd.n1592 gnd.n1246 585
R2258 gnd.n6152 gnd.n1246 585
R2259 gnd.n5602 gnd.n5601 585
R2260 gnd.n5603 gnd.n5602 585
R2261 gnd.n5600 gnd.n1596 585
R2262 gnd.n5563 gnd.n1596 585
R2263 gnd.n1604 gnd.n1597 585
R2264 gnd.n5595 gnd.n1604 585
R2265 gnd.n5582 gnd.n1616 585
R2266 gnd.n5561 gnd.n1616 585
R2267 gnd.n5584 gnd.n5583 585
R2268 gnd.n5585 gnd.n5584 585
R2269 gnd.n1617 gnd.n1615 585
R2270 gnd.n5577 gnd.n1615 585
R2271 gnd.n5540 gnd.n5539 585
R2272 gnd.n5539 gnd.n5538 585
R2273 gnd.n5541 gnd.n1630 585
R2274 gnd.n5555 gnd.n1630 585
R2275 gnd.n5542 gnd.n1642 585
R2276 gnd.n1680 gnd.n1642 585
R2277 gnd.n5544 gnd.n5543 585
R2278 gnd.n5545 gnd.n5544 585
R2279 gnd.n1643 gnd.n1641 585
R2280 gnd.n5468 gnd.n1641 585
R2281 gnd.n5473 gnd.n1662 585
R2282 gnd.n5485 gnd.n1662 585
R2283 gnd.n5474 gnd.n1672 585
R2284 gnd.n1672 gnd.n1658 585
R2285 gnd.n5476 gnd.n5475 585
R2286 gnd.n5477 gnd.n5476 585
R2287 gnd.n1673 gnd.n1671 585
R2288 gnd.n1714 gnd.n1671 585
R2289 gnd.n5437 gnd.n5436 585
R2290 gnd.n5436 gnd.n5435 585
R2291 gnd.n5438 gnd.n1695 585
R2292 gnd.n5452 gnd.n1695 585
R2293 gnd.n5439 gnd.n1707 585
R2294 gnd.n5423 gnd.n1707 585
R2295 gnd.n5441 gnd.n5440 585
R2296 gnd.n5442 gnd.n5441 585
R2297 gnd.n1708 gnd.n1706 585
R2298 gnd.n5411 gnd.n1706 585
R2299 gnd.n5387 gnd.n5386 585
R2300 gnd.n5386 gnd.n5385 585
R2301 gnd.n5388 gnd.n1733 585
R2302 gnd.n5402 gnd.n1733 585
R2303 gnd.n5389 gnd.n1745 585
R2304 gnd.n5373 gnd.n1745 585
R2305 gnd.n5391 gnd.n5390 585
R2306 gnd.n5392 gnd.n5391 585
R2307 gnd.n1746 gnd.n1744 585
R2308 gnd.n5366 gnd.n1744 585
R2309 gnd.n3607 gnd.n3606 585
R2310 gnd.n3606 gnd.n3605 585
R2311 gnd.n3595 gnd.n1769 585
R2312 gnd.n5357 gnd.n1769 585
R2313 gnd.n1804 gnd.n1803 585
R2314 gnd.n1804 gnd.n1766 585
R2315 gnd.n5329 gnd.n5328 585
R2316 gnd.n5328 gnd.n5327 585
R2317 gnd.n5330 gnd.n1799 585
R2318 gnd.n1805 gnd.n1799 585
R2319 gnd.n5332 gnd.n5331 585
R2320 gnd.n5333 gnd.n5332 585
R2321 gnd.n1792 gnd.n1791 585
R2322 gnd.n1795 gnd.n1792 585
R2323 gnd.n5343 gnd.n5342 585
R2324 gnd.n5342 gnd.n5341 585
R2325 gnd.n5344 gnd.n1786 585
R2326 gnd.n1786 gnd.n1784 585
R2327 gnd.n5346 gnd.n5345 585
R2328 gnd.n5347 gnd.n5346 585
R2329 gnd.n1787 gnd.n1785 585
R2330 gnd.n3548 gnd.n1785 585
R2331 gnd.n3628 gnd.n3627 585
R2332 gnd.n3629 gnd.n3628 585
R2333 gnd.n3393 gnd.n3392 585
R2334 gnd.n3630 gnd.n3393 585
R2335 gnd.n3639 gnd.n3638 585
R2336 gnd.n3638 gnd.n3637 585
R2337 gnd.n3640 gnd.n3388 585
R2338 gnd.n3388 gnd.n3387 585
R2339 gnd.n3642 gnd.n3641 585
R2340 gnd.n3643 gnd.n3642 585
R2341 gnd.n3374 gnd.n3373 585
R2342 gnd.n3377 gnd.n3374 585
R2343 gnd.n3651 gnd.n3650 585
R2344 gnd.n3650 gnd.n3649 585
R2345 gnd.n3652 gnd.n3369 585
R2346 gnd.n3369 gnd.n3368 585
R2347 gnd.n3654 gnd.n3653 585
R2348 gnd.n3655 gnd.n3654 585
R2349 gnd.n3355 gnd.n3354 585
R2350 gnd.n3365 gnd.n3355 585
R2351 gnd.n3663 gnd.n3662 585
R2352 gnd.n3662 gnd.n3661 585
R2353 gnd.n3664 gnd.n3350 585
R2354 gnd.n3350 gnd.n3349 585
R2355 gnd.n3666 gnd.n3665 585
R2356 gnd.n3667 gnd.n3666 585
R2357 gnd.n3336 gnd.n3335 585
R2358 gnd.n3339 gnd.n3336 585
R2359 gnd.n3675 gnd.n3674 585
R2360 gnd.n3674 gnd.n3673 585
R2361 gnd.n3676 gnd.n3331 585
R2362 gnd.n3331 gnd.n3330 585
R2363 gnd.n3678 gnd.n3677 585
R2364 gnd.n3679 gnd.n3678 585
R2365 gnd.n3317 gnd.n3316 585
R2366 gnd.n3327 gnd.n3317 585
R2367 gnd.n3687 gnd.n3686 585
R2368 gnd.n3686 gnd.n3685 585
R2369 gnd.n3688 gnd.n3312 585
R2370 gnd.n3312 gnd.n3311 585
R2371 gnd.n3690 gnd.n3689 585
R2372 gnd.n3691 gnd.n3690 585
R2373 gnd.n3298 gnd.n3297 585
R2374 gnd.n3301 gnd.n3298 585
R2375 gnd.n3699 gnd.n3698 585
R2376 gnd.n3698 gnd.n3697 585
R2377 gnd.n3700 gnd.n3291 585
R2378 gnd.n3291 gnd.n3289 585
R2379 gnd.n3702 gnd.n3701 585
R2380 gnd.n3703 gnd.n3702 585
R2381 gnd.n3293 gnd.n3290 585
R2382 gnd.n3290 gnd.n3286 585
R2383 gnd.n3292 gnd.n3277 585
R2384 gnd.n3709 gnd.n3277 585
R2385 gnd.n3429 gnd.n3271 585
R2386 gnd.n3429 gnd.n3202 585
R2387 gnd.n3431 gnd.n3430 585
R2388 gnd.n3433 gnd.n3432 585
R2389 gnd.n3435 gnd.n3434 585
R2390 gnd.n3439 gnd.n3427 585
R2391 gnd.n3441 gnd.n3440 585
R2392 gnd.n3443 gnd.n3442 585
R2393 gnd.n3445 gnd.n3444 585
R2394 gnd.n3449 gnd.n3425 585
R2395 gnd.n3451 gnd.n3450 585
R2396 gnd.n3453 gnd.n3452 585
R2397 gnd.n3455 gnd.n3454 585
R2398 gnd.n3459 gnd.n3423 585
R2399 gnd.n3461 gnd.n3460 585
R2400 gnd.n3463 gnd.n3462 585
R2401 gnd.n3465 gnd.n3464 585
R2402 gnd.n3420 gnd.n3419 585
R2403 gnd.n3469 gnd.n3421 585
R2404 gnd.n3470 gnd.n3416 585
R2405 gnd.n3471 gnd.n3201 585
R2406 gnd.n3833 gnd.n3201 585
R2407 gnd.n6155 gnd.n6154 585
R2408 gnd.n5679 gnd.n1239 585
R2409 gnd.n5681 gnd.n5680 585
R2410 gnd.n5677 gnd.n5665 585
R2411 gnd.n5688 gnd.n5664 585
R2412 gnd.n5689 gnd.n5662 585
R2413 gnd.n5661 gnd.n5654 585
R2414 gnd.n5696 gnd.n5653 585
R2415 gnd.n5697 gnd.n5652 585
R2416 gnd.n5650 gnd.n5642 585
R2417 gnd.n5704 gnd.n5641 585
R2418 gnd.n5705 gnd.n5639 585
R2419 gnd.n5638 gnd.n5631 585
R2420 gnd.n5712 gnd.n5630 585
R2421 gnd.n5713 gnd.n5629 585
R2422 gnd.n5627 gnd.n5619 585
R2423 gnd.n5720 gnd.n5618 585
R2424 gnd.n5721 gnd.n5616 585
R2425 gnd.n5615 gnd.n5614 585
R2426 gnd.n5615 gnd.n1253 585
R2427 gnd.n6153 gnd.n1242 585
R2428 gnd.n6153 gnd.n6152 585
R2429 gnd.n5565 gnd.n1241 585
R2430 gnd.n5603 gnd.n1241 585
R2431 gnd.n5569 gnd.n5564 585
R2432 gnd.n5564 gnd.n5563 585
R2433 gnd.n5570 gnd.n1602 585
R2434 gnd.n5595 gnd.n1602 585
R2435 gnd.n5571 gnd.n5562 585
R2436 gnd.n5562 gnd.n5561 585
R2437 gnd.n1623 gnd.n1613 585
R2438 gnd.n5585 gnd.n1613 585
R2439 gnd.n5576 gnd.n5575 585
R2440 gnd.n5577 gnd.n5576 585
R2441 gnd.n1622 gnd.n1621 585
R2442 gnd.n5538 gnd.n1621 585
R2443 gnd.n5557 gnd.n5556 585
R2444 gnd.n5556 gnd.n5555 585
R2445 gnd.n1626 gnd.n1625 585
R2446 gnd.n1680 gnd.n1626 585
R2447 gnd.n1685 gnd.n1639 585
R2448 gnd.n5545 gnd.n1639 585
R2449 gnd.n5467 gnd.n5466 585
R2450 gnd.n5468 gnd.n5467 585
R2451 gnd.n1684 gnd.n1660 585
R2452 gnd.n5485 gnd.n1660 585
R2453 gnd.n5461 gnd.n5460 585
R2454 gnd.n5460 gnd.n1658 585
R2455 gnd.n5459 gnd.n1669 585
R2456 gnd.n5477 gnd.n1669 585
R2457 gnd.n5458 gnd.n1688 585
R2458 gnd.n1714 gnd.n1688 585
R2459 gnd.n1692 gnd.n1687 585
R2460 gnd.n5435 gnd.n1692 585
R2461 gnd.n5454 gnd.n5453 585
R2462 gnd.n5453 gnd.n5452 585
R2463 gnd.n1691 gnd.n1690 585
R2464 gnd.n5423 gnd.n1691 585
R2465 gnd.n1727 gnd.n1704 585
R2466 gnd.n5442 gnd.n1704 585
R2467 gnd.n5410 gnd.n5409 585
R2468 gnd.n5411 gnd.n5410 585
R2469 gnd.n1726 gnd.n1725 585
R2470 gnd.n5385 gnd.n1725 585
R2471 gnd.n5404 gnd.n5403 585
R2472 gnd.n5403 gnd.n5402 585
R2473 gnd.n1730 gnd.n1729 585
R2474 gnd.n5373 gnd.n1730 585
R2475 gnd.n1762 gnd.n1742 585
R2476 gnd.n5392 gnd.n1742 585
R2477 gnd.n5365 gnd.n5364 585
R2478 gnd.n5366 gnd.n5365 585
R2479 gnd.n1761 gnd.n1760 585
R2480 gnd.n3605 gnd.n1760 585
R2481 gnd.n5359 gnd.n5358 585
R2482 gnd.n5358 gnd.n5357 585
R2483 gnd.n1765 gnd.n1764 585
R2484 gnd.n1766 gnd.n1765 585
R2485 gnd.n3536 gnd.n1807 585
R2486 gnd.n5327 gnd.n1807 585
R2487 gnd.n3537 gnd.n3535 585
R2488 gnd.n3535 gnd.n1805 585
R2489 gnd.n3533 gnd.n1798 585
R2490 gnd.n5333 gnd.n1798 585
R2491 gnd.n3541 gnd.n3532 585
R2492 gnd.n3532 gnd.n1795 585
R2493 gnd.n3542 gnd.n1794 585
R2494 gnd.n5341 gnd.n1794 585
R2495 gnd.n3544 gnd.n3543 585
R2496 gnd.n3543 gnd.n1784 585
R2497 gnd.n3545 gnd.n1783 585
R2498 gnd.n5347 gnd.n1783 585
R2499 gnd.n3547 gnd.n3546 585
R2500 gnd.n3548 gnd.n3547 585
R2501 gnd.n3401 gnd.n3400 585
R2502 gnd.n3629 gnd.n3400 585
R2503 gnd.n3525 gnd.n3398 585
R2504 gnd.n3630 gnd.n3398 585
R2505 gnd.n3524 gnd.n3395 585
R2506 gnd.n3637 gnd.n3395 585
R2507 gnd.n3523 gnd.n3522 585
R2508 gnd.n3522 gnd.n3387 585
R2509 gnd.n3403 gnd.n3386 585
R2510 gnd.n3643 gnd.n3386 585
R2511 gnd.n3518 gnd.n3517 585
R2512 gnd.n3517 gnd.n3377 585
R2513 gnd.n3516 gnd.n3376 585
R2514 gnd.n3649 gnd.n3376 585
R2515 gnd.n3515 gnd.n3514 585
R2516 gnd.n3514 gnd.n3368 585
R2517 gnd.n3405 gnd.n3367 585
R2518 gnd.n3655 gnd.n3367 585
R2519 gnd.n3510 gnd.n3509 585
R2520 gnd.n3509 gnd.n3365 585
R2521 gnd.n3508 gnd.n3357 585
R2522 gnd.n3661 gnd.n3357 585
R2523 gnd.n3507 gnd.n3506 585
R2524 gnd.n3506 gnd.n3349 585
R2525 gnd.n3407 gnd.n3348 585
R2526 gnd.n3667 gnd.n3348 585
R2527 gnd.n3502 gnd.n3501 585
R2528 gnd.n3501 gnd.n3339 585
R2529 gnd.n3500 gnd.n3338 585
R2530 gnd.n3673 gnd.n3338 585
R2531 gnd.n3499 gnd.n3498 585
R2532 gnd.n3498 gnd.n3330 585
R2533 gnd.n3409 gnd.n3329 585
R2534 gnd.n3679 gnd.n3329 585
R2535 gnd.n3494 gnd.n3493 585
R2536 gnd.n3493 gnd.n3327 585
R2537 gnd.n3492 gnd.n3319 585
R2538 gnd.n3685 gnd.n3319 585
R2539 gnd.n3491 gnd.n3490 585
R2540 gnd.n3490 gnd.n3311 585
R2541 gnd.n3411 gnd.n3310 585
R2542 gnd.n3691 gnd.n3310 585
R2543 gnd.n3486 gnd.n3485 585
R2544 gnd.n3485 gnd.n3301 585
R2545 gnd.n3484 gnd.n3300 585
R2546 gnd.n3697 gnd.n3300 585
R2547 gnd.n3483 gnd.n3482 585
R2548 gnd.n3482 gnd.n3289 585
R2549 gnd.n3413 gnd.n3288 585
R2550 gnd.n3703 gnd.n3288 585
R2551 gnd.n3478 gnd.n3477 585
R2552 gnd.n3477 gnd.n3286 585
R2553 gnd.n3476 gnd.n3276 585
R2554 gnd.n3709 gnd.n3276 585
R2555 gnd.n3475 gnd.n3474 585
R2556 gnd.n3474 gnd.n3202 585
R2557 gnd.n5220 gnd.n5219 585
R2558 gnd.n5221 gnd.n5220 585
R2559 gnd.n3895 gnd.n3894 585
R2560 gnd.n3901 gnd.n3894 585
R2561 gnd.n5195 gnd.n3913 585
R2562 gnd.n3913 gnd.n3900 585
R2563 gnd.n5197 gnd.n5196 585
R2564 gnd.n5198 gnd.n5197 585
R2565 gnd.n3914 gnd.n3912 585
R2566 gnd.n3912 gnd.n3908 585
R2567 gnd.n4929 gnd.n4928 585
R2568 gnd.n4928 gnd.n4927 585
R2569 gnd.n3919 gnd.n3918 585
R2570 gnd.n4898 gnd.n3919 585
R2571 gnd.n4918 gnd.n4917 585
R2572 gnd.n4917 gnd.n4916 585
R2573 gnd.n3926 gnd.n3925 585
R2574 gnd.n4904 gnd.n3926 585
R2575 gnd.n4874 gnd.n3946 585
R2576 gnd.n3946 gnd.n3945 585
R2577 gnd.n4876 gnd.n4875 585
R2578 gnd.n4877 gnd.n4876 585
R2579 gnd.n3947 gnd.n3944 585
R2580 gnd.n3955 gnd.n3944 585
R2581 gnd.n4852 gnd.n3967 585
R2582 gnd.n3967 gnd.n3954 585
R2583 gnd.n4854 gnd.n4853 585
R2584 gnd.n4855 gnd.n4854 585
R2585 gnd.n3968 gnd.n3966 585
R2586 gnd.n3966 gnd.n3962 585
R2587 gnd.n4840 gnd.n4839 585
R2588 gnd.n4839 gnd.n4838 585
R2589 gnd.n3973 gnd.n3972 585
R2590 gnd.n3983 gnd.n3973 585
R2591 gnd.n4829 gnd.n4828 585
R2592 gnd.n4828 gnd.n4827 585
R2593 gnd.n3980 gnd.n3979 585
R2594 gnd.n4815 gnd.n3980 585
R2595 gnd.n4789 gnd.n4001 585
R2596 gnd.n4001 gnd.n3990 585
R2597 gnd.n4791 gnd.n4790 585
R2598 gnd.n4792 gnd.n4791 585
R2599 gnd.n4002 gnd.n4000 585
R2600 gnd.n4010 gnd.n4000 585
R2601 gnd.n4767 gnd.n4022 585
R2602 gnd.n4022 gnd.n4009 585
R2603 gnd.n4769 gnd.n4768 585
R2604 gnd.n4770 gnd.n4769 585
R2605 gnd.n4023 gnd.n4021 585
R2606 gnd.n4021 gnd.n4017 585
R2607 gnd.n4755 gnd.n4754 585
R2608 gnd.n4754 gnd.n4753 585
R2609 gnd.n4028 gnd.n4027 585
R2610 gnd.n4037 gnd.n4028 585
R2611 gnd.n4744 gnd.n4743 585
R2612 gnd.n4743 gnd.n4742 585
R2613 gnd.n4035 gnd.n4034 585
R2614 gnd.n4730 gnd.n4035 585
R2615 gnd.n4168 gnd.n4167 585
R2616 gnd.n4168 gnd.n4044 585
R2617 gnd.n4687 gnd.n4686 585
R2618 gnd.n4686 gnd.n4685 585
R2619 gnd.n4688 gnd.n4162 585
R2620 gnd.n4173 gnd.n4162 585
R2621 gnd.n4690 gnd.n4689 585
R2622 gnd.n4691 gnd.n4690 585
R2623 gnd.n4163 gnd.n4161 585
R2624 gnd.n4186 gnd.n4161 585
R2625 gnd.n4146 gnd.n4145 585
R2626 gnd.n4149 gnd.n4146 585
R2627 gnd.n4701 gnd.n4700 585
R2628 gnd.n4700 gnd.n4699 585
R2629 gnd.n4702 gnd.n4140 585
R2630 gnd.n4661 gnd.n4140 585
R2631 gnd.n4704 gnd.n4703 585
R2632 gnd.n4705 gnd.n4704 585
R2633 gnd.n4141 gnd.n4139 585
R2634 gnd.n4200 gnd.n4139 585
R2635 gnd.n4653 gnd.n4652 585
R2636 gnd.n4652 gnd.n4651 585
R2637 gnd.n4197 gnd.n4196 585
R2638 gnd.n4635 gnd.n4197 585
R2639 gnd.n4622 gnd.n4216 585
R2640 gnd.n4216 gnd.n4215 585
R2641 gnd.n4624 gnd.n4623 585
R2642 gnd.n4625 gnd.n4624 585
R2643 gnd.n4217 gnd.n4214 585
R2644 gnd.n4223 gnd.n4214 585
R2645 gnd.n4603 gnd.n4602 585
R2646 gnd.n4604 gnd.n4603 585
R2647 gnd.n4234 gnd.n4233 585
R2648 gnd.n4233 gnd.n4229 585
R2649 gnd.n4593 gnd.n4592 585
R2650 gnd.n4594 gnd.n4593 585
R2651 gnd.n4244 gnd.n4243 585
R2652 gnd.n4249 gnd.n4243 585
R2653 gnd.n4571 gnd.n4262 585
R2654 gnd.n4262 gnd.n4248 585
R2655 gnd.n4573 gnd.n4572 585
R2656 gnd.n4574 gnd.n4573 585
R2657 gnd.n4263 gnd.n4261 585
R2658 gnd.n4261 gnd.n4257 585
R2659 gnd.n4562 gnd.n4561 585
R2660 gnd.n4563 gnd.n4562 585
R2661 gnd.n4270 gnd.n4269 585
R2662 gnd.n4274 gnd.n4269 585
R2663 gnd.n4539 gnd.n4291 585
R2664 gnd.n4291 gnd.n4273 585
R2665 gnd.n4541 gnd.n4540 585
R2666 gnd.n4542 gnd.n4541 585
R2667 gnd.n4292 gnd.n4290 585
R2668 gnd.n4290 gnd.n4281 585
R2669 gnd.n4534 gnd.n4533 585
R2670 gnd.n4533 gnd.n4532 585
R2671 gnd.n4339 gnd.n4338 585
R2672 gnd.n4340 gnd.n4339 585
R2673 gnd.n4493 gnd.n4492 585
R2674 gnd.n4494 gnd.n4493 585
R2675 gnd.n4349 gnd.n4348 585
R2676 gnd.n4348 gnd.n4347 585
R2677 gnd.n4488 gnd.n4487 585
R2678 gnd.n4487 gnd.n4486 585
R2679 gnd.n4352 gnd.n4351 585
R2680 gnd.n4353 gnd.n4352 585
R2681 gnd.n4477 gnd.n4476 585
R2682 gnd.n4478 gnd.n4477 585
R2683 gnd.n4360 gnd.n4359 585
R2684 gnd.n4469 gnd.n4359 585
R2685 gnd.n4472 gnd.n4471 585
R2686 gnd.n4471 gnd.n4470 585
R2687 gnd.n4363 gnd.n4362 585
R2688 gnd.n4364 gnd.n4363 585
R2689 gnd.n4458 gnd.n4457 585
R2690 gnd.n4456 gnd.n4382 585
R2691 gnd.n4455 gnd.n4381 585
R2692 gnd.n4460 gnd.n4381 585
R2693 gnd.n4454 gnd.n4453 585
R2694 gnd.n4452 gnd.n4451 585
R2695 gnd.n4450 gnd.n4449 585
R2696 gnd.n4448 gnd.n4447 585
R2697 gnd.n4446 gnd.n4445 585
R2698 gnd.n4444 gnd.n4443 585
R2699 gnd.n4442 gnd.n4441 585
R2700 gnd.n4440 gnd.n4439 585
R2701 gnd.n4438 gnd.n4437 585
R2702 gnd.n4436 gnd.n4435 585
R2703 gnd.n4434 gnd.n4433 585
R2704 gnd.n4432 gnd.n4431 585
R2705 gnd.n4430 gnd.n4429 585
R2706 gnd.n4428 gnd.n4427 585
R2707 gnd.n4426 gnd.n4425 585
R2708 gnd.n4424 gnd.n4423 585
R2709 gnd.n4422 gnd.n4421 585
R2710 gnd.n4420 gnd.n4419 585
R2711 gnd.n4418 gnd.n4417 585
R2712 gnd.n4416 gnd.n4415 585
R2713 gnd.n4414 gnd.n4413 585
R2714 gnd.n4412 gnd.n4411 585
R2715 gnd.n4369 gnd.n4368 585
R2716 gnd.n4463 gnd.n4462 585
R2717 gnd.n5224 gnd.n5223 585
R2718 gnd.n5226 gnd.n5225 585
R2719 gnd.n5228 gnd.n5227 585
R2720 gnd.n5230 gnd.n5229 585
R2721 gnd.n5232 gnd.n5231 585
R2722 gnd.n5234 gnd.n5233 585
R2723 gnd.n5236 gnd.n5235 585
R2724 gnd.n5238 gnd.n5237 585
R2725 gnd.n5240 gnd.n5239 585
R2726 gnd.n5242 gnd.n5241 585
R2727 gnd.n5244 gnd.n5243 585
R2728 gnd.n5246 gnd.n5245 585
R2729 gnd.n5248 gnd.n5247 585
R2730 gnd.n5250 gnd.n5249 585
R2731 gnd.n5252 gnd.n5251 585
R2732 gnd.n5254 gnd.n5253 585
R2733 gnd.n5256 gnd.n5255 585
R2734 gnd.n5258 gnd.n5257 585
R2735 gnd.n5260 gnd.n5259 585
R2736 gnd.n5262 gnd.n5261 585
R2737 gnd.n5264 gnd.n5263 585
R2738 gnd.n5266 gnd.n5265 585
R2739 gnd.n5268 gnd.n5267 585
R2740 gnd.n5270 gnd.n5269 585
R2741 gnd.n5272 gnd.n5271 585
R2742 gnd.n5273 gnd.n3862 585
R2743 gnd.n5274 gnd.n3150 585
R2744 gnd.n5312 gnd.n3150 585
R2745 gnd.n5222 gnd.n3892 585
R2746 gnd.n5222 gnd.n5221 585
R2747 gnd.n4891 gnd.n3891 585
R2748 gnd.n3901 gnd.n3891 585
R2749 gnd.n4893 gnd.n4892 585
R2750 gnd.n4892 gnd.n3900 585
R2751 gnd.n4894 gnd.n3910 585
R2752 gnd.n5198 gnd.n3910 585
R2753 gnd.n4896 gnd.n4895 585
R2754 gnd.n4895 gnd.n3908 585
R2755 gnd.n4897 gnd.n3921 585
R2756 gnd.n4927 gnd.n3921 585
R2757 gnd.n4900 gnd.n4899 585
R2758 gnd.n4899 gnd.n4898 585
R2759 gnd.n4901 gnd.n3928 585
R2760 gnd.n4916 gnd.n3928 585
R2761 gnd.n4903 gnd.n4902 585
R2762 gnd.n4904 gnd.n4903 585
R2763 gnd.n3938 gnd.n3937 585
R2764 gnd.n3945 gnd.n3937 585
R2765 gnd.n4879 gnd.n4878 585
R2766 gnd.n4878 gnd.n4877 585
R2767 gnd.n3941 gnd.n3940 585
R2768 gnd.n3955 gnd.n3941 585
R2769 gnd.n4805 gnd.n4804 585
R2770 gnd.n4804 gnd.n3954 585
R2771 gnd.n4806 gnd.n3964 585
R2772 gnd.n4855 gnd.n3964 585
R2773 gnd.n4808 gnd.n4807 585
R2774 gnd.n4807 gnd.n3962 585
R2775 gnd.n4809 gnd.n3975 585
R2776 gnd.n4838 gnd.n3975 585
R2777 gnd.n4811 gnd.n4810 585
R2778 gnd.n4810 gnd.n3983 585
R2779 gnd.n4812 gnd.n3982 585
R2780 gnd.n4827 gnd.n3982 585
R2781 gnd.n4814 gnd.n4813 585
R2782 gnd.n4815 gnd.n4814 585
R2783 gnd.n3994 gnd.n3993 585
R2784 gnd.n3993 gnd.n3990 585
R2785 gnd.n4794 gnd.n4793 585
R2786 gnd.n4793 gnd.n4792 585
R2787 gnd.n3997 gnd.n3996 585
R2788 gnd.n4010 gnd.n3997 585
R2789 gnd.n4718 gnd.n4717 585
R2790 gnd.n4717 gnd.n4009 585
R2791 gnd.n4719 gnd.n4019 585
R2792 gnd.n4770 gnd.n4019 585
R2793 gnd.n4721 gnd.n4720 585
R2794 gnd.n4720 gnd.n4017 585
R2795 gnd.n4722 gnd.n4030 585
R2796 gnd.n4753 gnd.n4030 585
R2797 gnd.n4724 gnd.n4723 585
R2798 gnd.n4723 gnd.n4037 585
R2799 gnd.n4725 gnd.n4036 585
R2800 gnd.n4742 gnd.n4036 585
R2801 gnd.n4727 gnd.n4726 585
R2802 gnd.n4730 gnd.n4727 585
R2803 gnd.n4047 gnd.n4046 585
R2804 gnd.n4046 gnd.n4044 585
R2805 gnd.n4170 gnd.n4169 585
R2806 gnd.n4685 gnd.n4169 585
R2807 gnd.n4172 gnd.n4171 585
R2808 gnd.n4173 gnd.n4172 585
R2809 gnd.n4183 gnd.n4159 585
R2810 gnd.n4691 gnd.n4159 585
R2811 gnd.n4185 gnd.n4184 585
R2812 gnd.n4186 gnd.n4185 585
R2813 gnd.n4182 gnd.n4181 585
R2814 gnd.n4182 gnd.n4149 585
R2815 gnd.n4180 gnd.n4147 585
R2816 gnd.n4699 gnd.n4147 585
R2817 gnd.n4136 gnd.n4134 585
R2818 gnd.n4661 gnd.n4136 585
R2819 gnd.n4707 gnd.n4706 585
R2820 gnd.n4706 gnd.n4705 585
R2821 gnd.n4135 gnd.n4133 585
R2822 gnd.n4200 gnd.n4135 585
R2823 gnd.n4632 gnd.n4199 585
R2824 gnd.n4651 gnd.n4199 585
R2825 gnd.n4634 gnd.n4633 585
R2826 gnd.n4635 gnd.n4634 585
R2827 gnd.n4209 gnd.n4208 585
R2828 gnd.n4215 gnd.n4208 585
R2829 gnd.n4627 gnd.n4626 585
R2830 gnd.n4626 gnd.n4625 585
R2831 gnd.n4212 gnd.n4211 585
R2832 gnd.n4223 gnd.n4212 585
R2833 gnd.n4512 gnd.n4231 585
R2834 gnd.n4604 gnd.n4231 585
R2835 gnd.n4514 gnd.n4513 585
R2836 gnd.n4513 gnd.n4229 585
R2837 gnd.n4515 gnd.n4242 585
R2838 gnd.n4594 gnd.n4242 585
R2839 gnd.n4517 gnd.n4516 585
R2840 gnd.n4517 gnd.n4249 585
R2841 gnd.n4519 gnd.n4518 585
R2842 gnd.n4518 gnd.n4248 585
R2843 gnd.n4520 gnd.n4259 585
R2844 gnd.n4574 gnd.n4259 585
R2845 gnd.n4522 gnd.n4521 585
R2846 gnd.n4521 gnd.n4257 585
R2847 gnd.n4523 gnd.n4268 585
R2848 gnd.n4563 gnd.n4268 585
R2849 gnd.n4525 gnd.n4524 585
R2850 gnd.n4525 gnd.n4274 585
R2851 gnd.n4527 gnd.n4526 585
R2852 gnd.n4526 gnd.n4273 585
R2853 gnd.n4528 gnd.n4289 585
R2854 gnd.n4542 gnd.n4289 585
R2855 gnd.n4529 gnd.n4342 585
R2856 gnd.n4342 gnd.n4281 585
R2857 gnd.n4531 gnd.n4530 585
R2858 gnd.n4532 gnd.n4531 585
R2859 gnd.n4343 gnd.n4341 585
R2860 gnd.n4341 gnd.n4340 585
R2861 gnd.n4496 gnd.n4495 585
R2862 gnd.n4495 gnd.n4494 585
R2863 gnd.n4346 gnd.n4345 585
R2864 gnd.n4347 gnd.n4346 585
R2865 gnd.n4485 gnd.n4484 585
R2866 gnd.n4486 gnd.n4485 585
R2867 gnd.n4355 gnd.n4354 585
R2868 gnd.n4354 gnd.n4353 585
R2869 gnd.n4480 gnd.n4479 585
R2870 gnd.n4479 gnd.n4478 585
R2871 gnd.n4358 gnd.n4357 585
R2872 gnd.n4469 gnd.n4358 585
R2873 gnd.n4468 gnd.n4467 585
R2874 gnd.n4470 gnd.n4468 585
R2875 gnd.n4366 gnd.n4365 585
R2876 gnd.n4365 gnd.n4364 585
R2877 gnd.n245 gnd.n244 585
R2878 gnd.n248 gnd.n245 585
R2879 gnd.n7893 gnd.n7892 585
R2880 gnd.n7892 gnd.n7891 585
R2881 gnd.n7894 gnd.n240 585
R2882 gnd.n240 gnd.n239 585
R2883 gnd.n7896 gnd.n7895 585
R2884 gnd.n7897 gnd.n7896 585
R2885 gnd.n225 gnd.n224 585
R2886 gnd.n229 gnd.n225 585
R2887 gnd.n7905 gnd.n7904 585
R2888 gnd.n7904 gnd.n7903 585
R2889 gnd.n7906 gnd.n220 585
R2890 gnd.n226 gnd.n220 585
R2891 gnd.n7908 gnd.n7907 585
R2892 gnd.n7909 gnd.n7908 585
R2893 gnd.n207 gnd.n206 585
R2894 gnd.n210 gnd.n207 585
R2895 gnd.n7917 gnd.n7916 585
R2896 gnd.n7916 gnd.n7915 585
R2897 gnd.n7918 gnd.n202 585
R2898 gnd.n7741 gnd.n202 585
R2899 gnd.n7920 gnd.n7919 585
R2900 gnd.n7921 gnd.n7920 585
R2901 gnd.n187 gnd.n186 585
R2902 gnd.n198 gnd.n187 585
R2903 gnd.n7929 gnd.n7928 585
R2904 gnd.n7928 gnd.n7927 585
R2905 gnd.n7930 gnd.n182 585
R2906 gnd.n188 gnd.n182 585
R2907 gnd.n7932 gnd.n7931 585
R2908 gnd.n7933 gnd.n7932 585
R2909 gnd.n169 gnd.n168 585
R2910 gnd.n172 gnd.n169 585
R2911 gnd.n7941 gnd.n7940 585
R2912 gnd.n7940 gnd.n7939 585
R2913 gnd.n7942 gnd.n164 585
R2914 gnd.n164 gnd.n163 585
R2915 gnd.n7944 gnd.n7943 585
R2916 gnd.n7945 gnd.n7944 585
R2917 gnd.n149 gnd.n148 585
R2918 gnd.n160 gnd.n149 585
R2919 gnd.n7953 gnd.n7952 585
R2920 gnd.n7952 gnd.n7951 585
R2921 gnd.n7954 gnd.n144 585
R2922 gnd.n150 gnd.n144 585
R2923 gnd.n7956 gnd.n7955 585
R2924 gnd.n7957 gnd.n7956 585
R2925 gnd.n132 gnd.n131 585
R2926 gnd.n135 gnd.n132 585
R2927 gnd.n7965 gnd.n7964 585
R2928 gnd.n7964 gnd.n7963 585
R2929 gnd.n7966 gnd.n126 585
R2930 gnd.n126 gnd.n124 585
R2931 gnd.n7968 gnd.n7967 585
R2932 gnd.n7969 gnd.n7968 585
R2933 gnd.n127 gnd.n125 585
R2934 gnd.n125 gnd.n121 585
R2935 gnd.n7575 gnd.n7574 585
R2936 gnd.n7574 gnd.n106 585
R2937 gnd.n7573 gnd.n107 585
R2938 gnd.n7977 gnd.n107 585
R2939 gnd.n7572 gnd.n7571 585
R2940 gnd.n7571 gnd.n7570 585
R2941 gnd.n357 gnd.n355 585
R2942 gnd.n358 gnd.n357 585
R2943 gnd.n7563 gnd.n7562 585
R2944 gnd.n7562 gnd.n7561 585
R2945 gnd.n363 gnd.n362 585
R2946 gnd.n7553 gnd.n363 585
R2947 gnd.n7529 gnd.n7528 585
R2948 gnd.n7528 gnd.n368 585
R2949 gnd.n7530 gnd.n378 585
R2950 gnd.n7545 gnd.n378 585
R2951 gnd.n7532 gnd.n7531 585
R2952 gnd.n7531 gnd.n376 585
R2953 gnd.n7533 gnd.n387 585
R2954 gnd.n7519 gnd.n387 585
R2955 gnd.n7535 gnd.n7534 585
R2956 gnd.n7536 gnd.n7535 585
R2957 gnd.n388 gnd.n386 585
R2958 gnd.n7508 gnd.n386 585
R2959 gnd.n7481 gnd.n7480 585
R2960 gnd.n7480 gnd.n403 585
R2961 gnd.n7482 gnd.n414 585
R2962 gnd.n7497 gnd.n414 585
R2963 gnd.n7483 gnd.n425 585
R2964 gnd.n7471 gnd.n425 585
R2965 gnd.n7485 gnd.n7484 585
R2966 gnd.n7486 gnd.n7485 585
R2967 gnd.n426 gnd.n424 585
R2968 gnd.n7457 gnd.n424 585
R2969 gnd.n7433 gnd.n7432 585
R2970 gnd.n7432 gnd.n438 585
R2971 gnd.n7434 gnd.n449 585
R2972 gnd.n7448 gnd.n449 585
R2973 gnd.n7435 gnd.n461 585
R2974 gnd.n7424 gnd.n461 585
R2975 gnd.n7437 gnd.n7436 585
R2976 gnd.n7438 gnd.n7437 585
R2977 gnd.n462 gnd.n460 585
R2978 gnd.n7420 gnd.n460 585
R2979 gnd.n7396 gnd.n7395 585
R2980 gnd.n7395 gnd.n7394 585
R2981 gnd.n7397 gnd.n479 585
R2982 gnd.n7411 gnd.n479 585
R2983 gnd.n7398 gnd.n491 585
R2984 gnd.n7338 gnd.n491 585
R2985 gnd.n7400 gnd.n7399 585
R2986 gnd.n7401 gnd.n7400 585
R2987 gnd.n492 gnd.n490 585
R2988 gnd.n7371 gnd.n490 585
R2989 gnd.n7347 gnd.n7346 585
R2990 gnd.n7346 gnd.n504 585
R2991 gnd.n7348 gnd.n515 585
R2992 gnd.n7362 gnd.n515 585
R2993 gnd.n7349 gnd.n527 585
R2994 gnd.n7333 gnd.n527 585
R2995 gnd.n7351 gnd.n7350 585
R2996 gnd.n7352 gnd.n7351 585
R2997 gnd.n528 gnd.n526 585
R2998 gnd.n7329 gnd.n526 585
R2999 gnd.n561 gnd.n560 585
R3000 gnd.n560 gnd.n559 585
R3001 gnd.n558 gnd.n545 585
R3002 gnd.n7320 gnd.n545 585
R3003 gnd.n7307 gnd.n556 585
R3004 gnd.n7302 gnd.n556 585
R3005 gnd.n7309 gnd.n7308 585
R3006 gnd.n7310 gnd.n7309 585
R3007 gnd.n686 gnd.n555 585
R3008 gnd.n7151 gnd.n687 585
R3009 gnd.n7150 gnd.n688 585
R3010 gnd.n695 gnd.n689 585
R3011 gnd.n7143 gnd.n696 585
R3012 gnd.n7142 gnd.n697 585
R3013 gnd.n699 gnd.n698 585
R3014 gnd.n7135 gnd.n705 585
R3015 gnd.n7134 gnd.n706 585
R3016 gnd.n713 gnd.n707 585
R3017 gnd.n7127 gnd.n714 585
R3018 gnd.n7126 gnd.n715 585
R3019 gnd.n717 gnd.n716 585
R3020 gnd.n7119 gnd.n723 585
R3021 gnd.n7118 gnd.n724 585
R3022 gnd.n733 gnd.n725 585
R3023 gnd.n7111 gnd.n734 585
R3024 gnd.n7110 gnd.n7107 585
R3025 gnd.n735 gnd.n609 585
R3026 gnd.n7274 gnd.n609 585
R3027 gnd.n7723 gnd.n7722 585
R3028 gnd.n7716 gnd.n7669 585
R3029 gnd.n7718 gnd.n7717 585
R3030 gnd.n7715 gnd.n7714 585
R3031 gnd.n7713 gnd.n7712 585
R3032 gnd.n7706 gnd.n7671 585
R3033 gnd.n7708 gnd.n7707 585
R3034 gnd.n7705 gnd.n7704 585
R3035 gnd.n7703 gnd.n7702 585
R3036 gnd.n7696 gnd.n7673 585
R3037 gnd.n7698 gnd.n7697 585
R3038 gnd.n7695 gnd.n7694 585
R3039 gnd.n7693 gnd.n7692 585
R3040 gnd.n7686 gnd.n7675 585
R3041 gnd.n7688 gnd.n7687 585
R3042 gnd.n7685 gnd.n7684 585
R3043 gnd.n7683 gnd.n7682 585
R3044 gnd.n7679 gnd.n7678 585
R3045 gnd.n7677 gnd.n255 585
R3046 gnd.n7883 gnd.n255 585
R3047 gnd.n7725 gnd.n7724 585
R3048 gnd.n7724 gnd.n248 585
R3049 gnd.n7726 gnd.n247 585
R3050 gnd.n7891 gnd.n247 585
R3051 gnd.n7728 gnd.n7727 585
R3052 gnd.n7727 gnd.n239 585
R3053 gnd.n7729 gnd.n238 585
R3054 gnd.n7897 gnd.n238 585
R3055 gnd.n7731 gnd.n7730 585
R3056 gnd.n7730 gnd.n229 585
R3057 gnd.n7732 gnd.n228 585
R3058 gnd.n7903 gnd.n228 585
R3059 gnd.n7734 gnd.n7733 585
R3060 gnd.n7733 gnd.n226 585
R3061 gnd.n7735 gnd.n219 585
R3062 gnd.n7909 gnd.n219 585
R3063 gnd.n7737 gnd.n7736 585
R3064 gnd.n7736 gnd.n210 585
R3065 gnd.n7738 gnd.n209 585
R3066 gnd.n7915 gnd.n209 585
R3067 gnd.n7740 gnd.n7739 585
R3068 gnd.n7741 gnd.n7740 585
R3069 gnd.n7610 gnd.n200 585
R3070 gnd.n7921 gnd.n200 585
R3071 gnd.n7653 gnd.n7652 585
R3072 gnd.n7652 gnd.n198 585
R3073 gnd.n7651 gnd.n190 585
R3074 gnd.n7927 gnd.n190 585
R3075 gnd.n7650 gnd.n7649 585
R3076 gnd.n7649 gnd.n188 585
R3077 gnd.n7612 gnd.n181 585
R3078 gnd.n7933 gnd.n181 585
R3079 gnd.n7645 gnd.n7644 585
R3080 gnd.n7644 gnd.n172 585
R3081 gnd.n7643 gnd.n171 585
R3082 gnd.n7939 gnd.n171 585
R3083 gnd.n7642 gnd.n7641 585
R3084 gnd.n7641 gnd.n163 585
R3085 gnd.n7614 gnd.n162 585
R3086 gnd.n7945 gnd.n162 585
R3087 gnd.n7637 gnd.n7636 585
R3088 gnd.n7636 gnd.n160 585
R3089 gnd.n7635 gnd.n152 585
R3090 gnd.n7951 gnd.n152 585
R3091 gnd.n7634 gnd.n7633 585
R3092 gnd.n7633 gnd.n150 585
R3093 gnd.n7616 gnd.n143 585
R3094 gnd.n7957 gnd.n143 585
R3095 gnd.n7629 gnd.n7628 585
R3096 gnd.n7628 gnd.n135 585
R3097 gnd.n7627 gnd.n134 585
R3098 gnd.n7963 gnd.n134 585
R3099 gnd.n7626 gnd.n7625 585
R3100 gnd.n7625 gnd.n124 585
R3101 gnd.n7618 gnd.n123 585
R3102 gnd.n7969 gnd.n123 585
R3103 gnd.n7621 gnd.n7620 585
R3104 gnd.n7620 gnd.n121 585
R3105 gnd.n104 gnd.n103 585
R3106 gnd.n106 gnd.n104 585
R3107 gnd.n7979 gnd.n7978 585
R3108 gnd.n7978 gnd.n7977 585
R3109 gnd.n7980 gnd.n102 585
R3110 gnd.n7570 gnd.n102 585
R3111 gnd.n365 gnd.n100 585
R3112 gnd.n365 gnd.n358 585
R3113 gnd.n372 gnd.n366 585
R3114 gnd.n7561 gnd.n366 585
R3115 gnd.n7552 gnd.n7551 585
R3116 gnd.n7553 gnd.n7552 585
R3117 gnd.n371 gnd.n370 585
R3118 gnd.n370 gnd.n368 585
R3119 gnd.n7547 gnd.n7546 585
R3120 gnd.n7546 gnd.n7545 585
R3121 gnd.n375 gnd.n374 585
R3122 gnd.n376 gnd.n375 585
R3123 gnd.n7502 gnd.n395 585
R3124 gnd.n7519 gnd.n395 585
R3125 gnd.n407 gnd.n385 585
R3126 gnd.n7536 gnd.n385 585
R3127 gnd.n7507 gnd.n7506 585
R3128 gnd.n7508 gnd.n7507 585
R3129 gnd.n406 gnd.n405 585
R3130 gnd.n405 gnd.n403 585
R3131 gnd.n7499 gnd.n7498 585
R3132 gnd.n7498 gnd.n7497 585
R3133 gnd.n410 gnd.n409 585
R3134 gnd.n7471 gnd.n410 585
R3135 gnd.n442 gnd.n423 585
R3136 gnd.n7486 gnd.n423 585
R3137 gnd.n7456 gnd.n7455 585
R3138 gnd.n7457 gnd.n7456 585
R3139 gnd.n441 gnd.n440 585
R3140 gnd.n440 gnd.n438 585
R3141 gnd.n7450 gnd.n7449 585
R3142 gnd.n7449 gnd.n7448 585
R3143 gnd.n445 gnd.n444 585
R3144 gnd.n7424 gnd.n445 585
R3145 gnd.n473 gnd.n458 585
R3146 gnd.n7438 gnd.n458 585
R3147 gnd.n7419 gnd.n7418 585
R3148 gnd.n7420 gnd.n7419 585
R3149 gnd.n472 gnd.n471 585
R3150 gnd.n7394 gnd.n471 585
R3151 gnd.n7413 gnd.n7412 585
R3152 gnd.n7412 gnd.n7411 585
R3153 gnd.n476 gnd.n475 585
R3154 gnd.n7338 gnd.n476 585
R3155 gnd.n508 gnd.n488 585
R3156 gnd.n7401 gnd.n488 585
R3157 gnd.n7370 gnd.n7369 585
R3158 gnd.n7371 gnd.n7370 585
R3159 gnd.n507 gnd.n506 585
R3160 gnd.n506 gnd.n504 585
R3161 gnd.n7364 gnd.n7363 585
R3162 gnd.n7363 gnd.n7362 585
R3163 gnd.n511 gnd.n510 585
R3164 gnd.n7333 gnd.n511 585
R3165 gnd.n539 gnd.n524 585
R3166 gnd.n7352 gnd.n524 585
R3167 gnd.n7328 gnd.n7327 585
R3168 gnd.n7329 gnd.n7328 585
R3169 gnd.n538 gnd.n537 585
R3170 gnd.n559 gnd.n537 585
R3171 gnd.n7322 gnd.n7321 585
R3172 gnd.n7321 gnd.n7320 585
R3173 gnd.n542 gnd.n541 585
R3174 gnd.n7302 gnd.n542 585
R3175 gnd.n7099 gnd.n553 585
R3176 gnd.n7310 gnd.n553 585
R3177 gnd.n5207 gnd.n3842 585
R3178 gnd.n3842 gnd.n3149 585
R3179 gnd.n5208 gnd.n3903 585
R3180 gnd.n3903 gnd.n3893 585
R3181 gnd.n5210 gnd.n5209 585
R3182 gnd.n5211 gnd.n5210 585
R3183 gnd.n3904 gnd.n3902 585
R3184 gnd.n3911 gnd.n3902 585
R3185 gnd.n5201 gnd.n5200 585
R3186 gnd.n5200 gnd.n5199 585
R3187 gnd.n3907 gnd.n3906 585
R3188 gnd.n4926 gnd.n3907 585
R3189 gnd.n4912 gnd.n3930 585
R3190 gnd.n3930 gnd.n3920 585
R3191 gnd.n4914 gnd.n4913 585
R3192 gnd.n4915 gnd.n4914 585
R3193 gnd.n3931 gnd.n3929 585
R3194 gnd.n3929 gnd.n3927 585
R3195 gnd.n4907 gnd.n4906 585
R3196 gnd.n4906 gnd.n4905 585
R3197 gnd.n3934 gnd.n3933 585
R3198 gnd.n3943 gnd.n3934 585
R3199 gnd.n4863 gnd.n3957 585
R3200 gnd.n3957 gnd.n3942 585
R3201 gnd.n4865 gnd.n4864 585
R3202 gnd.n4866 gnd.n4865 585
R3203 gnd.n3958 gnd.n3956 585
R3204 gnd.n3965 gnd.n3956 585
R3205 gnd.n4858 gnd.n4857 585
R3206 gnd.n4857 gnd.n4856 585
R3207 gnd.n3961 gnd.n3960 585
R3208 gnd.n4837 gnd.n3961 585
R3209 gnd.n4823 gnd.n3985 585
R3210 gnd.n3985 gnd.n3974 585
R3211 gnd.n4825 gnd.n4824 585
R3212 gnd.n4826 gnd.n4825 585
R3213 gnd.n3986 gnd.n3984 585
R3214 gnd.n3984 gnd.n3981 585
R3215 gnd.n4818 gnd.n4817 585
R3216 gnd.n4817 gnd.n4816 585
R3217 gnd.n3989 gnd.n3988 585
R3218 gnd.n3999 gnd.n3989 585
R3219 gnd.n4778 gnd.n4012 585
R3220 gnd.n4012 gnd.n3998 585
R3221 gnd.n4780 gnd.n4779 585
R3222 gnd.n4781 gnd.n4780 585
R3223 gnd.n4013 gnd.n4011 585
R3224 gnd.n4020 gnd.n4011 585
R3225 gnd.n4773 gnd.n4772 585
R3226 gnd.n4772 gnd.n4771 585
R3227 gnd.n4016 gnd.n4015 585
R3228 gnd.n4752 gnd.n4016 585
R3229 gnd.n4738 gnd.n4039 585
R3230 gnd.n4039 gnd.n4029 585
R3231 gnd.n4740 gnd.n4739 585
R3232 gnd.n4741 gnd.n4740 585
R3233 gnd.n4040 gnd.n4038 585
R3234 gnd.n4729 gnd.n4038 585
R3235 gnd.n4733 gnd.n4732 585
R3236 gnd.n4732 gnd.n4731 585
R3237 gnd.n4043 gnd.n4042 585
R3238 gnd.n4684 gnd.n4043 585
R3239 gnd.n4177 gnd.n4176 585
R3240 gnd.n4178 gnd.n4177 585
R3241 gnd.n4157 gnd.n4156 585
R3242 gnd.n4160 gnd.n4157 585
R3243 gnd.n4694 gnd.n4693 585
R3244 gnd.n4693 gnd.n4692 585
R3245 gnd.n4695 gnd.n4151 585
R3246 gnd.n4187 gnd.n4151 585
R3247 gnd.n4697 gnd.n4696 585
R3248 gnd.n4698 gnd.n4697 585
R3249 gnd.n4152 gnd.n4150 585
R3250 gnd.n4662 gnd.n4150 585
R3251 gnd.n4646 gnd.n4645 585
R3252 gnd.n4645 gnd.n4138 585
R3253 gnd.n4647 gnd.n4202 585
R3254 gnd.n4202 gnd.n4137 585
R3255 gnd.n4649 gnd.n4648 585
R3256 gnd.n4650 gnd.n4649 585
R3257 gnd.n4203 gnd.n4201 585
R3258 gnd.n4201 gnd.n4198 585
R3259 gnd.n4638 gnd.n4637 585
R3260 gnd.n4637 gnd.n4636 585
R3261 gnd.n4206 gnd.n4205 585
R3262 gnd.n4213 gnd.n4206 585
R3263 gnd.n4612 gnd.n4611 585
R3264 gnd.n4613 gnd.n4612 585
R3265 gnd.n4225 gnd.n4224 585
R3266 gnd.n4232 gnd.n4224 585
R3267 gnd.n4607 gnd.n4606 585
R3268 gnd.n4606 gnd.n4605 585
R3269 gnd.n4228 gnd.n4227 585
R3270 gnd.n4595 gnd.n4228 585
R3271 gnd.n4582 gnd.n4252 585
R3272 gnd.n4252 gnd.n4251 585
R3273 gnd.n4584 gnd.n4583 585
R3274 gnd.n4585 gnd.n4584 585
R3275 gnd.n4253 gnd.n4250 585
R3276 gnd.n4260 gnd.n4250 585
R3277 gnd.n4577 gnd.n4576 585
R3278 gnd.n4576 gnd.n4575 585
R3279 gnd.n4256 gnd.n4255 585
R3280 gnd.n4564 gnd.n4256 585
R3281 gnd.n4551 gnd.n4277 585
R3282 gnd.n4277 gnd.n4276 585
R3283 gnd.n4553 gnd.n4552 585
R3284 gnd.n4554 gnd.n4553 585
R3285 gnd.n4547 gnd.n4275 585
R3286 gnd.n4546 gnd.n4545 585
R3287 gnd.n4280 gnd.n4279 585
R3288 gnd.n4543 gnd.n4280 585
R3289 gnd.n4302 gnd.n4301 585
R3290 gnd.n4305 gnd.n4304 585
R3291 gnd.n4303 gnd.n4298 585
R3292 gnd.n4310 gnd.n4309 585
R3293 gnd.n4312 gnd.n4311 585
R3294 gnd.n4315 gnd.n4314 585
R3295 gnd.n4313 gnd.n4296 585
R3296 gnd.n4320 gnd.n4319 585
R3297 gnd.n4322 gnd.n4321 585
R3298 gnd.n4325 gnd.n4324 585
R3299 gnd.n4323 gnd.n4294 585
R3300 gnd.n4330 gnd.n4329 585
R3301 gnd.n4334 gnd.n4331 585
R3302 gnd.n4335 gnd.n4272 585
R3303 gnd.n5213 gnd.n3857 585
R3304 gnd.n5280 gnd.n5279 585
R3305 gnd.n5282 gnd.n5281 585
R3306 gnd.n5284 gnd.n5283 585
R3307 gnd.n5286 gnd.n5285 585
R3308 gnd.n5288 gnd.n5287 585
R3309 gnd.n5290 gnd.n5289 585
R3310 gnd.n5292 gnd.n5291 585
R3311 gnd.n5294 gnd.n5293 585
R3312 gnd.n5296 gnd.n5295 585
R3313 gnd.n5298 gnd.n5297 585
R3314 gnd.n5300 gnd.n5299 585
R3315 gnd.n5302 gnd.n5301 585
R3316 gnd.n5305 gnd.n5304 585
R3317 gnd.n5303 gnd.n3845 585
R3318 gnd.n5309 gnd.n3843 585
R3319 gnd.n5311 gnd.n5310 585
R3320 gnd.n5312 gnd.n5311 585
R3321 gnd.n5214 gnd.n3898 585
R3322 gnd.n5214 gnd.n3149 585
R3323 gnd.n5216 gnd.n5215 585
R3324 gnd.n5215 gnd.n3893 585
R3325 gnd.n5212 gnd.n3897 585
R3326 gnd.n5212 gnd.n5211 585
R3327 gnd.n5191 gnd.n3899 585
R3328 gnd.n3911 gnd.n3899 585
R3329 gnd.n5190 gnd.n3909 585
R3330 gnd.n5199 gnd.n3909 585
R3331 gnd.n4925 gnd.n3916 585
R3332 gnd.n4926 gnd.n4925 585
R3333 gnd.n4924 gnd.n4923 585
R3334 gnd.n4924 gnd.n3920 585
R3335 gnd.n4922 gnd.n3922 585
R3336 gnd.n4915 gnd.n3922 585
R3337 gnd.n3935 gnd.n3923 585
R3338 gnd.n3935 gnd.n3927 585
R3339 gnd.n4871 gnd.n3936 585
R3340 gnd.n4905 gnd.n3936 585
R3341 gnd.n4870 gnd.n4869 585
R3342 gnd.n4869 gnd.n3943 585
R3343 gnd.n4868 gnd.n3951 585
R3344 gnd.n4868 gnd.n3942 585
R3345 gnd.n4867 gnd.n3953 585
R3346 gnd.n4867 gnd.n4866 585
R3347 gnd.n4846 gnd.n3952 585
R3348 gnd.n3965 gnd.n3952 585
R3349 gnd.n4845 gnd.n3963 585
R3350 gnd.n4856 gnd.n3963 585
R3351 gnd.n4836 gnd.n3970 585
R3352 gnd.n4837 gnd.n4836 585
R3353 gnd.n4835 gnd.n4834 585
R3354 gnd.n4835 gnd.n3974 585
R3355 gnd.n4833 gnd.n3976 585
R3356 gnd.n4826 gnd.n3976 585
R3357 gnd.n3991 gnd.n3977 585
R3358 gnd.n3991 gnd.n3981 585
R3359 gnd.n4786 gnd.n3992 585
R3360 gnd.n4816 gnd.n3992 585
R3361 gnd.n4785 gnd.n4784 585
R3362 gnd.n4784 gnd.n3999 585
R3363 gnd.n4783 gnd.n4006 585
R3364 gnd.n4783 gnd.n3998 585
R3365 gnd.n4782 gnd.n4008 585
R3366 gnd.n4782 gnd.n4781 585
R3367 gnd.n4761 gnd.n4007 585
R3368 gnd.n4020 gnd.n4007 585
R3369 gnd.n4760 gnd.n4018 585
R3370 gnd.n4771 gnd.n4018 585
R3371 gnd.n4751 gnd.n4025 585
R3372 gnd.n4752 gnd.n4751 585
R3373 gnd.n4750 gnd.n4749 585
R3374 gnd.n4750 gnd.n4029 585
R3375 gnd.n4748 gnd.n4031 585
R3376 gnd.n4741 gnd.n4031 585
R3377 gnd.n4728 gnd.n4032 585
R3378 gnd.n4729 gnd.n4728 585
R3379 gnd.n4681 gnd.n4045 585
R3380 gnd.n4731 gnd.n4045 585
R3381 gnd.n4683 gnd.n4682 585
R3382 gnd.n4684 gnd.n4683 585
R3383 gnd.n4676 gnd.n4179 585
R3384 gnd.n4179 gnd.n4178 585
R3385 gnd.n4674 gnd.n4673 585
R3386 gnd.n4673 gnd.n4160 585
R3387 gnd.n4671 gnd.n4158 585
R3388 gnd.n4692 gnd.n4158 585
R3389 gnd.n4189 gnd.n4188 585
R3390 gnd.n4188 gnd.n4187 585
R3391 gnd.n4665 gnd.n4148 585
R3392 gnd.n4698 gnd.n4148 585
R3393 gnd.n4664 gnd.n4663 585
R3394 gnd.n4663 gnd.n4662 585
R3395 gnd.n4660 gnd.n4191 585
R3396 gnd.n4660 gnd.n4138 585
R3397 gnd.n4659 gnd.n4658 585
R3398 gnd.n4659 gnd.n4137 585
R3399 gnd.n4194 gnd.n4193 585
R3400 gnd.n4650 gnd.n4193 585
R3401 gnd.n4618 gnd.n4617 585
R3402 gnd.n4617 gnd.n4198 585
R3403 gnd.n4619 gnd.n4207 585
R3404 gnd.n4636 gnd.n4207 585
R3405 gnd.n4616 gnd.n4615 585
R3406 gnd.n4615 gnd.n4213 585
R3407 gnd.n4614 gnd.n4221 585
R3408 gnd.n4614 gnd.n4613 585
R3409 gnd.n4599 gnd.n4222 585
R3410 gnd.n4232 gnd.n4222 585
R3411 gnd.n4598 gnd.n4230 585
R3412 gnd.n4605 gnd.n4230 585
R3413 gnd.n4597 gnd.n4596 585
R3414 gnd.n4596 gnd.n4595 585
R3415 gnd.n4241 gnd.n4238 585
R3416 gnd.n4251 gnd.n4241 585
R3417 gnd.n4587 gnd.n4586 585
R3418 gnd.n4586 gnd.n4585 585
R3419 gnd.n4247 gnd.n4246 585
R3420 gnd.n4260 gnd.n4247 585
R3421 gnd.n4567 gnd.n4258 585
R3422 gnd.n4575 gnd.n4258 585
R3423 gnd.n4566 gnd.n4565 585
R3424 gnd.n4565 gnd.n4564 585
R3425 gnd.n4267 gnd.n4265 585
R3426 gnd.n4276 gnd.n4267 585
R3427 gnd.n4556 gnd.n4555 585
R3428 gnd.n4555 gnd.n4554 585
R3429 gnd.n6788 gnd.n6510 585
R3430 gnd.n6510 gnd.n840 585
R3431 gnd.n6790 gnd.n6789 585
R3432 gnd.n6791 gnd.n6790 585
R3433 gnd.n6511 gnd.n6509 585
R3434 gnd.n6509 gnd.n849 585
R3435 gnd.n6659 gnd.n6658 585
R3436 gnd.n6660 gnd.n6659 585
R3437 gnd.n6657 gnd.n6584 585
R3438 gnd.n6652 gnd.n6584 585
R3439 gnd.n6656 gnd.n6655 585
R3440 gnd.n6655 gnd.n6654 585
R3441 gnd.n6586 gnd.n6585 585
R3442 gnd.n6586 gnd.n855 585
R3443 gnd.n6644 gnd.n6643 585
R3444 gnd.n6645 gnd.n6644 585
R3445 gnd.n6642 gnd.n6591 585
R3446 gnd.n6591 gnd.n864 585
R3447 gnd.n6641 gnd.n6640 585
R3448 gnd.n6640 gnd.n862 585
R3449 gnd.n6639 gnd.n6592 585
R3450 gnd.n6639 gnd.n6638 585
R3451 gnd.n6626 gnd.n6593 585
R3452 gnd.n6594 gnd.n6593 585
R3453 gnd.n6627 gnd.n6602 585
R3454 gnd.n6602 gnd.n870 585
R3455 gnd.n6629 gnd.n6628 585
R3456 gnd.n6630 gnd.n6629 585
R3457 gnd.n6625 gnd.n6601 585
R3458 gnd.n6601 gnd.n6599 585
R3459 gnd.n6624 gnd.n6623 585
R3460 gnd.n6623 gnd.n877 585
R3461 gnd.n6622 gnd.n6603 585
R3462 gnd.n6622 gnd.n6621 585
R3463 gnd.n6607 gnd.n6606 585
R3464 gnd.n6608 gnd.n6607 585
R3465 gnd.n6605 gnd.n6604 585
R3466 gnd.n6604 gnd.n884 585
R3467 gnd.n968 gnd.n967 585
R3468 gnd.n6858 gnd.n968 585
R3469 gnd.n6861 gnd.n6860 585
R3470 gnd.n6860 gnd.n6859 585
R3471 gnd.n6862 gnd.n964 585
R3472 gnd.n964 gnd.n891 585
R3473 gnd.n6864 gnd.n6863 585
R3474 gnd.n6865 gnd.n6864 585
R3475 gnd.n966 gnd.n963 585
R3476 gnd.n963 gnd.n961 585
R3477 gnd.n965 gnd.n952 585
R3478 gnd.n6871 gnd.n952 585
R3479 gnd.n6874 gnd.n951 585
R3480 gnd.n6874 gnd.n6873 585
R3481 gnd.n6876 gnd.n6875 585
R3482 gnd.n6875 gnd.n905 585
R3483 gnd.n6877 gnd.n949 585
R3484 gnd.n949 gnd.n948 585
R3485 gnd.n6879 gnd.n6878 585
R3486 gnd.n6880 gnd.n6879 585
R3487 gnd.n950 gnd.n947 585
R3488 gnd.n947 gnd.n912 585
R3489 gnd.n939 gnd.n938 585
R3490 gnd.n6886 gnd.n939 585
R3491 gnd.n6890 gnd.n6889 585
R3492 gnd.n6889 gnd.n6888 585
R3493 gnd.n6891 gnd.n936 585
R3494 gnd.n936 gnd.n919 585
R3495 gnd.n6893 gnd.n6892 585
R3496 gnd.n6894 gnd.n6893 585
R3497 gnd.n937 gnd.n935 585
R3498 gnd.n935 gnd.n927 585
R3499 gnd.n6445 gnd.n925 585
R3500 gnd.n6900 gnd.n925 585
R3501 gnd.n6447 gnd.n6446 585
R3502 gnd.n6448 gnd.n6447 585
R3503 gnd.n6444 gnd.n1004 585
R3504 gnd.n1004 gnd.n1003 585
R3505 gnd.n6443 gnd.n6442 585
R3506 gnd.n6442 gnd.n6441 585
R3507 gnd.n1006 gnd.n1005 585
R3508 gnd.n1006 gnd.n985 585
R3509 gnd.n6429 gnd.n1013 585
R3510 gnd.n1013 gnd.n984 585
R3511 gnd.n6431 gnd.n6430 585
R3512 gnd.n6432 gnd.n6431 585
R3513 gnd.n6428 gnd.n1012 585
R3514 gnd.n1012 gnd.n995 585
R3515 gnd.n6427 gnd.n6426 585
R3516 gnd.n6426 gnd.n993 585
R3517 gnd.n6425 gnd.n1014 585
R3518 gnd.n6425 gnd.n6424 585
R3519 gnd.n6377 gnd.n1015 585
R3520 gnd.n6394 gnd.n1015 585
R3521 gnd.n6379 gnd.n6378 585
R3522 gnd.n6378 gnd.n1024 585
R3523 gnd.n6380 gnd.n1046 585
R3524 gnd.n1046 gnd.n1023 585
R3525 gnd.n6382 gnd.n6381 585
R3526 gnd.n6383 gnd.n6382 585
R3527 gnd.n6376 gnd.n1045 585
R3528 gnd.n1045 gnd.n1034 585
R3529 gnd.n6375 gnd.n6374 585
R3530 gnd.n6374 gnd.n1032 585
R3531 gnd.n6373 gnd.n1047 585
R3532 gnd.n6373 gnd.n6372 585
R3533 gnd.n6361 gnd.n1048 585
R3534 gnd.n1054 gnd.n1048 585
R3535 gnd.n6363 gnd.n6362 585
R3536 gnd.n6364 gnd.n6363 585
R3537 gnd.n6360 gnd.n1056 585
R3538 gnd.n1062 gnd.n1056 585
R3539 gnd.n6359 gnd.n6358 585
R3540 gnd.n6358 gnd.n6357 585
R3541 gnd.n1058 gnd.n1057 585
R3542 gnd.n5948 gnd.n1058 585
R3543 gnd.n5966 gnd.n5803 585
R3544 gnd.n5803 gnd.n1071 585
R3545 gnd.n5968 gnd.n5967 585
R3546 gnd.n5969 gnd.n5968 585
R3547 gnd.n5965 gnd.n5802 585
R3548 gnd.n5802 gnd.n5800 585
R3549 gnd.n5964 gnd.n1080 585
R3550 gnd.n6332 gnd.n1080 585
R3551 gnd.n5963 gnd.n5962 585
R3552 gnd.n5962 gnd.n1079 585
R3553 gnd.n5961 gnd.n5804 585
R3554 gnd.n5961 gnd.n5960 585
R3555 gnd.n5939 gnd.n5805 585
R3556 gnd.n5805 gnd.n1088 585
R3557 gnd.n5941 gnd.n5940 585
R3558 gnd.n5942 gnd.n5941 585
R3559 gnd.n5938 gnd.n5812 585
R3560 gnd.n5812 gnd.n5811 585
R3561 gnd.n5937 gnd.n5936 585
R3562 gnd.n5936 gnd.n1095 585
R3563 gnd.n5935 gnd.n5813 585
R3564 gnd.n5935 gnd.n5934 585
R3565 gnd.n5922 gnd.n5814 585
R3566 gnd.n5816 gnd.n5814 585
R3567 gnd.n5923 gnd.n5824 585
R3568 gnd.n5824 gnd.n1102 585
R3569 gnd.n5925 gnd.n5924 585
R3570 gnd.n5926 gnd.n5925 585
R3571 gnd.n5921 gnd.n5823 585
R3572 gnd.n5823 gnd.n5822 585
R3573 gnd.n5920 gnd.n5919 585
R3574 gnd.n5919 gnd.n5918 585
R3575 gnd.n5826 gnd.n5825 585
R3576 gnd.n5828 gnd.n5826 585
R3577 gnd.n5907 gnd.n5835 585
R3578 gnd.n5835 gnd.n1116 585
R3579 gnd.n5909 gnd.n5908 585
R3580 gnd.n5910 gnd.n5909 585
R3581 gnd.n5906 gnd.n5834 585
R3582 gnd.n5834 gnd.n5833 585
R3583 gnd.n5905 gnd.n5904 585
R3584 gnd.n5904 gnd.n1123 585
R3585 gnd.n5903 gnd.n5836 585
R3586 gnd.n5903 gnd.n5902 585
R3587 gnd.n5889 gnd.n5837 585
R3588 gnd.n5839 gnd.n5837 585
R3589 gnd.n5890 gnd.n5847 585
R3590 gnd.n5847 gnd.n1130 585
R3591 gnd.n5892 gnd.n5891 585
R3592 gnd.n5893 gnd.n5892 585
R3593 gnd.n5888 gnd.n5846 585
R3594 gnd.n5846 gnd.n5845 585
R3595 gnd.n5887 gnd.n5886 585
R3596 gnd.n5886 gnd.n1137 585
R3597 gnd.n5885 gnd.n5848 585
R3598 gnd.n5885 gnd.n5884 585
R3599 gnd.n5868 gnd.n5849 585
R3600 gnd.n5850 gnd.n5849 585
R3601 gnd.n5870 gnd.n5869 585
R3602 gnd.n5869 gnd.n1145 585
R3603 gnd.n5871 gnd.n5865 585
R3604 gnd.n5865 gnd.n1143 585
R3605 gnd.n5873 gnd.n5872 585
R3606 gnd.n5874 gnd.n5873 585
R3607 gnd.n5867 gnd.n5864 585
R3608 gnd.n5864 gnd.n1153 585
R3609 gnd.n5866 gnd.n1433 585
R3610 gnd.n1433 gnd.n1151 585
R3611 gnd.n6024 gnd.n1432 585
R3612 gnd.n6024 gnd.n6023 585
R3613 gnd.n6026 gnd.n6025 585
R3614 gnd.n6025 gnd.n1160 585
R3615 gnd.n6027 gnd.n1327 585
R3616 gnd.n1327 gnd.n1326 585
R3617 gnd.n6029 gnd.n6028 585
R3618 gnd.n6030 gnd.n6029 585
R3619 gnd.n1431 gnd.n1325 585
R3620 gnd.n1325 gnd.n1167 585
R3621 gnd.n1429 gnd.n1428 585
R3622 gnd.n1426 gnd.n1348 585
R3623 gnd.n1425 gnd.n1424 585
R3624 gnd.n1425 gnd.n1174 585
R3625 gnd.n1423 gnd.n1349 585
R3626 gnd.n1422 gnd.n1421 585
R3627 gnd.n1419 gnd.n1350 585
R3628 gnd.n1417 gnd.n1416 585
R3629 gnd.n1415 gnd.n1351 585
R3630 gnd.n1414 gnd.n1413 585
R3631 gnd.n1411 gnd.n1352 585
R3632 gnd.n1409 gnd.n1408 585
R3633 gnd.n1407 gnd.n1353 585
R3634 gnd.n1406 gnd.n1405 585
R3635 gnd.n1403 gnd.n1354 585
R3636 gnd.n1401 gnd.n1400 585
R3637 gnd.n1399 gnd.n1355 585
R3638 gnd.n1398 gnd.n1397 585
R3639 gnd.n1395 gnd.n1356 585
R3640 gnd.n1393 gnd.n1392 585
R3641 gnd.n1391 gnd.n1357 585
R3642 gnd.n1390 gnd.n1389 585
R3643 gnd.n1387 gnd.n1358 585
R3644 gnd.n1385 gnd.n1384 585
R3645 gnd.n1383 gnd.n1359 585
R3646 gnd.n1382 gnd.n1381 585
R3647 gnd.n1379 gnd.n1360 585
R3648 gnd.n1377 gnd.n1376 585
R3649 gnd.n1375 gnd.n1361 585
R3650 gnd.n1374 gnd.n1373 585
R3651 gnd.n1371 gnd.n1370 585
R3652 gnd.n1369 gnd.n1368 585
R3653 gnd.n1367 gnd.n1302 585
R3654 gnd.n6100 gnd.n6099 585
R3655 gnd.n6097 gnd.n1301 585
R3656 gnd.n6095 gnd.n6094 585
R3657 gnd.n6093 gnd.n1304 585
R3658 gnd.n6091 gnd.n6090 585
R3659 gnd.n6088 gnd.n1307 585
R3660 gnd.n6086 gnd.n6085 585
R3661 gnd.n6084 gnd.n1308 585
R3662 gnd.n6083 gnd.n6082 585
R3663 gnd.n6080 gnd.n1309 585
R3664 gnd.n6078 gnd.n6077 585
R3665 gnd.n6076 gnd.n1310 585
R3666 gnd.n6075 gnd.n6074 585
R3667 gnd.n6072 gnd.n1311 585
R3668 gnd.n6070 gnd.n6069 585
R3669 gnd.n6068 gnd.n1312 585
R3670 gnd.n6067 gnd.n6066 585
R3671 gnd.n6064 gnd.n1313 585
R3672 gnd.n6062 gnd.n6061 585
R3673 gnd.n6060 gnd.n1314 585
R3674 gnd.n6059 gnd.n6058 585
R3675 gnd.n6056 gnd.n1315 585
R3676 gnd.n6054 gnd.n6053 585
R3677 gnd.n6052 gnd.n1316 585
R3678 gnd.n6051 gnd.n6050 585
R3679 gnd.n6048 gnd.n1317 585
R3680 gnd.n6046 gnd.n6045 585
R3681 gnd.n6044 gnd.n1318 585
R3682 gnd.n6043 gnd.n6042 585
R3683 gnd.n6040 gnd.n1319 585
R3684 gnd.n6038 gnd.n6037 585
R3685 gnd.n6036 gnd.n1320 585
R3686 gnd.n6035 gnd.n6034 585
R3687 gnd.n6669 gnd.n6668 585
R3688 gnd.n6670 gnd.n6581 585
R3689 gnd.n6672 gnd.n6671 585
R3690 gnd.n6674 gnd.n6579 585
R3691 gnd.n6676 gnd.n6675 585
R3692 gnd.n6677 gnd.n6578 585
R3693 gnd.n6679 gnd.n6678 585
R3694 gnd.n6681 gnd.n6576 585
R3695 gnd.n6683 gnd.n6682 585
R3696 gnd.n6684 gnd.n6575 585
R3697 gnd.n6686 gnd.n6685 585
R3698 gnd.n6688 gnd.n6573 585
R3699 gnd.n6690 gnd.n6689 585
R3700 gnd.n6691 gnd.n6572 585
R3701 gnd.n6693 gnd.n6692 585
R3702 gnd.n6695 gnd.n6570 585
R3703 gnd.n6697 gnd.n6696 585
R3704 gnd.n6698 gnd.n6569 585
R3705 gnd.n6700 gnd.n6699 585
R3706 gnd.n6702 gnd.n6567 585
R3707 gnd.n6704 gnd.n6703 585
R3708 gnd.n6705 gnd.n6566 585
R3709 gnd.n6707 gnd.n6706 585
R3710 gnd.n6709 gnd.n6564 585
R3711 gnd.n6711 gnd.n6710 585
R3712 gnd.n6712 gnd.n6563 585
R3713 gnd.n6714 gnd.n6713 585
R3714 gnd.n6716 gnd.n6561 585
R3715 gnd.n6718 gnd.n6717 585
R3716 gnd.n6720 gnd.n6558 585
R3717 gnd.n6722 gnd.n6721 585
R3718 gnd.n6724 gnd.n6557 585
R3719 gnd.n6725 gnd.n6532 585
R3720 gnd.n6728 gnd.n639 585
R3721 gnd.n6730 gnd.n6729 585
R3722 gnd.n6732 gnd.n6555 585
R3723 gnd.n6734 gnd.n6733 585
R3724 gnd.n6736 gnd.n6552 585
R3725 gnd.n6738 gnd.n6737 585
R3726 gnd.n6740 gnd.n6550 585
R3727 gnd.n6742 gnd.n6741 585
R3728 gnd.n6743 gnd.n6549 585
R3729 gnd.n6745 gnd.n6744 585
R3730 gnd.n6747 gnd.n6547 585
R3731 gnd.n6749 gnd.n6748 585
R3732 gnd.n6750 gnd.n6546 585
R3733 gnd.n6752 gnd.n6751 585
R3734 gnd.n6754 gnd.n6544 585
R3735 gnd.n6756 gnd.n6755 585
R3736 gnd.n6757 gnd.n6543 585
R3737 gnd.n6759 gnd.n6758 585
R3738 gnd.n6761 gnd.n6541 585
R3739 gnd.n6763 gnd.n6762 585
R3740 gnd.n6764 gnd.n6540 585
R3741 gnd.n6766 gnd.n6765 585
R3742 gnd.n6768 gnd.n6538 585
R3743 gnd.n6770 gnd.n6769 585
R3744 gnd.n6771 gnd.n6537 585
R3745 gnd.n6773 gnd.n6772 585
R3746 gnd.n6775 gnd.n6535 585
R3747 gnd.n6777 gnd.n6776 585
R3748 gnd.n6778 gnd.n6534 585
R3749 gnd.n6780 gnd.n6779 585
R3750 gnd.n6782 gnd.n6533 585
R3751 gnd.n6783 gnd.n6531 585
R3752 gnd.n6786 gnd.n6785 585
R3753 gnd.n6667 gnd.n6665 585
R3754 gnd.n6667 gnd.n840 585
R3755 gnd.n6664 gnd.n6508 585
R3756 gnd.n6791 gnd.n6508 585
R3757 gnd.n6663 gnd.n6662 585
R3758 gnd.n6662 gnd.n849 585
R3759 gnd.n6661 gnd.n6582 585
R3760 gnd.n6661 gnd.n6660 585
R3761 gnd.n6649 gnd.n6583 585
R3762 gnd.n6652 gnd.n6583 585
R3763 gnd.n6651 gnd.n6650 585
R3764 gnd.n6654 gnd.n6651 585
R3765 gnd.n6648 gnd.n6587 585
R3766 gnd.n6587 gnd.n855 585
R3767 gnd.n6647 gnd.n6646 585
R3768 gnd.n6646 gnd.n6645 585
R3769 gnd.n6589 gnd.n6588 585
R3770 gnd.n6589 gnd.n864 585
R3771 gnd.n6635 gnd.n6596 585
R3772 gnd.n6596 gnd.n862 585
R3773 gnd.n6637 gnd.n6636 585
R3774 gnd.n6638 gnd.n6637 585
R3775 gnd.n6634 gnd.n6595 585
R3776 gnd.n6595 gnd.n6594 585
R3777 gnd.n6633 gnd.n6632 585
R3778 gnd.n6632 gnd.n870 585
R3779 gnd.n6631 gnd.n6597 585
R3780 gnd.n6631 gnd.n6630 585
R3781 gnd.n6616 gnd.n6598 585
R3782 gnd.n6599 gnd.n6598 585
R3783 gnd.n6617 gnd.n6610 585
R3784 gnd.n6610 gnd.n877 585
R3785 gnd.n6619 gnd.n6618 585
R3786 gnd.n6621 gnd.n6619 585
R3787 gnd.n6615 gnd.n6609 585
R3788 gnd.n6609 gnd.n6608 585
R3789 gnd.n6614 gnd.n6613 585
R3790 gnd.n6613 gnd.n884 585
R3791 gnd.n6612 gnd.n970 585
R3792 gnd.n6858 gnd.n970 585
R3793 gnd.n6611 gnd.n969 585
R3794 gnd.n6859 gnd.n969 585
R3795 gnd.n960 gnd.n959 585
R3796 gnd.n960 gnd.n891 585
R3797 gnd.n6867 gnd.n6866 585
R3798 gnd.n6866 gnd.n6865 585
R3799 gnd.n6868 gnd.n955 585
R3800 gnd.n961 gnd.n955 585
R3801 gnd.n6870 gnd.n6869 585
R3802 gnd.n6871 gnd.n6870 585
R3803 gnd.n958 gnd.n953 585
R3804 gnd.n6873 gnd.n953 585
R3805 gnd.n957 gnd.n956 585
R3806 gnd.n956 gnd.n905 585
R3807 gnd.n945 gnd.n944 585
R3808 gnd.n948 gnd.n945 585
R3809 gnd.n6882 gnd.n6881 585
R3810 gnd.n6881 gnd.n6880 585
R3811 gnd.n6883 gnd.n942 585
R3812 gnd.n942 gnd.n912 585
R3813 gnd.n6885 gnd.n6884 585
R3814 gnd.n6886 gnd.n6885 585
R3815 gnd.n943 gnd.n940 585
R3816 gnd.n6888 gnd.n940 585
R3817 gnd.n933 gnd.n932 585
R3818 gnd.n933 gnd.n919 585
R3819 gnd.n6896 gnd.n6895 585
R3820 gnd.n6895 gnd.n6894 585
R3821 gnd.n6897 gnd.n930 585
R3822 gnd.n930 gnd.n927 585
R3823 gnd.n6899 gnd.n6898 585
R3824 gnd.n6900 gnd.n6899 585
R3825 gnd.n931 gnd.n929 585
R3826 gnd.n6448 gnd.n929 585
R3827 gnd.n6437 gnd.n1008 585
R3828 gnd.n1008 gnd.n1003 585
R3829 gnd.n6439 gnd.n6438 585
R3830 gnd.n6441 gnd.n6439 585
R3831 gnd.n6436 gnd.n1007 585
R3832 gnd.n1007 gnd.n985 585
R3833 gnd.n6435 gnd.n6434 585
R3834 gnd.n6434 gnd.n984 585
R3835 gnd.n6433 gnd.n1009 585
R3836 gnd.n6433 gnd.n6432 585
R3837 gnd.n6388 gnd.n1010 585
R3838 gnd.n1010 gnd.n995 585
R3839 gnd.n6390 gnd.n6389 585
R3840 gnd.n6389 gnd.n993 585
R3841 gnd.n6391 gnd.n1016 585
R3842 gnd.n6424 gnd.n1016 585
R3843 gnd.n6393 gnd.n6392 585
R3844 gnd.n6394 gnd.n6393 585
R3845 gnd.n6387 gnd.n1041 585
R3846 gnd.n1041 gnd.n1024 585
R3847 gnd.n6386 gnd.n6385 585
R3848 gnd.n6385 gnd.n1023 585
R3849 gnd.n6384 gnd.n1042 585
R3850 gnd.n6384 gnd.n6383 585
R3851 gnd.n6368 gnd.n1043 585
R3852 gnd.n1043 gnd.n1034 585
R3853 gnd.n6369 gnd.n1051 585
R3854 gnd.n1051 gnd.n1032 585
R3855 gnd.n6371 gnd.n6370 585
R3856 gnd.n6372 gnd.n6371 585
R3857 gnd.n6367 gnd.n1050 585
R3858 gnd.n1054 gnd.n1050 585
R3859 gnd.n6366 gnd.n6365 585
R3860 gnd.n6365 gnd.n6364 585
R3861 gnd.n1053 gnd.n1052 585
R3862 gnd.n1062 gnd.n1053 585
R3863 gnd.n5946 gnd.n1060 585
R3864 gnd.n6357 gnd.n1060 585
R3865 gnd.n5949 gnd.n5947 585
R3866 gnd.n5949 gnd.n5948 585
R3867 gnd.n5951 gnd.n5950 585
R3868 gnd.n5950 gnd.n1071 585
R3869 gnd.n5952 gnd.n5801 585
R3870 gnd.n5969 gnd.n5801 585
R3871 gnd.n5954 gnd.n5953 585
R3872 gnd.n5953 gnd.n5800 585
R3873 gnd.n5955 gnd.n1082 585
R3874 gnd.n6332 gnd.n1082 585
R3875 gnd.n5956 gnd.n5807 585
R3876 gnd.n5807 gnd.n1079 585
R3877 gnd.n5958 gnd.n5957 585
R3878 gnd.n5960 gnd.n5958 585
R3879 gnd.n5945 gnd.n5806 585
R3880 gnd.n5806 gnd.n1088 585
R3881 gnd.n5944 gnd.n5943 585
R3882 gnd.n5943 gnd.n5942 585
R3883 gnd.n5809 gnd.n5808 585
R3884 gnd.n5811 gnd.n5809 585
R3885 gnd.n5931 gnd.n5818 585
R3886 gnd.n5818 gnd.n1095 585
R3887 gnd.n5933 gnd.n5932 585
R3888 gnd.n5934 gnd.n5933 585
R3889 gnd.n5930 gnd.n5817 585
R3890 gnd.n5817 gnd.n5816 585
R3891 gnd.n5929 gnd.n5928 585
R3892 gnd.n5928 gnd.n1102 585
R3893 gnd.n5927 gnd.n5819 585
R3894 gnd.n5927 gnd.n5926 585
R3895 gnd.n5915 gnd.n5820 585
R3896 gnd.n5822 gnd.n5820 585
R3897 gnd.n5917 gnd.n5916 585
R3898 gnd.n5918 gnd.n5917 585
R3899 gnd.n5914 gnd.n5829 585
R3900 gnd.n5829 gnd.n5828 585
R3901 gnd.n5913 gnd.n5912 585
R3902 gnd.n5912 gnd.n1116 585
R3903 gnd.n5911 gnd.n5830 585
R3904 gnd.n5911 gnd.n5910 585
R3905 gnd.n5898 gnd.n5831 585
R3906 gnd.n5833 gnd.n5831 585
R3907 gnd.n5899 gnd.n5841 585
R3908 gnd.n5841 gnd.n1123 585
R3909 gnd.n5901 gnd.n5900 585
R3910 gnd.n5902 gnd.n5901 585
R3911 gnd.n5897 gnd.n5840 585
R3912 gnd.n5840 gnd.n5839 585
R3913 gnd.n5896 gnd.n5895 585
R3914 gnd.n5895 gnd.n1130 585
R3915 gnd.n5894 gnd.n5842 585
R3916 gnd.n5894 gnd.n5893 585
R3917 gnd.n5880 gnd.n5843 585
R3918 gnd.n5845 gnd.n5843 585
R3919 gnd.n5881 gnd.n5852 585
R3920 gnd.n5852 gnd.n1137 585
R3921 gnd.n5883 gnd.n5882 585
R3922 gnd.n5884 gnd.n5883 585
R3923 gnd.n5879 gnd.n5851 585
R3924 gnd.n5851 gnd.n5850 585
R3925 gnd.n5878 gnd.n5877 585
R3926 gnd.n5877 gnd.n1145 585
R3927 gnd.n5876 gnd.n5853 585
R3928 gnd.n5876 gnd.n1143 585
R3929 gnd.n5875 gnd.n5862 585
R3930 gnd.n5875 gnd.n5874 585
R3931 gnd.n5861 gnd.n5854 585
R3932 gnd.n5854 gnd.n1153 585
R3933 gnd.n5860 gnd.n5859 585
R3934 gnd.n5859 gnd.n1151 585
R3935 gnd.n5858 gnd.n1434 585
R3936 gnd.n6023 gnd.n1434 585
R3937 gnd.n5857 gnd.n5856 585
R3938 gnd.n5856 gnd.n1160 585
R3939 gnd.n5855 gnd.n1322 585
R3940 gnd.n1326 gnd.n1322 585
R3941 gnd.n6031 gnd.n1323 585
R3942 gnd.n6031 gnd.n6030 585
R3943 gnd.n6032 gnd.n1321 585
R3944 gnd.n6032 gnd.n1167 585
R3945 gnd.n6151 gnd.n6150 585
R3946 gnd.n6152 gnd.n6151 585
R3947 gnd.n1249 gnd.n1247 585
R3948 gnd.n5603 gnd.n1247 585
R3949 gnd.n5592 gnd.n1606 585
R3950 gnd.n5563 gnd.n1606 585
R3951 gnd.n5594 gnd.n5593 585
R3952 gnd.n5595 gnd.n5594 585
R3953 gnd.n1607 gnd.n1605 585
R3954 gnd.n5561 gnd.n1605 585
R3955 gnd.n5587 gnd.n5586 585
R3956 gnd.n5586 gnd.n5585 585
R3957 gnd.n1610 gnd.n1609 585
R3958 gnd.n5577 gnd.n1610 585
R3959 gnd.n5552 gnd.n1632 585
R3960 gnd.n5538 gnd.n1632 585
R3961 gnd.n5554 gnd.n5553 585
R3962 gnd.n5555 gnd.n5554 585
R3963 gnd.n1633 gnd.n1631 585
R3964 gnd.n1680 gnd.n1631 585
R3965 gnd.n5547 gnd.n5546 585
R3966 gnd.n5546 gnd.n5545 585
R3967 gnd.n1636 gnd.n1635 585
R3968 gnd.n5468 gnd.n1636 585
R3969 gnd.n5484 gnd.n5483 585
R3970 gnd.n5485 gnd.n5484 585
R3971 gnd.n1664 gnd.n1663 585
R3972 gnd.n1663 gnd.n1658 585
R3973 gnd.n5479 gnd.n5478 585
R3974 gnd.n5478 gnd.n5477 585
R3975 gnd.n1667 gnd.n1666 585
R3976 gnd.n1714 gnd.n1667 585
R3977 gnd.n5449 gnd.n1697 585
R3978 gnd.n5435 gnd.n1697 585
R3979 gnd.n5451 gnd.n5450 585
R3980 gnd.n5452 gnd.n5451 585
R3981 gnd.n1698 gnd.n1696 585
R3982 gnd.n5423 gnd.n1696 585
R3983 gnd.n5444 gnd.n5443 585
R3984 gnd.n5443 gnd.n5442 585
R3985 gnd.n1701 gnd.n1700 585
R3986 gnd.n5411 gnd.n1701 585
R3987 gnd.n5399 gnd.n1735 585
R3988 gnd.n5385 gnd.n1735 585
R3989 gnd.n5401 gnd.n5400 585
R3990 gnd.n5402 gnd.n5401 585
R3991 gnd.n1736 gnd.n1734 585
R3992 gnd.n5373 gnd.n1734 585
R3993 gnd.n5394 gnd.n5393 585
R3994 gnd.n5393 gnd.n5392 585
R3995 gnd.n1739 gnd.n1738 585
R3996 gnd.n5366 gnd.n1739 585
R3997 gnd.n5354 gnd.n1771 585
R3998 gnd.n3605 gnd.n1771 585
R3999 gnd.n5356 gnd.n5355 585
R4000 gnd.n5357 gnd.n5356 585
R4001 gnd.n1772 gnd.n1770 585
R4002 gnd.n1770 gnd.n1766 585
R4003 gnd.n5326 gnd.n5325 585
R4004 gnd.n5327 gnd.n5326 585
R4005 gnd.n5324 gnd.n1796 585
R4006 gnd.n1805 gnd.n1796 585
R4007 gnd.n5335 gnd.n5334 585
R4008 gnd.n5334 gnd.n5333 585
R4009 gnd.n5337 gnd.n5336 585
R4010 gnd.n5337 gnd.n1795 585
R4011 gnd.n5340 gnd.n5339 585
R4012 gnd.n5341 gnd.n5340 585
R4013 gnd.n5338 gnd.n1781 585
R4014 gnd.n1784 gnd.n1781 585
R4015 gnd.n5349 gnd.n5348 585
R4016 gnd.n5348 gnd.n5347 585
R4017 gnd.n5350 gnd.n1780 585
R4018 gnd.n3548 gnd.n1780 585
R4019 gnd.n3396 gnd.n1779 585
R4020 gnd.n3629 gnd.n3396 585
R4021 gnd.n3634 gnd.n3631 585
R4022 gnd.n3631 gnd.n3630 585
R4023 gnd.n3636 gnd.n3635 585
R4024 gnd.n3637 gnd.n3636 585
R4025 gnd.n3384 gnd.n3383 585
R4026 gnd.n3387 gnd.n3384 585
R4027 gnd.n3645 gnd.n3644 585
R4028 gnd.n3644 gnd.n3643 585
R4029 gnd.n3646 gnd.n3378 585
R4030 gnd.n3378 gnd.n3377 585
R4031 gnd.n3648 gnd.n3647 585
R4032 gnd.n3649 gnd.n3648 585
R4033 gnd.n3364 gnd.n3363 585
R4034 gnd.n3368 gnd.n3364 585
R4035 gnd.n3657 gnd.n3656 585
R4036 gnd.n3656 gnd.n3655 585
R4037 gnd.n3658 gnd.n3358 585
R4038 gnd.n3365 gnd.n3358 585
R4039 gnd.n3660 gnd.n3659 585
R4040 gnd.n3661 gnd.n3660 585
R4041 gnd.n3346 gnd.n3345 585
R4042 gnd.n3349 gnd.n3346 585
R4043 gnd.n3669 gnd.n3668 585
R4044 gnd.n3668 gnd.n3667 585
R4045 gnd.n3670 gnd.n3340 585
R4046 gnd.n3340 gnd.n3339 585
R4047 gnd.n3672 gnd.n3671 585
R4048 gnd.n3673 gnd.n3672 585
R4049 gnd.n3326 gnd.n3325 585
R4050 gnd.n3330 gnd.n3326 585
R4051 gnd.n3681 gnd.n3680 585
R4052 gnd.n3680 gnd.n3679 585
R4053 gnd.n3682 gnd.n3320 585
R4054 gnd.n3327 gnd.n3320 585
R4055 gnd.n3684 gnd.n3683 585
R4056 gnd.n3685 gnd.n3684 585
R4057 gnd.n3308 gnd.n3307 585
R4058 gnd.n3311 gnd.n3308 585
R4059 gnd.n3693 gnd.n3692 585
R4060 gnd.n3692 gnd.n3691 585
R4061 gnd.n3694 gnd.n3302 585
R4062 gnd.n3302 gnd.n3301 585
R4063 gnd.n3696 gnd.n3695 585
R4064 gnd.n3697 gnd.n3696 585
R4065 gnd.n3285 gnd.n3284 585
R4066 gnd.n3289 gnd.n3285 585
R4067 gnd.n3705 gnd.n3704 585
R4068 gnd.n3704 gnd.n3703 585
R4069 gnd.n3706 gnd.n3278 585
R4070 gnd.n3286 gnd.n3278 585
R4071 gnd.n3708 gnd.n3707 585
R4072 gnd.n3709 gnd.n3708 585
R4073 gnd.n3279 gnd.n3205 585
R4074 gnd.n3205 gnd.n3202 585
R4075 gnd.n3831 gnd.n3830 585
R4076 gnd.n3829 gnd.n3204 585
R4077 gnd.n3828 gnd.n3203 585
R4078 gnd.n3833 gnd.n3203 585
R4079 gnd.n3827 gnd.n3826 585
R4080 gnd.n3825 gnd.n3824 585
R4081 gnd.n3823 gnd.n3822 585
R4082 gnd.n3821 gnd.n3820 585
R4083 gnd.n3819 gnd.n3818 585
R4084 gnd.n3817 gnd.n3816 585
R4085 gnd.n3815 gnd.n3814 585
R4086 gnd.n3813 gnd.n3812 585
R4087 gnd.n3811 gnd.n3810 585
R4088 gnd.n3809 gnd.n3808 585
R4089 gnd.n3807 gnd.n3806 585
R4090 gnd.n3805 gnd.n3804 585
R4091 gnd.n3803 gnd.n3802 585
R4092 gnd.n3801 gnd.n3800 585
R4093 gnd.n3799 gnd.n3798 585
R4094 gnd.n3796 gnd.n3795 585
R4095 gnd.n3794 gnd.n3793 585
R4096 gnd.n3792 gnd.n3791 585
R4097 gnd.n3790 gnd.n3789 585
R4098 gnd.n3788 gnd.n3787 585
R4099 gnd.n3786 gnd.n3785 585
R4100 gnd.n3784 gnd.n3783 585
R4101 gnd.n3782 gnd.n3781 585
R4102 gnd.n3780 gnd.n3779 585
R4103 gnd.n3778 gnd.n3777 585
R4104 gnd.n3776 gnd.n3775 585
R4105 gnd.n3774 gnd.n3773 585
R4106 gnd.n3772 gnd.n3771 585
R4107 gnd.n3770 gnd.n3769 585
R4108 gnd.n3768 gnd.n3767 585
R4109 gnd.n3766 gnd.n3765 585
R4110 gnd.n3764 gnd.n3763 585
R4111 gnd.n3762 gnd.n3761 585
R4112 gnd.n3760 gnd.n3759 585
R4113 gnd.n3758 gnd.n3757 585
R4114 gnd.n3756 gnd.n3755 585
R4115 gnd.n3754 gnd.n3753 585
R4116 gnd.n3752 gnd.n3751 585
R4117 gnd.n3750 gnd.n3749 585
R4118 gnd.n3748 gnd.n3747 585
R4119 gnd.n3746 gnd.n3745 585
R4120 gnd.n3744 gnd.n3743 585
R4121 gnd.n3742 gnd.n3741 585
R4122 gnd.n3740 gnd.n3739 585
R4123 gnd.n3738 gnd.n3737 585
R4124 gnd.n3736 gnd.n3735 585
R4125 gnd.n3734 gnd.n3733 585
R4126 gnd.n3732 gnd.n3731 585
R4127 gnd.n3730 gnd.n3729 585
R4128 gnd.n3728 gnd.n3727 585
R4129 gnd.n3726 gnd.n3725 585
R4130 gnd.n3724 gnd.n3723 585
R4131 gnd.n3722 gnd.n3721 585
R4132 gnd.n3720 gnd.n3719 585
R4133 gnd.n3718 gnd.n3717 585
R4134 gnd.n3274 gnd.n3267 585
R4135 gnd.n1589 gnd.n1588 585
R4136 gnd.n1586 gnd.n1482 585
R4137 gnd.n1585 gnd.n1584 585
R4138 gnd.n1578 gnd.n1484 585
R4139 gnd.n1580 gnd.n1579 585
R4140 gnd.n1576 gnd.n1486 585
R4141 gnd.n1575 gnd.n1574 585
R4142 gnd.n1568 gnd.n1488 585
R4143 gnd.n1570 gnd.n1569 585
R4144 gnd.n1566 gnd.n1490 585
R4145 gnd.n1565 gnd.n1564 585
R4146 gnd.n1558 gnd.n1492 585
R4147 gnd.n1560 gnd.n1559 585
R4148 gnd.n1556 gnd.n1494 585
R4149 gnd.n1555 gnd.n1554 585
R4150 gnd.n1548 gnd.n1496 585
R4151 gnd.n1550 gnd.n1549 585
R4152 gnd.n1546 gnd.n1498 585
R4153 gnd.n1545 gnd.n1544 585
R4154 gnd.n1538 gnd.n1500 585
R4155 gnd.n1540 gnd.n1539 585
R4156 gnd.n1536 gnd.n1504 585
R4157 gnd.n1535 gnd.n1534 585
R4158 gnd.n1528 gnd.n1506 585
R4159 gnd.n1530 gnd.n1529 585
R4160 gnd.n1526 gnd.n1508 585
R4161 gnd.n1525 gnd.n1524 585
R4162 gnd.n1518 gnd.n1510 585
R4163 gnd.n1520 gnd.n1519 585
R4164 gnd.n1516 gnd.n1513 585
R4165 gnd.n1515 gnd.n1297 585
R4166 gnd.n6102 gnd.n1293 585
R4167 gnd.n6104 gnd.n6103 585
R4168 gnd.n6106 gnd.n1291 585
R4169 gnd.n6108 gnd.n6107 585
R4170 gnd.n6109 gnd.n1286 585
R4171 gnd.n6111 gnd.n6110 585
R4172 gnd.n6113 gnd.n1284 585
R4173 gnd.n6115 gnd.n6114 585
R4174 gnd.n6117 gnd.n1277 585
R4175 gnd.n6119 gnd.n6118 585
R4176 gnd.n6121 gnd.n1275 585
R4177 gnd.n6123 gnd.n6122 585
R4178 gnd.n6124 gnd.n1270 585
R4179 gnd.n6126 gnd.n6125 585
R4180 gnd.n6128 gnd.n1268 585
R4181 gnd.n6130 gnd.n6129 585
R4182 gnd.n6131 gnd.n1263 585
R4183 gnd.n6133 gnd.n6132 585
R4184 gnd.n6135 gnd.n1261 585
R4185 gnd.n6137 gnd.n6136 585
R4186 gnd.n6138 gnd.n1255 585
R4187 gnd.n6140 gnd.n6139 585
R4188 gnd.n6142 gnd.n1254 585
R4189 gnd.n6143 gnd.n1252 585
R4190 gnd.n6146 gnd.n6145 585
R4191 gnd.n6147 gnd.n1248 585
R4192 gnd.n1253 gnd.n1248 585
R4193 gnd.n5606 gnd.n1244 585
R4194 gnd.n6152 gnd.n1244 585
R4195 gnd.n5605 gnd.n5604 585
R4196 gnd.n5604 gnd.n5603 585
R4197 gnd.n1594 gnd.n1593 585
R4198 gnd.n5563 gnd.n1594 585
R4199 gnd.n5597 gnd.n5596 585
R4200 gnd.n5596 gnd.n5595 585
R4201 gnd.n1600 gnd.n1599 585
R4202 gnd.n5561 gnd.n1600 585
R4203 gnd.n5580 gnd.n1612 585
R4204 gnd.n5585 gnd.n1612 585
R4205 gnd.n5579 gnd.n5578 585
R4206 gnd.n5578 gnd.n5577 585
R4207 gnd.n1620 gnd.n1619 585
R4208 gnd.n5538 gnd.n1620 585
R4209 gnd.n1679 gnd.n1628 585
R4210 gnd.n5555 gnd.n1628 585
R4211 gnd.n1682 gnd.n1681 585
R4212 gnd.n1681 gnd.n1680 585
R4213 gnd.n1683 gnd.n1638 585
R4214 gnd.n5545 gnd.n1638 585
R4215 gnd.n5470 gnd.n5469 585
R4216 gnd.n5469 gnd.n5468 585
R4217 gnd.n5471 gnd.n1659 585
R4218 gnd.n5485 gnd.n1659 585
R4219 gnd.n1678 gnd.n1677 585
R4220 gnd.n1677 gnd.n1658 585
R4221 gnd.n5416 gnd.n1668 585
R4222 gnd.n5477 gnd.n1668 585
R4223 gnd.n5418 gnd.n5417 585
R4224 gnd.n5417 gnd.n1714 585
R4225 gnd.n5419 gnd.n1713 585
R4226 gnd.n5435 gnd.n1713 585
R4227 gnd.n5420 gnd.n1693 585
R4228 gnd.n5452 gnd.n1693 585
R4229 gnd.n5422 gnd.n5421 585
R4230 gnd.n5423 gnd.n5422 585
R4231 gnd.n5414 gnd.n1703 585
R4232 gnd.n5442 gnd.n1703 585
R4233 gnd.n5413 gnd.n5412 585
R4234 gnd.n5412 gnd.n5411 585
R4235 gnd.n1724 gnd.n1722 585
R4236 gnd.n5385 gnd.n1724 585
R4237 gnd.n5370 gnd.n1731 585
R4238 gnd.n5402 gnd.n1731 585
R4239 gnd.n5372 gnd.n5371 585
R4240 gnd.n5373 gnd.n5372 585
R4241 gnd.n5369 gnd.n1741 585
R4242 gnd.n5392 gnd.n1741 585
R4243 gnd.n5368 gnd.n5367 585
R4244 gnd.n5367 gnd.n5366 585
R4245 gnd.n1759 gnd.n1757 585
R4246 gnd.n3605 gnd.n1759 585
R4247 gnd.n3610 gnd.n1767 585
R4248 gnd.n5357 gnd.n1767 585
R4249 gnd.n3612 gnd.n3611 585
R4250 gnd.n3611 gnd.n1766 585
R4251 gnd.n3613 gnd.n1806 585
R4252 gnd.n5327 gnd.n1806 585
R4253 gnd.n3615 gnd.n3614 585
R4254 gnd.n3614 gnd.n1805 585
R4255 gnd.n3616 gnd.n1797 585
R4256 gnd.n5333 gnd.n1797 585
R4257 gnd.n3618 gnd.n3617 585
R4258 gnd.n3617 gnd.n1795 585
R4259 gnd.n3619 gnd.n1793 585
R4260 gnd.n5341 gnd.n1793 585
R4261 gnd.n3621 gnd.n3620 585
R4262 gnd.n3620 gnd.n1784 585
R4263 gnd.n3622 gnd.n1782 585
R4264 gnd.n5347 gnd.n1782 585
R4265 gnd.n3624 gnd.n3623 585
R4266 gnd.n3623 gnd.n3548 585
R4267 gnd.n3625 gnd.n3399 585
R4268 gnd.n3629 gnd.n3399 585
R4269 gnd.n3592 gnd.n3397 585
R4270 gnd.n3630 gnd.n3397 585
R4271 gnd.n3591 gnd.n3394 585
R4272 gnd.n3637 gnd.n3394 585
R4273 gnd.n3590 gnd.n3589 585
R4274 gnd.n3589 gnd.n3387 585
R4275 gnd.n3588 gnd.n3385 585
R4276 gnd.n3643 gnd.n3385 585
R4277 gnd.n3587 gnd.n3586 585
R4278 gnd.n3586 gnd.n3377 585
R4279 gnd.n3584 gnd.n3375 585
R4280 gnd.n3649 gnd.n3375 585
R4281 gnd.n3583 gnd.n3582 585
R4282 gnd.n3582 gnd.n3368 585
R4283 gnd.n3581 gnd.n3366 585
R4284 gnd.n3655 gnd.n3366 585
R4285 gnd.n3580 gnd.n3579 585
R4286 gnd.n3579 gnd.n3365 585
R4287 gnd.n3577 gnd.n3356 585
R4288 gnd.n3661 gnd.n3356 585
R4289 gnd.n3576 gnd.n3575 585
R4290 gnd.n3575 gnd.n3349 585
R4291 gnd.n3574 gnd.n3347 585
R4292 gnd.n3667 gnd.n3347 585
R4293 gnd.n3573 gnd.n3572 585
R4294 gnd.n3572 gnd.n3339 585
R4295 gnd.n3570 gnd.n3337 585
R4296 gnd.n3673 gnd.n3337 585
R4297 gnd.n3569 gnd.n3568 585
R4298 gnd.n3568 gnd.n3330 585
R4299 gnd.n3567 gnd.n3328 585
R4300 gnd.n3679 gnd.n3328 585
R4301 gnd.n3566 gnd.n3565 585
R4302 gnd.n3565 gnd.n3327 585
R4303 gnd.n3563 gnd.n3318 585
R4304 gnd.n3685 gnd.n3318 585
R4305 gnd.n3562 gnd.n3561 585
R4306 gnd.n3561 gnd.n3311 585
R4307 gnd.n3560 gnd.n3309 585
R4308 gnd.n3691 gnd.n3309 585
R4309 gnd.n3559 gnd.n3558 585
R4310 gnd.n3558 gnd.n3301 585
R4311 gnd.n3556 gnd.n3299 585
R4312 gnd.n3697 gnd.n3299 585
R4313 gnd.n3555 gnd.n3554 585
R4314 gnd.n3554 gnd.n3289 585
R4315 gnd.n3553 gnd.n3287 585
R4316 gnd.n3703 gnd.n3287 585
R4317 gnd.n3552 gnd.n3275 585
R4318 gnd.n3286 gnd.n3275 585
R4319 gnd.n3710 gnd.n3273 585
R4320 gnd.n3710 gnd.n3709 585
R4321 gnd.n3712 gnd.n3711 585
R4322 gnd.n3711 gnd.n3202 585
R4323 gnd.n7888 gnd.n249 585
R4324 gnd.n249 gnd.n248 585
R4325 gnd.n7890 gnd.n7889 585
R4326 gnd.n7891 gnd.n7890 585
R4327 gnd.n236 gnd.n235 585
R4328 gnd.n239 gnd.n236 585
R4329 gnd.n7899 gnd.n7898 585
R4330 gnd.n7898 gnd.n7897 585
R4331 gnd.n7900 gnd.n230 585
R4332 gnd.n230 gnd.n229 585
R4333 gnd.n7902 gnd.n7901 585
R4334 gnd.n7903 gnd.n7902 585
R4335 gnd.n217 gnd.n216 585
R4336 gnd.n226 gnd.n217 585
R4337 gnd.n7911 gnd.n7910 585
R4338 gnd.n7910 gnd.n7909 585
R4339 gnd.n7912 gnd.n211 585
R4340 gnd.n211 gnd.n210 585
R4341 gnd.n7914 gnd.n7913 585
R4342 gnd.n7915 gnd.n7914 585
R4343 gnd.n197 gnd.n196 585
R4344 gnd.n7741 gnd.n197 585
R4345 gnd.n7923 gnd.n7922 585
R4346 gnd.n7922 gnd.n7921 585
R4347 gnd.n7924 gnd.n191 585
R4348 gnd.n198 gnd.n191 585
R4349 gnd.n7926 gnd.n7925 585
R4350 gnd.n7927 gnd.n7926 585
R4351 gnd.n179 gnd.n178 585
R4352 gnd.n188 gnd.n179 585
R4353 gnd.n7935 gnd.n7934 585
R4354 gnd.n7934 gnd.n7933 585
R4355 gnd.n7936 gnd.n173 585
R4356 gnd.n173 gnd.n172 585
R4357 gnd.n7938 gnd.n7937 585
R4358 gnd.n7939 gnd.n7938 585
R4359 gnd.n159 gnd.n158 585
R4360 gnd.n163 gnd.n159 585
R4361 gnd.n7947 gnd.n7946 585
R4362 gnd.n7946 gnd.n7945 585
R4363 gnd.n7948 gnd.n153 585
R4364 gnd.n160 gnd.n153 585
R4365 gnd.n7950 gnd.n7949 585
R4366 gnd.n7951 gnd.n7950 585
R4367 gnd.n141 gnd.n140 585
R4368 gnd.n150 gnd.n141 585
R4369 gnd.n7959 gnd.n7958 585
R4370 gnd.n7958 gnd.n7957 585
R4371 gnd.n7960 gnd.n136 585
R4372 gnd.n136 gnd.n135 585
R4373 gnd.n7962 gnd.n7961 585
R4374 gnd.n7963 gnd.n7962 585
R4375 gnd.n120 gnd.n118 585
R4376 gnd.n124 gnd.n120 585
R4377 gnd.n7971 gnd.n7970 585
R4378 gnd.n7970 gnd.n7969 585
R4379 gnd.n119 gnd.n111 585
R4380 gnd.n121 gnd.n119 585
R4381 gnd.n7974 gnd.n109 585
R4382 gnd.n109 gnd.n106 585
R4383 gnd.n7976 gnd.n7975 585
R4384 gnd.n7977 gnd.n7976 585
R4385 gnd.n7555 gnd.n108 585
R4386 gnd.n7570 gnd.n108 585
R4387 gnd.n7557 gnd.n7556 585
R4388 gnd.n7557 gnd.n358 585
R4389 gnd.n7560 gnd.n7559 585
R4390 gnd.n7561 gnd.n7560 585
R4391 gnd.n7558 gnd.n7554 585
R4392 gnd.n7554 gnd.n7553 585
R4393 gnd.n7542 gnd.n367 585
R4394 gnd.n368 gnd.n367 585
R4395 gnd.n7544 gnd.n7543 585
R4396 gnd.n7545 gnd.n7544 585
R4397 gnd.n7541 gnd.n7540 585
R4398 gnd.n7541 gnd.n376 585
R4399 gnd.n7539 gnd.n379 585
R4400 gnd.n7519 gnd.n379 585
R4401 gnd.n7538 gnd.n7537 585
R4402 gnd.n7537 gnd.n7536 585
R4403 gnd.n382 gnd.n380 585
R4404 gnd.n7508 gnd.n382 585
R4405 gnd.n7494 gnd.n416 585
R4406 gnd.n416 gnd.n403 585
R4407 gnd.n7496 gnd.n7495 585
R4408 gnd.n7497 gnd.n7496 585
R4409 gnd.n417 gnd.n415 585
R4410 gnd.n7471 gnd.n415 585
R4411 gnd.n7488 gnd.n7487 585
R4412 gnd.n7487 gnd.n7486 585
R4413 gnd.n420 gnd.n419 585
R4414 gnd.n7457 gnd.n420 585
R4415 gnd.n7445 gnd.n451 585
R4416 gnd.n451 gnd.n438 585
R4417 gnd.n7447 gnd.n7446 585
R4418 gnd.n7448 gnd.n7447 585
R4419 gnd.n452 gnd.n450 585
R4420 gnd.n7424 gnd.n450 585
R4421 gnd.n7440 gnd.n7439 585
R4422 gnd.n7439 gnd.n7438 585
R4423 gnd.n455 gnd.n454 585
R4424 gnd.n7420 gnd.n455 585
R4425 gnd.n7408 gnd.n481 585
R4426 gnd.n7394 gnd.n481 585
R4427 gnd.n7410 gnd.n7409 585
R4428 gnd.n7411 gnd.n7410 585
R4429 gnd.n482 gnd.n480 585
R4430 gnd.n7338 gnd.n480 585
R4431 gnd.n7403 gnd.n7402 585
R4432 gnd.n7402 gnd.n7401 585
R4433 gnd.n485 gnd.n484 585
R4434 gnd.n7371 gnd.n485 585
R4435 gnd.n7359 gnd.n517 585
R4436 gnd.n517 gnd.n504 585
R4437 gnd.n7361 gnd.n7360 585
R4438 gnd.n7362 gnd.n7361 585
R4439 gnd.n518 gnd.n516 585
R4440 gnd.n7333 gnd.n516 585
R4441 gnd.n7354 gnd.n7353 585
R4442 gnd.n7353 gnd.n7352 585
R4443 gnd.n521 gnd.n520 585
R4444 gnd.n7329 gnd.n521 585
R4445 gnd.n7317 gnd.n547 585
R4446 gnd.n559 gnd.n547 585
R4447 gnd.n7319 gnd.n7318 585
R4448 gnd.n7320 gnd.n7319 585
R4449 gnd.n548 gnd.n546 585
R4450 gnd.n7302 gnd.n546 585
R4451 gnd.n7312 gnd.n7311 585
R4452 gnd.n7311 gnd.n7310 585
R4453 gnd.n611 gnd.n550 585
R4454 gnd.n7272 gnd.n7271 585
R4455 gnd.n7270 gnd.n610 585
R4456 gnd.n7274 gnd.n610 585
R4457 gnd.n7269 gnd.n7268 585
R4458 gnd.n7267 gnd.n7266 585
R4459 gnd.n7265 gnd.n7264 585
R4460 gnd.n7263 gnd.n7262 585
R4461 gnd.n7261 gnd.n7260 585
R4462 gnd.n7259 gnd.n7258 585
R4463 gnd.n7257 gnd.n7256 585
R4464 gnd.n7255 gnd.n7254 585
R4465 gnd.n7253 gnd.n7252 585
R4466 gnd.n7251 gnd.n7250 585
R4467 gnd.n7249 gnd.n7248 585
R4468 gnd.n7247 gnd.n7246 585
R4469 gnd.n7245 gnd.n7244 585
R4470 gnd.n7243 gnd.n7242 585
R4471 gnd.n7241 gnd.n7240 585
R4472 gnd.n7238 gnd.n7237 585
R4473 gnd.n7236 gnd.n7235 585
R4474 gnd.n7234 gnd.n7233 585
R4475 gnd.n7232 gnd.n7231 585
R4476 gnd.n7230 gnd.n7229 585
R4477 gnd.n7228 gnd.n7227 585
R4478 gnd.n7226 gnd.n7225 585
R4479 gnd.n7224 gnd.n7223 585
R4480 gnd.n7221 gnd.n7220 585
R4481 gnd.n7219 gnd.n7218 585
R4482 gnd.n7217 gnd.n7216 585
R4483 gnd.n7215 gnd.n7214 585
R4484 gnd.n7213 gnd.n7212 585
R4485 gnd.n7211 gnd.n7210 585
R4486 gnd.n7209 gnd.n7208 585
R4487 gnd.n7207 gnd.n7206 585
R4488 gnd.n7205 gnd.n7204 585
R4489 gnd.n7203 gnd.n7202 585
R4490 gnd.n7201 gnd.n7200 585
R4491 gnd.n7199 gnd.n7198 585
R4492 gnd.n7197 gnd.n7196 585
R4493 gnd.n7195 gnd.n7194 585
R4494 gnd.n7193 gnd.n7192 585
R4495 gnd.n7191 gnd.n7190 585
R4496 gnd.n7189 gnd.n7188 585
R4497 gnd.n7187 gnd.n7186 585
R4498 gnd.n7185 gnd.n7184 585
R4499 gnd.n7183 gnd.n7182 585
R4500 gnd.n7181 gnd.n7180 585
R4501 gnd.n7179 gnd.n7178 585
R4502 gnd.n7177 gnd.n7176 585
R4503 gnd.n7175 gnd.n7174 585
R4504 gnd.n7173 gnd.n7172 585
R4505 gnd.n7171 gnd.n7170 585
R4506 gnd.n7169 gnd.n7168 585
R4507 gnd.n7167 gnd.n7166 585
R4508 gnd.n7165 gnd.n7164 585
R4509 gnd.n7163 gnd.n7162 585
R4510 gnd.n674 gnd.n673 585
R4511 gnd.n7759 gnd.n349 585
R4512 gnd.n7767 gnd.n7766 585
R4513 gnd.n7769 gnd.n7768 585
R4514 gnd.n7771 gnd.n7770 585
R4515 gnd.n7773 gnd.n7772 585
R4516 gnd.n7775 gnd.n7774 585
R4517 gnd.n7777 gnd.n7776 585
R4518 gnd.n7779 gnd.n7778 585
R4519 gnd.n7781 gnd.n7780 585
R4520 gnd.n7783 gnd.n7782 585
R4521 gnd.n7785 gnd.n7784 585
R4522 gnd.n7787 gnd.n7786 585
R4523 gnd.n7789 gnd.n7788 585
R4524 gnd.n7791 gnd.n7790 585
R4525 gnd.n7793 gnd.n7792 585
R4526 gnd.n7795 gnd.n7794 585
R4527 gnd.n7797 gnd.n7796 585
R4528 gnd.n7799 gnd.n7798 585
R4529 gnd.n7801 gnd.n7800 585
R4530 gnd.n7804 gnd.n7803 585
R4531 gnd.n7802 gnd.n329 585
R4532 gnd.n7809 gnd.n7808 585
R4533 gnd.n7811 gnd.n7810 585
R4534 gnd.n7813 gnd.n7812 585
R4535 gnd.n7815 gnd.n7814 585
R4536 gnd.n7817 gnd.n7816 585
R4537 gnd.n7819 gnd.n7818 585
R4538 gnd.n7821 gnd.n7820 585
R4539 gnd.n7823 gnd.n7822 585
R4540 gnd.n7825 gnd.n7824 585
R4541 gnd.n7827 gnd.n7826 585
R4542 gnd.n7829 gnd.n7828 585
R4543 gnd.n7831 gnd.n7830 585
R4544 gnd.n7833 gnd.n7832 585
R4545 gnd.n7835 gnd.n7834 585
R4546 gnd.n7837 gnd.n7836 585
R4547 gnd.n7839 gnd.n7838 585
R4548 gnd.n7841 gnd.n7840 585
R4549 gnd.n7843 gnd.n7842 585
R4550 gnd.n7845 gnd.n7844 585
R4551 gnd.n7847 gnd.n7846 585
R4552 gnd.n7852 gnd.n7851 585
R4553 gnd.n7854 gnd.n7853 585
R4554 gnd.n7856 gnd.n7855 585
R4555 gnd.n7858 gnd.n7857 585
R4556 gnd.n7860 gnd.n7859 585
R4557 gnd.n7862 gnd.n7861 585
R4558 gnd.n7864 gnd.n7863 585
R4559 gnd.n7866 gnd.n7865 585
R4560 gnd.n7868 gnd.n7867 585
R4561 gnd.n7870 gnd.n7869 585
R4562 gnd.n7872 gnd.n7871 585
R4563 gnd.n7874 gnd.n7873 585
R4564 gnd.n7876 gnd.n7875 585
R4565 gnd.n7878 gnd.n7877 585
R4566 gnd.n7879 gnd.n293 585
R4567 gnd.n7881 gnd.n7880 585
R4568 gnd.n254 gnd.n253 585
R4569 gnd.n7885 gnd.n7884 585
R4570 gnd.n7884 gnd.n7883 585
R4571 gnd.n7761 gnd.n7760 585
R4572 gnd.n7760 gnd.n248 585
R4573 gnd.n7758 gnd.n246 585
R4574 gnd.n7891 gnd.n246 585
R4575 gnd.n7757 gnd.n7756 585
R4576 gnd.n7756 gnd.n239 585
R4577 gnd.n7755 gnd.n237 585
R4578 gnd.n7897 gnd.n237 585
R4579 gnd.n7754 gnd.n7753 585
R4580 gnd.n7753 gnd.n229 585
R4581 gnd.n7751 gnd.n227 585
R4582 gnd.n7903 gnd.n227 585
R4583 gnd.n7750 gnd.n7749 585
R4584 gnd.n7749 gnd.n226 585
R4585 gnd.n7748 gnd.n218 585
R4586 gnd.n7909 gnd.n218 585
R4587 gnd.n7747 gnd.n7746 585
R4588 gnd.n7746 gnd.n210 585
R4589 gnd.n7744 gnd.n208 585
R4590 gnd.n7915 gnd.n208 585
R4591 gnd.n7743 gnd.n7742 585
R4592 gnd.n7742 gnd.n7741 585
R4593 gnd.n7609 gnd.n199 585
R4594 gnd.n7921 gnd.n199 585
R4595 gnd.n7608 gnd.n7607 585
R4596 gnd.n7607 gnd.n198 585
R4597 gnd.n7605 gnd.n189 585
R4598 gnd.n7927 gnd.n189 585
R4599 gnd.n7604 gnd.n7603 585
R4600 gnd.n7603 gnd.n188 585
R4601 gnd.n7602 gnd.n180 585
R4602 gnd.n7933 gnd.n180 585
R4603 gnd.n7601 gnd.n7600 585
R4604 gnd.n7600 gnd.n172 585
R4605 gnd.n7598 gnd.n170 585
R4606 gnd.n7939 gnd.n170 585
R4607 gnd.n7597 gnd.n7596 585
R4608 gnd.n7596 gnd.n163 585
R4609 gnd.n7595 gnd.n161 585
R4610 gnd.n7945 gnd.n161 585
R4611 gnd.n7594 gnd.n7593 585
R4612 gnd.n7593 gnd.n160 585
R4613 gnd.n7591 gnd.n151 585
R4614 gnd.n7951 gnd.n151 585
R4615 gnd.n7590 gnd.n7589 585
R4616 gnd.n7589 gnd.n150 585
R4617 gnd.n7588 gnd.n142 585
R4618 gnd.n7957 gnd.n142 585
R4619 gnd.n7587 gnd.n7586 585
R4620 gnd.n7586 gnd.n135 585
R4621 gnd.n7584 gnd.n133 585
R4622 gnd.n7963 gnd.n133 585
R4623 gnd.n7583 gnd.n7582 585
R4624 gnd.n7582 gnd.n124 585
R4625 gnd.n7581 gnd.n122 585
R4626 gnd.n7969 gnd.n122 585
R4627 gnd.n7580 gnd.n7579 585
R4628 gnd.n7579 gnd.n121 585
R4629 gnd.n7578 gnd.n353 585
R4630 gnd.n7578 gnd.n106 585
R4631 gnd.n7567 gnd.n105 585
R4632 gnd.n7977 gnd.n105 585
R4633 gnd.n7569 gnd.n7568 585
R4634 gnd.n7570 gnd.n7569 585
R4635 gnd.n7566 gnd.n359 585
R4636 gnd.n359 gnd.n358 585
R4637 gnd.n364 gnd.n360 585
R4638 gnd.n7561 gnd.n364 585
R4639 gnd.n7524 gnd.n369 585
R4640 gnd.n7553 gnd.n369 585
R4641 gnd.n7526 gnd.n7525 585
R4642 gnd.n7525 gnd.n368 585
R4643 gnd.n7523 gnd.n377 585
R4644 gnd.n7545 gnd.n377 585
R4645 gnd.n7522 gnd.n7521 585
R4646 gnd.n7521 gnd.n376 585
R4647 gnd.n7520 gnd.n393 585
R4648 gnd.n7520 gnd.n7519 585
R4649 gnd.n7475 gnd.n384 585
R4650 gnd.n7536 gnd.n384 585
R4651 gnd.n7476 gnd.n404 585
R4652 gnd.n7508 gnd.n404 585
R4653 gnd.n7478 gnd.n7477 585
R4654 gnd.n7477 gnd.n403 585
R4655 gnd.n7474 gnd.n412 585
R4656 gnd.n7497 gnd.n412 585
R4657 gnd.n7473 gnd.n7472 585
R4658 gnd.n7472 gnd.n7471 585
R4659 gnd.n431 gnd.n422 585
R4660 gnd.n7486 gnd.n422 585
R4661 gnd.n7428 gnd.n439 585
R4662 gnd.n7457 gnd.n439 585
R4663 gnd.n7430 gnd.n7429 585
R4664 gnd.n7429 gnd.n438 585
R4665 gnd.n7427 gnd.n447 585
R4666 gnd.n7448 gnd.n447 585
R4667 gnd.n7426 gnd.n7425 585
R4668 gnd.n7425 gnd.n7424 585
R4669 gnd.n7423 gnd.n457 585
R4670 gnd.n7438 gnd.n457 585
R4671 gnd.n7422 gnd.n7421 585
R4672 gnd.n7421 gnd.n7420 585
R4673 gnd.n469 gnd.n467 585
R4674 gnd.n7394 gnd.n469 585
R4675 gnd.n7337 gnd.n478 585
R4676 gnd.n7411 gnd.n478 585
R4677 gnd.n7340 gnd.n7339 585
R4678 gnd.n7339 gnd.n7338 585
R4679 gnd.n7341 gnd.n487 585
R4680 gnd.n7401 gnd.n487 585
R4681 gnd.n7342 gnd.n505 585
R4682 gnd.n7371 gnd.n505 585
R4683 gnd.n7344 gnd.n7343 585
R4684 gnd.n7343 gnd.n504 585
R4685 gnd.n7336 gnd.n513 585
R4686 gnd.n7362 gnd.n513 585
R4687 gnd.n7335 gnd.n7334 585
R4688 gnd.n7334 gnd.n7333 585
R4689 gnd.n7332 gnd.n523 585
R4690 gnd.n7352 gnd.n523 585
R4691 gnd.n7331 gnd.n7330 585
R4692 gnd.n7330 gnd.n7329 585
R4693 gnd.n535 gnd.n533 585
R4694 gnd.n559 gnd.n535 585
R4695 gnd.n7304 gnd.n543 585
R4696 gnd.n7320 gnd.n543 585
R4697 gnd.n7305 gnd.n7303 585
R4698 gnd.n7303 gnd.n7302 585
R4699 gnd.n564 gnd.n552 585
R4700 gnd.n7310 gnd.n552 585
R4701 gnd.n5322 gnd.n5321 585
R4702 gnd.n5323 gnd.n5322 585
R4703 gnd.n2436 gnd.n398 585
R4704 gnd.n398 gnd.n397 585
R4705 gnd.n7517 gnd.n7516 585
R4706 gnd.n7518 gnd.n7517 585
R4707 gnd.n399 gnd.n396 585
R4708 gnd.n396 gnd.n394 585
R4709 gnd.n7512 gnd.n7511 585
R4710 gnd.n7511 gnd.n383 585
R4711 gnd.n7510 gnd.n401 585
R4712 gnd.n7510 gnd.n7509 585
R4713 gnd.n7466 gnd.n402 585
R4714 gnd.n413 gnd.n402 585
R4715 gnd.n7467 gnd.n433 585
R4716 gnd.n433 gnd.n411 585
R4717 gnd.n7469 gnd.n7468 585
R4718 gnd.n7470 gnd.n7469 585
R4719 gnd.n434 gnd.n432 585
R4720 gnd.n432 gnd.n421 585
R4721 gnd.n7460 gnd.n7459 585
R4722 gnd.n7459 gnd.n7458 585
R4723 gnd.n437 gnd.n436 585
R4724 gnd.n448 gnd.n437 585
R4725 gnd.n7386 gnd.n7385 585
R4726 gnd.n7386 gnd.n446 585
R4727 gnd.n7387 gnd.n7382 585
R4728 gnd.n7387 gnd.n459 585
R4729 gnd.n7389 gnd.n7388 585
R4730 gnd.n7388 gnd.n456 585
R4731 gnd.n7390 gnd.n498 585
R4732 gnd.n498 gnd.n470 585
R4733 gnd.n7392 gnd.n7391 585
R4734 gnd.n7393 gnd.n7392 585
R4735 gnd.n499 gnd.n497 585
R4736 gnd.n497 gnd.n477 585
R4737 gnd.n7376 gnd.n7375 585
R4738 gnd.n7375 gnd.n489 585
R4739 gnd.n7374 gnd.n501 585
R4740 gnd.n7374 gnd.n486 585
R4741 gnd.n7373 gnd.n503 585
R4742 gnd.n7373 gnd.n7372 585
R4743 gnd.n7291 gnd.n502 585
R4744 gnd.n514 gnd.n502 585
R4745 gnd.n7292 gnd.n7285 585
R4746 gnd.n7285 gnd.n512 585
R4747 gnd.n7294 gnd.n7293 585
R4748 gnd.n7294 gnd.n525 585
R4749 gnd.n7295 gnd.n7284 585
R4750 gnd.n7295 gnd.n522 585
R4751 gnd.n7297 gnd.n7296 585
R4752 gnd.n7296 gnd.n536 585
R4753 gnd.n7298 gnd.n566 585
R4754 gnd.n566 gnd.n544 585
R4755 gnd.n7300 gnd.n7299 585
R4756 gnd.n7301 gnd.n7300 585
R4757 gnd.n567 gnd.n565 585
R4758 gnd.n565 gnd.n554 585
R4759 gnd.n7278 gnd.n7277 585
R4760 gnd.n7277 gnd.n551 585
R4761 gnd.n7276 gnd.n569 585
R4762 gnd.n7276 gnd.n7275 585
R4763 gnd.n7073 gnd.n570 585
R4764 gnd.n571 gnd.n570 585
R4765 gnd.n7074 gnd.n780 585
R4766 gnd.n780 gnd.n778 585
R4767 gnd.n7076 gnd.n7075 585
R4768 gnd.n7077 gnd.n7076 585
R4769 gnd.n781 gnd.n779 585
R4770 gnd.n779 gnd.n747 585
R4771 gnd.n7067 gnd.n746 585
R4772 gnd.n7094 gnd.n746 585
R4773 gnd.n7066 gnd.n7065 585
R4774 gnd.n7065 gnd.n745 585
R4775 gnd.n7064 gnd.n783 585
R4776 gnd.n7064 gnd.n7063 585
R4777 gnd.n7052 gnd.n784 585
R4778 gnd.n785 gnd.n784 585
R4779 gnd.n7054 gnd.n7053 585
R4780 gnd.n7055 gnd.n7054 585
R4781 gnd.n795 gnd.n794 585
R4782 gnd.n794 gnd.n792 585
R4783 gnd.n7046 gnd.n7045 585
R4784 gnd.n7045 gnd.n7044 585
R4785 gnd.n798 gnd.n797 585
R4786 gnd.n807 gnd.n798 585
R4787 gnd.n7035 gnd.n7034 585
R4788 gnd.n7036 gnd.n7035 585
R4789 gnd.n809 gnd.n808 585
R4790 gnd.n808 gnd.n805 585
R4791 gnd.n7030 gnd.n7029 585
R4792 gnd.n7029 gnd.n7028 585
R4793 gnd.n812 gnd.n811 585
R4794 gnd.n813 gnd.n812 585
R4795 gnd.n7019 gnd.n7018 585
R4796 gnd.n7020 gnd.n7019 585
R4797 gnd.n823 gnd.n822 585
R4798 gnd.n822 gnd.n820 585
R4799 gnd.n7014 gnd.n7013 585
R4800 gnd.n7013 gnd.n7012 585
R4801 gnd.n826 gnd.n825 585
R4802 gnd.n827 gnd.n826 585
R4803 gnd.n7003 gnd.n7002 585
R4804 gnd.n7004 gnd.n7003 585
R4805 gnd.n836 gnd.n835 585
R4806 gnd.n842 gnd.n835 585
R4807 gnd.n6998 gnd.n6997 585
R4808 gnd.n6997 gnd.n6996 585
R4809 gnd.n839 gnd.n838 585
R4810 gnd.n6792 gnd.n839 585
R4811 gnd.n6987 gnd.n6986 585
R4812 gnd.n6988 gnd.n6987 585
R4813 gnd.n851 gnd.n850 585
R4814 gnd.n6653 gnd.n850 585
R4815 gnd.n6982 gnd.n6981 585
R4816 gnd.n6981 gnd.n6980 585
R4817 gnd.n854 gnd.n853 585
R4818 gnd.n6590 gnd.n854 585
R4819 gnd.n6971 gnd.n6970 585
R4820 gnd.n6972 gnd.n6971 585
R4821 gnd.n866 gnd.n865 585
R4822 gnd.n6638 gnd.n865 585
R4823 gnd.n6966 gnd.n6965 585
R4824 gnd.n6965 gnd.n6964 585
R4825 gnd.n869 gnd.n868 585
R4826 gnd.n6600 gnd.n869 585
R4827 gnd.n6955 gnd.n6954 585
R4828 gnd.n6956 gnd.n6955 585
R4829 gnd.n880 gnd.n879 585
R4830 gnd.n6620 gnd.n879 585
R4831 gnd.n6950 gnd.n6949 585
R4832 gnd.n6949 gnd.n6948 585
R4833 gnd.n883 gnd.n882 585
R4834 gnd.n6857 gnd.n883 585
R4835 gnd.n6939 gnd.n6938 585
R4836 gnd.n6940 gnd.n6939 585
R4837 gnd.n894 gnd.n893 585
R4838 gnd.n962 gnd.n893 585
R4839 gnd.n6934 gnd.n6933 585
R4840 gnd.n6933 gnd.n6932 585
R4841 gnd.n897 gnd.n896 585
R4842 gnd.n6872 gnd.n897 585
R4843 gnd.n6923 gnd.n6922 585
R4844 gnd.n6924 gnd.n6923 585
R4845 gnd.n907 gnd.n906 585
R4846 gnd.n946 gnd.n906 585
R4847 gnd.n6918 gnd.n6917 585
R4848 gnd.n6917 gnd.n6916 585
R4849 gnd.n910 gnd.n909 585
R4850 gnd.n6887 gnd.n910 585
R4851 gnd.n6907 gnd.n6906 585
R4852 gnd.n6908 gnd.n6907 585
R4853 gnd.n921 gnd.n920 585
R4854 gnd.n934 gnd.n920 585
R4855 gnd.n6902 gnd.n6901 585
R4856 gnd.n6901 gnd.n6900 585
R4857 gnd.n924 gnd.n923 585
R4858 gnd.n6449 gnd.n924 585
R4859 gnd.n6469 gnd.n988 585
R4860 gnd.n6440 gnd.n988 585
R4861 gnd.n6471 gnd.n6470 585
R4862 gnd.n6472 gnd.n6471 585
R4863 gnd.n989 gnd.n987 585
R4864 gnd.n1011 gnd.n987 585
R4865 gnd.n6464 gnd.n6463 585
R4866 gnd.n6463 gnd.n6462 585
R4867 gnd.n992 gnd.n991 585
R4868 gnd.n6423 gnd.n992 585
R4869 gnd.n6411 gnd.n1027 585
R4870 gnd.n6395 gnd.n1027 585
R4871 gnd.n6413 gnd.n6412 585
R4872 gnd.n6414 gnd.n6413 585
R4873 gnd.n1028 gnd.n1026 585
R4874 gnd.n1044 gnd.n1026 585
R4875 gnd.n6406 gnd.n6405 585
R4876 gnd.n6405 gnd.n6404 585
R4877 gnd.n1031 gnd.n1030 585
R4878 gnd.n1049 gnd.n1031 585
R4879 gnd.n6353 gnd.n1065 585
R4880 gnd.n1065 gnd.n1055 585
R4881 gnd.n6355 gnd.n6354 585
R4882 gnd.n6356 gnd.n6355 585
R4883 gnd.n1066 gnd.n1064 585
R4884 gnd.n1064 gnd.n1059 585
R4885 gnd.n6348 gnd.n6347 585
R4886 gnd.n6347 gnd.n6346 585
R4887 gnd.n1069 gnd.n1068 585
R4888 gnd.n5970 gnd.n1069 585
R4889 gnd.n6331 gnd.n6330 585
R4890 gnd.n6332 gnd.n6331 585
R4891 gnd.n1084 gnd.n1083 585
R4892 gnd.n5959 gnd.n1083 585
R4893 gnd.n6326 gnd.n6325 585
R4894 gnd.n6325 gnd.n6324 585
R4895 gnd.n1087 gnd.n1086 585
R4896 gnd.n5810 gnd.n1087 585
R4897 gnd.n6315 gnd.n6314 585
R4898 gnd.n6316 gnd.n6315 585
R4899 gnd.n1098 gnd.n1097 585
R4900 gnd.n5815 gnd.n1097 585
R4901 gnd.n6310 gnd.n6309 585
R4902 gnd.n6309 gnd.n6308 585
R4903 gnd.n1101 gnd.n1100 585
R4904 gnd.n5821 gnd.n1101 585
R4905 gnd.n6299 gnd.n6298 585
R4906 gnd.n6300 gnd.n6299 585
R4907 gnd.n1111 gnd.n1110 585
R4908 gnd.n5827 gnd.n1110 585
R4909 gnd.n6294 gnd.n6293 585
R4910 gnd.n6293 gnd.n6292 585
R4911 gnd.n1114 gnd.n1113 585
R4912 gnd.n5832 gnd.n1114 585
R4913 gnd.n6283 gnd.n6282 585
R4914 gnd.n6284 gnd.n6283 585
R4915 gnd.n1125 gnd.n1124 585
R4916 gnd.n5838 gnd.n1124 585
R4917 gnd.n6278 gnd.n6277 585
R4918 gnd.n6277 gnd.n6276 585
R4919 gnd.n1128 gnd.n1127 585
R4920 gnd.n5844 gnd.n1128 585
R4921 gnd.n6267 gnd.n6266 585
R4922 gnd.n6268 gnd.n6267 585
R4923 gnd.n1139 gnd.n1138 585
R4924 gnd.n5850 gnd.n1138 585
R4925 gnd.n6262 gnd.n6261 585
R4926 gnd.n6261 gnd.n6260 585
R4927 gnd.n1142 gnd.n1141 585
R4928 gnd.n5863 gnd.n1142 585
R4929 gnd.n6251 gnd.n6250 585
R4930 gnd.n6252 gnd.n6251 585
R4931 gnd.n1155 gnd.n1154 585
R4932 gnd.n6022 gnd.n1154 585
R4933 gnd.n6246 gnd.n6245 585
R4934 gnd.n6245 gnd.n6244 585
R4935 gnd.n1158 gnd.n1157 585
R4936 gnd.n1324 gnd.n1158 585
R4937 gnd.n6235 gnd.n6234 585
R4938 gnd.n6236 gnd.n6235 585
R4939 gnd.n1169 gnd.n1168 585
R4940 gnd.n1439 gnd.n1168 585
R4941 gnd.n6230 gnd.n6229 585
R4942 gnd.n6229 gnd.n6228 585
R4943 gnd.n1172 gnd.n1171 585
R4944 gnd.n1182 gnd.n1172 585
R4945 gnd.n6219 gnd.n6218 585
R4946 gnd.n6220 gnd.n6219 585
R4947 gnd.n1184 gnd.n1183 585
R4948 gnd.n1183 gnd.n1180 585
R4949 gnd.n6214 gnd.n6213 585
R4950 gnd.n6213 gnd.n6212 585
R4951 gnd.n1187 gnd.n1186 585
R4952 gnd.n1196 gnd.n1187 585
R4953 gnd.n6203 gnd.n6202 585
R4954 gnd.n6204 gnd.n6203 585
R4955 gnd.n1198 gnd.n1197 585
R4956 gnd.n1197 gnd.n1194 585
R4957 gnd.n6198 gnd.n6197 585
R4958 gnd.n6197 gnd.n6196 585
R4959 gnd.n1201 gnd.n1200 585
R4960 gnd.n1202 gnd.n1201 585
R4961 gnd.n6187 gnd.n6186 585
R4962 gnd.n6188 gnd.n6187 585
R4963 gnd.n1212 gnd.n1211 585
R4964 gnd.n1211 gnd.n1209 585
R4965 gnd.n6182 gnd.n6181 585
R4966 gnd.n6181 gnd.n6180 585
R4967 gnd.n1215 gnd.n1214 585
R4968 gnd.n1216 gnd.n1215 585
R4969 gnd.n6171 gnd.n6170 585
R4970 gnd.n6172 gnd.n6171 585
R4971 gnd.n1225 gnd.n1224 585
R4972 gnd.n1231 gnd.n1224 585
R4973 gnd.n6166 gnd.n6165 585
R4974 gnd.n6165 gnd.n6164 585
R4975 gnd.n1228 gnd.n1227 585
R4976 gnd.n1229 gnd.n1228 585
R4977 gnd.n5516 gnd.n5515 585
R4978 gnd.n5516 gnd.n1456 585
R4979 gnd.n5520 gnd.n5519 585
R4980 gnd.n5519 gnd.n5518 585
R4981 gnd.n5521 gnd.n5509 585
R4982 gnd.n5517 gnd.n5509 585
R4983 gnd.n5524 gnd.n5522 585
R4984 gnd.n5524 gnd.n5523 585
R4985 gnd.n5525 gnd.n5508 585
R4986 gnd.n5525 gnd.n1245 585
R4987 gnd.n5527 gnd.n5526 585
R4988 gnd.n5526 gnd.n1243 585
R4989 gnd.n5528 gnd.n5503 585
R4990 gnd.n5503 gnd.n1595 585
R4991 gnd.n5530 gnd.n5529 585
R4992 gnd.n5530 gnd.n1603 585
R4993 gnd.n5531 gnd.n5502 585
R4994 gnd.n5531 gnd.n1601 585
R4995 gnd.n5533 gnd.n5532 585
R4996 gnd.n5532 gnd.n1614 585
R4997 gnd.n5534 gnd.n1649 585
R4998 gnd.n1649 gnd.n1611 585
R4999 gnd.n5536 gnd.n5535 585
R5000 gnd.n5537 gnd.n5536 585
R5001 gnd.n1650 gnd.n1648 585
R5002 gnd.n1648 gnd.n1629 585
R5003 gnd.n5496 gnd.n5495 585
R5004 gnd.n5495 gnd.n1627 585
R5005 gnd.n5494 gnd.n1652 585
R5006 gnd.n5494 gnd.n1640 585
R5007 gnd.n5493 gnd.n5492 585
R5008 gnd.n5493 gnd.n1637 585
R5009 gnd.n1654 gnd.n1653 585
R5010 gnd.n1661 gnd.n1653 585
R5011 gnd.n5488 gnd.n5487 585
R5012 gnd.n5487 gnd.n5486 585
R5013 gnd.n1657 gnd.n1656 585
R5014 gnd.n1670 gnd.n1657 585
R5015 gnd.n5431 gnd.n1717 585
R5016 gnd.n1717 gnd.n1716 585
R5017 gnd.n5433 gnd.n5432 585
R5018 gnd.n5434 gnd.n5433 585
R5019 gnd.n1718 gnd.n1715 585
R5020 gnd.n1715 gnd.n1694 585
R5021 gnd.n5426 gnd.n5425 585
R5022 gnd.n5425 gnd.n5424 585
R5023 gnd.n1721 gnd.n1720 585
R5024 gnd.n1721 gnd.n1705 585
R5025 gnd.n5381 gnd.n1752 585
R5026 gnd.n1752 gnd.n1702 585
R5027 gnd.n5383 gnd.n5382 585
R5028 gnd.n5384 gnd.n5383 585
R5029 gnd.n1753 gnd.n1751 585
R5030 gnd.n1751 gnd.n1732 585
R5031 gnd.n5376 gnd.n5375 585
R5032 gnd.n5375 gnd.n5374 585
R5033 gnd.n1756 gnd.n1755 585
R5034 gnd.n1756 gnd.n1743 585
R5035 gnd.n3598 gnd.n3596 585
R5036 gnd.n3596 gnd.n1740 585
R5037 gnd.n3603 gnd.n3602 585
R5038 gnd.n3604 gnd.n3603 585
R5039 gnd.n3597 gnd.n1809 585
R5040 gnd.n1809 gnd.n1768 585
R5041 gnd.n7093 gnd.n7092 585
R5042 gnd.n7094 gnd.n7093 585
R5043 gnd.n750 gnd.n748 585
R5044 gnd.n748 gnd.n745 585
R5045 gnd.n6810 gnd.n786 585
R5046 gnd.n7063 gnd.n786 585
R5047 gnd.n6813 gnd.n6809 585
R5048 gnd.n6809 gnd.n785 585
R5049 gnd.n6814 gnd.n793 585
R5050 gnd.n7055 gnd.n793 585
R5051 gnd.n6815 gnd.n6808 585
R5052 gnd.n6808 gnd.n792 585
R5053 gnd.n6806 gnd.n799 585
R5054 gnd.n7044 gnd.n799 585
R5055 gnd.n6819 gnd.n6805 585
R5056 gnd.n6805 gnd.n807 585
R5057 gnd.n6820 gnd.n806 585
R5058 gnd.n7036 gnd.n806 585
R5059 gnd.n6821 gnd.n6804 585
R5060 gnd.n6804 gnd.n805 585
R5061 gnd.n6802 gnd.n814 585
R5062 gnd.n7028 gnd.n814 585
R5063 gnd.n6825 gnd.n6801 585
R5064 gnd.n6801 gnd.n813 585
R5065 gnd.n6826 gnd.n821 585
R5066 gnd.n7020 gnd.n821 585
R5067 gnd.n6827 gnd.n6800 585
R5068 gnd.n6800 gnd.n820 585
R5069 gnd.n6798 gnd.n828 585
R5070 gnd.n7012 gnd.n828 585
R5071 gnd.n6831 gnd.n6797 585
R5072 gnd.n6797 gnd.n827 585
R5073 gnd.n6832 gnd.n834 585
R5074 gnd.n7004 gnd.n834 585
R5075 gnd.n6833 gnd.n6796 585
R5076 gnd.n6796 gnd.n842 585
R5077 gnd.n6794 gnd.n841 585
R5078 gnd.n6996 gnd.n841 585
R5079 gnd.n6837 gnd.n6793 585
R5080 gnd.n6793 gnd.n6792 585
R5081 gnd.n6838 gnd.n848 585
R5082 gnd.n6988 gnd.n848 585
R5083 gnd.n6839 gnd.n6507 585
R5084 gnd.n6653 gnd.n6507 585
R5085 gnd.n6505 gnd.n856 585
R5086 gnd.n6980 gnd.n856 585
R5087 gnd.n6843 gnd.n6504 585
R5088 gnd.n6590 gnd.n6504 585
R5089 gnd.n6844 gnd.n863 585
R5090 gnd.n6972 gnd.n863 585
R5091 gnd.n6845 gnd.n6503 585
R5092 gnd.n6638 gnd.n6503 585
R5093 gnd.n6501 gnd.n871 585
R5094 gnd.n6964 gnd.n871 585
R5095 gnd.n6849 gnd.n6500 585
R5096 gnd.n6600 gnd.n6500 585
R5097 gnd.n6850 gnd.n878 585
R5098 gnd.n6956 gnd.n878 585
R5099 gnd.n6851 gnd.n6499 585
R5100 gnd.n6620 gnd.n6499 585
R5101 gnd.n972 gnd.n885 585
R5102 gnd.n6948 gnd.n885 585
R5103 gnd.n6856 gnd.n6855 585
R5104 gnd.n6857 gnd.n6856 585
R5105 gnd.n971 gnd.n892 585
R5106 gnd.n6940 gnd.n892 585
R5107 gnd.n6495 gnd.n6494 585
R5108 gnd.n6494 gnd.n962 585
R5109 gnd.n6493 gnd.n898 585
R5110 gnd.n6932 gnd.n898 585
R5111 gnd.n6492 gnd.n954 585
R5112 gnd.n6872 gnd.n954 585
R5113 gnd.n974 gnd.n904 585
R5114 gnd.n6924 gnd.n904 585
R5115 gnd.n6488 gnd.n6487 585
R5116 gnd.n6487 gnd.n946 585
R5117 gnd.n6486 gnd.n911 585
R5118 gnd.n6916 gnd.n911 585
R5119 gnd.n6485 gnd.n941 585
R5120 gnd.n6887 gnd.n941 585
R5121 gnd.n976 gnd.n918 585
R5122 gnd.n6908 gnd.n918 585
R5123 gnd.n6481 gnd.n6480 585
R5124 gnd.n6480 gnd.n934 585
R5125 gnd.n6479 gnd.n926 585
R5126 gnd.n6900 gnd.n926 585
R5127 gnd.n6478 gnd.n979 585
R5128 gnd.n6449 gnd.n979 585
R5129 gnd.n983 gnd.n978 585
R5130 gnd.n6440 gnd.n983 585
R5131 gnd.n6474 gnd.n6473 585
R5132 gnd.n6473 gnd.n6472 585
R5133 gnd.n982 gnd.n981 585
R5134 gnd.n1011 gnd.n982 585
R5135 gnd.n1019 gnd.n994 585
R5136 gnd.n6462 gnd.n994 585
R5137 gnd.n6422 gnd.n6421 585
R5138 gnd.n6423 gnd.n6422 585
R5139 gnd.n1018 gnd.n1017 585
R5140 gnd.n6395 gnd.n1017 585
R5141 gnd.n6416 gnd.n6415 585
R5142 gnd.n6415 gnd.n6414 585
R5143 gnd.n1022 gnd.n1021 585
R5144 gnd.n1044 gnd.n1022 585
R5145 gnd.n5978 gnd.n1033 585
R5146 gnd.n6404 gnd.n1033 585
R5147 gnd.n5979 gnd.n5976 585
R5148 gnd.n5976 gnd.n1049 585
R5149 gnd.n5980 gnd.n5975 585
R5150 gnd.n5975 gnd.n1055 585
R5151 gnd.n5973 gnd.n1061 585
R5152 gnd.n6356 gnd.n1061 585
R5153 gnd.n5984 gnd.n5972 585
R5154 gnd.n5972 gnd.n1059 585
R5155 gnd.n5985 gnd.n1070 585
R5156 gnd.n6346 gnd.n1070 585
R5157 gnd.n5986 gnd.n5971 585
R5158 gnd.n5971 gnd.n5970 585
R5159 gnd.n5798 gnd.n1081 585
R5160 gnd.n6332 gnd.n1081 585
R5161 gnd.n5990 gnd.n5797 585
R5162 gnd.n5959 gnd.n5797 585
R5163 gnd.n5991 gnd.n1089 585
R5164 gnd.n6324 gnd.n1089 585
R5165 gnd.n5992 gnd.n5796 585
R5166 gnd.n5810 gnd.n5796 585
R5167 gnd.n5794 gnd.n1096 585
R5168 gnd.n6316 gnd.n1096 585
R5169 gnd.n5996 gnd.n5793 585
R5170 gnd.n5815 gnd.n5793 585
R5171 gnd.n5997 gnd.n1103 585
R5172 gnd.n6308 gnd.n1103 585
R5173 gnd.n5998 gnd.n5792 585
R5174 gnd.n5821 gnd.n5792 585
R5175 gnd.n5790 gnd.n1109 585
R5176 gnd.n6300 gnd.n1109 585
R5177 gnd.n6002 gnd.n5789 585
R5178 gnd.n5827 gnd.n5789 585
R5179 gnd.n6003 gnd.n1115 585
R5180 gnd.n6292 gnd.n1115 585
R5181 gnd.n6004 gnd.n5788 585
R5182 gnd.n5832 gnd.n5788 585
R5183 gnd.n5786 gnd.n1122 585
R5184 gnd.n6284 gnd.n1122 585
R5185 gnd.n6008 gnd.n5785 585
R5186 gnd.n5838 gnd.n5785 585
R5187 gnd.n6009 gnd.n1129 585
R5188 gnd.n6276 gnd.n1129 585
R5189 gnd.n6010 gnd.n5784 585
R5190 gnd.n5844 gnd.n5784 585
R5191 gnd.n5782 gnd.n1136 585
R5192 gnd.n6268 gnd.n1136 585
R5193 gnd.n6014 gnd.n5781 585
R5194 gnd.n5850 gnd.n5781 585
R5195 gnd.n6015 gnd.n1144 585
R5196 gnd.n6260 gnd.n1144 585
R5197 gnd.n6016 gnd.n5780 585
R5198 gnd.n5863 gnd.n5780 585
R5199 gnd.n1436 gnd.n1152 585
R5200 gnd.n6252 gnd.n1152 585
R5201 gnd.n6021 gnd.n6020 585
R5202 gnd.n6022 gnd.n6021 585
R5203 gnd.n1435 gnd.n1159 585
R5204 gnd.n6244 gnd.n1159 585
R5205 gnd.n5776 gnd.n5775 585
R5206 gnd.n5775 gnd.n1324 585
R5207 gnd.n5774 gnd.n1166 585
R5208 gnd.n6236 gnd.n1166 585
R5209 gnd.n5773 gnd.n1440 585
R5210 gnd.n1440 gnd.n1439 585
R5211 gnd.n1438 gnd.n1173 585
R5212 gnd.n6228 gnd.n1173 585
R5213 gnd.n5769 gnd.n5768 585
R5214 gnd.n5768 gnd.n1182 585
R5215 gnd.n5767 gnd.n1181 585
R5216 gnd.n6220 gnd.n1181 585
R5217 gnd.n5766 gnd.n1443 585
R5218 gnd.n1443 gnd.n1180 585
R5219 gnd.n1442 gnd.n1188 585
R5220 gnd.n6212 gnd.n1188 585
R5221 gnd.n5762 gnd.n5761 585
R5222 gnd.n5761 gnd.n1196 585
R5223 gnd.n5760 gnd.n1195 585
R5224 gnd.n6204 gnd.n1195 585
R5225 gnd.n5759 gnd.n1446 585
R5226 gnd.n1446 gnd.n1194 585
R5227 gnd.n1445 gnd.n1203 585
R5228 gnd.n6196 gnd.n1203 585
R5229 gnd.n5755 gnd.n5754 585
R5230 gnd.n5754 gnd.n1202 585
R5231 gnd.n5753 gnd.n1210 585
R5232 gnd.n6188 gnd.n1210 585
R5233 gnd.n5752 gnd.n1449 585
R5234 gnd.n1449 gnd.n1209 585
R5235 gnd.n1448 gnd.n1217 585
R5236 gnd.n6180 gnd.n1217 585
R5237 gnd.n5748 gnd.n5747 585
R5238 gnd.n5747 gnd.n1216 585
R5239 gnd.n5746 gnd.n1223 585
R5240 gnd.n6172 gnd.n1223 585
R5241 gnd.n5745 gnd.n1452 585
R5242 gnd.n1452 gnd.n1231 585
R5243 gnd.n1451 gnd.n1230 585
R5244 gnd.n6164 gnd.n1230 585
R5245 gnd.n5741 gnd.n5740 585
R5246 gnd.n1455 gnd.n1454 585
R5247 gnd.n5737 gnd.n5736 585
R5248 gnd.n5738 gnd.n5737 585
R5249 gnd.n1472 gnd.n1471 585
R5250 gnd.n5732 gnd.n1474 585
R5251 gnd.n5731 gnd.n1475 585
R5252 gnd.n5730 gnd.n1476 585
R5253 gnd.n1478 gnd.n1477 585
R5254 gnd.n5725 gnd.n5610 585
R5255 gnd.n5724 gnd.n5611 585
R5256 gnd.n5621 gnd.n5612 585
R5257 gnd.n5717 gnd.n5622 585
R5258 gnd.n5716 gnd.n5623 585
R5259 gnd.n5625 gnd.n5624 585
R5260 gnd.n5709 gnd.n5633 585
R5261 gnd.n5708 gnd.n5634 585
R5262 gnd.n5644 gnd.n5635 585
R5263 gnd.n5701 gnd.n5645 585
R5264 gnd.n5700 gnd.n5646 585
R5265 gnd.n5648 gnd.n5647 585
R5266 gnd.n5693 gnd.n5656 585
R5267 gnd.n5692 gnd.n5657 585
R5268 gnd.n5667 gnd.n5658 585
R5269 gnd.n5685 gnd.n5668 585
R5270 gnd.n5684 gnd.n5669 585
R5271 gnd.n5675 gnd.n5674 585
R5272 gnd.n1468 gnd.n1234 585
R5273 gnd.n6158 gnd.n1235 585
R5274 gnd.n6159 gnd.n1232 585
R5275 gnd.n7096 gnd.n7095 585
R5276 gnd.n7095 gnd.n7094 585
R5277 gnd.n743 gnd.n742 585
R5278 gnd.n745 gnd.n743 585
R5279 gnd.n7062 gnd.n7061 585
R5280 gnd.n7063 gnd.n7062 585
R5281 gnd.n788 gnd.n787 585
R5282 gnd.n787 gnd.n785 585
R5283 gnd.n7057 gnd.n7056 585
R5284 gnd.n7056 gnd.n7055 585
R5285 gnd.n791 gnd.n790 585
R5286 gnd.n792 gnd.n791 585
R5287 gnd.n7043 gnd.n7042 585
R5288 gnd.n7044 gnd.n7043 585
R5289 gnd.n801 gnd.n800 585
R5290 gnd.n807 gnd.n800 585
R5291 gnd.n7038 gnd.n7037 585
R5292 gnd.n7037 gnd.n7036 585
R5293 gnd.n804 gnd.n803 585
R5294 gnd.n805 gnd.n804 585
R5295 gnd.n7027 gnd.n7026 585
R5296 gnd.n7028 gnd.n7027 585
R5297 gnd.n816 gnd.n815 585
R5298 gnd.n815 gnd.n813 585
R5299 gnd.n7022 gnd.n7021 585
R5300 gnd.n7021 gnd.n7020 585
R5301 gnd.n819 gnd.n818 585
R5302 gnd.n820 gnd.n819 585
R5303 gnd.n7011 gnd.n7010 585
R5304 gnd.n7012 gnd.n7011 585
R5305 gnd.n830 gnd.n829 585
R5306 gnd.n829 gnd.n827 585
R5307 gnd.n7006 gnd.n7005 585
R5308 gnd.n7005 gnd.n7004 585
R5309 gnd.n833 gnd.n832 585
R5310 gnd.n842 gnd.n833 585
R5311 gnd.n6995 gnd.n6994 585
R5312 gnd.n6996 gnd.n6995 585
R5313 gnd.n844 gnd.n843 585
R5314 gnd.n6792 gnd.n843 585
R5315 gnd.n6990 gnd.n6989 585
R5316 gnd.n6989 gnd.n6988 585
R5317 gnd.n847 gnd.n846 585
R5318 gnd.n6653 gnd.n847 585
R5319 gnd.n6979 gnd.n6978 585
R5320 gnd.n6980 gnd.n6979 585
R5321 gnd.n858 gnd.n857 585
R5322 gnd.n6590 gnd.n857 585
R5323 gnd.n6974 gnd.n6973 585
R5324 gnd.n6973 gnd.n6972 585
R5325 gnd.n861 gnd.n860 585
R5326 gnd.n6638 gnd.n861 585
R5327 gnd.n6963 gnd.n6962 585
R5328 gnd.n6964 gnd.n6963 585
R5329 gnd.n873 gnd.n872 585
R5330 gnd.n6600 gnd.n872 585
R5331 gnd.n6958 gnd.n6957 585
R5332 gnd.n6957 gnd.n6956 585
R5333 gnd.n876 gnd.n875 585
R5334 gnd.n6620 gnd.n876 585
R5335 gnd.n6947 gnd.n6946 585
R5336 gnd.n6948 gnd.n6947 585
R5337 gnd.n887 gnd.n886 585
R5338 gnd.n6857 gnd.n886 585
R5339 gnd.n6942 gnd.n6941 585
R5340 gnd.n6941 gnd.n6940 585
R5341 gnd.n890 gnd.n889 585
R5342 gnd.n962 gnd.n890 585
R5343 gnd.n6931 gnd.n6930 585
R5344 gnd.n6932 gnd.n6931 585
R5345 gnd.n900 gnd.n899 585
R5346 gnd.n6872 gnd.n899 585
R5347 gnd.n6926 gnd.n6925 585
R5348 gnd.n6925 gnd.n6924 585
R5349 gnd.n903 gnd.n902 585
R5350 gnd.n946 gnd.n903 585
R5351 gnd.n6915 gnd.n6914 585
R5352 gnd.n6916 gnd.n6915 585
R5353 gnd.n914 gnd.n913 585
R5354 gnd.n6887 gnd.n913 585
R5355 gnd.n6910 gnd.n6909 585
R5356 gnd.n6909 gnd.n6908 585
R5357 gnd.n917 gnd.n916 585
R5358 gnd.n934 gnd.n917 585
R5359 gnd.n6451 gnd.n928 585
R5360 gnd.n6900 gnd.n928 585
R5361 gnd.n6454 gnd.n6450 585
R5362 gnd.n6450 gnd.n6449 585
R5363 gnd.n6455 gnd.n1002 585
R5364 gnd.n6440 gnd.n1002 585
R5365 gnd.n6456 gnd.n986 585
R5366 gnd.n6472 gnd.n986 585
R5367 gnd.n999 gnd.n997 585
R5368 gnd.n1011 gnd.n997 585
R5369 gnd.n6461 gnd.n6460 585
R5370 gnd.n6462 gnd.n6461 585
R5371 gnd.n998 gnd.n996 585
R5372 gnd.n6423 gnd.n996 585
R5373 gnd.n6397 gnd.n6396 585
R5374 gnd.n6396 gnd.n6395 585
R5375 gnd.n6398 gnd.n1025 585
R5376 gnd.n6414 gnd.n1025 585
R5377 gnd.n1038 gnd.n1036 585
R5378 gnd.n1044 gnd.n1036 585
R5379 gnd.n6403 gnd.n6402 585
R5380 gnd.n6404 gnd.n6403 585
R5381 gnd.n1037 gnd.n1035 585
R5382 gnd.n1049 gnd.n1035 585
R5383 gnd.n6339 gnd.n6338 585
R5384 gnd.n6338 gnd.n1055 585
R5385 gnd.n6340 gnd.n1063 585
R5386 gnd.n6356 gnd.n1063 585
R5387 gnd.n1075 gnd.n1073 585
R5388 gnd.n1073 gnd.n1059 585
R5389 gnd.n6345 gnd.n6344 585
R5390 gnd.n6346 gnd.n6345 585
R5391 gnd.n1074 gnd.n1072 585
R5392 gnd.n5970 gnd.n1072 585
R5393 gnd.n6334 gnd.n6333 585
R5394 gnd.n6333 gnd.n6332 585
R5395 gnd.n1078 gnd.n1077 585
R5396 gnd.n5959 gnd.n1078 585
R5397 gnd.n6323 gnd.n6322 585
R5398 gnd.n6324 gnd.n6323 585
R5399 gnd.n1091 gnd.n1090 585
R5400 gnd.n5810 gnd.n1090 585
R5401 gnd.n6318 gnd.n6317 585
R5402 gnd.n6317 gnd.n6316 585
R5403 gnd.n1094 gnd.n1093 585
R5404 gnd.n5815 gnd.n1094 585
R5405 gnd.n6307 gnd.n6306 585
R5406 gnd.n6308 gnd.n6307 585
R5407 gnd.n1105 gnd.n1104 585
R5408 gnd.n5821 gnd.n1104 585
R5409 gnd.n6302 gnd.n6301 585
R5410 gnd.n6301 gnd.n6300 585
R5411 gnd.n1108 gnd.n1107 585
R5412 gnd.n5827 gnd.n1108 585
R5413 gnd.n6291 gnd.n6290 585
R5414 gnd.n6292 gnd.n6291 585
R5415 gnd.n1118 gnd.n1117 585
R5416 gnd.n5832 gnd.n1117 585
R5417 gnd.n6286 gnd.n6285 585
R5418 gnd.n6285 gnd.n6284 585
R5419 gnd.n1121 gnd.n1120 585
R5420 gnd.n5838 gnd.n1121 585
R5421 gnd.n6275 gnd.n6274 585
R5422 gnd.n6276 gnd.n6275 585
R5423 gnd.n1132 gnd.n1131 585
R5424 gnd.n5844 gnd.n1131 585
R5425 gnd.n6270 gnd.n6269 585
R5426 gnd.n6269 gnd.n6268 585
R5427 gnd.n1135 gnd.n1134 585
R5428 gnd.n5850 gnd.n1135 585
R5429 gnd.n6259 gnd.n6258 585
R5430 gnd.n6260 gnd.n6259 585
R5431 gnd.n1147 gnd.n1146 585
R5432 gnd.n5863 gnd.n1146 585
R5433 gnd.n6254 gnd.n6253 585
R5434 gnd.n6253 gnd.n6252 585
R5435 gnd.n1150 gnd.n1149 585
R5436 gnd.n6022 gnd.n1150 585
R5437 gnd.n6243 gnd.n6242 585
R5438 gnd.n6244 gnd.n6243 585
R5439 gnd.n1162 gnd.n1161 585
R5440 gnd.n1324 gnd.n1161 585
R5441 gnd.n6238 gnd.n6237 585
R5442 gnd.n6237 gnd.n6236 585
R5443 gnd.n1165 gnd.n1164 585
R5444 gnd.n1439 gnd.n1165 585
R5445 gnd.n6227 gnd.n6226 585
R5446 gnd.n6228 gnd.n6227 585
R5447 gnd.n1176 gnd.n1175 585
R5448 gnd.n1182 gnd.n1175 585
R5449 gnd.n6222 gnd.n6221 585
R5450 gnd.n6221 gnd.n6220 585
R5451 gnd.n1179 gnd.n1178 585
R5452 gnd.n1180 gnd.n1179 585
R5453 gnd.n6211 gnd.n6210 585
R5454 gnd.n6212 gnd.n6211 585
R5455 gnd.n1190 gnd.n1189 585
R5456 gnd.n1196 gnd.n1189 585
R5457 gnd.n6206 gnd.n6205 585
R5458 gnd.n6205 gnd.n6204 585
R5459 gnd.n1193 gnd.n1192 585
R5460 gnd.n1194 gnd.n1193 585
R5461 gnd.n6195 gnd.n6194 585
R5462 gnd.n6196 gnd.n6195 585
R5463 gnd.n1205 gnd.n1204 585
R5464 gnd.n1204 gnd.n1202 585
R5465 gnd.n6190 gnd.n6189 585
R5466 gnd.n6189 gnd.n6188 585
R5467 gnd.n1208 gnd.n1207 585
R5468 gnd.n1209 gnd.n1208 585
R5469 gnd.n6179 gnd.n6178 585
R5470 gnd.n6180 gnd.n6179 585
R5471 gnd.n1219 gnd.n1218 585
R5472 gnd.n1218 gnd.n1216 585
R5473 gnd.n6174 gnd.n6173 585
R5474 gnd.n6173 gnd.n6172 585
R5475 gnd.n1222 gnd.n1221 585
R5476 gnd.n1231 gnd.n1222 585
R5477 gnd.n6163 gnd.n6162 585
R5478 gnd.n6164 gnd.n6163 585
R5479 gnd.n7114 gnd.n728 585
R5480 gnd.n7078 gnd.n728 585
R5481 gnd.n7115 gnd.n727 585
R5482 gnd.n773 gnd.n721 585
R5483 gnd.n7122 gnd.n720 585
R5484 gnd.n7123 gnd.n719 585
R5485 gnd.n770 gnd.n711 585
R5486 gnd.n7130 gnd.n710 585
R5487 gnd.n7131 gnd.n709 585
R5488 gnd.n768 gnd.n703 585
R5489 gnd.n7138 gnd.n702 585
R5490 gnd.n7139 gnd.n701 585
R5491 gnd.n765 gnd.n693 585
R5492 gnd.n7146 gnd.n692 585
R5493 gnd.n7147 gnd.n691 585
R5494 gnd.n763 gnd.n683 585
R5495 gnd.n7154 gnd.n682 585
R5496 gnd.n7155 gnd.n681 585
R5497 gnd.n7156 gnd.n680 585
R5498 gnd.n7080 gnd.n679 585
R5499 gnd.n7082 gnd.n7081 585
R5500 gnd.n7083 gnd.n757 585
R5501 gnd.n760 gnd.n755 585
R5502 gnd.n7087 gnd.n754 585
R5503 gnd.n7088 gnd.n753 585
R5504 gnd.n7089 gnd.n749 585
R5505 gnd.n744 gnd.n740 585
R5506 gnd.n7103 gnd.n739 585
R5507 gnd.n7104 gnd.n738 585
R5508 gnd.n775 gnd.n737 585
R5509 gnd.n6785 gnd.n6510 482.89
R5510 gnd.n6668 gnd.n6667 482.89
R5511 gnd.n6034 gnd.n6032 482.89
R5512 gnd.n1428 gnd.n1325 482.89
R5513 gnd.n1305 gnd.t156 443.966
R5514 gnd.n6559 gnd.t176 443.966
R5515 gnd.n1362 gnd.t204 443.966
R5516 gnd.n6553 gnd.t105 443.966
R5517 gnd.n2947 gnd.n1934 440.005
R5518 gnd.n5670 gnd.t134 371.625
R5519 gnd.n7108 gnd.t94 371.625
R5520 gnd.n1237 gnd.t123 371.625
R5521 gnd.n629 gnd.t182 371.625
R5522 gnd.n652 gnd.t185 371.625
R5523 gnd.n675 gnd.t147 371.625
R5524 gnd.n350 gnd.t112 371.625
R5525 gnd.n330 gnd.t120 371.625
R5526 gnd.n7848 gnd.t144 371.625
R5527 gnd.n7667 gnd.t191 371.625
R5528 gnd.n3224 gnd.t138 371.625
R5529 gnd.n3246 gnd.t160 371.625
R5530 gnd.n3268 gnd.t179 371.625
R5531 gnd.n3417 gnd.t130 371.625
R5532 gnd.n1281 gnd.t153 371.625
R5533 gnd.n1480 gnd.t170 371.625
R5534 gnd.n1502 gnd.t198 371.625
R5535 gnd.n729 gnd.t98 371.625
R5536 gnd.n4332 gnd.t116 323.425
R5537 gnd.n3858 gnd.t166 323.425
R5538 gnd.n5180 gnd.n5154 289.615
R5539 gnd.n5148 gnd.n5122 289.615
R5540 gnd.n5116 gnd.n5090 289.615
R5541 gnd.n5085 gnd.n5059 289.615
R5542 gnd.n5053 gnd.n5027 289.615
R5543 gnd.n5021 gnd.n4995 289.615
R5544 gnd.n4989 gnd.n4963 289.615
R5545 gnd.n4958 gnd.n4932 289.615
R5546 gnd.n4406 gnd.t90 279.217
R5547 gnd.n3884 gnd.t194 279.217
R5548 gnd.n1334 gnd.t190 260.649
R5549 gnd.n6523 gnd.t104 260.649
R5550 gnd.n1427 gnd.n1174 256.663
R5551 gnd.n1420 gnd.n1174 256.663
R5552 gnd.n1418 gnd.n1174 256.663
R5553 gnd.n1412 gnd.n1174 256.663
R5554 gnd.n1410 gnd.n1174 256.663
R5555 gnd.n1404 gnd.n1174 256.663
R5556 gnd.n1402 gnd.n1174 256.663
R5557 gnd.n1396 gnd.n1174 256.663
R5558 gnd.n1394 gnd.n1174 256.663
R5559 gnd.n1388 gnd.n1174 256.663
R5560 gnd.n1386 gnd.n1174 256.663
R5561 gnd.n1380 gnd.n1174 256.663
R5562 gnd.n1378 gnd.n1174 256.663
R5563 gnd.n1372 gnd.n1174 256.663
R5564 gnd.n1365 gnd.n1174 256.663
R5565 gnd.n1366 gnd.n1174 256.663
R5566 gnd.n6100 gnd.n1303 256.663
R5567 gnd.n6098 gnd.n1174 256.663
R5568 gnd.n6096 gnd.n1174 256.663
R5569 gnd.n6089 gnd.n1174 256.663
R5570 gnd.n6087 gnd.n1174 256.663
R5571 gnd.n6081 gnd.n1174 256.663
R5572 gnd.n6079 gnd.n1174 256.663
R5573 gnd.n6073 gnd.n1174 256.663
R5574 gnd.n6071 gnd.n1174 256.663
R5575 gnd.n6065 gnd.n1174 256.663
R5576 gnd.n6063 gnd.n1174 256.663
R5577 gnd.n6057 gnd.n1174 256.663
R5578 gnd.n6055 gnd.n1174 256.663
R5579 gnd.n6049 gnd.n1174 256.663
R5580 gnd.n6047 gnd.n1174 256.663
R5581 gnd.n6041 gnd.n1174 256.663
R5582 gnd.n6039 gnd.n1174 256.663
R5583 gnd.n6033 gnd.n1174 256.663
R5584 gnd.n6666 gnd.n6532 256.663
R5585 gnd.n6673 gnd.n6532 256.663
R5586 gnd.n6580 gnd.n6532 256.663
R5587 gnd.n6680 gnd.n6532 256.663
R5588 gnd.n6577 gnd.n6532 256.663
R5589 gnd.n6687 gnd.n6532 256.663
R5590 gnd.n6574 gnd.n6532 256.663
R5591 gnd.n6694 gnd.n6532 256.663
R5592 gnd.n6571 gnd.n6532 256.663
R5593 gnd.n6701 gnd.n6532 256.663
R5594 gnd.n6568 gnd.n6532 256.663
R5595 gnd.n6708 gnd.n6532 256.663
R5596 gnd.n6565 gnd.n6532 256.663
R5597 gnd.n6715 gnd.n6532 256.663
R5598 gnd.n6562 gnd.n6532 256.663
R5599 gnd.n6723 gnd.n6532 256.663
R5600 gnd.n6726 gnd.n639 256.663
R5601 gnd.n6727 gnd.n6532 256.663
R5602 gnd.n6731 gnd.n6532 256.663
R5603 gnd.n6556 gnd.n6532 256.663
R5604 gnd.n6739 gnd.n6532 256.663
R5605 gnd.n6551 gnd.n6532 256.663
R5606 gnd.n6746 gnd.n6532 256.663
R5607 gnd.n6548 gnd.n6532 256.663
R5608 gnd.n6753 gnd.n6532 256.663
R5609 gnd.n6545 gnd.n6532 256.663
R5610 gnd.n6760 gnd.n6532 256.663
R5611 gnd.n6542 gnd.n6532 256.663
R5612 gnd.n6767 gnd.n6532 256.663
R5613 gnd.n6539 gnd.n6532 256.663
R5614 gnd.n6774 gnd.n6532 256.663
R5615 gnd.n6536 gnd.n6532 256.663
R5616 gnd.n6781 gnd.n6532 256.663
R5617 gnd.n6784 gnd.n6532 256.663
R5618 gnd.n3833 gnd.n3192 242.672
R5619 gnd.n3833 gnd.n3193 242.672
R5620 gnd.n3833 gnd.n3194 242.672
R5621 gnd.n3833 gnd.n3195 242.672
R5622 gnd.n3833 gnd.n3196 242.672
R5623 gnd.n3833 gnd.n3197 242.672
R5624 gnd.n3833 gnd.n3198 242.672
R5625 gnd.n3833 gnd.n3199 242.672
R5626 gnd.n3833 gnd.n3200 242.672
R5627 gnd.n1253 gnd.n1240 242.672
R5628 gnd.n5678 gnd.n1253 242.672
R5629 gnd.n5663 gnd.n1253 242.672
R5630 gnd.n5660 gnd.n1253 242.672
R5631 gnd.n5651 gnd.n1253 242.672
R5632 gnd.n5640 gnd.n1253 242.672
R5633 gnd.n5637 gnd.n1253 242.672
R5634 gnd.n5628 gnd.n1253 242.672
R5635 gnd.n5617 gnd.n1253 242.672
R5636 gnd.n4460 gnd.n4459 242.672
R5637 gnd.n4460 gnd.n4370 242.672
R5638 gnd.n4460 gnd.n4371 242.672
R5639 gnd.n4460 gnd.n4372 242.672
R5640 gnd.n4460 gnd.n4373 242.672
R5641 gnd.n4460 gnd.n4374 242.672
R5642 gnd.n4460 gnd.n4375 242.672
R5643 gnd.n4460 gnd.n4376 242.672
R5644 gnd.n4460 gnd.n4377 242.672
R5645 gnd.n4460 gnd.n4378 242.672
R5646 gnd.n4460 gnd.n4379 242.672
R5647 gnd.n4460 gnd.n4380 242.672
R5648 gnd.n4461 gnd.n4460 242.672
R5649 gnd.n5312 gnd.n3163 242.672
R5650 gnd.n5312 gnd.n3162 242.672
R5651 gnd.n5312 gnd.n3161 242.672
R5652 gnd.n5312 gnd.n3160 242.672
R5653 gnd.n5312 gnd.n3159 242.672
R5654 gnd.n5312 gnd.n3158 242.672
R5655 gnd.n5312 gnd.n3157 242.672
R5656 gnd.n5312 gnd.n3156 242.672
R5657 gnd.n5312 gnd.n3155 242.672
R5658 gnd.n5312 gnd.n3154 242.672
R5659 gnd.n5312 gnd.n3153 242.672
R5660 gnd.n5312 gnd.n3152 242.672
R5661 gnd.n5312 gnd.n3151 242.672
R5662 gnd.n7274 gnd.n600 242.672
R5663 gnd.n7274 gnd.n601 242.672
R5664 gnd.n7274 gnd.n602 242.672
R5665 gnd.n7274 gnd.n603 242.672
R5666 gnd.n7274 gnd.n604 242.672
R5667 gnd.n7274 gnd.n605 242.672
R5668 gnd.n7274 gnd.n606 242.672
R5669 gnd.n7274 gnd.n607 242.672
R5670 gnd.n7274 gnd.n608 242.672
R5671 gnd.n7883 gnd.n264 242.672
R5672 gnd.n7883 gnd.n263 242.672
R5673 gnd.n7883 gnd.n262 242.672
R5674 gnd.n7883 gnd.n261 242.672
R5675 gnd.n7883 gnd.n260 242.672
R5676 gnd.n7883 gnd.n259 242.672
R5677 gnd.n7883 gnd.n258 242.672
R5678 gnd.n7883 gnd.n257 242.672
R5679 gnd.n7883 gnd.n256 242.672
R5680 gnd.n4544 gnd.n4543 242.672
R5681 gnd.n4543 gnd.n4282 242.672
R5682 gnd.n4543 gnd.n4283 242.672
R5683 gnd.n4543 gnd.n4284 242.672
R5684 gnd.n4543 gnd.n4285 242.672
R5685 gnd.n4543 gnd.n4286 242.672
R5686 gnd.n4543 gnd.n4287 242.672
R5687 gnd.n4543 gnd.n4288 242.672
R5688 gnd.n5312 gnd.n3834 242.672
R5689 gnd.n5312 gnd.n3835 242.672
R5690 gnd.n5312 gnd.n3836 242.672
R5691 gnd.n5312 gnd.n3837 242.672
R5692 gnd.n5312 gnd.n3838 242.672
R5693 gnd.n5312 gnd.n3839 242.672
R5694 gnd.n5312 gnd.n3840 242.672
R5695 gnd.n5312 gnd.n3841 242.672
R5696 gnd.n3833 gnd.n3832 242.672
R5697 gnd.n3833 gnd.n3164 242.672
R5698 gnd.n3833 gnd.n3165 242.672
R5699 gnd.n3833 gnd.n3166 242.672
R5700 gnd.n3833 gnd.n3167 242.672
R5701 gnd.n3833 gnd.n3168 242.672
R5702 gnd.n3833 gnd.n3169 242.672
R5703 gnd.n3833 gnd.n3170 242.672
R5704 gnd.n3833 gnd.n3171 242.672
R5705 gnd.n3833 gnd.n3172 242.672
R5706 gnd.n3833 gnd.n3173 242.672
R5707 gnd.n3833 gnd.n3174 242.672
R5708 gnd.n3833 gnd.n3175 242.672
R5709 gnd.n3833 gnd.n3176 242.672
R5710 gnd.n3833 gnd.n3177 242.672
R5711 gnd.n3833 gnd.n3178 242.672
R5712 gnd.n3833 gnd.n3179 242.672
R5713 gnd.n3833 gnd.n3180 242.672
R5714 gnd.n3833 gnd.n3181 242.672
R5715 gnd.n3833 gnd.n3182 242.672
R5716 gnd.n3833 gnd.n3183 242.672
R5717 gnd.n3833 gnd.n3184 242.672
R5718 gnd.n3833 gnd.n3185 242.672
R5719 gnd.n3833 gnd.n3186 242.672
R5720 gnd.n3833 gnd.n3187 242.672
R5721 gnd.n3833 gnd.n3188 242.672
R5722 gnd.n3833 gnd.n3189 242.672
R5723 gnd.n3833 gnd.n3190 242.672
R5724 gnd.n3833 gnd.n3191 242.672
R5725 gnd.n1587 gnd.n1253 242.672
R5726 gnd.n1483 gnd.n1253 242.672
R5727 gnd.n1577 gnd.n1253 242.672
R5728 gnd.n1487 gnd.n1253 242.672
R5729 gnd.n1567 gnd.n1253 242.672
R5730 gnd.n1491 gnd.n1253 242.672
R5731 gnd.n1557 gnd.n1253 242.672
R5732 gnd.n1495 gnd.n1253 242.672
R5733 gnd.n1547 gnd.n1253 242.672
R5734 gnd.n1499 gnd.n1253 242.672
R5735 gnd.n1537 gnd.n1253 242.672
R5736 gnd.n1505 gnd.n1253 242.672
R5737 gnd.n1527 gnd.n1253 242.672
R5738 gnd.n1509 gnd.n1253 242.672
R5739 gnd.n1517 gnd.n1253 242.672
R5740 gnd.n1514 gnd.n1253 242.672
R5741 gnd.n6101 gnd.n1299 242.672
R5742 gnd.n1298 gnd.n1253 242.672
R5743 gnd.n6105 gnd.n1253 242.672
R5744 gnd.n1292 gnd.n1253 242.672
R5745 gnd.n6112 gnd.n1253 242.672
R5746 gnd.n1285 gnd.n1253 242.672
R5747 gnd.n6120 gnd.n1253 242.672
R5748 gnd.n1276 gnd.n1253 242.672
R5749 gnd.n6127 gnd.n1253 242.672
R5750 gnd.n1269 gnd.n1253 242.672
R5751 gnd.n6134 gnd.n1253 242.672
R5752 gnd.n1262 gnd.n1253 242.672
R5753 gnd.n6141 gnd.n1253 242.672
R5754 gnd.n6144 gnd.n1253 242.672
R5755 gnd.n7274 gnd.n7273 242.672
R5756 gnd.n7274 gnd.n572 242.672
R5757 gnd.n7274 gnd.n573 242.672
R5758 gnd.n7274 gnd.n574 242.672
R5759 gnd.n7274 gnd.n575 242.672
R5760 gnd.n7274 gnd.n576 242.672
R5761 gnd.n7274 gnd.n577 242.672
R5762 gnd.n7274 gnd.n578 242.672
R5763 gnd.n7274 gnd.n579 242.672
R5764 gnd.n7274 gnd.n580 242.672
R5765 gnd.n7274 gnd.n581 242.672
R5766 gnd.n7274 gnd.n582 242.672
R5767 gnd.n7274 gnd.n583 242.672
R5768 gnd.n7222 gnd.n640 242.672
R5769 gnd.n7274 gnd.n584 242.672
R5770 gnd.n7274 gnd.n585 242.672
R5771 gnd.n7274 gnd.n586 242.672
R5772 gnd.n7274 gnd.n587 242.672
R5773 gnd.n7274 gnd.n588 242.672
R5774 gnd.n7274 gnd.n589 242.672
R5775 gnd.n7274 gnd.n590 242.672
R5776 gnd.n7274 gnd.n591 242.672
R5777 gnd.n7274 gnd.n592 242.672
R5778 gnd.n7274 gnd.n593 242.672
R5779 gnd.n7274 gnd.n594 242.672
R5780 gnd.n7274 gnd.n595 242.672
R5781 gnd.n7274 gnd.n596 242.672
R5782 gnd.n7274 gnd.n597 242.672
R5783 gnd.n7274 gnd.n598 242.672
R5784 gnd.n7274 gnd.n599 242.672
R5785 gnd.n7883 gnd.n265 242.672
R5786 gnd.n7883 gnd.n266 242.672
R5787 gnd.n7883 gnd.n267 242.672
R5788 gnd.n7883 gnd.n268 242.672
R5789 gnd.n7883 gnd.n269 242.672
R5790 gnd.n7883 gnd.n270 242.672
R5791 gnd.n7883 gnd.n271 242.672
R5792 gnd.n7883 gnd.n272 242.672
R5793 gnd.n7883 gnd.n273 242.672
R5794 gnd.n7883 gnd.n274 242.672
R5795 gnd.n7883 gnd.n275 242.672
R5796 gnd.n7883 gnd.n276 242.672
R5797 gnd.n7883 gnd.n277 242.672
R5798 gnd.n7883 gnd.n278 242.672
R5799 gnd.n7883 gnd.n279 242.672
R5800 gnd.n7883 gnd.n280 242.672
R5801 gnd.n7883 gnd.n281 242.672
R5802 gnd.n7883 gnd.n282 242.672
R5803 gnd.n7883 gnd.n283 242.672
R5804 gnd.n7883 gnd.n284 242.672
R5805 gnd.n7883 gnd.n285 242.672
R5806 gnd.n7883 gnd.n286 242.672
R5807 gnd.n7883 gnd.n287 242.672
R5808 gnd.n7883 gnd.n288 242.672
R5809 gnd.n7883 gnd.n289 242.672
R5810 gnd.n7883 gnd.n290 242.672
R5811 gnd.n7883 gnd.n291 242.672
R5812 gnd.n7883 gnd.n292 242.672
R5813 gnd.n7883 gnd.n7882 242.672
R5814 gnd.n5739 gnd.n5738 242.672
R5815 gnd.n5738 gnd.n1457 242.672
R5816 gnd.n5738 gnd.n1458 242.672
R5817 gnd.n5738 gnd.n1459 242.672
R5818 gnd.n5738 gnd.n1460 242.672
R5819 gnd.n5738 gnd.n1461 242.672
R5820 gnd.n5738 gnd.n1462 242.672
R5821 gnd.n5738 gnd.n1463 242.672
R5822 gnd.n5738 gnd.n1464 242.672
R5823 gnd.n5738 gnd.n1465 242.672
R5824 gnd.n5738 gnd.n1466 242.672
R5825 gnd.n5738 gnd.n1467 242.672
R5826 gnd.n5738 gnd.n1469 242.672
R5827 gnd.n5738 gnd.n1470 242.672
R5828 gnd.n7078 gnd.n774 242.672
R5829 gnd.n7078 gnd.n772 242.672
R5830 gnd.n7078 gnd.n771 242.672
R5831 gnd.n7078 gnd.n769 242.672
R5832 gnd.n7078 gnd.n767 242.672
R5833 gnd.n7078 gnd.n766 242.672
R5834 gnd.n7078 gnd.n764 242.672
R5835 gnd.n7078 gnd.n762 242.672
R5836 gnd.n7079 gnd.n7078 242.672
R5837 gnd.n7078 gnd.n758 242.672
R5838 gnd.n7078 gnd.n761 242.672
R5839 gnd.n7078 gnd.n759 242.672
R5840 gnd.n7078 gnd.n777 242.672
R5841 gnd.n7078 gnd.n776 242.672
R5842 gnd.n7884 gnd.n254 240.244
R5843 gnd.n7881 gnd.n293 240.244
R5844 gnd.n7877 gnd.n7876 240.244
R5845 gnd.n7873 gnd.n7872 240.244
R5846 gnd.n7869 gnd.n7868 240.244
R5847 gnd.n7865 gnd.n7864 240.244
R5848 gnd.n7861 gnd.n7860 240.244
R5849 gnd.n7857 gnd.n7856 240.244
R5850 gnd.n7853 gnd.n7852 240.244
R5851 gnd.n7846 gnd.n7845 240.244
R5852 gnd.n7842 gnd.n7841 240.244
R5853 gnd.n7838 gnd.n7837 240.244
R5854 gnd.n7834 gnd.n7833 240.244
R5855 gnd.n7830 gnd.n7829 240.244
R5856 gnd.n7826 gnd.n7825 240.244
R5857 gnd.n7822 gnd.n7821 240.244
R5858 gnd.n7818 gnd.n7817 240.244
R5859 gnd.n7814 gnd.n7813 240.244
R5860 gnd.n7810 gnd.n7809 240.244
R5861 gnd.n7803 gnd.n7802 240.244
R5862 gnd.n7800 gnd.n7799 240.244
R5863 gnd.n7796 gnd.n7795 240.244
R5864 gnd.n7792 gnd.n7791 240.244
R5865 gnd.n7788 gnd.n7787 240.244
R5866 gnd.n7784 gnd.n7783 240.244
R5867 gnd.n7780 gnd.n7779 240.244
R5868 gnd.n7776 gnd.n7775 240.244
R5869 gnd.n7772 gnd.n7771 240.244
R5870 gnd.n7768 gnd.n7767 240.244
R5871 gnd.n7303 gnd.n552 240.244
R5872 gnd.n7303 gnd.n543 240.244
R5873 gnd.n543 gnd.n535 240.244
R5874 gnd.n7330 gnd.n535 240.244
R5875 gnd.n7330 gnd.n523 240.244
R5876 gnd.n7334 gnd.n523 240.244
R5877 gnd.n7334 gnd.n513 240.244
R5878 gnd.n7343 gnd.n513 240.244
R5879 gnd.n7343 gnd.n505 240.244
R5880 gnd.n505 gnd.n487 240.244
R5881 gnd.n7339 gnd.n487 240.244
R5882 gnd.n7339 gnd.n478 240.244
R5883 gnd.n478 gnd.n469 240.244
R5884 gnd.n7421 gnd.n469 240.244
R5885 gnd.n7421 gnd.n457 240.244
R5886 gnd.n7425 gnd.n457 240.244
R5887 gnd.n7425 gnd.n447 240.244
R5888 gnd.n7429 gnd.n447 240.244
R5889 gnd.n7429 gnd.n439 240.244
R5890 gnd.n439 gnd.n422 240.244
R5891 gnd.n7472 gnd.n422 240.244
R5892 gnd.n7472 gnd.n412 240.244
R5893 gnd.n7477 gnd.n412 240.244
R5894 gnd.n7477 gnd.n404 240.244
R5895 gnd.n404 gnd.n384 240.244
R5896 gnd.n7520 gnd.n384 240.244
R5897 gnd.n7521 gnd.n7520 240.244
R5898 gnd.n7521 gnd.n377 240.244
R5899 gnd.n7525 gnd.n377 240.244
R5900 gnd.n7525 gnd.n369 240.244
R5901 gnd.n369 gnd.n364 240.244
R5902 gnd.n364 gnd.n359 240.244
R5903 gnd.n7569 gnd.n359 240.244
R5904 gnd.n7569 gnd.n105 240.244
R5905 gnd.n7578 gnd.n105 240.244
R5906 gnd.n7579 gnd.n7578 240.244
R5907 gnd.n7579 gnd.n122 240.244
R5908 gnd.n7582 gnd.n122 240.244
R5909 gnd.n7582 gnd.n133 240.244
R5910 gnd.n7586 gnd.n133 240.244
R5911 gnd.n7586 gnd.n142 240.244
R5912 gnd.n7589 gnd.n142 240.244
R5913 gnd.n7589 gnd.n151 240.244
R5914 gnd.n7593 gnd.n151 240.244
R5915 gnd.n7593 gnd.n161 240.244
R5916 gnd.n7596 gnd.n161 240.244
R5917 gnd.n7596 gnd.n170 240.244
R5918 gnd.n7600 gnd.n170 240.244
R5919 gnd.n7600 gnd.n180 240.244
R5920 gnd.n7603 gnd.n180 240.244
R5921 gnd.n7603 gnd.n189 240.244
R5922 gnd.n7607 gnd.n189 240.244
R5923 gnd.n7607 gnd.n199 240.244
R5924 gnd.n7742 gnd.n199 240.244
R5925 gnd.n7742 gnd.n208 240.244
R5926 gnd.n7746 gnd.n208 240.244
R5927 gnd.n7746 gnd.n218 240.244
R5928 gnd.n7749 gnd.n218 240.244
R5929 gnd.n7749 gnd.n227 240.244
R5930 gnd.n7753 gnd.n227 240.244
R5931 gnd.n7753 gnd.n237 240.244
R5932 gnd.n7756 gnd.n237 240.244
R5933 gnd.n7756 gnd.n246 240.244
R5934 gnd.n7760 gnd.n246 240.244
R5935 gnd.n7272 gnd.n610 240.244
R5936 gnd.n7268 gnd.n610 240.244
R5937 gnd.n7266 gnd.n7265 240.244
R5938 gnd.n7262 gnd.n7261 240.244
R5939 gnd.n7258 gnd.n7257 240.244
R5940 gnd.n7254 gnd.n7253 240.244
R5941 gnd.n7250 gnd.n7249 240.244
R5942 gnd.n7246 gnd.n7245 240.244
R5943 gnd.n7242 gnd.n7241 240.244
R5944 gnd.n7237 gnd.n7236 240.244
R5945 gnd.n7233 gnd.n7232 240.244
R5946 gnd.n7229 gnd.n7228 240.244
R5947 gnd.n7225 gnd.n7224 240.244
R5948 gnd.n7220 gnd.n7219 240.244
R5949 gnd.n7216 gnd.n7215 240.244
R5950 gnd.n7212 gnd.n7211 240.244
R5951 gnd.n7208 gnd.n7207 240.244
R5952 gnd.n7204 gnd.n7203 240.244
R5953 gnd.n7200 gnd.n7199 240.244
R5954 gnd.n7196 gnd.n7195 240.244
R5955 gnd.n7192 gnd.n7191 240.244
R5956 gnd.n7188 gnd.n7187 240.244
R5957 gnd.n7184 gnd.n7183 240.244
R5958 gnd.n7180 gnd.n7179 240.244
R5959 gnd.n7176 gnd.n7175 240.244
R5960 gnd.n7172 gnd.n7171 240.244
R5961 gnd.n7168 gnd.n7167 240.244
R5962 gnd.n7164 gnd.n7163 240.244
R5963 gnd.n7311 gnd.n546 240.244
R5964 gnd.n7319 gnd.n546 240.244
R5965 gnd.n7319 gnd.n547 240.244
R5966 gnd.n547 gnd.n521 240.244
R5967 gnd.n7353 gnd.n521 240.244
R5968 gnd.n7353 gnd.n516 240.244
R5969 gnd.n7361 gnd.n516 240.244
R5970 gnd.n7361 gnd.n517 240.244
R5971 gnd.n517 gnd.n485 240.244
R5972 gnd.n7402 gnd.n485 240.244
R5973 gnd.n7402 gnd.n480 240.244
R5974 gnd.n7410 gnd.n480 240.244
R5975 gnd.n7410 gnd.n481 240.244
R5976 gnd.n481 gnd.n455 240.244
R5977 gnd.n7439 gnd.n455 240.244
R5978 gnd.n7439 gnd.n450 240.244
R5979 gnd.n7447 gnd.n450 240.244
R5980 gnd.n7447 gnd.n451 240.244
R5981 gnd.n451 gnd.n420 240.244
R5982 gnd.n7487 gnd.n420 240.244
R5983 gnd.n7487 gnd.n415 240.244
R5984 gnd.n7496 gnd.n415 240.244
R5985 gnd.n7496 gnd.n416 240.244
R5986 gnd.n416 gnd.n382 240.244
R5987 gnd.n7537 gnd.n382 240.244
R5988 gnd.n7537 gnd.n379 240.244
R5989 gnd.n7541 gnd.n379 240.244
R5990 gnd.n7544 gnd.n7541 240.244
R5991 gnd.n7544 gnd.n367 240.244
R5992 gnd.n7554 gnd.n367 240.244
R5993 gnd.n7560 gnd.n7554 240.244
R5994 gnd.n7560 gnd.n7557 240.244
R5995 gnd.n7557 gnd.n108 240.244
R5996 gnd.n7976 gnd.n108 240.244
R5997 gnd.n7976 gnd.n109 240.244
R5998 gnd.n119 gnd.n109 240.244
R5999 gnd.n7970 gnd.n119 240.244
R6000 gnd.n7970 gnd.n120 240.244
R6001 gnd.n7962 gnd.n120 240.244
R6002 gnd.n7962 gnd.n136 240.244
R6003 gnd.n7958 gnd.n136 240.244
R6004 gnd.n7958 gnd.n141 240.244
R6005 gnd.n7950 gnd.n141 240.244
R6006 gnd.n7950 gnd.n153 240.244
R6007 gnd.n7946 gnd.n153 240.244
R6008 gnd.n7946 gnd.n159 240.244
R6009 gnd.n7938 gnd.n159 240.244
R6010 gnd.n7938 gnd.n173 240.244
R6011 gnd.n7934 gnd.n173 240.244
R6012 gnd.n7934 gnd.n179 240.244
R6013 gnd.n7926 gnd.n179 240.244
R6014 gnd.n7926 gnd.n191 240.244
R6015 gnd.n7922 gnd.n191 240.244
R6016 gnd.n7922 gnd.n197 240.244
R6017 gnd.n7914 gnd.n197 240.244
R6018 gnd.n7914 gnd.n211 240.244
R6019 gnd.n7910 gnd.n211 240.244
R6020 gnd.n7910 gnd.n217 240.244
R6021 gnd.n7902 gnd.n217 240.244
R6022 gnd.n7902 gnd.n230 240.244
R6023 gnd.n7898 gnd.n230 240.244
R6024 gnd.n7898 gnd.n236 240.244
R6025 gnd.n7890 gnd.n236 240.244
R6026 gnd.n7890 gnd.n249 240.244
R6027 gnd.n6145 gnd.n1248 240.244
R6028 gnd.n6143 gnd.n6142 240.244
R6029 gnd.n6140 gnd.n1255 240.244
R6030 gnd.n6136 gnd.n6135 240.244
R6031 gnd.n6133 gnd.n1263 240.244
R6032 gnd.n6129 gnd.n6128 240.244
R6033 gnd.n6126 gnd.n1270 240.244
R6034 gnd.n6122 gnd.n6121 240.244
R6035 gnd.n6119 gnd.n1277 240.244
R6036 gnd.n6114 gnd.n6113 240.244
R6037 gnd.n6111 gnd.n1286 240.244
R6038 gnd.n6107 gnd.n6106 240.244
R6039 gnd.n6104 gnd.n1293 240.244
R6040 gnd.n1516 gnd.n1515 240.244
R6041 gnd.n1519 gnd.n1518 240.244
R6042 gnd.n1526 gnd.n1525 240.244
R6043 gnd.n1529 gnd.n1528 240.244
R6044 gnd.n1536 gnd.n1535 240.244
R6045 gnd.n1539 gnd.n1538 240.244
R6046 gnd.n1546 gnd.n1545 240.244
R6047 gnd.n1549 gnd.n1548 240.244
R6048 gnd.n1556 gnd.n1555 240.244
R6049 gnd.n1559 gnd.n1558 240.244
R6050 gnd.n1566 gnd.n1565 240.244
R6051 gnd.n1569 gnd.n1568 240.244
R6052 gnd.n1576 gnd.n1575 240.244
R6053 gnd.n1579 gnd.n1578 240.244
R6054 gnd.n1586 gnd.n1585 240.244
R6055 gnd.n3711 gnd.n3710 240.244
R6056 gnd.n3710 gnd.n3275 240.244
R6057 gnd.n3287 gnd.n3275 240.244
R6058 gnd.n3554 gnd.n3287 240.244
R6059 gnd.n3554 gnd.n3299 240.244
R6060 gnd.n3558 gnd.n3299 240.244
R6061 gnd.n3558 gnd.n3309 240.244
R6062 gnd.n3561 gnd.n3309 240.244
R6063 gnd.n3561 gnd.n3318 240.244
R6064 gnd.n3565 gnd.n3318 240.244
R6065 gnd.n3565 gnd.n3328 240.244
R6066 gnd.n3568 gnd.n3328 240.244
R6067 gnd.n3568 gnd.n3337 240.244
R6068 gnd.n3572 gnd.n3337 240.244
R6069 gnd.n3572 gnd.n3347 240.244
R6070 gnd.n3575 gnd.n3347 240.244
R6071 gnd.n3575 gnd.n3356 240.244
R6072 gnd.n3579 gnd.n3356 240.244
R6073 gnd.n3579 gnd.n3366 240.244
R6074 gnd.n3582 gnd.n3366 240.244
R6075 gnd.n3582 gnd.n3375 240.244
R6076 gnd.n3586 gnd.n3375 240.244
R6077 gnd.n3586 gnd.n3385 240.244
R6078 gnd.n3589 gnd.n3385 240.244
R6079 gnd.n3589 gnd.n3394 240.244
R6080 gnd.n3397 gnd.n3394 240.244
R6081 gnd.n3399 gnd.n3397 240.244
R6082 gnd.n3623 gnd.n3399 240.244
R6083 gnd.n3623 gnd.n1782 240.244
R6084 gnd.n3620 gnd.n1782 240.244
R6085 gnd.n3620 gnd.n1793 240.244
R6086 gnd.n3617 gnd.n1793 240.244
R6087 gnd.n3617 gnd.n1797 240.244
R6088 gnd.n3614 gnd.n1797 240.244
R6089 gnd.n3614 gnd.n1806 240.244
R6090 gnd.n3611 gnd.n1806 240.244
R6091 gnd.n3611 gnd.n1767 240.244
R6092 gnd.n1767 gnd.n1759 240.244
R6093 gnd.n5367 gnd.n1759 240.244
R6094 gnd.n5367 gnd.n1741 240.244
R6095 gnd.n5372 gnd.n1741 240.244
R6096 gnd.n5372 gnd.n1731 240.244
R6097 gnd.n1731 gnd.n1724 240.244
R6098 gnd.n5412 gnd.n1724 240.244
R6099 gnd.n5412 gnd.n1703 240.244
R6100 gnd.n5422 gnd.n1703 240.244
R6101 gnd.n5422 gnd.n1693 240.244
R6102 gnd.n1713 gnd.n1693 240.244
R6103 gnd.n5417 gnd.n1713 240.244
R6104 gnd.n5417 gnd.n1668 240.244
R6105 gnd.n1677 gnd.n1668 240.244
R6106 gnd.n1677 gnd.n1659 240.244
R6107 gnd.n5469 gnd.n1659 240.244
R6108 gnd.n5469 gnd.n1638 240.244
R6109 gnd.n1681 gnd.n1638 240.244
R6110 gnd.n1681 gnd.n1628 240.244
R6111 gnd.n1628 gnd.n1620 240.244
R6112 gnd.n5578 gnd.n1620 240.244
R6113 gnd.n5578 gnd.n1612 240.244
R6114 gnd.n1612 gnd.n1600 240.244
R6115 gnd.n5596 gnd.n1600 240.244
R6116 gnd.n5596 gnd.n1594 240.244
R6117 gnd.n5604 gnd.n1594 240.244
R6118 gnd.n5604 gnd.n1244 240.244
R6119 gnd.n3204 gnd.n3203 240.244
R6120 gnd.n3826 gnd.n3203 240.244
R6121 gnd.n3824 gnd.n3823 240.244
R6122 gnd.n3820 gnd.n3819 240.244
R6123 gnd.n3816 gnd.n3815 240.244
R6124 gnd.n3812 gnd.n3811 240.244
R6125 gnd.n3808 gnd.n3807 240.244
R6126 gnd.n3804 gnd.n3803 240.244
R6127 gnd.n3800 gnd.n3799 240.244
R6128 gnd.n3795 gnd.n3794 240.244
R6129 gnd.n3791 gnd.n3790 240.244
R6130 gnd.n3787 gnd.n3786 240.244
R6131 gnd.n3783 gnd.n3782 240.244
R6132 gnd.n3779 gnd.n3778 240.244
R6133 gnd.n3775 gnd.n3774 240.244
R6134 gnd.n3771 gnd.n3770 240.244
R6135 gnd.n3767 gnd.n3766 240.244
R6136 gnd.n3763 gnd.n3762 240.244
R6137 gnd.n3759 gnd.n3758 240.244
R6138 gnd.n3755 gnd.n3754 240.244
R6139 gnd.n3751 gnd.n3750 240.244
R6140 gnd.n3747 gnd.n3746 240.244
R6141 gnd.n3743 gnd.n3742 240.244
R6142 gnd.n3739 gnd.n3738 240.244
R6143 gnd.n3735 gnd.n3734 240.244
R6144 gnd.n3731 gnd.n3730 240.244
R6145 gnd.n3727 gnd.n3726 240.244
R6146 gnd.n3723 gnd.n3722 240.244
R6147 gnd.n3719 gnd.n3718 240.244
R6148 gnd.n3708 gnd.n3205 240.244
R6149 gnd.n3708 gnd.n3278 240.244
R6150 gnd.n3704 gnd.n3278 240.244
R6151 gnd.n3704 gnd.n3285 240.244
R6152 gnd.n3696 gnd.n3285 240.244
R6153 gnd.n3696 gnd.n3302 240.244
R6154 gnd.n3692 gnd.n3302 240.244
R6155 gnd.n3692 gnd.n3308 240.244
R6156 gnd.n3684 gnd.n3308 240.244
R6157 gnd.n3684 gnd.n3320 240.244
R6158 gnd.n3680 gnd.n3320 240.244
R6159 gnd.n3680 gnd.n3326 240.244
R6160 gnd.n3672 gnd.n3326 240.244
R6161 gnd.n3672 gnd.n3340 240.244
R6162 gnd.n3668 gnd.n3340 240.244
R6163 gnd.n3668 gnd.n3346 240.244
R6164 gnd.n3660 gnd.n3346 240.244
R6165 gnd.n3660 gnd.n3358 240.244
R6166 gnd.n3656 gnd.n3358 240.244
R6167 gnd.n3656 gnd.n3364 240.244
R6168 gnd.n3648 gnd.n3364 240.244
R6169 gnd.n3648 gnd.n3378 240.244
R6170 gnd.n3644 gnd.n3378 240.244
R6171 gnd.n3644 gnd.n3384 240.244
R6172 gnd.n3636 gnd.n3384 240.244
R6173 gnd.n3636 gnd.n3631 240.244
R6174 gnd.n3631 gnd.n3396 240.244
R6175 gnd.n3396 gnd.n1780 240.244
R6176 gnd.n5348 gnd.n1780 240.244
R6177 gnd.n5348 gnd.n1781 240.244
R6178 gnd.n5340 gnd.n1781 240.244
R6179 gnd.n5340 gnd.n5337 240.244
R6180 gnd.n5337 gnd.n5334 240.244
R6181 gnd.n5334 gnd.n1796 240.244
R6182 gnd.n5326 gnd.n1796 240.244
R6183 gnd.n5326 gnd.n1770 240.244
R6184 gnd.n5356 gnd.n1770 240.244
R6185 gnd.n5356 gnd.n1771 240.244
R6186 gnd.n1771 gnd.n1739 240.244
R6187 gnd.n5393 gnd.n1739 240.244
R6188 gnd.n5393 gnd.n1734 240.244
R6189 gnd.n5401 gnd.n1734 240.244
R6190 gnd.n5401 gnd.n1735 240.244
R6191 gnd.n1735 gnd.n1701 240.244
R6192 gnd.n5443 gnd.n1701 240.244
R6193 gnd.n5443 gnd.n1696 240.244
R6194 gnd.n5451 gnd.n1696 240.244
R6195 gnd.n5451 gnd.n1697 240.244
R6196 gnd.n1697 gnd.n1667 240.244
R6197 gnd.n5478 gnd.n1667 240.244
R6198 gnd.n5478 gnd.n1663 240.244
R6199 gnd.n5484 gnd.n1663 240.244
R6200 gnd.n5484 gnd.n1636 240.244
R6201 gnd.n5546 gnd.n1636 240.244
R6202 gnd.n5546 gnd.n1631 240.244
R6203 gnd.n5554 gnd.n1631 240.244
R6204 gnd.n5554 gnd.n1632 240.244
R6205 gnd.n1632 gnd.n1610 240.244
R6206 gnd.n5586 gnd.n1610 240.244
R6207 gnd.n5586 gnd.n1605 240.244
R6208 gnd.n5594 gnd.n1605 240.244
R6209 gnd.n5594 gnd.n1606 240.244
R6210 gnd.n1606 gnd.n1247 240.244
R6211 gnd.n6151 gnd.n1247 240.244
R6212 gnd.n5311 gnd.n3843 240.244
R6213 gnd.n5304 gnd.n5303 240.244
R6214 gnd.n5301 gnd.n5300 240.244
R6215 gnd.n5297 gnd.n5296 240.244
R6216 gnd.n5293 gnd.n5292 240.244
R6217 gnd.n5289 gnd.n5288 240.244
R6218 gnd.n5285 gnd.n5284 240.244
R6219 gnd.n5281 gnd.n5280 240.244
R6220 gnd.n4555 gnd.n4267 240.244
R6221 gnd.n4565 gnd.n4267 240.244
R6222 gnd.n4565 gnd.n4258 240.244
R6223 gnd.n4258 gnd.n4247 240.244
R6224 gnd.n4586 gnd.n4247 240.244
R6225 gnd.n4586 gnd.n4241 240.244
R6226 gnd.n4596 gnd.n4241 240.244
R6227 gnd.n4596 gnd.n4230 240.244
R6228 gnd.n4230 gnd.n4222 240.244
R6229 gnd.n4614 gnd.n4222 240.244
R6230 gnd.n4615 gnd.n4614 240.244
R6231 gnd.n4615 gnd.n4207 240.244
R6232 gnd.n4617 gnd.n4207 240.244
R6233 gnd.n4617 gnd.n4193 240.244
R6234 gnd.n4659 gnd.n4193 240.244
R6235 gnd.n4660 gnd.n4659 240.244
R6236 gnd.n4663 gnd.n4660 240.244
R6237 gnd.n4663 gnd.n4148 240.244
R6238 gnd.n4188 gnd.n4148 240.244
R6239 gnd.n4188 gnd.n4158 240.244
R6240 gnd.n4673 gnd.n4158 240.244
R6241 gnd.n4673 gnd.n4179 240.244
R6242 gnd.n4683 gnd.n4179 240.244
R6243 gnd.n4683 gnd.n4045 240.244
R6244 gnd.n4728 gnd.n4045 240.244
R6245 gnd.n4728 gnd.n4031 240.244
R6246 gnd.n4750 gnd.n4031 240.244
R6247 gnd.n4751 gnd.n4750 240.244
R6248 gnd.n4751 gnd.n4018 240.244
R6249 gnd.n4018 gnd.n4007 240.244
R6250 gnd.n4782 gnd.n4007 240.244
R6251 gnd.n4783 gnd.n4782 240.244
R6252 gnd.n4784 gnd.n4783 240.244
R6253 gnd.n4784 gnd.n3992 240.244
R6254 gnd.n3992 gnd.n3991 240.244
R6255 gnd.n3991 gnd.n3976 240.244
R6256 gnd.n4835 gnd.n3976 240.244
R6257 gnd.n4836 gnd.n4835 240.244
R6258 gnd.n4836 gnd.n3963 240.244
R6259 gnd.n3963 gnd.n3952 240.244
R6260 gnd.n4867 gnd.n3952 240.244
R6261 gnd.n4868 gnd.n4867 240.244
R6262 gnd.n4869 gnd.n4868 240.244
R6263 gnd.n4869 gnd.n3936 240.244
R6264 gnd.n3936 gnd.n3935 240.244
R6265 gnd.n3935 gnd.n3922 240.244
R6266 gnd.n4924 gnd.n3922 240.244
R6267 gnd.n4925 gnd.n4924 240.244
R6268 gnd.n4925 gnd.n3909 240.244
R6269 gnd.n3909 gnd.n3899 240.244
R6270 gnd.n5212 gnd.n3899 240.244
R6271 gnd.n5215 gnd.n5212 240.244
R6272 gnd.n5215 gnd.n5214 240.244
R6273 gnd.n4545 gnd.n4280 240.244
R6274 gnd.n4301 gnd.n4280 240.244
R6275 gnd.n4304 gnd.n4303 240.244
R6276 gnd.n4311 gnd.n4310 240.244
R6277 gnd.n4314 gnd.n4313 240.244
R6278 gnd.n4321 gnd.n4320 240.244
R6279 gnd.n4324 gnd.n4323 240.244
R6280 gnd.n4331 gnd.n4330 240.244
R6281 gnd.n4553 gnd.n4277 240.244
R6282 gnd.n4277 gnd.n4256 240.244
R6283 gnd.n4576 gnd.n4256 240.244
R6284 gnd.n4576 gnd.n4250 240.244
R6285 gnd.n4584 gnd.n4250 240.244
R6286 gnd.n4584 gnd.n4252 240.244
R6287 gnd.n4252 gnd.n4228 240.244
R6288 gnd.n4606 gnd.n4228 240.244
R6289 gnd.n4606 gnd.n4224 240.244
R6290 gnd.n4612 gnd.n4224 240.244
R6291 gnd.n4612 gnd.n4206 240.244
R6292 gnd.n4637 gnd.n4206 240.244
R6293 gnd.n4637 gnd.n4201 240.244
R6294 gnd.n4649 gnd.n4201 240.244
R6295 gnd.n4649 gnd.n4202 240.244
R6296 gnd.n4645 gnd.n4202 240.244
R6297 gnd.n4645 gnd.n4150 240.244
R6298 gnd.n4697 gnd.n4150 240.244
R6299 gnd.n4697 gnd.n4151 240.244
R6300 gnd.n4693 gnd.n4151 240.244
R6301 gnd.n4693 gnd.n4157 240.244
R6302 gnd.n4177 gnd.n4157 240.244
R6303 gnd.n4177 gnd.n4043 240.244
R6304 gnd.n4732 gnd.n4043 240.244
R6305 gnd.n4732 gnd.n4038 240.244
R6306 gnd.n4740 gnd.n4038 240.244
R6307 gnd.n4740 gnd.n4039 240.244
R6308 gnd.n4039 gnd.n4016 240.244
R6309 gnd.n4772 gnd.n4016 240.244
R6310 gnd.n4772 gnd.n4011 240.244
R6311 gnd.n4780 gnd.n4011 240.244
R6312 gnd.n4780 gnd.n4012 240.244
R6313 gnd.n4012 gnd.n3989 240.244
R6314 gnd.n4817 gnd.n3989 240.244
R6315 gnd.n4817 gnd.n3984 240.244
R6316 gnd.n4825 gnd.n3984 240.244
R6317 gnd.n4825 gnd.n3985 240.244
R6318 gnd.n3985 gnd.n3961 240.244
R6319 gnd.n4857 gnd.n3961 240.244
R6320 gnd.n4857 gnd.n3956 240.244
R6321 gnd.n4865 gnd.n3956 240.244
R6322 gnd.n4865 gnd.n3957 240.244
R6323 gnd.n3957 gnd.n3934 240.244
R6324 gnd.n4906 gnd.n3934 240.244
R6325 gnd.n4906 gnd.n3929 240.244
R6326 gnd.n4914 gnd.n3929 240.244
R6327 gnd.n4914 gnd.n3930 240.244
R6328 gnd.n3930 gnd.n3907 240.244
R6329 gnd.n5200 gnd.n3907 240.244
R6330 gnd.n5200 gnd.n3902 240.244
R6331 gnd.n5210 gnd.n3902 240.244
R6332 gnd.n5210 gnd.n3903 240.244
R6333 gnd.n3903 gnd.n3842 240.244
R6334 gnd.n7678 gnd.n255 240.244
R6335 gnd.n7684 gnd.n7683 240.244
R6336 gnd.n7687 gnd.n7686 240.244
R6337 gnd.n7694 gnd.n7693 240.244
R6338 gnd.n7697 gnd.n7696 240.244
R6339 gnd.n7704 gnd.n7703 240.244
R6340 gnd.n7707 gnd.n7706 240.244
R6341 gnd.n7714 gnd.n7713 240.244
R6342 gnd.n7717 gnd.n7716 240.244
R6343 gnd.n553 gnd.n542 240.244
R6344 gnd.n7321 gnd.n542 240.244
R6345 gnd.n7321 gnd.n537 240.244
R6346 gnd.n7328 gnd.n537 240.244
R6347 gnd.n7328 gnd.n524 240.244
R6348 gnd.n524 gnd.n511 240.244
R6349 gnd.n7363 gnd.n511 240.244
R6350 gnd.n7363 gnd.n506 240.244
R6351 gnd.n7370 gnd.n506 240.244
R6352 gnd.n7370 gnd.n488 240.244
R6353 gnd.n488 gnd.n476 240.244
R6354 gnd.n7412 gnd.n476 240.244
R6355 gnd.n7412 gnd.n471 240.244
R6356 gnd.n7419 gnd.n471 240.244
R6357 gnd.n7419 gnd.n458 240.244
R6358 gnd.n458 gnd.n445 240.244
R6359 gnd.n7449 gnd.n445 240.244
R6360 gnd.n7449 gnd.n440 240.244
R6361 gnd.n7456 gnd.n440 240.244
R6362 gnd.n7456 gnd.n423 240.244
R6363 gnd.n423 gnd.n410 240.244
R6364 gnd.n7498 gnd.n410 240.244
R6365 gnd.n7498 gnd.n405 240.244
R6366 gnd.n7507 gnd.n405 240.244
R6367 gnd.n7507 gnd.n385 240.244
R6368 gnd.n395 gnd.n385 240.244
R6369 gnd.n395 gnd.n375 240.244
R6370 gnd.n7546 gnd.n375 240.244
R6371 gnd.n7546 gnd.n370 240.244
R6372 gnd.n7552 gnd.n370 240.244
R6373 gnd.n7552 gnd.n366 240.244
R6374 gnd.n366 gnd.n365 240.244
R6375 gnd.n365 gnd.n102 240.244
R6376 gnd.n7978 gnd.n102 240.244
R6377 gnd.n7978 gnd.n104 240.244
R6378 gnd.n7620 gnd.n104 240.244
R6379 gnd.n7620 gnd.n123 240.244
R6380 gnd.n7625 gnd.n123 240.244
R6381 gnd.n7625 gnd.n134 240.244
R6382 gnd.n7628 gnd.n134 240.244
R6383 gnd.n7628 gnd.n143 240.244
R6384 gnd.n7633 gnd.n143 240.244
R6385 gnd.n7633 gnd.n152 240.244
R6386 gnd.n7636 gnd.n152 240.244
R6387 gnd.n7636 gnd.n162 240.244
R6388 gnd.n7641 gnd.n162 240.244
R6389 gnd.n7641 gnd.n171 240.244
R6390 gnd.n7644 gnd.n171 240.244
R6391 gnd.n7644 gnd.n181 240.244
R6392 gnd.n7649 gnd.n181 240.244
R6393 gnd.n7649 gnd.n190 240.244
R6394 gnd.n7652 gnd.n190 240.244
R6395 gnd.n7652 gnd.n200 240.244
R6396 gnd.n7740 gnd.n200 240.244
R6397 gnd.n7740 gnd.n209 240.244
R6398 gnd.n7736 gnd.n209 240.244
R6399 gnd.n7736 gnd.n219 240.244
R6400 gnd.n7733 gnd.n219 240.244
R6401 gnd.n7733 gnd.n228 240.244
R6402 gnd.n7730 gnd.n228 240.244
R6403 gnd.n7730 gnd.n238 240.244
R6404 gnd.n7727 gnd.n238 240.244
R6405 gnd.n7727 gnd.n247 240.244
R6406 gnd.n7724 gnd.n247 240.244
R6407 gnd.n688 gnd.n687 240.244
R6408 gnd.n696 gnd.n695 240.244
R6409 gnd.n698 gnd.n697 240.244
R6410 gnd.n706 gnd.n705 240.244
R6411 gnd.n714 gnd.n713 240.244
R6412 gnd.n716 gnd.n715 240.244
R6413 gnd.n724 gnd.n723 240.244
R6414 gnd.n734 gnd.n733 240.244
R6415 gnd.n7107 gnd.n609 240.244
R6416 gnd.n7309 gnd.n556 240.244
R6417 gnd.n556 gnd.n545 240.244
R6418 gnd.n560 gnd.n545 240.244
R6419 gnd.n560 gnd.n526 240.244
R6420 gnd.n7351 gnd.n526 240.244
R6421 gnd.n7351 gnd.n527 240.244
R6422 gnd.n527 gnd.n515 240.244
R6423 gnd.n7346 gnd.n515 240.244
R6424 gnd.n7346 gnd.n490 240.244
R6425 gnd.n7400 gnd.n490 240.244
R6426 gnd.n7400 gnd.n491 240.244
R6427 gnd.n491 gnd.n479 240.244
R6428 gnd.n7395 gnd.n479 240.244
R6429 gnd.n7395 gnd.n460 240.244
R6430 gnd.n7437 gnd.n460 240.244
R6431 gnd.n7437 gnd.n461 240.244
R6432 gnd.n461 gnd.n449 240.244
R6433 gnd.n7432 gnd.n449 240.244
R6434 gnd.n7432 gnd.n424 240.244
R6435 gnd.n7485 gnd.n424 240.244
R6436 gnd.n7485 gnd.n425 240.244
R6437 gnd.n425 gnd.n414 240.244
R6438 gnd.n7480 gnd.n414 240.244
R6439 gnd.n7480 gnd.n386 240.244
R6440 gnd.n7535 gnd.n386 240.244
R6441 gnd.n7535 gnd.n387 240.244
R6442 gnd.n7531 gnd.n387 240.244
R6443 gnd.n7531 gnd.n378 240.244
R6444 gnd.n7528 gnd.n378 240.244
R6445 gnd.n7528 gnd.n363 240.244
R6446 gnd.n7562 gnd.n363 240.244
R6447 gnd.n7562 gnd.n357 240.244
R6448 gnd.n7571 gnd.n357 240.244
R6449 gnd.n7571 gnd.n107 240.244
R6450 gnd.n7574 gnd.n107 240.244
R6451 gnd.n7574 gnd.n125 240.244
R6452 gnd.n7968 gnd.n125 240.244
R6453 gnd.n7968 gnd.n126 240.244
R6454 gnd.n7964 gnd.n126 240.244
R6455 gnd.n7964 gnd.n132 240.244
R6456 gnd.n7956 gnd.n132 240.244
R6457 gnd.n7956 gnd.n144 240.244
R6458 gnd.n7952 gnd.n144 240.244
R6459 gnd.n7952 gnd.n149 240.244
R6460 gnd.n7944 gnd.n149 240.244
R6461 gnd.n7944 gnd.n164 240.244
R6462 gnd.n7940 gnd.n164 240.244
R6463 gnd.n7940 gnd.n169 240.244
R6464 gnd.n7932 gnd.n169 240.244
R6465 gnd.n7932 gnd.n182 240.244
R6466 gnd.n7928 gnd.n182 240.244
R6467 gnd.n7928 gnd.n187 240.244
R6468 gnd.n7920 gnd.n187 240.244
R6469 gnd.n7920 gnd.n202 240.244
R6470 gnd.n7916 gnd.n202 240.244
R6471 gnd.n7916 gnd.n207 240.244
R6472 gnd.n7908 gnd.n207 240.244
R6473 gnd.n7908 gnd.n220 240.244
R6474 gnd.n7904 gnd.n220 240.244
R6475 gnd.n7904 gnd.n225 240.244
R6476 gnd.n7896 gnd.n225 240.244
R6477 gnd.n7896 gnd.n240 240.244
R6478 gnd.n7892 gnd.n240 240.244
R6479 gnd.n7892 gnd.n245 240.244
R6480 gnd.n3862 gnd.n3150 240.244
R6481 gnd.n5271 gnd.n5270 240.244
R6482 gnd.n5267 gnd.n5266 240.244
R6483 gnd.n5263 gnd.n5262 240.244
R6484 gnd.n5259 gnd.n5258 240.244
R6485 gnd.n5255 gnd.n5254 240.244
R6486 gnd.n5251 gnd.n5250 240.244
R6487 gnd.n5247 gnd.n5246 240.244
R6488 gnd.n5243 gnd.n5242 240.244
R6489 gnd.n5239 gnd.n5238 240.244
R6490 gnd.n5235 gnd.n5234 240.244
R6491 gnd.n5231 gnd.n5230 240.244
R6492 gnd.n5227 gnd.n5226 240.244
R6493 gnd.n4468 gnd.n4365 240.244
R6494 gnd.n4468 gnd.n4358 240.244
R6495 gnd.n4479 gnd.n4358 240.244
R6496 gnd.n4479 gnd.n4354 240.244
R6497 gnd.n4485 gnd.n4354 240.244
R6498 gnd.n4485 gnd.n4346 240.244
R6499 gnd.n4495 gnd.n4346 240.244
R6500 gnd.n4495 gnd.n4341 240.244
R6501 gnd.n4531 gnd.n4341 240.244
R6502 gnd.n4531 gnd.n4342 240.244
R6503 gnd.n4342 gnd.n4289 240.244
R6504 gnd.n4526 gnd.n4289 240.244
R6505 gnd.n4526 gnd.n4525 240.244
R6506 gnd.n4525 gnd.n4268 240.244
R6507 gnd.n4521 gnd.n4268 240.244
R6508 gnd.n4521 gnd.n4259 240.244
R6509 gnd.n4518 gnd.n4259 240.244
R6510 gnd.n4518 gnd.n4517 240.244
R6511 gnd.n4517 gnd.n4242 240.244
R6512 gnd.n4513 gnd.n4242 240.244
R6513 gnd.n4513 gnd.n4231 240.244
R6514 gnd.n4231 gnd.n4212 240.244
R6515 gnd.n4626 gnd.n4212 240.244
R6516 gnd.n4626 gnd.n4208 240.244
R6517 gnd.n4634 gnd.n4208 240.244
R6518 gnd.n4634 gnd.n4199 240.244
R6519 gnd.n4199 gnd.n4135 240.244
R6520 gnd.n4706 gnd.n4135 240.244
R6521 gnd.n4706 gnd.n4136 240.244
R6522 gnd.n4147 gnd.n4136 240.244
R6523 gnd.n4182 gnd.n4147 240.244
R6524 gnd.n4185 gnd.n4182 240.244
R6525 gnd.n4185 gnd.n4159 240.244
R6526 gnd.n4172 gnd.n4159 240.244
R6527 gnd.n4172 gnd.n4169 240.244
R6528 gnd.n4169 gnd.n4046 240.244
R6529 gnd.n4727 gnd.n4046 240.244
R6530 gnd.n4727 gnd.n4036 240.244
R6531 gnd.n4723 gnd.n4036 240.244
R6532 gnd.n4723 gnd.n4030 240.244
R6533 gnd.n4720 gnd.n4030 240.244
R6534 gnd.n4720 gnd.n4019 240.244
R6535 gnd.n4717 gnd.n4019 240.244
R6536 gnd.n4717 gnd.n3997 240.244
R6537 gnd.n4793 gnd.n3997 240.244
R6538 gnd.n4793 gnd.n3993 240.244
R6539 gnd.n4814 gnd.n3993 240.244
R6540 gnd.n4814 gnd.n3982 240.244
R6541 gnd.n4810 gnd.n3982 240.244
R6542 gnd.n4810 gnd.n3975 240.244
R6543 gnd.n4807 gnd.n3975 240.244
R6544 gnd.n4807 gnd.n3964 240.244
R6545 gnd.n4804 gnd.n3964 240.244
R6546 gnd.n4804 gnd.n3941 240.244
R6547 gnd.n4878 gnd.n3941 240.244
R6548 gnd.n4878 gnd.n3937 240.244
R6549 gnd.n4903 gnd.n3937 240.244
R6550 gnd.n4903 gnd.n3928 240.244
R6551 gnd.n4899 gnd.n3928 240.244
R6552 gnd.n4899 gnd.n3921 240.244
R6553 gnd.n4895 gnd.n3921 240.244
R6554 gnd.n4895 gnd.n3910 240.244
R6555 gnd.n4892 gnd.n3910 240.244
R6556 gnd.n4892 gnd.n3891 240.244
R6557 gnd.n5222 gnd.n3891 240.244
R6558 gnd.n4382 gnd.n4381 240.244
R6559 gnd.n4453 gnd.n4381 240.244
R6560 gnd.n4451 gnd.n4450 240.244
R6561 gnd.n4447 gnd.n4446 240.244
R6562 gnd.n4443 gnd.n4442 240.244
R6563 gnd.n4439 gnd.n4438 240.244
R6564 gnd.n4435 gnd.n4434 240.244
R6565 gnd.n4431 gnd.n4430 240.244
R6566 gnd.n4427 gnd.n4426 240.244
R6567 gnd.n4423 gnd.n4422 240.244
R6568 gnd.n4419 gnd.n4418 240.244
R6569 gnd.n4415 gnd.n4414 240.244
R6570 gnd.n4411 gnd.n4369 240.244
R6571 gnd.n4471 gnd.n4363 240.244
R6572 gnd.n4471 gnd.n4359 240.244
R6573 gnd.n4477 gnd.n4359 240.244
R6574 gnd.n4477 gnd.n4352 240.244
R6575 gnd.n4487 gnd.n4352 240.244
R6576 gnd.n4487 gnd.n4348 240.244
R6577 gnd.n4493 gnd.n4348 240.244
R6578 gnd.n4493 gnd.n4339 240.244
R6579 gnd.n4533 gnd.n4339 240.244
R6580 gnd.n4533 gnd.n4290 240.244
R6581 gnd.n4541 gnd.n4290 240.244
R6582 gnd.n4541 gnd.n4291 240.244
R6583 gnd.n4291 gnd.n4269 240.244
R6584 gnd.n4562 gnd.n4269 240.244
R6585 gnd.n4562 gnd.n4261 240.244
R6586 gnd.n4573 gnd.n4261 240.244
R6587 gnd.n4573 gnd.n4262 240.244
R6588 gnd.n4262 gnd.n4243 240.244
R6589 gnd.n4593 gnd.n4243 240.244
R6590 gnd.n4593 gnd.n4233 240.244
R6591 gnd.n4603 gnd.n4233 240.244
R6592 gnd.n4603 gnd.n4214 240.244
R6593 gnd.n4624 gnd.n4214 240.244
R6594 gnd.n4624 gnd.n4216 240.244
R6595 gnd.n4216 gnd.n4197 240.244
R6596 gnd.n4652 gnd.n4197 240.244
R6597 gnd.n4652 gnd.n4139 240.244
R6598 gnd.n4704 gnd.n4139 240.244
R6599 gnd.n4704 gnd.n4140 240.244
R6600 gnd.n4700 gnd.n4140 240.244
R6601 gnd.n4700 gnd.n4146 240.244
R6602 gnd.n4161 gnd.n4146 240.244
R6603 gnd.n4690 gnd.n4161 240.244
R6604 gnd.n4690 gnd.n4162 240.244
R6605 gnd.n4686 gnd.n4162 240.244
R6606 gnd.n4686 gnd.n4168 240.244
R6607 gnd.n4168 gnd.n4035 240.244
R6608 gnd.n4743 gnd.n4035 240.244
R6609 gnd.n4743 gnd.n4028 240.244
R6610 gnd.n4754 gnd.n4028 240.244
R6611 gnd.n4754 gnd.n4021 240.244
R6612 gnd.n4769 gnd.n4021 240.244
R6613 gnd.n4769 gnd.n4022 240.244
R6614 gnd.n4022 gnd.n4000 240.244
R6615 gnd.n4791 gnd.n4000 240.244
R6616 gnd.n4791 gnd.n4001 240.244
R6617 gnd.n4001 gnd.n3980 240.244
R6618 gnd.n4828 gnd.n3980 240.244
R6619 gnd.n4828 gnd.n3973 240.244
R6620 gnd.n4839 gnd.n3973 240.244
R6621 gnd.n4839 gnd.n3966 240.244
R6622 gnd.n4854 gnd.n3966 240.244
R6623 gnd.n4854 gnd.n3967 240.244
R6624 gnd.n3967 gnd.n3944 240.244
R6625 gnd.n4876 gnd.n3944 240.244
R6626 gnd.n4876 gnd.n3946 240.244
R6627 gnd.n3946 gnd.n3926 240.244
R6628 gnd.n4917 gnd.n3926 240.244
R6629 gnd.n4917 gnd.n3919 240.244
R6630 gnd.n4928 gnd.n3919 240.244
R6631 gnd.n4928 gnd.n3912 240.244
R6632 gnd.n5197 gnd.n3912 240.244
R6633 gnd.n5197 gnd.n3913 240.244
R6634 gnd.n3913 gnd.n3894 240.244
R6635 gnd.n5220 gnd.n3894 240.244
R6636 gnd.n5616 gnd.n5615 240.244
R6637 gnd.n5627 gnd.n5618 240.244
R6638 gnd.n5630 gnd.n5629 240.244
R6639 gnd.n5639 gnd.n5638 240.244
R6640 gnd.n5650 gnd.n5641 240.244
R6641 gnd.n5653 gnd.n5652 240.244
R6642 gnd.n5662 gnd.n5661 240.244
R6643 gnd.n5677 gnd.n5664 240.244
R6644 gnd.n5680 gnd.n5679 240.244
R6645 gnd.n3474 gnd.n3276 240.244
R6646 gnd.n3477 gnd.n3276 240.244
R6647 gnd.n3477 gnd.n3288 240.244
R6648 gnd.n3482 gnd.n3288 240.244
R6649 gnd.n3482 gnd.n3300 240.244
R6650 gnd.n3485 gnd.n3300 240.244
R6651 gnd.n3485 gnd.n3310 240.244
R6652 gnd.n3490 gnd.n3310 240.244
R6653 gnd.n3490 gnd.n3319 240.244
R6654 gnd.n3493 gnd.n3319 240.244
R6655 gnd.n3493 gnd.n3329 240.244
R6656 gnd.n3498 gnd.n3329 240.244
R6657 gnd.n3498 gnd.n3338 240.244
R6658 gnd.n3501 gnd.n3338 240.244
R6659 gnd.n3501 gnd.n3348 240.244
R6660 gnd.n3506 gnd.n3348 240.244
R6661 gnd.n3506 gnd.n3357 240.244
R6662 gnd.n3509 gnd.n3357 240.244
R6663 gnd.n3509 gnd.n3367 240.244
R6664 gnd.n3514 gnd.n3367 240.244
R6665 gnd.n3514 gnd.n3376 240.244
R6666 gnd.n3517 gnd.n3376 240.244
R6667 gnd.n3517 gnd.n3386 240.244
R6668 gnd.n3522 gnd.n3386 240.244
R6669 gnd.n3522 gnd.n3395 240.244
R6670 gnd.n3398 gnd.n3395 240.244
R6671 gnd.n3400 gnd.n3398 240.244
R6672 gnd.n3547 gnd.n3400 240.244
R6673 gnd.n3547 gnd.n1783 240.244
R6674 gnd.n3543 gnd.n1783 240.244
R6675 gnd.n3543 gnd.n1794 240.244
R6676 gnd.n3532 gnd.n1794 240.244
R6677 gnd.n3532 gnd.n1798 240.244
R6678 gnd.n3535 gnd.n1798 240.244
R6679 gnd.n3535 gnd.n1807 240.244
R6680 gnd.n1807 gnd.n1765 240.244
R6681 gnd.n5358 gnd.n1765 240.244
R6682 gnd.n5358 gnd.n1760 240.244
R6683 gnd.n5365 gnd.n1760 240.244
R6684 gnd.n5365 gnd.n1742 240.244
R6685 gnd.n1742 gnd.n1730 240.244
R6686 gnd.n5403 gnd.n1730 240.244
R6687 gnd.n5403 gnd.n1725 240.244
R6688 gnd.n5410 gnd.n1725 240.244
R6689 gnd.n5410 gnd.n1704 240.244
R6690 gnd.n1704 gnd.n1691 240.244
R6691 gnd.n5453 gnd.n1691 240.244
R6692 gnd.n5453 gnd.n1692 240.244
R6693 gnd.n1692 gnd.n1688 240.244
R6694 gnd.n1688 gnd.n1669 240.244
R6695 gnd.n5460 gnd.n1669 240.244
R6696 gnd.n5460 gnd.n1660 240.244
R6697 gnd.n5467 gnd.n1660 240.244
R6698 gnd.n5467 gnd.n1639 240.244
R6699 gnd.n1639 gnd.n1626 240.244
R6700 gnd.n5556 gnd.n1626 240.244
R6701 gnd.n5556 gnd.n1621 240.244
R6702 gnd.n5576 gnd.n1621 240.244
R6703 gnd.n5576 gnd.n1613 240.244
R6704 gnd.n5562 gnd.n1613 240.244
R6705 gnd.n5562 gnd.n1602 240.244
R6706 gnd.n5564 gnd.n1602 240.244
R6707 gnd.n5564 gnd.n1241 240.244
R6708 gnd.n6153 gnd.n1241 240.244
R6709 gnd.n3434 gnd.n3433 240.244
R6710 gnd.n3440 gnd.n3439 240.244
R6711 gnd.n3444 gnd.n3443 240.244
R6712 gnd.n3450 gnd.n3449 240.244
R6713 gnd.n3454 gnd.n3453 240.244
R6714 gnd.n3460 gnd.n3459 240.244
R6715 gnd.n3464 gnd.n3463 240.244
R6716 gnd.n3421 gnd.n3420 240.244
R6717 gnd.n3416 gnd.n3201 240.244
R6718 gnd.n3429 gnd.n3277 240.244
R6719 gnd.n3290 gnd.n3277 240.244
R6720 gnd.n3702 gnd.n3290 240.244
R6721 gnd.n3702 gnd.n3291 240.244
R6722 gnd.n3698 gnd.n3291 240.244
R6723 gnd.n3698 gnd.n3298 240.244
R6724 gnd.n3690 gnd.n3298 240.244
R6725 gnd.n3690 gnd.n3312 240.244
R6726 gnd.n3686 gnd.n3312 240.244
R6727 gnd.n3686 gnd.n3317 240.244
R6728 gnd.n3678 gnd.n3317 240.244
R6729 gnd.n3678 gnd.n3331 240.244
R6730 gnd.n3674 gnd.n3331 240.244
R6731 gnd.n3674 gnd.n3336 240.244
R6732 gnd.n3666 gnd.n3336 240.244
R6733 gnd.n3666 gnd.n3350 240.244
R6734 gnd.n3662 gnd.n3350 240.244
R6735 gnd.n3662 gnd.n3355 240.244
R6736 gnd.n3654 gnd.n3355 240.244
R6737 gnd.n3654 gnd.n3369 240.244
R6738 gnd.n3650 gnd.n3369 240.244
R6739 gnd.n3650 gnd.n3374 240.244
R6740 gnd.n3642 gnd.n3374 240.244
R6741 gnd.n3642 gnd.n3388 240.244
R6742 gnd.n3638 gnd.n3388 240.244
R6743 gnd.n3638 gnd.n3393 240.244
R6744 gnd.n3628 gnd.n3393 240.244
R6745 gnd.n3628 gnd.n1785 240.244
R6746 gnd.n5346 gnd.n1785 240.244
R6747 gnd.n5346 gnd.n1786 240.244
R6748 gnd.n5342 gnd.n1786 240.244
R6749 gnd.n5342 gnd.n1792 240.244
R6750 gnd.n5332 gnd.n1792 240.244
R6751 gnd.n5332 gnd.n1799 240.244
R6752 gnd.n5328 gnd.n1799 240.244
R6753 gnd.n5328 gnd.n1804 240.244
R6754 gnd.n1804 gnd.n1769 240.244
R6755 gnd.n3606 gnd.n1769 240.244
R6756 gnd.n3606 gnd.n1744 240.244
R6757 gnd.n5391 gnd.n1744 240.244
R6758 gnd.n5391 gnd.n1745 240.244
R6759 gnd.n1745 gnd.n1733 240.244
R6760 gnd.n5386 gnd.n1733 240.244
R6761 gnd.n5386 gnd.n1706 240.244
R6762 gnd.n5441 gnd.n1706 240.244
R6763 gnd.n5441 gnd.n1707 240.244
R6764 gnd.n1707 gnd.n1695 240.244
R6765 gnd.n5436 gnd.n1695 240.244
R6766 gnd.n5436 gnd.n1671 240.244
R6767 gnd.n5476 gnd.n1671 240.244
R6768 gnd.n5476 gnd.n1672 240.244
R6769 gnd.n1672 gnd.n1662 240.244
R6770 gnd.n1662 gnd.n1641 240.244
R6771 gnd.n5544 gnd.n1641 240.244
R6772 gnd.n5544 gnd.n1642 240.244
R6773 gnd.n1642 gnd.n1630 240.244
R6774 gnd.n5539 gnd.n1630 240.244
R6775 gnd.n5539 gnd.n1615 240.244
R6776 gnd.n5584 gnd.n1615 240.244
R6777 gnd.n5584 gnd.n1616 240.244
R6778 gnd.n1616 gnd.n1604 240.244
R6779 gnd.n1604 gnd.n1596 240.244
R6780 gnd.n5602 gnd.n1596 240.244
R6781 gnd.n5602 gnd.n1246 240.244
R6782 gnd.n2940 gnd.n1935 240.244
R6783 gnd.n2940 gnd.n1938 240.244
R6784 gnd.n2936 gnd.n1938 240.244
R6785 gnd.n2936 gnd.n1940 240.244
R6786 gnd.n2932 gnd.n1940 240.244
R6787 gnd.n2932 gnd.n1946 240.244
R6788 gnd.n2928 gnd.n1946 240.244
R6789 gnd.n2928 gnd.n1948 240.244
R6790 gnd.n2924 gnd.n1948 240.244
R6791 gnd.n2924 gnd.n1954 240.244
R6792 gnd.n2920 gnd.n1954 240.244
R6793 gnd.n2920 gnd.n1956 240.244
R6794 gnd.n2916 gnd.n1956 240.244
R6795 gnd.n2916 gnd.n1962 240.244
R6796 gnd.n2912 gnd.n1962 240.244
R6797 gnd.n2912 gnd.n1964 240.244
R6798 gnd.n2908 gnd.n1964 240.244
R6799 gnd.n2908 gnd.n1970 240.244
R6800 gnd.n2904 gnd.n1970 240.244
R6801 gnd.n2904 gnd.n1972 240.244
R6802 gnd.n2900 gnd.n1972 240.244
R6803 gnd.n2900 gnd.n1978 240.244
R6804 gnd.n2896 gnd.n1978 240.244
R6805 gnd.n2896 gnd.n1980 240.244
R6806 gnd.n2892 gnd.n1980 240.244
R6807 gnd.n2892 gnd.n1986 240.244
R6808 gnd.n2888 gnd.n1986 240.244
R6809 gnd.n2888 gnd.n1988 240.244
R6810 gnd.n2884 gnd.n1988 240.244
R6811 gnd.n2884 gnd.n1994 240.244
R6812 gnd.n2880 gnd.n1994 240.244
R6813 gnd.n2880 gnd.n1996 240.244
R6814 gnd.n2876 gnd.n1996 240.244
R6815 gnd.n2876 gnd.n2002 240.244
R6816 gnd.n2872 gnd.n2002 240.244
R6817 gnd.n2872 gnd.n2004 240.244
R6818 gnd.n2868 gnd.n2004 240.244
R6819 gnd.n2868 gnd.n2010 240.244
R6820 gnd.n2864 gnd.n2010 240.244
R6821 gnd.n2864 gnd.n2012 240.244
R6822 gnd.n2860 gnd.n2012 240.244
R6823 gnd.n2860 gnd.n2018 240.244
R6824 gnd.n2856 gnd.n2018 240.244
R6825 gnd.n2856 gnd.n2020 240.244
R6826 gnd.n2852 gnd.n2020 240.244
R6827 gnd.n2852 gnd.n2026 240.244
R6828 gnd.n2848 gnd.n2026 240.244
R6829 gnd.n2848 gnd.n2028 240.244
R6830 gnd.n2844 gnd.n2028 240.244
R6831 gnd.n2844 gnd.n2034 240.244
R6832 gnd.n2840 gnd.n2034 240.244
R6833 gnd.n2840 gnd.n2036 240.244
R6834 gnd.n2836 gnd.n2036 240.244
R6835 gnd.n2836 gnd.n2042 240.244
R6836 gnd.n2832 gnd.n2042 240.244
R6837 gnd.n2832 gnd.n2044 240.244
R6838 gnd.n2828 gnd.n2044 240.244
R6839 gnd.n2828 gnd.n2050 240.244
R6840 gnd.n2824 gnd.n2050 240.244
R6841 gnd.n2824 gnd.n2052 240.244
R6842 gnd.n2820 gnd.n2052 240.244
R6843 gnd.n2820 gnd.n2058 240.244
R6844 gnd.n2816 gnd.n2058 240.244
R6845 gnd.n2816 gnd.n2060 240.244
R6846 gnd.n2812 gnd.n2060 240.244
R6847 gnd.n2812 gnd.n2066 240.244
R6848 gnd.n2808 gnd.n2066 240.244
R6849 gnd.n2808 gnd.n2068 240.244
R6850 gnd.n2804 gnd.n2068 240.244
R6851 gnd.n2804 gnd.n2074 240.244
R6852 gnd.n2800 gnd.n2074 240.244
R6853 gnd.n2800 gnd.n2076 240.244
R6854 gnd.n2796 gnd.n2076 240.244
R6855 gnd.n2796 gnd.n2082 240.244
R6856 gnd.n2792 gnd.n2082 240.244
R6857 gnd.n2792 gnd.n2084 240.244
R6858 gnd.n2788 gnd.n2084 240.244
R6859 gnd.n2788 gnd.n2090 240.244
R6860 gnd.n2784 gnd.n2090 240.244
R6861 gnd.n2784 gnd.n2092 240.244
R6862 gnd.n2780 gnd.n2092 240.244
R6863 gnd.n2780 gnd.n2098 240.244
R6864 gnd.n2776 gnd.n2098 240.244
R6865 gnd.n2776 gnd.n2100 240.244
R6866 gnd.n2772 gnd.n2100 240.244
R6867 gnd.n2772 gnd.n2106 240.244
R6868 gnd.n2768 gnd.n2106 240.244
R6869 gnd.n2768 gnd.n2108 240.244
R6870 gnd.n2764 gnd.n2108 240.244
R6871 gnd.n2764 gnd.n2114 240.244
R6872 gnd.n2760 gnd.n2114 240.244
R6873 gnd.n2760 gnd.n2116 240.244
R6874 gnd.n2756 gnd.n2116 240.244
R6875 gnd.n2756 gnd.n2122 240.244
R6876 gnd.n2752 gnd.n2122 240.244
R6877 gnd.n2752 gnd.n2124 240.244
R6878 gnd.n2748 gnd.n2124 240.244
R6879 gnd.n2748 gnd.n2130 240.244
R6880 gnd.n2744 gnd.n2130 240.244
R6881 gnd.n2744 gnd.n2132 240.244
R6882 gnd.n2740 gnd.n2132 240.244
R6883 gnd.n2740 gnd.n2138 240.244
R6884 gnd.n2736 gnd.n2138 240.244
R6885 gnd.n2736 gnd.n2140 240.244
R6886 gnd.n2732 gnd.n2140 240.244
R6887 gnd.n2732 gnd.n2146 240.244
R6888 gnd.n2728 gnd.n2146 240.244
R6889 gnd.n2728 gnd.n2148 240.244
R6890 gnd.n2724 gnd.n2148 240.244
R6891 gnd.n2724 gnd.n2154 240.244
R6892 gnd.n2720 gnd.n2154 240.244
R6893 gnd.n2720 gnd.n2156 240.244
R6894 gnd.n2716 gnd.n2156 240.244
R6895 gnd.n2716 gnd.n2162 240.244
R6896 gnd.n2712 gnd.n2162 240.244
R6897 gnd.n2712 gnd.n2164 240.244
R6898 gnd.n2708 gnd.n2164 240.244
R6899 gnd.n2708 gnd.n2170 240.244
R6900 gnd.n2704 gnd.n2170 240.244
R6901 gnd.n2704 gnd.n2172 240.244
R6902 gnd.n2700 gnd.n2172 240.244
R6903 gnd.n2700 gnd.n2178 240.244
R6904 gnd.n2696 gnd.n2178 240.244
R6905 gnd.n2696 gnd.n2180 240.244
R6906 gnd.n2692 gnd.n2180 240.244
R6907 gnd.n2692 gnd.n2186 240.244
R6908 gnd.n2688 gnd.n2186 240.244
R6909 gnd.n2688 gnd.n2188 240.244
R6910 gnd.n2684 gnd.n2188 240.244
R6911 gnd.n2684 gnd.n2194 240.244
R6912 gnd.n2680 gnd.n2194 240.244
R6913 gnd.n2680 gnd.n2196 240.244
R6914 gnd.n2676 gnd.n2196 240.244
R6915 gnd.n2676 gnd.n2202 240.244
R6916 gnd.n2672 gnd.n2202 240.244
R6917 gnd.n2672 gnd.n2204 240.244
R6918 gnd.n2668 gnd.n2204 240.244
R6919 gnd.n2668 gnd.n2210 240.244
R6920 gnd.n2664 gnd.n2210 240.244
R6921 gnd.n2664 gnd.n2212 240.244
R6922 gnd.n2660 gnd.n2212 240.244
R6923 gnd.n2660 gnd.n2218 240.244
R6924 gnd.n2656 gnd.n2218 240.244
R6925 gnd.n2656 gnd.n2220 240.244
R6926 gnd.n2652 gnd.n2220 240.244
R6927 gnd.n2652 gnd.n2226 240.244
R6928 gnd.n2648 gnd.n2226 240.244
R6929 gnd.n2648 gnd.n2228 240.244
R6930 gnd.n2644 gnd.n2228 240.244
R6931 gnd.n2644 gnd.n2234 240.244
R6932 gnd.n2640 gnd.n2234 240.244
R6933 gnd.n2640 gnd.n2236 240.244
R6934 gnd.n2636 gnd.n2236 240.244
R6935 gnd.n2636 gnd.n2242 240.244
R6936 gnd.n2632 gnd.n2242 240.244
R6937 gnd.n2632 gnd.n2244 240.244
R6938 gnd.n2628 gnd.n2244 240.244
R6939 gnd.n2628 gnd.n2250 240.244
R6940 gnd.n2624 gnd.n2250 240.244
R6941 gnd.n2624 gnd.n2252 240.244
R6942 gnd.n2620 gnd.n2252 240.244
R6943 gnd.n2620 gnd.n2258 240.244
R6944 gnd.n2616 gnd.n2258 240.244
R6945 gnd.n2616 gnd.n2260 240.244
R6946 gnd.n2612 gnd.n2260 240.244
R6947 gnd.n2612 gnd.n2266 240.244
R6948 gnd.n2608 gnd.n2266 240.244
R6949 gnd.n2271 gnd.n2268 240.244
R6950 gnd.n2601 gnd.n2271 240.244
R6951 gnd.n2601 gnd.n2274 240.244
R6952 gnd.n2597 gnd.n2274 240.244
R6953 gnd.n2597 gnd.n2277 240.244
R6954 gnd.n2593 gnd.n2277 240.244
R6955 gnd.n2593 gnd.n2283 240.244
R6956 gnd.n2589 gnd.n2283 240.244
R6957 gnd.n2589 gnd.n2285 240.244
R6958 gnd.n2585 gnd.n2285 240.244
R6959 gnd.n2585 gnd.n2291 240.244
R6960 gnd.n2581 gnd.n2291 240.244
R6961 gnd.n2581 gnd.n2293 240.244
R6962 gnd.n2577 gnd.n2293 240.244
R6963 gnd.n2577 gnd.n2299 240.244
R6964 gnd.n2573 gnd.n2299 240.244
R6965 gnd.n2573 gnd.n2301 240.244
R6966 gnd.n2569 gnd.n2301 240.244
R6967 gnd.n2569 gnd.n2307 240.244
R6968 gnd.n2565 gnd.n2307 240.244
R6969 gnd.n2565 gnd.n2309 240.244
R6970 gnd.n2561 gnd.n2309 240.244
R6971 gnd.n2561 gnd.n2315 240.244
R6972 gnd.n2557 gnd.n2315 240.244
R6973 gnd.n2557 gnd.n2317 240.244
R6974 gnd.n2553 gnd.n2317 240.244
R6975 gnd.n2553 gnd.n2323 240.244
R6976 gnd.n2549 gnd.n2323 240.244
R6977 gnd.n2549 gnd.n2325 240.244
R6978 gnd.n2545 gnd.n2325 240.244
R6979 gnd.n2545 gnd.n2331 240.244
R6980 gnd.n2541 gnd.n2331 240.244
R6981 gnd.n2541 gnd.n2333 240.244
R6982 gnd.n2537 gnd.n2333 240.244
R6983 gnd.n2537 gnd.n2339 240.244
R6984 gnd.n2533 gnd.n2339 240.244
R6985 gnd.n2533 gnd.n2341 240.244
R6986 gnd.n2529 gnd.n2341 240.244
R6987 gnd.n2529 gnd.n2347 240.244
R6988 gnd.n2525 gnd.n2347 240.244
R6989 gnd.n2525 gnd.n2349 240.244
R6990 gnd.n2521 gnd.n2349 240.244
R6991 gnd.n2521 gnd.n2355 240.244
R6992 gnd.n2517 gnd.n2355 240.244
R6993 gnd.n2517 gnd.n2357 240.244
R6994 gnd.n2513 gnd.n2357 240.244
R6995 gnd.n2513 gnd.n2363 240.244
R6996 gnd.n2509 gnd.n2363 240.244
R6997 gnd.n2509 gnd.n2365 240.244
R6998 gnd.n2505 gnd.n2365 240.244
R6999 gnd.n2505 gnd.n2371 240.244
R7000 gnd.n2501 gnd.n2371 240.244
R7001 gnd.n2501 gnd.n2373 240.244
R7002 gnd.n2497 gnd.n2373 240.244
R7003 gnd.n2497 gnd.n2379 240.244
R7004 gnd.n2493 gnd.n2379 240.244
R7005 gnd.n2493 gnd.n2381 240.244
R7006 gnd.n2489 gnd.n2381 240.244
R7007 gnd.n2489 gnd.n2387 240.244
R7008 gnd.n2485 gnd.n2387 240.244
R7009 gnd.n2485 gnd.n2389 240.244
R7010 gnd.n2481 gnd.n2389 240.244
R7011 gnd.n2481 gnd.n2395 240.244
R7012 gnd.n2477 gnd.n2395 240.244
R7013 gnd.n2477 gnd.n2397 240.244
R7014 gnd.n2473 gnd.n2397 240.244
R7015 gnd.n2473 gnd.n2403 240.244
R7016 gnd.n2469 gnd.n2403 240.244
R7017 gnd.n2469 gnd.n2405 240.244
R7018 gnd.n2465 gnd.n2405 240.244
R7019 gnd.n2465 gnd.n2411 240.244
R7020 gnd.n2461 gnd.n2411 240.244
R7021 gnd.n2461 gnd.n2413 240.244
R7022 gnd.n2457 gnd.n2413 240.244
R7023 gnd.n2457 gnd.n2419 240.244
R7024 gnd.n2453 gnd.n2419 240.244
R7025 gnd.n2453 gnd.n2421 240.244
R7026 gnd.n2449 gnd.n2421 240.244
R7027 gnd.n2449 gnd.n2427 240.244
R7028 gnd.n2445 gnd.n2427 240.244
R7029 gnd.n2445 gnd.n2429 240.244
R7030 gnd.n2441 gnd.n2429 240.244
R7031 gnd.n2441 gnd.n2438 240.244
R7032 gnd.n2438 gnd.n398 240.244
R7033 gnd.n3603 gnd.n1809 240.244
R7034 gnd.n3603 gnd.n3596 240.244
R7035 gnd.n3596 gnd.n1756 240.244
R7036 gnd.n5375 gnd.n1756 240.244
R7037 gnd.n5375 gnd.n1751 240.244
R7038 gnd.n5383 gnd.n1751 240.244
R7039 gnd.n5383 gnd.n1752 240.244
R7040 gnd.n1752 gnd.n1721 240.244
R7041 gnd.n5425 gnd.n1721 240.244
R7042 gnd.n5425 gnd.n1715 240.244
R7043 gnd.n5433 gnd.n1715 240.244
R7044 gnd.n5433 gnd.n1717 240.244
R7045 gnd.n1717 gnd.n1657 240.244
R7046 gnd.n5487 gnd.n1657 240.244
R7047 gnd.n5487 gnd.n1653 240.244
R7048 gnd.n5493 gnd.n1653 240.244
R7049 gnd.n5494 gnd.n5493 240.244
R7050 gnd.n5495 gnd.n5494 240.244
R7051 gnd.n5495 gnd.n1648 240.244
R7052 gnd.n5536 gnd.n1648 240.244
R7053 gnd.n5536 gnd.n1649 240.244
R7054 gnd.n5532 gnd.n1649 240.244
R7055 gnd.n5532 gnd.n5531 240.244
R7056 gnd.n5531 gnd.n5530 240.244
R7057 gnd.n5530 gnd.n5503 240.244
R7058 gnd.n5526 gnd.n5503 240.244
R7059 gnd.n5526 gnd.n5525 240.244
R7060 gnd.n5525 gnd.n5524 240.244
R7061 gnd.n5524 gnd.n5509 240.244
R7062 gnd.n5519 gnd.n5509 240.244
R7063 gnd.n5519 gnd.n5516 240.244
R7064 gnd.n5516 gnd.n1228 240.244
R7065 gnd.n6165 gnd.n1228 240.244
R7066 gnd.n6165 gnd.n1224 240.244
R7067 gnd.n6171 gnd.n1224 240.244
R7068 gnd.n6171 gnd.n1215 240.244
R7069 gnd.n6181 gnd.n1215 240.244
R7070 gnd.n6181 gnd.n1211 240.244
R7071 gnd.n6187 gnd.n1211 240.244
R7072 gnd.n6187 gnd.n1201 240.244
R7073 gnd.n6197 gnd.n1201 240.244
R7074 gnd.n6197 gnd.n1197 240.244
R7075 gnd.n6203 gnd.n1197 240.244
R7076 gnd.n6203 gnd.n1187 240.244
R7077 gnd.n6213 gnd.n1187 240.244
R7078 gnd.n6213 gnd.n1183 240.244
R7079 gnd.n6219 gnd.n1183 240.244
R7080 gnd.n6219 gnd.n1172 240.244
R7081 gnd.n6229 gnd.n1172 240.244
R7082 gnd.n6229 gnd.n1168 240.244
R7083 gnd.n6235 gnd.n1168 240.244
R7084 gnd.n6235 gnd.n1158 240.244
R7085 gnd.n6245 gnd.n1158 240.244
R7086 gnd.n6245 gnd.n1154 240.244
R7087 gnd.n6251 gnd.n1154 240.244
R7088 gnd.n6251 gnd.n1142 240.244
R7089 gnd.n6261 gnd.n1142 240.244
R7090 gnd.n6261 gnd.n1138 240.244
R7091 gnd.n6267 gnd.n1138 240.244
R7092 gnd.n6267 gnd.n1128 240.244
R7093 gnd.n6277 gnd.n1128 240.244
R7094 gnd.n6277 gnd.n1124 240.244
R7095 gnd.n6283 gnd.n1124 240.244
R7096 gnd.n6283 gnd.n1114 240.244
R7097 gnd.n6293 gnd.n1114 240.244
R7098 gnd.n6293 gnd.n1110 240.244
R7099 gnd.n6299 gnd.n1110 240.244
R7100 gnd.n6299 gnd.n1101 240.244
R7101 gnd.n6309 gnd.n1101 240.244
R7102 gnd.n6309 gnd.n1097 240.244
R7103 gnd.n6315 gnd.n1097 240.244
R7104 gnd.n6315 gnd.n1087 240.244
R7105 gnd.n6325 gnd.n1087 240.244
R7106 gnd.n6325 gnd.n1083 240.244
R7107 gnd.n6331 gnd.n1083 240.244
R7108 gnd.n6331 gnd.n1069 240.244
R7109 gnd.n6347 gnd.n1069 240.244
R7110 gnd.n6347 gnd.n1064 240.244
R7111 gnd.n6355 gnd.n1064 240.244
R7112 gnd.n6355 gnd.n1065 240.244
R7113 gnd.n1065 gnd.n1031 240.244
R7114 gnd.n6405 gnd.n1031 240.244
R7115 gnd.n6405 gnd.n1026 240.244
R7116 gnd.n6413 gnd.n1026 240.244
R7117 gnd.n6413 gnd.n1027 240.244
R7118 gnd.n1027 gnd.n992 240.244
R7119 gnd.n6463 gnd.n992 240.244
R7120 gnd.n6463 gnd.n987 240.244
R7121 gnd.n6471 gnd.n987 240.244
R7122 gnd.n6471 gnd.n988 240.244
R7123 gnd.n988 gnd.n924 240.244
R7124 gnd.n6901 gnd.n924 240.244
R7125 gnd.n6901 gnd.n920 240.244
R7126 gnd.n6907 gnd.n920 240.244
R7127 gnd.n6907 gnd.n910 240.244
R7128 gnd.n6917 gnd.n910 240.244
R7129 gnd.n6917 gnd.n906 240.244
R7130 gnd.n6923 gnd.n906 240.244
R7131 gnd.n6923 gnd.n897 240.244
R7132 gnd.n6933 gnd.n897 240.244
R7133 gnd.n6933 gnd.n893 240.244
R7134 gnd.n6939 gnd.n893 240.244
R7135 gnd.n6939 gnd.n883 240.244
R7136 gnd.n6949 gnd.n883 240.244
R7137 gnd.n6949 gnd.n879 240.244
R7138 gnd.n6955 gnd.n879 240.244
R7139 gnd.n6955 gnd.n869 240.244
R7140 gnd.n6965 gnd.n869 240.244
R7141 gnd.n6965 gnd.n865 240.244
R7142 gnd.n6971 gnd.n865 240.244
R7143 gnd.n6971 gnd.n854 240.244
R7144 gnd.n6981 gnd.n854 240.244
R7145 gnd.n6981 gnd.n850 240.244
R7146 gnd.n6987 gnd.n850 240.244
R7147 gnd.n6987 gnd.n839 240.244
R7148 gnd.n6997 gnd.n839 240.244
R7149 gnd.n6997 gnd.n835 240.244
R7150 gnd.n7003 gnd.n835 240.244
R7151 gnd.n7003 gnd.n826 240.244
R7152 gnd.n7013 gnd.n826 240.244
R7153 gnd.n7013 gnd.n822 240.244
R7154 gnd.n7019 gnd.n822 240.244
R7155 gnd.n7019 gnd.n812 240.244
R7156 gnd.n7029 gnd.n812 240.244
R7157 gnd.n7029 gnd.n808 240.244
R7158 gnd.n7035 gnd.n808 240.244
R7159 gnd.n7035 gnd.n798 240.244
R7160 gnd.n7045 gnd.n798 240.244
R7161 gnd.n7045 gnd.n794 240.244
R7162 gnd.n7054 gnd.n794 240.244
R7163 gnd.n7054 gnd.n784 240.244
R7164 gnd.n7064 gnd.n784 240.244
R7165 gnd.n7065 gnd.n7064 240.244
R7166 gnd.n7065 gnd.n746 240.244
R7167 gnd.n779 gnd.n746 240.244
R7168 gnd.n7076 gnd.n779 240.244
R7169 gnd.n7076 gnd.n780 240.244
R7170 gnd.n780 gnd.n570 240.244
R7171 gnd.n7276 gnd.n570 240.244
R7172 gnd.n7277 gnd.n7276 240.244
R7173 gnd.n7277 gnd.n565 240.244
R7174 gnd.n7300 gnd.n565 240.244
R7175 gnd.n7300 gnd.n566 240.244
R7176 gnd.n7296 gnd.n566 240.244
R7177 gnd.n7296 gnd.n7295 240.244
R7178 gnd.n7295 gnd.n7294 240.244
R7179 gnd.n7294 gnd.n7285 240.244
R7180 gnd.n7285 gnd.n502 240.244
R7181 gnd.n7373 gnd.n502 240.244
R7182 gnd.n7374 gnd.n7373 240.244
R7183 gnd.n7375 gnd.n7374 240.244
R7184 gnd.n7375 gnd.n497 240.244
R7185 gnd.n7392 gnd.n497 240.244
R7186 gnd.n7392 gnd.n498 240.244
R7187 gnd.n7388 gnd.n498 240.244
R7188 gnd.n7388 gnd.n7387 240.244
R7189 gnd.n7387 gnd.n7386 240.244
R7190 gnd.n7386 gnd.n437 240.244
R7191 gnd.n7459 gnd.n437 240.244
R7192 gnd.n7459 gnd.n432 240.244
R7193 gnd.n7469 gnd.n432 240.244
R7194 gnd.n7469 gnd.n433 240.244
R7195 gnd.n433 gnd.n402 240.244
R7196 gnd.n7510 gnd.n402 240.244
R7197 gnd.n7511 gnd.n7510 240.244
R7198 gnd.n7511 gnd.n396 240.244
R7199 gnd.n7517 gnd.n396 240.244
R7200 gnd.n2946 gnd.n1933 240.244
R7201 gnd.n2950 gnd.n1933 240.244
R7202 gnd.n2950 gnd.n1929 240.244
R7203 gnd.n2956 gnd.n1929 240.244
R7204 gnd.n2956 gnd.n1927 240.244
R7205 gnd.n2960 gnd.n1927 240.244
R7206 gnd.n2960 gnd.n1923 240.244
R7207 gnd.n2966 gnd.n1923 240.244
R7208 gnd.n2966 gnd.n1921 240.244
R7209 gnd.n2970 gnd.n1921 240.244
R7210 gnd.n2970 gnd.n1917 240.244
R7211 gnd.n2976 gnd.n1917 240.244
R7212 gnd.n2976 gnd.n1915 240.244
R7213 gnd.n2980 gnd.n1915 240.244
R7214 gnd.n2980 gnd.n1911 240.244
R7215 gnd.n2986 gnd.n1911 240.244
R7216 gnd.n2986 gnd.n1909 240.244
R7217 gnd.n2990 gnd.n1909 240.244
R7218 gnd.n2990 gnd.n1905 240.244
R7219 gnd.n2996 gnd.n1905 240.244
R7220 gnd.n2996 gnd.n1903 240.244
R7221 gnd.n3000 gnd.n1903 240.244
R7222 gnd.n3000 gnd.n1899 240.244
R7223 gnd.n3006 gnd.n1899 240.244
R7224 gnd.n3006 gnd.n1897 240.244
R7225 gnd.n3010 gnd.n1897 240.244
R7226 gnd.n3010 gnd.n1893 240.244
R7227 gnd.n3016 gnd.n1893 240.244
R7228 gnd.n3016 gnd.n1891 240.244
R7229 gnd.n3020 gnd.n1891 240.244
R7230 gnd.n3020 gnd.n1887 240.244
R7231 gnd.n3026 gnd.n1887 240.244
R7232 gnd.n3026 gnd.n1885 240.244
R7233 gnd.n3030 gnd.n1885 240.244
R7234 gnd.n3030 gnd.n1881 240.244
R7235 gnd.n3036 gnd.n1881 240.244
R7236 gnd.n3036 gnd.n1879 240.244
R7237 gnd.n3040 gnd.n1879 240.244
R7238 gnd.n3040 gnd.n1875 240.244
R7239 gnd.n3046 gnd.n1875 240.244
R7240 gnd.n3046 gnd.n1873 240.244
R7241 gnd.n3050 gnd.n1873 240.244
R7242 gnd.n3050 gnd.n1869 240.244
R7243 gnd.n3056 gnd.n1869 240.244
R7244 gnd.n3056 gnd.n1867 240.244
R7245 gnd.n3060 gnd.n1867 240.244
R7246 gnd.n3060 gnd.n1863 240.244
R7247 gnd.n3066 gnd.n1863 240.244
R7248 gnd.n3066 gnd.n1861 240.244
R7249 gnd.n3070 gnd.n1861 240.244
R7250 gnd.n3070 gnd.n1857 240.244
R7251 gnd.n3076 gnd.n1857 240.244
R7252 gnd.n3076 gnd.n1855 240.244
R7253 gnd.n3080 gnd.n1855 240.244
R7254 gnd.n3080 gnd.n1851 240.244
R7255 gnd.n3086 gnd.n1851 240.244
R7256 gnd.n3086 gnd.n1849 240.244
R7257 gnd.n3090 gnd.n1849 240.244
R7258 gnd.n3090 gnd.n1845 240.244
R7259 gnd.n3096 gnd.n1845 240.244
R7260 gnd.n3096 gnd.n1843 240.244
R7261 gnd.n3100 gnd.n1843 240.244
R7262 gnd.n3100 gnd.n1839 240.244
R7263 gnd.n3106 gnd.n1839 240.244
R7264 gnd.n3106 gnd.n1837 240.244
R7265 gnd.n3110 gnd.n1837 240.244
R7266 gnd.n3110 gnd.n1833 240.244
R7267 gnd.n3116 gnd.n1833 240.244
R7268 gnd.n3116 gnd.n1831 240.244
R7269 gnd.n3120 gnd.n1831 240.244
R7270 gnd.n3120 gnd.n1827 240.244
R7271 gnd.n3126 gnd.n1827 240.244
R7272 gnd.n3126 gnd.n1825 240.244
R7273 gnd.n3130 gnd.n1825 240.244
R7274 gnd.n3130 gnd.n1821 240.244
R7275 gnd.n3136 gnd.n1821 240.244
R7276 gnd.n3136 gnd.n1819 240.244
R7277 gnd.n3140 gnd.n1819 240.244
R7278 gnd.n3140 gnd.n1815 240.244
R7279 gnd.n3146 gnd.n1815 240.244
R7280 gnd.n3146 gnd.n1813 240.244
R7281 gnd.n5316 gnd.n1813 240.244
R7282 gnd.n5316 gnd.n1808 240.244
R7283 gnd.n5322 gnd.n1808 240.244
R7284 gnd.n1452 gnd.n1230 240.244
R7285 gnd.n1452 gnd.n1223 240.244
R7286 gnd.n5747 gnd.n1223 240.244
R7287 gnd.n5747 gnd.n1217 240.244
R7288 gnd.n1449 gnd.n1217 240.244
R7289 gnd.n1449 gnd.n1210 240.244
R7290 gnd.n5754 gnd.n1210 240.244
R7291 gnd.n5754 gnd.n1203 240.244
R7292 gnd.n1446 gnd.n1203 240.244
R7293 gnd.n1446 gnd.n1195 240.244
R7294 gnd.n5761 gnd.n1195 240.244
R7295 gnd.n5761 gnd.n1188 240.244
R7296 gnd.n1443 gnd.n1188 240.244
R7297 gnd.n1443 gnd.n1181 240.244
R7298 gnd.n5768 gnd.n1181 240.244
R7299 gnd.n5768 gnd.n1173 240.244
R7300 gnd.n1440 gnd.n1173 240.244
R7301 gnd.n1440 gnd.n1166 240.244
R7302 gnd.n5775 gnd.n1166 240.244
R7303 gnd.n5775 gnd.n1159 240.244
R7304 gnd.n6021 gnd.n1159 240.244
R7305 gnd.n6021 gnd.n1152 240.244
R7306 gnd.n5780 gnd.n1152 240.244
R7307 gnd.n5780 gnd.n1144 240.244
R7308 gnd.n5781 gnd.n1144 240.244
R7309 gnd.n5781 gnd.n1136 240.244
R7310 gnd.n5784 gnd.n1136 240.244
R7311 gnd.n5784 gnd.n1129 240.244
R7312 gnd.n5785 gnd.n1129 240.244
R7313 gnd.n5785 gnd.n1122 240.244
R7314 gnd.n5788 gnd.n1122 240.244
R7315 gnd.n5788 gnd.n1115 240.244
R7316 gnd.n5789 gnd.n1115 240.244
R7317 gnd.n5789 gnd.n1109 240.244
R7318 gnd.n5792 gnd.n1109 240.244
R7319 gnd.n5792 gnd.n1103 240.244
R7320 gnd.n5793 gnd.n1103 240.244
R7321 gnd.n5793 gnd.n1096 240.244
R7322 gnd.n5796 gnd.n1096 240.244
R7323 gnd.n5796 gnd.n1089 240.244
R7324 gnd.n5797 gnd.n1089 240.244
R7325 gnd.n5797 gnd.n1081 240.244
R7326 gnd.n5971 gnd.n1081 240.244
R7327 gnd.n5971 gnd.n1070 240.244
R7328 gnd.n5972 gnd.n1070 240.244
R7329 gnd.n5972 gnd.n1061 240.244
R7330 gnd.n5975 gnd.n1061 240.244
R7331 gnd.n5976 gnd.n5975 240.244
R7332 gnd.n5976 gnd.n1033 240.244
R7333 gnd.n1033 gnd.n1022 240.244
R7334 gnd.n6415 gnd.n1022 240.244
R7335 gnd.n6415 gnd.n1017 240.244
R7336 gnd.n6422 gnd.n1017 240.244
R7337 gnd.n6422 gnd.n994 240.244
R7338 gnd.n994 gnd.n982 240.244
R7339 gnd.n6473 gnd.n982 240.244
R7340 gnd.n6473 gnd.n983 240.244
R7341 gnd.n983 gnd.n979 240.244
R7342 gnd.n979 gnd.n926 240.244
R7343 gnd.n6480 gnd.n926 240.244
R7344 gnd.n6480 gnd.n918 240.244
R7345 gnd.n941 gnd.n918 240.244
R7346 gnd.n941 gnd.n911 240.244
R7347 gnd.n6487 gnd.n911 240.244
R7348 gnd.n6487 gnd.n904 240.244
R7349 gnd.n954 gnd.n904 240.244
R7350 gnd.n954 gnd.n898 240.244
R7351 gnd.n6494 gnd.n898 240.244
R7352 gnd.n6494 gnd.n892 240.244
R7353 gnd.n6856 gnd.n892 240.244
R7354 gnd.n6856 gnd.n885 240.244
R7355 gnd.n6499 gnd.n885 240.244
R7356 gnd.n6499 gnd.n878 240.244
R7357 gnd.n6500 gnd.n878 240.244
R7358 gnd.n6500 gnd.n871 240.244
R7359 gnd.n6503 gnd.n871 240.244
R7360 gnd.n6503 gnd.n863 240.244
R7361 gnd.n6504 gnd.n863 240.244
R7362 gnd.n6504 gnd.n856 240.244
R7363 gnd.n6507 gnd.n856 240.244
R7364 gnd.n6507 gnd.n848 240.244
R7365 gnd.n6793 gnd.n848 240.244
R7366 gnd.n6793 gnd.n841 240.244
R7367 gnd.n6796 gnd.n841 240.244
R7368 gnd.n6796 gnd.n834 240.244
R7369 gnd.n6797 gnd.n834 240.244
R7370 gnd.n6797 gnd.n828 240.244
R7371 gnd.n6800 gnd.n828 240.244
R7372 gnd.n6800 gnd.n821 240.244
R7373 gnd.n6801 gnd.n821 240.244
R7374 gnd.n6801 gnd.n814 240.244
R7375 gnd.n6804 gnd.n814 240.244
R7376 gnd.n6804 gnd.n806 240.244
R7377 gnd.n6805 gnd.n806 240.244
R7378 gnd.n6805 gnd.n799 240.244
R7379 gnd.n6808 gnd.n799 240.244
R7380 gnd.n6808 gnd.n793 240.244
R7381 gnd.n6809 gnd.n793 240.244
R7382 gnd.n6809 gnd.n786 240.244
R7383 gnd.n786 gnd.n748 240.244
R7384 gnd.n7093 gnd.n748 240.244
R7385 gnd.n5737 gnd.n1455 240.244
R7386 gnd.n5737 gnd.n1471 240.244
R7387 gnd.n1475 gnd.n1474 240.244
R7388 gnd.n1477 gnd.n1476 240.244
R7389 gnd.n5611 gnd.n5610 240.244
R7390 gnd.n5622 gnd.n5621 240.244
R7391 gnd.n5624 gnd.n5623 240.244
R7392 gnd.n5634 gnd.n5633 240.244
R7393 gnd.n5645 gnd.n5644 240.244
R7394 gnd.n5647 gnd.n5646 240.244
R7395 gnd.n5657 gnd.n5656 240.244
R7396 gnd.n5668 gnd.n5667 240.244
R7397 gnd.n5674 gnd.n5669 240.244
R7398 gnd.n1468 gnd.n1235 240.244
R7399 gnd.n6163 gnd.n1222 240.244
R7400 gnd.n6173 gnd.n1222 240.244
R7401 gnd.n6173 gnd.n1218 240.244
R7402 gnd.n6179 gnd.n1218 240.244
R7403 gnd.n6179 gnd.n1208 240.244
R7404 gnd.n6189 gnd.n1208 240.244
R7405 gnd.n6189 gnd.n1204 240.244
R7406 gnd.n6195 gnd.n1204 240.244
R7407 gnd.n6195 gnd.n1193 240.244
R7408 gnd.n6205 gnd.n1193 240.244
R7409 gnd.n6205 gnd.n1189 240.244
R7410 gnd.n6211 gnd.n1189 240.244
R7411 gnd.n6211 gnd.n1179 240.244
R7412 gnd.n6221 gnd.n1179 240.244
R7413 gnd.n6221 gnd.n1175 240.244
R7414 gnd.n6227 gnd.n1175 240.244
R7415 gnd.n6227 gnd.n1165 240.244
R7416 gnd.n6237 gnd.n1165 240.244
R7417 gnd.n6237 gnd.n1161 240.244
R7418 gnd.n6243 gnd.n1161 240.244
R7419 gnd.n6243 gnd.n1150 240.244
R7420 gnd.n6253 gnd.n1150 240.244
R7421 gnd.n6253 gnd.n1146 240.244
R7422 gnd.n6259 gnd.n1146 240.244
R7423 gnd.n6259 gnd.n1135 240.244
R7424 gnd.n6269 gnd.n1135 240.244
R7425 gnd.n6269 gnd.n1131 240.244
R7426 gnd.n6275 gnd.n1131 240.244
R7427 gnd.n6275 gnd.n1121 240.244
R7428 gnd.n6285 gnd.n1121 240.244
R7429 gnd.n6285 gnd.n1117 240.244
R7430 gnd.n6291 gnd.n1117 240.244
R7431 gnd.n6291 gnd.n1108 240.244
R7432 gnd.n6301 gnd.n1108 240.244
R7433 gnd.n6301 gnd.n1104 240.244
R7434 gnd.n6307 gnd.n1104 240.244
R7435 gnd.n6307 gnd.n1094 240.244
R7436 gnd.n6317 gnd.n1094 240.244
R7437 gnd.n6317 gnd.n1090 240.244
R7438 gnd.n6323 gnd.n1090 240.244
R7439 gnd.n6323 gnd.n1078 240.244
R7440 gnd.n6333 gnd.n1078 240.244
R7441 gnd.n6333 gnd.n1072 240.244
R7442 gnd.n6345 gnd.n1072 240.244
R7443 gnd.n6345 gnd.n1073 240.244
R7444 gnd.n1073 gnd.n1063 240.244
R7445 gnd.n6338 gnd.n1063 240.244
R7446 gnd.n6338 gnd.n1035 240.244
R7447 gnd.n6403 gnd.n1035 240.244
R7448 gnd.n6403 gnd.n1036 240.244
R7449 gnd.n1036 gnd.n1025 240.244
R7450 gnd.n6396 gnd.n1025 240.244
R7451 gnd.n6396 gnd.n996 240.244
R7452 gnd.n6461 gnd.n996 240.244
R7453 gnd.n6461 gnd.n997 240.244
R7454 gnd.n997 gnd.n986 240.244
R7455 gnd.n1002 gnd.n986 240.244
R7456 gnd.n6450 gnd.n1002 240.244
R7457 gnd.n6450 gnd.n928 240.244
R7458 gnd.n928 gnd.n917 240.244
R7459 gnd.n6909 gnd.n917 240.244
R7460 gnd.n6909 gnd.n913 240.244
R7461 gnd.n6915 gnd.n913 240.244
R7462 gnd.n6915 gnd.n903 240.244
R7463 gnd.n6925 gnd.n903 240.244
R7464 gnd.n6925 gnd.n899 240.244
R7465 gnd.n6931 gnd.n899 240.244
R7466 gnd.n6931 gnd.n890 240.244
R7467 gnd.n6941 gnd.n890 240.244
R7468 gnd.n6941 gnd.n886 240.244
R7469 gnd.n6947 gnd.n886 240.244
R7470 gnd.n6947 gnd.n876 240.244
R7471 gnd.n6957 gnd.n876 240.244
R7472 gnd.n6957 gnd.n872 240.244
R7473 gnd.n6963 gnd.n872 240.244
R7474 gnd.n6963 gnd.n861 240.244
R7475 gnd.n6973 gnd.n861 240.244
R7476 gnd.n6973 gnd.n857 240.244
R7477 gnd.n6979 gnd.n857 240.244
R7478 gnd.n6979 gnd.n847 240.244
R7479 gnd.n6989 gnd.n847 240.244
R7480 gnd.n6989 gnd.n843 240.244
R7481 gnd.n6995 gnd.n843 240.244
R7482 gnd.n6995 gnd.n833 240.244
R7483 gnd.n7005 gnd.n833 240.244
R7484 gnd.n7005 gnd.n829 240.244
R7485 gnd.n7011 gnd.n829 240.244
R7486 gnd.n7011 gnd.n819 240.244
R7487 gnd.n7021 gnd.n819 240.244
R7488 gnd.n7021 gnd.n815 240.244
R7489 gnd.n7027 gnd.n815 240.244
R7490 gnd.n7027 gnd.n804 240.244
R7491 gnd.n7037 gnd.n804 240.244
R7492 gnd.n7037 gnd.n800 240.244
R7493 gnd.n7043 gnd.n800 240.244
R7494 gnd.n7043 gnd.n791 240.244
R7495 gnd.n7056 gnd.n791 240.244
R7496 gnd.n7056 gnd.n787 240.244
R7497 gnd.n7062 gnd.n787 240.244
R7498 gnd.n7062 gnd.n743 240.244
R7499 gnd.n7095 gnd.n743 240.244
R7500 gnd.n754 gnd.n753 240.244
R7501 gnd.n760 gnd.n757 240.244
R7502 gnd.n7081 gnd.n7080 240.244
R7503 gnd.n681 gnd.n680 240.244
R7504 gnd.n763 gnd.n682 240.244
R7505 gnd.n692 gnd.n691 240.244
R7506 gnd.n765 gnd.n701 240.244
R7507 gnd.n768 gnd.n702 240.244
R7508 gnd.n710 gnd.n709 240.244
R7509 gnd.n770 gnd.n719 240.244
R7510 gnd.n773 gnd.n720 240.244
R7511 gnd.n728 gnd.n727 240.244
R7512 gnd.n775 gnd.n728 240.244
R7513 gnd.n739 gnd.n738 240.244
R7514 gnd.n1334 gnd.n1333 240.132
R7515 gnd.n6523 gnd.n6522 240.132
R7516 gnd.n2939 gnd.n1934 225.874
R7517 gnd.n2939 gnd.n2938 225.874
R7518 gnd.n2938 gnd.n2937 225.874
R7519 gnd.n2937 gnd.n1939 225.874
R7520 gnd.n2931 gnd.n1939 225.874
R7521 gnd.n2931 gnd.n2930 225.874
R7522 gnd.n2930 gnd.n2929 225.874
R7523 gnd.n2929 gnd.n1947 225.874
R7524 gnd.n2923 gnd.n1947 225.874
R7525 gnd.n2923 gnd.n2922 225.874
R7526 gnd.n2922 gnd.n2921 225.874
R7527 gnd.n2921 gnd.n1955 225.874
R7528 gnd.n2915 gnd.n1955 225.874
R7529 gnd.n2915 gnd.n2914 225.874
R7530 gnd.n2914 gnd.n2913 225.874
R7531 gnd.n2913 gnd.n1963 225.874
R7532 gnd.n2907 gnd.n1963 225.874
R7533 gnd.n2907 gnd.n2906 225.874
R7534 gnd.n2906 gnd.n2905 225.874
R7535 gnd.n2905 gnd.n1971 225.874
R7536 gnd.n2899 gnd.n1971 225.874
R7537 gnd.n2899 gnd.n2898 225.874
R7538 gnd.n2898 gnd.n2897 225.874
R7539 gnd.n2897 gnd.n1979 225.874
R7540 gnd.n2891 gnd.n1979 225.874
R7541 gnd.n2891 gnd.n2890 225.874
R7542 gnd.n2890 gnd.n2889 225.874
R7543 gnd.n2889 gnd.n1987 225.874
R7544 gnd.n2883 gnd.n1987 225.874
R7545 gnd.n2883 gnd.n2882 225.874
R7546 gnd.n2882 gnd.n2881 225.874
R7547 gnd.n2881 gnd.n1995 225.874
R7548 gnd.n2875 gnd.n1995 225.874
R7549 gnd.n2875 gnd.n2874 225.874
R7550 gnd.n2874 gnd.n2873 225.874
R7551 gnd.n2873 gnd.n2003 225.874
R7552 gnd.n2867 gnd.n2003 225.874
R7553 gnd.n2867 gnd.n2866 225.874
R7554 gnd.n2866 gnd.n2865 225.874
R7555 gnd.n2865 gnd.n2011 225.874
R7556 gnd.n2859 gnd.n2011 225.874
R7557 gnd.n2859 gnd.n2858 225.874
R7558 gnd.n2858 gnd.n2857 225.874
R7559 gnd.n2857 gnd.n2019 225.874
R7560 gnd.n2851 gnd.n2019 225.874
R7561 gnd.n2851 gnd.n2850 225.874
R7562 gnd.n2850 gnd.n2849 225.874
R7563 gnd.n2849 gnd.n2027 225.874
R7564 gnd.n2843 gnd.n2027 225.874
R7565 gnd.n2843 gnd.n2842 225.874
R7566 gnd.n2842 gnd.n2841 225.874
R7567 gnd.n2841 gnd.n2035 225.874
R7568 gnd.n2835 gnd.n2035 225.874
R7569 gnd.n2835 gnd.n2834 225.874
R7570 gnd.n2834 gnd.n2833 225.874
R7571 gnd.n2833 gnd.n2043 225.874
R7572 gnd.n2827 gnd.n2043 225.874
R7573 gnd.n2827 gnd.n2826 225.874
R7574 gnd.n2826 gnd.n2825 225.874
R7575 gnd.n2825 gnd.n2051 225.874
R7576 gnd.n2819 gnd.n2051 225.874
R7577 gnd.n2819 gnd.n2818 225.874
R7578 gnd.n2818 gnd.n2817 225.874
R7579 gnd.n2817 gnd.n2059 225.874
R7580 gnd.n2811 gnd.n2059 225.874
R7581 gnd.n2811 gnd.n2810 225.874
R7582 gnd.n2810 gnd.n2809 225.874
R7583 gnd.n2809 gnd.n2067 225.874
R7584 gnd.n2803 gnd.n2067 225.874
R7585 gnd.n2803 gnd.n2802 225.874
R7586 gnd.n2802 gnd.n2801 225.874
R7587 gnd.n2801 gnd.n2075 225.874
R7588 gnd.n2795 gnd.n2075 225.874
R7589 gnd.n2795 gnd.n2794 225.874
R7590 gnd.n2794 gnd.n2793 225.874
R7591 gnd.n2793 gnd.n2083 225.874
R7592 gnd.n2787 gnd.n2083 225.874
R7593 gnd.n2787 gnd.n2786 225.874
R7594 gnd.n2786 gnd.n2785 225.874
R7595 gnd.n2785 gnd.n2091 225.874
R7596 gnd.n2779 gnd.n2091 225.874
R7597 gnd.n2779 gnd.n2778 225.874
R7598 gnd.n2778 gnd.n2777 225.874
R7599 gnd.n2777 gnd.n2099 225.874
R7600 gnd.n2771 gnd.n2099 225.874
R7601 gnd.n2771 gnd.n2770 225.874
R7602 gnd.n2770 gnd.n2769 225.874
R7603 gnd.n2769 gnd.n2107 225.874
R7604 gnd.n2763 gnd.n2107 225.874
R7605 gnd.n2763 gnd.n2762 225.874
R7606 gnd.n2762 gnd.n2761 225.874
R7607 gnd.n2761 gnd.n2115 225.874
R7608 gnd.n2755 gnd.n2115 225.874
R7609 gnd.n2755 gnd.n2754 225.874
R7610 gnd.n2754 gnd.n2753 225.874
R7611 gnd.n2753 gnd.n2123 225.874
R7612 gnd.n2747 gnd.n2123 225.874
R7613 gnd.n2747 gnd.n2746 225.874
R7614 gnd.n2746 gnd.n2745 225.874
R7615 gnd.n2745 gnd.n2131 225.874
R7616 gnd.n2739 gnd.n2131 225.874
R7617 gnd.n2739 gnd.n2738 225.874
R7618 gnd.n2738 gnd.n2737 225.874
R7619 gnd.n2737 gnd.n2139 225.874
R7620 gnd.n2731 gnd.n2139 225.874
R7621 gnd.n2731 gnd.n2730 225.874
R7622 gnd.n2730 gnd.n2729 225.874
R7623 gnd.n2729 gnd.n2147 225.874
R7624 gnd.n2723 gnd.n2147 225.874
R7625 gnd.n2723 gnd.n2722 225.874
R7626 gnd.n2722 gnd.n2721 225.874
R7627 gnd.n2721 gnd.n2155 225.874
R7628 gnd.n2715 gnd.n2155 225.874
R7629 gnd.n2715 gnd.n2714 225.874
R7630 gnd.n2714 gnd.n2713 225.874
R7631 gnd.n2713 gnd.n2163 225.874
R7632 gnd.n2707 gnd.n2163 225.874
R7633 gnd.n2707 gnd.n2706 225.874
R7634 gnd.n2706 gnd.n2705 225.874
R7635 gnd.n2705 gnd.n2171 225.874
R7636 gnd.n2699 gnd.n2171 225.874
R7637 gnd.n2699 gnd.n2698 225.874
R7638 gnd.n2698 gnd.n2697 225.874
R7639 gnd.n2697 gnd.n2179 225.874
R7640 gnd.n2691 gnd.n2179 225.874
R7641 gnd.n2691 gnd.n2690 225.874
R7642 gnd.n2690 gnd.n2689 225.874
R7643 gnd.n2689 gnd.n2187 225.874
R7644 gnd.n2683 gnd.n2187 225.874
R7645 gnd.n2683 gnd.n2682 225.874
R7646 gnd.n2682 gnd.n2681 225.874
R7647 gnd.n2681 gnd.n2195 225.874
R7648 gnd.n2675 gnd.n2195 225.874
R7649 gnd.n2675 gnd.n2674 225.874
R7650 gnd.n2674 gnd.n2673 225.874
R7651 gnd.n2673 gnd.n2203 225.874
R7652 gnd.n2667 gnd.n2203 225.874
R7653 gnd.n2667 gnd.n2666 225.874
R7654 gnd.n2666 gnd.n2665 225.874
R7655 gnd.n2665 gnd.n2211 225.874
R7656 gnd.n2659 gnd.n2211 225.874
R7657 gnd.n2659 gnd.n2658 225.874
R7658 gnd.n2658 gnd.n2657 225.874
R7659 gnd.n2657 gnd.n2219 225.874
R7660 gnd.n2651 gnd.n2219 225.874
R7661 gnd.n2651 gnd.n2650 225.874
R7662 gnd.n2650 gnd.n2649 225.874
R7663 gnd.n2649 gnd.n2227 225.874
R7664 gnd.n2643 gnd.n2227 225.874
R7665 gnd.n2643 gnd.n2642 225.874
R7666 gnd.n2642 gnd.n2641 225.874
R7667 gnd.n2641 gnd.n2235 225.874
R7668 gnd.n2635 gnd.n2235 225.874
R7669 gnd.n2635 gnd.n2634 225.874
R7670 gnd.n2634 gnd.n2633 225.874
R7671 gnd.n2633 gnd.n2243 225.874
R7672 gnd.n2627 gnd.n2243 225.874
R7673 gnd.n2627 gnd.n2626 225.874
R7674 gnd.n2626 gnd.n2625 225.874
R7675 gnd.n2625 gnd.n2251 225.874
R7676 gnd.n2619 gnd.n2251 225.874
R7677 gnd.n2619 gnd.n2618 225.874
R7678 gnd.n2618 gnd.n2617 225.874
R7679 gnd.n2617 gnd.n2259 225.874
R7680 gnd.n2611 gnd.n2259 225.874
R7681 gnd.n2611 gnd.n2610 225.874
R7682 gnd.n2610 gnd.n2609 225.874
R7683 gnd.n4406 gnd.t93 224.174
R7684 gnd.n3884 gnd.t196 224.174
R7685 gnd.n640 gnd.n583 199.319
R7686 gnd.n640 gnd.n584 199.319
R7687 gnd.n1299 gnd.n1298 199.319
R7688 gnd.n1514 gnd.n1299 199.319
R7689 gnd.n1335 gnd.n1332 186.49
R7690 gnd.n6524 gnd.n6521 186.49
R7691 gnd.n5181 gnd.n5180 185
R7692 gnd.n5179 gnd.n5178 185
R7693 gnd.n5158 gnd.n5157 185
R7694 gnd.n5173 gnd.n5172 185
R7695 gnd.n5171 gnd.n5170 185
R7696 gnd.n5162 gnd.n5161 185
R7697 gnd.n5165 gnd.n5164 185
R7698 gnd.n5149 gnd.n5148 185
R7699 gnd.n5147 gnd.n5146 185
R7700 gnd.n5126 gnd.n5125 185
R7701 gnd.n5141 gnd.n5140 185
R7702 gnd.n5139 gnd.n5138 185
R7703 gnd.n5130 gnd.n5129 185
R7704 gnd.n5133 gnd.n5132 185
R7705 gnd.n5117 gnd.n5116 185
R7706 gnd.n5115 gnd.n5114 185
R7707 gnd.n5094 gnd.n5093 185
R7708 gnd.n5109 gnd.n5108 185
R7709 gnd.n5107 gnd.n5106 185
R7710 gnd.n5098 gnd.n5097 185
R7711 gnd.n5101 gnd.n5100 185
R7712 gnd.n5086 gnd.n5085 185
R7713 gnd.n5084 gnd.n5083 185
R7714 gnd.n5063 gnd.n5062 185
R7715 gnd.n5078 gnd.n5077 185
R7716 gnd.n5076 gnd.n5075 185
R7717 gnd.n5067 gnd.n5066 185
R7718 gnd.n5070 gnd.n5069 185
R7719 gnd.n5054 gnd.n5053 185
R7720 gnd.n5052 gnd.n5051 185
R7721 gnd.n5031 gnd.n5030 185
R7722 gnd.n5046 gnd.n5045 185
R7723 gnd.n5044 gnd.n5043 185
R7724 gnd.n5035 gnd.n5034 185
R7725 gnd.n5038 gnd.n5037 185
R7726 gnd.n5022 gnd.n5021 185
R7727 gnd.n5020 gnd.n5019 185
R7728 gnd.n4999 gnd.n4998 185
R7729 gnd.n5014 gnd.n5013 185
R7730 gnd.n5012 gnd.n5011 185
R7731 gnd.n5003 gnd.n5002 185
R7732 gnd.n5006 gnd.n5005 185
R7733 gnd.n4990 gnd.n4989 185
R7734 gnd.n4988 gnd.n4987 185
R7735 gnd.n4967 gnd.n4966 185
R7736 gnd.n4982 gnd.n4981 185
R7737 gnd.n4980 gnd.n4979 185
R7738 gnd.n4971 gnd.n4970 185
R7739 gnd.n4974 gnd.n4973 185
R7740 gnd.n4959 gnd.n4958 185
R7741 gnd.n4957 gnd.n4956 185
R7742 gnd.n4936 gnd.n4935 185
R7743 gnd.n4951 gnd.n4950 185
R7744 gnd.n4949 gnd.n4948 185
R7745 gnd.n4940 gnd.n4939 185
R7746 gnd.n4943 gnd.n4942 185
R7747 gnd.n4407 gnd.t92 178.987
R7748 gnd.n3885 gnd.t197 178.987
R7749 gnd.n1 gnd.t64 170.774
R7750 gnd.n9 gnd.t82 170.103
R7751 gnd.n8 gnd.t415 170.103
R7752 gnd.n7 gnd.t13 170.103
R7753 gnd.n6 gnd.t84 170.103
R7754 gnd.n5 gnd.t53 170.103
R7755 gnd.n4 gnd.t74 170.103
R7756 gnd.n3 gnd.t72 170.103
R7757 gnd.n2 gnd.t58 170.103
R7758 gnd.n1 gnd.t86 170.103
R7759 gnd.n6783 gnd.n6782 163.367
R7760 gnd.n6780 gnd.n6534 163.367
R7761 gnd.n6776 gnd.n6775 163.367
R7762 gnd.n6773 gnd.n6537 163.367
R7763 gnd.n6769 gnd.n6768 163.367
R7764 gnd.n6766 gnd.n6540 163.367
R7765 gnd.n6762 gnd.n6761 163.367
R7766 gnd.n6759 gnd.n6543 163.367
R7767 gnd.n6755 gnd.n6754 163.367
R7768 gnd.n6752 gnd.n6546 163.367
R7769 gnd.n6748 gnd.n6747 163.367
R7770 gnd.n6745 gnd.n6549 163.367
R7771 gnd.n6741 gnd.n6740 163.367
R7772 gnd.n6738 gnd.n6552 163.367
R7773 gnd.n6733 gnd.n6732 163.367
R7774 gnd.n6730 gnd.n6728 163.367
R7775 gnd.n6725 gnd.n6724 163.367
R7776 gnd.n6722 gnd.n6558 163.367
R7777 gnd.n6717 gnd.n6716 163.367
R7778 gnd.n6714 gnd.n6563 163.367
R7779 gnd.n6710 gnd.n6709 163.367
R7780 gnd.n6707 gnd.n6566 163.367
R7781 gnd.n6703 gnd.n6702 163.367
R7782 gnd.n6700 gnd.n6569 163.367
R7783 gnd.n6696 gnd.n6695 163.367
R7784 gnd.n6693 gnd.n6572 163.367
R7785 gnd.n6689 gnd.n6688 163.367
R7786 gnd.n6686 gnd.n6575 163.367
R7787 gnd.n6682 gnd.n6681 163.367
R7788 gnd.n6679 gnd.n6578 163.367
R7789 gnd.n6675 gnd.n6674 163.367
R7790 gnd.n6672 gnd.n6581 163.367
R7791 gnd.n6032 gnd.n6031 163.367
R7792 gnd.n6031 gnd.n1322 163.367
R7793 gnd.n5856 gnd.n1322 163.367
R7794 gnd.n5856 gnd.n1434 163.367
R7795 gnd.n5859 gnd.n1434 163.367
R7796 gnd.n5859 gnd.n5854 163.367
R7797 gnd.n5875 gnd.n5854 163.367
R7798 gnd.n5876 gnd.n5875 163.367
R7799 gnd.n5877 gnd.n5876 163.367
R7800 gnd.n5877 gnd.n5851 163.367
R7801 gnd.n5883 gnd.n5851 163.367
R7802 gnd.n5883 gnd.n5852 163.367
R7803 gnd.n5852 gnd.n5843 163.367
R7804 gnd.n5894 gnd.n5843 163.367
R7805 gnd.n5895 gnd.n5894 163.367
R7806 gnd.n5895 gnd.n5840 163.367
R7807 gnd.n5901 gnd.n5840 163.367
R7808 gnd.n5901 gnd.n5841 163.367
R7809 gnd.n5841 gnd.n5831 163.367
R7810 gnd.n5911 gnd.n5831 163.367
R7811 gnd.n5912 gnd.n5911 163.367
R7812 gnd.n5912 gnd.n5829 163.367
R7813 gnd.n5917 gnd.n5829 163.367
R7814 gnd.n5917 gnd.n5820 163.367
R7815 gnd.n5927 gnd.n5820 163.367
R7816 gnd.n5928 gnd.n5927 163.367
R7817 gnd.n5928 gnd.n5817 163.367
R7818 gnd.n5933 gnd.n5817 163.367
R7819 gnd.n5933 gnd.n5818 163.367
R7820 gnd.n5818 gnd.n5809 163.367
R7821 gnd.n5943 gnd.n5809 163.367
R7822 gnd.n5943 gnd.n5806 163.367
R7823 gnd.n5958 gnd.n5806 163.367
R7824 gnd.n5958 gnd.n5807 163.367
R7825 gnd.n5807 gnd.n1082 163.367
R7826 gnd.n5953 gnd.n1082 163.367
R7827 gnd.n5953 gnd.n5801 163.367
R7828 gnd.n5950 gnd.n5801 163.367
R7829 gnd.n5950 gnd.n5949 163.367
R7830 gnd.n5949 gnd.n1060 163.367
R7831 gnd.n1060 gnd.n1053 163.367
R7832 gnd.n6365 gnd.n1053 163.367
R7833 gnd.n6365 gnd.n1050 163.367
R7834 gnd.n6371 gnd.n1050 163.367
R7835 gnd.n6371 gnd.n1051 163.367
R7836 gnd.n1051 gnd.n1043 163.367
R7837 gnd.n6384 gnd.n1043 163.367
R7838 gnd.n6385 gnd.n6384 163.367
R7839 gnd.n6385 gnd.n1041 163.367
R7840 gnd.n6393 gnd.n1041 163.367
R7841 gnd.n6393 gnd.n1016 163.367
R7842 gnd.n6389 gnd.n1016 163.367
R7843 gnd.n6389 gnd.n1010 163.367
R7844 gnd.n6433 gnd.n1010 163.367
R7845 gnd.n6434 gnd.n6433 163.367
R7846 gnd.n6434 gnd.n1007 163.367
R7847 gnd.n6439 gnd.n1007 163.367
R7848 gnd.n6439 gnd.n1008 163.367
R7849 gnd.n1008 gnd.n929 163.367
R7850 gnd.n6899 gnd.n929 163.367
R7851 gnd.n6899 gnd.n930 163.367
R7852 gnd.n6895 gnd.n930 163.367
R7853 gnd.n6895 gnd.n933 163.367
R7854 gnd.n940 gnd.n933 163.367
R7855 gnd.n6885 gnd.n940 163.367
R7856 gnd.n6885 gnd.n942 163.367
R7857 gnd.n6881 gnd.n942 163.367
R7858 gnd.n6881 gnd.n945 163.367
R7859 gnd.n956 gnd.n945 163.367
R7860 gnd.n956 gnd.n953 163.367
R7861 gnd.n6870 gnd.n953 163.367
R7862 gnd.n6870 gnd.n955 163.367
R7863 gnd.n6866 gnd.n955 163.367
R7864 gnd.n6866 gnd.n960 163.367
R7865 gnd.n969 gnd.n960 163.367
R7866 gnd.n970 gnd.n969 163.367
R7867 gnd.n6613 gnd.n970 163.367
R7868 gnd.n6613 gnd.n6609 163.367
R7869 gnd.n6619 gnd.n6609 163.367
R7870 gnd.n6619 gnd.n6610 163.367
R7871 gnd.n6610 gnd.n6598 163.367
R7872 gnd.n6631 gnd.n6598 163.367
R7873 gnd.n6632 gnd.n6631 163.367
R7874 gnd.n6632 gnd.n6595 163.367
R7875 gnd.n6637 gnd.n6595 163.367
R7876 gnd.n6637 gnd.n6596 163.367
R7877 gnd.n6596 gnd.n6589 163.367
R7878 gnd.n6646 gnd.n6589 163.367
R7879 gnd.n6646 gnd.n6587 163.367
R7880 gnd.n6651 gnd.n6587 163.367
R7881 gnd.n6651 gnd.n6583 163.367
R7882 gnd.n6661 gnd.n6583 163.367
R7883 gnd.n6662 gnd.n6661 163.367
R7884 gnd.n6662 gnd.n6508 163.367
R7885 gnd.n6667 gnd.n6508 163.367
R7886 gnd.n1426 gnd.n1425 163.367
R7887 gnd.n1425 gnd.n1349 163.367
R7888 gnd.n1421 gnd.n1419 163.367
R7889 gnd.n1417 gnd.n1351 163.367
R7890 gnd.n1413 gnd.n1411 163.367
R7891 gnd.n1409 gnd.n1353 163.367
R7892 gnd.n1405 gnd.n1403 163.367
R7893 gnd.n1401 gnd.n1355 163.367
R7894 gnd.n1397 gnd.n1395 163.367
R7895 gnd.n1393 gnd.n1357 163.367
R7896 gnd.n1389 gnd.n1387 163.367
R7897 gnd.n1385 gnd.n1359 163.367
R7898 gnd.n1381 gnd.n1379 163.367
R7899 gnd.n1377 gnd.n1361 163.367
R7900 gnd.n1373 gnd.n1371 163.367
R7901 gnd.n1368 gnd.n1367 163.367
R7902 gnd.n6099 gnd.n6097 163.367
R7903 gnd.n6095 gnd.n1304 163.367
R7904 gnd.n6090 gnd.n6088 163.367
R7905 gnd.n6086 gnd.n1308 163.367
R7906 gnd.n6082 gnd.n6080 163.367
R7907 gnd.n6078 gnd.n1310 163.367
R7908 gnd.n6074 gnd.n6072 163.367
R7909 gnd.n6070 gnd.n1312 163.367
R7910 gnd.n6066 gnd.n6064 163.367
R7911 gnd.n6062 gnd.n1314 163.367
R7912 gnd.n6058 gnd.n6056 163.367
R7913 gnd.n6054 gnd.n1316 163.367
R7914 gnd.n6050 gnd.n6048 163.367
R7915 gnd.n6046 gnd.n1318 163.367
R7916 gnd.n6042 gnd.n6040 163.367
R7917 gnd.n6038 gnd.n1320 163.367
R7918 gnd.n6029 gnd.n1325 163.367
R7919 gnd.n6029 gnd.n1327 163.367
R7920 gnd.n6025 gnd.n1327 163.367
R7921 gnd.n6025 gnd.n6024 163.367
R7922 gnd.n6024 gnd.n1433 163.367
R7923 gnd.n5864 gnd.n1433 163.367
R7924 gnd.n5873 gnd.n5864 163.367
R7925 gnd.n5873 gnd.n5865 163.367
R7926 gnd.n5869 gnd.n5865 163.367
R7927 gnd.n5869 gnd.n5849 163.367
R7928 gnd.n5885 gnd.n5849 163.367
R7929 gnd.n5886 gnd.n5885 163.367
R7930 gnd.n5886 gnd.n5846 163.367
R7931 gnd.n5892 gnd.n5846 163.367
R7932 gnd.n5892 gnd.n5847 163.367
R7933 gnd.n5847 gnd.n5837 163.367
R7934 gnd.n5903 gnd.n5837 163.367
R7935 gnd.n5904 gnd.n5903 163.367
R7936 gnd.n5904 gnd.n5834 163.367
R7937 gnd.n5909 gnd.n5834 163.367
R7938 gnd.n5909 gnd.n5835 163.367
R7939 gnd.n5835 gnd.n5826 163.367
R7940 gnd.n5919 gnd.n5826 163.367
R7941 gnd.n5919 gnd.n5823 163.367
R7942 gnd.n5925 gnd.n5823 163.367
R7943 gnd.n5925 gnd.n5824 163.367
R7944 gnd.n5824 gnd.n5814 163.367
R7945 gnd.n5935 gnd.n5814 163.367
R7946 gnd.n5936 gnd.n5935 163.367
R7947 gnd.n5936 gnd.n5812 163.367
R7948 gnd.n5941 gnd.n5812 163.367
R7949 gnd.n5941 gnd.n5805 163.367
R7950 gnd.n5961 gnd.n5805 163.367
R7951 gnd.n5962 gnd.n5961 163.367
R7952 gnd.n5962 gnd.n1080 163.367
R7953 gnd.n5802 gnd.n1080 163.367
R7954 gnd.n5968 gnd.n5802 163.367
R7955 gnd.n5968 gnd.n5803 163.367
R7956 gnd.n5803 gnd.n1058 163.367
R7957 gnd.n6358 gnd.n1058 163.367
R7958 gnd.n6358 gnd.n1056 163.367
R7959 gnd.n6363 gnd.n1056 163.367
R7960 gnd.n6363 gnd.n1048 163.367
R7961 gnd.n6373 gnd.n1048 163.367
R7962 gnd.n6374 gnd.n6373 163.367
R7963 gnd.n6374 gnd.n1045 163.367
R7964 gnd.n6382 gnd.n1045 163.367
R7965 gnd.n6382 gnd.n1046 163.367
R7966 gnd.n6378 gnd.n1046 163.367
R7967 gnd.n6378 gnd.n1015 163.367
R7968 gnd.n6425 gnd.n1015 163.367
R7969 gnd.n6426 gnd.n6425 163.367
R7970 gnd.n6426 gnd.n1012 163.367
R7971 gnd.n6431 gnd.n1012 163.367
R7972 gnd.n6431 gnd.n1013 163.367
R7973 gnd.n1013 gnd.n1006 163.367
R7974 gnd.n6442 gnd.n1006 163.367
R7975 gnd.n6442 gnd.n1004 163.367
R7976 gnd.n6447 gnd.n1004 163.367
R7977 gnd.n6447 gnd.n925 163.367
R7978 gnd.n935 gnd.n925 163.367
R7979 gnd.n6893 gnd.n935 163.367
R7980 gnd.n6893 gnd.n936 163.367
R7981 gnd.n6889 gnd.n936 163.367
R7982 gnd.n6889 gnd.n939 163.367
R7983 gnd.n947 gnd.n939 163.367
R7984 gnd.n6879 gnd.n947 163.367
R7985 gnd.n6879 gnd.n949 163.367
R7986 gnd.n6875 gnd.n949 163.367
R7987 gnd.n6875 gnd.n6874 163.367
R7988 gnd.n6874 gnd.n952 163.367
R7989 gnd.n963 gnd.n952 163.367
R7990 gnd.n6864 gnd.n963 163.367
R7991 gnd.n6864 gnd.n964 163.367
R7992 gnd.n6860 gnd.n964 163.367
R7993 gnd.n6860 gnd.n968 163.367
R7994 gnd.n6604 gnd.n968 163.367
R7995 gnd.n6607 gnd.n6604 163.367
R7996 gnd.n6622 gnd.n6607 163.367
R7997 gnd.n6623 gnd.n6622 163.367
R7998 gnd.n6623 gnd.n6601 163.367
R7999 gnd.n6629 gnd.n6601 163.367
R8000 gnd.n6629 gnd.n6602 163.367
R8001 gnd.n6602 gnd.n6593 163.367
R8002 gnd.n6639 gnd.n6593 163.367
R8003 gnd.n6640 gnd.n6639 163.367
R8004 gnd.n6640 gnd.n6591 163.367
R8005 gnd.n6644 gnd.n6591 163.367
R8006 gnd.n6644 gnd.n6586 163.367
R8007 gnd.n6655 gnd.n6586 163.367
R8008 gnd.n6655 gnd.n6584 163.367
R8009 gnd.n6659 gnd.n6584 163.367
R8010 gnd.n6659 gnd.n6509 163.367
R8011 gnd.n6790 gnd.n6509 163.367
R8012 gnd.n6790 gnd.n6510 163.367
R8013 gnd.n6530 gnd.n6529 156.462
R8014 gnd.n5121 gnd.n5089 153.042
R8015 gnd.n5185 gnd.n5184 152.079
R8016 gnd.n5153 gnd.n5152 152.079
R8017 gnd.n5121 gnd.n5120 152.079
R8018 gnd.n1340 gnd.n1339 152
R8019 gnd.n1341 gnd.n1330 152
R8020 gnd.n1343 gnd.n1342 152
R8021 gnd.n1345 gnd.n1328 152
R8022 gnd.n1347 gnd.n1346 152
R8023 gnd.n6528 gnd.n6512 152
R8024 gnd.n6520 gnd.n6513 152
R8025 gnd.n6519 gnd.n6518 152
R8026 gnd.n6517 gnd.n6514 152
R8027 gnd.n6515 gnd.t102 150.546
R8028 gnd.t78 gnd.n5163 147.661
R8029 gnd.t60 gnd.n5131 147.661
R8030 gnd.t80 gnd.n5099 147.661
R8031 gnd.t5 gnd.n5068 147.661
R8032 gnd.t410 gnd.n5036 147.661
R8033 gnd.t408 gnd.n5004 147.661
R8034 gnd.t45 gnd.n4972 147.661
R8035 gnd.t412 gnd.n4941 147.661
R8036 gnd.n6727 gnd.n6726 143.351
R8037 gnd.n1366 gnd.n1303 143.351
R8038 gnd.n6098 gnd.n1303 143.351
R8039 gnd.n7222 gnd.n639 138.177
R8040 gnd.n6101 gnd.n6100 138.177
R8041 gnd.n1337 gnd.t163 130.484
R8042 gnd.n1346 gnd.t188 126.766
R8043 gnd.n1344 gnd.t109 126.766
R8044 gnd.n1330 gnd.t173 126.766
R8045 gnd.n1338 gnd.t141 126.766
R8046 gnd.n6516 gnd.t87 126.766
R8047 gnd.n6518 gnd.t201 126.766
R8048 gnd.n6527 gnd.t150 126.766
R8049 gnd.n6529 gnd.t127 126.766
R8050 gnd.n5180 gnd.n5179 104.615
R8051 gnd.n5179 gnd.n5157 104.615
R8052 gnd.n5172 gnd.n5157 104.615
R8053 gnd.n5172 gnd.n5171 104.615
R8054 gnd.n5171 gnd.n5161 104.615
R8055 gnd.n5164 gnd.n5161 104.615
R8056 gnd.n5148 gnd.n5147 104.615
R8057 gnd.n5147 gnd.n5125 104.615
R8058 gnd.n5140 gnd.n5125 104.615
R8059 gnd.n5140 gnd.n5139 104.615
R8060 gnd.n5139 gnd.n5129 104.615
R8061 gnd.n5132 gnd.n5129 104.615
R8062 gnd.n5116 gnd.n5115 104.615
R8063 gnd.n5115 gnd.n5093 104.615
R8064 gnd.n5108 gnd.n5093 104.615
R8065 gnd.n5108 gnd.n5107 104.615
R8066 gnd.n5107 gnd.n5097 104.615
R8067 gnd.n5100 gnd.n5097 104.615
R8068 gnd.n5085 gnd.n5084 104.615
R8069 gnd.n5084 gnd.n5062 104.615
R8070 gnd.n5077 gnd.n5062 104.615
R8071 gnd.n5077 gnd.n5076 104.615
R8072 gnd.n5076 gnd.n5066 104.615
R8073 gnd.n5069 gnd.n5066 104.615
R8074 gnd.n5053 gnd.n5052 104.615
R8075 gnd.n5052 gnd.n5030 104.615
R8076 gnd.n5045 gnd.n5030 104.615
R8077 gnd.n5045 gnd.n5044 104.615
R8078 gnd.n5044 gnd.n5034 104.615
R8079 gnd.n5037 gnd.n5034 104.615
R8080 gnd.n5021 gnd.n5020 104.615
R8081 gnd.n5020 gnd.n4998 104.615
R8082 gnd.n5013 gnd.n4998 104.615
R8083 gnd.n5013 gnd.n5012 104.615
R8084 gnd.n5012 gnd.n5002 104.615
R8085 gnd.n5005 gnd.n5002 104.615
R8086 gnd.n4989 gnd.n4988 104.615
R8087 gnd.n4988 gnd.n4966 104.615
R8088 gnd.n4981 gnd.n4966 104.615
R8089 gnd.n4981 gnd.n4980 104.615
R8090 gnd.n4980 gnd.n4970 104.615
R8091 gnd.n4973 gnd.n4970 104.615
R8092 gnd.n4958 gnd.n4957 104.615
R8093 gnd.n4957 gnd.n4935 104.615
R8094 gnd.n4950 gnd.n4935 104.615
R8095 gnd.n4950 gnd.n4949 104.615
R8096 gnd.n4949 gnd.n4939 104.615
R8097 gnd.n4942 gnd.n4939 104.615
R8098 gnd.n4332 gnd.t119 100.632
R8099 gnd.n3858 gnd.t168 100.632
R8100 gnd.n7882 gnd.n7881 99.6594
R8101 gnd.n7877 gnd.n292 99.6594
R8102 gnd.n7873 gnd.n291 99.6594
R8103 gnd.n7869 gnd.n290 99.6594
R8104 gnd.n7865 gnd.n289 99.6594
R8105 gnd.n7861 gnd.n288 99.6594
R8106 gnd.n7857 gnd.n287 99.6594
R8107 gnd.n7853 gnd.n286 99.6594
R8108 gnd.n7846 gnd.n285 99.6594
R8109 gnd.n7842 gnd.n284 99.6594
R8110 gnd.n7838 gnd.n283 99.6594
R8111 gnd.n7834 gnd.n282 99.6594
R8112 gnd.n7830 gnd.n281 99.6594
R8113 gnd.n7826 gnd.n280 99.6594
R8114 gnd.n7822 gnd.n279 99.6594
R8115 gnd.n7818 gnd.n278 99.6594
R8116 gnd.n7814 gnd.n277 99.6594
R8117 gnd.n7810 gnd.n276 99.6594
R8118 gnd.n7802 gnd.n275 99.6594
R8119 gnd.n7800 gnd.n274 99.6594
R8120 gnd.n7796 gnd.n273 99.6594
R8121 gnd.n7792 gnd.n272 99.6594
R8122 gnd.n7788 gnd.n271 99.6594
R8123 gnd.n7784 gnd.n270 99.6594
R8124 gnd.n7780 gnd.n269 99.6594
R8125 gnd.n7776 gnd.n268 99.6594
R8126 gnd.n7772 gnd.n267 99.6594
R8127 gnd.n7768 gnd.n266 99.6594
R8128 gnd.n7759 gnd.n265 99.6594
R8129 gnd.n7273 gnd.n550 99.6594
R8130 gnd.n7268 gnd.n572 99.6594
R8131 gnd.n7265 gnd.n573 99.6594
R8132 gnd.n7261 gnd.n574 99.6594
R8133 gnd.n7257 gnd.n575 99.6594
R8134 gnd.n7253 gnd.n576 99.6594
R8135 gnd.n7249 gnd.n577 99.6594
R8136 gnd.n7245 gnd.n578 99.6594
R8137 gnd.n7241 gnd.n579 99.6594
R8138 gnd.n7236 gnd.n580 99.6594
R8139 gnd.n7232 gnd.n581 99.6594
R8140 gnd.n7228 gnd.n582 99.6594
R8141 gnd.n7224 gnd.n583 99.6594
R8142 gnd.n7219 gnd.n585 99.6594
R8143 gnd.n7215 gnd.n586 99.6594
R8144 gnd.n7211 gnd.n587 99.6594
R8145 gnd.n7207 gnd.n588 99.6594
R8146 gnd.n7203 gnd.n589 99.6594
R8147 gnd.n7199 gnd.n590 99.6594
R8148 gnd.n7195 gnd.n591 99.6594
R8149 gnd.n7191 gnd.n592 99.6594
R8150 gnd.n7187 gnd.n593 99.6594
R8151 gnd.n7183 gnd.n594 99.6594
R8152 gnd.n7179 gnd.n595 99.6594
R8153 gnd.n7175 gnd.n596 99.6594
R8154 gnd.n7171 gnd.n597 99.6594
R8155 gnd.n7167 gnd.n598 99.6594
R8156 gnd.n7163 gnd.n599 99.6594
R8157 gnd.n6144 gnd.n6143 99.6594
R8158 gnd.n6141 gnd.n6140 99.6594
R8159 gnd.n6136 gnd.n1262 99.6594
R8160 gnd.n6134 gnd.n6133 99.6594
R8161 gnd.n6129 gnd.n1269 99.6594
R8162 gnd.n6127 gnd.n6126 99.6594
R8163 gnd.n6122 gnd.n1276 99.6594
R8164 gnd.n6120 gnd.n6119 99.6594
R8165 gnd.n6114 gnd.n1285 99.6594
R8166 gnd.n6112 gnd.n6111 99.6594
R8167 gnd.n6107 gnd.n1292 99.6594
R8168 gnd.n6105 gnd.n6104 99.6594
R8169 gnd.n1515 gnd.n1514 99.6594
R8170 gnd.n1519 gnd.n1517 99.6594
R8171 gnd.n1525 gnd.n1509 99.6594
R8172 gnd.n1529 gnd.n1527 99.6594
R8173 gnd.n1535 gnd.n1505 99.6594
R8174 gnd.n1539 gnd.n1537 99.6594
R8175 gnd.n1545 gnd.n1499 99.6594
R8176 gnd.n1549 gnd.n1547 99.6594
R8177 gnd.n1555 gnd.n1495 99.6594
R8178 gnd.n1559 gnd.n1557 99.6594
R8179 gnd.n1565 gnd.n1491 99.6594
R8180 gnd.n1569 gnd.n1567 99.6594
R8181 gnd.n1575 gnd.n1487 99.6594
R8182 gnd.n1579 gnd.n1577 99.6594
R8183 gnd.n1585 gnd.n1483 99.6594
R8184 gnd.n1588 gnd.n1587 99.6594
R8185 gnd.n3832 gnd.n3831 99.6594
R8186 gnd.n3826 gnd.n3164 99.6594
R8187 gnd.n3823 gnd.n3165 99.6594
R8188 gnd.n3819 gnd.n3166 99.6594
R8189 gnd.n3815 gnd.n3167 99.6594
R8190 gnd.n3811 gnd.n3168 99.6594
R8191 gnd.n3807 gnd.n3169 99.6594
R8192 gnd.n3803 gnd.n3170 99.6594
R8193 gnd.n3799 gnd.n3171 99.6594
R8194 gnd.n3794 gnd.n3172 99.6594
R8195 gnd.n3790 gnd.n3173 99.6594
R8196 gnd.n3786 gnd.n3174 99.6594
R8197 gnd.n3782 gnd.n3175 99.6594
R8198 gnd.n3778 gnd.n3176 99.6594
R8199 gnd.n3774 gnd.n3177 99.6594
R8200 gnd.n3770 gnd.n3178 99.6594
R8201 gnd.n3766 gnd.n3179 99.6594
R8202 gnd.n3762 gnd.n3180 99.6594
R8203 gnd.n3758 gnd.n3181 99.6594
R8204 gnd.n3754 gnd.n3182 99.6594
R8205 gnd.n3750 gnd.n3183 99.6594
R8206 gnd.n3746 gnd.n3184 99.6594
R8207 gnd.n3742 gnd.n3185 99.6594
R8208 gnd.n3738 gnd.n3186 99.6594
R8209 gnd.n3734 gnd.n3187 99.6594
R8210 gnd.n3730 gnd.n3188 99.6594
R8211 gnd.n3726 gnd.n3189 99.6594
R8212 gnd.n3722 gnd.n3190 99.6594
R8213 gnd.n3718 gnd.n3191 99.6594
R8214 gnd.n5303 gnd.n3841 99.6594
R8215 gnd.n5301 gnd.n3840 99.6594
R8216 gnd.n5297 gnd.n3839 99.6594
R8217 gnd.n5293 gnd.n3838 99.6594
R8218 gnd.n5289 gnd.n3837 99.6594
R8219 gnd.n5285 gnd.n3836 99.6594
R8220 gnd.n5281 gnd.n3835 99.6594
R8221 gnd.n5213 gnd.n3834 99.6594
R8222 gnd.n4544 gnd.n4275 99.6594
R8223 gnd.n4301 gnd.n4282 99.6594
R8224 gnd.n4303 gnd.n4283 99.6594
R8225 gnd.n4311 gnd.n4284 99.6594
R8226 gnd.n4313 gnd.n4285 99.6594
R8227 gnd.n4321 gnd.n4286 99.6594
R8228 gnd.n4323 gnd.n4287 99.6594
R8229 gnd.n4331 gnd.n4288 99.6594
R8230 gnd.n7683 gnd.n256 99.6594
R8231 gnd.n7687 gnd.n257 99.6594
R8232 gnd.n7693 gnd.n258 99.6594
R8233 gnd.n7697 gnd.n259 99.6594
R8234 gnd.n7703 gnd.n260 99.6594
R8235 gnd.n7707 gnd.n261 99.6594
R8236 gnd.n7713 gnd.n262 99.6594
R8237 gnd.n7717 gnd.n263 99.6594
R8238 gnd.n7723 gnd.n264 99.6594
R8239 gnd.n600 gnd.n555 99.6594
R8240 gnd.n688 gnd.n601 99.6594
R8241 gnd.n696 gnd.n602 99.6594
R8242 gnd.n698 gnd.n603 99.6594
R8243 gnd.n706 gnd.n604 99.6594
R8244 gnd.n714 gnd.n605 99.6594
R8245 gnd.n716 gnd.n606 99.6594
R8246 gnd.n724 gnd.n607 99.6594
R8247 gnd.n734 gnd.n608 99.6594
R8248 gnd.n5271 gnd.n3151 99.6594
R8249 gnd.n5267 gnd.n3152 99.6594
R8250 gnd.n5263 gnd.n3153 99.6594
R8251 gnd.n5259 gnd.n3154 99.6594
R8252 gnd.n5255 gnd.n3155 99.6594
R8253 gnd.n5251 gnd.n3156 99.6594
R8254 gnd.n5247 gnd.n3157 99.6594
R8255 gnd.n5243 gnd.n3158 99.6594
R8256 gnd.n5239 gnd.n3159 99.6594
R8257 gnd.n5235 gnd.n3160 99.6594
R8258 gnd.n5231 gnd.n3161 99.6594
R8259 gnd.n5227 gnd.n3162 99.6594
R8260 gnd.n5223 gnd.n3163 99.6594
R8261 gnd.n4459 gnd.n4458 99.6594
R8262 gnd.n4453 gnd.n4370 99.6594
R8263 gnd.n4450 gnd.n4371 99.6594
R8264 gnd.n4446 gnd.n4372 99.6594
R8265 gnd.n4442 gnd.n4373 99.6594
R8266 gnd.n4438 gnd.n4374 99.6594
R8267 gnd.n4434 gnd.n4375 99.6594
R8268 gnd.n4430 gnd.n4376 99.6594
R8269 gnd.n4426 gnd.n4377 99.6594
R8270 gnd.n4422 gnd.n4378 99.6594
R8271 gnd.n4418 gnd.n4379 99.6594
R8272 gnd.n4414 gnd.n4380 99.6594
R8273 gnd.n4461 gnd.n4369 99.6594
R8274 gnd.n5618 gnd.n5617 99.6594
R8275 gnd.n5629 gnd.n5628 99.6594
R8276 gnd.n5638 gnd.n5637 99.6594
R8277 gnd.n5641 gnd.n5640 99.6594
R8278 gnd.n5652 gnd.n5651 99.6594
R8279 gnd.n5661 gnd.n5660 99.6594
R8280 gnd.n5664 gnd.n5663 99.6594
R8281 gnd.n5680 gnd.n5678 99.6594
R8282 gnd.n6154 gnd.n1240 99.6594
R8283 gnd.n3430 gnd.n3192 99.6594
R8284 gnd.n3434 gnd.n3193 99.6594
R8285 gnd.n3440 gnd.n3194 99.6594
R8286 gnd.n3444 gnd.n3195 99.6594
R8287 gnd.n3450 gnd.n3196 99.6594
R8288 gnd.n3454 gnd.n3197 99.6594
R8289 gnd.n3460 gnd.n3198 99.6594
R8290 gnd.n3464 gnd.n3199 99.6594
R8291 gnd.n3421 gnd.n3200 99.6594
R8292 gnd.n3433 gnd.n3192 99.6594
R8293 gnd.n3439 gnd.n3193 99.6594
R8294 gnd.n3443 gnd.n3194 99.6594
R8295 gnd.n3449 gnd.n3195 99.6594
R8296 gnd.n3453 gnd.n3196 99.6594
R8297 gnd.n3459 gnd.n3197 99.6594
R8298 gnd.n3463 gnd.n3198 99.6594
R8299 gnd.n3420 gnd.n3199 99.6594
R8300 gnd.n3416 gnd.n3200 99.6594
R8301 gnd.n5679 gnd.n1240 99.6594
R8302 gnd.n5678 gnd.n5677 99.6594
R8303 gnd.n5663 gnd.n5662 99.6594
R8304 gnd.n5660 gnd.n5653 99.6594
R8305 gnd.n5651 gnd.n5650 99.6594
R8306 gnd.n5640 gnd.n5639 99.6594
R8307 gnd.n5637 gnd.n5630 99.6594
R8308 gnd.n5628 gnd.n5627 99.6594
R8309 gnd.n5617 gnd.n5616 99.6594
R8310 gnd.n4459 gnd.n4382 99.6594
R8311 gnd.n4451 gnd.n4370 99.6594
R8312 gnd.n4447 gnd.n4371 99.6594
R8313 gnd.n4443 gnd.n4372 99.6594
R8314 gnd.n4439 gnd.n4373 99.6594
R8315 gnd.n4435 gnd.n4374 99.6594
R8316 gnd.n4431 gnd.n4375 99.6594
R8317 gnd.n4427 gnd.n4376 99.6594
R8318 gnd.n4423 gnd.n4377 99.6594
R8319 gnd.n4419 gnd.n4378 99.6594
R8320 gnd.n4415 gnd.n4379 99.6594
R8321 gnd.n4411 gnd.n4380 99.6594
R8322 gnd.n4462 gnd.n4461 99.6594
R8323 gnd.n5226 gnd.n3163 99.6594
R8324 gnd.n5230 gnd.n3162 99.6594
R8325 gnd.n5234 gnd.n3161 99.6594
R8326 gnd.n5238 gnd.n3160 99.6594
R8327 gnd.n5242 gnd.n3159 99.6594
R8328 gnd.n5246 gnd.n3158 99.6594
R8329 gnd.n5250 gnd.n3157 99.6594
R8330 gnd.n5254 gnd.n3156 99.6594
R8331 gnd.n5258 gnd.n3155 99.6594
R8332 gnd.n5262 gnd.n3154 99.6594
R8333 gnd.n5266 gnd.n3153 99.6594
R8334 gnd.n5270 gnd.n3152 99.6594
R8335 gnd.n3862 gnd.n3151 99.6594
R8336 gnd.n687 gnd.n600 99.6594
R8337 gnd.n695 gnd.n601 99.6594
R8338 gnd.n697 gnd.n602 99.6594
R8339 gnd.n705 gnd.n603 99.6594
R8340 gnd.n713 gnd.n604 99.6594
R8341 gnd.n715 gnd.n605 99.6594
R8342 gnd.n723 gnd.n606 99.6594
R8343 gnd.n733 gnd.n607 99.6594
R8344 gnd.n7107 gnd.n608 99.6594
R8345 gnd.n7716 gnd.n264 99.6594
R8346 gnd.n7714 gnd.n263 99.6594
R8347 gnd.n7706 gnd.n262 99.6594
R8348 gnd.n7704 gnd.n261 99.6594
R8349 gnd.n7696 gnd.n260 99.6594
R8350 gnd.n7694 gnd.n259 99.6594
R8351 gnd.n7686 gnd.n258 99.6594
R8352 gnd.n7684 gnd.n257 99.6594
R8353 gnd.n7678 gnd.n256 99.6594
R8354 gnd.n4545 gnd.n4544 99.6594
R8355 gnd.n4304 gnd.n4282 99.6594
R8356 gnd.n4310 gnd.n4283 99.6594
R8357 gnd.n4314 gnd.n4284 99.6594
R8358 gnd.n4320 gnd.n4285 99.6594
R8359 gnd.n4324 gnd.n4286 99.6594
R8360 gnd.n4330 gnd.n4287 99.6594
R8361 gnd.n4288 gnd.n4272 99.6594
R8362 gnd.n5280 gnd.n3834 99.6594
R8363 gnd.n5284 gnd.n3835 99.6594
R8364 gnd.n5288 gnd.n3836 99.6594
R8365 gnd.n5292 gnd.n3837 99.6594
R8366 gnd.n5296 gnd.n3838 99.6594
R8367 gnd.n5300 gnd.n3839 99.6594
R8368 gnd.n5304 gnd.n3840 99.6594
R8369 gnd.n3843 gnd.n3841 99.6594
R8370 gnd.n3832 gnd.n3204 99.6594
R8371 gnd.n3824 gnd.n3164 99.6594
R8372 gnd.n3820 gnd.n3165 99.6594
R8373 gnd.n3816 gnd.n3166 99.6594
R8374 gnd.n3812 gnd.n3167 99.6594
R8375 gnd.n3808 gnd.n3168 99.6594
R8376 gnd.n3804 gnd.n3169 99.6594
R8377 gnd.n3800 gnd.n3170 99.6594
R8378 gnd.n3795 gnd.n3171 99.6594
R8379 gnd.n3791 gnd.n3172 99.6594
R8380 gnd.n3787 gnd.n3173 99.6594
R8381 gnd.n3783 gnd.n3174 99.6594
R8382 gnd.n3779 gnd.n3175 99.6594
R8383 gnd.n3775 gnd.n3176 99.6594
R8384 gnd.n3771 gnd.n3177 99.6594
R8385 gnd.n3767 gnd.n3178 99.6594
R8386 gnd.n3763 gnd.n3179 99.6594
R8387 gnd.n3759 gnd.n3180 99.6594
R8388 gnd.n3755 gnd.n3181 99.6594
R8389 gnd.n3751 gnd.n3182 99.6594
R8390 gnd.n3747 gnd.n3183 99.6594
R8391 gnd.n3743 gnd.n3184 99.6594
R8392 gnd.n3739 gnd.n3185 99.6594
R8393 gnd.n3735 gnd.n3186 99.6594
R8394 gnd.n3731 gnd.n3187 99.6594
R8395 gnd.n3727 gnd.n3188 99.6594
R8396 gnd.n3723 gnd.n3189 99.6594
R8397 gnd.n3719 gnd.n3190 99.6594
R8398 gnd.n3274 gnd.n3191 99.6594
R8399 gnd.n1587 gnd.n1586 99.6594
R8400 gnd.n1578 gnd.n1483 99.6594
R8401 gnd.n1577 gnd.n1576 99.6594
R8402 gnd.n1568 gnd.n1487 99.6594
R8403 gnd.n1567 gnd.n1566 99.6594
R8404 gnd.n1558 gnd.n1491 99.6594
R8405 gnd.n1557 gnd.n1556 99.6594
R8406 gnd.n1548 gnd.n1495 99.6594
R8407 gnd.n1547 gnd.n1546 99.6594
R8408 gnd.n1538 gnd.n1499 99.6594
R8409 gnd.n1537 gnd.n1536 99.6594
R8410 gnd.n1528 gnd.n1505 99.6594
R8411 gnd.n1527 gnd.n1526 99.6594
R8412 gnd.n1518 gnd.n1509 99.6594
R8413 gnd.n1517 gnd.n1516 99.6594
R8414 gnd.n1298 gnd.n1293 99.6594
R8415 gnd.n6106 gnd.n6105 99.6594
R8416 gnd.n1292 gnd.n1286 99.6594
R8417 gnd.n6113 gnd.n6112 99.6594
R8418 gnd.n1285 gnd.n1277 99.6594
R8419 gnd.n6121 gnd.n6120 99.6594
R8420 gnd.n1276 gnd.n1270 99.6594
R8421 gnd.n6128 gnd.n6127 99.6594
R8422 gnd.n1269 gnd.n1263 99.6594
R8423 gnd.n6135 gnd.n6134 99.6594
R8424 gnd.n1262 gnd.n1255 99.6594
R8425 gnd.n6142 gnd.n6141 99.6594
R8426 gnd.n6145 gnd.n6144 99.6594
R8427 gnd.n7273 gnd.n7272 99.6594
R8428 gnd.n7266 gnd.n572 99.6594
R8429 gnd.n7262 gnd.n573 99.6594
R8430 gnd.n7258 gnd.n574 99.6594
R8431 gnd.n7254 gnd.n575 99.6594
R8432 gnd.n7250 gnd.n576 99.6594
R8433 gnd.n7246 gnd.n577 99.6594
R8434 gnd.n7242 gnd.n578 99.6594
R8435 gnd.n7237 gnd.n579 99.6594
R8436 gnd.n7233 gnd.n580 99.6594
R8437 gnd.n7229 gnd.n581 99.6594
R8438 gnd.n7225 gnd.n582 99.6594
R8439 gnd.n7220 gnd.n584 99.6594
R8440 gnd.n7216 gnd.n585 99.6594
R8441 gnd.n7212 gnd.n586 99.6594
R8442 gnd.n7208 gnd.n587 99.6594
R8443 gnd.n7204 gnd.n588 99.6594
R8444 gnd.n7200 gnd.n589 99.6594
R8445 gnd.n7196 gnd.n590 99.6594
R8446 gnd.n7192 gnd.n591 99.6594
R8447 gnd.n7188 gnd.n592 99.6594
R8448 gnd.n7184 gnd.n593 99.6594
R8449 gnd.n7180 gnd.n594 99.6594
R8450 gnd.n7176 gnd.n595 99.6594
R8451 gnd.n7172 gnd.n596 99.6594
R8452 gnd.n7168 gnd.n597 99.6594
R8453 gnd.n7164 gnd.n598 99.6594
R8454 gnd.n673 gnd.n599 99.6594
R8455 gnd.n7767 gnd.n265 99.6594
R8456 gnd.n7771 gnd.n266 99.6594
R8457 gnd.n7775 gnd.n267 99.6594
R8458 gnd.n7779 gnd.n268 99.6594
R8459 gnd.n7783 gnd.n269 99.6594
R8460 gnd.n7787 gnd.n270 99.6594
R8461 gnd.n7791 gnd.n271 99.6594
R8462 gnd.n7795 gnd.n272 99.6594
R8463 gnd.n7799 gnd.n273 99.6594
R8464 gnd.n7803 gnd.n274 99.6594
R8465 gnd.n7809 gnd.n275 99.6594
R8466 gnd.n7813 gnd.n276 99.6594
R8467 gnd.n7817 gnd.n277 99.6594
R8468 gnd.n7821 gnd.n278 99.6594
R8469 gnd.n7825 gnd.n279 99.6594
R8470 gnd.n7829 gnd.n280 99.6594
R8471 gnd.n7833 gnd.n281 99.6594
R8472 gnd.n7837 gnd.n282 99.6594
R8473 gnd.n7841 gnd.n283 99.6594
R8474 gnd.n7845 gnd.n284 99.6594
R8475 gnd.n7852 gnd.n285 99.6594
R8476 gnd.n7856 gnd.n286 99.6594
R8477 gnd.n7860 gnd.n287 99.6594
R8478 gnd.n7864 gnd.n288 99.6594
R8479 gnd.n7868 gnd.n289 99.6594
R8480 gnd.n7872 gnd.n290 99.6594
R8481 gnd.n7876 gnd.n291 99.6594
R8482 gnd.n293 gnd.n292 99.6594
R8483 gnd.n7882 gnd.n254 99.6594
R8484 gnd.n5740 gnd.n5739 99.6594
R8485 gnd.n1471 gnd.n1457 99.6594
R8486 gnd.n1475 gnd.n1458 99.6594
R8487 gnd.n1477 gnd.n1459 99.6594
R8488 gnd.n5611 gnd.n1460 99.6594
R8489 gnd.n5622 gnd.n1461 99.6594
R8490 gnd.n5624 gnd.n1462 99.6594
R8491 gnd.n5634 gnd.n1463 99.6594
R8492 gnd.n5645 gnd.n1464 99.6594
R8493 gnd.n5647 gnd.n1465 99.6594
R8494 gnd.n5657 gnd.n1466 99.6594
R8495 gnd.n5668 gnd.n1467 99.6594
R8496 gnd.n5674 gnd.n1469 99.6594
R8497 gnd.n1470 gnd.n1235 99.6594
R8498 gnd.n5739 gnd.n1455 99.6594
R8499 gnd.n1474 gnd.n1457 99.6594
R8500 gnd.n1476 gnd.n1458 99.6594
R8501 gnd.n5610 gnd.n1459 99.6594
R8502 gnd.n5621 gnd.n1460 99.6594
R8503 gnd.n5623 gnd.n1461 99.6594
R8504 gnd.n5633 gnd.n1462 99.6594
R8505 gnd.n5644 gnd.n1463 99.6594
R8506 gnd.n5646 gnd.n1464 99.6594
R8507 gnd.n5656 gnd.n1465 99.6594
R8508 gnd.n5667 gnd.n1466 99.6594
R8509 gnd.n5669 gnd.n1467 99.6594
R8510 gnd.n1469 gnd.n1468 99.6594
R8511 gnd.n1470 gnd.n1232 99.6594
R8512 gnd.n759 gnd.n753 99.6594
R8513 gnd.n761 gnd.n760 99.6594
R8514 gnd.n7081 gnd.n758 99.6594
R8515 gnd.n7079 gnd.n680 99.6594
R8516 gnd.n762 gnd.n682 99.6594
R8517 gnd.n764 gnd.n691 99.6594
R8518 gnd.n766 gnd.n765 99.6594
R8519 gnd.n767 gnd.n702 99.6594
R8520 gnd.n769 gnd.n709 99.6594
R8521 gnd.n771 gnd.n770 99.6594
R8522 gnd.n772 gnd.n720 99.6594
R8523 gnd.n774 gnd.n727 99.6594
R8524 gnd.n776 gnd.n775 99.6594
R8525 gnd.n777 gnd.n739 99.6594
R8526 gnd.n774 gnd.n773 99.6594
R8527 gnd.n772 gnd.n719 99.6594
R8528 gnd.n771 gnd.n710 99.6594
R8529 gnd.n769 gnd.n768 99.6594
R8530 gnd.n767 gnd.n701 99.6594
R8531 gnd.n766 gnd.n692 99.6594
R8532 gnd.n764 gnd.n763 99.6594
R8533 gnd.n762 gnd.n681 99.6594
R8534 gnd.n7080 gnd.n7079 99.6594
R8535 gnd.n758 gnd.n757 99.6594
R8536 gnd.n761 gnd.n754 99.6594
R8537 gnd.n759 gnd.n749 99.6594
R8538 gnd.n777 gnd.n744 99.6594
R8539 gnd.n776 gnd.n738 99.6594
R8540 gnd.n5670 gnd.t137 98.63
R8541 gnd.n7108 gnd.t97 98.63
R8542 gnd.n1237 gnd.t125 98.63
R8543 gnd.n629 gnd.t184 98.63
R8544 gnd.n652 gnd.t187 98.63
R8545 gnd.n675 gnd.t149 98.63
R8546 gnd.n350 gnd.t114 98.63
R8547 gnd.n330 gnd.t121 98.63
R8548 gnd.n7848 gnd.t145 98.63
R8549 gnd.n7667 gnd.t192 98.63
R8550 gnd.n3224 gnd.t140 98.63
R8551 gnd.n3246 gnd.t162 98.63
R8552 gnd.n3268 gnd.t181 98.63
R8553 gnd.n3417 gnd.t133 98.63
R8554 gnd.n1281 gnd.t154 98.63
R8555 gnd.n1480 gnd.t171 98.63
R8556 gnd.n1502 gnd.t199 98.63
R8557 gnd.n729 gnd.t100 98.63
R8558 gnd.n1305 gnd.t159 92.8196
R8559 gnd.n6559 gnd.t177 92.8196
R8560 gnd.n1362 gnd.t206 92.8118
R8561 gnd.n6553 gnd.t107 92.8118
R8562 gnd.n2275 gnd.n2267 84.8607
R8563 gnd.n2600 gnd.n2275 84.8607
R8564 gnd.n2600 gnd.n2599 84.8607
R8565 gnd.n2599 gnd.n2598 84.8607
R8566 gnd.n2598 gnd.n2276 84.8607
R8567 gnd.n2592 gnd.n2276 84.8607
R8568 gnd.n2592 gnd.n2591 84.8607
R8569 gnd.n2591 gnd.n2590 84.8607
R8570 gnd.n2590 gnd.n2284 84.8607
R8571 gnd.n2584 gnd.n2284 84.8607
R8572 gnd.n2584 gnd.n2583 84.8607
R8573 gnd.n2583 gnd.n2582 84.8607
R8574 gnd.n2582 gnd.n2292 84.8607
R8575 gnd.n2576 gnd.n2292 84.8607
R8576 gnd.n2576 gnd.n2575 84.8607
R8577 gnd.n2575 gnd.n2574 84.8607
R8578 gnd.n2574 gnd.n2300 84.8607
R8579 gnd.n2568 gnd.n2300 84.8607
R8580 gnd.n2568 gnd.n2567 84.8607
R8581 gnd.n2567 gnd.n2566 84.8607
R8582 gnd.n2566 gnd.n2308 84.8607
R8583 gnd.n2560 gnd.n2308 84.8607
R8584 gnd.n2560 gnd.n2559 84.8607
R8585 gnd.n2559 gnd.n2558 84.8607
R8586 gnd.n2558 gnd.n2316 84.8607
R8587 gnd.n2552 gnd.n2316 84.8607
R8588 gnd.n2552 gnd.n2551 84.8607
R8589 gnd.n2551 gnd.n2550 84.8607
R8590 gnd.n2550 gnd.n2324 84.8607
R8591 gnd.n2544 gnd.n2324 84.8607
R8592 gnd.n2544 gnd.n2543 84.8607
R8593 gnd.n2543 gnd.n2542 84.8607
R8594 gnd.n2542 gnd.n2332 84.8607
R8595 gnd.n2536 gnd.n2332 84.8607
R8596 gnd.n2536 gnd.n2535 84.8607
R8597 gnd.n2535 gnd.n2534 84.8607
R8598 gnd.n2534 gnd.n2340 84.8607
R8599 gnd.n2528 gnd.n2340 84.8607
R8600 gnd.n2528 gnd.n2527 84.8607
R8601 gnd.n2527 gnd.n2526 84.8607
R8602 gnd.n2526 gnd.n2348 84.8607
R8603 gnd.n2520 gnd.n2348 84.8607
R8604 gnd.n2520 gnd.n2519 84.8607
R8605 gnd.n2519 gnd.n2518 84.8607
R8606 gnd.n2518 gnd.n2356 84.8607
R8607 gnd.n2512 gnd.n2356 84.8607
R8608 gnd.n2512 gnd.n2511 84.8607
R8609 gnd.n2511 gnd.n2510 84.8607
R8610 gnd.n2510 gnd.n2364 84.8607
R8611 gnd.n2504 gnd.n2364 84.8607
R8612 gnd.n2504 gnd.n2503 84.8607
R8613 gnd.n2503 gnd.n2502 84.8607
R8614 gnd.n2502 gnd.n2372 84.8607
R8615 gnd.n2496 gnd.n2372 84.8607
R8616 gnd.n2496 gnd.n2495 84.8607
R8617 gnd.n2495 gnd.n2494 84.8607
R8618 gnd.n2494 gnd.n2380 84.8607
R8619 gnd.n2488 gnd.n2380 84.8607
R8620 gnd.n2488 gnd.n2487 84.8607
R8621 gnd.n2487 gnd.n2486 84.8607
R8622 gnd.n2486 gnd.n2388 84.8607
R8623 gnd.n2480 gnd.n2388 84.8607
R8624 gnd.n2480 gnd.n2479 84.8607
R8625 gnd.n2479 gnd.n2478 84.8607
R8626 gnd.n2478 gnd.n2396 84.8607
R8627 gnd.n2472 gnd.n2396 84.8607
R8628 gnd.n2472 gnd.n2471 84.8607
R8629 gnd.n2471 gnd.n2470 84.8607
R8630 gnd.n2470 gnd.n2404 84.8607
R8631 gnd.n2464 gnd.n2404 84.8607
R8632 gnd.n2464 gnd.n2463 84.8607
R8633 gnd.n2463 gnd.n2462 84.8607
R8634 gnd.n2462 gnd.n2412 84.8607
R8635 gnd.n2456 gnd.n2412 84.8607
R8636 gnd.n2456 gnd.n2455 84.8607
R8637 gnd.n2455 gnd.n2454 84.8607
R8638 gnd.n2454 gnd.n2420 84.8607
R8639 gnd.n2448 gnd.n2420 84.8607
R8640 gnd.n2448 gnd.n2447 84.8607
R8641 gnd.n2447 gnd.n2446 84.8607
R8642 gnd.n2446 gnd.n2428 84.8607
R8643 gnd.n2440 gnd.n2428 84.8607
R8644 gnd.n2440 gnd.n2439 84.8607
R8645 gnd.n1337 gnd.n1336 81.8399
R8646 gnd.n4333 gnd.t118 74.8376
R8647 gnd.n3859 gnd.t169 74.8376
R8648 gnd.n1306 gnd.t158 72.8438
R8649 gnd.n6560 gnd.t178 72.8438
R8650 gnd.n1338 gnd.n1331 72.8411
R8651 gnd.n1344 gnd.n1329 72.8411
R8652 gnd.n6527 gnd.n6526 72.8411
R8653 gnd.n5671 gnd.t136 72.836
R8654 gnd.n1363 gnd.t205 72.836
R8655 gnd.n6554 gnd.t108 72.836
R8656 gnd.n7109 gnd.t96 72.836
R8657 gnd.n1238 gnd.t126 72.836
R8658 gnd.n630 gnd.t183 72.836
R8659 gnd.n653 gnd.t186 72.836
R8660 gnd.n676 gnd.t148 72.836
R8661 gnd.n351 gnd.t115 72.836
R8662 gnd.n331 gnd.t122 72.836
R8663 gnd.n7849 gnd.t146 72.836
R8664 gnd.n7668 gnd.t193 72.836
R8665 gnd.n3225 gnd.t139 72.836
R8666 gnd.n3247 gnd.t161 72.836
R8667 gnd.n3269 gnd.t180 72.836
R8668 gnd.n3418 gnd.t132 72.836
R8669 gnd.n1282 gnd.t155 72.836
R8670 gnd.n1481 gnd.t172 72.836
R8671 gnd.n1503 gnd.t200 72.836
R8672 gnd.n730 gnd.t101 72.836
R8673 gnd.n6784 gnd.n6783 71.676
R8674 gnd.n6781 gnd.n6780 71.676
R8675 gnd.n6776 gnd.n6536 71.676
R8676 gnd.n6774 gnd.n6773 71.676
R8677 gnd.n6769 gnd.n6539 71.676
R8678 gnd.n6767 gnd.n6766 71.676
R8679 gnd.n6762 gnd.n6542 71.676
R8680 gnd.n6760 gnd.n6759 71.676
R8681 gnd.n6755 gnd.n6545 71.676
R8682 gnd.n6753 gnd.n6752 71.676
R8683 gnd.n6748 gnd.n6548 71.676
R8684 gnd.n6746 gnd.n6745 71.676
R8685 gnd.n6741 gnd.n6551 71.676
R8686 gnd.n6739 gnd.n6738 71.676
R8687 gnd.n6733 gnd.n6556 71.676
R8688 gnd.n6731 gnd.n6730 71.676
R8689 gnd.n6726 gnd.n6725 71.676
R8690 gnd.n6723 gnd.n6722 71.676
R8691 gnd.n6717 gnd.n6562 71.676
R8692 gnd.n6715 gnd.n6714 71.676
R8693 gnd.n6710 gnd.n6565 71.676
R8694 gnd.n6708 gnd.n6707 71.676
R8695 gnd.n6703 gnd.n6568 71.676
R8696 gnd.n6701 gnd.n6700 71.676
R8697 gnd.n6696 gnd.n6571 71.676
R8698 gnd.n6694 gnd.n6693 71.676
R8699 gnd.n6689 gnd.n6574 71.676
R8700 gnd.n6687 gnd.n6686 71.676
R8701 gnd.n6682 gnd.n6577 71.676
R8702 gnd.n6680 gnd.n6679 71.676
R8703 gnd.n6675 gnd.n6580 71.676
R8704 gnd.n6673 gnd.n6672 71.676
R8705 gnd.n6668 gnd.n6666 71.676
R8706 gnd.n1428 gnd.n1427 71.676
R8707 gnd.n1420 gnd.n1349 71.676
R8708 gnd.n1419 gnd.n1418 71.676
R8709 gnd.n1412 gnd.n1351 71.676
R8710 gnd.n1411 gnd.n1410 71.676
R8711 gnd.n1404 gnd.n1353 71.676
R8712 gnd.n1403 gnd.n1402 71.676
R8713 gnd.n1396 gnd.n1355 71.676
R8714 gnd.n1395 gnd.n1394 71.676
R8715 gnd.n1388 gnd.n1357 71.676
R8716 gnd.n1387 gnd.n1386 71.676
R8717 gnd.n1380 gnd.n1359 71.676
R8718 gnd.n1379 gnd.n1378 71.676
R8719 gnd.n1372 gnd.n1361 71.676
R8720 gnd.n1371 gnd.n1365 71.676
R8721 gnd.n1367 gnd.n1366 71.676
R8722 gnd.n6097 gnd.n6096 71.676
R8723 gnd.n6089 gnd.n1304 71.676
R8724 gnd.n6088 gnd.n6087 71.676
R8725 gnd.n6081 gnd.n1308 71.676
R8726 gnd.n6080 gnd.n6079 71.676
R8727 gnd.n6073 gnd.n1310 71.676
R8728 gnd.n6072 gnd.n6071 71.676
R8729 gnd.n6065 gnd.n1312 71.676
R8730 gnd.n6064 gnd.n6063 71.676
R8731 gnd.n6057 gnd.n1314 71.676
R8732 gnd.n6056 gnd.n6055 71.676
R8733 gnd.n6049 gnd.n1316 71.676
R8734 gnd.n6048 gnd.n6047 71.676
R8735 gnd.n6041 gnd.n1318 71.676
R8736 gnd.n6040 gnd.n6039 71.676
R8737 gnd.n6033 gnd.n1320 71.676
R8738 gnd.n1427 gnd.n1426 71.676
R8739 gnd.n1421 gnd.n1420 71.676
R8740 gnd.n1418 gnd.n1417 71.676
R8741 gnd.n1413 gnd.n1412 71.676
R8742 gnd.n1410 gnd.n1409 71.676
R8743 gnd.n1405 gnd.n1404 71.676
R8744 gnd.n1402 gnd.n1401 71.676
R8745 gnd.n1397 gnd.n1396 71.676
R8746 gnd.n1394 gnd.n1393 71.676
R8747 gnd.n1389 gnd.n1388 71.676
R8748 gnd.n1386 gnd.n1385 71.676
R8749 gnd.n1381 gnd.n1380 71.676
R8750 gnd.n1378 gnd.n1377 71.676
R8751 gnd.n1373 gnd.n1372 71.676
R8752 gnd.n1368 gnd.n1365 71.676
R8753 gnd.n6099 gnd.n6098 71.676
R8754 gnd.n6096 gnd.n6095 71.676
R8755 gnd.n6090 gnd.n6089 71.676
R8756 gnd.n6087 gnd.n6086 71.676
R8757 gnd.n6082 gnd.n6081 71.676
R8758 gnd.n6079 gnd.n6078 71.676
R8759 gnd.n6074 gnd.n6073 71.676
R8760 gnd.n6071 gnd.n6070 71.676
R8761 gnd.n6066 gnd.n6065 71.676
R8762 gnd.n6063 gnd.n6062 71.676
R8763 gnd.n6058 gnd.n6057 71.676
R8764 gnd.n6055 gnd.n6054 71.676
R8765 gnd.n6050 gnd.n6049 71.676
R8766 gnd.n6047 gnd.n6046 71.676
R8767 gnd.n6042 gnd.n6041 71.676
R8768 gnd.n6039 gnd.n6038 71.676
R8769 gnd.n6034 gnd.n6033 71.676
R8770 gnd.n6666 gnd.n6581 71.676
R8771 gnd.n6674 gnd.n6673 71.676
R8772 gnd.n6580 gnd.n6578 71.676
R8773 gnd.n6681 gnd.n6680 71.676
R8774 gnd.n6577 gnd.n6575 71.676
R8775 gnd.n6688 gnd.n6687 71.676
R8776 gnd.n6574 gnd.n6572 71.676
R8777 gnd.n6695 gnd.n6694 71.676
R8778 gnd.n6571 gnd.n6569 71.676
R8779 gnd.n6702 gnd.n6701 71.676
R8780 gnd.n6568 gnd.n6566 71.676
R8781 gnd.n6709 gnd.n6708 71.676
R8782 gnd.n6565 gnd.n6563 71.676
R8783 gnd.n6716 gnd.n6715 71.676
R8784 gnd.n6562 gnd.n6558 71.676
R8785 gnd.n6724 gnd.n6723 71.676
R8786 gnd.n6728 gnd.n6727 71.676
R8787 gnd.n6732 gnd.n6731 71.676
R8788 gnd.n6556 gnd.n6552 71.676
R8789 gnd.n6740 gnd.n6739 71.676
R8790 gnd.n6551 gnd.n6549 71.676
R8791 gnd.n6747 gnd.n6746 71.676
R8792 gnd.n6548 gnd.n6546 71.676
R8793 gnd.n6754 gnd.n6753 71.676
R8794 gnd.n6545 gnd.n6543 71.676
R8795 gnd.n6761 gnd.n6760 71.676
R8796 gnd.n6542 gnd.n6540 71.676
R8797 gnd.n6768 gnd.n6767 71.676
R8798 gnd.n6539 gnd.n6537 71.676
R8799 gnd.n6775 gnd.n6774 71.676
R8800 gnd.n6536 gnd.n6534 71.676
R8801 gnd.n6782 gnd.n6781 71.676
R8802 gnd.n6785 gnd.n6784 71.676
R8803 gnd.n10 gnd.t11 69.1507
R8804 gnd.n18 gnd.t21 68.4792
R8805 gnd.n17 gnd.t76 68.4792
R8806 gnd.n16 gnd.t62 68.4792
R8807 gnd.n15 gnd.t33 68.4792
R8808 gnd.n14 gnd.t56 68.4792
R8809 gnd.n13 gnd.t49 68.4792
R8810 gnd.n12 gnd.t24 68.4792
R8811 gnd.n11 gnd.t35 68.4792
R8812 gnd.n10 gnd.t7 68.4792
R8813 gnd.n4460 gnd.n4364 64.369
R8814 gnd.n6092 gnd.n1306 59.5399
R8815 gnd.n6719 gnd.n6560 59.5399
R8816 gnd.n1364 gnd.n1363 59.5399
R8817 gnd.n6735 gnd.n6554 59.5399
R8818 gnd.n1430 gnd.n1347 59.1804
R8819 gnd.n4111 gnd.t358 56.407
R8820 gnd.n4052 gnd.t384 56.407
R8821 gnd.n4071 gnd.t335 56.407
R8822 gnd.n4091 gnd.t228 56.407
R8823 gnd.n80 gnd.t328 56.407
R8824 gnd.n21 gnd.t245 56.407
R8825 gnd.n40 gnd.t314 56.407
R8826 gnd.n60 gnd.t371 56.407
R8827 gnd.n4128 gnd.t388 55.8337
R8828 gnd.n4069 gnd.t218 55.8337
R8829 gnd.n4088 gnd.t232 55.8337
R8830 gnd.n4108 gnd.t300 55.8337
R8831 gnd.n97 gnd.t331 55.8337
R8832 gnd.n38 gnd.t243 55.8337
R8833 gnd.n57 gnd.t383 55.8337
R8834 gnd.n77 gnd.t375 55.8337
R8835 gnd.n1335 gnd.n1334 54.358
R8836 gnd.n6524 gnd.n6523 54.358
R8837 gnd.n4111 gnd.n4110 53.0052
R8838 gnd.n4113 gnd.n4112 53.0052
R8839 gnd.n4115 gnd.n4114 53.0052
R8840 gnd.n4117 gnd.n4116 53.0052
R8841 gnd.n4119 gnd.n4118 53.0052
R8842 gnd.n4121 gnd.n4120 53.0052
R8843 gnd.n4123 gnd.n4122 53.0052
R8844 gnd.n4125 gnd.n4124 53.0052
R8845 gnd.n4127 gnd.n4126 53.0052
R8846 gnd.n4052 gnd.n4051 53.0052
R8847 gnd.n4054 gnd.n4053 53.0052
R8848 gnd.n4056 gnd.n4055 53.0052
R8849 gnd.n4058 gnd.n4057 53.0052
R8850 gnd.n4060 gnd.n4059 53.0052
R8851 gnd.n4062 gnd.n4061 53.0052
R8852 gnd.n4064 gnd.n4063 53.0052
R8853 gnd.n4066 gnd.n4065 53.0052
R8854 gnd.n4068 gnd.n4067 53.0052
R8855 gnd.n4071 gnd.n4070 53.0052
R8856 gnd.n4073 gnd.n4072 53.0052
R8857 gnd.n4075 gnd.n4074 53.0052
R8858 gnd.n4077 gnd.n4076 53.0052
R8859 gnd.n4079 gnd.n4078 53.0052
R8860 gnd.n4081 gnd.n4080 53.0052
R8861 gnd.n4083 gnd.n4082 53.0052
R8862 gnd.n4085 gnd.n4084 53.0052
R8863 gnd.n4087 gnd.n4086 53.0052
R8864 gnd.n4091 gnd.n4090 53.0052
R8865 gnd.n4093 gnd.n4092 53.0052
R8866 gnd.n4095 gnd.n4094 53.0052
R8867 gnd.n4097 gnd.n4096 53.0052
R8868 gnd.n4099 gnd.n4098 53.0052
R8869 gnd.n4101 gnd.n4100 53.0052
R8870 gnd.n4103 gnd.n4102 53.0052
R8871 gnd.n4105 gnd.n4104 53.0052
R8872 gnd.n4107 gnd.n4106 53.0052
R8873 gnd.n96 gnd.n95 53.0052
R8874 gnd.n94 gnd.n93 53.0052
R8875 gnd.n92 gnd.n91 53.0052
R8876 gnd.n90 gnd.n89 53.0052
R8877 gnd.n88 gnd.n87 53.0052
R8878 gnd.n86 gnd.n85 53.0052
R8879 gnd.n84 gnd.n83 53.0052
R8880 gnd.n82 gnd.n81 53.0052
R8881 gnd.n80 gnd.n79 53.0052
R8882 gnd.n37 gnd.n36 53.0052
R8883 gnd.n35 gnd.n34 53.0052
R8884 gnd.n33 gnd.n32 53.0052
R8885 gnd.n31 gnd.n30 53.0052
R8886 gnd.n29 gnd.n28 53.0052
R8887 gnd.n27 gnd.n26 53.0052
R8888 gnd.n25 gnd.n24 53.0052
R8889 gnd.n23 gnd.n22 53.0052
R8890 gnd.n21 gnd.n20 53.0052
R8891 gnd.n56 gnd.n55 53.0052
R8892 gnd.n54 gnd.n53 53.0052
R8893 gnd.n52 gnd.n51 53.0052
R8894 gnd.n50 gnd.n49 53.0052
R8895 gnd.n48 gnd.n47 53.0052
R8896 gnd.n46 gnd.n45 53.0052
R8897 gnd.n44 gnd.n43 53.0052
R8898 gnd.n42 gnd.n41 53.0052
R8899 gnd.n40 gnd.n39 53.0052
R8900 gnd.n76 gnd.n75 53.0052
R8901 gnd.n74 gnd.n73 53.0052
R8902 gnd.n72 gnd.n71 53.0052
R8903 gnd.n70 gnd.n69 53.0052
R8904 gnd.n68 gnd.n67 53.0052
R8905 gnd.n66 gnd.n65 53.0052
R8906 gnd.n64 gnd.n63 53.0052
R8907 gnd.n62 gnd.n61 53.0052
R8908 gnd.n60 gnd.n59 53.0052
R8909 gnd.n6515 gnd.n6514 52.4801
R8910 gnd.n5164 gnd.t78 52.3082
R8911 gnd.n5132 gnd.t60 52.3082
R8912 gnd.n5100 gnd.t80 52.3082
R8913 gnd.n5069 gnd.t5 52.3082
R8914 gnd.n5037 gnd.t410 52.3082
R8915 gnd.n5005 gnd.t408 52.3082
R8916 gnd.n4973 gnd.t45 52.3082
R8917 gnd.n4942 gnd.t412 52.3082
R8918 gnd.n3833 gnd.n3202 51.6227
R8919 gnd.n7883 gnd.n248 51.6227
R8920 gnd.n4994 gnd.n4962 51.4173
R8921 gnd.n2439 gnd.n201 50.9166
R8922 gnd.n5058 gnd.n5057 50.455
R8923 gnd.n5026 gnd.n5025 50.455
R8924 gnd.n4994 gnd.n4993 50.455
R8925 gnd.n4407 gnd.n4406 45.1884
R8926 gnd.n3885 gnd.n3884 45.1884
R8927 gnd.n6787 gnd.n6530 44.3322
R8928 gnd.n1338 gnd.n1337 44.3189
R8929 gnd.n5672 gnd.n5671 42.4732
R8930 gnd.n731 gnd.n730 42.4732
R8931 gnd.n7110 gnd.n7109 42.2793
R8932 gnd.n4408 gnd.n4407 42.2793
R8933 gnd.n3886 gnd.n3885 42.2793
R8934 gnd.n4334 gnd.n4333 42.2793
R8935 gnd.n5279 gnd.n3859 42.2793
R8936 gnd.n1239 gnd.n1238 42.2793
R8937 gnd.n7239 gnd.n630 42.2793
R8938 gnd.n7202 gnd.n653 42.2793
R8939 gnd.n7162 gnd.n676 42.2793
R8940 gnd.n7766 gnd.n351 42.2793
R8941 gnd.n7808 gnd.n331 42.2793
R8942 gnd.n7850 gnd.n7849 42.2793
R8943 gnd.n7669 gnd.n7668 42.2793
R8944 gnd.n3797 gnd.n3225 42.2793
R8945 gnd.n3757 gnd.n3247 42.2793
R8946 gnd.n3717 gnd.n3269 42.2793
R8947 gnd.n3470 gnd.n3418 42.2793
R8948 gnd.n6116 gnd.n1282 42.2793
R8949 gnd.n1482 gnd.n1481 42.2793
R8950 gnd.n1504 gnd.n1503 42.2793
R8951 gnd.n1336 gnd.n1335 41.6274
R8952 gnd.n6525 gnd.n6524 41.6274
R8953 gnd.n1345 gnd.n1344 40.8975
R8954 gnd.n6528 gnd.n6527 40.8975
R8955 gnd.n1344 gnd.n1343 35.055
R8956 gnd.n1339 gnd.n1338 35.055
R8957 gnd.n6517 gnd.n6516 35.055
R8958 gnd.n6527 gnd.n6513 35.055
R8959 gnd.n2948 gnd.n2947 31.9958
R8960 gnd.n2949 gnd.n2948 31.9958
R8961 gnd.n2949 gnd.n1928 31.9958
R8962 gnd.n2957 gnd.n1928 31.9958
R8963 gnd.n2958 gnd.n2957 31.9958
R8964 gnd.n2959 gnd.n2958 31.9958
R8965 gnd.n2959 gnd.n1922 31.9958
R8966 gnd.n2967 gnd.n1922 31.9958
R8967 gnd.n2968 gnd.n2967 31.9958
R8968 gnd.n2969 gnd.n2968 31.9958
R8969 gnd.n2969 gnd.n1916 31.9958
R8970 gnd.n2977 gnd.n1916 31.9958
R8971 gnd.n2978 gnd.n2977 31.9958
R8972 gnd.n2979 gnd.n2978 31.9958
R8973 gnd.n2979 gnd.n1910 31.9958
R8974 gnd.n2987 gnd.n1910 31.9958
R8975 gnd.n2988 gnd.n2987 31.9958
R8976 gnd.n2989 gnd.n2988 31.9958
R8977 gnd.n2989 gnd.n1904 31.9958
R8978 gnd.n2997 gnd.n1904 31.9958
R8979 gnd.n2998 gnd.n2997 31.9958
R8980 gnd.n2999 gnd.n2998 31.9958
R8981 gnd.n2999 gnd.n1898 31.9958
R8982 gnd.n3007 gnd.n1898 31.9958
R8983 gnd.n3008 gnd.n3007 31.9958
R8984 gnd.n3009 gnd.n3008 31.9958
R8985 gnd.n3009 gnd.n1892 31.9958
R8986 gnd.n3017 gnd.n1892 31.9958
R8987 gnd.n3018 gnd.n3017 31.9958
R8988 gnd.n3019 gnd.n3018 31.9958
R8989 gnd.n3019 gnd.n1886 31.9958
R8990 gnd.n3027 gnd.n1886 31.9958
R8991 gnd.n3028 gnd.n3027 31.9958
R8992 gnd.n3029 gnd.n3028 31.9958
R8993 gnd.n3029 gnd.n1880 31.9958
R8994 gnd.n3037 gnd.n1880 31.9958
R8995 gnd.n3038 gnd.n3037 31.9958
R8996 gnd.n3039 gnd.n3038 31.9958
R8997 gnd.n3039 gnd.n1874 31.9958
R8998 gnd.n3047 gnd.n1874 31.9958
R8999 gnd.n3048 gnd.n3047 31.9958
R9000 gnd.n3049 gnd.n3048 31.9958
R9001 gnd.n3049 gnd.n1868 31.9958
R9002 gnd.n3057 gnd.n1868 31.9958
R9003 gnd.n3058 gnd.n3057 31.9958
R9004 gnd.n3059 gnd.n3058 31.9958
R9005 gnd.n3059 gnd.n1862 31.9958
R9006 gnd.n3067 gnd.n1862 31.9958
R9007 gnd.n3068 gnd.n3067 31.9958
R9008 gnd.n3069 gnd.n3068 31.9958
R9009 gnd.n3069 gnd.n1856 31.9958
R9010 gnd.n3077 gnd.n1856 31.9958
R9011 gnd.n3078 gnd.n3077 31.9958
R9012 gnd.n3079 gnd.n3078 31.9958
R9013 gnd.n3079 gnd.n1850 31.9958
R9014 gnd.n3087 gnd.n1850 31.9958
R9015 gnd.n3088 gnd.n3087 31.9958
R9016 gnd.n3089 gnd.n3088 31.9958
R9017 gnd.n3089 gnd.n1844 31.9958
R9018 gnd.n3097 gnd.n1844 31.9958
R9019 gnd.n3098 gnd.n3097 31.9958
R9020 gnd.n3099 gnd.n3098 31.9958
R9021 gnd.n3099 gnd.n1838 31.9958
R9022 gnd.n3107 gnd.n1838 31.9958
R9023 gnd.n3108 gnd.n3107 31.9958
R9024 gnd.n3109 gnd.n3108 31.9958
R9025 gnd.n3109 gnd.n1832 31.9958
R9026 gnd.n3117 gnd.n1832 31.9958
R9027 gnd.n3118 gnd.n3117 31.9958
R9028 gnd.n3119 gnd.n3118 31.9958
R9029 gnd.n3119 gnd.n1826 31.9958
R9030 gnd.n3127 gnd.n1826 31.9958
R9031 gnd.n3128 gnd.n3127 31.9958
R9032 gnd.n3129 gnd.n3128 31.9958
R9033 gnd.n3129 gnd.n1820 31.9958
R9034 gnd.n3137 gnd.n1820 31.9958
R9035 gnd.n3138 gnd.n3137 31.9958
R9036 gnd.n3139 gnd.n3138 31.9958
R9037 gnd.n3139 gnd.n1814 31.9958
R9038 gnd.n3147 gnd.n1814 31.9958
R9039 gnd.n3148 gnd.n3147 31.9958
R9040 gnd.n5315 gnd.n3148 31.9958
R9041 gnd.n5315 gnd.n5314 31.9958
R9042 gnd.n4470 gnd.n4364 31.8661
R9043 gnd.n4470 gnd.n4469 31.8661
R9044 gnd.n4478 gnd.n4353 31.8661
R9045 gnd.n4486 gnd.n4353 31.8661
R9046 gnd.n4486 gnd.n4347 31.8661
R9047 gnd.n4494 gnd.n4347 31.8661
R9048 gnd.n4494 gnd.n4340 31.8661
R9049 gnd.n4532 gnd.n4340 31.8661
R9050 gnd.n4542 gnd.n4273 31.8661
R9051 gnd.n3709 gnd.n3202 31.8661
R9052 gnd.n3703 gnd.n3286 31.8661
R9053 gnd.n3703 gnd.n3289 31.8661
R9054 gnd.n3697 gnd.n3289 31.8661
R9055 gnd.n3697 gnd.n3301 31.8661
R9056 gnd.n3691 gnd.n3311 31.8661
R9057 gnd.n3685 gnd.n3311 31.8661
R9058 gnd.n3679 gnd.n3327 31.8661
R9059 gnd.n3679 gnd.n3330 31.8661
R9060 gnd.n3673 gnd.n3339 31.8661
R9061 gnd.n3667 gnd.n3349 31.8661
R9062 gnd.n3661 gnd.n3349 31.8661
R9063 gnd.n3655 gnd.n3365 31.8661
R9064 gnd.n3655 gnd.n3368 31.8661
R9065 gnd.n3649 gnd.n3377 31.8661
R9066 gnd.n3643 gnd.n3387 31.8661
R9067 gnd.n3637 gnd.n3387 31.8661
R9068 gnd.n3630 gnd.n3629 31.8661
R9069 gnd.n3629 gnd.n3548 31.8661
R9070 gnd.n5347 gnd.n1784 31.8661
R9071 gnd.n5341 gnd.n1795 31.8661
R9072 gnd.n5333 gnd.n1795 31.8661
R9073 gnd.n5327 gnd.n1805 31.8661
R9074 gnd.n5357 gnd.n1766 31.8661
R9075 gnd.n5523 gnd.n1245 31.8661
R9076 gnd.n5518 gnd.n5517 31.8661
R9077 gnd.n5518 gnd.n1456 31.8661
R9078 gnd.n6164 gnd.n1229 31.8661
R9079 gnd.n6164 gnd.n1231 31.8661
R9080 gnd.n6172 gnd.n1216 31.8661
R9081 gnd.n6180 gnd.n1216 31.8661
R9082 gnd.n6180 gnd.n1209 31.8661
R9083 gnd.n6188 gnd.n1209 31.8661
R9084 gnd.n6196 gnd.n1202 31.8661
R9085 gnd.n6196 gnd.n1194 31.8661
R9086 gnd.n6204 gnd.n1194 31.8661
R9087 gnd.n6204 gnd.n1196 31.8661
R9088 gnd.n6212 gnd.n1180 31.8661
R9089 gnd.n6220 gnd.n1180 31.8661
R9090 gnd.n6220 gnd.n1182 31.8661
R9091 gnd.n6996 gnd.n842 31.8661
R9092 gnd.n7012 gnd.n827 31.8661
R9093 gnd.n7012 gnd.n820 31.8661
R9094 gnd.n7020 gnd.n820 31.8661
R9095 gnd.n7028 gnd.n813 31.8661
R9096 gnd.n7028 gnd.n805 31.8661
R9097 gnd.n7036 gnd.n805 31.8661
R9098 gnd.n7036 gnd.n807 31.8661
R9099 gnd.n7044 gnd.n792 31.8661
R9100 gnd.n7055 gnd.n792 31.8661
R9101 gnd.n7055 gnd.n785 31.8661
R9102 gnd.n7063 gnd.n785 31.8661
R9103 gnd.n7094 gnd.n745 31.8661
R9104 gnd.n7094 gnd.n747 31.8661
R9105 gnd.n7077 gnd.n778 31.8661
R9106 gnd.n778 gnd.n571 31.8661
R9107 gnd.n7275 gnd.n551 31.8661
R9108 gnd.n7545 gnd.n376 31.8661
R9109 gnd.n7553 gnd.n368 31.8661
R9110 gnd.n7561 gnd.n358 31.8661
R9111 gnd.n7570 gnd.n358 31.8661
R9112 gnd.n7977 gnd.n106 31.8661
R9113 gnd.n7969 gnd.n121 31.8661
R9114 gnd.n7969 gnd.n124 31.8661
R9115 gnd.n7963 gnd.n135 31.8661
R9116 gnd.n7957 gnd.n135 31.8661
R9117 gnd.n7951 gnd.n150 31.8661
R9118 gnd.n7945 gnd.n160 31.8661
R9119 gnd.n7945 gnd.n163 31.8661
R9120 gnd.n7939 gnd.n172 31.8661
R9121 gnd.n7933 gnd.n172 31.8661
R9122 gnd.n7927 gnd.n188 31.8661
R9123 gnd.n7921 gnd.n198 31.8661
R9124 gnd.n7915 gnd.n210 31.8661
R9125 gnd.n7909 gnd.n210 31.8661
R9126 gnd.n7903 gnd.n226 31.8661
R9127 gnd.n7903 gnd.n229 31.8661
R9128 gnd.n7897 gnd.n229 31.8661
R9129 gnd.n7897 gnd.n239 31.8661
R9130 gnd.n7891 gnd.n248 31.8661
R9131 gnd.n5347 gnd.t265 31.5474
R9132 gnd.t213 gnd.n106 31.5474
R9133 gnd.n6669 gnd.n6665 31.3761
R9134 gnd.n6035 gnd.n1321 31.3761
R9135 gnd.n3649 gnd.t256 30.9101
R9136 gnd.n6228 gnd.n1174 30.9101
R9137 gnd.n7951 gnd.t246 30.9101
R9138 gnd.n1439 gnd.t189 30.5915
R9139 gnd.n5313 gnd.n5312 30.2728
R9140 gnd.n3673 gnd.t238 30.2728
R9141 gnd.n7927 gnd.t347 30.2728
R9142 gnd.n3709 gnd.t131 28.3609
R9143 gnd.n7891 gnd.t113 28.3609
R9144 gnd.n5313 gnd.n3149 27.0862
R9145 gnd.n1182 gnd.t85 27.0862
R9146 gnd.t75 gnd.n827 27.0862
R9147 gnd.n7004 gnd.t128 26.1303
R9148 gnd.n5671 gnd.n5670 25.7944
R9149 gnd.n7109 gnd.n7108 25.7944
R9150 gnd.n4333 gnd.n4332 25.7944
R9151 gnd.n3859 gnd.n3858 25.7944
R9152 gnd.n1238 gnd.n1237 25.7944
R9153 gnd.n630 gnd.n629 25.7944
R9154 gnd.n653 gnd.n652 25.7944
R9155 gnd.n676 gnd.n675 25.7944
R9156 gnd.n351 gnd.n350 25.7944
R9157 gnd.n331 gnd.n330 25.7944
R9158 gnd.n7849 gnd.n7848 25.7944
R9159 gnd.n7668 gnd.n7667 25.7944
R9160 gnd.n3225 gnd.n3224 25.7944
R9161 gnd.n3247 gnd.n3246 25.7944
R9162 gnd.n3269 gnd.n3268 25.7944
R9163 gnd.n3418 gnd.n3417 25.7944
R9164 gnd.n1282 gnd.n1281 25.7944
R9165 gnd.n1481 gnd.n1480 25.7944
R9166 gnd.n1503 gnd.n1502 25.7944
R9167 gnd.n730 gnd.n729 25.7944
R9168 gnd.n4554 gnd.n4274 24.8557
R9169 gnd.n4564 gnd.n4257 24.8557
R9170 gnd.n4260 gnd.n4248 24.8557
R9171 gnd.n4585 gnd.n4249 24.8557
R9172 gnd.n4595 gnd.n4229 24.8557
R9173 gnd.n4605 gnd.n4604 24.8557
R9174 gnd.n4215 gnd.n4213 24.8557
R9175 gnd.n4636 gnd.n4635 24.8557
R9176 gnd.n4651 gnd.n4198 24.8557
R9177 gnd.n4705 gnd.n4137 24.8557
R9178 gnd.n4661 gnd.n4138 24.8557
R9179 gnd.n4698 gnd.n4149 24.8557
R9180 gnd.n4187 gnd.n4186 24.8557
R9181 gnd.n4692 gnd.n4691 24.8557
R9182 gnd.n4173 gnd.n4160 24.8557
R9183 gnd.n4731 gnd.n4730 24.8557
R9184 gnd.n4741 gnd.n4037 24.8557
R9185 gnd.n4753 gnd.n4029 24.8557
R9186 gnd.n4752 gnd.n4017 24.8557
R9187 gnd.n4771 gnd.n4770 24.8557
R9188 gnd.n4781 gnd.n4010 24.8557
R9189 gnd.n4792 gnd.n3998 24.8557
R9190 gnd.n4816 gnd.n4815 24.8557
R9191 gnd.n4827 gnd.n3981 24.8557
R9192 gnd.n4826 gnd.n3983 24.8557
R9193 gnd.n4838 gnd.n3974 24.8557
R9194 gnd.n4856 gnd.n4855 24.8557
R9195 gnd.n3965 gnd.n3954 24.8557
R9196 gnd.n4877 gnd.n3942 24.8557
R9197 gnd.n4905 gnd.n4904 24.8557
R9198 gnd.n4916 gnd.n3927 24.8557
R9199 gnd.n4927 gnd.n3920 24.8557
R9200 gnd.n4926 gnd.n3908 24.8557
R9201 gnd.n5199 gnd.n5198 24.8557
R9202 gnd.n5221 gnd.n3893 24.8557
R9203 gnd.n1231 gnd.t135 24.537
R9204 gnd.n6212 gnd.t10 24.537
R9205 gnd.n7020 gnd.t81 24.537
R9206 gnd.t99 gnd.n745 24.537
R9207 gnd.n7741 gnd.n201 24.537
R9208 gnd.n3605 gnd.n1768 24.2183
R9209 gnd.n5392 gnd.n1740 24.2183
R9210 gnd.n5373 gnd.n1743 24.2183
R9211 gnd.n5385 gnd.n1732 24.2183
R9212 gnd.n5442 gnd.n1702 24.2183
R9213 gnd.n5423 gnd.n1705 24.2183
R9214 gnd.n5435 gnd.n1694 24.2183
R9215 gnd.n5434 gnd.n1714 24.2183
R9216 gnd.n1670 gnd.n1658 24.2183
R9217 gnd.n5468 gnd.n1661 24.2183
R9218 gnd.n5545 gnd.n1637 24.2183
R9219 gnd.n5555 gnd.n1627 24.2183
R9220 gnd.n5538 gnd.n1629 24.2183
R9221 gnd.n5585 gnd.n1611 24.2183
R9222 gnd.n5561 gnd.n1614 24.2183
R9223 gnd.n5595 gnd.n1601 24.2183
R9224 gnd.n5563 gnd.n1603 24.2183
R9225 gnd.n5603 gnd.n1595 24.2183
R9226 gnd.n6152 gnd.n1243 24.2183
R9227 gnd.n7310 gnd.n554 24.2183
R9228 gnd.n7302 gnd.n7301 24.2183
R9229 gnd.n7320 gnd.n544 24.2183
R9230 gnd.n559 gnd.n536 24.2183
R9231 gnd.n7329 gnd.n522 24.2183
R9232 gnd.n7352 gnd.n525 24.2183
R9233 gnd.n7362 gnd.n514 24.2183
R9234 gnd.n7372 gnd.n504 24.2183
R9235 gnd.n7401 gnd.n489 24.2183
R9236 gnd.n7338 gnd.n477 24.2183
R9237 gnd.n7394 gnd.n470 24.2183
R9238 gnd.n7438 gnd.n459 24.2183
R9239 gnd.n7424 gnd.n446 24.2183
R9240 gnd.n7458 gnd.n438 24.2183
R9241 gnd.n7457 gnd.n421 24.2183
R9242 gnd.n7471 gnd.n411 24.2183
R9243 gnd.n7509 gnd.n403 24.2183
R9244 gnd.n7508 gnd.n383 24.2183
R9245 gnd.n7519 gnd.n7518 24.2183
R9246 gnd.n5738 gnd.n1229 23.8997
R9247 gnd.n7078 gnd.n747 23.8997
R9248 gnd.n4575 gnd.t411 23.2624
R9249 gnd.t217 gnd.n3301 23.2624
R9250 gnd.n5384 gnd.t235 23.2624
R9251 gnd.n5577 gnd.t227 23.2624
R9252 gnd.n7333 gnd.t244 23.2624
R9253 gnd.n7470 gnd.t291 23.2624
R9254 gnd.n226 gnd.t242 23.2624
R9255 gnd.n4276 gnd.t117 22.6251
R9256 gnd.t225 gnd.n3339 22.6251
R9257 gnd.n5477 gnd.t301 22.6251
R9258 gnd.n5486 gnd.t322 22.6251
R9259 gnd.n7393 gnd.t261 22.6251
R9260 gnd.n7420 gnd.t215 22.6251
R9261 gnd.n188 gnd.t263 22.6251
R9262 gnd.n5323 gnd.t307 22.3064
R9263 gnd.n397 gnd.t223 22.3064
R9264 gnd.t211 gnd.n3377 21.9878
R9265 gnd.n5402 gnd.t221 21.9878
R9266 gnd.n7497 gnd.t294 21.9878
R9267 gnd.n150 gnd.t311 21.9878
R9268 gnd.n6030 gnd.n1167 21.6691
R9269 gnd.n5893 gnd.n5845 21.6691
R9270 gnd.n5910 gnd.n5833 21.6691
R9271 gnd.n5918 gnd.n5828 21.6691
R9272 gnd.n5926 gnd.n1102 21.6691
R9273 gnd.n5934 gnd.n1095 21.6691
R9274 gnd.n5942 gnd.n1088 21.6691
R9275 gnd.n6332 gnd.n1079 21.6691
R9276 gnd.n6383 gnd.n1023 21.6691
R9277 gnd.n6900 gnd.n927 21.6691
R9278 gnd.n6888 gnd.n919 21.6691
R9279 gnd.n6880 gnd.n912 21.6691
R9280 gnd.n6873 gnd.n905 21.6691
R9281 gnd.n6865 gnd.n961 21.6691
R9282 gnd.n6859 gnd.n6858 21.6691
R9283 gnd.n6630 gnd.n6599 21.6691
R9284 gnd.n6638 gnd.n862 21.6691
R9285 gnd.n6645 gnd.n855 21.6691
R9286 gnd.t4 gnd.n4281 21.3504
R9287 gnd.t219 gnd.n1784 21.3504
R9288 gnd.n1805 gnd.t283 21.3504
R9289 gnd.n7553 gnd.t240 21.3504
R9290 gnd.n7977 gnd.t209 21.3504
R9291 gnd.t142 gnd.n1153 21.0318
R9292 gnd.t40 gnd.n3955 20.7131
R9293 gnd.n3630 gnd.t269 20.7131
R9294 gnd.t229 gnd.n124 20.7131
R9295 gnd.n5863 gnd.n1143 20.3945
R9296 gnd.n5844 gnd.n1137 20.3945
R9297 gnd.n6600 gnd.n870 20.3945
R9298 gnd.t69 gnd.n3990 20.0758
R9299 gnd.n3365 gnd.t253 20.0758
R9300 gnd.n5839 gnd.t34 20.0758
R9301 gnd.n6621 gnd.t12 20.0758
R9302 gnd.t271 gnd.n163 20.0758
R9303 gnd.n1306 gnd.n1305 19.9763
R9304 gnd.n6560 gnd.n6559 19.9763
R9305 gnd.n1363 gnd.n1362 19.9763
R9306 gnd.n6554 gnd.n6553 19.9763
R9307 gnd.n1333 gnd.t111 19.8005
R9308 gnd.n1333 gnd.t175 19.8005
R9309 gnd.n1332 gnd.t143 19.8005
R9310 gnd.n1332 gnd.t165 19.8005
R9311 gnd.n6522 gnd.t89 19.8005
R9312 gnd.n6522 gnd.t203 19.8005
R9313 gnd.n6521 gnd.t152 19.8005
R9314 gnd.n6521 gnd.t129 19.8005
R9315 gnd.n5517 gnd.n1253 19.7572
R9316 gnd.n7274 gnd.n571 19.7572
R9317 gnd.n1329 gnd.n1328 19.5087
R9318 gnd.n1342 gnd.n1329 19.5087
R9319 gnd.n1340 gnd.n1331 19.5087
R9320 gnd.n6526 gnd.n6520 19.5087
R9321 gnd.n4742 gnd.t30 19.4385
R9322 gnd.n3327 gnd.t278 19.4385
R9323 gnd.n6188 gnd.t63 19.4385
R9324 gnd.n7044 gnd.t20 19.4385
R9325 gnd.n7741 gnd.t233 19.4385
R9326 gnd.n6162 gnd.n1221 19.3944
R9327 gnd.n6174 gnd.n1221 19.3944
R9328 gnd.n6174 gnd.n1219 19.3944
R9329 gnd.n6178 gnd.n1219 19.3944
R9330 gnd.n6178 gnd.n1207 19.3944
R9331 gnd.n6190 gnd.n1207 19.3944
R9332 gnd.n6190 gnd.n1205 19.3944
R9333 gnd.n6194 gnd.n1205 19.3944
R9334 gnd.n6194 gnd.n1192 19.3944
R9335 gnd.n6206 gnd.n1192 19.3944
R9336 gnd.n6206 gnd.n1190 19.3944
R9337 gnd.n6210 gnd.n1190 19.3944
R9338 gnd.n6210 gnd.n1178 19.3944
R9339 gnd.n6222 gnd.n1178 19.3944
R9340 gnd.n6222 gnd.n1176 19.3944
R9341 gnd.n6226 gnd.n1176 19.3944
R9342 gnd.n6226 gnd.n1164 19.3944
R9343 gnd.n6238 gnd.n1164 19.3944
R9344 gnd.n6238 gnd.n1162 19.3944
R9345 gnd.n6242 gnd.n1162 19.3944
R9346 gnd.n6242 gnd.n1149 19.3944
R9347 gnd.n6254 gnd.n1149 19.3944
R9348 gnd.n6254 gnd.n1147 19.3944
R9349 gnd.n6258 gnd.n1147 19.3944
R9350 gnd.n6258 gnd.n1134 19.3944
R9351 gnd.n6270 gnd.n1134 19.3944
R9352 gnd.n6270 gnd.n1132 19.3944
R9353 gnd.n6274 gnd.n1132 19.3944
R9354 gnd.n6274 gnd.n1120 19.3944
R9355 gnd.n6286 gnd.n1120 19.3944
R9356 gnd.n6286 gnd.n1118 19.3944
R9357 gnd.n6290 gnd.n1118 19.3944
R9358 gnd.n6290 gnd.n1107 19.3944
R9359 gnd.n6302 gnd.n1107 19.3944
R9360 gnd.n6302 gnd.n1105 19.3944
R9361 gnd.n6306 gnd.n1105 19.3944
R9362 gnd.n6306 gnd.n1093 19.3944
R9363 gnd.n6318 gnd.n1093 19.3944
R9364 gnd.n6318 gnd.n1091 19.3944
R9365 gnd.n6322 gnd.n1091 19.3944
R9366 gnd.n6322 gnd.n1077 19.3944
R9367 gnd.n6334 gnd.n1077 19.3944
R9368 gnd.n6334 gnd.n1074 19.3944
R9369 gnd.n6344 gnd.n1074 19.3944
R9370 gnd.n6344 gnd.n1075 19.3944
R9371 gnd.n6340 gnd.n1075 19.3944
R9372 gnd.n6340 gnd.n6339 19.3944
R9373 gnd.n6339 gnd.n1037 19.3944
R9374 gnd.n6402 gnd.n1037 19.3944
R9375 gnd.n6402 gnd.n1038 19.3944
R9376 gnd.n6398 gnd.n1038 19.3944
R9377 gnd.n6398 gnd.n6397 19.3944
R9378 gnd.n6397 gnd.n998 19.3944
R9379 gnd.n6460 gnd.n998 19.3944
R9380 gnd.n6460 gnd.n999 19.3944
R9381 gnd.n6456 gnd.n999 19.3944
R9382 gnd.n6456 gnd.n6455 19.3944
R9383 gnd.n6455 gnd.n6454 19.3944
R9384 gnd.n6454 gnd.n6451 19.3944
R9385 gnd.n6451 gnd.n916 19.3944
R9386 gnd.n6910 gnd.n916 19.3944
R9387 gnd.n6910 gnd.n914 19.3944
R9388 gnd.n6914 gnd.n914 19.3944
R9389 gnd.n6914 gnd.n902 19.3944
R9390 gnd.n6926 gnd.n902 19.3944
R9391 gnd.n6926 gnd.n900 19.3944
R9392 gnd.n6930 gnd.n900 19.3944
R9393 gnd.n6930 gnd.n889 19.3944
R9394 gnd.n6942 gnd.n889 19.3944
R9395 gnd.n6942 gnd.n887 19.3944
R9396 gnd.n6946 gnd.n887 19.3944
R9397 gnd.n6946 gnd.n875 19.3944
R9398 gnd.n6958 gnd.n875 19.3944
R9399 gnd.n6958 gnd.n873 19.3944
R9400 gnd.n6962 gnd.n873 19.3944
R9401 gnd.n6962 gnd.n860 19.3944
R9402 gnd.n6974 gnd.n860 19.3944
R9403 gnd.n6974 gnd.n858 19.3944
R9404 gnd.n6978 gnd.n858 19.3944
R9405 gnd.n6978 gnd.n846 19.3944
R9406 gnd.n6990 gnd.n846 19.3944
R9407 gnd.n6990 gnd.n844 19.3944
R9408 gnd.n6994 gnd.n844 19.3944
R9409 gnd.n6994 gnd.n832 19.3944
R9410 gnd.n7006 gnd.n832 19.3944
R9411 gnd.n7006 gnd.n830 19.3944
R9412 gnd.n7010 gnd.n830 19.3944
R9413 gnd.n7010 gnd.n818 19.3944
R9414 gnd.n7022 gnd.n818 19.3944
R9415 gnd.n7022 gnd.n816 19.3944
R9416 gnd.n7026 gnd.n816 19.3944
R9417 gnd.n7026 gnd.n803 19.3944
R9418 gnd.n7038 gnd.n803 19.3944
R9419 gnd.n7038 gnd.n801 19.3944
R9420 gnd.n7042 gnd.n801 19.3944
R9421 gnd.n7042 gnd.n790 19.3944
R9422 gnd.n7057 gnd.n790 19.3944
R9423 gnd.n7057 gnd.n788 19.3944
R9424 gnd.n7061 gnd.n788 19.3944
R9425 gnd.n7061 gnd.n742 19.3944
R9426 gnd.n7096 gnd.n742 19.3944
R9427 gnd.n5675 gnd.n1234 19.3944
R9428 gnd.n6158 gnd.n1234 19.3944
R9429 gnd.n6159 gnd.n6158 19.3944
R9430 gnd.n5741 gnd.n1454 19.3944
R9431 gnd.n5736 gnd.n1454 19.3944
R9432 gnd.n5736 gnd.n1472 19.3944
R9433 gnd.n5732 gnd.n1472 19.3944
R9434 gnd.n5732 gnd.n5731 19.3944
R9435 gnd.n5731 gnd.n5730 19.3944
R9436 gnd.n5730 gnd.n1478 19.3944
R9437 gnd.n5725 gnd.n1478 19.3944
R9438 gnd.n5725 gnd.n5724 19.3944
R9439 gnd.n5724 gnd.n5612 19.3944
R9440 gnd.n5717 gnd.n5612 19.3944
R9441 gnd.n5717 gnd.n5716 19.3944
R9442 gnd.n5716 gnd.n5625 19.3944
R9443 gnd.n5709 gnd.n5625 19.3944
R9444 gnd.n5709 gnd.n5708 19.3944
R9445 gnd.n5708 gnd.n5635 19.3944
R9446 gnd.n5701 gnd.n5635 19.3944
R9447 gnd.n5701 gnd.n5700 19.3944
R9448 gnd.n5700 gnd.n5648 19.3944
R9449 gnd.n5693 gnd.n5648 19.3944
R9450 gnd.n5693 gnd.n5692 19.3944
R9451 gnd.n5692 gnd.n5658 19.3944
R9452 gnd.n5685 gnd.n5658 19.3944
R9453 gnd.n5685 gnd.n5684 19.3944
R9454 gnd.n7151 gnd.n686 19.3944
R9455 gnd.n7151 gnd.n7150 19.3944
R9456 gnd.n7150 gnd.n689 19.3944
R9457 gnd.n7143 gnd.n689 19.3944
R9458 gnd.n7143 gnd.n7142 19.3944
R9459 gnd.n7142 gnd.n699 19.3944
R9460 gnd.n7135 gnd.n699 19.3944
R9461 gnd.n7135 gnd.n7134 19.3944
R9462 gnd.n7134 gnd.n707 19.3944
R9463 gnd.n7127 gnd.n707 19.3944
R9464 gnd.n7127 gnd.n7126 19.3944
R9465 gnd.n7126 gnd.n717 19.3944
R9466 gnd.n7119 gnd.n717 19.3944
R9467 gnd.n7119 gnd.n7118 19.3944
R9468 gnd.n7118 gnd.n725 19.3944
R9469 gnd.n7111 gnd.n725 19.3944
R9470 gnd.n4457 gnd.n4456 19.3944
R9471 gnd.n4456 gnd.n4455 19.3944
R9472 gnd.n4455 gnd.n4454 19.3944
R9473 gnd.n4454 gnd.n4452 19.3944
R9474 gnd.n4452 gnd.n4449 19.3944
R9475 gnd.n4449 gnd.n4448 19.3944
R9476 gnd.n4448 gnd.n4445 19.3944
R9477 gnd.n4445 gnd.n4444 19.3944
R9478 gnd.n4444 gnd.n4441 19.3944
R9479 gnd.n4441 gnd.n4440 19.3944
R9480 gnd.n4440 gnd.n4437 19.3944
R9481 gnd.n4437 gnd.n4436 19.3944
R9482 gnd.n4436 gnd.n4433 19.3944
R9483 gnd.n4433 gnd.n4432 19.3944
R9484 gnd.n4432 gnd.n4429 19.3944
R9485 gnd.n4429 gnd.n4428 19.3944
R9486 gnd.n4428 gnd.n4425 19.3944
R9487 gnd.n4425 gnd.n4424 19.3944
R9488 gnd.n4424 gnd.n4421 19.3944
R9489 gnd.n4421 gnd.n4420 19.3944
R9490 gnd.n4420 gnd.n4417 19.3944
R9491 gnd.n4417 gnd.n4416 19.3944
R9492 gnd.n4413 gnd.n4412 19.3944
R9493 gnd.n4412 gnd.n4368 19.3944
R9494 gnd.n4463 gnd.n4368 19.3944
R9495 gnd.n5229 gnd.n5228 19.3944
R9496 gnd.n5228 gnd.n5225 19.3944
R9497 gnd.n5225 gnd.n5224 19.3944
R9498 gnd.n5274 gnd.n5273 19.3944
R9499 gnd.n5273 gnd.n5272 19.3944
R9500 gnd.n5272 gnd.n5269 19.3944
R9501 gnd.n5269 gnd.n5268 19.3944
R9502 gnd.n5268 gnd.n5265 19.3944
R9503 gnd.n5265 gnd.n5264 19.3944
R9504 gnd.n5264 gnd.n5261 19.3944
R9505 gnd.n5261 gnd.n5260 19.3944
R9506 gnd.n5260 gnd.n5257 19.3944
R9507 gnd.n5257 gnd.n5256 19.3944
R9508 gnd.n5256 gnd.n5253 19.3944
R9509 gnd.n5253 gnd.n5252 19.3944
R9510 gnd.n5252 gnd.n5249 19.3944
R9511 gnd.n5249 gnd.n5248 19.3944
R9512 gnd.n5248 gnd.n5245 19.3944
R9513 gnd.n5245 gnd.n5244 19.3944
R9514 gnd.n5244 gnd.n5241 19.3944
R9515 gnd.n5241 gnd.n5240 19.3944
R9516 gnd.n5240 gnd.n5237 19.3944
R9517 gnd.n5237 gnd.n5236 19.3944
R9518 gnd.n5236 gnd.n5233 19.3944
R9519 gnd.n5233 gnd.n5232 19.3944
R9520 gnd.n4556 gnd.n4265 19.3944
R9521 gnd.n4566 gnd.n4265 19.3944
R9522 gnd.n4567 gnd.n4566 19.3944
R9523 gnd.n4567 gnd.n4246 19.3944
R9524 gnd.n4587 gnd.n4246 19.3944
R9525 gnd.n4587 gnd.n4238 19.3944
R9526 gnd.n4597 gnd.n4238 19.3944
R9527 gnd.n4598 gnd.n4597 19.3944
R9528 gnd.n4599 gnd.n4598 19.3944
R9529 gnd.n4599 gnd.n4221 19.3944
R9530 gnd.n4616 gnd.n4221 19.3944
R9531 gnd.n4619 gnd.n4616 19.3944
R9532 gnd.n4619 gnd.n4618 19.3944
R9533 gnd.n4618 gnd.n4194 19.3944
R9534 gnd.n4658 gnd.n4194 19.3944
R9535 gnd.n4658 gnd.n4191 19.3944
R9536 gnd.n4664 gnd.n4191 19.3944
R9537 gnd.n4665 gnd.n4664 19.3944
R9538 gnd.n4665 gnd.n4189 19.3944
R9539 gnd.n4671 gnd.n4189 19.3944
R9540 gnd.n4674 gnd.n4671 19.3944
R9541 gnd.n4676 gnd.n4674 19.3944
R9542 gnd.n4682 gnd.n4676 19.3944
R9543 gnd.n4682 gnd.n4681 19.3944
R9544 gnd.n4681 gnd.n4032 19.3944
R9545 gnd.n4748 gnd.n4032 19.3944
R9546 gnd.n4749 gnd.n4748 19.3944
R9547 gnd.n4749 gnd.n4025 19.3944
R9548 gnd.n4760 gnd.n4025 19.3944
R9549 gnd.n4761 gnd.n4760 19.3944
R9550 gnd.n4761 gnd.n4008 19.3944
R9551 gnd.n4008 gnd.n4006 19.3944
R9552 gnd.n4785 gnd.n4006 19.3944
R9553 gnd.n4786 gnd.n4785 19.3944
R9554 gnd.n4786 gnd.n3977 19.3944
R9555 gnd.n4833 gnd.n3977 19.3944
R9556 gnd.n4834 gnd.n4833 19.3944
R9557 gnd.n4834 gnd.n3970 19.3944
R9558 gnd.n4845 gnd.n3970 19.3944
R9559 gnd.n4846 gnd.n4845 19.3944
R9560 gnd.n4846 gnd.n3953 19.3944
R9561 gnd.n3953 gnd.n3951 19.3944
R9562 gnd.n4870 gnd.n3951 19.3944
R9563 gnd.n4871 gnd.n4870 19.3944
R9564 gnd.n4871 gnd.n3923 19.3944
R9565 gnd.n4922 gnd.n3923 19.3944
R9566 gnd.n4923 gnd.n4922 19.3944
R9567 gnd.n4923 gnd.n3916 19.3944
R9568 gnd.n5190 gnd.n3916 19.3944
R9569 gnd.n5191 gnd.n5190 19.3944
R9570 gnd.n5191 gnd.n3897 19.3944
R9571 gnd.n5216 gnd.n3897 19.3944
R9572 gnd.n5216 gnd.n3898 19.3944
R9573 gnd.n4547 gnd.n4546 19.3944
R9574 gnd.n4546 gnd.n4279 19.3944
R9575 gnd.n4302 gnd.n4279 19.3944
R9576 gnd.n4305 gnd.n4302 19.3944
R9577 gnd.n4305 gnd.n4298 19.3944
R9578 gnd.n4309 gnd.n4298 19.3944
R9579 gnd.n4312 gnd.n4309 19.3944
R9580 gnd.n4315 gnd.n4312 19.3944
R9581 gnd.n4315 gnd.n4296 19.3944
R9582 gnd.n4319 gnd.n4296 19.3944
R9583 gnd.n4322 gnd.n4319 19.3944
R9584 gnd.n4325 gnd.n4322 19.3944
R9585 gnd.n4325 gnd.n4294 19.3944
R9586 gnd.n4329 gnd.n4294 19.3944
R9587 gnd.n4552 gnd.n4551 19.3944
R9588 gnd.n4551 gnd.n4255 19.3944
R9589 gnd.n4577 gnd.n4255 19.3944
R9590 gnd.n4577 gnd.n4253 19.3944
R9591 gnd.n4583 gnd.n4253 19.3944
R9592 gnd.n4583 gnd.n4582 19.3944
R9593 gnd.n4582 gnd.n4227 19.3944
R9594 gnd.n4607 gnd.n4227 19.3944
R9595 gnd.n4607 gnd.n4225 19.3944
R9596 gnd.n4611 gnd.n4225 19.3944
R9597 gnd.n4611 gnd.n4205 19.3944
R9598 gnd.n4638 gnd.n4205 19.3944
R9599 gnd.n4638 gnd.n4203 19.3944
R9600 gnd.n4648 gnd.n4203 19.3944
R9601 gnd.n4648 gnd.n4647 19.3944
R9602 gnd.n4647 gnd.n4646 19.3944
R9603 gnd.n4646 gnd.n4152 19.3944
R9604 gnd.n4696 gnd.n4152 19.3944
R9605 gnd.n4696 gnd.n4695 19.3944
R9606 gnd.n4695 gnd.n4694 19.3944
R9607 gnd.n4694 gnd.n4156 19.3944
R9608 gnd.n4176 gnd.n4156 19.3944
R9609 gnd.n4176 gnd.n4042 19.3944
R9610 gnd.n4733 gnd.n4042 19.3944
R9611 gnd.n4733 gnd.n4040 19.3944
R9612 gnd.n4739 gnd.n4040 19.3944
R9613 gnd.n4739 gnd.n4738 19.3944
R9614 gnd.n4738 gnd.n4015 19.3944
R9615 gnd.n4773 gnd.n4015 19.3944
R9616 gnd.n4773 gnd.n4013 19.3944
R9617 gnd.n4779 gnd.n4013 19.3944
R9618 gnd.n4779 gnd.n4778 19.3944
R9619 gnd.n4778 gnd.n3988 19.3944
R9620 gnd.n4818 gnd.n3988 19.3944
R9621 gnd.n4818 gnd.n3986 19.3944
R9622 gnd.n4824 gnd.n3986 19.3944
R9623 gnd.n4824 gnd.n4823 19.3944
R9624 gnd.n4823 gnd.n3960 19.3944
R9625 gnd.n4858 gnd.n3960 19.3944
R9626 gnd.n4858 gnd.n3958 19.3944
R9627 gnd.n4864 gnd.n3958 19.3944
R9628 gnd.n4864 gnd.n4863 19.3944
R9629 gnd.n4863 gnd.n3933 19.3944
R9630 gnd.n4907 gnd.n3933 19.3944
R9631 gnd.n4907 gnd.n3931 19.3944
R9632 gnd.n4913 gnd.n3931 19.3944
R9633 gnd.n4913 gnd.n4912 19.3944
R9634 gnd.n4912 gnd.n3906 19.3944
R9635 gnd.n5201 gnd.n3906 19.3944
R9636 gnd.n5201 gnd.n3904 19.3944
R9637 gnd.n5209 gnd.n3904 19.3944
R9638 gnd.n5209 gnd.n5208 19.3944
R9639 gnd.n5208 gnd.n5207 19.3944
R9640 gnd.n5310 gnd.n5309 19.3944
R9641 gnd.n5309 gnd.n3845 19.3944
R9642 gnd.n5305 gnd.n3845 19.3944
R9643 gnd.n5305 gnd.n5302 19.3944
R9644 gnd.n5302 gnd.n5299 19.3944
R9645 gnd.n5299 gnd.n5298 19.3944
R9646 gnd.n5298 gnd.n5295 19.3944
R9647 gnd.n5295 gnd.n5294 19.3944
R9648 gnd.n5294 gnd.n5291 19.3944
R9649 gnd.n5291 gnd.n5290 19.3944
R9650 gnd.n5290 gnd.n5287 19.3944
R9651 gnd.n5287 gnd.n5286 19.3944
R9652 gnd.n5286 gnd.n5283 19.3944
R9653 gnd.n5283 gnd.n5282 19.3944
R9654 gnd.n4467 gnd.n4366 19.3944
R9655 gnd.n4467 gnd.n4357 19.3944
R9656 gnd.n4480 gnd.n4357 19.3944
R9657 gnd.n4480 gnd.n4355 19.3944
R9658 gnd.n4484 gnd.n4355 19.3944
R9659 gnd.n4484 gnd.n4345 19.3944
R9660 gnd.n4496 gnd.n4345 19.3944
R9661 gnd.n4496 gnd.n4343 19.3944
R9662 gnd.n4530 gnd.n4343 19.3944
R9663 gnd.n4530 gnd.n4529 19.3944
R9664 gnd.n4529 gnd.n4528 19.3944
R9665 gnd.n4528 gnd.n4527 19.3944
R9666 gnd.n4527 gnd.n4524 19.3944
R9667 gnd.n4524 gnd.n4523 19.3944
R9668 gnd.n4523 gnd.n4522 19.3944
R9669 gnd.n4522 gnd.n4520 19.3944
R9670 gnd.n4520 gnd.n4519 19.3944
R9671 gnd.n4519 gnd.n4516 19.3944
R9672 gnd.n4516 gnd.n4515 19.3944
R9673 gnd.n4515 gnd.n4514 19.3944
R9674 gnd.n4514 gnd.n4512 19.3944
R9675 gnd.n4512 gnd.n4211 19.3944
R9676 gnd.n4627 gnd.n4211 19.3944
R9677 gnd.n4627 gnd.n4209 19.3944
R9678 gnd.n4633 gnd.n4209 19.3944
R9679 gnd.n4633 gnd.n4632 19.3944
R9680 gnd.n4632 gnd.n4133 19.3944
R9681 gnd.n4707 gnd.n4133 19.3944
R9682 gnd.n4707 gnd.n4134 19.3944
R9683 gnd.n4181 gnd.n4180 19.3944
R9684 gnd.n4184 gnd.n4183 19.3944
R9685 gnd.n4171 gnd.n4170 19.3944
R9686 gnd.n4726 gnd.n4047 19.3944
R9687 gnd.n4726 gnd.n4725 19.3944
R9688 gnd.n4725 gnd.n4724 19.3944
R9689 gnd.n4724 gnd.n4722 19.3944
R9690 gnd.n4722 gnd.n4721 19.3944
R9691 gnd.n4721 gnd.n4719 19.3944
R9692 gnd.n4719 gnd.n4718 19.3944
R9693 gnd.n4718 gnd.n3996 19.3944
R9694 gnd.n4794 gnd.n3996 19.3944
R9695 gnd.n4794 gnd.n3994 19.3944
R9696 gnd.n4813 gnd.n3994 19.3944
R9697 gnd.n4813 gnd.n4812 19.3944
R9698 gnd.n4812 gnd.n4811 19.3944
R9699 gnd.n4811 gnd.n4809 19.3944
R9700 gnd.n4809 gnd.n4808 19.3944
R9701 gnd.n4808 gnd.n4806 19.3944
R9702 gnd.n4806 gnd.n4805 19.3944
R9703 gnd.n4805 gnd.n3940 19.3944
R9704 gnd.n4879 gnd.n3940 19.3944
R9705 gnd.n4879 gnd.n3938 19.3944
R9706 gnd.n4902 gnd.n3938 19.3944
R9707 gnd.n4902 gnd.n4901 19.3944
R9708 gnd.n4901 gnd.n4900 19.3944
R9709 gnd.n4900 gnd.n4897 19.3944
R9710 gnd.n4897 gnd.n4896 19.3944
R9711 gnd.n4896 gnd.n4894 19.3944
R9712 gnd.n4894 gnd.n4893 19.3944
R9713 gnd.n4893 gnd.n4891 19.3944
R9714 gnd.n4891 gnd.n3892 19.3944
R9715 gnd.n4472 gnd.n4362 19.3944
R9716 gnd.n4472 gnd.n4360 19.3944
R9717 gnd.n4476 gnd.n4360 19.3944
R9718 gnd.n4476 gnd.n4351 19.3944
R9719 gnd.n4488 gnd.n4351 19.3944
R9720 gnd.n4488 gnd.n4349 19.3944
R9721 gnd.n4492 gnd.n4349 19.3944
R9722 gnd.n4492 gnd.n4338 19.3944
R9723 gnd.n4534 gnd.n4338 19.3944
R9724 gnd.n4534 gnd.n4292 19.3944
R9725 gnd.n4540 gnd.n4292 19.3944
R9726 gnd.n4540 gnd.n4539 19.3944
R9727 gnd.n4539 gnd.n4270 19.3944
R9728 gnd.n4561 gnd.n4270 19.3944
R9729 gnd.n4561 gnd.n4263 19.3944
R9730 gnd.n4572 gnd.n4263 19.3944
R9731 gnd.n4572 gnd.n4571 19.3944
R9732 gnd.n4571 gnd.n4244 19.3944
R9733 gnd.n4592 gnd.n4244 19.3944
R9734 gnd.n4592 gnd.n4234 19.3944
R9735 gnd.n4602 gnd.n4234 19.3944
R9736 gnd.n4602 gnd.n4217 19.3944
R9737 gnd.n4623 gnd.n4217 19.3944
R9738 gnd.n4623 gnd.n4622 19.3944
R9739 gnd.n4622 gnd.n4196 19.3944
R9740 gnd.n4653 gnd.n4196 19.3944
R9741 gnd.n4653 gnd.n4141 19.3944
R9742 gnd.n4703 gnd.n4141 19.3944
R9743 gnd.n4703 gnd.n4702 19.3944
R9744 gnd.n4702 gnd.n4701 19.3944
R9745 gnd.n4701 gnd.n4145 19.3944
R9746 gnd.n4163 gnd.n4145 19.3944
R9747 gnd.n4689 gnd.n4163 19.3944
R9748 gnd.n4689 gnd.n4688 19.3944
R9749 gnd.n4688 gnd.n4687 19.3944
R9750 gnd.n4687 gnd.n4167 19.3944
R9751 gnd.n4167 gnd.n4034 19.3944
R9752 gnd.n4744 gnd.n4034 19.3944
R9753 gnd.n4744 gnd.n4027 19.3944
R9754 gnd.n4755 gnd.n4027 19.3944
R9755 gnd.n4755 gnd.n4023 19.3944
R9756 gnd.n4768 gnd.n4023 19.3944
R9757 gnd.n4768 gnd.n4767 19.3944
R9758 gnd.n4767 gnd.n4002 19.3944
R9759 gnd.n4790 gnd.n4002 19.3944
R9760 gnd.n4790 gnd.n4789 19.3944
R9761 gnd.n4789 gnd.n3979 19.3944
R9762 gnd.n4829 gnd.n3979 19.3944
R9763 gnd.n4829 gnd.n3972 19.3944
R9764 gnd.n4840 gnd.n3972 19.3944
R9765 gnd.n4840 gnd.n3968 19.3944
R9766 gnd.n4853 gnd.n3968 19.3944
R9767 gnd.n4853 gnd.n4852 19.3944
R9768 gnd.n4852 gnd.n3947 19.3944
R9769 gnd.n4875 gnd.n3947 19.3944
R9770 gnd.n4875 gnd.n4874 19.3944
R9771 gnd.n4874 gnd.n3925 19.3944
R9772 gnd.n4918 gnd.n3925 19.3944
R9773 gnd.n4918 gnd.n3918 19.3944
R9774 gnd.n4929 gnd.n3918 19.3944
R9775 gnd.n4929 gnd.n3914 19.3944
R9776 gnd.n5196 gnd.n3914 19.3944
R9777 gnd.n5196 gnd.n5195 19.3944
R9778 gnd.n5195 gnd.n3895 19.3944
R9779 gnd.n5219 gnd.n3895 19.3944
R9780 gnd.n5721 gnd.n5614 19.3944
R9781 gnd.n5721 gnd.n5720 19.3944
R9782 gnd.n5720 gnd.n5619 19.3944
R9783 gnd.n5713 gnd.n5619 19.3944
R9784 gnd.n5713 gnd.n5712 19.3944
R9785 gnd.n5712 gnd.n5631 19.3944
R9786 gnd.n5705 gnd.n5631 19.3944
R9787 gnd.n5705 gnd.n5704 19.3944
R9788 gnd.n5704 gnd.n5642 19.3944
R9789 gnd.n5697 gnd.n5642 19.3944
R9790 gnd.n5697 gnd.n5696 19.3944
R9791 gnd.n5696 gnd.n5654 19.3944
R9792 gnd.n5689 gnd.n5654 19.3944
R9793 gnd.n5689 gnd.n5688 19.3944
R9794 gnd.n5688 gnd.n5665 19.3944
R9795 gnd.n5681 gnd.n5665 19.3944
R9796 gnd.n3602 gnd.n3597 19.3944
R9797 gnd.n3602 gnd.n3598 19.3944
R9798 gnd.n3598 gnd.n1755 19.3944
R9799 gnd.n5376 gnd.n1755 19.3944
R9800 gnd.n5376 gnd.n1753 19.3944
R9801 gnd.n5382 gnd.n1753 19.3944
R9802 gnd.n5382 gnd.n5381 19.3944
R9803 gnd.n5381 gnd.n1720 19.3944
R9804 gnd.n5426 gnd.n1720 19.3944
R9805 gnd.n5426 gnd.n1718 19.3944
R9806 gnd.n5432 gnd.n1718 19.3944
R9807 gnd.n5432 gnd.n5431 19.3944
R9808 gnd.n5431 gnd.n1656 19.3944
R9809 gnd.n5488 gnd.n1656 19.3944
R9810 gnd.n5488 gnd.n1654 19.3944
R9811 gnd.n5492 gnd.n1654 19.3944
R9812 gnd.n5492 gnd.n1652 19.3944
R9813 gnd.n5496 gnd.n1652 19.3944
R9814 gnd.n5496 gnd.n1650 19.3944
R9815 gnd.n5535 gnd.n1650 19.3944
R9816 gnd.n5535 gnd.n5534 19.3944
R9817 gnd.n5534 gnd.n5533 19.3944
R9818 gnd.n5533 gnd.n5502 19.3944
R9819 gnd.n5529 gnd.n5502 19.3944
R9820 gnd.n5529 gnd.n5528 19.3944
R9821 gnd.n5528 gnd.n5527 19.3944
R9822 gnd.n5527 gnd.n5508 19.3944
R9823 gnd.n5522 gnd.n5508 19.3944
R9824 gnd.n5522 gnd.n5521 19.3944
R9825 gnd.n5521 gnd.n5520 19.3944
R9826 gnd.n5520 gnd.n5515 19.3944
R9827 gnd.n5515 gnd.n1227 19.3944
R9828 gnd.n6166 gnd.n1227 19.3944
R9829 gnd.n6166 gnd.n1225 19.3944
R9830 gnd.n6170 gnd.n1225 19.3944
R9831 gnd.n6170 gnd.n1214 19.3944
R9832 gnd.n6182 gnd.n1214 19.3944
R9833 gnd.n6182 gnd.n1212 19.3944
R9834 gnd.n6186 gnd.n1212 19.3944
R9835 gnd.n6186 gnd.n1200 19.3944
R9836 gnd.n6198 gnd.n1200 19.3944
R9837 gnd.n6198 gnd.n1198 19.3944
R9838 gnd.n6202 gnd.n1198 19.3944
R9839 gnd.n6202 gnd.n1186 19.3944
R9840 gnd.n6214 gnd.n1186 19.3944
R9841 gnd.n6214 gnd.n1184 19.3944
R9842 gnd.n6218 gnd.n1184 19.3944
R9843 gnd.n6218 gnd.n1171 19.3944
R9844 gnd.n6230 gnd.n1171 19.3944
R9845 gnd.n6230 gnd.n1169 19.3944
R9846 gnd.n6234 gnd.n1169 19.3944
R9847 gnd.n6234 gnd.n1157 19.3944
R9848 gnd.n6246 gnd.n1157 19.3944
R9849 gnd.n6246 gnd.n1155 19.3944
R9850 gnd.n6250 gnd.n1155 19.3944
R9851 gnd.n6250 gnd.n1141 19.3944
R9852 gnd.n6262 gnd.n1141 19.3944
R9853 gnd.n6262 gnd.n1139 19.3944
R9854 gnd.n6266 gnd.n1139 19.3944
R9855 gnd.n6266 gnd.n1127 19.3944
R9856 gnd.n6278 gnd.n1127 19.3944
R9857 gnd.n6278 gnd.n1125 19.3944
R9858 gnd.n6282 gnd.n1125 19.3944
R9859 gnd.n6282 gnd.n1113 19.3944
R9860 gnd.n6294 gnd.n1113 19.3944
R9861 gnd.n6294 gnd.n1111 19.3944
R9862 gnd.n6298 gnd.n1111 19.3944
R9863 gnd.n6298 gnd.n1100 19.3944
R9864 gnd.n6310 gnd.n1100 19.3944
R9865 gnd.n6310 gnd.n1098 19.3944
R9866 gnd.n6314 gnd.n1098 19.3944
R9867 gnd.n6314 gnd.n1086 19.3944
R9868 gnd.n6326 gnd.n1086 19.3944
R9869 gnd.n6326 gnd.n1084 19.3944
R9870 gnd.n6330 gnd.n1084 19.3944
R9871 gnd.n6330 gnd.n1068 19.3944
R9872 gnd.n6348 gnd.n1068 19.3944
R9873 gnd.n6348 gnd.n1066 19.3944
R9874 gnd.n6354 gnd.n1066 19.3944
R9875 gnd.n6354 gnd.n6353 19.3944
R9876 gnd.n6353 gnd.n1030 19.3944
R9877 gnd.n6406 gnd.n1030 19.3944
R9878 gnd.n6406 gnd.n1028 19.3944
R9879 gnd.n6412 gnd.n1028 19.3944
R9880 gnd.n6412 gnd.n6411 19.3944
R9881 gnd.n6411 gnd.n991 19.3944
R9882 gnd.n6464 gnd.n991 19.3944
R9883 gnd.n6464 gnd.n989 19.3944
R9884 gnd.n6470 gnd.n989 19.3944
R9885 gnd.n6470 gnd.n6469 19.3944
R9886 gnd.n6469 gnd.n923 19.3944
R9887 gnd.n6902 gnd.n923 19.3944
R9888 gnd.n6902 gnd.n921 19.3944
R9889 gnd.n6906 gnd.n921 19.3944
R9890 gnd.n6906 gnd.n909 19.3944
R9891 gnd.n6918 gnd.n909 19.3944
R9892 gnd.n6918 gnd.n907 19.3944
R9893 gnd.n6922 gnd.n907 19.3944
R9894 gnd.n6922 gnd.n896 19.3944
R9895 gnd.n6934 gnd.n896 19.3944
R9896 gnd.n6934 gnd.n894 19.3944
R9897 gnd.n6938 gnd.n894 19.3944
R9898 gnd.n6938 gnd.n882 19.3944
R9899 gnd.n6950 gnd.n882 19.3944
R9900 gnd.n6950 gnd.n880 19.3944
R9901 gnd.n6954 gnd.n880 19.3944
R9902 gnd.n6954 gnd.n868 19.3944
R9903 gnd.n6966 gnd.n868 19.3944
R9904 gnd.n6966 gnd.n866 19.3944
R9905 gnd.n6970 gnd.n866 19.3944
R9906 gnd.n6970 gnd.n853 19.3944
R9907 gnd.n6982 gnd.n853 19.3944
R9908 gnd.n6982 gnd.n851 19.3944
R9909 gnd.n6986 gnd.n851 19.3944
R9910 gnd.n6986 gnd.n838 19.3944
R9911 gnd.n6998 gnd.n838 19.3944
R9912 gnd.n6998 gnd.n836 19.3944
R9913 gnd.n7002 gnd.n836 19.3944
R9914 gnd.n7002 gnd.n825 19.3944
R9915 gnd.n7014 gnd.n825 19.3944
R9916 gnd.n7014 gnd.n823 19.3944
R9917 gnd.n7018 gnd.n823 19.3944
R9918 gnd.n7018 gnd.n811 19.3944
R9919 gnd.n7030 gnd.n811 19.3944
R9920 gnd.n7030 gnd.n809 19.3944
R9921 gnd.n7034 gnd.n809 19.3944
R9922 gnd.n7034 gnd.n797 19.3944
R9923 gnd.n7046 gnd.n797 19.3944
R9924 gnd.n7046 gnd.n795 19.3944
R9925 gnd.n7053 gnd.n795 19.3944
R9926 gnd.n7053 gnd.n7052 19.3944
R9927 gnd.n7052 gnd.n783 19.3944
R9928 gnd.n7066 gnd.n783 19.3944
R9929 gnd.n7067 gnd.n7066 19.3944
R9930 gnd.n7067 gnd.n781 19.3944
R9931 gnd.n7075 gnd.n781 19.3944
R9932 gnd.n7075 gnd.n7074 19.3944
R9933 gnd.n7074 gnd.n7073 19.3944
R9934 gnd.n7073 gnd.n569 19.3944
R9935 gnd.n7278 gnd.n569 19.3944
R9936 gnd.n7278 gnd.n567 19.3944
R9937 gnd.n7299 gnd.n567 19.3944
R9938 gnd.n7299 gnd.n7298 19.3944
R9939 gnd.n7298 gnd.n7297 19.3944
R9940 gnd.n7297 gnd.n7284 19.3944
R9941 gnd.n7293 gnd.n7284 19.3944
R9942 gnd.n7293 gnd.n7292 19.3944
R9943 gnd.n7292 gnd.n7291 19.3944
R9944 gnd.n7291 gnd.n503 19.3944
R9945 gnd.n503 gnd.n501 19.3944
R9946 gnd.n7376 gnd.n501 19.3944
R9947 gnd.n7376 gnd.n499 19.3944
R9948 gnd.n7391 gnd.n499 19.3944
R9949 gnd.n7391 gnd.n7390 19.3944
R9950 gnd.n7390 gnd.n7389 19.3944
R9951 gnd.n7389 gnd.n7382 19.3944
R9952 gnd.n7385 gnd.n7382 19.3944
R9953 gnd.n7385 gnd.n436 19.3944
R9954 gnd.n7460 gnd.n436 19.3944
R9955 gnd.n7460 gnd.n434 19.3944
R9956 gnd.n7468 gnd.n434 19.3944
R9957 gnd.n7468 gnd.n7467 19.3944
R9958 gnd.n7467 gnd.n7466 19.3944
R9959 gnd.n7466 gnd.n401 19.3944
R9960 gnd.n7512 gnd.n401 19.3944
R9961 gnd.n7512 gnd.n399 19.3944
R9962 gnd.n7516 gnd.n399 19.3944
R9963 gnd.n2604 gnd.n2603 19.3944
R9964 gnd.n2603 gnd.n2602 19.3944
R9965 gnd.n2602 gnd.n2273 19.3944
R9966 gnd.n2596 gnd.n2273 19.3944
R9967 gnd.n2596 gnd.n2595 19.3944
R9968 gnd.n2595 gnd.n2594 19.3944
R9969 gnd.n2594 gnd.n2282 19.3944
R9970 gnd.n2588 gnd.n2282 19.3944
R9971 gnd.n2588 gnd.n2587 19.3944
R9972 gnd.n2587 gnd.n2586 19.3944
R9973 gnd.n2586 gnd.n2290 19.3944
R9974 gnd.n2580 gnd.n2290 19.3944
R9975 gnd.n2580 gnd.n2579 19.3944
R9976 gnd.n2579 gnd.n2578 19.3944
R9977 gnd.n2578 gnd.n2298 19.3944
R9978 gnd.n2572 gnd.n2298 19.3944
R9979 gnd.n2572 gnd.n2571 19.3944
R9980 gnd.n2571 gnd.n2570 19.3944
R9981 gnd.n2570 gnd.n2306 19.3944
R9982 gnd.n2564 gnd.n2306 19.3944
R9983 gnd.n2564 gnd.n2563 19.3944
R9984 gnd.n2563 gnd.n2562 19.3944
R9985 gnd.n2562 gnd.n2314 19.3944
R9986 gnd.n2556 gnd.n2314 19.3944
R9987 gnd.n2556 gnd.n2555 19.3944
R9988 gnd.n2555 gnd.n2554 19.3944
R9989 gnd.n2554 gnd.n2322 19.3944
R9990 gnd.n2548 gnd.n2322 19.3944
R9991 gnd.n2548 gnd.n2547 19.3944
R9992 gnd.n2547 gnd.n2546 19.3944
R9993 gnd.n2546 gnd.n2330 19.3944
R9994 gnd.n2540 gnd.n2330 19.3944
R9995 gnd.n2540 gnd.n2539 19.3944
R9996 gnd.n2539 gnd.n2538 19.3944
R9997 gnd.n2538 gnd.n2338 19.3944
R9998 gnd.n2532 gnd.n2338 19.3944
R9999 gnd.n2532 gnd.n2531 19.3944
R10000 gnd.n2531 gnd.n2530 19.3944
R10001 gnd.n2530 gnd.n2346 19.3944
R10002 gnd.n2524 gnd.n2346 19.3944
R10003 gnd.n2524 gnd.n2523 19.3944
R10004 gnd.n2523 gnd.n2522 19.3944
R10005 gnd.n2522 gnd.n2354 19.3944
R10006 gnd.n2516 gnd.n2354 19.3944
R10007 gnd.n2516 gnd.n2515 19.3944
R10008 gnd.n2515 gnd.n2514 19.3944
R10009 gnd.n2514 gnd.n2362 19.3944
R10010 gnd.n2508 gnd.n2362 19.3944
R10011 gnd.n2508 gnd.n2507 19.3944
R10012 gnd.n2507 gnd.n2506 19.3944
R10013 gnd.n2506 gnd.n2370 19.3944
R10014 gnd.n2500 gnd.n2370 19.3944
R10015 gnd.n2500 gnd.n2499 19.3944
R10016 gnd.n2499 gnd.n2498 19.3944
R10017 gnd.n2498 gnd.n2378 19.3944
R10018 gnd.n2492 gnd.n2378 19.3944
R10019 gnd.n2492 gnd.n2491 19.3944
R10020 gnd.n2491 gnd.n2490 19.3944
R10021 gnd.n2490 gnd.n2386 19.3944
R10022 gnd.n2484 gnd.n2386 19.3944
R10023 gnd.n2484 gnd.n2483 19.3944
R10024 gnd.n2483 gnd.n2482 19.3944
R10025 gnd.n2482 gnd.n2394 19.3944
R10026 gnd.n2476 gnd.n2394 19.3944
R10027 gnd.n2476 gnd.n2475 19.3944
R10028 gnd.n2475 gnd.n2474 19.3944
R10029 gnd.n2474 gnd.n2402 19.3944
R10030 gnd.n2468 gnd.n2402 19.3944
R10031 gnd.n2468 gnd.n2467 19.3944
R10032 gnd.n2467 gnd.n2466 19.3944
R10033 gnd.n2466 gnd.n2410 19.3944
R10034 gnd.n2460 gnd.n2410 19.3944
R10035 gnd.n2460 gnd.n2459 19.3944
R10036 gnd.n2459 gnd.n2458 19.3944
R10037 gnd.n2458 gnd.n2418 19.3944
R10038 gnd.n2452 gnd.n2418 19.3944
R10039 gnd.n2452 gnd.n2451 19.3944
R10040 gnd.n2451 gnd.n2450 19.3944
R10041 gnd.n2450 gnd.n2426 19.3944
R10042 gnd.n2444 gnd.n2426 19.3944
R10043 gnd.n2444 gnd.n2443 19.3944
R10044 gnd.n2443 gnd.n2442 19.3944
R10045 gnd.n2442 gnd.n2437 19.3944
R10046 gnd.n2437 gnd.n2436 19.3944
R10047 gnd.n2942 gnd.n2941 19.3944
R10048 gnd.n2941 gnd.n1937 19.3944
R10049 gnd.n2935 gnd.n1937 19.3944
R10050 gnd.n2935 gnd.n2934 19.3944
R10051 gnd.n2934 gnd.n2933 19.3944
R10052 gnd.n2933 gnd.n1945 19.3944
R10053 gnd.n2927 gnd.n1945 19.3944
R10054 gnd.n2927 gnd.n2926 19.3944
R10055 gnd.n2926 gnd.n2925 19.3944
R10056 gnd.n2925 gnd.n1953 19.3944
R10057 gnd.n2919 gnd.n1953 19.3944
R10058 gnd.n2919 gnd.n2918 19.3944
R10059 gnd.n2918 gnd.n2917 19.3944
R10060 gnd.n2917 gnd.n1961 19.3944
R10061 gnd.n2911 gnd.n1961 19.3944
R10062 gnd.n2911 gnd.n2910 19.3944
R10063 gnd.n2910 gnd.n2909 19.3944
R10064 gnd.n2909 gnd.n1969 19.3944
R10065 gnd.n2903 gnd.n1969 19.3944
R10066 gnd.n2903 gnd.n2902 19.3944
R10067 gnd.n2902 gnd.n2901 19.3944
R10068 gnd.n2901 gnd.n1977 19.3944
R10069 gnd.n2895 gnd.n1977 19.3944
R10070 gnd.n2895 gnd.n2894 19.3944
R10071 gnd.n2894 gnd.n2893 19.3944
R10072 gnd.n2893 gnd.n1985 19.3944
R10073 gnd.n2887 gnd.n1985 19.3944
R10074 gnd.n2887 gnd.n2886 19.3944
R10075 gnd.n2886 gnd.n2885 19.3944
R10076 gnd.n2885 gnd.n1993 19.3944
R10077 gnd.n2879 gnd.n1993 19.3944
R10078 gnd.n2879 gnd.n2878 19.3944
R10079 gnd.n2878 gnd.n2877 19.3944
R10080 gnd.n2877 gnd.n2001 19.3944
R10081 gnd.n2871 gnd.n2001 19.3944
R10082 gnd.n2871 gnd.n2870 19.3944
R10083 gnd.n2870 gnd.n2869 19.3944
R10084 gnd.n2869 gnd.n2009 19.3944
R10085 gnd.n2863 gnd.n2009 19.3944
R10086 gnd.n2863 gnd.n2862 19.3944
R10087 gnd.n2862 gnd.n2861 19.3944
R10088 gnd.n2861 gnd.n2017 19.3944
R10089 gnd.n2855 gnd.n2017 19.3944
R10090 gnd.n2855 gnd.n2854 19.3944
R10091 gnd.n2854 gnd.n2853 19.3944
R10092 gnd.n2853 gnd.n2025 19.3944
R10093 gnd.n2847 gnd.n2025 19.3944
R10094 gnd.n2847 gnd.n2846 19.3944
R10095 gnd.n2846 gnd.n2845 19.3944
R10096 gnd.n2845 gnd.n2033 19.3944
R10097 gnd.n2839 gnd.n2033 19.3944
R10098 gnd.n2839 gnd.n2838 19.3944
R10099 gnd.n2838 gnd.n2837 19.3944
R10100 gnd.n2837 gnd.n2041 19.3944
R10101 gnd.n2831 gnd.n2041 19.3944
R10102 gnd.n2831 gnd.n2830 19.3944
R10103 gnd.n2830 gnd.n2829 19.3944
R10104 gnd.n2829 gnd.n2049 19.3944
R10105 gnd.n2823 gnd.n2049 19.3944
R10106 gnd.n2823 gnd.n2822 19.3944
R10107 gnd.n2822 gnd.n2821 19.3944
R10108 gnd.n2821 gnd.n2057 19.3944
R10109 gnd.n2815 gnd.n2057 19.3944
R10110 gnd.n2815 gnd.n2814 19.3944
R10111 gnd.n2814 gnd.n2813 19.3944
R10112 gnd.n2813 gnd.n2065 19.3944
R10113 gnd.n2807 gnd.n2065 19.3944
R10114 gnd.n2807 gnd.n2806 19.3944
R10115 gnd.n2806 gnd.n2805 19.3944
R10116 gnd.n2805 gnd.n2073 19.3944
R10117 gnd.n2799 gnd.n2073 19.3944
R10118 gnd.n2799 gnd.n2798 19.3944
R10119 gnd.n2798 gnd.n2797 19.3944
R10120 gnd.n2797 gnd.n2081 19.3944
R10121 gnd.n2791 gnd.n2081 19.3944
R10122 gnd.n2791 gnd.n2790 19.3944
R10123 gnd.n2790 gnd.n2789 19.3944
R10124 gnd.n2789 gnd.n2089 19.3944
R10125 gnd.n2783 gnd.n2089 19.3944
R10126 gnd.n2783 gnd.n2782 19.3944
R10127 gnd.n2782 gnd.n2781 19.3944
R10128 gnd.n2781 gnd.n2097 19.3944
R10129 gnd.n2775 gnd.n2097 19.3944
R10130 gnd.n2775 gnd.n2774 19.3944
R10131 gnd.n2774 gnd.n2773 19.3944
R10132 gnd.n2773 gnd.n2105 19.3944
R10133 gnd.n2767 gnd.n2105 19.3944
R10134 gnd.n2767 gnd.n2766 19.3944
R10135 gnd.n2766 gnd.n2765 19.3944
R10136 gnd.n2765 gnd.n2113 19.3944
R10137 gnd.n2759 gnd.n2113 19.3944
R10138 gnd.n2759 gnd.n2758 19.3944
R10139 gnd.n2758 gnd.n2757 19.3944
R10140 gnd.n2757 gnd.n2121 19.3944
R10141 gnd.n2751 gnd.n2121 19.3944
R10142 gnd.n2751 gnd.n2750 19.3944
R10143 gnd.n2750 gnd.n2749 19.3944
R10144 gnd.n2749 gnd.n2129 19.3944
R10145 gnd.n2743 gnd.n2129 19.3944
R10146 gnd.n2743 gnd.n2742 19.3944
R10147 gnd.n2742 gnd.n2741 19.3944
R10148 gnd.n2741 gnd.n2137 19.3944
R10149 gnd.n2735 gnd.n2137 19.3944
R10150 gnd.n2735 gnd.n2734 19.3944
R10151 gnd.n2734 gnd.n2733 19.3944
R10152 gnd.n2733 gnd.n2145 19.3944
R10153 gnd.n2727 gnd.n2145 19.3944
R10154 gnd.n2727 gnd.n2726 19.3944
R10155 gnd.n2726 gnd.n2725 19.3944
R10156 gnd.n2725 gnd.n2153 19.3944
R10157 gnd.n2719 gnd.n2153 19.3944
R10158 gnd.n2719 gnd.n2718 19.3944
R10159 gnd.n2718 gnd.n2717 19.3944
R10160 gnd.n2717 gnd.n2161 19.3944
R10161 gnd.n2711 gnd.n2161 19.3944
R10162 gnd.n2711 gnd.n2710 19.3944
R10163 gnd.n2710 gnd.n2709 19.3944
R10164 gnd.n2709 gnd.n2169 19.3944
R10165 gnd.n2703 gnd.n2169 19.3944
R10166 gnd.n2703 gnd.n2702 19.3944
R10167 gnd.n2702 gnd.n2701 19.3944
R10168 gnd.n2701 gnd.n2177 19.3944
R10169 gnd.n2695 gnd.n2177 19.3944
R10170 gnd.n2695 gnd.n2694 19.3944
R10171 gnd.n2694 gnd.n2693 19.3944
R10172 gnd.n2693 gnd.n2185 19.3944
R10173 gnd.n2687 gnd.n2185 19.3944
R10174 gnd.n2687 gnd.n2686 19.3944
R10175 gnd.n2686 gnd.n2685 19.3944
R10176 gnd.n2685 gnd.n2193 19.3944
R10177 gnd.n2679 gnd.n2193 19.3944
R10178 gnd.n2679 gnd.n2678 19.3944
R10179 gnd.n2678 gnd.n2677 19.3944
R10180 gnd.n2677 gnd.n2201 19.3944
R10181 gnd.n2671 gnd.n2201 19.3944
R10182 gnd.n2671 gnd.n2670 19.3944
R10183 gnd.n2670 gnd.n2669 19.3944
R10184 gnd.n2669 gnd.n2209 19.3944
R10185 gnd.n2663 gnd.n2209 19.3944
R10186 gnd.n2663 gnd.n2662 19.3944
R10187 gnd.n2662 gnd.n2661 19.3944
R10188 gnd.n2661 gnd.n2217 19.3944
R10189 gnd.n2655 gnd.n2217 19.3944
R10190 gnd.n2655 gnd.n2654 19.3944
R10191 gnd.n2654 gnd.n2653 19.3944
R10192 gnd.n2653 gnd.n2225 19.3944
R10193 gnd.n2647 gnd.n2225 19.3944
R10194 gnd.n2647 gnd.n2646 19.3944
R10195 gnd.n2646 gnd.n2645 19.3944
R10196 gnd.n2645 gnd.n2233 19.3944
R10197 gnd.n2639 gnd.n2233 19.3944
R10198 gnd.n2639 gnd.n2638 19.3944
R10199 gnd.n2638 gnd.n2637 19.3944
R10200 gnd.n2637 gnd.n2241 19.3944
R10201 gnd.n2631 gnd.n2241 19.3944
R10202 gnd.n2631 gnd.n2630 19.3944
R10203 gnd.n2630 gnd.n2629 19.3944
R10204 gnd.n2629 gnd.n2249 19.3944
R10205 gnd.n2623 gnd.n2249 19.3944
R10206 gnd.n2623 gnd.n2622 19.3944
R10207 gnd.n2622 gnd.n2621 19.3944
R10208 gnd.n2621 gnd.n2257 19.3944
R10209 gnd.n2615 gnd.n2257 19.3944
R10210 gnd.n2615 gnd.n2614 19.3944
R10211 gnd.n2614 gnd.n2613 19.3944
R10212 gnd.n2613 gnd.n2265 19.3944
R10213 gnd.n2607 gnd.n2265 19.3944
R10214 gnd.n7271 gnd.n611 19.3944
R10215 gnd.n7271 gnd.n7270 19.3944
R10216 gnd.n7270 gnd.n7269 19.3944
R10217 gnd.n7269 gnd.n7267 19.3944
R10218 gnd.n7267 gnd.n7264 19.3944
R10219 gnd.n7264 gnd.n7263 19.3944
R10220 gnd.n7263 gnd.n7260 19.3944
R10221 gnd.n7260 gnd.n7259 19.3944
R10222 gnd.n7259 gnd.n7256 19.3944
R10223 gnd.n7256 gnd.n7255 19.3944
R10224 gnd.n7255 gnd.n7252 19.3944
R10225 gnd.n7252 gnd.n7251 19.3944
R10226 gnd.n7251 gnd.n7248 19.3944
R10227 gnd.n7248 gnd.n7247 19.3944
R10228 gnd.n7247 gnd.n7244 19.3944
R10229 gnd.n7244 gnd.n7243 19.3944
R10230 gnd.n7243 gnd.n7240 19.3944
R10231 gnd.n7238 gnd.n7235 19.3944
R10232 gnd.n7235 gnd.n7234 19.3944
R10233 gnd.n7234 gnd.n7231 19.3944
R10234 gnd.n7231 gnd.n7230 19.3944
R10235 gnd.n7230 gnd.n7227 19.3944
R10236 gnd.n7227 gnd.n7226 19.3944
R10237 gnd.n7226 gnd.n7223 19.3944
R10238 gnd.n7221 gnd.n7218 19.3944
R10239 gnd.n7218 gnd.n7217 19.3944
R10240 gnd.n7217 gnd.n7214 19.3944
R10241 gnd.n7214 gnd.n7213 19.3944
R10242 gnd.n7213 gnd.n7210 19.3944
R10243 gnd.n7210 gnd.n7209 19.3944
R10244 gnd.n7209 gnd.n7206 19.3944
R10245 gnd.n7206 gnd.n7205 19.3944
R10246 gnd.n7201 gnd.n7198 19.3944
R10247 gnd.n7198 gnd.n7197 19.3944
R10248 gnd.n7197 gnd.n7194 19.3944
R10249 gnd.n7194 gnd.n7193 19.3944
R10250 gnd.n7193 gnd.n7190 19.3944
R10251 gnd.n7190 gnd.n7189 19.3944
R10252 gnd.n7189 gnd.n7186 19.3944
R10253 gnd.n7186 gnd.n7185 19.3944
R10254 gnd.n7185 gnd.n7182 19.3944
R10255 gnd.n7182 gnd.n7181 19.3944
R10256 gnd.n7181 gnd.n7178 19.3944
R10257 gnd.n7178 gnd.n7177 19.3944
R10258 gnd.n7177 gnd.n7174 19.3944
R10259 gnd.n7174 gnd.n7173 19.3944
R10260 gnd.n7173 gnd.n7170 19.3944
R10261 gnd.n7170 gnd.n7169 19.3944
R10262 gnd.n7169 gnd.n7166 19.3944
R10263 gnd.n7166 gnd.n7165 19.3944
R10264 gnd.n7305 gnd.n564 19.3944
R10265 gnd.n7305 gnd.n7304 19.3944
R10266 gnd.n7304 gnd.n533 19.3944
R10267 gnd.n7331 gnd.n533 19.3944
R10268 gnd.n7332 gnd.n7331 19.3944
R10269 gnd.n7335 gnd.n7332 19.3944
R10270 gnd.n7336 gnd.n7335 19.3944
R10271 gnd.n7344 gnd.n7336 19.3944
R10272 gnd.n7344 gnd.n7342 19.3944
R10273 gnd.n7342 gnd.n7341 19.3944
R10274 gnd.n7341 gnd.n7340 19.3944
R10275 gnd.n7340 gnd.n7337 19.3944
R10276 gnd.n7337 gnd.n467 19.3944
R10277 gnd.n7422 gnd.n467 19.3944
R10278 gnd.n7423 gnd.n7422 19.3944
R10279 gnd.n7426 gnd.n7423 19.3944
R10280 gnd.n7427 gnd.n7426 19.3944
R10281 gnd.n7430 gnd.n7427 19.3944
R10282 gnd.n7430 gnd.n7428 19.3944
R10283 gnd.n7428 gnd.n431 19.3944
R10284 gnd.n7473 gnd.n431 19.3944
R10285 gnd.n7474 gnd.n7473 19.3944
R10286 gnd.n7478 gnd.n7474 19.3944
R10287 gnd.n7478 gnd.n7476 19.3944
R10288 gnd.n7476 gnd.n7475 19.3944
R10289 gnd.n7475 gnd.n393 19.3944
R10290 gnd.n7522 gnd.n393 19.3944
R10291 gnd.n7523 gnd.n7522 19.3944
R10292 gnd.n7526 gnd.n7523 19.3944
R10293 gnd.n7526 gnd.n7524 19.3944
R10294 gnd.n7524 gnd.n360 19.3944
R10295 gnd.n7566 gnd.n360 19.3944
R10296 gnd.n7568 gnd.n7566 19.3944
R10297 gnd.n7568 gnd.n7567 19.3944
R10298 gnd.n7567 gnd.n353 19.3944
R10299 gnd.n7580 gnd.n353 19.3944
R10300 gnd.n7581 gnd.n7580 19.3944
R10301 gnd.n7583 gnd.n7581 19.3944
R10302 gnd.n7584 gnd.n7583 19.3944
R10303 gnd.n7587 gnd.n7584 19.3944
R10304 gnd.n7588 gnd.n7587 19.3944
R10305 gnd.n7590 gnd.n7588 19.3944
R10306 gnd.n7591 gnd.n7590 19.3944
R10307 gnd.n7594 gnd.n7591 19.3944
R10308 gnd.n7595 gnd.n7594 19.3944
R10309 gnd.n7597 gnd.n7595 19.3944
R10310 gnd.n7598 gnd.n7597 19.3944
R10311 gnd.n7601 gnd.n7598 19.3944
R10312 gnd.n7602 gnd.n7601 19.3944
R10313 gnd.n7604 gnd.n7602 19.3944
R10314 gnd.n7605 gnd.n7604 19.3944
R10315 gnd.n7608 gnd.n7605 19.3944
R10316 gnd.n7609 gnd.n7608 19.3944
R10317 gnd.n7743 gnd.n7609 19.3944
R10318 gnd.n7744 gnd.n7743 19.3944
R10319 gnd.n7747 gnd.n7744 19.3944
R10320 gnd.n7748 gnd.n7747 19.3944
R10321 gnd.n7750 gnd.n7748 19.3944
R10322 gnd.n7751 gnd.n7750 19.3944
R10323 gnd.n7754 gnd.n7751 19.3944
R10324 gnd.n7755 gnd.n7754 19.3944
R10325 gnd.n7757 gnd.n7755 19.3944
R10326 gnd.n7758 gnd.n7757 19.3944
R10327 gnd.n7761 gnd.n7758 19.3944
R10328 gnd.n7308 gnd.n7307 19.3944
R10329 gnd.n7307 gnd.n558 19.3944
R10330 gnd.n561 gnd.n558 19.3944
R10331 gnd.n561 gnd.n528 19.3944
R10332 gnd.n7350 gnd.n528 19.3944
R10333 gnd.n7350 gnd.n7349 19.3944
R10334 gnd.n7349 gnd.n7348 19.3944
R10335 gnd.n7348 gnd.n7347 19.3944
R10336 gnd.n7347 gnd.n492 19.3944
R10337 gnd.n7399 gnd.n492 19.3944
R10338 gnd.n7399 gnd.n7398 19.3944
R10339 gnd.n7398 gnd.n7397 19.3944
R10340 gnd.n7397 gnd.n7396 19.3944
R10341 gnd.n7396 gnd.n462 19.3944
R10342 gnd.n7436 gnd.n462 19.3944
R10343 gnd.n7436 gnd.n7435 19.3944
R10344 gnd.n7435 gnd.n7434 19.3944
R10345 gnd.n7434 gnd.n7433 19.3944
R10346 gnd.n7433 gnd.n426 19.3944
R10347 gnd.n7484 gnd.n426 19.3944
R10348 gnd.n7484 gnd.n7483 19.3944
R10349 gnd.n7483 gnd.n7482 19.3944
R10350 gnd.n7482 gnd.n7481 19.3944
R10351 gnd.n7481 gnd.n388 19.3944
R10352 gnd.n7534 gnd.n388 19.3944
R10353 gnd.n7534 gnd.n7533 19.3944
R10354 gnd.n7533 gnd.n7532 19.3944
R10355 gnd.n7532 gnd.n7530 19.3944
R10356 gnd.n7530 gnd.n7529 19.3944
R10357 gnd.n7529 gnd.n362 19.3944
R10358 gnd.n7563 gnd.n362 19.3944
R10359 gnd.n7563 gnd.n355 19.3944
R10360 gnd.n7572 gnd.n355 19.3944
R10361 gnd.n7573 gnd.n7572 19.3944
R10362 gnd.n7575 gnd.n7573 19.3944
R10363 gnd.n7575 gnd.n127 19.3944
R10364 gnd.n7967 gnd.n127 19.3944
R10365 gnd.n7967 gnd.n7966 19.3944
R10366 gnd.n7966 gnd.n7965 19.3944
R10367 gnd.n7965 gnd.n131 19.3944
R10368 gnd.n7955 gnd.n131 19.3944
R10369 gnd.n7955 gnd.n7954 19.3944
R10370 gnd.n7954 gnd.n7953 19.3944
R10371 gnd.n7953 gnd.n148 19.3944
R10372 gnd.n7943 gnd.n148 19.3944
R10373 gnd.n7943 gnd.n7942 19.3944
R10374 gnd.n7942 gnd.n7941 19.3944
R10375 gnd.n7941 gnd.n168 19.3944
R10376 gnd.n7931 gnd.n168 19.3944
R10377 gnd.n7931 gnd.n7930 19.3944
R10378 gnd.n7930 gnd.n7929 19.3944
R10379 gnd.n7929 gnd.n186 19.3944
R10380 gnd.n7919 gnd.n186 19.3944
R10381 gnd.n7919 gnd.n7918 19.3944
R10382 gnd.n7918 gnd.n7917 19.3944
R10383 gnd.n7917 gnd.n206 19.3944
R10384 gnd.n7907 gnd.n206 19.3944
R10385 gnd.n7907 gnd.n7906 19.3944
R10386 gnd.n7906 gnd.n7905 19.3944
R10387 gnd.n7905 gnd.n224 19.3944
R10388 gnd.n7895 gnd.n224 19.3944
R10389 gnd.n7895 gnd.n7894 19.3944
R10390 gnd.n7894 gnd.n7893 19.3944
R10391 gnd.n7893 gnd.n244 19.3944
R10392 gnd.n7804 gnd.n329 19.3944
R10393 gnd.n7804 gnd.n7801 19.3944
R10394 gnd.n7801 gnd.n7798 19.3944
R10395 gnd.n7798 gnd.n7797 19.3944
R10396 gnd.n7797 gnd.n7794 19.3944
R10397 gnd.n7794 gnd.n7793 19.3944
R10398 gnd.n7793 gnd.n7790 19.3944
R10399 gnd.n7790 gnd.n7789 19.3944
R10400 gnd.n7789 gnd.n7786 19.3944
R10401 gnd.n7786 gnd.n7785 19.3944
R10402 gnd.n7785 gnd.n7782 19.3944
R10403 gnd.n7782 gnd.n7781 19.3944
R10404 gnd.n7781 gnd.n7778 19.3944
R10405 gnd.n7778 gnd.n7777 19.3944
R10406 gnd.n7777 gnd.n7774 19.3944
R10407 gnd.n7774 gnd.n7773 19.3944
R10408 gnd.n7773 gnd.n7770 19.3944
R10409 gnd.n7770 gnd.n7769 19.3944
R10410 gnd.n7847 gnd.n7844 19.3944
R10411 gnd.n7844 gnd.n7843 19.3944
R10412 gnd.n7843 gnd.n7840 19.3944
R10413 gnd.n7840 gnd.n7839 19.3944
R10414 gnd.n7839 gnd.n7836 19.3944
R10415 gnd.n7836 gnd.n7835 19.3944
R10416 gnd.n7835 gnd.n7832 19.3944
R10417 gnd.n7832 gnd.n7831 19.3944
R10418 gnd.n7831 gnd.n7828 19.3944
R10419 gnd.n7828 gnd.n7827 19.3944
R10420 gnd.n7827 gnd.n7824 19.3944
R10421 gnd.n7824 gnd.n7823 19.3944
R10422 gnd.n7823 gnd.n7820 19.3944
R10423 gnd.n7820 gnd.n7819 19.3944
R10424 gnd.n7819 gnd.n7816 19.3944
R10425 gnd.n7816 gnd.n7815 19.3944
R10426 gnd.n7815 gnd.n7812 19.3944
R10427 gnd.n7812 gnd.n7811 19.3944
R10428 gnd.n7885 gnd.n253 19.3944
R10429 gnd.n7880 gnd.n253 19.3944
R10430 gnd.n7880 gnd.n7879 19.3944
R10431 gnd.n7879 gnd.n7878 19.3944
R10432 gnd.n7878 gnd.n7875 19.3944
R10433 gnd.n7875 gnd.n7874 19.3944
R10434 gnd.n7874 gnd.n7871 19.3944
R10435 gnd.n7871 gnd.n7870 19.3944
R10436 gnd.n7870 gnd.n7867 19.3944
R10437 gnd.n7867 gnd.n7866 19.3944
R10438 gnd.n7866 gnd.n7863 19.3944
R10439 gnd.n7863 gnd.n7862 19.3944
R10440 gnd.n7862 gnd.n7859 19.3944
R10441 gnd.n7859 gnd.n7858 19.3944
R10442 gnd.n7858 gnd.n7855 19.3944
R10443 gnd.n7855 gnd.n7854 19.3944
R10444 gnd.n7854 gnd.n7851 19.3944
R10445 gnd.n7679 gnd.n7677 19.3944
R10446 gnd.n7682 gnd.n7679 19.3944
R10447 gnd.n7685 gnd.n7682 19.3944
R10448 gnd.n7688 gnd.n7685 19.3944
R10449 gnd.n7688 gnd.n7675 19.3944
R10450 gnd.n7692 gnd.n7675 19.3944
R10451 gnd.n7695 gnd.n7692 19.3944
R10452 gnd.n7698 gnd.n7695 19.3944
R10453 gnd.n7698 gnd.n7673 19.3944
R10454 gnd.n7702 gnd.n7673 19.3944
R10455 gnd.n7705 gnd.n7702 19.3944
R10456 gnd.n7708 gnd.n7705 19.3944
R10457 gnd.n7708 gnd.n7671 19.3944
R10458 gnd.n7712 gnd.n7671 19.3944
R10459 gnd.n7715 gnd.n7712 19.3944
R10460 gnd.n7718 gnd.n7715 19.3944
R10461 gnd.n7099 gnd.n541 19.3944
R10462 gnd.n7322 gnd.n541 19.3944
R10463 gnd.n7322 gnd.n538 19.3944
R10464 gnd.n7327 gnd.n538 19.3944
R10465 gnd.n7327 gnd.n539 19.3944
R10466 gnd.n539 gnd.n510 19.3944
R10467 gnd.n7364 gnd.n510 19.3944
R10468 gnd.n7364 gnd.n507 19.3944
R10469 gnd.n7369 gnd.n507 19.3944
R10470 gnd.n7369 gnd.n508 19.3944
R10471 gnd.n508 gnd.n475 19.3944
R10472 gnd.n7413 gnd.n475 19.3944
R10473 gnd.n7413 gnd.n472 19.3944
R10474 gnd.n7418 gnd.n472 19.3944
R10475 gnd.n7418 gnd.n473 19.3944
R10476 gnd.n473 gnd.n444 19.3944
R10477 gnd.n7450 gnd.n444 19.3944
R10478 gnd.n7450 gnd.n441 19.3944
R10479 gnd.n7455 gnd.n441 19.3944
R10480 gnd.n7455 gnd.n442 19.3944
R10481 gnd.n442 gnd.n409 19.3944
R10482 gnd.n7499 gnd.n409 19.3944
R10483 gnd.n7499 gnd.n406 19.3944
R10484 gnd.n7506 gnd.n406 19.3944
R10485 gnd.n7506 gnd.n407 19.3944
R10486 gnd.n7502 gnd.n407 19.3944
R10487 gnd.n7502 gnd.n374 19.3944
R10488 gnd.n7547 gnd.n374 19.3944
R10489 gnd.n7547 gnd.n371 19.3944
R10490 gnd.n7551 gnd.n371 19.3944
R10491 gnd.n7551 gnd.n372 19.3944
R10492 gnd.n372 gnd.n100 19.3944
R10493 gnd.n7980 gnd.n100 19.3944
R10494 gnd.n7980 gnd.n7979 19.3944
R10495 gnd.n7979 gnd.n103 19.3944
R10496 gnd.n7621 gnd.n103 19.3944
R10497 gnd.n7621 gnd.n7618 19.3944
R10498 gnd.n7626 gnd.n7618 19.3944
R10499 gnd.n7627 gnd.n7626 19.3944
R10500 gnd.n7629 gnd.n7627 19.3944
R10501 gnd.n7629 gnd.n7616 19.3944
R10502 gnd.n7634 gnd.n7616 19.3944
R10503 gnd.n7635 gnd.n7634 19.3944
R10504 gnd.n7637 gnd.n7635 19.3944
R10505 gnd.n7637 gnd.n7614 19.3944
R10506 gnd.n7642 gnd.n7614 19.3944
R10507 gnd.n7643 gnd.n7642 19.3944
R10508 gnd.n7645 gnd.n7643 19.3944
R10509 gnd.n7645 gnd.n7612 19.3944
R10510 gnd.n7650 gnd.n7612 19.3944
R10511 gnd.n7651 gnd.n7650 19.3944
R10512 gnd.n7653 gnd.n7651 19.3944
R10513 gnd.n7653 gnd.n7610 19.3944
R10514 gnd.n7739 gnd.n7610 19.3944
R10515 gnd.n7739 gnd.n7738 19.3944
R10516 gnd.n7738 gnd.n7737 19.3944
R10517 gnd.n7737 gnd.n7735 19.3944
R10518 gnd.n7735 gnd.n7734 19.3944
R10519 gnd.n7734 gnd.n7732 19.3944
R10520 gnd.n7732 gnd.n7731 19.3944
R10521 gnd.n7731 gnd.n7729 19.3944
R10522 gnd.n7729 gnd.n7728 19.3944
R10523 gnd.n7728 gnd.n7726 19.3944
R10524 gnd.n7726 gnd.n7725 19.3944
R10525 gnd.n7312 gnd.n548 19.3944
R10526 gnd.n7318 gnd.n548 19.3944
R10527 gnd.n7318 gnd.n7317 19.3944
R10528 gnd.n7317 gnd.n520 19.3944
R10529 gnd.n7354 gnd.n520 19.3944
R10530 gnd.n7354 gnd.n518 19.3944
R10531 gnd.n7360 gnd.n518 19.3944
R10532 gnd.n7360 gnd.n7359 19.3944
R10533 gnd.n7359 gnd.n484 19.3944
R10534 gnd.n7403 gnd.n484 19.3944
R10535 gnd.n7403 gnd.n482 19.3944
R10536 gnd.n7409 gnd.n482 19.3944
R10537 gnd.n7409 gnd.n7408 19.3944
R10538 gnd.n7408 gnd.n454 19.3944
R10539 gnd.n7440 gnd.n454 19.3944
R10540 gnd.n7440 gnd.n452 19.3944
R10541 gnd.n7446 gnd.n452 19.3944
R10542 gnd.n7446 gnd.n7445 19.3944
R10543 gnd.n7445 gnd.n419 19.3944
R10544 gnd.n7488 gnd.n419 19.3944
R10545 gnd.n7488 gnd.n417 19.3944
R10546 gnd.n7495 gnd.n417 19.3944
R10547 gnd.n7495 gnd.n7494 19.3944
R10548 gnd.n7494 gnd.n380 19.3944
R10549 gnd.n7538 gnd.n380 19.3944
R10550 gnd.n7539 gnd.n7538 19.3944
R10551 gnd.n7540 gnd.n7539 19.3944
R10552 gnd.n7543 gnd.n7542 19.3944
R10553 gnd.n7559 gnd.n7558 19.3944
R10554 gnd.n7556 gnd.n7555 19.3944
R10555 gnd.n7975 gnd.n7974 19.3944
R10556 gnd.n7971 gnd.n111 19.3944
R10557 gnd.n7971 gnd.n118 19.3944
R10558 gnd.n7961 gnd.n118 19.3944
R10559 gnd.n7961 gnd.n7960 19.3944
R10560 gnd.n7960 gnd.n7959 19.3944
R10561 gnd.n7959 gnd.n140 19.3944
R10562 gnd.n7949 gnd.n140 19.3944
R10563 gnd.n7949 gnd.n7948 19.3944
R10564 gnd.n7948 gnd.n7947 19.3944
R10565 gnd.n7947 gnd.n158 19.3944
R10566 gnd.n7937 gnd.n158 19.3944
R10567 gnd.n7937 gnd.n7936 19.3944
R10568 gnd.n7936 gnd.n7935 19.3944
R10569 gnd.n7935 gnd.n178 19.3944
R10570 gnd.n7925 gnd.n178 19.3944
R10571 gnd.n7925 gnd.n7924 19.3944
R10572 gnd.n7924 gnd.n7923 19.3944
R10573 gnd.n7923 gnd.n196 19.3944
R10574 gnd.n7913 gnd.n196 19.3944
R10575 gnd.n7913 gnd.n7912 19.3944
R10576 gnd.n7912 gnd.n7911 19.3944
R10577 gnd.n7911 gnd.n216 19.3944
R10578 gnd.n7901 gnd.n216 19.3944
R10579 gnd.n7901 gnd.n7900 19.3944
R10580 gnd.n7900 gnd.n7899 19.3944
R10581 gnd.n7899 gnd.n235 19.3944
R10582 gnd.n7889 gnd.n235 19.3944
R10583 gnd.n7889 gnd.n7888 19.3944
R10584 gnd.n3830 gnd.n3829 19.3944
R10585 gnd.n3829 gnd.n3828 19.3944
R10586 gnd.n3828 gnd.n3827 19.3944
R10587 gnd.n3827 gnd.n3825 19.3944
R10588 gnd.n3825 gnd.n3822 19.3944
R10589 gnd.n3822 gnd.n3821 19.3944
R10590 gnd.n3821 gnd.n3818 19.3944
R10591 gnd.n3818 gnd.n3817 19.3944
R10592 gnd.n3817 gnd.n3814 19.3944
R10593 gnd.n3814 gnd.n3813 19.3944
R10594 gnd.n3813 gnd.n3810 19.3944
R10595 gnd.n3810 gnd.n3809 19.3944
R10596 gnd.n3809 gnd.n3806 19.3944
R10597 gnd.n3806 gnd.n3805 19.3944
R10598 gnd.n3805 gnd.n3802 19.3944
R10599 gnd.n3802 gnd.n3801 19.3944
R10600 gnd.n3801 gnd.n3798 19.3944
R10601 gnd.n3796 gnd.n3793 19.3944
R10602 gnd.n3793 gnd.n3792 19.3944
R10603 gnd.n3792 gnd.n3789 19.3944
R10604 gnd.n3789 gnd.n3788 19.3944
R10605 gnd.n3788 gnd.n3785 19.3944
R10606 gnd.n3785 gnd.n3784 19.3944
R10607 gnd.n3784 gnd.n3781 19.3944
R10608 gnd.n3781 gnd.n3780 19.3944
R10609 gnd.n3780 gnd.n3777 19.3944
R10610 gnd.n3777 gnd.n3776 19.3944
R10611 gnd.n3776 gnd.n3773 19.3944
R10612 gnd.n3773 gnd.n3772 19.3944
R10613 gnd.n3772 gnd.n3769 19.3944
R10614 gnd.n3769 gnd.n3768 19.3944
R10615 gnd.n3768 gnd.n3765 19.3944
R10616 gnd.n3765 gnd.n3764 19.3944
R10617 gnd.n3764 gnd.n3761 19.3944
R10618 gnd.n3761 gnd.n3760 19.3944
R10619 gnd.n3756 gnd.n3753 19.3944
R10620 gnd.n3753 gnd.n3752 19.3944
R10621 gnd.n3752 gnd.n3749 19.3944
R10622 gnd.n3749 gnd.n3748 19.3944
R10623 gnd.n3748 gnd.n3745 19.3944
R10624 gnd.n3745 gnd.n3744 19.3944
R10625 gnd.n3744 gnd.n3741 19.3944
R10626 gnd.n3741 gnd.n3740 19.3944
R10627 gnd.n3740 gnd.n3737 19.3944
R10628 gnd.n3737 gnd.n3736 19.3944
R10629 gnd.n3736 gnd.n3733 19.3944
R10630 gnd.n3733 gnd.n3732 19.3944
R10631 gnd.n3732 gnd.n3729 19.3944
R10632 gnd.n3729 gnd.n3728 19.3944
R10633 gnd.n3728 gnd.n3725 19.3944
R10634 gnd.n3725 gnd.n3724 19.3944
R10635 gnd.n3724 gnd.n3721 19.3944
R10636 gnd.n3721 gnd.n3720 19.3944
R10637 gnd.n3432 gnd.n3431 19.3944
R10638 gnd.n3435 gnd.n3432 19.3944
R10639 gnd.n3435 gnd.n3427 19.3944
R10640 gnd.n3441 gnd.n3427 19.3944
R10641 gnd.n3442 gnd.n3441 19.3944
R10642 gnd.n3445 gnd.n3442 19.3944
R10643 gnd.n3445 gnd.n3425 19.3944
R10644 gnd.n3451 gnd.n3425 19.3944
R10645 gnd.n3452 gnd.n3451 19.3944
R10646 gnd.n3455 gnd.n3452 19.3944
R10647 gnd.n3455 gnd.n3423 19.3944
R10648 gnd.n3461 gnd.n3423 19.3944
R10649 gnd.n3462 gnd.n3461 19.3944
R10650 gnd.n3465 gnd.n3462 19.3944
R10651 gnd.n3465 gnd.n3419 19.3944
R10652 gnd.n3469 gnd.n3419 19.3944
R10653 gnd.n3476 gnd.n3475 19.3944
R10654 gnd.n3478 gnd.n3476 19.3944
R10655 gnd.n3478 gnd.n3413 19.3944
R10656 gnd.n3483 gnd.n3413 19.3944
R10657 gnd.n3484 gnd.n3483 19.3944
R10658 gnd.n3486 gnd.n3484 19.3944
R10659 gnd.n3486 gnd.n3411 19.3944
R10660 gnd.n3491 gnd.n3411 19.3944
R10661 gnd.n3492 gnd.n3491 19.3944
R10662 gnd.n3494 gnd.n3492 19.3944
R10663 gnd.n3494 gnd.n3409 19.3944
R10664 gnd.n3499 gnd.n3409 19.3944
R10665 gnd.n3500 gnd.n3499 19.3944
R10666 gnd.n3502 gnd.n3500 19.3944
R10667 gnd.n3502 gnd.n3407 19.3944
R10668 gnd.n3507 gnd.n3407 19.3944
R10669 gnd.n3508 gnd.n3507 19.3944
R10670 gnd.n3510 gnd.n3508 19.3944
R10671 gnd.n3510 gnd.n3405 19.3944
R10672 gnd.n3515 gnd.n3405 19.3944
R10673 gnd.n3516 gnd.n3515 19.3944
R10674 gnd.n3518 gnd.n3516 19.3944
R10675 gnd.n3518 gnd.n3403 19.3944
R10676 gnd.n3523 gnd.n3403 19.3944
R10677 gnd.n3524 gnd.n3523 19.3944
R10678 gnd.n3525 gnd.n3524 19.3944
R10679 gnd.n3525 gnd.n3401 19.3944
R10680 gnd.n3546 gnd.n3401 19.3944
R10681 gnd.n3546 gnd.n3545 19.3944
R10682 gnd.n3545 gnd.n3544 19.3944
R10683 gnd.n3544 gnd.n3542 19.3944
R10684 gnd.n3542 gnd.n3541 19.3944
R10685 gnd.n3541 gnd.n3533 19.3944
R10686 gnd.n3537 gnd.n3533 19.3944
R10687 gnd.n3537 gnd.n3536 19.3944
R10688 gnd.n3536 gnd.n1764 19.3944
R10689 gnd.n5359 gnd.n1764 19.3944
R10690 gnd.n5359 gnd.n1761 19.3944
R10691 gnd.n5364 gnd.n1761 19.3944
R10692 gnd.n5364 gnd.n1762 19.3944
R10693 gnd.n1762 gnd.n1729 19.3944
R10694 gnd.n5404 gnd.n1729 19.3944
R10695 gnd.n5404 gnd.n1726 19.3944
R10696 gnd.n5409 gnd.n1726 19.3944
R10697 gnd.n5409 gnd.n1727 19.3944
R10698 gnd.n1727 gnd.n1690 19.3944
R10699 gnd.n5454 gnd.n1690 19.3944
R10700 gnd.n5454 gnd.n1687 19.3944
R10701 gnd.n5458 gnd.n1687 19.3944
R10702 gnd.n5459 gnd.n5458 19.3944
R10703 gnd.n5461 gnd.n5459 19.3944
R10704 gnd.n5461 gnd.n1684 19.3944
R10705 gnd.n5466 gnd.n1684 19.3944
R10706 gnd.n5466 gnd.n1685 19.3944
R10707 gnd.n1685 gnd.n1625 19.3944
R10708 gnd.n5557 gnd.n1625 19.3944
R10709 gnd.n5557 gnd.n1622 19.3944
R10710 gnd.n5575 gnd.n1622 19.3944
R10711 gnd.n5575 gnd.n1623 19.3944
R10712 gnd.n5571 gnd.n1623 19.3944
R10713 gnd.n5571 gnd.n5570 19.3944
R10714 gnd.n5570 gnd.n5569 19.3944
R10715 gnd.n5569 gnd.n5565 19.3944
R10716 gnd.n5565 gnd.n1242 19.3944
R10717 gnd.n3712 gnd.n3273 19.3944
R10718 gnd.n3552 gnd.n3273 19.3944
R10719 gnd.n3553 gnd.n3552 19.3944
R10720 gnd.n3555 gnd.n3553 19.3944
R10721 gnd.n3556 gnd.n3555 19.3944
R10722 gnd.n3559 gnd.n3556 19.3944
R10723 gnd.n3560 gnd.n3559 19.3944
R10724 gnd.n3562 gnd.n3560 19.3944
R10725 gnd.n3563 gnd.n3562 19.3944
R10726 gnd.n3566 gnd.n3563 19.3944
R10727 gnd.n3567 gnd.n3566 19.3944
R10728 gnd.n3569 gnd.n3567 19.3944
R10729 gnd.n3570 gnd.n3569 19.3944
R10730 gnd.n3573 gnd.n3570 19.3944
R10731 gnd.n3574 gnd.n3573 19.3944
R10732 gnd.n3576 gnd.n3574 19.3944
R10733 gnd.n3577 gnd.n3576 19.3944
R10734 gnd.n3580 gnd.n3577 19.3944
R10735 gnd.n3581 gnd.n3580 19.3944
R10736 gnd.n3583 gnd.n3581 19.3944
R10737 gnd.n3584 gnd.n3583 19.3944
R10738 gnd.n3587 gnd.n3584 19.3944
R10739 gnd.n3588 gnd.n3587 19.3944
R10740 gnd.n3590 gnd.n3588 19.3944
R10741 gnd.n3591 gnd.n3590 19.3944
R10742 gnd.n3592 gnd.n3591 19.3944
R10743 gnd.n3625 gnd.n3592 19.3944
R10744 gnd.n3625 gnd.n3624 19.3944
R10745 gnd.n3624 gnd.n3622 19.3944
R10746 gnd.n3622 gnd.n3621 19.3944
R10747 gnd.n3621 gnd.n3619 19.3944
R10748 gnd.n3619 gnd.n3618 19.3944
R10749 gnd.n3618 gnd.n3616 19.3944
R10750 gnd.n3616 gnd.n3615 19.3944
R10751 gnd.n3615 gnd.n3613 19.3944
R10752 gnd.n3613 gnd.n3612 19.3944
R10753 gnd.n3612 gnd.n3610 19.3944
R10754 gnd.n3610 gnd.n1757 19.3944
R10755 gnd.n5368 gnd.n1757 19.3944
R10756 gnd.n5369 gnd.n5368 19.3944
R10757 gnd.n5371 gnd.n5369 19.3944
R10758 gnd.n5371 gnd.n5370 19.3944
R10759 gnd.n5370 gnd.n1722 19.3944
R10760 gnd.n5413 gnd.n1722 19.3944
R10761 gnd.n5414 gnd.n5413 19.3944
R10762 gnd.n5421 gnd.n5414 19.3944
R10763 gnd.n5421 gnd.n5420 19.3944
R10764 gnd.n5420 gnd.n5419 19.3944
R10765 gnd.n5419 gnd.n5418 19.3944
R10766 gnd.n5418 gnd.n5416 19.3944
R10767 gnd.n5416 gnd.n1678 19.3944
R10768 gnd.n5471 gnd.n1678 19.3944
R10769 gnd.n5471 gnd.n5470 19.3944
R10770 gnd.n5470 gnd.n1683 19.3944
R10771 gnd.n1683 gnd.n1682 19.3944
R10772 gnd.n1682 gnd.n1679 19.3944
R10773 gnd.n1679 gnd.n1619 19.3944
R10774 gnd.n5579 gnd.n1619 19.3944
R10775 gnd.n5580 gnd.n5579 19.3944
R10776 gnd.n5580 gnd.n1599 19.3944
R10777 gnd.n5597 gnd.n1599 19.3944
R10778 gnd.n5597 gnd.n1593 19.3944
R10779 gnd.n5605 gnd.n1593 19.3944
R10780 gnd.n5606 gnd.n5605 19.3944
R10781 gnd.n3292 gnd.n3271 19.3944
R10782 gnd.n3293 gnd.n3292 19.3944
R10783 gnd.n3701 gnd.n3293 19.3944
R10784 gnd.n3701 gnd.n3700 19.3944
R10785 gnd.n3700 gnd.n3699 19.3944
R10786 gnd.n3699 gnd.n3297 19.3944
R10787 gnd.n3689 gnd.n3297 19.3944
R10788 gnd.n3689 gnd.n3688 19.3944
R10789 gnd.n3688 gnd.n3687 19.3944
R10790 gnd.n3687 gnd.n3316 19.3944
R10791 gnd.n3677 gnd.n3316 19.3944
R10792 gnd.n3677 gnd.n3676 19.3944
R10793 gnd.n3676 gnd.n3675 19.3944
R10794 gnd.n3675 gnd.n3335 19.3944
R10795 gnd.n3665 gnd.n3335 19.3944
R10796 gnd.n3665 gnd.n3664 19.3944
R10797 gnd.n3664 gnd.n3663 19.3944
R10798 gnd.n3663 gnd.n3354 19.3944
R10799 gnd.n3653 gnd.n3354 19.3944
R10800 gnd.n3653 gnd.n3652 19.3944
R10801 gnd.n3652 gnd.n3651 19.3944
R10802 gnd.n3651 gnd.n3373 19.3944
R10803 gnd.n3641 gnd.n3373 19.3944
R10804 gnd.n3641 gnd.n3640 19.3944
R10805 gnd.n3640 gnd.n3639 19.3944
R10806 gnd.n3639 gnd.n3392 19.3944
R10807 gnd.n3627 gnd.n3392 19.3944
R10808 gnd.n3627 gnd.n1787 19.3944
R10809 gnd.n5345 gnd.n1787 19.3944
R10810 gnd.n5345 gnd.n5344 19.3944
R10811 gnd.n5344 gnd.n5343 19.3944
R10812 gnd.n5343 gnd.n1791 19.3944
R10813 gnd.n5331 gnd.n1791 19.3944
R10814 gnd.n5331 gnd.n5330 19.3944
R10815 gnd.n5330 gnd.n5329 19.3944
R10816 gnd.n5329 gnd.n1803 19.3944
R10817 gnd.n3595 gnd.n1803 19.3944
R10818 gnd.n3607 gnd.n3595 19.3944
R10819 gnd.n3607 gnd.n1746 19.3944
R10820 gnd.n5390 gnd.n1746 19.3944
R10821 gnd.n5390 gnd.n5389 19.3944
R10822 gnd.n5389 gnd.n5388 19.3944
R10823 gnd.n5388 gnd.n5387 19.3944
R10824 gnd.n5387 gnd.n1708 19.3944
R10825 gnd.n5440 gnd.n1708 19.3944
R10826 gnd.n5440 gnd.n5439 19.3944
R10827 gnd.n5439 gnd.n5438 19.3944
R10828 gnd.n5438 gnd.n5437 19.3944
R10829 gnd.n5437 gnd.n1673 19.3944
R10830 gnd.n5475 gnd.n1673 19.3944
R10831 gnd.n5475 gnd.n5474 19.3944
R10832 gnd.n5474 gnd.n5473 19.3944
R10833 gnd.n5473 gnd.n1643 19.3944
R10834 gnd.n5543 gnd.n1643 19.3944
R10835 gnd.n5543 gnd.n5542 19.3944
R10836 gnd.n5542 gnd.n5541 19.3944
R10837 gnd.n5541 gnd.n5540 19.3944
R10838 gnd.n5540 gnd.n1617 19.3944
R10839 gnd.n5583 gnd.n1617 19.3944
R10840 gnd.n5583 gnd.n5582 19.3944
R10841 gnd.n5582 gnd.n1597 19.3944
R10842 gnd.n5600 gnd.n1597 19.3944
R10843 gnd.n5601 gnd.n5600 19.3944
R10844 gnd.n5601 gnd.n1592 19.3944
R10845 gnd.n6147 gnd.n6146 19.3944
R10846 gnd.n6146 gnd.n1252 19.3944
R10847 gnd.n1254 gnd.n1252 19.3944
R10848 gnd.n6139 gnd.n1254 19.3944
R10849 gnd.n6139 gnd.n6138 19.3944
R10850 gnd.n6138 gnd.n6137 19.3944
R10851 gnd.n6137 gnd.n1261 19.3944
R10852 gnd.n6132 gnd.n1261 19.3944
R10853 gnd.n6132 gnd.n6131 19.3944
R10854 gnd.n6131 gnd.n6130 19.3944
R10855 gnd.n6130 gnd.n1268 19.3944
R10856 gnd.n6125 gnd.n1268 19.3944
R10857 gnd.n6125 gnd.n6124 19.3944
R10858 gnd.n6124 gnd.n6123 19.3944
R10859 gnd.n6123 gnd.n1275 19.3944
R10860 gnd.n6118 gnd.n1275 19.3944
R10861 gnd.n6118 gnd.n6117 19.3944
R10862 gnd.n1540 gnd.n1500 19.3944
R10863 gnd.n1544 gnd.n1500 19.3944
R10864 gnd.n1544 gnd.n1498 19.3944
R10865 gnd.n1550 gnd.n1498 19.3944
R10866 gnd.n1550 gnd.n1496 19.3944
R10867 gnd.n1554 gnd.n1496 19.3944
R10868 gnd.n1554 gnd.n1494 19.3944
R10869 gnd.n1560 gnd.n1494 19.3944
R10870 gnd.n1560 gnd.n1492 19.3944
R10871 gnd.n1564 gnd.n1492 19.3944
R10872 gnd.n1564 gnd.n1490 19.3944
R10873 gnd.n1570 gnd.n1490 19.3944
R10874 gnd.n1570 gnd.n1488 19.3944
R10875 gnd.n1574 gnd.n1488 19.3944
R10876 gnd.n1574 gnd.n1486 19.3944
R10877 gnd.n1580 gnd.n1486 19.3944
R10878 gnd.n1580 gnd.n1484 19.3944
R10879 gnd.n1584 gnd.n1484 19.3944
R10880 gnd.n1513 gnd.n1297 19.3944
R10881 gnd.n1520 gnd.n1513 19.3944
R10882 gnd.n1520 gnd.n1510 19.3944
R10883 gnd.n1524 gnd.n1510 19.3944
R10884 gnd.n1524 gnd.n1508 19.3944
R10885 gnd.n1530 gnd.n1508 19.3944
R10886 gnd.n1530 gnd.n1506 19.3944
R10887 gnd.n1534 gnd.n1506 19.3944
R10888 gnd.n6115 gnd.n1284 19.3944
R10889 gnd.n6110 gnd.n1284 19.3944
R10890 gnd.n6110 gnd.n6109 19.3944
R10891 gnd.n6109 gnd.n6108 19.3944
R10892 gnd.n6108 gnd.n1291 19.3944
R10893 gnd.n6103 gnd.n1291 19.3944
R10894 gnd.n6103 gnd.n6102 19.3944
R10895 gnd.n3707 gnd.n3279 19.3944
R10896 gnd.n3707 gnd.n3706 19.3944
R10897 gnd.n3706 gnd.n3705 19.3944
R10898 gnd.n3705 gnd.n3284 19.3944
R10899 gnd.n3695 gnd.n3284 19.3944
R10900 gnd.n3695 gnd.n3694 19.3944
R10901 gnd.n3694 gnd.n3693 19.3944
R10902 gnd.n3693 gnd.n3307 19.3944
R10903 gnd.n3683 gnd.n3307 19.3944
R10904 gnd.n3683 gnd.n3682 19.3944
R10905 gnd.n3682 gnd.n3681 19.3944
R10906 gnd.n3681 gnd.n3325 19.3944
R10907 gnd.n3671 gnd.n3325 19.3944
R10908 gnd.n3671 gnd.n3670 19.3944
R10909 gnd.n3670 gnd.n3669 19.3944
R10910 gnd.n3669 gnd.n3345 19.3944
R10911 gnd.n3659 gnd.n3345 19.3944
R10912 gnd.n3659 gnd.n3658 19.3944
R10913 gnd.n3658 gnd.n3657 19.3944
R10914 gnd.n3657 gnd.n3363 19.3944
R10915 gnd.n3647 gnd.n3363 19.3944
R10916 gnd.n3647 gnd.n3646 19.3944
R10917 gnd.n3646 gnd.n3645 19.3944
R10918 gnd.n3645 gnd.n3383 19.3944
R10919 gnd.n3635 gnd.n3383 19.3944
R10920 gnd.n3635 gnd.n3634 19.3944
R10921 gnd.n3634 gnd.n1779 19.3944
R10922 gnd.n5350 gnd.n5349 19.3944
R10923 gnd.n5339 gnd.n5338 19.3944
R10924 gnd.n5336 gnd.n5335 19.3944
R10925 gnd.n5325 gnd.n5324 19.3944
R10926 gnd.n5355 gnd.n1772 19.3944
R10927 gnd.n5355 gnd.n5354 19.3944
R10928 gnd.n5354 gnd.n1738 19.3944
R10929 gnd.n5394 gnd.n1738 19.3944
R10930 gnd.n5394 gnd.n1736 19.3944
R10931 gnd.n5400 gnd.n1736 19.3944
R10932 gnd.n5400 gnd.n5399 19.3944
R10933 gnd.n5399 gnd.n1700 19.3944
R10934 gnd.n5444 gnd.n1700 19.3944
R10935 gnd.n5444 gnd.n1698 19.3944
R10936 gnd.n5450 gnd.n1698 19.3944
R10937 gnd.n5450 gnd.n5449 19.3944
R10938 gnd.n5449 gnd.n1666 19.3944
R10939 gnd.n5479 gnd.n1666 19.3944
R10940 gnd.n5479 gnd.n1664 19.3944
R10941 gnd.n5483 gnd.n1664 19.3944
R10942 gnd.n5483 gnd.n1635 19.3944
R10943 gnd.n5547 gnd.n1635 19.3944
R10944 gnd.n5547 gnd.n1633 19.3944
R10945 gnd.n5553 gnd.n1633 19.3944
R10946 gnd.n5553 gnd.n5552 19.3944
R10947 gnd.n5552 gnd.n1609 19.3944
R10948 gnd.n5587 gnd.n1609 19.3944
R10949 gnd.n5587 gnd.n1607 19.3944
R10950 gnd.n5593 gnd.n1607 19.3944
R10951 gnd.n5593 gnd.n5592 19.3944
R10952 gnd.n5592 gnd.n1249 19.3944
R10953 gnd.n6150 gnd.n1249 19.3944
R10954 gnd.n2945 gnd.n1932 19.3944
R10955 gnd.n2951 gnd.n1932 19.3944
R10956 gnd.n2951 gnd.n1930 19.3944
R10957 gnd.n2955 gnd.n1930 19.3944
R10958 gnd.n2955 gnd.n1926 19.3944
R10959 gnd.n2961 gnd.n1926 19.3944
R10960 gnd.n2961 gnd.n1924 19.3944
R10961 gnd.n2965 gnd.n1924 19.3944
R10962 gnd.n2965 gnd.n1920 19.3944
R10963 gnd.n2971 gnd.n1920 19.3944
R10964 gnd.n2971 gnd.n1918 19.3944
R10965 gnd.n2975 gnd.n1918 19.3944
R10966 gnd.n2975 gnd.n1914 19.3944
R10967 gnd.n2981 gnd.n1914 19.3944
R10968 gnd.n2981 gnd.n1912 19.3944
R10969 gnd.n2985 gnd.n1912 19.3944
R10970 gnd.n2985 gnd.n1908 19.3944
R10971 gnd.n2991 gnd.n1908 19.3944
R10972 gnd.n2991 gnd.n1906 19.3944
R10973 gnd.n2995 gnd.n1906 19.3944
R10974 gnd.n2995 gnd.n1902 19.3944
R10975 gnd.n3001 gnd.n1902 19.3944
R10976 gnd.n3001 gnd.n1900 19.3944
R10977 gnd.n3005 gnd.n1900 19.3944
R10978 gnd.n3005 gnd.n1896 19.3944
R10979 gnd.n3011 gnd.n1896 19.3944
R10980 gnd.n3011 gnd.n1894 19.3944
R10981 gnd.n3015 gnd.n1894 19.3944
R10982 gnd.n3015 gnd.n1890 19.3944
R10983 gnd.n3021 gnd.n1890 19.3944
R10984 gnd.n3021 gnd.n1888 19.3944
R10985 gnd.n3025 gnd.n1888 19.3944
R10986 gnd.n3025 gnd.n1884 19.3944
R10987 gnd.n3031 gnd.n1884 19.3944
R10988 gnd.n3031 gnd.n1882 19.3944
R10989 gnd.n3035 gnd.n1882 19.3944
R10990 gnd.n3035 gnd.n1878 19.3944
R10991 gnd.n3041 gnd.n1878 19.3944
R10992 gnd.n3041 gnd.n1876 19.3944
R10993 gnd.n3045 gnd.n1876 19.3944
R10994 gnd.n3045 gnd.n1872 19.3944
R10995 gnd.n3051 gnd.n1872 19.3944
R10996 gnd.n3051 gnd.n1870 19.3944
R10997 gnd.n3055 gnd.n1870 19.3944
R10998 gnd.n3055 gnd.n1866 19.3944
R10999 gnd.n3061 gnd.n1866 19.3944
R11000 gnd.n3061 gnd.n1864 19.3944
R11001 gnd.n3065 gnd.n1864 19.3944
R11002 gnd.n3065 gnd.n1860 19.3944
R11003 gnd.n3071 gnd.n1860 19.3944
R11004 gnd.n3071 gnd.n1858 19.3944
R11005 gnd.n3075 gnd.n1858 19.3944
R11006 gnd.n3075 gnd.n1854 19.3944
R11007 gnd.n3081 gnd.n1854 19.3944
R11008 gnd.n3081 gnd.n1852 19.3944
R11009 gnd.n3085 gnd.n1852 19.3944
R11010 gnd.n3085 gnd.n1848 19.3944
R11011 gnd.n3091 gnd.n1848 19.3944
R11012 gnd.n3091 gnd.n1846 19.3944
R11013 gnd.n3095 gnd.n1846 19.3944
R11014 gnd.n3095 gnd.n1842 19.3944
R11015 gnd.n3101 gnd.n1842 19.3944
R11016 gnd.n3101 gnd.n1840 19.3944
R11017 gnd.n3105 gnd.n1840 19.3944
R11018 gnd.n3105 gnd.n1836 19.3944
R11019 gnd.n3111 gnd.n1836 19.3944
R11020 gnd.n3111 gnd.n1834 19.3944
R11021 gnd.n3115 gnd.n1834 19.3944
R11022 gnd.n3115 gnd.n1830 19.3944
R11023 gnd.n3121 gnd.n1830 19.3944
R11024 gnd.n3121 gnd.n1828 19.3944
R11025 gnd.n3125 gnd.n1828 19.3944
R11026 gnd.n3125 gnd.n1824 19.3944
R11027 gnd.n3131 gnd.n1824 19.3944
R11028 gnd.n3131 gnd.n1822 19.3944
R11029 gnd.n3135 gnd.n1822 19.3944
R11030 gnd.n3135 gnd.n1818 19.3944
R11031 gnd.n3141 gnd.n1818 19.3944
R11032 gnd.n3141 gnd.n1816 19.3944
R11033 gnd.n3145 gnd.n1816 19.3944
R11034 gnd.n3145 gnd.n1812 19.3944
R11035 gnd.n5317 gnd.n1812 19.3944
R11036 gnd.n5317 gnd.n1810 19.3944
R11037 gnd.n5321 gnd.n1810 19.3944
R11038 gnd.n5745 gnd.n1451 19.3944
R11039 gnd.n5746 gnd.n5745 19.3944
R11040 gnd.n5748 gnd.n5746 19.3944
R11041 gnd.n5748 gnd.n1448 19.3944
R11042 gnd.n5752 gnd.n1448 19.3944
R11043 gnd.n5753 gnd.n5752 19.3944
R11044 gnd.n5755 gnd.n5753 19.3944
R11045 gnd.n5755 gnd.n1445 19.3944
R11046 gnd.n5759 gnd.n1445 19.3944
R11047 gnd.n5760 gnd.n5759 19.3944
R11048 gnd.n5762 gnd.n5760 19.3944
R11049 gnd.n5762 gnd.n1442 19.3944
R11050 gnd.n5766 gnd.n1442 19.3944
R11051 gnd.n5767 gnd.n5766 19.3944
R11052 gnd.n5769 gnd.n5767 19.3944
R11053 gnd.n5769 gnd.n1438 19.3944
R11054 gnd.n5773 gnd.n1438 19.3944
R11055 gnd.n5774 gnd.n5773 19.3944
R11056 gnd.n5776 gnd.n5774 19.3944
R11057 gnd.n5776 gnd.n1435 19.3944
R11058 gnd.n6020 gnd.n1435 19.3944
R11059 gnd.n6020 gnd.n1436 19.3944
R11060 gnd.n6016 gnd.n1436 19.3944
R11061 gnd.n6016 gnd.n6015 19.3944
R11062 gnd.n6015 gnd.n6014 19.3944
R11063 gnd.n6014 gnd.n5782 19.3944
R11064 gnd.n6010 gnd.n5782 19.3944
R11065 gnd.n6010 gnd.n6009 19.3944
R11066 gnd.n6009 gnd.n6008 19.3944
R11067 gnd.n6008 gnd.n5786 19.3944
R11068 gnd.n6004 gnd.n5786 19.3944
R11069 gnd.n6004 gnd.n6003 19.3944
R11070 gnd.n6003 gnd.n6002 19.3944
R11071 gnd.n6002 gnd.n5790 19.3944
R11072 gnd.n5998 gnd.n5790 19.3944
R11073 gnd.n5998 gnd.n5997 19.3944
R11074 gnd.n5997 gnd.n5996 19.3944
R11075 gnd.n5996 gnd.n5794 19.3944
R11076 gnd.n5992 gnd.n5794 19.3944
R11077 gnd.n5992 gnd.n5991 19.3944
R11078 gnd.n5991 gnd.n5990 19.3944
R11079 gnd.n5990 gnd.n5798 19.3944
R11080 gnd.n5986 gnd.n5798 19.3944
R11081 gnd.n5986 gnd.n5985 19.3944
R11082 gnd.n5985 gnd.n5984 19.3944
R11083 gnd.n5984 gnd.n5973 19.3944
R11084 gnd.n5980 gnd.n5973 19.3944
R11085 gnd.n5980 gnd.n5979 19.3944
R11086 gnd.n5979 gnd.n5978 19.3944
R11087 gnd.n5978 gnd.n1021 19.3944
R11088 gnd.n6416 gnd.n1021 19.3944
R11089 gnd.n6416 gnd.n1018 19.3944
R11090 gnd.n6421 gnd.n1018 19.3944
R11091 gnd.n6421 gnd.n1019 19.3944
R11092 gnd.n1019 gnd.n981 19.3944
R11093 gnd.n6474 gnd.n981 19.3944
R11094 gnd.n6474 gnd.n978 19.3944
R11095 gnd.n6478 gnd.n978 19.3944
R11096 gnd.n6479 gnd.n6478 19.3944
R11097 gnd.n6481 gnd.n6479 19.3944
R11098 gnd.n6481 gnd.n976 19.3944
R11099 gnd.n6485 gnd.n976 19.3944
R11100 gnd.n6486 gnd.n6485 19.3944
R11101 gnd.n6488 gnd.n6486 19.3944
R11102 gnd.n6488 gnd.n974 19.3944
R11103 gnd.n6492 gnd.n974 19.3944
R11104 gnd.n6493 gnd.n6492 19.3944
R11105 gnd.n6495 gnd.n6493 19.3944
R11106 gnd.n6495 gnd.n971 19.3944
R11107 gnd.n6855 gnd.n971 19.3944
R11108 gnd.n6855 gnd.n972 19.3944
R11109 gnd.n6851 gnd.n972 19.3944
R11110 gnd.n6851 gnd.n6850 19.3944
R11111 gnd.n6850 gnd.n6849 19.3944
R11112 gnd.n6849 gnd.n6501 19.3944
R11113 gnd.n6845 gnd.n6501 19.3944
R11114 gnd.n6845 gnd.n6844 19.3944
R11115 gnd.n6844 gnd.n6843 19.3944
R11116 gnd.n6843 gnd.n6505 19.3944
R11117 gnd.n6839 gnd.n6505 19.3944
R11118 gnd.n6839 gnd.n6838 19.3944
R11119 gnd.n6838 gnd.n6837 19.3944
R11120 gnd.n6837 gnd.n6794 19.3944
R11121 gnd.n6833 gnd.n6794 19.3944
R11122 gnd.n6833 gnd.n6832 19.3944
R11123 gnd.n6832 gnd.n6831 19.3944
R11124 gnd.n6831 gnd.n6798 19.3944
R11125 gnd.n6827 gnd.n6798 19.3944
R11126 gnd.n6827 gnd.n6826 19.3944
R11127 gnd.n6826 gnd.n6825 19.3944
R11128 gnd.n6825 gnd.n6802 19.3944
R11129 gnd.n6821 gnd.n6802 19.3944
R11130 gnd.n6821 gnd.n6820 19.3944
R11131 gnd.n6820 gnd.n6819 19.3944
R11132 gnd.n6819 gnd.n6806 19.3944
R11133 gnd.n6815 gnd.n6806 19.3944
R11134 gnd.n6815 gnd.n6814 19.3944
R11135 gnd.n6814 gnd.n6813 19.3944
R11136 gnd.n6813 gnd.n6810 19.3944
R11137 gnd.n6810 gnd.n750 19.3944
R11138 gnd.n7092 gnd.n750 19.3944
R11139 gnd.n7089 gnd.n7088 19.3944
R11140 gnd.n7088 gnd.n7087 19.3944
R11141 gnd.n7087 gnd.n755 19.3944
R11142 gnd.n7083 gnd.n755 19.3944
R11143 gnd.n7083 gnd.n7082 19.3944
R11144 gnd.n7082 gnd.n679 19.3944
R11145 gnd.n7156 gnd.n679 19.3944
R11146 gnd.n7156 gnd.n7155 19.3944
R11147 gnd.n7155 gnd.n7154 19.3944
R11148 gnd.n7154 gnd.n683 19.3944
R11149 gnd.n7147 gnd.n683 19.3944
R11150 gnd.n7147 gnd.n7146 19.3944
R11151 gnd.n7146 gnd.n693 19.3944
R11152 gnd.n7139 gnd.n693 19.3944
R11153 gnd.n7139 gnd.n7138 19.3944
R11154 gnd.n7138 gnd.n703 19.3944
R11155 gnd.n7131 gnd.n703 19.3944
R11156 gnd.n7131 gnd.n7130 19.3944
R11157 gnd.n7130 gnd.n711 19.3944
R11158 gnd.n7123 gnd.n711 19.3944
R11159 gnd.n7123 gnd.n7122 19.3944
R11160 gnd.n7122 gnd.n721 19.3944
R11161 gnd.n7115 gnd.n721 19.3944
R11162 gnd.n7115 gnd.n7114 19.3944
R11163 gnd.n7104 gnd.n737 19.3944
R11164 gnd.n7104 gnd.n7103 19.3944
R11165 gnd.n7103 gnd.n740 19.3944
R11166 gnd.n1431 gnd.n1430 19.2005
R11167 gnd.n6788 gnd.n6787 19.2005
R11168 gnd.n5314 gnd.n5313 19.1977
R11169 gnd.n5838 gnd.n1130 19.1199
R11170 gnd.n6357 gnd.n6356 19.1199
R11171 gnd.n1011 gnd.n984 19.1199
R11172 gnd.n6620 gnd.n877 19.1199
R11173 gnd.n4699 gnd.t14 18.8012
R11174 gnd.n4684 gnd.t59 18.8012
R11175 gnd.n5884 gnd.t57 18.8012
R11176 gnd.n6594 gnd.t61 18.8012
R11177 gnd.n4543 gnd.n4542 18.4825
R11178 gnd.n7223 gnd.n7222 18.4247
R11179 gnd.n6102 gnd.n6101 18.4247
R11180 gnd.n7111 gnd.n7110 18.2308
R11181 gnd.n5681 gnd.n1239 18.2308
R11182 gnd.n7718 gnd.n7669 18.2308
R11183 gnd.n3470 gnd.n3469 18.2308
R11184 gnd.t41 gnd.n4223 18.1639
R11185 gnd.n1326 gnd.n1324 17.8452
R11186 gnd.n5832 gnd.n1123 17.8452
R11187 gnd.n1054 gnd.n1049 17.8452
R11188 gnd.n6423 gnd.n993 17.8452
R11189 gnd.n6857 gnd.n884 17.8452
R11190 gnd.n6792 gnd.n849 17.8452
R11191 gnd.n4251 gnd.t16 17.5266
R11192 gnd.n5816 gnd.t27 17.2079
R11193 gnd.n948 gnd.t26 17.2079
R11194 gnd.n4650 gnd.t31 16.8893
R11195 gnd.n7205 gnd.n7202 16.6793
R11196 gnd.n7811 gnd.n7808 16.6793
R11197 gnd.n3760 gnd.n3757 16.6793
R11198 gnd.n1534 gnd.n1504 16.6793
R11199 gnd.n5827 gnd.n1116 16.5706
R11200 gnd.n5811 gnd.t51 16.5706
R11201 gnd.n1044 gnd.n1034 16.5706
R11202 gnd.n6414 gnd.n1024 16.5706
R11203 gnd.n6886 gnd.t38 16.5706
R11204 gnd.n962 gnd.n891 16.5706
R11205 gnd.n4478 gnd.t91 16.2519
R11206 gnd.n4178 gnd.t42 16.2519
R11207 gnd.n5960 gnd.t0 15.9333
R11208 gnd.n6894 gnd.t9 15.9333
R11209 gnd.n5165 gnd.n5163 15.6674
R11210 gnd.n5133 gnd.n5131 15.6674
R11211 gnd.n5101 gnd.n5099 15.6674
R11212 gnd.n5070 gnd.n5068 15.6674
R11213 gnd.n5038 gnd.n5036 15.6674
R11214 gnd.n5006 gnd.n5004 15.6674
R11215 gnd.n4974 gnd.n4972 15.6674
R11216 gnd.n4943 gnd.n4941 15.6674
R11217 gnd.n4469 gnd.t91 15.6146
R11218 gnd.t195 gnd.n3900 15.6146
R11219 gnd.t167 gnd.n3901 15.6146
R11220 gnd.n7162 gnd.n674 15.3217
R11221 gnd.n7766 gnd.n349 15.3217
R11222 gnd.n3717 gnd.n3267 15.3217
R11223 gnd.n1589 gnd.n1482 15.3217
R11224 gnd.n6292 gnd.n1116 15.296
R11225 gnd.n5822 gnd.n5821 15.296
R11226 gnd.n5800 gnd.t28 15.296
R11227 gnd.n6404 gnd.n1034 15.296
R11228 gnd.n6395 gnd.n1024 15.296
R11229 gnd.n6448 gnd.t36 15.296
R11230 gnd.n6872 gnd.n6871 15.296
R11231 gnd.n6940 gnd.n891 15.296
R11232 gnd.t106 gnd.n6653 15.296
R11233 gnd.n6516 gnd.n6515 15.0827
R11234 gnd.n1336 gnd.n1331 15.0481
R11235 gnd.n6526 gnd.n6525 15.0481
R11236 gnd.n4837 gnd.t70 14.9773
R11237 gnd.n5948 gnd.t47 14.6587
R11238 gnd.t46 gnd.n985 14.6587
R11239 gnd.n6590 gnd.t103 14.6587
R11240 gnd.t409 gnd.n3943 14.34
R11241 gnd.n4915 gnd.t68 14.34
R11242 gnd.n6023 gnd.t6 14.34
R11243 gnd.n6652 gnd.t414 14.34
R11244 gnd.n6284 gnd.n1123 14.0214
R11245 gnd.n5816 gnd.n5815 14.0214
R11246 gnd.n6364 gnd.t1 14.0214
R11247 gnd.n1055 gnd.n1054 14.0214
R11248 gnd.n6462 gnd.n993 14.0214
R11249 gnd.t66 gnd.n995 14.0214
R11250 gnd.n948 gnd.n946 14.0214
R11251 gnd.n6948 gnd.n884 14.0214
R11252 gnd.n6988 gnd.n849 14.0214
R11253 gnd.n4625 gnd.t79 13.7027
R11254 gnd.n6346 gnd.t73 13.7027
R11255 gnd.n6440 gnd.t55 13.7027
R11256 gnd.n4335 gnd.n4334 13.5763
R11257 gnd.n5279 gnd.n3857 13.5763
R11258 gnd.n4543 gnd.n4281 13.384
R11259 gnd.t413 gnd.n1032 13.384
R11260 gnd.n6394 gnd.t2 13.384
R11261 gnd.n1347 gnd.n1328 13.1884
R11262 gnd.n1342 gnd.n1341 13.1884
R11263 gnd.n1341 gnd.n1340 13.1884
R11264 gnd.n6519 gnd.n6514 13.1884
R11265 gnd.n6520 gnd.n6519 13.1884
R11266 gnd.n1343 gnd.n1330 13.146
R11267 gnd.n1339 gnd.n1330 13.146
R11268 gnd.n6518 gnd.n6517 13.146
R11269 gnd.n6518 gnd.n6513 13.146
R11270 gnd.n3604 gnd.t251 13.0654
R11271 gnd.n394 gnd.t259 13.0654
R11272 gnd.n5166 gnd.n5162 12.8005
R11273 gnd.n5134 gnd.n5130 12.8005
R11274 gnd.n5102 gnd.n5098 12.8005
R11275 gnd.n5071 gnd.n5067 12.8005
R11276 gnd.n5039 gnd.n5035 12.8005
R11277 gnd.n5007 gnd.n5003 12.8005
R11278 gnd.n4975 gnd.n4971 12.8005
R11279 gnd.n4944 gnd.n4940 12.8005
R11280 gnd.n6252 gnd.n1151 12.7467
R11281 gnd.n5850 gnd.t164 12.7467
R11282 gnd.n6276 gnd.n1130 12.7467
R11283 gnd.n6357 gnd.n1059 12.7467
R11284 gnd.n6472 gnd.n984 12.7467
R11285 gnd.n6956 gnd.n877 12.7467
R11286 gnd.n6791 gnd.t151 12.7467
R11287 gnd.n3685 gnd.t278 12.4281
R11288 gnd.n5424 gnd.t287 12.4281
R11289 gnd.n1680 gnd.t309 12.4281
R11290 gnd.t63 gnd.n1202 12.4281
R11291 gnd.n807 gnd.t20 12.4281
R11292 gnd.n7371 gnd.t248 12.4281
R11293 gnd.t207 gnd.n448 12.4281
R11294 gnd.n7915 gnd.t233 12.4281
R11295 gnd.n4334 gnd.n4329 12.4126
R11296 gnd.n5282 gnd.n5279 12.4126
R11297 gnd.n1430 gnd.n1429 12.1761
R11298 gnd.n6787 gnd.n6786 12.1761
R11299 gnd.n5523 gnd.n1253 12.1094
R11300 gnd.n6244 gnd.t110 12.1094
R11301 gnd.n7275 gnd.n7274 12.1094
R11302 gnd.n5170 gnd.n5169 12.0247
R11303 gnd.n5138 gnd.n5137 12.0247
R11304 gnd.n5106 gnd.n5105 12.0247
R11305 gnd.n5075 gnd.n5074 12.0247
R11306 gnd.n5043 gnd.n5042 12.0247
R11307 gnd.n5011 gnd.n5010 12.0247
R11308 gnd.n4979 gnd.n4978 12.0247
R11309 gnd.n4948 gnd.n4947 12.0247
R11310 gnd.n3661 gnd.t253 11.7908
R11311 gnd.n5452 gnd.t287 11.7908
R11312 gnd.t309 gnd.n1640 11.7908
R11313 gnd.t248 gnd.n486 11.7908
R11314 gnd.n7448 gnd.t207 11.7908
R11315 gnd.n7939 gnd.t271 11.7908
R11316 gnd.n6260 gnd.n1143 11.4721
R11317 gnd.n6268 gnd.n1137 11.4721
R11318 gnd.n5960 gnd.n5959 11.4721
R11319 gnd.n5970 gnd.n5969 11.4721
R11320 gnd.n6449 gnd.n1003 11.4721
R11321 gnd.n6894 gnd.n934 11.4721
R11322 gnd.n6964 gnd.n870 11.4721
R11323 gnd.n6972 gnd.n864 11.4721
R11324 gnd.n5173 gnd.n5160 11.249
R11325 gnd.n5141 gnd.n5128 11.249
R11326 gnd.n5109 gnd.n5096 11.249
R11327 gnd.n5078 gnd.n5065 11.249
R11328 gnd.n5046 gnd.n5033 11.249
R11329 gnd.n5014 gnd.n5001 11.249
R11330 gnd.n4982 gnd.n4969 11.249
R11331 gnd.n4951 gnd.n4938 11.249
R11332 gnd.n4613 gnd.t79 11.1535
R11333 gnd.n3637 gnd.t269 11.1535
R11334 gnd.n5366 gnd.t251 11.1535
R11335 gnd.n5811 gnd.t23 11.1535
R11336 gnd.t83 gnd.n6886 11.1535
R11337 gnd.n7536 gnd.t259 11.1535
R11338 gnd.n7963 gnd.t229 11.1535
R11339 gnd.n7165 gnd.n7162 10.6672
R11340 gnd.n7769 gnd.n7766 10.6672
R11341 gnd.n3720 gnd.n3717 10.6672
R11342 gnd.n1584 gnd.n1482 10.6672
R11343 gnd.n6721 gnd.n6557 10.6151
R11344 gnd.n6721 gnd.n6720 10.6151
R11345 gnd.n6718 gnd.n6561 10.6151
R11346 gnd.n6713 gnd.n6561 10.6151
R11347 gnd.n6713 gnd.n6712 10.6151
R11348 gnd.n6712 gnd.n6711 10.6151
R11349 gnd.n6711 gnd.n6564 10.6151
R11350 gnd.n6706 gnd.n6564 10.6151
R11351 gnd.n6706 gnd.n6705 10.6151
R11352 gnd.n6705 gnd.n6704 10.6151
R11353 gnd.n6704 gnd.n6567 10.6151
R11354 gnd.n6699 gnd.n6567 10.6151
R11355 gnd.n6699 gnd.n6698 10.6151
R11356 gnd.n6698 gnd.n6697 10.6151
R11357 gnd.n6697 gnd.n6570 10.6151
R11358 gnd.n6692 gnd.n6570 10.6151
R11359 gnd.n6692 gnd.n6691 10.6151
R11360 gnd.n6691 gnd.n6690 10.6151
R11361 gnd.n6690 gnd.n6573 10.6151
R11362 gnd.n6685 gnd.n6573 10.6151
R11363 gnd.n6685 gnd.n6684 10.6151
R11364 gnd.n6684 gnd.n6683 10.6151
R11365 gnd.n6683 gnd.n6576 10.6151
R11366 gnd.n6678 gnd.n6576 10.6151
R11367 gnd.n6678 gnd.n6677 10.6151
R11368 gnd.n6677 gnd.n6676 10.6151
R11369 gnd.n6676 gnd.n6579 10.6151
R11370 gnd.n6671 gnd.n6579 10.6151
R11371 gnd.n6671 gnd.n6670 10.6151
R11372 gnd.n6670 gnd.n6669 10.6151
R11373 gnd.n1323 gnd.n1321 10.6151
R11374 gnd.n5855 gnd.n1323 10.6151
R11375 gnd.n5857 gnd.n5855 10.6151
R11376 gnd.n5858 gnd.n5857 10.6151
R11377 gnd.n5860 gnd.n5858 10.6151
R11378 gnd.n5861 gnd.n5860 10.6151
R11379 gnd.n5862 gnd.n5861 10.6151
R11380 gnd.n5862 gnd.n5853 10.6151
R11381 gnd.n5878 gnd.n5853 10.6151
R11382 gnd.n5879 gnd.n5878 10.6151
R11383 gnd.n5882 gnd.n5879 10.6151
R11384 gnd.n5882 gnd.n5881 10.6151
R11385 gnd.n5881 gnd.n5880 10.6151
R11386 gnd.n5880 gnd.n5842 10.6151
R11387 gnd.n5896 gnd.n5842 10.6151
R11388 gnd.n5897 gnd.n5896 10.6151
R11389 gnd.n5900 gnd.n5897 10.6151
R11390 gnd.n5900 gnd.n5899 10.6151
R11391 gnd.n5899 gnd.n5898 10.6151
R11392 gnd.n5898 gnd.n5830 10.6151
R11393 gnd.n5913 gnd.n5830 10.6151
R11394 gnd.n5914 gnd.n5913 10.6151
R11395 gnd.n5916 gnd.n5914 10.6151
R11396 gnd.n5916 gnd.n5915 10.6151
R11397 gnd.n5915 gnd.n5819 10.6151
R11398 gnd.n5929 gnd.n5819 10.6151
R11399 gnd.n5930 gnd.n5929 10.6151
R11400 gnd.n5932 gnd.n5930 10.6151
R11401 gnd.n5932 gnd.n5931 10.6151
R11402 gnd.n5931 gnd.n5808 10.6151
R11403 gnd.n5944 gnd.n5808 10.6151
R11404 gnd.n5945 gnd.n5944 10.6151
R11405 gnd.n5957 gnd.n5945 10.6151
R11406 gnd.n5957 gnd.n5956 10.6151
R11407 gnd.n5956 gnd.n5955 10.6151
R11408 gnd.n5955 gnd.n5954 10.6151
R11409 gnd.n5954 gnd.n5952 10.6151
R11410 gnd.n5952 gnd.n5951 10.6151
R11411 gnd.n5951 gnd.n5947 10.6151
R11412 gnd.n5947 gnd.n5946 10.6151
R11413 gnd.n5946 gnd.n1052 10.6151
R11414 gnd.n6366 gnd.n1052 10.6151
R11415 gnd.n6367 gnd.n6366 10.6151
R11416 gnd.n6370 gnd.n6367 10.6151
R11417 gnd.n6370 gnd.n6369 10.6151
R11418 gnd.n6369 gnd.n6368 10.6151
R11419 gnd.n6368 gnd.n1042 10.6151
R11420 gnd.n6386 gnd.n1042 10.6151
R11421 gnd.n6387 gnd.n6386 10.6151
R11422 gnd.n6392 gnd.n6387 10.6151
R11423 gnd.n6392 gnd.n6391 10.6151
R11424 gnd.n6391 gnd.n6390 10.6151
R11425 gnd.n6390 gnd.n6388 10.6151
R11426 gnd.n6388 gnd.n1009 10.6151
R11427 gnd.n6435 gnd.n1009 10.6151
R11428 gnd.n6436 gnd.n6435 10.6151
R11429 gnd.n6438 gnd.n6436 10.6151
R11430 gnd.n6438 gnd.n6437 10.6151
R11431 gnd.n6437 gnd.n931 10.6151
R11432 gnd.n6898 gnd.n931 10.6151
R11433 gnd.n6898 gnd.n6897 10.6151
R11434 gnd.n6897 gnd.n6896 10.6151
R11435 gnd.n6896 gnd.n932 10.6151
R11436 gnd.n943 gnd.n932 10.6151
R11437 gnd.n6884 gnd.n943 10.6151
R11438 gnd.n6884 gnd.n6883 10.6151
R11439 gnd.n6883 gnd.n6882 10.6151
R11440 gnd.n6882 gnd.n944 10.6151
R11441 gnd.n957 gnd.n944 10.6151
R11442 gnd.n958 gnd.n957 10.6151
R11443 gnd.n6869 gnd.n958 10.6151
R11444 gnd.n6869 gnd.n6868 10.6151
R11445 gnd.n6868 gnd.n6867 10.6151
R11446 gnd.n6867 gnd.n959 10.6151
R11447 gnd.n6611 gnd.n959 10.6151
R11448 gnd.n6612 gnd.n6611 10.6151
R11449 gnd.n6614 gnd.n6612 10.6151
R11450 gnd.n6615 gnd.n6614 10.6151
R11451 gnd.n6618 gnd.n6615 10.6151
R11452 gnd.n6618 gnd.n6617 10.6151
R11453 gnd.n6617 gnd.n6616 10.6151
R11454 gnd.n6616 gnd.n6597 10.6151
R11455 gnd.n6633 gnd.n6597 10.6151
R11456 gnd.n6634 gnd.n6633 10.6151
R11457 gnd.n6636 gnd.n6634 10.6151
R11458 gnd.n6636 gnd.n6635 10.6151
R11459 gnd.n6635 gnd.n6588 10.6151
R11460 gnd.n6647 gnd.n6588 10.6151
R11461 gnd.n6648 gnd.n6647 10.6151
R11462 gnd.n6650 gnd.n6648 10.6151
R11463 gnd.n6650 gnd.n6649 10.6151
R11464 gnd.n6649 gnd.n6582 10.6151
R11465 gnd.n6663 gnd.n6582 10.6151
R11466 gnd.n6664 gnd.n6663 10.6151
R11467 gnd.n6665 gnd.n6664 10.6151
R11468 gnd.n6094 gnd.n1301 10.6151
R11469 gnd.n6094 gnd.n6093 10.6151
R11470 gnd.n6091 gnd.n1307 10.6151
R11471 gnd.n6085 gnd.n1307 10.6151
R11472 gnd.n6085 gnd.n6084 10.6151
R11473 gnd.n6084 gnd.n6083 10.6151
R11474 gnd.n6083 gnd.n1309 10.6151
R11475 gnd.n6077 gnd.n1309 10.6151
R11476 gnd.n6077 gnd.n6076 10.6151
R11477 gnd.n6076 gnd.n6075 10.6151
R11478 gnd.n6075 gnd.n1311 10.6151
R11479 gnd.n6069 gnd.n1311 10.6151
R11480 gnd.n6069 gnd.n6068 10.6151
R11481 gnd.n6068 gnd.n6067 10.6151
R11482 gnd.n6067 gnd.n1313 10.6151
R11483 gnd.n6061 gnd.n1313 10.6151
R11484 gnd.n6061 gnd.n6060 10.6151
R11485 gnd.n6060 gnd.n6059 10.6151
R11486 gnd.n6059 gnd.n1315 10.6151
R11487 gnd.n6053 gnd.n1315 10.6151
R11488 gnd.n6053 gnd.n6052 10.6151
R11489 gnd.n6052 gnd.n6051 10.6151
R11490 gnd.n6051 gnd.n1317 10.6151
R11491 gnd.n6045 gnd.n1317 10.6151
R11492 gnd.n6045 gnd.n6044 10.6151
R11493 gnd.n6044 gnd.n6043 10.6151
R11494 gnd.n6043 gnd.n1319 10.6151
R11495 gnd.n6037 gnd.n1319 10.6151
R11496 gnd.n6037 gnd.n6036 10.6151
R11497 gnd.n6036 gnd.n6035 10.6151
R11498 gnd.n1429 gnd.n1348 10.6151
R11499 gnd.n1424 gnd.n1348 10.6151
R11500 gnd.n1424 gnd.n1423 10.6151
R11501 gnd.n1423 gnd.n1422 10.6151
R11502 gnd.n1422 gnd.n1350 10.6151
R11503 gnd.n1416 gnd.n1350 10.6151
R11504 gnd.n1416 gnd.n1415 10.6151
R11505 gnd.n1415 gnd.n1414 10.6151
R11506 gnd.n1414 gnd.n1352 10.6151
R11507 gnd.n1408 gnd.n1352 10.6151
R11508 gnd.n1408 gnd.n1407 10.6151
R11509 gnd.n1407 gnd.n1406 10.6151
R11510 gnd.n1406 gnd.n1354 10.6151
R11511 gnd.n1400 gnd.n1354 10.6151
R11512 gnd.n1400 gnd.n1399 10.6151
R11513 gnd.n1399 gnd.n1398 10.6151
R11514 gnd.n1398 gnd.n1356 10.6151
R11515 gnd.n1392 gnd.n1356 10.6151
R11516 gnd.n1392 gnd.n1391 10.6151
R11517 gnd.n1391 gnd.n1390 10.6151
R11518 gnd.n1390 gnd.n1358 10.6151
R11519 gnd.n1384 gnd.n1358 10.6151
R11520 gnd.n1384 gnd.n1383 10.6151
R11521 gnd.n1383 gnd.n1382 10.6151
R11522 gnd.n1382 gnd.n1360 10.6151
R11523 gnd.n1376 gnd.n1360 10.6151
R11524 gnd.n1376 gnd.n1375 10.6151
R11525 gnd.n1375 gnd.n1374 10.6151
R11526 gnd.n1370 gnd.n1369 10.6151
R11527 gnd.n1369 gnd.n1302 10.6151
R11528 gnd.n6786 gnd.n6531 10.6151
R11529 gnd.n6533 gnd.n6531 10.6151
R11530 gnd.n6779 gnd.n6533 10.6151
R11531 gnd.n6779 gnd.n6778 10.6151
R11532 gnd.n6778 gnd.n6777 10.6151
R11533 gnd.n6777 gnd.n6535 10.6151
R11534 gnd.n6772 gnd.n6535 10.6151
R11535 gnd.n6772 gnd.n6771 10.6151
R11536 gnd.n6771 gnd.n6770 10.6151
R11537 gnd.n6770 gnd.n6538 10.6151
R11538 gnd.n6765 gnd.n6538 10.6151
R11539 gnd.n6765 gnd.n6764 10.6151
R11540 gnd.n6764 gnd.n6763 10.6151
R11541 gnd.n6763 gnd.n6541 10.6151
R11542 gnd.n6758 gnd.n6541 10.6151
R11543 gnd.n6758 gnd.n6757 10.6151
R11544 gnd.n6757 gnd.n6756 10.6151
R11545 gnd.n6756 gnd.n6544 10.6151
R11546 gnd.n6751 gnd.n6544 10.6151
R11547 gnd.n6751 gnd.n6750 10.6151
R11548 gnd.n6750 gnd.n6749 10.6151
R11549 gnd.n6749 gnd.n6547 10.6151
R11550 gnd.n6744 gnd.n6547 10.6151
R11551 gnd.n6744 gnd.n6743 10.6151
R11552 gnd.n6743 gnd.n6742 10.6151
R11553 gnd.n6742 gnd.n6550 10.6151
R11554 gnd.n6737 gnd.n6550 10.6151
R11555 gnd.n6737 gnd.n6736 10.6151
R11556 gnd.n6734 gnd.n6555 10.6151
R11557 gnd.n6729 gnd.n6555 10.6151
R11558 gnd.n6028 gnd.n1431 10.6151
R11559 gnd.n6028 gnd.n6027 10.6151
R11560 gnd.n6027 gnd.n6026 10.6151
R11561 gnd.n6026 gnd.n1432 10.6151
R11562 gnd.n5866 gnd.n1432 10.6151
R11563 gnd.n5867 gnd.n5866 10.6151
R11564 gnd.n5872 gnd.n5867 10.6151
R11565 gnd.n5872 gnd.n5871 10.6151
R11566 gnd.n5871 gnd.n5870 10.6151
R11567 gnd.n5870 gnd.n5868 10.6151
R11568 gnd.n5868 gnd.n5848 10.6151
R11569 gnd.n5887 gnd.n5848 10.6151
R11570 gnd.n5888 gnd.n5887 10.6151
R11571 gnd.n5891 gnd.n5888 10.6151
R11572 gnd.n5891 gnd.n5890 10.6151
R11573 gnd.n5890 gnd.n5889 10.6151
R11574 gnd.n5889 gnd.n5836 10.6151
R11575 gnd.n5905 gnd.n5836 10.6151
R11576 gnd.n5906 gnd.n5905 10.6151
R11577 gnd.n5908 gnd.n5906 10.6151
R11578 gnd.n5908 gnd.n5907 10.6151
R11579 gnd.n5907 gnd.n5825 10.6151
R11580 gnd.n5920 gnd.n5825 10.6151
R11581 gnd.n5921 gnd.n5920 10.6151
R11582 gnd.n5924 gnd.n5921 10.6151
R11583 gnd.n5924 gnd.n5923 10.6151
R11584 gnd.n5923 gnd.n5922 10.6151
R11585 gnd.n5922 gnd.n5813 10.6151
R11586 gnd.n5937 gnd.n5813 10.6151
R11587 gnd.n5938 gnd.n5937 10.6151
R11588 gnd.n5940 gnd.n5938 10.6151
R11589 gnd.n5940 gnd.n5939 10.6151
R11590 gnd.n5939 gnd.n5804 10.6151
R11591 gnd.n5963 gnd.n5804 10.6151
R11592 gnd.n5964 gnd.n5963 10.6151
R11593 gnd.n5965 gnd.n5964 10.6151
R11594 gnd.n5967 gnd.n5965 10.6151
R11595 gnd.n5967 gnd.n5966 10.6151
R11596 gnd.n5966 gnd.n1057 10.6151
R11597 gnd.n6359 gnd.n1057 10.6151
R11598 gnd.n6360 gnd.n6359 10.6151
R11599 gnd.n6362 gnd.n6360 10.6151
R11600 gnd.n6362 gnd.n6361 10.6151
R11601 gnd.n6361 gnd.n1047 10.6151
R11602 gnd.n6375 gnd.n1047 10.6151
R11603 gnd.n6376 gnd.n6375 10.6151
R11604 gnd.n6381 gnd.n6376 10.6151
R11605 gnd.n6381 gnd.n6380 10.6151
R11606 gnd.n6380 gnd.n6379 10.6151
R11607 gnd.n6379 gnd.n6377 10.6151
R11608 gnd.n6377 gnd.n1014 10.6151
R11609 gnd.n6427 gnd.n1014 10.6151
R11610 gnd.n6428 gnd.n6427 10.6151
R11611 gnd.n6430 gnd.n6428 10.6151
R11612 gnd.n6430 gnd.n6429 10.6151
R11613 gnd.n6429 gnd.n1005 10.6151
R11614 gnd.n6443 gnd.n1005 10.6151
R11615 gnd.n6444 gnd.n6443 10.6151
R11616 gnd.n6446 gnd.n6444 10.6151
R11617 gnd.n6446 gnd.n6445 10.6151
R11618 gnd.n6445 gnd.n937 10.6151
R11619 gnd.n6892 gnd.n937 10.6151
R11620 gnd.n6892 gnd.n6891 10.6151
R11621 gnd.n6891 gnd.n6890 10.6151
R11622 gnd.n6890 gnd.n938 10.6151
R11623 gnd.n950 gnd.n938 10.6151
R11624 gnd.n6878 gnd.n950 10.6151
R11625 gnd.n6878 gnd.n6877 10.6151
R11626 gnd.n6877 gnd.n6876 10.6151
R11627 gnd.n6876 gnd.n951 10.6151
R11628 gnd.n965 gnd.n951 10.6151
R11629 gnd.n966 gnd.n965 10.6151
R11630 gnd.n6863 gnd.n966 10.6151
R11631 gnd.n6863 gnd.n6862 10.6151
R11632 gnd.n6862 gnd.n6861 10.6151
R11633 gnd.n6861 gnd.n967 10.6151
R11634 gnd.n6605 gnd.n967 10.6151
R11635 gnd.n6606 gnd.n6605 10.6151
R11636 gnd.n6606 gnd.n6603 10.6151
R11637 gnd.n6624 gnd.n6603 10.6151
R11638 gnd.n6625 gnd.n6624 10.6151
R11639 gnd.n6628 gnd.n6625 10.6151
R11640 gnd.n6628 gnd.n6627 10.6151
R11641 gnd.n6627 gnd.n6626 10.6151
R11642 gnd.n6626 gnd.n6592 10.6151
R11643 gnd.n6641 gnd.n6592 10.6151
R11644 gnd.n6642 gnd.n6641 10.6151
R11645 gnd.n6643 gnd.n6642 10.6151
R11646 gnd.n6643 gnd.n6585 10.6151
R11647 gnd.n6656 gnd.n6585 10.6151
R11648 gnd.n6657 gnd.n6656 10.6151
R11649 gnd.n6658 gnd.n6657 10.6151
R11650 gnd.n6658 gnd.n6511 10.6151
R11651 gnd.n6789 gnd.n6511 10.6151
R11652 gnd.n6789 gnd.n6788 10.6151
R11653 gnd.n4532 gnd.t4 10.5161
R11654 gnd.n3945 gnd.t409 10.5161
R11655 gnd.n4898 gnd.t68 10.5161
R11656 gnd.n5341 gnd.t219 10.5161
R11657 gnd.n5333 gnd.t283 10.5161
R11658 gnd.n6300 gnd.t71 10.5161
R11659 gnd.n6932 gnd.t32 10.5161
R11660 gnd.n7561 gnd.t240 10.5161
R11661 gnd.n7570 gnd.t209 10.5161
R11662 gnd.n5174 gnd.n5158 10.4732
R11663 gnd.n5142 gnd.n5126 10.4732
R11664 gnd.n5110 gnd.n5094 10.4732
R11665 gnd.n5079 gnd.n5063 10.4732
R11666 gnd.n5047 gnd.n5031 10.4732
R11667 gnd.n5015 gnd.n4999 10.4732
R11668 gnd.n4983 gnd.n4967 10.4732
R11669 gnd.n4952 gnd.n4936 10.4732
R11670 gnd.n6260 gnd.n1145 10.1975
R11671 gnd.n5959 gnd.n1079 10.1975
R11672 gnd.n5970 gnd.n5800 10.1975
R11673 gnd.n6449 gnd.n6448 10.1975
R11674 gnd.n934 gnd.n927 10.1975
R11675 gnd.n6972 gnd.n862 10.1975
R11676 gnd.t70 gnd.n3962 9.87883
R11677 gnd.n3643 gnd.t211 9.87883
R11678 gnd.n7957 gnd.t311 9.87883
R11679 gnd.n5178 gnd.n5177 9.69747
R11680 gnd.n5146 gnd.n5145 9.69747
R11681 gnd.n5114 gnd.n5113 9.69747
R11682 gnd.n5083 gnd.n5082 9.69747
R11683 gnd.n5051 gnd.n5050 9.69747
R11684 gnd.n5019 gnd.n5018 9.69747
R11685 gnd.n4987 gnd.n4986 9.69747
R11686 gnd.n4956 gnd.n4955 9.69747
R11687 gnd.n5184 gnd.n5183 9.45567
R11688 gnd.n5152 gnd.n5151 9.45567
R11689 gnd.n5120 gnd.n5119 9.45567
R11690 gnd.n5089 gnd.n5088 9.45567
R11691 gnd.n5057 gnd.n5056 9.45567
R11692 gnd.n5025 gnd.n5024 9.45567
R11693 gnd.n4993 gnd.n4992 9.45567
R11694 gnd.n4962 gnd.n4961 9.45567
R11695 gnd.n7202 gnd.n7201 9.30959
R11696 gnd.n7808 gnd.n329 9.30959
R11697 gnd.n3757 gnd.n3756 9.30959
R11698 gnd.n1540 gnd.n1504 9.30959
R11699 gnd.n5183 gnd.n5182 9.3005
R11700 gnd.n5156 gnd.n5155 9.3005
R11701 gnd.n5177 gnd.n5176 9.3005
R11702 gnd.n5175 gnd.n5174 9.3005
R11703 gnd.n5160 gnd.n5159 9.3005
R11704 gnd.n5169 gnd.n5168 9.3005
R11705 gnd.n5167 gnd.n5166 9.3005
R11706 gnd.n5151 gnd.n5150 9.3005
R11707 gnd.n5124 gnd.n5123 9.3005
R11708 gnd.n5145 gnd.n5144 9.3005
R11709 gnd.n5143 gnd.n5142 9.3005
R11710 gnd.n5128 gnd.n5127 9.3005
R11711 gnd.n5137 gnd.n5136 9.3005
R11712 gnd.n5135 gnd.n5134 9.3005
R11713 gnd.n5119 gnd.n5118 9.3005
R11714 gnd.n5092 gnd.n5091 9.3005
R11715 gnd.n5113 gnd.n5112 9.3005
R11716 gnd.n5111 gnd.n5110 9.3005
R11717 gnd.n5096 gnd.n5095 9.3005
R11718 gnd.n5105 gnd.n5104 9.3005
R11719 gnd.n5103 gnd.n5102 9.3005
R11720 gnd.n5088 gnd.n5087 9.3005
R11721 gnd.n5061 gnd.n5060 9.3005
R11722 gnd.n5082 gnd.n5081 9.3005
R11723 gnd.n5080 gnd.n5079 9.3005
R11724 gnd.n5065 gnd.n5064 9.3005
R11725 gnd.n5074 gnd.n5073 9.3005
R11726 gnd.n5072 gnd.n5071 9.3005
R11727 gnd.n5056 gnd.n5055 9.3005
R11728 gnd.n5029 gnd.n5028 9.3005
R11729 gnd.n5050 gnd.n5049 9.3005
R11730 gnd.n5048 gnd.n5047 9.3005
R11731 gnd.n5033 gnd.n5032 9.3005
R11732 gnd.n5042 gnd.n5041 9.3005
R11733 gnd.n5040 gnd.n5039 9.3005
R11734 gnd.n5024 gnd.n5023 9.3005
R11735 gnd.n4997 gnd.n4996 9.3005
R11736 gnd.n5018 gnd.n5017 9.3005
R11737 gnd.n5016 gnd.n5015 9.3005
R11738 gnd.n5001 gnd.n5000 9.3005
R11739 gnd.n5010 gnd.n5009 9.3005
R11740 gnd.n5008 gnd.n5007 9.3005
R11741 gnd.n4992 gnd.n4991 9.3005
R11742 gnd.n4965 gnd.n4964 9.3005
R11743 gnd.n4986 gnd.n4985 9.3005
R11744 gnd.n4984 gnd.n4983 9.3005
R11745 gnd.n4969 gnd.n4968 9.3005
R11746 gnd.n4978 gnd.n4977 9.3005
R11747 gnd.n4976 gnd.n4975 9.3005
R11748 gnd.n4961 gnd.n4960 9.3005
R11749 gnd.n4934 gnd.n4933 9.3005
R11750 gnd.n4955 gnd.n4954 9.3005
R11751 gnd.n4953 gnd.n4952 9.3005
R11752 gnd.n4938 gnd.n4937 9.3005
R11753 gnd.n4947 gnd.n4946 9.3005
R11754 gnd.n4945 gnd.n4944 9.3005
R11755 gnd.n5309 gnd.n5308 9.3005
R11756 gnd.n5307 gnd.n3845 9.3005
R11757 gnd.n5306 gnd.n5305 9.3005
R11758 gnd.n5302 gnd.n3846 9.3005
R11759 gnd.n5299 gnd.n3847 9.3005
R11760 gnd.n5298 gnd.n3848 9.3005
R11761 gnd.n5295 gnd.n3849 9.3005
R11762 gnd.n5294 gnd.n3850 9.3005
R11763 gnd.n5291 gnd.n3851 9.3005
R11764 gnd.n5290 gnd.n3852 9.3005
R11765 gnd.n5287 gnd.n3853 9.3005
R11766 gnd.n5286 gnd.n3854 9.3005
R11767 gnd.n5283 gnd.n3855 9.3005
R11768 gnd.n5282 gnd.n3856 9.3005
R11769 gnd.n5279 gnd.n5278 9.3005
R11770 gnd.n5277 gnd.n3857 9.3005
R11771 gnd.n5310 gnd.n3844 9.3005
R11772 gnd.n4551 gnd.n4550 9.3005
R11773 gnd.n4255 gnd.n4254 9.3005
R11774 gnd.n4578 gnd.n4577 9.3005
R11775 gnd.n4579 gnd.n4253 9.3005
R11776 gnd.n4583 gnd.n4580 9.3005
R11777 gnd.n4582 gnd.n4581 9.3005
R11778 gnd.n4227 gnd.n4226 9.3005
R11779 gnd.n4608 gnd.n4607 9.3005
R11780 gnd.n4609 gnd.n4225 9.3005
R11781 gnd.n4611 gnd.n4610 9.3005
R11782 gnd.n4205 gnd.n4204 9.3005
R11783 gnd.n4639 gnd.n4638 9.3005
R11784 gnd.n4640 gnd.n4203 9.3005
R11785 gnd.n4648 gnd.n4641 9.3005
R11786 gnd.n4647 gnd.n4642 9.3005
R11787 gnd.n4646 gnd.n4644 9.3005
R11788 gnd.n4643 gnd.n4152 9.3005
R11789 gnd.n4696 gnd.n4153 9.3005
R11790 gnd.n4695 gnd.n4154 9.3005
R11791 gnd.n4694 gnd.n4155 9.3005
R11792 gnd.n4174 gnd.n4156 9.3005
R11793 gnd.n4176 gnd.n4175 9.3005
R11794 gnd.n4042 gnd.n4041 9.3005
R11795 gnd.n4734 gnd.n4733 9.3005
R11796 gnd.n4735 gnd.n4040 9.3005
R11797 gnd.n4739 gnd.n4736 9.3005
R11798 gnd.n4738 gnd.n4737 9.3005
R11799 gnd.n4015 gnd.n4014 9.3005
R11800 gnd.n4774 gnd.n4773 9.3005
R11801 gnd.n4775 gnd.n4013 9.3005
R11802 gnd.n4779 gnd.n4776 9.3005
R11803 gnd.n4778 gnd.n4777 9.3005
R11804 gnd.n3988 gnd.n3987 9.3005
R11805 gnd.n4819 gnd.n4818 9.3005
R11806 gnd.n4820 gnd.n3986 9.3005
R11807 gnd.n4824 gnd.n4821 9.3005
R11808 gnd.n4823 gnd.n4822 9.3005
R11809 gnd.n3960 gnd.n3959 9.3005
R11810 gnd.n4859 gnd.n4858 9.3005
R11811 gnd.n4860 gnd.n3958 9.3005
R11812 gnd.n4864 gnd.n4861 9.3005
R11813 gnd.n4863 gnd.n4862 9.3005
R11814 gnd.n3933 gnd.n3932 9.3005
R11815 gnd.n4908 gnd.n4907 9.3005
R11816 gnd.n4909 gnd.n3931 9.3005
R11817 gnd.n4913 gnd.n4910 9.3005
R11818 gnd.n4912 gnd.n4911 9.3005
R11819 gnd.n3906 gnd.n3905 9.3005
R11820 gnd.n5202 gnd.n5201 9.3005
R11821 gnd.n5203 gnd.n3904 9.3005
R11822 gnd.n5209 gnd.n5204 9.3005
R11823 gnd.n5208 gnd.n5205 9.3005
R11824 gnd.n5207 gnd.n5206 9.3005
R11825 gnd.n4552 gnd.n4549 9.3005
R11826 gnd.n4334 gnd.n4293 9.3005
R11827 gnd.n4329 gnd.n4328 9.3005
R11828 gnd.n4327 gnd.n4294 9.3005
R11829 gnd.n4326 gnd.n4325 9.3005
R11830 gnd.n4322 gnd.n4295 9.3005
R11831 gnd.n4319 gnd.n4318 9.3005
R11832 gnd.n4317 gnd.n4296 9.3005
R11833 gnd.n4316 gnd.n4315 9.3005
R11834 gnd.n4312 gnd.n4297 9.3005
R11835 gnd.n4309 gnd.n4308 9.3005
R11836 gnd.n4307 gnd.n4298 9.3005
R11837 gnd.n4306 gnd.n4305 9.3005
R11838 gnd.n4302 gnd.n4300 9.3005
R11839 gnd.n4299 gnd.n4279 9.3005
R11840 gnd.n4546 gnd.n4278 9.3005
R11841 gnd.n4548 gnd.n4547 9.3005
R11842 gnd.n4336 gnd.n4335 9.3005
R11843 gnd.n4559 gnd.n4265 9.3005
R11844 gnd.n4566 gnd.n4266 9.3005
R11845 gnd.n4568 gnd.n4567 9.3005
R11846 gnd.n4569 gnd.n4246 9.3005
R11847 gnd.n4588 gnd.n4587 9.3005
R11848 gnd.n4590 gnd.n4238 9.3005
R11849 gnd.n4597 gnd.n4240 9.3005
R11850 gnd.n4598 gnd.n4235 9.3005
R11851 gnd.n4600 gnd.n4599 9.3005
R11852 gnd.n4236 gnd.n4221 9.3005
R11853 gnd.n4616 gnd.n4219 9.3005
R11854 gnd.n4620 gnd.n4619 9.3005
R11855 gnd.n4618 gnd.n4195 9.3005
R11856 gnd.n4655 gnd.n4194 9.3005
R11857 gnd.n4658 gnd.n4657 9.3005
R11858 gnd.n4191 gnd.n4190 9.3005
R11859 gnd.n4664 gnd.n4192 9.3005
R11860 gnd.n4666 gnd.n4665 9.3005
R11861 gnd.n4668 gnd.n4189 9.3005
R11862 gnd.n4671 gnd.n4670 9.3005
R11863 gnd.n4674 gnd.n4672 9.3005
R11864 gnd.n4676 gnd.n4675 9.3005
R11865 gnd.n4682 gnd.n4677 9.3005
R11866 gnd.n4681 gnd.n4680 9.3005
R11867 gnd.n4033 gnd.n4032 9.3005
R11868 gnd.n4748 gnd.n4747 9.3005
R11869 gnd.n4749 gnd.n4026 9.3005
R11870 gnd.n4757 gnd.n4025 9.3005
R11871 gnd.n4760 gnd.n4759 9.3005
R11872 gnd.n4762 gnd.n4761 9.3005
R11873 gnd.n4765 gnd.n4008 9.3005
R11874 gnd.n4763 gnd.n4006 9.3005
R11875 gnd.n4785 gnd.n4004 9.3005
R11876 gnd.n4787 gnd.n4786 9.3005
R11877 gnd.n3978 gnd.n3977 9.3005
R11878 gnd.n4833 gnd.n4832 9.3005
R11879 gnd.n4834 gnd.n3971 9.3005
R11880 gnd.n4842 gnd.n3970 9.3005
R11881 gnd.n4845 gnd.n4844 9.3005
R11882 gnd.n4847 gnd.n4846 9.3005
R11883 gnd.n4850 gnd.n3953 9.3005
R11884 gnd.n4848 gnd.n3951 9.3005
R11885 gnd.n4870 gnd.n3949 9.3005
R11886 gnd.n4872 gnd.n4871 9.3005
R11887 gnd.n3924 gnd.n3923 9.3005
R11888 gnd.n4922 gnd.n4921 9.3005
R11889 gnd.n4923 gnd.n3917 9.3005
R11890 gnd.n4931 gnd.n3916 9.3005
R11891 gnd.n5190 gnd.n5189 9.3005
R11892 gnd.n5192 gnd.n5191 9.3005
R11893 gnd.n5193 gnd.n3897 9.3005
R11894 gnd.n5217 gnd.n5216 9.3005
R11895 gnd.n3898 gnd.n3860 9.3005
R11896 gnd.n4557 gnd.n4556 9.3005
R11897 gnd.n5273 gnd.n3861 9.3005
R11898 gnd.n5272 gnd.n3863 9.3005
R11899 gnd.n5269 gnd.n3864 9.3005
R11900 gnd.n5268 gnd.n3865 9.3005
R11901 gnd.n5265 gnd.n3866 9.3005
R11902 gnd.n5264 gnd.n3867 9.3005
R11903 gnd.n5261 gnd.n3868 9.3005
R11904 gnd.n5260 gnd.n3869 9.3005
R11905 gnd.n5257 gnd.n3870 9.3005
R11906 gnd.n5256 gnd.n3871 9.3005
R11907 gnd.n5253 gnd.n3872 9.3005
R11908 gnd.n5252 gnd.n3873 9.3005
R11909 gnd.n5249 gnd.n3874 9.3005
R11910 gnd.n5248 gnd.n3875 9.3005
R11911 gnd.n5245 gnd.n3876 9.3005
R11912 gnd.n5244 gnd.n3877 9.3005
R11913 gnd.n5241 gnd.n3878 9.3005
R11914 gnd.n5240 gnd.n3879 9.3005
R11915 gnd.n5237 gnd.n3880 9.3005
R11916 gnd.n5236 gnd.n3881 9.3005
R11917 gnd.n5233 gnd.n3882 9.3005
R11918 gnd.n5232 gnd.n3883 9.3005
R11919 gnd.n5229 gnd.n3887 9.3005
R11920 gnd.n5228 gnd.n3888 9.3005
R11921 gnd.n5225 gnd.n3889 9.3005
R11922 gnd.n5224 gnd.n3890 9.3005
R11923 gnd.n5275 gnd.n5274 9.3005
R11924 gnd.n4726 gnd.n4710 9.3005
R11925 gnd.n4725 gnd.n4711 9.3005
R11926 gnd.n4724 gnd.n4712 9.3005
R11927 gnd.n4722 gnd.n4713 9.3005
R11928 gnd.n4721 gnd.n4714 9.3005
R11929 gnd.n4719 gnd.n4715 9.3005
R11930 gnd.n4718 gnd.n4716 9.3005
R11931 gnd.n3996 gnd.n3995 9.3005
R11932 gnd.n4795 gnd.n4794 9.3005
R11933 gnd.n4796 gnd.n3994 9.3005
R11934 gnd.n4813 gnd.n4797 9.3005
R11935 gnd.n4812 gnd.n4798 9.3005
R11936 gnd.n4811 gnd.n4799 9.3005
R11937 gnd.n4809 gnd.n4800 9.3005
R11938 gnd.n4808 gnd.n4801 9.3005
R11939 gnd.n4806 gnd.n4802 9.3005
R11940 gnd.n4805 gnd.n4803 9.3005
R11941 gnd.n3940 gnd.n3939 9.3005
R11942 gnd.n4880 gnd.n4879 9.3005
R11943 gnd.n4881 gnd.n3938 9.3005
R11944 gnd.n4902 gnd.n4882 9.3005
R11945 gnd.n4901 gnd.n4883 9.3005
R11946 gnd.n4900 gnd.n4884 9.3005
R11947 gnd.n4897 gnd.n4885 9.3005
R11948 gnd.n4896 gnd.n4886 9.3005
R11949 gnd.n4894 gnd.n4887 9.3005
R11950 gnd.n4893 gnd.n4888 9.3005
R11951 gnd.n4891 gnd.n4890 9.3005
R11952 gnd.n4889 gnd.n3892 9.3005
R11953 gnd.n4467 gnd.n4466 9.3005
R11954 gnd.n4357 gnd.n4356 9.3005
R11955 gnd.n4481 gnd.n4480 9.3005
R11956 gnd.n4482 gnd.n4355 9.3005
R11957 gnd.n4484 gnd.n4483 9.3005
R11958 gnd.n4345 gnd.n4344 9.3005
R11959 gnd.n4497 gnd.n4496 9.3005
R11960 gnd.n4498 gnd.n4343 9.3005
R11961 gnd.n4530 gnd.n4499 9.3005
R11962 gnd.n4529 gnd.n4500 9.3005
R11963 gnd.n4528 gnd.n4501 9.3005
R11964 gnd.n4527 gnd.n4502 9.3005
R11965 gnd.n4524 gnd.n4503 9.3005
R11966 gnd.n4523 gnd.n4504 9.3005
R11967 gnd.n4522 gnd.n4505 9.3005
R11968 gnd.n4520 gnd.n4506 9.3005
R11969 gnd.n4519 gnd.n4507 9.3005
R11970 gnd.n4516 gnd.n4508 9.3005
R11971 gnd.n4515 gnd.n4509 9.3005
R11972 gnd.n4514 gnd.n4510 9.3005
R11973 gnd.n4512 gnd.n4511 9.3005
R11974 gnd.n4211 gnd.n4210 9.3005
R11975 gnd.n4628 gnd.n4627 9.3005
R11976 gnd.n4629 gnd.n4209 9.3005
R11977 gnd.n4633 gnd.n4630 9.3005
R11978 gnd.n4632 gnd.n4631 9.3005
R11979 gnd.n4133 gnd.n4132 9.3005
R11980 gnd.n4708 gnd.n4707 9.3005
R11981 gnd.n4465 gnd.n4366 9.3005
R11982 gnd.n4368 gnd.n4367 9.3005
R11983 gnd.n4412 gnd.n4410 9.3005
R11984 gnd.n4413 gnd.n4409 9.3005
R11985 gnd.n4416 gnd.n4405 9.3005
R11986 gnd.n4417 gnd.n4404 9.3005
R11987 gnd.n4420 gnd.n4403 9.3005
R11988 gnd.n4421 gnd.n4402 9.3005
R11989 gnd.n4424 gnd.n4401 9.3005
R11990 gnd.n4425 gnd.n4400 9.3005
R11991 gnd.n4428 gnd.n4399 9.3005
R11992 gnd.n4429 gnd.n4398 9.3005
R11993 gnd.n4432 gnd.n4397 9.3005
R11994 gnd.n4433 gnd.n4396 9.3005
R11995 gnd.n4436 gnd.n4395 9.3005
R11996 gnd.n4437 gnd.n4394 9.3005
R11997 gnd.n4440 gnd.n4393 9.3005
R11998 gnd.n4441 gnd.n4392 9.3005
R11999 gnd.n4444 gnd.n4391 9.3005
R12000 gnd.n4445 gnd.n4390 9.3005
R12001 gnd.n4448 gnd.n4389 9.3005
R12002 gnd.n4449 gnd.n4388 9.3005
R12003 gnd.n4452 gnd.n4387 9.3005
R12004 gnd.n4454 gnd.n4386 9.3005
R12005 gnd.n4455 gnd.n4385 9.3005
R12006 gnd.n4456 gnd.n4384 9.3005
R12007 gnd.n4457 gnd.n4383 9.3005
R12008 gnd.n4464 gnd.n4463 9.3005
R12009 gnd.n4473 gnd.n4472 9.3005
R12010 gnd.n4474 gnd.n4360 9.3005
R12011 gnd.n4476 gnd.n4475 9.3005
R12012 gnd.n4351 gnd.n4350 9.3005
R12013 gnd.n4489 gnd.n4488 9.3005
R12014 gnd.n4490 gnd.n4349 9.3005
R12015 gnd.n4492 gnd.n4491 9.3005
R12016 gnd.n4338 gnd.n4337 9.3005
R12017 gnd.n4535 gnd.n4534 9.3005
R12018 gnd.n4536 gnd.n4292 9.3005
R12019 gnd.n4540 gnd.n4538 9.3005
R12020 gnd.n4539 gnd.n4271 9.3005
R12021 gnd.n4558 gnd.n4270 9.3005
R12022 gnd.n4561 gnd.n4560 9.3005
R12023 gnd.n4264 gnd.n4263 9.3005
R12024 gnd.n4572 gnd.n4570 9.3005
R12025 gnd.n4571 gnd.n4245 9.3005
R12026 gnd.n4589 gnd.n4244 9.3005
R12027 gnd.n4592 gnd.n4591 9.3005
R12028 gnd.n4239 gnd.n4234 9.3005
R12029 gnd.n4602 gnd.n4601 9.3005
R12030 gnd.n4237 gnd.n4217 9.3005
R12031 gnd.n4623 gnd.n4218 9.3005
R12032 gnd.n4622 gnd.n4621 9.3005
R12033 gnd.n4220 gnd.n4196 9.3005
R12034 gnd.n4654 gnd.n4653 9.3005
R12035 gnd.n4656 gnd.n4141 9.3005
R12036 gnd.n4703 gnd.n4142 9.3005
R12037 gnd.n4702 gnd.n4143 9.3005
R12038 gnd.n4701 gnd.n4144 9.3005
R12039 gnd.n4667 gnd.n4145 9.3005
R12040 gnd.n4669 gnd.n4163 9.3005
R12041 gnd.n4689 gnd.n4164 9.3005
R12042 gnd.n4688 gnd.n4165 9.3005
R12043 gnd.n4687 gnd.n4166 9.3005
R12044 gnd.n4678 gnd.n4167 9.3005
R12045 gnd.n4679 gnd.n4034 9.3005
R12046 gnd.n4745 gnd.n4744 9.3005
R12047 gnd.n4746 gnd.n4027 9.3005
R12048 gnd.n4756 gnd.n4755 9.3005
R12049 gnd.n4758 gnd.n4023 9.3005
R12050 gnd.n4768 gnd.n4024 9.3005
R12051 gnd.n4767 gnd.n4766 9.3005
R12052 gnd.n4764 gnd.n4002 9.3005
R12053 gnd.n4790 gnd.n4003 9.3005
R12054 gnd.n4789 gnd.n4788 9.3005
R12055 gnd.n4005 gnd.n3979 9.3005
R12056 gnd.n4830 gnd.n4829 9.3005
R12057 gnd.n4831 gnd.n3972 9.3005
R12058 gnd.n4841 gnd.n4840 9.3005
R12059 gnd.n4843 gnd.n3968 9.3005
R12060 gnd.n4853 gnd.n3969 9.3005
R12061 gnd.n4852 gnd.n4851 9.3005
R12062 gnd.n4849 gnd.n3947 9.3005
R12063 gnd.n4875 gnd.n3948 9.3005
R12064 gnd.n4874 gnd.n4873 9.3005
R12065 gnd.n3950 gnd.n3925 9.3005
R12066 gnd.n4919 gnd.n4918 9.3005
R12067 gnd.n4920 gnd.n3918 9.3005
R12068 gnd.n4930 gnd.n4929 9.3005
R12069 gnd.n5188 gnd.n3914 9.3005
R12070 gnd.n5196 gnd.n3915 9.3005
R12071 gnd.n5195 gnd.n5194 9.3005
R12072 gnd.n3896 gnd.n3895 9.3005
R12073 gnd.n5219 gnd.n5218 9.3005
R12074 gnd.n4362 gnd.n4361 9.3005
R12075 gnd.n2943 gnd.n2942 9.3005
R12076 gnd.n2941 gnd.n1936 9.3005
R12077 gnd.n1941 gnd.n1937 9.3005
R12078 gnd.n2935 gnd.n1942 9.3005
R12079 gnd.n2934 gnd.n1943 9.3005
R12080 gnd.n2933 gnd.n1944 9.3005
R12081 gnd.n1949 gnd.n1945 9.3005
R12082 gnd.n2927 gnd.n1950 9.3005
R12083 gnd.n2926 gnd.n1951 9.3005
R12084 gnd.n2925 gnd.n1952 9.3005
R12085 gnd.n1957 gnd.n1953 9.3005
R12086 gnd.n2919 gnd.n1958 9.3005
R12087 gnd.n2918 gnd.n1959 9.3005
R12088 gnd.n2917 gnd.n1960 9.3005
R12089 gnd.n1965 gnd.n1961 9.3005
R12090 gnd.n2911 gnd.n1966 9.3005
R12091 gnd.n2910 gnd.n1967 9.3005
R12092 gnd.n2909 gnd.n1968 9.3005
R12093 gnd.n1973 gnd.n1969 9.3005
R12094 gnd.n2903 gnd.n1974 9.3005
R12095 gnd.n2902 gnd.n1975 9.3005
R12096 gnd.n2901 gnd.n1976 9.3005
R12097 gnd.n1981 gnd.n1977 9.3005
R12098 gnd.n2895 gnd.n1982 9.3005
R12099 gnd.n2894 gnd.n1983 9.3005
R12100 gnd.n2893 gnd.n1984 9.3005
R12101 gnd.n1989 gnd.n1985 9.3005
R12102 gnd.n2887 gnd.n1990 9.3005
R12103 gnd.n2886 gnd.n1991 9.3005
R12104 gnd.n2885 gnd.n1992 9.3005
R12105 gnd.n1997 gnd.n1993 9.3005
R12106 gnd.n2879 gnd.n1998 9.3005
R12107 gnd.n2878 gnd.n1999 9.3005
R12108 gnd.n2877 gnd.n2000 9.3005
R12109 gnd.n2005 gnd.n2001 9.3005
R12110 gnd.n2871 gnd.n2006 9.3005
R12111 gnd.n2870 gnd.n2007 9.3005
R12112 gnd.n2869 gnd.n2008 9.3005
R12113 gnd.n2013 gnd.n2009 9.3005
R12114 gnd.n2863 gnd.n2014 9.3005
R12115 gnd.n2862 gnd.n2015 9.3005
R12116 gnd.n2861 gnd.n2016 9.3005
R12117 gnd.n2021 gnd.n2017 9.3005
R12118 gnd.n2855 gnd.n2022 9.3005
R12119 gnd.n2854 gnd.n2023 9.3005
R12120 gnd.n2853 gnd.n2024 9.3005
R12121 gnd.n2029 gnd.n2025 9.3005
R12122 gnd.n2847 gnd.n2030 9.3005
R12123 gnd.n2846 gnd.n2031 9.3005
R12124 gnd.n2845 gnd.n2032 9.3005
R12125 gnd.n2037 gnd.n2033 9.3005
R12126 gnd.n2839 gnd.n2038 9.3005
R12127 gnd.n2838 gnd.n2039 9.3005
R12128 gnd.n2837 gnd.n2040 9.3005
R12129 gnd.n2045 gnd.n2041 9.3005
R12130 gnd.n2831 gnd.n2046 9.3005
R12131 gnd.n2830 gnd.n2047 9.3005
R12132 gnd.n2829 gnd.n2048 9.3005
R12133 gnd.n2053 gnd.n2049 9.3005
R12134 gnd.n2823 gnd.n2054 9.3005
R12135 gnd.n2822 gnd.n2055 9.3005
R12136 gnd.n2821 gnd.n2056 9.3005
R12137 gnd.n2061 gnd.n2057 9.3005
R12138 gnd.n2815 gnd.n2062 9.3005
R12139 gnd.n2814 gnd.n2063 9.3005
R12140 gnd.n2813 gnd.n2064 9.3005
R12141 gnd.n2069 gnd.n2065 9.3005
R12142 gnd.n2807 gnd.n2070 9.3005
R12143 gnd.n2806 gnd.n2071 9.3005
R12144 gnd.n2805 gnd.n2072 9.3005
R12145 gnd.n2077 gnd.n2073 9.3005
R12146 gnd.n2799 gnd.n2078 9.3005
R12147 gnd.n2798 gnd.n2079 9.3005
R12148 gnd.n2797 gnd.n2080 9.3005
R12149 gnd.n2085 gnd.n2081 9.3005
R12150 gnd.n2791 gnd.n2086 9.3005
R12151 gnd.n2790 gnd.n2087 9.3005
R12152 gnd.n2789 gnd.n2088 9.3005
R12153 gnd.n2093 gnd.n2089 9.3005
R12154 gnd.n2783 gnd.n2094 9.3005
R12155 gnd.n2782 gnd.n2095 9.3005
R12156 gnd.n2781 gnd.n2096 9.3005
R12157 gnd.n2101 gnd.n2097 9.3005
R12158 gnd.n2775 gnd.n2102 9.3005
R12159 gnd.n2774 gnd.n2103 9.3005
R12160 gnd.n2773 gnd.n2104 9.3005
R12161 gnd.n2109 gnd.n2105 9.3005
R12162 gnd.n2767 gnd.n2110 9.3005
R12163 gnd.n2766 gnd.n2111 9.3005
R12164 gnd.n2765 gnd.n2112 9.3005
R12165 gnd.n2117 gnd.n2113 9.3005
R12166 gnd.n2759 gnd.n2118 9.3005
R12167 gnd.n2758 gnd.n2119 9.3005
R12168 gnd.n2757 gnd.n2120 9.3005
R12169 gnd.n2125 gnd.n2121 9.3005
R12170 gnd.n2751 gnd.n2126 9.3005
R12171 gnd.n2750 gnd.n2127 9.3005
R12172 gnd.n2749 gnd.n2128 9.3005
R12173 gnd.n2133 gnd.n2129 9.3005
R12174 gnd.n2743 gnd.n2134 9.3005
R12175 gnd.n2742 gnd.n2135 9.3005
R12176 gnd.n2741 gnd.n2136 9.3005
R12177 gnd.n2141 gnd.n2137 9.3005
R12178 gnd.n2735 gnd.n2142 9.3005
R12179 gnd.n2734 gnd.n2143 9.3005
R12180 gnd.n2733 gnd.n2144 9.3005
R12181 gnd.n2149 gnd.n2145 9.3005
R12182 gnd.n2727 gnd.n2150 9.3005
R12183 gnd.n2726 gnd.n2151 9.3005
R12184 gnd.n2725 gnd.n2152 9.3005
R12185 gnd.n2157 gnd.n2153 9.3005
R12186 gnd.n2719 gnd.n2158 9.3005
R12187 gnd.n2718 gnd.n2159 9.3005
R12188 gnd.n2717 gnd.n2160 9.3005
R12189 gnd.n2165 gnd.n2161 9.3005
R12190 gnd.n2711 gnd.n2166 9.3005
R12191 gnd.n2710 gnd.n2167 9.3005
R12192 gnd.n2709 gnd.n2168 9.3005
R12193 gnd.n2173 gnd.n2169 9.3005
R12194 gnd.n2703 gnd.n2174 9.3005
R12195 gnd.n2702 gnd.n2175 9.3005
R12196 gnd.n2701 gnd.n2176 9.3005
R12197 gnd.n2181 gnd.n2177 9.3005
R12198 gnd.n2695 gnd.n2182 9.3005
R12199 gnd.n2694 gnd.n2183 9.3005
R12200 gnd.n2693 gnd.n2184 9.3005
R12201 gnd.n2189 gnd.n2185 9.3005
R12202 gnd.n2687 gnd.n2190 9.3005
R12203 gnd.n2686 gnd.n2191 9.3005
R12204 gnd.n2685 gnd.n2192 9.3005
R12205 gnd.n2197 gnd.n2193 9.3005
R12206 gnd.n2679 gnd.n2198 9.3005
R12207 gnd.n2678 gnd.n2199 9.3005
R12208 gnd.n2677 gnd.n2200 9.3005
R12209 gnd.n2205 gnd.n2201 9.3005
R12210 gnd.n2671 gnd.n2206 9.3005
R12211 gnd.n2670 gnd.n2207 9.3005
R12212 gnd.n2669 gnd.n2208 9.3005
R12213 gnd.n2213 gnd.n2209 9.3005
R12214 gnd.n2663 gnd.n2214 9.3005
R12215 gnd.n2662 gnd.n2215 9.3005
R12216 gnd.n2661 gnd.n2216 9.3005
R12217 gnd.n2221 gnd.n2217 9.3005
R12218 gnd.n2655 gnd.n2222 9.3005
R12219 gnd.n2654 gnd.n2223 9.3005
R12220 gnd.n2653 gnd.n2224 9.3005
R12221 gnd.n2229 gnd.n2225 9.3005
R12222 gnd.n2647 gnd.n2230 9.3005
R12223 gnd.n2646 gnd.n2231 9.3005
R12224 gnd.n2645 gnd.n2232 9.3005
R12225 gnd.n2237 gnd.n2233 9.3005
R12226 gnd.n2639 gnd.n2238 9.3005
R12227 gnd.n2638 gnd.n2239 9.3005
R12228 gnd.n2637 gnd.n2240 9.3005
R12229 gnd.n2245 gnd.n2241 9.3005
R12230 gnd.n2631 gnd.n2246 9.3005
R12231 gnd.n2630 gnd.n2247 9.3005
R12232 gnd.n2629 gnd.n2248 9.3005
R12233 gnd.n2253 gnd.n2249 9.3005
R12234 gnd.n2623 gnd.n2254 9.3005
R12235 gnd.n2622 gnd.n2255 9.3005
R12236 gnd.n2621 gnd.n2256 9.3005
R12237 gnd.n2261 gnd.n2257 9.3005
R12238 gnd.n2615 gnd.n2262 9.3005
R12239 gnd.n2614 gnd.n2263 9.3005
R12240 gnd.n2613 gnd.n2264 9.3005
R12241 gnd.n2269 gnd.n2265 9.3005
R12242 gnd.n2607 gnd.n2606 9.3005
R12243 gnd.n2603 gnd.n2270 9.3005
R12244 gnd.n2602 gnd.n2272 9.3005
R12245 gnd.n2278 gnd.n2273 9.3005
R12246 gnd.n2596 gnd.n2279 9.3005
R12247 gnd.n2595 gnd.n2280 9.3005
R12248 gnd.n2594 gnd.n2281 9.3005
R12249 gnd.n2286 gnd.n2282 9.3005
R12250 gnd.n2588 gnd.n2287 9.3005
R12251 gnd.n2587 gnd.n2288 9.3005
R12252 gnd.n2586 gnd.n2289 9.3005
R12253 gnd.n2294 gnd.n2290 9.3005
R12254 gnd.n2580 gnd.n2295 9.3005
R12255 gnd.n2579 gnd.n2296 9.3005
R12256 gnd.n2578 gnd.n2297 9.3005
R12257 gnd.n2302 gnd.n2298 9.3005
R12258 gnd.n2572 gnd.n2303 9.3005
R12259 gnd.n2571 gnd.n2304 9.3005
R12260 gnd.n2570 gnd.n2305 9.3005
R12261 gnd.n2310 gnd.n2306 9.3005
R12262 gnd.n2564 gnd.n2311 9.3005
R12263 gnd.n2563 gnd.n2312 9.3005
R12264 gnd.n2562 gnd.n2313 9.3005
R12265 gnd.n2318 gnd.n2314 9.3005
R12266 gnd.n2556 gnd.n2319 9.3005
R12267 gnd.n2555 gnd.n2320 9.3005
R12268 gnd.n2554 gnd.n2321 9.3005
R12269 gnd.n2326 gnd.n2322 9.3005
R12270 gnd.n2548 gnd.n2327 9.3005
R12271 gnd.n2547 gnd.n2328 9.3005
R12272 gnd.n2546 gnd.n2329 9.3005
R12273 gnd.n2334 gnd.n2330 9.3005
R12274 gnd.n2540 gnd.n2335 9.3005
R12275 gnd.n2539 gnd.n2336 9.3005
R12276 gnd.n2538 gnd.n2337 9.3005
R12277 gnd.n2342 gnd.n2338 9.3005
R12278 gnd.n2532 gnd.n2343 9.3005
R12279 gnd.n2531 gnd.n2344 9.3005
R12280 gnd.n2530 gnd.n2345 9.3005
R12281 gnd.n2350 gnd.n2346 9.3005
R12282 gnd.n2524 gnd.n2351 9.3005
R12283 gnd.n2523 gnd.n2352 9.3005
R12284 gnd.n2522 gnd.n2353 9.3005
R12285 gnd.n2358 gnd.n2354 9.3005
R12286 gnd.n2516 gnd.n2359 9.3005
R12287 gnd.n2515 gnd.n2360 9.3005
R12288 gnd.n2514 gnd.n2361 9.3005
R12289 gnd.n2366 gnd.n2362 9.3005
R12290 gnd.n2508 gnd.n2367 9.3005
R12291 gnd.n2507 gnd.n2368 9.3005
R12292 gnd.n2506 gnd.n2369 9.3005
R12293 gnd.n2374 gnd.n2370 9.3005
R12294 gnd.n2500 gnd.n2375 9.3005
R12295 gnd.n2499 gnd.n2376 9.3005
R12296 gnd.n2498 gnd.n2377 9.3005
R12297 gnd.n2382 gnd.n2378 9.3005
R12298 gnd.n2492 gnd.n2383 9.3005
R12299 gnd.n2491 gnd.n2384 9.3005
R12300 gnd.n2490 gnd.n2385 9.3005
R12301 gnd.n2390 gnd.n2386 9.3005
R12302 gnd.n2484 gnd.n2391 9.3005
R12303 gnd.n2483 gnd.n2392 9.3005
R12304 gnd.n2482 gnd.n2393 9.3005
R12305 gnd.n2398 gnd.n2394 9.3005
R12306 gnd.n2476 gnd.n2399 9.3005
R12307 gnd.n2475 gnd.n2400 9.3005
R12308 gnd.n2474 gnd.n2401 9.3005
R12309 gnd.n2406 gnd.n2402 9.3005
R12310 gnd.n2468 gnd.n2407 9.3005
R12311 gnd.n2467 gnd.n2408 9.3005
R12312 gnd.n2466 gnd.n2409 9.3005
R12313 gnd.n2414 gnd.n2410 9.3005
R12314 gnd.n2460 gnd.n2415 9.3005
R12315 gnd.n2459 gnd.n2416 9.3005
R12316 gnd.n2458 gnd.n2417 9.3005
R12317 gnd.n2422 gnd.n2418 9.3005
R12318 gnd.n2452 gnd.n2423 9.3005
R12319 gnd.n2451 gnd.n2424 9.3005
R12320 gnd.n2450 gnd.n2425 9.3005
R12321 gnd.n2430 gnd.n2426 9.3005
R12322 gnd.n2444 gnd.n2431 9.3005
R12323 gnd.n2443 gnd.n2432 9.3005
R12324 gnd.n2442 gnd.n2433 9.3005
R12325 gnd.n2437 gnd.n2434 9.3005
R12326 gnd.n2436 gnd.n2435 9.3005
R12327 gnd.n2605 gnd.n2604 9.3005
R12328 gnd.n7981 gnd.n7980 9.3005
R12329 gnd.n7979 gnd.n101 9.3005
R12330 gnd.n7619 gnd.n103 9.3005
R12331 gnd.n7622 gnd.n7621 9.3005
R12332 gnd.n7623 gnd.n7618 9.3005
R12333 gnd.n7626 gnd.n7624 9.3005
R12334 gnd.n7627 gnd.n7617 9.3005
R12335 gnd.n7630 gnd.n7629 9.3005
R12336 gnd.n7631 gnd.n7616 9.3005
R12337 gnd.n7634 gnd.n7632 9.3005
R12338 gnd.n7635 gnd.n7615 9.3005
R12339 gnd.n7638 gnd.n7637 9.3005
R12340 gnd.n7639 gnd.n7614 9.3005
R12341 gnd.n7642 gnd.n7640 9.3005
R12342 gnd.n7643 gnd.n7613 9.3005
R12343 gnd.n7646 gnd.n7645 9.3005
R12344 gnd.n7647 gnd.n7612 9.3005
R12345 gnd.n7650 gnd.n7648 9.3005
R12346 gnd.n7651 gnd.n7611 9.3005
R12347 gnd.n7654 gnd.n7653 9.3005
R12348 gnd.n7655 gnd.n7610 9.3005
R12349 gnd.n7739 gnd.n7656 9.3005
R12350 gnd.n7738 gnd.n7657 9.3005
R12351 gnd.n7737 gnd.n7658 9.3005
R12352 gnd.n7735 gnd.n7659 9.3005
R12353 gnd.n7734 gnd.n7660 9.3005
R12354 gnd.n7732 gnd.n7661 9.3005
R12355 gnd.n7731 gnd.n7662 9.3005
R12356 gnd.n7729 gnd.n7663 9.3005
R12357 gnd.n7728 gnd.n7664 9.3005
R12358 gnd.n7726 gnd.n7665 9.3005
R12359 gnd.n7725 gnd.n7666 9.3005
R12360 gnd.n7680 gnd.n7679 9.3005
R12361 gnd.n7682 gnd.n7681 9.3005
R12362 gnd.n7685 gnd.n7676 9.3005
R12363 gnd.n7689 gnd.n7688 9.3005
R12364 gnd.n7690 gnd.n7675 9.3005
R12365 gnd.n7692 gnd.n7691 9.3005
R12366 gnd.n7695 gnd.n7674 9.3005
R12367 gnd.n7699 gnd.n7698 9.3005
R12368 gnd.n7700 gnd.n7673 9.3005
R12369 gnd.n7702 gnd.n7701 9.3005
R12370 gnd.n7705 gnd.n7672 9.3005
R12371 gnd.n7709 gnd.n7708 9.3005
R12372 gnd.n7710 gnd.n7671 9.3005
R12373 gnd.n7712 gnd.n7711 9.3005
R12374 gnd.n7715 gnd.n7670 9.3005
R12375 gnd.n7719 gnd.n7718 9.3005
R12376 gnd.n7720 gnd.n7669 9.3005
R12377 gnd.n7722 gnd.n7721 9.3005
R12378 gnd.n7677 gnd.n352 9.3005
R12379 gnd.n253 gnd.n252 9.3005
R12380 gnd.n7880 gnd.n294 9.3005
R12381 gnd.n7879 gnd.n295 9.3005
R12382 gnd.n7878 gnd.n296 9.3005
R12383 gnd.n7875 gnd.n297 9.3005
R12384 gnd.n7874 gnd.n298 9.3005
R12385 gnd.n7871 gnd.n299 9.3005
R12386 gnd.n7870 gnd.n300 9.3005
R12387 gnd.n7867 gnd.n301 9.3005
R12388 gnd.n7866 gnd.n302 9.3005
R12389 gnd.n7863 gnd.n303 9.3005
R12390 gnd.n7862 gnd.n304 9.3005
R12391 gnd.n7859 gnd.n305 9.3005
R12392 gnd.n7858 gnd.n306 9.3005
R12393 gnd.n7855 gnd.n307 9.3005
R12394 gnd.n7854 gnd.n308 9.3005
R12395 gnd.n7851 gnd.n309 9.3005
R12396 gnd.n7847 gnd.n310 9.3005
R12397 gnd.n7844 gnd.n311 9.3005
R12398 gnd.n7843 gnd.n312 9.3005
R12399 gnd.n7840 gnd.n313 9.3005
R12400 gnd.n7839 gnd.n314 9.3005
R12401 gnd.n7836 gnd.n315 9.3005
R12402 gnd.n7835 gnd.n316 9.3005
R12403 gnd.n7832 gnd.n317 9.3005
R12404 gnd.n7831 gnd.n318 9.3005
R12405 gnd.n7828 gnd.n319 9.3005
R12406 gnd.n7827 gnd.n320 9.3005
R12407 gnd.n7824 gnd.n321 9.3005
R12408 gnd.n7823 gnd.n322 9.3005
R12409 gnd.n7820 gnd.n323 9.3005
R12410 gnd.n7819 gnd.n324 9.3005
R12411 gnd.n7816 gnd.n325 9.3005
R12412 gnd.n7815 gnd.n326 9.3005
R12413 gnd.n7812 gnd.n327 9.3005
R12414 gnd.n7811 gnd.n328 9.3005
R12415 gnd.n7808 gnd.n7807 9.3005
R12416 gnd.n7806 gnd.n329 9.3005
R12417 gnd.n7805 gnd.n7804 9.3005
R12418 gnd.n7801 gnd.n332 9.3005
R12419 gnd.n7798 gnd.n333 9.3005
R12420 gnd.n7797 gnd.n334 9.3005
R12421 gnd.n7794 gnd.n335 9.3005
R12422 gnd.n7793 gnd.n336 9.3005
R12423 gnd.n7790 gnd.n337 9.3005
R12424 gnd.n7789 gnd.n338 9.3005
R12425 gnd.n7786 gnd.n339 9.3005
R12426 gnd.n7785 gnd.n340 9.3005
R12427 gnd.n7782 gnd.n341 9.3005
R12428 gnd.n7781 gnd.n342 9.3005
R12429 gnd.n7778 gnd.n343 9.3005
R12430 gnd.n7777 gnd.n344 9.3005
R12431 gnd.n7774 gnd.n345 9.3005
R12432 gnd.n7773 gnd.n346 9.3005
R12433 gnd.n7770 gnd.n347 9.3005
R12434 gnd.n7769 gnd.n348 9.3005
R12435 gnd.n7766 gnd.n7765 9.3005
R12436 gnd.n7764 gnd.n349 9.3005
R12437 gnd.n7886 gnd.n7885 9.3005
R12438 gnd.n7307 gnd.n7306 9.3005
R12439 gnd.n563 gnd.n558 9.3005
R12440 gnd.n562 gnd.n561 9.3005
R12441 gnd.n534 gnd.n528 9.3005
R12442 gnd.n7350 gnd.n529 9.3005
R12443 gnd.n7349 gnd.n530 9.3005
R12444 gnd.n7348 gnd.n531 9.3005
R12445 gnd.n7347 gnd.n7345 9.3005
R12446 gnd.n532 gnd.n492 9.3005
R12447 gnd.n7399 gnd.n493 9.3005
R12448 gnd.n7398 gnd.n494 9.3005
R12449 gnd.n7397 gnd.n495 9.3005
R12450 gnd.n7396 gnd.n496 9.3005
R12451 gnd.n468 gnd.n462 9.3005
R12452 gnd.n7436 gnd.n463 9.3005
R12453 gnd.n7435 gnd.n464 9.3005
R12454 gnd.n7434 gnd.n465 9.3005
R12455 gnd.n7433 gnd.n7431 9.3005
R12456 gnd.n466 gnd.n426 9.3005
R12457 gnd.n7484 gnd.n427 9.3005
R12458 gnd.n7483 gnd.n428 9.3005
R12459 gnd.n7482 gnd.n429 9.3005
R12460 gnd.n7481 gnd.n7479 9.3005
R12461 gnd.n430 gnd.n388 9.3005
R12462 gnd.n7534 gnd.n389 9.3005
R12463 gnd.n7533 gnd.n390 9.3005
R12464 gnd.n7532 gnd.n391 9.3005
R12465 gnd.n7530 gnd.n392 9.3005
R12466 gnd.n7529 gnd.n7527 9.3005
R12467 gnd.n362 gnd.n361 9.3005
R12468 gnd.n7564 gnd.n7563 9.3005
R12469 gnd.n7565 gnd.n355 9.3005
R12470 gnd.n7572 gnd.n356 9.3005
R12471 gnd.n7573 gnd.n354 9.3005
R12472 gnd.n7576 gnd.n7575 9.3005
R12473 gnd.n7577 gnd.n127 9.3005
R12474 gnd.n7967 gnd.n128 9.3005
R12475 gnd.n7966 gnd.n129 9.3005
R12476 gnd.n7965 gnd.n130 9.3005
R12477 gnd.n7585 gnd.n131 9.3005
R12478 gnd.n7955 gnd.n145 9.3005
R12479 gnd.n7954 gnd.n146 9.3005
R12480 gnd.n7953 gnd.n147 9.3005
R12481 gnd.n7592 gnd.n148 9.3005
R12482 gnd.n7943 gnd.n165 9.3005
R12483 gnd.n7942 gnd.n166 9.3005
R12484 gnd.n7941 gnd.n167 9.3005
R12485 gnd.n7599 gnd.n168 9.3005
R12486 gnd.n7931 gnd.n183 9.3005
R12487 gnd.n7930 gnd.n184 9.3005
R12488 gnd.n7929 gnd.n185 9.3005
R12489 gnd.n7606 gnd.n186 9.3005
R12490 gnd.n7919 gnd.n203 9.3005
R12491 gnd.n7918 gnd.n204 9.3005
R12492 gnd.n7917 gnd.n205 9.3005
R12493 gnd.n7745 gnd.n206 9.3005
R12494 gnd.n7907 gnd.n221 9.3005
R12495 gnd.n7906 gnd.n222 9.3005
R12496 gnd.n7905 gnd.n223 9.3005
R12497 gnd.n7752 gnd.n224 9.3005
R12498 gnd.n7895 gnd.n241 9.3005
R12499 gnd.n7894 gnd.n242 9.3005
R12500 gnd.n7893 gnd.n243 9.3005
R12501 gnd.n7762 gnd.n244 9.3005
R12502 gnd.n7308 gnd.n557 9.3005
R12503 gnd.n7306 gnd.n7305 9.3005
R12504 gnd.n7304 gnd.n563 9.3005
R12505 gnd.n562 gnd.n533 9.3005
R12506 gnd.n7331 gnd.n534 9.3005
R12507 gnd.n7332 gnd.n529 9.3005
R12508 gnd.n7335 gnd.n530 9.3005
R12509 gnd.n7336 gnd.n531 9.3005
R12510 gnd.n7345 gnd.n7344 9.3005
R12511 gnd.n7342 gnd.n532 9.3005
R12512 gnd.n7341 gnd.n493 9.3005
R12513 gnd.n7340 gnd.n494 9.3005
R12514 gnd.n7337 gnd.n495 9.3005
R12515 gnd.n496 gnd.n467 9.3005
R12516 gnd.n7422 gnd.n468 9.3005
R12517 gnd.n7423 gnd.n463 9.3005
R12518 gnd.n7426 gnd.n464 9.3005
R12519 gnd.n7427 gnd.n465 9.3005
R12520 gnd.n7431 gnd.n7430 9.3005
R12521 gnd.n7428 gnd.n466 9.3005
R12522 gnd.n431 gnd.n427 9.3005
R12523 gnd.n7473 gnd.n428 9.3005
R12524 gnd.n7474 gnd.n429 9.3005
R12525 gnd.n7479 gnd.n7478 9.3005
R12526 gnd.n7476 gnd.n430 9.3005
R12527 gnd.n7475 gnd.n389 9.3005
R12528 gnd.n393 gnd.n390 9.3005
R12529 gnd.n7522 gnd.n391 9.3005
R12530 gnd.n7523 gnd.n392 9.3005
R12531 gnd.n7527 gnd.n7526 9.3005
R12532 gnd.n7524 gnd.n361 9.3005
R12533 gnd.n7564 gnd.n360 9.3005
R12534 gnd.n7566 gnd.n7565 9.3005
R12535 gnd.n7568 gnd.n356 9.3005
R12536 gnd.n7567 gnd.n354 9.3005
R12537 gnd.n7576 gnd.n353 9.3005
R12538 gnd.n7580 gnd.n7577 9.3005
R12539 gnd.n7581 gnd.n128 9.3005
R12540 gnd.n7583 gnd.n129 9.3005
R12541 gnd.n7584 gnd.n130 9.3005
R12542 gnd.n7587 gnd.n7585 9.3005
R12543 gnd.n7588 gnd.n145 9.3005
R12544 gnd.n7590 gnd.n146 9.3005
R12545 gnd.n7591 gnd.n147 9.3005
R12546 gnd.n7594 gnd.n7592 9.3005
R12547 gnd.n7595 gnd.n165 9.3005
R12548 gnd.n7597 gnd.n166 9.3005
R12549 gnd.n7598 gnd.n167 9.3005
R12550 gnd.n7601 gnd.n7599 9.3005
R12551 gnd.n7602 gnd.n183 9.3005
R12552 gnd.n7604 gnd.n184 9.3005
R12553 gnd.n7605 gnd.n185 9.3005
R12554 gnd.n7608 gnd.n7606 9.3005
R12555 gnd.n7609 gnd.n203 9.3005
R12556 gnd.n7743 gnd.n204 9.3005
R12557 gnd.n7744 gnd.n205 9.3005
R12558 gnd.n7747 gnd.n7745 9.3005
R12559 gnd.n7748 gnd.n221 9.3005
R12560 gnd.n7750 gnd.n222 9.3005
R12561 gnd.n7751 gnd.n223 9.3005
R12562 gnd.n7754 gnd.n7752 9.3005
R12563 gnd.n7755 gnd.n241 9.3005
R12564 gnd.n7757 gnd.n242 9.3005
R12565 gnd.n7758 gnd.n243 9.3005
R12566 gnd.n7762 gnd.n7761 9.3005
R12567 gnd.n564 gnd.n557 9.3005
R12568 gnd.n7162 gnd.n7161 9.3005
R12569 gnd.n7165 gnd.n672 9.3005
R12570 gnd.n7166 gnd.n671 9.3005
R12571 gnd.n7169 gnd.n670 9.3005
R12572 gnd.n7170 gnd.n669 9.3005
R12573 gnd.n7173 gnd.n668 9.3005
R12574 gnd.n7174 gnd.n667 9.3005
R12575 gnd.n7177 gnd.n666 9.3005
R12576 gnd.n7178 gnd.n665 9.3005
R12577 gnd.n7181 gnd.n664 9.3005
R12578 gnd.n7182 gnd.n663 9.3005
R12579 gnd.n7185 gnd.n662 9.3005
R12580 gnd.n7186 gnd.n661 9.3005
R12581 gnd.n7189 gnd.n660 9.3005
R12582 gnd.n7190 gnd.n659 9.3005
R12583 gnd.n7193 gnd.n658 9.3005
R12584 gnd.n7194 gnd.n657 9.3005
R12585 gnd.n7197 gnd.n656 9.3005
R12586 gnd.n7198 gnd.n655 9.3005
R12587 gnd.n7201 gnd.n654 9.3005
R12588 gnd.n7205 gnd.n650 9.3005
R12589 gnd.n7206 gnd.n649 9.3005
R12590 gnd.n7209 gnd.n648 9.3005
R12591 gnd.n7210 gnd.n647 9.3005
R12592 gnd.n7213 gnd.n646 9.3005
R12593 gnd.n7214 gnd.n645 9.3005
R12594 gnd.n7217 gnd.n644 9.3005
R12595 gnd.n7218 gnd.n643 9.3005
R12596 gnd.n7221 gnd.n642 9.3005
R12597 gnd.n7223 gnd.n638 9.3005
R12598 gnd.n7226 gnd.n637 9.3005
R12599 gnd.n7227 gnd.n636 9.3005
R12600 gnd.n7230 gnd.n635 9.3005
R12601 gnd.n7231 gnd.n634 9.3005
R12602 gnd.n7234 gnd.n633 9.3005
R12603 gnd.n7235 gnd.n632 9.3005
R12604 gnd.n7238 gnd.n631 9.3005
R12605 gnd.n7240 gnd.n628 9.3005
R12606 gnd.n7243 gnd.n627 9.3005
R12607 gnd.n7244 gnd.n626 9.3005
R12608 gnd.n7247 gnd.n625 9.3005
R12609 gnd.n7248 gnd.n624 9.3005
R12610 gnd.n7251 gnd.n623 9.3005
R12611 gnd.n7252 gnd.n622 9.3005
R12612 gnd.n7255 gnd.n621 9.3005
R12613 gnd.n7256 gnd.n620 9.3005
R12614 gnd.n7259 gnd.n619 9.3005
R12615 gnd.n7260 gnd.n618 9.3005
R12616 gnd.n7263 gnd.n617 9.3005
R12617 gnd.n7264 gnd.n616 9.3005
R12618 gnd.n7267 gnd.n615 9.3005
R12619 gnd.n7269 gnd.n614 9.3005
R12620 gnd.n7270 gnd.n613 9.3005
R12621 gnd.n7271 gnd.n612 9.3005
R12622 gnd.n611 gnd.n549 9.3005
R12623 gnd.n7202 gnd.n651 9.3005
R12624 gnd.n7160 gnd.n674 9.3005
R12625 gnd.n7314 gnd.n548 9.3005
R12626 gnd.n7318 gnd.n7315 9.3005
R12627 gnd.n7317 gnd.n7316 9.3005
R12628 gnd.n520 gnd.n519 9.3005
R12629 gnd.n7355 gnd.n7354 9.3005
R12630 gnd.n7356 gnd.n518 9.3005
R12631 gnd.n7360 gnd.n7357 9.3005
R12632 gnd.n7359 gnd.n7358 9.3005
R12633 gnd.n484 gnd.n483 9.3005
R12634 gnd.n7404 gnd.n7403 9.3005
R12635 gnd.n7405 gnd.n482 9.3005
R12636 gnd.n7409 gnd.n7406 9.3005
R12637 gnd.n7408 gnd.n7407 9.3005
R12638 gnd.n454 gnd.n453 9.3005
R12639 gnd.n7441 gnd.n7440 9.3005
R12640 gnd.n7442 gnd.n452 9.3005
R12641 gnd.n7446 gnd.n7443 9.3005
R12642 gnd.n7445 gnd.n7444 9.3005
R12643 gnd.n419 gnd.n418 9.3005
R12644 gnd.n7489 gnd.n7488 9.3005
R12645 gnd.n7490 gnd.n417 9.3005
R12646 gnd.n7495 gnd.n7491 9.3005
R12647 gnd.n7494 gnd.n7493 9.3005
R12648 gnd.n7492 gnd.n380 9.3005
R12649 gnd.n7538 gnd.n381 9.3005
R12650 gnd.n7539 gnd.n113 9.3005
R12651 gnd.n118 gnd.n112 9.3005
R12652 gnd.n7961 gnd.n137 9.3005
R12653 gnd.n7960 gnd.n138 9.3005
R12654 gnd.n7959 gnd.n139 9.3005
R12655 gnd.n154 gnd.n140 9.3005
R12656 gnd.n7949 gnd.n155 9.3005
R12657 gnd.n7948 gnd.n156 9.3005
R12658 gnd.n7947 gnd.n157 9.3005
R12659 gnd.n174 gnd.n158 9.3005
R12660 gnd.n7937 gnd.n175 9.3005
R12661 gnd.n7936 gnd.n176 9.3005
R12662 gnd.n7935 gnd.n177 9.3005
R12663 gnd.n192 gnd.n178 9.3005
R12664 gnd.n7925 gnd.n193 9.3005
R12665 gnd.n7924 gnd.n194 9.3005
R12666 gnd.n7923 gnd.n195 9.3005
R12667 gnd.n212 gnd.n196 9.3005
R12668 gnd.n7913 gnd.n213 9.3005
R12669 gnd.n7912 gnd.n214 9.3005
R12670 gnd.n7911 gnd.n215 9.3005
R12671 gnd.n231 gnd.n216 9.3005
R12672 gnd.n7901 gnd.n232 9.3005
R12673 gnd.n7900 gnd.n233 9.3005
R12674 gnd.n7899 gnd.n234 9.3005
R12675 gnd.n250 gnd.n235 9.3005
R12676 gnd.n7889 gnd.n251 9.3005
R12677 gnd.n7888 gnd.n7887 9.3005
R12678 gnd.n7313 gnd.n7312 9.3005
R12679 gnd.n7972 gnd.n7971 9.3005
R12680 gnd.n3602 gnd.n3601 9.3005
R12681 gnd.n3600 gnd.n3598 9.3005
R12682 gnd.n1755 gnd.n1754 9.3005
R12683 gnd.n5377 gnd.n5376 9.3005
R12684 gnd.n5378 gnd.n1753 9.3005
R12685 gnd.n5382 gnd.n5379 9.3005
R12686 gnd.n5381 gnd.n5380 9.3005
R12687 gnd.n1720 gnd.n1719 9.3005
R12688 gnd.n5427 gnd.n5426 9.3005
R12689 gnd.n5428 gnd.n1718 9.3005
R12690 gnd.n5432 gnd.n5429 9.3005
R12691 gnd.n5431 gnd.n5430 9.3005
R12692 gnd.n1656 gnd.n1655 9.3005
R12693 gnd.n5489 gnd.n5488 9.3005
R12694 gnd.n5490 gnd.n1654 9.3005
R12695 gnd.n5492 gnd.n5491 9.3005
R12696 gnd.n1652 gnd.n1651 9.3005
R12697 gnd.n5497 gnd.n5496 9.3005
R12698 gnd.n5498 gnd.n1650 9.3005
R12699 gnd.n5535 gnd.n5499 9.3005
R12700 gnd.n5534 gnd.n5500 9.3005
R12701 gnd.n5533 gnd.n5501 9.3005
R12702 gnd.n5504 gnd.n5502 9.3005
R12703 gnd.n5529 gnd.n5505 9.3005
R12704 gnd.n5528 gnd.n5506 9.3005
R12705 gnd.n5527 gnd.n5507 9.3005
R12706 gnd.n5510 gnd.n5508 9.3005
R12707 gnd.n5522 gnd.n5511 9.3005
R12708 gnd.n5521 gnd.n5512 9.3005
R12709 gnd.n5520 gnd.n5513 9.3005
R12710 gnd.n5515 gnd.n5514 9.3005
R12711 gnd.n1227 gnd.n1226 9.3005
R12712 gnd.n6167 gnd.n6166 9.3005
R12713 gnd.n6168 gnd.n1225 9.3005
R12714 gnd.n6170 gnd.n6169 9.3005
R12715 gnd.n1214 gnd.n1213 9.3005
R12716 gnd.n6183 gnd.n6182 9.3005
R12717 gnd.n6184 gnd.n1212 9.3005
R12718 gnd.n6186 gnd.n6185 9.3005
R12719 gnd.n1200 gnd.n1199 9.3005
R12720 gnd.n6199 gnd.n6198 9.3005
R12721 gnd.n6200 gnd.n1198 9.3005
R12722 gnd.n6202 gnd.n6201 9.3005
R12723 gnd.n1186 gnd.n1185 9.3005
R12724 gnd.n6215 gnd.n6214 9.3005
R12725 gnd.n6216 gnd.n1184 9.3005
R12726 gnd.n6218 gnd.n6217 9.3005
R12727 gnd.n1171 gnd.n1170 9.3005
R12728 gnd.n6231 gnd.n6230 9.3005
R12729 gnd.n6232 gnd.n1169 9.3005
R12730 gnd.n6234 gnd.n6233 9.3005
R12731 gnd.n1157 gnd.n1156 9.3005
R12732 gnd.n6247 gnd.n6246 9.3005
R12733 gnd.n6248 gnd.n1155 9.3005
R12734 gnd.n6250 gnd.n6249 9.3005
R12735 gnd.n1141 gnd.n1140 9.3005
R12736 gnd.n6263 gnd.n6262 9.3005
R12737 gnd.n6264 gnd.n1139 9.3005
R12738 gnd.n6266 gnd.n6265 9.3005
R12739 gnd.n1127 gnd.n1126 9.3005
R12740 gnd.n6279 gnd.n6278 9.3005
R12741 gnd.n6280 gnd.n1125 9.3005
R12742 gnd.n6282 gnd.n6281 9.3005
R12743 gnd.n1113 gnd.n1112 9.3005
R12744 gnd.n6295 gnd.n6294 9.3005
R12745 gnd.n6296 gnd.n1111 9.3005
R12746 gnd.n6298 gnd.n6297 9.3005
R12747 gnd.n1100 gnd.n1099 9.3005
R12748 gnd.n6311 gnd.n6310 9.3005
R12749 gnd.n6312 gnd.n1098 9.3005
R12750 gnd.n6314 gnd.n6313 9.3005
R12751 gnd.n1086 gnd.n1085 9.3005
R12752 gnd.n6327 gnd.n6326 9.3005
R12753 gnd.n6328 gnd.n1084 9.3005
R12754 gnd.n6330 gnd.n6329 9.3005
R12755 gnd.n1068 gnd.n1067 9.3005
R12756 gnd.n6349 gnd.n6348 9.3005
R12757 gnd.n6350 gnd.n1066 9.3005
R12758 gnd.n6354 gnd.n6351 9.3005
R12759 gnd.n6353 gnd.n6352 9.3005
R12760 gnd.n1030 gnd.n1029 9.3005
R12761 gnd.n6407 gnd.n6406 9.3005
R12762 gnd.n6408 gnd.n1028 9.3005
R12763 gnd.n6412 gnd.n6409 9.3005
R12764 gnd.n6411 gnd.n6410 9.3005
R12765 gnd.n991 gnd.n990 9.3005
R12766 gnd.n6465 gnd.n6464 9.3005
R12767 gnd.n6466 gnd.n989 9.3005
R12768 gnd.n6470 gnd.n6467 9.3005
R12769 gnd.n6469 gnd.n6468 9.3005
R12770 gnd.n923 gnd.n922 9.3005
R12771 gnd.n6903 gnd.n6902 9.3005
R12772 gnd.n6904 gnd.n921 9.3005
R12773 gnd.n6906 gnd.n6905 9.3005
R12774 gnd.n909 gnd.n908 9.3005
R12775 gnd.n6919 gnd.n6918 9.3005
R12776 gnd.n6920 gnd.n907 9.3005
R12777 gnd.n6922 gnd.n6921 9.3005
R12778 gnd.n896 gnd.n895 9.3005
R12779 gnd.n6935 gnd.n6934 9.3005
R12780 gnd.n6936 gnd.n894 9.3005
R12781 gnd.n6938 gnd.n6937 9.3005
R12782 gnd.n882 gnd.n881 9.3005
R12783 gnd.n6951 gnd.n6950 9.3005
R12784 gnd.n6952 gnd.n880 9.3005
R12785 gnd.n6954 gnd.n6953 9.3005
R12786 gnd.n868 gnd.n867 9.3005
R12787 gnd.n6967 gnd.n6966 9.3005
R12788 gnd.n6968 gnd.n866 9.3005
R12789 gnd.n6970 gnd.n6969 9.3005
R12790 gnd.n853 gnd.n852 9.3005
R12791 gnd.n6983 gnd.n6982 9.3005
R12792 gnd.n6984 gnd.n851 9.3005
R12793 gnd.n6986 gnd.n6985 9.3005
R12794 gnd.n838 gnd.n837 9.3005
R12795 gnd.n6999 gnd.n6998 9.3005
R12796 gnd.n7000 gnd.n836 9.3005
R12797 gnd.n7002 gnd.n7001 9.3005
R12798 gnd.n825 gnd.n824 9.3005
R12799 gnd.n7015 gnd.n7014 9.3005
R12800 gnd.n7016 gnd.n823 9.3005
R12801 gnd.n7018 gnd.n7017 9.3005
R12802 gnd.n811 gnd.n810 9.3005
R12803 gnd.n7031 gnd.n7030 9.3005
R12804 gnd.n7032 gnd.n809 9.3005
R12805 gnd.n7034 gnd.n7033 9.3005
R12806 gnd.n797 gnd.n796 9.3005
R12807 gnd.n7047 gnd.n7046 9.3005
R12808 gnd.n7048 gnd.n795 9.3005
R12809 gnd.n7053 gnd.n7049 9.3005
R12810 gnd.n7052 gnd.n7051 9.3005
R12811 gnd.n7050 gnd.n783 9.3005
R12812 gnd.n7066 gnd.n782 9.3005
R12813 gnd.n7068 gnd.n7067 9.3005
R12814 gnd.n7069 gnd.n781 9.3005
R12815 gnd.n7075 gnd.n7070 9.3005
R12816 gnd.n7074 gnd.n7071 9.3005
R12817 gnd.n7073 gnd.n7072 9.3005
R12818 gnd.n569 gnd.n568 9.3005
R12819 gnd.n7279 gnd.n7278 9.3005
R12820 gnd.n7280 gnd.n567 9.3005
R12821 gnd.n7299 gnd.n7281 9.3005
R12822 gnd.n7298 gnd.n7282 9.3005
R12823 gnd.n7297 gnd.n7283 9.3005
R12824 gnd.n7286 gnd.n7284 9.3005
R12825 gnd.n7293 gnd.n7287 9.3005
R12826 gnd.n7292 gnd.n7288 9.3005
R12827 gnd.n7291 gnd.n7290 9.3005
R12828 gnd.n7289 gnd.n503 9.3005
R12829 gnd.n501 gnd.n500 9.3005
R12830 gnd.n7377 gnd.n7376 9.3005
R12831 gnd.n7378 gnd.n499 9.3005
R12832 gnd.n7391 gnd.n7379 9.3005
R12833 gnd.n7390 gnd.n7380 9.3005
R12834 gnd.n7389 gnd.n7381 9.3005
R12835 gnd.n7383 gnd.n7382 9.3005
R12836 gnd.n7385 gnd.n7384 9.3005
R12837 gnd.n436 gnd.n435 9.3005
R12838 gnd.n7461 gnd.n7460 9.3005
R12839 gnd.n7462 gnd.n434 9.3005
R12840 gnd.n7468 gnd.n7463 9.3005
R12841 gnd.n7467 gnd.n7464 9.3005
R12842 gnd.n7466 gnd.n7465 9.3005
R12843 gnd.n401 gnd.n400 9.3005
R12844 gnd.n7513 gnd.n7512 9.3005
R12845 gnd.n7514 gnd.n399 9.3005
R12846 gnd.n7516 gnd.n7515 9.3005
R12847 gnd.n3599 gnd.n3597 9.3005
R12848 gnd.n3541 gnd.n3540 9.3005
R12849 gnd.n3476 gnd.n3414 9.3005
R12850 gnd.n3479 gnd.n3478 9.3005
R12851 gnd.n3480 gnd.n3413 9.3005
R12852 gnd.n3483 gnd.n3481 9.3005
R12853 gnd.n3484 gnd.n3412 9.3005
R12854 gnd.n3487 gnd.n3486 9.3005
R12855 gnd.n3488 gnd.n3411 9.3005
R12856 gnd.n3491 gnd.n3489 9.3005
R12857 gnd.n3492 gnd.n3410 9.3005
R12858 gnd.n3495 gnd.n3494 9.3005
R12859 gnd.n3496 gnd.n3409 9.3005
R12860 gnd.n3499 gnd.n3497 9.3005
R12861 gnd.n3500 gnd.n3408 9.3005
R12862 gnd.n3503 gnd.n3502 9.3005
R12863 gnd.n3504 gnd.n3407 9.3005
R12864 gnd.n3507 gnd.n3505 9.3005
R12865 gnd.n3508 gnd.n3406 9.3005
R12866 gnd.n3511 gnd.n3510 9.3005
R12867 gnd.n3512 gnd.n3405 9.3005
R12868 gnd.n3515 gnd.n3513 9.3005
R12869 gnd.n3516 gnd.n3404 9.3005
R12870 gnd.n3519 gnd.n3518 9.3005
R12871 gnd.n3520 gnd.n3403 9.3005
R12872 gnd.n3523 gnd.n3521 9.3005
R12873 gnd.n3524 gnd.n3402 9.3005
R12874 gnd.n3526 gnd.n3525 9.3005
R12875 gnd.n3527 gnd.n3401 9.3005
R12876 gnd.n3546 gnd.n3528 9.3005
R12877 gnd.n3545 gnd.n3529 9.3005
R12878 gnd.n3544 gnd.n3530 9.3005
R12879 gnd.n3542 gnd.n3531 9.3005
R12880 gnd.n3475 gnd.n3473 9.3005
R12881 gnd.n3469 gnd.n3468 9.3005
R12882 gnd.n3467 gnd.n3419 9.3005
R12883 gnd.n3466 gnd.n3465 9.3005
R12884 gnd.n3462 gnd.n3422 9.3005
R12885 gnd.n3461 gnd.n3458 9.3005
R12886 gnd.n3457 gnd.n3423 9.3005
R12887 gnd.n3456 gnd.n3455 9.3005
R12888 gnd.n3452 gnd.n3424 9.3005
R12889 gnd.n3451 gnd.n3448 9.3005
R12890 gnd.n3447 gnd.n3425 9.3005
R12891 gnd.n3446 gnd.n3445 9.3005
R12892 gnd.n3442 gnd.n3426 9.3005
R12893 gnd.n3441 gnd.n3438 9.3005
R12894 gnd.n3437 gnd.n3427 9.3005
R12895 gnd.n3436 gnd.n3435 9.3005
R12896 gnd.n3432 gnd.n3428 9.3005
R12897 gnd.n3431 gnd.n3270 9.3005
R12898 gnd.n3470 gnd.n3415 9.3005
R12899 gnd.n3472 gnd.n3471 9.3005
R12900 gnd.n6102 gnd.n1296 9.3005
R12901 gnd.n6103 gnd.n1295 9.3005
R12902 gnd.n1294 gnd.n1291 9.3005
R12903 gnd.n6108 gnd.n1290 9.3005
R12904 gnd.n6109 gnd.n1289 9.3005
R12905 gnd.n6110 gnd.n1288 9.3005
R12906 gnd.n1287 gnd.n1284 9.3005
R12907 gnd.n6115 gnd.n1283 9.3005
R12908 gnd.n6117 gnd.n1280 9.3005
R12909 gnd.n6118 gnd.n1279 9.3005
R12910 gnd.n1278 gnd.n1275 9.3005
R12911 gnd.n6123 gnd.n1274 9.3005
R12912 gnd.n6124 gnd.n1273 9.3005
R12913 gnd.n6125 gnd.n1272 9.3005
R12914 gnd.n1271 gnd.n1268 9.3005
R12915 gnd.n6130 gnd.n1267 9.3005
R12916 gnd.n6131 gnd.n1266 9.3005
R12917 gnd.n6132 gnd.n1265 9.3005
R12918 gnd.n1264 gnd.n1261 9.3005
R12919 gnd.n6137 gnd.n1260 9.3005
R12920 gnd.n6138 gnd.n1259 9.3005
R12921 gnd.n6139 gnd.n1258 9.3005
R12922 gnd.n1257 gnd.n1254 9.3005
R12923 gnd.n1256 gnd.n1252 9.3005
R12924 gnd.n6146 gnd.n1251 9.3005
R12925 gnd.n6148 gnd.n6147 9.3005
R12926 gnd.n1513 gnd.n1512 9.3005
R12927 gnd.n1521 gnd.n1520 9.3005
R12928 gnd.n1522 gnd.n1510 9.3005
R12929 gnd.n1524 gnd.n1523 9.3005
R12930 gnd.n1508 gnd.n1507 9.3005
R12931 gnd.n1531 gnd.n1530 9.3005
R12932 gnd.n1532 gnd.n1506 9.3005
R12933 gnd.n1534 gnd.n1533 9.3005
R12934 gnd.n1504 gnd.n1501 9.3005
R12935 gnd.n1541 gnd.n1540 9.3005
R12936 gnd.n1542 gnd.n1500 9.3005
R12937 gnd.n1544 gnd.n1543 9.3005
R12938 gnd.n1498 gnd.n1497 9.3005
R12939 gnd.n1551 gnd.n1550 9.3005
R12940 gnd.n1552 gnd.n1496 9.3005
R12941 gnd.n1554 gnd.n1553 9.3005
R12942 gnd.n1494 gnd.n1493 9.3005
R12943 gnd.n1561 gnd.n1560 9.3005
R12944 gnd.n1562 gnd.n1492 9.3005
R12945 gnd.n1564 gnd.n1563 9.3005
R12946 gnd.n1490 gnd.n1489 9.3005
R12947 gnd.n1571 gnd.n1570 9.3005
R12948 gnd.n1572 gnd.n1488 9.3005
R12949 gnd.n1574 gnd.n1573 9.3005
R12950 gnd.n1486 gnd.n1485 9.3005
R12951 gnd.n1581 gnd.n1580 9.3005
R12952 gnd.n1582 gnd.n1484 9.3005
R12953 gnd.n1584 gnd.n1583 9.3005
R12954 gnd.n1482 gnd.n1479 9.3005
R12955 gnd.n1590 gnd.n1589 9.3005
R12956 gnd.n1511 gnd.n1297 9.3005
R12957 gnd.n3292 gnd.n3272 9.3005
R12958 gnd.n3551 gnd.n3293 9.3005
R12959 gnd.n3701 gnd.n3294 9.3005
R12960 gnd.n3700 gnd.n3295 9.3005
R12961 gnd.n3699 gnd.n3296 9.3005
R12962 gnd.n3557 gnd.n3297 9.3005
R12963 gnd.n3689 gnd.n3313 9.3005
R12964 gnd.n3688 gnd.n3314 9.3005
R12965 gnd.n3687 gnd.n3315 9.3005
R12966 gnd.n3564 gnd.n3316 9.3005
R12967 gnd.n3677 gnd.n3332 9.3005
R12968 gnd.n3676 gnd.n3333 9.3005
R12969 gnd.n3675 gnd.n3334 9.3005
R12970 gnd.n3571 gnd.n3335 9.3005
R12971 gnd.n3665 gnd.n3351 9.3005
R12972 gnd.n3664 gnd.n3352 9.3005
R12973 gnd.n3663 gnd.n3353 9.3005
R12974 gnd.n3578 gnd.n3354 9.3005
R12975 gnd.n3653 gnd.n3370 9.3005
R12976 gnd.n3652 gnd.n3371 9.3005
R12977 gnd.n3651 gnd.n3372 9.3005
R12978 gnd.n3585 gnd.n3373 9.3005
R12979 gnd.n3641 gnd.n3389 9.3005
R12980 gnd.n3640 gnd.n3390 9.3005
R12981 gnd.n3639 gnd.n3391 9.3005
R12982 gnd.n3549 gnd.n3392 9.3005
R12983 gnd.n3627 gnd.n3626 9.3005
R12984 gnd.n3550 gnd.n1787 9.3005
R12985 gnd.n5345 gnd.n1788 9.3005
R12986 gnd.n5344 gnd.n1789 9.3005
R12987 gnd.n5343 gnd.n1790 9.3005
R12988 gnd.n3593 gnd.n1791 9.3005
R12989 gnd.n5331 gnd.n1800 9.3005
R12990 gnd.n5330 gnd.n1801 9.3005
R12991 gnd.n5329 gnd.n1802 9.3005
R12992 gnd.n3594 gnd.n1803 9.3005
R12993 gnd.n3609 gnd.n3595 9.3005
R12994 gnd.n3608 gnd.n3607 9.3005
R12995 gnd.n1758 gnd.n1746 9.3005
R12996 gnd.n5390 gnd.n1747 9.3005
R12997 gnd.n5389 gnd.n1748 9.3005
R12998 gnd.n5388 gnd.n1749 9.3005
R12999 gnd.n5387 gnd.n1750 9.3005
R13000 gnd.n1723 gnd.n1708 9.3005
R13001 gnd.n5440 gnd.n1709 9.3005
R13002 gnd.n5439 gnd.n1710 9.3005
R13003 gnd.n5438 gnd.n1711 9.3005
R13004 gnd.n5437 gnd.n1712 9.3005
R13005 gnd.n5415 gnd.n1673 9.3005
R13006 gnd.n5475 gnd.n1674 9.3005
R13007 gnd.n5474 gnd.n1675 9.3005
R13008 gnd.n5473 gnd.n5472 9.3005
R13009 gnd.n1676 gnd.n1643 9.3005
R13010 gnd.n5543 gnd.n1644 9.3005
R13011 gnd.n5542 gnd.n1645 9.3005
R13012 gnd.n5541 gnd.n1646 9.3005
R13013 gnd.n5540 gnd.n1647 9.3005
R13014 gnd.n1618 gnd.n1617 9.3005
R13015 gnd.n5583 gnd.n5581 9.3005
R13016 gnd.n5582 gnd.n1598 9.3005
R13017 gnd.n5598 gnd.n1597 9.3005
R13018 gnd.n5600 gnd.n5599 9.3005
R13019 gnd.n5601 gnd.n1591 9.3005
R13020 gnd.n5607 gnd.n1592 9.3005
R13021 gnd.n3713 gnd.n3271 9.3005
R13022 gnd.n3273 gnd.n3272 9.3005
R13023 gnd.n3552 gnd.n3551 9.3005
R13024 gnd.n3553 gnd.n3294 9.3005
R13025 gnd.n3555 gnd.n3295 9.3005
R13026 gnd.n3556 gnd.n3296 9.3005
R13027 gnd.n3559 gnd.n3557 9.3005
R13028 gnd.n3560 gnd.n3313 9.3005
R13029 gnd.n3562 gnd.n3314 9.3005
R13030 gnd.n3563 gnd.n3315 9.3005
R13031 gnd.n3566 gnd.n3564 9.3005
R13032 gnd.n3567 gnd.n3332 9.3005
R13033 gnd.n3569 gnd.n3333 9.3005
R13034 gnd.n3570 gnd.n3334 9.3005
R13035 gnd.n3573 gnd.n3571 9.3005
R13036 gnd.n3574 gnd.n3351 9.3005
R13037 gnd.n3576 gnd.n3352 9.3005
R13038 gnd.n3577 gnd.n3353 9.3005
R13039 gnd.n3580 gnd.n3578 9.3005
R13040 gnd.n3581 gnd.n3370 9.3005
R13041 gnd.n3583 gnd.n3371 9.3005
R13042 gnd.n3584 gnd.n3372 9.3005
R13043 gnd.n3587 gnd.n3585 9.3005
R13044 gnd.n3588 gnd.n3389 9.3005
R13045 gnd.n3590 gnd.n3390 9.3005
R13046 gnd.n3591 gnd.n3391 9.3005
R13047 gnd.n3592 gnd.n3549 9.3005
R13048 gnd.n3626 gnd.n3625 9.3005
R13049 gnd.n3624 gnd.n3550 9.3005
R13050 gnd.n3622 gnd.n1788 9.3005
R13051 gnd.n3621 gnd.n1789 9.3005
R13052 gnd.n3619 gnd.n1790 9.3005
R13053 gnd.n3618 gnd.n3593 9.3005
R13054 gnd.n3616 gnd.n1800 9.3005
R13055 gnd.n3615 gnd.n1801 9.3005
R13056 gnd.n3613 gnd.n1802 9.3005
R13057 gnd.n3612 gnd.n3594 9.3005
R13058 gnd.n3610 gnd.n3609 9.3005
R13059 gnd.n3608 gnd.n1757 9.3005
R13060 gnd.n5368 gnd.n1758 9.3005
R13061 gnd.n5369 gnd.n1747 9.3005
R13062 gnd.n5371 gnd.n1748 9.3005
R13063 gnd.n5370 gnd.n1749 9.3005
R13064 gnd.n1750 gnd.n1722 9.3005
R13065 gnd.n5413 gnd.n1723 9.3005
R13066 gnd.n5414 gnd.n1709 9.3005
R13067 gnd.n5421 gnd.n1710 9.3005
R13068 gnd.n5420 gnd.n1711 9.3005
R13069 gnd.n5419 gnd.n1712 9.3005
R13070 gnd.n5418 gnd.n5415 9.3005
R13071 gnd.n5416 gnd.n1674 9.3005
R13072 gnd.n1678 gnd.n1675 9.3005
R13073 gnd.n5472 gnd.n5471 9.3005
R13074 gnd.n5470 gnd.n1676 9.3005
R13075 gnd.n1683 gnd.n1644 9.3005
R13076 gnd.n1682 gnd.n1645 9.3005
R13077 gnd.n1679 gnd.n1646 9.3005
R13078 gnd.n1647 gnd.n1619 9.3005
R13079 gnd.n5579 gnd.n1618 9.3005
R13080 gnd.n5581 gnd.n5580 9.3005
R13081 gnd.n1599 gnd.n1598 9.3005
R13082 gnd.n5598 gnd.n5597 9.3005
R13083 gnd.n5599 gnd.n1593 9.3005
R13084 gnd.n5605 gnd.n1591 9.3005
R13085 gnd.n5607 gnd.n5606 9.3005
R13086 gnd.n3713 gnd.n3712 9.3005
R13087 gnd.n3717 gnd.n3716 9.3005
R13088 gnd.n3720 gnd.n3266 9.3005
R13089 gnd.n3721 gnd.n3265 9.3005
R13090 gnd.n3724 gnd.n3264 9.3005
R13091 gnd.n3725 gnd.n3263 9.3005
R13092 gnd.n3728 gnd.n3262 9.3005
R13093 gnd.n3729 gnd.n3261 9.3005
R13094 gnd.n3732 gnd.n3260 9.3005
R13095 gnd.n3733 gnd.n3259 9.3005
R13096 gnd.n3736 gnd.n3258 9.3005
R13097 gnd.n3737 gnd.n3257 9.3005
R13098 gnd.n3740 gnd.n3256 9.3005
R13099 gnd.n3741 gnd.n3255 9.3005
R13100 gnd.n3744 gnd.n3254 9.3005
R13101 gnd.n3745 gnd.n3253 9.3005
R13102 gnd.n3748 gnd.n3252 9.3005
R13103 gnd.n3749 gnd.n3251 9.3005
R13104 gnd.n3752 gnd.n3250 9.3005
R13105 gnd.n3753 gnd.n3249 9.3005
R13106 gnd.n3756 gnd.n3248 9.3005
R13107 gnd.n3760 gnd.n3244 9.3005
R13108 gnd.n3761 gnd.n3243 9.3005
R13109 gnd.n3764 gnd.n3242 9.3005
R13110 gnd.n3765 gnd.n3241 9.3005
R13111 gnd.n3768 gnd.n3240 9.3005
R13112 gnd.n3769 gnd.n3239 9.3005
R13113 gnd.n3772 gnd.n3238 9.3005
R13114 gnd.n3773 gnd.n3237 9.3005
R13115 gnd.n3776 gnd.n3236 9.3005
R13116 gnd.n3777 gnd.n3235 9.3005
R13117 gnd.n3780 gnd.n3234 9.3005
R13118 gnd.n3781 gnd.n3233 9.3005
R13119 gnd.n3784 gnd.n3232 9.3005
R13120 gnd.n3785 gnd.n3231 9.3005
R13121 gnd.n3788 gnd.n3230 9.3005
R13122 gnd.n3789 gnd.n3229 9.3005
R13123 gnd.n3792 gnd.n3228 9.3005
R13124 gnd.n3793 gnd.n3227 9.3005
R13125 gnd.n3796 gnd.n3226 9.3005
R13126 gnd.n3798 gnd.n3223 9.3005
R13127 gnd.n3801 gnd.n3222 9.3005
R13128 gnd.n3802 gnd.n3221 9.3005
R13129 gnd.n3805 gnd.n3220 9.3005
R13130 gnd.n3806 gnd.n3219 9.3005
R13131 gnd.n3809 gnd.n3218 9.3005
R13132 gnd.n3810 gnd.n3217 9.3005
R13133 gnd.n3813 gnd.n3216 9.3005
R13134 gnd.n3814 gnd.n3215 9.3005
R13135 gnd.n3817 gnd.n3214 9.3005
R13136 gnd.n3818 gnd.n3213 9.3005
R13137 gnd.n3821 gnd.n3212 9.3005
R13138 gnd.n3822 gnd.n3211 9.3005
R13139 gnd.n3825 gnd.n3210 9.3005
R13140 gnd.n3827 gnd.n3209 9.3005
R13141 gnd.n3828 gnd.n3208 9.3005
R13142 gnd.n3829 gnd.n3207 9.3005
R13143 gnd.n3830 gnd.n3206 9.3005
R13144 gnd.n3757 gnd.n3245 9.3005
R13145 gnd.n3715 gnd.n3267 9.3005
R13146 gnd.n3707 gnd.n3281 9.3005
R13147 gnd.n3706 gnd.n3282 9.3005
R13148 gnd.n3705 gnd.n3283 9.3005
R13149 gnd.n3303 gnd.n3284 9.3005
R13150 gnd.n3695 gnd.n3304 9.3005
R13151 gnd.n3694 gnd.n3305 9.3005
R13152 gnd.n3693 gnd.n3306 9.3005
R13153 gnd.n3321 gnd.n3307 9.3005
R13154 gnd.n3683 gnd.n3322 9.3005
R13155 gnd.n3682 gnd.n3323 9.3005
R13156 gnd.n3681 gnd.n3324 9.3005
R13157 gnd.n3341 gnd.n3325 9.3005
R13158 gnd.n3671 gnd.n3342 9.3005
R13159 gnd.n3670 gnd.n3343 9.3005
R13160 gnd.n3669 gnd.n3344 9.3005
R13161 gnd.n3359 gnd.n3345 9.3005
R13162 gnd.n3659 gnd.n3360 9.3005
R13163 gnd.n3658 gnd.n3361 9.3005
R13164 gnd.n3657 gnd.n3362 9.3005
R13165 gnd.n3379 gnd.n3363 9.3005
R13166 gnd.n3647 gnd.n3380 9.3005
R13167 gnd.n3646 gnd.n3381 9.3005
R13168 gnd.n3645 gnd.n3382 9.3005
R13169 gnd.n3632 gnd.n3383 9.3005
R13170 gnd.n3635 gnd.n3633 9.3005
R13171 gnd.n3634 gnd.n1773 9.3005
R13172 gnd.n5354 gnd.n5353 9.3005
R13173 gnd.n1738 gnd.n1737 9.3005
R13174 gnd.n5395 gnd.n5394 9.3005
R13175 gnd.n5396 gnd.n1736 9.3005
R13176 gnd.n5400 gnd.n5397 9.3005
R13177 gnd.n5399 gnd.n5398 9.3005
R13178 gnd.n1700 gnd.n1699 9.3005
R13179 gnd.n5445 gnd.n5444 9.3005
R13180 gnd.n5446 gnd.n1698 9.3005
R13181 gnd.n5450 gnd.n5447 9.3005
R13182 gnd.n5449 gnd.n5448 9.3005
R13183 gnd.n1666 gnd.n1665 9.3005
R13184 gnd.n5480 gnd.n5479 9.3005
R13185 gnd.n5481 gnd.n1664 9.3005
R13186 gnd.n5483 gnd.n5482 9.3005
R13187 gnd.n1635 gnd.n1634 9.3005
R13188 gnd.n5548 gnd.n5547 9.3005
R13189 gnd.n5549 gnd.n1633 9.3005
R13190 gnd.n5553 gnd.n5550 9.3005
R13191 gnd.n5552 gnd.n5551 9.3005
R13192 gnd.n1609 gnd.n1608 9.3005
R13193 gnd.n5588 gnd.n5587 9.3005
R13194 gnd.n5589 gnd.n1607 9.3005
R13195 gnd.n5593 gnd.n5590 9.3005
R13196 gnd.n5592 gnd.n5591 9.3005
R13197 gnd.n1250 gnd.n1249 9.3005
R13198 gnd.n6150 gnd.n6149 9.3005
R13199 gnd.n3280 gnd.n3279 9.3005
R13200 gnd.n5355 gnd.n5352 9.3005
R13201 gnd.n5319 gnd.n1810 9.3005
R13202 gnd.n5318 gnd.n5317 9.3005
R13203 gnd.n1812 gnd.n1811 9.3005
R13204 gnd.n3145 gnd.n3144 9.3005
R13205 gnd.n3143 gnd.n1816 9.3005
R13206 gnd.n3142 gnd.n3141 9.3005
R13207 gnd.n1818 gnd.n1817 9.3005
R13208 gnd.n3135 gnd.n3134 9.3005
R13209 gnd.n3133 gnd.n1822 9.3005
R13210 gnd.n3132 gnd.n3131 9.3005
R13211 gnd.n1824 gnd.n1823 9.3005
R13212 gnd.n3125 gnd.n3124 9.3005
R13213 gnd.n3123 gnd.n1828 9.3005
R13214 gnd.n3122 gnd.n3121 9.3005
R13215 gnd.n1830 gnd.n1829 9.3005
R13216 gnd.n3115 gnd.n3114 9.3005
R13217 gnd.n3113 gnd.n1834 9.3005
R13218 gnd.n3112 gnd.n3111 9.3005
R13219 gnd.n1836 gnd.n1835 9.3005
R13220 gnd.n3105 gnd.n3104 9.3005
R13221 gnd.n3103 gnd.n1840 9.3005
R13222 gnd.n3102 gnd.n3101 9.3005
R13223 gnd.n1842 gnd.n1841 9.3005
R13224 gnd.n3095 gnd.n3094 9.3005
R13225 gnd.n3093 gnd.n1846 9.3005
R13226 gnd.n3092 gnd.n3091 9.3005
R13227 gnd.n1848 gnd.n1847 9.3005
R13228 gnd.n3085 gnd.n3084 9.3005
R13229 gnd.n3083 gnd.n1852 9.3005
R13230 gnd.n3082 gnd.n3081 9.3005
R13231 gnd.n1854 gnd.n1853 9.3005
R13232 gnd.n3075 gnd.n3074 9.3005
R13233 gnd.n3073 gnd.n1858 9.3005
R13234 gnd.n3072 gnd.n3071 9.3005
R13235 gnd.n1860 gnd.n1859 9.3005
R13236 gnd.n3065 gnd.n3064 9.3005
R13237 gnd.n3063 gnd.n1864 9.3005
R13238 gnd.n3062 gnd.n3061 9.3005
R13239 gnd.n1866 gnd.n1865 9.3005
R13240 gnd.n3055 gnd.n3054 9.3005
R13241 gnd.n3053 gnd.n1870 9.3005
R13242 gnd.n3052 gnd.n3051 9.3005
R13243 gnd.n1872 gnd.n1871 9.3005
R13244 gnd.n3045 gnd.n3044 9.3005
R13245 gnd.n3043 gnd.n1876 9.3005
R13246 gnd.n3042 gnd.n3041 9.3005
R13247 gnd.n1878 gnd.n1877 9.3005
R13248 gnd.n3035 gnd.n3034 9.3005
R13249 gnd.n3033 gnd.n1882 9.3005
R13250 gnd.n3032 gnd.n3031 9.3005
R13251 gnd.n1884 gnd.n1883 9.3005
R13252 gnd.n3025 gnd.n3024 9.3005
R13253 gnd.n3023 gnd.n1888 9.3005
R13254 gnd.n3022 gnd.n3021 9.3005
R13255 gnd.n1890 gnd.n1889 9.3005
R13256 gnd.n3015 gnd.n3014 9.3005
R13257 gnd.n3013 gnd.n1894 9.3005
R13258 gnd.n3012 gnd.n3011 9.3005
R13259 gnd.n1896 gnd.n1895 9.3005
R13260 gnd.n3005 gnd.n3004 9.3005
R13261 gnd.n3003 gnd.n1900 9.3005
R13262 gnd.n3002 gnd.n3001 9.3005
R13263 gnd.n1902 gnd.n1901 9.3005
R13264 gnd.n2995 gnd.n2994 9.3005
R13265 gnd.n2993 gnd.n1906 9.3005
R13266 gnd.n2992 gnd.n2991 9.3005
R13267 gnd.n1908 gnd.n1907 9.3005
R13268 gnd.n2985 gnd.n2984 9.3005
R13269 gnd.n2983 gnd.n1912 9.3005
R13270 gnd.n2982 gnd.n2981 9.3005
R13271 gnd.n1914 gnd.n1913 9.3005
R13272 gnd.n2975 gnd.n2974 9.3005
R13273 gnd.n2973 gnd.n1918 9.3005
R13274 gnd.n2972 gnd.n2971 9.3005
R13275 gnd.n1920 gnd.n1919 9.3005
R13276 gnd.n2965 gnd.n2964 9.3005
R13277 gnd.n2963 gnd.n1924 9.3005
R13278 gnd.n2962 gnd.n2961 9.3005
R13279 gnd.n1926 gnd.n1925 9.3005
R13280 gnd.n2955 gnd.n2954 9.3005
R13281 gnd.n2953 gnd.n1930 9.3005
R13282 gnd.n2952 gnd.n2951 9.3005
R13283 gnd.n1932 gnd.n1931 9.3005
R13284 gnd.n2945 gnd.n2944 9.3005
R13285 gnd.n5321 gnd.n5320 9.3005
R13286 gnd.n7098 gnd.n740 9.3005
R13287 gnd.n1221 gnd.n1220 9.3005
R13288 gnd.n6175 gnd.n6174 9.3005
R13289 gnd.n6176 gnd.n1219 9.3005
R13290 gnd.n6178 gnd.n6177 9.3005
R13291 gnd.n1207 gnd.n1206 9.3005
R13292 gnd.n6191 gnd.n6190 9.3005
R13293 gnd.n6192 gnd.n1205 9.3005
R13294 gnd.n6194 gnd.n6193 9.3005
R13295 gnd.n1192 gnd.n1191 9.3005
R13296 gnd.n6207 gnd.n6206 9.3005
R13297 gnd.n6208 gnd.n1190 9.3005
R13298 gnd.n6210 gnd.n6209 9.3005
R13299 gnd.n1178 gnd.n1177 9.3005
R13300 gnd.n6223 gnd.n6222 9.3005
R13301 gnd.n6224 gnd.n1176 9.3005
R13302 gnd.n6226 gnd.n6225 9.3005
R13303 gnd.n1164 gnd.n1163 9.3005
R13304 gnd.n6239 gnd.n6238 9.3005
R13305 gnd.n6240 gnd.n1162 9.3005
R13306 gnd.n6242 gnd.n6241 9.3005
R13307 gnd.n1149 gnd.n1148 9.3005
R13308 gnd.n6255 gnd.n6254 9.3005
R13309 gnd.n6256 gnd.n1147 9.3005
R13310 gnd.n6258 gnd.n6257 9.3005
R13311 gnd.n1134 gnd.n1133 9.3005
R13312 gnd.n6271 gnd.n6270 9.3005
R13313 gnd.n6272 gnd.n1132 9.3005
R13314 gnd.n6274 gnd.n6273 9.3005
R13315 gnd.n1120 gnd.n1119 9.3005
R13316 gnd.n6287 gnd.n6286 9.3005
R13317 gnd.n6288 gnd.n1118 9.3005
R13318 gnd.n6290 gnd.n6289 9.3005
R13319 gnd.n1107 gnd.n1106 9.3005
R13320 gnd.n6303 gnd.n6302 9.3005
R13321 gnd.n6304 gnd.n1105 9.3005
R13322 gnd.n6306 gnd.n6305 9.3005
R13323 gnd.n1093 gnd.n1092 9.3005
R13324 gnd.n6319 gnd.n6318 9.3005
R13325 gnd.n6320 gnd.n1091 9.3005
R13326 gnd.n6322 gnd.n6321 9.3005
R13327 gnd.n1077 gnd.n1076 9.3005
R13328 gnd.n6335 gnd.n6334 9.3005
R13329 gnd.n6336 gnd.n1074 9.3005
R13330 gnd.n6344 gnd.n6343 9.3005
R13331 gnd.n6342 gnd.n1075 9.3005
R13332 gnd.n6341 gnd.n6340 9.3005
R13333 gnd.n6339 gnd.n6337 9.3005
R13334 gnd.n1039 gnd.n1037 9.3005
R13335 gnd.n6402 gnd.n6401 9.3005
R13336 gnd.n6400 gnd.n1038 9.3005
R13337 gnd.n6399 gnd.n6398 9.3005
R13338 gnd.n6397 gnd.n1040 9.3005
R13339 gnd.n1000 gnd.n998 9.3005
R13340 gnd.n6460 gnd.n6459 9.3005
R13341 gnd.n6458 gnd.n999 9.3005
R13342 gnd.n6457 gnd.n6456 9.3005
R13343 gnd.n6455 gnd.n1001 9.3005
R13344 gnd.n6454 gnd.n6453 9.3005
R13345 gnd.n6452 gnd.n6451 9.3005
R13346 gnd.n916 gnd.n915 9.3005
R13347 gnd.n6911 gnd.n6910 9.3005
R13348 gnd.n6912 gnd.n914 9.3005
R13349 gnd.n6914 gnd.n6913 9.3005
R13350 gnd.n902 gnd.n901 9.3005
R13351 gnd.n6927 gnd.n6926 9.3005
R13352 gnd.n6928 gnd.n900 9.3005
R13353 gnd.n6930 gnd.n6929 9.3005
R13354 gnd.n889 gnd.n888 9.3005
R13355 gnd.n6943 gnd.n6942 9.3005
R13356 gnd.n6944 gnd.n887 9.3005
R13357 gnd.n6946 gnd.n6945 9.3005
R13358 gnd.n875 gnd.n874 9.3005
R13359 gnd.n6959 gnd.n6958 9.3005
R13360 gnd.n6960 gnd.n873 9.3005
R13361 gnd.n6962 gnd.n6961 9.3005
R13362 gnd.n860 gnd.n859 9.3005
R13363 gnd.n6975 gnd.n6974 9.3005
R13364 gnd.n6976 gnd.n858 9.3005
R13365 gnd.n6978 gnd.n6977 9.3005
R13366 gnd.n846 gnd.n845 9.3005
R13367 gnd.n6991 gnd.n6990 9.3005
R13368 gnd.n6992 gnd.n844 9.3005
R13369 gnd.n6994 gnd.n6993 9.3005
R13370 gnd.n832 gnd.n831 9.3005
R13371 gnd.n7007 gnd.n7006 9.3005
R13372 gnd.n7008 gnd.n830 9.3005
R13373 gnd.n7010 gnd.n7009 9.3005
R13374 gnd.n818 gnd.n817 9.3005
R13375 gnd.n7023 gnd.n7022 9.3005
R13376 gnd.n7024 gnd.n816 9.3005
R13377 gnd.n7026 gnd.n7025 9.3005
R13378 gnd.n803 gnd.n802 9.3005
R13379 gnd.n7039 gnd.n7038 9.3005
R13380 gnd.n7040 gnd.n801 9.3005
R13381 gnd.n7042 gnd.n7041 9.3005
R13382 gnd.n790 gnd.n789 9.3005
R13383 gnd.n7058 gnd.n7057 9.3005
R13384 gnd.n7059 gnd.n788 9.3005
R13385 gnd.n7061 gnd.n7060 9.3005
R13386 gnd.n742 gnd.n741 9.3005
R13387 gnd.n7097 gnd.n7096 9.3005
R13388 gnd.n6162 gnd.n6161 9.3005
R13389 gnd.n6160 gnd.n6159 9.3005
R13390 gnd.n3539 gnd.n3533 9.3005
R13391 gnd.n3538 gnd.n3537 9.3005
R13392 gnd.n3536 gnd.n3534 9.3005
R13393 gnd.n1764 gnd.n1763 9.3005
R13394 gnd.n5360 gnd.n5359 9.3005
R13395 gnd.n5361 gnd.n1761 9.3005
R13396 gnd.n5364 gnd.n5363 9.3005
R13397 gnd.n5362 gnd.n1762 9.3005
R13398 gnd.n1729 gnd.n1728 9.3005
R13399 gnd.n5405 gnd.n5404 9.3005
R13400 gnd.n5406 gnd.n1726 9.3005
R13401 gnd.n5409 gnd.n5408 9.3005
R13402 gnd.n5407 gnd.n1727 9.3005
R13403 gnd.n1690 gnd.n1689 9.3005
R13404 gnd.n5455 gnd.n5454 9.3005
R13405 gnd.n5456 gnd.n1687 9.3005
R13406 gnd.n5458 gnd.n5457 9.3005
R13407 gnd.n5459 gnd.n1686 9.3005
R13408 gnd.n5462 gnd.n5461 9.3005
R13409 gnd.n5463 gnd.n1684 9.3005
R13410 gnd.n5466 gnd.n5465 9.3005
R13411 gnd.n5464 gnd.n1685 9.3005
R13412 gnd.n1625 gnd.n1624 9.3005
R13413 gnd.n5558 gnd.n5557 9.3005
R13414 gnd.n5559 gnd.n1622 9.3005
R13415 gnd.n5575 gnd.n5574 9.3005
R13416 gnd.n5573 gnd.n1623 9.3005
R13417 gnd.n5572 gnd.n5571 9.3005
R13418 gnd.n5570 gnd.n5560 9.3005
R13419 gnd.n5569 gnd.n5568 9.3005
R13420 gnd.n5567 gnd.n5565 9.3005
R13421 gnd.n5566 gnd.n1242 9.3005
R13422 gnd.n5722 gnd.n5721 9.3005
R13423 gnd.n5720 gnd.n5719 9.3005
R13424 gnd.n5620 gnd.n5619 9.3005
R13425 gnd.n5714 gnd.n5713 9.3005
R13426 gnd.n5712 gnd.n5711 9.3005
R13427 gnd.n5632 gnd.n5631 9.3005
R13428 gnd.n5706 gnd.n5705 9.3005
R13429 gnd.n5704 gnd.n5703 9.3005
R13430 gnd.n5643 gnd.n5642 9.3005
R13431 gnd.n5698 gnd.n5697 9.3005
R13432 gnd.n5696 gnd.n5695 9.3005
R13433 gnd.n5655 gnd.n5654 9.3005
R13434 gnd.n5690 gnd.n5689 9.3005
R13435 gnd.n5688 gnd.n5687 9.3005
R13436 gnd.n5666 gnd.n5665 9.3005
R13437 gnd.n5682 gnd.n5681 9.3005
R13438 gnd.n5673 gnd.n1239 9.3005
R13439 gnd.n6156 gnd.n6155 9.3005
R13440 gnd.n5614 gnd.n5609 9.3005
R13441 gnd.n6158 gnd.n6157 9.3005
R13442 gnd.n1236 gnd.n1234 9.3005
R13443 gnd.n5676 gnd.n5675 9.3005
R13444 gnd.n5684 gnd.n5683 9.3005
R13445 gnd.n5686 gnd.n5685 9.3005
R13446 gnd.n5659 gnd.n5658 9.3005
R13447 gnd.n5692 gnd.n5691 9.3005
R13448 gnd.n5694 gnd.n5693 9.3005
R13449 gnd.n5649 gnd.n5648 9.3005
R13450 gnd.n5700 gnd.n5699 9.3005
R13451 gnd.n5702 gnd.n5701 9.3005
R13452 gnd.n5636 gnd.n5635 9.3005
R13453 gnd.n5708 gnd.n5707 9.3005
R13454 gnd.n5710 gnd.n5709 9.3005
R13455 gnd.n5626 gnd.n5625 9.3005
R13456 gnd.n5716 gnd.n5715 9.3005
R13457 gnd.n5718 gnd.n5717 9.3005
R13458 gnd.n5613 gnd.n5612 9.3005
R13459 gnd.n5724 gnd.n5723 9.3005
R13460 gnd.n5726 gnd.n5725 9.3005
R13461 gnd.n5727 gnd.n1478 9.3005
R13462 gnd.n5730 gnd.n5729 9.3005
R13463 gnd.n5731 gnd.n1473 9.3005
R13464 gnd.n5733 gnd.n5732 9.3005
R13465 gnd.n5734 gnd.n1472 9.3005
R13466 gnd.n5736 gnd.n5735 9.3005
R13467 gnd.n1454 gnd.n1453 9.3005
R13468 gnd.n5742 gnd.n5741 9.3005
R13469 gnd.n5745 gnd.n5744 9.3005
R13470 gnd.n5746 gnd.n1450 9.3005
R13471 gnd.n5749 gnd.n5748 9.3005
R13472 gnd.n5750 gnd.n1448 9.3005
R13473 gnd.n5752 gnd.n5751 9.3005
R13474 gnd.n5753 gnd.n1447 9.3005
R13475 gnd.n5756 gnd.n5755 9.3005
R13476 gnd.n5757 gnd.n1445 9.3005
R13477 gnd.n5759 gnd.n5758 9.3005
R13478 gnd.n5760 gnd.n1444 9.3005
R13479 gnd.n5763 gnd.n5762 9.3005
R13480 gnd.n5764 gnd.n1442 9.3005
R13481 gnd.n5766 gnd.n5765 9.3005
R13482 gnd.n5767 gnd.n1441 9.3005
R13483 gnd.n5770 gnd.n5769 9.3005
R13484 gnd.n5771 gnd.n1438 9.3005
R13485 gnd.n5773 gnd.n5772 9.3005
R13486 gnd.n5774 gnd.n1437 9.3005
R13487 gnd.n5777 gnd.n5776 9.3005
R13488 gnd.n5778 gnd.n1435 9.3005
R13489 gnd.n6020 gnd.n6019 9.3005
R13490 gnd.n6018 gnd.n1436 9.3005
R13491 gnd.n6017 gnd.n6016 9.3005
R13492 gnd.n6015 gnd.n5779 9.3005
R13493 gnd.n6014 gnd.n6013 9.3005
R13494 gnd.n6012 gnd.n5782 9.3005
R13495 gnd.n6011 gnd.n6010 9.3005
R13496 gnd.n6009 gnd.n5783 9.3005
R13497 gnd.n6008 gnd.n6007 9.3005
R13498 gnd.n6006 gnd.n5786 9.3005
R13499 gnd.n6005 gnd.n6004 9.3005
R13500 gnd.n6003 gnd.n5787 9.3005
R13501 gnd.n6002 gnd.n6001 9.3005
R13502 gnd.n6000 gnd.n5790 9.3005
R13503 gnd.n5999 gnd.n5998 9.3005
R13504 gnd.n5997 gnd.n5791 9.3005
R13505 gnd.n5996 gnd.n5995 9.3005
R13506 gnd.n5994 gnd.n5794 9.3005
R13507 gnd.n5993 gnd.n5992 9.3005
R13508 gnd.n5991 gnd.n5795 9.3005
R13509 gnd.n5990 gnd.n5989 9.3005
R13510 gnd.n5988 gnd.n5798 9.3005
R13511 gnd.n5987 gnd.n5986 9.3005
R13512 gnd.n5985 gnd.n5799 9.3005
R13513 gnd.n5984 gnd.n5983 9.3005
R13514 gnd.n5982 gnd.n5973 9.3005
R13515 gnd.n5981 gnd.n5980 9.3005
R13516 gnd.n5979 gnd.n5974 9.3005
R13517 gnd.n5978 gnd.n5977 9.3005
R13518 gnd.n1021 gnd.n1020 9.3005
R13519 gnd.n6417 gnd.n6416 9.3005
R13520 gnd.n6418 gnd.n1018 9.3005
R13521 gnd.n6421 gnd.n6420 9.3005
R13522 gnd.n6419 gnd.n1019 9.3005
R13523 gnd.n981 gnd.n980 9.3005
R13524 gnd.n6475 gnd.n6474 9.3005
R13525 gnd.n6476 gnd.n978 9.3005
R13526 gnd.n6478 gnd.n6477 9.3005
R13527 gnd.n6479 gnd.n977 9.3005
R13528 gnd.n6482 gnd.n6481 9.3005
R13529 gnd.n6483 gnd.n976 9.3005
R13530 gnd.n6485 gnd.n6484 9.3005
R13531 gnd.n6486 gnd.n975 9.3005
R13532 gnd.n6489 gnd.n6488 9.3005
R13533 gnd.n6490 gnd.n974 9.3005
R13534 gnd.n6492 gnd.n6491 9.3005
R13535 gnd.n6493 gnd.n973 9.3005
R13536 gnd.n6496 gnd.n6495 9.3005
R13537 gnd.n6497 gnd.n971 9.3005
R13538 gnd.n6855 gnd.n6854 9.3005
R13539 gnd.n6853 gnd.n972 9.3005
R13540 gnd.n6852 gnd.n6851 9.3005
R13541 gnd.n6850 gnd.n6498 9.3005
R13542 gnd.n6849 gnd.n6848 9.3005
R13543 gnd.n6847 gnd.n6501 9.3005
R13544 gnd.n6846 gnd.n6845 9.3005
R13545 gnd.n6844 gnd.n6502 9.3005
R13546 gnd.n6843 gnd.n6842 9.3005
R13547 gnd.n6841 gnd.n6505 9.3005
R13548 gnd.n6840 gnd.n6839 9.3005
R13549 gnd.n6838 gnd.n6506 9.3005
R13550 gnd.n6837 gnd.n6836 9.3005
R13551 gnd.n6835 gnd.n6794 9.3005
R13552 gnd.n6834 gnd.n6833 9.3005
R13553 gnd.n6832 gnd.n6795 9.3005
R13554 gnd.n6831 gnd.n6830 9.3005
R13555 gnd.n6829 gnd.n6798 9.3005
R13556 gnd.n6828 gnd.n6827 9.3005
R13557 gnd.n6826 gnd.n6799 9.3005
R13558 gnd.n6825 gnd.n6824 9.3005
R13559 gnd.n6823 gnd.n6802 9.3005
R13560 gnd.n6822 gnd.n6821 9.3005
R13561 gnd.n6820 gnd.n6803 9.3005
R13562 gnd.n6819 gnd.n6818 9.3005
R13563 gnd.n6817 gnd.n6806 9.3005
R13564 gnd.n6816 gnd.n6815 9.3005
R13565 gnd.n6814 gnd.n6807 9.3005
R13566 gnd.n6813 gnd.n6812 9.3005
R13567 gnd.n6811 gnd.n6810 9.3005
R13568 gnd.n751 gnd.n750 9.3005
R13569 gnd.n7092 gnd.n7091 9.3005
R13570 gnd.n5743 gnd.n1451 9.3005
R13571 gnd.n7088 gnd.n752 9.3005
R13572 gnd.n7087 gnd.n7086 9.3005
R13573 gnd.n7085 gnd.n755 9.3005
R13574 gnd.n7084 gnd.n7083 9.3005
R13575 gnd.n7082 gnd.n756 9.3005
R13576 gnd.n679 gnd.n677 9.3005
R13577 gnd.n7090 gnd.n7089 9.3005
R13578 gnd.n7112 gnd.n7111 9.3005
R13579 gnd.n726 gnd.n725 9.3005
R13580 gnd.n7118 gnd.n7117 9.3005
R13581 gnd.n7120 gnd.n7119 9.3005
R13582 gnd.n718 gnd.n717 9.3005
R13583 gnd.n7126 gnd.n7125 9.3005
R13584 gnd.n7128 gnd.n7127 9.3005
R13585 gnd.n708 gnd.n707 9.3005
R13586 gnd.n7134 gnd.n7133 9.3005
R13587 gnd.n7136 gnd.n7135 9.3005
R13588 gnd.n700 gnd.n699 9.3005
R13589 gnd.n7142 gnd.n7141 9.3005
R13590 gnd.n7144 gnd.n7143 9.3005
R13591 gnd.n690 gnd.n689 9.3005
R13592 gnd.n7150 gnd.n7149 9.3005
R13593 gnd.n7152 gnd.n7151 9.3005
R13594 gnd.n686 gnd.n684 9.3005
R13595 gnd.n7110 gnd.n7106 9.3005
R13596 gnd.n736 gnd.n735 9.3005
R13597 gnd.n7157 gnd.n7156 9.3005
R13598 gnd.n7155 gnd.n678 9.3005
R13599 gnd.n7154 gnd.n7153 9.3005
R13600 gnd.n685 gnd.n683 9.3005
R13601 gnd.n7148 gnd.n7147 9.3005
R13602 gnd.n7146 gnd.n7145 9.3005
R13603 gnd.n694 gnd.n693 9.3005
R13604 gnd.n7140 gnd.n7139 9.3005
R13605 gnd.n7138 gnd.n7137 9.3005
R13606 gnd.n704 gnd.n703 9.3005
R13607 gnd.n7132 gnd.n7131 9.3005
R13608 gnd.n7130 gnd.n7129 9.3005
R13609 gnd.n712 gnd.n711 9.3005
R13610 gnd.n7124 gnd.n7123 9.3005
R13611 gnd.n7122 gnd.n7121 9.3005
R13612 gnd.n722 gnd.n721 9.3005
R13613 gnd.n7116 gnd.n7115 9.3005
R13614 gnd.n7114 gnd.n7113 9.3005
R13615 gnd.n737 gnd.n732 9.3005
R13616 gnd.n7105 gnd.n7104 9.3005
R13617 gnd.n7103 gnd.n7102 9.3005
R13618 gnd.n541 gnd.n540 9.3005
R13619 gnd.n7323 gnd.n7322 9.3005
R13620 gnd.n7324 gnd.n538 9.3005
R13621 gnd.n7327 gnd.n7326 9.3005
R13622 gnd.n7325 gnd.n539 9.3005
R13623 gnd.n510 gnd.n509 9.3005
R13624 gnd.n7365 gnd.n7364 9.3005
R13625 gnd.n7366 gnd.n507 9.3005
R13626 gnd.n7369 gnd.n7368 9.3005
R13627 gnd.n7367 gnd.n508 9.3005
R13628 gnd.n475 gnd.n474 9.3005
R13629 gnd.n7414 gnd.n7413 9.3005
R13630 gnd.n7415 gnd.n472 9.3005
R13631 gnd.n7418 gnd.n7417 9.3005
R13632 gnd.n7416 gnd.n473 9.3005
R13633 gnd.n444 gnd.n443 9.3005
R13634 gnd.n7451 gnd.n7450 9.3005
R13635 gnd.n7452 gnd.n441 9.3005
R13636 gnd.n7455 gnd.n7454 9.3005
R13637 gnd.n7453 gnd.n442 9.3005
R13638 gnd.n409 gnd.n408 9.3005
R13639 gnd.n7500 gnd.n7499 9.3005
R13640 gnd.n7501 gnd.n406 9.3005
R13641 gnd.n7506 gnd.n7505 9.3005
R13642 gnd.n7504 gnd.n407 9.3005
R13643 gnd.n7503 gnd.n7502 9.3005
R13644 gnd.n374 gnd.n373 9.3005
R13645 gnd.n7548 gnd.n7547 9.3005
R13646 gnd.n7549 gnd.n371 9.3005
R13647 gnd.n7551 gnd.n7550 9.3005
R13648 gnd.n372 gnd.n99 9.3005
R13649 gnd.n7100 gnd.n7099 9.3005
R13650 gnd.n7982 gnd.n100 9.3005
R13651 gnd.t18 gnd.n4009 9.24152
R13652 gnd.n3911 gnd.t195 9.24152
R13653 gnd.n5211 gnd.t167 9.24152
R13654 gnd.n3667 gnd.t225 9.24152
R13655 gnd.n5327 gnd.n5323 9.24152
R13656 gnd.n397 gnd.n368 9.24152
R13657 gnd.n7933 gnd.t263 9.24152
R13658 gnd.t407 gnd.t18 8.92286
R13659 gnd.n6022 gnd.t174 8.92286
R13660 gnd.n6252 gnd.n1153 8.92286
R13661 gnd.t164 gnd.n1145 8.92286
R13662 gnd.n6268 gnd.t19 8.92286
R13663 gnd.n5942 gnd.n5810 8.92286
R13664 gnd.n5948 gnd.n1059 8.92286
R13665 gnd.n6472 gnd.n985 8.92286
R13666 gnd.n6888 gnd.n6887 8.92286
R13667 gnd.n6964 gnd.t65 8.92286
R13668 gnd.n6980 gnd.n855 8.92286
R13669 gnd.t151 gnd.n840 8.92286
R13670 gnd.n5181 gnd.n5156 8.92171
R13671 gnd.n5149 gnd.n5124 8.92171
R13672 gnd.n5117 gnd.n5092 8.92171
R13673 gnd.n5086 gnd.n5061 8.92171
R13674 gnd.n5054 gnd.n5029 8.92171
R13675 gnd.n5022 gnd.n4997 8.92171
R13676 gnd.n4990 gnd.n4965 8.92171
R13677 gnd.n4959 gnd.n4934 8.92171
R13678 gnd.n6530 gnd.n6512 8.72777
R13679 gnd.n4685 gnd.t42 8.60421
R13680 gnd.n3691 gnd.t217 8.60421
R13681 gnd.n7909 gnd.t242 8.60421
R13682 gnd.n4089 gnd.n4069 8.43656
R13683 gnd.n58 gnd.n38 8.43656
R13684 gnd.n5182 gnd.n5154 8.14595
R13685 gnd.n5150 gnd.n5122 8.14595
R13686 gnd.n5118 gnd.n5090 8.14595
R13687 gnd.n5087 gnd.n5059 8.14595
R13688 gnd.n5055 gnd.n5027 8.14595
R13689 gnd.n5023 gnd.n4995 8.14595
R13690 gnd.n4991 gnd.n4963 8.14595
R13691 gnd.n4960 gnd.n4932 8.14595
R13692 gnd.n3540 gnd.n0 8.10675
R13693 gnd.n7983 gnd.n7982 8.10675
R13694 gnd.n5187 gnd.n5186 7.97301
R13695 gnd.t31 gnd.n4200 7.9669
R13696 gnd.n5738 gnd.n1456 7.9669
R13697 gnd.n7078 gnd.n7077 7.9669
R13698 gnd.n7983 gnd.n98 7.95236
R13699 gnd.n7110 gnd.n735 7.75808
R13700 gnd.n6155 gnd.n1239 7.75808
R13701 gnd.n7722 gnd.n7669 7.75808
R13702 gnd.n3471 gnd.n3470 7.75808
R13703 gnd.n5357 gnd.n1768 7.64824
R13704 gnd.n3605 gnd.n3604 7.64824
R13705 gnd.n5366 gnd.n1740 7.64824
R13706 gnd.n5392 gnd.n1743 7.64824
R13707 gnd.n5374 gnd.n5373 7.64824
R13708 gnd.n5402 gnd.n1732 7.64824
R13709 gnd.n5385 gnd.n5384 7.64824
R13710 gnd.n5411 gnd.n1702 7.64824
R13711 gnd.n5442 gnd.n1705 7.64824
R13712 gnd.n5424 gnd.n5423 7.64824
R13713 gnd.n5452 gnd.n1694 7.64824
R13714 gnd.n5435 gnd.n5434 7.64824
R13715 gnd.n1716 gnd.n1714 7.64824
R13716 gnd.n5477 gnd.n1670 7.64824
R13717 gnd.n5486 gnd.n1658 7.64824
R13718 gnd.n5485 gnd.n1661 7.64824
R13719 gnd.n5468 gnd.n1637 7.64824
R13720 gnd.n5545 gnd.n1640 7.64824
R13721 gnd.n1680 gnd.n1627 7.64824
R13722 gnd.n5555 gnd.n1629 7.64824
R13723 gnd.n5538 gnd.n5537 7.64824
R13724 gnd.n5577 gnd.n1611 7.64824
R13725 gnd.n5585 gnd.n1614 7.64824
R13726 gnd.n5561 gnd.n1601 7.64824
R13727 gnd.n5595 gnd.n1603 7.64824
R13728 gnd.n5603 gnd.n1243 7.64824
R13729 gnd.n6152 gnd.n1245 7.64824
R13730 gnd.n6244 gnd.n1160 7.64824
R13731 gnd.n5934 gnd.n5815 7.64824
R13732 gnd.n1062 gnd.t1 7.64824
R13733 gnd.n6364 gnd.n1055 7.64824
R13734 gnd.n6462 gnd.n995 7.64824
R13735 gnd.n6432 gnd.t66 7.64824
R13736 gnd.n6880 gnd.n946 7.64824
R13737 gnd.n7310 gnd.n551 7.64824
R13738 gnd.n7302 gnd.n554 7.64824
R13739 gnd.n559 gnd.n544 7.64824
R13740 gnd.n7329 gnd.n536 7.64824
R13741 gnd.n7352 gnd.n522 7.64824
R13742 gnd.n7333 gnd.n525 7.64824
R13743 gnd.n7362 gnd.n512 7.64824
R13744 gnd.n514 gnd.n504 7.64824
R13745 gnd.n7372 gnd.n7371 7.64824
R13746 gnd.n7401 gnd.n486 7.64824
R13747 gnd.n7338 gnd.n489 7.64824
R13748 gnd.n7411 gnd.n477 7.64824
R13749 gnd.n7394 gnd.n7393 7.64824
R13750 gnd.n7420 gnd.n470 7.64824
R13751 gnd.n7438 gnd.n456 7.64824
R13752 gnd.n7424 gnd.n459 7.64824
R13753 gnd.n7448 gnd.n446 7.64824
R13754 gnd.n448 gnd.n438 7.64824
R13755 gnd.n7458 gnd.n7457 7.64824
R13756 gnd.n7486 gnd.n421 7.64824
R13757 gnd.n7471 gnd.n7470 7.64824
R13758 gnd.n7497 gnd.n411 7.64824
R13759 gnd.n413 gnd.n403 7.64824
R13760 gnd.n7509 gnd.n7508 7.64824
R13761 gnd.n7536 gnd.n383 7.64824
R13762 gnd.n7519 gnd.n394 7.64824
R13763 gnd.n7518 gnd.n376 7.64824
R13764 gnd.n4130 gnd.n4129 7.53171
R13765 gnd.n4594 gnd.t16 7.32958
R13766 gnd.n6172 gnd.t135 7.32958
R13767 gnd.n1196 gnd.t10 7.32958
R13768 gnd.t6 gnd.n1160 7.32958
R13769 gnd.n6660 gnd.t414 7.32958
R13770 gnd.t81 gnd.n813 7.32958
R13771 gnd.n7063 gnd.t99 7.32958
R13772 gnd.n7921 gnd.n201 7.32958
R13773 gnd.n1346 gnd.n1345 7.30353
R13774 gnd.n6529 gnd.n6528 7.30353
R13775 gnd.n4554 gnd.n4273 7.01093
R13776 gnd.n4276 gnd.n4274 7.01093
R13777 gnd.n4564 gnd.n4563 7.01093
R13778 gnd.n4575 gnd.n4257 7.01093
R13779 gnd.n4574 gnd.n4260 7.01093
R13780 gnd.n4585 gnd.n4248 7.01093
R13781 gnd.n4251 gnd.n4249 7.01093
R13782 gnd.n4595 gnd.n4594 7.01093
R13783 gnd.n4605 gnd.n4229 7.01093
R13784 gnd.n4604 gnd.n4232 7.01093
R13785 gnd.n4613 gnd.n4223 7.01093
R13786 gnd.n4625 gnd.n4213 7.01093
R13787 gnd.n4635 gnd.n4198 7.01093
R13788 gnd.n4651 gnd.n4650 7.01093
R13789 gnd.n4200 gnd.n4137 7.01093
R13790 gnd.n4705 gnd.n4138 7.01093
R13791 gnd.n4699 gnd.n4698 7.01093
R13792 gnd.n4187 gnd.n4149 7.01093
R13793 gnd.n4691 gnd.n4160 7.01093
R13794 gnd.n4178 gnd.n4173 7.01093
R13795 gnd.n4685 gnd.n4684 7.01093
R13796 gnd.n4731 gnd.n4044 7.01093
R13797 gnd.n4730 gnd.n4729 7.01093
R13798 gnd.n4742 gnd.n4741 7.01093
R13799 gnd.n4037 gnd.n4029 7.01093
R13800 gnd.n4771 gnd.n4017 7.01093
R13801 gnd.n4770 gnd.n4020 7.01093
R13802 gnd.n4781 gnd.n4009 7.01093
R13803 gnd.n4010 gnd.n3998 7.01093
R13804 gnd.n4792 gnd.n3999 7.01093
R13805 gnd.n4816 gnd.n3990 7.01093
R13806 gnd.n4815 gnd.n3981 7.01093
R13807 gnd.n4838 gnd.n4837 7.01093
R13808 gnd.n4856 gnd.n3962 7.01093
R13809 gnd.n4855 gnd.n3965 7.01093
R13810 gnd.n4866 gnd.n3954 7.01093
R13811 gnd.n3955 gnd.n3942 7.01093
R13812 gnd.n4877 gnd.n3943 7.01093
R13813 gnd.n4904 gnd.n3927 7.01093
R13814 gnd.n4916 gnd.n4915 7.01093
R13815 gnd.n4898 gnd.n3920 7.01093
R13816 gnd.n4927 gnd.n4926 7.01093
R13817 gnd.n5199 gnd.n3908 7.01093
R13818 gnd.n5198 gnd.n3911 7.01093
R13819 gnd.n5211 gnd.n3900 7.01093
R13820 gnd.n3901 gnd.n3893 7.01093
R13821 gnd.n5221 gnd.n3149 7.01093
R13822 gnd.n6276 gnd.t39 7.01093
R13823 gnd.t47 gnd.n1071 7.01093
R13824 gnd.n6441 gnd.t46 7.01093
R13825 gnd.n6956 gnd.t29 7.01093
R13826 gnd.n4232 gnd.t41 6.69227
R13827 gnd.n4020 gnd.t407 6.69227
R13828 gnd.n4905 gnd.t43 6.69227
R13829 gnd.n5969 gnd.t73 6.69227
R13830 gnd.t55 gnd.n1003 6.69227
R13831 gnd.n6720 gnd.n6719 6.5566
R13832 gnd.n6093 gnd.n6092 6.5566
R13833 gnd.n1370 gnd.n1364 6.5566
R13834 gnd.n6735 gnd.n6734 6.5566
R13835 gnd.n6236 gnd.n1167 6.37362
R13836 gnd.t174 gnd.t157 6.37362
R13837 gnd.n5926 gnd.n5821 6.37362
R13838 gnd.n6332 gnd.t28 6.37362
R13839 gnd.n6404 gnd.n1032 6.37362
R13840 gnd.n6395 gnd.n6394 6.37362
R13841 gnd.n6900 gnd.t36 6.37362
R13842 gnd.n6873 gnd.n6872 6.37362
R13843 gnd.n6980 gnd.t88 6.37362
R13844 gnd.n6654 gnd.t88 6.37362
R13845 gnd.n6996 gnd.n840 6.37362
R13846 gnd.n5675 gnd.n5672 6.20656
R13847 gnd.n737 gnd.n731 6.20656
R13848 gnd.t44 gnd.n4661 6.05496
R13849 gnd.n4662 gnd.t14 6.05496
R13850 gnd.t59 gnd.n4044 6.05496
R13851 gnd.t54 gnd.n4826 6.05496
R13852 gnd.n5822 gnd.t71 6.05496
R13853 gnd.t48 gnd.t413 6.05496
R13854 gnd.t2 gnd.t52 6.05496
R13855 gnd.n6871 gnd.t32 6.05496
R13856 gnd.n5184 gnd.n5154 5.81868
R13857 gnd.n5152 gnd.n5122 5.81868
R13858 gnd.n5120 gnd.n5090 5.81868
R13859 gnd.n5089 gnd.n5059 5.81868
R13860 gnd.n5057 gnd.n5027 5.81868
R13861 gnd.n5025 gnd.n4995 5.81868
R13862 gnd.n4993 gnd.n4963 5.81868
R13863 gnd.n4962 gnd.n4932 5.81868
R13864 gnd.t103 gnd.n864 5.73631
R13865 gnd.n6557 gnd.n639 5.62001
R13866 gnd.n6100 gnd.n1301 5.62001
R13867 gnd.n6100 gnd.n1302 5.62001
R13868 gnd.n6729 gnd.n639 5.62001
R13869 gnd.n4413 gnd.n4408 5.4308
R13870 gnd.n5229 gnd.n3886 5.4308
R13871 gnd.n4729 gnd.t30 5.41765
R13872 gnd.t67 gnd.n4752 5.41765
R13873 gnd.t77 gnd.n3974 5.41765
R13874 gnd.n6284 gnd.t3 5.09899
R13875 gnd.n5828 gnd.n5827 5.09899
R13876 gnd.n6383 gnd.n1044 5.09899
R13877 gnd.n6414 gnd.n1023 5.09899
R13878 gnd.n6865 gnd.n962 5.09899
R13879 gnd.n6948 gnd.t25 5.09899
R13880 gnd.n5182 gnd.n5181 5.04292
R13881 gnd.n5150 gnd.n5149 5.04292
R13882 gnd.n5118 gnd.n5117 5.04292
R13883 gnd.n5087 gnd.n5086 5.04292
R13884 gnd.n5055 gnd.n5054 5.04292
R13885 gnd.n5023 gnd.n5022 5.04292
R13886 gnd.n4991 gnd.n4990 5.04292
R13887 gnd.n4960 gnd.n4959 5.04292
R13888 gnd.n4692 gnd.t15 4.78034
R13889 gnd.n3999 gnd.t69 4.78034
R13890 gnd.n6228 gnd.t85 4.78034
R13891 gnd.n6532 gnd.t128 4.78034
R13892 gnd.n7004 gnd.t75 4.78034
R13893 gnd.n4134 gnd.n4131 4.74817
R13894 gnd.n4184 gnd.n4050 4.74817
R13895 gnd.n4171 gnd.n4049 4.74817
R13896 gnd.n4048 gnd.n4047 4.74817
R13897 gnd.n4180 gnd.n4131 4.74817
R13898 gnd.n4181 gnd.n4050 4.74817
R13899 gnd.n4183 gnd.n4049 4.74817
R13900 gnd.n4170 gnd.n4048 4.74817
R13901 gnd.n7543 gnd.n117 4.74817
R13902 gnd.n7558 gnd.n116 4.74817
R13903 gnd.n7556 gnd.n115 4.74817
R13904 gnd.n7975 gnd.n110 4.74817
R13905 gnd.n7973 gnd.n111 4.74817
R13906 gnd.n7540 gnd.n117 4.74817
R13907 gnd.n7542 gnd.n116 4.74817
R13908 gnd.n7559 gnd.n115 4.74817
R13909 gnd.n7555 gnd.n110 4.74817
R13910 gnd.n7974 gnd.n7973 4.74817
R13911 gnd.n5351 gnd.n5350 4.74817
R13912 gnd.n5338 gnd.n1778 4.74817
R13913 gnd.n5336 gnd.n1777 4.74817
R13914 gnd.n5324 gnd.n1776 4.74817
R13915 gnd.n1775 gnd.n1772 4.74817
R13916 gnd.n5351 gnd.n1779 4.74817
R13917 gnd.n5349 gnd.n1778 4.74817
R13918 gnd.n5339 gnd.n1777 4.74817
R13919 gnd.n5335 gnd.n1776 4.74817
R13920 gnd.n5325 gnd.n1775 4.74817
R13921 gnd.n4129 gnd.n4128 4.74296
R13922 gnd.n98 gnd.n97 4.74296
R13923 gnd.n4089 gnd.n4088 4.7074
R13924 gnd.n4109 gnd.n4108 4.7074
R13925 gnd.n58 gnd.n57 4.7074
R13926 gnd.n78 gnd.n77 4.7074
R13927 gnd.n4129 gnd.n4109 4.65959
R13928 gnd.n98 gnd.n78 4.65959
R13929 gnd.n7222 gnd.n641 4.6132
R13930 gnd.n6101 gnd.n1300 4.6132
R13931 gnd.n6324 gnd.t0 4.46168
R13932 gnd.n6908 gnd.t9 4.46168
R13933 gnd.n6988 gnd.t202 4.46168
R13934 gnd.n6525 gnd.n6512 4.46111
R13935 gnd.n5167 gnd.n5163 4.38594
R13936 gnd.n5135 gnd.n5131 4.38594
R13937 gnd.n5103 gnd.n5099 4.38594
R13938 gnd.n5072 gnd.n5068 4.38594
R13939 gnd.n5040 gnd.n5036 4.38594
R13940 gnd.n5008 gnd.n5004 4.38594
R13941 gnd.n4976 gnd.n4972 4.38594
R13942 gnd.n4945 gnd.n4941 4.38594
R13943 gnd.n5178 gnd.n5156 4.26717
R13944 gnd.n5146 gnd.n5124 4.26717
R13945 gnd.n5114 gnd.n5092 4.26717
R13946 gnd.n5083 gnd.n5061 4.26717
R13947 gnd.n5051 gnd.n5029 4.26717
R13948 gnd.n5019 gnd.n4997 4.26717
R13949 gnd.n4987 gnd.n4965 4.26717
R13950 gnd.n4956 gnd.n4934 4.26717
R13951 gnd.n4636 gnd.t17 4.14303
R13952 gnd.n4866 gnd.t40 4.14303
R13953 gnd.t124 gnd.n1595 4.14303
R13954 gnd.n7301 gnd.t95 4.14303
R13955 gnd.n5186 gnd.n5185 4.08274
R13956 gnd.n6719 gnd.n6718 4.05904
R13957 gnd.n6092 gnd.n6091 4.05904
R13958 gnd.n1374 gnd.n1364 4.05904
R13959 gnd.n6736 gnd.n6735 4.05904
R13960 gnd.n19 gnd.n9 3.99943
R13961 gnd.n6030 gnd.n1324 3.82437
R13962 gnd.t157 gnd.n1151 3.82437
R13963 gnd.n5833 gnd.n5832 3.82437
R13964 gnd.n5918 gnd.t8 3.82437
R13965 gnd.n6308 gnd.n1102 3.82437
R13966 gnd.n6372 gnd.n1049 3.82437
R13967 gnd.n6424 gnd.n6423 3.82437
R13968 gnd.n6924 gnd.n905 3.82437
R13969 gnd.n961 gnd.t22 3.82437
R13970 gnd.n6858 gnd.n6857 3.82437
R13971 gnd.n6654 gnd.t106 3.82437
R13972 gnd.n6792 gnd.n6791 3.82437
R13973 gnd.n4709 gnd.n4130 3.81325
R13974 gnd.n4109 gnd.n4089 3.72967
R13975 gnd.n78 gnd.n58 3.72967
R13976 gnd.n5186 gnd.n5058 3.70378
R13977 gnd.n19 gnd.n18 3.60163
R13978 gnd.n3286 gnd.t131 3.50571
R13979 gnd.n5563 gnd.t124 3.50571
R13980 gnd.n7320 gnd.t95 3.50571
R13981 gnd.t113 gnd.n239 3.50571
R13982 gnd.n5177 gnd.n5158 3.49141
R13983 gnd.n5145 gnd.n5126 3.49141
R13984 gnd.n5113 gnd.n5094 3.49141
R13985 gnd.n5082 gnd.n5063 3.49141
R13986 gnd.n5050 gnd.n5031 3.49141
R13987 gnd.n5018 gnd.n4999 3.49141
R13988 gnd.n4986 gnd.n4967 3.49141
R13989 gnd.n4955 gnd.n4936 3.49141
R13990 gnd.n7240 gnd.n7239 3.29747
R13991 gnd.n7239 gnd.n7238 3.29747
R13992 gnd.n7850 gnd.n7847 3.29747
R13993 gnd.n7851 gnd.n7850 3.29747
R13994 gnd.n3798 gnd.n3797 3.29747
R13995 gnd.n3797 gnd.n3796 3.29747
R13996 gnd.n6117 gnd.n6116 3.29747
R13997 gnd.n6116 gnd.n6115 3.29747
R13998 gnd.n5910 gnd.t37 3.18706
R13999 gnd.n6292 gnd.t37 3.18706
R14000 gnd.n6940 gnd.t50 3.18706
R14001 gnd.n6859 gnd.t50 3.18706
R14002 gnd.n6660 gnd.t202 3.18706
R14003 gnd.n4215 gnd.t17 2.8684
R14004 gnd.n5850 gnd.t57 2.8684
R14005 gnd.n6638 gnd.t61 2.8684
R14006 gnd.n4110 gnd.t333 2.82907
R14007 gnd.n4110 gnd.t406 2.82907
R14008 gnd.n4112 gnd.t288 2.82907
R14009 gnd.n4112 gnd.t389 2.82907
R14010 gnd.n4114 gnd.t222 2.82907
R14011 gnd.n4114 gnd.t362 2.82907
R14012 gnd.n4116 gnd.t393 2.82907
R14013 gnd.n4116 gnd.t285 2.82907
R14014 gnd.n4118 gnd.t320 2.82907
R14015 gnd.n4118 gnd.t297 2.82907
R14016 gnd.n4120 gnd.t296 2.82907
R14017 gnd.n4120 gnd.t266 2.82907
R14018 gnd.n4122 gnd.t305 2.82907
R14019 gnd.n4122 gnd.t349 2.82907
R14020 gnd.n4124 gnd.t356 2.82907
R14021 gnd.n4124 gnd.t306 2.82907
R14022 gnd.n4126 gnd.t342 2.82907
R14023 gnd.n4126 gnd.t239 2.82907
R14024 gnd.n4051 gnd.t339 2.82907
R14025 gnd.n4051 gnd.t359 2.82907
R14026 gnd.n4053 gnd.t372 2.82907
R14027 gnd.n4053 gnd.t396 2.82907
R14028 gnd.n4055 gnd.t329 2.82907
R14029 gnd.n4055 gnd.t345 2.82907
R14030 gnd.n4057 gnd.t360 2.82907
R14031 gnd.n4057 gnd.t252 2.82907
R14032 gnd.n4059 gnd.t344 2.82907
R14033 gnd.n4059 gnd.t338 2.82907
R14034 gnd.n4061 gnd.t379 2.82907
R14035 gnd.n4061 gnd.t374 2.82907
R14036 gnd.n4063 gnd.t275 2.82907
R14037 gnd.n4063 gnd.t353 2.82907
R14038 gnd.n4065 gnd.t394 2.82907
R14039 gnd.n4065 gnd.t254 2.82907
R14040 gnd.n4067 gnd.t279 2.82907
R14041 gnd.n4067 gnd.t369 2.82907
R14042 gnd.n4070 gnd.t323 2.82907
R14043 gnd.n4070 gnd.t310 2.82907
R14044 gnd.n4072 gnd.t290 2.82907
R14045 gnd.n4072 gnd.t336 2.82907
R14046 gnd.n4074 gnd.t280 2.82907
R14047 gnd.n4074 gnd.t324 2.82907
R14048 gnd.n4076 gnd.t326 2.82907
R14049 gnd.n4076 gnd.t299 2.82907
R14050 gnd.n4078 gnd.t220 2.82907
R14051 gnd.n4078 gnd.t284 2.82907
R14052 gnd.n4080 gnd.t270 2.82907
R14053 gnd.n4080 gnd.t327 2.82907
R14054 gnd.n4082 gnd.t257 2.82907
R14055 gnd.n4082 gnd.t212 2.82907
R14056 gnd.n4084 gnd.t231 2.82907
R14057 gnd.n4084 gnd.t281 2.82907
R14058 gnd.n4086 gnd.t282 2.82907
R14059 gnd.n4086 gnd.t250 2.82907
R14060 gnd.n4090 gnd.t381 2.82907
R14061 gnd.n4090 gnd.t318 2.82907
R14062 gnd.n4092 gnd.t352 2.82907
R14063 gnd.n4092 gnd.t302 2.82907
R14064 gnd.n4094 gnd.t332 2.82907
R14065 gnd.n4094 gnd.t236 2.82907
R14066 gnd.n4096 gnd.t308 2.82907
R14067 gnd.n4096 gnd.t350 2.82907
R14068 gnd.n4098 gnd.t370 2.82907
R14069 gnd.n4098 gnd.t357 2.82907
R14070 gnd.n4100 gnd.t354 2.82907
R14071 gnd.n4100 gnd.t343 2.82907
R14072 gnd.n4102 gnd.t361 2.82907
R14073 gnd.n4102 gnd.t401 2.82907
R14074 gnd.n4104 gnd.t226 2.82907
R14075 gnd.n4104 gnd.t363 2.82907
R14076 gnd.n4106 gnd.t395 2.82907
R14077 gnd.n4106 gnd.t337 2.82907
R14078 gnd.n95 gnd.t348 2.82907
R14079 gnd.n95 gnd.t234 2.82907
R14080 gnd.n93 gnd.t378 2.82907
R14081 gnd.n93 gnd.t264 2.82907
R14082 gnd.n91 gnd.t312 2.82907
R14083 gnd.n91 gnd.t365 2.82907
R14084 gnd.n89 gnd.t387 2.82907
R14085 gnd.n89 gnd.t400 2.82907
R14086 gnd.n87 gnd.t403 2.82907
R14087 gnd.n87 gnd.t277 2.82907
R14088 gnd.n85 gnd.t397 2.82907
R14089 gnd.n85 gnd.t355 2.82907
R14090 gnd.n83 gnd.t330 2.82907
R14091 gnd.n83 gnd.t385 2.82907
R14092 gnd.n81 gnd.t351 2.82907
R14093 gnd.n81 gnd.t398 2.82907
R14094 gnd.n79 gnd.t368 2.82907
R14095 gnd.n79 gnd.t262 2.82907
R14096 gnd.n36 gnd.t377 2.82907
R14097 gnd.n36 gnd.t303 2.82907
R14098 gnd.n34 gnd.t272 2.82907
R14099 gnd.n34 gnd.t404 2.82907
R14100 gnd.n32 gnd.t386 2.82907
R14101 gnd.n32 gnd.t255 2.82907
R14102 gnd.n30 gnd.t214 2.82907
R14103 gnd.n30 gnd.t237 2.82907
R14104 gnd.n28 gnd.t366 2.82907
R14105 gnd.n28 gnd.t210 2.82907
R14106 gnd.n26 gnd.t319 2.82907
R14107 gnd.n26 gnd.t392 2.82907
R14108 gnd.n24 gnd.t380 2.82907
R14109 gnd.n24 gnd.t304 2.82907
R14110 gnd.n22 gnd.t274 2.82907
R14111 gnd.n22 gnd.t208 2.82907
R14112 gnd.n20 gnd.t391 2.82907
R14113 gnd.n20 gnd.t367 2.82907
R14114 gnd.n55 gnd.t390 2.82907
R14115 gnd.n55 gnd.t405 2.82907
R14116 gnd.n53 gnd.t402 2.82907
R14117 gnd.n53 gnd.t382 2.82907
R14118 gnd.n51 gnd.t373 2.82907
R14119 gnd.n51 gnd.t273 2.82907
R14120 gnd.n49 gnd.t293 2.82907
R14121 gnd.n49 gnd.t230 2.82907
R14122 gnd.n47 gnd.t241 2.82907
R14123 gnd.n47 gnd.t258 2.82907
R14124 gnd.n45 gnd.t260 2.82907
R14125 gnd.n45 gnd.t289 2.82907
R14126 gnd.n43 gnd.t292 2.82907
R14127 gnd.n43 gnd.t315 2.82907
R14128 gnd.n41 gnd.t313 2.82907
R14129 gnd.n41 gnd.t267 2.82907
R14130 gnd.n39 gnd.t268 2.82907
R14131 gnd.n39 gnd.t286 2.82907
R14132 gnd.n75 gnd.t399 2.82907
R14133 gnd.n75 gnd.t334 2.82907
R14134 gnd.n73 gnd.t276 2.82907
R14135 gnd.n73 gnd.t341 2.82907
R14136 gnd.n71 gnd.t364 2.82907
R14137 gnd.n71 gnd.t247 2.82907
R14138 gnd.n69 gnd.t298 2.82907
R14139 gnd.n69 gnd.t321 2.82907
R14140 gnd.n67 gnd.t325 2.82907
R14141 gnd.n67 gnd.t346 2.82907
R14142 gnd.n65 gnd.t316 2.82907
R14143 gnd.n65 gnd.t224 2.82907
R14144 gnd.n63 gnd.t376 2.82907
R14145 gnd.n63 gnd.t295 2.82907
R14146 gnd.n61 gnd.t216 2.82907
R14147 gnd.n61 gnd.t317 2.82907
R14148 gnd.n59 gnd.t249 2.82907
R14149 gnd.n59 gnd.t340 2.82907
R14150 gnd.n5174 gnd.n5173 2.71565
R14151 gnd.n5142 gnd.n5141 2.71565
R14152 gnd.n5110 gnd.n5109 2.71565
R14153 gnd.n5079 gnd.n5078 2.71565
R14154 gnd.n5047 gnd.n5046 2.71565
R14155 gnd.n5015 gnd.n5014 2.71565
R14156 gnd.n4983 gnd.n4982 2.71565
R14157 gnd.n4952 gnd.n4951 2.71565
R14158 gnd.n6023 gnd.n6022 2.54975
R14159 gnd.n5839 gnd.n5838 2.54975
R14160 gnd.n5902 gnd.t3 2.54975
R14161 gnd.n6316 gnd.n1095 2.54975
R14162 gnd.n6316 gnd.t51 2.54975
R14163 gnd.n6356 gnd.n1062 2.54975
R14164 gnd.n6432 gnd.n1011 2.54975
R14165 gnd.n6916 gnd.t38 2.54975
R14166 gnd.n6916 gnd.n912 2.54975
R14167 gnd.n6608 gnd.t25 2.54975
R14168 gnd.n6621 gnd.n6620 2.54975
R14169 gnd.n6653 gnd.n6652 2.54975
R14170 gnd.n4709 gnd.n4131 2.27742
R14171 gnd.n4709 gnd.n4050 2.27742
R14172 gnd.n4709 gnd.n4049 2.27742
R14173 gnd.n4709 gnd.n4048 2.27742
R14174 gnd.n7972 gnd.n117 2.27742
R14175 gnd.n7972 gnd.n116 2.27742
R14176 gnd.n7972 gnd.n115 2.27742
R14177 gnd.n7972 gnd.n110 2.27742
R14178 gnd.n7973 gnd.n7972 2.27742
R14179 gnd.n5352 gnd.n5351 2.27742
R14180 gnd.n5352 gnd.n1778 2.27742
R14181 gnd.n5352 gnd.n1777 2.27742
R14182 gnd.n5352 gnd.n1776 2.27742
R14183 gnd.n5352 gnd.n1775 2.27742
R14184 gnd.n4563 gnd.t117 2.23109
R14185 gnd.n4186 gnd.t15 2.23109
R14186 gnd.n5374 gnd.t221 2.23109
R14187 gnd.n6372 gnd.t48 2.23109
R14188 gnd.n6424 gnd.t52 2.23109
R14189 gnd.t294 gnd.n413 2.23109
R14190 gnd.n5170 gnd.n5160 1.93989
R14191 gnd.n5138 gnd.n5128 1.93989
R14192 gnd.n5106 gnd.n5096 1.93989
R14193 gnd.n5075 gnd.n5065 1.93989
R14194 gnd.n5043 gnd.n5033 1.93989
R14195 gnd.n5011 gnd.n5001 1.93989
R14196 gnd.n4979 gnd.n4969 1.93989
R14197 gnd.n4948 gnd.n4938 1.93989
R14198 gnd.n1326 gnd.t110 1.91244
R14199 gnd.n5893 gnd.t39 1.91244
R14200 gnd.n6599 gnd.t29 1.91244
R14201 gnd.t411 gnd.n4574 1.59378
R14202 gnd.n4753 gnd.t67 1.59378
R14203 gnd.n3983 gnd.t77 1.59378
R14204 gnd.t238 gnd.n3330 1.59378
R14205 gnd.n1716 gnd.t301 1.59378
R14206 gnd.t322 gnd.n5485 1.59378
R14207 gnd.n5902 gnd.t34 1.59378
R14208 gnd.t23 gnd.n5810 1.59378
R14209 gnd.n6887 gnd.t83 1.59378
R14210 gnd.n6608 gnd.t12 1.59378
R14211 gnd.n7411 gnd.t261 1.59378
R14212 gnd.t215 gnd.n456 1.59378
R14213 gnd.n198 gnd.t347 1.59378
R14214 gnd.n6236 gnd.t189 1.27512
R14215 gnd.n5874 gnd.n5863 1.27512
R14216 gnd.n5884 gnd.t19 1.27512
R14217 gnd.n5845 gnd.n5844 1.27512
R14218 gnd.n6300 gnd.t8 1.27512
R14219 gnd.n6324 gnd.n1088 1.27512
R14220 gnd.n6346 gnd.n1071 1.27512
R14221 gnd.n6441 gnd.n6440 1.27512
R14222 gnd.n6908 gnd.n919 1.27512
R14223 gnd.n6932 gnd.t22 1.27512
R14224 gnd.n6630 gnd.n6600 1.27512
R14225 gnd.n6594 gnd.t65 1.27512
R14226 gnd.n6645 gnd.n6590 1.27512
R14227 gnd.n4416 gnd.n4408 1.16414
R14228 gnd.n5232 gnd.n3886 1.16414
R14229 gnd.n5169 gnd.n5162 1.16414
R14230 gnd.n5137 gnd.n5130 1.16414
R14231 gnd.n5105 gnd.n5098 1.16414
R14232 gnd.n5074 gnd.n5067 1.16414
R14233 gnd.n5042 gnd.n5035 1.16414
R14234 gnd.n5010 gnd.n5003 1.16414
R14235 gnd.n4978 gnd.n4971 1.16414
R14236 gnd.n4947 gnd.n4940 1.16414
R14237 gnd.n7222 gnd.n7221 0.970197
R14238 gnd.n6101 gnd.n1297 0.970197
R14239 gnd.n5153 gnd.n5121 0.962709
R14240 gnd.n5185 gnd.n5153 0.962709
R14241 gnd.n5026 gnd.n4994 0.962709
R14242 gnd.n5058 gnd.n5026 0.962709
R14243 gnd.n4662 gnd.t44 0.956468
R14244 gnd.n4827 gnd.t54 0.956468
R14245 gnd.t256 gnd.n3368 0.956468
R14246 gnd.n5411 gnd.t235 0.956468
R14247 gnd.n5537 gnd.t227 0.956468
R14248 gnd.n1439 gnd.n1174 0.956468
R14249 gnd.n6532 gnd.n842 0.956468
R14250 gnd.t244 gnd.n512 0.956468
R14251 gnd.n7486 gnd.t291 0.956468
R14252 gnd.n160 gnd.t246 0.956468
R14253 gnd gnd.n0 0.70738
R14254 gnd.n2 gnd.n1 0.672012
R14255 gnd.n3 gnd.n2 0.672012
R14256 gnd.n4 gnd.n3 0.672012
R14257 gnd.n5 gnd.n4 0.672012
R14258 gnd.n6 gnd.n5 0.672012
R14259 gnd.n7 gnd.n6 0.672012
R14260 gnd.n8 gnd.n7 0.672012
R14261 gnd.n9 gnd.n8 0.672012
R14262 gnd.n11 gnd.n10 0.672012
R14263 gnd.n12 gnd.n11 0.672012
R14264 gnd.n13 gnd.n12 0.672012
R14265 gnd.n14 gnd.n13 0.672012
R14266 gnd.n15 gnd.n14 0.672012
R14267 gnd.n16 gnd.n15 0.672012
R14268 gnd.n17 gnd.n16 0.672012
R14269 gnd.n18 gnd.n17 0.672012
R14270 gnd.n5874 gnd.t142 0.637812
R14271 gnd.n6308 gnd.t27 0.637812
R14272 gnd.n6924 gnd.t26 0.637812
R14273 gnd.n7984 gnd.n7983 0.637193
R14274 gnd.n4128 gnd.n4127 0.573776
R14275 gnd.n4127 gnd.n4125 0.573776
R14276 gnd.n4125 gnd.n4123 0.573776
R14277 gnd.n4123 gnd.n4121 0.573776
R14278 gnd.n4121 gnd.n4119 0.573776
R14279 gnd.n4119 gnd.n4117 0.573776
R14280 gnd.n4117 gnd.n4115 0.573776
R14281 gnd.n4115 gnd.n4113 0.573776
R14282 gnd.n4113 gnd.n4111 0.573776
R14283 gnd.n4069 gnd.n4068 0.573776
R14284 gnd.n4068 gnd.n4066 0.573776
R14285 gnd.n4066 gnd.n4064 0.573776
R14286 gnd.n4064 gnd.n4062 0.573776
R14287 gnd.n4062 gnd.n4060 0.573776
R14288 gnd.n4060 gnd.n4058 0.573776
R14289 gnd.n4058 gnd.n4056 0.573776
R14290 gnd.n4056 gnd.n4054 0.573776
R14291 gnd.n4054 gnd.n4052 0.573776
R14292 gnd.n4088 gnd.n4087 0.573776
R14293 gnd.n4087 gnd.n4085 0.573776
R14294 gnd.n4085 gnd.n4083 0.573776
R14295 gnd.n4083 gnd.n4081 0.573776
R14296 gnd.n4081 gnd.n4079 0.573776
R14297 gnd.n4079 gnd.n4077 0.573776
R14298 gnd.n4077 gnd.n4075 0.573776
R14299 gnd.n4075 gnd.n4073 0.573776
R14300 gnd.n4073 gnd.n4071 0.573776
R14301 gnd.n4108 gnd.n4107 0.573776
R14302 gnd.n4107 gnd.n4105 0.573776
R14303 gnd.n4105 gnd.n4103 0.573776
R14304 gnd.n4103 gnd.n4101 0.573776
R14305 gnd.n4101 gnd.n4099 0.573776
R14306 gnd.n4099 gnd.n4097 0.573776
R14307 gnd.n4097 gnd.n4095 0.573776
R14308 gnd.n4095 gnd.n4093 0.573776
R14309 gnd.n4093 gnd.n4091 0.573776
R14310 gnd.n82 gnd.n80 0.573776
R14311 gnd.n84 gnd.n82 0.573776
R14312 gnd.n86 gnd.n84 0.573776
R14313 gnd.n88 gnd.n86 0.573776
R14314 gnd.n90 gnd.n88 0.573776
R14315 gnd.n92 gnd.n90 0.573776
R14316 gnd.n94 gnd.n92 0.573776
R14317 gnd.n96 gnd.n94 0.573776
R14318 gnd.n97 gnd.n96 0.573776
R14319 gnd.n23 gnd.n21 0.573776
R14320 gnd.n25 gnd.n23 0.573776
R14321 gnd.n27 gnd.n25 0.573776
R14322 gnd.n29 gnd.n27 0.573776
R14323 gnd.n31 gnd.n29 0.573776
R14324 gnd.n33 gnd.n31 0.573776
R14325 gnd.n35 gnd.n33 0.573776
R14326 gnd.n37 gnd.n35 0.573776
R14327 gnd.n38 gnd.n37 0.573776
R14328 gnd.n42 gnd.n40 0.573776
R14329 gnd.n44 gnd.n42 0.573776
R14330 gnd.n46 gnd.n44 0.573776
R14331 gnd.n48 gnd.n46 0.573776
R14332 gnd.n50 gnd.n48 0.573776
R14333 gnd.n52 gnd.n50 0.573776
R14334 gnd.n54 gnd.n52 0.573776
R14335 gnd.n56 gnd.n54 0.573776
R14336 gnd.n57 gnd.n56 0.573776
R14337 gnd.n62 gnd.n60 0.573776
R14338 gnd.n64 gnd.n62 0.573776
R14339 gnd.n66 gnd.n64 0.573776
R14340 gnd.n68 gnd.n66 0.573776
R14341 gnd.n70 gnd.n68 0.573776
R14342 gnd.n72 gnd.n70 0.573776
R14343 gnd.n74 gnd.n72 0.573776
R14344 gnd.n76 gnd.n74 0.573776
R14345 gnd.n77 gnd.n76 0.573776
R14346 gnd.n4889 gnd.n3890 0.486781
R14347 gnd.n4465 gnd.n4464 0.48678
R14348 gnd.n5206 gnd.n3844 0.480683
R14349 gnd.n4549 gnd.n4548 0.480683
R14350 gnd.n2944 gnd.n2943 0.480683
R14351 gnd.n2606 gnd.n2605 0.480683
R14352 gnd.n7721 gnd.n7666 0.477634
R14353 gnd.n3473 gnd.n3472 0.477634
R14354 gnd.n7098 gnd.n7097 0.451719
R14355 gnd.n6161 gnd.n6160 0.451719
R14356 gnd.n5743 gnd.n5742 0.451719
R14357 gnd.n7091 gnd.n7090 0.451719
R14358 gnd.n7887 gnd.n7886 0.442573
R14359 gnd.n7313 gnd.n549 0.442573
R14360 gnd.n6149 gnd.n6148 0.442573
R14361 gnd.n3280 gnd.n3206 0.442573
R14362 gnd.n7972 gnd.n114 0.420375
R14363 gnd.n5352 gnd.n1774 0.420375
R14364 gnd.n5684 gnd.n5672 0.388379
R14365 gnd.n5166 gnd.n5165 0.388379
R14366 gnd.n5134 gnd.n5133 0.388379
R14367 gnd.n5102 gnd.n5101 0.388379
R14368 gnd.n5071 gnd.n5070 0.388379
R14369 gnd.n5039 gnd.n5038 0.388379
R14370 gnd.n5007 gnd.n5006 0.388379
R14371 gnd.n4975 gnd.n4974 0.388379
R14372 gnd.n4944 gnd.n4943 0.388379
R14373 gnd.n7114 gnd.n731 0.388379
R14374 gnd.n7984 gnd.n19 0.374463
R14375 gnd gnd.n7984 0.367492
R14376 gnd.n3945 gnd.t43 0.319156
R14377 gnd.n3548 gnd.t265 0.319156
R14378 gnd.t307 gnd.n1766 0.319156
R14379 gnd.n7545 gnd.t223 0.319156
R14380 gnd.n121 gnd.t213 0.319156
R14381 gnd.n4383 gnd.n4361 0.311721
R14382 gnd.n7763 gnd.n352 0.293183
R14383 gnd.n3714 gnd.n3270 0.293183
R14384 gnd.n2435 gnd.n114 0.282512
R14385 gnd.n5320 gnd.n1774 0.282512
R14386 gnd.n5277 gnd.n5276 0.268793
R14387 gnd.n7764 gnd.n7763 0.258122
R14388 gnd.n7160 gnd.n7159 0.258122
R14389 gnd.n5608 gnd.n1590 0.258122
R14390 gnd.n3715 gnd.n3714 0.258122
R14391 gnd.n5566 gnd.n1233 0.247451
R14392 gnd.n7101 gnd.n7100 0.247451
R14393 gnd.n5276 gnd.n5275 0.241354
R14394 gnd.n641 gnd.n638 0.229039
R14395 gnd.n642 gnd.n641 0.229039
R14396 gnd.n1300 gnd.n1296 0.229039
R14397 gnd.n1511 gnd.n1300 0.229039
R14398 gnd.n4130 gnd.n0 0.210825
R14399 gnd.n4537 gnd.n4336 0.206293
R14400 gnd.n7515 gnd.n114 0.198671
R14401 gnd.n3599 gnd.n1774 0.198671
R14402 gnd.n5183 gnd.n5155 0.155672
R14403 gnd.n5176 gnd.n5155 0.155672
R14404 gnd.n5176 gnd.n5175 0.155672
R14405 gnd.n5175 gnd.n5159 0.155672
R14406 gnd.n5168 gnd.n5159 0.155672
R14407 gnd.n5168 gnd.n5167 0.155672
R14408 gnd.n5151 gnd.n5123 0.155672
R14409 gnd.n5144 gnd.n5123 0.155672
R14410 gnd.n5144 gnd.n5143 0.155672
R14411 gnd.n5143 gnd.n5127 0.155672
R14412 gnd.n5136 gnd.n5127 0.155672
R14413 gnd.n5136 gnd.n5135 0.155672
R14414 gnd.n5119 gnd.n5091 0.155672
R14415 gnd.n5112 gnd.n5091 0.155672
R14416 gnd.n5112 gnd.n5111 0.155672
R14417 gnd.n5111 gnd.n5095 0.155672
R14418 gnd.n5104 gnd.n5095 0.155672
R14419 gnd.n5104 gnd.n5103 0.155672
R14420 gnd.n5088 gnd.n5060 0.155672
R14421 gnd.n5081 gnd.n5060 0.155672
R14422 gnd.n5081 gnd.n5080 0.155672
R14423 gnd.n5080 gnd.n5064 0.155672
R14424 gnd.n5073 gnd.n5064 0.155672
R14425 gnd.n5073 gnd.n5072 0.155672
R14426 gnd.n5056 gnd.n5028 0.155672
R14427 gnd.n5049 gnd.n5028 0.155672
R14428 gnd.n5049 gnd.n5048 0.155672
R14429 gnd.n5048 gnd.n5032 0.155672
R14430 gnd.n5041 gnd.n5032 0.155672
R14431 gnd.n5041 gnd.n5040 0.155672
R14432 gnd.n5024 gnd.n4996 0.155672
R14433 gnd.n5017 gnd.n4996 0.155672
R14434 gnd.n5017 gnd.n5016 0.155672
R14435 gnd.n5016 gnd.n5000 0.155672
R14436 gnd.n5009 gnd.n5000 0.155672
R14437 gnd.n5009 gnd.n5008 0.155672
R14438 gnd.n4992 gnd.n4964 0.155672
R14439 gnd.n4985 gnd.n4964 0.155672
R14440 gnd.n4985 gnd.n4984 0.155672
R14441 gnd.n4984 gnd.n4968 0.155672
R14442 gnd.n4977 gnd.n4968 0.155672
R14443 gnd.n4977 gnd.n4976 0.155672
R14444 gnd.n4961 gnd.n4933 0.155672
R14445 gnd.n4954 gnd.n4933 0.155672
R14446 gnd.n4954 gnd.n4953 0.155672
R14447 gnd.n4953 gnd.n4937 0.155672
R14448 gnd.n4946 gnd.n4937 0.155672
R14449 gnd.n4946 gnd.n4945 0.155672
R14450 gnd.n5308 gnd.n3844 0.152939
R14451 gnd.n5308 gnd.n5307 0.152939
R14452 gnd.n5307 gnd.n5306 0.152939
R14453 gnd.n5306 gnd.n3846 0.152939
R14454 gnd.n3847 gnd.n3846 0.152939
R14455 gnd.n3848 gnd.n3847 0.152939
R14456 gnd.n3849 gnd.n3848 0.152939
R14457 gnd.n3850 gnd.n3849 0.152939
R14458 gnd.n3851 gnd.n3850 0.152939
R14459 gnd.n3852 gnd.n3851 0.152939
R14460 gnd.n3853 gnd.n3852 0.152939
R14461 gnd.n3854 gnd.n3853 0.152939
R14462 gnd.n3855 gnd.n3854 0.152939
R14463 gnd.n3856 gnd.n3855 0.152939
R14464 gnd.n5278 gnd.n3856 0.152939
R14465 gnd.n5278 gnd.n5277 0.152939
R14466 gnd.n4550 gnd.n4549 0.152939
R14467 gnd.n4550 gnd.n4254 0.152939
R14468 gnd.n4578 gnd.n4254 0.152939
R14469 gnd.n4579 gnd.n4578 0.152939
R14470 gnd.n4580 gnd.n4579 0.152939
R14471 gnd.n4581 gnd.n4580 0.152939
R14472 gnd.n4581 gnd.n4226 0.152939
R14473 gnd.n4608 gnd.n4226 0.152939
R14474 gnd.n4609 gnd.n4608 0.152939
R14475 gnd.n4610 gnd.n4609 0.152939
R14476 gnd.n4610 gnd.n4204 0.152939
R14477 gnd.n4639 gnd.n4204 0.152939
R14478 gnd.n4640 gnd.n4639 0.152939
R14479 gnd.n4641 gnd.n4640 0.152939
R14480 gnd.n4642 gnd.n4641 0.152939
R14481 gnd.n4644 gnd.n4642 0.152939
R14482 gnd.n4644 gnd.n4643 0.152939
R14483 gnd.n4643 gnd.n4153 0.152939
R14484 gnd.n4154 gnd.n4153 0.152939
R14485 gnd.n4155 gnd.n4154 0.152939
R14486 gnd.n4174 gnd.n4155 0.152939
R14487 gnd.n4175 gnd.n4174 0.152939
R14488 gnd.n4175 gnd.n4041 0.152939
R14489 gnd.n4734 gnd.n4041 0.152939
R14490 gnd.n4735 gnd.n4734 0.152939
R14491 gnd.n4736 gnd.n4735 0.152939
R14492 gnd.n4737 gnd.n4736 0.152939
R14493 gnd.n4737 gnd.n4014 0.152939
R14494 gnd.n4774 gnd.n4014 0.152939
R14495 gnd.n4775 gnd.n4774 0.152939
R14496 gnd.n4776 gnd.n4775 0.152939
R14497 gnd.n4777 gnd.n4776 0.152939
R14498 gnd.n4777 gnd.n3987 0.152939
R14499 gnd.n4819 gnd.n3987 0.152939
R14500 gnd.n4820 gnd.n4819 0.152939
R14501 gnd.n4821 gnd.n4820 0.152939
R14502 gnd.n4822 gnd.n4821 0.152939
R14503 gnd.n4822 gnd.n3959 0.152939
R14504 gnd.n4859 gnd.n3959 0.152939
R14505 gnd.n4860 gnd.n4859 0.152939
R14506 gnd.n4861 gnd.n4860 0.152939
R14507 gnd.n4862 gnd.n4861 0.152939
R14508 gnd.n4862 gnd.n3932 0.152939
R14509 gnd.n4908 gnd.n3932 0.152939
R14510 gnd.n4909 gnd.n4908 0.152939
R14511 gnd.n4910 gnd.n4909 0.152939
R14512 gnd.n4911 gnd.n4910 0.152939
R14513 gnd.n4911 gnd.n3905 0.152939
R14514 gnd.n5202 gnd.n3905 0.152939
R14515 gnd.n5203 gnd.n5202 0.152939
R14516 gnd.n5204 gnd.n5203 0.152939
R14517 gnd.n5205 gnd.n5204 0.152939
R14518 gnd.n5206 gnd.n5205 0.152939
R14519 gnd.n4548 gnd.n4278 0.152939
R14520 gnd.n4299 gnd.n4278 0.152939
R14521 gnd.n4300 gnd.n4299 0.152939
R14522 gnd.n4306 gnd.n4300 0.152939
R14523 gnd.n4307 gnd.n4306 0.152939
R14524 gnd.n4308 gnd.n4307 0.152939
R14525 gnd.n4308 gnd.n4297 0.152939
R14526 gnd.n4316 gnd.n4297 0.152939
R14527 gnd.n4317 gnd.n4316 0.152939
R14528 gnd.n4318 gnd.n4317 0.152939
R14529 gnd.n4318 gnd.n4295 0.152939
R14530 gnd.n4326 gnd.n4295 0.152939
R14531 gnd.n4327 gnd.n4326 0.152939
R14532 gnd.n4328 gnd.n4327 0.152939
R14533 gnd.n4328 gnd.n4293 0.152939
R14534 gnd.n4336 gnd.n4293 0.152939
R14535 gnd.n5275 gnd.n3861 0.152939
R14536 gnd.n3863 gnd.n3861 0.152939
R14537 gnd.n3864 gnd.n3863 0.152939
R14538 gnd.n3865 gnd.n3864 0.152939
R14539 gnd.n3866 gnd.n3865 0.152939
R14540 gnd.n3867 gnd.n3866 0.152939
R14541 gnd.n3868 gnd.n3867 0.152939
R14542 gnd.n3869 gnd.n3868 0.152939
R14543 gnd.n3870 gnd.n3869 0.152939
R14544 gnd.n3871 gnd.n3870 0.152939
R14545 gnd.n3872 gnd.n3871 0.152939
R14546 gnd.n3873 gnd.n3872 0.152939
R14547 gnd.n3874 gnd.n3873 0.152939
R14548 gnd.n3875 gnd.n3874 0.152939
R14549 gnd.n3876 gnd.n3875 0.152939
R14550 gnd.n3877 gnd.n3876 0.152939
R14551 gnd.n3878 gnd.n3877 0.152939
R14552 gnd.n3879 gnd.n3878 0.152939
R14553 gnd.n3880 gnd.n3879 0.152939
R14554 gnd.n3881 gnd.n3880 0.152939
R14555 gnd.n3882 gnd.n3881 0.152939
R14556 gnd.n3883 gnd.n3882 0.152939
R14557 gnd.n3887 gnd.n3883 0.152939
R14558 gnd.n3888 gnd.n3887 0.152939
R14559 gnd.n3889 gnd.n3888 0.152939
R14560 gnd.n3890 gnd.n3889 0.152939
R14561 gnd.n4711 gnd.n4710 0.152939
R14562 gnd.n4712 gnd.n4711 0.152939
R14563 gnd.n4713 gnd.n4712 0.152939
R14564 gnd.n4714 gnd.n4713 0.152939
R14565 gnd.n4715 gnd.n4714 0.152939
R14566 gnd.n4716 gnd.n4715 0.152939
R14567 gnd.n4716 gnd.n3995 0.152939
R14568 gnd.n4795 gnd.n3995 0.152939
R14569 gnd.n4796 gnd.n4795 0.152939
R14570 gnd.n4797 gnd.n4796 0.152939
R14571 gnd.n4798 gnd.n4797 0.152939
R14572 gnd.n4799 gnd.n4798 0.152939
R14573 gnd.n4800 gnd.n4799 0.152939
R14574 gnd.n4801 gnd.n4800 0.152939
R14575 gnd.n4802 gnd.n4801 0.152939
R14576 gnd.n4803 gnd.n4802 0.152939
R14577 gnd.n4803 gnd.n3939 0.152939
R14578 gnd.n4880 gnd.n3939 0.152939
R14579 gnd.n4881 gnd.n4880 0.152939
R14580 gnd.n4882 gnd.n4881 0.152939
R14581 gnd.n4883 gnd.n4882 0.152939
R14582 gnd.n4884 gnd.n4883 0.152939
R14583 gnd.n4885 gnd.n4884 0.152939
R14584 gnd.n4886 gnd.n4885 0.152939
R14585 gnd.n4887 gnd.n4886 0.152939
R14586 gnd.n4888 gnd.n4887 0.152939
R14587 gnd.n4890 gnd.n4888 0.152939
R14588 gnd.n4890 gnd.n4889 0.152939
R14589 gnd.n4466 gnd.n4465 0.152939
R14590 gnd.n4466 gnd.n4356 0.152939
R14591 gnd.n4481 gnd.n4356 0.152939
R14592 gnd.n4482 gnd.n4481 0.152939
R14593 gnd.n4483 gnd.n4482 0.152939
R14594 gnd.n4483 gnd.n4344 0.152939
R14595 gnd.n4497 gnd.n4344 0.152939
R14596 gnd.n4498 gnd.n4497 0.152939
R14597 gnd.n4499 gnd.n4498 0.152939
R14598 gnd.n4500 gnd.n4499 0.152939
R14599 gnd.n4501 gnd.n4500 0.152939
R14600 gnd.n4502 gnd.n4501 0.152939
R14601 gnd.n4503 gnd.n4502 0.152939
R14602 gnd.n4504 gnd.n4503 0.152939
R14603 gnd.n4505 gnd.n4504 0.152939
R14604 gnd.n4506 gnd.n4505 0.152939
R14605 gnd.n4507 gnd.n4506 0.152939
R14606 gnd.n4508 gnd.n4507 0.152939
R14607 gnd.n4509 gnd.n4508 0.152939
R14608 gnd.n4510 gnd.n4509 0.152939
R14609 gnd.n4511 gnd.n4510 0.152939
R14610 gnd.n4511 gnd.n4210 0.152939
R14611 gnd.n4628 gnd.n4210 0.152939
R14612 gnd.n4629 gnd.n4628 0.152939
R14613 gnd.n4630 gnd.n4629 0.152939
R14614 gnd.n4631 gnd.n4630 0.152939
R14615 gnd.n4631 gnd.n4132 0.152939
R14616 gnd.n4708 gnd.n4132 0.152939
R14617 gnd.n4384 gnd.n4383 0.152939
R14618 gnd.n4385 gnd.n4384 0.152939
R14619 gnd.n4386 gnd.n4385 0.152939
R14620 gnd.n4387 gnd.n4386 0.152939
R14621 gnd.n4388 gnd.n4387 0.152939
R14622 gnd.n4389 gnd.n4388 0.152939
R14623 gnd.n4390 gnd.n4389 0.152939
R14624 gnd.n4391 gnd.n4390 0.152939
R14625 gnd.n4392 gnd.n4391 0.152939
R14626 gnd.n4393 gnd.n4392 0.152939
R14627 gnd.n4394 gnd.n4393 0.152939
R14628 gnd.n4395 gnd.n4394 0.152939
R14629 gnd.n4396 gnd.n4395 0.152939
R14630 gnd.n4397 gnd.n4396 0.152939
R14631 gnd.n4398 gnd.n4397 0.152939
R14632 gnd.n4399 gnd.n4398 0.152939
R14633 gnd.n4400 gnd.n4399 0.152939
R14634 gnd.n4401 gnd.n4400 0.152939
R14635 gnd.n4402 gnd.n4401 0.152939
R14636 gnd.n4403 gnd.n4402 0.152939
R14637 gnd.n4404 gnd.n4403 0.152939
R14638 gnd.n4405 gnd.n4404 0.152939
R14639 gnd.n4409 gnd.n4405 0.152939
R14640 gnd.n4410 gnd.n4409 0.152939
R14641 gnd.n4410 gnd.n4367 0.152939
R14642 gnd.n4464 gnd.n4367 0.152939
R14643 gnd.n2943 gnd.n1936 0.152939
R14644 gnd.n1941 gnd.n1936 0.152939
R14645 gnd.n1942 gnd.n1941 0.152939
R14646 gnd.n1943 gnd.n1942 0.152939
R14647 gnd.n1944 gnd.n1943 0.152939
R14648 gnd.n1949 gnd.n1944 0.152939
R14649 gnd.n1950 gnd.n1949 0.152939
R14650 gnd.n1951 gnd.n1950 0.152939
R14651 gnd.n1952 gnd.n1951 0.152939
R14652 gnd.n1957 gnd.n1952 0.152939
R14653 gnd.n1958 gnd.n1957 0.152939
R14654 gnd.n1959 gnd.n1958 0.152939
R14655 gnd.n1960 gnd.n1959 0.152939
R14656 gnd.n1965 gnd.n1960 0.152939
R14657 gnd.n1966 gnd.n1965 0.152939
R14658 gnd.n1967 gnd.n1966 0.152939
R14659 gnd.n1968 gnd.n1967 0.152939
R14660 gnd.n1973 gnd.n1968 0.152939
R14661 gnd.n1974 gnd.n1973 0.152939
R14662 gnd.n1975 gnd.n1974 0.152939
R14663 gnd.n1976 gnd.n1975 0.152939
R14664 gnd.n1981 gnd.n1976 0.152939
R14665 gnd.n1982 gnd.n1981 0.152939
R14666 gnd.n1983 gnd.n1982 0.152939
R14667 gnd.n1984 gnd.n1983 0.152939
R14668 gnd.n1989 gnd.n1984 0.152939
R14669 gnd.n1990 gnd.n1989 0.152939
R14670 gnd.n1991 gnd.n1990 0.152939
R14671 gnd.n1992 gnd.n1991 0.152939
R14672 gnd.n1997 gnd.n1992 0.152939
R14673 gnd.n1998 gnd.n1997 0.152939
R14674 gnd.n1999 gnd.n1998 0.152939
R14675 gnd.n2000 gnd.n1999 0.152939
R14676 gnd.n2005 gnd.n2000 0.152939
R14677 gnd.n2006 gnd.n2005 0.152939
R14678 gnd.n2007 gnd.n2006 0.152939
R14679 gnd.n2008 gnd.n2007 0.152939
R14680 gnd.n2013 gnd.n2008 0.152939
R14681 gnd.n2014 gnd.n2013 0.152939
R14682 gnd.n2015 gnd.n2014 0.152939
R14683 gnd.n2016 gnd.n2015 0.152939
R14684 gnd.n2021 gnd.n2016 0.152939
R14685 gnd.n2022 gnd.n2021 0.152939
R14686 gnd.n2023 gnd.n2022 0.152939
R14687 gnd.n2024 gnd.n2023 0.152939
R14688 gnd.n2029 gnd.n2024 0.152939
R14689 gnd.n2030 gnd.n2029 0.152939
R14690 gnd.n2031 gnd.n2030 0.152939
R14691 gnd.n2032 gnd.n2031 0.152939
R14692 gnd.n2037 gnd.n2032 0.152939
R14693 gnd.n2038 gnd.n2037 0.152939
R14694 gnd.n2039 gnd.n2038 0.152939
R14695 gnd.n2040 gnd.n2039 0.152939
R14696 gnd.n2045 gnd.n2040 0.152939
R14697 gnd.n2046 gnd.n2045 0.152939
R14698 gnd.n2047 gnd.n2046 0.152939
R14699 gnd.n2048 gnd.n2047 0.152939
R14700 gnd.n2053 gnd.n2048 0.152939
R14701 gnd.n2054 gnd.n2053 0.152939
R14702 gnd.n2055 gnd.n2054 0.152939
R14703 gnd.n2056 gnd.n2055 0.152939
R14704 gnd.n2061 gnd.n2056 0.152939
R14705 gnd.n2062 gnd.n2061 0.152939
R14706 gnd.n2063 gnd.n2062 0.152939
R14707 gnd.n2064 gnd.n2063 0.152939
R14708 gnd.n2069 gnd.n2064 0.152939
R14709 gnd.n2070 gnd.n2069 0.152939
R14710 gnd.n2071 gnd.n2070 0.152939
R14711 gnd.n2072 gnd.n2071 0.152939
R14712 gnd.n2077 gnd.n2072 0.152939
R14713 gnd.n2078 gnd.n2077 0.152939
R14714 gnd.n2079 gnd.n2078 0.152939
R14715 gnd.n2080 gnd.n2079 0.152939
R14716 gnd.n2085 gnd.n2080 0.152939
R14717 gnd.n2086 gnd.n2085 0.152939
R14718 gnd.n2087 gnd.n2086 0.152939
R14719 gnd.n2088 gnd.n2087 0.152939
R14720 gnd.n2093 gnd.n2088 0.152939
R14721 gnd.n2094 gnd.n2093 0.152939
R14722 gnd.n2095 gnd.n2094 0.152939
R14723 gnd.n2096 gnd.n2095 0.152939
R14724 gnd.n2101 gnd.n2096 0.152939
R14725 gnd.n2102 gnd.n2101 0.152939
R14726 gnd.n2103 gnd.n2102 0.152939
R14727 gnd.n2104 gnd.n2103 0.152939
R14728 gnd.n2109 gnd.n2104 0.152939
R14729 gnd.n2110 gnd.n2109 0.152939
R14730 gnd.n2111 gnd.n2110 0.152939
R14731 gnd.n2112 gnd.n2111 0.152939
R14732 gnd.n2117 gnd.n2112 0.152939
R14733 gnd.n2118 gnd.n2117 0.152939
R14734 gnd.n2119 gnd.n2118 0.152939
R14735 gnd.n2120 gnd.n2119 0.152939
R14736 gnd.n2125 gnd.n2120 0.152939
R14737 gnd.n2126 gnd.n2125 0.152939
R14738 gnd.n2127 gnd.n2126 0.152939
R14739 gnd.n2128 gnd.n2127 0.152939
R14740 gnd.n2133 gnd.n2128 0.152939
R14741 gnd.n2134 gnd.n2133 0.152939
R14742 gnd.n2135 gnd.n2134 0.152939
R14743 gnd.n2136 gnd.n2135 0.152939
R14744 gnd.n2141 gnd.n2136 0.152939
R14745 gnd.n2142 gnd.n2141 0.152939
R14746 gnd.n2143 gnd.n2142 0.152939
R14747 gnd.n2144 gnd.n2143 0.152939
R14748 gnd.n2149 gnd.n2144 0.152939
R14749 gnd.n2150 gnd.n2149 0.152939
R14750 gnd.n2151 gnd.n2150 0.152939
R14751 gnd.n2152 gnd.n2151 0.152939
R14752 gnd.n2157 gnd.n2152 0.152939
R14753 gnd.n2158 gnd.n2157 0.152939
R14754 gnd.n2159 gnd.n2158 0.152939
R14755 gnd.n2160 gnd.n2159 0.152939
R14756 gnd.n2165 gnd.n2160 0.152939
R14757 gnd.n2166 gnd.n2165 0.152939
R14758 gnd.n2167 gnd.n2166 0.152939
R14759 gnd.n2168 gnd.n2167 0.152939
R14760 gnd.n2173 gnd.n2168 0.152939
R14761 gnd.n2174 gnd.n2173 0.152939
R14762 gnd.n2175 gnd.n2174 0.152939
R14763 gnd.n2176 gnd.n2175 0.152939
R14764 gnd.n2181 gnd.n2176 0.152939
R14765 gnd.n2182 gnd.n2181 0.152939
R14766 gnd.n2183 gnd.n2182 0.152939
R14767 gnd.n2184 gnd.n2183 0.152939
R14768 gnd.n2189 gnd.n2184 0.152939
R14769 gnd.n2190 gnd.n2189 0.152939
R14770 gnd.n2191 gnd.n2190 0.152939
R14771 gnd.n2192 gnd.n2191 0.152939
R14772 gnd.n2197 gnd.n2192 0.152939
R14773 gnd.n2198 gnd.n2197 0.152939
R14774 gnd.n2199 gnd.n2198 0.152939
R14775 gnd.n2200 gnd.n2199 0.152939
R14776 gnd.n2205 gnd.n2200 0.152939
R14777 gnd.n2206 gnd.n2205 0.152939
R14778 gnd.n2207 gnd.n2206 0.152939
R14779 gnd.n2208 gnd.n2207 0.152939
R14780 gnd.n2213 gnd.n2208 0.152939
R14781 gnd.n2214 gnd.n2213 0.152939
R14782 gnd.n2215 gnd.n2214 0.152939
R14783 gnd.n2216 gnd.n2215 0.152939
R14784 gnd.n2221 gnd.n2216 0.152939
R14785 gnd.n2222 gnd.n2221 0.152939
R14786 gnd.n2223 gnd.n2222 0.152939
R14787 gnd.n2224 gnd.n2223 0.152939
R14788 gnd.n2229 gnd.n2224 0.152939
R14789 gnd.n2230 gnd.n2229 0.152939
R14790 gnd.n2231 gnd.n2230 0.152939
R14791 gnd.n2232 gnd.n2231 0.152939
R14792 gnd.n2237 gnd.n2232 0.152939
R14793 gnd.n2238 gnd.n2237 0.152939
R14794 gnd.n2239 gnd.n2238 0.152939
R14795 gnd.n2240 gnd.n2239 0.152939
R14796 gnd.n2245 gnd.n2240 0.152939
R14797 gnd.n2246 gnd.n2245 0.152939
R14798 gnd.n2247 gnd.n2246 0.152939
R14799 gnd.n2248 gnd.n2247 0.152939
R14800 gnd.n2253 gnd.n2248 0.152939
R14801 gnd.n2254 gnd.n2253 0.152939
R14802 gnd.n2255 gnd.n2254 0.152939
R14803 gnd.n2256 gnd.n2255 0.152939
R14804 gnd.n2261 gnd.n2256 0.152939
R14805 gnd.n2262 gnd.n2261 0.152939
R14806 gnd.n2263 gnd.n2262 0.152939
R14807 gnd.n2264 gnd.n2263 0.152939
R14808 gnd.n2269 gnd.n2264 0.152939
R14809 gnd.n2606 gnd.n2269 0.152939
R14810 gnd.n2605 gnd.n2270 0.152939
R14811 gnd.n2272 gnd.n2270 0.152939
R14812 gnd.n2278 gnd.n2272 0.152939
R14813 gnd.n2279 gnd.n2278 0.152939
R14814 gnd.n2280 gnd.n2279 0.152939
R14815 gnd.n2281 gnd.n2280 0.152939
R14816 gnd.n2286 gnd.n2281 0.152939
R14817 gnd.n2287 gnd.n2286 0.152939
R14818 gnd.n2288 gnd.n2287 0.152939
R14819 gnd.n2289 gnd.n2288 0.152939
R14820 gnd.n2294 gnd.n2289 0.152939
R14821 gnd.n2295 gnd.n2294 0.152939
R14822 gnd.n2296 gnd.n2295 0.152939
R14823 gnd.n2297 gnd.n2296 0.152939
R14824 gnd.n2302 gnd.n2297 0.152939
R14825 gnd.n2303 gnd.n2302 0.152939
R14826 gnd.n2304 gnd.n2303 0.152939
R14827 gnd.n2305 gnd.n2304 0.152939
R14828 gnd.n2310 gnd.n2305 0.152939
R14829 gnd.n2311 gnd.n2310 0.152939
R14830 gnd.n2312 gnd.n2311 0.152939
R14831 gnd.n2313 gnd.n2312 0.152939
R14832 gnd.n2318 gnd.n2313 0.152939
R14833 gnd.n2319 gnd.n2318 0.152939
R14834 gnd.n2320 gnd.n2319 0.152939
R14835 gnd.n2321 gnd.n2320 0.152939
R14836 gnd.n2326 gnd.n2321 0.152939
R14837 gnd.n2327 gnd.n2326 0.152939
R14838 gnd.n2328 gnd.n2327 0.152939
R14839 gnd.n2329 gnd.n2328 0.152939
R14840 gnd.n2334 gnd.n2329 0.152939
R14841 gnd.n2335 gnd.n2334 0.152939
R14842 gnd.n2336 gnd.n2335 0.152939
R14843 gnd.n2337 gnd.n2336 0.152939
R14844 gnd.n2342 gnd.n2337 0.152939
R14845 gnd.n2343 gnd.n2342 0.152939
R14846 gnd.n2344 gnd.n2343 0.152939
R14847 gnd.n2345 gnd.n2344 0.152939
R14848 gnd.n2350 gnd.n2345 0.152939
R14849 gnd.n2351 gnd.n2350 0.152939
R14850 gnd.n2352 gnd.n2351 0.152939
R14851 gnd.n2353 gnd.n2352 0.152939
R14852 gnd.n2358 gnd.n2353 0.152939
R14853 gnd.n2359 gnd.n2358 0.152939
R14854 gnd.n2360 gnd.n2359 0.152939
R14855 gnd.n2361 gnd.n2360 0.152939
R14856 gnd.n2366 gnd.n2361 0.152939
R14857 gnd.n2367 gnd.n2366 0.152939
R14858 gnd.n2368 gnd.n2367 0.152939
R14859 gnd.n2369 gnd.n2368 0.152939
R14860 gnd.n2374 gnd.n2369 0.152939
R14861 gnd.n2375 gnd.n2374 0.152939
R14862 gnd.n2376 gnd.n2375 0.152939
R14863 gnd.n2377 gnd.n2376 0.152939
R14864 gnd.n2382 gnd.n2377 0.152939
R14865 gnd.n2383 gnd.n2382 0.152939
R14866 gnd.n2384 gnd.n2383 0.152939
R14867 gnd.n2385 gnd.n2384 0.152939
R14868 gnd.n2390 gnd.n2385 0.152939
R14869 gnd.n2391 gnd.n2390 0.152939
R14870 gnd.n2392 gnd.n2391 0.152939
R14871 gnd.n2393 gnd.n2392 0.152939
R14872 gnd.n2398 gnd.n2393 0.152939
R14873 gnd.n2399 gnd.n2398 0.152939
R14874 gnd.n2400 gnd.n2399 0.152939
R14875 gnd.n2401 gnd.n2400 0.152939
R14876 gnd.n2406 gnd.n2401 0.152939
R14877 gnd.n2407 gnd.n2406 0.152939
R14878 gnd.n2408 gnd.n2407 0.152939
R14879 gnd.n2409 gnd.n2408 0.152939
R14880 gnd.n2414 gnd.n2409 0.152939
R14881 gnd.n2415 gnd.n2414 0.152939
R14882 gnd.n2416 gnd.n2415 0.152939
R14883 gnd.n2417 gnd.n2416 0.152939
R14884 gnd.n2422 gnd.n2417 0.152939
R14885 gnd.n2423 gnd.n2422 0.152939
R14886 gnd.n2424 gnd.n2423 0.152939
R14887 gnd.n2425 gnd.n2424 0.152939
R14888 gnd.n2430 gnd.n2425 0.152939
R14889 gnd.n2431 gnd.n2430 0.152939
R14890 gnd.n2432 gnd.n2431 0.152939
R14891 gnd.n2433 gnd.n2432 0.152939
R14892 gnd.n2434 gnd.n2433 0.152939
R14893 gnd.n2435 gnd.n2434 0.152939
R14894 gnd.n7972 gnd.n112 0.152939
R14895 gnd.n137 gnd.n112 0.152939
R14896 gnd.n138 gnd.n137 0.152939
R14897 gnd.n139 gnd.n138 0.152939
R14898 gnd.n154 gnd.n139 0.152939
R14899 gnd.n155 gnd.n154 0.152939
R14900 gnd.n156 gnd.n155 0.152939
R14901 gnd.n157 gnd.n156 0.152939
R14902 gnd.n174 gnd.n157 0.152939
R14903 gnd.n175 gnd.n174 0.152939
R14904 gnd.n176 gnd.n175 0.152939
R14905 gnd.n177 gnd.n176 0.152939
R14906 gnd.n192 gnd.n177 0.152939
R14907 gnd.n193 gnd.n192 0.152939
R14908 gnd.n194 gnd.n193 0.152939
R14909 gnd.n195 gnd.n194 0.152939
R14910 gnd.n212 gnd.n195 0.152939
R14911 gnd.n213 gnd.n212 0.152939
R14912 gnd.n214 gnd.n213 0.152939
R14913 gnd.n215 gnd.n214 0.152939
R14914 gnd.n231 gnd.n215 0.152939
R14915 gnd.n232 gnd.n231 0.152939
R14916 gnd.n233 gnd.n232 0.152939
R14917 gnd.n234 gnd.n233 0.152939
R14918 gnd.n250 gnd.n234 0.152939
R14919 gnd.n251 gnd.n250 0.152939
R14920 gnd.n7887 gnd.n251 0.152939
R14921 gnd.n7981 gnd.n101 0.152939
R14922 gnd.n7619 gnd.n101 0.152939
R14923 gnd.n7622 gnd.n7619 0.152939
R14924 gnd.n7623 gnd.n7622 0.152939
R14925 gnd.n7624 gnd.n7623 0.152939
R14926 gnd.n7624 gnd.n7617 0.152939
R14927 gnd.n7630 gnd.n7617 0.152939
R14928 gnd.n7631 gnd.n7630 0.152939
R14929 gnd.n7632 gnd.n7631 0.152939
R14930 gnd.n7632 gnd.n7615 0.152939
R14931 gnd.n7638 gnd.n7615 0.152939
R14932 gnd.n7639 gnd.n7638 0.152939
R14933 gnd.n7640 gnd.n7639 0.152939
R14934 gnd.n7640 gnd.n7613 0.152939
R14935 gnd.n7646 gnd.n7613 0.152939
R14936 gnd.n7647 gnd.n7646 0.152939
R14937 gnd.n7648 gnd.n7647 0.152939
R14938 gnd.n7648 gnd.n7611 0.152939
R14939 gnd.n7654 gnd.n7611 0.152939
R14940 gnd.n7655 gnd.n7654 0.152939
R14941 gnd.n7656 gnd.n7655 0.152939
R14942 gnd.n7657 gnd.n7656 0.152939
R14943 gnd.n7658 gnd.n7657 0.152939
R14944 gnd.n7659 gnd.n7658 0.152939
R14945 gnd.n7660 gnd.n7659 0.152939
R14946 gnd.n7661 gnd.n7660 0.152939
R14947 gnd.n7662 gnd.n7661 0.152939
R14948 gnd.n7663 gnd.n7662 0.152939
R14949 gnd.n7664 gnd.n7663 0.152939
R14950 gnd.n7665 gnd.n7664 0.152939
R14951 gnd.n7666 gnd.n7665 0.152939
R14952 gnd.n7680 gnd.n352 0.152939
R14953 gnd.n7681 gnd.n7680 0.152939
R14954 gnd.n7681 gnd.n7676 0.152939
R14955 gnd.n7689 gnd.n7676 0.152939
R14956 gnd.n7690 gnd.n7689 0.152939
R14957 gnd.n7691 gnd.n7690 0.152939
R14958 gnd.n7691 gnd.n7674 0.152939
R14959 gnd.n7699 gnd.n7674 0.152939
R14960 gnd.n7700 gnd.n7699 0.152939
R14961 gnd.n7701 gnd.n7700 0.152939
R14962 gnd.n7701 gnd.n7672 0.152939
R14963 gnd.n7709 gnd.n7672 0.152939
R14964 gnd.n7710 gnd.n7709 0.152939
R14965 gnd.n7711 gnd.n7710 0.152939
R14966 gnd.n7711 gnd.n7670 0.152939
R14967 gnd.n7719 gnd.n7670 0.152939
R14968 gnd.n7720 gnd.n7719 0.152939
R14969 gnd.n7721 gnd.n7720 0.152939
R14970 gnd.n7886 gnd.n252 0.152939
R14971 gnd.n294 gnd.n252 0.152939
R14972 gnd.n295 gnd.n294 0.152939
R14973 gnd.n296 gnd.n295 0.152939
R14974 gnd.n297 gnd.n296 0.152939
R14975 gnd.n298 gnd.n297 0.152939
R14976 gnd.n299 gnd.n298 0.152939
R14977 gnd.n300 gnd.n299 0.152939
R14978 gnd.n301 gnd.n300 0.152939
R14979 gnd.n302 gnd.n301 0.152939
R14980 gnd.n303 gnd.n302 0.152939
R14981 gnd.n304 gnd.n303 0.152939
R14982 gnd.n305 gnd.n304 0.152939
R14983 gnd.n306 gnd.n305 0.152939
R14984 gnd.n307 gnd.n306 0.152939
R14985 gnd.n308 gnd.n307 0.152939
R14986 gnd.n309 gnd.n308 0.152939
R14987 gnd.n310 gnd.n309 0.152939
R14988 gnd.n311 gnd.n310 0.152939
R14989 gnd.n312 gnd.n311 0.152939
R14990 gnd.n313 gnd.n312 0.152939
R14991 gnd.n314 gnd.n313 0.152939
R14992 gnd.n315 gnd.n314 0.152939
R14993 gnd.n316 gnd.n315 0.152939
R14994 gnd.n317 gnd.n316 0.152939
R14995 gnd.n318 gnd.n317 0.152939
R14996 gnd.n319 gnd.n318 0.152939
R14997 gnd.n320 gnd.n319 0.152939
R14998 gnd.n321 gnd.n320 0.152939
R14999 gnd.n322 gnd.n321 0.152939
R15000 gnd.n323 gnd.n322 0.152939
R15001 gnd.n324 gnd.n323 0.152939
R15002 gnd.n325 gnd.n324 0.152939
R15003 gnd.n326 gnd.n325 0.152939
R15004 gnd.n327 gnd.n326 0.152939
R15005 gnd.n328 gnd.n327 0.152939
R15006 gnd.n7807 gnd.n328 0.152939
R15007 gnd.n7807 gnd.n7806 0.152939
R15008 gnd.n7806 gnd.n7805 0.152939
R15009 gnd.n7805 gnd.n332 0.152939
R15010 gnd.n333 gnd.n332 0.152939
R15011 gnd.n334 gnd.n333 0.152939
R15012 gnd.n335 gnd.n334 0.152939
R15013 gnd.n336 gnd.n335 0.152939
R15014 gnd.n337 gnd.n336 0.152939
R15015 gnd.n338 gnd.n337 0.152939
R15016 gnd.n339 gnd.n338 0.152939
R15017 gnd.n340 gnd.n339 0.152939
R15018 gnd.n341 gnd.n340 0.152939
R15019 gnd.n342 gnd.n341 0.152939
R15020 gnd.n343 gnd.n342 0.152939
R15021 gnd.n344 gnd.n343 0.152939
R15022 gnd.n345 gnd.n344 0.152939
R15023 gnd.n346 gnd.n345 0.152939
R15024 gnd.n347 gnd.n346 0.152939
R15025 gnd.n348 gnd.n347 0.152939
R15026 gnd.n7765 gnd.n348 0.152939
R15027 gnd.n7765 gnd.n7764 0.152939
R15028 gnd.n612 gnd.n549 0.152939
R15029 gnd.n613 gnd.n612 0.152939
R15030 gnd.n614 gnd.n613 0.152939
R15031 gnd.n615 gnd.n614 0.152939
R15032 gnd.n616 gnd.n615 0.152939
R15033 gnd.n617 gnd.n616 0.152939
R15034 gnd.n618 gnd.n617 0.152939
R15035 gnd.n619 gnd.n618 0.152939
R15036 gnd.n620 gnd.n619 0.152939
R15037 gnd.n621 gnd.n620 0.152939
R15038 gnd.n622 gnd.n621 0.152939
R15039 gnd.n623 gnd.n622 0.152939
R15040 gnd.n624 gnd.n623 0.152939
R15041 gnd.n625 gnd.n624 0.152939
R15042 gnd.n626 gnd.n625 0.152939
R15043 gnd.n627 gnd.n626 0.152939
R15044 gnd.n628 gnd.n627 0.152939
R15045 gnd.n631 gnd.n628 0.152939
R15046 gnd.n632 gnd.n631 0.152939
R15047 gnd.n633 gnd.n632 0.152939
R15048 gnd.n634 gnd.n633 0.152939
R15049 gnd.n635 gnd.n634 0.152939
R15050 gnd.n636 gnd.n635 0.152939
R15051 gnd.n637 gnd.n636 0.152939
R15052 gnd.n638 gnd.n637 0.152939
R15053 gnd.n643 gnd.n642 0.152939
R15054 gnd.n644 gnd.n643 0.152939
R15055 gnd.n645 gnd.n644 0.152939
R15056 gnd.n646 gnd.n645 0.152939
R15057 gnd.n647 gnd.n646 0.152939
R15058 gnd.n648 gnd.n647 0.152939
R15059 gnd.n649 gnd.n648 0.152939
R15060 gnd.n650 gnd.n649 0.152939
R15061 gnd.n651 gnd.n650 0.152939
R15062 gnd.n654 gnd.n651 0.152939
R15063 gnd.n655 gnd.n654 0.152939
R15064 gnd.n656 gnd.n655 0.152939
R15065 gnd.n657 gnd.n656 0.152939
R15066 gnd.n658 gnd.n657 0.152939
R15067 gnd.n659 gnd.n658 0.152939
R15068 gnd.n660 gnd.n659 0.152939
R15069 gnd.n661 gnd.n660 0.152939
R15070 gnd.n662 gnd.n661 0.152939
R15071 gnd.n663 gnd.n662 0.152939
R15072 gnd.n664 gnd.n663 0.152939
R15073 gnd.n665 gnd.n664 0.152939
R15074 gnd.n666 gnd.n665 0.152939
R15075 gnd.n667 gnd.n666 0.152939
R15076 gnd.n668 gnd.n667 0.152939
R15077 gnd.n669 gnd.n668 0.152939
R15078 gnd.n670 gnd.n669 0.152939
R15079 gnd.n671 gnd.n670 0.152939
R15080 gnd.n672 gnd.n671 0.152939
R15081 gnd.n7161 gnd.n672 0.152939
R15082 gnd.n7161 gnd.n7160 0.152939
R15083 gnd.n7314 gnd.n7313 0.152939
R15084 gnd.n7315 gnd.n7314 0.152939
R15085 gnd.n7316 gnd.n7315 0.152939
R15086 gnd.n7316 gnd.n519 0.152939
R15087 gnd.n7355 gnd.n519 0.152939
R15088 gnd.n7356 gnd.n7355 0.152939
R15089 gnd.n7357 gnd.n7356 0.152939
R15090 gnd.n7358 gnd.n7357 0.152939
R15091 gnd.n7358 gnd.n483 0.152939
R15092 gnd.n7404 gnd.n483 0.152939
R15093 gnd.n7405 gnd.n7404 0.152939
R15094 gnd.n7406 gnd.n7405 0.152939
R15095 gnd.n7407 gnd.n7406 0.152939
R15096 gnd.n7407 gnd.n453 0.152939
R15097 gnd.n7441 gnd.n453 0.152939
R15098 gnd.n7442 gnd.n7441 0.152939
R15099 gnd.n7443 gnd.n7442 0.152939
R15100 gnd.n7444 gnd.n7443 0.152939
R15101 gnd.n7444 gnd.n418 0.152939
R15102 gnd.n7489 gnd.n418 0.152939
R15103 gnd.n7490 gnd.n7489 0.152939
R15104 gnd.n7491 gnd.n7490 0.152939
R15105 gnd.n7493 gnd.n7491 0.152939
R15106 gnd.n7493 gnd.n7492 0.152939
R15107 gnd.n7492 gnd.n381 0.152939
R15108 gnd.n381 gnd.n113 0.152939
R15109 gnd.n7972 gnd.n113 0.152939
R15110 gnd.n3601 gnd.n3599 0.152939
R15111 gnd.n3601 gnd.n3600 0.152939
R15112 gnd.n3600 gnd.n1754 0.152939
R15113 gnd.n5377 gnd.n1754 0.152939
R15114 gnd.n5378 gnd.n5377 0.152939
R15115 gnd.n5379 gnd.n5378 0.152939
R15116 gnd.n5380 gnd.n5379 0.152939
R15117 gnd.n5380 gnd.n1719 0.152939
R15118 gnd.n5427 gnd.n1719 0.152939
R15119 gnd.n5428 gnd.n5427 0.152939
R15120 gnd.n5429 gnd.n5428 0.152939
R15121 gnd.n5430 gnd.n5429 0.152939
R15122 gnd.n5430 gnd.n1655 0.152939
R15123 gnd.n5489 gnd.n1655 0.152939
R15124 gnd.n5490 gnd.n5489 0.152939
R15125 gnd.n5491 gnd.n5490 0.152939
R15126 gnd.n5491 gnd.n1651 0.152939
R15127 gnd.n5497 gnd.n1651 0.152939
R15128 gnd.n5498 gnd.n5497 0.152939
R15129 gnd.n5499 gnd.n5498 0.152939
R15130 gnd.n5500 gnd.n5499 0.152939
R15131 gnd.n5501 gnd.n5500 0.152939
R15132 gnd.n5504 gnd.n5501 0.152939
R15133 gnd.n5505 gnd.n5504 0.152939
R15134 gnd.n5506 gnd.n5505 0.152939
R15135 gnd.n5507 gnd.n5506 0.152939
R15136 gnd.n5510 gnd.n5507 0.152939
R15137 gnd.n5511 gnd.n5510 0.152939
R15138 gnd.n5512 gnd.n5511 0.152939
R15139 gnd.n5513 gnd.n5512 0.152939
R15140 gnd.n5514 gnd.n5513 0.152939
R15141 gnd.n5514 gnd.n1226 0.152939
R15142 gnd.n6167 gnd.n1226 0.152939
R15143 gnd.n6168 gnd.n6167 0.152939
R15144 gnd.n6169 gnd.n6168 0.152939
R15145 gnd.n6169 gnd.n1213 0.152939
R15146 gnd.n6183 gnd.n1213 0.152939
R15147 gnd.n6184 gnd.n6183 0.152939
R15148 gnd.n6185 gnd.n6184 0.152939
R15149 gnd.n6185 gnd.n1199 0.152939
R15150 gnd.n6199 gnd.n1199 0.152939
R15151 gnd.n6200 gnd.n6199 0.152939
R15152 gnd.n6201 gnd.n6200 0.152939
R15153 gnd.n6201 gnd.n1185 0.152939
R15154 gnd.n6215 gnd.n1185 0.152939
R15155 gnd.n6216 gnd.n6215 0.152939
R15156 gnd.n6217 gnd.n6216 0.152939
R15157 gnd.n6217 gnd.n1170 0.152939
R15158 gnd.n6231 gnd.n1170 0.152939
R15159 gnd.n6232 gnd.n6231 0.152939
R15160 gnd.n6233 gnd.n6232 0.152939
R15161 gnd.n6233 gnd.n1156 0.152939
R15162 gnd.n6247 gnd.n1156 0.152939
R15163 gnd.n6248 gnd.n6247 0.152939
R15164 gnd.n6249 gnd.n6248 0.152939
R15165 gnd.n6249 gnd.n1140 0.152939
R15166 gnd.n6263 gnd.n1140 0.152939
R15167 gnd.n6264 gnd.n6263 0.152939
R15168 gnd.n6265 gnd.n6264 0.152939
R15169 gnd.n6265 gnd.n1126 0.152939
R15170 gnd.n6279 gnd.n1126 0.152939
R15171 gnd.n6280 gnd.n6279 0.152939
R15172 gnd.n6281 gnd.n6280 0.152939
R15173 gnd.n6281 gnd.n1112 0.152939
R15174 gnd.n6295 gnd.n1112 0.152939
R15175 gnd.n6296 gnd.n6295 0.152939
R15176 gnd.n6297 gnd.n6296 0.152939
R15177 gnd.n6297 gnd.n1099 0.152939
R15178 gnd.n6311 gnd.n1099 0.152939
R15179 gnd.n6312 gnd.n6311 0.152939
R15180 gnd.n6313 gnd.n6312 0.152939
R15181 gnd.n6313 gnd.n1085 0.152939
R15182 gnd.n6327 gnd.n1085 0.152939
R15183 gnd.n6328 gnd.n6327 0.152939
R15184 gnd.n6329 gnd.n6328 0.152939
R15185 gnd.n6329 gnd.n1067 0.152939
R15186 gnd.n6349 gnd.n1067 0.152939
R15187 gnd.n6350 gnd.n6349 0.152939
R15188 gnd.n6351 gnd.n6350 0.152939
R15189 gnd.n6352 gnd.n6351 0.152939
R15190 gnd.n6352 gnd.n1029 0.152939
R15191 gnd.n6407 gnd.n1029 0.152939
R15192 gnd.n6408 gnd.n6407 0.152939
R15193 gnd.n6409 gnd.n6408 0.152939
R15194 gnd.n6410 gnd.n6409 0.152939
R15195 gnd.n6410 gnd.n990 0.152939
R15196 gnd.n6465 gnd.n990 0.152939
R15197 gnd.n6466 gnd.n6465 0.152939
R15198 gnd.n6467 gnd.n6466 0.152939
R15199 gnd.n6468 gnd.n6467 0.152939
R15200 gnd.n6468 gnd.n922 0.152939
R15201 gnd.n6903 gnd.n922 0.152939
R15202 gnd.n6904 gnd.n6903 0.152939
R15203 gnd.n6905 gnd.n6904 0.152939
R15204 gnd.n6905 gnd.n908 0.152939
R15205 gnd.n6919 gnd.n908 0.152939
R15206 gnd.n6920 gnd.n6919 0.152939
R15207 gnd.n6921 gnd.n6920 0.152939
R15208 gnd.n6921 gnd.n895 0.152939
R15209 gnd.n6935 gnd.n895 0.152939
R15210 gnd.n6936 gnd.n6935 0.152939
R15211 gnd.n6937 gnd.n6936 0.152939
R15212 gnd.n6937 gnd.n881 0.152939
R15213 gnd.n6951 gnd.n881 0.152939
R15214 gnd.n6952 gnd.n6951 0.152939
R15215 gnd.n6953 gnd.n6952 0.152939
R15216 gnd.n6953 gnd.n867 0.152939
R15217 gnd.n6967 gnd.n867 0.152939
R15218 gnd.n6968 gnd.n6967 0.152939
R15219 gnd.n6969 gnd.n6968 0.152939
R15220 gnd.n6969 gnd.n852 0.152939
R15221 gnd.n6983 gnd.n852 0.152939
R15222 gnd.n6984 gnd.n6983 0.152939
R15223 gnd.n6985 gnd.n6984 0.152939
R15224 gnd.n6985 gnd.n837 0.152939
R15225 gnd.n6999 gnd.n837 0.152939
R15226 gnd.n7000 gnd.n6999 0.152939
R15227 gnd.n7001 gnd.n7000 0.152939
R15228 gnd.n7001 gnd.n824 0.152939
R15229 gnd.n7015 gnd.n824 0.152939
R15230 gnd.n7016 gnd.n7015 0.152939
R15231 gnd.n7017 gnd.n7016 0.152939
R15232 gnd.n7017 gnd.n810 0.152939
R15233 gnd.n7031 gnd.n810 0.152939
R15234 gnd.n7032 gnd.n7031 0.152939
R15235 gnd.n7033 gnd.n7032 0.152939
R15236 gnd.n7033 gnd.n796 0.152939
R15237 gnd.n7047 gnd.n796 0.152939
R15238 gnd.n7048 gnd.n7047 0.152939
R15239 gnd.n7049 gnd.n7048 0.152939
R15240 gnd.n7051 gnd.n7049 0.152939
R15241 gnd.n7051 gnd.n7050 0.152939
R15242 gnd.n7050 gnd.n782 0.152939
R15243 gnd.n7068 gnd.n782 0.152939
R15244 gnd.n7069 gnd.n7068 0.152939
R15245 gnd.n7070 gnd.n7069 0.152939
R15246 gnd.n7071 gnd.n7070 0.152939
R15247 gnd.n7072 gnd.n7071 0.152939
R15248 gnd.n7072 gnd.n568 0.152939
R15249 gnd.n7279 gnd.n568 0.152939
R15250 gnd.n7280 gnd.n7279 0.152939
R15251 gnd.n7281 gnd.n7280 0.152939
R15252 gnd.n7282 gnd.n7281 0.152939
R15253 gnd.n7283 gnd.n7282 0.152939
R15254 gnd.n7286 gnd.n7283 0.152939
R15255 gnd.n7287 gnd.n7286 0.152939
R15256 gnd.n7288 gnd.n7287 0.152939
R15257 gnd.n7290 gnd.n7288 0.152939
R15258 gnd.n7290 gnd.n7289 0.152939
R15259 gnd.n7289 gnd.n500 0.152939
R15260 gnd.n7377 gnd.n500 0.152939
R15261 gnd.n7378 gnd.n7377 0.152939
R15262 gnd.n7379 gnd.n7378 0.152939
R15263 gnd.n7380 gnd.n7379 0.152939
R15264 gnd.n7381 gnd.n7380 0.152939
R15265 gnd.n7383 gnd.n7381 0.152939
R15266 gnd.n7384 gnd.n7383 0.152939
R15267 gnd.n7384 gnd.n435 0.152939
R15268 gnd.n7461 gnd.n435 0.152939
R15269 gnd.n7462 gnd.n7461 0.152939
R15270 gnd.n7463 gnd.n7462 0.152939
R15271 gnd.n7464 gnd.n7463 0.152939
R15272 gnd.n7465 gnd.n7464 0.152939
R15273 gnd.n7465 gnd.n400 0.152939
R15274 gnd.n7513 gnd.n400 0.152939
R15275 gnd.n7514 gnd.n7513 0.152939
R15276 gnd.n7515 gnd.n7514 0.152939
R15277 gnd.n3473 gnd.n3414 0.152939
R15278 gnd.n3479 gnd.n3414 0.152939
R15279 gnd.n3480 gnd.n3479 0.152939
R15280 gnd.n3481 gnd.n3480 0.152939
R15281 gnd.n3481 gnd.n3412 0.152939
R15282 gnd.n3487 gnd.n3412 0.152939
R15283 gnd.n3488 gnd.n3487 0.152939
R15284 gnd.n3489 gnd.n3488 0.152939
R15285 gnd.n3489 gnd.n3410 0.152939
R15286 gnd.n3495 gnd.n3410 0.152939
R15287 gnd.n3496 gnd.n3495 0.152939
R15288 gnd.n3497 gnd.n3496 0.152939
R15289 gnd.n3497 gnd.n3408 0.152939
R15290 gnd.n3503 gnd.n3408 0.152939
R15291 gnd.n3504 gnd.n3503 0.152939
R15292 gnd.n3505 gnd.n3504 0.152939
R15293 gnd.n3505 gnd.n3406 0.152939
R15294 gnd.n3511 gnd.n3406 0.152939
R15295 gnd.n3512 gnd.n3511 0.152939
R15296 gnd.n3513 gnd.n3512 0.152939
R15297 gnd.n3513 gnd.n3404 0.152939
R15298 gnd.n3519 gnd.n3404 0.152939
R15299 gnd.n3520 gnd.n3519 0.152939
R15300 gnd.n3521 gnd.n3520 0.152939
R15301 gnd.n3521 gnd.n3402 0.152939
R15302 gnd.n3526 gnd.n3402 0.152939
R15303 gnd.n3527 gnd.n3526 0.152939
R15304 gnd.n3528 gnd.n3527 0.152939
R15305 gnd.n3529 gnd.n3528 0.152939
R15306 gnd.n3530 gnd.n3529 0.152939
R15307 gnd.n3531 gnd.n3530 0.152939
R15308 gnd.n3428 gnd.n3270 0.152939
R15309 gnd.n3436 gnd.n3428 0.152939
R15310 gnd.n3437 gnd.n3436 0.152939
R15311 gnd.n3438 gnd.n3437 0.152939
R15312 gnd.n3438 gnd.n3426 0.152939
R15313 gnd.n3446 gnd.n3426 0.152939
R15314 gnd.n3447 gnd.n3446 0.152939
R15315 gnd.n3448 gnd.n3447 0.152939
R15316 gnd.n3448 gnd.n3424 0.152939
R15317 gnd.n3456 gnd.n3424 0.152939
R15318 gnd.n3457 gnd.n3456 0.152939
R15319 gnd.n3458 gnd.n3457 0.152939
R15320 gnd.n3458 gnd.n3422 0.152939
R15321 gnd.n3466 gnd.n3422 0.152939
R15322 gnd.n3467 gnd.n3466 0.152939
R15323 gnd.n3468 gnd.n3467 0.152939
R15324 gnd.n3468 gnd.n3415 0.152939
R15325 gnd.n3472 gnd.n3415 0.152939
R15326 gnd.n5353 gnd.n5352 0.152939
R15327 gnd.n5353 gnd.n1737 0.152939
R15328 gnd.n5395 gnd.n1737 0.152939
R15329 gnd.n5396 gnd.n5395 0.152939
R15330 gnd.n5397 gnd.n5396 0.152939
R15331 gnd.n5398 gnd.n5397 0.152939
R15332 gnd.n5398 gnd.n1699 0.152939
R15333 gnd.n5445 gnd.n1699 0.152939
R15334 gnd.n5446 gnd.n5445 0.152939
R15335 gnd.n5447 gnd.n5446 0.152939
R15336 gnd.n5448 gnd.n5447 0.152939
R15337 gnd.n5448 gnd.n1665 0.152939
R15338 gnd.n5480 gnd.n1665 0.152939
R15339 gnd.n5481 gnd.n5480 0.152939
R15340 gnd.n5482 gnd.n5481 0.152939
R15341 gnd.n5482 gnd.n1634 0.152939
R15342 gnd.n5548 gnd.n1634 0.152939
R15343 gnd.n5549 gnd.n5548 0.152939
R15344 gnd.n5550 gnd.n5549 0.152939
R15345 gnd.n5551 gnd.n5550 0.152939
R15346 gnd.n5551 gnd.n1608 0.152939
R15347 gnd.n5588 gnd.n1608 0.152939
R15348 gnd.n5589 gnd.n5588 0.152939
R15349 gnd.n5590 gnd.n5589 0.152939
R15350 gnd.n5591 gnd.n5590 0.152939
R15351 gnd.n5591 gnd.n1250 0.152939
R15352 gnd.n6149 gnd.n1250 0.152939
R15353 gnd.n6148 gnd.n1251 0.152939
R15354 gnd.n1256 gnd.n1251 0.152939
R15355 gnd.n1257 gnd.n1256 0.152939
R15356 gnd.n1258 gnd.n1257 0.152939
R15357 gnd.n1259 gnd.n1258 0.152939
R15358 gnd.n1260 gnd.n1259 0.152939
R15359 gnd.n1264 gnd.n1260 0.152939
R15360 gnd.n1265 gnd.n1264 0.152939
R15361 gnd.n1266 gnd.n1265 0.152939
R15362 gnd.n1267 gnd.n1266 0.152939
R15363 gnd.n1271 gnd.n1267 0.152939
R15364 gnd.n1272 gnd.n1271 0.152939
R15365 gnd.n1273 gnd.n1272 0.152939
R15366 gnd.n1274 gnd.n1273 0.152939
R15367 gnd.n1278 gnd.n1274 0.152939
R15368 gnd.n1279 gnd.n1278 0.152939
R15369 gnd.n1280 gnd.n1279 0.152939
R15370 gnd.n1283 gnd.n1280 0.152939
R15371 gnd.n1287 gnd.n1283 0.152939
R15372 gnd.n1288 gnd.n1287 0.152939
R15373 gnd.n1289 gnd.n1288 0.152939
R15374 gnd.n1290 gnd.n1289 0.152939
R15375 gnd.n1294 gnd.n1290 0.152939
R15376 gnd.n1295 gnd.n1294 0.152939
R15377 gnd.n1296 gnd.n1295 0.152939
R15378 gnd.n1512 gnd.n1511 0.152939
R15379 gnd.n1521 gnd.n1512 0.152939
R15380 gnd.n1522 gnd.n1521 0.152939
R15381 gnd.n1523 gnd.n1522 0.152939
R15382 gnd.n1523 gnd.n1507 0.152939
R15383 gnd.n1531 gnd.n1507 0.152939
R15384 gnd.n1532 gnd.n1531 0.152939
R15385 gnd.n1533 gnd.n1532 0.152939
R15386 gnd.n1533 gnd.n1501 0.152939
R15387 gnd.n1541 gnd.n1501 0.152939
R15388 gnd.n1542 gnd.n1541 0.152939
R15389 gnd.n1543 gnd.n1542 0.152939
R15390 gnd.n1543 gnd.n1497 0.152939
R15391 gnd.n1551 gnd.n1497 0.152939
R15392 gnd.n1552 gnd.n1551 0.152939
R15393 gnd.n1553 gnd.n1552 0.152939
R15394 gnd.n1553 gnd.n1493 0.152939
R15395 gnd.n1561 gnd.n1493 0.152939
R15396 gnd.n1562 gnd.n1561 0.152939
R15397 gnd.n1563 gnd.n1562 0.152939
R15398 gnd.n1563 gnd.n1489 0.152939
R15399 gnd.n1571 gnd.n1489 0.152939
R15400 gnd.n1572 gnd.n1571 0.152939
R15401 gnd.n1573 gnd.n1572 0.152939
R15402 gnd.n1573 gnd.n1485 0.152939
R15403 gnd.n1581 gnd.n1485 0.152939
R15404 gnd.n1582 gnd.n1581 0.152939
R15405 gnd.n1583 gnd.n1582 0.152939
R15406 gnd.n1583 gnd.n1479 0.152939
R15407 gnd.n1590 gnd.n1479 0.152939
R15408 gnd.n3207 gnd.n3206 0.152939
R15409 gnd.n3208 gnd.n3207 0.152939
R15410 gnd.n3209 gnd.n3208 0.152939
R15411 gnd.n3210 gnd.n3209 0.152939
R15412 gnd.n3211 gnd.n3210 0.152939
R15413 gnd.n3212 gnd.n3211 0.152939
R15414 gnd.n3213 gnd.n3212 0.152939
R15415 gnd.n3214 gnd.n3213 0.152939
R15416 gnd.n3215 gnd.n3214 0.152939
R15417 gnd.n3216 gnd.n3215 0.152939
R15418 gnd.n3217 gnd.n3216 0.152939
R15419 gnd.n3218 gnd.n3217 0.152939
R15420 gnd.n3219 gnd.n3218 0.152939
R15421 gnd.n3220 gnd.n3219 0.152939
R15422 gnd.n3221 gnd.n3220 0.152939
R15423 gnd.n3222 gnd.n3221 0.152939
R15424 gnd.n3223 gnd.n3222 0.152939
R15425 gnd.n3226 gnd.n3223 0.152939
R15426 gnd.n3227 gnd.n3226 0.152939
R15427 gnd.n3228 gnd.n3227 0.152939
R15428 gnd.n3229 gnd.n3228 0.152939
R15429 gnd.n3230 gnd.n3229 0.152939
R15430 gnd.n3231 gnd.n3230 0.152939
R15431 gnd.n3232 gnd.n3231 0.152939
R15432 gnd.n3233 gnd.n3232 0.152939
R15433 gnd.n3234 gnd.n3233 0.152939
R15434 gnd.n3235 gnd.n3234 0.152939
R15435 gnd.n3236 gnd.n3235 0.152939
R15436 gnd.n3237 gnd.n3236 0.152939
R15437 gnd.n3238 gnd.n3237 0.152939
R15438 gnd.n3239 gnd.n3238 0.152939
R15439 gnd.n3240 gnd.n3239 0.152939
R15440 gnd.n3241 gnd.n3240 0.152939
R15441 gnd.n3242 gnd.n3241 0.152939
R15442 gnd.n3243 gnd.n3242 0.152939
R15443 gnd.n3244 gnd.n3243 0.152939
R15444 gnd.n3245 gnd.n3244 0.152939
R15445 gnd.n3248 gnd.n3245 0.152939
R15446 gnd.n3249 gnd.n3248 0.152939
R15447 gnd.n3250 gnd.n3249 0.152939
R15448 gnd.n3251 gnd.n3250 0.152939
R15449 gnd.n3252 gnd.n3251 0.152939
R15450 gnd.n3253 gnd.n3252 0.152939
R15451 gnd.n3254 gnd.n3253 0.152939
R15452 gnd.n3255 gnd.n3254 0.152939
R15453 gnd.n3256 gnd.n3255 0.152939
R15454 gnd.n3257 gnd.n3256 0.152939
R15455 gnd.n3258 gnd.n3257 0.152939
R15456 gnd.n3259 gnd.n3258 0.152939
R15457 gnd.n3260 gnd.n3259 0.152939
R15458 gnd.n3261 gnd.n3260 0.152939
R15459 gnd.n3262 gnd.n3261 0.152939
R15460 gnd.n3263 gnd.n3262 0.152939
R15461 gnd.n3264 gnd.n3263 0.152939
R15462 gnd.n3265 gnd.n3264 0.152939
R15463 gnd.n3266 gnd.n3265 0.152939
R15464 gnd.n3716 gnd.n3266 0.152939
R15465 gnd.n3716 gnd.n3715 0.152939
R15466 gnd.n3281 gnd.n3280 0.152939
R15467 gnd.n3282 gnd.n3281 0.152939
R15468 gnd.n3283 gnd.n3282 0.152939
R15469 gnd.n3303 gnd.n3283 0.152939
R15470 gnd.n3304 gnd.n3303 0.152939
R15471 gnd.n3305 gnd.n3304 0.152939
R15472 gnd.n3306 gnd.n3305 0.152939
R15473 gnd.n3321 gnd.n3306 0.152939
R15474 gnd.n3322 gnd.n3321 0.152939
R15475 gnd.n3323 gnd.n3322 0.152939
R15476 gnd.n3324 gnd.n3323 0.152939
R15477 gnd.n3341 gnd.n3324 0.152939
R15478 gnd.n3342 gnd.n3341 0.152939
R15479 gnd.n3343 gnd.n3342 0.152939
R15480 gnd.n3344 gnd.n3343 0.152939
R15481 gnd.n3359 gnd.n3344 0.152939
R15482 gnd.n3360 gnd.n3359 0.152939
R15483 gnd.n3361 gnd.n3360 0.152939
R15484 gnd.n3362 gnd.n3361 0.152939
R15485 gnd.n3379 gnd.n3362 0.152939
R15486 gnd.n3380 gnd.n3379 0.152939
R15487 gnd.n3381 gnd.n3380 0.152939
R15488 gnd.n3382 gnd.n3381 0.152939
R15489 gnd.n3632 gnd.n3382 0.152939
R15490 gnd.n3633 gnd.n3632 0.152939
R15491 gnd.n3633 gnd.n1773 0.152939
R15492 gnd.n5352 gnd.n1773 0.152939
R15493 gnd.n2944 gnd.n1931 0.152939
R15494 gnd.n2952 gnd.n1931 0.152939
R15495 gnd.n2953 gnd.n2952 0.152939
R15496 gnd.n2954 gnd.n2953 0.152939
R15497 gnd.n2954 gnd.n1925 0.152939
R15498 gnd.n2962 gnd.n1925 0.152939
R15499 gnd.n2963 gnd.n2962 0.152939
R15500 gnd.n2964 gnd.n2963 0.152939
R15501 gnd.n2964 gnd.n1919 0.152939
R15502 gnd.n2972 gnd.n1919 0.152939
R15503 gnd.n2973 gnd.n2972 0.152939
R15504 gnd.n2974 gnd.n2973 0.152939
R15505 gnd.n2974 gnd.n1913 0.152939
R15506 gnd.n2982 gnd.n1913 0.152939
R15507 gnd.n2983 gnd.n2982 0.152939
R15508 gnd.n2984 gnd.n2983 0.152939
R15509 gnd.n2984 gnd.n1907 0.152939
R15510 gnd.n2992 gnd.n1907 0.152939
R15511 gnd.n2993 gnd.n2992 0.152939
R15512 gnd.n2994 gnd.n2993 0.152939
R15513 gnd.n2994 gnd.n1901 0.152939
R15514 gnd.n3002 gnd.n1901 0.152939
R15515 gnd.n3003 gnd.n3002 0.152939
R15516 gnd.n3004 gnd.n3003 0.152939
R15517 gnd.n3004 gnd.n1895 0.152939
R15518 gnd.n3012 gnd.n1895 0.152939
R15519 gnd.n3013 gnd.n3012 0.152939
R15520 gnd.n3014 gnd.n3013 0.152939
R15521 gnd.n3014 gnd.n1889 0.152939
R15522 gnd.n3022 gnd.n1889 0.152939
R15523 gnd.n3023 gnd.n3022 0.152939
R15524 gnd.n3024 gnd.n3023 0.152939
R15525 gnd.n3024 gnd.n1883 0.152939
R15526 gnd.n3032 gnd.n1883 0.152939
R15527 gnd.n3033 gnd.n3032 0.152939
R15528 gnd.n3034 gnd.n3033 0.152939
R15529 gnd.n3034 gnd.n1877 0.152939
R15530 gnd.n3042 gnd.n1877 0.152939
R15531 gnd.n3043 gnd.n3042 0.152939
R15532 gnd.n3044 gnd.n3043 0.152939
R15533 gnd.n3044 gnd.n1871 0.152939
R15534 gnd.n3052 gnd.n1871 0.152939
R15535 gnd.n3053 gnd.n3052 0.152939
R15536 gnd.n3054 gnd.n3053 0.152939
R15537 gnd.n3054 gnd.n1865 0.152939
R15538 gnd.n3062 gnd.n1865 0.152939
R15539 gnd.n3063 gnd.n3062 0.152939
R15540 gnd.n3064 gnd.n3063 0.152939
R15541 gnd.n3064 gnd.n1859 0.152939
R15542 gnd.n3072 gnd.n1859 0.152939
R15543 gnd.n3073 gnd.n3072 0.152939
R15544 gnd.n3074 gnd.n3073 0.152939
R15545 gnd.n3074 gnd.n1853 0.152939
R15546 gnd.n3082 gnd.n1853 0.152939
R15547 gnd.n3083 gnd.n3082 0.152939
R15548 gnd.n3084 gnd.n3083 0.152939
R15549 gnd.n3084 gnd.n1847 0.152939
R15550 gnd.n3092 gnd.n1847 0.152939
R15551 gnd.n3093 gnd.n3092 0.152939
R15552 gnd.n3094 gnd.n3093 0.152939
R15553 gnd.n3094 gnd.n1841 0.152939
R15554 gnd.n3102 gnd.n1841 0.152939
R15555 gnd.n3103 gnd.n3102 0.152939
R15556 gnd.n3104 gnd.n3103 0.152939
R15557 gnd.n3104 gnd.n1835 0.152939
R15558 gnd.n3112 gnd.n1835 0.152939
R15559 gnd.n3113 gnd.n3112 0.152939
R15560 gnd.n3114 gnd.n3113 0.152939
R15561 gnd.n3114 gnd.n1829 0.152939
R15562 gnd.n3122 gnd.n1829 0.152939
R15563 gnd.n3123 gnd.n3122 0.152939
R15564 gnd.n3124 gnd.n3123 0.152939
R15565 gnd.n3124 gnd.n1823 0.152939
R15566 gnd.n3132 gnd.n1823 0.152939
R15567 gnd.n3133 gnd.n3132 0.152939
R15568 gnd.n3134 gnd.n3133 0.152939
R15569 gnd.n3134 gnd.n1817 0.152939
R15570 gnd.n3142 gnd.n1817 0.152939
R15571 gnd.n3143 gnd.n3142 0.152939
R15572 gnd.n3144 gnd.n3143 0.152939
R15573 gnd.n3144 gnd.n1811 0.152939
R15574 gnd.n5318 gnd.n1811 0.152939
R15575 gnd.n5319 gnd.n5318 0.152939
R15576 gnd.n5320 gnd.n5319 0.152939
R15577 gnd.n6161 gnd.n1220 0.152939
R15578 gnd.n6175 gnd.n1220 0.152939
R15579 gnd.n6176 gnd.n6175 0.152939
R15580 gnd.n6177 gnd.n6176 0.152939
R15581 gnd.n6177 gnd.n1206 0.152939
R15582 gnd.n6191 gnd.n1206 0.152939
R15583 gnd.n6192 gnd.n6191 0.152939
R15584 gnd.n6193 gnd.n6192 0.152939
R15585 gnd.n6193 gnd.n1191 0.152939
R15586 gnd.n6207 gnd.n1191 0.152939
R15587 gnd.n6208 gnd.n6207 0.152939
R15588 gnd.n6209 gnd.n6208 0.152939
R15589 gnd.n6209 gnd.n1177 0.152939
R15590 gnd.n6223 gnd.n1177 0.152939
R15591 gnd.n6224 gnd.n6223 0.152939
R15592 gnd.n6225 gnd.n6224 0.152939
R15593 gnd.n6225 gnd.n1163 0.152939
R15594 gnd.n6239 gnd.n1163 0.152939
R15595 gnd.n6240 gnd.n6239 0.152939
R15596 gnd.n6241 gnd.n6240 0.152939
R15597 gnd.n6241 gnd.n1148 0.152939
R15598 gnd.n6255 gnd.n1148 0.152939
R15599 gnd.n6256 gnd.n6255 0.152939
R15600 gnd.n6257 gnd.n6256 0.152939
R15601 gnd.n6257 gnd.n1133 0.152939
R15602 gnd.n6271 gnd.n1133 0.152939
R15603 gnd.n6272 gnd.n6271 0.152939
R15604 gnd.n6273 gnd.n6272 0.152939
R15605 gnd.n6273 gnd.n1119 0.152939
R15606 gnd.n6287 gnd.n1119 0.152939
R15607 gnd.n6288 gnd.n6287 0.152939
R15608 gnd.n6289 gnd.n6288 0.152939
R15609 gnd.n6289 gnd.n1106 0.152939
R15610 gnd.n6303 gnd.n1106 0.152939
R15611 gnd.n6304 gnd.n6303 0.152939
R15612 gnd.n6305 gnd.n6304 0.152939
R15613 gnd.n6305 gnd.n1092 0.152939
R15614 gnd.n6319 gnd.n1092 0.152939
R15615 gnd.n6320 gnd.n6319 0.152939
R15616 gnd.n6321 gnd.n6320 0.152939
R15617 gnd.n6321 gnd.n1076 0.152939
R15618 gnd.n6335 gnd.n1076 0.152939
R15619 gnd.n6336 gnd.n6335 0.152939
R15620 gnd.n6343 gnd.n6336 0.152939
R15621 gnd.n6343 gnd.n6342 0.152939
R15622 gnd.n6342 gnd.n6341 0.152939
R15623 gnd.n6341 gnd.n6337 0.152939
R15624 gnd.n6337 gnd.n1039 0.152939
R15625 gnd.n6401 gnd.n1039 0.152939
R15626 gnd.n6401 gnd.n6400 0.152939
R15627 gnd.n6400 gnd.n6399 0.152939
R15628 gnd.n6399 gnd.n1040 0.152939
R15629 gnd.n1040 gnd.n1000 0.152939
R15630 gnd.n6459 gnd.n1000 0.152939
R15631 gnd.n6459 gnd.n6458 0.152939
R15632 gnd.n6458 gnd.n6457 0.152939
R15633 gnd.n6457 gnd.n1001 0.152939
R15634 gnd.n6453 gnd.n1001 0.152939
R15635 gnd.n6453 gnd.n6452 0.152939
R15636 gnd.n6452 gnd.n915 0.152939
R15637 gnd.n6911 gnd.n915 0.152939
R15638 gnd.n6912 gnd.n6911 0.152939
R15639 gnd.n6913 gnd.n6912 0.152939
R15640 gnd.n6913 gnd.n901 0.152939
R15641 gnd.n6927 gnd.n901 0.152939
R15642 gnd.n6928 gnd.n6927 0.152939
R15643 gnd.n6929 gnd.n6928 0.152939
R15644 gnd.n6929 gnd.n888 0.152939
R15645 gnd.n6943 gnd.n888 0.152939
R15646 gnd.n6944 gnd.n6943 0.152939
R15647 gnd.n6945 gnd.n6944 0.152939
R15648 gnd.n6945 gnd.n874 0.152939
R15649 gnd.n6959 gnd.n874 0.152939
R15650 gnd.n6960 gnd.n6959 0.152939
R15651 gnd.n6961 gnd.n6960 0.152939
R15652 gnd.n6961 gnd.n859 0.152939
R15653 gnd.n6975 gnd.n859 0.152939
R15654 gnd.n6976 gnd.n6975 0.152939
R15655 gnd.n6977 gnd.n6976 0.152939
R15656 gnd.n6977 gnd.n845 0.152939
R15657 gnd.n6991 gnd.n845 0.152939
R15658 gnd.n6992 gnd.n6991 0.152939
R15659 gnd.n6993 gnd.n6992 0.152939
R15660 gnd.n6993 gnd.n831 0.152939
R15661 gnd.n7007 gnd.n831 0.152939
R15662 gnd.n7008 gnd.n7007 0.152939
R15663 gnd.n7009 gnd.n7008 0.152939
R15664 gnd.n7009 gnd.n817 0.152939
R15665 gnd.n7023 gnd.n817 0.152939
R15666 gnd.n7024 gnd.n7023 0.152939
R15667 gnd.n7025 gnd.n7024 0.152939
R15668 gnd.n7025 gnd.n802 0.152939
R15669 gnd.n7039 gnd.n802 0.152939
R15670 gnd.n7040 gnd.n7039 0.152939
R15671 gnd.n7041 gnd.n7040 0.152939
R15672 gnd.n7041 gnd.n789 0.152939
R15673 gnd.n7058 gnd.n789 0.152939
R15674 gnd.n7059 gnd.n7058 0.152939
R15675 gnd.n7060 gnd.n7059 0.152939
R15676 gnd.n7060 gnd.n741 0.152939
R15677 gnd.n7097 gnd.n741 0.152939
R15678 gnd.n3539 gnd.n3538 0.152939
R15679 gnd.n3538 gnd.n3534 0.152939
R15680 gnd.n3534 gnd.n1763 0.152939
R15681 gnd.n5360 gnd.n1763 0.152939
R15682 gnd.n5361 gnd.n5360 0.152939
R15683 gnd.n5363 gnd.n5361 0.152939
R15684 gnd.n5363 gnd.n5362 0.152939
R15685 gnd.n5362 gnd.n1728 0.152939
R15686 gnd.n5405 gnd.n1728 0.152939
R15687 gnd.n5406 gnd.n5405 0.152939
R15688 gnd.n5408 gnd.n5406 0.152939
R15689 gnd.n5408 gnd.n5407 0.152939
R15690 gnd.n5407 gnd.n1689 0.152939
R15691 gnd.n5455 gnd.n1689 0.152939
R15692 gnd.n5456 gnd.n5455 0.152939
R15693 gnd.n5457 gnd.n5456 0.152939
R15694 gnd.n5457 gnd.n1686 0.152939
R15695 gnd.n5462 gnd.n1686 0.152939
R15696 gnd.n5463 gnd.n5462 0.152939
R15697 gnd.n5465 gnd.n5463 0.152939
R15698 gnd.n5465 gnd.n5464 0.152939
R15699 gnd.n5464 gnd.n1624 0.152939
R15700 gnd.n5558 gnd.n1624 0.152939
R15701 gnd.n5559 gnd.n5558 0.152939
R15702 gnd.n5574 gnd.n5559 0.152939
R15703 gnd.n5574 gnd.n5573 0.152939
R15704 gnd.n5573 gnd.n5572 0.152939
R15705 gnd.n5572 gnd.n5560 0.152939
R15706 gnd.n5568 gnd.n5560 0.152939
R15707 gnd.n5568 gnd.n5567 0.152939
R15708 gnd.n5567 gnd.n5566 0.152939
R15709 gnd.n5742 gnd.n1453 0.152939
R15710 gnd.n5735 gnd.n1453 0.152939
R15711 gnd.n5735 gnd.n5734 0.152939
R15712 gnd.n5734 gnd.n5733 0.152939
R15713 gnd.n5733 gnd.n1473 0.152939
R15714 gnd.n5729 gnd.n1473 0.152939
R15715 gnd.n5744 gnd.n5743 0.152939
R15716 gnd.n5744 gnd.n1450 0.152939
R15717 gnd.n5749 gnd.n1450 0.152939
R15718 gnd.n5750 gnd.n5749 0.152939
R15719 gnd.n5751 gnd.n5750 0.152939
R15720 gnd.n5751 gnd.n1447 0.152939
R15721 gnd.n5756 gnd.n1447 0.152939
R15722 gnd.n5757 gnd.n5756 0.152939
R15723 gnd.n5758 gnd.n5757 0.152939
R15724 gnd.n5758 gnd.n1444 0.152939
R15725 gnd.n5763 gnd.n1444 0.152939
R15726 gnd.n5764 gnd.n5763 0.152939
R15727 gnd.n5765 gnd.n5764 0.152939
R15728 gnd.n5765 gnd.n1441 0.152939
R15729 gnd.n5770 gnd.n1441 0.152939
R15730 gnd.n5771 gnd.n5770 0.152939
R15731 gnd.n5772 gnd.n5771 0.152939
R15732 gnd.n5772 gnd.n1437 0.152939
R15733 gnd.n5777 gnd.n1437 0.152939
R15734 gnd.n5778 gnd.n5777 0.152939
R15735 gnd.n6019 gnd.n5778 0.152939
R15736 gnd.n6019 gnd.n6018 0.152939
R15737 gnd.n6018 gnd.n6017 0.152939
R15738 gnd.n6017 gnd.n5779 0.152939
R15739 gnd.n6013 gnd.n5779 0.152939
R15740 gnd.n6013 gnd.n6012 0.152939
R15741 gnd.n6012 gnd.n6011 0.152939
R15742 gnd.n6011 gnd.n5783 0.152939
R15743 gnd.n6007 gnd.n5783 0.152939
R15744 gnd.n6007 gnd.n6006 0.152939
R15745 gnd.n6006 gnd.n6005 0.152939
R15746 gnd.n6005 gnd.n5787 0.152939
R15747 gnd.n6001 gnd.n5787 0.152939
R15748 gnd.n6001 gnd.n6000 0.152939
R15749 gnd.n6000 gnd.n5999 0.152939
R15750 gnd.n5999 gnd.n5791 0.152939
R15751 gnd.n5995 gnd.n5791 0.152939
R15752 gnd.n5995 gnd.n5994 0.152939
R15753 gnd.n5994 gnd.n5993 0.152939
R15754 gnd.n5993 gnd.n5795 0.152939
R15755 gnd.n5989 gnd.n5795 0.152939
R15756 gnd.n5989 gnd.n5988 0.152939
R15757 gnd.n5988 gnd.n5987 0.152939
R15758 gnd.n5987 gnd.n5799 0.152939
R15759 gnd.n5983 gnd.n5799 0.152939
R15760 gnd.n5983 gnd.n5982 0.152939
R15761 gnd.n5982 gnd.n5981 0.152939
R15762 gnd.n5981 gnd.n5974 0.152939
R15763 gnd.n5977 gnd.n5974 0.152939
R15764 gnd.n5977 gnd.n1020 0.152939
R15765 gnd.n6417 gnd.n1020 0.152939
R15766 gnd.n6418 gnd.n6417 0.152939
R15767 gnd.n6420 gnd.n6418 0.152939
R15768 gnd.n6420 gnd.n6419 0.152939
R15769 gnd.n6419 gnd.n980 0.152939
R15770 gnd.n6475 gnd.n980 0.152939
R15771 gnd.n6476 gnd.n6475 0.152939
R15772 gnd.n6477 gnd.n6476 0.152939
R15773 gnd.n6477 gnd.n977 0.152939
R15774 gnd.n6482 gnd.n977 0.152939
R15775 gnd.n6483 gnd.n6482 0.152939
R15776 gnd.n6484 gnd.n6483 0.152939
R15777 gnd.n6484 gnd.n975 0.152939
R15778 gnd.n6489 gnd.n975 0.152939
R15779 gnd.n6490 gnd.n6489 0.152939
R15780 gnd.n6491 gnd.n6490 0.152939
R15781 gnd.n6491 gnd.n973 0.152939
R15782 gnd.n6496 gnd.n973 0.152939
R15783 gnd.n6497 gnd.n6496 0.152939
R15784 gnd.n6854 gnd.n6497 0.152939
R15785 gnd.n6854 gnd.n6853 0.152939
R15786 gnd.n6853 gnd.n6852 0.152939
R15787 gnd.n6852 gnd.n6498 0.152939
R15788 gnd.n6848 gnd.n6498 0.152939
R15789 gnd.n6848 gnd.n6847 0.152939
R15790 gnd.n6847 gnd.n6846 0.152939
R15791 gnd.n6846 gnd.n6502 0.152939
R15792 gnd.n6842 gnd.n6502 0.152939
R15793 gnd.n6842 gnd.n6841 0.152939
R15794 gnd.n6841 gnd.n6840 0.152939
R15795 gnd.n6840 gnd.n6506 0.152939
R15796 gnd.n6836 gnd.n6506 0.152939
R15797 gnd.n6836 gnd.n6835 0.152939
R15798 gnd.n6835 gnd.n6834 0.152939
R15799 gnd.n6834 gnd.n6795 0.152939
R15800 gnd.n6830 gnd.n6795 0.152939
R15801 gnd.n6830 gnd.n6829 0.152939
R15802 gnd.n6829 gnd.n6828 0.152939
R15803 gnd.n6828 gnd.n6799 0.152939
R15804 gnd.n6824 gnd.n6799 0.152939
R15805 gnd.n6824 gnd.n6823 0.152939
R15806 gnd.n6823 gnd.n6822 0.152939
R15807 gnd.n6822 gnd.n6803 0.152939
R15808 gnd.n6818 gnd.n6803 0.152939
R15809 gnd.n6818 gnd.n6817 0.152939
R15810 gnd.n6817 gnd.n6816 0.152939
R15811 gnd.n6816 gnd.n6807 0.152939
R15812 gnd.n6812 gnd.n6807 0.152939
R15813 gnd.n6812 gnd.n6811 0.152939
R15814 gnd.n6811 gnd.n751 0.152939
R15815 gnd.n7091 gnd.n751 0.152939
R15816 gnd.n7090 gnd.n752 0.152939
R15817 gnd.n7086 gnd.n752 0.152939
R15818 gnd.n7086 gnd.n7085 0.152939
R15819 gnd.n7085 gnd.n7084 0.152939
R15820 gnd.n7084 gnd.n756 0.152939
R15821 gnd.n756 gnd.n677 0.152939
R15822 gnd.n7100 gnd.n540 0.152939
R15823 gnd.n7323 gnd.n540 0.152939
R15824 gnd.n7324 gnd.n7323 0.152939
R15825 gnd.n7326 gnd.n7324 0.152939
R15826 gnd.n7326 gnd.n7325 0.152939
R15827 gnd.n7325 gnd.n509 0.152939
R15828 gnd.n7365 gnd.n509 0.152939
R15829 gnd.n7366 gnd.n7365 0.152939
R15830 gnd.n7368 gnd.n7366 0.152939
R15831 gnd.n7368 gnd.n7367 0.152939
R15832 gnd.n7367 gnd.n474 0.152939
R15833 gnd.n7414 gnd.n474 0.152939
R15834 gnd.n7415 gnd.n7414 0.152939
R15835 gnd.n7417 gnd.n7415 0.152939
R15836 gnd.n7417 gnd.n7416 0.152939
R15837 gnd.n7416 gnd.n443 0.152939
R15838 gnd.n7451 gnd.n443 0.152939
R15839 gnd.n7452 gnd.n7451 0.152939
R15840 gnd.n7454 gnd.n7452 0.152939
R15841 gnd.n7454 gnd.n7453 0.152939
R15842 gnd.n7453 gnd.n408 0.152939
R15843 gnd.n7500 gnd.n408 0.152939
R15844 gnd.n7501 gnd.n7500 0.152939
R15845 gnd.n7505 gnd.n7501 0.152939
R15846 gnd.n7505 gnd.n7504 0.152939
R15847 gnd.n7504 gnd.n7503 0.152939
R15848 gnd.n7503 gnd.n373 0.152939
R15849 gnd.n7548 gnd.n373 0.152939
R15850 gnd.n7549 gnd.n7548 0.152939
R15851 gnd.n7550 gnd.n7549 0.152939
R15852 gnd.n7550 gnd.n99 0.152939
R15853 gnd.n7982 gnd.n7981 0.145814
R15854 gnd.n3540 gnd.n3531 0.145814
R15855 gnd.n3540 gnd.n3539 0.145814
R15856 gnd.n7982 gnd.n99 0.145814
R15857 gnd.n5729 gnd.n5728 0.128549
R15858 gnd.n7158 gnd.n677 0.128549
R15859 gnd.n4710 gnd.n4709 0.0767195
R15860 gnd.n4709 gnd.n4708 0.0767195
R15861 gnd.n5728 gnd.n5608 0.063
R15862 gnd.n7159 gnd.n7158 0.063
R15863 gnd.n5276 gnd.n3860 0.0477147
R15864 gnd.n4473 gnd.n4361 0.0442063
R15865 gnd.n4474 gnd.n4473 0.0442063
R15866 gnd.n4475 gnd.n4474 0.0442063
R15867 gnd.n4475 gnd.n4350 0.0442063
R15868 gnd.n4489 gnd.n4350 0.0442063
R15869 gnd.n4490 gnd.n4489 0.0442063
R15870 gnd.n4491 gnd.n4490 0.0442063
R15871 gnd.n4491 gnd.n4337 0.0442063
R15872 gnd.n4535 gnd.n4337 0.0442063
R15873 gnd.n4536 gnd.n4535 0.0442063
R15874 gnd.n7159 gnd.n557 0.0416005
R15875 gnd.n7763 gnd.n7762 0.0416005
R15876 gnd.n3714 gnd.n3713 0.0416005
R15877 gnd.n5608 gnd.n5607 0.0416005
R15878 gnd.n4538 gnd.n4271 0.0344674
R15879 gnd.n7306 gnd.n557 0.0344674
R15880 gnd.n7306 gnd.n563 0.0344674
R15881 gnd.n563 gnd.n562 0.0344674
R15882 gnd.n562 gnd.n534 0.0344674
R15883 gnd.n534 gnd.n529 0.0344674
R15884 gnd.n530 gnd.n529 0.0344674
R15885 gnd.n531 gnd.n530 0.0344674
R15886 gnd.n7345 gnd.n531 0.0344674
R15887 gnd.n7345 gnd.n532 0.0344674
R15888 gnd.n532 gnd.n493 0.0344674
R15889 gnd.n494 gnd.n493 0.0344674
R15890 gnd.n495 gnd.n494 0.0344674
R15891 gnd.n496 gnd.n495 0.0344674
R15892 gnd.n496 gnd.n468 0.0344674
R15893 gnd.n468 gnd.n463 0.0344674
R15894 gnd.n464 gnd.n463 0.0344674
R15895 gnd.n465 gnd.n464 0.0344674
R15896 gnd.n7431 gnd.n465 0.0344674
R15897 gnd.n7431 gnd.n466 0.0344674
R15898 gnd.n466 gnd.n427 0.0344674
R15899 gnd.n428 gnd.n427 0.0344674
R15900 gnd.n429 gnd.n428 0.0344674
R15901 gnd.n7479 gnd.n429 0.0344674
R15902 gnd.n7479 gnd.n430 0.0344674
R15903 gnd.n430 gnd.n389 0.0344674
R15904 gnd.n390 gnd.n389 0.0344674
R15905 gnd.n391 gnd.n390 0.0344674
R15906 gnd.n392 gnd.n391 0.0344674
R15907 gnd.n7527 gnd.n392 0.0344674
R15908 gnd.n7527 gnd.n361 0.0344674
R15909 gnd.n7564 gnd.n361 0.0344674
R15910 gnd.n7565 gnd.n7564 0.0344674
R15911 gnd.n7565 gnd.n356 0.0344674
R15912 gnd.n356 gnd.n354 0.0344674
R15913 gnd.n7576 gnd.n354 0.0344674
R15914 gnd.n7577 gnd.n7576 0.0344674
R15915 gnd.n7577 gnd.n128 0.0344674
R15916 gnd.n129 gnd.n128 0.0344674
R15917 gnd.n130 gnd.n129 0.0344674
R15918 gnd.n7585 gnd.n130 0.0344674
R15919 gnd.n7585 gnd.n145 0.0344674
R15920 gnd.n146 gnd.n145 0.0344674
R15921 gnd.n147 gnd.n146 0.0344674
R15922 gnd.n7592 gnd.n147 0.0344674
R15923 gnd.n7592 gnd.n165 0.0344674
R15924 gnd.n166 gnd.n165 0.0344674
R15925 gnd.n167 gnd.n166 0.0344674
R15926 gnd.n7599 gnd.n167 0.0344674
R15927 gnd.n7599 gnd.n183 0.0344674
R15928 gnd.n184 gnd.n183 0.0344674
R15929 gnd.n185 gnd.n184 0.0344674
R15930 gnd.n7606 gnd.n185 0.0344674
R15931 gnd.n7606 gnd.n203 0.0344674
R15932 gnd.n204 gnd.n203 0.0344674
R15933 gnd.n205 gnd.n204 0.0344674
R15934 gnd.n7745 gnd.n205 0.0344674
R15935 gnd.n7745 gnd.n221 0.0344674
R15936 gnd.n222 gnd.n221 0.0344674
R15937 gnd.n223 gnd.n222 0.0344674
R15938 gnd.n7752 gnd.n223 0.0344674
R15939 gnd.n7752 gnd.n241 0.0344674
R15940 gnd.n242 gnd.n241 0.0344674
R15941 gnd.n243 gnd.n242 0.0344674
R15942 gnd.n7762 gnd.n243 0.0344674
R15943 gnd.n3713 gnd.n3272 0.0344674
R15944 gnd.n3551 gnd.n3272 0.0344674
R15945 gnd.n3551 gnd.n3294 0.0344674
R15946 gnd.n3295 gnd.n3294 0.0344674
R15947 gnd.n3296 gnd.n3295 0.0344674
R15948 gnd.n3557 gnd.n3296 0.0344674
R15949 gnd.n3557 gnd.n3313 0.0344674
R15950 gnd.n3314 gnd.n3313 0.0344674
R15951 gnd.n3315 gnd.n3314 0.0344674
R15952 gnd.n3564 gnd.n3315 0.0344674
R15953 gnd.n3564 gnd.n3332 0.0344674
R15954 gnd.n3333 gnd.n3332 0.0344674
R15955 gnd.n3334 gnd.n3333 0.0344674
R15956 gnd.n3571 gnd.n3334 0.0344674
R15957 gnd.n3571 gnd.n3351 0.0344674
R15958 gnd.n3352 gnd.n3351 0.0344674
R15959 gnd.n3353 gnd.n3352 0.0344674
R15960 gnd.n3578 gnd.n3353 0.0344674
R15961 gnd.n3578 gnd.n3370 0.0344674
R15962 gnd.n3371 gnd.n3370 0.0344674
R15963 gnd.n3372 gnd.n3371 0.0344674
R15964 gnd.n3585 gnd.n3372 0.0344674
R15965 gnd.n3585 gnd.n3389 0.0344674
R15966 gnd.n3390 gnd.n3389 0.0344674
R15967 gnd.n3391 gnd.n3390 0.0344674
R15968 gnd.n3549 gnd.n3391 0.0344674
R15969 gnd.n3626 gnd.n3549 0.0344674
R15970 gnd.n3626 gnd.n3550 0.0344674
R15971 gnd.n3550 gnd.n1788 0.0344674
R15972 gnd.n1789 gnd.n1788 0.0344674
R15973 gnd.n1790 gnd.n1789 0.0344674
R15974 gnd.n3593 gnd.n1790 0.0344674
R15975 gnd.n3593 gnd.n1800 0.0344674
R15976 gnd.n1801 gnd.n1800 0.0344674
R15977 gnd.n1802 gnd.n1801 0.0344674
R15978 gnd.n3594 gnd.n1802 0.0344674
R15979 gnd.n3609 gnd.n3594 0.0344674
R15980 gnd.n3609 gnd.n3608 0.0344674
R15981 gnd.n3608 gnd.n1758 0.0344674
R15982 gnd.n1758 gnd.n1747 0.0344674
R15983 gnd.n1748 gnd.n1747 0.0344674
R15984 gnd.n1749 gnd.n1748 0.0344674
R15985 gnd.n1750 gnd.n1749 0.0344674
R15986 gnd.n1750 gnd.n1723 0.0344674
R15987 gnd.n1723 gnd.n1709 0.0344674
R15988 gnd.n1710 gnd.n1709 0.0344674
R15989 gnd.n1711 gnd.n1710 0.0344674
R15990 gnd.n1712 gnd.n1711 0.0344674
R15991 gnd.n5415 gnd.n1712 0.0344674
R15992 gnd.n5415 gnd.n1674 0.0344674
R15993 gnd.n1675 gnd.n1674 0.0344674
R15994 gnd.n5472 gnd.n1675 0.0344674
R15995 gnd.n5472 gnd.n1676 0.0344674
R15996 gnd.n1676 gnd.n1644 0.0344674
R15997 gnd.n1645 gnd.n1644 0.0344674
R15998 gnd.n1646 gnd.n1645 0.0344674
R15999 gnd.n1647 gnd.n1646 0.0344674
R16000 gnd.n1647 gnd.n1618 0.0344674
R16001 gnd.n5581 gnd.n1618 0.0344674
R16002 gnd.n5581 gnd.n1598 0.0344674
R16003 gnd.n5598 gnd.n1598 0.0344674
R16004 gnd.n5599 gnd.n5598 0.0344674
R16005 gnd.n5599 gnd.n1591 0.0344674
R16006 gnd.n5607 gnd.n1591 0.0344674
R16007 gnd.n5727 gnd.n5726 0.0343753
R16008 gnd.n7157 gnd.n678 0.0343753
R16009 gnd.n6157 gnd.n1233 0.0296328
R16010 gnd.n7102 gnd.n7101 0.0296328
R16011 gnd.n4558 gnd.n4557 0.0269946
R16012 gnd.n4560 gnd.n4559 0.0269946
R16013 gnd.n4266 gnd.n4264 0.0269946
R16014 gnd.n4570 gnd.n4568 0.0269946
R16015 gnd.n4569 gnd.n4245 0.0269946
R16016 gnd.n4589 gnd.n4588 0.0269946
R16017 gnd.n4591 gnd.n4590 0.0269946
R16018 gnd.n4240 gnd.n4239 0.0269946
R16019 gnd.n4601 gnd.n4235 0.0269946
R16020 gnd.n4600 gnd.n4237 0.0269946
R16021 gnd.n4236 gnd.n4218 0.0269946
R16022 gnd.n4621 gnd.n4219 0.0269946
R16023 gnd.n4620 gnd.n4220 0.0269946
R16024 gnd.n4654 gnd.n4195 0.0269946
R16025 gnd.n4656 gnd.n4655 0.0269946
R16026 gnd.n4657 gnd.n4142 0.0269946
R16027 gnd.n4190 gnd.n4143 0.0269946
R16028 gnd.n4192 gnd.n4144 0.0269946
R16029 gnd.n4667 gnd.n4666 0.0269946
R16030 gnd.n4669 gnd.n4668 0.0269946
R16031 gnd.n4670 gnd.n4164 0.0269946
R16032 gnd.n4672 gnd.n4165 0.0269946
R16033 gnd.n4675 gnd.n4166 0.0269946
R16034 gnd.n4678 gnd.n4677 0.0269946
R16035 gnd.n4680 gnd.n4679 0.0269946
R16036 gnd.n4745 gnd.n4033 0.0269946
R16037 gnd.n4747 gnd.n4746 0.0269946
R16038 gnd.n4756 gnd.n4026 0.0269946
R16039 gnd.n4758 gnd.n4757 0.0269946
R16040 gnd.n4759 gnd.n4024 0.0269946
R16041 gnd.n4766 gnd.n4762 0.0269946
R16042 gnd.n4765 gnd.n4764 0.0269946
R16043 gnd.n4763 gnd.n4003 0.0269946
R16044 gnd.n4788 gnd.n4004 0.0269946
R16045 gnd.n4787 gnd.n4005 0.0269946
R16046 gnd.n4830 gnd.n3978 0.0269946
R16047 gnd.n4832 gnd.n4831 0.0269946
R16048 gnd.n4841 gnd.n3971 0.0269946
R16049 gnd.n4843 gnd.n4842 0.0269946
R16050 gnd.n4844 gnd.n3969 0.0269946
R16051 gnd.n4851 gnd.n4847 0.0269946
R16052 gnd.n4850 gnd.n4849 0.0269946
R16053 gnd.n4848 gnd.n3948 0.0269946
R16054 gnd.n4873 gnd.n3949 0.0269946
R16055 gnd.n4872 gnd.n3950 0.0269946
R16056 gnd.n4919 gnd.n3924 0.0269946
R16057 gnd.n4921 gnd.n4920 0.0269946
R16058 gnd.n4930 gnd.n3917 0.0269946
R16059 gnd.n5189 gnd.n3915 0.0269946
R16060 gnd.n5194 gnd.n5192 0.0269946
R16061 gnd.n5193 gnd.n3896 0.0269946
R16062 gnd.n5218 gnd.n5217 0.0269946
R16063 gnd.n5723 gnd.n5609 0.022519
R16064 gnd.n5722 gnd.n5613 0.022519
R16065 gnd.n5719 gnd.n5718 0.022519
R16066 gnd.n5715 gnd.n5620 0.022519
R16067 gnd.n5714 gnd.n5626 0.022519
R16068 gnd.n5711 gnd.n5710 0.022519
R16069 gnd.n5707 gnd.n5632 0.022519
R16070 gnd.n5706 gnd.n5636 0.022519
R16071 gnd.n5703 gnd.n5702 0.022519
R16072 gnd.n5699 gnd.n5643 0.022519
R16073 gnd.n5698 gnd.n5649 0.022519
R16074 gnd.n5695 gnd.n5694 0.022519
R16075 gnd.n5691 gnd.n5655 0.022519
R16076 gnd.n5690 gnd.n5659 0.022519
R16077 gnd.n5687 gnd.n5686 0.022519
R16078 gnd.n5683 gnd.n5666 0.022519
R16079 gnd.n5682 gnd.n5676 0.022519
R16080 gnd.n5673 gnd.n1236 0.022519
R16081 gnd.n6157 gnd.n6156 0.022519
R16082 gnd.n7153 gnd.n684 0.022519
R16083 gnd.n7152 gnd.n685 0.022519
R16084 gnd.n7149 gnd.n7148 0.022519
R16085 gnd.n7145 gnd.n690 0.022519
R16086 gnd.n7144 gnd.n694 0.022519
R16087 gnd.n7141 gnd.n7140 0.022519
R16088 gnd.n7137 gnd.n700 0.022519
R16089 gnd.n7136 gnd.n704 0.022519
R16090 gnd.n7133 gnd.n7132 0.022519
R16091 gnd.n7129 gnd.n708 0.022519
R16092 gnd.n7128 gnd.n712 0.022519
R16093 gnd.n7125 gnd.n7124 0.022519
R16094 gnd.n7121 gnd.n718 0.022519
R16095 gnd.n7120 gnd.n722 0.022519
R16096 gnd.n7117 gnd.n7116 0.022519
R16097 gnd.n7113 gnd.n726 0.022519
R16098 gnd.n7112 gnd.n732 0.022519
R16099 gnd.n7106 gnd.n7105 0.022519
R16100 gnd.n7102 gnd.n736 0.022519
R16101 gnd.n7101 gnd.n7098 0.0218415
R16102 gnd.n6160 gnd.n1233 0.0218415
R16103 gnd.n4538 gnd.n4537 0.0202011
R16104 gnd.n4537 gnd.n4536 0.0148637
R16105 gnd.n5187 gnd.n4931 0.0144266
R16106 gnd.n5188 gnd.n5187 0.0130679
R16107 gnd.n5726 gnd.n5609 0.0123564
R16108 gnd.n5723 gnd.n5722 0.0123564
R16109 gnd.n5719 gnd.n5613 0.0123564
R16110 gnd.n5718 gnd.n5620 0.0123564
R16111 gnd.n5715 gnd.n5714 0.0123564
R16112 gnd.n5711 gnd.n5626 0.0123564
R16113 gnd.n5710 gnd.n5632 0.0123564
R16114 gnd.n5707 gnd.n5706 0.0123564
R16115 gnd.n5703 gnd.n5636 0.0123564
R16116 gnd.n5702 gnd.n5643 0.0123564
R16117 gnd.n5699 gnd.n5698 0.0123564
R16118 gnd.n5695 gnd.n5649 0.0123564
R16119 gnd.n5694 gnd.n5655 0.0123564
R16120 gnd.n5691 gnd.n5690 0.0123564
R16121 gnd.n5687 gnd.n5659 0.0123564
R16122 gnd.n5686 gnd.n5666 0.0123564
R16123 gnd.n5683 gnd.n5682 0.0123564
R16124 gnd.n5676 gnd.n5673 0.0123564
R16125 gnd.n6156 gnd.n1236 0.0123564
R16126 gnd.n684 gnd.n678 0.0123564
R16127 gnd.n7153 gnd.n7152 0.0123564
R16128 gnd.n7149 gnd.n685 0.0123564
R16129 gnd.n7148 gnd.n690 0.0123564
R16130 gnd.n7145 gnd.n7144 0.0123564
R16131 gnd.n7141 gnd.n694 0.0123564
R16132 gnd.n7140 gnd.n700 0.0123564
R16133 gnd.n7137 gnd.n7136 0.0123564
R16134 gnd.n7133 gnd.n704 0.0123564
R16135 gnd.n7132 gnd.n708 0.0123564
R16136 gnd.n7129 gnd.n7128 0.0123564
R16137 gnd.n7125 gnd.n712 0.0123564
R16138 gnd.n7124 gnd.n718 0.0123564
R16139 gnd.n7121 gnd.n7120 0.0123564
R16140 gnd.n7117 gnd.n722 0.0123564
R16141 gnd.n7116 gnd.n726 0.0123564
R16142 gnd.n7113 gnd.n7112 0.0123564
R16143 gnd.n7106 gnd.n732 0.0123564
R16144 gnd.n7105 gnd.n736 0.0123564
R16145 gnd.n4557 gnd.n4271 0.00797283
R16146 gnd.n4559 gnd.n4558 0.00797283
R16147 gnd.n4560 gnd.n4266 0.00797283
R16148 gnd.n4568 gnd.n4264 0.00797283
R16149 gnd.n4570 gnd.n4569 0.00797283
R16150 gnd.n4588 gnd.n4245 0.00797283
R16151 gnd.n4590 gnd.n4589 0.00797283
R16152 gnd.n4591 gnd.n4240 0.00797283
R16153 gnd.n4239 gnd.n4235 0.00797283
R16154 gnd.n4601 gnd.n4600 0.00797283
R16155 gnd.n4237 gnd.n4236 0.00797283
R16156 gnd.n4219 gnd.n4218 0.00797283
R16157 gnd.n4621 gnd.n4620 0.00797283
R16158 gnd.n4220 gnd.n4195 0.00797283
R16159 gnd.n4655 gnd.n4654 0.00797283
R16160 gnd.n4657 gnd.n4656 0.00797283
R16161 gnd.n4190 gnd.n4142 0.00797283
R16162 gnd.n4192 gnd.n4143 0.00797283
R16163 gnd.n4666 gnd.n4144 0.00797283
R16164 gnd.n4668 gnd.n4667 0.00797283
R16165 gnd.n4670 gnd.n4669 0.00797283
R16166 gnd.n4672 gnd.n4164 0.00797283
R16167 gnd.n4675 gnd.n4165 0.00797283
R16168 gnd.n4677 gnd.n4166 0.00797283
R16169 gnd.n4680 gnd.n4678 0.00797283
R16170 gnd.n4679 gnd.n4033 0.00797283
R16171 gnd.n4747 gnd.n4745 0.00797283
R16172 gnd.n4746 gnd.n4026 0.00797283
R16173 gnd.n4757 gnd.n4756 0.00797283
R16174 gnd.n4759 gnd.n4758 0.00797283
R16175 gnd.n4762 gnd.n4024 0.00797283
R16176 gnd.n4766 gnd.n4765 0.00797283
R16177 gnd.n4764 gnd.n4763 0.00797283
R16178 gnd.n4004 gnd.n4003 0.00797283
R16179 gnd.n4788 gnd.n4787 0.00797283
R16180 gnd.n4005 gnd.n3978 0.00797283
R16181 gnd.n4832 gnd.n4830 0.00797283
R16182 gnd.n4831 gnd.n3971 0.00797283
R16183 gnd.n4842 gnd.n4841 0.00797283
R16184 gnd.n4844 gnd.n4843 0.00797283
R16185 gnd.n4847 gnd.n3969 0.00797283
R16186 gnd.n4851 gnd.n4850 0.00797283
R16187 gnd.n4849 gnd.n4848 0.00797283
R16188 gnd.n3949 gnd.n3948 0.00797283
R16189 gnd.n4873 gnd.n4872 0.00797283
R16190 gnd.n3950 gnd.n3924 0.00797283
R16191 gnd.n4921 gnd.n4919 0.00797283
R16192 gnd.n4920 gnd.n3917 0.00797283
R16193 gnd.n4931 gnd.n4930 0.00797283
R16194 gnd.n5189 gnd.n5188 0.00797283
R16195 gnd.n5192 gnd.n3915 0.00797283
R16196 gnd.n5194 gnd.n5193 0.00797283
R16197 gnd.n5217 gnd.n3896 0.00797283
R16198 gnd.n5218 gnd.n3860 0.00797283
R16199 gnd.n5728 gnd.n5727 0.00592005
R16200 gnd.n7158 gnd.n7157 0.00592005
R16201 plus.n53 plus.t20 323.478
R16202 plus.n11 plus.t15 323.478
R16203 plus.n52 plus.t19 297.12
R16204 plus.n56 plus.t26 297.12
R16205 plus.n58 plus.t25 297.12
R16206 plus.n62 plus.t27 297.12
R16207 plus.n64 plus.t9 297.12
R16208 plus.n68 plus.t7 297.12
R16209 plus.n70 plus.t14 297.12
R16210 plus.n74 plus.t12 297.12
R16211 plus.n76 plus.t28 297.12
R16212 plus.n80 plus.t10 297.12
R16213 plus.n82 plus.t8 297.12
R16214 plus.n40 plus.t21 297.12
R16215 plus.n38 plus.t22 297.12
R16216 plus.n2 plus.t16 297.12
R16217 plus.n32 plus.t17 297.12
R16218 plus.n4 plus.t11 297.12
R16219 plus.n26 plus.t5 297.12
R16220 plus.n6 plus.t6 297.12
R16221 plus.n20 plus.t23 297.12
R16222 plus.n8 plus.t24 297.12
R16223 plus.n14 plus.t18 297.12
R16224 plus.n10 plus.t13 297.12
R16225 plus.n86 plus.t2 243.97
R16226 plus.n86 plus.n85 223.454
R16227 plus.n88 plus.n87 223.454
R16228 plus.n83 plus.n82 161.3
R16229 plus.n81 plus.n42 161.3
R16230 plus.n80 plus.n79 161.3
R16231 plus.n78 plus.n43 161.3
R16232 plus.n77 plus.n76 161.3
R16233 plus.n75 plus.n44 161.3
R16234 plus.n74 plus.n73 161.3
R16235 plus.n72 plus.n45 161.3
R16236 plus.n71 plus.n70 161.3
R16237 plus.n69 plus.n46 161.3
R16238 plus.n68 plus.n67 161.3
R16239 plus.n66 plus.n47 161.3
R16240 plus.n65 plus.n64 161.3
R16241 plus.n63 plus.n48 161.3
R16242 plus.n62 plus.n61 161.3
R16243 plus.n60 plus.n49 161.3
R16244 plus.n59 plus.n58 161.3
R16245 plus.n57 plus.n50 161.3
R16246 plus.n56 plus.n55 161.3
R16247 plus.n54 plus.n51 161.3
R16248 plus.n13 plus.n12 161.3
R16249 plus.n14 plus.n9 161.3
R16250 plus.n16 plus.n15 161.3
R16251 plus.n17 plus.n8 161.3
R16252 plus.n19 plus.n18 161.3
R16253 plus.n20 plus.n7 161.3
R16254 plus.n22 plus.n21 161.3
R16255 plus.n23 plus.n6 161.3
R16256 plus.n25 plus.n24 161.3
R16257 plus.n26 plus.n5 161.3
R16258 plus.n28 plus.n27 161.3
R16259 plus.n29 plus.n4 161.3
R16260 plus.n31 plus.n30 161.3
R16261 plus.n32 plus.n3 161.3
R16262 plus.n34 plus.n33 161.3
R16263 plus.n35 plus.n2 161.3
R16264 plus.n37 plus.n36 161.3
R16265 plus.n38 plus.n1 161.3
R16266 plus.n39 plus.n0 161.3
R16267 plus.n41 plus.n40 161.3
R16268 plus.n82 plus.n81 46.0096
R16269 plus.n40 plus.n39 46.0096
R16270 plus.n54 plus.n53 45.0871
R16271 plus.n12 plus.n11 45.0871
R16272 plus.n52 plus.n51 41.6278
R16273 plus.n80 plus.n43 41.6278
R16274 plus.n38 plus.n37 41.6278
R16275 plus.n13 plus.n10 41.6278
R16276 plus.n57 plus.n56 37.246
R16277 plus.n76 plus.n75 37.246
R16278 plus.n33 plus.n2 37.246
R16279 plus.n15 plus.n14 37.246
R16280 plus.n84 plus.n83 33.1766
R16281 plus.n58 plus.n49 32.8641
R16282 plus.n74 plus.n45 32.8641
R16283 plus.n32 plus.n31 32.8641
R16284 plus.n19 plus.n8 32.8641
R16285 plus.n63 plus.n62 28.4823
R16286 plus.n70 plus.n69 28.4823
R16287 plus.n27 plus.n4 28.4823
R16288 plus.n21 plus.n20 28.4823
R16289 plus.n64 plus.n47 24.1005
R16290 plus.n68 plus.n47 24.1005
R16291 plus.n26 plus.n25 24.1005
R16292 plus.n25 plus.n6 24.1005
R16293 plus.n85 plus.t3 19.8005
R16294 plus.n85 plus.t1 19.8005
R16295 plus.n87 plus.t4 19.8005
R16296 plus.n87 plus.t0 19.8005
R16297 plus.n64 plus.n63 19.7187
R16298 plus.n69 plus.n68 19.7187
R16299 plus.n27 plus.n26 19.7187
R16300 plus.n21 plus.n6 19.7187
R16301 plus.n62 plus.n49 15.3369
R16302 plus.n70 plus.n45 15.3369
R16303 plus.n31 plus.n4 15.3369
R16304 plus.n20 plus.n19 15.3369
R16305 plus plus.n89 15.1953
R16306 plus.n53 plus.n52 14.1472
R16307 plus.n11 plus.n10 14.1472
R16308 plus.n84 plus.n41 11.8774
R16309 plus.n58 plus.n57 10.955
R16310 plus.n75 plus.n74 10.955
R16311 plus.n33 plus.n32 10.955
R16312 plus.n15 plus.n8 10.955
R16313 plus.n56 plus.n51 6.57323
R16314 plus.n76 plus.n43 6.57323
R16315 plus.n37 plus.n2 6.57323
R16316 plus.n14 plus.n13 6.57323
R16317 plus.n89 plus.n88 5.40567
R16318 plus.n81 plus.n80 2.19141
R16319 plus.n39 plus.n38 2.19141
R16320 plus.n89 plus.n84 1.188
R16321 plus.n88 plus.n86 0.716017
R16322 plus.n55 plus.n54 0.189894
R16323 plus.n55 plus.n50 0.189894
R16324 plus.n59 plus.n50 0.189894
R16325 plus.n60 plus.n59 0.189894
R16326 plus.n61 plus.n60 0.189894
R16327 plus.n61 plus.n48 0.189894
R16328 plus.n65 plus.n48 0.189894
R16329 plus.n66 plus.n65 0.189894
R16330 plus.n67 plus.n66 0.189894
R16331 plus.n67 plus.n46 0.189894
R16332 plus.n71 plus.n46 0.189894
R16333 plus.n72 plus.n71 0.189894
R16334 plus.n73 plus.n72 0.189894
R16335 plus.n73 plus.n44 0.189894
R16336 plus.n77 plus.n44 0.189894
R16337 plus.n78 plus.n77 0.189894
R16338 plus.n79 plus.n78 0.189894
R16339 plus.n79 plus.n42 0.189894
R16340 plus.n83 plus.n42 0.189894
R16341 plus.n41 plus.n0 0.189894
R16342 plus.n1 plus.n0 0.189894
R16343 plus.n36 plus.n1 0.189894
R16344 plus.n36 plus.n35 0.189894
R16345 plus.n35 plus.n34 0.189894
R16346 plus.n34 plus.n3 0.189894
R16347 plus.n30 plus.n3 0.189894
R16348 plus.n30 plus.n29 0.189894
R16349 plus.n29 plus.n28 0.189894
R16350 plus.n28 plus.n5 0.189894
R16351 plus.n24 plus.n5 0.189894
R16352 plus.n24 plus.n23 0.189894
R16353 plus.n23 plus.n22 0.189894
R16354 plus.n22 plus.n7 0.189894
R16355 plus.n18 plus.n7 0.189894
R16356 plus.n18 plus.n17 0.189894
R16357 plus.n17 plus.n16 0.189894
R16358 plus.n16 plus.n9 0.189894
R16359 plus.n12 plus.n9 0.189894
R16360 a_n3827_n3924.n9 a_n3827_n3924.t45 214.994
R16361 a_n3827_n3924.n5 a_n3827_n3924.t52 214.786
R16362 a_n3827_n3924.n5 a_n3827_n3924.t57 214.321
R16363 a_n3827_n3924.n5 a_n3827_n3924.t4 214.321
R16364 a_n3827_n3924.n5 a_n3827_n3924.t53 214.321
R16365 a_n3827_n3924.n7 a_n3827_n3924.t41 214.321
R16366 a_n3827_n3924.n7 a_n3827_n3924.t49 214.321
R16367 a_n3827_n3924.n8 a_n3827_n3924.t48 214.321
R16368 a_n3827_n3924.n9 a_n3827_n3924.t42 214.321
R16369 a_n3827_n3924.n9 a_n3827_n3924.t54 214.321
R16370 a_n3827_n3924.n1 a_n3827_n3924.t21 55.8337
R16371 a_n3827_n3924.n1 a_n3827_n3924.t55 55.8337
R16372 a_n3827_n3924.n11 a_n3827_n3924.t34 55.8337
R16373 a_n3827_n3924.n0 a_n3827_n3924.t11 55.8335
R16374 a_n3827_n3924.n10 a_n3827_n3924.t46 55.8335
R16375 a_n3827_n3924.n4 a_n3827_n3924.t3 55.8335
R16376 a_n3827_n3924.n4 a_n3827_n3924.t15 55.8335
R16377 a_n3827_n3924.n3 a_n3827_n3924.t12 55.8335
R16378 a_n3827_n3924.n0 a_n3827_n3924.n27 53.0052
R16379 a_n3827_n3924.n0 a_n3827_n3924.n28 53.0052
R16380 a_n3827_n3924.n0 a_n3827_n3924.n29 53.0052
R16381 a_n3827_n3924.n1 a_n3827_n3924.n30 53.0052
R16382 a_n3827_n3924.n1 a_n3827_n3924.n31 53.0052
R16383 a_n3827_n3924.n1 a_n3827_n3924.n32 53.0052
R16384 a_n3827_n3924.n6 a_n3827_n3924.n12 53.0052
R16385 a_n3827_n3924.n6 a_n3827_n3924.n13 53.0052
R16386 a_n3827_n3924.n11 a_n3827_n3924.n14 53.0052
R16387 a_n3827_n3924.n10 a_n3827_n3924.n25 53.0051
R16388 a_n3827_n3924.n2 a_n3827_n3924.n24 53.0051
R16389 a_n3827_n3924.n2 a_n3827_n3924.n23 53.0051
R16390 a_n3827_n3924.n2 a_n3827_n3924.n22 53.0051
R16391 a_n3827_n3924.n2 a_n3827_n3924.n21 53.0051
R16392 a_n3827_n3924.n4 a_n3827_n3924.n20 53.0051
R16393 a_n3827_n3924.n4 a_n3827_n3924.n19 53.0051
R16394 a_n3827_n3924.n4 a_n3827_n3924.n18 53.0051
R16395 a_n3827_n3924.n3 a_n3827_n3924.n17 53.0051
R16396 a_n3827_n3924.n3 a_n3827_n3924.n16 53.0051
R16397 a_n3827_n3924.n33 a_n3827_n3924.n1 53.0051
R16398 a_n3827_n3924.n15 a_n3827_n3924.n11 12.1986
R16399 a_n3827_n3924.n0 a_n3827_n3924.n26 12.1986
R16400 a_n3827_n3924.n3 a_n3827_n3924.n15 5.11903
R16401 a_n3827_n3924.n26 a_n3827_n3924.n10 5.11903
R16402 a_n3827_n3924.n27 a_n3827_n3924.t6 2.82907
R16403 a_n3827_n3924.n27 a_n3827_n3924.t20 2.82907
R16404 a_n3827_n3924.n28 a_n3827_n3924.t25 2.82907
R16405 a_n3827_n3924.n28 a_n3827_n3924.t10 2.82907
R16406 a_n3827_n3924.n29 a_n3827_n3924.t23 2.82907
R16407 a_n3827_n3924.n29 a_n3827_n3924.t16 2.82907
R16408 a_n3827_n3924.n30 a_n3827_n3924.t9 2.82907
R16409 a_n3827_n3924.n30 a_n3827_n3924.t13 2.82907
R16410 a_n3827_n3924.n31 a_n3827_n3924.t7 2.82907
R16411 a_n3827_n3924.n31 a_n3827_n3924.t5 2.82907
R16412 a_n3827_n3924.n32 a_n3827_n3924.t44 2.82907
R16413 a_n3827_n3924.n32 a_n3827_n3924.t1 2.82907
R16414 a_n3827_n3924.n12 a_n3827_n3924.t31 2.82907
R16415 a_n3827_n3924.n12 a_n3827_n3924.t43 2.82907
R16416 a_n3827_n3924.n13 a_n3827_n3924.t56 2.82907
R16417 a_n3827_n3924.n13 a_n3827_n3924.t38 2.82907
R16418 a_n3827_n3924.n14 a_n3827_n3924.t36 2.82907
R16419 a_n3827_n3924.n14 a_n3827_n3924.t2 2.82907
R16420 a_n3827_n3924.n25 a_n3827_n3924.t29 2.82907
R16421 a_n3827_n3924.n25 a_n3827_n3924.t37 2.82907
R16422 a_n3827_n3924.n24 a_n3827_n3924.t33 2.82907
R16423 a_n3827_n3924.n24 a_n3827_n3924.t39 2.82907
R16424 a_n3827_n3924.n23 a_n3827_n3924.t35 2.82907
R16425 a_n3827_n3924.n23 a_n3827_n3924.t30 2.82907
R16426 a_n3827_n3924.n22 a_n3827_n3924.t51 2.82907
R16427 a_n3827_n3924.n22 a_n3827_n3924.t40 2.82907
R16428 a_n3827_n3924.n21 a_n3827_n3924.t47 2.82907
R16429 a_n3827_n3924.n21 a_n3827_n3924.t50 2.82907
R16430 a_n3827_n3924.n20 a_n3827_n3924.t26 2.82907
R16431 a_n3827_n3924.n20 a_n3827_n3924.t28 2.82907
R16432 a_n3827_n3924.n19 a_n3827_n3924.t22 2.82907
R16433 a_n3827_n3924.n19 a_n3827_n3924.t19 2.82907
R16434 a_n3827_n3924.n18 a_n3827_n3924.t8 2.82907
R16435 a_n3827_n3924.n18 a_n3827_n3924.t14 2.82907
R16436 a_n3827_n3924.n17 a_n3827_n3924.t18 2.82907
R16437 a_n3827_n3924.n17 a_n3827_n3924.t17 2.82907
R16438 a_n3827_n3924.n16 a_n3827_n3924.t24 2.82907
R16439 a_n3827_n3924.n16 a_n3827_n3924.t27 2.82907
R16440 a_n3827_n3924.t0 a_n3827_n3924.n33 2.82907
R16441 a_n3827_n3924.n33 a_n3827_n3924.t32 2.82907
R16442 a_n3827_n3924.n1 a_n3827_n3924.n0 2.66429
R16443 a_n3827_n3924.n7 a_n3827_n3924.n5 2.22216
R16444 a_n3827_n3924.n2 a_n3827_n3924.n4 2.01128
R16445 a_n3827_n3924.n26 a_n3827_n3924.n5 1.95694
R16446 a_n3827_n3924.n15 a_n3827_n3924.n9 1.95694
R16447 a_n3827_n3924.n4 a_n3827_n3924.n3 1.77636
R16448 a_n3827_n3924.n10 a_n3827_n3924.n2 1.77636
R16449 a_n3827_n3924.n1 a_n3827_n3924.n6 1.56731
R16450 a_n3827_n3924.n8 a_n3827_n3924.n7 1.34352
R16451 a_n3827_n3924.n9 a_n3827_n3924.n8 1.34352
R16452 a_n3827_n3924.n11 a_n3827_n3924.n6 1.3324
R16453 a_n7636_8799.n99 a_n7636_8799.t58 485.149
R16454 a_n7636_8799.n121 a_n7636_8799.t61 485.149
R16455 a_n7636_8799.n144 a_n7636_8799.t76 485.149
R16456 a_n7636_8799.n31 a_n7636_8799.t87 485.149
R16457 a_n7636_8799.n53 a_n7636_8799.t94 485.149
R16458 a_n7636_8799.n76 a_n7636_8799.t75 485.149
R16459 a_n7636_8799.n114 a_n7636_8799.t50 464.166
R16460 a_n7636_8799.n113 a_n7636_8799.t49 464.166
R16461 a_n7636_8799.n95 a_n7636_8799.t80 464.166
R16462 a_n7636_8799.n107 a_n7636_8799.t57 464.166
R16463 a_n7636_8799.n106 a_n7636_8799.t51 464.166
R16464 a_n7636_8799.n98 a_n7636_8799.t84 464.166
R16465 a_n7636_8799.n100 a_n7636_8799.t67 464.166
R16466 a_n7636_8799.n136 a_n7636_8799.t53 464.166
R16467 a_n7636_8799.n135 a_n7636_8799.t52 464.166
R16468 a_n7636_8799.n117 a_n7636_8799.t91 464.166
R16469 a_n7636_8799.n129 a_n7636_8799.t60 464.166
R16470 a_n7636_8799.n128 a_n7636_8799.t56 464.166
R16471 a_n7636_8799.n120 a_n7636_8799.t92 464.166
R16472 a_n7636_8799.n122 a_n7636_8799.t74 464.166
R16473 a_n7636_8799.n159 a_n7636_8799.t73 464.166
R16474 a_n7636_8799.n158 a_n7636_8799.t79 464.166
R16475 a_n7636_8799.n140 a_n7636_8799.t55 464.166
R16476 a_n7636_8799.n152 a_n7636_8799.t90 464.166
R16477 a_n7636_8799.n151 a_n7636_8799.t63 464.166
R16478 a_n7636_8799.n143 a_n7636_8799.t85 464.166
R16479 a_n7636_8799.n145 a_n7636_8799.t59 464.166
R16480 a_n7636_8799.n32 a_n7636_8799.t88 464.166
R16481 a_n7636_8799.n34 a_n7636_8799.t66 464.166
R16482 a_n7636_8799.n38 a_n7636_8799.t78 464.166
R16483 a_n7636_8799.n39 a_n7636_8799.t86 464.166
R16484 a_n7636_8799.n27 a_n7636_8799.t64 464.166
R16485 a_n7636_8799.n45 a_n7636_8799.t65 464.166
R16486 a_n7636_8799.n46 a_n7636_8799.t77 464.166
R16487 a_n7636_8799.n54 a_n7636_8799.t95 464.166
R16488 a_n7636_8799.n56 a_n7636_8799.t71 464.166
R16489 a_n7636_8799.n60 a_n7636_8799.t83 464.166
R16490 a_n7636_8799.n61 a_n7636_8799.t93 464.166
R16491 a_n7636_8799.n49 a_n7636_8799.t69 464.166
R16492 a_n7636_8799.n67 a_n7636_8799.t70 464.166
R16493 a_n7636_8799.n68 a_n7636_8799.t81 464.166
R16494 a_n7636_8799.n77 a_n7636_8799.t68 464.166
R16495 a_n7636_8799.n79 a_n7636_8799.t82 464.166
R16496 a_n7636_8799.n83 a_n7636_8799.t62 464.166
R16497 a_n7636_8799.n84 a_n7636_8799.t89 464.166
R16498 a_n7636_8799.n72 a_n7636_8799.t54 464.166
R16499 a_n7636_8799.n90 a_n7636_8799.t48 464.166
R16500 a_n7636_8799.n91 a_n7636_8799.t72 464.166
R16501 a_n7636_8799.n102 a_n7636_8799.n101 161.3
R16502 a_n7636_8799.n103 a_n7636_8799.n98 161.3
R16503 a_n7636_8799.n105 a_n7636_8799.n104 161.3
R16504 a_n7636_8799.n106 a_n7636_8799.n97 161.3
R16505 a_n7636_8799.n107 a_n7636_8799.n96 161.3
R16506 a_n7636_8799.n109 a_n7636_8799.n108 161.3
R16507 a_n7636_8799.n110 a_n7636_8799.n95 161.3
R16508 a_n7636_8799.n112 a_n7636_8799.n111 161.3
R16509 a_n7636_8799.n113 a_n7636_8799.n94 161.3
R16510 a_n7636_8799.n115 a_n7636_8799.n114 161.3
R16511 a_n7636_8799.n124 a_n7636_8799.n123 161.3
R16512 a_n7636_8799.n125 a_n7636_8799.n120 161.3
R16513 a_n7636_8799.n127 a_n7636_8799.n126 161.3
R16514 a_n7636_8799.n128 a_n7636_8799.n119 161.3
R16515 a_n7636_8799.n129 a_n7636_8799.n118 161.3
R16516 a_n7636_8799.n131 a_n7636_8799.n130 161.3
R16517 a_n7636_8799.n132 a_n7636_8799.n117 161.3
R16518 a_n7636_8799.n134 a_n7636_8799.n133 161.3
R16519 a_n7636_8799.n135 a_n7636_8799.n116 161.3
R16520 a_n7636_8799.n137 a_n7636_8799.n136 161.3
R16521 a_n7636_8799.n147 a_n7636_8799.n146 161.3
R16522 a_n7636_8799.n148 a_n7636_8799.n143 161.3
R16523 a_n7636_8799.n150 a_n7636_8799.n149 161.3
R16524 a_n7636_8799.n151 a_n7636_8799.n142 161.3
R16525 a_n7636_8799.n152 a_n7636_8799.n141 161.3
R16526 a_n7636_8799.n154 a_n7636_8799.n153 161.3
R16527 a_n7636_8799.n155 a_n7636_8799.n140 161.3
R16528 a_n7636_8799.n157 a_n7636_8799.n156 161.3
R16529 a_n7636_8799.n158 a_n7636_8799.n139 161.3
R16530 a_n7636_8799.n160 a_n7636_8799.n159 161.3
R16531 a_n7636_8799.n47 a_n7636_8799.n46 161.3
R16532 a_n7636_8799.n45 a_n7636_8799.n26 161.3
R16533 a_n7636_8799.n44 a_n7636_8799.n43 161.3
R16534 a_n7636_8799.n42 a_n7636_8799.n27 161.3
R16535 a_n7636_8799.n41 a_n7636_8799.n40 161.3
R16536 a_n7636_8799.n39 a_n7636_8799.n28 161.3
R16537 a_n7636_8799.n38 a_n7636_8799.n37 161.3
R16538 a_n7636_8799.n36 a_n7636_8799.n29 161.3
R16539 a_n7636_8799.n35 a_n7636_8799.n34 161.3
R16540 a_n7636_8799.n33 a_n7636_8799.n30 161.3
R16541 a_n7636_8799.n69 a_n7636_8799.n68 161.3
R16542 a_n7636_8799.n67 a_n7636_8799.n48 161.3
R16543 a_n7636_8799.n66 a_n7636_8799.n65 161.3
R16544 a_n7636_8799.n64 a_n7636_8799.n49 161.3
R16545 a_n7636_8799.n63 a_n7636_8799.n62 161.3
R16546 a_n7636_8799.n61 a_n7636_8799.n50 161.3
R16547 a_n7636_8799.n60 a_n7636_8799.n59 161.3
R16548 a_n7636_8799.n58 a_n7636_8799.n51 161.3
R16549 a_n7636_8799.n57 a_n7636_8799.n56 161.3
R16550 a_n7636_8799.n55 a_n7636_8799.n52 161.3
R16551 a_n7636_8799.n92 a_n7636_8799.n91 161.3
R16552 a_n7636_8799.n90 a_n7636_8799.n71 161.3
R16553 a_n7636_8799.n89 a_n7636_8799.n88 161.3
R16554 a_n7636_8799.n87 a_n7636_8799.n72 161.3
R16555 a_n7636_8799.n86 a_n7636_8799.n85 161.3
R16556 a_n7636_8799.n84 a_n7636_8799.n73 161.3
R16557 a_n7636_8799.n83 a_n7636_8799.n82 161.3
R16558 a_n7636_8799.n81 a_n7636_8799.n74 161.3
R16559 a_n7636_8799.n80 a_n7636_8799.n79 161.3
R16560 a_n7636_8799.n78 a_n7636_8799.n75 161.3
R16561 a_n7636_8799.n16 a_n7636_8799.n14 98.9633
R16562 a_n7636_8799.n5 a_n7636_8799.n3 98.9631
R16563 a_n7636_8799.n24 a_n7636_8799.n23 98.6055
R16564 a_n7636_8799.n22 a_n7636_8799.n21 98.6055
R16565 a_n7636_8799.n20 a_n7636_8799.n19 98.6055
R16566 a_n7636_8799.n18 a_n7636_8799.n17 98.6055
R16567 a_n7636_8799.n16 a_n7636_8799.n15 98.6055
R16568 a_n7636_8799.n5 a_n7636_8799.n4 98.6055
R16569 a_n7636_8799.n7 a_n7636_8799.n6 98.6055
R16570 a_n7636_8799.n9 a_n7636_8799.n8 98.6055
R16571 a_n7636_8799.n11 a_n7636_8799.n10 98.6055
R16572 a_n7636_8799.n13 a_n7636_8799.n12 98.6055
R16573 a_n7636_8799.n166 a_n7636_8799.n164 81.3764
R16574 a_n7636_8799.n178 a_n7636_8799.n176 81.3764
R16575 a_n7636_8799.n2 a_n7636_8799.n0 81.3764
R16576 a_n7636_8799.n183 a_n7636_8799.n182 80.9326
R16577 a_n7636_8799.n175 a_n7636_8799.n174 80.9324
R16578 a_n7636_8799.n173 a_n7636_8799.n172 80.9324
R16579 a_n7636_8799.n171 a_n7636_8799.n170 80.9324
R16580 a_n7636_8799.n168 a_n7636_8799.n167 80.9324
R16581 a_n7636_8799.n166 a_n7636_8799.n165 80.9324
R16582 a_n7636_8799.n178 a_n7636_8799.n177 80.9324
R16583 a_n7636_8799.n180 a_n7636_8799.n179 80.9324
R16584 a_n7636_8799.n2 a_n7636_8799.n1 80.9324
R16585 a_n7636_8799.n102 a_n7636_8799.n99 70.4033
R16586 a_n7636_8799.n124 a_n7636_8799.n121 70.4033
R16587 a_n7636_8799.n147 a_n7636_8799.n144 70.4033
R16588 a_n7636_8799.n31 a_n7636_8799.n30 70.4033
R16589 a_n7636_8799.n53 a_n7636_8799.n52 70.4033
R16590 a_n7636_8799.n76 a_n7636_8799.n75 70.4033
R16591 a_n7636_8799.n114 a_n7636_8799.n113 48.2005
R16592 a_n7636_8799.n107 a_n7636_8799.n106 48.2005
R16593 a_n7636_8799.n136 a_n7636_8799.n135 48.2005
R16594 a_n7636_8799.n129 a_n7636_8799.n128 48.2005
R16595 a_n7636_8799.n159 a_n7636_8799.n158 48.2005
R16596 a_n7636_8799.n152 a_n7636_8799.n151 48.2005
R16597 a_n7636_8799.n39 a_n7636_8799.n38 48.2005
R16598 a_n7636_8799.n46 a_n7636_8799.n45 48.2005
R16599 a_n7636_8799.n61 a_n7636_8799.n60 48.2005
R16600 a_n7636_8799.n68 a_n7636_8799.n67 48.2005
R16601 a_n7636_8799.n84 a_n7636_8799.n83 48.2005
R16602 a_n7636_8799.n91 a_n7636_8799.n90 48.2005
R16603 a_n7636_8799.n112 a_n7636_8799.n95 37.246
R16604 a_n7636_8799.n101 a_n7636_8799.n98 37.246
R16605 a_n7636_8799.n134 a_n7636_8799.n117 37.246
R16606 a_n7636_8799.n123 a_n7636_8799.n120 37.246
R16607 a_n7636_8799.n157 a_n7636_8799.n140 37.246
R16608 a_n7636_8799.n146 a_n7636_8799.n143 37.246
R16609 a_n7636_8799.n34 a_n7636_8799.n33 37.246
R16610 a_n7636_8799.n44 a_n7636_8799.n27 37.246
R16611 a_n7636_8799.n56 a_n7636_8799.n55 37.246
R16612 a_n7636_8799.n66 a_n7636_8799.n49 37.246
R16613 a_n7636_8799.n79 a_n7636_8799.n78 37.246
R16614 a_n7636_8799.n89 a_n7636_8799.n72 37.246
R16615 a_n7636_8799.n108 a_n7636_8799.n95 35.7853
R16616 a_n7636_8799.n105 a_n7636_8799.n98 35.7853
R16617 a_n7636_8799.n130 a_n7636_8799.n117 35.7853
R16618 a_n7636_8799.n127 a_n7636_8799.n120 35.7853
R16619 a_n7636_8799.n153 a_n7636_8799.n140 35.7853
R16620 a_n7636_8799.n150 a_n7636_8799.n143 35.7853
R16621 a_n7636_8799.n34 a_n7636_8799.n29 35.7853
R16622 a_n7636_8799.n40 a_n7636_8799.n27 35.7853
R16623 a_n7636_8799.n56 a_n7636_8799.n51 35.7853
R16624 a_n7636_8799.n62 a_n7636_8799.n49 35.7853
R16625 a_n7636_8799.n79 a_n7636_8799.n74 35.7853
R16626 a_n7636_8799.n85 a_n7636_8799.n72 35.7853
R16627 a_n7636_8799.n25 a_n7636_8799.n13 34.1553
R16628 a_n7636_8799.n181 a_n7636_8799.n175 33.4185
R16629 a_n7636_8799.n100 a_n7636_8799.n99 20.9576
R16630 a_n7636_8799.n122 a_n7636_8799.n121 20.9576
R16631 a_n7636_8799.n145 a_n7636_8799.n144 20.9576
R16632 a_n7636_8799.n32 a_n7636_8799.n31 20.9576
R16633 a_n7636_8799.n54 a_n7636_8799.n53 20.9576
R16634 a_n7636_8799.n77 a_n7636_8799.n76 20.9576
R16635 a_n7636_8799.n25 a_n7636_8799.n24 20.7339
R16636 a_n7636_8799.n108 a_n7636_8799.n107 12.4157
R16637 a_n7636_8799.n106 a_n7636_8799.n105 12.4157
R16638 a_n7636_8799.n130 a_n7636_8799.n129 12.4157
R16639 a_n7636_8799.n128 a_n7636_8799.n127 12.4157
R16640 a_n7636_8799.n153 a_n7636_8799.n152 12.4157
R16641 a_n7636_8799.n151 a_n7636_8799.n150 12.4157
R16642 a_n7636_8799.n38 a_n7636_8799.n29 12.4157
R16643 a_n7636_8799.n40 a_n7636_8799.n39 12.4157
R16644 a_n7636_8799.n60 a_n7636_8799.n51 12.4157
R16645 a_n7636_8799.n62 a_n7636_8799.n61 12.4157
R16646 a_n7636_8799.n83 a_n7636_8799.n74 12.4157
R16647 a_n7636_8799.n85 a_n7636_8799.n84 12.4157
R16648 a_n7636_8799.n169 a_n7636_8799.n163 12.3339
R16649 a_n7636_8799.n163 a_n7636_8799.n25 11.4887
R16650 a_n7636_8799.n113 a_n7636_8799.n112 10.955
R16651 a_n7636_8799.n101 a_n7636_8799.n100 10.955
R16652 a_n7636_8799.n135 a_n7636_8799.n134 10.955
R16653 a_n7636_8799.n123 a_n7636_8799.n122 10.955
R16654 a_n7636_8799.n158 a_n7636_8799.n157 10.955
R16655 a_n7636_8799.n146 a_n7636_8799.n145 10.955
R16656 a_n7636_8799.n33 a_n7636_8799.n32 10.955
R16657 a_n7636_8799.n45 a_n7636_8799.n44 10.955
R16658 a_n7636_8799.n55 a_n7636_8799.n54 10.955
R16659 a_n7636_8799.n67 a_n7636_8799.n66 10.955
R16660 a_n7636_8799.n78 a_n7636_8799.n77 10.955
R16661 a_n7636_8799.n90 a_n7636_8799.n89 10.955
R16662 a_n7636_8799.n138 a_n7636_8799.n115 9.05164
R16663 a_n7636_8799.n70 a_n7636_8799.n47 9.05164
R16664 a_n7636_8799.n162 a_n7636_8799.n93 7.2142
R16665 a_n7636_8799.n162 a_n7636_8799.n161 6.79277
R16666 a_n7636_8799.n138 a_n7636_8799.n137 4.94368
R16667 a_n7636_8799.n161 a_n7636_8799.n160 4.94368
R16668 a_n7636_8799.n70 a_n7636_8799.n69 4.94368
R16669 a_n7636_8799.n93 a_n7636_8799.n92 4.94368
R16670 a_n7636_8799.n161 a_n7636_8799.n138 4.10845
R16671 a_n7636_8799.n93 a_n7636_8799.n70 4.10845
R16672 a_n7636_8799.n23 a_n7636_8799.t43 3.61217
R16673 a_n7636_8799.n23 a_n7636_8799.t33 3.61217
R16674 a_n7636_8799.n21 a_n7636_8799.t0 3.61217
R16675 a_n7636_8799.n21 a_n7636_8799.t36 3.61217
R16676 a_n7636_8799.n19 a_n7636_8799.t37 3.61217
R16677 a_n7636_8799.n19 a_n7636_8799.t45 3.61217
R16678 a_n7636_8799.n17 a_n7636_8799.t38 3.61217
R16679 a_n7636_8799.n17 a_n7636_8799.t1 3.61217
R16680 a_n7636_8799.n15 a_n7636_8799.t41 3.61217
R16681 a_n7636_8799.n15 a_n7636_8799.t35 3.61217
R16682 a_n7636_8799.n14 a_n7636_8799.t5 3.61217
R16683 a_n7636_8799.n14 a_n7636_8799.t44 3.61217
R16684 a_n7636_8799.n3 a_n7636_8799.t47 3.61217
R16685 a_n7636_8799.n3 a_n7636_8799.t3 3.61217
R16686 a_n7636_8799.n4 a_n7636_8799.t4 3.61217
R16687 a_n7636_8799.n4 a_n7636_8799.t32 3.61217
R16688 a_n7636_8799.n6 a_n7636_8799.t31 3.61217
R16689 a_n7636_8799.n6 a_n7636_8799.t46 3.61217
R16690 a_n7636_8799.n8 a_n7636_8799.t39 3.61217
R16691 a_n7636_8799.n8 a_n7636_8799.t2 3.61217
R16692 a_n7636_8799.n10 a_n7636_8799.t42 3.61217
R16693 a_n7636_8799.n10 a_n7636_8799.t30 3.61217
R16694 a_n7636_8799.n12 a_n7636_8799.t34 3.61217
R16695 a_n7636_8799.n12 a_n7636_8799.t40 3.61217
R16696 a_n7636_8799.n163 a_n7636_8799.n162 3.4105
R16697 a_n7636_8799.n176 a_n7636_8799.t21 2.82907
R16698 a_n7636_8799.n176 a_n7636_8799.t19 2.82907
R16699 a_n7636_8799.n177 a_n7636_8799.t10 2.82907
R16700 a_n7636_8799.n177 a_n7636_8799.t16 2.82907
R16701 a_n7636_8799.n179 a_n7636_8799.t28 2.82907
R16702 a_n7636_8799.n179 a_n7636_8799.t11 2.82907
R16703 a_n7636_8799.n1 a_n7636_8799.t18 2.82907
R16704 a_n7636_8799.n1 a_n7636_8799.t17 2.82907
R16705 a_n7636_8799.n0 a_n7636_8799.t13 2.82907
R16706 a_n7636_8799.n0 a_n7636_8799.t12 2.82907
R16707 a_n7636_8799.n174 a_n7636_8799.t24 2.82907
R16708 a_n7636_8799.n174 a_n7636_8799.t26 2.82907
R16709 a_n7636_8799.n172 a_n7636_8799.t22 2.82907
R16710 a_n7636_8799.n172 a_n7636_8799.t6 2.82907
R16711 a_n7636_8799.n170 a_n7636_8799.t27 2.82907
R16712 a_n7636_8799.n170 a_n7636_8799.t20 2.82907
R16713 a_n7636_8799.n167 a_n7636_8799.t7 2.82907
R16714 a_n7636_8799.n167 a_n7636_8799.t25 2.82907
R16715 a_n7636_8799.n165 a_n7636_8799.t8 2.82907
R16716 a_n7636_8799.n165 a_n7636_8799.t9 2.82907
R16717 a_n7636_8799.n164 a_n7636_8799.t14 2.82907
R16718 a_n7636_8799.n164 a_n7636_8799.t15 2.82907
R16719 a_n7636_8799.n183 a_n7636_8799.t23 2.82907
R16720 a_n7636_8799.t29 a_n7636_8799.n183 2.82907
R16721 a_n7636_8799.n168 a_n7636_8799.n166 0.444466
R16722 a_n7636_8799.n173 a_n7636_8799.n171 0.444466
R16723 a_n7636_8799.n175 a_n7636_8799.n173 0.444466
R16724 a_n7636_8799.n182 a_n7636_8799.n2 0.444466
R16725 a_n7636_8799.n180 a_n7636_8799.n178 0.444466
R16726 a_n7636_8799.n18 a_n7636_8799.n16 0.358259
R16727 a_n7636_8799.n20 a_n7636_8799.n18 0.358259
R16728 a_n7636_8799.n22 a_n7636_8799.n20 0.358259
R16729 a_n7636_8799.n24 a_n7636_8799.n22 0.358259
R16730 a_n7636_8799.n13 a_n7636_8799.n11 0.358259
R16731 a_n7636_8799.n11 a_n7636_8799.n9 0.358259
R16732 a_n7636_8799.n9 a_n7636_8799.n7 0.358259
R16733 a_n7636_8799.n7 a_n7636_8799.n5 0.358259
R16734 a_n7636_8799.n169 a_n7636_8799.n168 0.222483
R16735 a_n7636_8799.n171 a_n7636_8799.n169 0.222483
R16736 a_n7636_8799.n182 a_n7636_8799.n181 0.222483
R16737 a_n7636_8799.n181 a_n7636_8799.n180 0.222483
R16738 a_n7636_8799.n115 a_n7636_8799.n94 0.189894
R16739 a_n7636_8799.n111 a_n7636_8799.n94 0.189894
R16740 a_n7636_8799.n111 a_n7636_8799.n110 0.189894
R16741 a_n7636_8799.n110 a_n7636_8799.n109 0.189894
R16742 a_n7636_8799.n109 a_n7636_8799.n96 0.189894
R16743 a_n7636_8799.n97 a_n7636_8799.n96 0.189894
R16744 a_n7636_8799.n104 a_n7636_8799.n97 0.189894
R16745 a_n7636_8799.n104 a_n7636_8799.n103 0.189894
R16746 a_n7636_8799.n103 a_n7636_8799.n102 0.189894
R16747 a_n7636_8799.n137 a_n7636_8799.n116 0.189894
R16748 a_n7636_8799.n133 a_n7636_8799.n116 0.189894
R16749 a_n7636_8799.n133 a_n7636_8799.n132 0.189894
R16750 a_n7636_8799.n132 a_n7636_8799.n131 0.189894
R16751 a_n7636_8799.n131 a_n7636_8799.n118 0.189894
R16752 a_n7636_8799.n119 a_n7636_8799.n118 0.189894
R16753 a_n7636_8799.n126 a_n7636_8799.n119 0.189894
R16754 a_n7636_8799.n126 a_n7636_8799.n125 0.189894
R16755 a_n7636_8799.n125 a_n7636_8799.n124 0.189894
R16756 a_n7636_8799.n160 a_n7636_8799.n139 0.189894
R16757 a_n7636_8799.n156 a_n7636_8799.n139 0.189894
R16758 a_n7636_8799.n156 a_n7636_8799.n155 0.189894
R16759 a_n7636_8799.n155 a_n7636_8799.n154 0.189894
R16760 a_n7636_8799.n154 a_n7636_8799.n141 0.189894
R16761 a_n7636_8799.n142 a_n7636_8799.n141 0.189894
R16762 a_n7636_8799.n149 a_n7636_8799.n142 0.189894
R16763 a_n7636_8799.n149 a_n7636_8799.n148 0.189894
R16764 a_n7636_8799.n148 a_n7636_8799.n147 0.189894
R16765 a_n7636_8799.n35 a_n7636_8799.n30 0.189894
R16766 a_n7636_8799.n36 a_n7636_8799.n35 0.189894
R16767 a_n7636_8799.n37 a_n7636_8799.n36 0.189894
R16768 a_n7636_8799.n37 a_n7636_8799.n28 0.189894
R16769 a_n7636_8799.n41 a_n7636_8799.n28 0.189894
R16770 a_n7636_8799.n42 a_n7636_8799.n41 0.189894
R16771 a_n7636_8799.n43 a_n7636_8799.n42 0.189894
R16772 a_n7636_8799.n43 a_n7636_8799.n26 0.189894
R16773 a_n7636_8799.n47 a_n7636_8799.n26 0.189894
R16774 a_n7636_8799.n57 a_n7636_8799.n52 0.189894
R16775 a_n7636_8799.n58 a_n7636_8799.n57 0.189894
R16776 a_n7636_8799.n59 a_n7636_8799.n58 0.189894
R16777 a_n7636_8799.n59 a_n7636_8799.n50 0.189894
R16778 a_n7636_8799.n63 a_n7636_8799.n50 0.189894
R16779 a_n7636_8799.n64 a_n7636_8799.n63 0.189894
R16780 a_n7636_8799.n65 a_n7636_8799.n64 0.189894
R16781 a_n7636_8799.n65 a_n7636_8799.n48 0.189894
R16782 a_n7636_8799.n69 a_n7636_8799.n48 0.189894
R16783 a_n7636_8799.n80 a_n7636_8799.n75 0.189894
R16784 a_n7636_8799.n81 a_n7636_8799.n80 0.189894
R16785 a_n7636_8799.n82 a_n7636_8799.n81 0.189894
R16786 a_n7636_8799.n82 a_n7636_8799.n73 0.189894
R16787 a_n7636_8799.n86 a_n7636_8799.n73 0.189894
R16788 a_n7636_8799.n87 a_n7636_8799.n86 0.189894
R16789 a_n7636_8799.n88 a_n7636_8799.n87 0.189894
R16790 a_n7636_8799.n88 a_n7636_8799.n71 0.189894
R16791 a_n7636_8799.n92 a_n7636_8799.n71 0.189894
R16792 a_n2982_13878.n125 a_n2982_13878.t94 512.366
R16793 a_n2982_13878.n115 a_n2982_13878.t83 512.366
R16794 a_n2982_13878.n126 a_n2982_13878.t72 512.366
R16795 a_n2982_13878.n123 a_n2982_13878.t102 512.366
R16796 a_n2982_13878.n116 a_n2982_13878.t91 512.366
R16797 a_n2982_13878.n124 a_n2982_13878.t90 512.366
R16798 a_n2982_13878.n121 a_n2982_13878.t98 512.366
R16799 a_n2982_13878.n117 a_n2982_13878.t81 512.366
R16800 a_n2982_13878.n122 a_n2982_13878.t82 512.366
R16801 a_n2982_13878.n119 a_n2982_13878.t85 512.366
R16802 a_n2982_13878.n118 a_n2982_13878.t96 512.366
R16803 a_n2982_13878.n120 a_n2982_13878.t111 512.366
R16804 a_n2982_13878.n31 a_n2982_13878.t110 538.698
R16805 a_n2982_13878.n134 a_n2982_13878.t87 512.366
R16806 a_n2982_13878.n133 a_n2982_13878.t92 512.366
R16807 a_n2982_13878.n86 a_n2982_13878.t80 512.366
R16808 a_n2982_13878.n132 a_n2982_13878.t97 512.366
R16809 a_n2982_13878.n131 a_n2982_13878.t106 512.366
R16810 a_n2982_13878.n87 a_n2982_13878.t107 512.366
R16811 a_n2982_13878.n130 a_n2982_13878.t74 512.366
R16812 a_n2982_13878.n129 a_n2982_13878.t89 512.366
R16813 a_n2982_13878.n88 a_n2982_13878.t77 512.366
R16814 a_n2982_13878.n128 a_n2982_13878.t84 512.366
R16815 a_n2982_13878.n33 a_n2982_13878.t18 538.699
R16816 a_n2982_13878.n135 a_n2982_13878.t32 512.366
R16817 a_n2982_13878.n83 a_n2982_13878.t50 512.366
R16818 a_n2982_13878.n38 a_n2982_13878.t44 538.698
R16819 a_n2982_13878.n153 a_n2982_13878.t6 512.366
R16820 a_n2982_13878.n152 a_n2982_13878.t10 512.366
R16821 a_n2982_13878.n84 a_n2982_13878.t46 512.366
R16822 a_n2982_13878.n151 a_n2982_13878.t24 512.366
R16823 a_n2982_13878.n150 a_n2982_13878.t48 512.366
R16824 a_n2982_13878.n85 a_n2982_13878.t52 512.366
R16825 a_n2982_13878.n149 a_n2982_13878.t16 512.366
R16826 a_n2982_13878.n148 a_n2982_13878.t12 512.366
R16827 a_n2982_13878.n19 a_n2982_13878.t8 538.698
R16828 a_n2982_13878.n108 a_n2982_13878.t26 512.366
R16829 a_n2982_13878.n97 a_n2982_13878.t36 512.366
R16830 a_n2982_13878.n109 a_n2982_13878.t14 512.366
R16831 a_n2982_13878.n96 a_n2982_13878.t22 512.366
R16832 a_n2982_13878.n110 a_n2982_13878.t20 512.366
R16833 a_n2982_13878.n111 a_n2982_13878.t38 512.366
R16834 a_n2982_13878.n95 a_n2982_13878.t40 512.366
R16835 a_n2982_13878.n112 a_n2982_13878.t30 512.366
R16836 a_n2982_13878.n94 a_n2982_13878.t34 512.366
R16837 a_n2982_13878.n113 a_n2982_13878.t42 512.366
R16838 a_n2982_13878.n25 a_n2982_13878.t109 538.698
R16839 a_n2982_13878.n102 a_n2982_13878.t78 512.366
R16840 a_n2982_13878.n101 a_n2982_13878.t79 512.366
R16841 a_n2982_13878.n103 a_n2982_13878.t104 512.366
R16842 a_n2982_13878.n100 a_n2982_13878.t105 512.366
R16843 a_n2982_13878.n104 a_n2982_13878.t76 512.366
R16844 a_n2982_13878.n105 a_n2982_13878.t100 512.366
R16845 a_n2982_13878.n99 a_n2982_13878.t101 512.366
R16846 a_n2982_13878.n106 a_n2982_13878.t73 512.366
R16847 a_n2982_13878.n98 a_n2982_13878.t86 512.366
R16848 a_n2982_13878.n107 a_n2982_13878.t95 512.366
R16849 a_n2982_13878.n5 a_n2982_13878.n82 70.1674
R16850 a_n2982_13878.n7 a_n2982_13878.n80 70.1674
R16851 a_n2982_13878.n9 a_n2982_13878.n78 70.1674
R16852 a_n2982_13878.n12 a_n2982_13878.n76 70.1674
R16853 a_n2982_13878.n58 a_n2982_13878.n26 70.5844
R16854 a_n2982_13878.n50 a_n2982_13878.n32 44.5605
R16855 a_n2982_13878.n148 a_n2982_13878.n50 21.3688
R16856 a_n2982_13878.n49 a_n2982_13878.n34 80.4688
R16857 a_n2982_13878.n49 a_n2982_13878.n149 0.365327
R16858 a_n2982_13878.n35 a_n2982_13878.n48 75.0448
R16859 a_n2982_13878.n47 a_n2982_13878.n35 70.1674
R16860 a_n2982_13878.n151 a_n2982_13878.n47 20.9683
R16861 a_n2982_13878.n37 a_n2982_13878.n46 70.3058
R16862 a_n2982_13878.n46 a_n2982_13878.n84 20.6913
R16863 a_n2982_13878.n45 a_n2982_13878.n37 75.3623
R16864 a_n2982_13878.n152 a_n2982_13878.n45 10.5784
R16865 a_n2982_13878.n36 a_n2982_13878.n38 44.7878
R16866 a_n2982_13878.n33 a_n2982_13878.n32 44.7878
R16867 a_n2982_13878.n33 a_n2982_13878.n135 14.1664
R16868 a_n2982_13878.n26 a_n2982_13878.n57 70.1674
R16869 a_n2982_13878.n57 a_n2982_13878.n88 20.9683
R16870 a_n2982_13878.n56 a_n2982_13878.n27 74.73
R16871 a_n2982_13878.n129 a_n2982_13878.n56 11.843
R16872 a_n2982_13878.n55 a_n2982_13878.n27 80.4688
R16873 a_n2982_13878.n55 a_n2982_13878.n130 0.365327
R16874 a_n2982_13878.n28 a_n2982_13878.n54 75.0448
R16875 a_n2982_13878.n53 a_n2982_13878.n28 70.1674
R16876 a_n2982_13878.n132 a_n2982_13878.n53 20.9683
R16877 a_n2982_13878.n30 a_n2982_13878.n52 70.3058
R16878 a_n2982_13878.n52 a_n2982_13878.n86 20.6913
R16879 a_n2982_13878.n51 a_n2982_13878.n30 75.3623
R16880 a_n2982_13878.n133 a_n2982_13878.n51 10.5784
R16881 a_n2982_13878.n29 a_n2982_13878.n31 44.7878
R16882 a_n2982_13878.n15 a_n2982_13878.n74 70.5844
R16883 a_n2982_13878.n21 a_n2982_13878.n66 70.5844
R16884 a_n2982_13878.n65 a_n2982_13878.n21 70.1674
R16885 a_n2982_13878.n65 a_n2982_13878.n98 20.9683
R16886 a_n2982_13878.n20 a_n2982_13878.n64 74.73
R16887 a_n2982_13878.n106 a_n2982_13878.n64 11.843
R16888 a_n2982_13878.n63 a_n2982_13878.n20 80.4688
R16889 a_n2982_13878.n63 a_n2982_13878.n99 0.365327
R16890 a_n2982_13878.n22 a_n2982_13878.n62 75.0448
R16891 a_n2982_13878.n61 a_n2982_13878.n22 70.1674
R16892 a_n2982_13878.n61 a_n2982_13878.n100 20.9683
R16893 a_n2982_13878.n23 a_n2982_13878.n60 70.3058
R16894 a_n2982_13878.n103 a_n2982_13878.n60 20.6913
R16895 a_n2982_13878.n59 a_n2982_13878.n23 75.3623
R16896 a_n2982_13878.n59 a_n2982_13878.n101 10.5784
R16897 a_n2982_13878.n25 a_n2982_13878.n24 44.7878
R16898 a_n2982_13878.n73 a_n2982_13878.n15 70.1674
R16899 a_n2982_13878.n73 a_n2982_13878.n94 20.9683
R16900 a_n2982_13878.n14 a_n2982_13878.n72 74.73
R16901 a_n2982_13878.n112 a_n2982_13878.n72 11.843
R16902 a_n2982_13878.n71 a_n2982_13878.n14 80.4688
R16903 a_n2982_13878.n71 a_n2982_13878.n95 0.365327
R16904 a_n2982_13878.n16 a_n2982_13878.n70 75.0448
R16905 a_n2982_13878.n69 a_n2982_13878.n16 70.1674
R16906 a_n2982_13878.n69 a_n2982_13878.n96 20.9683
R16907 a_n2982_13878.n17 a_n2982_13878.n68 70.3058
R16908 a_n2982_13878.n109 a_n2982_13878.n68 20.6913
R16909 a_n2982_13878.n67 a_n2982_13878.n17 75.3623
R16910 a_n2982_13878.n67 a_n2982_13878.n97 10.5784
R16911 a_n2982_13878.n19 a_n2982_13878.n18 44.7878
R16912 a_n2982_13878.n120 a_n2982_13878.n76 20.9683
R16913 a_n2982_13878.n75 a_n2982_13878.n13 75.0448
R16914 a_n2982_13878.n75 a_n2982_13878.n118 11.2134
R16915 a_n2982_13878.n13 a_n2982_13878.n119 161.3
R16916 a_n2982_13878.n122 a_n2982_13878.n78 20.9683
R16917 a_n2982_13878.n77 a_n2982_13878.n10 75.0448
R16918 a_n2982_13878.n77 a_n2982_13878.n117 11.2134
R16919 a_n2982_13878.n10 a_n2982_13878.n121 161.3
R16920 a_n2982_13878.n124 a_n2982_13878.n80 20.9683
R16921 a_n2982_13878.n79 a_n2982_13878.n8 75.0448
R16922 a_n2982_13878.n79 a_n2982_13878.n116 11.2134
R16923 a_n2982_13878.n8 a_n2982_13878.n123 161.3
R16924 a_n2982_13878.n126 a_n2982_13878.n82 20.9683
R16925 a_n2982_13878.n81 a_n2982_13878.n6 75.0448
R16926 a_n2982_13878.n81 a_n2982_13878.n115 11.2134
R16927 a_n2982_13878.n6 a_n2982_13878.n125 161.3
R16928 a_n2982_13878.n3 a_n2982_13878.n145 81.3764
R16929 a_n2982_13878.n4 a_n2982_13878.n139 81.3764
R16930 a_n2982_13878.n0 a_n2982_13878.n136 81.3764
R16931 a_n2982_13878.n3 a_n2982_13878.n146 80.9324
R16932 a_n2982_13878.n2 a_n2982_13878.n147 80.9324
R16933 a_n2982_13878.n2 a_n2982_13878.n144 80.9324
R16934 a_n2982_13878.n2 a_n2982_13878.n143 80.9324
R16935 a_n2982_13878.n1 a_n2982_13878.n142 80.9324
R16936 a_n2982_13878.n4 a_n2982_13878.n140 80.9324
R16937 a_n2982_13878.n0 a_n2982_13878.n141 80.9324
R16938 a_n2982_13878.n0 a_n2982_13878.n138 80.9324
R16939 a_n2982_13878.n0 a_n2982_13878.n137 80.9324
R16940 a_n2982_13878.n44 a_n2982_13878.t19 74.6477
R16941 a_n2982_13878.n39 a_n2982_13878.t9 74.6477
R16942 a_n2982_13878.n43 a_n2982_13878.t45 74.2899
R16943 a_n2982_13878.n41 a_n2982_13878.t29 74.2897
R16944 a_n2982_13878.n44 a_n2982_13878.n155 70.6783
R16945 a_n2982_13878.n44 a_n2982_13878.n156 70.6783
R16946 a_n2982_13878.n42 a_n2982_13878.n157 70.6783
R16947 a_n2982_13878.n42 a_n2982_13878.n158 70.6783
R16948 a_n2982_13878.n41 a_n2982_13878.n93 70.6783
R16949 a_n2982_13878.n40 a_n2982_13878.n92 70.6783
R16950 a_n2982_13878.n40 a_n2982_13878.n91 70.6783
R16951 a_n2982_13878.n39 a_n2982_13878.n90 70.6783
R16952 a_n2982_13878.n39 a_n2982_13878.n89 70.6783
R16953 a_n2982_13878.n159 a_n2982_13878.n43 70.6782
R16954 a_n2982_13878.n125 a_n2982_13878.n115 48.2005
R16955 a_n2982_13878.t99 a_n2982_13878.n82 533.335
R16956 a_n2982_13878.n123 a_n2982_13878.n116 48.2005
R16957 a_n2982_13878.t108 a_n2982_13878.n80 533.335
R16958 a_n2982_13878.n121 a_n2982_13878.n117 48.2005
R16959 a_n2982_13878.t93 a_n2982_13878.n78 533.335
R16960 a_n2982_13878.n119 a_n2982_13878.n118 48.2005
R16961 a_n2982_13878.t88 a_n2982_13878.n76 533.335
R16962 a_n2982_13878.n134 a_n2982_13878.n133 48.2005
R16963 a_n2982_13878.n53 a_n2982_13878.n131 20.9683
R16964 a_n2982_13878.n130 a_n2982_13878.n87 48.2005
R16965 a_n2982_13878.n128 a_n2982_13878.n57 20.9683
R16966 a_n2982_13878.n135 a_n2982_13878.n83 48.2005
R16967 a_n2982_13878.n153 a_n2982_13878.n152 48.2005
R16968 a_n2982_13878.n47 a_n2982_13878.n150 20.9683
R16969 a_n2982_13878.n149 a_n2982_13878.n85 48.2005
R16970 a_n2982_13878.n108 a_n2982_13878.n97 48.2005
R16971 a_n2982_13878.n110 a_n2982_13878.n69 20.9683
R16972 a_n2982_13878.n111 a_n2982_13878.n95 48.2005
R16973 a_n2982_13878.n113 a_n2982_13878.n73 20.9683
R16974 a_n2982_13878.n102 a_n2982_13878.n101 48.2005
R16975 a_n2982_13878.n104 a_n2982_13878.n61 20.9683
R16976 a_n2982_13878.n105 a_n2982_13878.n99 48.2005
R16977 a_n2982_13878.n107 a_n2982_13878.n65 20.9683
R16978 a_n2982_13878.n132 a_n2982_13878.n52 21.4216
R16979 a_n2982_13878.n151 a_n2982_13878.n46 21.4216
R16980 a_n2982_13878.n96 a_n2982_13878.n68 21.4216
R16981 a_n2982_13878.n100 a_n2982_13878.n60 21.4216
R16982 a_n2982_13878.n58 a_n2982_13878.t103 532.5
R16983 a_n2982_13878.t28 a_n2982_13878.n74 532.5
R16984 a_n2982_13878.t75 a_n2982_13878.n66 532.5
R16985 a_n2982_13878.n1 a_n2982_13878.n0 32.6799
R16986 a_n2982_13878.n56 a_n2982_13878.n88 34.4824
R16987 a_n2982_13878.n50 a_n2982_13878.n83 20.5623
R16988 a_n2982_13878.n94 a_n2982_13878.n72 34.4824
R16989 a_n2982_13878.n98 a_n2982_13878.n64 34.4824
R16990 a_n2982_13878.n126 a_n2982_13878.n81 35.3134
R16991 a_n2982_13878.n124 a_n2982_13878.n79 35.3134
R16992 a_n2982_13878.n122 a_n2982_13878.n77 35.3134
R16993 a_n2982_13878.n120 a_n2982_13878.n75 35.3134
R16994 a_n2982_13878.n131 a_n2982_13878.n54 35.3134
R16995 a_n2982_13878.n54 a_n2982_13878.n87 11.2134
R16996 a_n2982_13878.n150 a_n2982_13878.n48 35.3134
R16997 a_n2982_13878.n48 a_n2982_13878.n85 11.2134
R16998 a_n2982_13878.n70 a_n2982_13878.n110 35.3134
R16999 a_n2982_13878.n111 a_n2982_13878.n70 11.2134
R17000 a_n2982_13878.n62 a_n2982_13878.n104 35.3134
R17001 a_n2982_13878.n105 a_n2982_13878.n62 11.2134
R17002 a_n2982_13878.n32 a_n2982_13878.n2 23.891
R17003 a_n2982_13878.n51 a_n2982_13878.n86 36.139
R17004 a_n2982_13878.n45 a_n2982_13878.n84 36.139
R17005 a_n2982_13878.n109 a_n2982_13878.n67 36.139
R17006 a_n2982_13878.n103 a_n2982_13878.n59 36.139
R17007 a_n2982_13878.n24 a_n2982_13878.n11 13.9285
R17008 a_n2982_13878.n26 a_n2982_13878.n127 13.724
R17009 a_n2982_13878.n154 a_n2982_13878.n36 12.4191
R17010 a_n2982_13878.n127 a_n2982_13878.n5 11.2486
R17011 a_n2982_13878.n13 a_n2982_13878.n11 11.2486
R17012 a_n2982_13878.n114 a_n2982_13878.n41 10.5745
R17013 a_n2982_13878.n114 a_n2982_13878.n15 8.58383
R17014 a_n2982_13878.n43 a_n2982_13878.n154 6.7311
R17015 a_n2982_13878.n127 a_n2982_13878.n114 5.3452
R17016 a_n2982_13878.n32 a_n2982_13878.n29 3.94368
R17017 a_n2982_13878.n18 a_n2982_13878.n21 3.94368
R17018 a_n2982_13878.n155 a_n2982_13878.t51 3.61217
R17019 a_n2982_13878.n155 a_n2982_13878.t33 3.61217
R17020 a_n2982_13878.n156 a_n2982_13878.t17 3.61217
R17021 a_n2982_13878.n156 a_n2982_13878.t13 3.61217
R17022 a_n2982_13878.n157 a_n2982_13878.t49 3.61217
R17023 a_n2982_13878.n157 a_n2982_13878.t53 3.61217
R17024 a_n2982_13878.n158 a_n2982_13878.t47 3.61217
R17025 a_n2982_13878.n158 a_n2982_13878.t25 3.61217
R17026 a_n2982_13878.n93 a_n2982_13878.t35 3.61217
R17027 a_n2982_13878.n93 a_n2982_13878.t43 3.61217
R17028 a_n2982_13878.n92 a_n2982_13878.t41 3.61217
R17029 a_n2982_13878.n92 a_n2982_13878.t31 3.61217
R17030 a_n2982_13878.n91 a_n2982_13878.t21 3.61217
R17031 a_n2982_13878.n91 a_n2982_13878.t39 3.61217
R17032 a_n2982_13878.n90 a_n2982_13878.t15 3.61217
R17033 a_n2982_13878.n90 a_n2982_13878.t23 3.61217
R17034 a_n2982_13878.n89 a_n2982_13878.t27 3.61217
R17035 a_n2982_13878.n89 a_n2982_13878.t37 3.61217
R17036 a_n2982_13878.t7 a_n2982_13878.n159 3.61217
R17037 a_n2982_13878.n159 a_n2982_13878.t11 3.61217
R17038 a_n2982_13878.n145 a_n2982_13878.t1 2.82907
R17039 a_n2982_13878.n145 a_n2982_13878.t70 2.82907
R17040 a_n2982_13878.n146 a_n2982_13878.t55 2.82907
R17041 a_n2982_13878.n146 a_n2982_13878.t65 2.82907
R17042 a_n2982_13878.n147 a_n2982_13878.t64 2.82907
R17043 a_n2982_13878.n147 a_n2982_13878.t0 2.82907
R17044 a_n2982_13878.n144 a_n2982_13878.t61 2.82907
R17045 a_n2982_13878.n144 a_n2982_13878.t54 2.82907
R17046 a_n2982_13878.n143 a_n2982_13878.t2 2.82907
R17047 a_n2982_13878.n143 a_n2982_13878.t71 2.82907
R17048 a_n2982_13878.n142 a_n2982_13878.t57 2.82907
R17049 a_n2982_13878.n142 a_n2982_13878.t59 2.82907
R17050 a_n2982_13878.n139 a_n2982_13878.t60 2.82907
R17051 a_n2982_13878.n139 a_n2982_13878.t66 2.82907
R17052 a_n2982_13878.n140 a_n2982_13878.t62 2.82907
R17053 a_n2982_13878.n140 a_n2982_13878.t4 2.82907
R17054 a_n2982_13878.n141 a_n2982_13878.t5 2.82907
R17055 a_n2982_13878.n141 a_n2982_13878.t56 2.82907
R17056 a_n2982_13878.n138 a_n2982_13878.t63 2.82907
R17057 a_n2982_13878.n138 a_n2982_13878.t58 2.82907
R17058 a_n2982_13878.n137 a_n2982_13878.t68 2.82907
R17059 a_n2982_13878.n137 a_n2982_13878.t69 2.82907
R17060 a_n2982_13878.n136 a_n2982_13878.t3 2.82907
R17061 a_n2982_13878.n136 a_n2982_13878.t67 2.82907
R17062 a_n2982_13878.n31 a_n2982_13878.n134 14.1668
R17063 a_n2982_13878.n128 a_n2982_13878.n58 22.3251
R17064 a_n2982_13878.n38 a_n2982_13878.n153 14.1668
R17065 a_n2982_13878.n108 a_n2982_13878.n19 14.1668
R17066 a_n2982_13878.n74 a_n2982_13878.n113 22.3251
R17067 a_n2982_13878.n102 a_n2982_13878.n25 14.1668
R17068 a_n2982_13878.n66 a_n2982_13878.n107 22.3251
R17069 a_n2982_13878.n154 a_n2982_13878.n11 1.30542
R17070 a_n2982_13878.n8 a_n2982_13878.n9 1.04595
R17071 a_n2982_13878.n55 a_n2982_13878.n129 47.835
R17072 a_n2982_13878.n49 a_n2982_13878.n148 47.835
R17073 a_n2982_13878.n112 a_n2982_13878.n71 47.835
R17074 a_n2982_13878.n106 a_n2982_13878.n63 47.835
R17075 a_n2982_13878.n0 a_n2982_13878.n4 1.3324
R17076 a_n2982_13878.n27 a_n2982_13878.n26 1.13686
R17077 a_n2982_13878.n21 a_n2982_13878.n20 1.13686
R17078 a_n2982_13878.n15 a_n2982_13878.n14 1.13686
R17079 a_n2982_13878.n32 a_n2982_13878.n34 1.09898
R17080 a_n2982_13878.n43 a_n2982_13878.n42 1.07378
R17081 a_n2982_13878.n40 a_n2982_13878.n39 1.07378
R17082 a_n2982_13878.n2 a_n2982_13878.n3 0.888431
R17083 a_n2982_13878.n2 a_n2982_13878.n1 0.888431
R17084 a_n2982_13878.n37 a_n2982_13878.n36 0.758076
R17085 a_n2982_13878.n37 a_n2982_13878.n35 0.758076
R17086 a_n2982_13878.n35 a_n2982_13878.n34 0.758076
R17087 a_n2982_13878.n30 a_n2982_13878.n29 0.758076
R17088 a_n2982_13878.n30 a_n2982_13878.n28 0.758076
R17089 a_n2982_13878.n28 a_n2982_13878.n27 0.758076
R17090 a_n2982_13878.n23 a_n2982_13878.n24 0.758076
R17091 a_n2982_13878.n22 a_n2982_13878.n23 0.758076
R17092 a_n2982_13878.n20 a_n2982_13878.n22 0.758076
R17093 a_n2982_13878.n17 a_n2982_13878.n18 0.758076
R17094 a_n2982_13878.n16 a_n2982_13878.n17 0.758076
R17095 a_n2982_13878.n14 a_n2982_13878.n16 0.758076
R17096 a_n2982_13878.n13 a_n2982_13878.n12 0.758076
R17097 a_n2982_13878.n10 a_n2982_13878.n9 0.758076
R17098 a_n2982_13878.n8 a_n2982_13878.n7 0.758076
R17099 a_n2982_13878.n6 a_n2982_13878.n5 0.758076
R17100 a_n2982_13878.n42 a_n2982_13878.n44 0.716017
R17101 a_n2982_13878.n41 a_n2982_13878.n40 0.716017
R17102 a_n2982_13878.n10 a_n2982_13878.n12 0.67853
R17103 a_n2982_13878.n6 a_n2982_13878.n7 0.67853
R17104 a_n2804_13878.n29 a_n2804_13878.n28 98.9632
R17105 a_n2804_13878.n2 a_n2804_13878.n0 98.7517
R17106 a_n2804_13878.n22 a_n2804_13878.n21 98.6055
R17107 a_n2804_13878.n24 a_n2804_13878.n23 98.6055
R17108 a_n2804_13878.n26 a_n2804_13878.n25 98.6055
R17109 a_n2804_13878.n28 a_n2804_13878.n27 98.6055
R17110 a_n2804_13878.n10 a_n2804_13878.n9 98.6055
R17111 a_n2804_13878.n8 a_n2804_13878.n7 98.6055
R17112 a_n2804_13878.n6 a_n2804_13878.n5 98.6055
R17113 a_n2804_13878.n4 a_n2804_13878.n3 98.6055
R17114 a_n2804_13878.n2 a_n2804_13878.n1 98.6055
R17115 a_n2804_13878.n20 a_n2804_13878.n19 98.6054
R17116 a_n2804_13878.n12 a_n2804_13878.t30 74.6477
R17117 a_n2804_13878.n17 a_n2804_13878.t31 74.2899
R17118 a_n2804_13878.n14 a_n2804_13878.t28 74.2899
R17119 a_n2804_13878.n13 a_n2804_13878.t2 74.2899
R17120 a_n2804_13878.n16 a_n2804_13878.n15 70.6783
R17121 a_n2804_13878.n12 a_n2804_13878.n11 70.6783
R17122 a_n2804_13878.n18 a_n2804_13878.n10 15.7159
R17123 a_n2804_13878.n20 a_n2804_13878.n18 12.6495
R17124 a_n2804_13878.n18 a_n2804_13878.n17 8.38735
R17125 a_n2804_13878.n19 a_n2804_13878.t10 3.61217
R17126 a_n2804_13878.n19 a_n2804_13878.t19 3.61217
R17127 a_n2804_13878.n21 a_n2804_13878.t23 3.61217
R17128 a_n2804_13878.n21 a_n2804_13878.t9 3.61217
R17129 a_n2804_13878.n23 a_n2804_13878.t13 3.61217
R17130 a_n2804_13878.n23 a_n2804_13878.t14 3.61217
R17131 a_n2804_13878.n25 a_n2804_13878.t24 3.61217
R17132 a_n2804_13878.n25 a_n2804_13878.t25 3.61217
R17133 a_n2804_13878.n27 a_n2804_13878.t3 3.61217
R17134 a_n2804_13878.n27 a_n2804_13878.t15 3.61217
R17135 a_n2804_13878.n15 a_n2804_13878.t27 3.61217
R17136 a_n2804_13878.n15 a_n2804_13878.t1 3.61217
R17137 a_n2804_13878.n11 a_n2804_13878.t0 3.61217
R17138 a_n2804_13878.n11 a_n2804_13878.t29 3.61217
R17139 a_n2804_13878.n9 a_n2804_13878.t16 3.61217
R17140 a_n2804_13878.n9 a_n2804_13878.t4 3.61217
R17141 a_n2804_13878.n7 a_n2804_13878.t21 3.61217
R17142 a_n2804_13878.n7 a_n2804_13878.t6 3.61217
R17143 a_n2804_13878.n5 a_n2804_13878.t5 3.61217
R17144 a_n2804_13878.n5 a_n2804_13878.t8 3.61217
R17145 a_n2804_13878.n3 a_n2804_13878.t18 3.61217
R17146 a_n2804_13878.n3 a_n2804_13878.t11 3.61217
R17147 a_n2804_13878.n1 a_n2804_13878.t22 3.61217
R17148 a_n2804_13878.n1 a_n2804_13878.t12 3.61217
R17149 a_n2804_13878.n0 a_n2804_13878.t7 3.61217
R17150 a_n2804_13878.n0 a_n2804_13878.t17 3.61217
R17151 a_n2804_13878.n29 a_n2804_13878.t20 3.61217
R17152 a_n2804_13878.t26 a_n2804_13878.n29 3.61217
R17153 a_n2804_13878.n13 a_n2804_13878.n12 0.358259
R17154 a_n2804_13878.n16 a_n2804_13878.n14 0.358259
R17155 a_n2804_13878.n17 a_n2804_13878.n16 0.358259
R17156 a_n2804_13878.n28 a_n2804_13878.n26 0.358259
R17157 a_n2804_13878.n26 a_n2804_13878.n24 0.358259
R17158 a_n2804_13878.n24 a_n2804_13878.n22 0.358259
R17159 a_n2804_13878.n22 a_n2804_13878.n20 0.358259
R17160 a_n2804_13878.n4 a_n2804_13878.n2 0.146627
R17161 a_n2804_13878.n6 a_n2804_13878.n4 0.146627
R17162 a_n2804_13878.n8 a_n2804_13878.n6 0.146627
R17163 a_n2804_13878.n10 a_n2804_13878.n8 0.146627
R17164 a_n2804_13878.n14 a_n2804_13878.n13 0.101793
R17165 vdd.n291 vdd.n255 756.745
R17166 vdd.n244 vdd.n208 756.745
R17167 vdd.n201 vdd.n165 756.745
R17168 vdd.n154 vdd.n118 756.745
R17169 vdd.n112 vdd.n76 756.745
R17170 vdd.n65 vdd.n29 756.745
R17171 vdd.n1561 vdd.n1525 756.745
R17172 vdd.n1608 vdd.n1572 756.745
R17173 vdd.n1471 vdd.n1435 756.745
R17174 vdd.n1518 vdd.n1482 756.745
R17175 vdd.n1382 vdd.n1346 756.745
R17176 vdd.n1429 vdd.n1393 756.745
R17177 vdd.n1105 vdd.t71 640.208
R17178 vdd.n800 vdd.t116 640.208
R17179 vdd.n1109 vdd.t113 640.208
R17180 vdd.n791 vdd.t134 640.208
R17181 vdd.n686 vdd.t89 640.208
R17182 vdd.n2437 vdd.t131 640.208
R17183 vdd.n622 vdd.t82 640.208
R17184 vdd.n2434 vdd.t123 640.208
R17185 vdd.n589 vdd.t67 640.208
R17186 vdd.n861 vdd.t127 640.208
R17187 vdd.n1775 vdd.t104 592.009
R17188 vdd.n1813 vdd.t93 592.009
R17189 vdd.n1709 vdd.t107 592.009
R17190 vdd.n1976 vdd.t97 592.009
R17191 vdd.n1038 vdd.t75 592.009
R17192 vdd.n998 vdd.t79 592.009
R17193 vdd.n3180 vdd.t100 592.009
R17194 vdd.n405 vdd.t137 592.009
R17195 vdd.n365 vdd.t140 592.009
R17196 vdd.n557 vdd.t110 592.009
R17197 vdd.n3076 vdd.t120 592.009
R17198 vdd.n2983 vdd.t85 592.009
R17199 vdd.n292 vdd.n291 585
R17200 vdd.n290 vdd.n257 585
R17201 vdd.n289 vdd.n288 585
R17202 vdd.n260 vdd.n258 585
R17203 vdd.n283 vdd.n282 585
R17204 vdd.n281 vdd.n280 585
R17205 vdd.n264 vdd.n263 585
R17206 vdd.n275 vdd.n274 585
R17207 vdd.n273 vdd.n272 585
R17208 vdd.n268 vdd.n267 585
R17209 vdd.n245 vdd.n244 585
R17210 vdd.n243 vdd.n210 585
R17211 vdd.n242 vdd.n241 585
R17212 vdd.n213 vdd.n211 585
R17213 vdd.n236 vdd.n235 585
R17214 vdd.n234 vdd.n233 585
R17215 vdd.n217 vdd.n216 585
R17216 vdd.n228 vdd.n227 585
R17217 vdd.n226 vdd.n225 585
R17218 vdd.n221 vdd.n220 585
R17219 vdd.n202 vdd.n201 585
R17220 vdd.n200 vdd.n167 585
R17221 vdd.n199 vdd.n198 585
R17222 vdd.n170 vdd.n168 585
R17223 vdd.n193 vdd.n192 585
R17224 vdd.n191 vdd.n190 585
R17225 vdd.n174 vdd.n173 585
R17226 vdd.n185 vdd.n184 585
R17227 vdd.n183 vdd.n182 585
R17228 vdd.n178 vdd.n177 585
R17229 vdd.n155 vdd.n154 585
R17230 vdd.n153 vdd.n120 585
R17231 vdd.n152 vdd.n151 585
R17232 vdd.n123 vdd.n121 585
R17233 vdd.n146 vdd.n145 585
R17234 vdd.n144 vdd.n143 585
R17235 vdd.n127 vdd.n126 585
R17236 vdd.n138 vdd.n137 585
R17237 vdd.n136 vdd.n135 585
R17238 vdd.n131 vdd.n130 585
R17239 vdd.n113 vdd.n112 585
R17240 vdd.n111 vdd.n78 585
R17241 vdd.n110 vdd.n109 585
R17242 vdd.n81 vdd.n79 585
R17243 vdd.n104 vdd.n103 585
R17244 vdd.n102 vdd.n101 585
R17245 vdd.n85 vdd.n84 585
R17246 vdd.n96 vdd.n95 585
R17247 vdd.n94 vdd.n93 585
R17248 vdd.n89 vdd.n88 585
R17249 vdd.n66 vdd.n65 585
R17250 vdd.n64 vdd.n31 585
R17251 vdd.n63 vdd.n62 585
R17252 vdd.n34 vdd.n32 585
R17253 vdd.n57 vdd.n56 585
R17254 vdd.n55 vdd.n54 585
R17255 vdd.n38 vdd.n37 585
R17256 vdd.n49 vdd.n48 585
R17257 vdd.n47 vdd.n46 585
R17258 vdd.n42 vdd.n41 585
R17259 vdd.n1562 vdd.n1561 585
R17260 vdd.n1560 vdd.n1527 585
R17261 vdd.n1559 vdd.n1558 585
R17262 vdd.n1530 vdd.n1528 585
R17263 vdd.n1553 vdd.n1552 585
R17264 vdd.n1551 vdd.n1550 585
R17265 vdd.n1534 vdd.n1533 585
R17266 vdd.n1545 vdd.n1544 585
R17267 vdd.n1543 vdd.n1542 585
R17268 vdd.n1538 vdd.n1537 585
R17269 vdd.n1609 vdd.n1608 585
R17270 vdd.n1607 vdd.n1574 585
R17271 vdd.n1606 vdd.n1605 585
R17272 vdd.n1577 vdd.n1575 585
R17273 vdd.n1600 vdd.n1599 585
R17274 vdd.n1598 vdd.n1597 585
R17275 vdd.n1581 vdd.n1580 585
R17276 vdd.n1592 vdd.n1591 585
R17277 vdd.n1590 vdd.n1589 585
R17278 vdd.n1585 vdd.n1584 585
R17279 vdd.n1472 vdd.n1471 585
R17280 vdd.n1470 vdd.n1437 585
R17281 vdd.n1469 vdd.n1468 585
R17282 vdd.n1440 vdd.n1438 585
R17283 vdd.n1463 vdd.n1462 585
R17284 vdd.n1461 vdd.n1460 585
R17285 vdd.n1444 vdd.n1443 585
R17286 vdd.n1455 vdd.n1454 585
R17287 vdd.n1453 vdd.n1452 585
R17288 vdd.n1448 vdd.n1447 585
R17289 vdd.n1519 vdd.n1518 585
R17290 vdd.n1517 vdd.n1484 585
R17291 vdd.n1516 vdd.n1515 585
R17292 vdd.n1487 vdd.n1485 585
R17293 vdd.n1510 vdd.n1509 585
R17294 vdd.n1508 vdd.n1507 585
R17295 vdd.n1491 vdd.n1490 585
R17296 vdd.n1502 vdd.n1501 585
R17297 vdd.n1500 vdd.n1499 585
R17298 vdd.n1495 vdd.n1494 585
R17299 vdd.n1383 vdd.n1382 585
R17300 vdd.n1381 vdd.n1348 585
R17301 vdd.n1380 vdd.n1379 585
R17302 vdd.n1351 vdd.n1349 585
R17303 vdd.n1374 vdd.n1373 585
R17304 vdd.n1372 vdd.n1371 585
R17305 vdd.n1355 vdd.n1354 585
R17306 vdd.n1366 vdd.n1365 585
R17307 vdd.n1364 vdd.n1363 585
R17308 vdd.n1359 vdd.n1358 585
R17309 vdd.n1430 vdd.n1429 585
R17310 vdd.n1428 vdd.n1395 585
R17311 vdd.n1427 vdd.n1426 585
R17312 vdd.n1398 vdd.n1396 585
R17313 vdd.n1421 vdd.n1420 585
R17314 vdd.n1419 vdd.n1418 585
R17315 vdd.n1402 vdd.n1401 585
R17316 vdd.n1413 vdd.n1412 585
R17317 vdd.n1411 vdd.n1410 585
R17318 vdd.n1406 vdd.n1405 585
R17319 vdd.n3296 vdd.n330 515.122
R17320 vdd.n3178 vdd.n328 515.122
R17321 vdd.n515 vdd.n478 515.122
R17322 vdd.n3114 vdd.n479 515.122
R17323 vdd.n1971 vdd.n1320 515.122
R17324 vdd.n1974 vdd.n1973 515.122
R17325 vdd.n1682 vdd.n1646 515.122
R17326 vdd.n1878 vdd.n1647 515.122
R17327 vdd.n269 vdd.t201 329.043
R17328 vdd.n222 vdd.t209 329.043
R17329 vdd.n179 vdd.t198 329.043
R17330 vdd.n132 vdd.t206 329.043
R17331 vdd.n90 vdd.t178 329.043
R17332 vdd.n43 vdd.t183 329.043
R17333 vdd.n1539 vdd.t176 329.043
R17334 vdd.n1586 vdd.t162 329.043
R17335 vdd.n1449 vdd.t171 329.043
R17336 vdd.n1496 vdd.t151 329.043
R17337 vdd.n1360 vdd.t184 329.043
R17338 vdd.n1407 vdd.t179 329.043
R17339 vdd.n1775 vdd.t106 319.788
R17340 vdd.n1813 vdd.t96 319.788
R17341 vdd.n1709 vdd.t109 319.788
R17342 vdd.n1976 vdd.t98 319.788
R17343 vdd.n1038 vdd.t77 319.788
R17344 vdd.n998 vdd.t80 319.788
R17345 vdd.n3180 vdd.t102 319.788
R17346 vdd.n405 vdd.t138 319.788
R17347 vdd.n365 vdd.t141 319.788
R17348 vdd.n557 vdd.t112 319.788
R17349 vdd.n3076 vdd.t122 319.788
R17350 vdd.n2983 vdd.t88 319.788
R17351 vdd.n1776 vdd.t105 303.69
R17352 vdd.n1814 vdd.t95 303.69
R17353 vdd.n1710 vdd.t108 303.69
R17354 vdd.n1977 vdd.t99 303.69
R17355 vdd.n1039 vdd.t78 303.69
R17356 vdd.n999 vdd.t81 303.69
R17357 vdd.n3181 vdd.t103 303.69
R17358 vdd.n406 vdd.t139 303.69
R17359 vdd.n366 vdd.t142 303.69
R17360 vdd.n558 vdd.t111 303.69
R17361 vdd.n3077 vdd.t121 303.69
R17362 vdd.n2984 vdd.t87 303.69
R17363 vdd.n2704 vdd.n750 279.512
R17364 vdd.n2944 vdd.n599 279.512
R17365 vdd.n2881 vdd.n596 279.512
R17366 vdd.n2636 vdd.n2635 279.512
R17367 vdd.n2397 vdd.n788 279.512
R17368 vdd.n2328 vdd.n2327 279.512
R17369 vdd.n1145 vdd.n1144 279.512
R17370 vdd.n2122 vdd.n928 279.512
R17371 vdd.n2860 vdd.n597 279.512
R17372 vdd.n2947 vdd.n2946 279.512
R17373 vdd.n2509 vdd.n2432 279.512
R17374 vdd.n2440 vdd.n746 279.512
R17375 vdd.n2325 vdd.n798 279.512
R17376 vdd.n796 vdd.n770 279.512
R17377 vdd.n1270 vdd.n965 279.512
R17378 vdd.n1070 vdd.n923 279.512
R17379 vdd.n2120 vdd.n931 254.619
R17380 vdd.n3112 vdd.n484 254.619
R17381 vdd.n2862 vdd.n597 185
R17382 vdd.n2945 vdd.n597 185
R17383 vdd.n2864 vdd.n2863 185
R17384 vdd.n2863 vdd.n595 185
R17385 vdd.n2865 vdd.n629 185
R17386 vdd.n2875 vdd.n629 185
R17387 vdd.n2866 vdd.n638 185
R17388 vdd.n638 vdd.n636 185
R17389 vdd.n2868 vdd.n2867 185
R17390 vdd.n2869 vdd.n2868 185
R17391 vdd.n2821 vdd.n637 185
R17392 vdd.n637 vdd.n633 185
R17393 vdd.n2820 vdd.n2819 185
R17394 vdd.n2819 vdd.n2818 185
R17395 vdd.n640 vdd.n639 185
R17396 vdd.n641 vdd.n640 185
R17397 vdd.n2811 vdd.n2810 185
R17398 vdd.n2812 vdd.n2811 185
R17399 vdd.n2809 vdd.n649 185
R17400 vdd.n654 vdd.n649 185
R17401 vdd.n2808 vdd.n2807 185
R17402 vdd.n2807 vdd.n2806 185
R17403 vdd.n651 vdd.n650 185
R17404 vdd.n660 vdd.n651 185
R17405 vdd.n2799 vdd.n2798 185
R17406 vdd.n2800 vdd.n2799 185
R17407 vdd.n2797 vdd.n661 185
R17408 vdd.n667 vdd.n661 185
R17409 vdd.n2796 vdd.n2795 185
R17410 vdd.n2795 vdd.n2794 185
R17411 vdd.n663 vdd.n662 185
R17412 vdd.n664 vdd.n663 185
R17413 vdd.n2787 vdd.n2786 185
R17414 vdd.n2788 vdd.n2787 185
R17415 vdd.n2785 vdd.n674 185
R17416 vdd.n674 vdd.n671 185
R17417 vdd.n2784 vdd.n2783 185
R17418 vdd.n2783 vdd.n2782 185
R17419 vdd.n676 vdd.n675 185
R17420 vdd.n677 vdd.n676 185
R17421 vdd.n2775 vdd.n2774 185
R17422 vdd.n2776 vdd.n2775 185
R17423 vdd.n2773 vdd.n685 185
R17424 vdd.n691 vdd.n685 185
R17425 vdd.n2772 vdd.n2771 185
R17426 vdd.n2771 vdd.n2770 185
R17427 vdd.n2761 vdd.n688 185
R17428 vdd.n698 vdd.n688 185
R17429 vdd.n2763 vdd.n2762 185
R17430 vdd.n2764 vdd.n2763 185
R17431 vdd.n2760 vdd.n699 185
R17432 vdd.n699 vdd.n695 185
R17433 vdd.n2759 vdd.n2758 185
R17434 vdd.n2758 vdd.n2757 185
R17435 vdd.n701 vdd.n700 185
R17436 vdd.n702 vdd.n701 185
R17437 vdd.n2750 vdd.n2749 185
R17438 vdd.n2751 vdd.n2750 185
R17439 vdd.n2748 vdd.n710 185
R17440 vdd.n715 vdd.n710 185
R17441 vdd.n2747 vdd.n2746 185
R17442 vdd.n2746 vdd.n2745 185
R17443 vdd.n712 vdd.n711 185
R17444 vdd.n721 vdd.n712 185
R17445 vdd.n2738 vdd.n2737 185
R17446 vdd.n2739 vdd.n2738 185
R17447 vdd.n2736 vdd.n722 185
R17448 vdd.n2612 vdd.n722 185
R17449 vdd.n2735 vdd.n2734 185
R17450 vdd.n2734 vdd.n2733 185
R17451 vdd.n724 vdd.n723 185
R17452 vdd.n2618 vdd.n724 185
R17453 vdd.n2726 vdd.n2725 185
R17454 vdd.n2727 vdd.n2726 185
R17455 vdd.n2724 vdd.n733 185
R17456 vdd.n733 vdd.n730 185
R17457 vdd.n2723 vdd.n2722 185
R17458 vdd.n2722 vdd.n2721 185
R17459 vdd.n735 vdd.n734 185
R17460 vdd.n736 vdd.n735 185
R17461 vdd.n2714 vdd.n2713 185
R17462 vdd.n2715 vdd.n2714 185
R17463 vdd.n2712 vdd.n744 185
R17464 vdd.n2630 vdd.n744 185
R17465 vdd.n2711 vdd.n2710 185
R17466 vdd.n2710 vdd.n2709 185
R17467 vdd.n746 vdd.n745 185
R17468 vdd.n747 vdd.n746 185
R17469 vdd.n2441 vdd.n2440 185
R17470 vdd.n2443 vdd.n2442 185
R17471 vdd.n2445 vdd.n2444 185
R17472 vdd.n2447 vdd.n2446 185
R17473 vdd.n2449 vdd.n2448 185
R17474 vdd.n2451 vdd.n2450 185
R17475 vdd.n2453 vdd.n2452 185
R17476 vdd.n2455 vdd.n2454 185
R17477 vdd.n2457 vdd.n2456 185
R17478 vdd.n2459 vdd.n2458 185
R17479 vdd.n2461 vdd.n2460 185
R17480 vdd.n2463 vdd.n2462 185
R17481 vdd.n2465 vdd.n2464 185
R17482 vdd.n2467 vdd.n2466 185
R17483 vdd.n2469 vdd.n2468 185
R17484 vdd.n2471 vdd.n2470 185
R17485 vdd.n2473 vdd.n2472 185
R17486 vdd.n2475 vdd.n2474 185
R17487 vdd.n2477 vdd.n2476 185
R17488 vdd.n2479 vdd.n2478 185
R17489 vdd.n2481 vdd.n2480 185
R17490 vdd.n2483 vdd.n2482 185
R17491 vdd.n2485 vdd.n2484 185
R17492 vdd.n2487 vdd.n2486 185
R17493 vdd.n2489 vdd.n2488 185
R17494 vdd.n2491 vdd.n2490 185
R17495 vdd.n2493 vdd.n2492 185
R17496 vdd.n2495 vdd.n2494 185
R17497 vdd.n2497 vdd.n2496 185
R17498 vdd.n2499 vdd.n2498 185
R17499 vdd.n2501 vdd.n2500 185
R17500 vdd.n2503 vdd.n2502 185
R17501 vdd.n2505 vdd.n2504 185
R17502 vdd.n2507 vdd.n2506 185
R17503 vdd.n2508 vdd.n2432 185
R17504 vdd.n2702 vdd.n2432 185
R17505 vdd.n2948 vdd.n2947 185
R17506 vdd.n2949 vdd.n588 185
R17507 vdd.n2951 vdd.n2950 185
R17508 vdd.n2953 vdd.n586 185
R17509 vdd.n2955 vdd.n2954 185
R17510 vdd.n2956 vdd.n585 185
R17511 vdd.n2958 vdd.n2957 185
R17512 vdd.n2960 vdd.n583 185
R17513 vdd.n2962 vdd.n2961 185
R17514 vdd.n2963 vdd.n582 185
R17515 vdd.n2965 vdd.n2964 185
R17516 vdd.n2967 vdd.n580 185
R17517 vdd.n2969 vdd.n2968 185
R17518 vdd.n2970 vdd.n579 185
R17519 vdd.n2972 vdd.n2971 185
R17520 vdd.n2974 vdd.n578 185
R17521 vdd.n2975 vdd.n576 185
R17522 vdd.n2978 vdd.n2977 185
R17523 vdd.n577 vdd.n575 185
R17524 vdd.n2834 vdd.n2833 185
R17525 vdd.n2836 vdd.n2835 185
R17526 vdd.n2838 vdd.n2830 185
R17527 vdd.n2840 vdd.n2839 185
R17528 vdd.n2841 vdd.n2829 185
R17529 vdd.n2843 vdd.n2842 185
R17530 vdd.n2845 vdd.n2827 185
R17531 vdd.n2847 vdd.n2846 185
R17532 vdd.n2848 vdd.n2826 185
R17533 vdd.n2850 vdd.n2849 185
R17534 vdd.n2852 vdd.n2824 185
R17535 vdd.n2854 vdd.n2853 185
R17536 vdd.n2855 vdd.n2823 185
R17537 vdd.n2857 vdd.n2856 185
R17538 vdd.n2859 vdd.n2822 185
R17539 vdd.n2861 vdd.n2860 185
R17540 vdd.n2860 vdd.n484 185
R17541 vdd.n2946 vdd.n592 185
R17542 vdd.n2946 vdd.n2945 185
R17543 vdd.n2563 vdd.n594 185
R17544 vdd.n595 vdd.n594 185
R17545 vdd.n2564 vdd.n628 185
R17546 vdd.n2875 vdd.n628 185
R17547 vdd.n2566 vdd.n2565 185
R17548 vdd.n2565 vdd.n636 185
R17549 vdd.n2567 vdd.n635 185
R17550 vdd.n2869 vdd.n635 185
R17551 vdd.n2569 vdd.n2568 185
R17552 vdd.n2568 vdd.n633 185
R17553 vdd.n2570 vdd.n643 185
R17554 vdd.n2818 vdd.n643 185
R17555 vdd.n2572 vdd.n2571 185
R17556 vdd.n2571 vdd.n641 185
R17557 vdd.n2573 vdd.n648 185
R17558 vdd.n2812 vdd.n648 185
R17559 vdd.n2575 vdd.n2574 185
R17560 vdd.n2574 vdd.n654 185
R17561 vdd.n2576 vdd.n653 185
R17562 vdd.n2806 vdd.n653 185
R17563 vdd.n2578 vdd.n2577 185
R17564 vdd.n2577 vdd.n660 185
R17565 vdd.n2579 vdd.n659 185
R17566 vdd.n2800 vdd.n659 185
R17567 vdd.n2581 vdd.n2580 185
R17568 vdd.n2580 vdd.n667 185
R17569 vdd.n2582 vdd.n666 185
R17570 vdd.n2794 vdd.n666 185
R17571 vdd.n2584 vdd.n2583 185
R17572 vdd.n2583 vdd.n664 185
R17573 vdd.n2585 vdd.n673 185
R17574 vdd.n2788 vdd.n673 185
R17575 vdd.n2587 vdd.n2586 185
R17576 vdd.n2586 vdd.n671 185
R17577 vdd.n2588 vdd.n679 185
R17578 vdd.n2782 vdd.n679 185
R17579 vdd.n2590 vdd.n2589 185
R17580 vdd.n2589 vdd.n677 185
R17581 vdd.n2591 vdd.n684 185
R17582 vdd.n2776 vdd.n684 185
R17583 vdd.n2593 vdd.n2592 185
R17584 vdd.n2592 vdd.n691 185
R17585 vdd.n2594 vdd.n690 185
R17586 vdd.n2770 vdd.n690 185
R17587 vdd.n2596 vdd.n2595 185
R17588 vdd.n2595 vdd.n698 185
R17589 vdd.n2597 vdd.n697 185
R17590 vdd.n2764 vdd.n697 185
R17591 vdd.n2599 vdd.n2598 185
R17592 vdd.n2598 vdd.n695 185
R17593 vdd.n2600 vdd.n704 185
R17594 vdd.n2757 vdd.n704 185
R17595 vdd.n2602 vdd.n2601 185
R17596 vdd.n2601 vdd.n702 185
R17597 vdd.n2603 vdd.n709 185
R17598 vdd.n2751 vdd.n709 185
R17599 vdd.n2605 vdd.n2604 185
R17600 vdd.n2604 vdd.n715 185
R17601 vdd.n2606 vdd.n714 185
R17602 vdd.n2745 vdd.n714 185
R17603 vdd.n2608 vdd.n2607 185
R17604 vdd.n2607 vdd.n721 185
R17605 vdd.n2609 vdd.n720 185
R17606 vdd.n2739 vdd.n720 185
R17607 vdd.n2611 vdd.n2610 185
R17608 vdd.n2612 vdd.n2611 185
R17609 vdd.n2512 vdd.n726 185
R17610 vdd.n2733 vdd.n726 185
R17611 vdd.n2620 vdd.n2619 185
R17612 vdd.n2619 vdd.n2618 185
R17613 vdd.n2621 vdd.n732 185
R17614 vdd.n2727 vdd.n732 185
R17615 vdd.n2623 vdd.n2622 185
R17616 vdd.n2622 vdd.n730 185
R17617 vdd.n2624 vdd.n738 185
R17618 vdd.n2721 vdd.n738 185
R17619 vdd.n2626 vdd.n2625 185
R17620 vdd.n2625 vdd.n736 185
R17621 vdd.n2627 vdd.n743 185
R17622 vdd.n2715 vdd.n743 185
R17623 vdd.n2629 vdd.n2628 185
R17624 vdd.n2630 vdd.n2629 185
R17625 vdd.n2511 vdd.n749 185
R17626 vdd.n2709 vdd.n749 185
R17627 vdd.n2510 vdd.n2509 185
R17628 vdd.n2509 vdd.n747 185
R17629 vdd.n1971 vdd.n1970 185
R17630 vdd.n1972 vdd.n1971 185
R17631 vdd.n1321 vdd.n1319 185
R17632 vdd.n1963 vdd.n1319 185
R17633 vdd.n1966 vdd.n1965 185
R17634 vdd.n1965 vdd.n1964 185
R17635 vdd.n1324 vdd.n1323 185
R17636 vdd.n1325 vdd.n1324 185
R17637 vdd.n1952 vdd.n1951 185
R17638 vdd.n1953 vdd.n1952 185
R17639 vdd.n1333 vdd.n1332 185
R17640 vdd.n1944 vdd.n1332 185
R17641 vdd.n1947 vdd.n1946 185
R17642 vdd.n1946 vdd.n1945 185
R17643 vdd.n1336 vdd.n1335 185
R17644 vdd.n1343 vdd.n1336 185
R17645 vdd.n1935 vdd.n1934 185
R17646 vdd.n1936 vdd.n1935 185
R17647 vdd.n1345 vdd.n1344 185
R17648 vdd.n1344 vdd.n1342 185
R17649 vdd.n1930 vdd.n1929 185
R17650 vdd.n1929 vdd.n1928 185
R17651 vdd.n1618 vdd.n1617 185
R17652 vdd.n1619 vdd.n1618 185
R17653 vdd.n1919 vdd.n1918 185
R17654 vdd.n1920 vdd.n1919 185
R17655 vdd.n1626 vdd.n1625 185
R17656 vdd.n1910 vdd.n1625 185
R17657 vdd.n1913 vdd.n1912 185
R17658 vdd.n1912 vdd.n1911 185
R17659 vdd.n1629 vdd.n1628 185
R17660 vdd.n1635 vdd.n1629 185
R17661 vdd.n1901 vdd.n1900 185
R17662 vdd.n1902 vdd.n1901 185
R17663 vdd.n1637 vdd.n1636 185
R17664 vdd.n1893 vdd.n1636 185
R17665 vdd.n1896 vdd.n1895 185
R17666 vdd.n1895 vdd.n1894 185
R17667 vdd.n1640 vdd.n1639 185
R17668 vdd.n1641 vdd.n1640 185
R17669 vdd.n1884 vdd.n1883 185
R17670 vdd.n1885 vdd.n1884 185
R17671 vdd.n1648 vdd.n1647 185
R17672 vdd.n1683 vdd.n1647 185
R17673 vdd.n1879 vdd.n1878 185
R17674 vdd.n1651 vdd.n1650 185
R17675 vdd.n1875 vdd.n1874 185
R17676 vdd.n1876 vdd.n1875 185
R17677 vdd.n1685 vdd.n1684 185
R17678 vdd.n1870 vdd.n1687 185
R17679 vdd.n1869 vdd.n1688 185
R17680 vdd.n1868 vdd.n1689 185
R17681 vdd.n1691 vdd.n1690 185
R17682 vdd.n1864 vdd.n1693 185
R17683 vdd.n1863 vdd.n1694 185
R17684 vdd.n1862 vdd.n1695 185
R17685 vdd.n1697 vdd.n1696 185
R17686 vdd.n1858 vdd.n1699 185
R17687 vdd.n1857 vdd.n1700 185
R17688 vdd.n1856 vdd.n1701 185
R17689 vdd.n1703 vdd.n1702 185
R17690 vdd.n1852 vdd.n1705 185
R17691 vdd.n1851 vdd.n1706 185
R17692 vdd.n1850 vdd.n1707 185
R17693 vdd.n1711 vdd.n1708 185
R17694 vdd.n1846 vdd.n1713 185
R17695 vdd.n1845 vdd.n1714 185
R17696 vdd.n1844 vdd.n1715 185
R17697 vdd.n1717 vdd.n1716 185
R17698 vdd.n1840 vdd.n1719 185
R17699 vdd.n1839 vdd.n1720 185
R17700 vdd.n1838 vdd.n1721 185
R17701 vdd.n1723 vdd.n1722 185
R17702 vdd.n1834 vdd.n1725 185
R17703 vdd.n1833 vdd.n1726 185
R17704 vdd.n1832 vdd.n1727 185
R17705 vdd.n1729 vdd.n1728 185
R17706 vdd.n1828 vdd.n1731 185
R17707 vdd.n1827 vdd.n1732 185
R17708 vdd.n1826 vdd.n1733 185
R17709 vdd.n1735 vdd.n1734 185
R17710 vdd.n1822 vdd.n1737 185
R17711 vdd.n1821 vdd.n1738 185
R17712 vdd.n1820 vdd.n1739 185
R17713 vdd.n1741 vdd.n1740 185
R17714 vdd.n1816 vdd.n1743 185
R17715 vdd.n1815 vdd.n1812 185
R17716 vdd.n1811 vdd.n1744 185
R17717 vdd.n1746 vdd.n1745 185
R17718 vdd.n1807 vdd.n1748 185
R17719 vdd.n1806 vdd.n1749 185
R17720 vdd.n1805 vdd.n1750 185
R17721 vdd.n1752 vdd.n1751 185
R17722 vdd.n1801 vdd.n1754 185
R17723 vdd.n1800 vdd.n1755 185
R17724 vdd.n1799 vdd.n1756 185
R17725 vdd.n1758 vdd.n1757 185
R17726 vdd.n1795 vdd.n1760 185
R17727 vdd.n1794 vdd.n1761 185
R17728 vdd.n1793 vdd.n1762 185
R17729 vdd.n1764 vdd.n1763 185
R17730 vdd.n1789 vdd.n1766 185
R17731 vdd.n1788 vdd.n1767 185
R17732 vdd.n1787 vdd.n1768 185
R17733 vdd.n1770 vdd.n1769 185
R17734 vdd.n1783 vdd.n1772 185
R17735 vdd.n1782 vdd.n1773 185
R17736 vdd.n1781 vdd.n1774 185
R17737 vdd.n1778 vdd.n1682 185
R17738 vdd.n1876 vdd.n1682 185
R17739 vdd.n1975 vdd.n1974 185
R17740 vdd.n1979 vdd.n1315 185
R17741 vdd.n1314 vdd.n1308 185
R17742 vdd.n1312 vdd.n1311 185
R17743 vdd.n1310 vdd.n1069 185
R17744 vdd.n1983 vdd.n1066 185
R17745 vdd.n1985 vdd.n1984 185
R17746 vdd.n1987 vdd.n1064 185
R17747 vdd.n1989 vdd.n1988 185
R17748 vdd.n1990 vdd.n1059 185
R17749 vdd.n1992 vdd.n1991 185
R17750 vdd.n1994 vdd.n1057 185
R17751 vdd.n1996 vdd.n1995 185
R17752 vdd.n1997 vdd.n1052 185
R17753 vdd.n1999 vdd.n1998 185
R17754 vdd.n2001 vdd.n1050 185
R17755 vdd.n2003 vdd.n2002 185
R17756 vdd.n2004 vdd.n1046 185
R17757 vdd.n2006 vdd.n2005 185
R17758 vdd.n2008 vdd.n1043 185
R17759 vdd.n2010 vdd.n2009 185
R17760 vdd.n1044 vdd.n1037 185
R17761 vdd.n2014 vdd.n1041 185
R17762 vdd.n2015 vdd.n1033 185
R17763 vdd.n2017 vdd.n2016 185
R17764 vdd.n2019 vdd.n1031 185
R17765 vdd.n2021 vdd.n2020 185
R17766 vdd.n2022 vdd.n1026 185
R17767 vdd.n2024 vdd.n2023 185
R17768 vdd.n2026 vdd.n1024 185
R17769 vdd.n2028 vdd.n2027 185
R17770 vdd.n2029 vdd.n1019 185
R17771 vdd.n2031 vdd.n2030 185
R17772 vdd.n2033 vdd.n1017 185
R17773 vdd.n2035 vdd.n2034 185
R17774 vdd.n2036 vdd.n1012 185
R17775 vdd.n2038 vdd.n2037 185
R17776 vdd.n2040 vdd.n1010 185
R17777 vdd.n2042 vdd.n2041 185
R17778 vdd.n2043 vdd.n1006 185
R17779 vdd.n2045 vdd.n2044 185
R17780 vdd.n2047 vdd.n1003 185
R17781 vdd.n2049 vdd.n2048 185
R17782 vdd.n1004 vdd.n997 185
R17783 vdd.n2053 vdd.n1001 185
R17784 vdd.n2054 vdd.n993 185
R17785 vdd.n2056 vdd.n2055 185
R17786 vdd.n2058 vdd.n991 185
R17787 vdd.n2060 vdd.n2059 185
R17788 vdd.n2061 vdd.n986 185
R17789 vdd.n2063 vdd.n2062 185
R17790 vdd.n2065 vdd.n984 185
R17791 vdd.n2067 vdd.n2066 185
R17792 vdd.n2068 vdd.n979 185
R17793 vdd.n2070 vdd.n2069 185
R17794 vdd.n2072 vdd.n977 185
R17795 vdd.n2074 vdd.n2073 185
R17796 vdd.n2075 vdd.n975 185
R17797 vdd.n2077 vdd.n2076 185
R17798 vdd.n2080 vdd.n2079 185
R17799 vdd.n2082 vdd.n2081 185
R17800 vdd.n2084 vdd.n973 185
R17801 vdd.n2086 vdd.n2085 185
R17802 vdd.n1320 vdd.n972 185
R17803 vdd.n1973 vdd.n1318 185
R17804 vdd.n1973 vdd.n1972 185
R17805 vdd.n1328 vdd.n1317 185
R17806 vdd.n1963 vdd.n1317 185
R17807 vdd.n1962 vdd.n1961 185
R17808 vdd.n1964 vdd.n1962 185
R17809 vdd.n1327 vdd.n1326 185
R17810 vdd.n1326 vdd.n1325 185
R17811 vdd.n1955 vdd.n1954 185
R17812 vdd.n1954 vdd.n1953 185
R17813 vdd.n1331 vdd.n1330 185
R17814 vdd.n1944 vdd.n1331 185
R17815 vdd.n1943 vdd.n1942 185
R17816 vdd.n1945 vdd.n1943 185
R17817 vdd.n1338 vdd.n1337 185
R17818 vdd.n1343 vdd.n1337 185
R17819 vdd.n1938 vdd.n1937 185
R17820 vdd.n1937 vdd.n1936 185
R17821 vdd.n1341 vdd.n1340 185
R17822 vdd.n1342 vdd.n1341 185
R17823 vdd.n1927 vdd.n1926 185
R17824 vdd.n1928 vdd.n1927 185
R17825 vdd.n1621 vdd.n1620 185
R17826 vdd.n1620 vdd.n1619 185
R17827 vdd.n1922 vdd.n1921 185
R17828 vdd.n1921 vdd.n1920 185
R17829 vdd.n1624 vdd.n1623 185
R17830 vdd.n1910 vdd.n1624 185
R17831 vdd.n1909 vdd.n1908 185
R17832 vdd.n1911 vdd.n1909 185
R17833 vdd.n1631 vdd.n1630 185
R17834 vdd.n1635 vdd.n1630 185
R17835 vdd.n1904 vdd.n1903 185
R17836 vdd.n1903 vdd.n1902 185
R17837 vdd.n1634 vdd.n1633 185
R17838 vdd.n1893 vdd.n1634 185
R17839 vdd.n1892 vdd.n1891 185
R17840 vdd.n1894 vdd.n1892 185
R17841 vdd.n1643 vdd.n1642 185
R17842 vdd.n1642 vdd.n1641 185
R17843 vdd.n1887 vdd.n1886 185
R17844 vdd.n1886 vdd.n1885 185
R17845 vdd.n1646 vdd.n1645 185
R17846 vdd.n1683 vdd.n1646 185
R17847 vdd.n790 vdd.n788 185
R17848 vdd.n2326 vdd.n788 185
R17849 vdd.n2248 vdd.n808 185
R17850 vdd.n808 vdd.n795 185
R17851 vdd.n2250 vdd.n2249 185
R17852 vdd.n2251 vdd.n2250 185
R17853 vdd.n2247 vdd.n807 185
R17854 vdd.n1189 vdd.n807 185
R17855 vdd.n2246 vdd.n2245 185
R17856 vdd.n2245 vdd.n2244 185
R17857 vdd.n810 vdd.n809 185
R17858 vdd.n811 vdd.n810 185
R17859 vdd.n2235 vdd.n2234 185
R17860 vdd.n2236 vdd.n2235 185
R17861 vdd.n2233 vdd.n821 185
R17862 vdd.n821 vdd.n818 185
R17863 vdd.n2232 vdd.n2231 185
R17864 vdd.n2231 vdd.n2230 185
R17865 vdd.n823 vdd.n822 185
R17866 vdd.n1215 vdd.n823 185
R17867 vdd.n2223 vdd.n2222 185
R17868 vdd.n2224 vdd.n2223 185
R17869 vdd.n2221 vdd.n831 185
R17870 vdd.n836 vdd.n831 185
R17871 vdd.n2220 vdd.n2219 185
R17872 vdd.n2219 vdd.n2218 185
R17873 vdd.n833 vdd.n832 185
R17874 vdd.n842 vdd.n833 185
R17875 vdd.n2211 vdd.n2210 185
R17876 vdd.n2212 vdd.n2211 185
R17877 vdd.n2209 vdd.n843 185
R17878 vdd.n1227 vdd.n843 185
R17879 vdd.n2208 vdd.n2207 185
R17880 vdd.n2207 vdd.n2206 185
R17881 vdd.n845 vdd.n844 185
R17882 vdd.n846 vdd.n845 185
R17883 vdd.n2199 vdd.n2198 185
R17884 vdd.n2200 vdd.n2199 185
R17885 vdd.n2197 vdd.n855 185
R17886 vdd.n855 vdd.n852 185
R17887 vdd.n2196 vdd.n2195 185
R17888 vdd.n2195 vdd.n2194 185
R17889 vdd.n857 vdd.n856 185
R17890 vdd.n866 vdd.n857 185
R17891 vdd.n2186 vdd.n2185 185
R17892 vdd.n2187 vdd.n2186 185
R17893 vdd.n2184 vdd.n867 185
R17894 vdd.n873 vdd.n867 185
R17895 vdd.n2183 vdd.n2182 185
R17896 vdd.n2182 vdd.n2181 185
R17897 vdd.n869 vdd.n868 185
R17898 vdd.n870 vdd.n869 185
R17899 vdd.n2174 vdd.n2173 185
R17900 vdd.n2175 vdd.n2174 185
R17901 vdd.n2172 vdd.n880 185
R17902 vdd.n880 vdd.n877 185
R17903 vdd.n2171 vdd.n2170 185
R17904 vdd.n2170 vdd.n2169 185
R17905 vdd.n882 vdd.n881 185
R17906 vdd.n883 vdd.n882 185
R17907 vdd.n2162 vdd.n2161 185
R17908 vdd.n2163 vdd.n2162 185
R17909 vdd.n2160 vdd.n891 185
R17910 vdd.n896 vdd.n891 185
R17911 vdd.n2159 vdd.n2158 185
R17912 vdd.n2158 vdd.n2157 185
R17913 vdd.n893 vdd.n892 185
R17914 vdd.n902 vdd.n893 185
R17915 vdd.n2150 vdd.n2149 185
R17916 vdd.n2151 vdd.n2150 185
R17917 vdd.n2148 vdd.n903 185
R17918 vdd.n909 vdd.n903 185
R17919 vdd.n2147 vdd.n2146 185
R17920 vdd.n2146 vdd.n2145 185
R17921 vdd.n905 vdd.n904 185
R17922 vdd.n906 vdd.n905 185
R17923 vdd.n2138 vdd.n2137 185
R17924 vdd.n2139 vdd.n2138 185
R17925 vdd.n2136 vdd.n916 185
R17926 vdd.n916 vdd.n913 185
R17927 vdd.n2135 vdd.n2134 185
R17928 vdd.n2134 vdd.n2133 185
R17929 vdd.n918 vdd.n917 185
R17930 vdd.n927 vdd.n918 185
R17931 vdd.n2126 vdd.n2125 185
R17932 vdd.n2127 vdd.n2126 185
R17933 vdd.n2124 vdd.n928 185
R17934 vdd.n928 vdd.n924 185
R17935 vdd.n2123 vdd.n2122 185
R17936 vdd.n930 vdd.n929 185
R17937 vdd.n2119 vdd.n2118 185
R17938 vdd.n2120 vdd.n2119 185
R17939 vdd.n2117 vdd.n966 185
R17940 vdd.n2116 vdd.n2115 185
R17941 vdd.n2114 vdd.n2113 185
R17942 vdd.n2112 vdd.n2111 185
R17943 vdd.n2110 vdd.n2109 185
R17944 vdd.n2108 vdd.n2107 185
R17945 vdd.n2106 vdd.n2105 185
R17946 vdd.n2104 vdd.n2103 185
R17947 vdd.n2102 vdd.n2101 185
R17948 vdd.n2100 vdd.n2099 185
R17949 vdd.n2098 vdd.n2097 185
R17950 vdd.n2096 vdd.n2095 185
R17951 vdd.n2094 vdd.n2093 185
R17952 vdd.n2092 vdd.n2091 185
R17953 vdd.n2090 vdd.n2089 185
R17954 vdd.n1111 vdd.n967 185
R17955 vdd.n1113 vdd.n1112 185
R17956 vdd.n1115 vdd.n1114 185
R17957 vdd.n1117 vdd.n1116 185
R17958 vdd.n1119 vdd.n1118 185
R17959 vdd.n1121 vdd.n1120 185
R17960 vdd.n1123 vdd.n1122 185
R17961 vdd.n1125 vdd.n1124 185
R17962 vdd.n1127 vdd.n1126 185
R17963 vdd.n1129 vdd.n1128 185
R17964 vdd.n1131 vdd.n1130 185
R17965 vdd.n1133 vdd.n1132 185
R17966 vdd.n1135 vdd.n1134 185
R17967 vdd.n1137 vdd.n1136 185
R17968 vdd.n1140 vdd.n1139 185
R17969 vdd.n1142 vdd.n1141 185
R17970 vdd.n1144 vdd.n1143 185
R17971 vdd.n2329 vdd.n2328 185
R17972 vdd.n2331 vdd.n2330 185
R17973 vdd.n2333 vdd.n2332 185
R17974 vdd.n2336 vdd.n2335 185
R17975 vdd.n2338 vdd.n2337 185
R17976 vdd.n2340 vdd.n2339 185
R17977 vdd.n2342 vdd.n2341 185
R17978 vdd.n2344 vdd.n2343 185
R17979 vdd.n2346 vdd.n2345 185
R17980 vdd.n2348 vdd.n2347 185
R17981 vdd.n2350 vdd.n2349 185
R17982 vdd.n2352 vdd.n2351 185
R17983 vdd.n2354 vdd.n2353 185
R17984 vdd.n2356 vdd.n2355 185
R17985 vdd.n2358 vdd.n2357 185
R17986 vdd.n2360 vdd.n2359 185
R17987 vdd.n2362 vdd.n2361 185
R17988 vdd.n2364 vdd.n2363 185
R17989 vdd.n2366 vdd.n2365 185
R17990 vdd.n2368 vdd.n2367 185
R17991 vdd.n2370 vdd.n2369 185
R17992 vdd.n2372 vdd.n2371 185
R17993 vdd.n2374 vdd.n2373 185
R17994 vdd.n2376 vdd.n2375 185
R17995 vdd.n2378 vdd.n2377 185
R17996 vdd.n2380 vdd.n2379 185
R17997 vdd.n2382 vdd.n2381 185
R17998 vdd.n2384 vdd.n2383 185
R17999 vdd.n2386 vdd.n2385 185
R18000 vdd.n2388 vdd.n2387 185
R18001 vdd.n2390 vdd.n2389 185
R18002 vdd.n2392 vdd.n2391 185
R18003 vdd.n2394 vdd.n2393 185
R18004 vdd.n2395 vdd.n789 185
R18005 vdd.n2397 vdd.n2396 185
R18006 vdd.n2398 vdd.n2397 185
R18007 vdd.n2327 vdd.n793 185
R18008 vdd.n2327 vdd.n2326 185
R18009 vdd.n1187 vdd.n794 185
R18010 vdd.n795 vdd.n794 185
R18011 vdd.n1188 vdd.n805 185
R18012 vdd.n2251 vdd.n805 185
R18013 vdd.n1191 vdd.n1190 185
R18014 vdd.n1190 vdd.n1189 185
R18015 vdd.n1192 vdd.n812 185
R18016 vdd.n2244 vdd.n812 185
R18017 vdd.n1194 vdd.n1193 185
R18018 vdd.n1193 vdd.n811 185
R18019 vdd.n1195 vdd.n819 185
R18020 vdd.n2236 vdd.n819 185
R18021 vdd.n1197 vdd.n1196 185
R18022 vdd.n1196 vdd.n818 185
R18023 vdd.n1198 vdd.n824 185
R18024 vdd.n2230 vdd.n824 185
R18025 vdd.n1217 vdd.n1216 185
R18026 vdd.n1216 vdd.n1215 185
R18027 vdd.n1218 vdd.n829 185
R18028 vdd.n2224 vdd.n829 185
R18029 vdd.n1220 vdd.n1219 185
R18030 vdd.n1219 vdd.n836 185
R18031 vdd.n1221 vdd.n834 185
R18032 vdd.n2218 vdd.n834 185
R18033 vdd.n1223 vdd.n1222 185
R18034 vdd.n1222 vdd.n842 185
R18035 vdd.n1224 vdd.n840 185
R18036 vdd.n2212 vdd.n840 185
R18037 vdd.n1226 vdd.n1225 185
R18038 vdd.n1227 vdd.n1226 185
R18039 vdd.n1186 vdd.n847 185
R18040 vdd.n2206 vdd.n847 185
R18041 vdd.n1185 vdd.n1184 185
R18042 vdd.n1184 vdd.n846 185
R18043 vdd.n1183 vdd.n853 185
R18044 vdd.n2200 vdd.n853 185
R18045 vdd.n1182 vdd.n1181 185
R18046 vdd.n1181 vdd.n852 185
R18047 vdd.n1180 vdd.n858 185
R18048 vdd.n2194 vdd.n858 185
R18049 vdd.n1179 vdd.n1178 185
R18050 vdd.n1178 vdd.n866 185
R18051 vdd.n1177 vdd.n864 185
R18052 vdd.n2187 vdd.n864 185
R18053 vdd.n1176 vdd.n1175 185
R18054 vdd.n1175 vdd.n873 185
R18055 vdd.n1174 vdd.n871 185
R18056 vdd.n2181 vdd.n871 185
R18057 vdd.n1173 vdd.n1172 185
R18058 vdd.n1172 vdd.n870 185
R18059 vdd.n1171 vdd.n878 185
R18060 vdd.n2175 vdd.n878 185
R18061 vdd.n1170 vdd.n1169 185
R18062 vdd.n1169 vdd.n877 185
R18063 vdd.n1168 vdd.n884 185
R18064 vdd.n2169 vdd.n884 185
R18065 vdd.n1167 vdd.n1166 185
R18066 vdd.n1166 vdd.n883 185
R18067 vdd.n1165 vdd.n889 185
R18068 vdd.n2163 vdd.n889 185
R18069 vdd.n1164 vdd.n1163 185
R18070 vdd.n1163 vdd.n896 185
R18071 vdd.n1162 vdd.n894 185
R18072 vdd.n2157 vdd.n894 185
R18073 vdd.n1161 vdd.n1160 185
R18074 vdd.n1160 vdd.n902 185
R18075 vdd.n1159 vdd.n900 185
R18076 vdd.n2151 vdd.n900 185
R18077 vdd.n1158 vdd.n1157 185
R18078 vdd.n1157 vdd.n909 185
R18079 vdd.n1156 vdd.n907 185
R18080 vdd.n2145 vdd.n907 185
R18081 vdd.n1155 vdd.n1154 185
R18082 vdd.n1154 vdd.n906 185
R18083 vdd.n1153 vdd.n914 185
R18084 vdd.n2139 vdd.n914 185
R18085 vdd.n1152 vdd.n1151 185
R18086 vdd.n1151 vdd.n913 185
R18087 vdd.n1150 vdd.n919 185
R18088 vdd.n2133 vdd.n919 185
R18089 vdd.n1149 vdd.n1148 185
R18090 vdd.n1148 vdd.n927 185
R18091 vdd.n1147 vdd.n925 185
R18092 vdd.n2127 vdd.n925 185
R18093 vdd.n1146 vdd.n1145 185
R18094 vdd.n1145 vdd.n924 185
R18095 vdd.n3296 vdd.n3295 185
R18096 vdd.n3297 vdd.n3296 185
R18097 vdd.n325 vdd.n324 185
R18098 vdd.n3298 vdd.n325 185
R18099 vdd.n3301 vdd.n3300 185
R18100 vdd.n3300 vdd.n3299 185
R18101 vdd.n3302 vdd.n319 185
R18102 vdd.n319 vdd.n318 185
R18103 vdd.n3304 vdd.n3303 185
R18104 vdd.n3305 vdd.n3304 185
R18105 vdd.n314 vdd.n313 185
R18106 vdd.n3306 vdd.n314 185
R18107 vdd.n3309 vdd.n3308 185
R18108 vdd.n3308 vdd.n3307 185
R18109 vdd.n3310 vdd.n309 185
R18110 vdd.n309 vdd.n308 185
R18111 vdd.n3312 vdd.n3311 185
R18112 vdd.n3313 vdd.n3312 185
R18113 vdd.n303 vdd.n301 185
R18114 vdd.n3314 vdd.n303 185
R18115 vdd.n3317 vdd.n3316 185
R18116 vdd.n3316 vdd.n3315 185
R18117 vdd.n302 vdd.n300 185
R18118 vdd.n304 vdd.n302 185
R18119 vdd.n3153 vdd.n3152 185
R18120 vdd.n3154 vdd.n3153 185
R18121 vdd.n458 vdd.n457 185
R18122 vdd.n457 vdd.n456 185
R18123 vdd.n3148 vdd.n3147 185
R18124 vdd.n3147 vdd.n3146 185
R18125 vdd.n461 vdd.n460 185
R18126 vdd.n467 vdd.n461 185
R18127 vdd.n3137 vdd.n3136 185
R18128 vdd.n3138 vdd.n3137 185
R18129 vdd.n469 vdd.n468 185
R18130 vdd.n3129 vdd.n468 185
R18131 vdd.n3132 vdd.n3131 185
R18132 vdd.n3131 vdd.n3130 185
R18133 vdd.n472 vdd.n471 185
R18134 vdd.n473 vdd.n472 185
R18135 vdd.n3120 vdd.n3119 185
R18136 vdd.n3121 vdd.n3120 185
R18137 vdd.n480 vdd.n479 185
R18138 vdd.n516 vdd.n479 185
R18139 vdd.n3115 vdd.n3114 185
R18140 vdd.n483 vdd.n482 185
R18141 vdd.n3111 vdd.n3110 185
R18142 vdd.n3112 vdd.n3111 185
R18143 vdd.n518 vdd.n517 185
R18144 vdd.n522 vdd.n521 185
R18145 vdd.n3106 vdd.n523 185
R18146 vdd.n3105 vdd.n3104 185
R18147 vdd.n3103 vdd.n3102 185
R18148 vdd.n3101 vdd.n3100 185
R18149 vdd.n3099 vdd.n3098 185
R18150 vdd.n3097 vdd.n3096 185
R18151 vdd.n3095 vdd.n3094 185
R18152 vdd.n3093 vdd.n3092 185
R18153 vdd.n3091 vdd.n3090 185
R18154 vdd.n3089 vdd.n3088 185
R18155 vdd.n3087 vdd.n3086 185
R18156 vdd.n3085 vdd.n3084 185
R18157 vdd.n3083 vdd.n3082 185
R18158 vdd.n3081 vdd.n3080 185
R18159 vdd.n3079 vdd.n3078 185
R18160 vdd.n3070 vdd.n536 185
R18161 vdd.n3072 vdd.n3071 185
R18162 vdd.n3069 vdd.n3068 185
R18163 vdd.n3067 vdd.n3066 185
R18164 vdd.n3065 vdd.n3064 185
R18165 vdd.n3063 vdd.n3062 185
R18166 vdd.n3061 vdd.n3060 185
R18167 vdd.n3059 vdd.n3058 185
R18168 vdd.n3057 vdd.n3056 185
R18169 vdd.n3055 vdd.n3054 185
R18170 vdd.n3053 vdd.n3052 185
R18171 vdd.n3051 vdd.n3050 185
R18172 vdd.n3049 vdd.n3048 185
R18173 vdd.n3047 vdd.n3046 185
R18174 vdd.n3045 vdd.n3044 185
R18175 vdd.n3043 vdd.n3042 185
R18176 vdd.n3041 vdd.n3040 185
R18177 vdd.n3039 vdd.n3038 185
R18178 vdd.n3037 vdd.n3036 185
R18179 vdd.n3035 vdd.n3034 185
R18180 vdd.n3033 vdd.n3032 185
R18181 vdd.n3031 vdd.n3030 185
R18182 vdd.n3024 vdd.n556 185
R18183 vdd.n3026 vdd.n3025 185
R18184 vdd.n3023 vdd.n3022 185
R18185 vdd.n3021 vdd.n3020 185
R18186 vdd.n3019 vdd.n3018 185
R18187 vdd.n3017 vdd.n3016 185
R18188 vdd.n3015 vdd.n3014 185
R18189 vdd.n3013 vdd.n3012 185
R18190 vdd.n3011 vdd.n3010 185
R18191 vdd.n3009 vdd.n3008 185
R18192 vdd.n3007 vdd.n3006 185
R18193 vdd.n3005 vdd.n3004 185
R18194 vdd.n3003 vdd.n3002 185
R18195 vdd.n3001 vdd.n3000 185
R18196 vdd.n2999 vdd.n2998 185
R18197 vdd.n2997 vdd.n2996 185
R18198 vdd.n2995 vdd.n2994 185
R18199 vdd.n2993 vdd.n2992 185
R18200 vdd.n2991 vdd.n2990 185
R18201 vdd.n2989 vdd.n2988 185
R18202 vdd.n2987 vdd.n2986 185
R18203 vdd.n2982 vdd.n515 185
R18204 vdd.n3112 vdd.n515 185
R18205 vdd.n3179 vdd.n3178 185
R18206 vdd.n3183 vdd.n440 185
R18207 vdd.n3185 vdd.n3184 185
R18208 vdd.n3187 vdd.n438 185
R18209 vdd.n3189 vdd.n3188 185
R18210 vdd.n3190 vdd.n433 185
R18211 vdd.n3192 vdd.n3191 185
R18212 vdd.n3194 vdd.n431 185
R18213 vdd.n3196 vdd.n3195 185
R18214 vdd.n3197 vdd.n426 185
R18215 vdd.n3199 vdd.n3198 185
R18216 vdd.n3201 vdd.n424 185
R18217 vdd.n3203 vdd.n3202 185
R18218 vdd.n3204 vdd.n419 185
R18219 vdd.n3206 vdd.n3205 185
R18220 vdd.n3208 vdd.n417 185
R18221 vdd.n3210 vdd.n3209 185
R18222 vdd.n3211 vdd.n413 185
R18223 vdd.n3213 vdd.n3212 185
R18224 vdd.n3215 vdd.n410 185
R18225 vdd.n3217 vdd.n3216 185
R18226 vdd.n411 vdd.n404 185
R18227 vdd.n3221 vdd.n408 185
R18228 vdd.n3222 vdd.n400 185
R18229 vdd.n3224 vdd.n3223 185
R18230 vdd.n3226 vdd.n398 185
R18231 vdd.n3228 vdd.n3227 185
R18232 vdd.n3229 vdd.n393 185
R18233 vdd.n3231 vdd.n3230 185
R18234 vdd.n3233 vdd.n391 185
R18235 vdd.n3235 vdd.n3234 185
R18236 vdd.n3236 vdd.n386 185
R18237 vdd.n3238 vdd.n3237 185
R18238 vdd.n3240 vdd.n384 185
R18239 vdd.n3242 vdd.n3241 185
R18240 vdd.n3243 vdd.n379 185
R18241 vdd.n3245 vdd.n3244 185
R18242 vdd.n3247 vdd.n377 185
R18243 vdd.n3249 vdd.n3248 185
R18244 vdd.n3250 vdd.n373 185
R18245 vdd.n3252 vdd.n3251 185
R18246 vdd.n3254 vdd.n370 185
R18247 vdd.n3256 vdd.n3255 185
R18248 vdd.n371 vdd.n364 185
R18249 vdd.n3260 vdd.n368 185
R18250 vdd.n3261 vdd.n360 185
R18251 vdd.n3263 vdd.n3262 185
R18252 vdd.n3265 vdd.n358 185
R18253 vdd.n3267 vdd.n3266 185
R18254 vdd.n3268 vdd.n353 185
R18255 vdd.n3270 vdd.n3269 185
R18256 vdd.n3272 vdd.n351 185
R18257 vdd.n3274 vdd.n3273 185
R18258 vdd.n3275 vdd.n346 185
R18259 vdd.n3277 vdd.n3276 185
R18260 vdd.n3279 vdd.n344 185
R18261 vdd.n3281 vdd.n3280 185
R18262 vdd.n3282 vdd.n338 185
R18263 vdd.n3284 vdd.n3283 185
R18264 vdd.n3286 vdd.n337 185
R18265 vdd.n3287 vdd.n336 185
R18266 vdd.n3290 vdd.n3289 185
R18267 vdd.n3291 vdd.n334 185
R18268 vdd.n3292 vdd.n330 185
R18269 vdd.n3174 vdd.n328 185
R18270 vdd.n3297 vdd.n328 185
R18271 vdd.n3173 vdd.n327 185
R18272 vdd.n3298 vdd.n327 185
R18273 vdd.n3172 vdd.n326 185
R18274 vdd.n3299 vdd.n326 185
R18275 vdd.n446 vdd.n445 185
R18276 vdd.n445 vdd.n318 185
R18277 vdd.n3168 vdd.n317 185
R18278 vdd.n3305 vdd.n317 185
R18279 vdd.n3167 vdd.n316 185
R18280 vdd.n3306 vdd.n316 185
R18281 vdd.n3166 vdd.n315 185
R18282 vdd.n3307 vdd.n315 185
R18283 vdd.n449 vdd.n448 185
R18284 vdd.n448 vdd.n308 185
R18285 vdd.n3162 vdd.n307 185
R18286 vdd.n3313 vdd.n307 185
R18287 vdd.n3161 vdd.n306 185
R18288 vdd.n3314 vdd.n306 185
R18289 vdd.n3160 vdd.n305 185
R18290 vdd.n3315 vdd.n305 185
R18291 vdd.n455 vdd.n451 185
R18292 vdd.n455 vdd.n304 185
R18293 vdd.n3156 vdd.n3155 185
R18294 vdd.n3155 vdd.n3154 185
R18295 vdd.n454 vdd.n453 185
R18296 vdd.n456 vdd.n454 185
R18297 vdd.n3145 vdd.n3144 185
R18298 vdd.n3146 vdd.n3145 185
R18299 vdd.n463 vdd.n462 185
R18300 vdd.n467 vdd.n462 185
R18301 vdd.n3140 vdd.n3139 185
R18302 vdd.n3139 vdd.n3138 185
R18303 vdd.n466 vdd.n465 185
R18304 vdd.n3129 vdd.n466 185
R18305 vdd.n3128 vdd.n3127 185
R18306 vdd.n3130 vdd.n3128 185
R18307 vdd.n475 vdd.n474 185
R18308 vdd.n474 vdd.n473 185
R18309 vdd.n3123 vdd.n3122 185
R18310 vdd.n3122 vdd.n3121 185
R18311 vdd.n478 vdd.n477 185
R18312 vdd.n516 vdd.n478 185
R18313 vdd.n2705 vdd.n2704 185
R18314 vdd.n752 vdd.n751 185
R18315 vdd.n2701 vdd.n2700 185
R18316 vdd.n2702 vdd.n2701 185
R18317 vdd.n2699 vdd.n2433 185
R18318 vdd.n2698 vdd.n2697 185
R18319 vdd.n2696 vdd.n2695 185
R18320 vdd.n2694 vdd.n2693 185
R18321 vdd.n2692 vdd.n2691 185
R18322 vdd.n2690 vdd.n2689 185
R18323 vdd.n2688 vdd.n2687 185
R18324 vdd.n2686 vdd.n2685 185
R18325 vdd.n2684 vdd.n2683 185
R18326 vdd.n2682 vdd.n2681 185
R18327 vdd.n2680 vdd.n2679 185
R18328 vdd.n2678 vdd.n2677 185
R18329 vdd.n2676 vdd.n2675 185
R18330 vdd.n2674 vdd.n2673 185
R18331 vdd.n2672 vdd.n2671 185
R18332 vdd.n2670 vdd.n2669 185
R18333 vdd.n2668 vdd.n2667 185
R18334 vdd.n2666 vdd.n2665 185
R18335 vdd.n2664 vdd.n2663 185
R18336 vdd.n2662 vdd.n2661 185
R18337 vdd.n2660 vdd.n2659 185
R18338 vdd.n2658 vdd.n2657 185
R18339 vdd.n2656 vdd.n2655 185
R18340 vdd.n2654 vdd.n2653 185
R18341 vdd.n2652 vdd.n2651 185
R18342 vdd.n2650 vdd.n2649 185
R18343 vdd.n2648 vdd.n2647 185
R18344 vdd.n2646 vdd.n2645 185
R18345 vdd.n2644 vdd.n2643 185
R18346 vdd.n2641 vdd.n2640 185
R18347 vdd.n2639 vdd.n2638 185
R18348 vdd.n2637 vdd.n2636 185
R18349 vdd.n2881 vdd.n2880 185
R18350 vdd.n2883 vdd.n624 185
R18351 vdd.n2885 vdd.n2884 185
R18352 vdd.n2887 vdd.n621 185
R18353 vdd.n2889 vdd.n2888 185
R18354 vdd.n2891 vdd.n619 185
R18355 vdd.n2893 vdd.n2892 185
R18356 vdd.n2894 vdd.n618 185
R18357 vdd.n2896 vdd.n2895 185
R18358 vdd.n2898 vdd.n616 185
R18359 vdd.n2900 vdd.n2899 185
R18360 vdd.n2901 vdd.n615 185
R18361 vdd.n2903 vdd.n2902 185
R18362 vdd.n2905 vdd.n613 185
R18363 vdd.n2907 vdd.n2906 185
R18364 vdd.n2908 vdd.n612 185
R18365 vdd.n2910 vdd.n2909 185
R18366 vdd.n2912 vdd.n520 185
R18367 vdd.n2914 vdd.n2913 185
R18368 vdd.n2916 vdd.n610 185
R18369 vdd.n2918 vdd.n2917 185
R18370 vdd.n2919 vdd.n609 185
R18371 vdd.n2921 vdd.n2920 185
R18372 vdd.n2923 vdd.n607 185
R18373 vdd.n2925 vdd.n2924 185
R18374 vdd.n2926 vdd.n606 185
R18375 vdd.n2928 vdd.n2927 185
R18376 vdd.n2930 vdd.n604 185
R18377 vdd.n2932 vdd.n2931 185
R18378 vdd.n2933 vdd.n603 185
R18379 vdd.n2935 vdd.n2934 185
R18380 vdd.n2937 vdd.n602 185
R18381 vdd.n2938 vdd.n601 185
R18382 vdd.n2941 vdd.n2940 185
R18383 vdd.n2942 vdd.n599 185
R18384 vdd.n599 vdd.n484 185
R18385 vdd.n2879 vdd.n596 185
R18386 vdd.n2945 vdd.n596 185
R18387 vdd.n2878 vdd.n2877 185
R18388 vdd.n2877 vdd.n595 185
R18389 vdd.n2876 vdd.n626 185
R18390 vdd.n2876 vdd.n2875 185
R18391 vdd.n2519 vdd.n627 185
R18392 vdd.n636 vdd.n627 185
R18393 vdd.n2520 vdd.n634 185
R18394 vdd.n2869 vdd.n634 185
R18395 vdd.n2522 vdd.n2521 185
R18396 vdd.n2521 vdd.n633 185
R18397 vdd.n2523 vdd.n642 185
R18398 vdd.n2818 vdd.n642 185
R18399 vdd.n2525 vdd.n2524 185
R18400 vdd.n2524 vdd.n641 185
R18401 vdd.n2526 vdd.n647 185
R18402 vdd.n2812 vdd.n647 185
R18403 vdd.n2528 vdd.n2527 185
R18404 vdd.n2527 vdd.n654 185
R18405 vdd.n2529 vdd.n652 185
R18406 vdd.n2806 vdd.n652 185
R18407 vdd.n2531 vdd.n2530 185
R18408 vdd.n2530 vdd.n660 185
R18409 vdd.n2532 vdd.n658 185
R18410 vdd.n2800 vdd.n658 185
R18411 vdd.n2534 vdd.n2533 185
R18412 vdd.n2533 vdd.n667 185
R18413 vdd.n2535 vdd.n665 185
R18414 vdd.n2794 vdd.n665 185
R18415 vdd.n2537 vdd.n2536 185
R18416 vdd.n2536 vdd.n664 185
R18417 vdd.n2538 vdd.n672 185
R18418 vdd.n2788 vdd.n672 185
R18419 vdd.n2540 vdd.n2539 185
R18420 vdd.n2539 vdd.n671 185
R18421 vdd.n2541 vdd.n678 185
R18422 vdd.n2782 vdd.n678 185
R18423 vdd.n2543 vdd.n2542 185
R18424 vdd.n2542 vdd.n677 185
R18425 vdd.n2544 vdd.n683 185
R18426 vdd.n2776 vdd.n683 185
R18427 vdd.n2546 vdd.n2545 185
R18428 vdd.n2545 vdd.n691 185
R18429 vdd.n2547 vdd.n689 185
R18430 vdd.n2770 vdd.n689 185
R18431 vdd.n2549 vdd.n2548 185
R18432 vdd.n2548 vdd.n698 185
R18433 vdd.n2550 vdd.n696 185
R18434 vdd.n2764 vdd.n696 185
R18435 vdd.n2552 vdd.n2551 185
R18436 vdd.n2551 vdd.n695 185
R18437 vdd.n2553 vdd.n703 185
R18438 vdd.n2757 vdd.n703 185
R18439 vdd.n2555 vdd.n2554 185
R18440 vdd.n2554 vdd.n702 185
R18441 vdd.n2556 vdd.n708 185
R18442 vdd.n2751 vdd.n708 185
R18443 vdd.n2558 vdd.n2557 185
R18444 vdd.n2557 vdd.n715 185
R18445 vdd.n2559 vdd.n713 185
R18446 vdd.n2745 vdd.n713 185
R18447 vdd.n2561 vdd.n2560 185
R18448 vdd.n2560 vdd.n721 185
R18449 vdd.n2562 vdd.n719 185
R18450 vdd.n2739 vdd.n719 185
R18451 vdd.n2614 vdd.n2613 185
R18452 vdd.n2613 vdd.n2612 185
R18453 vdd.n2615 vdd.n725 185
R18454 vdd.n2733 vdd.n725 185
R18455 vdd.n2617 vdd.n2616 185
R18456 vdd.n2618 vdd.n2617 185
R18457 vdd.n2518 vdd.n731 185
R18458 vdd.n2727 vdd.n731 185
R18459 vdd.n2517 vdd.n2516 185
R18460 vdd.n2516 vdd.n730 185
R18461 vdd.n2515 vdd.n737 185
R18462 vdd.n2721 vdd.n737 185
R18463 vdd.n2514 vdd.n2513 185
R18464 vdd.n2513 vdd.n736 185
R18465 vdd.n2436 vdd.n742 185
R18466 vdd.n2715 vdd.n742 185
R18467 vdd.n2632 vdd.n2631 185
R18468 vdd.n2631 vdd.n2630 185
R18469 vdd.n2633 vdd.n748 185
R18470 vdd.n2709 vdd.n748 185
R18471 vdd.n2635 vdd.n2634 185
R18472 vdd.n2635 vdd.n747 185
R18473 vdd.n2706 vdd.n750 185
R18474 vdd.n750 vdd.n747 185
R18475 vdd.n2708 vdd.n2707 185
R18476 vdd.n2709 vdd.n2708 185
R18477 vdd.n741 vdd.n740 185
R18478 vdd.n2630 vdd.n741 185
R18479 vdd.n2717 vdd.n2716 185
R18480 vdd.n2716 vdd.n2715 185
R18481 vdd.n2718 vdd.n739 185
R18482 vdd.n739 vdd.n736 185
R18483 vdd.n2720 vdd.n2719 185
R18484 vdd.n2721 vdd.n2720 185
R18485 vdd.n729 vdd.n728 185
R18486 vdd.n730 vdd.n729 185
R18487 vdd.n2729 vdd.n2728 185
R18488 vdd.n2728 vdd.n2727 185
R18489 vdd.n2730 vdd.n727 185
R18490 vdd.n2618 vdd.n727 185
R18491 vdd.n2732 vdd.n2731 185
R18492 vdd.n2733 vdd.n2732 185
R18493 vdd.n718 vdd.n717 185
R18494 vdd.n2612 vdd.n718 185
R18495 vdd.n2741 vdd.n2740 185
R18496 vdd.n2740 vdd.n2739 185
R18497 vdd.n2742 vdd.n716 185
R18498 vdd.n721 vdd.n716 185
R18499 vdd.n2744 vdd.n2743 185
R18500 vdd.n2745 vdd.n2744 185
R18501 vdd.n707 vdd.n706 185
R18502 vdd.n715 vdd.n707 185
R18503 vdd.n2753 vdd.n2752 185
R18504 vdd.n2752 vdd.n2751 185
R18505 vdd.n2754 vdd.n705 185
R18506 vdd.n705 vdd.n702 185
R18507 vdd.n2756 vdd.n2755 185
R18508 vdd.n2757 vdd.n2756 185
R18509 vdd.n694 vdd.n693 185
R18510 vdd.n695 vdd.n694 185
R18511 vdd.n2766 vdd.n2765 185
R18512 vdd.n2765 vdd.n2764 185
R18513 vdd.n2767 vdd.n692 185
R18514 vdd.n698 vdd.n692 185
R18515 vdd.n2769 vdd.n2768 185
R18516 vdd.n2770 vdd.n2769 185
R18517 vdd.n682 vdd.n681 185
R18518 vdd.n691 vdd.n682 185
R18519 vdd.n2778 vdd.n2777 185
R18520 vdd.n2777 vdd.n2776 185
R18521 vdd.n2779 vdd.n680 185
R18522 vdd.n680 vdd.n677 185
R18523 vdd.n2781 vdd.n2780 185
R18524 vdd.n2782 vdd.n2781 185
R18525 vdd.n670 vdd.n669 185
R18526 vdd.n671 vdd.n670 185
R18527 vdd.n2790 vdd.n2789 185
R18528 vdd.n2789 vdd.n2788 185
R18529 vdd.n2791 vdd.n668 185
R18530 vdd.n668 vdd.n664 185
R18531 vdd.n2793 vdd.n2792 185
R18532 vdd.n2794 vdd.n2793 185
R18533 vdd.n657 vdd.n656 185
R18534 vdd.n667 vdd.n657 185
R18535 vdd.n2802 vdd.n2801 185
R18536 vdd.n2801 vdd.n2800 185
R18537 vdd.n2803 vdd.n655 185
R18538 vdd.n660 vdd.n655 185
R18539 vdd.n2805 vdd.n2804 185
R18540 vdd.n2806 vdd.n2805 185
R18541 vdd.n646 vdd.n645 185
R18542 vdd.n654 vdd.n646 185
R18543 vdd.n2814 vdd.n2813 185
R18544 vdd.n2813 vdd.n2812 185
R18545 vdd.n2815 vdd.n644 185
R18546 vdd.n644 vdd.n641 185
R18547 vdd.n2817 vdd.n2816 185
R18548 vdd.n2818 vdd.n2817 185
R18549 vdd.n632 vdd.n631 185
R18550 vdd.n633 vdd.n632 185
R18551 vdd.n2871 vdd.n2870 185
R18552 vdd.n2870 vdd.n2869 185
R18553 vdd.n2872 vdd.n630 185
R18554 vdd.n636 vdd.n630 185
R18555 vdd.n2874 vdd.n2873 185
R18556 vdd.n2875 vdd.n2874 185
R18557 vdd.n600 vdd.n598 185
R18558 vdd.n598 vdd.n595 185
R18559 vdd.n2944 vdd.n2943 185
R18560 vdd.n2945 vdd.n2944 185
R18561 vdd.n2325 vdd.n2324 185
R18562 vdd.n2326 vdd.n2325 185
R18563 vdd.n799 vdd.n797 185
R18564 vdd.n797 vdd.n795 185
R18565 vdd.n2240 vdd.n806 185
R18566 vdd.n2251 vdd.n806 185
R18567 vdd.n2241 vdd.n815 185
R18568 vdd.n1189 vdd.n815 185
R18569 vdd.n2243 vdd.n2242 185
R18570 vdd.n2244 vdd.n2243 185
R18571 vdd.n2239 vdd.n814 185
R18572 vdd.n814 vdd.n811 185
R18573 vdd.n2238 vdd.n2237 185
R18574 vdd.n2237 vdd.n2236 185
R18575 vdd.n817 vdd.n816 185
R18576 vdd.n818 vdd.n817 185
R18577 vdd.n2229 vdd.n2228 185
R18578 vdd.n2230 vdd.n2229 185
R18579 vdd.n2227 vdd.n826 185
R18580 vdd.n1215 vdd.n826 185
R18581 vdd.n2226 vdd.n2225 185
R18582 vdd.n2225 vdd.n2224 185
R18583 vdd.n828 vdd.n827 185
R18584 vdd.n836 vdd.n828 185
R18585 vdd.n2217 vdd.n2216 185
R18586 vdd.n2218 vdd.n2217 185
R18587 vdd.n2215 vdd.n837 185
R18588 vdd.n842 vdd.n837 185
R18589 vdd.n2214 vdd.n2213 185
R18590 vdd.n2213 vdd.n2212 185
R18591 vdd.n839 vdd.n838 185
R18592 vdd.n1227 vdd.n839 185
R18593 vdd.n2205 vdd.n2204 185
R18594 vdd.n2206 vdd.n2205 185
R18595 vdd.n2203 vdd.n849 185
R18596 vdd.n849 vdd.n846 185
R18597 vdd.n2202 vdd.n2201 185
R18598 vdd.n2201 vdd.n2200 185
R18599 vdd.n851 vdd.n850 185
R18600 vdd.n852 vdd.n851 185
R18601 vdd.n2193 vdd.n2192 185
R18602 vdd.n2194 vdd.n2193 185
R18603 vdd.n2190 vdd.n860 185
R18604 vdd.n866 vdd.n860 185
R18605 vdd.n2189 vdd.n2188 185
R18606 vdd.n2188 vdd.n2187 185
R18607 vdd.n863 vdd.n862 185
R18608 vdd.n873 vdd.n863 185
R18609 vdd.n2180 vdd.n2179 185
R18610 vdd.n2181 vdd.n2180 185
R18611 vdd.n2178 vdd.n874 185
R18612 vdd.n874 vdd.n870 185
R18613 vdd.n2177 vdd.n2176 185
R18614 vdd.n2176 vdd.n2175 185
R18615 vdd.n876 vdd.n875 185
R18616 vdd.n877 vdd.n876 185
R18617 vdd.n2168 vdd.n2167 185
R18618 vdd.n2169 vdd.n2168 185
R18619 vdd.n2166 vdd.n886 185
R18620 vdd.n886 vdd.n883 185
R18621 vdd.n2165 vdd.n2164 185
R18622 vdd.n2164 vdd.n2163 185
R18623 vdd.n888 vdd.n887 185
R18624 vdd.n896 vdd.n888 185
R18625 vdd.n2156 vdd.n2155 185
R18626 vdd.n2157 vdd.n2156 185
R18627 vdd.n2154 vdd.n897 185
R18628 vdd.n902 vdd.n897 185
R18629 vdd.n2153 vdd.n2152 185
R18630 vdd.n2152 vdd.n2151 185
R18631 vdd.n899 vdd.n898 185
R18632 vdd.n909 vdd.n899 185
R18633 vdd.n2144 vdd.n2143 185
R18634 vdd.n2145 vdd.n2144 185
R18635 vdd.n2142 vdd.n910 185
R18636 vdd.n910 vdd.n906 185
R18637 vdd.n2141 vdd.n2140 185
R18638 vdd.n2140 vdd.n2139 185
R18639 vdd.n912 vdd.n911 185
R18640 vdd.n913 vdd.n912 185
R18641 vdd.n2132 vdd.n2131 185
R18642 vdd.n2133 vdd.n2132 185
R18643 vdd.n2130 vdd.n921 185
R18644 vdd.n927 vdd.n921 185
R18645 vdd.n2129 vdd.n2128 185
R18646 vdd.n2128 vdd.n2127 185
R18647 vdd.n923 vdd.n922 185
R18648 vdd.n924 vdd.n923 185
R18649 vdd.n2256 vdd.n770 185
R18650 vdd.n2398 vdd.n770 185
R18651 vdd.n2258 vdd.n2257 185
R18652 vdd.n2260 vdd.n2259 185
R18653 vdd.n2262 vdd.n2261 185
R18654 vdd.n2264 vdd.n2263 185
R18655 vdd.n2266 vdd.n2265 185
R18656 vdd.n2268 vdd.n2267 185
R18657 vdd.n2270 vdd.n2269 185
R18658 vdd.n2272 vdd.n2271 185
R18659 vdd.n2274 vdd.n2273 185
R18660 vdd.n2276 vdd.n2275 185
R18661 vdd.n2278 vdd.n2277 185
R18662 vdd.n2280 vdd.n2279 185
R18663 vdd.n2282 vdd.n2281 185
R18664 vdd.n2284 vdd.n2283 185
R18665 vdd.n2286 vdd.n2285 185
R18666 vdd.n2288 vdd.n2287 185
R18667 vdd.n2290 vdd.n2289 185
R18668 vdd.n2292 vdd.n2291 185
R18669 vdd.n2294 vdd.n2293 185
R18670 vdd.n2296 vdd.n2295 185
R18671 vdd.n2298 vdd.n2297 185
R18672 vdd.n2300 vdd.n2299 185
R18673 vdd.n2302 vdd.n2301 185
R18674 vdd.n2304 vdd.n2303 185
R18675 vdd.n2306 vdd.n2305 185
R18676 vdd.n2308 vdd.n2307 185
R18677 vdd.n2310 vdd.n2309 185
R18678 vdd.n2312 vdd.n2311 185
R18679 vdd.n2314 vdd.n2313 185
R18680 vdd.n2316 vdd.n2315 185
R18681 vdd.n2318 vdd.n2317 185
R18682 vdd.n2320 vdd.n2319 185
R18683 vdd.n2322 vdd.n2321 185
R18684 vdd.n2323 vdd.n798 185
R18685 vdd.n2255 vdd.n796 185
R18686 vdd.n2326 vdd.n796 185
R18687 vdd.n2254 vdd.n2253 185
R18688 vdd.n2253 vdd.n795 185
R18689 vdd.n2252 vdd.n803 185
R18690 vdd.n2252 vdd.n2251 185
R18691 vdd.n1205 vdd.n804 185
R18692 vdd.n1189 vdd.n804 185
R18693 vdd.n1206 vdd.n813 185
R18694 vdd.n2244 vdd.n813 185
R18695 vdd.n1208 vdd.n1207 185
R18696 vdd.n1207 vdd.n811 185
R18697 vdd.n1209 vdd.n820 185
R18698 vdd.n2236 vdd.n820 185
R18699 vdd.n1211 vdd.n1210 185
R18700 vdd.n1210 vdd.n818 185
R18701 vdd.n1212 vdd.n825 185
R18702 vdd.n2230 vdd.n825 185
R18703 vdd.n1214 vdd.n1213 185
R18704 vdd.n1215 vdd.n1214 185
R18705 vdd.n1204 vdd.n830 185
R18706 vdd.n2224 vdd.n830 185
R18707 vdd.n1203 vdd.n1202 185
R18708 vdd.n1202 vdd.n836 185
R18709 vdd.n1201 vdd.n835 185
R18710 vdd.n2218 vdd.n835 185
R18711 vdd.n1200 vdd.n1199 185
R18712 vdd.n1199 vdd.n842 185
R18713 vdd.n1108 vdd.n841 185
R18714 vdd.n2212 vdd.n841 185
R18715 vdd.n1229 vdd.n1228 185
R18716 vdd.n1228 vdd.n1227 185
R18717 vdd.n1230 vdd.n848 185
R18718 vdd.n2206 vdd.n848 185
R18719 vdd.n1232 vdd.n1231 185
R18720 vdd.n1231 vdd.n846 185
R18721 vdd.n1233 vdd.n854 185
R18722 vdd.n2200 vdd.n854 185
R18723 vdd.n1235 vdd.n1234 185
R18724 vdd.n1234 vdd.n852 185
R18725 vdd.n1236 vdd.n859 185
R18726 vdd.n2194 vdd.n859 185
R18727 vdd.n1238 vdd.n1237 185
R18728 vdd.n1237 vdd.n866 185
R18729 vdd.n1239 vdd.n865 185
R18730 vdd.n2187 vdd.n865 185
R18731 vdd.n1241 vdd.n1240 185
R18732 vdd.n1240 vdd.n873 185
R18733 vdd.n1242 vdd.n872 185
R18734 vdd.n2181 vdd.n872 185
R18735 vdd.n1244 vdd.n1243 185
R18736 vdd.n1243 vdd.n870 185
R18737 vdd.n1245 vdd.n879 185
R18738 vdd.n2175 vdd.n879 185
R18739 vdd.n1247 vdd.n1246 185
R18740 vdd.n1246 vdd.n877 185
R18741 vdd.n1248 vdd.n885 185
R18742 vdd.n2169 vdd.n885 185
R18743 vdd.n1250 vdd.n1249 185
R18744 vdd.n1249 vdd.n883 185
R18745 vdd.n1251 vdd.n890 185
R18746 vdd.n2163 vdd.n890 185
R18747 vdd.n1253 vdd.n1252 185
R18748 vdd.n1252 vdd.n896 185
R18749 vdd.n1254 vdd.n895 185
R18750 vdd.n2157 vdd.n895 185
R18751 vdd.n1256 vdd.n1255 185
R18752 vdd.n1255 vdd.n902 185
R18753 vdd.n1257 vdd.n901 185
R18754 vdd.n2151 vdd.n901 185
R18755 vdd.n1259 vdd.n1258 185
R18756 vdd.n1258 vdd.n909 185
R18757 vdd.n1260 vdd.n908 185
R18758 vdd.n2145 vdd.n908 185
R18759 vdd.n1262 vdd.n1261 185
R18760 vdd.n1261 vdd.n906 185
R18761 vdd.n1263 vdd.n915 185
R18762 vdd.n2139 vdd.n915 185
R18763 vdd.n1265 vdd.n1264 185
R18764 vdd.n1264 vdd.n913 185
R18765 vdd.n1266 vdd.n920 185
R18766 vdd.n2133 vdd.n920 185
R18767 vdd.n1268 vdd.n1267 185
R18768 vdd.n1267 vdd.n927 185
R18769 vdd.n1269 vdd.n926 185
R18770 vdd.n2127 vdd.n926 185
R18771 vdd.n1271 vdd.n1270 185
R18772 vdd.n1270 vdd.n924 185
R18773 vdd.n1071 vdd.n1070 185
R18774 vdd.n1073 vdd.n1072 185
R18775 vdd.n1075 vdd.n1074 185
R18776 vdd.n1077 vdd.n1076 185
R18777 vdd.n1079 vdd.n1078 185
R18778 vdd.n1081 vdd.n1080 185
R18779 vdd.n1083 vdd.n1082 185
R18780 vdd.n1085 vdd.n1084 185
R18781 vdd.n1087 vdd.n1086 185
R18782 vdd.n1089 vdd.n1088 185
R18783 vdd.n1091 vdd.n1090 185
R18784 vdd.n1093 vdd.n1092 185
R18785 vdd.n1095 vdd.n1094 185
R18786 vdd.n1097 vdd.n1096 185
R18787 vdd.n1099 vdd.n1098 185
R18788 vdd.n1101 vdd.n1100 185
R18789 vdd.n1103 vdd.n1102 185
R18790 vdd.n1305 vdd.n1104 185
R18791 vdd.n1304 vdd.n1303 185
R18792 vdd.n1302 vdd.n1301 185
R18793 vdd.n1300 vdd.n1299 185
R18794 vdd.n1298 vdd.n1297 185
R18795 vdd.n1296 vdd.n1295 185
R18796 vdd.n1294 vdd.n1293 185
R18797 vdd.n1292 vdd.n1291 185
R18798 vdd.n1290 vdd.n1289 185
R18799 vdd.n1288 vdd.n1287 185
R18800 vdd.n1286 vdd.n1285 185
R18801 vdd.n1284 vdd.n1283 185
R18802 vdd.n1282 vdd.n1281 185
R18803 vdd.n1280 vdd.n1279 185
R18804 vdd.n1278 vdd.n1277 185
R18805 vdd.n1276 vdd.n1275 185
R18806 vdd.n1274 vdd.n1273 185
R18807 vdd.n1272 vdd.n965 185
R18808 vdd.n2120 vdd.n965 185
R18809 vdd.n291 vdd.n290 171.744
R18810 vdd.n290 vdd.n289 171.744
R18811 vdd.n289 vdd.n258 171.744
R18812 vdd.n282 vdd.n258 171.744
R18813 vdd.n282 vdd.n281 171.744
R18814 vdd.n281 vdd.n263 171.744
R18815 vdd.n274 vdd.n263 171.744
R18816 vdd.n274 vdd.n273 171.744
R18817 vdd.n273 vdd.n267 171.744
R18818 vdd.n244 vdd.n243 171.744
R18819 vdd.n243 vdd.n242 171.744
R18820 vdd.n242 vdd.n211 171.744
R18821 vdd.n235 vdd.n211 171.744
R18822 vdd.n235 vdd.n234 171.744
R18823 vdd.n234 vdd.n216 171.744
R18824 vdd.n227 vdd.n216 171.744
R18825 vdd.n227 vdd.n226 171.744
R18826 vdd.n226 vdd.n220 171.744
R18827 vdd.n201 vdd.n200 171.744
R18828 vdd.n200 vdd.n199 171.744
R18829 vdd.n199 vdd.n168 171.744
R18830 vdd.n192 vdd.n168 171.744
R18831 vdd.n192 vdd.n191 171.744
R18832 vdd.n191 vdd.n173 171.744
R18833 vdd.n184 vdd.n173 171.744
R18834 vdd.n184 vdd.n183 171.744
R18835 vdd.n183 vdd.n177 171.744
R18836 vdd.n154 vdd.n153 171.744
R18837 vdd.n153 vdd.n152 171.744
R18838 vdd.n152 vdd.n121 171.744
R18839 vdd.n145 vdd.n121 171.744
R18840 vdd.n145 vdd.n144 171.744
R18841 vdd.n144 vdd.n126 171.744
R18842 vdd.n137 vdd.n126 171.744
R18843 vdd.n137 vdd.n136 171.744
R18844 vdd.n136 vdd.n130 171.744
R18845 vdd.n112 vdd.n111 171.744
R18846 vdd.n111 vdd.n110 171.744
R18847 vdd.n110 vdd.n79 171.744
R18848 vdd.n103 vdd.n79 171.744
R18849 vdd.n103 vdd.n102 171.744
R18850 vdd.n102 vdd.n84 171.744
R18851 vdd.n95 vdd.n84 171.744
R18852 vdd.n95 vdd.n94 171.744
R18853 vdd.n94 vdd.n88 171.744
R18854 vdd.n65 vdd.n64 171.744
R18855 vdd.n64 vdd.n63 171.744
R18856 vdd.n63 vdd.n32 171.744
R18857 vdd.n56 vdd.n32 171.744
R18858 vdd.n56 vdd.n55 171.744
R18859 vdd.n55 vdd.n37 171.744
R18860 vdd.n48 vdd.n37 171.744
R18861 vdd.n48 vdd.n47 171.744
R18862 vdd.n47 vdd.n41 171.744
R18863 vdd.n1561 vdd.n1560 171.744
R18864 vdd.n1560 vdd.n1559 171.744
R18865 vdd.n1559 vdd.n1528 171.744
R18866 vdd.n1552 vdd.n1528 171.744
R18867 vdd.n1552 vdd.n1551 171.744
R18868 vdd.n1551 vdd.n1533 171.744
R18869 vdd.n1544 vdd.n1533 171.744
R18870 vdd.n1544 vdd.n1543 171.744
R18871 vdd.n1543 vdd.n1537 171.744
R18872 vdd.n1608 vdd.n1607 171.744
R18873 vdd.n1607 vdd.n1606 171.744
R18874 vdd.n1606 vdd.n1575 171.744
R18875 vdd.n1599 vdd.n1575 171.744
R18876 vdd.n1599 vdd.n1598 171.744
R18877 vdd.n1598 vdd.n1580 171.744
R18878 vdd.n1591 vdd.n1580 171.744
R18879 vdd.n1591 vdd.n1590 171.744
R18880 vdd.n1590 vdd.n1584 171.744
R18881 vdd.n1471 vdd.n1470 171.744
R18882 vdd.n1470 vdd.n1469 171.744
R18883 vdd.n1469 vdd.n1438 171.744
R18884 vdd.n1462 vdd.n1438 171.744
R18885 vdd.n1462 vdd.n1461 171.744
R18886 vdd.n1461 vdd.n1443 171.744
R18887 vdd.n1454 vdd.n1443 171.744
R18888 vdd.n1454 vdd.n1453 171.744
R18889 vdd.n1453 vdd.n1447 171.744
R18890 vdd.n1518 vdd.n1517 171.744
R18891 vdd.n1517 vdd.n1516 171.744
R18892 vdd.n1516 vdd.n1485 171.744
R18893 vdd.n1509 vdd.n1485 171.744
R18894 vdd.n1509 vdd.n1508 171.744
R18895 vdd.n1508 vdd.n1490 171.744
R18896 vdd.n1501 vdd.n1490 171.744
R18897 vdd.n1501 vdd.n1500 171.744
R18898 vdd.n1500 vdd.n1494 171.744
R18899 vdd.n1382 vdd.n1381 171.744
R18900 vdd.n1381 vdd.n1380 171.744
R18901 vdd.n1380 vdd.n1349 171.744
R18902 vdd.n1373 vdd.n1349 171.744
R18903 vdd.n1373 vdd.n1372 171.744
R18904 vdd.n1372 vdd.n1354 171.744
R18905 vdd.n1365 vdd.n1354 171.744
R18906 vdd.n1365 vdd.n1364 171.744
R18907 vdd.n1364 vdd.n1358 171.744
R18908 vdd.n1429 vdd.n1428 171.744
R18909 vdd.n1428 vdd.n1427 171.744
R18910 vdd.n1427 vdd.n1396 171.744
R18911 vdd.n1420 vdd.n1396 171.744
R18912 vdd.n1420 vdd.n1419 171.744
R18913 vdd.n1419 vdd.n1401 171.744
R18914 vdd.n1412 vdd.n1401 171.744
R18915 vdd.n1412 vdd.n1411 171.744
R18916 vdd.n1411 vdd.n1405 171.744
R18917 vdd.n3289 vdd.n334 146.341
R18918 vdd.n3287 vdd.n3286 146.341
R18919 vdd.n3284 vdd.n338 146.341
R18920 vdd.n3280 vdd.n3279 146.341
R18921 vdd.n3277 vdd.n346 146.341
R18922 vdd.n3273 vdd.n3272 146.341
R18923 vdd.n3270 vdd.n353 146.341
R18924 vdd.n3266 vdd.n3265 146.341
R18925 vdd.n3263 vdd.n360 146.341
R18926 vdd.n371 vdd.n368 146.341
R18927 vdd.n3255 vdd.n3254 146.341
R18928 vdd.n3252 vdd.n373 146.341
R18929 vdd.n3248 vdd.n3247 146.341
R18930 vdd.n3245 vdd.n379 146.341
R18931 vdd.n3241 vdd.n3240 146.341
R18932 vdd.n3238 vdd.n386 146.341
R18933 vdd.n3234 vdd.n3233 146.341
R18934 vdd.n3231 vdd.n393 146.341
R18935 vdd.n3227 vdd.n3226 146.341
R18936 vdd.n3224 vdd.n400 146.341
R18937 vdd.n411 vdd.n408 146.341
R18938 vdd.n3216 vdd.n3215 146.341
R18939 vdd.n3213 vdd.n413 146.341
R18940 vdd.n3209 vdd.n3208 146.341
R18941 vdd.n3206 vdd.n419 146.341
R18942 vdd.n3202 vdd.n3201 146.341
R18943 vdd.n3199 vdd.n426 146.341
R18944 vdd.n3195 vdd.n3194 146.341
R18945 vdd.n3192 vdd.n433 146.341
R18946 vdd.n3188 vdd.n3187 146.341
R18947 vdd.n3185 vdd.n440 146.341
R18948 vdd.n3122 vdd.n478 146.341
R18949 vdd.n3122 vdd.n474 146.341
R18950 vdd.n3128 vdd.n474 146.341
R18951 vdd.n3128 vdd.n466 146.341
R18952 vdd.n3139 vdd.n466 146.341
R18953 vdd.n3139 vdd.n462 146.341
R18954 vdd.n3145 vdd.n462 146.341
R18955 vdd.n3145 vdd.n454 146.341
R18956 vdd.n3155 vdd.n454 146.341
R18957 vdd.n3155 vdd.n455 146.341
R18958 vdd.n455 vdd.n305 146.341
R18959 vdd.n306 vdd.n305 146.341
R18960 vdd.n307 vdd.n306 146.341
R18961 vdd.n448 vdd.n307 146.341
R18962 vdd.n448 vdd.n315 146.341
R18963 vdd.n316 vdd.n315 146.341
R18964 vdd.n317 vdd.n316 146.341
R18965 vdd.n445 vdd.n317 146.341
R18966 vdd.n445 vdd.n326 146.341
R18967 vdd.n327 vdd.n326 146.341
R18968 vdd.n328 vdd.n327 146.341
R18969 vdd.n3111 vdd.n483 146.341
R18970 vdd.n3111 vdd.n517 146.341
R18971 vdd.n523 vdd.n522 146.341
R18972 vdd.n3104 vdd.n3103 146.341
R18973 vdd.n3100 vdd.n3099 146.341
R18974 vdd.n3096 vdd.n3095 146.341
R18975 vdd.n3092 vdd.n3091 146.341
R18976 vdd.n3088 vdd.n3087 146.341
R18977 vdd.n3084 vdd.n3083 146.341
R18978 vdd.n3080 vdd.n3079 146.341
R18979 vdd.n3071 vdd.n3070 146.341
R18980 vdd.n3068 vdd.n3067 146.341
R18981 vdd.n3064 vdd.n3063 146.341
R18982 vdd.n3060 vdd.n3059 146.341
R18983 vdd.n3056 vdd.n3055 146.341
R18984 vdd.n3052 vdd.n3051 146.341
R18985 vdd.n3048 vdd.n3047 146.341
R18986 vdd.n3044 vdd.n3043 146.341
R18987 vdd.n3040 vdd.n3039 146.341
R18988 vdd.n3036 vdd.n3035 146.341
R18989 vdd.n3032 vdd.n3031 146.341
R18990 vdd.n3025 vdd.n3024 146.341
R18991 vdd.n3022 vdd.n3021 146.341
R18992 vdd.n3018 vdd.n3017 146.341
R18993 vdd.n3014 vdd.n3013 146.341
R18994 vdd.n3010 vdd.n3009 146.341
R18995 vdd.n3006 vdd.n3005 146.341
R18996 vdd.n3002 vdd.n3001 146.341
R18997 vdd.n2998 vdd.n2997 146.341
R18998 vdd.n2994 vdd.n2993 146.341
R18999 vdd.n2990 vdd.n2989 146.341
R19000 vdd.n2986 vdd.n515 146.341
R19001 vdd.n3120 vdd.n479 146.341
R19002 vdd.n3120 vdd.n472 146.341
R19003 vdd.n3131 vdd.n472 146.341
R19004 vdd.n3131 vdd.n468 146.341
R19005 vdd.n3137 vdd.n468 146.341
R19006 vdd.n3137 vdd.n461 146.341
R19007 vdd.n3147 vdd.n461 146.341
R19008 vdd.n3147 vdd.n457 146.341
R19009 vdd.n3153 vdd.n457 146.341
R19010 vdd.n3153 vdd.n302 146.341
R19011 vdd.n3316 vdd.n302 146.341
R19012 vdd.n3316 vdd.n303 146.341
R19013 vdd.n3312 vdd.n303 146.341
R19014 vdd.n3312 vdd.n309 146.341
R19015 vdd.n3308 vdd.n309 146.341
R19016 vdd.n3308 vdd.n314 146.341
R19017 vdd.n3304 vdd.n314 146.341
R19018 vdd.n3304 vdd.n319 146.341
R19019 vdd.n3300 vdd.n319 146.341
R19020 vdd.n3300 vdd.n325 146.341
R19021 vdd.n3296 vdd.n325 146.341
R19022 vdd.n2085 vdd.n2084 146.341
R19023 vdd.n2082 vdd.n2079 146.341
R19024 vdd.n2077 vdd.n975 146.341
R19025 vdd.n2073 vdd.n2072 146.341
R19026 vdd.n2070 vdd.n979 146.341
R19027 vdd.n2066 vdd.n2065 146.341
R19028 vdd.n2063 vdd.n986 146.341
R19029 vdd.n2059 vdd.n2058 146.341
R19030 vdd.n2056 vdd.n993 146.341
R19031 vdd.n1004 vdd.n1001 146.341
R19032 vdd.n2048 vdd.n2047 146.341
R19033 vdd.n2045 vdd.n1006 146.341
R19034 vdd.n2041 vdd.n2040 146.341
R19035 vdd.n2038 vdd.n1012 146.341
R19036 vdd.n2034 vdd.n2033 146.341
R19037 vdd.n2031 vdd.n1019 146.341
R19038 vdd.n2027 vdd.n2026 146.341
R19039 vdd.n2024 vdd.n1026 146.341
R19040 vdd.n2020 vdd.n2019 146.341
R19041 vdd.n2017 vdd.n1033 146.341
R19042 vdd.n1044 vdd.n1041 146.341
R19043 vdd.n2009 vdd.n2008 146.341
R19044 vdd.n2006 vdd.n1046 146.341
R19045 vdd.n2002 vdd.n2001 146.341
R19046 vdd.n1999 vdd.n1052 146.341
R19047 vdd.n1995 vdd.n1994 146.341
R19048 vdd.n1992 vdd.n1059 146.341
R19049 vdd.n1988 vdd.n1987 146.341
R19050 vdd.n1985 vdd.n1066 146.341
R19051 vdd.n1312 vdd.n1310 146.341
R19052 vdd.n1315 vdd.n1314 146.341
R19053 vdd.n1886 vdd.n1646 146.341
R19054 vdd.n1886 vdd.n1642 146.341
R19055 vdd.n1892 vdd.n1642 146.341
R19056 vdd.n1892 vdd.n1634 146.341
R19057 vdd.n1903 vdd.n1634 146.341
R19058 vdd.n1903 vdd.n1630 146.341
R19059 vdd.n1909 vdd.n1630 146.341
R19060 vdd.n1909 vdd.n1624 146.341
R19061 vdd.n1921 vdd.n1624 146.341
R19062 vdd.n1921 vdd.n1620 146.341
R19063 vdd.n1927 vdd.n1620 146.341
R19064 vdd.n1927 vdd.n1341 146.341
R19065 vdd.n1937 vdd.n1341 146.341
R19066 vdd.n1937 vdd.n1337 146.341
R19067 vdd.n1943 vdd.n1337 146.341
R19068 vdd.n1943 vdd.n1331 146.341
R19069 vdd.n1954 vdd.n1331 146.341
R19070 vdd.n1954 vdd.n1326 146.341
R19071 vdd.n1962 vdd.n1326 146.341
R19072 vdd.n1962 vdd.n1317 146.341
R19073 vdd.n1973 vdd.n1317 146.341
R19074 vdd.n1875 vdd.n1651 146.341
R19075 vdd.n1875 vdd.n1684 146.341
R19076 vdd.n1688 vdd.n1687 146.341
R19077 vdd.n1690 vdd.n1689 146.341
R19078 vdd.n1694 vdd.n1693 146.341
R19079 vdd.n1696 vdd.n1695 146.341
R19080 vdd.n1700 vdd.n1699 146.341
R19081 vdd.n1702 vdd.n1701 146.341
R19082 vdd.n1706 vdd.n1705 146.341
R19083 vdd.n1708 vdd.n1707 146.341
R19084 vdd.n1714 vdd.n1713 146.341
R19085 vdd.n1716 vdd.n1715 146.341
R19086 vdd.n1720 vdd.n1719 146.341
R19087 vdd.n1722 vdd.n1721 146.341
R19088 vdd.n1726 vdd.n1725 146.341
R19089 vdd.n1728 vdd.n1727 146.341
R19090 vdd.n1732 vdd.n1731 146.341
R19091 vdd.n1734 vdd.n1733 146.341
R19092 vdd.n1738 vdd.n1737 146.341
R19093 vdd.n1740 vdd.n1739 146.341
R19094 vdd.n1812 vdd.n1743 146.341
R19095 vdd.n1745 vdd.n1744 146.341
R19096 vdd.n1749 vdd.n1748 146.341
R19097 vdd.n1751 vdd.n1750 146.341
R19098 vdd.n1755 vdd.n1754 146.341
R19099 vdd.n1757 vdd.n1756 146.341
R19100 vdd.n1761 vdd.n1760 146.341
R19101 vdd.n1763 vdd.n1762 146.341
R19102 vdd.n1767 vdd.n1766 146.341
R19103 vdd.n1769 vdd.n1768 146.341
R19104 vdd.n1773 vdd.n1772 146.341
R19105 vdd.n1774 vdd.n1682 146.341
R19106 vdd.n1884 vdd.n1647 146.341
R19107 vdd.n1884 vdd.n1640 146.341
R19108 vdd.n1895 vdd.n1640 146.341
R19109 vdd.n1895 vdd.n1636 146.341
R19110 vdd.n1901 vdd.n1636 146.341
R19111 vdd.n1901 vdd.n1629 146.341
R19112 vdd.n1912 vdd.n1629 146.341
R19113 vdd.n1912 vdd.n1625 146.341
R19114 vdd.n1919 vdd.n1625 146.341
R19115 vdd.n1919 vdd.n1618 146.341
R19116 vdd.n1929 vdd.n1618 146.341
R19117 vdd.n1929 vdd.n1344 146.341
R19118 vdd.n1935 vdd.n1344 146.341
R19119 vdd.n1935 vdd.n1336 146.341
R19120 vdd.n1946 vdd.n1336 146.341
R19121 vdd.n1946 vdd.n1332 146.341
R19122 vdd.n1952 vdd.n1332 146.341
R19123 vdd.n1952 vdd.n1324 146.341
R19124 vdd.n1965 vdd.n1324 146.341
R19125 vdd.n1965 vdd.n1319 146.341
R19126 vdd.n1971 vdd.n1319 146.341
R19127 vdd.n1105 vdd.t74 127.284
R19128 vdd.n800 vdd.t118 127.284
R19129 vdd.n1109 vdd.t115 127.284
R19130 vdd.n791 vdd.t135 127.284
R19131 vdd.n686 vdd.t91 127.284
R19132 vdd.n686 vdd.t92 127.284
R19133 vdd.n2437 vdd.t133 127.284
R19134 vdd.n622 vdd.t83 127.284
R19135 vdd.n2434 vdd.t126 127.284
R19136 vdd.n589 vdd.t69 127.284
R19137 vdd.n861 vdd.t129 127.284
R19138 vdd.n861 vdd.t130 127.284
R19139 vdd.n22 vdd.n20 117.314
R19140 vdd.n17 vdd.n15 117.314
R19141 vdd.n27 vdd.n26 116.927
R19142 vdd.n24 vdd.n23 116.927
R19143 vdd.n22 vdd.n21 116.927
R19144 vdd.n17 vdd.n16 116.927
R19145 vdd.n19 vdd.n18 116.927
R19146 vdd.n27 vdd.n25 116.927
R19147 vdd.n1106 vdd.t73 111.188
R19148 vdd.n801 vdd.t119 111.188
R19149 vdd.n1110 vdd.t114 111.188
R19150 vdd.n792 vdd.t136 111.188
R19151 vdd.n2438 vdd.t132 111.188
R19152 vdd.n623 vdd.t84 111.188
R19153 vdd.n2435 vdd.t125 111.188
R19154 vdd.n590 vdd.t70 111.188
R19155 vdd.n2708 vdd.n750 99.5127
R19156 vdd.n2708 vdd.n741 99.5127
R19157 vdd.n2716 vdd.n741 99.5127
R19158 vdd.n2716 vdd.n739 99.5127
R19159 vdd.n2720 vdd.n739 99.5127
R19160 vdd.n2720 vdd.n729 99.5127
R19161 vdd.n2728 vdd.n729 99.5127
R19162 vdd.n2728 vdd.n727 99.5127
R19163 vdd.n2732 vdd.n727 99.5127
R19164 vdd.n2732 vdd.n718 99.5127
R19165 vdd.n2740 vdd.n718 99.5127
R19166 vdd.n2740 vdd.n716 99.5127
R19167 vdd.n2744 vdd.n716 99.5127
R19168 vdd.n2744 vdd.n707 99.5127
R19169 vdd.n2752 vdd.n707 99.5127
R19170 vdd.n2752 vdd.n705 99.5127
R19171 vdd.n2756 vdd.n705 99.5127
R19172 vdd.n2756 vdd.n694 99.5127
R19173 vdd.n2765 vdd.n694 99.5127
R19174 vdd.n2765 vdd.n692 99.5127
R19175 vdd.n2769 vdd.n692 99.5127
R19176 vdd.n2769 vdd.n682 99.5127
R19177 vdd.n2777 vdd.n682 99.5127
R19178 vdd.n2777 vdd.n680 99.5127
R19179 vdd.n2781 vdd.n680 99.5127
R19180 vdd.n2781 vdd.n670 99.5127
R19181 vdd.n2789 vdd.n670 99.5127
R19182 vdd.n2789 vdd.n668 99.5127
R19183 vdd.n2793 vdd.n668 99.5127
R19184 vdd.n2793 vdd.n657 99.5127
R19185 vdd.n2801 vdd.n657 99.5127
R19186 vdd.n2801 vdd.n655 99.5127
R19187 vdd.n2805 vdd.n655 99.5127
R19188 vdd.n2805 vdd.n646 99.5127
R19189 vdd.n2813 vdd.n646 99.5127
R19190 vdd.n2813 vdd.n644 99.5127
R19191 vdd.n2817 vdd.n644 99.5127
R19192 vdd.n2817 vdd.n632 99.5127
R19193 vdd.n2870 vdd.n632 99.5127
R19194 vdd.n2870 vdd.n630 99.5127
R19195 vdd.n2874 vdd.n630 99.5127
R19196 vdd.n2874 vdd.n598 99.5127
R19197 vdd.n2944 vdd.n598 99.5127
R19198 vdd.n2940 vdd.n599 99.5127
R19199 vdd.n2938 vdd.n2937 99.5127
R19200 vdd.n2935 vdd.n603 99.5127
R19201 vdd.n2931 vdd.n2930 99.5127
R19202 vdd.n2928 vdd.n606 99.5127
R19203 vdd.n2924 vdd.n2923 99.5127
R19204 vdd.n2921 vdd.n609 99.5127
R19205 vdd.n2917 vdd.n2916 99.5127
R19206 vdd.n2914 vdd.n2912 99.5127
R19207 vdd.n2910 vdd.n612 99.5127
R19208 vdd.n2906 vdd.n2905 99.5127
R19209 vdd.n2903 vdd.n615 99.5127
R19210 vdd.n2899 vdd.n2898 99.5127
R19211 vdd.n2896 vdd.n618 99.5127
R19212 vdd.n2892 vdd.n2891 99.5127
R19213 vdd.n2889 vdd.n621 99.5127
R19214 vdd.n2884 vdd.n2883 99.5127
R19215 vdd.n2635 vdd.n748 99.5127
R19216 vdd.n2631 vdd.n748 99.5127
R19217 vdd.n2631 vdd.n742 99.5127
R19218 vdd.n2513 vdd.n742 99.5127
R19219 vdd.n2513 vdd.n737 99.5127
R19220 vdd.n2516 vdd.n737 99.5127
R19221 vdd.n2516 vdd.n731 99.5127
R19222 vdd.n2617 vdd.n731 99.5127
R19223 vdd.n2617 vdd.n725 99.5127
R19224 vdd.n2613 vdd.n725 99.5127
R19225 vdd.n2613 vdd.n719 99.5127
R19226 vdd.n2560 vdd.n719 99.5127
R19227 vdd.n2560 vdd.n713 99.5127
R19228 vdd.n2557 vdd.n713 99.5127
R19229 vdd.n2557 vdd.n708 99.5127
R19230 vdd.n2554 vdd.n708 99.5127
R19231 vdd.n2554 vdd.n703 99.5127
R19232 vdd.n2551 vdd.n703 99.5127
R19233 vdd.n2551 vdd.n696 99.5127
R19234 vdd.n2548 vdd.n696 99.5127
R19235 vdd.n2548 vdd.n689 99.5127
R19236 vdd.n2545 vdd.n689 99.5127
R19237 vdd.n2545 vdd.n683 99.5127
R19238 vdd.n2542 vdd.n683 99.5127
R19239 vdd.n2542 vdd.n678 99.5127
R19240 vdd.n2539 vdd.n678 99.5127
R19241 vdd.n2539 vdd.n672 99.5127
R19242 vdd.n2536 vdd.n672 99.5127
R19243 vdd.n2536 vdd.n665 99.5127
R19244 vdd.n2533 vdd.n665 99.5127
R19245 vdd.n2533 vdd.n658 99.5127
R19246 vdd.n2530 vdd.n658 99.5127
R19247 vdd.n2530 vdd.n652 99.5127
R19248 vdd.n2527 vdd.n652 99.5127
R19249 vdd.n2527 vdd.n647 99.5127
R19250 vdd.n2524 vdd.n647 99.5127
R19251 vdd.n2524 vdd.n642 99.5127
R19252 vdd.n2521 vdd.n642 99.5127
R19253 vdd.n2521 vdd.n634 99.5127
R19254 vdd.n634 vdd.n627 99.5127
R19255 vdd.n2876 vdd.n627 99.5127
R19256 vdd.n2877 vdd.n2876 99.5127
R19257 vdd.n2877 vdd.n596 99.5127
R19258 vdd.n2701 vdd.n752 99.5127
R19259 vdd.n2701 vdd.n2433 99.5127
R19260 vdd.n2697 vdd.n2696 99.5127
R19261 vdd.n2693 vdd.n2692 99.5127
R19262 vdd.n2689 vdd.n2688 99.5127
R19263 vdd.n2685 vdd.n2684 99.5127
R19264 vdd.n2681 vdd.n2680 99.5127
R19265 vdd.n2677 vdd.n2676 99.5127
R19266 vdd.n2673 vdd.n2672 99.5127
R19267 vdd.n2669 vdd.n2668 99.5127
R19268 vdd.n2665 vdd.n2664 99.5127
R19269 vdd.n2661 vdd.n2660 99.5127
R19270 vdd.n2657 vdd.n2656 99.5127
R19271 vdd.n2653 vdd.n2652 99.5127
R19272 vdd.n2649 vdd.n2648 99.5127
R19273 vdd.n2645 vdd.n2644 99.5127
R19274 vdd.n2640 vdd.n2639 99.5127
R19275 vdd.n2397 vdd.n789 99.5127
R19276 vdd.n2393 vdd.n2392 99.5127
R19277 vdd.n2389 vdd.n2388 99.5127
R19278 vdd.n2385 vdd.n2384 99.5127
R19279 vdd.n2381 vdd.n2380 99.5127
R19280 vdd.n2377 vdd.n2376 99.5127
R19281 vdd.n2373 vdd.n2372 99.5127
R19282 vdd.n2369 vdd.n2368 99.5127
R19283 vdd.n2365 vdd.n2364 99.5127
R19284 vdd.n2361 vdd.n2360 99.5127
R19285 vdd.n2357 vdd.n2356 99.5127
R19286 vdd.n2353 vdd.n2352 99.5127
R19287 vdd.n2349 vdd.n2348 99.5127
R19288 vdd.n2345 vdd.n2344 99.5127
R19289 vdd.n2341 vdd.n2340 99.5127
R19290 vdd.n2337 vdd.n2336 99.5127
R19291 vdd.n2332 vdd.n2331 99.5127
R19292 vdd.n1145 vdd.n925 99.5127
R19293 vdd.n1148 vdd.n925 99.5127
R19294 vdd.n1148 vdd.n919 99.5127
R19295 vdd.n1151 vdd.n919 99.5127
R19296 vdd.n1151 vdd.n914 99.5127
R19297 vdd.n1154 vdd.n914 99.5127
R19298 vdd.n1154 vdd.n907 99.5127
R19299 vdd.n1157 vdd.n907 99.5127
R19300 vdd.n1157 vdd.n900 99.5127
R19301 vdd.n1160 vdd.n900 99.5127
R19302 vdd.n1160 vdd.n894 99.5127
R19303 vdd.n1163 vdd.n894 99.5127
R19304 vdd.n1163 vdd.n889 99.5127
R19305 vdd.n1166 vdd.n889 99.5127
R19306 vdd.n1166 vdd.n884 99.5127
R19307 vdd.n1169 vdd.n884 99.5127
R19308 vdd.n1169 vdd.n878 99.5127
R19309 vdd.n1172 vdd.n878 99.5127
R19310 vdd.n1172 vdd.n871 99.5127
R19311 vdd.n1175 vdd.n871 99.5127
R19312 vdd.n1175 vdd.n864 99.5127
R19313 vdd.n1178 vdd.n864 99.5127
R19314 vdd.n1178 vdd.n858 99.5127
R19315 vdd.n1181 vdd.n858 99.5127
R19316 vdd.n1181 vdd.n853 99.5127
R19317 vdd.n1184 vdd.n853 99.5127
R19318 vdd.n1184 vdd.n847 99.5127
R19319 vdd.n1226 vdd.n847 99.5127
R19320 vdd.n1226 vdd.n840 99.5127
R19321 vdd.n1222 vdd.n840 99.5127
R19322 vdd.n1222 vdd.n834 99.5127
R19323 vdd.n1219 vdd.n834 99.5127
R19324 vdd.n1219 vdd.n829 99.5127
R19325 vdd.n1216 vdd.n829 99.5127
R19326 vdd.n1216 vdd.n824 99.5127
R19327 vdd.n1196 vdd.n824 99.5127
R19328 vdd.n1196 vdd.n819 99.5127
R19329 vdd.n1193 vdd.n819 99.5127
R19330 vdd.n1193 vdd.n812 99.5127
R19331 vdd.n1190 vdd.n812 99.5127
R19332 vdd.n1190 vdd.n805 99.5127
R19333 vdd.n805 vdd.n794 99.5127
R19334 vdd.n2327 vdd.n794 99.5127
R19335 vdd.n2119 vdd.n930 99.5127
R19336 vdd.n2119 vdd.n966 99.5127
R19337 vdd.n2115 vdd.n2114 99.5127
R19338 vdd.n2111 vdd.n2110 99.5127
R19339 vdd.n2107 vdd.n2106 99.5127
R19340 vdd.n2103 vdd.n2102 99.5127
R19341 vdd.n2099 vdd.n2098 99.5127
R19342 vdd.n2095 vdd.n2094 99.5127
R19343 vdd.n2091 vdd.n2090 99.5127
R19344 vdd.n1112 vdd.n1111 99.5127
R19345 vdd.n1116 vdd.n1115 99.5127
R19346 vdd.n1120 vdd.n1119 99.5127
R19347 vdd.n1124 vdd.n1123 99.5127
R19348 vdd.n1128 vdd.n1127 99.5127
R19349 vdd.n1132 vdd.n1131 99.5127
R19350 vdd.n1136 vdd.n1135 99.5127
R19351 vdd.n1141 vdd.n1140 99.5127
R19352 vdd.n2126 vdd.n928 99.5127
R19353 vdd.n2126 vdd.n918 99.5127
R19354 vdd.n2134 vdd.n918 99.5127
R19355 vdd.n2134 vdd.n916 99.5127
R19356 vdd.n2138 vdd.n916 99.5127
R19357 vdd.n2138 vdd.n905 99.5127
R19358 vdd.n2146 vdd.n905 99.5127
R19359 vdd.n2146 vdd.n903 99.5127
R19360 vdd.n2150 vdd.n903 99.5127
R19361 vdd.n2150 vdd.n893 99.5127
R19362 vdd.n2158 vdd.n893 99.5127
R19363 vdd.n2158 vdd.n891 99.5127
R19364 vdd.n2162 vdd.n891 99.5127
R19365 vdd.n2162 vdd.n882 99.5127
R19366 vdd.n2170 vdd.n882 99.5127
R19367 vdd.n2170 vdd.n880 99.5127
R19368 vdd.n2174 vdd.n880 99.5127
R19369 vdd.n2174 vdd.n869 99.5127
R19370 vdd.n2182 vdd.n869 99.5127
R19371 vdd.n2182 vdd.n867 99.5127
R19372 vdd.n2186 vdd.n867 99.5127
R19373 vdd.n2186 vdd.n857 99.5127
R19374 vdd.n2195 vdd.n857 99.5127
R19375 vdd.n2195 vdd.n855 99.5127
R19376 vdd.n2199 vdd.n855 99.5127
R19377 vdd.n2199 vdd.n845 99.5127
R19378 vdd.n2207 vdd.n845 99.5127
R19379 vdd.n2207 vdd.n843 99.5127
R19380 vdd.n2211 vdd.n843 99.5127
R19381 vdd.n2211 vdd.n833 99.5127
R19382 vdd.n2219 vdd.n833 99.5127
R19383 vdd.n2219 vdd.n831 99.5127
R19384 vdd.n2223 vdd.n831 99.5127
R19385 vdd.n2223 vdd.n823 99.5127
R19386 vdd.n2231 vdd.n823 99.5127
R19387 vdd.n2231 vdd.n821 99.5127
R19388 vdd.n2235 vdd.n821 99.5127
R19389 vdd.n2235 vdd.n810 99.5127
R19390 vdd.n2245 vdd.n810 99.5127
R19391 vdd.n2245 vdd.n807 99.5127
R19392 vdd.n2250 vdd.n807 99.5127
R19393 vdd.n2250 vdd.n808 99.5127
R19394 vdd.n808 vdd.n788 99.5127
R19395 vdd.n2860 vdd.n2859 99.5127
R19396 vdd.n2857 vdd.n2823 99.5127
R19397 vdd.n2853 vdd.n2852 99.5127
R19398 vdd.n2850 vdd.n2826 99.5127
R19399 vdd.n2846 vdd.n2845 99.5127
R19400 vdd.n2843 vdd.n2829 99.5127
R19401 vdd.n2839 vdd.n2838 99.5127
R19402 vdd.n2836 vdd.n2833 99.5127
R19403 vdd.n2977 vdd.n577 99.5127
R19404 vdd.n2975 vdd.n2974 99.5127
R19405 vdd.n2972 vdd.n579 99.5127
R19406 vdd.n2968 vdd.n2967 99.5127
R19407 vdd.n2965 vdd.n582 99.5127
R19408 vdd.n2961 vdd.n2960 99.5127
R19409 vdd.n2958 vdd.n585 99.5127
R19410 vdd.n2954 vdd.n2953 99.5127
R19411 vdd.n2951 vdd.n588 99.5127
R19412 vdd.n2509 vdd.n749 99.5127
R19413 vdd.n2629 vdd.n749 99.5127
R19414 vdd.n2629 vdd.n743 99.5127
R19415 vdd.n2625 vdd.n743 99.5127
R19416 vdd.n2625 vdd.n738 99.5127
R19417 vdd.n2622 vdd.n738 99.5127
R19418 vdd.n2622 vdd.n732 99.5127
R19419 vdd.n2619 vdd.n732 99.5127
R19420 vdd.n2619 vdd.n726 99.5127
R19421 vdd.n2611 vdd.n726 99.5127
R19422 vdd.n2611 vdd.n720 99.5127
R19423 vdd.n2607 vdd.n720 99.5127
R19424 vdd.n2607 vdd.n714 99.5127
R19425 vdd.n2604 vdd.n714 99.5127
R19426 vdd.n2604 vdd.n709 99.5127
R19427 vdd.n2601 vdd.n709 99.5127
R19428 vdd.n2601 vdd.n704 99.5127
R19429 vdd.n2598 vdd.n704 99.5127
R19430 vdd.n2598 vdd.n697 99.5127
R19431 vdd.n2595 vdd.n697 99.5127
R19432 vdd.n2595 vdd.n690 99.5127
R19433 vdd.n2592 vdd.n690 99.5127
R19434 vdd.n2592 vdd.n684 99.5127
R19435 vdd.n2589 vdd.n684 99.5127
R19436 vdd.n2589 vdd.n679 99.5127
R19437 vdd.n2586 vdd.n679 99.5127
R19438 vdd.n2586 vdd.n673 99.5127
R19439 vdd.n2583 vdd.n673 99.5127
R19440 vdd.n2583 vdd.n666 99.5127
R19441 vdd.n2580 vdd.n666 99.5127
R19442 vdd.n2580 vdd.n659 99.5127
R19443 vdd.n2577 vdd.n659 99.5127
R19444 vdd.n2577 vdd.n653 99.5127
R19445 vdd.n2574 vdd.n653 99.5127
R19446 vdd.n2574 vdd.n648 99.5127
R19447 vdd.n2571 vdd.n648 99.5127
R19448 vdd.n2571 vdd.n643 99.5127
R19449 vdd.n2568 vdd.n643 99.5127
R19450 vdd.n2568 vdd.n635 99.5127
R19451 vdd.n2565 vdd.n635 99.5127
R19452 vdd.n2565 vdd.n628 99.5127
R19453 vdd.n628 vdd.n594 99.5127
R19454 vdd.n2946 vdd.n594 99.5127
R19455 vdd.n2444 vdd.n2443 99.5127
R19456 vdd.n2448 vdd.n2447 99.5127
R19457 vdd.n2452 vdd.n2451 99.5127
R19458 vdd.n2456 vdd.n2455 99.5127
R19459 vdd.n2460 vdd.n2459 99.5127
R19460 vdd.n2464 vdd.n2463 99.5127
R19461 vdd.n2468 vdd.n2467 99.5127
R19462 vdd.n2472 vdd.n2471 99.5127
R19463 vdd.n2476 vdd.n2475 99.5127
R19464 vdd.n2480 vdd.n2479 99.5127
R19465 vdd.n2484 vdd.n2483 99.5127
R19466 vdd.n2488 vdd.n2487 99.5127
R19467 vdd.n2492 vdd.n2491 99.5127
R19468 vdd.n2496 vdd.n2495 99.5127
R19469 vdd.n2500 vdd.n2499 99.5127
R19470 vdd.n2504 vdd.n2503 99.5127
R19471 vdd.n2506 vdd.n2432 99.5127
R19472 vdd.n2710 vdd.n746 99.5127
R19473 vdd.n2710 vdd.n744 99.5127
R19474 vdd.n2714 vdd.n744 99.5127
R19475 vdd.n2714 vdd.n735 99.5127
R19476 vdd.n2722 vdd.n735 99.5127
R19477 vdd.n2722 vdd.n733 99.5127
R19478 vdd.n2726 vdd.n733 99.5127
R19479 vdd.n2726 vdd.n724 99.5127
R19480 vdd.n2734 vdd.n724 99.5127
R19481 vdd.n2734 vdd.n722 99.5127
R19482 vdd.n2738 vdd.n722 99.5127
R19483 vdd.n2738 vdd.n712 99.5127
R19484 vdd.n2746 vdd.n712 99.5127
R19485 vdd.n2746 vdd.n710 99.5127
R19486 vdd.n2750 vdd.n710 99.5127
R19487 vdd.n2750 vdd.n701 99.5127
R19488 vdd.n2758 vdd.n701 99.5127
R19489 vdd.n2758 vdd.n699 99.5127
R19490 vdd.n2763 vdd.n699 99.5127
R19491 vdd.n2763 vdd.n688 99.5127
R19492 vdd.n2771 vdd.n688 99.5127
R19493 vdd.n2771 vdd.n685 99.5127
R19494 vdd.n2775 vdd.n685 99.5127
R19495 vdd.n2775 vdd.n676 99.5127
R19496 vdd.n2783 vdd.n676 99.5127
R19497 vdd.n2783 vdd.n674 99.5127
R19498 vdd.n2787 vdd.n674 99.5127
R19499 vdd.n2787 vdd.n663 99.5127
R19500 vdd.n2795 vdd.n663 99.5127
R19501 vdd.n2795 vdd.n661 99.5127
R19502 vdd.n2799 vdd.n661 99.5127
R19503 vdd.n2799 vdd.n651 99.5127
R19504 vdd.n2807 vdd.n651 99.5127
R19505 vdd.n2807 vdd.n649 99.5127
R19506 vdd.n2811 vdd.n649 99.5127
R19507 vdd.n2811 vdd.n640 99.5127
R19508 vdd.n2819 vdd.n640 99.5127
R19509 vdd.n2819 vdd.n637 99.5127
R19510 vdd.n2868 vdd.n637 99.5127
R19511 vdd.n2868 vdd.n638 99.5127
R19512 vdd.n638 vdd.n629 99.5127
R19513 vdd.n2863 vdd.n629 99.5127
R19514 vdd.n2863 vdd.n597 99.5127
R19515 vdd.n2321 vdd.n2320 99.5127
R19516 vdd.n2317 vdd.n2316 99.5127
R19517 vdd.n2313 vdd.n2312 99.5127
R19518 vdd.n2309 vdd.n2308 99.5127
R19519 vdd.n2305 vdd.n2304 99.5127
R19520 vdd.n2301 vdd.n2300 99.5127
R19521 vdd.n2297 vdd.n2296 99.5127
R19522 vdd.n2293 vdd.n2292 99.5127
R19523 vdd.n2289 vdd.n2288 99.5127
R19524 vdd.n2285 vdd.n2284 99.5127
R19525 vdd.n2281 vdd.n2280 99.5127
R19526 vdd.n2277 vdd.n2276 99.5127
R19527 vdd.n2273 vdd.n2272 99.5127
R19528 vdd.n2269 vdd.n2268 99.5127
R19529 vdd.n2265 vdd.n2264 99.5127
R19530 vdd.n2261 vdd.n2260 99.5127
R19531 vdd.n2257 vdd.n770 99.5127
R19532 vdd.n1270 vdd.n926 99.5127
R19533 vdd.n1267 vdd.n926 99.5127
R19534 vdd.n1267 vdd.n920 99.5127
R19535 vdd.n1264 vdd.n920 99.5127
R19536 vdd.n1264 vdd.n915 99.5127
R19537 vdd.n1261 vdd.n915 99.5127
R19538 vdd.n1261 vdd.n908 99.5127
R19539 vdd.n1258 vdd.n908 99.5127
R19540 vdd.n1258 vdd.n901 99.5127
R19541 vdd.n1255 vdd.n901 99.5127
R19542 vdd.n1255 vdd.n895 99.5127
R19543 vdd.n1252 vdd.n895 99.5127
R19544 vdd.n1252 vdd.n890 99.5127
R19545 vdd.n1249 vdd.n890 99.5127
R19546 vdd.n1249 vdd.n885 99.5127
R19547 vdd.n1246 vdd.n885 99.5127
R19548 vdd.n1246 vdd.n879 99.5127
R19549 vdd.n1243 vdd.n879 99.5127
R19550 vdd.n1243 vdd.n872 99.5127
R19551 vdd.n1240 vdd.n872 99.5127
R19552 vdd.n1240 vdd.n865 99.5127
R19553 vdd.n1237 vdd.n865 99.5127
R19554 vdd.n1237 vdd.n859 99.5127
R19555 vdd.n1234 vdd.n859 99.5127
R19556 vdd.n1234 vdd.n854 99.5127
R19557 vdd.n1231 vdd.n854 99.5127
R19558 vdd.n1231 vdd.n848 99.5127
R19559 vdd.n1228 vdd.n848 99.5127
R19560 vdd.n1228 vdd.n841 99.5127
R19561 vdd.n1199 vdd.n841 99.5127
R19562 vdd.n1199 vdd.n835 99.5127
R19563 vdd.n1202 vdd.n835 99.5127
R19564 vdd.n1202 vdd.n830 99.5127
R19565 vdd.n1214 vdd.n830 99.5127
R19566 vdd.n1214 vdd.n825 99.5127
R19567 vdd.n1210 vdd.n825 99.5127
R19568 vdd.n1210 vdd.n820 99.5127
R19569 vdd.n1207 vdd.n820 99.5127
R19570 vdd.n1207 vdd.n813 99.5127
R19571 vdd.n813 vdd.n804 99.5127
R19572 vdd.n2252 vdd.n804 99.5127
R19573 vdd.n2253 vdd.n2252 99.5127
R19574 vdd.n2253 vdd.n796 99.5127
R19575 vdd.n1074 vdd.n1073 99.5127
R19576 vdd.n1078 vdd.n1077 99.5127
R19577 vdd.n1082 vdd.n1081 99.5127
R19578 vdd.n1086 vdd.n1085 99.5127
R19579 vdd.n1090 vdd.n1089 99.5127
R19580 vdd.n1094 vdd.n1093 99.5127
R19581 vdd.n1098 vdd.n1097 99.5127
R19582 vdd.n1102 vdd.n1101 99.5127
R19583 vdd.n1303 vdd.n1104 99.5127
R19584 vdd.n1301 vdd.n1300 99.5127
R19585 vdd.n1297 vdd.n1296 99.5127
R19586 vdd.n1293 vdd.n1292 99.5127
R19587 vdd.n1289 vdd.n1288 99.5127
R19588 vdd.n1285 vdd.n1284 99.5127
R19589 vdd.n1281 vdd.n1280 99.5127
R19590 vdd.n1277 vdd.n1276 99.5127
R19591 vdd.n1273 vdd.n965 99.5127
R19592 vdd.n2128 vdd.n923 99.5127
R19593 vdd.n2128 vdd.n921 99.5127
R19594 vdd.n2132 vdd.n921 99.5127
R19595 vdd.n2132 vdd.n912 99.5127
R19596 vdd.n2140 vdd.n912 99.5127
R19597 vdd.n2140 vdd.n910 99.5127
R19598 vdd.n2144 vdd.n910 99.5127
R19599 vdd.n2144 vdd.n899 99.5127
R19600 vdd.n2152 vdd.n899 99.5127
R19601 vdd.n2152 vdd.n897 99.5127
R19602 vdd.n2156 vdd.n897 99.5127
R19603 vdd.n2156 vdd.n888 99.5127
R19604 vdd.n2164 vdd.n888 99.5127
R19605 vdd.n2164 vdd.n886 99.5127
R19606 vdd.n2168 vdd.n886 99.5127
R19607 vdd.n2168 vdd.n876 99.5127
R19608 vdd.n2176 vdd.n876 99.5127
R19609 vdd.n2176 vdd.n874 99.5127
R19610 vdd.n2180 vdd.n874 99.5127
R19611 vdd.n2180 vdd.n863 99.5127
R19612 vdd.n2188 vdd.n863 99.5127
R19613 vdd.n2188 vdd.n860 99.5127
R19614 vdd.n2193 vdd.n860 99.5127
R19615 vdd.n2193 vdd.n851 99.5127
R19616 vdd.n2201 vdd.n851 99.5127
R19617 vdd.n2201 vdd.n849 99.5127
R19618 vdd.n2205 vdd.n849 99.5127
R19619 vdd.n2205 vdd.n839 99.5127
R19620 vdd.n2213 vdd.n839 99.5127
R19621 vdd.n2213 vdd.n837 99.5127
R19622 vdd.n2217 vdd.n837 99.5127
R19623 vdd.n2217 vdd.n828 99.5127
R19624 vdd.n2225 vdd.n828 99.5127
R19625 vdd.n2225 vdd.n826 99.5127
R19626 vdd.n2229 vdd.n826 99.5127
R19627 vdd.n2229 vdd.n817 99.5127
R19628 vdd.n2237 vdd.n817 99.5127
R19629 vdd.n2237 vdd.n814 99.5127
R19630 vdd.n2243 vdd.n814 99.5127
R19631 vdd.n2243 vdd.n815 99.5127
R19632 vdd.n815 vdd.n806 99.5127
R19633 vdd.n806 vdd.n797 99.5127
R19634 vdd.n2325 vdd.n797 99.5127
R19635 vdd.n9 vdd.n7 98.9633
R19636 vdd.n2 vdd.n0 98.9633
R19637 vdd.n9 vdd.n8 98.6055
R19638 vdd.n11 vdd.n10 98.6055
R19639 vdd.n13 vdd.n12 98.6055
R19640 vdd.n6 vdd.n5 98.6055
R19641 vdd.n4 vdd.n3 98.6055
R19642 vdd.n2 vdd.n1 98.6055
R19643 vdd.t201 vdd.n267 85.8723
R19644 vdd.t209 vdd.n220 85.8723
R19645 vdd.t198 vdd.n177 85.8723
R19646 vdd.t206 vdd.n130 85.8723
R19647 vdd.t178 vdd.n88 85.8723
R19648 vdd.t183 vdd.n41 85.8723
R19649 vdd.t176 vdd.n1537 85.8723
R19650 vdd.t162 vdd.n1584 85.8723
R19651 vdd.t171 vdd.n1447 85.8723
R19652 vdd.t151 vdd.n1494 85.8723
R19653 vdd.t184 vdd.n1358 85.8723
R19654 vdd.t179 vdd.n1405 85.8723
R19655 vdd.n687 vdd.n686 78.546
R19656 vdd.n2191 vdd.n861 78.546
R19657 vdd.n254 vdd.n253 75.1835
R19658 vdd.n252 vdd.n251 75.1835
R19659 vdd.n250 vdd.n249 75.1835
R19660 vdd.n164 vdd.n163 75.1835
R19661 vdd.n162 vdd.n161 75.1835
R19662 vdd.n160 vdd.n159 75.1835
R19663 vdd.n75 vdd.n74 75.1835
R19664 vdd.n73 vdd.n72 75.1835
R19665 vdd.n71 vdd.n70 75.1835
R19666 vdd.n1567 vdd.n1566 75.1835
R19667 vdd.n1569 vdd.n1568 75.1835
R19668 vdd.n1571 vdd.n1570 75.1835
R19669 vdd.n1477 vdd.n1476 75.1835
R19670 vdd.n1479 vdd.n1478 75.1835
R19671 vdd.n1481 vdd.n1480 75.1835
R19672 vdd.n1388 vdd.n1387 75.1835
R19673 vdd.n1390 vdd.n1389 75.1835
R19674 vdd.n1392 vdd.n1391 75.1835
R19675 vdd.n2702 vdd.n2415 72.8958
R19676 vdd.n2702 vdd.n2416 72.8958
R19677 vdd.n2702 vdd.n2417 72.8958
R19678 vdd.n2702 vdd.n2418 72.8958
R19679 vdd.n2702 vdd.n2419 72.8958
R19680 vdd.n2702 vdd.n2420 72.8958
R19681 vdd.n2702 vdd.n2421 72.8958
R19682 vdd.n2702 vdd.n2422 72.8958
R19683 vdd.n2702 vdd.n2423 72.8958
R19684 vdd.n2702 vdd.n2424 72.8958
R19685 vdd.n2702 vdd.n2425 72.8958
R19686 vdd.n2702 vdd.n2426 72.8958
R19687 vdd.n2702 vdd.n2427 72.8958
R19688 vdd.n2702 vdd.n2428 72.8958
R19689 vdd.n2702 vdd.n2429 72.8958
R19690 vdd.n2702 vdd.n2430 72.8958
R19691 vdd.n2702 vdd.n2431 72.8958
R19692 vdd.n593 vdd.n484 72.8958
R19693 vdd.n2952 vdd.n484 72.8958
R19694 vdd.n587 vdd.n484 72.8958
R19695 vdd.n2959 vdd.n484 72.8958
R19696 vdd.n584 vdd.n484 72.8958
R19697 vdd.n2966 vdd.n484 72.8958
R19698 vdd.n581 vdd.n484 72.8958
R19699 vdd.n2973 vdd.n484 72.8958
R19700 vdd.n2976 vdd.n484 72.8958
R19701 vdd.n2832 vdd.n484 72.8958
R19702 vdd.n2837 vdd.n484 72.8958
R19703 vdd.n2831 vdd.n484 72.8958
R19704 vdd.n2844 vdd.n484 72.8958
R19705 vdd.n2828 vdd.n484 72.8958
R19706 vdd.n2851 vdd.n484 72.8958
R19707 vdd.n2825 vdd.n484 72.8958
R19708 vdd.n2858 vdd.n484 72.8958
R19709 vdd.n2121 vdd.n2120 72.8958
R19710 vdd.n2120 vdd.n932 72.8958
R19711 vdd.n2120 vdd.n933 72.8958
R19712 vdd.n2120 vdd.n934 72.8958
R19713 vdd.n2120 vdd.n935 72.8958
R19714 vdd.n2120 vdd.n936 72.8958
R19715 vdd.n2120 vdd.n937 72.8958
R19716 vdd.n2120 vdd.n938 72.8958
R19717 vdd.n2120 vdd.n939 72.8958
R19718 vdd.n2120 vdd.n940 72.8958
R19719 vdd.n2120 vdd.n941 72.8958
R19720 vdd.n2120 vdd.n942 72.8958
R19721 vdd.n2120 vdd.n943 72.8958
R19722 vdd.n2120 vdd.n944 72.8958
R19723 vdd.n2120 vdd.n945 72.8958
R19724 vdd.n2120 vdd.n946 72.8958
R19725 vdd.n2120 vdd.n947 72.8958
R19726 vdd.n2398 vdd.n771 72.8958
R19727 vdd.n2398 vdd.n772 72.8958
R19728 vdd.n2398 vdd.n773 72.8958
R19729 vdd.n2398 vdd.n774 72.8958
R19730 vdd.n2398 vdd.n775 72.8958
R19731 vdd.n2398 vdd.n776 72.8958
R19732 vdd.n2398 vdd.n777 72.8958
R19733 vdd.n2398 vdd.n778 72.8958
R19734 vdd.n2398 vdd.n779 72.8958
R19735 vdd.n2398 vdd.n780 72.8958
R19736 vdd.n2398 vdd.n781 72.8958
R19737 vdd.n2398 vdd.n782 72.8958
R19738 vdd.n2398 vdd.n783 72.8958
R19739 vdd.n2398 vdd.n784 72.8958
R19740 vdd.n2398 vdd.n785 72.8958
R19741 vdd.n2398 vdd.n786 72.8958
R19742 vdd.n2398 vdd.n787 72.8958
R19743 vdd.n2703 vdd.n2702 72.8958
R19744 vdd.n2702 vdd.n2399 72.8958
R19745 vdd.n2702 vdd.n2400 72.8958
R19746 vdd.n2702 vdd.n2401 72.8958
R19747 vdd.n2702 vdd.n2402 72.8958
R19748 vdd.n2702 vdd.n2403 72.8958
R19749 vdd.n2702 vdd.n2404 72.8958
R19750 vdd.n2702 vdd.n2405 72.8958
R19751 vdd.n2702 vdd.n2406 72.8958
R19752 vdd.n2702 vdd.n2407 72.8958
R19753 vdd.n2702 vdd.n2408 72.8958
R19754 vdd.n2702 vdd.n2409 72.8958
R19755 vdd.n2702 vdd.n2410 72.8958
R19756 vdd.n2702 vdd.n2411 72.8958
R19757 vdd.n2702 vdd.n2412 72.8958
R19758 vdd.n2702 vdd.n2413 72.8958
R19759 vdd.n2702 vdd.n2414 72.8958
R19760 vdd.n2882 vdd.n484 72.8958
R19761 vdd.n625 vdd.n484 72.8958
R19762 vdd.n2890 vdd.n484 72.8958
R19763 vdd.n620 vdd.n484 72.8958
R19764 vdd.n2897 vdd.n484 72.8958
R19765 vdd.n617 vdd.n484 72.8958
R19766 vdd.n2904 vdd.n484 72.8958
R19767 vdd.n614 vdd.n484 72.8958
R19768 vdd.n2911 vdd.n484 72.8958
R19769 vdd.n2915 vdd.n484 72.8958
R19770 vdd.n611 vdd.n484 72.8958
R19771 vdd.n2922 vdd.n484 72.8958
R19772 vdd.n608 vdd.n484 72.8958
R19773 vdd.n2929 vdd.n484 72.8958
R19774 vdd.n605 vdd.n484 72.8958
R19775 vdd.n2936 vdd.n484 72.8958
R19776 vdd.n2939 vdd.n484 72.8958
R19777 vdd.n2398 vdd.n769 72.8958
R19778 vdd.n2398 vdd.n768 72.8958
R19779 vdd.n2398 vdd.n767 72.8958
R19780 vdd.n2398 vdd.n766 72.8958
R19781 vdd.n2398 vdd.n765 72.8958
R19782 vdd.n2398 vdd.n764 72.8958
R19783 vdd.n2398 vdd.n763 72.8958
R19784 vdd.n2398 vdd.n762 72.8958
R19785 vdd.n2398 vdd.n761 72.8958
R19786 vdd.n2398 vdd.n760 72.8958
R19787 vdd.n2398 vdd.n759 72.8958
R19788 vdd.n2398 vdd.n758 72.8958
R19789 vdd.n2398 vdd.n757 72.8958
R19790 vdd.n2398 vdd.n756 72.8958
R19791 vdd.n2398 vdd.n755 72.8958
R19792 vdd.n2398 vdd.n754 72.8958
R19793 vdd.n2398 vdd.n753 72.8958
R19794 vdd.n2120 vdd.n948 72.8958
R19795 vdd.n2120 vdd.n949 72.8958
R19796 vdd.n2120 vdd.n950 72.8958
R19797 vdd.n2120 vdd.n951 72.8958
R19798 vdd.n2120 vdd.n952 72.8958
R19799 vdd.n2120 vdd.n953 72.8958
R19800 vdd.n2120 vdd.n954 72.8958
R19801 vdd.n2120 vdd.n955 72.8958
R19802 vdd.n2120 vdd.n956 72.8958
R19803 vdd.n2120 vdd.n957 72.8958
R19804 vdd.n2120 vdd.n958 72.8958
R19805 vdd.n2120 vdd.n959 72.8958
R19806 vdd.n2120 vdd.n960 72.8958
R19807 vdd.n2120 vdd.n961 72.8958
R19808 vdd.n2120 vdd.n962 72.8958
R19809 vdd.n2120 vdd.n963 72.8958
R19810 vdd.n2120 vdd.n964 72.8958
R19811 vdd.n1877 vdd.n1876 66.2847
R19812 vdd.n1876 vdd.n1652 66.2847
R19813 vdd.n1876 vdd.n1653 66.2847
R19814 vdd.n1876 vdd.n1654 66.2847
R19815 vdd.n1876 vdd.n1655 66.2847
R19816 vdd.n1876 vdd.n1656 66.2847
R19817 vdd.n1876 vdd.n1657 66.2847
R19818 vdd.n1876 vdd.n1658 66.2847
R19819 vdd.n1876 vdd.n1659 66.2847
R19820 vdd.n1876 vdd.n1660 66.2847
R19821 vdd.n1876 vdd.n1661 66.2847
R19822 vdd.n1876 vdd.n1662 66.2847
R19823 vdd.n1876 vdd.n1663 66.2847
R19824 vdd.n1876 vdd.n1664 66.2847
R19825 vdd.n1876 vdd.n1665 66.2847
R19826 vdd.n1876 vdd.n1666 66.2847
R19827 vdd.n1876 vdd.n1667 66.2847
R19828 vdd.n1876 vdd.n1668 66.2847
R19829 vdd.n1876 vdd.n1669 66.2847
R19830 vdd.n1876 vdd.n1670 66.2847
R19831 vdd.n1876 vdd.n1671 66.2847
R19832 vdd.n1876 vdd.n1672 66.2847
R19833 vdd.n1876 vdd.n1673 66.2847
R19834 vdd.n1876 vdd.n1674 66.2847
R19835 vdd.n1876 vdd.n1675 66.2847
R19836 vdd.n1876 vdd.n1676 66.2847
R19837 vdd.n1876 vdd.n1677 66.2847
R19838 vdd.n1876 vdd.n1678 66.2847
R19839 vdd.n1876 vdd.n1679 66.2847
R19840 vdd.n1876 vdd.n1680 66.2847
R19841 vdd.n1876 vdd.n1681 66.2847
R19842 vdd.n1316 vdd.n931 66.2847
R19843 vdd.n1313 vdd.n931 66.2847
R19844 vdd.n1309 vdd.n931 66.2847
R19845 vdd.n1986 vdd.n931 66.2847
R19846 vdd.n1065 vdd.n931 66.2847
R19847 vdd.n1993 vdd.n931 66.2847
R19848 vdd.n1058 vdd.n931 66.2847
R19849 vdd.n2000 vdd.n931 66.2847
R19850 vdd.n1051 vdd.n931 66.2847
R19851 vdd.n2007 vdd.n931 66.2847
R19852 vdd.n1045 vdd.n931 66.2847
R19853 vdd.n1040 vdd.n931 66.2847
R19854 vdd.n2018 vdd.n931 66.2847
R19855 vdd.n1032 vdd.n931 66.2847
R19856 vdd.n2025 vdd.n931 66.2847
R19857 vdd.n1025 vdd.n931 66.2847
R19858 vdd.n2032 vdd.n931 66.2847
R19859 vdd.n1018 vdd.n931 66.2847
R19860 vdd.n2039 vdd.n931 66.2847
R19861 vdd.n1011 vdd.n931 66.2847
R19862 vdd.n2046 vdd.n931 66.2847
R19863 vdd.n1005 vdd.n931 66.2847
R19864 vdd.n1000 vdd.n931 66.2847
R19865 vdd.n2057 vdd.n931 66.2847
R19866 vdd.n992 vdd.n931 66.2847
R19867 vdd.n2064 vdd.n931 66.2847
R19868 vdd.n985 vdd.n931 66.2847
R19869 vdd.n2071 vdd.n931 66.2847
R19870 vdd.n978 vdd.n931 66.2847
R19871 vdd.n2078 vdd.n931 66.2847
R19872 vdd.n2083 vdd.n931 66.2847
R19873 vdd.n974 vdd.n931 66.2847
R19874 vdd.n3113 vdd.n3112 66.2847
R19875 vdd.n3112 vdd.n485 66.2847
R19876 vdd.n3112 vdd.n486 66.2847
R19877 vdd.n3112 vdd.n487 66.2847
R19878 vdd.n3112 vdd.n488 66.2847
R19879 vdd.n3112 vdd.n489 66.2847
R19880 vdd.n3112 vdd.n490 66.2847
R19881 vdd.n3112 vdd.n491 66.2847
R19882 vdd.n3112 vdd.n492 66.2847
R19883 vdd.n3112 vdd.n493 66.2847
R19884 vdd.n3112 vdd.n494 66.2847
R19885 vdd.n3112 vdd.n495 66.2847
R19886 vdd.n3112 vdd.n496 66.2847
R19887 vdd.n3112 vdd.n497 66.2847
R19888 vdd.n3112 vdd.n498 66.2847
R19889 vdd.n3112 vdd.n499 66.2847
R19890 vdd.n3112 vdd.n500 66.2847
R19891 vdd.n3112 vdd.n501 66.2847
R19892 vdd.n3112 vdd.n502 66.2847
R19893 vdd.n3112 vdd.n503 66.2847
R19894 vdd.n3112 vdd.n504 66.2847
R19895 vdd.n3112 vdd.n505 66.2847
R19896 vdd.n3112 vdd.n506 66.2847
R19897 vdd.n3112 vdd.n507 66.2847
R19898 vdd.n3112 vdd.n508 66.2847
R19899 vdd.n3112 vdd.n509 66.2847
R19900 vdd.n3112 vdd.n510 66.2847
R19901 vdd.n3112 vdd.n511 66.2847
R19902 vdd.n3112 vdd.n512 66.2847
R19903 vdd.n3112 vdd.n513 66.2847
R19904 vdd.n3112 vdd.n514 66.2847
R19905 vdd.n3177 vdd.n329 66.2847
R19906 vdd.n3186 vdd.n329 66.2847
R19907 vdd.n439 vdd.n329 66.2847
R19908 vdd.n3193 vdd.n329 66.2847
R19909 vdd.n432 vdd.n329 66.2847
R19910 vdd.n3200 vdd.n329 66.2847
R19911 vdd.n425 vdd.n329 66.2847
R19912 vdd.n3207 vdd.n329 66.2847
R19913 vdd.n418 vdd.n329 66.2847
R19914 vdd.n3214 vdd.n329 66.2847
R19915 vdd.n412 vdd.n329 66.2847
R19916 vdd.n407 vdd.n329 66.2847
R19917 vdd.n3225 vdd.n329 66.2847
R19918 vdd.n399 vdd.n329 66.2847
R19919 vdd.n3232 vdd.n329 66.2847
R19920 vdd.n392 vdd.n329 66.2847
R19921 vdd.n3239 vdd.n329 66.2847
R19922 vdd.n385 vdd.n329 66.2847
R19923 vdd.n3246 vdd.n329 66.2847
R19924 vdd.n378 vdd.n329 66.2847
R19925 vdd.n3253 vdd.n329 66.2847
R19926 vdd.n372 vdd.n329 66.2847
R19927 vdd.n367 vdd.n329 66.2847
R19928 vdd.n3264 vdd.n329 66.2847
R19929 vdd.n359 vdd.n329 66.2847
R19930 vdd.n3271 vdd.n329 66.2847
R19931 vdd.n352 vdd.n329 66.2847
R19932 vdd.n3278 vdd.n329 66.2847
R19933 vdd.n345 vdd.n329 66.2847
R19934 vdd.n3285 vdd.n329 66.2847
R19935 vdd.n3288 vdd.n329 66.2847
R19936 vdd.n333 vdd.n329 66.2847
R19937 vdd.n334 vdd.n333 52.4337
R19938 vdd.n3288 vdd.n3287 52.4337
R19939 vdd.n3285 vdd.n3284 52.4337
R19940 vdd.n3280 vdd.n345 52.4337
R19941 vdd.n3278 vdd.n3277 52.4337
R19942 vdd.n3273 vdd.n352 52.4337
R19943 vdd.n3271 vdd.n3270 52.4337
R19944 vdd.n3266 vdd.n359 52.4337
R19945 vdd.n3264 vdd.n3263 52.4337
R19946 vdd.n368 vdd.n367 52.4337
R19947 vdd.n3255 vdd.n372 52.4337
R19948 vdd.n3253 vdd.n3252 52.4337
R19949 vdd.n3248 vdd.n378 52.4337
R19950 vdd.n3246 vdd.n3245 52.4337
R19951 vdd.n3241 vdd.n385 52.4337
R19952 vdd.n3239 vdd.n3238 52.4337
R19953 vdd.n3234 vdd.n392 52.4337
R19954 vdd.n3232 vdd.n3231 52.4337
R19955 vdd.n3227 vdd.n399 52.4337
R19956 vdd.n3225 vdd.n3224 52.4337
R19957 vdd.n408 vdd.n407 52.4337
R19958 vdd.n3216 vdd.n412 52.4337
R19959 vdd.n3214 vdd.n3213 52.4337
R19960 vdd.n3209 vdd.n418 52.4337
R19961 vdd.n3207 vdd.n3206 52.4337
R19962 vdd.n3202 vdd.n425 52.4337
R19963 vdd.n3200 vdd.n3199 52.4337
R19964 vdd.n3195 vdd.n432 52.4337
R19965 vdd.n3193 vdd.n3192 52.4337
R19966 vdd.n3188 vdd.n439 52.4337
R19967 vdd.n3186 vdd.n3185 52.4337
R19968 vdd.n3178 vdd.n3177 52.4337
R19969 vdd.n3114 vdd.n3113 52.4337
R19970 vdd.n517 vdd.n485 52.4337
R19971 vdd.n523 vdd.n486 52.4337
R19972 vdd.n3103 vdd.n487 52.4337
R19973 vdd.n3099 vdd.n488 52.4337
R19974 vdd.n3095 vdd.n489 52.4337
R19975 vdd.n3091 vdd.n490 52.4337
R19976 vdd.n3087 vdd.n491 52.4337
R19977 vdd.n3083 vdd.n492 52.4337
R19978 vdd.n3079 vdd.n493 52.4337
R19979 vdd.n3071 vdd.n494 52.4337
R19980 vdd.n3067 vdd.n495 52.4337
R19981 vdd.n3063 vdd.n496 52.4337
R19982 vdd.n3059 vdd.n497 52.4337
R19983 vdd.n3055 vdd.n498 52.4337
R19984 vdd.n3051 vdd.n499 52.4337
R19985 vdd.n3047 vdd.n500 52.4337
R19986 vdd.n3043 vdd.n501 52.4337
R19987 vdd.n3039 vdd.n502 52.4337
R19988 vdd.n3035 vdd.n503 52.4337
R19989 vdd.n3031 vdd.n504 52.4337
R19990 vdd.n3025 vdd.n505 52.4337
R19991 vdd.n3021 vdd.n506 52.4337
R19992 vdd.n3017 vdd.n507 52.4337
R19993 vdd.n3013 vdd.n508 52.4337
R19994 vdd.n3009 vdd.n509 52.4337
R19995 vdd.n3005 vdd.n510 52.4337
R19996 vdd.n3001 vdd.n511 52.4337
R19997 vdd.n2997 vdd.n512 52.4337
R19998 vdd.n2993 vdd.n513 52.4337
R19999 vdd.n2989 vdd.n514 52.4337
R20000 vdd.n2085 vdd.n974 52.4337
R20001 vdd.n2083 vdd.n2082 52.4337
R20002 vdd.n2078 vdd.n2077 52.4337
R20003 vdd.n2073 vdd.n978 52.4337
R20004 vdd.n2071 vdd.n2070 52.4337
R20005 vdd.n2066 vdd.n985 52.4337
R20006 vdd.n2064 vdd.n2063 52.4337
R20007 vdd.n2059 vdd.n992 52.4337
R20008 vdd.n2057 vdd.n2056 52.4337
R20009 vdd.n1001 vdd.n1000 52.4337
R20010 vdd.n2048 vdd.n1005 52.4337
R20011 vdd.n2046 vdd.n2045 52.4337
R20012 vdd.n2041 vdd.n1011 52.4337
R20013 vdd.n2039 vdd.n2038 52.4337
R20014 vdd.n2034 vdd.n1018 52.4337
R20015 vdd.n2032 vdd.n2031 52.4337
R20016 vdd.n2027 vdd.n1025 52.4337
R20017 vdd.n2025 vdd.n2024 52.4337
R20018 vdd.n2020 vdd.n1032 52.4337
R20019 vdd.n2018 vdd.n2017 52.4337
R20020 vdd.n1041 vdd.n1040 52.4337
R20021 vdd.n2009 vdd.n1045 52.4337
R20022 vdd.n2007 vdd.n2006 52.4337
R20023 vdd.n2002 vdd.n1051 52.4337
R20024 vdd.n2000 vdd.n1999 52.4337
R20025 vdd.n1995 vdd.n1058 52.4337
R20026 vdd.n1993 vdd.n1992 52.4337
R20027 vdd.n1988 vdd.n1065 52.4337
R20028 vdd.n1986 vdd.n1985 52.4337
R20029 vdd.n1310 vdd.n1309 52.4337
R20030 vdd.n1314 vdd.n1313 52.4337
R20031 vdd.n1974 vdd.n1316 52.4337
R20032 vdd.n1878 vdd.n1877 52.4337
R20033 vdd.n1684 vdd.n1652 52.4337
R20034 vdd.n1688 vdd.n1653 52.4337
R20035 vdd.n1690 vdd.n1654 52.4337
R20036 vdd.n1694 vdd.n1655 52.4337
R20037 vdd.n1696 vdd.n1656 52.4337
R20038 vdd.n1700 vdd.n1657 52.4337
R20039 vdd.n1702 vdd.n1658 52.4337
R20040 vdd.n1706 vdd.n1659 52.4337
R20041 vdd.n1708 vdd.n1660 52.4337
R20042 vdd.n1714 vdd.n1661 52.4337
R20043 vdd.n1716 vdd.n1662 52.4337
R20044 vdd.n1720 vdd.n1663 52.4337
R20045 vdd.n1722 vdd.n1664 52.4337
R20046 vdd.n1726 vdd.n1665 52.4337
R20047 vdd.n1728 vdd.n1666 52.4337
R20048 vdd.n1732 vdd.n1667 52.4337
R20049 vdd.n1734 vdd.n1668 52.4337
R20050 vdd.n1738 vdd.n1669 52.4337
R20051 vdd.n1740 vdd.n1670 52.4337
R20052 vdd.n1812 vdd.n1671 52.4337
R20053 vdd.n1745 vdd.n1672 52.4337
R20054 vdd.n1749 vdd.n1673 52.4337
R20055 vdd.n1751 vdd.n1674 52.4337
R20056 vdd.n1755 vdd.n1675 52.4337
R20057 vdd.n1757 vdd.n1676 52.4337
R20058 vdd.n1761 vdd.n1677 52.4337
R20059 vdd.n1763 vdd.n1678 52.4337
R20060 vdd.n1767 vdd.n1679 52.4337
R20061 vdd.n1769 vdd.n1680 52.4337
R20062 vdd.n1773 vdd.n1681 52.4337
R20063 vdd.n1877 vdd.n1651 52.4337
R20064 vdd.n1687 vdd.n1652 52.4337
R20065 vdd.n1689 vdd.n1653 52.4337
R20066 vdd.n1693 vdd.n1654 52.4337
R20067 vdd.n1695 vdd.n1655 52.4337
R20068 vdd.n1699 vdd.n1656 52.4337
R20069 vdd.n1701 vdd.n1657 52.4337
R20070 vdd.n1705 vdd.n1658 52.4337
R20071 vdd.n1707 vdd.n1659 52.4337
R20072 vdd.n1713 vdd.n1660 52.4337
R20073 vdd.n1715 vdd.n1661 52.4337
R20074 vdd.n1719 vdd.n1662 52.4337
R20075 vdd.n1721 vdd.n1663 52.4337
R20076 vdd.n1725 vdd.n1664 52.4337
R20077 vdd.n1727 vdd.n1665 52.4337
R20078 vdd.n1731 vdd.n1666 52.4337
R20079 vdd.n1733 vdd.n1667 52.4337
R20080 vdd.n1737 vdd.n1668 52.4337
R20081 vdd.n1739 vdd.n1669 52.4337
R20082 vdd.n1743 vdd.n1670 52.4337
R20083 vdd.n1744 vdd.n1671 52.4337
R20084 vdd.n1748 vdd.n1672 52.4337
R20085 vdd.n1750 vdd.n1673 52.4337
R20086 vdd.n1754 vdd.n1674 52.4337
R20087 vdd.n1756 vdd.n1675 52.4337
R20088 vdd.n1760 vdd.n1676 52.4337
R20089 vdd.n1762 vdd.n1677 52.4337
R20090 vdd.n1766 vdd.n1678 52.4337
R20091 vdd.n1768 vdd.n1679 52.4337
R20092 vdd.n1772 vdd.n1680 52.4337
R20093 vdd.n1774 vdd.n1681 52.4337
R20094 vdd.n1316 vdd.n1315 52.4337
R20095 vdd.n1313 vdd.n1312 52.4337
R20096 vdd.n1309 vdd.n1066 52.4337
R20097 vdd.n1987 vdd.n1986 52.4337
R20098 vdd.n1065 vdd.n1059 52.4337
R20099 vdd.n1994 vdd.n1993 52.4337
R20100 vdd.n1058 vdd.n1052 52.4337
R20101 vdd.n2001 vdd.n2000 52.4337
R20102 vdd.n1051 vdd.n1046 52.4337
R20103 vdd.n2008 vdd.n2007 52.4337
R20104 vdd.n1045 vdd.n1044 52.4337
R20105 vdd.n1040 vdd.n1033 52.4337
R20106 vdd.n2019 vdd.n2018 52.4337
R20107 vdd.n1032 vdd.n1026 52.4337
R20108 vdd.n2026 vdd.n2025 52.4337
R20109 vdd.n1025 vdd.n1019 52.4337
R20110 vdd.n2033 vdd.n2032 52.4337
R20111 vdd.n1018 vdd.n1012 52.4337
R20112 vdd.n2040 vdd.n2039 52.4337
R20113 vdd.n1011 vdd.n1006 52.4337
R20114 vdd.n2047 vdd.n2046 52.4337
R20115 vdd.n1005 vdd.n1004 52.4337
R20116 vdd.n1000 vdd.n993 52.4337
R20117 vdd.n2058 vdd.n2057 52.4337
R20118 vdd.n992 vdd.n986 52.4337
R20119 vdd.n2065 vdd.n2064 52.4337
R20120 vdd.n985 vdd.n979 52.4337
R20121 vdd.n2072 vdd.n2071 52.4337
R20122 vdd.n978 vdd.n975 52.4337
R20123 vdd.n2079 vdd.n2078 52.4337
R20124 vdd.n2084 vdd.n2083 52.4337
R20125 vdd.n1320 vdd.n974 52.4337
R20126 vdd.n3113 vdd.n483 52.4337
R20127 vdd.n522 vdd.n485 52.4337
R20128 vdd.n3104 vdd.n486 52.4337
R20129 vdd.n3100 vdd.n487 52.4337
R20130 vdd.n3096 vdd.n488 52.4337
R20131 vdd.n3092 vdd.n489 52.4337
R20132 vdd.n3088 vdd.n490 52.4337
R20133 vdd.n3084 vdd.n491 52.4337
R20134 vdd.n3080 vdd.n492 52.4337
R20135 vdd.n3070 vdd.n493 52.4337
R20136 vdd.n3068 vdd.n494 52.4337
R20137 vdd.n3064 vdd.n495 52.4337
R20138 vdd.n3060 vdd.n496 52.4337
R20139 vdd.n3056 vdd.n497 52.4337
R20140 vdd.n3052 vdd.n498 52.4337
R20141 vdd.n3048 vdd.n499 52.4337
R20142 vdd.n3044 vdd.n500 52.4337
R20143 vdd.n3040 vdd.n501 52.4337
R20144 vdd.n3036 vdd.n502 52.4337
R20145 vdd.n3032 vdd.n503 52.4337
R20146 vdd.n3024 vdd.n504 52.4337
R20147 vdd.n3022 vdd.n505 52.4337
R20148 vdd.n3018 vdd.n506 52.4337
R20149 vdd.n3014 vdd.n507 52.4337
R20150 vdd.n3010 vdd.n508 52.4337
R20151 vdd.n3006 vdd.n509 52.4337
R20152 vdd.n3002 vdd.n510 52.4337
R20153 vdd.n2998 vdd.n511 52.4337
R20154 vdd.n2994 vdd.n512 52.4337
R20155 vdd.n2990 vdd.n513 52.4337
R20156 vdd.n2986 vdd.n514 52.4337
R20157 vdd.n3177 vdd.n440 52.4337
R20158 vdd.n3187 vdd.n3186 52.4337
R20159 vdd.n439 vdd.n433 52.4337
R20160 vdd.n3194 vdd.n3193 52.4337
R20161 vdd.n432 vdd.n426 52.4337
R20162 vdd.n3201 vdd.n3200 52.4337
R20163 vdd.n425 vdd.n419 52.4337
R20164 vdd.n3208 vdd.n3207 52.4337
R20165 vdd.n418 vdd.n413 52.4337
R20166 vdd.n3215 vdd.n3214 52.4337
R20167 vdd.n412 vdd.n411 52.4337
R20168 vdd.n407 vdd.n400 52.4337
R20169 vdd.n3226 vdd.n3225 52.4337
R20170 vdd.n399 vdd.n393 52.4337
R20171 vdd.n3233 vdd.n3232 52.4337
R20172 vdd.n392 vdd.n386 52.4337
R20173 vdd.n3240 vdd.n3239 52.4337
R20174 vdd.n385 vdd.n379 52.4337
R20175 vdd.n3247 vdd.n3246 52.4337
R20176 vdd.n378 vdd.n373 52.4337
R20177 vdd.n3254 vdd.n3253 52.4337
R20178 vdd.n372 vdd.n371 52.4337
R20179 vdd.n367 vdd.n360 52.4337
R20180 vdd.n3265 vdd.n3264 52.4337
R20181 vdd.n359 vdd.n353 52.4337
R20182 vdd.n3272 vdd.n3271 52.4337
R20183 vdd.n352 vdd.n346 52.4337
R20184 vdd.n3279 vdd.n3278 52.4337
R20185 vdd.n345 vdd.n338 52.4337
R20186 vdd.n3286 vdd.n3285 52.4337
R20187 vdd.n3289 vdd.n3288 52.4337
R20188 vdd.n333 vdd.n330 52.4337
R20189 vdd.t20 vdd.t33 51.4683
R20190 vdd.n250 vdd.n248 42.0461
R20191 vdd.n160 vdd.n158 42.0461
R20192 vdd.n71 vdd.n69 42.0461
R20193 vdd.n1567 vdd.n1565 42.0461
R20194 vdd.n1477 vdd.n1475 42.0461
R20195 vdd.n1388 vdd.n1386 42.0461
R20196 vdd.n296 vdd.n295 41.6884
R20197 vdd.n206 vdd.n205 41.6884
R20198 vdd.n117 vdd.n116 41.6884
R20199 vdd.n1613 vdd.n1612 41.6884
R20200 vdd.n1523 vdd.n1522 41.6884
R20201 vdd.n1434 vdd.n1433 41.6884
R20202 vdd.n1777 vdd.n1776 41.1157
R20203 vdd.n1815 vdd.n1814 41.1157
R20204 vdd.n1711 vdd.n1710 41.1157
R20205 vdd.n3182 vdd.n3181 41.1157
R20206 vdd.n3221 vdd.n406 41.1157
R20207 vdd.n3260 vdd.n366 41.1157
R20208 vdd.n2939 vdd.n2938 39.2114
R20209 vdd.n2936 vdd.n2935 39.2114
R20210 vdd.n2931 vdd.n605 39.2114
R20211 vdd.n2929 vdd.n2928 39.2114
R20212 vdd.n2924 vdd.n608 39.2114
R20213 vdd.n2922 vdd.n2921 39.2114
R20214 vdd.n2917 vdd.n611 39.2114
R20215 vdd.n2915 vdd.n2914 39.2114
R20216 vdd.n2911 vdd.n2910 39.2114
R20217 vdd.n2906 vdd.n614 39.2114
R20218 vdd.n2904 vdd.n2903 39.2114
R20219 vdd.n2899 vdd.n617 39.2114
R20220 vdd.n2897 vdd.n2896 39.2114
R20221 vdd.n2892 vdd.n620 39.2114
R20222 vdd.n2890 vdd.n2889 39.2114
R20223 vdd.n2884 vdd.n625 39.2114
R20224 vdd.n2882 vdd.n2881 39.2114
R20225 vdd.n2704 vdd.n2703 39.2114
R20226 vdd.n2433 vdd.n2399 39.2114
R20227 vdd.n2696 vdd.n2400 39.2114
R20228 vdd.n2692 vdd.n2401 39.2114
R20229 vdd.n2688 vdd.n2402 39.2114
R20230 vdd.n2684 vdd.n2403 39.2114
R20231 vdd.n2680 vdd.n2404 39.2114
R20232 vdd.n2676 vdd.n2405 39.2114
R20233 vdd.n2672 vdd.n2406 39.2114
R20234 vdd.n2668 vdd.n2407 39.2114
R20235 vdd.n2664 vdd.n2408 39.2114
R20236 vdd.n2660 vdd.n2409 39.2114
R20237 vdd.n2656 vdd.n2410 39.2114
R20238 vdd.n2652 vdd.n2411 39.2114
R20239 vdd.n2648 vdd.n2412 39.2114
R20240 vdd.n2644 vdd.n2413 39.2114
R20241 vdd.n2639 vdd.n2414 39.2114
R20242 vdd.n2393 vdd.n787 39.2114
R20243 vdd.n2389 vdd.n786 39.2114
R20244 vdd.n2385 vdd.n785 39.2114
R20245 vdd.n2381 vdd.n784 39.2114
R20246 vdd.n2377 vdd.n783 39.2114
R20247 vdd.n2373 vdd.n782 39.2114
R20248 vdd.n2369 vdd.n781 39.2114
R20249 vdd.n2365 vdd.n780 39.2114
R20250 vdd.n2361 vdd.n779 39.2114
R20251 vdd.n2357 vdd.n778 39.2114
R20252 vdd.n2353 vdd.n777 39.2114
R20253 vdd.n2349 vdd.n776 39.2114
R20254 vdd.n2345 vdd.n775 39.2114
R20255 vdd.n2341 vdd.n774 39.2114
R20256 vdd.n2337 vdd.n773 39.2114
R20257 vdd.n2332 vdd.n772 39.2114
R20258 vdd.n2328 vdd.n771 39.2114
R20259 vdd.n2122 vdd.n2121 39.2114
R20260 vdd.n966 vdd.n932 39.2114
R20261 vdd.n2114 vdd.n933 39.2114
R20262 vdd.n2110 vdd.n934 39.2114
R20263 vdd.n2106 vdd.n935 39.2114
R20264 vdd.n2102 vdd.n936 39.2114
R20265 vdd.n2098 vdd.n937 39.2114
R20266 vdd.n2094 vdd.n938 39.2114
R20267 vdd.n2090 vdd.n939 39.2114
R20268 vdd.n1112 vdd.n940 39.2114
R20269 vdd.n1116 vdd.n941 39.2114
R20270 vdd.n1120 vdd.n942 39.2114
R20271 vdd.n1124 vdd.n943 39.2114
R20272 vdd.n1128 vdd.n944 39.2114
R20273 vdd.n1132 vdd.n945 39.2114
R20274 vdd.n1136 vdd.n946 39.2114
R20275 vdd.n1141 vdd.n947 39.2114
R20276 vdd.n2858 vdd.n2857 39.2114
R20277 vdd.n2853 vdd.n2825 39.2114
R20278 vdd.n2851 vdd.n2850 39.2114
R20279 vdd.n2846 vdd.n2828 39.2114
R20280 vdd.n2844 vdd.n2843 39.2114
R20281 vdd.n2839 vdd.n2831 39.2114
R20282 vdd.n2837 vdd.n2836 39.2114
R20283 vdd.n2832 vdd.n577 39.2114
R20284 vdd.n2976 vdd.n2975 39.2114
R20285 vdd.n2973 vdd.n2972 39.2114
R20286 vdd.n2968 vdd.n581 39.2114
R20287 vdd.n2966 vdd.n2965 39.2114
R20288 vdd.n2961 vdd.n584 39.2114
R20289 vdd.n2959 vdd.n2958 39.2114
R20290 vdd.n2954 vdd.n587 39.2114
R20291 vdd.n2952 vdd.n2951 39.2114
R20292 vdd.n2947 vdd.n593 39.2114
R20293 vdd.n2440 vdd.n2415 39.2114
R20294 vdd.n2444 vdd.n2416 39.2114
R20295 vdd.n2448 vdd.n2417 39.2114
R20296 vdd.n2452 vdd.n2418 39.2114
R20297 vdd.n2456 vdd.n2419 39.2114
R20298 vdd.n2460 vdd.n2420 39.2114
R20299 vdd.n2464 vdd.n2421 39.2114
R20300 vdd.n2468 vdd.n2422 39.2114
R20301 vdd.n2472 vdd.n2423 39.2114
R20302 vdd.n2476 vdd.n2424 39.2114
R20303 vdd.n2480 vdd.n2425 39.2114
R20304 vdd.n2484 vdd.n2426 39.2114
R20305 vdd.n2488 vdd.n2427 39.2114
R20306 vdd.n2492 vdd.n2428 39.2114
R20307 vdd.n2496 vdd.n2429 39.2114
R20308 vdd.n2500 vdd.n2430 39.2114
R20309 vdd.n2504 vdd.n2431 39.2114
R20310 vdd.n2443 vdd.n2415 39.2114
R20311 vdd.n2447 vdd.n2416 39.2114
R20312 vdd.n2451 vdd.n2417 39.2114
R20313 vdd.n2455 vdd.n2418 39.2114
R20314 vdd.n2459 vdd.n2419 39.2114
R20315 vdd.n2463 vdd.n2420 39.2114
R20316 vdd.n2467 vdd.n2421 39.2114
R20317 vdd.n2471 vdd.n2422 39.2114
R20318 vdd.n2475 vdd.n2423 39.2114
R20319 vdd.n2479 vdd.n2424 39.2114
R20320 vdd.n2483 vdd.n2425 39.2114
R20321 vdd.n2487 vdd.n2426 39.2114
R20322 vdd.n2491 vdd.n2427 39.2114
R20323 vdd.n2495 vdd.n2428 39.2114
R20324 vdd.n2499 vdd.n2429 39.2114
R20325 vdd.n2503 vdd.n2430 39.2114
R20326 vdd.n2506 vdd.n2431 39.2114
R20327 vdd.n593 vdd.n588 39.2114
R20328 vdd.n2953 vdd.n2952 39.2114
R20329 vdd.n587 vdd.n585 39.2114
R20330 vdd.n2960 vdd.n2959 39.2114
R20331 vdd.n584 vdd.n582 39.2114
R20332 vdd.n2967 vdd.n2966 39.2114
R20333 vdd.n581 vdd.n579 39.2114
R20334 vdd.n2974 vdd.n2973 39.2114
R20335 vdd.n2977 vdd.n2976 39.2114
R20336 vdd.n2833 vdd.n2832 39.2114
R20337 vdd.n2838 vdd.n2837 39.2114
R20338 vdd.n2831 vdd.n2829 39.2114
R20339 vdd.n2845 vdd.n2844 39.2114
R20340 vdd.n2828 vdd.n2826 39.2114
R20341 vdd.n2852 vdd.n2851 39.2114
R20342 vdd.n2825 vdd.n2823 39.2114
R20343 vdd.n2859 vdd.n2858 39.2114
R20344 vdd.n2121 vdd.n930 39.2114
R20345 vdd.n2115 vdd.n932 39.2114
R20346 vdd.n2111 vdd.n933 39.2114
R20347 vdd.n2107 vdd.n934 39.2114
R20348 vdd.n2103 vdd.n935 39.2114
R20349 vdd.n2099 vdd.n936 39.2114
R20350 vdd.n2095 vdd.n937 39.2114
R20351 vdd.n2091 vdd.n938 39.2114
R20352 vdd.n1111 vdd.n939 39.2114
R20353 vdd.n1115 vdd.n940 39.2114
R20354 vdd.n1119 vdd.n941 39.2114
R20355 vdd.n1123 vdd.n942 39.2114
R20356 vdd.n1127 vdd.n943 39.2114
R20357 vdd.n1131 vdd.n944 39.2114
R20358 vdd.n1135 vdd.n945 39.2114
R20359 vdd.n1140 vdd.n946 39.2114
R20360 vdd.n1144 vdd.n947 39.2114
R20361 vdd.n2331 vdd.n771 39.2114
R20362 vdd.n2336 vdd.n772 39.2114
R20363 vdd.n2340 vdd.n773 39.2114
R20364 vdd.n2344 vdd.n774 39.2114
R20365 vdd.n2348 vdd.n775 39.2114
R20366 vdd.n2352 vdd.n776 39.2114
R20367 vdd.n2356 vdd.n777 39.2114
R20368 vdd.n2360 vdd.n778 39.2114
R20369 vdd.n2364 vdd.n779 39.2114
R20370 vdd.n2368 vdd.n780 39.2114
R20371 vdd.n2372 vdd.n781 39.2114
R20372 vdd.n2376 vdd.n782 39.2114
R20373 vdd.n2380 vdd.n783 39.2114
R20374 vdd.n2384 vdd.n784 39.2114
R20375 vdd.n2388 vdd.n785 39.2114
R20376 vdd.n2392 vdd.n786 39.2114
R20377 vdd.n789 vdd.n787 39.2114
R20378 vdd.n2703 vdd.n752 39.2114
R20379 vdd.n2697 vdd.n2399 39.2114
R20380 vdd.n2693 vdd.n2400 39.2114
R20381 vdd.n2689 vdd.n2401 39.2114
R20382 vdd.n2685 vdd.n2402 39.2114
R20383 vdd.n2681 vdd.n2403 39.2114
R20384 vdd.n2677 vdd.n2404 39.2114
R20385 vdd.n2673 vdd.n2405 39.2114
R20386 vdd.n2669 vdd.n2406 39.2114
R20387 vdd.n2665 vdd.n2407 39.2114
R20388 vdd.n2661 vdd.n2408 39.2114
R20389 vdd.n2657 vdd.n2409 39.2114
R20390 vdd.n2653 vdd.n2410 39.2114
R20391 vdd.n2649 vdd.n2411 39.2114
R20392 vdd.n2645 vdd.n2412 39.2114
R20393 vdd.n2640 vdd.n2413 39.2114
R20394 vdd.n2636 vdd.n2414 39.2114
R20395 vdd.n2883 vdd.n2882 39.2114
R20396 vdd.n625 vdd.n621 39.2114
R20397 vdd.n2891 vdd.n2890 39.2114
R20398 vdd.n620 vdd.n618 39.2114
R20399 vdd.n2898 vdd.n2897 39.2114
R20400 vdd.n617 vdd.n615 39.2114
R20401 vdd.n2905 vdd.n2904 39.2114
R20402 vdd.n614 vdd.n612 39.2114
R20403 vdd.n2912 vdd.n2911 39.2114
R20404 vdd.n2916 vdd.n2915 39.2114
R20405 vdd.n611 vdd.n609 39.2114
R20406 vdd.n2923 vdd.n2922 39.2114
R20407 vdd.n608 vdd.n606 39.2114
R20408 vdd.n2930 vdd.n2929 39.2114
R20409 vdd.n605 vdd.n603 39.2114
R20410 vdd.n2937 vdd.n2936 39.2114
R20411 vdd.n2940 vdd.n2939 39.2114
R20412 vdd.n798 vdd.n753 39.2114
R20413 vdd.n2320 vdd.n754 39.2114
R20414 vdd.n2316 vdd.n755 39.2114
R20415 vdd.n2312 vdd.n756 39.2114
R20416 vdd.n2308 vdd.n757 39.2114
R20417 vdd.n2304 vdd.n758 39.2114
R20418 vdd.n2300 vdd.n759 39.2114
R20419 vdd.n2296 vdd.n760 39.2114
R20420 vdd.n2292 vdd.n761 39.2114
R20421 vdd.n2288 vdd.n762 39.2114
R20422 vdd.n2284 vdd.n763 39.2114
R20423 vdd.n2280 vdd.n764 39.2114
R20424 vdd.n2276 vdd.n765 39.2114
R20425 vdd.n2272 vdd.n766 39.2114
R20426 vdd.n2268 vdd.n767 39.2114
R20427 vdd.n2264 vdd.n768 39.2114
R20428 vdd.n2260 vdd.n769 39.2114
R20429 vdd.n1070 vdd.n948 39.2114
R20430 vdd.n1074 vdd.n949 39.2114
R20431 vdd.n1078 vdd.n950 39.2114
R20432 vdd.n1082 vdd.n951 39.2114
R20433 vdd.n1086 vdd.n952 39.2114
R20434 vdd.n1090 vdd.n953 39.2114
R20435 vdd.n1094 vdd.n954 39.2114
R20436 vdd.n1098 vdd.n955 39.2114
R20437 vdd.n1102 vdd.n956 39.2114
R20438 vdd.n1303 vdd.n957 39.2114
R20439 vdd.n1300 vdd.n958 39.2114
R20440 vdd.n1296 vdd.n959 39.2114
R20441 vdd.n1292 vdd.n960 39.2114
R20442 vdd.n1288 vdd.n961 39.2114
R20443 vdd.n1284 vdd.n962 39.2114
R20444 vdd.n1280 vdd.n963 39.2114
R20445 vdd.n1276 vdd.n964 39.2114
R20446 vdd.n2257 vdd.n769 39.2114
R20447 vdd.n2261 vdd.n768 39.2114
R20448 vdd.n2265 vdd.n767 39.2114
R20449 vdd.n2269 vdd.n766 39.2114
R20450 vdd.n2273 vdd.n765 39.2114
R20451 vdd.n2277 vdd.n764 39.2114
R20452 vdd.n2281 vdd.n763 39.2114
R20453 vdd.n2285 vdd.n762 39.2114
R20454 vdd.n2289 vdd.n761 39.2114
R20455 vdd.n2293 vdd.n760 39.2114
R20456 vdd.n2297 vdd.n759 39.2114
R20457 vdd.n2301 vdd.n758 39.2114
R20458 vdd.n2305 vdd.n757 39.2114
R20459 vdd.n2309 vdd.n756 39.2114
R20460 vdd.n2313 vdd.n755 39.2114
R20461 vdd.n2317 vdd.n754 39.2114
R20462 vdd.n2321 vdd.n753 39.2114
R20463 vdd.n1073 vdd.n948 39.2114
R20464 vdd.n1077 vdd.n949 39.2114
R20465 vdd.n1081 vdd.n950 39.2114
R20466 vdd.n1085 vdd.n951 39.2114
R20467 vdd.n1089 vdd.n952 39.2114
R20468 vdd.n1093 vdd.n953 39.2114
R20469 vdd.n1097 vdd.n954 39.2114
R20470 vdd.n1101 vdd.n955 39.2114
R20471 vdd.n1104 vdd.n956 39.2114
R20472 vdd.n1301 vdd.n957 39.2114
R20473 vdd.n1297 vdd.n958 39.2114
R20474 vdd.n1293 vdd.n959 39.2114
R20475 vdd.n1289 vdd.n960 39.2114
R20476 vdd.n1285 vdd.n961 39.2114
R20477 vdd.n1281 vdd.n962 39.2114
R20478 vdd.n1277 vdd.n963 39.2114
R20479 vdd.n1273 vdd.n964 39.2114
R20480 vdd.n1978 vdd.n1977 37.2369
R20481 vdd.n2014 vdd.n1039 37.2369
R20482 vdd.n2053 vdd.n999 37.2369
R20483 vdd.n3030 vdd.n558 37.2369
R20484 vdd.n3078 vdd.n3077 37.2369
R20485 vdd.n2985 vdd.n2984 37.2369
R20486 vdd.n1107 vdd.n1106 30.449
R20487 vdd.n802 vdd.n801 30.449
R20488 vdd.n1138 vdd.n1110 30.449
R20489 vdd.n2334 vdd.n792 30.449
R20490 vdd.n2439 vdd.n2438 30.449
R20491 vdd.n2886 vdd.n623 30.449
R20492 vdd.n2642 vdd.n2435 30.449
R20493 vdd.n591 vdd.n590 30.449
R20494 vdd.n2124 vdd.n2123 29.8151
R20495 vdd.n2396 vdd.n790 29.8151
R20496 vdd.n2329 vdd.n793 29.8151
R20497 vdd.n1146 vdd.n1143 29.8151
R20498 vdd.n2637 vdd.n2634 29.8151
R20499 vdd.n2880 vdd.n2879 29.8151
R20500 vdd.n2706 vdd.n2705 29.8151
R20501 vdd.n2943 vdd.n2942 29.8151
R20502 vdd.n2862 vdd.n2861 29.8151
R20503 vdd.n2948 vdd.n592 29.8151
R20504 vdd.n2510 vdd.n2508 29.8151
R20505 vdd.n2441 vdd.n745 29.8151
R20506 vdd.n1071 vdd.n922 29.8151
R20507 vdd.n2324 vdd.n2323 29.8151
R20508 vdd.n2256 vdd.n2255 29.8151
R20509 vdd.n1272 vdd.n1271 29.8151
R20510 vdd.n1876 vdd.n1683 22.6735
R20511 vdd.n1972 vdd.n931 22.6735
R20512 vdd.n3112 vdd.n516 22.6735
R20513 vdd.n3297 vdd.n329 22.6735
R20514 vdd.n1887 vdd.n1645 19.3944
R20515 vdd.n1887 vdd.n1643 19.3944
R20516 vdd.n1891 vdd.n1643 19.3944
R20517 vdd.n1891 vdd.n1633 19.3944
R20518 vdd.n1904 vdd.n1633 19.3944
R20519 vdd.n1904 vdd.n1631 19.3944
R20520 vdd.n1908 vdd.n1631 19.3944
R20521 vdd.n1908 vdd.n1623 19.3944
R20522 vdd.n1922 vdd.n1623 19.3944
R20523 vdd.n1922 vdd.n1621 19.3944
R20524 vdd.n1926 vdd.n1621 19.3944
R20525 vdd.n1926 vdd.n1340 19.3944
R20526 vdd.n1938 vdd.n1340 19.3944
R20527 vdd.n1938 vdd.n1338 19.3944
R20528 vdd.n1942 vdd.n1338 19.3944
R20529 vdd.n1942 vdd.n1330 19.3944
R20530 vdd.n1955 vdd.n1330 19.3944
R20531 vdd.n1955 vdd.n1327 19.3944
R20532 vdd.n1961 vdd.n1327 19.3944
R20533 vdd.n1961 vdd.n1328 19.3944
R20534 vdd.n1328 vdd.n1318 19.3944
R20535 vdd.n1811 vdd.n1746 19.3944
R20536 vdd.n1807 vdd.n1746 19.3944
R20537 vdd.n1807 vdd.n1806 19.3944
R20538 vdd.n1806 vdd.n1805 19.3944
R20539 vdd.n1805 vdd.n1752 19.3944
R20540 vdd.n1801 vdd.n1752 19.3944
R20541 vdd.n1801 vdd.n1800 19.3944
R20542 vdd.n1800 vdd.n1799 19.3944
R20543 vdd.n1799 vdd.n1758 19.3944
R20544 vdd.n1795 vdd.n1758 19.3944
R20545 vdd.n1795 vdd.n1794 19.3944
R20546 vdd.n1794 vdd.n1793 19.3944
R20547 vdd.n1793 vdd.n1764 19.3944
R20548 vdd.n1789 vdd.n1764 19.3944
R20549 vdd.n1789 vdd.n1788 19.3944
R20550 vdd.n1788 vdd.n1787 19.3944
R20551 vdd.n1787 vdd.n1770 19.3944
R20552 vdd.n1783 vdd.n1770 19.3944
R20553 vdd.n1783 vdd.n1782 19.3944
R20554 vdd.n1782 vdd.n1781 19.3944
R20555 vdd.n1846 vdd.n1845 19.3944
R20556 vdd.n1845 vdd.n1844 19.3944
R20557 vdd.n1844 vdd.n1717 19.3944
R20558 vdd.n1840 vdd.n1717 19.3944
R20559 vdd.n1840 vdd.n1839 19.3944
R20560 vdd.n1839 vdd.n1838 19.3944
R20561 vdd.n1838 vdd.n1723 19.3944
R20562 vdd.n1834 vdd.n1723 19.3944
R20563 vdd.n1834 vdd.n1833 19.3944
R20564 vdd.n1833 vdd.n1832 19.3944
R20565 vdd.n1832 vdd.n1729 19.3944
R20566 vdd.n1828 vdd.n1729 19.3944
R20567 vdd.n1828 vdd.n1827 19.3944
R20568 vdd.n1827 vdd.n1826 19.3944
R20569 vdd.n1826 vdd.n1735 19.3944
R20570 vdd.n1822 vdd.n1735 19.3944
R20571 vdd.n1822 vdd.n1821 19.3944
R20572 vdd.n1821 vdd.n1820 19.3944
R20573 vdd.n1820 vdd.n1741 19.3944
R20574 vdd.n1816 vdd.n1741 19.3944
R20575 vdd.n1879 vdd.n1650 19.3944
R20576 vdd.n1874 vdd.n1650 19.3944
R20577 vdd.n1874 vdd.n1685 19.3944
R20578 vdd.n1870 vdd.n1685 19.3944
R20579 vdd.n1870 vdd.n1869 19.3944
R20580 vdd.n1869 vdd.n1868 19.3944
R20581 vdd.n1868 vdd.n1691 19.3944
R20582 vdd.n1864 vdd.n1691 19.3944
R20583 vdd.n1864 vdd.n1863 19.3944
R20584 vdd.n1863 vdd.n1862 19.3944
R20585 vdd.n1862 vdd.n1697 19.3944
R20586 vdd.n1858 vdd.n1697 19.3944
R20587 vdd.n1858 vdd.n1857 19.3944
R20588 vdd.n1857 vdd.n1856 19.3944
R20589 vdd.n1856 vdd.n1703 19.3944
R20590 vdd.n1852 vdd.n1703 19.3944
R20591 vdd.n1852 vdd.n1851 19.3944
R20592 vdd.n1851 vdd.n1850 19.3944
R20593 vdd.n2010 vdd.n1037 19.3944
R20594 vdd.n2010 vdd.n1043 19.3944
R20595 vdd.n2005 vdd.n1043 19.3944
R20596 vdd.n2005 vdd.n2004 19.3944
R20597 vdd.n2004 vdd.n2003 19.3944
R20598 vdd.n2003 vdd.n1050 19.3944
R20599 vdd.n1998 vdd.n1050 19.3944
R20600 vdd.n1998 vdd.n1997 19.3944
R20601 vdd.n1997 vdd.n1996 19.3944
R20602 vdd.n1996 vdd.n1057 19.3944
R20603 vdd.n1991 vdd.n1057 19.3944
R20604 vdd.n1991 vdd.n1990 19.3944
R20605 vdd.n1990 vdd.n1989 19.3944
R20606 vdd.n1989 vdd.n1064 19.3944
R20607 vdd.n1984 vdd.n1064 19.3944
R20608 vdd.n1984 vdd.n1983 19.3944
R20609 vdd.n1311 vdd.n1069 19.3944
R20610 vdd.n1979 vdd.n1308 19.3944
R20611 vdd.n2049 vdd.n997 19.3944
R20612 vdd.n2049 vdd.n1003 19.3944
R20613 vdd.n2044 vdd.n1003 19.3944
R20614 vdd.n2044 vdd.n2043 19.3944
R20615 vdd.n2043 vdd.n2042 19.3944
R20616 vdd.n2042 vdd.n1010 19.3944
R20617 vdd.n2037 vdd.n1010 19.3944
R20618 vdd.n2037 vdd.n2036 19.3944
R20619 vdd.n2036 vdd.n2035 19.3944
R20620 vdd.n2035 vdd.n1017 19.3944
R20621 vdd.n2030 vdd.n1017 19.3944
R20622 vdd.n2030 vdd.n2029 19.3944
R20623 vdd.n2029 vdd.n2028 19.3944
R20624 vdd.n2028 vdd.n1024 19.3944
R20625 vdd.n2023 vdd.n1024 19.3944
R20626 vdd.n2023 vdd.n2022 19.3944
R20627 vdd.n2022 vdd.n2021 19.3944
R20628 vdd.n2021 vdd.n1031 19.3944
R20629 vdd.n2016 vdd.n1031 19.3944
R20630 vdd.n2016 vdd.n2015 19.3944
R20631 vdd.n2086 vdd.n972 19.3944
R20632 vdd.n2086 vdd.n973 19.3944
R20633 vdd.n2081 vdd.n2080 19.3944
R20634 vdd.n2076 vdd.n2075 19.3944
R20635 vdd.n2075 vdd.n2074 19.3944
R20636 vdd.n2074 vdd.n977 19.3944
R20637 vdd.n2069 vdd.n977 19.3944
R20638 vdd.n2069 vdd.n2068 19.3944
R20639 vdd.n2068 vdd.n2067 19.3944
R20640 vdd.n2067 vdd.n984 19.3944
R20641 vdd.n2062 vdd.n984 19.3944
R20642 vdd.n2062 vdd.n2061 19.3944
R20643 vdd.n2061 vdd.n2060 19.3944
R20644 vdd.n2060 vdd.n991 19.3944
R20645 vdd.n2055 vdd.n991 19.3944
R20646 vdd.n2055 vdd.n2054 19.3944
R20647 vdd.n1883 vdd.n1648 19.3944
R20648 vdd.n1883 vdd.n1639 19.3944
R20649 vdd.n1896 vdd.n1639 19.3944
R20650 vdd.n1896 vdd.n1637 19.3944
R20651 vdd.n1900 vdd.n1637 19.3944
R20652 vdd.n1900 vdd.n1628 19.3944
R20653 vdd.n1913 vdd.n1628 19.3944
R20654 vdd.n1913 vdd.n1626 19.3944
R20655 vdd.n1918 vdd.n1626 19.3944
R20656 vdd.n1918 vdd.n1617 19.3944
R20657 vdd.n1930 vdd.n1617 19.3944
R20658 vdd.n1930 vdd.n1345 19.3944
R20659 vdd.n1934 vdd.n1345 19.3944
R20660 vdd.n1934 vdd.n1335 19.3944
R20661 vdd.n1947 vdd.n1335 19.3944
R20662 vdd.n1947 vdd.n1333 19.3944
R20663 vdd.n1951 vdd.n1333 19.3944
R20664 vdd.n1951 vdd.n1323 19.3944
R20665 vdd.n1966 vdd.n1323 19.3944
R20666 vdd.n1966 vdd.n1321 19.3944
R20667 vdd.n1970 vdd.n1321 19.3944
R20668 vdd.n3123 vdd.n477 19.3944
R20669 vdd.n3123 vdd.n475 19.3944
R20670 vdd.n3127 vdd.n475 19.3944
R20671 vdd.n3127 vdd.n465 19.3944
R20672 vdd.n3140 vdd.n465 19.3944
R20673 vdd.n3140 vdd.n463 19.3944
R20674 vdd.n3144 vdd.n463 19.3944
R20675 vdd.n3144 vdd.n453 19.3944
R20676 vdd.n3156 vdd.n453 19.3944
R20677 vdd.n3156 vdd.n451 19.3944
R20678 vdd.n3160 vdd.n451 19.3944
R20679 vdd.n3161 vdd.n3160 19.3944
R20680 vdd.n3162 vdd.n3161 19.3944
R20681 vdd.n3162 vdd.n449 19.3944
R20682 vdd.n3166 vdd.n449 19.3944
R20683 vdd.n3167 vdd.n3166 19.3944
R20684 vdd.n3168 vdd.n3167 19.3944
R20685 vdd.n3168 vdd.n446 19.3944
R20686 vdd.n3172 vdd.n446 19.3944
R20687 vdd.n3173 vdd.n3172 19.3944
R20688 vdd.n3174 vdd.n3173 19.3944
R20689 vdd.n3217 vdd.n404 19.3944
R20690 vdd.n3217 vdd.n410 19.3944
R20691 vdd.n3212 vdd.n410 19.3944
R20692 vdd.n3212 vdd.n3211 19.3944
R20693 vdd.n3211 vdd.n3210 19.3944
R20694 vdd.n3210 vdd.n417 19.3944
R20695 vdd.n3205 vdd.n417 19.3944
R20696 vdd.n3205 vdd.n3204 19.3944
R20697 vdd.n3204 vdd.n3203 19.3944
R20698 vdd.n3203 vdd.n424 19.3944
R20699 vdd.n3198 vdd.n424 19.3944
R20700 vdd.n3198 vdd.n3197 19.3944
R20701 vdd.n3197 vdd.n3196 19.3944
R20702 vdd.n3196 vdd.n431 19.3944
R20703 vdd.n3191 vdd.n431 19.3944
R20704 vdd.n3191 vdd.n3190 19.3944
R20705 vdd.n3190 vdd.n3189 19.3944
R20706 vdd.n3189 vdd.n438 19.3944
R20707 vdd.n3184 vdd.n438 19.3944
R20708 vdd.n3184 vdd.n3183 19.3944
R20709 vdd.n3256 vdd.n364 19.3944
R20710 vdd.n3256 vdd.n370 19.3944
R20711 vdd.n3251 vdd.n370 19.3944
R20712 vdd.n3251 vdd.n3250 19.3944
R20713 vdd.n3250 vdd.n3249 19.3944
R20714 vdd.n3249 vdd.n377 19.3944
R20715 vdd.n3244 vdd.n377 19.3944
R20716 vdd.n3244 vdd.n3243 19.3944
R20717 vdd.n3243 vdd.n3242 19.3944
R20718 vdd.n3242 vdd.n384 19.3944
R20719 vdd.n3237 vdd.n384 19.3944
R20720 vdd.n3237 vdd.n3236 19.3944
R20721 vdd.n3236 vdd.n3235 19.3944
R20722 vdd.n3235 vdd.n391 19.3944
R20723 vdd.n3230 vdd.n391 19.3944
R20724 vdd.n3230 vdd.n3229 19.3944
R20725 vdd.n3229 vdd.n3228 19.3944
R20726 vdd.n3228 vdd.n398 19.3944
R20727 vdd.n3223 vdd.n398 19.3944
R20728 vdd.n3223 vdd.n3222 19.3944
R20729 vdd.n3292 vdd.n3291 19.3944
R20730 vdd.n3291 vdd.n3290 19.3944
R20731 vdd.n3290 vdd.n336 19.3944
R20732 vdd.n337 vdd.n336 19.3944
R20733 vdd.n3283 vdd.n337 19.3944
R20734 vdd.n3283 vdd.n3282 19.3944
R20735 vdd.n3282 vdd.n3281 19.3944
R20736 vdd.n3281 vdd.n344 19.3944
R20737 vdd.n3276 vdd.n344 19.3944
R20738 vdd.n3276 vdd.n3275 19.3944
R20739 vdd.n3275 vdd.n3274 19.3944
R20740 vdd.n3274 vdd.n351 19.3944
R20741 vdd.n3269 vdd.n351 19.3944
R20742 vdd.n3269 vdd.n3268 19.3944
R20743 vdd.n3268 vdd.n3267 19.3944
R20744 vdd.n3267 vdd.n358 19.3944
R20745 vdd.n3262 vdd.n358 19.3944
R20746 vdd.n3262 vdd.n3261 19.3944
R20747 vdd.n3119 vdd.n480 19.3944
R20748 vdd.n3119 vdd.n471 19.3944
R20749 vdd.n3132 vdd.n471 19.3944
R20750 vdd.n3132 vdd.n469 19.3944
R20751 vdd.n3136 vdd.n469 19.3944
R20752 vdd.n3136 vdd.n460 19.3944
R20753 vdd.n3148 vdd.n460 19.3944
R20754 vdd.n3148 vdd.n458 19.3944
R20755 vdd.n3152 vdd.n458 19.3944
R20756 vdd.n3152 vdd.n300 19.3944
R20757 vdd.n3317 vdd.n300 19.3944
R20758 vdd.n3317 vdd.n301 19.3944
R20759 vdd.n3311 vdd.n301 19.3944
R20760 vdd.n3311 vdd.n3310 19.3944
R20761 vdd.n3310 vdd.n3309 19.3944
R20762 vdd.n3309 vdd.n313 19.3944
R20763 vdd.n3303 vdd.n313 19.3944
R20764 vdd.n3303 vdd.n3302 19.3944
R20765 vdd.n3302 vdd.n3301 19.3944
R20766 vdd.n3301 vdd.n324 19.3944
R20767 vdd.n3295 vdd.n324 19.3944
R20768 vdd.n3072 vdd.n536 19.3944
R20769 vdd.n3072 vdd.n3069 19.3944
R20770 vdd.n3069 vdd.n3066 19.3944
R20771 vdd.n3066 vdd.n3065 19.3944
R20772 vdd.n3065 vdd.n3062 19.3944
R20773 vdd.n3062 vdd.n3061 19.3944
R20774 vdd.n3061 vdd.n3058 19.3944
R20775 vdd.n3058 vdd.n3057 19.3944
R20776 vdd.n3057 vdd.n3054 19.3944
R20777 vdd.n3054 vdd.n3053 19.3944
R20778 vdd.n3053 vdd.n3050 19.3944
R20779 vdd.n3050 vdd.n3049 19.3944
R20780 vdd.n3049 vdd.n3046 19.3944
R20781 vdd.n3046 vdd.n3045 19.3944
R20782 vdd.n3045 vdd.n3042 19.3944
R20783 vdd.n3042 vdd.n3041 19.3944
R20784 vdd.n3041 vdd.n3038 19.3944
R20785 vdd.n3038 vdd.n3037 19.3944
R20786 vdd.n3037 vdd.n3034 19.3944
R20787 vdd.n3034 vdd.n3033 19.3944
R20788 vdd.n3115 vdd.n482 19.3944
R20789 vdd.n3110 vdd.n482 19.3944
R20790 vdd.n521 vdd.n518 19.3944
R20791 vdd.n3106 vdd.n3105 19.3944
R20792 vdd.n3105 vdd.n3102 19.3944
R20793 vdd.n3102 vdd.n3101 19.3944
R20794 vdd.n3101 vdd.n3098 19.3944
R20795 vdd.n3098 vdd.n3097 19.3944
R20796 vdd.n3097 vdd.n3094 19.3944
R20797 vdd.n3094 vdd.n3093 19.3944
R20798 vdd.n3093 vdd.n3090 19.3944
R20799 vdd.n3090 vdd.n3089 19.3944
R20800 vdd.n3089 vdd.n3086 19.3944
R20801 vdd.n3086 vdd.n3085 19.3944
R20802 vdd.n3085 vdd.n3082 19.3944
R20803 vdd.n3082 vdd.n3081 19.3944
R20804 vdd.n3026 vdd.n556 19.3944
R20805 vdd.n3026 vdd.n3023 19.3944
R20806 vdd.n3023 vdd.n3020 19.3944
R20807 vdd.n3020 vdd.n3019 19.3944
R20808 vdd.n3019 vdd.n3016 19.3944
R20809 vdd.n3016 vdd.n3015 19.3944
R20810 vdd.n3015 vdd.n3012 19.3944
R20811 vdd.n3012 vdd.n3011 19.3944
R20812 vdd.n3011 vdd.n3008 19.3944
R20813 vdd.n3008 vdd.n3007 19.3944
R20814 vdd.n3007 vdd.n3004 19.3944
R20815 vdd.n3004 vdd.n3003 19.3944
R20816 vdd.n3003 vdd.n3000 19.3944
R20817 vdd.n3000 vdd.n2999 19.3944
R20818 vdd.n2999 vdd.n2996 19.3944
R20819 vdd.n2996 vdd.n2995 19.3944
R20820 vdd.n2992 vdd.n2991 19.3944
R20821 vdd.n2988 vdd.n2987 19.3944
R20822 vdd.n1815 vdd.n1811 19.0066
R20823 vdd.n2014 vdd.n1037 19.0066
R20824 vdd.n3221 vdd.n404 19.0066
R20825 vdd.n3030 vdd.n556 19.0066
R20826 vdd.n1106 vdd.n1105 16.0975
R20827 vdd.n801 vdd.n800 16.0975
R20828 vdd.n1776 vdd.n1775 16.0975
R20829 vdd.n1814 vdd.n1813 16.0975
R20830 vdd.n1710 vdd.n1709 16.0975
R20831 vdd.n1977 vdd.n1976 16.0975
R20832 vdd.n1039 vdd.n1038 16.0975
R20833 vdd.n999 vdd.n998 16.0975
R20834 vdd.n1110 vdd.n1109 16.0975
R20835 vdd.n792 vdd.n791 16.0975
R20836 vdd.n2438 vdd.n2437 16.0975
R20837 vdd.n3181 vdd.n3180 16.0975
R20838 vdd.n406 vdd.n405 16.0975
R20839 vdd.n366 vdd.n365 16.0975
R20840 vdd.n558 vdd.n557 16.0975
R20841 vdd.n3077 vdd.n3076 16.0975
R20842 vdd.n623 vdd.n622 16.0975
R20843 vdd.n2435 vdd.n2434 16.0975
R20844 vdd.n2984 vdd.n2983 16.0975
R20845 vdd.n590 vdd.n589 16.0975
R20846 vdd.t33 vdd.n2398 15.4182
R20847 vdd.n2702 vdd.t20 15.4182
R20848 vdd.n28 vdd.n27 14.8792
R20849 vdd.n292 vdd.n257 13.1884
R20850 vdd.n245 vdd.n210 13.1884
R20851 vdd.n202 vdd.n167 13.1884
R20852 vdd.n155 vdd.n120 13.1884
R20853 vdd.n113 vdd.n78 13.1884
R20854 vdd.n66 vdd.n31 13.1884
R20855 vdd.n1562 vdd.n1527 13.1884
R20856 vdd.n1609 vdd.n1574 13.1884
R20857 vdd.n1472 vdd.n1437 13.1884
R20858 vdd.n1519 vdd.n1484 13.1884
R20859 vdd.n1383 vdd.n1348 13.1884
R20860 vdd.n1430 vdd.n1395 13.1884
R20861 vdd.n2120 vdd.n924 13.1509
R20862 vdd.n2945 vdd.n484 13.1509
R20863 vdd.n1846 vdd.n1711 12.9944
R20864 vdd.n1850 vdd.n1711 12.9944
R20865 vdd.n2053 vdd.n997 12.9944
R20866 vdd.n2054 vdd.n2053 12.9944
R20867 vdd.n3260 vdd.n364 12.9944
R20868 vdd.n3261 vdd.n3260 12.9944
R20869 vdd.n3078 vdd.n536 12.9944
R20870 vdd.n3081 vdd.n3078 12.9944
R20871 vdd.n293 vdd.n255 12.8005
R20872 vdd.n288 vdd.n259 12.8005
R20873 vdd.n246 vdd.n208 12.8005
R20874 vdd.n241 vdd.n212 12.8005
R20875 vdd.n203 vdd.n165 12.8005
R20876 vdd.n198 vdd.n169 12.8005
R20877 vdd.n156 vdd.n118 12.8005
R20878 vdd.n151 vdd.n122 12.8005
R20879 vdd.n114 vdd.n76 12.8005
R20880 vdd.n109 vdd.n80 12.8005
R20881 vdd.n67 vdd.n29 12.8005
R20882 vdd.n62 vdd.n33 12.8005
R20883 vdd.n1563 vdd.n1525 12.8005
R20884 vdd.n1558 vdd.n1529 12.8005
R20885 vdd.n1610 vdd.n1572 12.8005
R20886 vdd.n1605 vdd.n1576 12.8005
R20887 vdd.n1473 vdd.n1435 12.8005
R20888 vdd.n1468 vdd.n1439 12.8005
R20889 vdd.n1520 vdd.n1482 12.8005
R20890 vdd.n1515 vdd.n1486 12.8005
R20891 vdd.n1384 vdd.n1346 12.8005
R20892 vdd.n1379 vdd.n1350 12.8005
R20893 vdd.n1431 vdd.n1393 12.8005
R20894 vdd.n1426 vdd.n1397 12.8005
R20895 vdd.n287 vdd.n260 12.0247
R20896 vdd.n240 vdd.n213 12.0247
R20897 vdd.n197 vdd.n170 12.0247
R20898 vdd.n150 vdd.n123 12.0247
R20899 vdd.n108 vdd.n81 12.0247
R20900 vdd.n61 vdd.n34 12.0247
R20901 vdd.n1557 vdd.n1530 12.0247
R20902 vdd.n1604 vdd.n1577 12.0247
R20903 vdd.n1467 vdd.n1440 12.0247
R20904 vdd.n1514 vdd.n1487 12.0247
R20905 vdd.n1378 vdd.n1351 12.0247
R20906 vdd.n1425 vdd.n1398 12.0247
R20907 vdd.n1885 vdd.n1641 11.337
R20908 vdd.n1894 vdd.n1641 11.337
R20909 vdd.n1894 vdd.n1893 11.337
R20910 vdd.n1902 vdd.n1635 11.337
R20911 vdd.n1911 vdd.n1910 11.337
R20912 vdd.n1928 vdd.n1619 11.337
R20913 vdd.n1936 vdd.n1342 11.337
R20914 vdd.n1945 vdd.n1944 11.337
R20915 vdd.n1953 vdd.n1325 11.337
R20916 vdd.n1964 vdd.n1325 11.337
R20917 vdd.n1964 vdd.n1963 11.337
R20918 vdd.n3121 vdd.n473 11.337
R20919 vdd.n3130 vdd.n473 11.337
R20920 vdd.n3130 vdd.n3129 11.337
R20921 vdd.n3138 vdd.n467 11.337
R20922 vdd.n3154 vdd.n456 11.337
R20923 vdd.n3315 vdd.n304 11.337
R20924 vdd.n3313 vdd.n308 11.337
R20925 vdd.n3307 vdd.n3306 11.337
R20926 vdd.n3305 vdd.n318 11.337
R20927 vdd.n3299 vdd.n318 11.337
R20928 vdd.n3299 vdd.n3298 11.337
R20929 vdd.n284 vdd.n283 11.249
R20930 vdd.n237 vdd.n236 11.249
R20931 vdd.n194 vdd.n193 11.249
R20932 vdd.n147 vdd.n146 11.249
R20933 vdd.n105 vdd.n104 11.249
R20934 vdd.n58 vdd.n57 11.249
R20935 vdd.n1554 vdd.n1553 11.249
R20936 vdd.n1601 vdd.n1600 11.249
R20937 vdd.n1464 vdd.n1463 11.249
R20938 vdd.n1511 vdd.n1510 11.249
R20939 vdd.n1375 vdd.n1374 11.249
R20940 vdd.n1422 vdd.n1421 11.249
R20941 vdd.n1683 vdd.t94 10.7702
R20942 vdd.t101 vdd.n3297 10.7702
R20943 vdd.n269 vdd.n268 10.7238
R20944 vdd.n222 vdd.n221 10.7238
R20945 vdd.n179 vdd.n178 10.7238
R20946 vdd.n132 vdd.n131 10.7238
R20947 vdd.n90 vdd.n89 10.7238
R20948 vdd.n43 vdd.n42 10.7238
R20949 vdd.n1539 vdd.n1538 10.7238
R20950 vdd.n1586 vdd.n1585 10.7238
R20951 vdd.n1449 vdd.n1448 10.7238
R20952 vdd.n1496 vdd.n1495 10.7238
R20953 vdd.n1360 vdd.n1359 10.7238
R20954 vdd.n1407 vdd.n1406 10.7238
R20955 vdd.n2125 vdd.n2124 10.6151
R20956 vdd.n2125 vdd.n917 10.6151
R20957 vdd.n2135 vdd.n917 10.6151
R20958 vdd.n2136 vdd.n2135 10.6151
R20959 vdd.n2137 vdd.n2136 10.6151
R20960 vdd.n2137 vdd.n904 10.6151
R20961 vdd.n2147 vdd.n904 10.6151
R20962 vdd.n2148 vdd.n2147 10.6151
R20963 vdd.n2149 vdd.n2148 10.6151
R20964 vdd.n2149 vdd.n892 10.6151
R20965 vdd.n2159 vdd.n892 10.6151
R20966 vdd.n2160 vdd.n2159 10.6151
R20967 vdd.n2161 vdd.n2160 10.6151
R20968 vdd.n2161 vdd.n881 10.6151
R20969 vdd.n2171 vdd.n881 10.6151
R20970 vdd.n2172 vdd.n2171 10.6151
R20971 vdd.n2173 vdd.n2172 10.6151
R20972 vdd.n2173 vdd.n868 10.6151
R20973 vdd.n2183 vdd.n868 10.6151
R20974 vdd.n2184 vdd.n2183 10.6151
R20975 vdd.n2185 vdd.n2184 10.6151
R20976 vdd.n2185 vdd.n856 10.6151
R20977 vdd.n2196 vdd.n856 10.6151
R20978 vdd.n2197 vdd.n2196 10.6151
R20979 vdd.n2198 vdd.n2197 10.6151
R20980 vdd.n2198 vdd.n844 10.6151
R20981 vdd.n2208 vdd.n844 10.6151
R20982 vdd.n2209 vdd.n2208 10.6151
R20983 vdd.n2210 vdd.n2209 10.6151
R20984 vdd.n2210 vdd.n832 10.6151
R20985 vdd.n2220 vdd.n832 10.6151
R20986 vdd.n2221 vdd.n2220 10.6151
R20987 vdd.n2222 vdd.n2221 10.6151
R20988 vdd.n2222 vdd.n822 10.6151
R20989 vdd.n2232 vdd.n822 10.6151
R20990 vdd.n2233 vdd.n2232 10.6151
R20991 vdd.n2234 vdd.n2233 10.6151
R20992 vdd.n2234 vdd.n809 10.6151
R20993 vdd.n2246 vdd.n809 10.6151
R20994 vdd.n2247 vdd.n2246 10.6151
R20995 vdd.n2249 vdd.n2247 10.6151
R20996 vdd.n2249 vdd.n2248 10.6151
R20997 vdd.n2248 vdd.n790 10.6151
R20998 vdd.n2396 vdd.n2395 10.6151
R20999 vdd.n2395 vdd.n2394 10.6151
R21000 vdd.n2394 vdd.n2391 10.6151
R21001 vdd.n2391 vdd.n2390 10.6151
R21002 vdd.n2390 vdd.n2387 10.6151
R21003 vdd.n2387 vdd.n2386 10.6151
R21004 vdd.n2386 vdd.n2383 10.6151
R21005 vdd.n2383 vdd.n2382 10.6151
R21006 vdd.n2382 vdd.n2379 10.6151
R21007 vdd.n2379 vdd.n2378 10.6151
R21008 vdd.n2378 vdd.n2375 10.6151
R21009 vdd.n2375 vdd.n2374 10.6151
R21010 vdd.n2374 vdd.n2371 10.6151
R21011 vdd.n2371 vdd.n2370 10.6151
R21012 vdd.n2370 vdd.n2367 10.6151
R21013 vdd.n2367 vdd.n2366 10.6151
R21014 vdd.n2366 vdd.n2363 10.6151
R21015 vdd.n2363 vdd.n2362 10.6151
R21016 vdd.n2362 vdd.n2359 10.6151
R21017 vdd.n2359 vdd.n2358 10.6151
R21018 vdd.n2358 vdd.n2355 10.6151
R21019 vdd.n2355 vdd.n2354 10.6151
R21020 vdd.n2354 vdd.n2351 10.6151
R21021 vdd.n2351 vdd.n2350 10.6151
R21022 vdd.n2350 vdd.n2347 10.6151
R21023 vdd.n2347 vdd.n2346 10.6151
R21024 vdd.n2346 vdd.n2343 10.6151
R21025 vdd.n2343 vdd.n2342 10.6151
R21026 vdd.n2342 vdd.n2339 10.6151
R21027 vdd.n2339 vdd.n2338 10.6151
R21028 vdd.n2338 vdd.n2335 10.6151
R21029 vdd.n2333 vdd.n2330 10.6151
R21030 vdd.n2330 vdd.n2329 10.6151
R21031 vdd.n1147 vdd.n1146 10.6151
R21032 vdd.n1149 vdd.n1147 10.6151
R21033 vdd.n1150 vdd.n1149 10.6151
R21034 vdd.n1152 vdd.n1150 10.6151
R21035 vdd.n1153 vdd.n1152 10.6151
R21036 vdd.n1155 vdd.n1153 10.6151
R21037 vdd.n1156 vdd.n1155 10.6151
R21038 vdd.n1158 vdd.n1156 10.6151
R21039 vdd.n1159 vdd.n1158 10.6151
R21040 vdd.n1161 vdd.n1159 10.6151
R21041 vdd.n1162 vdd.n1161 10.6151
R21042 vdd.n1164 vdd.n1162 10.6151
R21043 vdd.n1165 vdd.n1164 10.6151
R21044 vdd.n1167 vdd.n1165 10.6151
R21045 vdd.n1168 vdd.n1167 10.6151
R21046 vdd.n1170 vdd.n1168 10.6151
R21047 vdd.n1171 vdd.n1170 10.6151
R21048 vdd.n1173 vdd.n1171 10.6151
R21049 vdd.n1174 vdd.n1173 10.6151
R21050 vdd.n1176 vdd.n1174 10.6151
R21051 vdd.n1177 vdd.n1176 10.6151
R21052 vdd.n1179 vdd.n1177 10.6151
R21053 vdd.n1180 vdd.n1179 10.6151
R21054 vdd.n1182 vdd.n1180 10.6151
R21055 vdd.n1183 vdd.n1182 10.6151
R21056 vdd.n1185 vdd.n1183 10.6151
R21057 vdd.n1186 vdd.n1185 10.6151
R21058 vdd.n1225 vdd.n1186 10.6151
R21059 vdd.n1225 vdd.n1224 10.6151
R21060 vdd.n1224 vdd.n1223 10.6151
R21061 vdd.n1223 vdd.n1221 10.6151
R21062 vdd.n1221 vdd.n1220 10.6151
R21063 vdd.n1220 vdd.n1218 10.6151
R21064 vdd.n1218 vdd.n1217 10.6151
R21065 vdd.n1217 vdd.n1198 10.6151
R21066 vdd.n1198 vdd.n1197 10.6151
R21067 vdd.n1197 vdd.n1195 10.6151
R21068 vdd.n1195 vdd.n1194 10.6151
R21069 vdd.n1194 vdd.n1192 10.6151
R21070 vdd.n1192 vdd.n1191 10.6151
R21071 vdd.n1191 vdd.n1188 10.6151
R21072 vdd.n1188 vdd.n1187 10.6151
R21073 vdd.n1187 vdd.n793 10.6151
R21074 vdd.n2123 vdd.n929 10.6151
R21075 vdd.n2118 vdd.n929 10.6151
R21076 vdd.n2118 vdd.n2117 10.6151
R21077 vdd.n2117 vdd.n2116 10.6151
R21078 vdd.n2116 vdd.n2113 10.6151
R21079 vdd.n2113 vdd.n2112 10.6151
R21080 vdd.n2112 vdd.n2109 10.6151
R21081 vdd.n2109 vdd.n2108 10.6151
R21082 vdd.n2108 vdd.n2105 10.6151
R21083 vdd.n2105 vdd.n2104 10.6151
R21084 vdd.n2104 vdd.n2101 10.6151
R21085 vdd.n2101 vdd.n2100 10.6151
R21086 vdd.n2100 vdd.n2097 10.6151
R21087 vdd.n2097 vdd.n2096 10.6151
R21088 vdd.n2096 vdd.n2093 10.6151
R21089 vdd.n2093 vdd.n2092 10.6151
R21090 vdd.n2092 vdd.n2089 10.6151
R21091 vdd.n2089 vdd.n967 10.6151
R21092 vdd.n1113 vdd.n967 10.6151
R21093 vdd.n1114 vdd.n1113 10.6151
R21094 vdd.n1117 vdd.n1114 10.6151
R21095 vdd.n1118 vdd.n1117 10.6151
R21096 vdd.n1121 vdd.n1118 10.6151
R21097 vdd.n1122 vdd.n1121 10.6151
R21098 vdd.n1125 vdd.n1122 10.6151
R21099 vdd.n1126 vdd.n1125 10.6151
R21100 vdd.n1129 vdd.n1126 10.6151
R21101 vdd.n1130 vdd.n1129 10.6151
R21102 vdd.n1133 vdd.n1130 10.6151
R21103 vdd.n1134 vdd.n1133 10.6151
R21104 vdd.n1137 vdd.n1134 10.6151
R21105 vdd.n1142 vdd.n1139 10.6151
R21106 vdd.n1143 vdd.n1142 10.6151
R21107 vdd.n2634 vdd.n2633 10.6151
R21108 vdd.n2633 vdd.n2632 10.6151
R21109 vdd.n2632 vdd.n2436 10.6151
R21110 vdd.n2514 vdd.n2436 10.6151
R21111 vdd.n2515 vdd.n2514 10.6151
R21112 vdd.n2517 vdd.n2515 10.6151
R21113 vdd.n2518 vdd.n2517 10.6151
R21114 vdd.n2616 vdd.n2518 10.6151
R21115 vdd.n2616 vdd.n2615 10.6151
R21116 vdd.n2615 vdd.n2614 10.6151
R21117 vdd.n2614 vdd.n2562 10.6151
R21118 vdd.n2562 vdd.n2561 10.6151
R21119 vdd.n2561 vdd.n2559 10.6151
R21120 vdd.n2559 vdd.n2558 10.6151
R21121 vdd.n2558 vdd.n2556 10.6151
R21122 vdd.n2556 vdd.n2555 10.6151
R21123 vdd.n2555 vdd.n2553 10.6151
R21124 vdd.n2553 vdd.n2552 10.6151
R21125 vdd.n2552 vdd.n2550 10.6151
R21126 vdd.n2550 vdd.n2549 10.6151
R21127 vdd.n2549 vdd.n2547 10.6151
R21128 vdd.n2547 vdd.n2546 10.6151
R21129 vdd.n2546 vdd.n2544 10.6151
R21130 vdd.n2544 vdd.n2543 10.6151
R21131 vdd.n2543 vdd.n2541 10.6151
R21132 vdd.n2541 vdd.n2540 10.6151
R21133 vdd.n2540 vdd.n2538 10.6151
R21134 vdd.n2538 vdd.n2537 10.6151
R21135 vdd.n2537 vdd.n2535 10.6151
R21136 vdd.n2535 vdd.n2534 10.6151
R21137 vdd.n2534 vdd.n2532 10.6151
R21138 vdd.n2532 vdd.n2531 10.6151
R21139 vdd.n2531 vdd.n2529 10.6151
R21140 vdd.n2529 vdd.n2528 10.6151
R21141 vdd.n2528 vdd.n2526 10.6151
R21142 vdd.n2526 vdd.n2525 10.6151
R21143 vdd.n2525 vdd.n2523 10.6151
R21144 vdd.n2523 vdd.n2522 10.6151
R21145 vdd.n2522 vdd.n2520 10.6151
R21146 vdd.n2520 vdd.n2519 10.6151
R21147 vdd.n2519 vdd.n626 10.6151
R21148 vdd.n2878 vdd.n626 10.6151
R21149 vdd.n2879 vdd.n2878 10.6151
R21150 vdd.n2705 vdd.n751 10.6151
R21151 vdd.n2700 vdd.n751 10.6151
R21152 vdd.n2700 vdd.n2699 10.6151
R21153 vdd.n2699 vdd.n2698 10.6151
R21154 vdd.n2698 vdd.n2695 10.6151
R21155 vdd.n2695 vdd.n2694 10.6151
R21156 vdd.n2694 vdd.n2691 10.6151
R21157 vdd.n2691 vdd.n2690 10.6151
R21158 vdd.n2690 vdd.n2687 10.6151
R21159 vdd.n2687 vdd.n2686 10.6151
R21160 vdd.n2686 vdd.n2683 10.6151
R21161 vdd.n2683 vdd.n2682 10.6151
R21162 vdd.n2682 vdd.n2679 10.6151
R21163 vdd.n2679 vdd.n2678 10.6151
R21164 vdd.n2678 vdd.n2675 10.6151
R21165 vdd.n2675 vdd.n2674 10.6151
R21166 vdd.n2674 vdd.n2671 10.6151
R21167 vdd.n2671 vdd.n2670 10.6151
R21168 vdd.n2670 vdd.n2667 10.6151
R21169 vdd.n2667 vdd.n2666 10.6151
R21170 vdd.n2666 vdd.n2663 10.6151
R21171 vdd.n2663 vdd.n2662 10.6151
R21172 vdd.n2662 vdd.n2659 10.6151
R21173 vdd.n2659 vdd.n2658 10.6151
R21174 vdd.n2658 vdd.n2655 10.6151
R21175 vdd.n2655 vdd.n2654 10.6151
R21176 vdd.n2654 vdd.n2651 10.6151
R21177 vdd.n2651 vdd.n2650 10.6151
R21178 vdd.n2650 vdd.n2647 10.6151
R21179 vdd.n2647 vdd.n2646 10.6151
R21180 vdd.n2646 vdd.n2643 10.6151
R21181 vdd.n2641 vdd.n2638 10.6151
R21182 vdd.n2638 vdd.n2637 10.6151
R21183 vdd.n2707 vdd.n2706 10.6151
R21184 vdd.n2707 vdd.n740 10.6151
R21185 vdd.n2717 vdd.n740 10.6151
R21186 vdd.n2718 vdd.n2717 10.6151
R21187 vdd.n2719 vdd.n2718 10.6151
R21188 vdd.n2719 vdd.n728 10.6151
R21189 vdd.n2729 vdd.n728 10.6151
R21190 vdd.n2730 vdd.n2729 10.6151
R21191 vdd.n2731 vdd.n2730 10.6151
R21192 vdd.n2731 vdd.n717 10.6151
R21193 vdd.n2741 vdd.n717 10.6151
R21194 vdd.n2742 vdd.n2741 10.6151
R21195 vdd.n2743 vdd.n2742 10.6151
R21196 vdd.n2743 vdd.n706 10.6151
R21197 vdd.n2753 vdd.n706 10.6151
R21198 vdd.n2754 vdd.n2753 10.6151
R21199 vdd.n2755 vdd.n2754 10.6151
R21200 vdd.n2755 vdd.n693 10.6151
R21201 vdd.n2766 vdd.n693 10.6151
R21202 vdd.n2767 vdd.n2766 10.6151
R21203 vdd.n2768 vdd.n2767 10.6151
R21204 vdd.n2768 vdd.n681 10.6151
R21205 vdd.n2778 vdd.n681 10.6151
R21206 vdd.n2779 vdd.n2778 10.6151
R21207 vdd.n2780 vdd.n2779 10.6151
R21208 vdd.n2780 vdd.n669 10.6151
R21209 vdd.n2790 vdd.n669 10.6151
R21210 vdd.n2791 vdd.n2790 10.6151
R21211 vdd.n2792 vdd.n2791 10.6151
R21212 vdd.n2792 vdd.n656 10.6151
R21213 vdd.n2802 vdd.n656 10.6151
R21214 vdd.n2803 vdd.n2802 10.6151
R21215 vdd.n2804 vdd.n2803 10.6151
R21216 vdd.n2804 vdd.n645 10.6151
R21217 vdd.n2814 vdd.n645 10.6151
R21218 vdd.n2815 vdd.n2814 10.6151
R21219 vdd.n2816 vdd.n2815 10.6151
R21220 vdd.n2816 vdd.n631 10.6151
R21221 vdd.n2871 vdd.n631 10.6151
R21222 vdd.n2872 vdd.n2871 10.6151
R21223 vdd.n2873 vdd.n2872 10.6151
R21224 vdd.n2873 vdd.n600 10.6151
R21225 vdd.n2943 vdd.n600 10.6151
R21226 vdd.n2942 vdd.n2941 10.6151
R21227 vdd.n2941 vdd.n601 10.6151
R21228 vdd.n602 vdd.n601 10.6151
R21229 vdd.n2934 vdd.n602 10.6151
R21230 vdd.n2934 vdd.n2933 10.6151
R21231 vdd.n2933 vdd.n2932 10.6151
R21232 vdd.n2932 vdd.n604 10.6151
R21233 vdd.n2927 vdd.n604 10.6151
R21234 vdd.n2927 vdd.n2926 10.6151
R21235 vdd.n2926 vdd.n2925 10.6151
R21236 vdd.n2925 vdd.n607 10.6151
R21237 vdd.n2920 vdd.n607 10.6151
R21238 vdd.n2920 vdd.n2919 10.6151
R21239 vdd.n2919 vdd.n2918 10.6151
R21240 vdd.n2918 vdd.n610 10.6151
R21241 vdd.n2913 vdd.n610 10.6151
R21242 vdd.n2913 vdd.n520 10.6151
R21243 vdd.n2909 vdd.n520 10.6151
R21244 vdd.n2909 vdd.n2908 10.6151
R21245 vdd.n2908 vdd.n2907 10.6151
R21246 vdd.n2907 vdd.n613 10.6151
R21247 vdd.n2902 vdd.n613 10.6151
R21248 vdd.n2902 vdd.n2901 10.6151
R21249 vdd.n2901 vdd.n2900 10.6151
R21250 vdd.n2900 vdd.n616 10.6151
R21251 vdd.n2895 vdd.n616 10.6151
R21252 vdd.n2895 vdd.n2894 10.6151
R21253 vdd.n2894 vdd.n2893 10.6151
R21254 vdd.n2893 vdd.n619 10.6151
R21255 vdd.n2888 vdd.n619 10.6151
R21256 vdd.n2888 vdd.n2887 10.6151
R21257 vdd.n2885 vdd.n624 10.6151
R21258 vdd.n2880 vdd.n624 10.6151
R21259 vdd.n2861 vdd.n2822 10.6151
R21260 vdd.n2856 vdd.n2822 10.6151
R21261 vdd.n2856 vdd.n2855 10.6151
R21262 vdd.n2855 vdd.n2854 10.6151
R21263 vdd.n2854 vdd.n2824 10.6151
R21264 vdd.n2849 vdd.n2824 10.6151
R21265 vdd.n2849 vdd.n2848 10.6151
R21266 vdd.n2848 vdd.n2847 10.6151
R21267 vdd.n2847 vdd.n2827 10.6151
R21268 vdd.n2842 vdd.n2827 10.6151
R21269 vdd.n2842 vdd.n2841 10.6151
R21270 vdd.n2841 vdd.n2840 10.6151
R21271 vdd.n2840 vdd.n2830 10.6151
R21272 vdd.n2835 vdd.n2830 10.6151
R21273 vdd.n2835 vdd.n2834 10.6151
R21274 vdd.n2834 vdd.n575 10.6151
R21275 vdd.n2978 vdd.n575 10.6151
R21276 vdd.n2978 vdd.n576 10.6151
R21277 vdd.n578 vdd.n576 10.6151
R21278 vdd.n2971 vdd.n578 10.6151
R21279 vdd.n2971 vdd.n2970 10.6151
R21280 vdd.n2970 vdd.n2969 10.6151
R21281 vdd.n2969 vdd.n580 10.6151
R21282 vdd.n2964 vdd.n580 10.6151
R21283 vdd.n2964 vdd.n2963 10.6151
R21284 vdd.n2963 vdd.n2962 10.6151
R21285 vdd.n2962 vdd.n583 10.6151
R21286 vdd.n2957 vdd.n583 10.6151
R21287 vdd.n2957 vdd.n2956 10.6151
R21288 vdd.n2956 vdd.n2955 10.6151
R21289 vdd.n2955 vdd.n586 10.6151
R21290 vdd.n2950 vdd.n2949 10.6151
R21291 vdd.n2949 vdd.n2948 10.6151
R21292 vdd.n2511 vdd.n2510 10.6151
R21293 vdd.n2628 vdd.n2511 10.6151
R21294 vdd.n2628 vdd.n2627 10.6151
R21295 vdd.n2627 vdd.n2626 10.6151
R21296 vdd.n2626 vdd.n2624 10.6151
R21297 vdd.n2624 vdd.n2623 10.6151
R21298 vdd.n2623 vdd.n2621 10.6151
R21299 vdd.n2621 vdd.n2620 10.6151
R21300 vdd.n2620 vdd.n2512 10.6151
R21301 vdd.n2610 vdd.n2512 10.6151
R21302 vdd.n2610 vdd.n2609 10.6151
R21303 vdd.n2609 vdd.n2608 10.6151
R21304 vdd.n2608 vdd.n2606 10.6151
R21305 vdd.n2606 vdd.n2605 10.6151
R21306 vdd.n2605 vdd.n2603 10.6151
R21307 vdd.n2603 vdd.n2602 10.6151
R21308 vdd.n2602 vdd.n2600 10.6151
R21309 vdd.n2600 vdd.n2599 10.6151
R21310 vdd.n2599 vdd.n2597 10.6151
R21311 vdd.n2597 vdd.n2596 10.6151
R21312 vdd.n2596 vdd.n2594 10.6151
R21313 vdd.n2594 vdd.n2593 10.6151
R21314 vdd.n2593 vdd.n2591 10.6151
R21315 vdd.n2591 vdd.n2590 10.6151
R21316 vdd.n2590 vdd.n2588 10.6151
R21317 vdd.n2588 vdd.n2587 10.6151
R21318 vdd.n2587 vdd.n2585 10.6151
R21319 vdd.n2585 vdd.n2584 10.6151
R21320 vdd.n2584 vdd.n2582 10.6151
R21321 vdd.n2582 vdd.n2581 10.6151
R21322 vdd.n2581 vdd.n2579 10.6151
R21323 vdd.n2579 vdd.n2578 10.6151
R21324 vdd.n2578 vdd.n2576 10.6151
R21325 vdd.n2576 vdd.n2575 10.6151
R21326 vdd.n2575 vdd.n2573 10.6151
R21327 vdd.n2573 vdd.n2572 10.6151
R21328 vdd.n2572 vdd.n2570 10.6151
R21329 vdd.n2570 vdd.n2569 10.6151
R21330 vdd.n2569 vdd.n2567 10.6151
R21331 vdd.n2567 vdd.n2566 10.6151
R21332 vdd.n2566 vdd.n2564 10.6151
R21333 vdd.n2564 vdd.n2563 10.6151
R21334 vdd.n2563 vdd.n592 10.6151
R21335 vdd.n2442 vdd.n2441 10.6151
R21336 vdd.n2445 vdd.n2442 10.6151
R21337 vdd.n2446 vdd.n2445 10.6151
R21338 vdd.n2449 vdd.n2446 10.6151
R21339 vdd.n2450 vdd.n2449 10.6151
R21340 vdd.n2453 vdd.n2450 10.6151
R21341 vdd.n2454 vdd.n2453 10.6151
R21342 vdd.n2457 vdd.n2454 10.6151
R21343 vdd.n2458 vdd.n2457 10.6151
R21344 vdd.n2461 vdd.n2458 10.6151
R21345 vdd.n2462 vdd.n2461 10.6151
R21346 vdd.n2465 vdd.n2462 10.6151
R21347 vdd.n2466 vdd.n2465 10.6151
R21348 vdd.n2469 vdd.n2466 10.6151
R21349 vdd.n2470 vdd.n2469 10.6151
R21350 vdd.n2473 vdd.n2470 10.6151
R21351 vdd.n2474 vdd.n2473 10.6151
R21352 vdd.n2477 vdd.n2474 10.6151
R21353 vdd.n2478 vdd.n2477 10.6151
R21354 vdd.n2481 vdd.n2478 10.6151
R21355 vdd.n2482 vdd.n2481 10.6151
R21356 vdd.n2485 vdd.n2482 10.6151
R21357 vdd.n2486 vdd.n2485 10.6151
R21358 vdd.n2489 vdd.n2486 10.6151
R21359 vdd.n2490 vdd.n2489 10.6151
R21360 vdd.n2493 vdd.n2490 10.6151
R21361 vdd.n2494 vdd.n2493 10.6151
R21362 vdd.n2497 vdd.n2494 10.6151
R21363 vdd.n2498 vdd.n2497 10.6151
R21364 vdd.n2501 vdd.n2498 10.6151
R21365 vdd.n2502 vdd.n2501 10.6151
R21366 vdd.n2507 vdd.n2505 10.6151
R21367 vdd.n2508 vdd.n2507 10.6151
R21368 vdd.n2711 vdd.n745 10.6151
R21369 vdd.n2712 vdd.n2711 10.6151
R21370 vdd.n2713 vdd.n2712 10.6151
R21371 vdd.n2713 vdd.n734 10.6151
R21372 vdd.n2723 vdd.n734 10.6151
R21373 vdd.n2724 vdd.n2723 10.6151
R21374 vdd.n2725 vdd.n2724 10.6151
R21375 vdd.n2725 vdd.n723 10.6151
R21376 vdd.n2735 vdd.n723 10.6151
R21377 vdd.n2736 vdd.n2735 10.6151
R21378 vdd.n2737 vdd.n2736 10.6151
R21379 vdd.n2737 vdd.n711 10.6151
R21380 vdd.n2747 vdd.n711 10.6151
R21381 vdd.n2748 vdd.n2747 10.6151
R21382 vdd.n2749 vdd.n2748 10.6151
R21383 vdd.n2749 vdd.n700 10.6151
R21384 vdd.n2759 vdd.n700 10.6151
R21385 vdd.n2760 vdd.n2759 10.6151
R21386 vdd.n2762 vdd.n2760 10.6151
R21387 vdd.n2762 vdd.n2761 10.6151
R21388 vdd.n2773 vdd.n2772 10.6151
R21389 vdd.n2774 vdd.n2773 10.6151
R21390 vdd.n2774 vdd.n675 10.6151
R21391 vdd.n2784 vdd.n675 10.6151
R21392 vdd.n2785 vdd.n2784 10.6151
R21393 vdd.n2786 vdd.n2785 10.6151
R21394 vdd.n2786 vdd.n662 10.6151
R21395 vdd.n2796 vdd.n662 10.6151
R21396 vdd.n2797 vdd.n2796 10.6151
R21397 vdd.n2798 vdd.n2797 10.6151
R21398 vdd.n2798 vdd.n650 10.6151
R21399 vdd.n2808 vdd.n650 10.6151
R21400 vdd.n2809 vdd.n2808 10.6151
R21401 vdd.n2810 vdd.n2809 10.6151
R21402 vdd.n2810 vdd.n639 10.6151
R21403 vdd.n2820 vdd.n639 10.6151
R21404 vdd.n2821 vdd.n2820 10.6151
R21405 vdd.n2867 vdd.n2821 10.6151
R21406 vdd.n2867 vdd.n2866 10.6151
R21407 vdd.n2866 vdd.n2865 10.6151
R21408 vdd.n2865 vdd.n2864 10.6151
R21409 vdd.n2864 vdd.n2862 10.6151
R21410 vdd.n2129 vdd.n922 10.6151
R21411 vdd.n2130 vdd.n2129 10.6151
R21412 vdd.n2131 vdd.n2130 10.6151
R21413 vdd.n2131 vdd.n911 10.6151
R21414 vdd.n2141 vdd.n911 10.6151
R21415 vdd.n2142 vdd.n2141 10.6151
R21416 vdd.n2143 vdd.n2142 10.6151
R21417 vdd.n2143 vdd.n898 10.6151
R21418 vdd.n2153 vdd.n898 10.6151
R21419 vdd.n2154 vdd.n2153 10.6151
R21420 vdd.n2155 vdd.n2154 10.6151
R21421 vdd.n2155 vdd.n887 10.6151
R21422 vdd.n2165 vdd.n887 10.6151
R21423 vdd.n2166 vdd.n2165 10.6151
R21424 vdd.n2167 vdd.n2166 10.6151
R21425 vdd.n2167 vdd.n875 10.6151
R21426 vdd.n2177 vdd.n875 10.6151
R21427 vdd.n2178 vdd.n2177 10.6151
R21428 vdd.n2179 vdd.n2178 10.6151
R21429 vdd.n2179 vdd.n862 10.6151
R21430 vdd.n2189 vdd.n862 10.6151
R21431 vdd.n2190 vdd.n2189 10.6151
R21432 vdd.n2192 vdd.n850 10.6151
R21433 vdd.n2202 vdd.n850 10.6151
R21434 vdd.n2203 vdd.n2202 10.6151
R21435 vdd.n2204 vdd.n2203 10.6151
R21436 vdd.n2204 vdd.n838 10.6151
R21437 vdd.n2214 vdd.n838 10.6151
R21438 vdd.n2215 vdd.n2214 10.6151
R21439 vdd.n2216 vdd.n2215 10.6151
R21440 vdd.n2216 vdd.n827 10.6151
R21441 vdd.n2226 vdd.n827 10.6151
R21442 vdd.n2227 vdd.n2226 10.6151
R21443 vdd.n2228 vdd.n2227 10.6151
R21444 vdd.n2228 vdd.n816 10.6151
R21445 vdd.n2238 vdd.n816 10.6151
R21446 vdd.n2239 vdd.n2238 10.6151
R21447 vdd.n2242 vdd.n2239 10.6151
R21448 vdd.n2242 vdd.n2241 10.6151
R21449 vdd.n2241 vdd.n2240 10.6151
R21450 vdd.n2240 vdd.n799 10.6151
R21451 vdd.n2324 vdd.n799 10.6151
R21452 vdd.n2323 vdd.n2322 10.6151
R21453 vdd.n2322 vdd.n2319 10.6151
R21454 vdd.n2319 vdd.n2318 10.6151
R21455 vdd.n2318 vdd.n2315 10.6151
R21456 vdd.n2315 vdd.n2314 10.6151
R21457 vdd.n2314 vdd.n2311 10.6151
R21458 vdd.n2311 vdd.n2310 10.6151
R21459 vdd.n2310 vdd.n2307 10.6151
R21460 vdd.n2307 vdd.n2306 10.6151
R21461 vdd.n2306 vdd.n2303 10.6151
R21462 vdd.n2303 vdd.n2302 10.6151
R21463 vdd.n2302 vdd.n2299 10.6151
R21464 vdd.n2299 vdd.n2298 10.6151
R21465 vdd.n2298 vdd.n2295 10.6151
R21466 vdd.n2295 vdd.n2294 10.6151
R21467 vdd.n2294 vdd.n2291 10.6151
R21468 vdd.n2291 vdd.n2290 10.6151
R21469 vdd.n2290 vdd.n2287 10.6151
R21470 vdd.n2287 vdd.n2286 10.6151
R21471 vdd.n2286 vdd.n2283 10.6151
R21472 vdd.n2283 vdd.n2282 10.6151
R21473 vdd.n2282 vdd.n2279 10.6151
R21474 vdd.n2279 vdd.n2278 10.6151
R21475 vdd.n2278 vdd.n2275 10.6151
R21476 vdd.n2275 vdd.n2274 10.6151
R21477 vdd.n2274 vdd.n2271 10.6151
R21478 vdd.n2271 vdd.n2270 10.6151
R21479 vdd.n2270 vdd.n2267 10.6151
R21480 vdd.n2267 vdd.n2266 10.6151
R21481 vdd.n2266 vdd.n2263 10.6151
R21482 vdd.n2263 vdd.n2262 10.6151
R21483 vdd.n2259 vdd.n2258 10.6151
R21484 vdd.n2258 vdd.n2256 10.6151
R21485 vdd.n1271 vdd.n1269 10.6151
R21486 vdd.n1269 vdd.n1268 10.6151
R21487 vdd.n1268 vdd.n1266 10.6151
R21488 vdd.n1266 vdd.n1265 10.6151
R21489 vdd.n1265 vdd.n1263 10.6151
R21490 vdd.n1263 vdd.n1262 10.6151
R21491 vdd.n1262 vdd.n1260 10.6151
R21492 vdd.n1260 vdd.n1259 10.6151
R21493 vdd.n1259 vdd.n1257 10.6151
R21494 vdd.n1257 vdd.n1256 10.6151
R21495 vdd.n1256 vdd.n1254 10.6151
R21496 vdd.n1254 vdd.n1253 10.6151
R21497 vdd.n1253 vdd.n1251 10.6151
R21498 vdd.n1251 vdd.n1250 10.6151
R21499 vdd.n1250 vdd.n1248 10.6151
R21500 vdd.n1248 vdd.n1247 10.6151
R21501 vdd.n1247 vdd.n1245 10.6151
R21502 vdd.n1245 vdd.n1244 10.6151
R21503 vdd.n1244 vdd.n1242 10.6151
R21504 vdd.n1242 vdd.n1241 10.6151
R21505 vdd.n1241 vdd.n1239 10.6151
R21506 vdd.n1239 vdd.n1238 10.6151
R21507 vdd.n1238 vdd.n1236 10.6151
R21508 vdd.n1236 vdd.n1235 10.6151
R21509 vdd.n1235 vdd.n1233 10.6151
R21510 vdd.n1233 vdd.n1232 10.6151
R21511 vdd.n1232 vdd.n1230 10.6151
R21512 vdd.n1230 vdd.n1229 10.6151
R21513 vdd.n1229 vdd.n1108 10.6151
R21514 vdd.n1200 vdd.n1108 10.6151
R21515 vdd.n1201 vdd.n1200 10.6151
R21516 vdd.n1203 vdd.n1201 10.6151
R21517 vdd.n1204 vdd.n1203 10.6151
R21518 vdd.n1213 vdd.n1204 10.6151
R21519 vdd.n1213 vdd.n1212 10.6151
R21520 vdd.n1212 vdd.n1211 10.6151
R21521 vdd.n1211 vdd.n1209 10.6151
R21522 vdd.n1209 vdd.n1208 10.6151
R21523 vdd.n1208 vdd.n1206 10.6151
R21524 vdd.n1206 vdd.n1205 10.6151
R21525 vdd.n1205 vdd.n803 10.6151
R21526 vdd.n2254 vdd.n803 10.6151
R21527 vdd.n2255 vdd.n2254 10.6151
R21528 vdd.n1072 vdd.n1071 10.6151
R21529 vdd.n1075 vdd.n1072 10.6151
R21530 vdd.n1076 vdd.n1075 10.6151
R21531 vdd.n1079 vdd.n1076 10.6151
R21532 vdd.n1080 vdd.n1079 10.6151
R21533 vdd.n1083 vdd.n1080 10.6151
R21534 vdd.n1084 vdd.n1083 10.6151
R21535 vdd.n1087 vdd.n1084 10.6151
R21536 vdd.n1088 vdd.n1087 10.6151
R21537 vdd.n1091 vdd.n1088 10.6151
R21538 vdd.n1092 vdd.n1091 10.6151
R21539 vdd.n1095 vdd.n1092 10.6151
R21540 vdd.n1096 vdd.n1095 10.6151
R21541 vdd.n1099 vdd.n1096 10.6151
R21542 vdd.n1100 vdd.n1099 10.6151
R21543 vdd.n1103 vdd.n1100 10.6151
R21544 vdd.n1305 vdd.n1103 10.6151
R21545 vdd.n1305 vdd.n1304 10.6151
R21546 vdd.n1304 vdd.n1302 10.6151
R21547 vdd.n1302 vdd.n1299 10.6151
R21548 vdd.n1299 vdd.n1298 10.6151
R21549 vdd.n1298 vdd.n1295 10.6151
R21550 vdd.n1295 vdd.n1294 10.6151
R21551 vdd.n1294 vdd.n1291 10.6151
R21552 vdd.n1291 vdd.n1290 10.6151
R21553 vdd.n1290 vdd.n1287 10.6151
R21554 vdd.n1287 vdd.n1286 10.6151
R21555 vdd.n1286 vdd.n1283 10.6151
R21556 vdd.n1283 vdd.n1282 10.6151
R21557 vdd.n1282 vdd.n1279 10.6151
R21558 vdd.n1279 vdd.n1278 10.6151
R21559 vdd.n1275 vdd.n1274 10.6151
R21560 vdd.n1274 vdd.n1272 10.6151
R21561 vdd.n280 vdd.n262 10.4732
R21562 vdd.n233 vdd.n215 10.4732
R21563 vdd.n190 vdd.n172 10.4732
R21564 vdd.n143 vdd.n125 10.4732
R21565 vdd.n101 vdd.n83 10.4732
R21566 vdd.n54 vdd.n36 10.4732
R21567 vdd.n1550 vdd.n1532 10.4732
R21568 vdd.n1597 vdd.n1579 10.4732
R21569 vdd.n1460 vdd.n1442 10.4732
R21570 vdd.n1507 vdd.n1489 10.4732
R21571 vdd.n1371 vdd.n1353 10.4732
R21572 vdd.n1418 vdd.n1400 10.4732
R21573 vdd.t188 vdd.n1343 10.3167
R21574 vdd.n3146 vdd.t156 10.3167
R21575 vdd.n1920 vdd.t168 10.09
R21576 vdd.n3314 vdd.t154 10.09
R21577 vdd.n2089 vdd.n2088 9.98956
R21578 vdd.n3108 vdd.n520 9.98956
R21579 vdd.n2979 vdd.n2978 9.98956
R21580 vdd.n1981 vdd.n1305 9.98956
R21581 vdd.n2326 vdd.t40 9.7499
R21582 vdd.t38 vdd.n747 9.7499
R21583 vdd.n279 vdd.n264 9.69747
R21584 vdd.n232 vdd.n217 9.69747
R21585 vdd.n189 vdd.n174 9.69747
R21586 vdd.n142 vdd.n127 9.69747
R21587 vdd.n100 vdd.n85 9.69747
R21588 vdd.n53 vdd.n38 9.69747
R21589 vdd.n1549 vdd.n1534 9.69747
R21590 vdd.n1596 vdd.n1581 9.69747
R21591 vdd.n1459 vdd.n1444 9.69747
R21592 vdd.n1506 vdd.n1491 9.69747
R21593 vdd.n1370 vdd.n1355 9.69747
R21594 vdd.n1417 vdd.n1402 9.69747
R21595 vdd.n295 vdd.n294 9.45567
R21596 vdd.n248 vdd.n247 9.45567
R21597 vdd.n205 vdd.n204 9.45567
R21598 vdd.n158 vdd.n157 9.45567
R21599 vdd.n116 vdd.n115 9.45567
R21600 vdd.n69 vdd.n68 9.45567
R21601 vdd.n1565 vdd.n1564 9.45567
R21602 vdd.n1612 vdd.n1611 9.45567
R21603 vdd.n1475 vdd.n1474 9.45567
R21604 vdd.n1522 vdd.n1521 9.45567
R21605 vdd.n1386 vdd.n1385 9.45567
R21606 vdd.n1433 vdd.n1432 9.45567
R21607 vdd.n2051 vdd.n997 9.3005
R21608 vdd.n2050 vdd.n2049 9.3005
R21609 vdd.n1003 vdd.n1002 9.3005
R21610 vdd.n2044 vdd.n1007 9.3005
R21611 vdd.n2043 vdd.n1008 9.3005
R21612 vdd.n2042 vdd.n1009 9.3005
R21613 vdd.n1013 vdd.n1010 9.3005
R21614 vdd.n2037 vdd.n1014 9.3005
R21615 vdd.n2036 vdd.n1015 9.3005
R21616 vdd.n2035 vdd.n1016 9.3005
R21617 vdd.n1020 vdd.n1017 9.3005
R21618 vdd.n2030 vdd.n1021 9.3005
R21619 vdd.n2029 vdd.n1022 9.3005
R21620 vdd.n2028 vdd.n1023 9.3005
R21621 vdd.n1027 vdd.n1024 9.3005
R21622 vdd.n2023 vdd.n1028 9.3005
R21623 vdd.n2022 vdd.n1029 9.3005
R21624 vdd.n2021 vdd.n1030 9.3005
R21625 vdd.n1034 vdd.n1031 9.3005
R21626 vdd.n2016 vdd.n1035 9.3005
R21627 vdd.n2015 vdd.n1036 9.3005
R21628 vdd.n2014 vdd.n2013 9.3005
R21629 vdd.n2012 vdd.n1037 9.3005
R21630 vdd.n2011 vdd.n2010 9.3005
R21631 vdd.n1043 vdd.n1042 9.3005
R21632 vdd.n2005 vdd.n1047 9.3005
R21633 vdd.n2004 vdd.n1048 9.3005
R21634 vdd.n2003 vdd.n1049 9.3005
R21635 vdd.n1053 vdd.n1050 9.3005
R21636 vdd.n1998 vdd.n1054 9.3005
R21637 vdd.n1997 vdd.n1055 9.3005
R21638 vdd.n1996 vdd.n1056 9.3005
R21639 vdd.n1060 vdd.n1057 9.3005
R21640 vdd.n1991 vdd.n1061 9.3005
R21641 vdd.n1990 vdd.n1062 9.3005
R21642 vdd.n1989 vdd.n1063 9.3005
R21643 vdd.n1067 vdd.n1064 9.3005
R21644 vdd.n1984 vdd.n1068 9.3005
R21645 vdd.n2053 vdd.n2052 9.3005
R21646 vdd.n2075 vdd.n968 9.3005
R21647 vdd.n2074 vdd.n976 9.3005
R21648 vdd.n980 vdd.n977 9.3005
R21649 vdd.n2069 vdd.n981 9.3005
R21650 vdd.n2068 vdd.n982 9.3005
R21651 vdd.n2067 vdd.n983 9.3005
R21652 vdd.n987 vdd.n984 9.3005
R21653 vdd.n2062 vdd.n988 9.3005
R21654 vdd.n2061 vdd.n989 9.3005
R21655 vdd.n2060 vdd.n990 9.3005
R21656 vdd.n994 vdd.n991 9.3005
R21657 vdd.n2055 vdd.n995 9.3005
R21658 vdd.n2054 vdd.n996 9.3005
R21659 vdd.n2087 vdd.n2086 9.3005
R21660 vdd.n972 vdd.n971 9.3005
R21661 vdd.n1931 vdd.n1930 9.3005
R21662 vdd.n1932 vdd.n1345 9.3005
R21663 vdd.n1934 vdd.n1933 9.3005
R21664 vdd.n1335 vdd.n1334 9.3005
R21665 vdd.n1948 vdd.n1947 9.3005
R21666 vdd.n1949 vdd.n1333 9.3005
R21667 vdd.n1951 vdd.n1950 9.3005
R21668 vdd.n1323 vdd.n1322 9.3005
R21669 vdd.n1967 vdd.n1966 9.3005
R21670 vdd.n1968 vdd.n1321 9.3005
R21671 vdd.n1970 vdd.n1969 9.3005
R21672 vdd.n271 vdd.n270 9.3005
R21673 vdd.n266 vdd.n265 9.3005
R21674 vdd.n277 vdd.n276 9.3005
R21675 vdd.n279 vdd.n278 9.3005
R21676 vdd.n262 vdd.n261 9.3005
R21677 vdd.n285 vdd.n284 9.3005
R21678 vdd.n287 vdd.n286 9.3005
R21679 vdd.n259 vdd.n256 9.3005
R21680 vdd.n294 vdd.n293 9.3005
R21681 vdd.n224 vdd.n223 9.3005
R21682 vdd.n219 vdd.n218 9.3005
R21683 vdd.n230 vdd.n229 9.3005
R21684 vdd.n232 vdd.n231 9.3005
R21685 vdd.n215 vdd.n214 9.3005
R21686 vdd.n238 vdd.n237 9.3005
R21687 vdd.n240 vdd.n239 9.3005
R21688 vdd.n212 vdd.n209 9.3005
R21689 vdd.n247 vdd.n246 9.3005
R21690 vdd.n181 vdd.n180 9.3005
R21691 vdd.n176 vdd.n175 9.3005
R21692 vdd.n187 vdd.n186 9.3005
R21693 vdd.n189 vdd.n188 9.3005
R21694 vdd.n172 vdd.n171 9.3005
R21695 vdd.n195 vdd.n194 9.3005
R21696 vdd.n197 vdd.n196 9.3005
R21697 vdd.n169 vdd.n166 9.3005
R21698 vdd.n204 vdd.n203 9.3005
R21699 vdd.n134 vdd.n133 9.3005
R21700 vdd.n129 vdd.n128 9.3005
R21701 vdd.n140 vdd.n139 9.3005
R21702 vdd.n142 vdd.n141 9.3005
R21703 vdd.n125 vdd.n124 9.3005
R21704 vdd.n148 vdd.n147 9.3005
R21705 vdd.n150 vdd.n149 9.3005
R21706 vdd.n122 vdd.n119 9.3005
R21707 vdd.n157 vdd.n156 9.3005
R21708 vdd.n92 vdd.n91 9.3005
R21709 vdd.n87 vdd.n86 9.3005
R21710 vdd.n98 vdd.n97 9.3005
R21711 vdd.n100 vdd.n99 9.3005
R21712 vdd.n83 vdd.n82 9.3005
R21713 vdd.n106 vdd.n105 9.3005
R21714 vdd.n108 vdd.n107 9.3005
R21715 vdd.n80 vdd.n77 9.3005
R21716 vdd.n115 vdd.n114 9.3005
R21717 vdd.n45 vdd.n44 9.3005
R21718 vdd.n40 vdd.n39 9.3005
R21719 vdd.n51 vdd.n50 9.3005
R21720 vdd.n53 vdd.n52 9.3005
R21721 vdd.n36 vdd.n35 9.3005
R21722 vdd.n59 vdd.n58 9.3005
R21723 vdd.n61 vdd.n60 9.3005
R21724 vdd.n33 vdd.n30 9.3005
R21725 vdd.n68 vdd.n67 9.3005
R21726 vdd.n3030 vdd.n3029 9.3005
R21727 vdd.n3033 vdd.n555 9.3005
R21728 vdd.n3034 vdd.n554 9.3005
R21729 vdd.n3037 vdd.n553 9.3005
R21730 vdd.n3038 vdd.n552 9.3005
R21731 vdd.n3041 vdd.n551 9.3005
R21732 vdd.n3042 vdd.n550 9.3005
R21733 vdd.n3045 vdd.n549 9.3005
R21734 vdd.n3046 vdd.n548 9.3005
R21735 vdd.n3049 vdd.n547 9.3005
R21736 vdd.n3050 vdd.n546 9.3005
R21737 vdd.n3053 vdd.n545 9.3005
R21738 vdd.n3054 vdd.n544 9.3005
R21739 vdd.n3057 vdd.n543 9.3005
R21740 vdd.n3058 vdd.n542 9.3005
R21741 vdd.n3061 vdd.n541 9.3005
R21742 vdd.n3062 vdd.n540 9.3005
R21743 vdd.n3065 vdd.n539 9.3005
R21744 vdd.n3066 vdd.n538 9.3005
R21745 vdd.n3069 vdd.n537 9.3005
R21746 vdd.n3073 vdd.n3072 9.3005
R21747 vdd.n3074 vdd.n536 9.3005
R21748 vdd.n3078 vdd.n3075 9.3005
R21749 vdd.n3081 vdd.n535 9.3005
R21750 vdd.n3082 vdd.n534 9.3005
R21751 vdd.n3085 vdd.n533 9.3005
R21752 vdd.n3086 vdd.n532 9.3005
R21753 vdd.n3089 vdd.n531 9.3005
R21754 vdd.n3090 vdd.n530 9.3005
R21755 vdd.n3093 vdd.n529 9.3005
R21756 vdd.n3094 vdd.n528 9.3005
R21757 vdd.n3097 vdd.n527 9.3005
R21758 vdd.n3098 vdd.n526 9.3005
R21759 vdd.n3101 vdd.n525 9.3005
R21760 vdd.n3102 vdd.n524 9.3005
R21761 vdd.n3105 vdd.n519 9.3005
R21762 vdd.n482 vdd.n481 9.3005
R21763 vdd.n3116 vdd.n3115 9.3005
R21764 vdd.n3119 vdd.n3118 9.3005
R21765 vdd.n471 vdd.n470 9.3005
R21766 vdd.n3133 vdd.n3132 9.3005
R21767 vdd.n3134 vdd.n469 9.3005
R21768 vdd.n3136 vdd.n3135 9.3005
R21769 vdd.n460 vdd.n459 9.3005
R21770 vdd.n3149 vdd.n3148 9.3005
R21771 vdd.n3150 vdd.n458 9.3005
R21772 vdd.n3152 vdd.n3151 9.3005
R21773 vdd.n300 vdd.n298 9.3005
R21774 vdd.n3117 vdd.n480 9.3005
R21775 vdd.n3318 vdd.n3317 9.3005
R21776 vdd.n301 vdd.n299 9.3005
R21777 vdd.n3311 vdd.n310 9.3005
R21778 vdd.n3310 vdd.n311 9.3005
R21779 vdd.n3309 vdd.n312 9.3005
R21780 vdd.n320 vdd.n313 9.3005
R21781 vdd.n3303 vdd.n321 9.3005
R21782 vdd.n3302 vdd.n322 9.3005
R21783 vdd.n3301 vdd.n323 9.3005
R21784 vdd.n331 vdd.n324 9.3005
R21785 vdd.n3295 vdd.n3294 9.3005
R21786 vdd.n3291 vdd.n332 9.3005
R21787 vdd.n3290 vdd.n335 9.3005
R21788 vdd.n339 vdd.n336 9.3005
R21789 vdd.n340 vdd.n337 9.3005
R21790 vdd.n3283 vdd.n341 9.3005
R21791 vdd.n3282 vdd.n342 9.3005
R21792 vdd.n3281 vdd.n343 9.3005
R21793 vdd.n347 vdd.n344 9.3005
R21794 vdd.n3276 vdd.n348 9.3005
R21795 vdd.n3275 vdd.n349 9.3005
R21796 vdd.n3274 vdd.n350 9.3005
R21797 vdd.n354 vdd.n351 9.3005
R21798 vdd.n3269 vdd.n355 9.3005
R21799 vdd.n3268 vdd.n356 9.3005
R21800 vdd.n3267 vdd.n357 9.3005
R21801 vdd.n361 vdd.n358 9.3005
R21802 vdd.n3262 vdd.n362 9.3005
R21803 vdd.n3261 vdd.n363 9.3005
R21804 vdd.n3260 vdd.n3259 9.3005
R21805 vdd.n3258 vdd.n364 9.3005
R21806 vdd.n3257 vdd.n3256 9.3005
R21807 vdd.n370 vdd.n369 9.3005
R21808 vdd.n3251 vdd.n374 9.3005
R21809 vdd.n3250 vdd.n375 9.3005
R21810 vdd.n3249 vdd.n376 9.3005
R21811 vdd.n380 vdd.n377 9.3005
R21812 vdd.n3244 vdd.n381 9.3005
R21813 vdd.n3243 vdd.n382 9.3005
R21814 vdd.n3242 vdd.n383 9.3005
R21815 vdd.n387 vdd.n384 9.3005
R21816 vdd.n3237 vdd.n388 9.3005
R21817 vdd.n3236 vdd.n389 9.3005
R21818 vdd.n3235 vdd.n390 9.3005
R21819 vdd.n394 vdd.n391 9.3005
R21820 vdd.n3230 vdd.n395 9.3005
R21821 vdd.n3229 vdd.n396 9.3005
R21822 vdd.n3228 vdd.n397 9.3005
R21823 vdd.n401 vdd.n398 9.3005
R21824 vdd.n3223 vdd.n402 9.3005
R21825 vdd.n3222 vdd.n403 9.3005
R21826 vdd.n3221 vdd.n3220 9.3005
R21827 vdd.n3219 vdd.n404 9.3005
R21828 vdd.n3218 vdd.n3217 9.3005
R21829 vdd.n410 vdd.n409 9.3005
R21830 vdd.n3212 vdd.n414 9.3005
R21831 vdd.n3211 vdd.n415 9.3005
R21832 vdd.n3210 vdd.n416 9.3005
R21833 vdd.n420 vdd.n417 9.3005
R21834 vdd.n3205 vdd.n421 9.3005
R21835 vdd.n3204 vdd.n422 9.3005
R21836 vdd.n3203 vdd.n423 9.3005
R21837 vdd.n427 vdd.n424 9.3005
R21838 vdd.n3198 vdd.n428 9.3005
R21839 vdd.n3197 vdd.n429 9.3005
R21840 vdd.n3196 vdd.n430 9.3005
R21841 vdd.n434 vdd.n431 9.3005
R21842 vdd.n3191 vdd.n435 9.3005
R21843 vdd.n3190 vdd.n436 9.3005
R21844 vdd.n3189 vdd.n437 9.3005
R21845 vdd.n441 vdd.n438 9.3005
R21846 vdd.n3184 vdd.n442 9.3005
R21847 vdd.n3183 vdd.n443 9.3005
R21848 vdd.n3179 vdd.n3176 9.3005
R21849 vdd.n3293 vdd.n3292 9.3005
R21850 vdd.n3124 vdd.n3123 9.3005
R21851 vdd.n3125 vdd.n475 9.3005
R21852 vdd.n3127 vdd.n3126 9.3005
R21853 vdd.n465 vdd.n464 9.3005
R21854 vdd.n3141 vdd.n3140 9.3005
R21855 vdd.n3142 vdd.n463 9.3005
R21856 vdd.n3144 vdd.n3143 9.3005
R21857 vdd.n453 vdd.n452 9.3005
R21858 vdd.n3157 vdd.n3156 9.3005
R21859 vdd.n3158 vdd.n451 9.3005
R21860 vdd.n3160 vdd.n3159 9.3005
R21861 vdd.n3161 vdd.n450 9.3005
R21862 vdd.n3163 vdd.n3162 9.3005
R21863 vdd.n3164 vdd.n449 9.3005
R21864 vdd.n3166 vdd.n3165 9.3005
R21865 vdd.n3167 vdd.n447 9.3005
R21866 vdd.n3169 vdd.n3168 9.3005
R21867 vdd.n3170 vdd.n446 9.3005
R21868 vdd.n3172 vdd.n3171 9.3005
R21869 vdd.n3173 vdd.n444 9.3005
R21870 vdd.n3175 vdd.n3174 9.3005
R21871 vdd.n477 vdd.n476 9.3005
R21872 vdd.n2982 vdd.n2981 9.3005
R21873 vdd.n2987 vdd.n2980 9.3005
R21874 vdd.n2996 vdd.n572 9.3005
R21875 vdd.n2999 vdd.n571 9.3005
R21876 vdd.n3000 vdd.n570 9.3005
R21877 vdd.n3003 vdd.n569 9.3005
R21878 vdd.n3004 vdd.n568 9.3005
R21879 vdd.n3007 vdd.n567 9.3005
R21880 vdd.n3008 vdd.n566 9.3005
R21881 vdd.n3011 vdd.n565 9.3005
R21882 vdd.n3012 vdd.n564 9.3005
R21883 vdd.n3015 vdd.n563 9.3005
R21884 vdd.n3016 vdd.n562 9.3005
R21885 vdd.n3019 vdd.n561 9.3005
R21886 vdd.n3020 vdd.n560 9.3005
R21887 vdd.n3023 vdd.n559 9.3005
R21888 vdd.n3027 vdd.n3026 9.3005
R21889 vdd.n3028 vdd.n556 9.3005
R21890 vdd.n1980 vdd.n1979 9.3005
R21891 vdd.n1975 vdd.n1307 9.3005
R21892 vdd.n1888 vdd.n1887 9.3005
R21893 vdd.n1889 vdd.n1643 9.3005
R21894 vdd.n1891 vdd.n1890 9.3005
R21895 vdd.n1633 vdd.n1632 9.3005
R21896 vdd.n1905 vdd.n1904 9.3005
R21897 vdd.n1906 vdd.n1631 9.3005
R21898 vdd.n1908 vdd.n1907 9.3005
R21899 vdd.n1623 vdd.n1622 9.3005
R21900 vdd.n1923 vdd.n1922 9.3005
R21901 vdd.n1924 vdd.n1621 9.3005
R21902 vdd.n1926 vdd.n1925 9.3005
R21903 vdd.n1340 vdd.n1339 9.3005
R21904 vdd.n1939 vdd.n1938 9.3005
R21905 vdd.n1940 vdd.n1338 9.3005
R21906 vdd.n1942 vdd.n1941 9.3005
R21907 vdd.n1330 vdd.n1329 9.3005
R21908 vdd.n1956 vdd.n1955 9.3005
R21909 vdd.n1957 vdd.n1327 9.3005
R21910 vdd.n1961 vdd.n1960 9.3005
R21911 vdd.n1959 vdd.n1328 9.3005
R21912 vdd.n1958 vdd.n1318 9.3005
R21913 vdd.n1645 vdd.n1644 9.3005
R21914 vdd.n1781 vdd.n1780 9.3005
R21915 vdd.n1782 vdd.n1771 9.3005
R21916 vdd.n1784 vdd.n1783 9.3005
R21917 vdd.n1785 vdd.n1770 9.3005
R21918 vdd.n1787 vdd.n1786 9.3005
R21919 vdd.n1788 vdd.n1765 9.3005
R21920 vdd.n1790 vdd.n1789 9.3005
R21921 vdd.n1791 vdd.n1764 9.3005
R21922 vdd.n1793 vdd.n1792 9.3005
R21923 vdd.n1794 vdd.n1759 9.3005
R21924 vdd.n1796 vdd.n1795 9.3005
R21925 vdd.n1797 vdd.n1758 9.3005
R21926 vdd.n1799 vdd.n1798 9.3005
R21927 vdd.n1800 vdd.n1753 9.3005
R21928 vdd.n1802 vdd.n1801 9.3005
R21929 vdd.n1803 vdd.n1752 9.3005
R21930 vdd.n1805 vdd.n1804 9.3005
R21931 vdd.n1806 vdd.n1747 9.3005
R21932 vdd.n1808 vdd.n1807 9.3005
R21933 vdd.n1809 vdd.n1746 9.3005
R21934 vdd.n1811 vdd.n1810 9.3005
R21935 vdd.n1815 vdd.n1742 9.3005
R21936 vdd.n1817 vdd.n1816 9.3005
R21937 vdd.n1818 vdd.n1741 9.3005
R21938 vdd.n1820 vdd.n1819 9.3005
R21939 vdd.n1821 vdd.n1736 9.3005
R21940 vdd.n1823 vdd.n1822 9.3005
R21941 vdd.n1824 vdd.n1735 9.3005
R21942 vdd.n1826 vdd.n1825 9.3005
R21943 vdd.n1827 vdd.n1730 9.3005
R21944 vdd.n1829 vdd.n1828 9.3005
R21945 vdd.n1830 vdd.n1729 9.3005
R21946 vdd.n1832 vdd.n1831 9.3005
R21947 vdd.n1833 vdd.n1724 9.3005
R21948 vdd.n1835 vdd.n1834 9.3005
R21949 vdd.n1836 vdd.n1723 9.3005
R21950 vdd.n1838 vdd.n1837 9.3005
R21951 vdd.n1839 vdd.n1718 9.3005
R21952 vdd.n1841 vdd.n1840 9.3005
R21953 vdd.n1842 vdd.n1717 9.3005
R21954 vdd.n1844 vdd.n1843 9.3005
R21955 vdd.n1845 vdd.n1712 9.3005
R21956 vdd.n1847 vdd.n1846 9.3005
R21957 vdd.n1848 vdd.n1711 9.3005
R21958 vdd.n1850 vdd.n1849 9.3005
R21959 vdd.n1851 vdd.n1704 9.3005
R21960 vdd.n1853 vdd.n1852 9.3005
R21961 vdd.n1854 vdd.n1703 9.3005
R21962 vdd.n1856 vdd.n1855 9.3005
R21963 vdd.n1857 vdd.n1698 9.3005
R21964 vdd.n1859 vdd.n1858 9.3005
R21965 vdd.n1860 vdd.n1697 9.3005
R21966 vdd.n1862 vdd.n1861 9.3005
R21967 vdd.n1863 vdd.n1692 9.3005
R21968 vdd.n1865 vdd.n1864 9.3005
R21969 vdd.n1866 vdd.n1691 9.3005
R21970 vdd.n1868 vdd.n1867 9.3005
R21971 vdd.n1869 vdd.n1686 9.3005
R21972 vdd.n1871 vdd.n1870 9.3005
R21973 vdd.n1872 vdd.n1685 9.3005
R21974 vdd.n1874 vdd.n1873 9.3005
R21975 vdd.n1650 vdd.n1649 9.3005
R21976 vdd.n1880 vdd.n1879 9.3005
R21977 vdd.n1779 vdd.n1778 9.3005
R21978 vdd.n1883 vdd.n1882 9.3005
R21979 vdd.n1639 vdd.n1638 9.3005
R21980 vdd.n1897 vdd.n1896 9.3005
R21981 vdd.n1898 vdd.n1637 9.3005
R21982 vdd.n1900 vdd.n1899 9.3005
R21983 vdd.n1628 vdd.n1627 9.3005
R21984 vdd.n1914 vdd.n1913 9.3005
R21985 vdd.n1915 vdd.n1626 9.3005
R21986 vdd.n1918 vdd.n1917 9.3005
R21987 vdd.n1916 vdd.n1617 9.3005
R21988 vdd.n1881 vdd.n1648 9.3005
R21989 vdd.n1541 vdd.n1540 9.3005
R21990 vdd.n1536 vdd.n1535 9.3005
R21991 vdd.n1547 vdd.n1546 9.3005
R21992 vdd.n1549 vdd.n1548 9.3005
R21993 vdd.n1532 vdd.n1531 9.3005
R21994 vdd.n1555 vdd.n1554 9.3005
R21995 vdd.n1557 vdd.n1556 9.3005
R21996 vdd.n1529 vdd.n1526 9.3005
R21997 vdd.n1564 vdd.n1563 9.3005
R21998 vdd.n1588 vdd.n1587 9.3005
R21999 vdd.n1583 vdd.n1582 9.3005
R22000 vdd.n1594 vdd.n1593 9.3005
R22001 vdd.n1596 vdd.n1595 9.3005
R22002 vdd.n1579 vdd.n1578 9.3005
R22003 vdd.n1602 vdd.n1601 9.3005
R22004 vdd.n1604 vdd.n1603 9.3005
R22005 vdd.n1576 vdd.n1573 9.3005
R22006 vdd.n1611 vdd.n1610 9.3005
R22007 vdd.n1451 vdd.n1450 9.3005
R22008 vdd.n1446 vdd.n1445 9.3005
R22009 vdd.n1457 vdd.n1456 9.3005
R22010 vdd.n1459 vdd.n1458 9.3005
R22011 vdd.n1442 vdd.n1441 9.3005
R22012 vdd.n1465 vdd.n1464 9.3005
R22013 vdd.n1467 vdd.n1466 9.3005
R22014 vdd.n1439 vdd.n1436 9.3005
R22015 vdd.n1474 vdd.n1473 9.3005
R22016 vdd.n1498 vdd.n1497 9.3005
R22017 vdd.n1493 vdd.n1492 9.3005
R22018 vdd.n1504 vdd.n1503 9.3005
R22019 vdd.n1506 vdd.n1505 9.3005
R22020 vdd.n1489 vdd.n1488 9.3005
R22021 vdd.n1512 vdd.n1511 9.3005
R22022 vdd.n1514 vdd.n1513 9.3005
R22023 vdd.n1486 vdd.n1483 9.3005
R22024 vdd.n1521 vdd.n1520 9.3005
R22025 vdd.n1362 vdd.n1361 9.3005
R22026 vdd.n1357 vdd.n1356 9.3005
R22027 vdd.n1368 vdd.n1367 9.3005
R22028 vdd.n1370 vdd.n1369 9.3005
R22029 vdd.n1353 vdd.n1352 9.3005
R22030 vdd.n1376 vdd.n1375 9.3005
R22031 vdd.n1378 vdd.n1377 9.3005
R22032 vdd.n1350 vdd.n1347 9.3005
R22033 vdd.n1385 vdd.n1384 9.3005
R22034 vdd.n1409 vdd.n1408 9.3005
R22035 vdd.n1404 vdd.n1403 9.3005
R22036 vdd.n1415 vdd.n1414 9.3005
R22037 vdd.n1417 vdd.n1416 9.3005
R22038 vdd.n1400 vdd.n1399 9.3005
R22039 vdd.n1423 vdd.n1422 9.3005
R22040 vdd.n1425 vdd.n1424 9.3005
R22041 vdd.n1397 vdd.n1394 9.3005
R22042 vdd.n1432 vdd.n1431 9.3005
R22043 vdd.n1893 vdd.t150 8.95635
R22044 vdd.t177 vdd.n3305 8.95635
R22045 vdd.n276 vdd.n275 8.92171
R22046 vdd.n229 vdd.n228 8.92171
R22047 vdd.n186 vdd.n185 8.92171
R22048 vdd.n139 vdd.n138 8.92171
R22049 vdd.n97 vdd.n96 8.92171
R22050 vdd.n50 vdd.n49 8.92171
R22051 vdd.n1546 vdd.n1545 8.92171
R22052 vdd.n1593 vdd.n1592 8.92171
R22053 vdd.n1456 vdd.n1455 8.92171
R22054 vdd.n1503 vdd.n1502 8.92171
R22055 vdd.n1367 vdd.n1366 8.92171
R22056 vdd.n1414 vdd.n1413 8.92171
R22057 vdd.n207 vdd.n117 8.81535
R22058 vdd.n1524 vdd.n1434 8.81535
R22059 vdd.n1920 vdd.t166 8.72962
R22060 vdd.t195 vdd.n3314 8.72962
R22061 vdd.n1343 vdd.t186 8.50289
R22062 vdd.n1972 vdd.t76 8.50289
R22063 vdd.n516 vdd.t86 8.50289
R22064 vdd.n3146 vdd.t173 8.50289
R22065 vdd.n28 vdd.n14 8.42249
R22066 vdd.n3320 vdd.n3319 8.16225
R22067 vdd.n1616 vdd.n1615 8.16225
R22068 vdd.n272 vdd.n266 8.14595
R22069 vdd.n225 vdd.n219 8.14595
R22070 vdd.n182 vdd.n176 8.14595
R22071 vdd.n135 vdd.n129 8.14595
R22072 vdd.n93 vdd.n87 8.14595
R22073 vdd.n46 vdd.n40 8.14595
R22074 vdd.n1542 vdd.n1536 8.14595
R22075 vdd.n1589 vdd.n1583 8.14595
R22076 vdd.n1452 vdd.n1446 8.14595
R22077 vdd.n1499 vdd.n1493 8.14595
R22078 vdd.n1363 vdd.n1357 8.14595
R22079 vdd.n1410 vdd.n1404 8.14595
R22080 vdd.n2127 vdd.n924 7.70933
R22081 vdd.n2127 vdd.n927 7.70933
R22082 vdd.n2133 vdd.n913 7.70933
R22083 vdd.n2139 vdd.n913 7.70933
R22084 vdd.n2139 vdd.n906 7.70933
R22085 vdd.n2145 vdd.n906 7.70933
R22086 vdd.n2145 vdd.n909 7.70933
R22087 vdd.n2151 vdd.n902 7.70933
R22088 vdd.n2157 vdd.n896 7.70933
R22089 vdd.n2163 vdd.n883 7.70933
R22090 vdd.n2169 vdd.n883 7.70933
R22091 vdd.n2175 vdd.n877 7.70933
R22092 vdd.n2181 vdd.n870 7.70933
R22093 vdd.n2181 vdd.n873 7.70933
R22094 vdd.n2187 vdd.n866 7.70933
R22095 vdd.n2194 vdd.n852 7.70933
R22096 vdd.n2200 vdd.n852 7.70933
R22097 vdd.n2206 vdd.n846 7.70933
R22098 vdd.n2212 vdd.n842 7.70933
R22099 vdd.n2218 vdd.n836 7.70933
R22100 vdd.n2236 vdd.n818 7.70933
R22101 vdd.n2236 vdd.n811 7.70933
R22102 vdd.n2244 vdd.n811 7.70933
R22103 vdd.n2326 vdd.n795 7.70933
R22104 vdd.n2709 vdd.n747 7.70933
R22105 vdd.n2721 vdd.n736 7.70933
R22106 vdd.n2721 vdd.n730 7.70933
R22107 vdd.n2727 vdd.n730 7.70933
R22108 vdd.n2739 vdd.n721 7.70933
R22109 vdd.n2745 vdd.n715 7.70933
R22110 vdd.n2757 vdd.n702 7.70933
R22111 vdd.n2764 vdd.n695 7.70933
R22112 vdd.n2764 vdd.n698 7.70933
R22113 vdd.n2770 vdd.n691 7.70933
R22114 vdd.n2776 vdd.n677 7.70933
R22115 vdd.n2782 vdd.n677 7.70933
R22116 vdd.n2788 vdd.n671 7.70933
R22117 vdd.n2794 vdd.n664 7.70933
R22118 vdd.n2794 vdd.n667 7.70933
R22119 vdd.n2800 vdd.n660 7.70933
R22120 vdd.n2806 vdd.n654 7.70933
R22121 vdd.n2812 vdd.n641 7.70933
R22122 vdd.n2818 vdd.n641 7.70933
R22123 vdd.n2818 vdd.n633 7.70933
R22124 vdd.n2869 vdd.n633 7.70933
R22125 vdd.n2869 vdd.n636 7.70933
R22126 vdd.n2875 vdd.n595 7.70933
R22127 vdd.n2945 vdd.n595 7.70933
R22128 vdd.n271 vdd.n268 7.3702
R22129 vdd.n224 vdd.n221 7.3702
R22130 vdd.n181 vdd.n178 7.3702
R22131 vdd.n134 vdd.n131 7.3702
R22132 vdd.n92 vdd.n89 7.3702
R22133 vdd.n45 vdd.n42 7.3702
R22134 vdd.n1541 vdd.n1538 7.3702
R22135 vdd.n1588 vdd.n1585 7.3702
R22136 vdd.n1451 vdd.n1448 7.3702
R22137 vdd.n1498 vdd.n1495 7.3702
R22138 vdd.n1362 vdd.n1359 7.3702
R22139 vdd.n1409 vdd.n1406 7.3702
R22140 vdd.n896 vdd.t58 7.36923
R22141 vdd.n2800 vdd.t35 7.36923
R22142 vdd.n2151 vdd.t10 7.1425
R22143 vdd.n1215 vdd.t6 7.1425
R22144 vdd.n2733 vdd.t9 7.1425
R22145 vdd.n654 vdd.t19 7.1425
R22146 vdd.n1816 vdd.n1815 6.98232
R22147 vdd.n2015 vdd.n2014 6.98232
R22148 vdd.n3222 vdd.n3221 6.98232
R22149 vdd.n3033 vdd.n3030 6.98232
R22150 vdd.n1215 vdd.t7 6.80241
R22151 vdd.n2733 vdd.t53 6.80241
R22152 vdd.n1953 vdd.t170 6.68904
R22153 vdd.n3129 vdd.t182 6.68904
R22154 vdd.t152 vdd.n1342 6.46231
R22155 vdd.n2175 vdd.t17 6.46231
R22156 vdd.t22 vdd.n846 6.46231
R22157 vdd.n2757 vdd.t27 6.46231
R22158 vdd.t45 vdd.n671 6.46231
R22159 vdd.n3154 vdd.t158 6.46231
R22160 vdd.n2251 vdd.t55 6.34895
R22161 vdd.n2630 vdd.t42 6.34895
R22162 vdd.n2772 vdd.n687 6.2444
R22163 vdd.n2191 vdd.n2190 6.2444
R22164 vdd.n1911 vdd.t148 6.23558
R22165 vdd.t180 vdd.n308 6.23558
R22166 vdd.n3320 vdd.n297 6.22547
R22167 vdd.n1615 vdd.n1614 6.22547
R22168 vdd.n2212 vdd.t50 5.89549
R22169 vdd.n715 vdd.t23 5.89549
R22170 vdd.n272 vdd.n271 5.81868
R22171 vdd.n225 vdd.n224 5.81868
R22172 vdd.n182 vdd.n181 5.81868
R22173 vdd.n135 vdd.n134 5.81868
R22174 vdd.n93 vdd.n92 5.81868
R22175 vdd.n46 vdd.n45 5.81868
R22176 vdd.n1542 vdd.n1541 5.81868
R22177 vdd.n1589 vdd.n1588 5.81868
R22178 vdd.n1452 vdd.n1451 5.81868
R22179 vdd.n1499 vdd.n1498 5.81868
R22180 vdd.n1363 vdd.n1362 5.81868
R22181 vdd.n1410 vdd.n1409 5.81868
R22182 vdd.n2334 vdd.n2333 5.77611
R22183 vdd.n1139 vdd.n1138 5.77611
R22184 vdd.n2642 vdd.n2641 5.77611
R22185 vdd.n2886 vdd.n2885 5.77611
R22186 vdd.n2950 vdd.n591 5.77611
R22187 vdd.n2505 vdd.n2439 5.77611
R22188 vdd.n2259 vdd.n802 5.77611
R22189 vdd.n1275 vdd.n1107 5.77611
R22190 vdd.n1778 vdd.n1777 5.62474
R22191 vdd.n1978 vdd.n1975 5.62474
R22192 vdd.n3182 vdd.n3179 5.62474
R22193 vdd.n2985 vdd.n2982 5.62474
R22194 vdd.n2187 vdd.t37 5.55539
R22195 vdd.n691 vdd.t13 5.55539
R22196 vdd.n1635 vdd.t148 5.10193
R22197 vdd.n3307 vdd.t180 5.10193
R22198 vdd.n275 vdd.n266 5.04292
R22199 vdd.n228 vdd.n219 5.04292
R22200 vdd.n185 vdd.n176 5.04292
R22201 vdd.n138 vdd.n129 5.04292
R22202 vdd.n96 vdd.n87 5.04292
R22203 vdd.n49 vdd.n40 5.04292
R22204 vdd.n1545 vdd.n1536 5.04292
R22205 vdd.n1592 vdd.n1583 5.04292
R22206 vdd.n1455 vdd.n1446 5.04292
R22207 vdd.n1502 vdd.n1493 5.04292
R22208 vdd.n1366 vdd.n1357 5.04292
R22209 vdd.n1413 vdd.n1404 5.04292
R22210 vdd.n1928 vdd.t152 4.8752
R22211 vdd.t16 vdd.t28 4.8752
R22212 vdd.t59 vdd.t5 4.8752
R22213 vdd.t158 vdd.n304 4.8752
R22214 vdd.n2335 vdd.n2334 4.83952
R22215 vdd.n1138 vdd.n1137 4.83952
R22216 vdd.n2643 vdd.n2642 4.83952
R22217 vdd.n2887 vdd.n2886 4.83952
R22218 vdd.n591 vdd.n586 4.83952
R22219 vdd.n2502 vdd.n2439 4.83952
R22220 vdd.n2262 vdd.n802 4.83952
R22221 vdd.n1278 vdd.n1107 4.83952
R22222 vdd.n1189 vdd.t25 4.76184
R22223 vdd.n2715 vdd.t11 4.76184
R22224 vdd.n1983 vdd.n1982 4.74817
R22225 vdd.n1311 vdd.n1306 4.74817
R22226 vdd.n973 vdd.n970 4.74817
R22227 vdd.n2076 vdd.n969 4.74817
R22228 vdd.n2081 vdd.n970 4.74817
R22229 vdd.n2080 vdd.n969 4.74817
R22230 vdd.n3110 vdd.n3109 4.74817
R22231 vdd.n3107 vdd.n3106 4.74817
R22232 vdd.n3107 vdd.n521 4.74817
R22233 vdd.n3109 vdd.n518 4.74817
R22234 vdd.n2992 vdd.n573 4.74817
R22235 vdd.n2988 vdd.n574 4.74817
R22236 vdd.n2991 vdd.n574 4.74817
R22237 vdd.n2995 vdd.n573 4.74817
R22238 vdd.n1982 vdd.n1069 4.74817
R22239 vdd.n1308 vdd.n1306 4.74817
R22240 vdd.n297 vdd.n296 4.7074
R22241 vdd.n207 vdd.n206 4.7074
R22242 vdd.n1614 vdd.n1613 4.7074
R22243 vdd.n1524 vdd.n1523 4.7074
R22244 vdd.n1944 vdd.t170 4.64847
R22245 vdd.t18 vdd.n877 4.64847
R22246 vdd.n2206 vdd.t57 4.64847
R22247 vdd.t48 vdd.n702 4.64847
R22248 vdd.n2788 vdd.t44 4.64847
R22249 vdd.n3138 vdd.t182 4.64847
R22250 vdd.n866 vdd.t128 4.53511
R22251 vdd.n2770 vdd.t90 4.53511
R22252 vdd.n2133 vdd.t72 4.42174
R22253 vdd.n1189 vdd.t117 4.42174
R22254 vdd.n2715 vdd.t124 4.42174
R22255 vdd.n636 vdd.t68 4.42174
R22256 vdd.n2761 vdd.n687 4.37123
R22257 vdd.n2192 vdd.n2191 4.37123
R22258 vdd.n2230 vdd.t46 4.30838
R22259 vdd.n2618 vdd.t31 4.30838
R22260 vdd.n276 vdd.n264 4.26717
R22261 vdd.n229 vdd.n217 4.26717
R22262 vdd.n186 vdd.n174 4.26717
R22263 vdd.n139 vdd.n127 4.26717
R22264 vdd.n97 vdd.n85 4.26717
R22265 vdd.n50 vdd.n38 4.26717
R22266 vdd.n1546 vdd.n1534 4.26717
R22267 vdd.n1593 vdd.n1581 4.26717
R22268 vdd.n1456 vdd.n1444 4.26717
R22269 vdd.n1503 vdd.n1491 4.26717
R22270 vdd.n1367 vdd.n1355 4.26717
R22271 vdd.n1414 vdd.n1402 4.26717
R22272 vdd.n297 vdd.n207 4.10845
R22273 vdd.n1614 vdd.n1524 4.10845
R22274 vdd.n253 vdd.t165 4.06363
R22275 vdd.n253 vdd.t191 4.06363
R22276 vdd.n251 vdd.t202 4.06363
R22277 vdd.n251 vdd.t208 4.06363
R22278 vdd.n249 vdd.t210 4.06363
R22279 vdd.n249 vdd.t172 4.06363
R22280 vdd.n163 vdd.t155 4.06363
R22281 vdd.n163 vdd.t181 4.06363
R22282 vdd.n161 vdd.t199 4.06363
R22283 vdd.n161 vdd.t203 4.06363
R22284 vdd.n159 vdd.t207 4.06363
R22285 vdd.n159 vdd.t157 4.06363
R22286 vdd.n74 vdd.t164 4.06363
R22287 vdd.n74 vdd.t200 4.06363
R22288 vdd.n72 vdd.t159 4.06363
R22289 vdd.n72 vdd.t196 4.06363
R22290 vdd.n70 vdd.t174 4.06363
R22291 vdd.n70 vdd.t204 4.06363
R22292 vdd.n1566 vdd.t194 4.06363
R22293 vdd.n1566 vdd.t193 4.06363
R22294 vdd.n1568 vdd.t175 4.06363
R22295 vdd.n1568 vdd.t163 4.06363
R22296 vdd.n1570 vdd.t161 4.06363
R22297 vdd.n1570 vdd.t192 4.06363
R22298 vdd.n1476 vdd.t189 4.06363
R22299 vdd.n1476 vdd.t187 4.06363
R22300 vdd.n1478 vdd.t167 4.06363
R22301 vdd.n1478 vdd.t153 4.06363
R22302 vdd.n1480 vdd.t149 4.06363
R22303 vdd.n1480 vdd.t185 4.06363
R22304 vdd.n1387 vdd.t205 4.06363
R22305 vdd.n1387 vdd.t211 4.06363
R22306 vdd.n1389 vdd.t197 4.06363
R22307 vdd.n1389 vdd.t160 4.06363
R22308 vdd.n1391 vdd.t190 4.06363
R22309 vdd.n1391 vdd.t169 4.06363
R22310 vdd.n902 vdd.t52 3.96828
R22311 vdd.n2224 vdd.t30 3.96828
R22312 vdd.n2612 vdd.t49 3.96828
R22313 vdd.n2806 vdd.t36 3.96828
R22314 vdd.n26 vdd.t144 3.9605
R22315 vdd.n26 vdd.t4 3.9605
R22316 vdd.n23 vdd.t0 3.9605
R22317 vdd.n23 vdd.t1 3.9605
R22318 vdd.n21 vdd.t3 3.9605
R22319 vdd.n21 vdd.t62 3.9605
R22320 vdd.n20 vdd.t2 3.9605
R22321 vdd.n20 vdd.t64 3.9605
R22322 vdd.n15 vdd.t66 3.9605
R22323 vdd.n15 vdd.t145 3.9605
R22324 vdd.n16 vdd.t147 3.9605
R22325 vdd.n16 vdd.t63 3.9605
R22326 vdd.n18 vdd.t146 3.9605
R22327 vdd.n18 vdd.t143 3.9605
R22328 vdd.n25 vdd.t65 3.9605
R22329 vdd.n25 vdd.t61 3.9605
R22330 vdd.n2157 vdd.t52 3.74155
R22331 vdd.n836 vdd.t30 3.74155
R22332 vdd.n2739 vdd.t49 3.74155
R22333 vdd.n660 vdd.t36 3.74155
R22334 vdd.n7 vdd.t60 3.61217
R22335 vdd.n7 vdd.t24 3.61217
R22336 vdd.n8 vdd.t32 3.61217
R22337 vdd.n8 vdd.t54 3.61217
R22338 vdd.n10 vdd.t43 3.61217
R22339 vdd.n10 vdd.t12 3.61217
R22340 vdd.n12 vdd.t21 3.61217
R22341 vdd.n12 vdd.t39 3.61217
R22342 vdd.n5 vdd.t41 3.61217
R22343 vdd.n5 vdd.t34 3.61217
R22344 vdd.n3 vdd.t26 3.61217
R22345 vdd.n3 vdd.t56 3.61217
R22346 vdd.n1 vdd.t8 3.61217
R22347 vdd.n1 vdd.t47 3.61217
R22348 vdd.n0 vdd.t51 3.61217
R22349 vdd.n0 vdd.t29 3.61217
R22350 vdd.n280 vdd.n279 3.49141
R22351 vdd.n233 vdd.n232 3.49141
R22352 vdd.n190 vdd.n189 3.49141
R22353 vdd.n143 vdd.n142 3.49141
R22354 vdd.n101 vdd.n100 3.49141
R22355 vdd.n54 vdd.n53 3.49141
R22356 vdd.n1550 vdd.n1549 3.49141
R22357 vdd.n1597 vdd.n1596 3.49141
R22358 vdd.n1460 vdd.n1459 3.49141
R22359 vdd.n1507 vdd.n1506 3.49141
R22360 vdd.n1371 vdd.n1370 3.49141
R22361 vdd.n1418 vdd.n1417 3.49141
R22362 vdd.t46 vdd.n818 3.40145
R22363 vdd.n2398 vdd.t40 3.40145
R22364 vdd.n2702 vdd.t38 3.40145
R22365 vdd.n2727 vdd.t31 3.40145
R22366 vdd.n927 vdd.t72 3.28809
R22367 vdd.n2251 vdd.t117 3.28809
R22368 vdd.n2630 vdd.t124 3.28809
R22369 vdd.n2875 vdd.t68 3.28809
R22370 vdd.n2169 vdd.t18 3.06136
R22371 vdd.n1227 vdd.t57 3.06136
R22372 vdd.n2751 vdd.t48 3.06136
R22373 vdd.t44 vdd.n664 3.06136
R22374 vdd.n2244 vdd.t25 2.94799
R22375 vdd.t11 vdd.n736 2.94799
R22376 vdd.n1945 vdd.t186 2.83463
R22377 vdd.n1963 vdd.t76 2.83463
R22378 vdd.n3121 vdd.t86 2.83463
R22379 vdd.n467 vdd.t173 2.83463
R22380 vdd.n283 vdd.n262 2.71565
R22381 vdd.n236 vdd.n215 2.71565
R22382 vdd.n193 vdd.n172 2.71565
R22383 vdd.n146 vdd.n125 2.71565
R22384 vdd.n104 vdd.n83 2.71565
R22385 vdd.n57 vdd.n36 2.71565
R22386 vdd.n1553 vdd.n1532 2.71565
R22387 vdd.n1600 vdd.n1579 2.71565
R22388 vdd.n1463 vdd.n1442 2.71565
R22389 vdd.n1510 vdd.n1489 2.71565
R22390 vdd.n1374 vdd.n1353 2.71565
R22391 vdd.n1421 vdd.n1400 2.71565
R22392 vdd.t166 vdd.n1619 2.6079
R22393 vdd.n3315 vdd.t195 2.6079
R22394 vdd.n2218 vdd.t28 2.49453
R22395 vdd.n721 vdd.t59 2.49453
R22396 vdd.n270 vdd.n269 2.4129
R22397 vdd.n223 vdd.n222 2.4129
R22398 vdd.n180 vdd.n179 2.4129
R22399 vdd.n133 vdd.n132 2.4129
R22400 vdd.n91 vdd.n90 2.4129
R22401 vdd.n44 vdd.n43 2.4129
R22402 vdd.n1540 vdd.n1539 2.4129
R22403 vdd.n1587 vdd.n1586 2.4129
R22404 vdd.n1450 vdd.n1449 2.4129
R22405 vdd.n1497 vdd.n1496 2.4129
R22406 vdd.n1361 vdd.n1360 2.4129
R22407 vdd.n1408 vdd.n1407 2.4129
R22408 vdd.n1902 vdd.t150 2.38117
R22409 vdd.n3306 vdd.t177 2.38117
R22410 vdd.n2088 vdd.n970 2.27742
R22411 vdd.n2088 vdd.n969 2.27742
R22412 vdd.n3108 vdd.n3107 2.27742
R22413 vdd.n3109 vdd.n3108 2.27742
R22414 vdd.n2979 vdd.n574 2.27742
R22415 vdd.n2979 vdd.n573 2.27742
R22416 vdd.n1982 vdd.n1981 2.27742
R22417 vdd.n1981 vdd.n1306 2.27742
R22418 vdd.n873 vdd.t37 2.15444
R22419 vdd.n2194 vdd.t15 2.15444
R22420 vdd.n698 vdd.t14 2.15444
R22421 vdd.n2776 vdd.t13 2.15444
R22422 vdd.n284 vdd.n260 1.93989
R22423 vdd.n237 vdd.n213 1.93989
R22424 vdd.n194 vdd.n170 1.93989
R22425 vdd.n147 vdd.n123 1.93989
R22426 vdd.n105 vdd.n81 1.93989
R22427 vdd.n58 vdd.n34 1.93989
R22428 vdd.n1554 vdd.n1530 1.93989
R22429 vdd.n1601 vdd.n1577 1.93989
R22430 vdd.n1464 vdd.n1440 1.93989
R22431 vdd.n1511 vdd.n1487 1.93989
R22432 vdd.n1375 vdd.n1351 1.93989
R22433 vdd.n1422 vdd.n1398 1.93989
R22434 vdd.n1227 vdd.t50 1.81434
R22435 vdd.n2751 vdd.t23 1.81434
R22436 vdd.t55 vdd.n795 1.36088
R22437 vdd.n2709 vdd.t42 1.36088
R22438 vdd.n1910 vdd.t168 1.24752
R22439 vdd.t17 vdd.n870 1.24752
R22440 vdd.n2200 vdd.t22 1.24752
R22441 vdd.t27 vdd.n695 1.24752
R22442 vdd.n2782 vdd.t45 1.24752
R22443 vdd.t154 vdd.n3313 1.24752
R22444 vdd.n295 vdd.n255 1.16414
R22445 vdd.n288 vdd.n287 1.16414
R22446 vdd.n248 vdd.n208 1.16414
R22447 vdd.n241 vdd.n240 1.16414
R22448 vdd.n205 vdd.n165 1.16414
R22449 vdd.n198 vdd.n197 1.16414
R22450 vdd.n158 vdd.n118 1.16414
R22451 vdd.n151 vdd.n150 1.16414
R22452 vdd.n116 vdd.n76 1.16414
R22453 vdd.n109 vdd.n108 1.16414
R22454 vdd.n69 vdd.n29 1.16414
R22455 vdd.n62 vdd.n61 1.16414
R22456 vdd.n1565 vdd.n1525 1.16414
R22457 vdd.n1558 vdd.n1557 1.16414
R22458 vdd.n1612 vdd.n1572 1.16414
R22459 vdd.n1605 vdd.n1604 1.16414
R22460 vdd.n1475 vdd.n1435 1.16414
R22461 vdd.n1468 vdd.n1467 1.16414
R22462 vdd.n1522 vdd.n1482 1.16414
R22463 vdd.n1515 vdd.n1514 1.16414
R22464 vdd.n1386 vdd.n1346 1.16414
R22465 vdd.n1379 vdd.n1378 1.16414
R22466 vdd.n1433 vdd.n1393 1.16414
R22467 vdd.n1426 vdd.n1425 1.16414
R22468 vdd.n1615 vdd.n28 1.06035
R22469 vdd vdd.n3320 1.05252
R22470 vdd.n1936 vdd.t188 1.02079
R22471 vdd.t128 vdd.t15 1.02079
R22472 vdd.t14 vdd.t90 1.02079
R22473 vdd.t156 vdd.n456 1.02079
R22474 vdd.n1781 vdd.n1777 0.970197
R22475 vdd.n1979 vdd.n1978 0.970197
R22476 vdd.n3183 vdd.n3182 0.970197
R22477 vdd.n2987 vdd.n2985 0.970197
R22478 vdd.n2224 vdd.t7 0.907421
R22479 vdd.n2612 vdd.t53 0.907421
R22480 vdd.n1885 vdd.t94 0.567326
R22481 vdd.n909 vdd.t10 0.567326
R22482 vdd.n2230 vdd.t6 0.567326
R22483 vdd.n2618 vdd.t9 0.567326
R22484 vdd.n2812 vdd.t19 0.567326
R22485 vdd.n3298 vdd.t101 0.567326
R22486 vdd.n1969 vdd.n971 0.537085
R22487 vdd.n3117 vdd.n3116 0.537085
R22488 vdd.n3294 vdd.n3293 0.537085
R22489 vdd.n3176 vdd.n3175 0.537085
R22490 vdd.n2981 vdd.n476 0.537085
R22491 vdd.n1958 vdd.n1307 0.537085
R22492 vdd.n1779 vdd.n1644 0.537085
R22493 vdd.n1881 vdd.n1880 0.537085
R22494 vdd.n4 vdd.n2 0.459552
R22495 vdd.n11 vdd.n9 0.459552
R22496 vdd.n293 vdd.n292 0.388379
R22497 vdd.n259 vdd.n257 0.388379
R22498 vdd.n246 vdd.n245 0.388379
R22499 vdd.n212 vdd.n210 0.388379
R22500 vdd.n203 vdd.n202 0.388379
R22501 vdd.n169 vdd.n167 0.388379
R22502 vdd.n156 vdd.n155 0.388379
R22503 vdd.n122 vdd.n120 0.388379
R22504 vdd.n114 vdd.n113 0.388379
R22505 vdd.n80 vdd.n78 0.388379
R22506 vdd.n67 vdd.n66 0.388379
R22507 vdd.n33 vdd.n31 0.388379
R22508 vdd.n1563 vdd.n1562 0.388379
R22509 vdd.n1529 vdd.n1527 0.388379
R22510 vdd.n1610 vdd.n1609 0.388379
R22511 vdd.n1576 vdd.n1574 0.388379
R22512 vdd.n1473 vdd.n1472 0.388379
R22513 vdd.n1439 vdd.n1437 0.388379
R22514 vdd.n1520 vdd.n1519 0.388379
R22515 vdd.n1486 vdd.n1484 0.388379
R22516 vdd.n1384 vdd.n1383 0.388379
R22517 vdd.n1350 vdd.n1348 0.388379
R22518 vdd.n1431 vdd.n1430 0.388379
R22519 vdd.n1397 vdd.n1395 0.388379
R22520 vdd.n19 vdd.n17 0.387128
R22521 vdd.n24 vdd.n22 0.387128
R22522 vdd.n6 vdd.n4 0.358259
R22523 vdd.n13 vdd.n11 0.358259
R22524 vdd.n252 vdd.n250 0.358259
R22525 vdd.n254 vdd.n252 0.358259
R22526 vdd.n296 vdd.n254 0.358259
R22527 vdd.n162 vdd.n160 0.358259
R22528 vdd.n164 vdd.n162 0.358259
R22529 vdd.n206 vdd.n164 0.358259
R22530 vdd.n73 vdd.n71 0.358259
R22531 vdd.n75 vdd.n73 0.358259
R22532 vdd.n117 vdd.n75 0.358259
R22533 vdd.n1613 vdd.n1571 0.358259
R22534 vdd.n1571 vdd.n1569 0.358259
R22535 vdd.n1569 vdd.n1567 0.358259
R22536 vdd.n1523 vdd.n1481 0.358259
R22537 vdd.n1481 vdd.n1479 0.358259
R22538 vdd.n1479 vdd.n1477 0.358259
R22539 vdd.n1434 vdd.n1392 0.358259
R22540 vdd.n1392 vdd.n1390 0.358259
R22541 vdd.n1390 vdd.n1388 0.358259
R22542 vdd.n2163 vdd.t58 0.340595
R22543 vdd.n842 vdd.t16 0.340595
R22544 vdd.n2745 vdd.t5 0.340595
R22545 vdd.n667 vdd.t35 0.340595
R22546 vdd.n14 vdd.n6 0.334552
R22547 vdd.n14 vdd.n13 0.334552
R22548 vdd.n27 vdd.n19 0.21707
R22549 vdd.n27 vdd.n24 0.21707
R22550 vdd.n294 vdd.n256 0.155672
R22551 vdd.n286 vdd.n256 0.155672
R22552 vdd.n286 vdd.n285 0.155672
R22553 vdd.n285 vdd.n261 0.155672
R22554 vdd.n278 vdd.n261 0.155672
R22555 vdd.n278 vdd.n277 0.155672
R22556 vdd.n277 vdd.n265 0.155672
R22557 vdd.n270 vdd.n265 0.155672
R22558 vdd.n247 vdd.n209 0.155672
R22559 vdd.n239 vdd.n209 0.155672
R22560 vdd.n239 vdd.n238 0.155672
R22561 vdd.n238 vdd.n214 0.155672
R22562 vdd.n231 vdd.n214 0.155672
R22563 vdd.n231 vdd.n230 0.155672
R22564 vdd.n230 vdd.n218 0.155672
R22565 vdd.n223 vdd.n218 0.155672
R22566 vdd.n204 vdd.n166 0.155672
R22567 vdd.n196 vdd.n166 0.155672
R22568 vdd.n196 vdd.n195 0.155672
R22569 vdd.n195 vdd.n171 0.155672
R22570 vdd.n188 vdd.n171 0.155672
R22571 vdd.n188 vdd.n187 0.155672
R22572 vdd.n187 vdd.n175 0.155672
R22573 vdd.n180 vdd.n175 0.155672
R22574 vdd.n157 vdd.n119 0.155672
R22575 vdd.n149 vdd.n119 0.155672
R22576 vdd.n149 vdd.n148 0.155672
R22577 vdd.n148 vdd.n124 0.155672
R22578 vdd.n141 vdd.n124 0.155672
R22579 vdd.n141 vdd.n140 0.155672
R22580 vdd.n140 vdd.n128 0.155672
R22581 vdd.n133 vdd.n128 0.155672
R22582 vdd.n115 vdd.n77 0.155672
R22583 vdd.n107 vdd.n77 0.155672
R22584 vdd.n107 vdd.n106 0.155672
R22585 vdd.n106 vdd.n82 0.155672
R22586 vdd.n99 vdd.n82 0.155672
R22587 vdd.n99 vdd.n98 0.155672
R22588 vdd.n98 vdd.n86 0.155672
R22589 vdd.n91 vdd.n86 0.155672
R22590 vdd.n68 vdd.n30 0.155672
R22591 vdd.n60 vdd.n30 0.155672
R22592 vdd.n60 vdd.n59 0.155672
R22593 vdd.n59 vdd.n35 0.155672
R22594 vdd.n52 vdd.n35 0.155672
R22595 vdd.n52 vdd.n51 0.155672
R22596 vdd.n51 vdd.n39 0.155672
R22597 vdd.n44 vdd.n39 0.155672
R22598 vdd.n1564 vdd.n1526 0.155672
R22599 vdd.n1556 vdd.n1526 0.155672
R22600 vdd.n1556 vdd.n1555 0.155672
R22601 vdd.n1555 vdd.n1531 0.155672
R22602 vdd.n1548 vdd.n1531 0.155672
R22603 vdd.n1548 vdd.n1547 0.155672
R22604 vdd.n1547 vdd.n1535 0.155672
R22605 vdd.n1540 vdd.n1535 0.155672
R22606 vdd.n1611 vdd.n1573 0.155672
R22607 vdd.n1603 vdd.n1573 0.155672
R22608 vdd.n1603 vdd.n1602 0.155672
R22609 vdd.n1602 vdd.n1578 0.155672
R22610 vdd.n1595 vdd.n1578 0.155672
R22611 vdd.n1595 vdd.n1594 0.155672
R22612 vdd.n1594 vdd.n1582 0.155672
R22613 vdd.n1587 vdd.n1582 0.155672
R22614 vdd.n1474 vdd.n1436 0.155672
R22615 vdd.n1466 vdd.n1436 0.155672
R22616 vdd.n1466 vdd.n1465 0.155672
R22617 vdd.n1465 vdd.n1441 0.155672
R22618 vdd.n1458 vdd.n1441 0.155672
R22619 vdd.n1458 vdd.n1457 0.155672
R22620 vdd.n1457 vdd.n1445 0.155672
R22621 vdd.n1450 vdd.n1445 0.155672
R22622 vdd.n1521 vdd.n1483 0.155672
R22623 vdd.n1513 vdd.n1483 0.155672
R22624 vdd.n1513 vdd.n1512 0.155672
R22625 vdd.n1512 vdd.n1488 0.155672
R22626 vdd.n1505 vdd.n1488 0.155672
R22627 vdd.n1505 vdd.n1504 0.155672
R22628 vdd.n1504 vdd.n1492 0.155672
R22629 vdd.n1497 vdd.n1492 0.155672
R22630 vdd.n1385 vdd.n1347 0.155672
R22631 vdd.n1377 vdd.n1347 0.155672
R22632 vdd.n1377 vdd.n1376 0.155672
R22633 vdd.n1376 vdd.n1352 0.155672
R22634 vdd.n1369 vdd.n1352 0.155672
R22635 vdd.n1369 vdd.n1368 0.155672
R22636 vdd.n1368 vdd.n1356 0.155672
R22637 vdd.n1361 vdd.n1356 0.155672
R22638 vdd.n1432 vdd.n1394 0.155672
R22639 vdd.n1424 vdd.n1394 0.155672
R22640 vdd.n1424 vdd.n1423 0.155672
R22641 vdd.n1423 vdd.n1399 0.155672
R22642 vdd.n1416 vdd.n1399 0.155672
R22643 vdd.n1416 vdd.n1415 0.155672
R22644 vdd.n1415 vdd.n1403 0.155672
R22645 vdd.n1408 vdd.n1403 0.155672
R22646 vdd.n976 vdd.n968 0.152939
R22647 vdd.n980 vdd.n976 0.152939
R22648 vdd.n981 vdd.n980 0.152939
R22649 vdd.n982 vdd.n981 0.152939
R22650 vdd.n983 vdd.n982 0.152939
R22651 vdd.n987 vdd.n983 0.152939
R22652 vdd.n988 vdd.n987 0.152939
R22653 vdd.n989 vdd.n988 0.152939
R22654 vdd.n990 vdd.n989 0.152939
R22655 vdd.n994 vdd.n990 0.152939
R22656 vdd.n995 vdd.n994 0.152939
R22657 vdd.n996 vdd.n995 0.152939
R22658 vdd.n2052 vdd.n996 0.152939
R22659 vdd.n2052 vdd.n2051 0.152939
R22660 vdd.n2051 vdd.n2050 0.152939
R22661 vdd.n2050 vdd.n1002 0.152939
R22662 vdd.n1007 vdd.n1002 0.152939
R22663 vdd.n1008 vdd.n1007 0.152939
R22664 vdd.n1009 vdd.n1008 0.152939
R22665 vdd.n1013 vdd.n1009 0.152939
R22666 vdd.n1014 vdd.n1013 0.152939
R22667 vdd.n1015 vdd.n1014 0.152939
R22668 vdd.n1016 vdd.n1015 0.152939
R22669 vdd.n1020 vdd.n1016 0.152939
R22670 vdd.n1021 vdd.n1020 0.152939
R22671 vdd.n1022 vdd.n1021 0.152939
R22672 vdd.n1023 vdd.n1022 0.152939
R22673 vdd.n1027 vdd.n1023 0.152939
R22674 vdd.n1028 vdd.n1027 0.152939
R22675 vdd.n1029 vdd.n1028 0.152939
R22676 vdd.n1030 vdd.n1029 0.152939
R22677 vdd.n1034 vdd.n1030 0.152939
R22678 vdd.n1035 vdd.n1034 0.152939
R22679 vdd.n1036 vdd.n1035 0.152939
R22680 vdd.n2013 vdd.n1036 0.152939
R22681 vdd.n2013 vdd.n2012 0.152939
R22682 vdd.n2012 vdd.n2011 0.152939
R22683 vdd.n2011 vdd.n1042 0.152939
R22684 vdd.n1047 vdd.n1042 0.152939
R22685 vdd.n1048 vdd.n1047 0.152939
R22686 vdd.n1049 vdd.n1048 0.152939
R22687 vdd.n1053 vdd.n1049 0.152939
R22688 vdd.n1054 vdd.n1053 0.152939
R22689 vdd.n1055 vdd.n1054 0.152939
R22690 vdd.n1056 vdd.n1055 0.152939
R22691 vdd.n1060 vdd.n1056 0.152939
R22692 vdd.n1061 vdd.n1060 0.152939
R22693 vdd.n1062 vdd.n1061 0.152939
R22694 vdd.n1063 vdd.n1062 0.152939
R22695 vdd.n1067 vdd.n1063 0.152939
R22696 vdd.n1068 vdd.n1067 0.152939
R22697 vdd.n2087 vdd.n971 0.152939
R22698 vdd.n1932 vdd.n1931 0.152939
R22699 vdd.n1933 vdd.n1932 0.152939
R22700 vdd.n1933 vdd.n1334 0.152939
R22701 vdd.n1948 vdd.n1334 0.152939
R22702 vdd.n1949 vdd.n1948 0.152939
R22703 vdd.n1950 vdd.n1949 0.152939
R22704 vdd.n1950 vdd.n1322 0.152939
R22705 vdd.n1967 vdd.n1322 0.152939
R22706 vdd.n1968 vdd.n1967 0.152939
R22707 vdd.n1969 vdd.n1968 0.152939
R22708 vdd.n524 vdd.n519 0.152939
R22709 vdd.n525 vdd.n524 0.152939
R22710 vdd.n526 vdd.n525 0.152939
R22711 vdd.n527 vdd.n526 0.152939
R22712 vdd.n528 vdd.n527 0.152939
R22713 vdd.n529 vdd.n528 0.152939
R22714 vdd.n530 vdd.n529 0.152939
R22715 vdd.n531 vdd.n530 0.152939
R22716 vdd.n532 vdd.n531 0.152939
R22717 vdd.n533 vdd.n532 0.152939
R22718 vdd.n534 vdd.n533 0.152939
R22719 vdd.n535 vdd.n534 0.152939
R22720 vdd.n3075 vdd.n535 0.152939
R22721 vdd.n3075 vdd.n3074 0.152939
R22722 vdd.n3074 vdd.n3073 0.152939
R22723 vdd.n3073 vdd.n537 0.152939
R22724 vdd.n538 vdd.n537 0.152939
R22725 vdd.n539 vdd.n538 0.152939
R22726 vdd.n540 vdd.n539 0.152939
R22727 vdd.n541 vdd.n540 0.152939
R22728 vdd.n542 vdd.n541 0.152939
R22729 vdd.n543 vdd.n542 0.152939
R22730 vdd.n544 vdd.n543 0.152939
R22731 vdd.n545 vdd.n544 0.152939
R22732 vdd.n546 vdd.n545 0.152939
R22733 vdd.n547 vdd.n546 0.152939
R22734 vdd.n548 vdd.n547 0.152939
R22735 vdd.n549 vdd.n548 0.152939
R22736 vdd.n550 vdd.n549 0.152939
R22737 vdd.n551 vdd.n550 0.152939
R22738 vdd.n552 vdd.n551 0.152939
R22739 vdd.n553 vdd.n552 0.152939
R22740 vdd.n554 vdd.n553 0.152939
R22741 vdd.n555 vdd.n554 0.152939
R22742 vdd.n3029 vdd.n555 0.152939
R22743 vdd.n3029 vdd.n3028 0.152939
R22744 vdd.n3028 vdd.n3027 0.152939
R22745 vdd.n3027 vdd.n559 0.152939
R22746 vdd.n560 vdd.n559 0.152939
R22747 vdd.n561 vdd.n560 0.152939
R22748 vdd.n562 vdd.n561 0.152939
R22749 vdd.n563 vdd.n562 0.152939
R22750 vdd.n564 vdd.n563 0.152939
R22751 vdd.n565 vdd.n564 0.152939
R22752 vdd.n566 vdd.n565 0.152939
R22753 vdd.n567 vdd.n566 0.152939
R22754 vdd.n568 vdd.n567 0.152939
R22755 vdd.n569 vdd.n568 0.152939
R22756 vdd.n570 vdd.n569 0.152939
R22757 vdd.n571 vdd.n570 0.152939
R22758 vdd.n572 vdd.n571 0.152939
R22759 vdd.n3116 vdd.n481 0.152939
R22760 vdd.n3118 vdd.n3117 0.152939
R22761 vdd.n3118 vdd.n470 0.152939
R22762 vdd.n3133 vdd.n470 0.152939
R22763 vdd.n3134 vdd.n3133 0.152939
R22764 vdd.n3135 vdd.n3134 0.152939
R22765 vdd.n3135 vdd.n459 0.152939
R22766 vdd.n3149 vdd.n459 0.152939
R22767 vdd.n3150 vdd.n3149 0.152939
R22768 vdd.n3151 vdd.n3150 0.152939
R22769 vdd.n3151 vdd.n298 0.152939
R22770 vdd.n3318 vdd.n299 0.152939
R22771 vdd.n310 vdd.n299 0.152939
R22772 vdd.n311 vdd.n310 0.152939
R22773 vdd.n312 vdd.n311 0.152939
R22774 vdd.n320 vdd.n312 0.152939
R22775 vdd.n321 vdd.n320 0.152939
R22776 vdd.n322 vdd.n321 0.152939
R22777 vdd.n323 vdd.n322 0.152939
R22778 vdd.n331 vdd.n323 0.152939
R22779 vdd.n3294 vdd.n331 0.152939
R22780 vdd.n3293 vdd.n332 0.152939
R22781 vdd.n335 vdd.n332 0.152939
R22782 vdd.n339 vdd.n335 0.152939
R22783 vdd.n340 vdd.n339 0.152939
R22784 vdd.n341 vdd.n340 0.152939
R22785 vdd.n342 vdd.n341 0.152939
R22786 vdd.n343 vdd.n342 0.152939
R22787 vdd.n347 vdd.n343 0.152939
R22788 vdd.n348 vdd.n347 0.152939
R22789 vdd.n349 vdd.n348 0.152939
R22790 vdd.n350 vdd.n349 0.152939
R22791 vdd.n354 vdd.n350 0.152939
R22792 vdd.n355 vdd.n354 0.152939
R22793 vdd.n356 vdd.n355 0.152939
R22794 vdd.n357 vdd.n356 0.152939
R22795 vdd.n361 vdd.n357 0.152939
R22796 vdd.n362 vdd.n361 0.152939
R22797 vdd.n363 vdd.n362 0.152939
R22798 vdd.n3259 vdd.n363 0.152939
R22799 vdd.n3259 vdd.n3258 0.152939
R22800 vdd.n3258 vdd.n3257 0.152939
R22801 vdd.n3257 vdd.n369 0.152939
R22802 vdd.n374 vdd.n369 0.152939
R22803 vdd.n375 vdd.n374 0.152939
R22804 vdd.n376 vdd.n375 0.152939
R22805 vdd.n380 vdd.n376 0.152939
R22806 vdd.n381 vdd.n380 0.152939
R22807 vdd.n382 vdd.n381 0.152939
R22808 vdd.n383 vdd.n382 0.152939
R22809 vdd.n387 vdd.n383 0.152939
R22810 vdd.n388 vdd.n387 0.152939
R22811 vdd.n389 vdd.n388 0.152939
R22812 vdd.n390 vdd.n389 0.152939
R22813 vdd.n394 vdd.n390 0.152939
R22814 vdd.n395 vdd.n394 0.152939
R22815 vdd.n396 vdd.n395 0.152939
R22816 vdd.n397 vdd.n396 0.152939
R22817 vdd.n401 vdd.n397 0.152939
R22818 vdd.n402 vdd.n401 0.152939
R22819 vdd.n403 vdd.n402 0.152939
R22820 vdd.n3220 vdd.n403 0.152939
R22821 vdd.n3220 vdd.n3219 0.152939
R22822 vdd.n3219 vdd.n3218 0.152939
R22823 vdd.n3218 vdd.n409 0.152939
R22824 vdd.n414 vdd.n409 0.152939
R22825 vdd.n415 vdd.n414 0.152939
R22826 vdd.n416 vdd.n415 0.152939
R22827 vdd.n420 vdd.n416 0.152939
R22828 vdd.n421 vdd.n420 0.152939
R22829 vdd.n422 vdd.n421 0.152939
R22830 vdd.n423 vdd.n422 0.152939
R22831 vdd.n427 vdd.n423 0.152939
R22832 vdd.n428 vdd.n427 0.152939
R22833 vdd.n429 vdd.n428 0.152939
R22834 vdd.n430 vdd.n429 0.152939
R22835 vdd.n434 vdd.n430 0.152939
R22836 vdd.n435 vdd.n434 0.152939
R22837 vdd.n436 vdd.n435 0.152939
R22838 vdd.n437 vdd.n436 0.152939
R22839 vdd.n441 vdd.n437 0.152939
R22840 vdd.n442 vdd.n441 0.152939
R22841 vdd.n443 vdd.n442 0.152939
R22842 vdd.n3176 vdd.n443 0.152939
R22843 vdd.n3124 vdd.n476 0.152939
R22844 vdd.n3125 vdd.n3124 0.152939
R22845 vdd.n3126 vdd.n3125 0.152939
R22846 vdd.n3126 vdd.n464 0.152939
R22847 vdd.n3141 vdd.n464 0.152939
R22848 vdd.n3142 vdd.n3141 0.152939
R22849 vdd.n3143 vdd.n3142 0.152939
R22850 vdd.n3143 vdd.n452 0.152939
R22851 vdd.n3157 vdd.n452 0.152939
R22852 vdd.n3158 vdd.n3157 0.152939
R22853 vdd.n3159 vdd.n3158 0.152939
R22854 vdd.n3159 vdd.n450 0.152939
R22855 vdd.n3163 vdd.n450 0.152939
R22856 vdd.n3164 vdd.n3163 0.152939
R22857 vdd.n3165 vdd.n3164 0.152939
R22858 vdd.n3165 vdd.n447 0.152939
R22859 vdd.n3169 vdd.n447 0.152939
R22860 vdd.n3170 vdd.n3169 0.152939
R22861 vdd.n3171 vdd.n3170 0.152939
R22862 vdd.n3171 vdd.n444 0.152939
R22863 vdd.n3175 vdd.n444 0.152939
R22864 vdd.n2981 vdd.n2980 0.152939
R22865 vdd.n1980 vdd.n1307 0.152939
R22866 vdd.n1888 vdd.n1644 0.152939
R22867 vdd.n1889 vdd.n1888 0.152939
R22868 vdd.n1890 vdd.n1889 0.152939
R22869 vdd.n1890 vdd.n1632 0.152939
R22870 vdd.n1905 vdd.n1632 0.152939
R22871 vdd.n1906 vdd.n1905 0.152939
R22872 vdd.n1907 vdd.n1906 0.152939
R22873 vdd.n1907 vdd.n1622 0.152939
R22874 vdd.n1923 vdd.n1622 0.152939
R22875 vdd.n1924 vdd.n1923 0.152939
R22876 vdd.n1925 vdd.n1924 0.152939
R22877 vdd.n1925 vdd.n1339 0.152939
R22878 vdd.n1939 vdd.n1339 0.152939
R22879 vdd.n1940 vdd.n1939 0.152939
R22880 vdd.n1941 vdd.n1940 0.152939
R22881 vdd.n1941 vdd.n1329 0.152939
R22882 vdd.n1956 vdd.n1329 0.152939
R22883 vdd.n1957 vdd.n1956 0.152939
R22884 vdd.n1960 vdd.n1957 0.152939
R22885 vdd.n1960 vdd.n1959 0.152939
R22886 vdd.n1959 vdd.n1958 0.152939
R22887 vdd.n1880 vdd.n1649 0.152939
R22888 vdd.n1873 vdd.n1649 0.152939
R22889 vdd.n1873 vdd.n1872 0.152939
R22890 vdd.n1872 vdd.n1871 0.152939
R22891 vdd.n1871 vdd.n1686 0.152939
R22892 vdd.n1867 vdd.n1686 0.152939
R22893 vdd.n1867 vdd.n1866 0.152939
R22894 vdd.n1866 vdd.n1865 0.152939
R22895 vdd.n1865 vdd.n1692 0.152939
R22896 vdd.n1861 vdd.n1692 0.152939
R22897 vdd.n1861 vdd.n1860 0.152939
R22898 vdd.n1860 vdd.n1859 0.152939
R22899 vdd.n1859 vdd.n1698 0.152939
R22900 vdd.n1855 vdd.n1698 0.152939
R22901 vdd.n1855 vdd.n1854 0.152939
R22902 vdd.n1854 vdd.n1853 0.152939
R22903 vdd.n1853 vdd.n1704 0.152939
R22904 vdd.n1849 vdd.n1704 0.152939
R22905 vdd.n1849 vdd.n1848 0.152939
R22906 vdd.n1848 vdd.n1847 0.152939
R22907 vdd.n1847 vdd.n1712 0.152939
R22908 vdd.n1843 vdd.n1712 0.152939
R22909 vdd.n1843 vdd.n1842 0.152939
R22910 vdd.n1842 vdd.n1841 0.152939
R22911 vdd.n1841 vdd.n1718 0.152939
R22912 vdd.n1837 vdd.n1718 0.152939
R22913 vdd.n1837 vdd.n1836 0.152939
R22914 vdd.n1836 vdd.n1835 0.152939
R22915 vdd.n1835 vdd.n1724 0.152939
R22916 vdd.n1831 vdd.n1724 0.152939
R22917 vdd.n1831 vdd.n1830 0.152939
R22918 vdd.n1830 vdd.n1829 0.152939
R22919 vdd.n1829 vdd.n1730 0.152939
R22920 vdd.n1825 vdd.n1730 0.152939
R22921 vdd.n1825 vdd.n1824 0.152939
R22922 vdd.n1824 vdd.n1823 0.152939
R22923 vdd.n1823 vdd.n1736 0.152939
R22924 vdd.n1819 vdd.n1736 0.152939
R22925 vdd.n1819 vdd.n1818 0.152939
R22926 vdd.n1818 vdd.n1817 0.152939
R22927 vdd.n1817 vdd.n1742 0.152939
R22928 vdd.n1810 vdd.n1742 0.152939
R22929 vdd.n1810 vdd.n1809 0.152939
R22930 vdd.n1809 vdd.n1808 0.152939
R22931 vdd.n1808 vdd.n1747 0.152939
R22932 vdd.n1804 vdd.n1747 0.152939
R22933 vdd.n1804 vdd.n1803 0.152939
R22934 vdd.n1803 vdd.n1802 0.152939
R22935 vdd.n1802 vdd.n1753 0.152939
R22936 vdd.n1798 vdd.n1753 0.152939
R22937 vdd.n1798 vdd.n1797 0.152939
R22938 vdd.n1797 vdd.n1796 0.152939
R22939 vdd.n1796 vdd.n1759 0.152939
R22940 vdd.n1792 vdd.n1759 0.152939
R22941 vdd.n1792 vdd.n1791 0.152939
R22942 vdd.n1791 vdd.n1790 0.152939
R22943 vdd.n1790 vdd.n1765 0.152939
R22944 vdd.n1786 vdd.n1765 0.152939
R22945 vdd.n1786 vdd.n1785 0.152939
R22946 vdd.n1785 vdd.n1784 0.152939
R22947 vdd.n1784 vdd.n1771 0.152939
R22948 vdd.n1780 vdd.n1771 0.152939
R22949 vdd.n1780 vdd.n1779 0.152939
R22950 vdd.n1882 vdd.n1881 0.152939
R22951 vdd.n1882 vdd.n1638 0.152939
R22952 vdd.n1897 vdd.n1638 0.152939
R22953 vdd.n1898 vdd.n1897 0.152939
R22954 vdd.n1899 vdd.n1898 0.152939
R22955 vdd.n1899 vdd.n1627 0.152939
R22956 vdd.n1914 vdd.n1627 0.152939
R22957 vdd.n1915 vdd.n1914 0.152939
R22958 vdd.n1917 vdd.n1915 0.152939
R22959 vdd.n1917 vdd.n1916 0.152939
R22960 vdd.n2088 vdd.n2087 0.110256
R22961 vdd.n3108 vdd.n481 0.110256
R22962 vdd.n2980 vdd.n2979 0.110256
R22963 vdd.n1981 vdd.n1980 0.110256
R22964 vdd.n1931 vdd.n1616 0.0695946
R22965 vdd.n3319 vdd.n298 0.0695946
R22966 vdd.n3319 vdd.n3318 0.0695946
R22967 vdd.n1916 vdd.n1616 0.0695946
R22968 vdd.n2088 vdd.n968 0.0431829
R22969 vdd.n1981 vdd.n1068 0.0431829
R22970 vdd.n3108 vdd.n519 0.0431829
R22971 vdd.n2979 vdd.n572 0.0431829
R22972 vdd vdd.n28 0.00833333
R22973 CSoutput.n19 CSoutput.t185 184.661
R22974 CSoutput.n78 CSoutput.n77 165.8
R22975 CSoutput.n76 CSoutput.n0 165.8
R22976 CSoutput.n75 CSoutput.n74 165.8
R22977 CSoutput.n73 CSoutput.n72 165.8
R22978 CSoutput.n71 CSoutput.n2 165.8
R22979 CSoutput.n69 CSoutput.n68 165.8
R22980 CSoutput.n67 CSoutput.n3 165.8
R22981 CSoutput.n66 CSoutput.n65 165.8
R22982 CSoutput.n63 CSoutput.n4 165.8
R22983 CSoutput.n61 CSoutput.n60 165.8
R22984 CSoutput.n59 CSoutput.n5 165.8
R22985 CSoutput.n58 CSoutput.n57 165.8
R22986 CSoutput.n55 CSoutput.n6 165.8
R22987 CSoutput.n54 CSoutput.n53 165.8
R22988 CSoutput.n52 CSoutput.n51 165.8
R22989 CSoutput.n50 CSoutput.n8 165.8
R22990 CSoutput.n48 CSoutput.n47 165.8
R22991 CSoutput.n46 CSoutput.n9 165.8
R22992 CSoutput.n45 CSoutput.n44 165.8
R22993 CSoutput.n42 CSoutput.n10 165.8
R22994 CSoutput.n41 CSoutput.n40 165.8
R22995 CSoutput.n39 CSoutput.n38 165.8
R22996 CSoutput.n37 CSoutput.n12 165.8
R22997 CSoutput.n35 CSoutput.n34 165.8
R22998 CSoutput.n33 CSoutput.n13 165.8
R22999 CSoutput.n32 CSoutput.n31 165.8
R23000 CSoutput.n29 CSoutput.n14 165.8
R23001 CSoutput.n28 CSoutput.n27 165.8
R23002 CSoutput.n26 CSoutput.n25 165.8
R23003 CSoutput.n24 CSoutput.n16 165.8
R23004 CSoutput.n22 CSoutput.n21 165.8
R23005 CSoutput.n20 CSoutput.n17 165.8
R23006 CSoutput.n77 CSoutput.t188 162.194
R23007 CSoutput.n18 CSoutput.t181 120.501
R23008 CSoutput.n23 CSoutput.t174 120.501
R23009 CSoutput.n15 CSoutput.t169 120.501
R23010 CSoutput.n30 CSoutput.t183 120.501
R23011 CSoutput.n36 CSoutput.t184 120.501
R23012 CSoutput.n11 CSoutput.t171 120.501
R23013 CSoutput.n43 CSoutput.t168 120.501
R23014 CSoutput.n49 CSoutput.t187 120.501
R23015 CSoutput.n7 CSoutput.t175 120.501
R23016 CSoutput.n56 CSoutput.t178 120.501
R23017 CSoutput.n62 CSoutput.t189 120.501
R23018 CSoutput.n64 CSoutput.t179 120.501
R23019 CSoutput.n70 CSoutput.t180 120.501
R23020 CSoutput.n1 CSoutput.t173 120.501
R23021 CSoutput.n270 CSoutput.n268 103.469
R23022 CSoutput.n262 CSoutput.n260 103.469
R23023 CSoutput.n255 CSoutput.n253 103.469
R23024 CSoutput.n96 CSoutput.n94 103.469
R23025 CSoutput.n88 CSoutput.n86 103.469
R23026 CSoutput.n81 CSoutput.n79 103.469
R23027 CSoutput.n272 CSoutput.n271 103.111
R23028 CSoutput.n270 CSoutput.n269 103.111
R23029 CSoutput.n266 CSoutput.n265 103.111
R23030 CSoutput.n264 CSoutput.n263 103.111
R23031 CSoutput.n262 CSoutput.n261 103.111
R23032 CSoutput.n259 CSoutput.n258 103.111
R23033 CSoutput.n257 CSoutput.n256 103.111
R23034 CSoutput.n255 CSoutput.n254 103.111
R23035 CSoutput.n96 CSoutput.n95 103.111
R23036 CSoutput.n98 CSoutput.n97 103.111
R23037 CSoutput.n100 CSoutput.n99 103.111
R23038 CSoutput.n88 CSoutput.n87 103.111
R23039 CSoutput.n90 CSoutput.n89 103.111
R23040 CSoutput.n92 CSoutput.n91 103.111
R23041 CSoutput.n81 CSoutput.n80 103.111
R23042 CSoutput.n83 CSoutput.n82 103.111
R23043 CSoutput.n85 CSoutput.n84 103.111
R23044 CSoutput.n274 CSoutput.n273 103.111
R23045 CSoutput.n318 CSoutput.n316 81.5057
R23046 CSoutput.n298 CSoutput.n296 81.5057
R23047 CSoutput.n279 CSoutput.n277 81.5057
R23048 CSoutput.n378 CSoutput.n376 81.5057
R23049 CSoutput.n358 CSoutput.n356 81.5057
R23050 CSoutput.n339 CSoutput.n337 81.5057
R23051 CSoutput.n334 CSoutput.n333 80.9324
R23052 CSoutput.n332 CSoutput.n331 80.9324
R23053 CSoutput.n330 CSoutput.n329 80.9324
R23054 CSoutput.n328 CSoutput.n327 80.9324
R23055 CSoutput.n326 CSoutput.n325 80.9324
R23056 CSoutput.n324 CSoutput.n323 80.9324
R23057 CSoutput.n322 CSoutput.n321 80.9324
R23058 CSoutput.n320 CSoutput.n319 80.9324
R23059 CSoutput.n318 CSoutput.n317 80.9324
R23060 CSoutput.n314 CSoutput.n313 80.9324
R23061 CSoutput.n312 CSoutput.n311 80.9324
R23062 CSoutput.n310 CSoutput.n309 80.9324
R23063 CSoutput.n308 CSoutput.n307 80.9324
R23064 CSoutput.n306 CSoutput.n305 80.9324
R23065 CSoutput.n304 CSoutput.n303 80.9324
R23066 CSoutput.n302 CSoutput.n301 80.9324
R23067 CSoutput.n300 CSoutput.n299 80.9324
R23068 CSoutput.n298 CSoutput.n297 80.9324
R23069 CSoutput.n295 CSoutput.n294 80.9324
R23070 CSoutput.n293 CSoutput.n292 80.9324
R23071 CSoutput.n291 CSoutput.n290 80.9324
R23072 CSoutput.n289 CSoutput.n288 80.9324
R23073 CSoutput.n287 CSoutput.n286 80.9324
R23074 CSoutput.n285 CSoutput.n284 80.9324
R23075 CSoutput.n283 CSoutput.n282 80.9324
R23076 CSoutput.n281 CSoutput.n280 80.9324
R23077 CSoutput.n279 CSoutput.n278 80.9324
R23078 CSoutput.n378 CSoutput.n377 80.9324
R23079 CSoutput.n380 CSoutput.n379 80.9324
R23080 CSoutput.n382 CSoutput.n381 80.9324
R23081 CSoutput.n384 CSoutput.n383 80.9324
R23082 CSoutput.n386 CSoutput.n385 80.9324
R23083 CSoutput.n388 CSoutput.n387 80.9324
R23084 CSoutput.n390 CSoutput.n389 80.9324
R23085 CSoutput.n392 CSoutput.n391 80.9324
R23086 CSoutput.n394 CSoutput.n393 80.9324
R23087 CSoutput.n358 CSoutput.n357 80.9324
R23088 CSoutput.n360 CSoutput.n359 80.9324
R23089 CSoutput.n362 CSoutput.n361 80.9324
R23090 CSoutput.n364 CSoutput.n363 80.9324
R23091 CSoutput.n366 CSoutput.n365 80.9324
R23092 CSoutput.n368 CSoutput.n367 80.9324
R23093 CSoutput.n370 CSoutput.n369 80.9324
R23094 CSoutput.n372 CSoutput.n371 80.9324
R23095 CSoutput.n374 CSoutput.n373 80.9324
R23096 CSoutput.n339 CSoutput.n338 80.9324
R23097 CSoutput.n341 CSoutput.n340 80.9324
R23098 CSoutput.n343 CSoutput.n342 80.9324
R23099 CSoutput.n345 CSoutput.n344 80.9324
R23100 CSoutput.n347 CSoutput.n346 80.9324
R23101 CSoutput.n349 CSoutput.n348 80.9324
R23102 CSoutput.n351 CSoutput.n350 80.9324
R23103 CSoutput.n353 CSoutput.n352 80.9324
R23104 CSoutput.n355 CSoutput.n354 80.9324
R23105 CSoutput.n25 CSoutput.n24 48.1486
R23106 CSoutput.n69 CSoutput.n3 48.1486
R23107 CSoutput.n38 CSoutput.n37 48.1486
R23108 CSoutput.n42 CSoutput.n41 48.1486
R23109 CSoutput.n51 CSoutput.n50 48.1486
R23110 CSoutput.n55 CSoutput.n54 48.1486
R23111 CSoutput.n22 CSoutput.n17 46.462
R23112 CSoutput.n72 CSoutput.n71 46.462
R23113 CSoutput.n20 CSoutput.n19 44.9055
R23114 CSoutput.n29 CSoutput.n28 43.7635
R23115 CSoutput.n65 CSoutput.n63 43.7635
R23116 CSoutput.n35 CSoutput.n13 41.7396
R23117 CSoutput.n57 CSoutput.n5 41.7396
R23118 CSoutput.n44 CSoutput.n9 37.0171
R23119 CSoutput.n48 CSoutput.n9 37.0171
R23120 CSoutput.n76 CSoutput.n75 34.9932
R23121 CSoutput.n31 CSoutput.n13 32.2947
R23122 CSoutput.n61 CSoutput.n5 32.2947
R23123 CSoutput.n30 CSoutput.n29 29.6014
R23124 CSoutput.n63 CSoutput.n62 29.6014
R23125 CSoutput.n19 CSoutput.n18 28.4085
R23126 CSoutput.n18 CSoutput.n17 25.1176
R23127 CSoutput.n72 CSoutput.n1 25.1176
R23128 CSoutput.n43 CSoutput.n42 22.0922
R23129 CSoutput.n50 CSoutput.n49 22.0922
R23130 CSoutput.n77 CSoutput.n76 21.8586
R23131 CSoutput.n37 CSoutput.n36 18.9681
R23132 CSoutput.n56 CSoutput.n55 18.9681
R23133 CSoutput.n25 CSoutput.n15 17.6292
R23134 CSoutput.n64 CSoutput.n3 17.6292
R23135 CSoutput.n24 CSoutput.n23 15.844
R23136 CSoutput.n70 CSoutput.n69 15.844
R23137 CSoutput.n38 CSoutput.n11 14.5051
R23138 CSoutput.n54 CSoutput.n7 14.5051
R23139 CSoutput.n397 CSoutput.n78 11.4982
R23140 CSoutput.n41 CSoutput.n11 11.3811
R23141 CSoutput.n51 CSoutput.n7 11.3811
R23142 CSoutput.n23 CSoutput.n22 10.0422
R23143 CSoutput.n71 CSoutput.n70 10.0422
R23144 CSoutput.n267 CSoutput.n259 9.25285
R23145 CSoutput.n93 CSoutput.n85 9.25285
R23146 CSoutput.n336 CSoutput.n276 9.09467
R23147 CSoutput.n315 CSoutput.n295 8.98182
R23148 CSoutput.n375 CSoutput.n355 8.98182
R23149 CSoutput.n28 CSoutput.n15 8.25698
R23150 CSoutput.n65 CSoutput.n64 8.25698
R23151 CSoutput.n276 CSoutput.n275 7.12641
R23152 CSoutput.n102 CSoutput.n101 7.12641
R23153 CSoutput.n36 CSoutput.n35 6.91809
R23154 CSoutput.n57 CSoutput.n56 6.91809
R23155 CSoutput.n336 CSoutput.n335 6.02792
R23156 CSoutput.n396 CSoutput.n395 6.02792
R23157 CSoutput.n397 CSoutput.n102 5.50223
R23158 CSoutput.n335 CSoutput.n334 5.25266
R23159 CSoutput.n315 CSoutput.n314 5.25266
R23160 CSoutput.n395 CSoutput.n394 5.25266
R23161 CSoutput.n375 CSoutput.n374 5.25266
R23162 CSoutput.n275 CSoutput.n274 5.1449
R23163 CSoutput.n267 CSoutput.n266 5.1449
R23164 CSoutput.n101 CSoutput.n100 5.1449
R23165 CSoutput.n93 CSoutput.n92 5.1449
R23166 CSoutput.n193 CSoutput.n146 4.5005
R23167 CSoutput.n162 CSoutput.n146 4.5005
R23168 CSoutput.n157 CSoutput.n141 4.5005
R23169 CSoutput.n157 CSoutput.n143 4.5005
R23170 CSoutput.n157 CSoutput.n140 4.5005
R23171 CSoutput.n157 CSoutput.n144 4.5005
R23172 CSoutput.n157 CSoutput.n139 4.5005
R23173 CSoutput.n157 CSoutput.t172 4.5005
R23174 CSoutput.n157 CSoutput.n138 4.5005
R23175 CSoutput.n157 CSoutput.n145 4.5005
R23176 CSoutput.n157 CSoutput.n146 4.5005
R23177 CSoutput.n155 CSoutput.n141 4.5005
R23178 CSoutput.n155 CSoutput.n143 4.5005
R23179 CSoutput.n155 CSoutput.n140 4.5005
R23180 CSoutput.n155 CSoutput.n144 4.5005
R23181 CSoutput.n155 CSoutput.n139 4.5005
R23182 CSoutput.n155 CSoutput.t172 4.5005
R23183 CSoutput.n155 CSoutput.n138 4.5005
R23184 CSoutput.n155 CSoutput.n145 4.5005
R23185 CSoutput.n155 CSoutput.n146 4.5005
R23186 CSoutput.n154 CSoutput.n141 4.5005
R23187 CSoutput.n154 CSoutput.n143 4.5005
R23188 CSoutput.n154 CSoutput.n140 4.5005
R23189 CSoutput.n154 CSoutput.n144 4.5005
R23190 CSoutput.n154 CSoutput.n139 4.5005
R23191 CSoutput.n154 CSoutput.t172 4.5005
R23192 CSoutput.n154 CSoutput.n138 4.5005
R23193 CSoutput.n154 CSoutput.n145 4.5005
R23194 CSoutput.n154 CSoutput.n146 4.5005
R23195 CSoutput.n239 CSoutput.n141 4.5005
R23196 CSoutput.n239 CSoutput.n143 4.5005
R23197 CSoutput.n239 CSoutput.n140 4.5005
R23198 CSoutput.n239 CSoutput.n144 4.5005
R23199 CSoutput.n239 CSoutput.n139 4.5005
R23200 CSoutput.n239 CSoutput.t172 4.5005
R23201 CSoutput.n239 CSoutput.n138 4.5005
R23202 CSoutput.n239 CSoutput.n145 4.5005
R23203 CSoutput.n239 CSoutput.n146 4.5005
R23204 CSoutput.n237 CSoutput.n141 4.5005
R23205 CSoutput.n237 CSoutput.n143 4.5005
R23206 CSoutput.n237 CSoutput.n140 4.5005
R23207 CSoutput.n237 CSoutput.n144 4.5005
R23208 CSoutput.n237 CSoutput.n139 4.5005
R23209 CSoutput.n237 CSoutput.t172 4.5005
R23210 CSoutput.n237 CSoutput.n138 4.5005
R23211 CSoutput.n237 CSoutput.n145 4.5005
R23212 CSoutput.n235 CSoutput.n141 4.5005
R23213 CSoutput.n235 CSoutput.n143 4.5005
R23214 CSoutput.n235 CSoutput.n140 4.5005
R23215 CSoutput.n235 CSoutput.n144 4.5005
R23216 CSoutput.n235 CSoutput.n139 4.5005
R23217 CSoutput.n235 CSoutput.t172 4.5005
R23218 CSoutput.n235 CSoutput.n138 4.5005
R23219 CSoutput.n235 CSoutput.n145 4.5005
R23220 CSoutput.n165 CSoutput.n141 4.5005
R23221 CSoutput.n165 CSoutput.n143 4.5005
R23222 CSoutput.n165 CSoutput.n140 4.5005
R23223 CSoutput.n165 CSoutput.n144 4.5005
R23224 CSoutput.n165 CSoutput.n139 4.5005
R23225 CSoutput.n165 CSoutput.t172 4.5005
R23226 CSoutput.n165 CSoutput.n138 4.5005
R23227 CSoutput.n165 CSoutput.n145 4.5005
R23228 CSoutput.n165 CSoutput.n146 4.5005
R23229 CSoutput.n164 CSoutput.n141 4.5005
R23230 CSoutput.n164 CSoutput.n143 4.5005
R23231 CSoutput.n164 CSoutput.n140 4.5005
R23232 CSoutput.n164 CSoutput.n144 4.5005
R23233 CSoutput.n164 CSoutput.n139 4.5005
R23234 CSoutput.n164 CSoutput.t172 4.5005
R23235 CSoutput.n164 CSoutput.n138 4.5005
R23236 CSoutput.n164 CSoutput.n145 4.5005
R23237 CSoutput.n164 CSoutput.n146 4.5005
R23238 CSoutput.n168 CSoutput.n141 4.5005
R23239 CSoutput.n168 CSoutput.n143 4.5005
R23240 CSoutput.n168 CSoutput.n140 4.5005
R23241 CSoutput.n168 CSoutput.n144 4.5005
R23242 CSoutput.n168 CSoutput.n139 4.5005
R23243 CSoutput.n168 CSoutput.t172 4.5005
R23244 CSoutput.n168 CSoutput.n138 4.5005
R23245 CSoutput.n168 CSoutput.n145 4.5005
R23246 CSoutput.n168 CSoutput.n146 4.5005
R23247 CSoutput.n167 CSoutput.n141 4.5005
R23248 CSoutput.n167 CSoutput.n143 4.5005
R23249 CSoutput.n167 CSoutput.n140 4.5005
R23250 CSoutput.n167 CSoutput.n144 4.5005
R23251 CSoutput.n167 CSoutput.n139 4.5005
R23252 CSoutput.n167 CSoutput.t172 4.5005
R23253 CSoutput.n167 CSoutput.n138 4.5005
R23254 CSoutput.n167 CSoutput.n145 4.5005
R23255 CSoutput.n167 CSoutput.n146 4.5005
R23256 CSoutput.n150 CSoutput.n141 4.5005
R23257 CSoutput.n150 CSoutput.n143 4.5005
R23258 CSoutput.n150 CSoutput.n140 4.5005
R23259 CSoutput.n150 CSoutput.n144 4.5005
R23260 CSoutput.n150 CSoutput.n139 4.5005
R23261 CSoutput.n150 CSoutput.t172 4.5005
R23262 CSoutput.n150 CSoutput.n138 4.5005
R23263 CSoutput.n150 CSoutput.n145 4.5005
R23264 CSoutput.n150 CSoutput.n146 4.5005
R23265 CSoutput.n242 CSoutput.n141 4.5005
R23266 CSoutput.n242 CSoutput.n143 4.5005
R23267 CSoutput.n242 CSoutput.n140 4.5005
R23268 CSoutput.n242 CSoutput.n144 4.5005
R23269 CSoutput.n242 CSoutput.n139 4.5005
R23270 CSoutput.n242 CSoutput.t172 4.5005
R23271 CSoutput.n242 CSoutput.n138 4.5005
R23272 CSoutput.n242 CSoutput.n145 4.5005
R23273 CSoutput.n242 CSoutput.n146 4.5005
R23274 CSoutput.n229 CSoutput.n200 4.5005
R23275 CSoutput.n229 CSoutput.n206 4.5005
R23276 CSoutput.n187 CSoutput.n176 4.5005
R23277 CSoutput.n187 CSoutput.n178 4.5005
R23278 CSoutput.n187 CSoutput.n175 4.5005
R23279 CSoutput.n187 CSoutput.n179 4.5005
R23280 CSoutput.n187 CSoutput.n174 4.5005
R23281 CSoutput.n187 CSoutput.t176 4.5005
R23282 CSoutput.n187 CSoutput.n173 4.5005
R23283 CSoutput.n187 CSoutput.n180 4.5005
R23284 CSoutput.n229 CSoutput.n187 4.5005
R23285 CSoutput.n208 CSoutput.n176 4.5005
R23286 CSoutput.n208 CSoutput.n178 4.5005
R23287 CSoutput.n208 CSoutput.n175 4.5005
R23288 CSoutput.n208 CSoutput.n179 4.5005
R23289 CSoutput.n208 CSoutput.n174 4.5005
R23290 CSoutput.n208 CSoutput.t176 4.5005
R23291 CSoutput.n208 CSoutput.n173 4.5005
R23292 CSoutput.n208 CSoutput.n180 4.5005
R23293 CSoutput.n229 CSoutput.n208 4.5005
R23294 CSoutput.n186 CSoutput.n176 4.5005
R23295 CSoutput.n186 CSoutput.n178 4.5005
R23296 CSoutput.n186 CSoutput.n175 4.5005
R23297 CSoutput.n186 CSoutput.n179 4.5005
R23298 CSoutput.n186 CSoutput.n174 4.5005
R23299 CSoutput.n186 CSoutput.t176 4.5005
R23300 CSoutput.n186 CSoutput.n173 4.5005
R23301 CSoutput.n186 CSoutput.n180 4.5005
R23302 CSoutput.n229 CSoutput.n186 4.5005
R23303 CSoutput.n210 CSoutput.n176 4.5005
R23304 CSoutput.n210 CSoutput.n178 4.5005
R23305 CSoutput.n210 CSoutput.n175 4.5005
R23306 CSoutput.n210 CSoutput.n179 4.5005
R23307 CSoutput.n210 CSoutput.n174 4.5005
R23308 CSoutput.n210 CSoutput.t176 4.5005
R23309 CSoutput.n210 CSoutput.n173 4.5005
R23310 CSoutput.n210 CSoutput.n180 4.5005
R23311 CSoutput.n229 CSoutput.n210 4.5005
R23312 CSoutput.n176 CSoutput.n171 4.5005
R23313 CSoutput.n178 CSoutput.n171 4.5005
R23314 CSoutput.n175 CSoutput.n171 4.5005
R23315 CSoutput.n179 CSoutput.n171 4.5005
R23316 CSoutput.n174 CSoutput.n171 4.5005
R23317 CSoutput.t176 CSoutput.n171 4.5005
R23318 CSoutput.n173 CSoutput.n171 4.5005
R23319 CSoutput.n180 CSoutput.n171 4.5005
R23320 CSoutput.n232 CSoutput.n176 4.5005
R23321 CSoutput.n232 CSoutput.n178 4.5005
R23322 CSoutput.n232 CSoutput.n175 4.5005
R23323 CSoutput.n232 CSoutput.n179 4.5005
R23324 CSoutput.n232 CSoutput.n174 4.5005
R23325 CSoutput.n232 CSoutput.t176 4.5005
R23326 CSoutput.n232 CSoutput.n173 4.5005
R23327 CSoutput.n232 CSoutput.n180 4.5005
R23328 CSoutput.n230 CSoutput.n176 4.5005
R23329 CSoutput.n230 CSoutput.n178 4.5005
R23330 CSoutput.n230 CSoutput.n175 4.5005
R23331 CSoutput.n230 CSoutput.n179 4.5005
R23332 CSoutput.n230 CSoutput.n174 4.5005
R23333 CSoutput.n230 CSoutput.t176 4.5005
R23334 CSoutput.n230 CSoutput.n173 4.5005
R23335 CSoutput.n230 CSoutput.n180 4.5005
R23336 CSoutput.n230 CSoutput.n229 4.5005
R23337 CSoutput.n212 CSoutput.n176 4.5005
R23338 CSoutput.n212 CSoutput.n178 4.5005
R23339 CSoutput.n212 CSoutput.n175 4.5005
R23340 CSoutput.n212 CSoutput.n179 4.5005
R23341 CSoutput.n212 CSoutput.n174 4.5005
R23342 CSoutput.n212 CSoutput.t176 4.5005
R23343 CSoutput.n212 CSoutput.n173 4.5005
R23344 CSoutput.n212 CSoutput.n180 4.5005
R23345 CSoutput.n229 CSoutput.n212 4.5005
R23346 CSoutput.n184 CSoutput.n176 4.5005
R23347 CSoutput.n184 CSoutput.n178 4.5005
R23348 CSoutput.n184 CSoutput.n175 4.5005
R23349 CSoutput.n184 CSoutput.n179 4.5005
R23350 CSoutput.n184 CSoutput.n174 4.5005
R23351 CSoutput.n184 CSoutput.t176 4.5005
R23352 CSoutput.n184 CSoutput.n173 4.5005
R23353 CSoutput.n184 CSoutput.n180 4.5005
R23354 CSoutput.n229 CSoutput.n184 4.5005
R23355 CSoutput.n214 CSoutput.n176 4.5005
R23356 CSoutput.n214 CSoutput.n178 4.5005
R23357 CSoutput.n214 CSoutput.n175 4.5005
R23358 CSoutput.n214 CSoutput.n179 4.5005
R23359 CSoutput.n214 CSoutput.n174 4.5005
R23360 CSoutput.n214 CSoutput.t176 4.5005
R23361 CSoutput.n214 CSoutput.n173 4.5005
R23362 CSoutput.n214 CSoutput.n180 4.5005
R23363 CSoutput.n229 CSoutput.n214 4.5005
R23364 CSoutput.n183 CSoutput.n176 4.5005
R23365 CSoutput.n183 CSoutput.n178 4.5005
R23366 CSoutput.n183 CSoutput.n175 4.5005
R23367 CSoutput.n183 CSoutput.n179 4.5005
R23368 CSoutput.n183 CSoutput.n174 4.5005
R23369 CSoutput.n183 CSoutput.t176 4.5005
R23370 CSoutput.n183 CSoutput.n173 4.5005
R23371 CSoutput.n183 CSoutput.n180 4.5005
R23372 CSoutput.n229 CSoutput.n183 4.5005
R23373 CSoutput.n228 CSoutput.n176 4.5005
R23374 CSoutput.n228 CSoutput.n178 4.5005
R23375 CSoutput.n228 CSoutput.n175 4.5005
R23376 CSoutput.n228 CSoutput.n179 4.5005
R23377 CSoutput.n228 CSoutput.n174 4.5005
R23378 CSoutput.n228 CSoutput.t176 4.5005
R23379 CSoutput.n228 CSoutput.n173 4.5005
R23380 CSoutput.n228 CSoutput.n180 4.5005
R23381 CSoutput.n229 CSoutput.n228 4.5005
R23382 CSoutput.n227 CSoutput.n112 4.5005
R23383 CSoutput.n128 CSoutput.n112 4.5005
R23384 CSoutput.n123 CSoutput.n107 4.5005
R23385 CSoutput.n123 CSoutput.n109 4.5005
R23386 CSoutput.n123 CSoutput.n106 4.5005
R23387 CSoutput.n123 CSoutput.n110 4.5005
R23388 CSoutput.n123 CSoutput.n105 4.5005
R23389 CSoutput.n123 CSoutput.t177 4.5005
R23390 CSoutput.n123 CSoutput.n104 4.5005
R23391 CSoutput.n123 CSoutput.n111 4.5005
R23392 CSoutput.n123 CSoutput.n112 4.5005
R23393 CSoutput.n121 CSoutput.n107 4.5005
R23394 CSoutput.n121 CSoutput.n109 4.5005
R23395 CSoutput.n121 CSoutput.n106 4.5005
R23396 CSoutput.n121 CSoutput.n110 4.5005
R23397 CSoutput.n121 CSoutput.n105 4.5005
R23398 CSoutput.n121 CSoutput.t177 4.5005
R23399 CSoutput.n121 CSoutput.n104 4.5005
R23400 CSoutput.n121 CSoutput.n111 4.5005
R23401 CSoutput.n121 CSoutput.n112 4.5005
R23402 CSoutput.n120 CSoutput.n107 4.5005
R23403 CSoutput.n120 CSoutput.n109 4.5005
R23404 CSoutput.n120 CSoutput.n106 4.5005
R23405 CSoutput.n120 CSoutput.n110 4.5005
R23406 CSoutput.n120 CSoutput.n105 4.5005
R23407 CSoutput.n120 CSoutput.t177 4.5005
R23408 CSoutput.n120 CSoutput.n104 4.5005
R23409 CSoutput.n120 CSoutput.n111 4.5005
R23410 CSoutput.n120 CSoutput.n112 4.5005
R23411 CSoutput.n249 CSoutput.n107 4.5005
R23412 CSoutput.n249 CSoutput.n109 4.5005
R23413 CSoutput.n249 CSoutput.n106 4.5005
R23414 CSoutput.n249 CSoutput.n110 4.5005
R23415 CSoutput.n249 CSoutput.n105 4.5005
R23416 CSoutput.n249 CSoutput.t177 4.5005
R23417 CSoutput.n249 CSoutput.n104 4.5005
R23418 CSoutput.n249 CSoutput.n111 4.5005
R23419 CSoutput.n249 CSoutput.n112 4.5005
R23420 CSoutput.n247 CSoutput.n107 4.5005
R23421 CSoutput.n247 CSoutput.n109 4.5005
R23422 CSoutput.n247 CSoutput.n106 4.5005
R23423 CSoutput.n247 CSoutput.n110 4.5005
R23424 CSoutput.n247 CSoutput.n105 4.5005
R23425 CSoutput.n247 CSoutput.t177 4.5005
R23426 CSoutput.n247 CSoutput.n104 4.5005
R23427 CSoutput.n247 CSoutput.n111 4.5005
R23428 CSoutput.n245 CSoutput.n107 4.5005
R23429 CSoutput.n245 CSoutput.n109 4.5005
R23430 CSoutput.n245 CSoutput.n106 4.5005
R23431 CSoutput.n245 CSoutput.n110 4.5005
R23432 CSoutput.n245 CSoutput.n105 4.5005
R23433 CSoutput.n245 CSoutput.t177 4.5005
R23434 CSoutput.n245 CSoutput.n104 4.5005
R23435 CSoutput.n245 CSoutput.n111 4.5005
R23436 CSoutput.n131 CSoutput.n107 4.5005
R23437 CSoutput.n131 CSoutput.n109 4.5005
R23438 CSoutput.n131 CSoutput.n106 4.5005
R23439 CSoutput.n131 CSoutput.n110 4.5005
R23440 CSoutput.n131 CSoutput.n105 4.5005
R23441 CSoutput.n131 CSoutput.t177 4.5005
R23442 CSoutput.n131 CSoutput.n104 4.5005
R23443 CSoutput.n131 CSoutput.n111 4.5005
R23444 CSoutput.n131 CSoutput.n112 4.5005
R23445 CSoutput.n130 CSoutput.n107 4.5005
R23446 CSoutput.n130 CSoutput.n109 4.5005
R23447 CSoutput.n130 CSoutput.n106 4.5005
R23448 CSoutput.n130 CSoutput.n110 4.5005
R23449 CSoutput.n130 CSoutput.n105 4.5005
R23450 CSoutput.n130 CSoutput.t177 4.5005
R23451 CSoutput.n130 CSoutput.n104 4.5005
R23452 CSoutput.n130 CSoutput.n111 4.5005
R23453 CSoutput.n130 CSoutput.n112 4.5005
R23454 CSoutput.n134 CSoutput.n107 4.5005
R23455 CSoutput.n134 CSoutput.n109 4.5005
R23456 CSoutput.n134 CSoutput.n106 4.5005
R23457 CSoutput.n134 CSoutput.n110 4.5005
R23458 CSoutput.n134 CSoutput.n105 4.5005
R23459 CSoutput.n134 CSoutput.t177 4.5005
R23460 CSoutput.n134 CSoutput.n104 4.5005
R23461 CSoutput.n134 CSoutput.n111 4.5005
R23462 CSoutput.n134 CSoutput.n112 4.5005
R23463 CSoutput.n133 CSoutput.n107 4.5005
R23464 CSoutput.n133 CSoutput.n109 4.5005
R23465 CSoutput.n133 CSoutput.n106 4.5005
R23466 CSoutput.n133 CSoutput.n110 4.5005
R23467 CSoutput.n133 CSoutput.n105 4.5005
R23468 CSoutput.n133 CSoutput.t177 4.5005
R23469 CSoutput.n133 CSoutput.n104 4.5005
R23470 CSoutput.n133 CSoutput.n111 4.5005
R23471 CSoutput.n133 CSoutput.n112 4.5005
R23472 CSoutput.n116 CSoutput.n107 4.5005
R23473 CSoutput.n116 CSoutput.n109 4.5005
R23474 CSoutput.n116 CSoutput.n106 4.5005
R23475 CSoutput.n116 CSoutput.n110 4.5005
R23476 CSoutput.n116 CSoutput.n105 4.5005
R23477 CSoutput.n116 CSoutput.t177 4.5005
R23478 CSoutput.n116 CSoutput.n104 4.5005
R23479 CSoutput.n116 CSoutput.n111 4.5005
R23480 CSoutput.n116 CSoutput.n112 4.5005
R23481 CSoutput.n252 CSoutput.n107 4.5005
R23482 CSoutput.n252 CSoutput.n109 4.5005
R23483 CSoutput.n252 CSoutput.n106 4.5005
R23484 CSoutput.n252 CSoutput.n110 4.5005
R23485 CSoutput.n252 CSoutput.n105 4.5005
R23486 CSoutput.n252 CSoutput.t177 4.5005
R23487 CSoutput.n252 CSoutput.n104 4.5005
R23488 CSoutput.n252 CSoutput.n111 4.5005
R23489 CSoutput.n252 CSoutput.n112 4.5005
R23490 CSoutput.n275 CSoutput.n267 4.10845
R23491 CSoutput.n101 CSoutput.n93 4.10845
R23492 CSoutput.n273 CSoutput.t148 4.06363
R23493 CSoutput.n273 CSoutput.t157 4.06363
R23494 CSoutput.n271 CSoutput.t164 4.06363
R23495 CSoutput.n271 CSoutput.t131 4.06363
R23496 CSoutput.n269 CSoutput.t135 4.06363
R23497 CSoutput.n269 CSoutput.t158 4.06363
R23498 CSoutput.n268 CSoutput.t165 4.06363
R23499 CSoutput.n268 CSoutput.t166 4.06363
R23500 CSoutput.n265 CSoutput.t141 4.06363
R23501 CSoutput.n265 CSoutput.t154 4.06363
R23502 CSoutput.n263 CSoutput.t159 4.06363
R23503 CSoutput.n263 CSoutput.t123 4.06363
R23504 CSoutput.n261 CSoutput.t124 4.06363
R23505 CSoutput.n261 CSoutput.t155 4.06363
R23506 CSoutput.n260 CSoutput.t162 4.06363
R23507 CSoutput.n260 CSoutput.t163 4.06363
R23508 CSoutput.n258 CSoutput.t156 4.06363
R23509 CSoutput.n258 CSoutput.t139 4.06363
R23510 CSoutput.n256 CSoutput.t152 4.06363
R23511 CSoutput.n256 CSoutput.t130 4.06363
R23512 CSoutput.n254 CSoutput.t160 4.06363
R23513 CSoutput.n254 CSoutput.t125 4.06363
R23514 CSoutput.n253 CSoutput.t142 4.06363
R23515 CSoutput.n253 CSoutput.t136 4.06363
R23516 CSoutput.n94 CSoutput.t150 4.06363
R23517 CSoutput.n94 CSoutput.t138 4.06363
R23518 CSoutput.n95 CSoutput.t129 4.06363
R23519 CSoutput.n95 CSoutput.t151 4.06363
R23520 CSoutput.n97 CSoutput.t149 4.06363
R23521 CSoutput.n97 CSoutput.t137 4.06363
R23522 CSoutput.n99 CSoutput.t128 4.06363
R23523 CSoutput.n99 CSoutput.t127 4.06363
R23524 CSoutput.n86 CSoutput.t145 4.06363
R23525 CSoutput.n86 CSoutput.t134 4.06363
R23526 CSoutput.n87 CSoutput.t122 4.06363
R23527 CSoutput.n87 CSoutput.t146 4.06363
R23528 CSoutput.n89 CSoutput.t144 4.06363
R23529 CSoutput.n89 CSoutput.t132 4.06363
R23530 CSoutput.n91 CSoutput.t121 4.06363
R23531 CSoutput.n91 CSoutput.t120 4.06363
R23532 CSoutput.n79 CSoutput.t167 4.06363
R23533 CSoutput.n79 CSoutput.t143 4.06363
R23534 CSoutput.n80 CSoutput.t126 4.06363
R23535 CSoutput.n80 CSoutput.t161 4.06363
R23536 CSoutput.n82 CSoutput.t133 4.06363
R23537 CSoutput.n82 CSoutput.t153 4.06363
R23538 CSoutput.n84 CSoutput.t140 4.06363
R23539 CSoutput.n84 CSoutput.t147 4.06363
R23540 CSoutput.n44 CSoutput.n43 3.79402
R23541 CSoutput.n49 CSoutput.n48 3.79402
R23542 CSoutput.n335 CSoutput.n315 3.72967
R23543 CSoutput.n395 CSoutput.n375 3.72967
R23544 CSoutput.n396 CSoutput.n336 3.71319
R23545 CSoutput.n397 CSoutput.n396 3.57343
R23546 CSoutput.n333 CSoutput.t48 2.82907
R23547 CSoutput.n333 CSoutput.t15 2.82907
R23548 CSoutput.n331 CSoutput.t118 2.82907
R23549 CSoutput.n331 CSoutput.t100 2.82907
R23550 CSoutput.n329 CSoutput.t22 2.82907
R23551 CSoutput.n329 CSoutput.t29 2.82907
R23552 CSoutput.n327 CSoutput.t13 2.82907
R23553 CSoutput.n327 CSoutput.t107 2.82907
R23554 CSoutput.n325 CSoutput.t69 2.82907
R23555 CSoutput.n325 CSoutput.t1 2.82907
R23556 CSoutput.n323 CSoutput.t111 2.82907
R23557 CSoutput.n323 CSoutput.t91 2.82907
R23558 CSoutput.n321 CSoutput.t49 2.82907
R23559 CSoutput.n321 CSoutput.t58 2.82907
R23560 CSoutput.n319 CSoutput.t0 2.82907
R23561 CSoutput.n319 CSoutput.t101 2.82907
R23562 CSoutput.n317 CSoutput.t92 2.82907
R23563 CSoutput.n317 CSoutput.t31 2.82907
R23564 CSoutput.n316 CSoutput.t16 2.82907
R23565 CSoutput.n316 CSoutput.t110 2.82907
R23566 CSoutput.n313 CSoutput.t119 2.82907
R23567 CSoutput.n313 CSoutput.t105 2.82907
R23568 CSoutput.n311 CSoutput.t104 2.82907
R23569 CSoutput.n311 CSoutput.t109 2.82907
R23570 CSoutput.n309 CSoutput.t30 2.82907
R23571 CSoutput.n309 CSoutput.t117 2.82907
R23572 CSoutput.n307 CSoutput.t9 2.82907
R23573 CSoutput.n307 CSoutput.t108 2.82907
R23574 CSoutput.n305 CSoutput.t24 2.82907
R23575 CSoutput.n305 CSoutput.t42 2.82907
R23576 CSoutput.n303 CSoutput.t40 2.82907
R23577 CSoutput.n303 CSoutput.t14 2.82907
R23578 CSoutput.n301 CSoutput.t55 2.82907
R23579 CSoutput.n301 CSoutput.t25 2.82907
R23580 CSoutput.n299 CSoutput.t26 2.82907
R23581 CSoutput.n299 CSoutput.t41 2.82907
R23582 CSoutput.n297 CSoutput.t39 2.82907
R23583 CSoutput.n297 CSoutput.t53 2.82907
R23584 CSoutput.n296 CSoutput.t54 2.82907
R23585 CSoutput.n296 CSoutput.t27 2.82907
R23586 CSoutput.n294 CSoutput.t68 2.82907
R23587 CSoutput.n294 CSoutput.t99 2.82907
R23588 CSoutput.n292 CSoutput.t76 2.82907
R23589 CSoutput.n292 CSoutput.t115 2.82907
R23590 CSoutput.n290 CSoutput.t17 2.82907
R23591 CSoutput.n290 CSoutput.t33 2.82907
R23592 CSoutput.n288 CSoutput.t59 2.82907
R23593 CSoutput.n288 CSoutput.t90 2.82907
R23594 CSoutput.n286 CSoutput.t80 2.82907
R23595 CSoutput.n286 CSoutput.t44 2.82907
R23596 CSoutput.n284 CSoutput.t6 2.82907
R23597 CSoutput.n284 CSoutput.t63 2.82907
R23598 CSoutput.n282 CSoutput.t43 2.82907
R23599 CSoutput.n282 CSoutput.t56 2.82907
R23600 CSoutput.n280 CSoutput.t57 2.82907
R23601 CSoutput.n280 CSoutput.t98 2.82907
R23602 CSoutput.n278 CSoutput.t75 2.82907
R23603 CSoutput.n278 CSoutput.t2 2.82907
R23604 CSoutput.n277 CSoutput.t95 2.82907
R23605 CSoutput.n277 CSoutput.t18 2.82907
R23606 CSoutput.n376 CSoutput.t86 2.82907
R23607 CSoutput.n376 CSoutput.t106 2.82907
R23608 CSoutput.n377 CSoutput.t114 2.82907
R23609 CSoutput.n377 CSoutput.t74 2.82907
R23610 CSoutput.n379 CSoutput.t79 2.82907
R23611 CSoutput.n379 CSoutput.t96 2.82907
R23612 CSoutput.n381 CSoutput.t20 2.82907
R23613 CSoutput.n381 CSoutput.t66 2.82907
R23614 CSoutput.n383 CSoutput.t73 2.82907
R23615 CSoutput.n383 CSoutput.t87 2.82907
R23616 CSoutput.n385 CSoutput.t97 2.82907
R23617 CSoutput.n385 CSoutput.t78 2.82907
R23618 CSoutput.n387 CSoutput.t83 2.82907
R23619 CSoutput.n387 CSoutput.t103 2.82907
R23620 CSoutput.n389 CSoutput.t21 2.82907
R23621 CSoutput.n389 CSoutput.t32 2.82907
R23622 CSoutput.n391 CSoutput.t93 2.82907
R23623 CSoutput.n391 CSoutput.t112 2.82907
R23624 CSoutput.n393 CSoutput.t3 2.82907
R23625 CSoutput.n393 CSoutput.t34 2.82907
R23626 CSoutput.n356 CSoutput.t51 2.82907
R23627 CSoutput.n356 CSoutput.t70 2.82907
R23628 CSoutput.n357 CSoutput.t71 2.82907
R23629 CSoutput.n357 CSoutput.t60 2.82907
R23630 CSoutput.n359 CSoutput.t61 2.82907
R23631 CSoutput.n359 CSoutput.t52 2.82907
R23632 CSoutput.n361 CSoutput.t45 2.82907
R23633 CSoutput.n361 CSoutput.t37 2.82907
R23634 CSoutput.n363 CSoutput.t38 2.82907
R23635 CSoutput.n363 CSoutput.t62 2.82907
R23636 CSoutput.n365 CSoutput.t64 2.82907
R23637 CSoutput.n365 CSoutput.t4 2.82907
R23638 CSoutput.n367 CSoutput.t5 2.82907
R23639 CSoutput.n367 CSoutput.t28 2.82907
R23640 CSoutput.n369 CSoutput.t35 2.82907
R23641 CSoutput.n369 CSoutput.t23 2.82907
R23642 CSoutput.n371 CSoutput.t19 2.82907
R23643 CSoutput.n371 CSoutput.t10 2.82907
R23644 CSoutput.n373 CSoutput.t11 2.82907
R23645 CSoutput.n373 CSoutput.t36 2.82907
R23646 CSoutput.n337 CSoutput.t65 2.82907
R23647 CSoutput.n337 CSoutput.t8 2.82907
R23648 CSoutput.n338 CSoutput.t47 2.82907
R23649 CSoutput.n338 CSoutput.t102 2.82907
R23650 CSoutput.n340 CSoutput.t12 2.82907
R23651 CSoutput.n340 CSoutput.t82 2.82907
R23652 CSoutput.n342 CSoutput.t81 2.82907
R23653 CSoutput.n342 CSoutput.t67 2.82907
R23654 CSoutput.n344 CSoutput.t85 2.82907
R23655 CSoutput.n344 CSoutput.t50 2.82907
R23656 CSoutput.n346 CSoutput.t77 2.82907
R23657 CSoutput.n346 CSoutput.t94 2.82907
R23658 CSoutput.n348 CSoutput.t116 2.82907
R23659 CSoutput.n348 CSoutput.t84 2.82907
R23660 CSoutput.n350 CSoutput.t89 2.82907
R23661 CSoutput.n350 CSoutput.t88 2.82907
R23662 CSoutput.n352 CSoutput.t72 2.82907
R23663 CSoutput.n352 CSoutput.t7 2.82907
R23664 CSoutput.n354 CSoutput.t46 2.82907
R23665 CSoutput.n354 CSoutput.t113 2.82907
R23666 CSoutput.n276 CSoutput.n102 2.57547
R23667 CSoutput.n75 CSoutput.n1 2.45513
R23668 CSoutput.n193 CSoutput.n191 2.251
R23669 CSoutput.n193 CSoutput.n190 2.251
R23670 CSoutput.n193 CSoutput.n189 2.251
R23671 CSoutput.n193 CSoutput.n188 2.251
R23672 CSoutput.n162 CSoutput.n161 2.251
R23673 CSoutput.n162 CSoutput.n160 2.251
R23674 CSoutput.n162 CSoutput.n159 2.251
R23675 CSoutput.n162 CSoutput.n158 2.251
R23676 CSoutput.n235 CSoutput.n234 2.251
R23677 CSoutput.n200 CSoutput.n198 2.251
R23678 CSoutput.n200 CSoutput.n197 2.251
R23679 CSoutput.n200 CSoutput.n196 2.251
R23680 CSoutput.n218 CSoutput.n200 2.251
R23681 CSoutput.n206 CSoutput.n205 2.251
R23682 CSoutput.n206 CSoutput.n204 2.251
R23683 CSoutput.n206 CSoutput.n203 2.251
R23684 CSoutput.n206 CSoutput.n202 2.251
R23685 CSoutput.n232 CSoutput.n172 2.251
R23686 CSoutput.n227 CSoutput.n225 2.251
R23687 CSoutput.n227 CSoutput.n224 2.251
R23688 CSoutput.n227 CSoutput.n223 2.251
R23689 CSoutput.n227 CSoutput.n222 2.251
R23690 CSoutput.n128 CSoutput.n127 2.251
R23691 CSoutput.n128 CSoutput.n126 2.251
R23692 CSoutput.n128 CSoutput.n125 2.251
R23693 CSoutput.n128 CSoutput.n124 2.251
R23694 CSoutput.n245 CSoutput.n244 2.251
R23695 CSoutput.n162 CSoutput.n142 2.2505
R23696 CSoutput.n157 CSoutput.n142 2.2505
R23697 CSoutput.n155 CSoutput.n142 2.2505
R23698 CSoutput.n154 CSoutput.n142 2.2505
R23699 CSoutput.n239 CSoutput.n142 2.2505
R23700 CSoutput.n237 CSoutput.n142 2.2505
R23701 CSoutput.n235 CSoutput.n142 2.2505
R23702 CSoutput.n165 CSoutput.n142 2.2505
R23703 CSoutput.n164 CSoutput.n142 2.2505
R23704 CSoutput.n168 CSoutput.n142 2.2505
R23705 CSoutput.n167 CSoutput.n142 2.2505
R23706 CSoutput.n150 CSoutput.n142 2.2505
R23707 CSoutput.n242 CSoutput.n142 2.2505
R23708 CSoutput.n242 CSoutput.n241 2.2505
R23709 CSoutput.n206 CSoutput.n177 2.2505
R23710 CSoutput.n187 CSoutput.n177 2.2505
R23711 CSoutput.n208 CSoutput.n177 2.2505
R23712 CSoutput.n186 CSoutput.n177 2.2505
R23713 CSoutput.n210 CSoutput.n177 2.2505
R23714 CSoutput.n177 CSoutput.n171 2.2505
R23715 CSoutput.n232 CSoutput.n177 2.2505
R23716 CSoutput.n230 CSoutput.n177 2.2505
R23717 CSoutput.n212 CSoutput.n177 2.2505
R23718 CSoutput.n184 CSoutput.n177 2.2505
R23719 CSoutput.n214 CSoutput.n177 2.2505
R23720 CSoutput.n183 CSoutput.n177 2.2505
R23721 CSoutput.n228 CSoutput.n177 2.2505
R23722 CSoutput.n228 CSoutput.n181 2.2505
R23723 CSoutput.n128 CSoutput.n108 2.2505
R23724 CSoutput.n123 CSoutput.n108 2.2505
R23725 CSoutput.n121 CSoutput.n108 2.2505
R23726 CSoutput.n120 CSoutput.n108 2.2505
R23727 CSoutput.n249 CSoutput.n108 2.2505
R23728 CSoutput.n247 CSoutput.n108 2.2505
R23729 CSoutput.n245 CSoutput.n108 2.2505
R23730 CSoutput.n131 CSoutput.n108 2.2505
R23731 CSoutput.n130 CSoutput.n108 2.2505
R23732 CSoutput.n134 CSoutput.n108 2.2505
R23733 CSoutput.n133 CSoutput.n108 2.2505
R23734 CSoutput.n116 CSoutput.n108 2.2505
R23735 CSoutput.n252 CSoutput.n108 2.2505
R23736 CSoutput.n252 CSoutput.n251 2.2505
R23737 CSoutput.n170 CSoutput.n163 2.25024
R23738 CSoutput.n170 CSoutput.n156 2.25024
R23739 CSoutput.n238 CSoutput.n170 2.25024
R23740 CSoutput.n170 CSoutput.n166 2.25024
R23741 CSoutput.n170 CSoutput.n169 2.25024
R23742 CSoutput.n170 CSoutput.n137 2.25024
R23743 CSoutput.n220 CSoutput.n217 2.25024
R23744 CSoutput.n220 CSoutput.n216 2.25024
R23745 CSoutput.n220 CSoutput.n215 2.25024
R23746 CSoutput.n220 CSoutput.n182 2.25024
R23747 CSoutput.n220 CSoutput.n219 2.25024
R23748 CSoutput.n221 CSoutput.n220 2.25024
R23749 CSoutput.n136 CSoutput.n129 2.25024
R23750 CSoutput.n136 CSoutput.n122 2.25024
R23751 CSoutput.n248 CSoutput.n136 2.25024
R23752 CSoutput.n136 CSoutput.n132 2.25024
R23753 CSoutput.n136 CSoutput.n135 2.25024
R23754 CSoutput.n136 CSoutput.n103 2.25024
R23755 CSoutput.n237 CSoutput.n147 1.50111
R23756 CSoutput.n185 CSoutput.n171 1.50111
R23757 CSoutput.n247 CSoutput.n113 1.50111
R23758 CSoutput.n193 CSoutput.n192 1.501
R23759 CSoutput.n200 CSoutput.n199 1.501
R23760 CSoutput.n227 CSoutput.n226 1.501
R23761 CSoutput.n241 CSoutput.n152 1.12536
R23762 CSoutput.n241 CSoutput.n153 1.12536
R23763 CSoutput.n241 CSoutput.n240 1.12536
R23764 CSoutput.n201 CSoutput.n181 1.12536
R23765 CSoutput.n207 CSoutput.n181 1.12536
R23766 CSoutput.n209 CSoutput.n181 1.12536
R23767 CSoutput.n251 CSoutput.n118 1.12536
R23768 CSoutput.n251 CSoutput.n119 1.12536
R23769 CSoutput.n251 CSoutput.n250 1.12536
R23770 CSoutput.n241 CSoutput.n148 1.12536
R23771 CSoutput.n241 CSoutput.n149 1.12536
R23772 CSoutput.n241 CSoutput.n151 1.12536
R23773 CSoutput.n231 CSoutput.n181 1.12536
R23774 CSoutput.n211 CSoutput.n181 1.12536
R23775 CSoutput.n213 CSoutput.n181 1.12536
R23776 CSoutput.n251 CSoutput.n114 1.12536
R23777 CSoutput.n251 CSoutput.n115 1.12536
R23778 CSoutput.n251 CSoutput.n117 1.12536
R23779 CSoutput.n31 CSoutput.n30 0.669944
R23780 CSoutput.n62 CSoutput.n61 0.669944
R23781 CSoutput.n320 CSoutput.n318 0.573776
R23782 CSoutput.n322 CSoutput.n320 0.573776
R23783 CSoutput.n324 CSoutput.n322 0.573776
R23784 CSoutput.n326 CSoutput.n324 0.573776
R23785 CSoutput.n328 CSoutput.n326 0.573776
R23786 CSoutput.n330 CSoutput.n328 0.573776
R23787 CSoutput.n332 CSoutput.n330 0.573776
R23788 CSoutput.n334 CSoutput.n332 0.573776
R23789 CSoutput.n300 CSoutput.n298 0.573776
R23790 CSoutput.n302 CSoutput.n300 0.573776
R23791 CSoutput.n304 CSoutput.n302 0.573776
R23792 CSoutput.n306 CSoutput.n304 0.573776
R23793 CSoutput.n308 CSoutput.n306 0.573776
R23794 CSoutput.n310 CSoutput.n308 0.573776
R23795 CSoutput.n312 CSoutput.n310 0.573776
R23796 CSoutput.n314 CSoutput.n312 0.573776
R23797 CSoutput.n281 CSoutput.n279 0.573776
R23798 CSoutput.n283 CSoutput.n281 0.573776
R23799 CSoutput.n285 CSoutput.n283 0.573776
R23800 CSoutput.n287 CSoutput.n285 0.573776
R23801 CSoutput.n289 CSoutput.n287 0.573776
R23802 CSoutput.n291 CSoutput.n289 0.573776
R23803 CSoutput.n293 CSoutput.n291 0.573776
R23804 CSoutput.n295 CSoutput.n293 0.573776
R23805 CSoutput.n394 CSoutput.n392 0.573776
R23806 CSoutput.n392 CSoutput.n390 0.573776
R23807 CSoutput.n390 CSoutput.n388 0.573776
R23808 CSoutput.n388 CSoutput.n386 0.573776
R23809 CSoutput.n386 CSoutput.n384 0.573776
R23810 CSoutput.n384 CSoutput.n382 0.573776
R23811 CSoutput.n382 CSoutput.n380 0.573776
R23812 CSoutput.n380 CSoutput.n378 0.573776
R23813 CSoutput.n374 CSoutput.n372 0.573776
R23814 CSoutput.n372 CSoutput.n370 0.573776
R23815 CSoutput.n370 CSoutput.n368 0.573776
R23816 CSoutput.n368 CSoutput.n366 0.573776
R23817 CSoutput.n366 CSoutput.n364 0.573776
R23818 CSoutput.n364 CSoutput.n362 0.573776
R23819 CSoutput.n362 CSoutput.n360 0.573776
R23820 CSoutput.n360 CSoutput.n358 0.573776
R23821 CSoutput.n355 CSoutput.n353 0.573776
R23822 CSoutput.n353 CSoutput.n351 0.573776
R23823 CSoutput.n351 CSoutput.n349 0.573776
R23824 CSoutput.n349 CSoutput.n347 0.573776
R23825 CSoutput.n347 CSoutput.n345 0.573776
R23826 CSoutput.n345 CSoutput.n343 0.573776
R23827 CSoutput.n343 CSoutput.n341 0.573776
R23828 CSoutput.n341 CSoutput.n339 0.573776
R23829 CSoutput.n397 CSoutput.n252 0.53442
R23830 CSoutput.n272 CSoutput.n270 0.358259
R23831 CSoutput.n274 CSoutput.n272 0.358259
R23832 CSoutput.n264 CSoutput.n262 0.358259
R23833 CSoutput.n266 CSoutput.n264 0.358259
R23834 CSoutput.n257 CSoutput.n255 0.358259
R23835 CSoutput.n259 CSoutput.n257 0.358259
R23836 CSoutput.n100 CSoutput.n98 0.358259
R23837 CSoutput.n98 CSoutput.n96 0.358259
R23838 CSoutput.n92 CSoutput.n90 0.358259
R23839 CSoutput.n90 CSoutput.n88 0.358259
R23840 CSoutput.n85 CSoutput.n83 0.358259
R23841 CSoutput.n83 CSoutput.n81 0.358259
R23842 CSoutput.n21 CSoutput.n20 0.169105
R23843 CSoutput.n21 CSoutput.n16 0.169105
R23844 CSoutput.n26 CSoutput.n16 0.169105
R23845 CSoutput.n27 CSoutput.n26 0.169105
R23846 CSoutput.n27 CSoutput.n14 0.169105
R23847 CSoutput.n32 CSoutput.n14 0.169105
R23848 CSoutput.n33 CSoutput.n32 0.169105
R23849 CSoutput.n34 CSoutput.n33 0.169105
R23850 CSoutput.n34 CSoutput.n12 0.169105
R23851 CSoutput.n39 CSoutput.n12 0.169105
R23852 CSoutput.n40 CSoutput.n39 0.169105
R23853 CSoutput.n40 CSoutput.n10 0.169105
R23854 CSoutput.n45 CSoutput.n10 0.169105
R23855 CSoutput.n46 CSoutput.n45 0.169105
R23856 CSoutput.n47 CSoutput.n46 0.169105
R23857 CSoutput.n47 CSoutput.n8 0.169105
R23858 CSoutput.n52 CSoutput.n8 0.169105
R23859 CSoutput.n53 CSoutput.n52 0.169105
R23860 CSoutput.n53 CSoutput.n6 0.169105
R23861 CSoutput.n58 CSoutput.n6 0.169105
R23862 CSoutput.n59 CSoutput.n58 0.169105
R23863 CSoutput.n60 CSoutput.n59 0.169105
R23864 CSoutput.n60 CSoutput.n4 0.169105
R23865 CSoutput.n66 CSoutput.n4 0.169105
R23866 CSoutput.n67 CSoutput.n66 0.169105
R23867 CSoutput.n68 CSoutput.n67 0.169105
R23868 CSoutput.n68 CSoutput.n2 0.169105
R23869 CSoutput.n73 CSoutput.n2 0.169105
R23870 CSoutput.n74 CSoutput.n73 0.169105
R23871 CSoutput.n74 CSoutput.n0 0.169105
R23872 CSoutput.n78 CSoutput.n0 0.169105
R23873 CSoutput.n195 CSoutput.n194 0.0910737
R23874 CSoutput.n246 CSoutput.n243 0.0723685
R23875 CSoutput.n200 CSoutput.n195 0.0522944
R23876 CSoutput.n243 CSoutput.n242 0.0499135
R23877 CSoutput.n194 CSoutput.n193 0.0499135
R23878 CSoutput.n228 CSoutput.n227 0.0464294
R23879 CSoutput.n236 CSoutput.n233 0.0391444
R23880 CSoutput.n195 CSoutput.t186 0.023435
R23881 CSoutput.n243 CSoutput.t170 0.02262
R23882 CSoutput.n194 CSoutput.t182 0.02262
R23883 CSoutput CSoutput.n397 0.0052
R23884 CSoutput.n165 CSoutput.n148 0.00365111
R23885 CSoutput.n168 CSoutput.n149 0.00365111
R23886 CSoutput.n151 CSoutput.n150 0.00365111
R23887 CSoutput.n193 CSoutput.n152 0.00365111
R23888 CSoutput.n157 CSoutput.n153 0.00365111
R23889 CSoutput.n240 CSoutput.n154 0.00365111
R23890 CSoutput.n231 CSoutput.n230 0.00365111
R23891 CSoutput.n211 CSoutput.n184 0.00365111
R23892 CSoutput.n213 CSoutput.n183 0.00365111
R23893 CSoutput.n201 CSoutput.n200 0.00365111
R23894 CSoutput.n207 CSoutput.n187 0.00365111
R23895 CSoutput.n209 CSoutput.n186 0.00365111
R23896 CSoutput.n131 CSoutput.n114 0.00365111
R23897 CSoutput.n134 CSoutput.n115 0.00365111
R23898 CSoutput.n117 CSoutput.n116 0.00365111
R23899 CSoutput.n227 CSoutput.n118 0.00365111
R23900 CSoutput.n123 CSoutput.n119 0.00365111
R23901 CSoutput.n250 CSoutput.n120 0.00365111
R23902 CSoutput.n162 CSoutput.n152 0.00340054
R23903 CSoutput.n155 CSoutput.n153 0.00340054
R23904 CSoutput.n240 CSoutput.n239 0.00340054
R23905 CSoutput.n235 CSoutput.n148 0.00340054
R23906 CSoutput.n164 CSoutput.n149 0.00340054
R23907 CSoutput.n167 CSoutput.n151 0.00340054
R23908 CSoutput.n206 CSoutput.n201 0.00340054
R23909 CSoutput.n208 CSoutput.n207 0.00340054
R23910 CSoutput.n210 CSoutput.n209 0.00340054
R23911 CSoutput.n232 CSoutput.n231 0.00340054
R23912 CSoutput.n212 CSoutput.n211 0.00340054
R23913 CSoutput.n214 CSoutput.n213 0.00340054
R23914 CSoutput.n128 CSoutput.n118 0.00340054
R23915 CSoutput.n121 CSoutput.n119 0.00340054
R23916 CSoutput.n250 CSoutput.n249 0.00340054
R23917 CSoutput.n245 CSoutput.n114 0.00340054
R23918 CSoutput.n130 CSoutput.n115 0.00340054
R23919 CSoutput.n133 CSoutput.n117 0.00340054
R23920 CSoutput.n163 CSoutput.n157 0.00252698
R23921 CSoutput.n156 CSoutput.n154 0.00252698
R23922 CSoutput.n238 CSoutput.n237 0.00252698
R23923 CSoutput.n166 CSoutput.n164 0.00252698
R23924 CSoutput.n169 CSoutput.n167 0.00252698
R23925 CSoutput.n242 CSoutput.n137 0.00252698
R23926 CSoutput.n163 CSoutput.n162 0.00252698
R23927 CSoutput.n156 CSoutput.n155 0.00252698
R23928 CSoutput.n239 CSoutput.n238 0.00252698
R23929 CSoutput.n166 CSoutput.n165 0.00252698
R23930 CSoutput.n169 CSoutput.n168 0.00252698
R23931 CSoutput.n150 CSoutput.n137 0.00252698
R23932 CSoutput.n217 CSoutput.n187 0.00252698
R23933 CSoutput.n216 CSoutput.n186 0.00252698
R23934 CSoutput.n215 CSoutput.n171 0.00252698
R23935 CSoutput.n212 CSoutput.n182 0.00252698
R23936 CSoutput.n219 CSoutput.n214 0.00252698
R23937 CSoutput.n228 CSoutput.n221 0.00252698
R23938 CSoutput.n217 CSoutput.n206 0.00252698
R23939 CSoutput.n216 CSoutput.n208 0.00252698
R23940 CSoutput.n215 CSoutput.n210 0.00252698
R23941 CSoutput.n230 CSoutput.n182 0.00252698
R23942 CSoutput.n219 CSoutput.n184 0.00252698
R23943 CSoutput.n221 CSoutput.n183 0.00252698
R23944 CSoutput.n129 CSoutput.n123 0.00252698
R23945 CSoutput.n122 CSoutput.n120 0.00252698
R23946 CSoutput.n248 CSoutput.n247 0.00252698
R23947 CSoutput.n132 CSoutput.n130 0.00252698
R23948 CSoutput.n135 CSoutput.n133 0.00252698
R23949 CSoutput.n252 CSoutput.n103 0.00252698
R23950 CSoutput.n129 CSoutput.n128 0.00252698
R23951 CSoutput.n122 CSoutput.n121 0.00252698
R23952 CSoutput.n249 CSoutput.n248 0.00252698
R23953 CSoutput.n132 CSoutput.n131 0.00252698
R23954 CSoutput.n135 CSoutput.n134 0.00252698
R23955 CSoutput.n116 CSoutput.n103 0.00252698
R23956 CSoutput.n237 CSoutput.n236 0.0020275
R23957 CSoutput.n236 CSoutput.n235 0.0020275
R23958 CSoutput.n233 CSoutput.n171 0.0020275
R23959 CSoutput.n233 CSoutput.n232 0.0020275
R23960 CSoutput.n247 CSoutput.n246 0.0020275
R23961 CSoutput.n246 CSoutput.n245 0.0020275
R23962 CSoutput.n147 CSoutput.n146 0.00166668
R23963 CSoutput.n229 CSoutput.n185 0.00166668
R23964 CSoutput.n113 CSoutput.n112 0.00166668
R23965 CSoutput.n251 CSoutput.n113 0.00133328
R23966 CSoutput.n185 CSoutput.n181 0.00133328
R23967 CSoutput.n241 CSoutput.n147 0.00133328
R23968 CSoutput.n244 CSoutput.n136 0.001
R23969 CSoutput.n222 CSoutput.n136 0.001
R23970 CSoutput.n124 CSoutput.n104 0.001
R23971 CSoutput.n223 CSoutput.n104 0.001
R23972 CSoutput.n125 CSoutput.n105 0.001
R23973 CSoutput.n224 CSoutput.n105 0.001
R23974 CSoutput.n126 CSoutput.n106 0.001
R23975 CSoutput.n225 CSoutput.n106 0.001
R23976 CSoutput.n127 CSoutput.n107 0.001
R23977 CSoutput.n226 CSoutput.n107 0.001
R23978 CSoutput.n220 CSoutput.n172 0.001
R23979 CSoutput.n220 CSoutput.n218 0.001
R23980 CSoutput.n202 CSoutput.n173 0.001
R23981 CSoutput.n196 CSoutput.n173 0.001
R23982 CSoutput.n203 CSoutput.n174 0.001
R23983 CSoutput.n197 CSoutput.n174 0.001
R23984 CSoutput.n204 CSoutput.n175 0.001
R23985 CSoutput.n198 CSoutput.n175 0.001
R23986 CSoutput.n205 CSoutput.n176 0.001
R23987 CSoutput.n199 CSoutput.n176 0.001
R23988 CSoutput.n234 CSoutput.n170 0.001
R23989 CSoutput.n188 CSoutput.n170 0.001
R23990 CSoutput.n158 CSoutput.n138 0.001
R23991 CSoutput.n189 CSoutput.n138 0.001
R23992 CSoutput.n159 CSoutput.n139 0.001
R23993 CSoutput.n190 CSoutput.n139 0.001
R23994 CSoutput.n160 CSoutput.n140 0.001
R23995 CSoutput.n191 CSoutput.n140 0.001
R23996 CSoutput.n161 CSoutput.n141 0.001
R23997 CSoutput.n192 CSoutput.n141 0.001
R23998 CSoutput.n192 CSoutput.n142 0.001
R23999 CSoutput.n191 CSoutput.n143 0.001
R24000 CSoutput.n190 CSoutput.n144 0.001
R24001 CSoutput.n189 CSoutput.t172 0.001
R24002 CSoutput.n188 CSoutput.n145 0.001
R24003 CSoutput.n161 CSoutput.n143 0.001
R24004 CSoutput.n160 CSoutput.n144 0.001
R24005 CSoutput.n159 CSoutput.t172 0.001
R24006 CSoutput.n158 CSoutput.n145 0.001
R24007 CSoutput.n234 CSoutput.n146 0.001
R24008 CSoutput.n199 CSoutput.n177 0.001
R24009 CSoutput.n198 CSoutput.n178 0.001
R24010 CSoutput.n197 CSoutput.n179 0.001
R24011 CSoutput.n196 CSoutput.t176 0.001
R24012 CSoutput.n218 CSoutput.n180 0.001
R24013 CSoutput.n205 CSoutput.n178 0.001
R24014 CSoutput.n204 CSoutput.n179 0.001
R24015 CSoutput.n203 CSoutput.t176 0.001
R24016 CSoutput.n202 CSoutput.n180 0.001
R24017 CSoutput.n229 CSoutput.n172 0.001
R24018 CSoutput.n226 CSoutput.n108 0.001
R24019 CSoutput.n225 CSoutput.n109 0.001
R24020 CSoutput.n224 CSoutput.n110 0.001
R24021 CSoutput.n223 CSoutput.t177 0.001
R24022 CSoutput.n222 CSoutput.n111 0.001
R24023 CSoutput.n127 CSoutput.n109 0.001
R24024 CSoutput.n126 CSoutput.n110 0.001
R24025 CSoutput.n125 CSoutput.t177 0.001
R24026 CSoutput.n124 CSoutput.n111 0.001
R24027 CSoutput.n244 CSoutput.n112 0.001
R24028 minus.n53 minus.t28 323.478
R24029 minus.n11 minus.t8 323.478
R24030 minus.n82 minus.t13 297.12
R24031 minus.n80 minus.t15 297.12
R24032 minus.n44 minus.t5 297.12
R24033 minus.n74 minus.t6 297.12
R24034 minus.n46 minus.t26 297.12
R24035 minus.n68 minus.t21 297.12
R24036 minus.n48 minus.t23 297.12
R24037 minus.n62 minus.t16 297.12
R24038 minus.n50 minus.t17 297.12
R24039 minus.n56 minus.t9 297.12
R24040 minus.n52 minus.t27 297.12
R24041 minus.n10 minus.t7 297.12
R24042 minus.n14 minus.t11 297.12
R24043 minus.n16 minus.t10 297.12
R24044 minus.n20 minus.t12 297.12
R24045 minus.n22 minus.t20 297.12
R24046 minus.n26 minus.t18 297.12
R24047 minus.n28 minus.t25 297.12
R24048 minus.n32 minus.t24 297.12
R24049 minus.n34 minus.t14 297.12
R24050 minus.n38 minus.t22 297.12
R24051 minus.n40 minus.t19 297.12
R24052 minus.n88 minus.t2 243.255
R24053 minus.n87 minus.n85 224.169
R24054 minus.n87 minus.n86 223.454
R24055 minus.n55 minus.n54 161.3
R24056 minus.n56 minus.n51 161.3
R24057 minus.n58 minus.n57 161.3
R24058 minus.n59 minus.n50 161.3
R24059 minus.n61 minus.n60 161.3
R24060 minus.n62 minus.n49 161.3
R24061 minus.n64 minus.n63 161.3
R24062 minus.n65 minus.n48 161.3
R24063 minus.n67 minus.n66 161.3
R24064 minus.n68 minus.n47 161.3
R24065 minus.n70 minus.n69 161.3
R24066 minus.n71 minus.n46 161.3
R24067 minus.n73 minus.n72 161.3
R24068 minus.n74 minus.n45 161.3
R24069 minus.n76 minus.n75 161.3
R24070 minus.n77 minus.n44 161.3
R24071 minus.n79 minus.n78 161.3
R24072 minus.n80 minus.n43 161.3
R24073 minus.n81 minus.n42 161.3
R24074 minus.n83 minus.n82 161.3
R24075 minus.n41 minus.n40 161.3
R24076 minus.n39 minus.n0 161.3
R24077 minus.n38 minus.n37 161.3
R24078 minus.n36 minus.n1 161.3
R24079 minus.n35 minus.n34 161.3
R24080 minus.n33 minus.n2 161.3
R24081 minus.n32 minus.n31 161.3
R24082 minus.n30 minus.n3 161.3
R24083 minus.n29 minus.n28 161.3
R24084 minus.n27 minus.n4 161.3
R24085 minus.n26 minus.n25 161.3
R24086 minus.n24 minus.n5 161.3
R24087 minus.n23 minus.n22 161.3
R24088 minus.n21 minus.n6 161.3
R24089 minus.n20 minus.n19 161.3
R24090 minus.n18 minus.n7 161.3
R24091 minus.n17 minus.n16 161.3
R24092 minus.n15 minus.n8 161.3
R24093 minus.n14 minus.n13 161.3
R24094 minus.n12 minus.n9 161.3
R24095 minus.n82 minus.n81 46.0096
R24096 minus.n40 minus.n39 46.0096
R24097 minus.n12 minus.n11 45.0871
R24098 minus.n54 minus.n53 45.0871
R24099 minus.n80 minus.n79 41.6278
R24100 minus.n55 minus.n52 41.6278
R24101 minus.n10 minus.n9 41.6278
R24102 minus.n38 minus.n1 41.6278
R24103 minus.n75 minus.n44 37.246
R24104 minus.n57 minus.n56 37.246
R24105 minus.n15 minus.n14 37.246
R24106 minus.n34 minus.n33 37.246
R24107 minus.n84 minus.n83 33.3925
R24108 minus.n74 minus.n73 32.8641
R24109 minus.n61 minus.n50 32.8641
R24110 minus.n16 minus.n7 32.8641
R24111 minus.n32 minus.n3 32.8641
R24112 minus.n69 minus.n46 28.4823
R24113 minus.n63 minus.n62 28.4823
R24114 minus.n21 minus.n20 28.4823
R24115 minus.n28 minus.n27 28.4823
R24116 minus.n68 minus.n67 24.1005
R24117 minus.n67 minus.n48 24.1005
R24118 minus.n22 minus.n5 24.1005
R24119 minus.n26 minus.n5 24.1005
R24120 minus.n86 minus.t4 19.8005
R24121 minus.n86 minus.t3 19.8005
R24122 minus.n85 minus.t1 19.8005
R24123 minus.n85 minus.t0 19.8005
R24124 minus.n69 minus.n68 19.7187
R24125 minus.n63 minus.n48 19.7187
R24126 minus.n22 minus.n21 19.7187
R24127 minus.n27 minus.n26 19.7187
R24128 minus.n73 minus.n46 15.3369
R24129 minus.n62 minus.n61 15.3369
R24130 minus.n20 minus.n7 15.3369
R24131 minus.n28 minus.n3 15.3369
R24132 minus.n53 minus.n52 14.1472
R24133 minus.n11 minus.n10 14.1472
R24134 minus.n84 minus.n41 12.0933
R24135 minus minus.n89 12.0331
R24136 minus.n75 minus.n74 10.955
R24137 minus.n57 minus.n50 10.955
R24138 minus.n16 minus.n15 10.955
R24139 minus.n33 minus.n32 10.955
R24140 minus.n79 minus.n44 6.57323
R24141 minus.n56 minus.n55 6.57323
R24142 minus.n14 minus.n9 6.57323
R24143 minus.n34 minus.n1 6.57323
R24144 minus.n89 minus.n88 4.80222
R24145 minus.n81 minus.n80 2.19141
R24146 minus.n39 minus.n38 2.19141
R24147 minus.n89 minus.n84 0.972091
R24148 minus.n88 minus.n87 0.716017
R24149 minus.n83 minus.n42 0.189894
R24150 minus.n43 minus.n42 0.189894
R24151 minus.n78 minus.n43 0.189894
R24152 minus.n78 minus.n77 0.189894
R24153 minus.n77 minus.n76 0.189894
R24154 minus.n76 minus.n45 0.189894
R24155 minus.n72 minus.n45 0.189894
R24156 minus.n72 minus.n71 0.189894
R24157 minus.n71 minus.n70 0.189894
R24158 minus.n70 minus.n47 0.189894
R24159 minus.n66 minus.n47 0.189894
R24160 minus.n66 minus.n65 0.189894
R24161 minus.n65 minus.n64 0.189894
R24162 minus.n64 minus.n49 0.189894
R24163 minus.n60 minus.n49 0.189894
R24164 minus.n60 minus.n59 0.189894
R24165 minus.n59 minus.n58 0.189894
R24166 minus.n58 minus.n51 0.189894
R24167 minus.n54 minus.n51 0.189894
R24168 minus.n13 minus.n12 0.189894
R24169 minus.n13 minus.n8 0.189894
R24170 minus.n17 minus.n8 0.189894
R24171 minus.n18 minus.n17 0.189894
R24172 minus.n19 minus.n18 0.189894
R24173 minus.n19 minus.n6 0.189894
R24174 minus.n23 minus.n6 0.189894
R24175 minus.n24 minus.n23 0.189894
R24176 minus.n25 minus.n24 0.189894
R24177 minus.n25 minus.n4 0.189894
R24178 minus.n29 minus.n4 0.189894
R24179 minus.n30 minus.n29 0.189894
R24180 minus.n31 minus.n30 0.189894
R24181 minus.n31 minus.n2 0.189894
R24182 minus.n35 minus.n2 0.189894
R24183 minus.n36 minus.n35 0.189894
R24184 minus.n37 minus.n36 0.189894
R24185 minus.n37 minus.n0 0.189894
R24186 minus.n41 minus.n0 0.189894
R24187 diffpairibias.n0 diffpairibias.t27 436.822
R24188 diffpairibias.n27 diffpairibias.t24 435.479
R24189 diffpairibias.n26 diffpairibias.t21 435.479
R24190 diffpairibias.n25 diffpairibias.t22 435.479
R24191 diffpairibias.n24 diffpairibias.t26 435.479
R24192 diffpairibias.n23 diffpairibias.t20 435.479
R24193 diffpairibias.n0 diffpairibias.t23 435.479
R24194 diffpairibias.n1 diffpairibias.t28 435.479
R24195 diffpairibias.n2 diffpairibias.t25 435.479
R24196 diffpairibias.n3 diffpairibias.t29 435.479
R24197 diffpairibias.n13 diffpairibias.t14 377.536
R24198 diffpairibias.n13 diffpairibias.t0 376.193
R24199 diffpairibias.n14 diffpairibias.t10 376.193
R24200 diffpairibias.n15 diffpairibias.t12 376.193
R24201 diffpairibias.n16 diffpairibias.t6 376.193
R24202 diffpairibias.n17 diffpairibias.t2 376.193
R24203 diffpairibias.n18 diffpairibias.t16 376.193
R24204 diffpairibias.n19 diffpairibias.t4 376.193
R24205 diffpairibias.n20 diffpairibias.t18 376.193
R24206 diffpairibias.n21 diffpairibias.t8 376.193
R24207 diffpairibias.n4 diffpairibias.t15 113.368
R24208 diffpairibias.n4 diffpairibias.t1 112.698
R24209 diffpairibias.n5 diffpairibias.t11 112.698
R24210 diffpairibias.n6 diffpairibias.t13 112.698
R24211 diffpairibias.n7 diffpairibias.t7 112.698
R24212 diffpairibias.n8 diffpairibias.t3 112.698
R24213 diffpairibias.n9 diffpairibias.t17 112.698
R24214 diffpairibias.n10 diffpairibias.t5 112.698
R24215 diffpairibias.n11 diffpairibias.t19 112.698
R24216 diffpairibias.n12 diffpairibias.t9 112.698
R24217 diffpairibias.n22 diffpairibias.n21 4.77242
R24218 diffpairibias.n22 diffpairibias.n12 4.30807
R24219 diffpairibias.n23 diffpairibias.n22 4.13945
R24220 diffpairibias.n21 diffpairibias.n20 1.34352
R24221 diffpairibias.n20 diffpairibias.n19 1.34352
R24222 diffpairibias.n19 diffpairibias.n18 1.34352
R24223 diffpairibias.n18 diffpairibias.n17 1.34352
R24224 diffpairibias.n17 diffpairibias.n16 1.34352
R24225 diffpairibias.n16 diffpairibias.n15 1.34352
R24226 diffpairibias.n15 diffpairibias.n14 1.34352
R24227 diffpairibias.n14 diffpairibias.n13 1.34352
R24228 diffpairibias.n3 diffpairibias.n2 1.34352
R24229 diffpairibias.n2 diffpairibias.n1 1.34352
R24230 diffpairibias.n1 diffpairibias.n0 1.34352
R24231 diffpairibias.n24 diffpairibias.n23 1.34352
R24232 diffpairibias.n25 diffpairibias.n24 1.34352
R24233 diffpairibias.n26 diffpairibias.n25 1.34352
R24234 diffpairibias.n27 diffpairibias.n26 1.34352
R24235 diffpairibias.n28 diffpairibias.n27 0.862419
R24236 diffpairibias diffpairibias.n28 0.684875
R24237 diffpairibias.n12 diffpairibias.n11 0.672012
R24238 diffpairibias.n11 diffpairibias.n10 0.672012
R24239 diffpairibias.n10 diffpairibias.n9 0.672012
R24240 diffpairibias.n9 diffpairibias.n8 0.672012
R24241 diffpairibias.n8 diffpairibias.n7 0.672012
R24242 diffpairibias.n7 diffpairibias.n6 0.672012
R24243 diffpairibias.n6 diffpairibias.n5 0.672012
R24244 diffpairibias.n5 diffpairibias.n4 0.672012
R24245 diffpairibias.n28 diffpairibias.n3 0.190907
R24246 a_n2982_8322.n12 a_n2982_8322.t3 74.6477
R24247 a_n2982_8322.n1 a_n2982_8322.t14 74.6477
R24248 a_n2982_8322.n28 a_n2982_8322.t29 74.6474
R24249 a_n2982_8322.n20 a_n2982_8322.t9 74.2899
R24250 a_n2982_8322.n13 a_n2982_8322.t1 74.2899
R24251 a_n2982_8322.n14 a_n2982_8322.t4 74.2899
R24252 a_n2982_8322.n17 a_n2982_8322.t5 74.2899
R24253 a_n2982_8322.n10 a_n2982_8322.t8 74.2899
R24254 a_n2982_8322.n28 a_n2982_8322.n27 70.6783
R24255 a_n2982_8322.n26 a_n2982_8322.n25 70.6783
R24256 a_n2982_8322.n24 a_n2982_8322.n23 70.6783
R24257 a_n2982_8322.n22 a_n2982_8322.n21 70.6783
R24258 a_n2982_8322.n12 a_n2982_8322.n11 70.6783
R24259 a_n2982_8322.n16 a_n2982_8322.n15 70.6783
R24260 a_n2982_8322.n1 a_n2982_8322.n0 70.6783
R24261 a_n2982_8322.n3 a_n2982_8322.n2 70.6783
R24262 a_n2982_8322.n5 a_n2982_8322.n4 70.6783
R24263 a_n2982_8322.n7 a_n2982_8322.n6 70.6783
R24264 a_n2982_8322.n9 a_n2982_8322.n8 70.6783
R24265 a_n2982_8322.n30 a_n2982_8322.n29 70.6782
R24266 a_n2982_8322.n18 a_n2982_8322.n10 24.9022
R24267 a_n2982_8322.n19 a_n2982_8322.t32 9.96358
R24268 a_n2982_8322.n18 a_n2982_8322.n17 8.38735
R24269 a_n2982_8322.n20 a_n2982_8322.n19 6.90998
R24270 a_n2982_8322.n19 a_n2982_8322.n18 5.3452
R24271 a_n2982_8322.n27 a_n2982_8322.t22 3.61217
R24272 a_n2982_8322.n27 a_n2982_8322.t18 3.61217
R24273 a_n2982_8322.n25 a_n2982_8322.t28 3.61217
R24274 a_n2982_8322.n25 a_n2982_8322.t16 3.61217
R24275 a_n2982_8322.n23 a_n2982_8322.t13 3.61217
R24276 a_n2982_8322.n23 a_n2982_8322.t12 3.61217
R24277 a_n2982_8322.n21 a_n2982_8322.t26 3.61217
R24278 a_n2982_8322.n21 a_n2982_8322.t25 3.61217
R24279 a_n2982_8322.n11 a_n2982_8322.t7 3.61217
R24280 a_n2982_8322.n11 a_n2982_8322.t6 3.61217
R24281 a_n2982_8322.n15 a_n2982_8322.t2 3.61217
R24282 a_n2982_8322.n15 a_n2982_8322.t0 3.61217
R24283 a_n2982_8322.n0 a_n2982_8322.t27 3.61217
R24284 a_n2982_8322.n0 a_n2982_8322.t23 3.61217
R24285 a_n2982_8322.n2 a_n2982_8322.t30 3.61217
R24286 a_n2982_8322.n2 a_n2982_8322.t20 3.61217
R24287 a_n2982_8322.n4 a_n2982_8322.t11 3.61217
R24288 a_n2982_8322.n4 a_n2982_8322.t10 3.61217
R24289 a_n2982_8322.n6 a_n2982_8322.t24 3.61217
R24290 a_n2982_8322.n6 a_n2982_8322.t17 3.61217
R24291 a_n2982_8322.n8 a_n2982_8322.t21 3.61217
R24292 a_n2982_8322.n8 a_n2982_8322.t19 3.61217
R24293 a_n2982_8322.n30 a_n2982_8322.t15 3.61217
R24294 a_n2982_8322.t31 a_n2982_8322.n30 3.61217
R24295 a_n2982_8322.n17 a_n2982_8322.n16 0.358259
R24296 a_n2982_8322.n16 a_n2982_8322.n14 0.358259
R24297 a_n2982_8322.n13 a_n2982_8322.n12 0.358259
R24298 a_n2982_8322.n10 a_n2982_8322.n9 0.358259
R24299 a_n2982_8322.n9 a_n2982_8322.n7 0.358259
R24300 a_n2982_8322.n7 a_n2982_8322.n5 0.358259
R24301 a_n2982_8322.n5 a_n2982_8322.n3 0.358259
R24302 a_n2982_8322.n3 a_n2982_8322.n1 0.358259
R24303 a_n2982_8322.n22 a_n2982_8322.n20 0.358259
R24304 a_n2982_8322.n24 a_n2982_8322.n22 0.358259
R24305 a_n2982_8322.n26 a_n2982_8322.n24 0.358259
R24306 a_n2982_8322.n29 a_n2982_8322.n26 0.358259
R24307 a_n2982_8322.n29 a_n2982_8322.n28 0.358259
R24308 a_n2982_8322.n14 a_n2982_8322.n13 0.101793
R24309 a_n2982_8322.t37 a_n2982_8322.t34 0.0788333
R24310 a_n2982_8322.t36 a_n2982_8322.t35 0.0788333
R24311 a_n2982_8322.t32 a_n2982_8322.t33 0.0788333
R24312 a_n2982_8322.t36 a_n2982_8322.t37 0.0318333
R24313 a_n2982_8322.t32 a_n2982_8322.t35 0.0318333
R24314 a_n2982_8322.t34 a_n2982_8322.t35 0.0318333
R24315 a_n2982_8322.t33 a_n2982_8322.t36 0.0318333
R24316 outputibias.n27 outputibias.n1 289.615
R24317 outputibias.n58 outputibias.n32 289.615
R24318 outputibias.n90 outputibias.n64 289.615
R24319 outputibias.n122 outputibias.n96 289.615
R24320 outputibias.n28 outputibias.n27 185
R24321 outputibias.n26 outputibias.n25 185
R24322 outputibias.n5 outputibias.n4 185
R24323 outputibias.n20 outputibias.n19 185
R24324 outputibias.n18 outputibias.n17 185
R24325 outputibias.n9 outputibias.n8 185
R24326 outputibias.n12 outputibias.n11 185
R24327 outputibias.n59 outputibias.n58 185
R24328 outputibias.n57 outputibias.n56 185
R24329 outputibias.n36 outputibias.n35 185
R24330 outputibias.n51 outputibias.n50 185
R24331 outputibias.n49 outputibias.n48 185
R24332 outputibias.n40 outputibias.n39 185
R24333 outputibias.n43 outputibias.n42 185
R24334 outputibias.n91 outputibias.n90 185
R24335 outputibias.n89 outputibias.n88 185
R24336 outputibias.n68 outputibias.n67 185
R24337 outputibias.n83 outputibias.n82 185
R24338 outputibias.n81 outputibias.n80 185
R24339 outputibias.n72 outputibias.n71 185
R24340 outputibias.n75 outputibias.n74 185
R24341 outputibias.n123 outputibias.n122 185
R24342 outputibias.n121 outputibias.n120 185
R24343 outputibias.n100 outputibias.n99 185
R24344 outputibias.n115 outputibias.n114 185
R24345 outputibias.n113 outputibias.n112 185
R24346 outputibias.n104 outputibias.n103 185
R24347 outputibias.n107 outputibias.n106 185
R24348 outputibias.n0 outputibias.t11 178.945
R24349 outputibias.n133 outputibias.t8 177.018
R24350 outputibias.n132 outputibias.t10 177.018
R24351 outputibias.n0 outputibias.t9 177.018
R24352 outputibias.t5 outputibias.n10 147.661
R24353 outputibias.t7 outputibias.n41 147.661
R24354 outputibias.t3 outputibias.n73 147.661
R24355 outputibias.t1 outputibias.n105 147.661
R24356 outputibias.n128 outputibias.t4 132.363
R24357 outputibias.n128 outputibias.t6 130.436
R24358 outputibias.n129 outputibias.t2 130.436
R24359 outputibias.n130 outputibias.t0 130.436
R24360 outputibias.n27 outputibias.n26 104.615
R24361 outputibias.n26 outputibias.n4 104.615
R24362 outputibias.n19 outputibias.n4 104.615
R24363 outputibias.n19 outputibias.n18 104.615
R24364 outputibias.n18 outputibias.n8 104.615
R24365 outputibias.n11 outputibias.n8 104.615
R24366 outputibias.n58 outputibias.n57 104.615
R24367 outputibias.n57 outputibias.n35 104.615
R24368 outputibias.n50 outputibias.n35 104.615
R24369 outputibias.n50 outputibias.n49 104.615
R24370 outputibias.n49 outputibias.n39 104.615
R24371 outputibias.n42 outputibias.n39 104.615
R24372 outputibias.n90 outputibias.n89 104.615
R24373 outputibias.n89 outputibias.n67 104.615
R24374 outputibias.n82 outputibias.n67 104.615
R24375 outputibias.n82 outputibias.n81 104.615
R24376 outputibias.n81 outputibias.n71 104.615
R24377 outputibias.n74 outputibias.n71 104.615
R24378 outputibias.n122 outputibias.n121 104.615
R24379 outputibias.n121 outputibias.n99 104.615
R24380 outputibias.n114 outputibias.n99 104.615
R24381 outputibias.n114 outputibias.n113 104.615
R24382 outputibias.n113 outputibias.n103 104.615
R24383 outputibias.n106 outputibias.n103 104.615
R24384 outputibias.n63 outputibias.n31 95.6354
R24385 outputibias.n63 outputibias.n62 94.6732
R24386 outputibias.n95 outputibias.n94 94.6732
R24387 outputibias.n127 outputibias.n126 94.6732
R24388 outputibias.n11 outputibias.t5 52.3082
R24389 outputibias.n42 outputibias.t7 52.3082
R24390 outputibias.n74 outputibias.t3 52.3082
R24391 outputibias.n106 outputibias.t1 52.3082
R24392 outputibias.n12 outputibias.n10 15.6674
R24393 outputibias.n43 outputibias.n41 15.6674
R24394 outputibias.n75 outputibias.n73 15.6674
R24395 outputibias.n107 outputibias.n105 15.6674
R24396 outputibias.n13 outputibias.n9 12.8005
R24397 outputibias.n44 outputibias.n40 12.8005
R24398 outputibias.n76 outputibias.n72 12.8005
R24399 outputibias.n108 outputibias.n104 12.8005
R24400 outputibias.n17 outputibias.n16 12.0247
R24401 outputibias.n48 outputibias.n47 12.0247
R24402 outputibias.n80 outputibias.n79 12.0247
R24403 outputibias.n112 outputibias.n111 12.0247
R24404 outputibias.n20 outputibias.n7 11.249
R24405 outputibias.n51 outputibias.n38 11.249
R24406 outputibias.n83 outputibias.n70 11.249
R24407 outputibias.n115 outputibias.n102 11.249
R24408 outputibias.n21 outputibias.n5 10.4732
R24409 outputibias.n52 outputibias.n36 10.4732
R24410 outputibias.n84 outputibias.n68 10.4732
R24411 outputibias.n116 outputibias.n100 10.4732
R24412 outputibias.n25 outputibias.n24 9.69747
R24413 outputibias.n56 outputibias.n55 9.69747
R24414 outputibias.n88 outputibias.n87 9.69747
R24415 outputibias.n120 outputibias.n119 9.69747
R24416 outputibias.n31 outputibias.n30 9.45567
R24417 outputibias.n62 outputibias.n61 9.45567
R24418 outputibias.n94 outputibias.n93 9.45567
R24419 outputibias.n126 outputibias.n125 9.45567
R24420 outputibias.n30 outputibias.n29 9.3005
R24421 outputibias.n3 outputibias.n2 9.3005
R24422 outputibias.n24 outputibias.n23 9.3005
R24423 outputibias.n22 outputibias.n21 9.3005
R24424 outputibias.n7 outputibias.n6 9.3005
R24425 outputibias.n16 outputibias.n15 9.3005
R24426 outputibias.n14 outputibias.n13 9.3005
R24427 outputibias.n61 outputibias.n60 9.3005
R24428 outputibias.n34 outputibias.n33 9.3005
R24429 outputibias.n55 outputibias.n54 9.3005
R24430 outputibias.n53 outputibias.n52 9.3005
R24431 outputibias.n38 outputibias.n37 9.3005
R24432 outputibias.n47 outputibias.n46 9.3005
R24433 outputibias.n45 outputibias.n44 9.3005
R24434 outputibias.n93 outputibias.n92 9.3005
R24435 outputibias.n66 outputibias.n65 9.3005
R24436 outputibias.n87 outputibias.n86 9.3005
R24437 outputibias.n85 outputibias.n84 9.3005
R24438 outputibias.n70 outputibias.n69 9.3005
R24439 outputibias.n79 outputibias.n78 9.3005
R24440 outputibias.n77 outputibias.n76 9.3005
R24441 outputibias.n125 outputibias.n124 9.3005
R24442 outputibias.n98 outputibias.n97 9.3005
R24443 outputibias.n119 outputibias.n118 9.3005
R24444 outputibias.n117 outputibias.n116 9.3005
R24445 outputibias.n102 outputibias.n101 9.3005
R24446 outputibias.n111 outputibias.n110 9.3005
R24447 outputibias.n109 outputibias.n108 9.3005
R24448 outputibias.n28 outputibias.n3 8.92171
R24449 outputibias.n59 outputibias.n34 8.92171
R24450 outputibias.n91 outputibias.n66 8.92171
R24451 outputibias.n123 outputibias.n98 8.92171
R24452 outputibias.n29 outputibias.n1 8.14595
R24453 outputibias.n60 outputibias.n32 8.14595
R24454 outputibias.n92 outputibias.n64 8.14595
R24455 outputibias.n124 outputibias.n96 8.14595
R24456 outputibias.n31 outputibias.n1 5.81868
R24457 outputibias.n62 outputibias.n32 5.81868
R24458 outputibias.n94 outputibias.n64 5.81868
R24459 outputibias.n126 outputibias.n96 5.81868
R24460 outputibias.n131 outputibias.n130 5.20947
R24461 outputibias.n29 outputibias.n28 5.04292
R24462 outputibias.n60 outputibias.n59 5.04292
R24463 outputibias.n92 outputibias.n91 5.04292
R24464 outputibias.n124 outputibias.n123 5.04292
R24465 outputibias.n131 outputibias.n127 4.42209
R24466 outputibias.n14 outputibias.n10 4.38594
R24467 outputibias.n45 outputibias.n41 4.38594
R24468 outputibias.n77 outputibias.n73 4.38594
R24469 outputibias.n109 outputibias.n105 4.38594
R24470 outputibias.n132 outputibias.n131 4.28454
R24471 outputibias.n25 outputibias.n3 4.26717
R24472 outputibias.n56 outputibias.n34 4.26717
R24473 outputibias.n88 outputibias.n66 4.26717
R24474 outputibias.n120 outputibias.n98 4.26717
R24475 outputibias.n24 outputibias.n5 3.49141
R24476 outputibias.n55 outputibias.n36 3.49141
R24477 outputibias.n87 outputibias.n68 3.49141
R24478 outputibias.n119 outputibias.n100 3.49141
R24479 outputibias.n21 outputibias.n20 2.71565
R24480 outputibias.n52 outputibias.n51 2.71565
R24481 outputibias.n84 outputibias.n83 2.71565
R24482 outputibias.n116 outputibias.n115 2.71565
R24483 outputibias.n17 outputibias.n7 1.93989
R24484 outputibias.n48 outputibias.n38 1.93989
R24485 outputibias.n80 outputibias.n70 1.93989
R24486 outputibias.n112 outputibias.n102 1.93989
R24487 outputibias.n130 outputibias.n129 1.9266
R24488 outputibias.n129 outputibias.n128 1.9266
R24489 outputibias.n133 outputibias.n132 1.92658
R24490 outputibias.n134 outputibias.n133 1.29913
R24491 outputibias.n16 outputibias.n9 1.16414
R24492 outputibias.n47 outputibias.n40 1.16414
R24493 outputibias.n79 outputibias.n72 1.16414
R24494 outputibias.n111 outputibias.n104 1.16414
R24495 outputibias.n127 outputibias.n95 0.962709
R24496 outputibias.n95 outputibias.n63 0.962709
R24497 outputibias.n13 outputibias.n12 0.388379
R24498 outputibias.n44 outputibias.n43 0.388379
R24499 outputibias.n76 outputibias.n75 0.388379
R24500 outputibias.n108 outputibias.n107 0.388379
R24501 outputibias.n134 outputibias.n0 0.337251
R24502 outputibias outputibias.n134 0.302375
R24503 outputibias.n30 outputibias.n2 0.155672
R24504 outputibias.n23 outputibias.n2 0.155672
R24505 outputibias.n23 outputibias.n22 0.155672
R24506 outputibias.n22 outputibias.n6 0.155672
R24507 outputibias.n15 outputibias.n6 0.155672
R24508 outputibias.n15 outputibias.n14 0.155672
R24509 outputibias.n61 outputibias.n33 0.155672
R24510 outputibias.n54 outputibias.n33 0.155672
R24511 outputibias.n54 outputibias.n53 0.155672
R24512 outputibias.n53 outputibias.n37 0.155672
R24513 outputibias.n46 outputibias.n37 0.155672
R24514 outputibias.n46 outputibias.n45 0.155672
R24515 outputibias.n93 outputibias.n65 0.155672
R24516 outputibias.n86 outputibias.n65 0.155672
R24517 outputibias.n86 outputibias.n85 0.155672
R24518 outputibias.n85 outputibias.n69 0.155672
R24519 outputibias.n78 outputibias.n69 0.155672
R24520 outputibias.n78 outputibias.n77 0.155672
R24521 outputibias.n125 outputibias.n97 0.155672
R24522 outputibias.n118 outputibias.n97 0.155672
R24523 outputibias.n118 outputibias.n117 0.155672
R24524 outputibias.n117 outputibias.n101 0.155672
R24525 outputibias.n110 outputibias.n101 0.155672
R24526 outputibias.n110 outputibias.n109 0.155672
R24527 output.n41 output.n15 289.615
R24528 output.n72 output.n46 289.615
R24529 output.n104 output.n78 289.615
R24530 output.n136 output.n110 289.615
R24531 output.n77 output.n45 197.26
R24532 output.n77 output.n76 196.298
R24533 output.n109 output.n108 196.298
R24534 output.n141 output.n140 196.298
R24535 output.n42 output.n41 185
R24536 output.n40 output.n39 185
R24537 output.n19 output.n18 185
R24538 output.n34 output.n33 185
R24539 output.n32 output.n31 185
R24540 output.n23 output.n22 185
R24541 output.n26 output.n25 185
R24542 output.n73 output.n72 185
R24543 output.n71 output.n70 185
R24544 output.n50 output.n49 185
R24545 output.n65 output.n64 185
R24546 output.n63 output.n62 185
R24547 output.n54 output.n53 185
R24548 output.n57 output.n56 185
R24549 output.n105 output.n104 185
R24550 output.n103 output.n102 185
R24551 output.n82 output.n81 185
R24552 output.n97 output.n96 185
R24553 output.n95 output.n94 185
R24554 output.n86 output.n85 185
R24555 output.n89 output.n88 185
R24556 output.n137 output.n136 185
R24557 output.n135 output.n134 185
R24558 output.n114 output.n113 185
R24559 output.n129 output.n128 185
R24560 output.n127 output.n126 185
R24561 output.n118 output.n117 185
R24562 output.n121 output.n120 185
R24563 output.t0 output.n24 147.661
R24564 output.t2 output.n55 147.661
R24565 output.t3 output.n87 147.661
R24566 output.t1 output.n119 147.661
R24567 output.n41 output.n40 104.615
R24568 output.n40 output.n18 104.615
R24569 output.n33 output.n18 104.615
R24570 output.n33 output.n32 104.615
R24571 output.n32 output.n22 104.615
R24572 output.n25 output.n22 104.615
R24573 output.n72 output.n71 104.615
R24574 output.n71 output.n49 104.615
R24575 output.n64 output.n49 104.615
R24576 output.n64 output.n63 104.615
R24577 output.n63 output.n53 104.615
R24578 output.n56 output.n53 104.615
R24579 output.n104 output.n103 104.615
R24580 output.n103 output.n81 104.615
R24581 output.n96 output.n81 104.615
R24582 output.n96 output.n95 104.615
R24583 output.n95 output.n85 104.615
R24584 output.n88 output.n85 104.615
R24585 output.n136 output.n135 104.615
R24586 output.n135 output.n113 104.615
R24587 output.n128 output.n113 104.615
R24588 output.n128 output.n127 104.615
R24589 output.n127 output.n117 104.615
R24590 output.n120 output.n117 104.615
R24591 output.n1 output.t5 77.056
R24592 output.n14 output.t7 76.6694
R24593 output.n1 output.n0 72.7095
R24594 output.n3 output.n2 72.7095
R24595 output.n5 output.n4 72.7095
R24596 output.n7 output.n6 72.7095
R24597 output.n9 output.n8 72.7095
R24598 output.n11 output.n10 72.7095
R24599 output.n13 output.n12 72.7095
R24600 output.n25 output.t0 52.3082
R24601 output.n56 output.t2 52.3082
R24602 output.n88 output.t3 52.3082
R24603 output.n120 output.t1 52.3082
R24604 output.n26 output.n24 15.6674
R24605 output.n57 output.n55 15.6674
R24606 output.n89 output.n87 15.6674
R24607 output.n121 output.n119 15.6674
R24608 output.n27 output.n23 12.8005
R24609 output.n58 output.n54 12.8005
R24610 output.n90 output.n86 12.8005
R24611 output.n122 output.n118 12.8005
R24612 output.n31 output.n30 12.0247
R24613 output.n62 output.n61 12.0247
R24614 output.n94 output.n93 12.0247
R24615 output.n126 output.n125 12.0247
R24616 output.n34 output.n21 11.249
R24617 output.n65 output.n52 11.249
R24618 output.n97 output.n84 11.249
R24619 output.n129 output.n116 11.249
R24620 output.n35 output.n19 10.4732
R24621 output.n66 output.n50 10.4732
R24622 output.n98 output.n82 10.4732
R24623 output.n130 output.n114 10.4732
R24624 output.n39 output.n38 9.69747
R24625 output.n70 output.n69 9.69747
R24626 output.n102 output.n101 9.69747
R24627 output.n134 output.n133 9.69747
R24628 output.n45 output.n44 9.45567
R24629 output.n76 output.n75 9.45567
R24630 output.n108 output.n107 9.45567
R24631 output.n140 output.n139 9.45567
R24632 output.n44 output.n43 9.3005
R24633 output.n17 output.n16 9.3005
R24634 output.n38 output.n37 9.3005
R24635 output.n36 output.n35 9.3005
R24636 output.n21 output.n20 9.3005
R24637 output.n30 output.n29 9.3005
R24638 output.n28 output.n27 9.3005
R24639 output.n75 output.n74 9.3005
R24640 output.n48 output.n47 9.3005
R24641 output.n69 output.n68 9.3005
R24642 output.n67 output.n66 9.3005
R24643 output.n52 output.n51 9.3005
R24644 output.n61 output.n60 9.3005
R24645 output.n59 output.n58 9.3005
R24646 output.n107 output.n106 9.3005
R24647 output.n80 output.n79 9.3005
R24648 output.n101 output.n100 9.3005
R24649 output.n99 output.n98 9.3005
R24650 output.n84 output.n83 9.3005
R24651 output.n93 output.n92 9.3005
R24652 output.n91 output.n90 9.3005
R24653 output.n139 output.n138 9.3005
R24654 output.n112 output.n111 9.3005
R24655 output.n133 output.n132 9.3005
R24656 output.n131 output.n130 9.3005
R24657 output.n116 output.n115 9.3005
R24658 output.n125 output.n124 9.3005
R24659 output.n123 output.n122 9.3005
R24660 output.n42 output.n17 8.92171
R24661 output.n73 output.n48 8.92171
R24662 output.n105 output.n80 8.92171
R24663 output.n137 output.n112 8.92171
R24664 output output.n141 8.15037
R24665 output.n43 output.n15 8.14595
R24666 output.n74 output.n46 8.14595
R24667 output.n106 output.n78 8.14595
R24668 output.n138 output.n110 8.14595
R24669 output.n45 output.n15 5.81868
R24670 output.n76 output.n46 5.81868
R24671 output.n108 output.n78 5.81868
R24672 output.n140 output.n110 5.81868
R24673 output.n43 output.n42 5.04292
R24674 output.n74 output.n73 5.04292
R24675 output.n106 output.n105 5.04292
R24676 output.n138 output.n137 5.04292
R24677 output.n28 output.n24 4.38594
R24678 output.n59 output.n55 4.38594
R24679 output.n91 output.n87 4.38594
R24680 output.n123 output.n119 4.38594
R24681 output.n39 output.n17 4.26717
R24682 output.n70 output.n48 4.26717
R24683 output.n102 output.n80 4.26717
R24684 output.n134 output.n112 4.26717
R24685 output.n0 output.t11 3.9605
R24686 output.n0 output.t16 3.9605
R24687 output.n2 output.t4 3.9605
R24688 output.n2 output.t12 3.9605
R24689 output.n4 output.t14 3.9605
R24690 output.n4 output.t13 3.9605
R24691 output.n6 output.t19 3.9605
R24692 output.n6 output.t6 3.9605
R24693 output.n8 output.t8 3.9605
R24694 output.n8 output.t17 3.9605
R24695 output.n10 output.t18 3.9605
R24696 output.n10 output.t9 3.9605
R24697 output.n12 output.t10 3.9605
R24698 output.n12 output.t15 3.9605
R24699 output.n38 output.n19 3.49141
R24700 output.n69 output.n50 3.49141
R24701 output.n101 output.n82 3.49141
R24702 output.n133 output.n114 3.49141
R24703 output.n35 output.n34 2.71565
R24704 output.n66 output.n65 2.71565
R24705 output.n98 output.n97 2.71565
R24706 output.n130 output.n129 2.71565
R24707 output.n31 output.n21 1.93989
R24708 output.n62 output.n52 1.93989
R24709 output.n94 output.n84 1.93989
R24710 output.n126 output.n116 1.93989
R24711 output.n30 output.n23 1.16414
R24712 output.n61 output.n54 1.16414
R24713 output.n93 output.n86 1.16414
R24714 output.n125 output.n118 1.16414
R24715 output.n141 output.n109 0.962709
R24716 output.n109 output.n77 0.962709
R24717 output.n27 output.n26 0.388379
R24718 output.n58 output.n57 0.388379
R24719 output.n90 output.n89 0.388379
R24720 output.n122 output.n121 0.388379
R24721 output.n14 output.n13 0.387128
R24722 output.n13 output.n11 0.387128
R24723 output.n11 output.n9 0.387128
R24724 output.n9 output.n7 0.387128
R24725 output.n7 output.n5 0.387128
R24726 output.n5 output.n3 0.387128
R24727 output.n3 output.n1 0.387128
R24728 output.n44 output.n16 0.155672
R24729 output.n37 output.n16 0.155672
R24730 output.n37 output.n36 0.155672
R24731 output.n36 output.n20 0.155672
R24732 output.n29 output.n20 0.155672
R24733 output.n29 output.n28 0.155672
R24734 output.n75 output.n47 0.155672
R24735 output.n68 output.n47 0.155672
R24736 output.n68 output.n67 0.155672
R24737 output.n67 output.n51 0.155672
R24738 output.n60 output.n51 0.155672
R24739 output.n60 output.n59 0.155672
R24740 output.n107 output.n79 0.155672
R24741 output.n100 output.n79 0.155672
R24742 output.n100 output.n99 0.155672
R24743 output.n99 output.n83 0.155672
R24744 output.n92 output.n83 0.155672
R24745 output.n92 output.n91 0.155672
R24746 output.n139 output.n111 0.155672
R24747 output.n132 output.n111 0.155672
R24748 output.n132 output.n131 0.155672
R24749 output.n131 output.n115 0.155672
R24750 output.n124 output.n115 0.155672
R24751 output.n124 output.n123 0.155672
R24752 output output.n14 0.126227
C0 commonsourceibias outputibias 0.003832f
C1 plus diffpairibias 4.56e-19
C2 vdd commonsourceibias 0.004218f
C3 CSoutput plus 0.91196f
C4 commonsourceibias diffpairibias 0.064336f
C5 CSoutput commonsourceibias 66.8263f
C6 minus plus 10.303599f
C7 minus commonsourceibias 0.337549f
C8 plus commonsourceibias 0.283677f
C9 output outputibias 2.34152f
C10 vdd output 7.23429f
C11 CSoutput output 6.13881f
C12 CSoutput outputibias 0.032386f
C13 vdd CSoutput 68.5846f
C14 minus diffpairibias 4.33e-19
C15 commonsourceibias output 0.006808f
C16 CSoutput minus 3.17016f
C17 vdd plus 0.080016f
C18 diffpairibias gnd 60.00273f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.223205p
C22 plus gnd 37.775303f
C23 minus gnd 31.29577f
C24 CSoutput gnd 0.144715p
C25 vdd gnd 0.449105p
C26 output.t5 gnd 0.464308f
C27 output.t11 gnd 0.044422f
C28 output.t16 gnd 0.044422f
C29 output.n0 gnd 0.364624f
C30 output.n1 gnd 0.614102f
C31 output.t4 gnd 0.044422f
C32 output.t12 gnd 0.044422f
C33 output.n2 gnd 0.364624f
C34 output.n3 gnd 0.350265f
C35 output.t14 gnd 0.044422f
C36 output.t13 gnd 0.044422f
C37 output.n4 gnd 0.364624f
C38 output.n5 gnd 0.350265f
C39 output.t19 gnd 0.044422f
C40 output.t6 gnd 0.044422f
C41 output.n6 gnd 0.364624f
C42 output.n7 gnd 0.350265f
C43 output.t8 gnd 0.044422f
C44 output.t17 gnd 0.044422f
C45 output.n8 gnd 0.364624f
C46 output.n9 gnd 0.350265f
C47 output.t18 gnd 0.044422f
C48 output.t9 gnd 0.044422f
C49 output.n10 gnd 0.364624f
C50 output.n11 gnd 0.350265f
C51 output.t10 gnd 0.044422f
C52 output.t15 gnd 0.044422f
C53 output.n12 gnd 0.364624f
C54 output.n13 gnd 0.350265f
C55 output.t7 gnd 0.462979f
C56 output.n14 gnd 0.28994f
C57 output.n15 gnd 0.015803f
C58 output.n16 gnd 0.011243f
C59 output.n17 gnd 0.006041f
C60 output.n18 gnd 0.01428f
C61 output.n19 gnd 0.006397f
C62 output.n20 gnd 0.011243f
C63 output.n21 gnd 0.006041f
C64 output.n22 gnd 0.01428f
C65 output.n23 gnd 0.006397f
C66 output.n24 gnd 0.048111f
C67 output.t0 gnd 0.023274f
C68 output.n25 gnd 0.01071f
C69 output.n26 gnd 0.008435f
C70 output.n27 gnd 0.006041f
C71 output.n28 gnd 0.267512f
C72 output.n29 gnd 0.011243f
C73 output.n30 gnd 0.006041f
C74 output.n31 gnd 0.006397f
C75 output.n32 gnd 0.01428f
C76 output.n33 gnd 0.01428f
C77 output.n34 gnd 0.006397f
C78 output.n35 gnd 0.006041f
C79 output.n36 gnd 0.011243f
C80 output.n37 gnd 0.011243f
C81 output.n38 gnd 0.006041f
C82 output.n39 gnd 0.006397f
C83 output.n40 gnd 0.01428f
C84 output.n41 gnd 0.030913f
C85 output.n42 gnd 0.006397f
C86 output.n43 gnd 0.006041f
C87 output.n44 gnd 0.025987f
C88 output.n45 gnd 0.097665f
C89 output.n46 gnd 0.015803f
C90 output.n47 gnd 0.011243f
C91 output.n48 gnd 0.006041f
C92 output.n49 gnd 0.01428f
C93 output.n50 gnd 0.006397f
C94 output.n51 gnd 0.011243f
C95 output.n52 gnd 0.006041f
C96 output.n53 gnd 0.01428f
C97 output.n54 gnd 0.006397f
C98 output.n55 gnd 0.048111f
C99 output.t2 gnd 0.023274f
C100 output.n56 gnd 0.01071f
C101 output.n57 gnd 0.008435f
C102 output.n58 gnd 0.006041f
C103 output.n59 gnd 0.267512f
C104 output.n60 gnd 0.011243f
C105 output.n61 gnd 0.006041f
C106 output.n62 gnd 0.006397f
C107 output.n63 gnd 0.01428f
C108 output.n64 gnd 0.01428f
C109 output.n65 gnd 0.006397f
C110 output.n66 gnd 0.006041f
C111 output.n67 gnd 0.011243f
C112 output.n68 gnd 0.011243f
C113 output.n69 gnd 0.006041f
C114 output.n70 gnd 0.006397f
C115 output.n71 gnd 0.01428f
C116 output.n72 gnd 0.030913f
C117 output.n73 gnd 0.006397f
C118 output.n74 gnd 0.006041f
C119 output.n75 gnd 0.025987f
C120 output.n76 gnd 0.09306f
C121 output.n77 gnd 1.65264f
C122 output.n78 gnd 0.015803f
C123 output.n79 gnd 0.011243f
C124 output.n80 gnd 0.006041f
C125 output.n81 gnd 0.01428f
C126 output.n82 gnd 0.006397f
C127 output.n83 gnd 0.011243f
C128 output.n84 gnd 0.006041f
C129 output.n85 gnd 0.01428f
C130 output.n86 gnd 0.006397f
C131 output.n87 gnd 0.048111f
C132 output.t3 gnd 0.023274f
C133 output.n88 gnd 0.01071f
C134 output.n89 gnd 0.008435f
C135 output.n90 gnd 0.006041f
C136 output.n91 gnd 0.267512f
C137 output.n92 gnd 0.011243f
C138 output.n93 gnd 0.006041f
C139 output.n94 gnd 0.006397f
C140 output.n95 gnd 0.01428f
C141 output.n96 gnd 0.01428f
C142 output.n97 gnd 0.006397f
C143 output.n98 gnd 0.006041f
C144 output.n99 gnd 0.011243f
C145 output.n100 gnd 0.011243f
C146 output.n101 gnd 0.006041f
C147 output.n102 gnd 0.006397f
C148 output.n103 gnd 0.01428f
C149 output.n104 gnd 0.030913f
C150 output.n105 gnd 0.006397f
C151 output.n106 gnd 0.006041f
C152 output.n107 gnd 0.025987f
C153 output.n108 gnd 0.09306f
C154 output.n109 gnd 0.713089f
C155 output.n110 gnd 0.015803f
C156 output.n111 gnd 0.011243f
C157 output.n112 gnd 0.006041f
C158 output.n113 gnd 0.01428f
C159 output.n114 gnd 0.006397f
C160 output.n115 gnd 0.011243f
C161 output.n116 gnd 0.006041f
C162 output.n117 gnd 0.01428f
C163 output.n118 gnd 0.006397f
C164 output.n119 gnd 0.048111f
C165 output.t1 gnd 0.023274f
C166 output.n120 gnd 0.01071f
C167 output.n121 gnd 0.008435f
C168 output.n122 gnd 0.006041f
C169 output.n123 gnd 0.267512f
C170 output.n124 gnd 0.011243f
C171 output.n125 gnd 0.006041f
C172 output.n126 gnd 0.006397f
C173 output.n127 gnd 0.01428f
C174 output.n128 gnd 0.01428f
C175 output.n129 gnd 0.006397f
C176 output.n130 gnd 0.006041f
C177 output.n131 gnd 0.011243f
C178 output.n132 gnd 0.011243f
C179 output.n133 gnd 0.006041f
C180 output.n134 gnd 0.006397f
C181 output.n135 gnd 0.01428f
C182 output.n136 gnd 0.030913f
C183 output.n137 gnd 0.006397f
C184 output.n138 gnd 0.006041f
C185 output.n139 gnd 0.025987f
C186 output.n140 gnd 0.09306f
C187 output.n141 gnd 1.67353f
C188 outputibias.t9 gnd 0.11477f
C189 outputibias.t11 gnd 0.115567f
C190 outputibias.n0 gnd 0.130108f
C191 outputibias.n1 gnd 0.001372f
C192 outputibias.n2 gnd 9.76e-19
C193 outputibias.n3 gnd 5.24e-19
C194 outputibias.n4 gnd 0.001239f
C195 outputibias.n5 gnd 5.55e-19
C196 outputibias.n6 gnd 9.76e-19
C197 outputibias.n7 gnd 5.24e-19
C198 outputibias.n8 gnd 0.001239f
C199 outputibias.n9 gnd 5.55e-19
C200 outputibias.n10 gnd 0.004176f
C201 outputibias.t5 gnd 0.00202f
C202 outputibias.n11 gnd 9.3e-19
C203 outputibias.n12 gnd 7.32e-19
C204 outputibias.n13 gnd 5.24e-19
C205 outputibias.n14 gnd 0.02322f
C206 outputibias.n15 gnd 9.76e-19
C207 outputibias.n16 gnd 5.24e-19
C208 outputibias.n17 gnd 5.55e-19
C209 outputibias.n18 gnd 0.001239f
C210 outputibias.n19 gnd 0.001239f
C211 outputibias.n20 gnd 5.55e-19
C212 outputibias.n21 gnd 5.24e-19
C213 outputibias.n22 gnd 9.76e-19
C214 outputibias.n23 gnd 9.76e-19
C215 outputibias.n24 gnd 5.24e-19
C216 outputibias.n25 gnd 5.55e-19
C217 outputibias.n26 gnd 0.001239f
C218 outputibias.n27 gnd 0.002683f
C219 outputibias.n28 gnd 5.55e-19
C220 outputibias.n29 gnd 5.24e-19
C221 outputibias.n30 gnd 0.002256f
C222 outputibias.n31 gnd 0.005781f
C223 outputibias.n32 gnd 0.001372f
C224 outputibias.n33 gnd 9.76e-19
C225 outputibias.n34 gnd 5.24e-19
C226 outputibias.n35 gnd 0.001239f
C227 outputibias.n36 gnd 5.55e-19
C228 outputibias.n37 gnd 9.76e-19
C229 outputibias.n38 gnd 5.24e-19
C230 outputibias.n39 gnd 0.001239f
C231 outputibias.n40 gnd 5.55e-19
C232 outputibias.n41 gnd 0.004176f
C233 outputibias.t7 gnd 0.00202f
C234 outputibias.n42 gnd 9.3e-19
C235 outputibias.n43 gnd 7.32e-19
C236 outputibias.n44 gnd 5.24e-19
C237 outputibias.n45 gnd 0.02322f
C238 outputibias.n46 gnd 9.76e-19
C239 outputibias.n47 gnd 5.24e-19
C240 outputibias.n48 gnd 5.55e-19
C241 outputibias.n49 gnd 0.001239f
C242 outputibias.n50 gnd 0.001239f
C243 outputibias.n51 gnd 5.55e-19
C244 outputibias.n52 gnd 5.24e-19
C245 outputibias.n53 gnd 9.76e-19
C246 outputibias.n54 gnd 9.76e-19
C247 outputibias.n55 gnd 5.24e-19
C248 outputibias.n56 gnd 5.55e-19
C249 outputibias.n57 gnd 0.001239f
C250 outputibias.n58 gnd 0.002683f
C251 outputibias.n59 gnd 5.55e-19
C252 outputibias.n60 gnd 5.24e-19
C253 outputibias.n61 gnd 0.002256f
C254 outputibias.n62 gnd 0.005197f
C255 outputibias.n63 gnd 0.121892f
C256 outputibias.n64 gnd 0.001372f
C257 outputibias.n65 gnd 9.76e-19
C258 outputibias.n66 gnd 5.24e-19
C259 outputibias.n67 gnd 0.001239f
C260 outputibias.n68 gnd 5.55e-19
C261 outputibias.n69 gnd 9.76e-19
C262 outputibias.n70 gnd 5.24e-19
C263 outputibias.n71 gnd 0.001239f
C264 outputibias.n72 gnd 5.55e-19
C265 outputibias.n73 gnd 0.004176f
C266 outputibias.t3 gnd 0.00202f
C267 outputibias.n74 gnd 9.3e-19
C268 outputibias.n75 gnd 7.32e-19
C269 outputibias.n76 gnd 5.24e-19
C270 outputibias.n77 gnd 0.02322f
C271 outputibias.n78 gnd 9.76e-19
C272 outputibias.n79 gnd 5.24e-19
C273 outputibias.n80 gnd 5.55e-19
C274 outputibias.n81 gnd 0.001239f
C275 outputibias.n82 gnd 0.001239f
C276 outputibias.n83 gnd 5.55e-19
C277 outputibias.n84 gnd 5.24e-19
C278 outputibias.n85 gnd 9.76e-19
C279 outputibias.n86 gnd 9.76e-19
C280 outputibias.n87 gnd 5.24e-19
C281 outputibias.n88 gnd 5.55e-19
C282 outputibias.n89 gnd 0.001239f
C283 outputibias.n90 gnd 0.002683f
C284 outputibias.n91 gnd 5.55e-19
C285 outputibias.n92 gnd 5.24e-19
C286 outputibias.n93 gnd 0.002256f
C287 outputibias.n94 gnd 0.005197f
C288 outputibias.n95 gnd 0.064513f
C289 outputibias.n96 gnd 0.001372f
C290 outputibias.n97 gnd 9.76e-19
C291 outputibias.n98 gnd 5.24e-19
C292 outputibias.n99 gnd 0.001239f
C293 outputibias.n100 gnd 5.55e-19
C294 outputibias.n101 gnd 9.76e-19
C295 outputibias.n102 gnd 5.24e-19
C296 outputibias.n103 gnd 0.001239f
C297 outputibias.n104 gnd 5.55e-19
C298 outputibias.n105 gnd 0.004176f
C299 outputibias.t1 gnd 0.00202f
C300 outputibias.n106 gnd 9.3e-19
C301 outputibias.n107 gnd 7.32e-19
C302 outputibias.n108 gnd 5.24e-19
C303 outputibias.n109 gnd 0.02322f
C304 outputibias.n110 gnd 9.76e-19
C305 outputibias.n111 gnd 5.24e-19
C306 outputibias.n112 gnd 5.55e-19
C307 outputibias.n113 gnd 0.001239f
C308 outputibias.n114 gnd 0.001239f
C309 outputibias.n115 gnd 5.55e-19
C310 outputibias.n116 gnd 5.24e-19
C311 outputibias.n117 gnd 9.76e-19
C312 outputibias.n118 gnd 9.76e-19
C313 outputibias.n119 gnd 5.24e-19
C314 outputibias.n120 gnd 5.55e-19
C315 outputibias.n121 gnd 0.001239f
C316 outputibias.n122 gnd 0.002683f
C317 outputibias.n123 gnd 5.55e-19
C318 outputibias.n124 gnd 5.24e-19
C319 outputibias.n125 gnd 0.002256f
C320 outputibias.n126 gnd 0.005197f
C321 outputibias.n127 gnd 0.084814f
C322 outputibias.t0 gnd 0.108319f
C323 outputibias.t2 gnd 0.108319f
C324 outputibias.t6 gnd 0.108319f
C325 outputibias.t4 gnd 0.109238f
C326 outputibias.n128 gnd 0.134674f
C327 outputibias.n129 gnd 0.07244f
C328 outputibias.n130 gnd 0.079818f
C329 outputibias.n131 gnd 0.164901f
C330 outputibias.t10 gnd 0.11477f
C331 outputibias.n132 gnd 0.067481f
C332 outputibias.t8 gnd 0.11477f
C333 outputibias.n133 gnd 0.065115f
C334 outputibias.n134 gnd 0.029159f
C335 a_n2982_8322.t15 gnd 0.100128f
C336 a_n2982_8322.t35 gnd 20.7724f
C337 a_n2982_8322.t34 gnd 20.6268f
C338 a_n2982_8322.t37 gnd 20.6268f
C339 a_n2982_8322.t36 gnd 20.7724f
C340 a_n2982_8322.t33 gnd 20.6268f
C341 a_n2982_8322.t32 gnd 30.221401f
C342 a_n2982_8322.t14 gnd 0.937544f
C343 a_n2982_8322.t27 gnd 0.100128f
C344 a_n2982_8322.t23 gnd 0.100128f
C345 a_n2982_8322.n0 gnd 0.705299f
C346 a_n2982_8322.n1 gnd 0.788068f
C347 a_n2982_8322.t30 gnd 0.100128f
C348 a_n2982_8322.t20 gnd 0.100128f
C349 a_n2982_8322.n2 gnd 0.705299f
C350 a_n2982_8322.n3 gnd 0.400407f
C351 a_n2982_8322.t11 gnd 0.100128f
C352 a_n2982_8322.t10 gnd 0.100128f
C353 a_n2982_8322.n4 gnd 0.705299f
C354 a_n2982_8322.n5 gnd 0.400407f
C355 a_n2982_8322.t24 gnd 0.100128f
C356 a_n2982_8322.t17 gnd 0.100128f
C357 a_n2982_8322.n6 gnd 0.705299f
C358 a_n2982_8322.n7 gnd 0.400407f
C359 a_n2982_8322.t21 gnd 0.100128f
C360 a_n2982_8322.t19 gnd 0.100128f
C361 a_n2982_8322.n8 gnd 0.705299f
C362 a_n2982_8322.n9 gnd 0.400407f
C363 a_n2982_8322.t8 gnd 0.935678f
C364 a_n2982_8322.n10 gnd 1.87079f
C365 a_n2982_8322.t3 gnd 0.937544f
C366 a_n2982_8322.t7 gnd 0.100128f
C367 a_n2982_8322.t6 gnd 0.100128f
C368 a_n2982_8322.n11 gnd 0.705299f
C369 a_n2982_8322.n12 gnd 0.788068f
C370 a_n2982_8322.t1 gnd 0.935678f
C371 a_n2982_8322.n13 gnd 0.396567f
C372 a_n2982_8322.t4 gnd 0.935678f
C373 a_n2982_8322.n14 gnd 0.396567f
C374 a_n2982_8322.t2 gnd 0.100128f
C375 a_n2982_8322.t0 gnd 0.100128f
C376 a_n2982_8322.n15 gnd 0.705299f
C377 a_n2982_8322.n16 gnd 0.400407f
C378 a_n2982_8322.t5 gnd 0.935678f
C379 a_n2982_8322.n17 gnd 1.47094f
C380 a_n2982_8322.n18 gnd 2.35059f
C381 a_n2982_8322.n19 gnd 3.83141f
C382 a_n2982_8322.t9 gnd 0.935678f
C383 a_n2982_8322.n20 gnd 1.11111f
C384 a_n2982_8322.t26 gnd 0.100128f
C385 a_n2982_8322.t25 gnd 0.100128f
C386 a_n2982_8322.n21 gnd 0.705299f
C387 a_n2982_8322.n22 gnd 0.400407f
C388 a_n2982_8322.t13 gnd 0.100128f
C389 a_n2982_8322.t12 gnd 0.100128f
C390 a_n2982_8322.n23 gnd 0.705299f
C391 a_n2982_8322.n24 gnd 0.400407f
C392 a_n2982_8322.t28 gnd 0.100128f
C393 a_n2982_8322.t16 gnd 0.100128f
C394 a_n2982_8322.n25 gnd 0.705299f
C395 a_n2982_8322.n26 gnd 0.400407f
C396 a_n2982_8322.t29 gnd 0.937542f
C397 a_n2982_8322.t22 gnd 0.100128f
C398 a_n2982_8322.t18 gnd 0.100128f
C399 a_n2982_8322.n27 gnd 0.705299f
C400 a_n2982_8322.n28 gnd 0.78807f
C401 a_n2982_8322.n29 gnd 0.400405f
C402 a_n2982_8322.n30 gnd 0.705301f
C403 a_n2982_8322.t31 gnd 0.100128f
C404 diffpairibias.t27 gnd 0.090128f
C405 diffpairibias.t23 gnd 0.08996f
C406 diffpairibias.n0 gnd 0.105991f
C407 diffpairibias.t28 gnd 0.08996f
C408 diffpairibias.n1 gnd 0.051736f
C409 diffpairibias.t25 gnd 0.08996f
C410 diffpairibias.n2 gnd 0.051736f
C411 diffpairibias.t29 gnd 0.08996f
C412 diffpairibias.n3 gnd 0.041084f
C413 diffpairibias.t15 gnd 0.086371f
C414 diffpairibias.t1 gnd 0.085993f
C415 diffpairibias.n4 gnd 0.13579f
C416 diffpairibias.t11 gnd 0.085993f
C417 diffpairibias.n5 gnd 0.072463f
C418 diffpairibias.t13 gnd 0.085993f
C419 diffpairibias.n6 gnd 0.072463f
C420 diffpairibias.t7 gnd 0.085993f
C421 diffpairibias.n7 gnd 0.072463f
C422 diffpairibias.t3 gnd 0.085993f
C423 diffpairibias.n8 gnd 0.072463f
C424 diffpairibias.t17 gnd 0.085993f
C425 diffpairibias.n9 gnd 0.072463f
C426 diffpairibias.t5 gnd 0.085993f
C427 diffpairibias.n10 gnd 0.072463f
C428 diffpairibias.t19 gnd 0.085993f
C429 diffpairibias.n11 gnd 0.072463f
C430 diffpairibias.t9 gnd 0.085993f
C431 diffpairibias.n12 gnd 0.102883f
C432 diffpairibias.t14 gnd 0.086899f
C433 diffpairibias.t0 gnd 0.086748f
C434 diffpairibias.n13 gnd 0.094648f
C435 diffpairibias.t10 gnd 0.086748f
C436 diffpairibias.n14 gnd 0.052262f
C437 diffpairibias.t12 gnd 0.086748f
C438 diffpairibias.n15 gnd 0.052262f
C439 diffpairibias.t6 gnd 0.086748f
C440 diffpairibias.n16 gnd 0.052262f
C441 diffpairibias.t2 gnd 0.086748f
C442 diffpairibias.n17 gnd 0.052262f
C443 diffpairibias.t16 gnd 0.086748f
C444 diffpairibias.n18 gnd 0.052262f
C445 diffpairibias.t4 gnd 0.086748f
C446 diffpairibias.n19 gnd 0.052262f
C447 diffpairibias.t18 gnd 0.086748f
C448 diffpairibias.n20 gnd 0.052262f
C449 diffpairibias.t8 gnd 0.086748f
C450 diffpairibias.n21 gnd 0.061849f
C451 diffpairibias.n22 gnd 0.233513f
C452 diffpairibias.t20 gnd 0.08996f
C453 diffpairibias.n23 gnd 0.051747f
C454 diffpairibias.t26 gnd 0.08996f
C455 diffpairibias.n24 gnd 0.051736f
C456 diffpairibias.t22 gnd 0.08996f
C457 diffpairibias.n25 gnd 0.051736f
C458 diffpairibias.t21 gnd 0.08996f
C459 diffpairibias.n26 gnd 0.051736f
C460 diffpairibias.t24 gnd 0.08996f
C461 diffpairibias.n27 gnd 0.04729f
C462 diffpairibias.n28 gnd 0.047711f
C463 minus.n0 gnd 0.031253f
C464 minus.n1 gnd 0.007092f
C465 minus.n2 gnd 0.031253f
C466 minus.n3 gnd 0.007092f
C467 minus.n4 gnd 0.031253f
C468 minus.n5 gnd 0.007092f
C469 minus.n6 gnd 0.031253f
C470 minus.n7 gnd 0.007092f
C471 minus.n8 gnd 0.031253f
C472 minus.n9 gnd 0.007092f
C473 minus.t8 gnd 0.458091f
C474 minus.t7 gnd 0.442045f
C475 minus.n10 gnd 0.202766f
C476 minus.n11 gnd 0.181989f
C477 minus.n12 gnd 0.134546f
C478 minus.n13 gnd 0.031253f
C479 minus.t11 gnd 0.442045f
C480 minus.n14 gnd 0.196371f
C481 minus.n15 gnd 0.007092f
C482 minus.t10 gnd 0.442045f
C483 minus.n16 gnd 0.196371f
C484 minus.n17 gnd 0.031253f
C485 minus.n18 gnd 0.031253f
C486 minus.n19 gnd 0.031253f
C487 minus.t12 gnd 0.442045f
C488 minus.n20 gnd 0.196371f
C489 minus.n21 gnd 0.007092f
C490 minus.t20 gnd 0.442045f
C491 minus.n22 gnd 0.196371f
C492 minus.n23 gnd 0.031253f
C493 minus.n24 gnd 0.031253f
C494 minus.n25 gnd 0.031253f
C495 minus.t18 gnd 0.442045f
C496 minus.n26 gnd 0.196371f
C497 minus.n27 gnd 0.007092f
C498 minus.t25 gnd 0.442045f
C499 minus.n28 gnd 0.196371f
C500 minus.n29 gnd 0.031253f
C501 minus.n30 gnd 0.031253f
C502 minus.n31 gnd 0.031253f
C503 minus.t24 gnd 0.442045f
C504 minus.n32 gnd 0.196371f
C505 minus.n33 gnd 0.007092f
C506 minus.t14 gnd 0.442045f
C507 minus.n34 gnd 0.196371f
C508 minus.n35 gnd 0.031253f
C509 minus.n36 gnd 0.031253f
C510 minus.n37 gnd 0.031253f
C511 minus.t22 gnd 0.442045f
C512 minus.n38 gnd 0.196371f
C513 minus.n39 gnd 0.007092f
C514 minus.t19 gnd 0.442045f
C515 minus.n40 gnd 0.19666f
C516 minus.n41 gnd 0.361941f
C517 minus.n42 gnd 0.031253f
C518 minus.t13 gnd 0.442045f
C519 minus.t15 gnd 0.442045f
C520 minus.n43 gnd 0.031253f
C521 minus.t5 gnd 0.442045f
C522 minus.n44 gnd 0.196371f
C523 minus.n45 gnd 0.031253f
C524 minus.t6 gnd 0.442045f
C525 minus.t26 gnd 0.442045f
C526 minus.n46 gnd 0.196371f
C527 minus.n47 gnd 0.031253f
C528 minus.t21 gnd 0.442045f
C529 minus.t23 gnd 0.442045f
C530 minus.n48 gnd 0.196371f
C531 minus.n49 gnd 0.031253f
C532 minus.t16 gnd 0.442045f
C533 minus.t17 gnd 0.442045f
C534 minus.n50 gnd 0.196371f
C535 minus.n51 gnd 0.031253f
C536 minus.t9 gnd 0.442045f
C537 minus.t27 gnd 0.442045f
C538 minus.n52 gnd 0.202766f
C539 minus.t28 gnd 0.458091f
C540 minus.n53 gnd 0.181989f
C541 minus.n54 gnd 0.134546f
C542 minus.n55 gnd 0.007092f
C543 minus.n56 gnd 0.196371f
C544 minus.n57 gnd 0.007092f
C545 minus.n58 gnd 0.031253f
C546 minus.n59 gnd 0.031253f
C547 minus.n60 gnd 0.031253f
C548 minus.n61 gnd 0.007092f
C549 minus.n62 gnd 0.196371f
C550 minus.n63 gnd 0.007092f
C551 minus.n64 gnd 0.031253f
C552 minus.n65 gnd 0.031253f
C553 minus.n66 gnd 0.031253f
C554 minus.n67 gnd 0.007092f
C555 minus.n68 gnd 0.196371f
C556 minus.n69 gnd 0.007092f
C557 minus.n70 gnd 0.031253f
C558 minus.n71 gnd 0.031253f
C559 minus.n72 gnd 0.031253f
C560 minus.n73 gnd 0.007092f
C561 minus.n74 gnd 0.196371f
C562 minus.n75 gnd 0.007092f
C563 minus.n76 gnd 0.031253f
C564 minus.n77 gnd 0.031253f
C565 minus.n78 gnd 0.031253f
C566 minus.n79 gnd 0.007092f
C567 minus.n80 gnd 0.196371f
C568 minus.n81 gnd 0.007092f
C569 minus.n82 gnd 0.19666f
C570 minus.n83 gnd 1.04701f
C571 minus.n84 gnd 1.56003f
C572 minus.t1 gnd 0.009634f
C573 minus.t0 gnd 0.009634f
C574 minus.n85 gnd 0.03168f
C575 minus.t4 gnd 0.009634f
C576 minus.t3 gnd 0.009634f
C577 minus.n86 gnd 0.031246f
C578 minus.n87 gnd 0.266671f
C579 minus.t2 gnd 0.053624f
C580 minus.n88 gnd 0.14552f
C581 minus.n89 gnd 2.31716f
C582 CSoutput.n0 gnd 0.038243f
C583 CSoutput.t173 gnd 0.252966f
C584 CSoutput.n1 gnd 0.114227f
C585 CSoutput.n2 gnd 0.038243f
C586 CSoutput.t180 gnd 0.252966f
C587 CSoutput.n3 gnd 0.03031f
C588 CSoutput.n4 gnd 0.038243f
C589 CSoutput.t189 gnd 0.252966f
C590 CSoutput.n5 gnd 0.026137f
C591 CSoutput.n6 gnd 0.038243f
C592 CSoutput.t178 gnd 0.252966f
C593 CSoutput.t175 gnd 0.252966f
C594 CSoutput.n7 gnd 0.112982f
C595 CSoutput.n8 gnd 0.038243f
C596 CSoutput.t187 gnd 0.252966f
C597 CSoutput.n9 gnd 0.02492f
C598 CSoutput.n10 gnd 0.038243f
C599 CSoutput.t168 gnd 0.252966f
C600 CSoutput.t171 gnd 0.252966f
C601 CSoutput.n11 gnd 0.112982f
C602 CSoutput.n12 gnd 0.038243f
C603 CSoutput.t184 gnd 0.252966f
C604 CSoutput.n13 gnd 0.026137f
C605 CSoutput.n14 gnd 0.038243f
C606 CSoutput.t183 gnd 0.252966f
C607 CSoutput.t169 gnd 0.252966f
C608 CSoutput.n15 gnd 0.112982f
C609 CSoutput.n16 gnd 0.038243f
C610 CSoutput.t174 gnd 0.252966f
C611 CSoutput.n17 gnd 0.027915f
C612 CSoutput.t185 gnd 0.302301f
C613 CSoutput.t181 gnd 0.252966f
C614 CSoutput.n18 gnd 0.144234f
C615 CSoutput.n19 gnd 0.139957f
C616 CSoutput.n20 gnd 0.162367f
C617 CSoutput.n21 gnd 0.038243f
C618 CSoutput.n22 gnd 0.031918f
C619 CSoutput.n23 gnd 0.112982f
C620 CSoutput.n24 gnd 0.030768f
C621 CSoutput.n25 gnd 0.03031f
C622 CSoutput.n26 gnd 0.038243f
C623 CSoutput.n27 gnd 0.038243f
C624 CSoutput.n28 gnd 0.031672f
C625 CSoutput.n29 gnd 0.026891f
C626 CSoutput.n30 gnd 0.115497f
C627 CSoutput.n31 gnd 0.027261f
C628 CSoutput.n32 gnd 0.038243f
C629 CSoutput.n33 gnd 0.038243f
C630 CSoutput.n34 gnd 0.038243f
C631 CSoutput.n35 gnd 0.031335f
C632 CSoutput.n36 gnd 0.112982f
C633 CSoutput.n37 gnd 0.029967f
C634 CSoutput.n38 gnd 0.031111f
C635 CSoutput.n39 gnd 0.038243f
C636 CSoutput.n40 gnd 0.038243f
C637 CSoutput.n41 gnd 0.031911f
C638 CSoutput.n42 gnd 0.029167f
C639 CSoutput.n43 gnd 0.112982f
C640 CSoutput.n44 gnd 0.029906f
C641 CSoutput.n45 gnd 0.038243f
C642 CSoutput.n46 gnd 0.038243f
C643 CSoutput.n47 gnd 0.038243f
C644 CSoutput.n48 gnd 0.029906f
C645 CSoutput.n49 gnd 0.112982f
C646 CSoutput.n50 gnd 0.029167f
C647 CSoutput.n51 gnd 0.031911f
C648 CSoutput.n52 gnd 0.038243f
C649 CSoutput.n53 gnd 0.038243f
C650 CSoutput.n54 gnd 0.031111f
C651 CSoutput.n55 gnd 0.029967f
C652 CSoutput.n56 gnd 0.112982f
C653 CSoutput.n57 gnd 0.031335f
C654 CSoutput.n58 gnd 0.038243f
C655 CSoutput.n59 gnd 0.038243f
C656 CSoutput.n60 gnd 0.038243f
C657 CSoutput.n61 gnd 0.027261f
C658 CSoutput.n62 gnd 0.115497f
C659 CSoutput.n63 gnd 0.026891f
C660 CSoutput.t179 gnd 0.252966f
C661 CSoutput.n64 gnd 0.112982f
C662 CSoutput.n65 gnd 0.031672f
C663 CSoutput.n66 gnd 0.038243f
C664 CSoutput.n67 gnd 0.038243f
C665 CSoutput.n68 gnd 0.038243f
C666 CSoutput.n69 gnd 0.030768f
C667 CSoutput.n70 gnd 0.112982f
C668 CSoutput.n71 gnd 0.031918f
C669 CSoutput.n72 gnd 0.027915f
C670 CSoutput.n73 gnd 0.038243f
C671 CSoutput.n74 gnd 0.038243f
C672 CSoutput.n75 gnd 0.02895f
C673 CSoutput.n76 gnd 0.017194f
C674 CSoutput.t188 gnd 0.284226f
C675 CSoutput.n77 gnd 0.141192f
C676 CSoutput.n78 gnd 0.577609f
C677 CSoutput.t167 gnd 0.047702f
C678 CSoutput.t143 gnd 0.047702f
C679 CSoutput.n79 gnd 0.369326f
C680 CSoutput.t126 gnd 0.047702f
C681 CSoutput.t161 gnd 0.047702f
C682 CSoutput.n80 gnd 0.368668f
C683 CSoutput.n81 gnd 0.374197f
C684 CSoutput.t133 gnd 0.047702f
C685 CSoutput.t153 gnd 0.047702f
C686 CSoutput.n82 gnd 0.368668f
C687 CSoutput.n83 gnd 0.184389f
C688 CSoutput.t140 gnd 0.047702f
C689 CSoutput.t147 gnd 0.047702f
C690 CSoutput.n84 gnd 0.368668f
C691 CSoutput.n85 gnd 0.338126f
C692 CSoutput.t145 gnd 0.047702f
C693 CSoutput.t134 gnd 0.047702f
C694 CSoutput.n86 gnd 0.369326f
C695 CSoutput.t122 gnd 0.047702f
C696 CSoutput.t146 gnd 0.047702f
C697 CSoutput.n87 gnd 0.368668f
C698 CSoutput.n88 gnd 0.374197f
C699 CSoutput.t144 gnd 0.047702f
C700 CSoutput.t132 gnd 0.047702f
C701 CSoutput.n89 gnd 0.368668f
C702 CSoutput.n90 gnd 0.184389f
C703 CSoutput.t121 gnd 0.047702f
C704 CSoutput.t120 gnd 0.047702f
C705 CSoutput.n91 gnd 0.368668f
C706 CSoutput.n92 gnd 0.27497f
C707 CSoutput.n93 gnd 0.346735f
C708 CSoutput.t150 gnd 0.047702f
C709 CSoutput.t138 gnd 0.047702f
C710 CSoutput.n94 gnd 0.369326f
C711 CSoutput.t129 gnd 0.047702f
C712 CSoutput.t151 gnd 0.047702f
C713 CSoutput.n95 gnd 0.368668f
C714 CSoutput.n96 gnd 0.374197f
C715 CSoutput.t149 gnd 0.047702f
C716 CSoutput.t137 gnd 0.047702f
C717 CSoutput.n97 gnd 0.368668f
C718 CSoutput.n98 gnd 0.184389f
C719 CSoutput.t128 gnd 0.047702f
C720 CSoutput.t127 gnd 0.047702f
C721 CSoutput.n99 gnd 0.368668f
C722 CSoutput.n100 gnd 0.27497f
C723 CSoutput.n101 gnd 0.387561f
C724 CSoutput.n102 gnd 8.072221f
C725 CSoutput.n104 gnd 0.676504f
C726 CSoutput.n105 gnd 0.507378f
C727 CSoutput.n106 gnd 0.676504f
C728 CSoutput.n107 gnd 0.676504f
C729 CSoutput.n108 gnd 1.82136f
C730 CSoutput.n109 gnd 0.676504f
C731 CSoutput.n110 gnd 0.676504f
C732 CSoutput.t177 gnd 0.84563f
C733 CSoutput.n111 gnd 0.676504f
C734 CSoutput.n112 gnd 0.676504f
C735 CSoutput.n116 gnd 0.676504f
C736 CSoutput.n120 gnd 0.676504f
C737 CSoutput.n121 gnd 0.676504f
C738 CSoutput.n123 gnd 0.676504f
C739 CSoutput.n128 gnd 0.676504f
C740 CSoutput.n130 gnd 0.676504f
C741 CSoutput.n131 gnd 0.676504f
C742 CSoutput.n133 gnd 0.676504f
C743 CSoutput.n134 gnd 0.676504f
C744 CSoutput.n136 gnd 0.676504f
C745 CSoutput.t170 gnd 11.3043f
C746 CSoutput.n138 gnd 0.676504f
C747 CSoutput.n139 gnd 0.507378f
C748 CSoutput.n140 gnd 0.676504f
C749 CSoutput.n141 gnd 0.676504f
C750 CSoutput.n142 gnd 1.82136f
C751 CSoutput.n143 gnd 0.676504f
C752 CSoutput.n144 gnd 0.676504f
C753 CSoutput.t172 gnd 0.84563f
C754 CSoutput.n145 gnd 0.676504f
C755 CSoutput.n146 gnd 0.676504f
C756 CSoutput.n150 gnd 0.676504f
C757 CSoutput.n154 gnd 0.676504f
C758 CSoutput.n155 gnd 0.676504f
C759 CSoutput.n157 gnd 0.676504f
C760 CSoutput.n162 gnd 0.676504f
C761 CSoutput.n164 gnd 0.676504f
C762 CSoutput.n165 gnd 0.676504f
C763 CSoutput.n167 gnd 0.676504f
C764 CSoutput.n168 gnd 0.676504f
C765 CSoutput.n170 gnd 0.676504f
C766 CSoutput.n171 gnd 0.507378f
C767 CSoutput.n173 gnd 0.676504f
C768 CSoutput.n174 gnd 0.507378f
C769 CSoutput.n175 gnd 0.676504f
C770 CSoutput.n176 gnd 0.676504f
C771 CSoutput.n177 gnd 1.82136f
C772 CSoutput.n178 gnd 0.676504f
C773 CSoutput.n179 gnd 0.676504f
C774 CSoutput.t176 gnd 0.84563f
C775 CSoutput.n180 gnd 0.676504f
C776 CSoutput.n181 gnd 1.82136f
C777 CSoutput.n183 gnd 0.676504f
C778 CSoutput.n184 gnd 0.676504f
C779 CSoutput.n186 gnd 0.676504f
C780 CSoutput.n187 gnd 0.676504f
C781 CSoutput.t186 gnd 11.120099f
C782 CSoutput.t182 gnd 11.3043f
C783 CSoutput.n193 gnd 2.12229f
C784 CSoutput.n194 gnd 8.645451f
C785 CSoutput.n195 gnd 9.007211f
C786 CSoutput.n200 gnd 2.29901f
C787 CSoutput.n206 gnd 0.676504f
C788 CSoutput.n208 gnd 0.676504f
C789 CSoutput.n210 gnd 0.676504f
C790 CSoutput.n212 gnd 0.676504f
C791 CSoutput.n214 gnd 0.676504f
C792 CSoutput.n220 gnd 0.676504f
C793 CSoutput.n227 gnd 1.24112f
C794 CSoutput.n228 gnd 1.24112f
C795 CSoutput.n229 gnd 0.676504f
C796 CSoutput.n230 gnd 0.676504f
C797 CSoutput.n232 gnd 0.507378f
C798 CSoutput.n233 gnd 0.434524f
C799 CSoutput.n235 gnd 0.507378f
C800 CSoutput.n236 gnd 0.434524f
C801 CSoutput.n237 gnd 0.507378f
C802 CSoutput.n239 gnd 0.676504f
C803 CSoutput.n241 gnd 1.82136f
C804 CSoutput.n242 gnd 2.12229f
C805 CSoutput.n243 gnd 7.95158f
C806 CSoutput.n245 gnd 0.507378f
C807 CSoutput.n246 gnd 1.30551f
C808 CSoutput.n247 gnd 0.507378f
C809 CSoutput.n249 gnd 0.676504f
C810 CSoutput.n251 gnd 1.82136f
C811 CSoutput.n252 gnd 3.96721f
C812 CSoutput.t142 gnd 0.047702f
C813 CSoutput.t136 gnd 0.047702f
C814 CSoutput.n253 gnd 0.369326f
C815 CSoutput.t160 gnd 0.047702f
C816 CSoutput.t125 gnd 0.047702f
C817 CSoutput.n254 gnd 0.368668f
C818 CSoutput.n255 gnd 0.374197f
C819 CSoutput.t152 gnd 0.047702f
C820 CSoutput.t130 gnd 0.047702f
C821 CSoutput.n256 gnd 0.368668f
C822 CSoutput.n257 gnd 0.184389f
C823 CSoutput.t156 gnd 0.047702f
C824 CSoutput.t139 gnd 0.047702f
C825 CSoutput.n258 gnd 0.368668f
C826 CSoutput.n259 gnd 0.338126f
C827 CSoutput.t162 gnd 0.047702f
C828 CSoutput.t163 gnd 0.047702f
C829 CSoutput.n260 gnd 0.369326f
C830 CSoutput.t124 gnd 0.047702f
C831 CSoutput.t155 gnd 0.047702f
C832 CSoutput.n261 gnd 0.368668f
C833 CSoutput.n262 gnd 0.374197f
C834 CSoutput.t159 gnd 0.047702f
C835 CSoutput.t123 gnd 0.047702f
C836 CSoutput.n263 gnd 0.368668f
C837 CSoutput.n264 gnd 0.184389f
C838 CSoutput.t141 gnd 0.047702f
C839 CSoutput.t154 gnd 0.047702f
C840 CSoutput.n265 gnd 0.368668f
C841 CSoutput.n266 gnd 0.27497f
C842 CSoutput.n267 gnd 0.346735f
C843 CSoutput.t165 gnd 0.047702f
C844 CSoutput.t166 gnd 0.047702f
C845 CSoutput.n268 gnd 0.369326f
C846 CSoutput.t135 gnd 0.047702f
C847 CSoutput.t158 gnd 0.047702f
C848 CSoutput.n269 gnd 0.368668f
C849 CSoutput.n270 gnd 0.374197f
C850 CSoutput.t164 gnd 0.047702f
C851 CSoutput.t131 gnd 0.047702f
C852 CSoutput.n271 gnd 0.368668f
C853 CSoutput.n272 gnd 0.184389f
C854 CSoutput.t148 gnd 0.047702f
C855 CSoutput.t157 gnd 0.047702f
C856 CSoutput.n273 gnd 0.368666f
C857 CSoutput.n274 gnd 0.274971f
C858 CSoutput.n275 gnd 0.387561f
C859 CSoutput.n276 gnd 11.1098f
C860 CSoutput.t95 gnd 0.041739f
C861 CSoutput.t18 gnd 0.041739f
C862 CSoutput.n277 gnd 0.370059f
C863 CSoutput.t75 gnd 0.041739f
C864 CSoutput.t2 gnd 0.041739f
C865 CSoutput.n278 gnd 0.368824f
C866 CSoutput.n279 gnd 0.343675f
C867 CSoutput.t57 gnd 0.041739f
C868 CSoutput.t98 gnd 0.041739f
C869 CSoutput.n280 gnd 0.368824f
C870 CSoutput.n281 gnd 0.169416f
C871 CSoutput.t43 gnd 0.041739f
C872 CSoutput.t56 gnd 0.041739f
C873 CSoutput.n282 gnd 0.368824f
C874 CSoutput.n283 gnd 0.169416f
C875 CSoutput.t6 gnd 0.041739f
C876 CSoutput.t63 gnd 0.041739f
C877 CSoutput.n284 gnd 0.368824f
C878 CSoutput.n285 gnd 0.169416f
C879 CSoutput.t80 gnd 0.041739f
C880 CSoutput.t44 gnd 0.041739f
C881 CSoutput.n286 gnd 0.368824f
C882 CSoutput.n287 gnd 0.169416f
C883 CSoutput.t59 gnd 0.041739f
C884 CSoutput.t90 gnd 0.041739f
C885 CSoutput.n288 gnd 0.368824f
C886 CSoutput.n289 gnd 0.169416f
C887 CSoutput.t17 gnd 0.041739f
C888 CSoutput.t33 gnd 0.041739f
C889 CSoutput.n290 gnd 0.368824f
C890 CSoutput.n291 gnd 0.169416f
C891 CSoutput.t76 gnd 0.041739f
C892 CSoutput.t115 gnd 0.041739f
C893 CSoutput.n292 gnd 0.368824f
C894 CSoutput.n293 gnd 0.169416f
C895 CSoutput.t68 gnd 0.041739f
C896 CSoutput.t99 gnd 0.041739f
C897 CSoutput.n294 gnd 0.368824f
C898 CSoutput.n295 gnd 0.312478f
C899 CSoutput.t54 gnd 0.041739f
C900 CSoutput.t27 gnd 0.041739f
C901 CSoutput.n296 gnd 0.370059f
C902 CSoutput.t39 gnd 0.041739f
C903 CSoutput.t53 gnd 0.041739f
C904 CSoutput.n297 gnd 0.368824f
C905 CSoutput.n298 gnd 0.343675f
C906 CSoutput.t26 gnd 0.041739f
C907 CSoutput.t41 gnd 0.041739f
C908 CSoutput.n299 gnd 0.368824f
C909 CSoutput.n300 gnd 0.169416f
C910 CSoutput.t55 gnd 0.041739f
C911 CSoutput.t25 gnd 0.041739f
C912 CSoutput.n301 gnd 0.368824f
C913 CSoutput.n302 gnd 0.169416f
C914 CSoutput.t40 gnd 0.041739f
C915 CSoutput.t14 gnd 0.041739f
C916 CSoutput.n303 gnd 0.368824f
C917 CSoutput.n304 gnd 0.169416f
C918 CSoutput.t24 gnd 0.041739f
C919 CSoutput.t42 gnd 0.041739f
C920 CSoutput.n305 gnd 0.368824f
C921 CSoutput.n306 gnd 0.169416f
C922 CSoutput.t9 gnd 0.041739f
C923 CSoutput.t108 gnd 0.041739f
C924 CSoutput.n307 gnd 0.368824f
C925 CSoutput.n308 gnd 0.169416f
C926 CSoutput.t30 gnd 0.041739f
C927 CSoutput.t117 gnd 0.041739f
C928 CSoutput.n309 gnd 0.368824f
C929 CSoutput.n310 gnd 0.169416f
C930 CSoutput.t104 gnd 0.041739f
C931 CSoutput.t109 gnd 0.041739f
C932 CSoutput.n311 gnd 0.368824f
C933 CSoutput.n312 gnd 0.169416f
C934 CSoutput.t119 gnd 0.041739f
C935 CSoutput.t105 gnd 0.041739f
C936 CSoutput.n313 gnd 0.368824f
C937 CSoutput.n314 gnd 0.257209f
C938 CSoutput.n315 gnd 0.324421f
C939 CSoutput.t16 gnd 0.041739f
C940 CSoutput.t110 gnd 0.041739f
C941 CSoutput.n316 gnd 0.370059f
C942 CSoutput.t92 gnd 0.041739f
C943 CSoutput.t31 gnd 0.041739f
C944 CSoutput.n317 gnd 0.368824f
C945 CSoutput.n318 gnd 0.343675f
C946 CSoutput.t0 gnd 0.041739f
C947 CSoutput.t101 gnd 0.041739f
C948 CSoutput.n319 gnd 0.368824f
C949 CSoutput.n320 gnd 0.169416f
C950 CSoutput.t49 gnd 0.041739f
C951 CSoutput.t58 gnd 0.041739f
C952 CSoutput.n321 gnd 0.368824f
C953 CSoutput.n322 gnd 0.169416f
C954 CSoutput.t111 gnd 0.041739f
C955 CSoutput.t91 gnd 0.041739f
C956 CSoutput.n323 gnd 0.368824f
C957 CSoutput.n324 gnd 0.169416f
C958 CSoutput.t69 gnd 0.041739f
C959 CSoutput.t1 gnd 0.041739f
C960 CSoutput.n325 gnd 0.368824f
C961 CSoutput.n326 gnd 0.169416f
C962 CSoutput.t13 gnd 0.041739f
C963 CSoutput.t107 gnd 0.041739f
C964 CSoutput.n327 gnd 0.368824f
C965 CSoutput.n328 gnd 0.169416f
C966 CSoutput.t22 gnd 0.041739f
C967 CSoutput.t29 gnd 0.041739f
C968 CSoutput.n329 gnd 0.368824f
C969 CSoutput.n330 gnd 0.169416f
C970 CSoutput.t118 gnd 0.041739f
C971 CSoutput.t100 gnd 0.041739f
C972 CSoutput.n331 gnd 0.368824f
C973 CSoutput.n332 gnd 0.169416f
C974 CSoutput.t48 gnd 0.041739f
C975 CSoutput.t15 gnd 0.041739f
C976 CSoutput.n333 gnd 0.368824f
C977 CSoutput.n334 gnd 0.257209f
C978 CSoutput.n335 gnd 0.348377f
C979 CSoutput.n336 gnd 11.808401f
C980 CSoutput.t65 gnd 0.041739f
C981 CSoutput.t8 gnd 0.041739f
C982 CSoutput.n337 gnd 0.370059f
C983 CSoutput.t47 gnd 0.041739f
C984 CSoutput.t102 gnd 0.041739f
C985 CSoutput.n338 gnd 0.368824f
C986 CSoutput.n339 gnd 0.343675f
C987 CSoutput.t12 gnd 0.041739f
C988 CSoutput.t82 gnd 0.041739f
C989 CSoutput.n340 gnd 0.368824f
C990 CSoutput.n341 gnd 0.169416f
C991 CSoutput.t81 gnd 0.041739f
C992 CSoutput.t67 gnd 0.041739f
C993 CSoutput.n342 gnd 0.368824f
C994 CSoutput.n343 gnd 0.169416f
C995 CSoutput.t85 gnd 0.041739f
C996 CSoutput.t50 gnd 0.041739f
C997 CSoutput.n344 gnd 0.368824f
C998 CSoutput.n345 gnd 0.169416f
C999 CSoutput.t77 gnd 0.041739f
C1000 CSoutput.t94 gnd 0.041739f
C1001 CSoutput.n346 gnd 0.368824f
C1002 CSoutput.n347 gnd 0.169416f
C1003 CSoutput.t116 gnd 0.041739f
C1004 CSoutput.t84 gnd 0.041739f
C1005 CSoutput.n348 gnd 0.368824f
C1006 CSoutput.n349 gnd 0.169416f
C1007 CSoutput.t89 gnd 0.041739f
C1008 CSoutput.t88 gnd 0.041739f
C1009 CSoutput.n350 gnd 0.368824f
C1010 CSoutput.n351 gnd 0.169416f
C1011 CSoutput.t72 gnd 0.041739f
C1012 CSoutput.t7 gnd 0.041739f
C1013 CSoutput.n352 gnd 0.368824f
C1014 CSoutput.n353 gnd 0.169416f
C1015 CSoutput.t46 gnd 0.041739f
C1016 CSoutput.t113 gnd 0.041739f
C1017 CSoutput.n354 gnd 0.368824f
C1018 CSoutput.n355 gnd 0.312478f
C1019 CSoutput.t51 gnd 0.041739f
C1020 CSoutput.t70 gnd 0.041739f
C1021 CSoutput.n356 gnd 0.370059f
C1022 CSoutput.t71 gnd 0.041739f
C1023 CSoutput.t60 gnd 0.041739f
C1024 CSoutput.n357 gnd 0.368824f
C1025 CSoutput.n358 gnd 0.343675f
C1026 CSoutput.t61 gnd 0.041739f
C1027 CSoutput.t52 gnd 0.041739f
C1028 CSoutput.n359 gnd 0.368824f
C1029 CSoutput.n360 gnd 0.169416f
C1030 CSoutput.t45 gnd 0.041739f
C1031 CSoutput.t37 gnd 0.041739f
C1032 CSoutput.n361 gnd 0.368824f
C1033 CSoutput.n362 gnd 0.169416f
C1034 CSoutput.t38 gnd 0.041739f
C1035 CSoutput.t62 gnd 0.041739f
C1036 CSoutput.n363 gnd 0.368824f
C1037 CSoutput.n364 gnd 0.169416f
C1038 CSoutput.t64 gnd 0.041739f
C1039 CSoutput.t4 gnd 0.041739f
C1040 CSoutput.n365 gnd 0.368824f
C1041 CSoutput.n366 gnd 0.169416f
C1042 CSoutput.t5 gnd 0.041739f
C1043 CSoutput.t28 gnd 0.041739f
C1044 CSoutput.n367 gnd 0.368824f
C1045 CSoutput.n368 gnd 0.169416f
C1046 CSoutput.t35 gnd 0.041739f
C1047 CSoutput.t23 gnd 0.041739f
C1048 CSoutput.n369 gnd 0.368824f
C1049 CSoutput.n370 gnd 0.169416f
C1050 CSoutput.t19 gnd 0.041739f
C1051 CSoutput.t10 gnd 0.041739f
C1052 CSoutput.n371 gnd 0.368824f
C1053 CSoutput.n372 gnd 0.169416f
C1054 CSoutput.t11 gnd 0.041739f
C1055 CSoutput.t36 gnd 0.041739f
C1056 CSoutput.n373 gnd 0.368824f
C1057 CSoutput.n374 gnd 0.257209f
C1058 CSoutput.n375 gnd 0.324421f
C1059 CSoutput.t86 gnd 0.041739f
C1060 CSoutput.t106 gnd 0.041739f
C1061 CSoutput.n376 gnd 0.370059f
C1062 CSoutput.t114 gnd 0.041739f
C1063 CSoutput.t74 gnd 0.041739f
C1064 CSoutput.n377 gnd 0.368824f
C1065 CSoutput.n378 gnd 0.343675f
C1066 CSoutput.t79 gnd 0.041739f
C1067 CSoutput.t96 gnd 0.041739f
C1068 CSoutput.n379 gnd 0.368824f
C1069 CSoutput.n380 gnd 0.169416f
C1070 CSoutput.t20 gnd 0.041739f
C1071 CSoutput.t66 gnd 0.041739f
C1072 CSoutput.n381 gnd 0.368824f
C1073 CSoutput.n382 gnd 0.169416f
C1074 CSoutput.t73 gnd 0.041739f
C1075 CSoutput.t87 gnd 0.041739f
C1076 CSoutput.n383 gnd 0.368824f
C1077 CSoutput.n384 gnd 0.169416f
C1078 CSoutput.t97 gnd 0.041739f
C1079 CSoutput.t78 gnd 0.041739f
C1080 CSoutput.n385 gnd 0.368824f
C1081 CSoutput.n386 gnd 0.169416f
C1082 CSoutput.t83 gnd 0.041739f
C1083 CSoutput.t103 gnd 0.041739f
C1084 CSoutput.n387 gnd 0.368824f
C1085 CSoutput.n388 gnd 0.169416f
C1086 CSoutput.t21 gnd 0.041739f
C1087 CSoutput.t32 gnd 0.041739f
C1088 CSoutput.n389 gnd 0.368824f
C1089 CSoutput.n390 gnd 0.169416f
C1090 CSoutput.t93 gnd 0.041739f
C1091 CSoutput.t112 gnd 0.041739f
C1092 CSoutput.n391 gnd 0.368824f
C1093 CSoutput.n392 gnd 0.169416f
C1094 CSoutput.t3 gnd 0.041739f
C1095 CSoutput.t34 gnd 0.041739f
C1096 CSoutput.n393 gnd 0.368824f
C1097 CSoutput.n394 gnd 0.257209f
C1098 CSoutput.n395 gnd 0.348377f
C1099 CSoutput.n396 gnd 7.15579f
C1100 CSoutput.n397 gnd 11.7809f
C1101 vdd.t51 gnd 0.029713f
C1102 vdd.t29 gnd 0.029713f
C1103 vdd.n0 gnd 0.234355f
C1104 vdd.t8 gnd 0.029713f
C1105 vdd.t47 gnd 0.029713f
C1106 vdd.n1 gnd 0.233968f
C1107 vdd.n2 gnd 0.215763f
C1108 vdd.t26 gnd 0.029713f
C1109 vdd.t56 gnd 0.029713f
C1110 vdd.n3 gnd 0.233968f
C1111 vdd.n4 gnd 0.10912f
C1112 vdd.t41 gnd 0.029713f
C1113 vdd.t34 gnd 0.029713f
C1114 vdd.n5 gnd 0.233968f
C1115 vdd.n6 gnd 0.102388f
C1116 vdd.t60 gnd 0.029713f
C1117 vdd.t24 gnd 0.029713f
C1118 vdd.n7 gnd 0.234355f
C1119 vdd.t32 gnd 0.029713f
C1120 vdd.t54 gnd 0.029713f
C1121 vdd.n8 gnd 0.233968f
C1122 vdd.n9 gnd 0.215763f
C1123 vdd.t43 gnd 0.029713f
C1124 vdd.t12 gnd 0.029713f
C1125 vdd.n10 gnd 0.233968f
C1126 vdd.n11 gnd 0.10912f
C1127 vdd.t21 gnd 0.029713f
C1128 vdd.t39 gnd 0.029713f
C1129 vdd.n12 gnd 0.233968f
C1130 vdd.n13 gnd 0.102388f
C1131 vdd.n14 gnd 0.072387f
C1132 vdd.t66 gnd 0.016507f
C1133 vdd.t145 gnd 0.016507f
C1134 vdd.n15 gnd 0.151944f
C1135 vdd.t147 gnd 0.016507f
C1136 vdd.t63 gnd 0.016507f
C1137 vdd.n16 gnd 0.1515f
C1138 vdd.n17 gnd 0.263657f
C1139 vdd.t146 gnd 0.016507f
C1140 vdd.t143 gnd 0.016507f
C1141 vdd.n18 gnd 0.1515f
C1142 vdd.n19 gnd 0.109078f
C1143 vdd.t2 gnd 0.016507f
C1144 vdd.t64 gnd 0.016507f
C1145 vdd.n20 gnd 0.151944f
C1146 vdd.t3 gnd 0.016507f
C1147 vdd.t62 gnd 0.016507f
C1148 vdd.n21 gnd 0.1515f
C1149 vdd.n22 gnd 0.263657f
C1150 vdd.t0 gnd 0.016507f
C1151 vdd.t1 gnd 0.016507f
C1152 vdd.n23 gnd 0.1515f
C1153 vdd.n24 gnd 0.109078f
C1154 vdd.t65 gnd 0.016507f
C1155 vdd.t61 gnd 0.016507f
C1156 vdd.n25 gnd 0.1515f
C1157 vdd.t144 gnd 0.016507f
C1158 vdd.t4 gnd 0.016507f
C1159 vdd.n26 gnd 0.1515f
C1160 vdd.n27 gnd 16.948801f
C1161 vdd.n28 gnd 6.76264f
C1162 vdd.n29 gnd 0.004502f
C1163 vdd.n30 gnd 0.004178f
C1164 vdd.n31 gnd 0.002311f
C1165 vdd.n32 gnd 0.005306f
C1166 vdd.n33 gnd 0.002245f
C1167 vdd.n34 gnd 0.002377f
C1168 vdd.n35 gnd 0.004178f
C1169 vdd.n36 gnd 0.002245f
C1170 vdd.n37 gnd 0.005306f
C1171 vdd.n38 gnd 0.002377f
C1172 vdd.n39 gnd 0.004178f
C1173 vdd.n40 gnd 0.002245f
C1174 vdd.n41 gnd 0.00398f
C1175 vdd.n42 gnd 0.003992f
C1176 vdd.t183 gnd 0.0114f
C1177 vdd.n43 gnd 0.025366f
C1178 vdd.n44 gnd 0.132009f
C1179 vdd.n45 gnd 0.002245f
C1180 vdd.n46 gnd 0.002377f
C1181 vdd.n47 gnd 0.005306f
C1182 vdd.n48 gnd 0.005306f
C1183 vdd.n49 gnd 0.002377f
C1184 vdd.n50 gnd 0.002245f
C1185 vdd.n51 gnd 0.004178f
C1186 vdd.n52 gnd 0.004178f
C1187 vdd.n53 gnd 0.002245f
C1188 vdd.n54 gnd 0.002377f
C1189 vdd.n55 gnd 0.005306f
C1190 vdd.n56 gnd 0.005306f
C1191 vdd.n57 gnd 0.002377f
C1192 vdd.n58 gnd 0.002245f
C1193 vdd.n59 gnd 0.004178f
C1194 vdd.n60 gnd 0.004178f
C1195 vdd.n61 gnd 0.002245f
C1196 vdd.n62 gnd 0.002377f
C1197 vdd.n63 gnd 0.005306f
C1198 vdd.n64 gnd 0.005306f
C1199 vdd.n65 gnd 0.012545f
C1200 vdd.n66 gnd 0.002311f
C1201 vdd.n67 gnd 0.002245f
C1202 vdd.n68 gnd 0.010799f
C1203 vdd.n69 gnd 0.007539f
C1204 vdd.t174 gnd 0.026412f
C1205 vdd.t204 gnd 0.026412f
C1206 vdd.n70 gnd 0.181521f
C1207 vdd.n71 gnd 0.142739f
C1208 vdd.t159 gnd 0.026412f
C1209 vdd.t196 gnd 0.026412f
C1210 vdd.n72 gnd 0.181521f
C1211 vdd.n73 gnd 0.115189f
C1212 vdd.t164 gnd 0.026412f
C1213 vdd.t200 gnd 0.026412f
C1214 vdd.n74 gnd 0.181521f
C1215 vdd.n75 gnd 0.115189f
C1216 vdd.n76 gnd 0.004502f
C1217 vdd.n77 gnd 0.004178f
C1218 vdd.n78 gnd 0.002311f
C1219 vdd.n79 gnd 0.005306f
C1220 vdd.n80 gnd 0.002245f
C1221 vdd.n81 gnd 0.002377f
C1222 vdd.n82 gnd 0.004178f
C1223 vdd.n83 gnd 0.002245f
C1224 vdd.n84 gnd 0.005306f
C1225 vdd.n85 gnd 0.002377f
C1226 vdd.n86 gnd 0.004178f
C1227 vdd.n87 gnd 0.002245f
C1228 vdd.n88 gnd 0.00398f
C1229 vdd.n89 gnd 0.003992f
C1230 vdd.t178 gnd 0.0114f
C1231 vdd.n90 gnd 0.025366f
C1232 vdd.n91 gnd 0.132009f
C1233 vdd.n92 gnd 0.002245f
C1234 vdd.n93 gnd 0.002377f
C1235 vdd.n94 gnd 0.005306f
C1236 vdd.n95 gnd 0.005306f
C1237 vdd.n96 gnd 0.002377f
C1238 vdd.n97 gnd 0.002245f
C1239 vdd.n98 gnd 0.004178f
C1240 vdd.n99 gnd 0.004178f
C1241 vdd.n100 gnd 0.002245f
C1242 vdd.n101 gnd 0.002377f
C1243 vdd.n102 gnd 0.005306f
C1244 vdd.n103 gnd 0.005306f
C1245 vdd.n104 gnd 0.002377f
C1246 vdd.n105 gnd 0.002245f
C1247 vdd.n106 gnd 0.004178f
C1248 vdd.n107 gnd 0.004178f
C1249 vdd.n108 gnd 0.002245f
C1250 vdd.n109 gnd 0.002377f
C1251 vdd.n110 gnd 0.005306f
C1252 vdd.n111 gnd 0.005306f
C1253 vdd.n112 gnd 0.012545f
C1254 vdd.n113 gnd 0.002311f
C1255 vdd.n114 gnd 0.002245f
C1256 vdd.n115 gnd 0.010799f
C1257 vdd.n116 gnd 0.007302f
C1258 vdd.n117 gnd 0.085702f
C1259 vdd.n118 gnd 0.004502f
C1260 vdd.n119 gnd 0.004178f
C1261 vdd.n120 gnd 0.002311f
C1262 vdd.n121 gnd 0.005306f
C1263 vdd.n122 gnd 0.002245f
C1264 vdd.n123 gnd 0.002377f
C1265 vdd.n124 gnd 0.004178f
C1266 vdd.n125 gnd 0.002245f
C1267 vdd.n126 gnd 0.005306f
C1268 vdd.n127 gnd 0.002377f
C1269 vdd.n128 gnd 0.004178f
C1270 vdd.n129 gnd 0.002245f
C1271 vdd.n130 gnd 0.00398f
C1272 vdd.n131 gnd 0.003992f
C1273 vdd.t206 gnd 0.0114f
C1274 vdd.n132 gnd 0.025366f
C1275 vdd.n133 gnd 0.132009f
C1276 vdd.n134 gnd 0.002245f
C1277 vdd.n135 gnd 0.002377f
C1278 vdd.n136 gnd 0.005306f
C1279 vdd.n137 gnd 0.005306f
C1280 vdd.n138 gnd 0.002377f
C1281 vdd.n139 gnd 0.002245f
C1282 vdd.n140 gnd 0.004178f
C1283 vdd.n141 gnd 0.004178f
C1284 vdd.n142 gnd 0.002245f
C1285 vdd.n143 gnd 0.002377f
C1286 vdd.n144 gnd 0.005306f
C1287 vdd.n145 gnd 0.005306f
C1288 vdd.n146 gnd 0.002377f
C1289 vdd.n147 gnd 0.002245f
C1290 vdd.n148 gnd 0.004178f
C1291 vdd.n149 gnd 0.004178f
C1292 vdd.n150 gnd 0.002245f
C1293 vdd.n151 gnd 0.002377f
C1294 vdd.n152 gnd 0.005306f
C1295 vdd.n153 gnd 0.005306f
C1296 vdd.n154 gnd 0.012545f
C1297 vdd.n155 gnd 0.002311f
C1298 vdd.n156 gnd 0.002245f
C1299 vdd.n157 gnd 0.010799f
C1300 vdd.n158 gnd 0.007539f
C1301 vdd.t207 gnd 0.026412f
C1302 vdd.t157 gnd 0.026412f
C1303 vdd.n159 gnd 0.181521f
C1304 vdd.n160 gnd 0.142739f
C1305 vdd.t199 gnd 0.026412f
C1306 vdd.t203 gnd 0.026412f
C1307 vdd.n161 gnd 0.181521f
C1308 vdd.n162 gnd 0.115189f
C1309 vdd.t155 gnd 0.026412f
C1310 vdd.t181 gnd 0.026412f
C1311 vdd.n163 gnd 0.181521f
C1312 vdd.n164 gnd 0.115189f
C1313 vdd.n165 gnd 0.004502f
C1314 vdd.n166 gnd 0.004178f
C1315 vdd.n167 gnd 0.002311f
C1316 vdd.n168 gnd 0.005306f
C1317 vdd.n169 gnd 0.002245f
C1318 vdd.n170 gnd 0.002377f
C1319 vdd.n171 gnd 0.004178f
C1320 vdd.n172 gnd 0.002245f
C1321 vdd.n173 gnd 0.005306f
C1322 vdd.n174 gnd 0.002377f
C1323 vdd.n175 gnd 0.004178f
C1324 vdd.n176 gnd 0.002245f
C1325 vdd.n177 gnd 0.00398f
C1326 vdd.n178 gnd 0.003992f
C1327 vdd.t198 gnd 0.0114f
C1328 vdd.n179 gnd 0.025366f
C1329 vdd.n180 gnd 0.132009f
C1330 vdd.n181 gnd 0.002245f
C1331 vdd.n182 gnd 0.002377f
C1332 vdd.n183 gnd 0.005306f
C1333 vdd.n184 gnd 0.005306f
C1334 vdd.n185 gnd 0.002377f
C1335 vdd.n186 gnd 0.002245f
C1336 vdd.n187 gnd 0.004178f
C1337 vdd.n188 gnd 0.004178f
C1338 vdd.n189 gnd 0.002245f
C1339 vdd.n190 gnd 0.002377f
C1340 vdd.n191 gnd 0.005306f
C1341 vdd.n192 gnd 0.005306f
C1342 vdd.n193 gnd 0.002377f
C1343 vdd.n194 gnd 0.002245f
C1344 vdd.n195 gnd 0.004178f
C1345 vdd.n196 gnd 0.004178f
C1346 vdd.n197 gnd 0.002245f
C1347 vdd.n198 gnd 0.002377f
C1348 vdd.n199 gnd 0.005306f
C1349 vdd.n200 gnd 0.005306f
C1350 vdd.n201 gnd 0.012545f
C1351 vdd.n202 gnd 0.002311f
C1352 vdd.n203 gnd 0.002245f
C1353 vdd.n204 gnd 0.010799f
C1354 vdd.n205 gnd 0.007302f
C1355 vdd.n206 gnd 0.050984f
C1356 vdd.n207 gnd 0.183708f
C1357 vdd.n208 gnd 0.004502f
C1358 vdd.n209 gnd 0.004178f
C1359 vdd.n210 gnd 0.002311f
C1360 vdd.n211 gnd 0.005306f
C1361 vdd.n212 gnd 0.002245f
C1362 vdd.n213 gnd 0.002377f
C1363 vdd.n214 gnd 0.004178f
C1364 vdd.n215 gnd 0.002245f
C1365 vdd.n216 gnd 0.005306f
C1366 vdd.n217 gnd 0.002377f
C1367 vdd.n218 gnd 0.004178f
C1368 vdd.n219 gnd 0.002245f
C1369 vdd.n220 gnd 0.00398f
C1370 vdd.n221 gnd 0.003992f
C1371 vdd.t209 gnd 0.0114f
C1372 vdd.n222 gnd 0.025366f
C1373 vdd.n223 gnd 0.132009f
C1374 vdd.n224 gnd 0.002245f
C1375 vdd.n225 gnd 0.002377f
C1376 vdd.n226 gnd 0.005306f
C1377 vdd.n227 gnd 0.005306f
C1378 vdd.n228 gnd 0.002377f
C1379 vdd.n229 gnd 0.002245f
C1380 vdd.n230 gnd 0.004178f
C1381 vdd.n231 gnd 0.004178f
C1382 vdd.n232 gnd 0.002245f
C1383 vdd.n233 gnd 0.002377f
C1384 vdd.n234 gnd 0.005306f
C1385 vdd.n235 gnd 0.005306f
C1386 vdd.n236 gnd 0.002377f
C1387 vdd.n237 gnd 0.002245f
C1388 vdd.n238 gnd 0.004178f
C1389 vdd.n239 gnd 0.004178f
C1390 vdd.n240 gnd 0.002245f
C1391 vdd.n241 gnd 0.002377f
C1392 vdd.n242 gnd 0.005306f
C1393 vdd.n243 gnd 0.005306f
C1394 vdd.n244 gnd 0.012545f
C1395 vdd.n245 gnd 0.002311f
C1396 vdd.n246 gnd 0.002245f
C1397 vdd.n247 gnd 0.010799f
C1398 vdd.n248 gnd 0.007539f
C1399 vdd.t210 gnd 0.026412f
C1400 vdd.t172 gnd 0.026412f
C1401 vdd.n249 gnd 0.181521f
C1402 vdd.n250 gnd 0.142739f
C1403 vdd.t202 gnd 0.026412f
C1404 vdd.t208 gnd 0.026412f
C1405 vdd.n251 gnd 0.181521f
C1406 vdd.n252 gnd 0.115189f
C1407 vdd.t165 gnd 0.026412f
C1408 vdd.t191 gnd 0.026412f
C1409 vdd.n253 gnd 0.181521f
C1410 vdd.n254 gnd 0.115189f
C1411 vdd.n255 gnd 0.004502f
C1412 vdd.n256 gnd 0.004178f
C1413 vdd.n257 gnd 0.002311f
C1414 vdd.n258 gnd 0.005306f
C1415 vdd.n259 gnd 0.002245f
C1416 vdd.n260 gnd 0.002377f
C1417 vdd.n261 gnd 0.004178f
C1418 vdd.n262 gnd 0.002245f
C1419 vdd.n263 gnd 0.005306f
C1420 vdd.n264 gnd 0.002377f
C1421 vdd.n265 gnd 0.004178f
C1422 vdd.n266 gnd 0.002245f
C1423 vdd.n267 gnd 0.00398f
C1424 vdd.n268 gnd 0.003992f
C1425 vdd.t201 gnd 0.0114f
C1426 vdd.n269 gnd 0.025366f
C1427 vdd.n270 gnd 0.132009f
C1428 vdd.n271 gnd 0.002245f
C1429 vdd.n272 gnd 0.002377f
C1430 vdd.n273 gnd 0.005306f
C1431 vdd.n274 gnd 0.005306f
C1432 vdd.n275 gnd 0.002377f
C1433 vdd.n276 gnd 0.002245f
C1434 vdd.n277 gnd 0.004178f
C1435 vdd.n278 gnd 0.004178f
C1436 vdd.n279 gnd 0.002245f
C1437 vdd.n280 gnd 0.002377f
C1438 vdd.n281 gnd 0.005306f
C1439 vdd.n282 gnd 0.005306f
C1440 vdd.n283 gnd 0.002377f
C1441 vdd.n284 gnd 0.002245f
C1442 vdd.n285 gnd 0.004178f
C1443 vdd.n286 gnd 0.004178f
C1444 vdd.n287 gnd 0.002245f
C1445 vdd.n288 gnd 0.002377f
C1446 vdd.n289 gnd 0.005306f
C1447 vdd.n290 gnd 0.005306f
C1448 vdd.n291 gnd 0.012545f
C1449 vdd.n292 gnd 0.002311f
C1450 vdd.n293 gnd 0.002245f
C1451 vdd.n294 gnd 0.010799f
C1452 vdd.n295 gnd 0.007302f
C1453 vdd.n296 gnd 0.050984f
C1454 vdd.n297 gnd 0.198842f
C1455 vdd.n298 gnd 0.006305f
C1456 vdd.n299 gnd 0.008204f
C1457 vdd.n300 gnd 0.006603f
C1458 vdd.n301 gnd 0.006603f
C1459 vdd.n302 gnd 0.008204f
C1460 vdd.n303 gnd 0.008204f
C1461 vdd.n304 gnd 0.599442f
C1462 vdd.n305 gnd 0.008204f
C1463 vdd.n306 gnd 0.008204f
C1464 vdd.n307 gnd 0.008204f
C1465 vdd.n308 gnd 0.649745f
C1466 vdd.n309 gnd 0.008204f
C1467 vdd.n310 gnd 0.008204f
C1468 vdd.n311 gnd 0.008204f
C1469 vdd.n312 gnd 0.008204f
C1470 vdd.n313 gnd 0.006603f
C1471 vdd.n314 gnd 0.008204f
C1472 vdd.t180 gnd 0.41919f
C1473 vdd.n315 gnd 0.008204f
C1474 vdd.n316 gnd 0.008204f
C1475 vdd.n317 gnd 0.008204f
C1476 vdd.n318 gnd 0.83838f
C1477 vdd.n319 gnd 0.008204f
C1478 vdd.n320 gnd 0.008204f
C1479 vdd.n321 gnd 0.008204f
C1480 vdd.n322 gnd 0.008204f
C1481 vdd.n323 gnd 0.008204f
C1482 vdd.n324 gnd 0.006603f
C1483 vdd.n325 gnd 0.008204f
C1484 vdd.n326 gnd 0.008204f
C1485 vdd.n327 gnd 0.008204f
C1486 vdd.n328 gnd 0.019993f
C1487 vdd.n329 gnd 2.00373f
C1488 vdd.n330 gnd 0.020451f
C1489 vdd.n331 gnd 0.008204f
C1490 vdd.n332 gnd 0.008204f
C1491 vdd.n334 gnd 0.008204f
C1492 vdd.n335 gnd 0.008204f
C1493 vdd.n336 gnd 0.006603f
C1494 vdd.n337 gnd 0.006603f
C1495 vdd.n338 gnd 0.008204f
C1496 vdd.n339 gnd 0.008204f
C1497 vdd.n340 gnd 0.008204f
C1498 vdd.n341 gnd 0.008204f
C1499 vdd.n342 gnd 0.008204f
C1500 vdd.n343 gnd 0.008204f
C1501 vdd.n344 gnd 0.006603f
C1502 vdd.n346 gnd 0.008204f
C1503 vdd.n347 gnd 0.008204f
C1504 vdd.n348 gnd 0.008204f
C1505 vdd.n349 gnd 0.008204f
C1506 vdd.n350 gnd 0.008204f
C1507 vdd.n351 gnd 0.006603f
C1508 vdd.n353 gnd 0.008204f
C1509 vdd.n354 gnd 0.008204f
C1510 vdd.n355 gnd 0.008204f
C1511 vdd.n356 gnd 0.008204f
C1512 vdd.n357 gnd 0.008204f
C1513 vdd.n358 gnd 0.006603f
C1514 vdd.n360 gnd 0.008204f
C1515 vdd.n361 gnd 0.008204f
C1516 vdd.n362 gnd 0.008204f
C1517 vdd.n363 gnd 0.008204f
C1518 vdd.n364 gnd 0.005514f
C1519 vdd.t142 gnd 0.100927f
C1520 vdd.t141 gnd 0.107863f
C1521 vdd.t140 gnd 0.13181f
C1522 vdd.n365 gnd 0.168961f
C1523 vdd.n366 gnd 0.142618f
C1524 vdd.n368 gnd 0.008204f
C1525 vdd.n369 gnd 0.008204f
C1526 vdd.n370 gnd 0.006603f
C1527 vdd.n371 gnd 0.008204f
C1528 vdd.n373 gnd 0.008204f
C1529 vdd.n374 gnd 0.008204f
C1530 vdd.n375 gnd 0.008204f
C1531 vdd.n376 gnd 0.008204f
C1532 vdd.n377 gnd 0.006603f
C1533 vdd.n379 gnd 0.008204f
C1534 vdd.n380 gnd 0.008204f
C1535 vdd.n381 gnd 0.008204f
C1536 vdd.n382 gnd 0.008204f
C1537 vdd.n383 gnd 0.008204f
C1538 vdd.n384 gnd 0.006603f
C1539 vdd.n386 gnd 0.008204f
C1540 vdd.n387 gnd 0.008204f
C1541 vdd.n388 gnd 0.008204f
C1542 vdd.n389 gnd 0.008204f
C1543 vdd.n390 gnd 0.008204f
C1544 vdd.n391 gnd 0.006603f
C1545 vdd.n393 gnd 0.008204f
C1546 vdd.n394 gnd 0.008204f
C1547 vdd.n395 gnd 0.008204f
C1548 vdd.n396 gnd 0.008204f
C1549 vdd.n397 gnd 0.008204f
C1550 vdd.n398 gnd 0.006603f
C1551 vdd.n400 gnd 0.008204f
C1552 vdd.n401 gnd 0.008204f
C1553 vdd.n402 gnd 0.008204f
C1554 vdd.n403 gnd 0.008204f
C1555 vdd.n404 gnd 0.006537f
C1556 vdd.t139 gnd 0.100927f
C1557 vdd.t138 gnd 0.107863f
C1558 vdd.t137 gnd 0.13181f
C1559 vdd.n405 gnd 0.168961f
C1560 vdd.n406 gnd 0.142618f
C1561 vdd.n408 gnd 0.008204f
C1562 vdd.n409 gnd 0.008204f
C1563 vdd.n410 gnd 0.006603f
C1564 vdd.n411 gnd 0.008204f
C1565 vdd.n413 gnd 0.008204f
C1566 vdd.n414 gnd 0.008204f
C1567 vdd.n415 gnd 0.008204f
C1568 vdd.n416 gnd 0.008204f
C1569 vdd.n417 gnd 0.006603f
C1570 vdd.n419 gnd 0.008204f
C1571 vdd.n420 gnd 0.008204f
C1572 vdd.n421 gnd 0.008204f
C1573 vdd.n422 gnd 0.008204f
C1574 vdd.n423 gnd 0.008204f
C1575 vdd.n424 gnd 0.006603f
C1576 vdd.n426 gnd 0.008204f
C1577 vdd.n427 gnd 0.008204f
C1578 vdd.n428 gnd 0.008204f
C1579 vdd.n429 gnd 0.008204f
C1580 vdd.n430 gnd 0.008204f
C1581 vdd.n431 gnd 0.006603f
C1582 vdd.n433 gnd 0.008204f
C1583 vdd.n434 gnd 0.008204f
C1584 vdd.n435 gnd 0.008204f
C1585 vdd.n436 gnd 0.008204f
C1586 vdd.n437 gnd 0.008204f
C1587 vdd.n438 gnd 0.006603f
C1588 vdd.n440 gnd 0.008204f
C1589 vdd.n441 gnd 0.008204f
C1590 vdd.n442 gnd 0.008204f
C1591 vdd.n443 gnd 0.008204f
C1592 vdd.n444 gnd 0.008204f
C1593 vdd.n445 gnd 0.008204f
C1594 vdd.n446 gnd 0.006603f
C1595 vdd.n447 gnd 0.008204f
C1596 vdd.n448 gnd 0.008204f
C1597 vdd.n449 gnd 0.006603f
C1598 vdd.n450 gnd 0.008204f
C1599 vdd.n451 gnd 0.006603f
C1600 vdd.n452 gnd 0.008204f
C1601 vdd.n453 gnd 0.006603f
C1602 vdd.n454 gnd 0.008204f
C1603 vdd.n455 gnd 0.008204f
C1604 vdd.n456 gnd 0.456917f
C1605 vdd.t158 gnd 0.41919f
C1606 vdd.n457 gnd 0.008204f
C1607 vdd.n458 gnd 0.006603f
C1608 vdd.n459 gnd 0.008204f
C1609 vdd.n460 gnd 0.006603f
C1610 vdd.n461 gnd 0.008204f
C1611 vdd.t173 gnd 0.41919f
C1612 vdd.n462 gnd 0.008204f
C1613 vdd.n463 gnd 0.006603f
C1614 vdd.n464 gnd 0.008204f
C1615 vdd.n465 gnd 0.006603f
C1616 vdd.n466 gnd 0.008204f
C1617 vdd.t182 gnd 0.41919f
C1618 vdd.n467 gnd 0.523988f
C1619 vdd.n468 gnd 0.008204f
C1620 vdd.n469 gnd 0.006603f
C1621 vdd.n470 gnd 0.008204f
C1622 vdd.n471 gnd 0.006603f
C1623 vdd.n472 gnd 0.008204f
C1624 vdd.n473 gnd 0.83838f
C1625 vdd.n474 gnd 0.008204f
C1626 vdd.n475 gnd 0.006603f
C1627 vdd.n476 gnd 0.019993f
C1628 vdd.n477 gnd 0.00548f
C1629 vdd.n478 gnd 0.019993f
C1630 vdd.t86 gnd 0.41919f
C1631 vdd.n479 gnd 0.019993f
C1632 vdd.n480 gnd 0.00548f
C1633 vdd.n481 gnd 0.007055f
C1634 vdd.n482 gnd 0.006603f
C1635 vdd.n483 gnd 0.008204f
C1636 vdd.n484 gnd 9.90127f
C1637 vdd.n515 gnd 0.020451f
C1638 vdd.n516 gnd 1.15277f
C1639 vdd.n517 gnd 0.008204f
C1640 vdd.n518 gnd 0.006603f
C1641 vdd.n519 gnd 0.00525f
C1642 vdd.n520 gnd 0.034447f
C1643 vdd.n521 gnd 0.006603f
C1644 vdd.n522 gnd 0.008204f
C1645 vdd.n523 gnd 0.008204f
C1646 vdd.n524 gnd 0.008204f
C1647 vdd.n525 gnd 0.008204f
C1648 vdd.n526 gnd 0.008204f
C1649 vdd.n527 gnd 0.008204f
C1650 vdd.n528 gnd 0.008204f
C1651 vdd.n529 gnd 0.008204f
C1652 vdd.n530 gnd 0.008204f
C1653 vdd.n531 gnd 0.008204f
C1654 vdd.n532 gnd 0.008204f
C1655 vdd.n533 gnd 0.008204f
C1656 vdd.n534 gnd 0.008204f
C1657 vdd.n535 gnd 0.008204f
C1658 vdd.n536 gnd 0.005514f
C1659 vdd.n537 gnd 0.008204f
C1660 vdd.n538 gnd 0.008204f
C1661 vdd.n539 gnd 0.008204f
C1662 vdd.n540 gnd 0.008204f
C1663 vdd.n541 gnd 0.008204f
C1664 vdd.n542 gnd 0.008204f
C1665 vdd.n543 gnd 0.008204f
C1666 vdd.n544 gnd 0.008204f
C1667 vdd.n545 gnd 0.008204f
C1668 vdd.n546 gnd 0.008204f
C1669 vdd.n547 gnd 0.008204f
C1670 vdd.n548 gnd 0.008204f
C1671 vdd.n549 gnd 0.008204f
C1672 vdd.n550 gnd 0.008204f
C1673 vdd.n551 gnd 0.008204f
C1674 vdd.n552 gnd 0.008204f
C1675 vdd.n553 gnd 0.008204f
C1676 vdd.n554 gnd 0.008204f
C1677 vdd.n555 gnd 0.008204f
C1678 vdd.n556 gnd 0.006537f
C1679 vdd.t111 gnd 0.100927f
C1680 vdd.t112 gnd 0.107863f
C1681 vdd.t110 gnd 0.13181f
C1682 vdd.n557 gnd 0.168961f
C1683 vdd.n558 gnd 0.141958f
C1684 vdd.n559 gnd 0.008204f
C1685 vdd.n560 gnd 0.008204f
C1686 vdd.n561 gnd 0.008204f
C1687 vdd.n562 gnd 0.008204f
C1688 vdd.n563 gnd 0.008204f
C1689 vdd.n564 gnd 0.008204f
C1690 vdd.n565 gnd 0.008204f
C1691 vdd.n566 gnd 0.008204f
C1692 vdd.n567 gnd 0.008204f
C1693 vdd.n568 gnd 0.008204f
C1694 vdd.n569 gnd 0.008204f
C1695 vdd.n570 gnd 0.008204f
C1696 vdd.n571 gnd 0.008204f
C1697 vdd.n572 gnd 0.00525f
C1698 vdd.n575 gnd 0.005579f
C1699 vdd.n576 gnd 0.005579f
C1700 vdd.n577 gnd 0.005579f
C1701 vdd.n578 gnd 0.005579f
C1702 vdd.n579 gnd 0.005579f
C1703 vdd.n580 gnd 0.005579f
C1704 vdd.n582 gnd 0.005579f
C1705 vdd.n583 gnd 0.005579f
C1706 vdd.n585 gnd 0.005579f
C1707 vdd.n586 gnd 0.004061f
C1708 vdd.n588 gnd 0.005579f
C1709 vdd.t70 gnd 0.225427f
C1710 vdd.t69 gnd 0.230753f
C1711 vdd.t67 gnd 0.147168f
C1712 vdd.n589 gnd 0.079536f
C1713 vdd.n590 gnd 0.045115f
C1714 vdd.n591 gnd 0.007973f
C1715 vdd.n592 gnd 0.012667f
C1716 vdd.n594 gnd 0.005579f
C1717 vdd.n595 gnd 0.570099f
C1718 vdd.n596 gnd 0.011945f
C1719 vdd.n597 gnd 0.011945f
C1720 vdd.n598 gnd 0.005579f
C1721 vdd.n599 gnd 0.012667f
C1722 vdd.n600 gnd 0.005579f
C1723 vdd.n601 gnd 0.005579f
C1724 vdd.n602 gnd 0.005579f
C1725 vdd.n603 gnd 0.005579f
C1726 vdd.n604 gnd 0.005579f
C1727 vdd.n606 gnd 0.005579f
C1728 vdd.n607 gnd 0.005579f
C1729 vdd.n609 gnd 0.005579f
C1730 vdd.n610 gnd 0.005579f
C1731 vdd.n612 gnd 0.005579f
C1732 vdd.n613 gnd 0.005579f
C1733 vdd.n615 gnd 0.005579f
C1734 vdd.n616 gnd 0.005579f
C1735 vdd.n618 gnd 0.005579f
C1736 vdd.n619 gnd 0.005579f
C1737 vdd.n621 gnd 0.005579f
C1738 vdd.t84 gnd 0.225427f
C1739 vdd.t83 gnd 0.230753f
C1740 vdd.t82 gnd 0.147168f
C1741 vdd.n622 gnd 0.079536f
C1742 vdd.n623 gnd 0.045115f
C1743 vdd.n624 gnd 0.005579f
C1744 vdd.n626 gnd 0.005579f
C1745 vdd.n627 gnd 0.005579f
C1746 vdd.t68 gnd 0.285049f
C1747 vdd.n628 gnd 0.005579f
C1748 vdd.n629 gnd 0.005579f
C1749 vdd.n630 gnd 0.005579f
C1750 vdd.n631 gnd 0.005579f
C1751 vdd.n632 gnd 0.005579f
C1752 vdd.n633 gnd 0.570099f
C1753 vdd.n634 gnd 0.005579f
C1754 vdd.n635 gnd 0.005579f
C1755 vdd.n636 gnd 0.448533f
C1756 vdd.n637 gnd 0.005579f
C1757 vdd.n638 gnd 0.005579f
C1758 vdd.n639 gnd 0.005579f
C1759 vdd.n640 gnd 0.005579f
C1760 vdd.n641 gnd 0.570099f
C1761 vdd.n642 gnd 0.005579f
C1762 vdd.n643 gnd 0.005579f
C1763 vdd.n644 gnd 0.005579f
C1764 vdd.n645 gnd 0.005579f
C1765 vdd.n646 gnd 0.005579f
C1766 vdd.t19 gnd 0.285049f
C1767 vdd.n647 gnd 0.005579f
C1768 vdd.n648 gnd 0.005579f
C1769 vdd.n649 gnd 0.005579f
C1770 vdd.n650 gnd 0.005579f
C1771 vdd.n651 gnd 0.005579f
C1772 vdd.t36 gnd 0.285049f
C1773 vdd.n652 gnd 0.005579f
C1774 vdd.n653 gnd 0.005579f
C1775 vdd.n654 gnd 0.549139f
C1776 vdd.n655 gnd 0.005579f
C1777 vdd.n656 gnd 0.005579f
C1778 vdd.n657 gnd 0.005579f
C1779 vdd.t35 gnd 0.285049f
C1780 vdd.n658 gnd 0.005579f
C1781 vdd.n659 gnd 0.005579f
C1782 vdd.n660 gnd 0.423382f
C1783 vdd.n661 gnd 0.005579f
C1784 vdd.n662 gnd 0.005579f
C1785 vdd.n663 gnd 0.005579f
C1786 vdd.n664 gnd 0.398231f
C1787 vdd.n665 gnd 0.005579f
C1788 vdd.n666 gnd 0.005579f
C1789 vdd.n667 gnd 0.297625f
C1790 vdd.n668 gnd 0.005579f
C1791 vdd.n669 gnd 0.005579f
C1792 vdd.n670 gnd 0.005579f
C1793 vdd.n671 gnd 0.523988f
C1794 vdd.n672 gnd 0.005579f
C1795 vdd.n673 gnd 0.005579f
C1796 vdd.t44 gnd 0.285049f
C1797 vdd.n674 gnd 0.005579f
C1798 vdd.n675 gnd 0.005579f
C1799 vdd.n676 gnd 0.005579f
C1800 vdd.n677 gnd 0.570099f
C1801 vdd.n678 gnd 0.005579f
C1802 vdd.n679 gnd 0.005579f
C1803 vdd.t45 gnd 0.285049f
C1804 vdd.n680 gnd 0.005579f
C1805 vdd.n681 gnd 0.005579f
C1806 vdd.n682 gnd 0.005579f
C1807 vdd.t13 gnd 0.285049f
C1808 vdd.n683 gnd 0.005579f
C1809 vdd.n684 gnd 0.005579f
C1810 vdd.n685 gnd 0.005579f
C1811 vdd.t91 gnd 0.230753f
C1812 vdd.t89 gnd 0.147168f
C1813 vdd.t92 gnd 0.230753f
C1814 vdd.n686 gnd 0.129693f
C1815 vdd.n687 gnd 0.01616f
C1816 vdd.n688 gnd 0.005579f
C1817 vdd.t90 gnd 0.205403f
C1818 vdd.n689 gnd 0.005579f
C1819 vdd.n690 gnd 0.005579f
C1820 vdd.n691 gnd 0.490452f
C1821 vdd.n692 gnd 0.005579f
C1822 vdd.n693 gnd 0.005579f
C1823 vdd.n694 gnd 0.005579f
C1824 vdd.n695 gnd 0.33116f
C1825 vdd.n696 gnd 0.005579f
C1826 vdd.n697 gnd 0.005579f
C1827 vdd.t14 gnd 0.117373f
C1828 vdd.n698 gnd 0.364695f
C1829 vdd.n699 gnd 0.005579f
C1830 vdd.n700 gnd 0.005579f
C1831 vdd.n701 gnd 0.005579f
C1832 vdd.n702 gnd 0.456917f
C1833 vdd.n703 gnd 0.005579f
C1834 vdd.n704 gnd 0.005579f
C1835 vdd.t27 gnd 0.285049f
C1836 vdd.n705 gnd 0.005579f
C1837 vdd.n706 gnd 0.005579f
C1838 vdd.n707 gnd 0.005579f
C1839 vdd.t23 gnd 0.285049f
C1840 vdd.n708 gnd 0.005579f
C1841 vdd.n709 gnd 0.005579f
C1842 vdd.t48 gnd 0.285049f
C1843 vdd.n710 gnd 0.005579f
C1844 vdd.n711 gnd 0.005579f
C1845 vdd.n712 gnd 0.005579f
C1846 vdd.t5 gnd 0.192827f
C1847 vdd.n713 gnd 0.005579f
C1848 vdd.n714 gnd 0.005579f
C1849 vdd.n715 gnd 0.503028f
C1850 vdd.n716 gnd 0.005579f
C1851 vdd.n717 gnd 0.005579f
C1852 vdd.n718 gnd 0.005579f
C1853 vdd.t49 gnd 0.285049f
C1854 vdd.n719 gnd 0.005579f
C1855 vdd.n720 gnd 0.005579f
C1856 vdd.t59 gnd 0.272474f
C1857 vdd.n721 gnd 0.377271f
C1858 vdd.n722 gnd 0.005579f
C1859 vdd.n723 gnd 0.005579f
C1860 vdd.n724 gnd 0.005579f
C1861 vdd.t9 gnd 0.285049f
C1862 vdd.n725 gnd 0.005579f
C1863 vdd.n726 gnd 0.005579f
C1864 vdd.t53 gnd 0.285049f
C1865 vdd.n727 gnd 0.005579f
C1866 vdd.n728 gnd 0.005579f
C1867 vdd.n729 gnd 0.005579f
C1868 vdd.n730 gnd 0.570099f
C1869 vdd.n731 gnd 0.005579f
C1870 vdd.n732 gnd 0.005579f
C1871 vdd.t31 gnd 0.285049f
C1872 vdd.n733 gnd 0.005579f
C1873 vdd.n734 gnd 0.005579f
C1874 vdd.n735 gnd 0.005579f
C1875 vdd.n736 gnd 0.394039f
C1876 vdd.n737 gnd 0.005579f
C1877 vdd.n738 gnd 0.005579f
C1878 vdd.n739 gnd 0.005579f
C1879 vdd.n740 gnd 0.005579f
C1880 vdd.n741 gnd 0.005579f
C1881 vdd.t124 gnd 0.285049f
C1882 vdd.n742 gnd 0.005579f
C1883 vdd.n743 gnd 0.005579f
C1884 vdd.t11 gnd 0.285049f
C1885 vdd.n744 gnd 0.005579f
C1886 vdd.n745 gnd 0.011945f
C1887 vdd.n746 gnd 0.011945f
C1888 vdd.n747 gnd 0.645553f
C1889 vdd.n748 gnd 0.005579f
C1890 vdd.n749 gnd 0.005579f
C1891 vdd.t42 gnd 0.285049f
C1892 vdd.n750 gnd 0.011945f
C1893 vdd.n751 gnd 0.005579f
C1894 vdd.n752 gnd 0.005579f
C1895 vdd.t40 gnd 0.486261f
C1896 vdd.n770 gnd 0.012667f
C1897 vdd.n788 gnd 0.011945f
C1898 vdd.n789 gnd 0.005579f
C1899 vdd.n790 gnd 0.011945f
C1900 vdd.t136 gnd 0.225427f
C1901 vdd.t135 gnd 0.230753f
C1902 vdd.t134 gnd 0.147168f
C1903 vdd.n791 gnd 0.079536f
C1904 vdd.n792 gnd 0.045115f
C1905 vdd.n793 gnd 0.012667f
C1906 vdd.n794 gnd 0.005579f
C1907 vdd.n795 gnd 0.335352f
C1908 vdd.n796 gnd 0.011945f
C1909 vdd.n797 gnd 0.005579f
C1910 vdd.n798 gnd 0.012667f
C1911 vdd.n799 gnd 0.005579f
C1912 vdd.t119 gnd 0.225427f
C1913 vdd.t118 gnd 0.230753f
C1914 vdd.t116 gnd 0.147168f
C1915 vdd.n800 gnd 0.079536f
C1916 vdd.n801 gnd 0.045115f
C1917 vdd.n802 gnd 0.007973f
C1918 vdd.n803 gnd 0.005579f
C1919 vdd.n804 gnd 0.005579f
C1920 vdd.t117 gnd 0.285049f
C1921 vdd.n805 gnd 0.005579f
C1922 vdd.t55 gnd 0.285049f
C1923 vdd.n806 gnd 0.005579f
C1924 vdd.n807 gnd 0.005579f
C1925 vdd.n808 gnd 0.005579f
C1926 vdd.n809 gnd 0.005579f
C1927 vdd.n810 gnd 0.005579f
C1928 vdd.n811 gnd 0.570099f
C1929 vdd.n812 gnd 0.005579f
C1930 vdd.n813 gnd 0.005579f
C1931 vdd.t25 gnd 0.285049f
C1932 vdd.n814 gnd 0.005579f
C1933 vdd.n815 gnd 0.005579f
C1934 vdd.n816 gnd 0.005579f
C1935 vdd.n817 gnd 0.005579f
C1936 vdd.n818 gnd 0.410806f
C1937 vdd.n819 gnd 0.005579f
C1938 vdd.n820 gnd 0.005579f
C1939 vdd.n821 gnd 0.005579f
C1940 vdd.n822 gnd 0.005579f
C1941 vdd.n823 gnd 0.005579f
C1942 vdd.t6 gnd 0.285049f
C1943 vdd.n824 gnd 0.005579f
C1944 vdd.n825 gnd 0.005579f
C1945 vdd.t46 gnd 0.285049f
C1946 vdd.n826 gnd 0.005579f
C1947 vdd.n827 gnd 0.005579f
C1948 vdd.n828 gnd 0.005579f
C1949 vdd.t30 gnd 0.285049f
C1950 vdd.n829 gnd 0.005579f
C1951 vdd.n830 gnd 0.005579f
C1952 vdd.t7 gnd 0.285049f
C1953 vdd.n831 gnd 0.005579f
C1954 vdd.n832 gnd 0.005579f
C1955 vdd.n833 gnd 0.005579f
C1956 vdd.t28 gnd 0.272474f
C1957 vdd.n834 gnd 0.005579f
C1958 vdd.n835 gnd 0.005579f
C1959 vdd.n836 gnd 0.423382f
C1960 vdd.n837 gnd 0.005579f
C1961 vdd.n838 gnd 0.005579f
C1962 vdd.n839 gnd 0.005579f
C1963 vdd.t50 gnd 0.285049f
C1964 vdd.n840 gnd 0.005579f
C1965 vdd.n841 gnd 0.005579f
C1966 vdd.t16 gnd 0.192827f
C1967 vdd.n842 gnd 0.297625f
C1968 vdd.n843 gnd 0.005579f
C1969 vdd.n844 gnd 0.005579f
C1970 vdd.n845 gnd 0.005579f
C1971 vdd.n846 gnd 0.523988f
C1972 vdd.n847 gnd 0.005579f
C1973 vdd.n848 gnd 0.005579f
C1974 vdd.t57 gnd 0.285049f
C1975 vdd.n849 gnd 0.005579f
C1976 vdd.n850 gnd 0.005579f
C1977 vdd.n851 gnd 0.005579f
C1978 vdd.n852 gnd 0.570099f
C1979 vdd.n853 gnd 0.005579f
C1980 vdd.n854 gnd 0.005579f
C1981 vdd.t22 gnd 0.285049f
C1982 vdd.n855 gnd 0.005579f
C1983 vdd.n856 gnd 0.005579f
C1984 vdd.n857 gnd 0.005579f
C1985 vdd.t15 gnd 0.117373f
C1986 vdd.n858 gnd 0.005579f
C1987 vdd.n859 gnd 0.005579f
C1988 vdd.n860 gnd 0.005579f
C1989 vdd.t129 gnd 0.230753f
C1990 vdd.t127 gnd 0.147168f
C1991 vdd.t130 gnd 0.230753f
C1992 vdd.n861 gnd 0.129693f
C1993 vdd.n862 gnd 0.005579f
C1994 vdd.n863 gnd 0.005579f
C1995 vdd.t37 gnd 0.285049f
C1996 vdd.n864 gnd 0.005579f
C1997 vdd.n865 gnd 0.005579f
C1998 vdd.t128 gnd 0.205403f
C1999 vdd.n866 gnd 0.452725f
C2000 vdd.n867 gnd 0.005579f
C2001 vdd.n868 gnd 0.005579f
C2002 vdd.n869 gnd 0.005579f
C2003 vdd.n870 gnd 0.33116f
C2004 vdd.n871 gnd 0.005579f
C2005 vdd.n872 gnd 0.005579f
C2006 vdd.n873 gnd 0.364695f
C2007 vdd.n874 gnd 0.005579f
C2008 vdd.n875 gnd 0.005579f
C2009 vdd.n876 gnd 0.005579f
C2010 vdd.n877 gnd 0.456917f
C2011 vdd.n878 gnd 0.005579f
C2012 vdd.n879 gnd 0.005579f
C2013 vdd.t17 gnd 0.285049f
C2014 vdd.n880 gnd 0.005579f
C2015 vdd.n881 gnd 0.005579f
C2016 vdd.n882 gnd 0.005579f
C2017 vdd.n883 gnd 0.570099f
C2018 vdd.n884 gnd 0.005579f
C2019 vdd.n885 gnd 0.005579f
C2020 vdd.t18 gnd 0.285049f
C2021 vdd.n886 gnd 0.005579f
C2022 vdd.n887 gnd 0.005579f
C2023 vdd.n888 gnd 0.005579f
C2024 vdd.t58 gnd 0.285049f
C2025 vdd.n889 gnd 0.005579f
C2026 vdd.n890 gnd 0.005579f
C2027 vdd.n891 gnd 0.005579f
C2028 vdd.n892 gnd 0.005579f
C2029 vdd.n893 gnd 0.005579f
C2030 vdd.t52 gnd 0.285049f
C2031 vdd.n894 gnd 0.005579f
C2032 vdd.n895 gnd 0.005579f
C2033 vdd.n896 gnd 0.557523f
C2034 vdd.n897 gnd 0.005579f
C2035 vdd.n898 gnd 0.005579f
C2036 vdd.n899 gnd 0.005579f
C2037 vdd.t10 gnd 0.285049f
C2038 vdd.n900 gnd 0.005579f
C2039 vdd.n901 gnd 0.005579f
C2040 vdd.n902 gnd 0.431766f
C2041 vdd.n903 gnd 0.005579f
C2042 vdd.n904 gnd 0.005579f
C2043 vdd.n905 gnd 0.005579f
C2044 vdd.n906 gnd 0.570099f
C2045 vdd.n907 gnd 0.005579f
C2046 vdd.n908 gnd 0.005579f
C2047 vdd.n909 gnd 0.306009f
C2048 vdd.n910 gnd 0.005579f
C2049 vdd.n911 gnd 0.005579f
C2050 vdd.n912 gnd 0.005579f
C2051 vdd.n913 gnd 0.570099f
C2052 vdd.n914 gnd 0.005579f
C2053 vdd.n915 gnd 0.005579f
C2054 vdd.n916 gnd 0.005579f
C2055 vdd.n917 gnd 0.005579f
C2056 vdd.n918 gnd 0.005579f
C2057 vdd.t72 gnd 0.285049f
C2058 vdd.n919 gnd 0.005579f
C2059 vdd.n920 gnd 0.005579f
C2060 vdd.n921 gnd 0.005579f
C2061 vdd.n922 gnd 0.011945f
C2062 vdd.n923 gnd 0.011945f
C2063 vdd.n924 gnd 0.77131f
C2064 vdd.n925 gnd 0.005579f
C2065 vdd.n926 gnd 0.005579f
C2066 vdd.n927 gnd 0.406614f
C2067 vdd.n928 gnd 0.011945f
C2068 vdd.n929 gnd 0.005579f
C2069 vdd.n930 gnd 0.005579f
C2070 vdd.n931 gnd 10.253401f
C2071 vdd.n965 gnd 0.012667f
C2072 vdd.n966 gnd 0.005579f
C2073 vdd.n967 gnd 0.005579f
C2074 vdd.n968 gnd 0.00525f
C2075 vdd.n971 gnd 0.020451f
C2076 vdd.n972 gnd 0.00548f
C2077 vdd.n973 gnd 0.006603f
C2078 vdd.n975 gnd 0.008204f
C2079 vdd.n976 gnd 0.008204f
C2080 vdd.n977 gnd 0.006603f
C2081 vdd.n979 gnd 0.008204f
C2082 vdd.n980 gnd 0.008204f
C2083 vdd.n981 gnd 0.008204f
C2084 vdd.n982 gnd 0.008204f
C2085 vdd.n983 gnd 0.008204f
C2086 vdd.n984 gnd 0.006603f
C2087 vdd.n986 gnd 0.008204f
C2088 vdd.n987 gnd 0.008204f
C2089 vdd.n988 gnd 0.008204f
C2090 vdd.n989 gnd 0.008204f
C2091 vdd.n990 gnd 0.008204f
C2092 vdd.n991 gnd 0.006603f
C2093 vdd.n993 gnd 0.008204f
C2094 vdd.n994 gnd 0.008204f
C2095 vdd.n995 gnd 0.008204f
C2096 vdd.n996 gnd 0.008204f
C2097 vdd.n997 gnd 0.005514f
C2098 vdd.t81 gnd 0.100927f
C2099 vdd.t80 gnd 0.107863f
C2100 vdd.t79 gnd 0.13181f
C2101 vdd.n998 gnd 0.168961f
C2102 vdd.n999 gnd 0.141958f
C2103 vdd.n1001 gnd 0.008204f
C2104 vdd.n1002 gnd 0.008204f
C2105 vdd.n1003 gnd 0.006603f
C2106 vdd.n1004 gnd 0.008204f
C2107 vdd.n1006 gnd 0.008204f
C2108 vdd.n1007 gnd 0.008204f
C2109 vdd.n1008 gnd 0.008204f
C2110 vdd.n1009 gnd 0.008204f
C2111 vdd.n1010 gnd 0.006603f
C2112 vdd.n1012 gnd 0.008204f
C2113 vdd.n1013 gnd 0.008204f
C2114 vdd.n1014 gnd 0.008204f
C2115 vdd.n1015 gnd 0.008204f
C2116 vdd.n1016 gnd 0.008204f
C2117 vdd.n1017 gnd 0.006603f
C2118 vdd.n1019 gnd 0.008204f
C2119 vdd.n1020 gnd 0.008204f
C2120 vdd.n1021 gnd 0.008204f
C2121 vdd.n1022 gnd 0.008204f
C2122 vdd.n1023 gnd 0.008204f
C2123 vdd.n1024 gnd 0.006603f
C2124 vdd.n1026 gnd 0.008204f
C2125 vdd.n1027 gnd 0.008204f
C2126 vdd.n1028 gnd 0.008204f
C2127 vdd.n1029 gnd 0.008204f
C2128 vdd.n1030 gnd 0.008204f
C2129 vdd.n1031 gnd 0.006603f
C2130 vdd.n1033 gnd 0.008204f
C2131 vdd.n1034 gnd 0.008204f
C2132 vdd.n1035 gnd 0.008204f
C2133 vdd.n1036 gnd 0.008204f
C2134 vdd.n1037 gnd 0.006537f
C2135 vdd.t78 gnd 0.100927f
C2136 vdd.t77 gnd 0.107863f
C2137 vdd.t75 gnd 0.13181f
C2138 vdd.n1038 gnd 0.168961f
C2139 vdd.n1039 gnd 0.141958f
C2140 vdd.n1041 gnd 0.008204f
C2141 vdd.n1042 gnd 0.008204f
C2142 vdd.n1043 gnd 0.006603f
C2143 vdd.n1044 gnd 0.008204f
C2144 vdd.n1046 gnd 0.008204f
C2145 vdd.n1047 gnd 0.008204f
C2146 vdd.n1048 gnd 0.008204f
C2147 vdd.n1049 gnd 0.008204f
C2148 vdd.n1050 gnd 0.006603f
C2149 vdd.n1052 gnd 0.008204f
C2150 vdd.n1053 gnd 0.008204f
C2151 vdd.n1054 gnd 0.008204f
C2152 vdd.n1055 gnd 0.008204f
C2153 vdd.n1056 gnd 0.008204f
C2154 vdd.n1057 gnd 0.006603f
C2155 vdd.n1059 gnd 0.008204f
C2156 vdd.n1060 gnd 0.008204f
C2157 vdd.n1061 gnd 0.008204f
C2158 vdd.n1062 gnd 0.008204f
C2159 vdd.n1063 gnd 0.008204f
C2160 vdd.n1064 gnd 0.006603f
C2161 vdd.n1066 gnd 0.008204f
C2162 vdd.n1067 gnd 0.008204f
C2163 vdd.n1068 gnd 0.00525f
C2164 vdd.n1069 gnd 0.006603f
C2165 vdd.n1070 gnd 0.012667f
C2166 vdd.n1071 gnd 0.012667f
C2167 vdd.n1072 gnd 0.005579f
C2168 vdd.n1073 gnd 0.005579f
C2169 vdd.n1074 gnd 0.005579f
C2170 vdd.n1075 gnd 0.005579f
C2171 vdd.n1076 gnd 0.005579f
C2172 vdd.n1077 gnd 0.005579f
C2173 vdd.n1078 gnd 0.005579f
C2174 vdd.n1079 gnd 0.005579f
C2175 vdd.n1080 gnd 0.005579f
C2176 vdd.n1081 gnd 0.005579f
C2177 vdd.n1082 gnd 0.005579f
C2178 vdd.n1083 gnd 0.005579f
C2179 vdd.n1084 gnd 0.005579f
C2180 vdd.n1085 gnd 0.005579f
C2181 vdd.n1086 gnd 0.005579f
C2182 vdd.n1087 gnd 0.005579f
C2183 vdd.n1088 gnd 0.005579f
C2184 vdd.n1089 gnd 0.005579f
C2185 vdd.n1090 gnd 0.005579f
C2186 vdd.n1091 gnd 0.005579f
C2187 vdd.n1092 gnd 0.005579f
C2188 vdd.n1093 gnd 0.005579f
C2189 vdd.n1094 gnd 0.005579f
C2190 vdd.n1095 gnd 0.005579f
C2191 vdd.n1096 gnd 0.005579f
C2192 vdd.n1097 gnd 0.005579f
C2193 vdd.n1098 gnd 0.005579f
C2194 vdd.n1099 gnd 0.005579f
C2195 vdd.n1100 gnd 0.005579f
C2196 vdd.n1101 gnd 0.005579f
C2197 vdd.n1102 gnd 0.005579f
C2198 vdd.n1103 gnd 0.005579f
C2199 vdd.n1104 gnd 0.005579f
C2200 vdd.t73 gnd 0.225427f
C2201 vdd.t74 gnd 0.230753f
C2202 vdd.t71 gnd 0.147168f
C2203 vdd.n1105 gnd 0.079536f
C2204 vdd.n1106 gnd 0.045115f
C2205 vdd.n1107 gnd 0.007973f
C2206 vdd.n1108 gnd 0.005579f
C2207 vdd.t114 gnd 0.225427f
C2208 vdd.t115 gnd 0.230753f
C2209 vdd.t113 gnd 0.147168f
C2210 vdd.n1109 gnd 0.079536f
C2211 vdd.n1110 gnd 0.045115f
C2212 vdd.n1111 gnd 0.005579f
C2213 vdd.n1112 gnd 0.005579f
C2214 vdd.n1113 gnd 0.005579f
C2215 vdd.n1114 gnd 0.005579f
C2216 vdd.n1115 gnd 0.005579f
C2217 vdd.n1116 gnd 0.005579f
C2218 vdd.n1117 gnd 0.005579f
C2219 vdd.n1118 gnd 0.005579f
C2220 vdd.n1119 gnd 0.005579f
C2221 vdd.n1120 gnd 0.005579f
C2222 vdd.n1121 gnd 0.005579f
C2223 vdd.n1122 gnd 0.005579f
C2224 vdd.n1123 gnd 0.005579f
C2225 vdd.n1124 gnd 0.005579f
C2226 vdd.n1125 gnd 0.005579f
C2227 vdd.n1126 gnd 0.005579f
C2228 vdd.n1127 gnd 0.005579f
C2229 vdd.n1128 gnd 0.005579f
C2230 vdd.n1129 gnd 0.005579f
C2231 vdd.n1130 gnd 0.005579f
C2232 vdd.n1131 gnd 0.005579f
C2233 vdd.n1132 gnd 0.005579f
C2234 vdd.n1133 gnd 0.005579f
C2235 vdd.n1134 gnd 0.005579f
C2236 vdd.n1135 gnd 0.005579f
C2237 vdd.n1136 gnd 0.005579f
C2238 vdd.n1137 gnd 0.004061f
C2239 vdd.n1138 gnd 0.007973f
C2240 vdd.n1139 gnd 0.004307f
C2241 vdd.n1140 gnd 0.005579f
C2242 vdd.n1141 gnd 0.005579f
C2243 vdd.n1142 gnd 0.005579f
C2244 vdd.n1143 gnd 0.012667f
C2245 vdd.n1144 gnd 0.012667f
C2246 vdd.n1145 gnd 0.011945f
C2247 vdd.n1146 gnd 0.011945f
C2248 vdd.n1147 gnd 0.005579f
C2249 vdd.n1148 gnd 0.005579f
C2250 vdd.n1149 gnd 0.005579f
C2251 vdd.n1150 gnd 0.005579f
C2252 vdd.n1151 gnd 0.005579f
C2253 vdd.n1152 gnd 0.005579f
C2254 vdd.n1153 gnd 0.005579f
C2255 vdd.n1154 gnd 0.005579f
C2256 vdd.n1155 gnd 0.005579f
C2257 vdd.n1156 gnd 0.005579f
C2258 vdd.n1157 gnd 0.005579f
C2259 vdd.n1158 gnd 0.005579f
C2260 vdd.n1159 gnd 0.005579f
C2261 vdd.n1160 gnd 0.005579f
C2262 vdd.n1161 gnd 0.005579f
C2263 vdd.n1162 gnd 0.005579f
C2264 vdd.n1163 gnd 0.005579f
C2265 vdd.n1164 gnd 0.005579f
C2266 vdd.n1165 gnd 0.005579f
C2267 vdd.n1166 gnd 0.005579f
C2268 vdd.n1167 gnd 0.005579f
C2269 vdd.n1168 gnd 0.005579f
C2270 vdd.n1169 gnd 0.005579f
C2271 vdd.n1170 gnd 0.005579f
C2272 vdd.n1171 gnd 0.005579f
C2273 vdd.n1172 gnd 0.005579f
C2274 vdd.n1173 gnd 0.005579f
C2275 vdd.n1174 gnd 0.005579f
C2276 vdd.n1175 gnd 0.005579f
C2277 vdd.n1176 gnd 0.005579f
C2278 vdd.n1177 gnd 0.005579f
C2279 vdd.n1178 gnd 0.005579f
C2280 vdd.n1179 gnd 0.005579f
C2281 vdd.n1180 gnd 0.005579f
C2282 vdd.n1181 gnd 0.005579f
C2283 vdd.n1182 gnd 0.005579f
C2284 vdd.n1183 gnd 0.005579f
C2285 vdd.n1184 gnd 0.005579f
C2286 vdd.n1185 gnd 0.005579f
C2287 vdd.n1186 gnd 0.005579f
C2288 vdd.n1187 gnd 0.005579f
C2289 vdd.n1188 gnd 0.005579f
C2290 vdd.n1189 gnd 0.339544f
C2291 vdd.n1190 gnd 0.005579f
C2292 vdd.n1191 gnd 0.005579f
C2293 vdd.n1192 gnd 0.005579f
C2294 vdd.n1193 gnd 0.005579f
C2295 vdd.n1194 gnd 0.005579f
C2296 vdd.n1195 gnd 0.005579f
C2297 vdd.n1196 gnd 0.005579f
C2298 vdd.n1197 gnd 0.005579f
C2299 vdd.n1198 gnd 0.005579f
C2300 vdd.n1199 gnd 0.005579f
C2301 vdd.n1200 gnd 0.005579f
C2302 vdd.n1201 gnd 0.005579f
C2303 vdd.n1202 gnd 0.005579f
C2304 vdd.n1203 gnd 0.005579f
C2305 vdd.n1204 gnd 0.005579f
C2306 vdd.n1205 gnd 0.005579f
C2307 vdd.n1206 gnd 0.005579f
C2308 vdd.n1207 gnd 0.005579f
C2309 vdd.n1208 gnd 0.005579f
C2310 vdd.n1209 gnd 0.005579f
C2311 vdd.n1210 gnd 0.005579f
C2312 vdd.n1211 gnd 0.005579f
C2313 vdd.n1212 gnd 0.005579f
C2314 vdd.n1213 gnd 0.005579f
C2315 vdd.n1214 gnd 0.005579f
C2316 vdd.n1215 gnd 0.515604f
C2317 vdd.n1216 gnd 0.005579f
C2318 vdd.n1217 gnd 0.005579f
C2319 vdd.n1218 gnd 0.005579f
C2320 vdd.n1219 gnd 0.005579f
C2321 vdd.n1220 gnd 0.005579f
C2322 vdd.n1221 gnd 0.005579f
C2323 vdd.n1222 gnd 0.005579f
C2324 vdd.n1223 gnd 0.005579f
C2325 vdd.n1224 gnd 0.005579f
C2326 vdd.n1225 gnd 0.005579f
C2327 vdd.n1226 gnd 0.005579f
C2328 vdd.n1227 gnd 0.180252f
C2329 vdd.n1228 gnd 0.005579f
C2330 vdd.n1229 gnd 0.005579f
C2331 vdd.n1230 gnd 0.005579f
C2332 vdd.n1231 gnd 0.005579f
C2333 vdd.n1232 gnd 0.005579f
C2334 vdd.n1233 gnd 0.005579f
C2335 vdd.n1234 gnd 0.005579f
C2336 vdd.n1235 gnd 0.005579f
C2337 vdd.n1236 gnd 0.005579f
C2338 vdd.n1237 gnd 0.005579f
C2339 vdd.n1238 gnd 0.005579f
C2340 vdd.n1239 gnd 0.005579f
C2341 vdd.n1240 gnd 0.005579f
C2342 vdd.n1241 gnd 0.005579f
C2343 vdd.n1242 gnd 0.005579f
C2344 vdd.n1243 gnd 0.005579f
C2345 vdd.n1244 gnd 0.005579f
C2346 vdd.n1245 gnd 0.005579f
C2347 vdd.n1246 gnd 0.005579f
C2348 vdd.n1247 gnd 0.005579f
C2349 vdd.n1248 gnd 0.005579f
C2350 vdd.n1249 gnd 0.005579f
C2351 vdd.n1250 gnd 0.005579f
C2352 vdd.n1251 gnd 0.005579f
C2353 vdd.n1252 gnd 0.005579f
C2354 vdd.n1253 gnd 0.005579f
C2355 vdd.n1254 gnd 0.005579f
C2356 vdd.n1255 gnd 0.005579f
C2357 vdd.n1256 gnd 0.005579f
C2358 vdd.n1257 gnd 0.005579f
C2359 vdd.n1258 gnd 0.005579f
C2360 vdd.n1259 gnd 0.005579f
C2361 vdd.n1260 gnd 0.005579f
C2362 vdd.n1261 gnd 0.005579f
C2363 vdd.n1262 gnd 0.005579f
C2364 vdd.n1263 gnd 0.005579f
C2365 vdd.n1264 gnd 0.005579f
C2366 vdd.n1265 gnd 0.005579f
C2367 vdd.n1266 gnd 0.005579f
C2368 vdd.n1267 gnd 0.005579f
C2369 vdd.n1268 gnd 0.005579f
C2370 vdd.n1269 gnd 0.005579f
C2371 vdd.n1270 gnd 0.011945f
C2372 vdd.n1271 gnd 0.011945f
C2373 vdd.n1272 gnd 0.012667f
C2374 vdd.n1273 gnd 0.005579f
C2375 vdd.n1274 gnd 0.005579f
C2376 vdd.n1275 gnd 0.004307f
C2377 vdd.n1276 gnd 0.005579f
C2378 vdd.n1277 gnd 0.005579f
C2379 vdd.n1278 gnd 0.004061f
C2380 vdd.n1279 gnd 0.005579f
C2381 vdd.n1280 gnd 0.005579f
C2382 vdd.n1281 gnd 0.005579f
C2383 vdd.n1282 gnd 0.005579f
C2384 vdd.n1283 gnd 0.005579f
C2385 vdd.n1284 gnd 0.005579f
C2386 vdd.n1285 gnd 0.005579f
C2387 vdd.n1286 gnd 0.005579f
C2388 vdd.n1287 gnd 0.005579f
C2389 vdd.n1288 gnd 0.005579f
C2390 vdd.n1289 gnd 0.005579f
C2391 vdd.n1290 gnd 0.005579f
C2392 vdd.n1291 gnd 0.005579f
C2393 vdd.n1292 gnd 0.005579f
C2394 vdd.n1293 gnd 0.005579f
C2395 vdd.n1294 gnd 0.005579f
C2396 vdd.n1295 gnd 0.005579f
C2397 vdd.n1296 gnd 0.005579f
C2398 vdd.n1297 gnd 0.005579f
C2399 vdd.n1298 gnd 0.005579f
C2400 vdd.n1299 gnd 0.005579f
C2401 vdd.n1300 gnd 0.005579f
C2402 vdd.n1301 gnd 0.005579f
C2403 vdd.n1302 gnd 0.005579f
C2404 vdd.n1303 gnd 0.005579f
C2405 vdd.n1304 gnd 0.005579f
C2406 vdd.n1305 gnd 0.03758f
C2407 vdd.n1307 gnd 0.020451f
C2408 vdd.n1308 gnd 0.006603f
C2409 vdd.n1310 gnd 0.008204f
C2410 vdd.n1311 gnd 0.006603f
C2411 vdd.n1312 gnd 0.008204f
C2412 vdd.n1314 gnd 0.008204f
C2413 vdd.n1315 gnd 0.008204f
C2414 vdd.n1317 gnd 0.008204f
C2415 vdd.n1318 gnd 0.00548f
C2416 vdd.t76 gnd 0.41919f
C2417 vdd.n1319 gnd 0.008204f
C2418 vdd.n1320 gnd 0.020451f
C2419 vdd.n1321 gnd 0.006603f
C2420 vdd.n1322 gnd 0.008204f
C2421 vdd.n1323 gnd 0.006603f
C2422 vdd.n1324 gnd 0.008204f
C2423 vdd.n1325 gnd 0.83838f
C2424 vdd.n1326 gnd 0.008204f
C2425 vdd.n1327 gnd 0.006603f
C2426 vdd.n1328 gnd 0.006603f
C2427 vdd.n1329 gnd 0.008204f
C2428 vdd.n1330 gnd 0.006603f
C2429 vdd.n1331 gnd 0.008204f
C2430 vdd.t170 gnd 0.41919f
C2431 vdd.n1332 gnd 0.008204f
C2432 vdd.n1333 gnd 0.006603f
C2433 vdd.n1334 gnd 0.008204f
C2434 vdd.n1335 gnd 0.006603f
C2435 vdd.n1336 gnd 0.008204f
C2436 vdd.t186 gnd 0.41919f
C2437 vdd.n1337 gnd 0.008204f
C2438 vdd.n1338 gnd 0.006603f
C2439 vdd.n1339 gnd 0.008204f
C2440 vdd.n1340 gnd 0.006603f
C2441 vdd.n1341 gnd 0.008204f
C2442 vdd.n1342 gnd 0.658129f
C2443 vdd.n1343 gnd 0.695856f
C2444 vdd.t188 gnd 0.41919f
C2445 vdd.n1344 gnd 0.008204f
C2446 vdd.n1345 gnd 0.006603f
C2447 vdd.n1346 gnd 0.004502f
C2448 vdd.n1347 gnd 0.004178f
C2449 vdd.n1348 gnd 0.002311f
C2450 vdd.n1349 gnd 0.005306f
C2451 vdd.n1350 gnd 0.002245f
C2452 vdd.n1351 gnd 0.002377f
C2453 vdd.n1352 gnd 0.004178f
C2454 vdd.n1353 gnd 0.002245f
C2455 vdd.n1354 gnd 0.005306f
C2456 vdd.n1355 gnd 0.002377f
C2457 vdd.n1356 gnd 0.004178f
C2458 vdd.n1357 gnd 0.002245f
C2459 vdd.n1358 gnd 0.00398f
C2460 vdd.n1359 gnd 0.003992f
C2461 vdd.t184 gnd 0.0114f
C2462 vdd.n1360 gnd 0.025366f
C2463 vdd.n1361 gnd 0.132009f
C2464 vdd.n1362 gnd 0.002245f
C2465 vdd.n1363 gnd 0.002377f
C2466 vdd.n1364 gnd 0.005306f
C2467 vdd.n1365 gnd 0.005306f
C2468 vdd.n1366 gnd 0.002377f
C2469 vdd.n1367 gnd 0.002245f
C2470 vdd.n1368 gnd 0.004178f
C2471 vdd.n1369 gnd 0.004178f
C2472 vdd.n1370 gnd 0.002245f
C2473 vdd.n1371 gnd 0.002377f
C2474 vdd.n1372 gnd 0.005306f
C2475 vdd.n1373 gnd 0.005306f
C2476 vdd.n1374 gnd 0.002377f
C2477 vdd.n1375 gnd 0.002245f
C2478 vdd.n1376 gnd 0.004178f
C2479 vdd.n1377 gnd 0.004178f
C2480 vdd.n1378 gnd 0.002245f
C2481 vdd.n1379 gnd 0.002377f
C2482 vdd.n1380 gnd 0.005306f
C2483 vdd.n1381 gnd 0.005306f
C2484 vdd.n1382 gnd 0.012545f
C2485 vdd.n1383 gnd 0.002311f
C2486 vdd.n1384 gnd 0.002245f
C2487 vdd.n1385 gnd 0.010799f
C2488 vdd.n1386 gnd 0.007539f
C2489 vdd.t205 gnd 0.026412f
C2490 vdd.t211 gnd 0.026412f
C2491 vdd.n1387 gnd 0.181521f
C2492 vdd.n1388 gnd 0.142739f
C2493 vdd.t197 gnd 0.026412f
C2494 vdd.t160 gnd 0.026412f
C2495 vdd.n1389 gnd 0.181521f
C2496 vdd.n1390 gnd 0.115189f
C2497 vdd.t190 gnd 0.026412f
C2498 vdd.t169 gnd 0.026412f
C2499 vdd.n1391 gnd 0.181521f
C2500 vdd.n1392 gnd 0.115189f
C2501 vdd.n1393 gnd 0.004502f
C2502 vdd.n1394 gnd 0.004178f
C2503 vdd.n1395 gnd 0.002311f
C2504 vdd.n1396 gnd 0.005306f
C2505 vdd.n1397 gnd 0.002245f
C2506 vdd.n1398 gnd 0.002377f
C2507 vdd.n1399 gnd 0.004178f
C2508 vdd.n1400 gnd 0.002245f
C2509 vdd.n1401 gnd 0.005306f
C2510 vdd.n1402 gnd 0.002377f
C2511 vdd.n1403 gnd 0.004178f
C2512 vdd.n1404 gnd 0.002245f
C2513 vdd.n1405 gnd 0.00398f
C2514 vdd.n1406 gnd 0.003992f
C2515 vdd.t179 gnd 0.0114f
C2516 vdd.n1407 gnd 0.025366f
C2517 vdd.n1408 gnd 0.132009f
C2518 vdd.n1409 gnd 0.002245f
C2519 vdd.n1410 gnd 0.002377f
C2520 vdd.n1411 gnd 0.005306f
C2521 vdd.n1412 gnd 0.005306f
C2522 vdd.n1413 gnd 0.002377f
C2523 vdd.n1414 gnd 0.002245f
C2524 vdd.n1415 gnd 0.004178f
C2525 vdd.n1416 gnd 0.004178f
C2526 vdd.n1417 gnd 0.002245f
C2527 vdd.n1418 gnd 0.002377f
C2528 vdd.n1419 gnd 0.005306f
C2529 vdd.n1420 gnd 0.005306f
C2530 vdd.n1421 gnd 0.002377f
C2531 vdd.n1422 gnd 0.002245f
C2532 vdd.n1423 gnd 0.004178f
C2533 vdd.n1424 gnd 0.004178f
C2534 vdd.n1425 gnd 0.002245f
C2535 vdd.n1426 gnd 0.002377f
C2536 vdd.n1427 gnd 0.005306f
C2537 vdd.n1428 gnd 0.005306f
C2538 vdd.n1429 gnd 0.012545f
C2539 vdd.n1430 gnd 0.002311f
C2540 vdd.n1431 gnd 0.002245f
C2541 vdd.n1432 gnd 0.010799f
C2542 vdd.n1433 gnd 0.007302f
C2543 vdd.n1434 gnd 0.085702f
C2544 vdd.n1435 gnd 0.004502f
C2545 vdd.n1436 gnd 0.004178f
C2546 vdd.n1437 gnd 0.002311f
C2547 vdd.n1438 gnd 0.005306f
C2548 vdd.n1439 gnd 0.002245f
C2549 vdd.n1440 gnd 0.002377f
C2550 vdd.n1441 gnd 0.004178f
C2551 vdd.n1442 gnd 0.002245f
C2552 vdd.n1443 gnd 0.005306f
C2553 vdd.n1444 gnd 0.002377f
C2554 vdd.n1445 gnd 0.004178f
C2555 vdd.n1446 gnd 0.002245f
C2556 vdd.n1447 gnd 0.00398f
C2557 vdd.n1448 gnd 0.003992f
C2558 vdd.t171 gnd 0.0114f
C2559 vdd.n1449 gnd 0.025366f
C2560 vdd.n1450 gnd 0.132009f
C2561 vdd.n1451 gnd 0.002245f
C2562 vdd.n1452 gnd 0.002377f
C2563 vdd.n1453 gnd 0.005306f
C2564 vdd.n1454 gnd 0.005306f
C2565 vdd.n1455 gnd 0.002377f
C2566 vdd.n1456 gnd 0.002245f
C2567 vdd.n1457 gnd 0.004178f
C2568 vdd.n1458 gnd 0.004178f
C2569 vdd.n1459 gnd 0.002245f
C2570 vdd.n1460 gnd 0.002377f
C2571 vdd.n1461 gnd 0.005306f
C2572 vdd.n1462 gnd 0.005306f
C2573 vdd.n1463 gnd 0.002377f
C2574 vdd.n1464 gnd 0.002245f
C2575 vdd.n1465 gnd 0.004178f
C2576 vdd.n1466 gnd 0.004178f
C2577 vdd.n1467 gnd 0.002245f
C2578 vdd.n1468 gnd 0.002377f
C2579 vdd.n1469 gnd 0.005306f
C2580 vdd.n1470 gnd 0.005306f
C2581 vdd.n1471 gnd 0.012545f
C2582 vdd.n1472 gnd 0.002311f
C2583 vdd.n1473 gnd 0.002245f
C2584 vdd.n1474 gnd 0.010799f
C2585 vdd.n1475 gnd 0.007539f
C2586 vdd.t189 gnd 0.026412f
C2587 vdd.t187 gnd 0.026412f
C2588 vdd.n1476 gnd 0.181521f
C2589 vdd.n1477 gnd 0.142739f
C2590 vdd.t167 gnd 0.026412f
C2591 vdd.t153 gnd 0.026412f
C2592 vdd.n1478 gnd 0.181521f
C2593 vdd.n1479 gnd 0.115189f
C2594 vdd.t149 gnd 0.026412f
C2595 vdd.t185 gnd 0.026412f
C2596 vdd.n1480 gnd 0.181521f
C2597 vdd.n1481 gnd 0.115189f
C2598 vdd.n1482 gnd 0.004502f
C2599 vdd.n1483 gnd 0.004178f
C2600 vdd.n1484 gnd 0.002311f
C2601 vdd.n1485 gnd 0.005306f
C2602 vdd.n1486 gnd 0.002245f
C2603 vdd.n1487 gnd 0.002377f
C2604 vdd.n1488 gnd 0.004178f
C2605 vdd.n1489 gnd 0.002245f
C2606 vdd.n1490 gnd 0.005306f
C2607 vdd.n1491 gnd 0.002377f
C2608 vdd.n1492 gnd 0.004178f
C2609 vdd.n1493 gnd 0.002245f
C2610 vdd.n1494 gnd 0.00398f
C2611 vdd.n1495 gnd 0.003992f
C2612 vdd.t151 gnd 0.0114f
C2613 vdd.n1496 gnd 0.025366f
C2614 vdd.n1497 gnd 0.132009f
C2615 vdd.n1498 gnd 0.002245f
C2616 vdd.n1499 gnd 0.002377f
C2617 vdd.n1500 gnd 0.005306f
C2618 vdd.n1501 gnd 0.005306f
C2619 vdd.n1502 gnd 0.002377f
C2620 vdd.n1503 gnd 0.002245f
C2621 vdd.n1504 gnd 0.004178f
C2622 vdd.n1505 gnd 0.004178f
C2623 vdd.n1506 gnd 0.002245f
C2624 vdd.n1507 gnd 0.002377f
C2625 vdd.n1508 gnd 0.005306f
C2626 vdd.n1509 gnd 0.005306f
C2627 vdd.n1510 gnd 0.002377f
C2628 vdd.n1511 gnd 0.002245f
C2629 vdd.n1512 gnd 0.004178f
C2630 vdd.n1513 gnd 0.004178f
C2631 vdd.n1514 gnd 0.002245f
C2632 vdd.n1515 gnd 0.002377f
C2633 vdd.n1516 gnd 0.005306f
C2634 vdd.n1517 gnd 0.005306f
C2635 vdd.n1518 gnd 0.012545f
C2636 vdd.n1519 gnd 0.002311f
C2637 vdd.n1520 gnd 0.002245f
C2638 vdd.n1521 gnd 0.010799f
C2639 vdd.n1522 gnd 0.007302f
C2640 vdd.n1523 gnd 0.050984f
C2641 vdd.n1524 gnd 0.183708f
C2642 vdd.n1525 gnd 0.004502f
C2643 vdd.n1526 gnd 0.004178f
C2644 vdd.n1527 gnd 0.002311f
C2645 vdd.n1528 gnd 0.005306f
C2646 vdd.n1529 gnd 0.002245f
C2647 vdd.n1530 gnd 0.002377f
C2648 vdd.n1531 gnd 0.004178f
C2649 vdd.n1532 gnd 0.002245f
C2650 vdd.n1533 gnd 0.005306f
C2651 vdd.n1534 gnd 0.002377f
C2652 vdd.n1535 gnd 0.004178f
C2653 vdd.n1536 gnd 0.002245f
C2654 vdd.n1537 gnd 0.00398f
C2655 vdd.n1538 gnd 0.003992f
C2656 vdd.t176 gnd 0.0114f
C2657 vdd.n1539 gnd 0.025366f
C2658 vdd.n1540 gnd 0.132009f
C2659 vdd.n1541 gnd 0.002245f
C2660 vdd.n1542 gnd 0.002377f
C2661 vdd.n1543 gnd 0.005306f
C2662 vdd.n1544 gnd 0.005306f
C2663 vdd.n1545 gnd 0.002377f
C2664 vdd.n1546 gnd 0.002245f
C2665 vdd.n1547 gnd 0.004178f
C2666 vdd.n1548 gnd 0.004178f
C2667 vdd.n1549 gnd 0.002245f
C2668 vdd.n1550 gnd 0.002377f
C2669 vdd.n1551 gnd 0.005306f
C2670 vdd.n1552 gnd 0.005306f
C2671 vdd.n1553 gnd 0.002377f
C2672 vdd.n1554 gnd 0.002245f
C2673 vdd.n1555 gnd 0.004178f
C2674 vdd.n1556 gnd 0.004178f
C2675 vdd.n1557 gnd 0.002245f
C2676 vdd.n1558 gnd 0.002377f
C2677 vdd.n1559 gnd 0.005306f
C2678 vdd.n1560 gnd 0.005306f
C2679 vdd.n1561 gnd 0.012545f
C2680 vdd.n1562 gnd 0.002311f
C2681 vdd.n1563 gnd 0.002245f
C2682 vdd.n1564 gnd 0.010799f
C2683 vdd.n1565 gnd 0.007539f
C2684 vdd.t194 gnd 0.026412f
C2685 vdd.t193 gnd 0.026412f
C2686 vdd.n1566 gnd 0.181521f
C2687 vdd.n1567 gnd 0.142739f
C2688 vdd.t175 gnd 0.026412f
C2689 vdd.t163 gnd 0.026412f
C2690 vdd.n1568 gnd 0.181521f
C2691 vdd.n1569 gnd 0.115189f
C2692 vdd.t161 gnd 0.026412f
C2693 vdd.t192 gnd 0.026412f
C2694 vdd.n1570 gnd 0.181521f
C2695 vdd.n1571 gnd 0.115189f
C2696 vdd.n1572 gnd 0.004502f
C2697 vdd.n1573 gnd 0.004178f
C2698 vdd.n1574 gnd 0.002311f
C2699 vdd.n1575 gnd 0.005306f
C2700 vdd.n1576 gnd 0.002245f
C2701 vdd.n1577 gnd 0.002377f
C2702 vdd.n1578 gnd 0.004178f
C2703 vdd.n1579 gnd 0.002245f
C2704 vdd.n1580 gnd 0.005306f
C2705 vdd.n1581 gnd 0.002377f
C2706 vdd.n1582 gnd 0.004178f
C2707 vdd.n1583 gnd 0.002245f
C2708 vdd.n1584 gnd 0.00398f
C2709 vdd.n1585 gnd 0.003992f
C2710 vdd.t162 gnd 0.0114f
C2711 vdd.n1586 gnd 0.025366f
C2712 vdd.n1587 gnd 0.132009f
C2713 vdd.n1588 gnd 0.002245f
C2714 vdd.n1589 gnd 0.002377f
C2715 vdd.n1590 gnd 0.005306f
C2716 vdd.n1591 gnd 0.005306f
C2717 vdd.n1592 gnd 0.002377f
C2718 vdd.n1593 gnd 0.002245f
C2719 vdd.n1594 gnd 0.004178f
C2720 vdd.n1595 gnd 0.004178f
C2721 vdd.n1596 gnd 0.002245f
C2722 vdd.n1597 gnd 0.002377f
C2723 vdd.n1598 gnd 0.005306f
C2724 vdd.n1599 gnd 0.005306f
C2725 vdd.n1600 gnd 0.002377f
C2726 vdd.n1601 gnd 0.002245f
C2727 vdd.n1602 gnd 0.004178f
C2728 vdd.n1603 gnd 0.004178f
C2729 vdd.n1604 gnd 0.002245f
C2730 vdd.n1605 gnd 0.002377f
C2731 vdd.n1606 gnd 0.005306f
C2732 vdd.n1607 gnd 0.005306f
C2733 vdd.n1608 gnd 0.012545f
C2734 vdd.n1609 gnd 0.002311f
C2735 vdd.n1610 gnd 0.002245f
C2736 vdd.n1611 gnd 0.010799f
C2737 vdd.n1612 gnd 0.007302f
C2738 vdd.n1613 gnd 0.050984f
C2739 vdd.n1614 gnd 0.198842f
C2740 vdd.n1615 gnd 1.96832f
C2741 vdd.n1616 gnd 0.483886f
C2742 vdd.n1617 gnd 0.006603f
C2743 vdd.n1618 gnd 0.008204f
C2744 vdd.n1619 gnd 0.515604f
C2745 vdd.n1620 gnd 0.008204f
C2746 vdd.n1621 gnd 0.006603f
C2747 vdd.n1622 gnd 0.008204f
C2748 vdd.n1623 gnd 0.006603f
C2749 vdd.n1624 gnd 0.008204f
C2750 vdd.t168 gnd 0.41919f
C2751 vdd.t166 gnd 0.41919f
C2752 vdd.n1625 gnd 0.008204f
C2753 vdd.n1626 gnd 0.006603f
C2754 vdd.n1627 gnd 0.008204f
C2755 vdd.n1628 gnd 0.006603f
C2756 vdd.n1629 gnd 0.008204f
C2757 vdd.t148 gnd 0.41919f
C2758 vdd.n1630 gnd 0.008204f
C2759 vdd.n1631 gnd 0.006603f
C2760 vdd.n1632 gnd 0.008204f
C2761 vdd.n1633 gnd 0.006603f
C2762 vdd.n1634 gnd 0.008204f
C2763 vdd.t150 gnd 0.41919f
C2764 vdd.n1635 gnd 0.607826f
C2765 vdd.n1636 gnd 0.008204f
C2766 vdd.n1637 gnd 0.006603f
C2767 vdd.n1638 gnd 0.008204f
C2768 vdd.n1639 gnd 0.006603f
C2769 vdd.n1640 gnd 0.008204f
C2770 vdd.n1641 gnd 0.83838f
C2771 vdd.n1642 gnd 0.008204f
C2772 vdd.n1643 gnd 0.006603f
C2773 vdd.n1644 gnd 0.019993f
C2774 vdd.n1645 gnd 0.00548f
C2775 vdd.n1646 gnd 0.019993f
C2776 vdd.t94 gnd 0.41919f
C2777 vdd.n1647 gnd 0.019993f
C2778 vdd.n1648 gnd 0.00548f
C2779 vdd.n1649 gnd 0.008204f
C2780 vdd.n1650 gnd 0.006603f
C2781 vdd.n1651 gnd 0.008204f
C2782 vdd.n1682 gnd 0.020451f
C2783 vdd.n1683 gnd 1.23661f
C2784 vdd.n1684 gnd 0.008204f
C2785 vdd.n1685 gnd 0.006603f
C2786 vdd.n1686 gnd 0.008204f
C2787 vdd.n1687 gnd 0.008204f
C2788 vdd.n1688 gnd 0.008204f
C2789 vdd.n1689 gnd 0.008204f
C2790 vdd.n1690 gnd 0.008204f
C2791 vdd.n1691 gnd 0.006603f
C2792 vdd.n1692 gnd 0.008204f
C2793 vdd.n1693 gnd 0.008204f
C2794 vdd.n1694 gnd 0.008204f
C2795 vdd.n1695 gnd 0.008204f
C2796 vdd.n1696 gnd 0.008204f
C2797 vdd.n1697 gnd 0.006603f
C2798 vdd.n1698 gnd 0.008204f
C2799 vdd.n1699 gnd 0.008204f
C2800 vdd.n1700 gnd 0.008204f
C2801 vdd.n1701 gnd 0.008204f
C2802 vdd.n1702 gnd 0.008204f
C2803 vdd.n1703 gnd 0.006603f
C2804 vdd.n1704 gnd 0.008204f
C2805 vdd.n1705 gnd 0.008204f
C2806 vdd.n1706 gnd 0.008204f
C2807 vdd.n1707 gnd 0.008204f
C2808 vdd.n1708 gnd 0.008204f
C2809 vdd.t108 gnd 0.100927f
C2810 vdd.t109 gnd 0.107863f
C2811 vdd.t107 gnd 0.13181f
C2812 vdd.n1709 gnd 0.168961f
C2813 vdd.n1710 gnd 0.142618f
C2814 vdd.n1711 gnd 0.01413f
C2815 vdd.n1712 gnd 0.008204f
C2816 vdd.n1713 gnd 0.008204f
C2817 vdd.n1714 gnd 0.008204f
C2818 vdd.n1715 gnd 0.008204f
C2819 vdd.n1716 gnd 0.008204f
C2820 vdd.n1717 gnd 0.006603f
C2821 vdd.n1718 gnd 0.008204f
C2822 vdd.n1719 gnd 0.008204f
C2823 vdd.n1720 gnd 0.008204f
C2824 vdd.n1721 gnd 0.008204f
C2825 vdd.n1722 gnd 0.008204f
C2826 vdd.n1723 gnd 0.006603f
C2827 vdd.n1724 gnd 0.008204f
C2828 vdd.n1725 gnd 0.008204f
C2829 vdd.n1726 gnd 0.008204f
C2830 vdd.n1727 gnd 0.008204f
C2831 vdd.n1728 gnd 0.008204f
C2832 vdd.n1729 gnd 0.006603f
C2833 vdd.n1730 gnd 0.008204f
C2834 vdd.n1731 gnd 0.008204f
C2835 vdd.n1732 gnd 0.008204f
C2836 vdd.n1733 gnd 0.008204f
C2837 vdd.n1734 gnd 0.008204f
C2838 vdd.n1735 gnd 0.006603f
C2839 vdd.n1736 gnd 0.008204f
C2840 vdd.n1737 gnd 0.008204f
C2841 vdd.n1738 gnd 0.008204f
C2842 vdd.n1739 gnd 0.008204f
C2843 vdd.n1740 gnd 0.008204f
C2844 vdd.n1741 gnd 0.006603f
C2845 vdd.n1742 gnd 0.008204f
C2846 vdd.n1743 gnd 0.008204f
C2847 vdd.n1744 gnd 0.008204f
C2848 vdd.n1745 gnd 0.008204f
C2849 vdd.n1746 gnd 0.006603f
C2850 vdd.n1747 gnd 0.008204f
C2851 vdd.n1748 gnd 0.008204f
C2852 vdd.n1749 gnd 0.008204f
C2853 vdd.n1750 gnd 0.008204f
C2854 vdd.n1751 gnd 0.008204f
C2855 vdd.n1752 gnd 0.006603f
C2856 vdd.n1753 gnd 0.008204f
C2857 vdd.n1754 gnd 0.008204f
C2858 vdd.n1755 gnd 0.008204f
C2859 vdd.n1756 gnd 0.008204f
C2860 vdd.n1757 gnd 0.008204f
C2861 vdd.n1758 gnd 0.006603f
C2862 vdd.n1759 gnd 0.008204f
C2863 vdd.n1760 gnd 0.008204f
C2864 vdd.n1761 gnd 0.008204f
C2865 vdd.n1762 gnd 0.008204f
C2866 vdd.n1763 gnd 0.008204f
C2867 vdd.n1764 gnd 0.006603f
C2868 vdd.n1765 gnd 0.008204f
C2869 vdd.n1766 gnd 0.008204f
C2870 vdd.n1767 gnd 0.008204f
C2871 vdd.n1768 gnd 0.008204f
C2872 vdd.n1769 gnd 0.008204f
C2873 vdd.n1770 gnd 0.006603f
C2874 vdd.n1771 gnd 0.008204f
C2875 vdd.n1772 gnd 0.008204f
C2876 vdd.n1773 gnd 0.008204f
C2877 vdd.n1774 gnd 0.008204f
C2878 vdd.t105 gnd 0.100927f
C2879 vdd.t106 gnd 0.107863f
C2880 vdd.t104 gnd 0.13181f
C2881 vdd.n1775 gnd 0.168961f
C2882 vdd.n1776 gnd 0.142618f
C2883 vdd.n1777 gnd 0.010829f
C2884 vdd.n1778 gnd 0.003136f
C2885 vdd.n1779 gnd 0.020451f
C2886 vdd.n1780 gnd 0.008204f
C2887 vdd.n1781 gnd 0.003467f
C2888 vdd.n1782 gnd 0.006603f
C2889 vdd.n1783 gnd 0.006603f
C2890 vdd.n1784 gnd 0.008204f
C2891 vdd.n1785 gnd 0.008204f
C2892 vdd.n1786 gnd 0.008204f
C2893 vdd.n1787 gnd 0.006603f
C2894 vdd.n1788 gnd 0.006603f
C2895 vdd.n1789 gnd 0.006603f
C2896 vdd.n1790 gnd 0.008204f
C2897 vdd.n1791 gnd 0.008204f
C2898 vdd.n1792 gnd 0.008204f
C2899 vdd.n1793 gnd 0.006603f
C2900 vdd.n1794 gnd 0.006603f
C2901 vdd.n1795 gnd 0.006603f
C2902 vdd.n1796 gnd 0.008204f
C2903 vdd.n1797 gnd 0.008204f
C2904 vdd.n1798 gnd 0.008204f
C2905 vdd.n1799 gnd 0.006603f
C2906 vdd.n1800 gnd 0.006603f
C2907 vdd.n1801 gnd 0.006603f
C2908 vdd.n1802 gnd 0.008204f
C2909 vdd.n1803 gnd 0.008204f
C2910 vdd.n1804 gnd 0.008204f
C2911 vdd.n1805 gnd 0.006603f
C2912 vdd.n1806 gnd 0.006603f
C2913 vdd.n1807 gnd 0.006603f
C2914 vdd.n1808 gnd 0.008204f
C2915 vdd.n1809 gnd 0.008204f
C2916 vdd.n1810 gnd 0.008204f
C2917 vdd.n1811 gnd 0.006537f
C2918 vdd.n1812 gnd 0.008204f
C2919 vdd.t95 gnd 0.100927f
C2920 vdd.t96 gnd 0.107863f
C2921 vdd.t93 gnd 0.13181f
C2922 vdd.n1813 gnd 0.168961f
C2923 vdd.n1814 gnd 0.142618f
C2924 vdd.n1815 gnd 0.01413f
C2925 vdd.n1816 gnd 0.00449f
C2926 vdd.n1817 gnd 0.008204f
C2927 vdd.n1818 gnd 0.008204f
C2928 vdd.n1819 gnd 0.008204f
C2929 vdd.n1820 gnd 0.006603f
C2930 vdd.n1821 gnd 0.006603f
C2931 vdd.n1822 gnd 0.006603f
C2932 vdd.n1823 gnd 0.008204f
C2933 vdd.n1824 gnd 0.008204f
C2934 vdd.n1825 gnd 0.008204f
C2935 vdd.n1826 gnd 0.006603f
C2936 vdd.n1827 gnd 0.006603f
C2937 vdd.n1828 gnd 0.006603f
C2938 vdd.n1829 gnd 0.008204f
C2939 vdd.n1830 gnd 0.008204f
C2940 vdd.n1831 gnd 0.008204f
C2941 vdd.n1832 gnd 0.006603f
C2942 vdd.n1833 gnd 0.006603f
C2943 vdd.n1834 gnd 0.006603f
C2944 vdd.n1835 gnd 0.008204f
C2945 vdd.n1836 gnd 0.008204f
C2946 vdd.n1837 gnd 0.008204f
C2947 vdd.n1838 gnd 0.006603f
C2948 vdd.n1839 gnd 0.006603f
C2949 vdd.n1840 gnd 0.006603f
C2950 vdd.n1841 gnd 0.008204f
C2951 vdd.n1842 gnd 0.008204f
C2952 vdd.n1843 gnd 0.008204f
C2953 vdd.n1844 gnd 0.006603f
C2954 vdd.n1845 gnd 0.006603f
C2955 vdd.n1846 gnd 0.005514f
C2956 vdd.n1847 gnd 0.008204f
C2957 vdd.n1848 gnd 0.008204f
C2958 vdd.n1849 gnd 0.008204f
C2959 vdd.n1850 gnd 0.005514f
C2960 vdd.n1851 gnd 0.006603f
C2961 vdd.n1852 gnd 0.006603f
C2962 vdd.n1853 gnd 0.008204f
C2963 vdd.n1854 gnd 0.008204f
C2964 vdd.n1855 gnd 0.008204f
C2965 vdd.n1856 gnd 0.006603f
C2966 vdd.n1857 gnd 0.006603f
C2967 vdd.n1858 gnd 0.006603f
C2968 vdd.n1859 gnd 0.008204f
C2969 vdd.n1860 gnd 0.008204f
C2970 vdd.n1861 gnd 0.008204f
C2971 vdd.n1862 gnd 0.006603f
C2972 vdd.n1863 gnd 0.006603f
C2973 vdd.n1864 gnd 0.006603f
C2974 vdd.n1865 gnd 0.008204f
C2975 vdd.n1866 gnd 0.008204f
C2976 vdd.n1867 gnd 0.008204f
C2977 vdd.n1868 gnd 0.006603f
C2978 vdd.n1869 gnd 0.006603f
C2979 vdd.n1870 gnd 0.006603f
C2980 vdd.n1871 gnd 0.008204f
C2981 vdd.n1872 gnd 0.008204f
C2982 vdd.n1873 gnd 0.008204f
C2983 vdd.n1874 gnd 0.006603f
C2984 vdd.n1875 gnd 0.008204f
C2985 vdd.n1876 gnd 2.00373f
C2986 vdd.n1878 gnd 0.020451f
C2987 vdd.n1879 gnd 0.00548f
C2988 vdd.n1880 gnd 0.020451f
C2989 vdd.n1881 gnd 0.019993f
C2990 vdd.n1882 gnd 0.008204f
C2991 vdd.n1883 gnd 0.006603f
C2992 vdd.n1884 gnd 0.008204f
C2993 vdd.n1885 gnd 0.44015f
C2994 vdd.n1886 gnd 0.008204f
C2995 vdd.n1887 gnd 0.006603f
C2996 vdd.n1888 gnd 0.008204f
C2997 vdd.n1889 gnd 0.008204f
C2998 vdd.n1890 gnd 0.008204f
C2999 vdd.n1891 gnd 0.006603f
C3000 vdd.n1892 gnd 0.008204f
C3001 vdd.n1893 gnd 0.75035f
C3002 vdd.n1894 gnd 0.83838f
C3003 vdd.n1895 gnd 0.008204f
C3004 vdd.n1896 gnd 0.006603f
C3005 vdd.n1897 gnd 0.008204f
C3006 vdd.n1898 gnd 0.008204f
C3007 vdd.n1899 gnd 0.008204f
C3008 vdd.n1900 gnd 0.006603f
C3009 vdd.n1901 gnd 0.008204f
C3010 vdd.n1902 gnd 0.50722f
C3011 vdd.n1903 gnd 0.008204f
C3012 vdd.n1904 gnd 0.006603f
C3013 vdd.n1905 gnd 0.008204f
C3014 vdd.n1906 gnd 0.008204f
C3015 vdd.n1907 gnd 0.008204f
C3016 vdd.n1908 gnd 0.006603f
C3017 vdd.n1909 gnd 0.008204f
C3018 vdd.n1910 gnd 0.465301f
C3019 vdd.n1911 gnd 0.649745f
C3020 vdd.n1912 gnd 0.008204f
C3021 vdd.n1913 gnd 0.006603f
C3022 vdd.n1914 gnd 0.008204f
C3023 vdd.n1915 gnd 0.008204f
C3024 vdd.n1916 gnd 0.006305f
C3025 vdd.n1917 gnd 0.008204f
C3026 vdd.n1918 gnd 0.006603f
C3027 vdd.n1919 gnd 0.008204f
C3028 vdd.n1920 gnd 0.695856f
C3029 vdd.n1921 gnd 0.008204f
C3030 vdd.n1922 gnd 0.006603f
C3031 vdd.n1923 gnd 0.008204f
C3032 vdd.n1924 gnd 0.008204f
C3033 vdd.n1925 gnd 0.008204f
C3034 vdd.n1926 gnd 0.006603f
C3035 vdd.n1927 gnd 0.008204f
C3036 vdd.t152 gnd 0.41919f
C3037 vdd.n1928 gnd 0.599442f
C3038 vdd.n1929 gnd 0.008204f
C3039 vdd.n1930 gnd 0.006603f
C3040 vdd.n1931 gnd 0.006305f
C3041 vdd.n1932 gnd 0.008204f
C3042 vdd.n1933 gnd 0.008204f
C3043 vdd.n1934 gnd 0.006603f
C3044 vdd.n1935 gnd 0.008204f
C3045 vdd.n1936 gnd 0.456917f
C3046 vdd.n1937 gnd 0.008204f
C3047 vdd.n1938 gnd 0.006603f
C3048 vdd.n1939 gnd 0.008204f
C3049 vdd.n1940 gnd 0.008204f
C3050 vdd.n1941 gnd 0.008204f
C3051 vdd.n1942 gnd 0.006603f
C3052 vdd.n1943 gnd 0.008204f
C3053 vdd.n1944 gnd 0.591058f
C3054 vdd.n1945 gnd 0.523988f
C3055 vdd.n1946 gnd 0.008204f
C3056 vdd.n1947 gnd 0.006603f
C3057 vdd.n1948 gnd 0.008204f
C3058 vdd.n1949 gnd 0.008204f
C3059 vdd.n1950 gnd 0.008204f
C3060 vdd.n1951 gnd 0.006603f
C3061 vdd.n1952 gnd 0.008204f
C3062 vdd.n1953 gnd 0.666512f
C3063 vdd.n1954 gnd 0.008204f
C3064 vdd.n1955 gnd 0.006603f
C3065 vdd.n1956 gnd 0.008204f
C3066 vdd.n1957 gnd 0.008204f
C3067 vdd.n1958 gnd 0.019993f
C3068 vdd.n1959 gnd 0.008204f
C3069 vdd.n1960 gnd 0.008204f
C3070 vdd.n1961 gnd 0.006603f
C3071 vdd.n1962 gnd 0.008204f
C3072 vdd.n1963 gnd 0.523988f
C3073 vdd.n1964 gnd 0.83838f
C3074 vdd.n1965 gnd 0.008204f
C3075 vdd.n1966 gnd 0.006603f
C3076 vdd.n1967 gnd 0.008204f
C3077 vdd.n1968 gnd 0.008204f
C3078 vdd.n1969 gnd 0.019993f
C3079 vdd.n1970 gnd 0.00548f
C3080 vdd.n1971 gnd 0.019993f
C3081 vdd.n1972 gnd 1.15277f
C3082 vdd.n1973 gnd 0.019993f
C3083 vdd.n1974 gnd 0.020451f
C3084 vdd.n1975 gnd 0.003136f
C3085 vdd.t99 gnd 0.100927f
C3086 vdd.t98 gnd 0.107863f
C3087 vdd.t97 gnd 0.13181f
C3088 vdd.n1976 gnd 0.168961f
C3089 vdd.n1977 gnd 0.141958f
C3090 vdd.n1978 gnd 0.010169f
C3091 vdd.n1979 gnd 0.003467f
C3092 vdd.n1980 gnd 0.007055f
C3093 vdd.n1981 gnd 0.870908f
C3094 vdd.n1983 gnd 0.006603f
C3095 vdd.n1984 gnd 0.006603f
C3096 vdd.n1985 gnd 0.008204f
C3097 vdd.n1987 gnd 0.008204f
C3098 vdd.n1988 gnd 0.008204f
C3099 vdd.n1989 gnd 0.006603f
C3100 vdd.n1990 gnd 0.006603f
C3101 vdd.n1991 gnd 0.006603f
C3102 vdd.n1992 gnd 0.008204f
C3103 vdd.n1994 gnd 0.008204f
C3104 vdd.n1995 gnd 0.008204f
C3105 vdd.n1996 gnd 0.006603f
C3106 vdd.n1997 gnd 0.006603f
C3107 vdd.n1998 gnd 0.006603f
C3108 vdd.n1999 gnd 0.008204f
C3109 vdd.n2001 gnd 0.008204f
C3110 vdd.n2002 gnd 0.008204f
C3111 vdd.n2003 gnd 0.006603f
C3112 vdd.n2004 gnd 0.006603f
C3113 vdd.n2005 gnd 0.006603f
C3114 vdd.n2006 gnd 0.008204f
C3115 vdd.n2008 gnd 0.008204f
C3116 vdd.n2009 gnd 0.008204f
C3117 vdd.n2010 gnd 0.006603f
C3118 vdd.n2011 gnd 0.008204f
C3119 vdd.n2012 gnd 0.008204f
C3120 vdd.n2013 gnd 0.008204f
C3121 vdd.n2014 gnd 0.01347f
C3122 vdd.n2015 gnd 0.00449f
C3123 vdd.n2016 gnd 0.006603f
C3124 vdd.n2017 gnd 0.008204f
C3125 vdd.n2019 gnd 0.008204f
C3126 vdd.n2020 gnd 0.008204f
C3127 vdd.n2021 gnd 0.006603f
C3128 vdd.n2022 gnd 0.006603f
C3129 vdd.n2023 gnd 0.006603f
C3130 vdd.n2024 gnd 0.008204f
C3131 vdd.n2026 gnd 0.008204f
C3132 vdd.n2027 gnd 0.008204f
C3133 vdd.n2028 gnd 0.006603f
C3134 vdd.n2029 gnd 0.006603f
C3135 vdd.n2030 gnd 0.006603f
C3136 vdd.n2031 gnd 0.008204f
C3137 vdd.n2033 gnd 0.008204f
C3138 vdd.n2034 gnd 0.008204f
C3139 vdd.n2035 gnd 0.006603f
C3140 vdd.n2036 gnd 0.006603f
C3141 vdd.n2037 gnd 0.006603f
C3142 vdd.n2038 gnd 0.008204f
C3143 vdd.n2040 gnd 0.008204f
C3144 vdd.n2041 gnd 0.008204f
C3145 vdd.n2042 gnd 0.006603f
C3146 vdd.n2043 gnd 0.006603f
C3147 vdd.n2044 gnd 0.006603f
C3148 vdd.n2045 gnd 0.008204f
C3149 vdd.n2047 gnd 0.008204f
C3150 vdd.n2048 gnd 0.008204f
C3151 vdd.n2049 gnd 0.006603f
C3152 vdd.n2050 gnd 0.008204f
C3153 vdd.n2051 gnd 0.008204f
C3154 vdd.n2052 gnd 0.008204f
C3155 vdd.n2053 gnd 0.01347f
C3156 vdd.n2054 gnd 0.005514f
C3157 vdd.n2055 gnd 0.006603f
C3158 vdd.n2056 gnd 0.008204f
C3159 vdd.n2058 gnd 0.008204f
C3160 vdd.n2059 gnd 0.008204f
C3161 vdd.n2060 gnd 0.006603f
C3162 vdd.n2061 gnd 0.006603f
C3163 vdd.n2062 gnd 0.006603f
C3164 vdd.n2063 gnd 0.008204f
C3165 vdd.n2065 gnd 0.008204f
C3166 vdd.n2066 gnd 0.008204f
C3167 vdd.n2067 gnd 0.006603f
C3168 vdd.n2068 gnd 0.006603f
C3169 vdd.n2069 gnd 0.006603f
C3170 vdd.n2070 gnd 0.008204f
C3171 vdd.n2072 gnd 0.008204f
C3172 vdd.n2073 gnd 0.008204f
C3173 vdd.n2074 gnd 0.006603f
C3174 vdd.n2075 gnd 0.006603f
C3175 vdd.n2076 gnd 0.006603f
C3176 vdd.n2077 gnd 0.008204f
C3177 vdd.n2079 gnd 0.008204f
C3178 vdd.n2080 gnd 0.006603f
C3179 vdd.n2081 gnd 0.006603f
C3180 vdd.n2082 gnd 0.008204f
C3181 vdd.n2084 gnd 0.008204f
C3182 vdd.n2085 gnd 0.008204f
C3183 vdd.n2086 gnd 0.006603f
C3184 vdd.n2087 gnd 0.007055f
C3185 vdd.n2088 gnd 0.870908f
C3186 vdd.n2089 gnd 0.03758f
C3187 vdd.n2090 gnd 0.005579f
C3188 vdd.n2091 gnd 0.005579f
C3189 vdd.n2092 gnd 0.005579f
C3190 vdd.n2093 gnd 0.005579f
C3191 vdd.n2094 gnd 0.005579f
C3192 vdd.n2095 gnd 0.005579f
C3193 vdd.n2096 gnd 0.005579f
C3194 vdd.n2097 gnd 0.005579f
C3195 vdd.n2098 gnd 0.005579f
C3196 vdd.n2099 gnd 0.005579f
C3197 vdd.n2100 gnd 0.005579f
C3198 vdd.n2101 gnd 0.005579f
C3199 vdd.n2102 gnd 0.005579f
C3200 vdd.n2103 gnd 0.005579f
C3201 vdd.n2104 gnd 0.005579f
C3202 vdd.n2105 gnd 0.005579f
C3203 vdd.n2106 gnd 0.005579f
C3204 vdd.n2107 gnd 0.005579f
C3205 vdd.n2108 gnd 0.005579f
C3206 vdd.n2109 gnd 0.005579f
C3207 vdd.n2110 gnd 0.005579f
C3208 vdd.n2111 gnd 0.005579f
C3209 vdd.n2112 gnd 0.005579f
C3210 vdd.n2113 gnd 0.005579f
C3211 vdd.n2114 gnd 0.005579f
C3212 vdd.n2115 gnd 0.005579f
C3213 vdd.n2116 gnd 0.005579f
C3214 vdd.n2117 gnd 0.005579f
C3215 vdd.n2118 gnd 0.005579f
C3216 vdd.n2119 gnd 0.005579f
C3217 vdd.n2120 gnd 9.90127f
C3218 vdd.n2122 gnd 0.012667f
C3219 vdd.n2123 gnd 0.012667f
C3220 vdd.n2124 gnd 0.011945f
C3221 vdd.n2125 gnd 0.005579f
C3222 vdd.n2126 gnd 0.005579f
C3223 vdd.n2127 gnd 0.570099f
C3224 vdd.n2128 gnd 0.005579f
C3225 vdd.n2129 gnd 0.005579f
C3226 vdd.n2130 gnd 0.005579f
C3227 vdd.n2131 gnd 0.005579f
C3228 vdd.n2132 gnd 0.005579f
C3229 vdd.n2133 gnd 0.448533f
C3230 vdd.n2134 gnd 0.005579f
C3231 vdd.n2135 gnd 0.005579f
C3232 vdd.n2136 gnd 0.005579f
C3233 vdd.n2137 gnd 0.005579f
C3234 vdd.n2138 gnd 0.005579f
C3235 vdd.n2139 gnd 0.570099f
C3236 vdd.n2140 gnd 0.005579f
C3237 vdd.n2141 gnd 0.005579f
C3238 vdd.n2142 gnd 0.005579f
C3239 vdd.n2143 gnd 0.005579f
C3240 vdd.n2144 gnd 0.005579f
C3241 vdd.n2145 gnd 0.570099f
C3242 vdd.n2146 gnd 0.005579f
C3243 vdd.n2147 gnd 0.005579f
C3244 vdd.n2148 gnd 0.005579f
C3245 vdd.n2149 gnd 0.005579f
C3246 vdd.n2150 gnd 0.005579f
C3247 vdd.n2151 gnd 0.549139f
C3248 vdd.n2152 gnd 0.005579f
C3249 vdd.n2153 gnd 0.005579f
C3250 vdd.n2154 gnd 0.005579f
C3251 vdd.n2155 gnd 0.005579f
C3252 vdd.n2156 gnd 0.005579f
C3253 vdd.n2157 gnd 0.423382f
C3254 vdd.n2158 gnd 0.005579f
C3255 vdd.n2159 gnd 0.005579f
C3256 vdd.n2160 gnd 0.005579f
C3257 vdd.n2161 gnd 0.005579f
C3258 vdd.n2162 gnd 0.005579f
C3259 vdd.n2163 gnd 0.297625f
C3260 vdd.n2164 gnd 0.005579f
C3261 vdd.n2165 gnd 0.005579f
C3262 vdd.n2166 gnd 0.005579f
C3263 vdd.n2167 gnd 0.005579f
C3264 vdd.n2168 gnd 0.005579f
C3265 vdd.n2169 gnd 0.398231f
C3266 vdd.n2170 gnd 0.005579f
C3267 vdd.n2171 gnd 0.005579f
C3268 vdd.n2172 gnd 0.005579f
C3269 vdd.n2173 gnd 0.005579f
C3270 vdd.n2174 gnd 0.005579f
C3271 vdd.n2175 gnd 0.523988f
C3272 vdd.n2176 gnd 0.005579f
C3273 vdd.n2177 gnd 0.005579f
C3274 vdd.n2178 gnd 0.005579f
C3275 vdd.n2179 gnd 0.005579f
C3276 vdd.n2180 gnd 0.005579f
C3277 vdd.n2181 gnd 0.570099f
C3278 vdd.n2182 gnd 0.005579f
C3279 vdd.n2183 gnd 0.005579f
C3280 vdd.n2184 gnd 0.005579f
C3281 vdd.n2185 gnd 0.005579f
C3282 vdd.n2186 gnd 0.005579f
C3283 vdd.n2187 gnd 0.490452f
C3284 vdd.n2188 gnd 0.005579f
C3285 vdd.n2189 gnd 0.005579f
C3286 vdd.n2190 gnd 0.00443f
C3287 vdd.n2191 gnd 0.01616f
C3288 vdd.n2192 gnd 0.003938f
C3289 vdd.n2193 gnd 0.005579f
C3290 vdd.n2194 gnd 0.364695f
C3291 vdd.n2195 gnd 0.005579f
C3292 vdd.n2196 gnd 0.005579f
C3293 vdd.n2197 gnd 0.005579f
C3294 vdd.n2198 gnd 0.005579f
C3295 vdd.n2199 gnd 0.005579f
C3296 vdd.n2200 gnd 0.33116f
C3297 vdd.n2201 gnd 0.005579f
C3298 vdd.n2202 gnd 0.005579f
C3299 vdd.n2203 gnd 0.005579f
C3300 vdd.n2204 gnd 0.005579f
C3301 vdd.n2205 gnd 0.005579f
C3302 vdd.n2206 gnd 0.456917f
C3303 vdd.n2207 gnd 0.005579f
C3304 vdd.n2208 gnd 0.005579f
C3305 vdd.n2209 gnd 0.005579f
C3306 vdd.n2210 gnd 0.005579f
C3307 vdd.n2211 gnd 0.005579f
C3308 vdd.n2212 gnd 0.503028f
C3309 vdd.n2213 gnd 0.005579f
C3310 vdd.n2214 gnd 0.005579f
C3311 vdd.n2215 gnd 0.005579f
C3312 vdd.n2216 gnd 0.005579f
C3313 vdd.n2217 gnd 0.005579f
C3314 vdd.n2218 gnd 0.377271f
C3315 vdd.n2219 gnd 0.005579f
C3316 vdd.n2220 gnd 0.005579f
C3317 vdd.n2221 gnd 0.005579f
C3318 vdd.n2222 gnd 0.005579f
C3319 vdd.n2223 gnd 0.005579f
C3320 vdd.n2224 gnd 0.180252f
C3321 vdd.n2225 gnd 0.005579f
C3322 vdd.n2226 gnd 0.005579f
C3323 vdd.n2227 gnd 0.005579f
C3324 vdd.n2228 gnd 0.005579f
C3325 vdd.n2229 gnd 0.005579f
C3326 vdd.n2230 gnd 0.180252f
C3327 vdd.n2231 gnd 0.005579f
C3328 vdd.n2232 gnd 0.005579f
C3329 vdd.n2233 gnd 0.005579f
C3330 vdd.n2234 gnd 0.005579f
C3331 vdd.n2235 gnd 0.005579f
C3332 vdd.n2236 gnd 0.570099f
C3333 vdd.n2237 gnd 0.005579f
C3334 vdd.n2238 gnd 0.005579f
C3335 vdd.n2239 gnd 0.005579f
C3336 vdd.n2240 gnd 0.005579f
C3337 vdd.n2241 gnd 0.005579f
C3338 vdd.n2242 gnd 0.005579f
C3339 vdd.n2243 gnd 0.005579f
C3340 vdd.n2244 gnd 0.394039f
C3341 vdd.n2245 gnd 0.005579f
C3342 vdd.n2246 gnd 0.005579f
C3343 vdd.n2247 gnd 0.005579f
C3344 vdd.n2248 gnd 0.005579f
C3345 vdd.n2249 gnd 0.005579f
C3346 vdd.n2250 gnd 0.005579f
C3347 vdd.n2251 gnd 0.356312f
C3348 vdd.n2252 gnd 0.005579f
C3349 vdd.n2253 gnd 0.005579f
C3350 vdd.n2254 gnd 0.005579f
C3351 vdd.n2255 gnd 0.012667f
C3352 vdd.n2256 gnd 0.011945f
C3353 vdd.n2257 gnd 0.005579f
C3354 vdd.n2258 gnd 0.005579f
C3355 vdd.n2259 gnd 0.004307f
C3356 vdd.n2260 gnd 0.005579f
C3357 vdd.n2261 gnd 0.005579f
C3358 vdd.n2262 gnd 0.004061f
C3359 vdd.n2263 gnd 0.005579f
C3360 vdd.n2264 gnd 0.005579f
C3361 vdd.n2265 gnd 0.005579f
C3362 vdd.n2266 gnd 0.005579f
C3363 vdd.n2267 gnd 0.005579f
C3364 vdd.n2268 gnd 0.005579f
C3365 vdd.n2269 gnd 0.005579f
C3366 vdd.n2270 gnd 0.005579f
C3367 vdd.n2271 gnd 0.005579f
C3368 vdd.n2272 gnd 0.005579f
C3369 vdd.n2273 gnd 0.005579f
C3370 vdd.n2274 gnd 0.005579f
C3371 vdd.n2275 gnd 0.005579f
C3372 vdd.n2276 gnd 0.005579f
C3373 vdd.n2277 gnd 0.005579f
C3374 vdd.n2278 gnd 0.005579f
C3375 vdd.n2279 gnd 0.005579f
C3376 vdd.n2280 gnd 0.005579f
C3377 vdd.n2281 gnd 0.005579f
C3378 vdd.n2282 gnd 0.005579f
C3379 vdd.n2283 gnd 0.005579f
C3380 vdd.n2284 gnd 0.005579f
C3381 vdd.n2285 gnd 0.005579f
C3382 vdd.n2286 gnd 0.005579f
C3383 vdd.n2287 gnd 0.005579f
C3384 vdd.n2288 gnd 0.005579f
C3385 vdd.n2289 gnd 0.005579f
C3386 vdd.n2290 gnd 0.005579f
C3387 vdd.n2291 gnd 0.005579f
C3388 vdd.n2292 gnd 0.005579f
C3389 vdd.n2293 gnd 0.005579f
C3390 vdd.n2294 gnd 0.005579f
C3391 vdd.n2295 gnd 0.005579f
C3392 vdd.n2296 gnd 0.005579f
C3393 vdd.n2297 gnd 0.005579f
C3394 vdd.n2298 gnd 0.005579f
C3395 vdd.n2299 gnd 0.005579f
C3396 vdd.n2300 gnd 0.005579f
C3397 vdd.n2301 gnd 0.005579f
C3398 vdd.n2302 gnd 0.005579f
C3399 vdd.n2303 gnd 0.005579f
C3400 vdd.n2304 gnd 0.005579f
C3401 vdd.n2305 gnd 0.005579f
C3402 vdd.n2306 gnd 0.005579f
C3403 vdd.n2307 gnd 0.005579f
C3404 vdd.n2308 gnd 0.005579f
C3405 vdd.n2309 gnd 0.005579f
C3406 vdd.n2310 gnd 0.005579f
C3407 vdd.n2311 gnd 0.005579f
C3408 vdd.n2312 gnd 0.005579f
C3409 vdd.n2313 gnd 0.005579f
C3410 vdd.n2314 gnd 0.005579f
C3411 vdd.n2315 gnd 0.005579f
C3412 vdd.n2316 gnd 0.005579f
C3413 vdd.n2317 gnd 0.005579f
C3414 vdd.n2318 gnd 0.005579f
C3415 vdd.n2319 gnd 0.005579f
C3416 vdd.n2320 gnd 0.005579f
C3417 vdd.n2321 gnd 0.005579f
C3418 vdd.n2322 gnd 0.005579f
C3419 vdd.n2323 gnd 0.012667f
C3420 vdd.n2324 gnd 0.011945f
C3421 vdd.n2325 gnd 0.011945f
C3422 vdd.n2326 gnd 0.645553f
C3423 vdd.n2327 gnd 0.011945f
C3424 vdd.n2328 gnd 0.012667f
C3425 vdd.n2329 gnd 0.011945f
C3426 vdd.n2330 gnd 0.005579f
C3427 vdd.n2331 gnd 0.005579f
C3428 vdd.n2332 gnd 0.005579f
C3429 vdd.n2333 gnd 0.004307f
C3430 vdd.n2334 gnd 0.007973f
C3431 vdd.n2335 gnd 0.004061f
C3432 vdd.n2336 gnd 0.005579f
C3433 vdd.n2337 gnd 0.005579f
C3434 vdd.n2338 gnd 0.005579f
C3435 vdd.n2339 gnd 0.005579f
C3436 vdd.n2340 gnd 0.005579f
C3437 vdd.n2341 gnd 0.005579f
C3438 vdd.n2342 gnd 0.005579f
C3439 vdd.n2343 gnd 0.005579f
C3440 vdd.n2344 gnd 0.005579f
C3441 vdd.n2345 gnd 0.005579f
C3442 vdd.n2346 gnd 0.005579f
C3443 vdd.n2347 gnd 0.005579f
C3444 vdd.n2348 gnd 0.005579f
C3445 vdd.n2349 gnd 0.005579f
C3446 vdd.n2350 gnd 0.005579f
C3447 vdd.n2351 gnd 0.005579f
C3448 vdd.n2352 gnd 0.005579f
C3449 vdd.n2353 gnd 0.005579f
C3450 vdd.n2354 gnd 0.005579f
C3451 vdd.n2355 gnd 0.005579f
C3452 vdd.n2356 gnd 0.005579f
C3453 vdd.n2357 gnd 0.005579f
C3454 vdd.n2358 gnd 0.005579f
C3455 vdd.n2359 gnd 0.005579f
C3456 vdd.n2360 gnd 0.005579f
C3457 vdd.n2361 gnd 0.005579f
C3458 vdd.n2362 gnd 0.005579f
C3459 vdd.n2363 gnd 0.005579f
C3460 vdd.n2364 gnd 0.005579f
C3461 vdd.n2365 gnd 0.005579f
C3462 vdd.n2366 gnd 0.005579f
C3463 vdd.n2367 gnd 0.005579f
C3464 vdd.n2368 gnd 0.005579f
C3465 vdd.n2369 gnd 0.005579f
C3466 vdd.n2370 gnd 0.005579f
C3467 vdd.n2371 gnd 0.005579f
C3468 vdd.n2372 gnd 0.005579f
C3469 vdd.n2373 gnd 0.005579f
C3470 vdd.n2374 gnd 0.005579f
C3471 vdd.n2375 gnd 0.005579f
C3472 vdd.n2376 gnd 0.005579f
C3473 vdd.n2377 gnd 0.005579f
C3474 vdd.n2378 gnd 0.005579f
C3475 vdd.n2379 gnd 0.005579f
C3476 vdd.n2380 gnd 0.005579f
C3477 vdd.n2381 gnd 0.005579f
C3478 vdd.n2382 gnd 0.005579f
C3479 vdd.n2383 gnd 0.005579f
C3480 vdd.n2384 gnd 0.005579f
C3481 vdd.n2385 gnd 0.005579f
C3482 vdd.n2386 gnd 0.005579f
C3483 vdd.n2387 gnd 0.005579f
C3484 vdd.n2388 gnd 0.005579f
C3485 vdd.n2389 gnd 0.005579f
C3486 vdd.n2390 gnd 0.005579f
C3487 vdd.n2391 gnd 0.005579f
C3488 vdd.n2392 gnd 0.005579f
C3489 vdd.n2393 gnd 0.005579f
C3490 vdd.n2394 gnd 0.005579f
C3491 vdd.n2395 gnd 0.005579f
C3492 vdd.n2396 gnd 0.012667f
C3493 vdd.n2397 gnd 0.012667f
C3494 vdd.n2398 gnd 0.695856f
C3495 vdd.t33 gnd 2.47322f
C3496 vdd.t20 gnd 2.47322f
C3497 vdd.n2432 gnd 0.012667f
C3498 vdd.t38 gnd 0.486261f
C3499 vdd.n2433 gnd 0.005579f
C3500 vdd.t125 gnd 0.225427f
C3501 vdd.t126 gnd 0.230753f
C3502 vdd.t123 gnd 0.147168f
C3503 vdd.n2434 gnd 0.079536f
C3504 vdd.n2435 gnd 0.045115f
C3505 vdd.n2436 gnd 0.005579f
C3506 vdd.t132 gnd 0.225427f
C3507 vdd.t133 gnd 0.230753f
C3508 vdd.t131 gnd 0.147168f
C3509 vdd.n2437 gnd 0.079536f
C3510 vdd.n2438 gnd 0.045115f
C3511 vdd.n2439 gnd 0.007973f
C3512 vdd.n2440 gnd 0.012667f
C3513 vdd.n2441 gnd 0.012667f
C3514 vdd.n2442 gnd 0.005579f
C3515 vdd.n2443 gnd 0.005579f
C3516 vdd.n2444 gnd 0.005579f
C3517 vdd.n2445 gnd 0.005579f
C3518 vdd.n2446 gnd 0.005579f
C3519 vdd.n2447 gnd 0.005579f
C3520 vdd.n2448 gnd 0.005579f
C3521 vdd.n2449 gnd 0.005579f
C3522 vdd.n2450 gnd 0.005579f
C3523 vdd.n2451 gnd 0.005579f
C3524 vdd.n2452 gnd 0.005579f
C3525 vdd.n2453 gnd 0.005579f
C3526 vdd.n2454 gnd 0.005579f
C3527 vdd.n2455 gnd 0.005579f
C3528 vdd.n2456 gnd 0.005579f
C3529 vdd.n2457 gnd 0.005579f
C3530 vdd.n2458 gnd 0.005579f
C3531 vdd.n2459 gnd 0.005579f
C3532 vdd.n2460 gnd 0.005579f
C3533 vdd.n2461 gnd 0.005579f
C3534 vdd.n2462 gnd 0.005579f
C3535 vdd.n2463 gnd 0.005579f
C3536 vdd.n2464 gnd 0.005579f
C3537 vdd.n2465 gnd 0.005579f
C3538 vdd.n2466 gnd 0.005579f
C3539 vdd.n2467 gnd 0.005579f
C3540 vdd.n2468 gnd 0.005579f
C3541 vdd.n2469 gnd 0.005579f
C3542 vdd.n2470 gnd 0.005579f
C3543 vdd.n2471 gnd 0.005579f
C3544 vdd.n2472 gnd 0.005579f
C3545 vdd.n2473 gnd 0.005579f
C3546 vdd.n2474 gnd 0.005579f
C3547 vdd.n2475 gnd 0.005579f
C3548 vdd.n2476 gnd 0.005579f
C3549 vdd.n2477 gnd 0.005579f
C3550 vdd.n2478 gnd 0.005579f
C3551 vdd.n2479 gnd 0.005579f
C3552 vdd.n2480 gnd 0.005579f
C3553 vdd.n2481 gnd 0.005579f
C3554 vdd.n2482 gnd 0.005579f
C3555 vdd.n2483 gnd 0.005579f
C3556 vdd.n2484 gnd 0.005579f
C3557 vdd.n2485 gnd 0.005579f
C3558 vdd.n2486 gnd 0.005579f
C3559 vdd.n2487 gnd 0.005579f
C3560 vdd.n2488 gnd 0.005579f
C3561 vdd.n2489 gnd 0.005579f
C3562 vdd.n2490 gnd 0.005579f
C3563 vdd.n2491 gnd 0.005579f
C3564 vdd.n2492 gnd 0.005579f
C3565 vdd.n2493 gnd 0.005579f
C3566 vdd.n2494 gnd 0.005579f
C3567 vdd.n2495 gnd 0.005579f
C3568 vdd.n2496 gnd 0.005579f
C3569 vdd.n2497 gnd 0.005579f
C3570 vdd.n2498 gnd 0.005579f
C3571 vdd.n2499 gnd 0.005579f
C3572 vdd.n2500 gnd 0.005579f
C3573 vdd.n2501 gnd 0.005579f
C3574 vdd.n2502 gnd 0.004061f
C3575 vdd.n2503 gnd 0.005579f
C3576 vdd.n2504 gnd 0.005579f
C3577 vdd.n2505 gnd 0.004307f
C3578 vdd.n2506 gnd 0.005579f
C3579 vdd.n2507 gnd 0.005579f
C3580 vdd.n2508 gnd 0.012667f
C3581 vdd.n2509 gnd 0.011945f
C3582 vdd.n2510 gnd 0.011945f
C3583 vdd.n2511 gnd 0.005579f
C3584 vdd.n2512 gnd 0.005579f
C3585 vdd.n2513 gnd 0.005579f
C3586 vdd.n2514 gnd 0.005579f
C3587 vdd.n2515 gnd 0.005579f
C3588 vdd.n2516 gnd 0.005579f
C3589 vdd.n2517 gnd 0.005579f
C3590 vdd.n2518 gnd 0.005579f
C3591 vdd.n2519 gnd 0.005579f
C3592 vdd.n2520 gnd 0.005579f
C3593 vdd.n2521 gnd 0.005579f
C3594 vdd.n2522 gnd 0.005579f
C3595 vdd.n2523 gnd 0.005579f
C3596 vdd.n2524 gnd 0.005579f
C3597 vdd.n2525 gnd 0.005579f
C3598 vdd.n2526 gnd 0.005579f
C3599 vdd.n2527 gnd 0.005579f
C3600 vdd.n2528 gnd 0.005579f
C3601 vdd.n2529 gnd 0.005579f
C3602 vdd.n2530 gnd 0.005579f
C3603 vdd.n2531 gnd 0.005579f
C3604 vdd.n2532 gnd 0.005579f
C3605 vdd.n2533 gnd 0.005579f
C3606 vdd.n2534 gnd 0.005579f
C3607 vdd.n2535 gnd 0.005579f
C3608 vdd.n2536 gnd 0.005579f
C3609 vdd.n2537 gnd 0.005579f
C3610 vdd.n2538 gnd 0.005579f
C3611 vdd.n2539 gnd 0.005579f
C3612 vdd.n2540 gnd 0.005579f
C3613 vdd.n2541 gnd 0.005579f
C3614 vdd.n2542 gnd 0.005579f
C3615 vdd.n2543 gnd 0.005579f
C3616 vdd.n2544 gnd 0.005579f
C3617 vdd.n2545 gnd 0.005579f
C3618 vdd.n2546 gnd 0.005579f
C3619 vdd.n2547 gnd 0.005579f
C3620 vdd.n2548 gnd 0.005579f
C3621 vdd.n2549 gnd 0.005579f
C3622 vdd.n2550 gnd 0.005579f
C3623 vdd.n2551 gnd 0.005579f
C3624 vdd.n2552 gnd 0.005579f
C3625 vdd.n2553 gnd 0.005579f
C3626 vdd.n2554 gnd 0.005579f
C3627 vdd.n2555 gnd 0.005579f
C3628 vdd.n2556 gnd 0.005579f
C3629 vdd.n2557 gnd 0.005579f
C3630 vdd.n2558 gnd 0.005579f
C3631 vdd.n2559 gnd 0.005579f
C3632 vdd.n2560 gnd 0.005579f
C3633 vdd.n2561 gnd 0.005579f
C3634 vdd.n2562 gnd 0.005579f
C3635 vdd.n2563 gnd 0.005579f
C3636 vdd.n2564 gnd 0.005579f
C3637 vdd.n2565 gnd 0.005579f
C3638 vdd.n2566 gnd 0.005579f
C3639 vdd.n2567 gnd 0.005579f
C3640 vdd.n2568 gnd 0.005579f
C3641 vdd.n2569 gnd 0.005579f
C3642 vdd.n2570 gnd 0.005579f
C3643 vdd.n2571 gnd 0.005579f
C3644 vdd.n2572 gnd 0.005579f
C3645 vdd.n2573 gnd 0.005579f
C3646 vdd.n2574 gnd 0.005579f
C3647 vdd.n2575 gnd 0.005579f
C3648 vdd.n2576 gnd 0.005579f
C3649 vdd.n2577 gnd 0.005579f
C3650 vdd.n2578 gnd 0.005579f
C3651 vdd.n2579 gnd 0.005579f
C3652 vdd.n2580 gnd 0.005579f
C3653 vdd.n2581 gnd 0.005579f
C3654 vdd.n2582 gnd 0.005579f
C3655 vdd.n2583 gnd 0.005579f
C3656 vdd.n2584 gnd 0.005579f
C3657 vdd.n2585 gnd 0.005579f
C3658 vdd.n2586 gnd 0.005579f
C3659 vdd.n2587 gnd 0.005579f
C3660 vdd.n2588 gnd 0.005579f
C3661 vdd.n2589 gnd 0.005579f
C3662 vdd.n2590 gnd 0.005579f
C3663 vdd.n2591 gnd 0.005579f
C3664 vdd.n2592 gnd 0.005579f
C3665 vdd.n2593 gnd 0.005579f
C3666 vdd.n2594 gnd 0.005579f
C3667 vdd.n2595 gnd 0.005579f
C3668 vdd.n2596 gnd 0.005579f
C3669 vdd.n2597 gnd 0.005579f
C3670 vdd.n2598 gnd 0.005579f
C3671 vdd.n2599 gnd 0.005579f
C3672 vdd.n2600 gnd 0.005579f
C3673 vdd.n2601 gnd 0.005579f
C3674 vdd.n2602 gnd 0.005579f
C3675 vdd.n2603 gnd 0.005579f
C3676 vdd.n2604 gnd 0.005579f
C3677 vdd.n2605 gnd 0.005579f
C3678 vdd.n2606 gnd 0.005579f
C3679 vdd.n2607 gnd 0.005579f
C3680 vdd.n2608 gnd 0.005579f
C3681 vdd.n2609 gnd 0.005579f
C3682 vdd.n2610 gnd 0.005579f
C3683 vdd.n2611 gnd 0.005579f
C3684 vdd.n2612 gnd 0.180252f
C3685 vdd.n2613 gnd 0.005579f
C3686 vdd.n2614 gnd 0.005579f
C3687 vdd.n2615 gnd 0.005579f
C3688 vdd.n2616 gnd 0.005579f
C3689 vdd.n2617 gnd 0.005579f
C3690 vdd.n2618 gnd 0.180252f
C3691 vdd.n2619 gnd 0.005579f
C3692 vdd.n2620 gnd 0.005579f
C3693 vdd.n2621 gnd 0.005579f
C3694 vdd.n2622 gnd 0.005579f
C3695 vdd.n2623 gnd 0.005579f
C3696 vdd.n2624 gnd 0.005579f
C3697 vdd.n2625 gnd 0.005579f
C3698 vdd.n2626 gnd 0.005579f
C3699 vdd.n2627 gnd 0.005579f
C3700 vdd.n2628 gnd 0.005579f
C3701 vdd.n2629 gnd 0.005579f
C3702 vdd.n2630 gnd 0.356312f
C3703 vdd.n2631 gnd 0.005579f
C3704 vdd.n2632 gnd 0.005579f
C3705 vdd.n2633 gnd 0.005579f
C3706 vdd.n2634 gnd 0.011945f
C3707 vdd.n2635 gnd 0.011945f
C3708 vdd.n2636 gnd 0.012667f
C3709 vdd.n2637 gnd 0.012667f
C3710 vdd.n2638 gnd 0.005579f
C3711 vdd.n2639 gnd 0.005579f
C3712 vdd.n2640 gnd 0.005579f
C3713 vdd.n2641 gnd 0.004307f
C3714 vdd.n2642 gnd 0.007973f
C3715 vdd.n2643 gnd 0.004061f
C3716 vdd.n2644 gnd 0.005579f
C3717 vdd.n2645 gnd 0.005579f
C3718 vdd.n2646 gnd 0.005579f
C3719 vdd.n2647 gnd 0.005579f
C3720 vdd.n2648 gnd 0.005579f
C3721 vdd.n2649 gnd 0.005579f
C3722 vdd.n2650 gnd 0.005579f
C3723 vdd.n2651 gnd 0.005579f
C3724 vdd.n2652 gnd 0.005579f
C3725 vdd.n2653 gnd 0.005579f
C3726 vdd.n2654 gnd 0.005579f
C3727 vdd.n2655 gnd 0.005579f
C3728 vdd.n2656 gnd 0.005579f
C3729 vdd.n2657 gnd 0.005579f
C3730 vdd.n2658 gnd 0.005579f
C3731 vdd.n2659 gnd 0.005579f
C3732 vdd.n2660 gnd 0.005579f
C3733 vdd.n2661 gnd 0.005579f
C3734 vdd.n2662 gnd 0.005579f
C3735 vdd.n2663 gnd 0.005579f
C3736 vdd.n2664 gnd 0.005579f
C3737 vdd.n2665 gnd 0.005579f
C3738 vdd.n2666 gnd 0.005579f
C3739 vdd.n2667 gnd 0.005579f
C3740 vdd.n2668 gnd 0.005579f
C3741 vdd.n2669 gnd 0.005579f
C3742 vdd.n2670 gnd 0.005579f
C3743 vdd.n2671 gnd 0.005579f
C3744 vdd.n2672 gnd 0.005579f
C3745 vdd.n2673 gnd 0.005579f
C3746 vdd.n2674 gnd 0.005579f
C3747 vdd.n2675 gnd 0.005579f
C3748 vdd.n2676 gnd 0.005579f
C3749 vdd.n2677 gnd 0.005579f
C3750 vdd.n2678 gnd 0.005579f
C3751 vdd.n2679 gnd 0.005579f
C3752 vdd.n2680 gnd 0.005579f
C3753 vdd.n2681 gnd 0.005579f
C3754 vdd.n2682 gnd 0.005579f
C3755 vdd.n2683 gnd 0.005579f
C3756 vdd.n2684 gnd 0.005579f
C3757 vdd.n2685 gnd 0.005579f
C3758 vdd.n2686 gnd 0.005579f
C3759 vdd.n2687 gnd 0.005579f
C3760 vdd.n2688 gnd 0.005579f
C3761 vdd.n2689 gnd 0.005579f
C3762 vdd.n2690 gnd 0.005579f
C3763 vdd.n2691 gnd 0.005579f
C3764 vdd.n2692 gnd 0.005579f
C3765 vdd.n2693 gnd 0.005579f
C3766 vdd.n2694 gnd 0.005579f
C3767 vdd.n2695 gnd 0.005579f
C3768 vdd.n2696 gnd 0.005579f
C3769 vdd.n2697 gnd 0.005579f
C3770 vdd.n2698 gnd 0.005579f
C3771 vdd.n2699 gnd 0.005579f
C3772 vdd.n2700 gnd 0.005579f
C3773 vdd.n2701 gnd 0.005579f
C3774 vdd.n2702 gnd 0.695856f
C3775 vdd.n2704 gnd 0.012667f
C3776 vdd.n2705 gnd 0.012667f
C3777 vdd.n2706 gnd 0.011945f
C3778 vdd.n2707 gnd 0.005579f
C3779 vdd.n2708 gnd 0.005579f
C3780 vdd.n2709 gnd 0.335352f
C3781 vdd.n2710 gnd 0.005579f
C3782 vdd.n2711 gnd 0.005579f
C3783 vdd.n2712 gnd 0.005579f
C3784 vdd.n2713 gnd 0.005579f
C3785 vdd.n2714 gnd 0.005579f
C3786 vdd.n2715 gnd 0.339544f
C3787 vdd.n2716 gnd 0.005579f
C3788 vdd.n2717 gnd 0.005579f
C3789 vdd.n2718 gnd 0.005579f
C3790 vdd.n2719 gnd 0.005579f
C3791 vdd.n2720 gnd 0.005579f
C3792 vdd.n2721 gnd 0.570099f
C3793 vdd.n2722 gnd 0.005579f
C3794 vdd.n2723 gnd 0.005579f
C3795 vdd.n2724 gnd 0.005579f
C3796 vdd.n2725 gnd 0.005579f
C3797 vdd.n2726 gnd 0.005579f
C3798 vdd.n2727 gnd 0.410806f
C3799 vdd.n2728 gnd 0.005579f
C3800 vdd.n2729 gnd 0.005579f
C3801 vdd.n2730 gnd 0.005579f
C3802 vdd.n2731 gnd 0.005579f
C3803 vdd.n2732 gnd 0.005579f
C3804 vdd.n2733 gnd 0.515604f
C3805 vdd.n2734 gnd 0.005579f
C3806 vdd.n2735 gnd 0.005579f
C3807 vdd.n2736 gnd 0.005579f
C3808 vdd.n2737 gnd 0.005579f
C3809 vdd.n2738 gnd 0.005579f
C3810 vdd.n2739 gnd 0.423382f
C3811 vdd.n2740 gnd 0.005579f
C3812 vdd.n2741 gnd 0.005579f
C3813 vdd.n2742 gnd 0.005579f
C3814 vdd.n2743 gnd 0.005579f
C3815 vdd.n2744 gnd 0.005579f
C3816 vdd.n2745 gnd 0.297625f
C3817 vdd.n2746 gnd 0.005579f
C3818 vdd.n2747 gnd 0.005579f
C3819 vdd.n2748 gnd 0.005579f
C3820 vdd.n2749 gnd 0.005579f
C3821 vdd.n2750 gnd 0.005579f
C3822 vdd.n2751 gnd 0.180252f
C3823 vdd.n2752 gnd 0.005579f
C3824 vdd.n2753 gnd 0.005579f
C3825 vdd.n2754 gnd 0.005579f
C3826 vdd.n2755 gnd 0.005579f
C3827 vdd.n2756 gnd 0.005579f
C3828 vdd.n2757 gnd 0.523988f
C3829 vdd.n2758 gnd 0.005579f
C3830 vdd.n2759 gnd 0.005579f
C3831 vdd.n2760 gnd 0.005579f
C3832 vdd.n2761 gnd 0.003938f
C3833 vdd.n2762 gnd 0.005579f
C3834 vdd.n2763 gnd 0.005579f
C3835 vdd.n2764 gnd 0.570099f
C3836 vdd.n2765 gnd 0.005579f
C3837 vdd.n2766 gnd 0.005579f
C3838 vdd.n2767 gnd 0.005579f
C3839 vdd.n2768 gnd 0.005579f
C3840 vdd.n2769 gnd 0.005579f
C3841 vdd.n2770 gnd 0.452725f
C3842 vdd.n2771 gnd 0.005579f
C3843 vdd.n2772 gnd 0.00443f
C3844 vdd.n2773 gnd 0.005579f
C3845 vdd.n2774 gnd 0.005579f
C3846 vdd.n2775 gnd 0.005579f
C3847 vdd.n2776 gnd 0.364695f
C3848 vdd.n2777 gnd 0.005579f
C3849 vdd.n2778 gnd 0.005579f
C3850 vdd.n2779 gnd 0.005579f
C3851 vdd.n2780 gnd 0.005579f
C3852 vdd.n2781 gnd 0.005579f
C3853 vdd.n2782 gnd 0.33116f
C3854 vdd.n2783 gnd 0.005579f
C3855 vdd.n2784 gnd 0.005579f
C3856 vdd.n2785 gnd 0.005579f
C3857 vdd.n2786 gnd 0.005579f
C3858 vdd.n2787 gnd 0.005579f
C3859 vdd.n2788 gnd 0.456917f
C3860 vdd.n2789 gnd 0.005579f
C3861 vdd.n2790 gnd 0.005579f
C3862 vdd.n2791 gnd 0.005579f
C3863 vdd.n2792 gnd 0.005579f
C3864 vdd.n2793 gnd 0.005579f
C3865 vdd.n2794 gnd 0.570099f
C3866 vdd.n2795 gnd 0.005579f
C3867 vdd.n2796 gnd 0.005579f
C3868 vdd.n2797 gnd 0.005579f
C3869 vdd.n2798 gnd 0.005579f
C3870 vdd.n2799 gnd 0.005579f
C3871 vdd.n2800 gnd 0.557523f
C3872 vdd.n2801 gnd 0.005579f
C3873 vdd.n2802 gnd 0.005579f
C3874 vdd.n2803 gnd 0.005579f
C3875 vdd.n2804 gnd 0.005579f
C3876 vdd.n2805 gnd 0.005579f
C3877 vdd.n2806 gnd 0.431766f
C3878 vdd.n2807 gnd 0.005579f
C3879 vdd.n2808 gnd 0.005579f
C3880 vdd.n2809 gnd 0.005579f
C3881 vdd.n2810 gnd 0.005579f
C3882 vdd.n2811 gnd 0.005579f
C3883 vdd.n2812 gnd 0.306009f
C3884 vdd.n2813 gnd 0.005579f
C3885 vdd.n2814 gnd 0.005579f
C3886 vdd.n2815 gnd 0.005579f
C3887 vdd.n2816 gnd 0.005579f
C3888 vdd.n2817 gnd 0.005579f
C3889 vdd.n2818 gnd 0.570099f
C3890 vdd.n2819 gnd 0.005579f
C3891 vdd.n2820 gnd 0.005579f
C3892 vdd.n2821 gnd 0.005579f
C3893 vdd.n2822 gnd 0.005579f
C3894 vdd.n2823 gnd 0.005579f
C3895 vdd.n2824 gnd 0.005579f
C3896 vdd.n2826 gnd 0.005579f
C3897 vdd.n2827 gnd 0.005579f
C3898 vdd.n2829 gnd 0.005579f
C3899 vdd.n2830 gnd 0.005579f
C3900 vdd.n2833 gnd 0.005579f
C3901 vdd.n2834 gnd 0.005579f
C3902 vdd.n2835 gnd 0.005579f
C3903 vdd.n2836 gnd 0.005579f
C3904 vdd.n2838 gnd 0.005579f
C3905 vdd.n2839 gnd 0.005579f
C3906 vdd.n2840 gnd 0.005579f
C3907 vdd.n2841 gnd 0.005579f
C3908 vdd.n2842 gnd 0.005579f
C3909 vdd.n2843 gnd 0.005579f
C3910 vdd.n2845 gnd 0.005579f
C3911 vdd.n2846 gnd 0.005579f
C3912 vdd.n2847 gnd 0.005579f
C3913 vdd.n2848 gnd 0.005579f
C3914 vdd.n2849 gnd 0.005579f
C3915 vdd.n2850 gnd 0.005579f
C3916 vdd.n2852 gnd 0.005579f
C3917 vdd.n2853 gnd 0.005579f
C3918 vdd.n2854 gnd 0.005579f
C3919 vdd.n2855 gnd 0.005579f
C3920 vdd.n2856 gnd 0.005579f
C3921 vdd.n2857 gnd 0.005579f
C3922 vdd.n2859 gnd 0.005579f
C3923 vdd.n2860 gnd 0.012667f
C3924 vdd.n2861 gnd 0.012667f
C3925 vdd.n2862 gnd 0.011945f
C3926 vdd.n2863 gnd 0.005579f
C3927 vdd.n2864 gnd 0.005579f
C3928 vdd.n2865 gnd 0.005579f
C3929 vdd.n2866 gnd 0.005579f
C3930 vdd.n2867 gnd 0.005579f
C3931 vdd.n2868 gnd 0.005579f
C3932 vdd.n2869 gnd 0.570099f
C3933 vdd.n2870 gnd 0.005579f
C3934 vdd.n2871 gnd 0.005579f
C3935 vdd.n2872 gnd 0.005579f
C3936 vdd.n2873 gnd 0.005579f
C3937 vdd.n2874 gnd 0.005579f
C3938 vdd.n2875 gnd 0.406614f
C3939 vdd.n2876 gnd 0.005579f
C3940 vdd.n2877 gnd 0.005579f
C3941 vdd.n2878 gnd 0.005579f
C3942 vdd.n2879 gnd 0.012667f
C3943 vdd.n2880 gnd 0.011945f
C3944 vdd.n2881 gnd 0.012667f
C3945 vdd.n2883 gnd 0.005579f
C3946 vdd.n2884 gnd 0.005579f
C3947 vdd.n2885 gnd 0.004307f
C3948 vdd.n2886 gnd 0.007973f
C3949 vdd.n2887 gnd 0.004061f
C3950 vdd.n2888 gnd 0.005579f
C3951 vdd.n2889 gnd 0.005579f
C3952 vdd.n2891 gnd 0.005579f
C3953 vdd.n2892 gnd 0.005579f
C3954 vdd.n2893 gnd 0.005579f
C3955 vdd.n2894 gnd 0.005579f
C3956 vdd.n2895 gnd 0.005579f
C3957 vdd.n2896 gnd 0.005579f
C3958 vdd.n2898 gnd 0.005579f
C3959 vdd.n2899 gnd 0.005579f
C3960 vdd.n2900 gnd 0.005579f
C3961 vdd.n2901 gnd 0.005579f
C3962 vdd.n2902 gnd 0.005579f
C3963 vdd.n2903 gnd 0.005579f
C3964 vdd.n2905 gnd 0.005579f
C3965 vdd.n2906 gnd 0.005579f
C3966 vdd.n2907 gnd 0.005579f
C3967 vdd.n2908 gnd 0.005579f
C3968 vdd.n2909 gnd 0.005579f
C3969 vdd.n2910 gnd 0.005579f
C3970 vdd.n2912 gnd 0.005579f
C3971 vdd.n2913 gnd 0.005579f
C3972 vdd.n2914 gnd 0.005579f
C3973 vdd.n2916 gnd 0.005579f
C3974 vdd.n2917 gnd 0.005579f
C3975 vdd.n2918 gnd 0.005579f
C3976 vdd.n2919 gnd 0.005579f
C3977 vdd.n2920 gnd 0.005579f
C3978 vdd.n2921 gnd 0.005579f
C3979 vdd.n2923 gnd 0.005579f
C3980 vdd.n2924 gnd 0.005579f
C3981 vdd.n2925 gnd 0.005579f
C3982 vdd.n2926 gnd 0.005579f
C3983 vdd.n2927 gnd 0.005579f
C3984 vdd.n2928 gnd 0.005579f
C3985 vdd.n2930 gnd 0.005579f
C3986 vdd.n2931 gnd 0.005579f
C3987 vdd.n2932 gnd 0.005579f
C3988 vdd.n2933 gnd 0.005579f
C3989 vdd.n2934 gnd 0.005579f
C3990 vdd.n2935 gnd 0.005579f
C3991 vdd.n2937 gnd 0.005579f
C3992 vdd.n2938 gnd 0.005579f
C3993 vdd.n2940 gnd 0.005579f
C3994 vdd.n2941 gnd 0.005579f
C3995 vdd.n2942 gnd 0.012667f
C3996 vdd.n2943 gnd 0.011945f
C3997 vdd.n2944 gnd 0.011945f
C3998 vdd.n2945 gnd 0.77131f
C3999 vdd.n2946 gnd 0.011945f
C4000 vdd.n2947 gnd 0.012667f
C4001 vdd.n2948 gnd 0.011945f
C4002 vdd.n2949 gnd 0.005579f
C4003 vdd.n2950 gnd 0.004307f
C4004 vdd.n2951 gnd 0.005579f
C4005 vdd.n2953 gnd 0.005579f
C4006 vdd.n2954 gnd 0.005579f
C4007 vdd.n2955 gnd 0.005579f
C4008 vdd.n2956 gnd 0.005579f
C4009 vdd.n2957 gnd 0.005579f
C4010 vdd.n2958 gnd 0.005579f
C4011 vdd.n2960 gnd 0.005579f
C4012 vdd.n2961 gnd 0.005579f
C4013 vdd.n2962 gnd 0.005579f
C4014 vdd.n2963 gnd 0.005579f
C4015 vdd.n2964 gnd 0.005579f
C4016 vdd.n2965 gnd 0.005579f
C4017 vdd.n2967 gnd 0.005579f
C4018 vdd.n2968 gnd 0.005579f
C4019 vdd.n2969 gnd 0.005579f
C4020 vdd.n2970 gnd 0.005579f
C4021 vdd.n2971 gnd 0.005579f
C4022 vdd.n2972 gnd 0.005579f
C4023 vdd.n2974 gnd 0.005579f
C4024 vdd.n2975 gnd 0.005579f
C4025 vdd.n2977 gnd 0.005579f
C4026 vdd.n2978 gnd 0.034447f
C4027 vdd.n2979 gnd 0.874042f
C4028 vdd.n2980 gnd 0.007055f
C4029 vdd.n2981 gnd 0.020451f
C4030 vdd.n2982 gnd 0.003136f
C4031 vdd.t87 gnd 0.100927f
C4032 vdd.t88 gnd 0.107863f
C4033 vdd.t85 gnd 0.13181f
C4034 vdd.n2983 gnd 0.168961f
C4035 vdd.n2984 gnd 0.141958f
C4036 vdd.n2985 gnd 0.010169f
C4037 vdd.n2986 gnd 0.008204f
C4038 vdd.n2987 gnd 0.003467f
C4039 vdd.n2988 gnd 0.006603f
C4040 vdd.n2989 gnd 0.008204f
C4041 vdd.n2990 gnd 0.008204f
C4042 vdd.n2991 gnd 0.006603f
C4043 vdd.n2992 gnd 0.006603f
C4044 vdd.n2993 gnd 0.008204f
C4045 vdd.n2994 gnd 0.008204f
C4046 vdd.n2995 gnd 0.006603f
C4047 vdd.n2996 gnd 0.006603f
C4048 vdd.n2997 gnd 0.008204f
C4049 vdd.n2998 gnd 0.008204f
C4050 vdd.n2999 gnd 0.006603f
C4051 vdd.n3000 gnd 0.006603f
C4052 vdd.n3001 gnd 0.008204f
C4053 vdd.n3002 gnd 0.008204f
C4054 vdd.n3003 gnd 0.006603f
C4055 vdd.n3004 gnd 0.006603f
C4056 vdd.n3005 gnd 0.008204f
C4057 vdd.n3006 gnd 0.008204f
C4058 vdd.n3007 gnd 0.006603f
C4059 vdd.n3008 gnd 0.006603f
C4060 vdd.n3009 gnd 0.008204f
C4061 vdd.n3010 gnd 0.008204f
C4062 vdd.n3011 gnd 0.006603f
C4063 vdd.n3012 gnd 0.006603f
C4064 vdd.n3013 gnd 0.008204f
C4065 vdd.n3014 gnd 0.008204f
C4066 vdd.n3015 gnd 0.006603f
C4067 vdd.n3016 gnd 0.006603f
C4068 vdd.n3017 gnd 0.008204f
C4069 vdd.n3018 gnd 0.008204f
C4070 vdd.n3019 gnd 0.006603f
C4071 vdd.n3020 gnd 0.006603f
C4072 vdd.n3021 gnd 0.008204f
C4073 vdd.n3022 gnd 0.008204f
C4074 vdd.n3023 gnd 0.006603f
C4075 vdd.n3024 gnd 0.008204f
C4076 vdd.n3025 gnd 0.008204f
C4077 vdd.n3026 gnd 0.006603f
C4078 vdd.n3027 gnd 0.008204f
C4079 vdd.n3028 gnd 0.008204f
C4080 vdd.n3029 gnd 0.008204f
C4081 vdd.n3030 gnd 0.01347f
C4082 vdd.n3031 gnd 0.008204f
C4083 vdd.n3032 gnd 0.008204f
C4084 vdd.n3033 gnd 0.00449f
C4085 vdd.n3034 gnd 0.006603f
C4086 vdd.n3035 gnd 0.008204f
C4087 vdd.n3036 gnd 0.008204f
C4088 vdd.n3037 gnd 0.006603f
C4089 vdd.n3038 gnd 0.006603f
C4090 vdd.n3039 gnd 0.008204f
C4091 vdd.n3040 gnd 0.008204f
C4092 vdd.n3041 gnd 0.006603f
C4093 vdd.n3042 gnd 0.006603f
C4094 vdd.n3043 gnd 0.008204f
C4095 vdd.n3044 gnd 0.008204f
C4096 vdd.n3045 gnd 0.006603f
C4097 vdd.n3046 gnd 0.006603f
C4098 vdd.n3047 gnd 0.008204f
C4099 vdd.n3048 gnd 0.008204f
C4100 vdd.n3049 gnd 0.006603f
C4101 vdd.n3050 gnd 0.006603f
C4102 vdd.n3051 gnd 0.008204f
C4103 vdd.n3052 gnd 0.008204f
C4104 vdd.n3053 gnd 0.006603f
C4105 vdd.n3054 gnd 0.006603f
C4106 vdd.n3055 gnd 0.008204f
C4107 vdd.n3056 gnd 0.008204f
C4108 vdd.n3057 gnd 0.006603f
C4109 vdd.n3058 gnd 0.006603f
C4110 vdd.n3059 gnd 0.008204f
C4111 vdd.n3060 gnd 0.008204f
C4112 vdd.n3061 gnd 0.006603f
C4113 vdd.n3062 gnd 0.006603f
C4114 vdd.n3063 gnd 0.008204f
C4115 vdd.n3064 gnd 0.008204f
C4116 vdd.n3065 gnd 0.006603f
C4117 vdd.n3066 gnd 0.006603f
C4118 vdd.n3067 gnd 0.008204f
C4119 vdd.n3068 gnd 0.008204f
C4120 vdd.n3069 gnd 0.006603f
C4121 vdd.n3070 gnd 0.008204f
C4122 vdd.n3071 gnd 0.008204f
C4123 vdd.n3072 gnd 0.006603f
C4124 vdd.n3073 gnd 0.008204f
C4125 vdd.n3074 gnd 0.008204f
C4126 vdd.n3075 gnd 0.008204f
C4127 vdd.t121 gnd 0.100927f
C4128 vdd.t122 gnd 0.107863f
C4129 vdd.t120 gnd 0.13181f
C4130 vdd.n3076 gnd 0.168961f
C4131 vdd.n3077 gnd 0.141958f
C4132 vdd.n3078 gnd 0.01347f
C4133 vdd.n3079 gnd 0.008204f
C4134 vdd.n3080 gnd 0.008204f
C4135 vdd.n3081 gnd 0.005514f
C4136 vdd.n3082 gnd 0.006603f
C4137 vdd.n3083 gnd 0.008204f
C4138 vdd.n3084 gnd 0.008204f
C4139 vdd.n3085 gnd 0.006603f
C4140 vdd.n3086 gnd 0.006603f
C4141 vdd.n3087 gnd 0.008204f
C4142 vdd.n3088 gnd 0.008204f
C4143 vdd.n3089 gnd 0.006603f
C4144 vdd.n3090 gnd 0.006603f
C4145 vdd.n3091 gnd 0.008204f
C4146 vdd.n3092 gnd 0.008204f
C4147 vdd.n3093 gnd 0.006603f
C4148 vdd.n3094 gnd 0.006603f
C4149 vdd.n3095 gnd 0.008204f
C4150 vdd.n3096 gnd 0.008204f
C4151 vdd.n3097 gnd 0.006603f
C4152 vdd.n3098 gnd 0.006603f
C4153 vdd.n3099 gnd 0.008204f
C4154 vdd.n3100 gnd 0.008204f
C4155 vdd.n3101 gnd 0.006603f
C4156 vdd.n3102 gnd 0.006603f
C4157 vdd.n3103 gnd 0.008204f
C4158 vdd.n3104 gnd 0.008204f
C4159 vdd.n3105 gnd 0.006603f
C4160 vdd.n3106 gnd 0.006603f
C4161 vdd.n3108 gnd 0.874042f
C4162 vdd.n3110 gnd 0.006603f
C4163 vdd.n3111 gnd 0.008204f
C4164 vdd.n3112 gnd 10.253401f
C4165 vdd.n3114 gnd 0.020451f
C4166 vdd.n3115 gnd 0.00548f
C4167 vdd.n3116 gnd 0.020451f
C4168 vdd.n3117 gnd 0.019993f
C4169 vdd.n3118 gnd 0.008204f
C4170 vdd.n3119 gnd 0.006603f
C4171 vdd.n3120 gnd 0.008204f
C4172 vdd.n3121 gnd 0.523988f
C4173 vdd.n3122 gnd 0.008204f
C4174 vdd.n3123 gnd 0.006603f
C4175 vdd.n3124 gnd 0.008204f
C4176 vdd.n3125 gnd 0.008204f
C4177 vdd.n3126 gnd 0.008204f
C4178 vdd.n3127 gnd 0.006603f
C4179 vdd.n3128 gnd 0.008204f
C4180 vdd.n3129 gnd 0.666512f
C4181 vdd.n3130 gnd 0.83838f
C4182 vdd.n3131 gnd 0.008204f
C4183 vdd.n3132 gnd 0.006603f
C4184 vdd.n3133 gnd 0.008204f
C4185 vdd.n3134 gnd 0.008204f
C4186 vdd.n3135 gnd 0.008204f
C4187 vdd.n3136 gnd 0.006603f
C4188 vdd.n3137 gnd 0.008204f
C4189 vdd.n3138 gnd 0.591058f
C4190 vdd.n3139 gnd 0.008204f
C4191 vdd.n3140 gnd 0.006603f
C4192 vdd.n3141 gnd 0.008204f
C4193 vdd.n3142 gnd 0.008204f
C4194 vdd.n3143 gnd 0.008204f
C4195 vdd.n3144 gnd 0.006603f
C4196 vdd.n3145 gnd 0.008204f
C4197 vdd.t156 gnd 0.41919f
C4198 vdd.n3146 gnd 0.695856f
C4199 vdd.n3147 gnd 0.008204f
C4200 vdd.n3148 gnd 0.006603f
C4201 vdd.n3149 gnd 0.008204f
C4202 vdd.n3150 gnd 0.008204f
C4203 vdd.n3151 gnd 0.008204f
C4204 vdd.n3152 gnd 0.006603f
C4205 vdd.n3153 gnd 0.008204f
C4206 vdd.n3154 gnd 0.658129f
C4207 vdd.n3155 gnd 0.008204f
C4208 vdd.n3156 gnd 0.006603f
C4209 vdd.n3157 gnd 0.008204f
C4210 vdd.n3158 gnd 0.008204f
C4211 vdd.n3159 gnd 0.008204f
C4212 vdd.n3160 gnd 0.006603f
C4213 vdd.n3161 gnd 0.006603f
C4214 vdd.n3162 gnd 0.006603f
C4215 vdd.n3163 gnd 0.008204f
C4216 vdd.n3164 gnd 0.008204f
C4217 vdd.n3165 gnd 0.008204f
C4218 vdd.n3166 gnd 0.006603f
C4219 vdd.n3167 gnd 0.006603f
C4220 vdd.n3168 gnd 0.006603f
C4221 vdd.n3169 gnd 0.008204f
C4222 vdd.n3170 gnd 0.008204f
C4223 vdd.n3171 gnd 0.008204f
C4224 vdd.n3172 gnd 0.006603f
C4225 vdd.n3173 gnd 0.006603f
C4226 vdd.n3174 gnd 0.00548f
C4227 vdd.n3175 gnd 0.019993f
C4228 vdd.n3176 gnd 0.020451f
C4229 vdd.n3178 gnd 0.020451f
C4230 vdd.n3179 gnd 0.003136f
C4231 vdd.t103 gnd 0.100927f
C4232 vdd.t102 gnd 0.107863f
C4233 vdd.t100 gnd 0.13181f
C4234 vdd.n3180 gnd 0.168961f
C4235 vdd.n3181 gnd 0.142618f
C4236 vdd.n3182 gnd 0.010829f
C4237 vdd.n3183 gnd 0.003467f
C4238 vdd.n3184 gnd 0.006603f
C4239 vdd.n3185 gnd 0.008204f
C4240 vdd.n3187 gnd 0.008204f
C4241 vdd.n3188 gnd 0.008204f
C4242 vdd.n3189 gnd 0.006603f
C4243 vdd.n3190 gnd 0.006603f
C4244 vdd.n3191 gnd 0.006603f
C4245 vdd.n3192 gnd 0.008204f
C4246 vdd.n3194 gnd 0.008204f
C4247 vdd.n3195 gnd 0.008204f
C4248 vdd.n3196 gnd 0.006603f
C4249 vdd.n3197 gnd 0.006603f
C4250 vdd.n3198 gnd 0.006603f
C4251 vdd.n3199 gnd 0.008204f
C4252 vdd.n3201 gnd 0.008204f
C4253 vdd.n3202 gnd 0.008204f
C4254 vdd.n3203 gnd 0.006603f
C4255 vdd.n3204 gnd 0.006603f
C4256 vdd.n3205 gnd 0.006603f
C4257 vdd.n3206 gnd 0.008204f
C4258 vdd.n3208 gnd 0.008204f
C4259 vdd.n3209 gnd 0.008204f
C4260 vdd.n3210 gnd 0.006603f
C4261 vdd.n3211 gnd 0.006603f
C4262 vdd.n3212 gnd 0.006603f
C4263 vdd.n3213 gnd 0.008204f
C4264 vdd.n3215 gnd 0.008204f
C4265 vdd.n3216 gnd 0.008204f
C4266 vdd.n3217 gnd 0.006603f
C4267 vdd.n3218 gnd 0.008204f
C4268 vdd.n3219 gnd 0.008204f
C4269 vdd.n3220 gnd 0.008204f
C4270 vdd.n3221 gnd 0.01413f
C4271 vdd.n3222 gnd 0.00449f
C4272 vdd.n3223 gnd 0.006603f
C4273 vdd.n3224 gnd 0.008204f
C4274 vdd.n3226 gnd 0.008204f
C4275 vdd.n3227 gnd 0.008204f
C4276 vdd.n3228 gnd 0.006603f
C4277 vdd.n3229 gnd 0.006603f
C4278 vdd.n3230 gnd 0.006603f
C4279 vdd.n3231 gnd 0.008204f
C4280 vdd.n3233 gnd 0.008204f
C4281 vdd.n3234 gnd 0.008204f
C4282 vdd.n3235 gnd 0.006603f
C4283 vdd.n3236 gnd 0.006603f
C4284 vdd.n3237 gnd 0.006603f
C4285 vdd.n3238 gnd 0.008204f
C4286 vdd.n3240 gnd 0.008204f
C4287 vdd.n3241 gnd 0.008204f
C4288 vdd.n3242 gnd 0.006603f
C4289 vdd.n3243 gnd 0.006603f
C4290 vdd.n3244 gnd 0.006603f
C4291 vdd.n3245 gnd 0.008204f
C4292 vdd.n3247 gnd 0.008204f
C4293 vdd.n3248 gnd 0.008204f
C4294 vdd.n3249 gnd 0.006603f
C4295 vdd.n3250 gnd 0.006603f
C4296 vdd.n3251 gnd 0.006603f
C4297 vdd.n3252 gnd 0.008204f
C4298 vdd.n3254 gnd 0.008204f
C4299 vdd.n3255 gnd 0.008204f
C4300 vdd.n3256 gnd 0.006603f
C4301 vdd.n3257 gnd 0.008204f
C4302 vdd.n3258 gnd 0.008204f
C4303 vdd.n3259 gnd 0.008204f
C4304 vdd.n3260 gnd 0.01413f
C4305 vdd.n3261 gnd 0.005514f
C4306 vdd.n3262 gnd 0.006603f
C4307 vdd.n3263 gnd 0.008204f
C4308 vdd.n3265 gnd 0.008204f
C4309 vdd.n3266 gnd 0.008204f
C4310 vdd.n3267 gnd 0.006603f
C4311 vdd.n3268 gnd 0.006603f
C4312 vdd.n3269 gnd 0.006603f
C4313 vdd.n3270 gnd 0.008204f
C4314 vdd.n3272 gnd 0.008204f
C4315 vdd.n3273 gnd 0.008204f
C4316 vdd.n3274 gnd 0.006603f
C4317 vdd.n3275 gnd 0.006603f
C4318 vdd.n3276 gnd 0.006603f
C4319 vdd.n3277 gnd 0.008204f
C4320 vdd.n3279 gnd 0.008204f
C4321 vdd.n3280 gnd 0.008204f
C4322 vdd.n3281 gnd 0.006603f
C4323 vdd.n3282 gnd 0.006603f
C4324 vdd.n3283 gnd 0.006603f
C4325 vdd.n3284 gnd 0.008204f
C4326 vdd.n3286 gnd 0.008204f
C4327 vdd.n3287 gnd 0.008204f
C4328 vdd.n3289 gnd 0.008204f
C4329 vdd.n3290 gnd 0.006603f
C4330 vdd.n3291 gnd 0.006603f
C4331 vdd.n3292 gnd 0.00548f
C4332 vdd.n3293 gnd 0.020451f
C4333 vdd.n3294 gnd 0.019993f
C4334 vdd.n3295 gnd 0.00548f
C4335 vdd.n3296 gnd 0.019993f
C4336 vdd.n3297 gnd 1.23661f
C4337 vdd.t101 gnd 0.41919f
C4338 vdd.n3298 gnd 0.44015f
C4339 vdd.n3299 gnd 0.83838f
C4340 vdd.n3300 gnd 0.008204f
C4341 vdd.n3301 gnd 0.006603f
C4342 vdd.n3302 gnd 0.006603f
C4343 vdd.n3303 gnd 0.006603f
C4344 vdd.n3304 gnd 0.008204f
C4345 vdd.n3305 gnd 0.75035f
C4346 vdd.t177 gnd 0.41919f
C4347 vdd.n3306 gnd 0.50722f
C4348 vdd.n3307 gnd 0.607826f
C4349 vdd.n3308 gnd 0.008204f
C4350 vdd.n3309 gnd 0.006603f
C4351 vdd.n3310 gnd 0.006603f
C4352 vdd.n3311 gnd 0.006603f
C4353 vdd.n3312 gnd 0.008204f
C4354 vdd.n3313 gnd 0.465301f
C4355 vdd.t154 gnd 0.41919f
C4356 vdd.n3314 gnd 0.695856f
C4357 vdd.t195 gnd 0.41919f
C4358 vdd.n3315 gnd 0.515604f
C4359 vdd.n3316 gnd 0.008204f
C4360 vdd.n3317 gnd 0.006603f
C4361 vdd.n3318 gnd 0.006305f
C4362 vdd.n3319 gnd 0.483886f
C4363 vdd.n3320 gnd 1.95934f
C4364 a_n2804_13878.t20 gnd 0.194878f
C4365 a_n2804_13878.t7 gnd 0.194878f
C4366 a_n2804_13878.t17 gnd 0.194878f
C4367 a_n2804_13878.n0 gnd 1.53612f
C4368 a_n2804_13878.t22 gnd 0.194878f
C4369 a_n2804_13878.t12 gnd 0.194878f
C4370 a_n2804_13878.n1 gnd 1.5345f
C4371 a_n2804_13878.n2 gnd 2.14416f
C4372 a_n2804_13878.t18 gnd 0.194878f
C4373 a_n2804_13878.t11 gnd 0.194878f
C4374 a_n2804_13878.n3 gnd 1.5345f
C4375 a_n2804_13878.n4 gnd 1.04587f
C4376 a_n2804_13878.t5 gnd 0.194878f
C4377 a_n2804_13878.t8 gnd 0.194878f
C4378 a_n2804_13878.n5 gnd 1.5345f
C4379 a_n2804_13878.n6 gnd 1.04587f
C4380 a_n2804_13878.t21 gnd 0.194878f
C4381 a_n2804_13878.t6 gnd 0.194878f
C4382 a_n2804_13878.n7 gnd 1.5345f
C4383 a_n2804_13878.n8 gnd 1.04587f
C4384 a_n2804_13878.t16 gnd 0.194878f
C4385 a_n2804_13878.t4 gnd 0.194878f
C4386 a_n2804_13878.n9 gnd 1.5345f
C4387 a_n2804_13878.n10 gnd 4.90989f
C4388 a_n2804_13878.t30 gnd 1.82474f
C4389 a_n2804_13878.t0 gnd 0.194878f
C4390 a_n2804_13878.t29 gnd 0.194878f
C4391 a_n2804_13878.n11 gnd 1.37272f
C4392 a_n2804_13878.n12 gnd 1.53381f
C4393 a_n2804_13878.t2 gnd 1.8211f
C4394 a_n2804_13878.n13 gnd 0.771835f
C4395 a_n2804_13878.t28 gnd 1.8211f
C4396 a_n2804_13878.n14 gnd 0.771835f
C4397 a_n2804_13878.t27 gnd 0.194878f
C4398 a_n2804_13878.t1 gnd 0.194878f
C4399 a_n2804_13878.n15 gnd 1.37272f
C4400 a_n2804_13878.n16 gnd 0.77931f
C4401 a_n2804_13878.t31 gnd 1.8211f
C4402 a_n2804_13878.n17 gnd 2.86287f
C4403 a_n2804_13878.n18 gnd 3.75497f
C4404 a_n2804_13878.t10 gnd 0.194878f
C4405 a_n2804_13878.t19 gnd 0.194878f
C4406 a_n2804_13878.n19 gnd 1.53449f
C4407 a_n2804_13878.n20 gnd 2.50654f
C4408 a_n2804_13878.t23 gnd 0.194878f
C4409 a_n2804_13878.t9 gnd 0.194878f
C4410 a_n2804_13878.n21 gnd 1.5345f
C4411 a_n2804_13878.n22 gnd 0.679894f
C4412 a_n2804_13878.t13 gnd 0.194878f
C4413 a_n2804_13878.t14 gnd 0.194878f
C4414 a_n2804_13878.n23 gnd 1.5345f
C4415 a_n2804_13878.n24 gnd 0.679894f
C4416 a_n2804_13878.t24 gnd 0.194878f
C4417 a_n2804_13878.t25 gnd 0.194878f
C4418 a_n2804_13878.n25 gnd 1.5345f
C4419 a_n2804_13878.n26 gnd 0.679894f
C4420 a_n2804_13878.t3 gnd 0.194878f
C4421 a_n2804_13878.t15 gnd 0.194878f
C4422 a_n2804_13878.n27 gnd 1.5345f
C4423 a_n2804_13878.n28 gnd 1.37932f
C4424 a_n2804_13878.n29 gnd 1.53704f
C4425 a_n2804_13878.t26 gnd 0.194878f
C4426 a_n2982_13878.n0 gnd 3.88594f
C4427 a_n2982_13878.n1 gnd 2.85743f
C4428 a_n2982_13878.n2 gnd 3.82475f
C4429 a_n2982_13878.n3 gnd 0.806598f
C4430 a_n2982_13878.n4 gnd 0.8066f
C4431 a_n2982_13878.n5 gnd 0.916876f
C4432 a_n2982_13878.n6 gnd 0.201555f
C4433 a_n2982_13878.n7 gnd 0.148449f
C4434 a_n2982_13878.n8 gnd 0.233314f
C4435 a_n2982_13878.n9 gnd 0.180209f
C4436 a_n2982_13878.n10 gnd 0.201555f
C4437 a_n2982_13878.n11 gnd 1.34265f
C4438 a_n2982_13878.n12 gnd 0.148449f
C4439 a_n2982_13878.n13 gnd 0.969982f
C4440 a_n2982_13878.n14 gnd 0.212423f
C4441 a_n2982_13878.n15 gnd 0.747657f
C4442 a_n2982_13878.n16 gnd 0.212423f
C4443 a_n2982_13878.n17 gnd 0.212423f
C4444 a_n2982_13878.n18 gnd 0.483791f
C4445 a_n2982_13878.n19 gnd 0.278519f
C4446 a_n2982_13878.n20 gnd 0.212423f
C4447 a_n2982_13878.n21 gnd 0.536897f
C4448 a_n2982_13878.n22 gnd 0.212423f
C4449 a_n2982_13878.n23 gnd 0.212423f
C4450 a_n2982_13878.n24 gnd 0.945129f
C4451 a_n2982_13878.n25 gnd 0.278519f
C4452 a_n2982_13878.n26 gnd 0.985614f
C4453 a_n2982_13878.n27 gnd 0.212423f
C4454 a_n2982_13878.n28 gnd 0.212423f
C4455 a_n2982_13878.n29 gnd 0.483791f
C4456 a_n2982_13878.n30 gnd 0.212423f
C4457 a_n2982_13878.n31 gnd 0.278519f
C4458 a_n2982_13878.n32 gnd 3.26746f
C4459 a_n2982_13878.n33 gnd 0.278518f
C4460 a_n2982_13878.n34 gnd 0.106212f
C4461 a_n2982_13878.n35 gnd 0.212423f
C4462 a_n2982_13878.n36 gnd 0.85592f
C4463 a_n2982_13878.n37 gnd 0.212423f
C4464 a_n2982_13878.n38 gnd 0.278519f
C4465 a_n2982_13878.n39 gnd 1.74886f
C4466 a_n2982_13878.n40 gnd 1.17841f
C4467 a_n2982_13878.n41 gnd 2.35355f
C4468 a_n2982_13878.n42 gnd 1.17841f
C4469 a_n2982_13878.n43 gnd 2.1518f
C4470 a_n2982_13878.n44 gnd 1.74886f
C4471 a_n2982_13878.n45 gnd 0.008523f
C4472 a_n2982_13878.n46 gnd 4.11e-19
C4473 a_n2982_13878.n48 gnd 0.008224f
C4474 a_n2982_13878.n49 gnd 0.011959f
C4475 a_n2982_13878.n50 gnd 0.004385f
C4476 a_n2982_13878.n51 gnd 0.008523f
C4477 a_n2982_13878.n52 gnd 4.11e-19
C4478 a_n2982_13878.n54 gnd 0.008224f
C4479 a_n2982_13878.n55 gnd 0.011959f
C4480 a_n2982_13878.n56 gnd 0.007912f
C4481 a_n2982_13878.n58 gnd 0.28176f
C4482 a_n2982_13878.n59 gnd 0.008523f
C4483 a_n2982_13878.n60 gnd 4.11e-19
C4484 a_n2982_13878.n62 gnd 0.008224f
C4485 a_n2982_13878.n63 gnd 0.011959f
C4486 a_n2982_13878.n64 gnd 0.007912f
C4487 a_n2982_13878.n66 gnd 0.28176f
C4488 a_n2982_13878.n67 gnd 0.008523f
C4489 a_n2982_13878.n68 gnd 4.11e-19
C4490 a_n2982_13878.n70 gnd 0.008224f
C4491 a_n2982_13878.n71 gnd 0.011959f
C4492 a_n2982_13878.n72 gnd 0.007912f
C4493 a_n2982_13878.n74 gnd 0.28176f
C4494 a_n2982_13878.n75 gnd 0.008224f
C4495 a_n2982_13878.n76 gnd 0.280611f
C4496 a_n2982_13878.n77 gnd 0.008224f
C4497 a_n2982_13878.n78 gnd 0.280611f
C4498 a_n2982_13878.n79 gnd 0.008224f
C4499 a_n2982_13878.n80 gnd 0.280611f
C4500 a_n2982_13878.n81 gnd 0.008224f
C4501 a_n2982_13878.n82 gnd 0.280611f
C4502 a_n2982_13878.n83 gnd 0.301308f
C4503 a_n2982_13878.t11 gnd 0.147339f
C4504 a_n2982_13878.t44 gnd 0.699618f
C4505 a_n2982_13878.t6 gnd 0.68535f
C4506 a_n2982_13878.t10 gnd 0.68535f
C4507 a_n2982_13878.t46 gnd 0.68535f
C4508 a_n2982_13878.n84 gnd 0.301188f
C4509 a_n2982_13878.t24 gnd 0.68535f
C4510 a_n2982_13878.t48 gnd 0.68535f
C4511 a_n2982_13878.t52 gnd 0.68535f
C4512 a_n2982_13878.n85 gnd 0.297497f
C4513 a_n2982_13878.t16 gnd 0.68535f
C4514 a_n2982_13878.t12 gnd 0.68535f
C4515 a_n2982_13878.t50 gnd 0.68535f
C4516 a_n2982_13878.t18 gnd 0.699618f
C4517 a_n2982_13878.t110 gnd 0.699618f
C4518 a_n2982_13878.t87 gnd 0.68535f
C4519 a_n2982_13878.t92 gnd 0.68535f
C4520 a_n2982_13878.t80 gnd 0.68535f
C4521 a_n2982_13878.n86 gnd 0.301188f
C4522 a_n2982_13878.t97 gnd 0.68535f
C4523 a_n2982_13878.t106 gnd 0.68535f
C4524 a_n2982_13878.t107 gnd 0.68535f
C4525 a_n2982_13878.n87 gnd 0.297497f
C4526 a_n2982_13878.t74 gnd 0.68535f
C4527 a_n2982_13878.t89 gnd 0.68535f
C4528 a_n2982_13878.t77 gnd 0.68535f
C4529 a_n2982_13878.n88 gnd 0.301308f
C4530 a_n2982_13878.t84 gnd 0.68535f
C4531 a_n2982_13878.t103 gnd 0.696376f
C4532 a_n2982_13878.t9 gnd 1.37961f
C4533 a_n2982_13878.t27 gnd 0.147339f
C4534 a_n2982_13878.t37 gnd 0.147339f
C4535 a_n2982_13878.n89 gnd 1.03786f
C4536 a_n2982_13878.t15 gnd 0.147339f
C4537 a_n2982_13878.t23 gnd 0.147339f
C4538 a_n2982_13878.n90 gnd 1.03786f
C4539 a_n2982_13878.t21 gnd 0.147339f
C4540 a_n2982_13878.t39 gnd 0.147339f
C4541 a_n2982_13878.n91 gnd 1.03786f
C4542 a_n2982_13878.t41 gnd 0.147339f
C4543 a_n2982_13878.t31 gnd 0.147339f
C4544 a_n2982_13878.n92 gnd 1.03786f
C4545 a_n2982_13878.t35 gnd 0.147339f
C4546 a_n2982_13878.t43 gnd 0.147339f
C4547 a_n2982_13878.n93 gnd 1.03786f
C4548 a_n2982_13878.t29 gnd 1.37686f
C4549 a_n2982_13878.t34 gnd 0.68535f
C4550 a_n2982_13878.n94 gnd 0.301308f
C4551 a_n2982_13878.t42 gnd 0.68535f
C4552 a_n2982_13878.t40 gnd 0.68535f
C4553 a_n2982_13878.n95 gnd 0.292258f
C4554 a_n2982_13878.t22 gnd 0.68535f
C4555 a_n2982_13878.n96 gnd 0.303898f
C4556 a_n2982_13878.t20 gnd 0.68535f
C4557 a_n2982_13878.t36 gnd 0.68535f
C4558 a_n2982_13878.n97 gnd 0.297169f
C4559 a_n2982_13878.t8 gnd 0.699618f
C4560 a_n2982_13878.t86 gnd 0.68535f
C4561 a_n2982_13878.n98 gnd 0.301308f
C4562 a_n2982_13878.t95 gnd 0.68535f
C4563 a_n2982_13878.t101 gnd 0.68535f
C4564 a_n2982_13878.n99 gnd 0.292258f
C4565 a_n2982_13878.t105 gnd 0.68535f
C4566 a_n2982_13878.n100 gnd 0.303898f
C4567 a_n2982_13878.t76 gnd 0.68535f
C4568 a_n2982_13878.t79 gnd 0.68535f
C4569 a_n2982_13878.n101 gnd 0.297169f
C4570 a_n2982_13878.t109 gnd 0.699618f
C4571 a_n2982_13878.t78 gnd 0.68535f
C4572 a_n2982_13878.n102 gnd 0.303453f
C4573 a_n2982_13878.t104 gnd 0.68535f
C4574 a_n2982_13878.n103 gnd 0.301188f
C4575 a_n2982_13878.n104 gnd 0.301323f
C4576 a_n2982_13878.t100 gnd 0.68535f
C4577 a_n2982_13878.n105 gnd 0.297497f
C4578 a_n2982_13878.t73 gnd 0.68535f
C4579 a_n2982_13878.n106 gnd 0.297752f
C4580 a_n2982_13878.n107 gnd 0.303454f
C4581 a_n2982_13878.t75 gnd 0.696376f
C4582 a_n2982_13878.t26 gnd 0.68535f
C4583 a_n2982_13878.n108 gnd 0.303453f
C4584 a_n2982_13878.t14 gnd 0.68535f
C4585 a_n2982_13878.n109 gnd 0.301188f
C4586 a_n2982_13878.n110 gnd 0.301323f
C4587 a_n2982_13878.t38 gnd 0.68535f
C4588 a_n2982_13878.n111 gnd 0.297497f
C4589 a_n2982_13878.t30 gnd 0.68535f
C4590 a_n2982_13878.n112 gnd 0.297752f
C4591 a_n2982_13878.n113 gnd 0.303454f
C4592 a_n2982_13878.t28 gnd 0.696376f
C4593 a_n2982_13878.n114 gnd 1.32692f
C4594 a_n2982_13878.t83 gnd 0.68535f
C4595 a_n2982_13878.n115 gnd 0.297497f
C4596 a_n2982_13878.t91 gnd 0.68535f
C4597 a_n2982_13878.n116 gnd 0.297497f
C4598 a_n2982_13878.t81 gnd 0.68535f
C4599 a_n2982_13878.n117 gnd 0.297497f
C4600 a_n2982_13878.t96 gnd 0.68535f
C4601 a_n2982_13878.n118 gnd 0.297497f
C4602 a_n2982_13878.t85 gnd 0.68535f
C4603 a_n2982_13878.n119 gnd 0.292094f
C4604 a_n2982_13878.t111 gnd 0.68535f
C4605 a_n2982_13878.n120 gnd 0.301323f
C4606 a_n2982_13878.t88 gnd 0.696834f
C4607 a_n2982_13878.t98 gnd 0.68535f
C4608 a_n2982_13878.n121 gnd 0.292094f
C4609 a_n2982_13878.t82 gnd 0.68535f
C4610 a_n2982_13878.n122 gnd 0.301323f
C4611 a_n2982_13878.t93 gnd 0.696834f
C4612 a_n2982_13878.t102 gnd 0.68535f
C4613 a_n2982_13878.n123 gnd 0.292094f
C4614 a_n2982_13878.t90 gnd 0.68535f
C4615 a_n2982_13878.n124 gnd 0.301323f
C4616 a_n2982_13878.t108 gnd 0.696834f
C4617 a_n2982_13878.t94 gnd 0.68535f
C4618 a_n2982_13878.n125 gnd 0.292094f
C4619 a_n2982_13878.t72 gnd 0.68535f
C4620 a_n2982_13878.n126 gnd 0.301323f
C4621 a_n2982_13878.t99 gnd 0.696834f
C4622 a_n2982_13878.n127 gnd 1.6691f
C4623 a_n2982_13878.n128 gnd 0.303454f
C4624 a_n2982_13878.n129 gnd 0.297752f
C4625 a_n2982_13878.n130 gnd 0.292258f
C4626 a_n2982_13878.n131 gnd 0.301323f
C4627 a_n2982_13878.n132 gnd 0.303898f
C4628 a_n2982_13878.n133 gnd 0.297169f
C4629 a_n2982_13878.n134 gnd 0.303453f
C4630 a_n2982_13878.t32 gnd 0.68535f
C4631 a_n2982_13878.n135 gnd 0.303454f
C4632 a_n2982_13878.t3 gnd 0.114597f
C4633 a_n2982_13878.t67 gnd 0.114597f
C4634 a_n2982_13878.n136 gnd 1.01487f
C4635 a_n2982_13878.t68 gnd 0.114597f
C4636 a_n2982_13878.t69 gnd 0.114597f
C4637 a_n2982_13878.n137 gnd 1.01262f
C4638 a_n2982_13878.t63 gnd 0.114597f
C4639 a_n2982_13878.t58 gnd 0.114597f
C4640 a_n2982_13878.n138 gnd 1.01262f
C4641 a_n2982_13878.t60 gnd 0.114597f
C4642 a_n2982_13878.t66 gnd 0.114597f
C4643 a_n2982_13878.n139 gnd 1.01487f
C4644 a_n2982_13878.t62 gnd 0.114597f
C4645 a_n2982_13878.t4 gnd 0.114597f
C4646 a_n2982_13878.n140 gnd 1.01262f
C4647 a_n2982_13878.t5 gnd 0.114597f
C4648 a_n2982_13878.t56 gnd 0.114597f
C4649 a_n2982_13878.n141 gnd 1.01262f
C4650 a_n2982_13878.t57 gnd 0.114597f
C4651 a_n2982_13878.t59 gnd 0.114597f
C4652 a_n2982_13878.n142 gnd 1.01262f
C4653 a_n2982_13878.t2 gnd 0.114597f
C4654 a_n2982_13878.t71 gnd 0.114597f
C4655 a_n2982_13878.n143 gnd 1.01262f
C4656 a_n2982_13878.t61 gnd 0.114597f
C4657 a_n2982_13878.t54 gnd 0.114597f
C4658 a_n2982_13878.n144 gnd 1.01262f
C4659 a_n2982_13878.t1 gnd 0.114597f
C4660 a_n2982_13878.t70 gnd 0.114597f
C4661 a_n2982_13878.n145 gnd 1.01487f
C4662 a_n2982_13878.t55 gnd 0.114597f
C4663 a_n2982_13878.t65 gnd 0.114597f
C4664 a_n2982_13878.n146 gnd 1.01262f
C4665 a_n2982_13878.t64 gnd 0.114597f
C4666 a_n2982_13878.t0 gnd 0.114597f
C4667 a_n2982_13878.n147 gnd 1.01262f
C4668 a_n2982_13878.n148 gnd 0.30128f
C4669 a_n2982_13878.n149 gnd 0.292258f
C4670 a_n2982_13878.n150 gnd 0.301323f
C4671 a_n2982_13878.n151 gnd 0.303898f
C4672 a_n2982_13878.n152 gnd 0.297169f
C4673 a_n2982_13878.n153 gnd 0.303453f
C4674 a_n2982_13878.n154 gnd 1.00893f
C4675 a_n2982_13878.t45 gnd 1.37686f
C4676 a_n2982_13878.t19 gnd 1.37961f
C4677 a_n2982_13878.t51 gnd 0.147339f
C4678 a_n2982_13878.t33 gnd 0.147339f
C4679 a_n2982_13878.n155 gnd 1.03786f
C4680 a_n2982_13878.t17 gnd 0.147339f
C4681 a_n2982_13878.t13 gnd 0.147339f
C4682 a_n2982_13878.n156 gnd 1.03786f
C4683 a_n2982_13878.t49 gnd 0.147339f
C4684 a_n2982_13878.t53 gnd 0.147339f
C4685 a_n2982_13878.n157 gnd 1.03786f
C4686 a_n2982_13878.t47 gnd 0.147339f
C4687 a_n2982_13878.t25 gnd 0.147339f
C4688 a_n2982_13878.n158 gnd 1.03786f
C4689 a_n2982_13878.n159 gnd 1.03786f
C4690 a_n2982_13878.t7 gnd 0.147339f
C4691 a_n7636_8799.t23 gnd 0.114884f
C4692 a_n7636_8799.t13 gnd 0.114884f
C4693 a_n7636_8799.t12 gnd 0.114884f
C4694 a_n7636_8799.n0 gnd 1.01741f
C4695 a_n7636_8799.t18 gnd 0.114884f
C4696 a_n7636_8799.t17 gnd 0.114884f
C4697 a_n7636_8799.n1 gnd 1.01515f
C4698 a_n7636_8799.n2 gnd 0.808618f
C4699 a_n7636_8799.t47 gnd 0.147708f
C4700 a_n7636_8799.t3 gnd 0.147708f
C4701 a_n7636_8799.n3 gnd 1.16499f
C4702 a_n7636_8799.t4 gnd 0.147708f
C4703 a_n7636_8799.t32 gnd 0.147708f
C4704 a_n7636_8799.n4 gnd 1.16307f
C4705 a_n7636_8799.n5 gnd 1.04546f
C4706 a_n7636_8799.t31 gnd 0.147708f
C4707 a_n7636_8799.t46 gnd 0.147708f
C4708 a_n7636_8799.n6 gnd 1.16307f
C4709 a_n7636_8799.n7 gnd 0.515326f
C4710 a_n7636_8799.t39 gnd 0.147708f
C4711 a_n7636_8799.t2 gnd 0.147708f
C4712 a_n7636_8799.n8 gnd 1.16307f
C4713 a_n7636_8799.n9 gnd 0.515326f
C4714 a_n7636_8799.t42 gnd 0.147708f
C4715 a_n7636_8799.t30 gnd 0.147708f
C4716 a_n7636_8799.n10 gnd 1.16307f
C4717 a_n7636_8799.n11 gnd 0.515326f
C4718 a_n7636_8799.t34 gnd 0.147708f
C4719 a_n7636_8799.t40 gnd 0.147708f
C4720 a_n7636_8799.n12 gnd 1.16307f
C4721 a_n7636_8799.n13 gnd 3.80462f
C4722 a_n7636_8799.t5 gnd 0.147708f
C4723 a_n7636_8799.t44 gnd 0.147708f
C4724 a_n7636_8799.n14 gnd 1.16499f
C4725 a_n7636_8799.t41 gnd 0.147708f
C4726 a_n7636_8799.t35 gnd 0.147708f
C4727 a_n7636_8799.n15 gnd 1.16307f
C4728 a_n7636_8799.n16 gnd 1.04546f
C4729 a_n7636_8799.t38 gnd 0.147708f
C4730 a_n7636_8799.t1 gnd 0.147708f
C4731 a_n7636_8799.n17 gnd 1.16307f
C4732 a_n7636_8799.n18 gnd 0.515326f
C4733 a_n7636_8799.t37 gnd 0.147708f
C4734 a_n7636_8799.t45 gnd 0.147708f
C4735 a_n7636_8799.n19 gnd 1.16307f
C4736 a_n7636_8799.n20 gnd 0.515326f
C4737 a_n7636_8799.t0 gnd 0.147708f
C4738 a_n7636_8799.t36 gnd 0.147708f
C4739 a_n7636_8799.n21 gnd 1.16307f
C4740 a_n7636_8799.n22 gnd 0.515326f
C4741 a_n7636_8799.t43 gnd 0.147708f
C4742 a_n7636_8799.t33 gnd 0.147708f
C4743 a_n7636_8799.n23 gnd 1.16307f
C4744 a_n7636_8799.n24 gnd 2.54343f
C4745 a_n7636_8799.n25 gnd 7.813859f
C4746 a_n7636_8799.n26 gnd 0.053239f
C4747 a_n7636_8799.t64 gnd 0.612465f
C4748 a_n7636_8799.n27 gnd 0.273539f
C4749 a_n7636_8799.n28 gnd 0.053239f
C4750 a_n7636_8799.n29 gnd 0.012081f
C4751 a_n7636_8799.t78 gnd 0.612465f
C4752 a_n7636_8799.n30 gnd 0.169503f
C4753 a_n7636_8799.t88 gnd 0.612465f
C4754 a_n7636_8799.t87 gnd 0.624057f
C4755 a_n7636_8799.n31 gnd 0.256755f
C4756 a_n7636_8799.n32 gnd 0.27042f
C4757 a_n7636_8799.n33 gnd 0.012081f
C4758 a_n7636_8799.t66 gnd 0.612465f
C4759 a_n7636_8799.n34 gnd 0.273539f
C4760 a_n7636_8799.n35 gnd 0.053239f
C4761 a_n7636_8799.n36 gnd 0.053239f
C4762 a_n7636_8799.n37 gnd 0.053239f
C4763 a_n7636_8799.n38 gnd 0.270749f
C4764 a_n7636_8799.t86 gnd 0.612465f
C4765 a_n7636_8799.n39 gnd 0.270749f
C4766 a_n7636_8799.n40 gnd 0.012081f
C4767 a_n7636_8799.n41 gnd 0.053239f
C4768 a_n7636_8799.n42 gnd 0.053239f
C4769 a_n7636_8799.n43 gnd 0.053239f
C4770 a_n7636_8799.n44 gnd 0.012081f
C4771 a_n7636_8799.t65 gnd 0.612465f
C4772 a_n7636_8799.n45 gnd 0.27042f
C4773 a_n7636_8799.t77 gnd 0.612465f
C4774 a_n7636_8799.n46 gnd 0.267958f
C4775 a_n7636_8799.n47 gnd 0.30294f
C4776 a_n7636_8799.n48 gnd 0.053239f
C4777 a_n7636_8799.t69 gnd 0.612465f
C4778 a_n7636_8799.n49 gnd 0.273539f
C4779 a_n7636_8799.n50 gnd 0.053239f
C4780 a_n7636_8799.n51 gnd 0.012081f
C4781 a_n7636_8799.t83 gnd 0.612465f
C4782 a_n7636_8799.n52 gnd 0.169503f
C4783 a_n7636_8799.t95 gnd 0.612465f
C4784 a_n7636_8799.t94 gnd 0.624057f
C4785 a_n7636_8799.n53 gnd 0.256755f
C4786 a_n7636_8799.n54 gnd 0.27042f
C4787 a_n7636_8799.n55 gnd 0.012081f
C4788 a_n7636_8799.t71 gnd 0.612465f
C4789 a_n7636_8799.n56 gnd 0.273539f
C4790 a_n7636_8799.n57 gnd 0.053239f
C4791 a_n7636_8799.n58 gnd 0.053239f
C4792 a_n7636_8799.n59 gnd 0.053239f
C4793 a_n7636_8799.n60 gnd 0.270749f
C4794 a_n7636_8799.t93 gnd 0.612465f
C4795 a_n7636_8799.n61 gnd 0.270749f
C4796 a_n7636_8799.n62 gnd 0.012081f
C4797 a_n7636_8799.n63 gnd 0.053239f
C4798 a_n7636_8799.n64 gnd 0.053239f
C4799 a_n7636_8799.n65 gnd 0.053239f
C4800 a_n7636_8799.n66 gnd 0.012081f
C4801 a_n7636_8799.t70 gnd 0.612465f
C4802 a_n7636_8799.n67 gnd 0.27042f
C4803 a_n7636_8799.t81 gnd 0.612465f
C4804 a_n7636_8799.n68 gnd 0.267958f
C4805 a_n7636_8799.n69 gnd 0.133864f
C4806 a_n7636_8799.n70 gnd 0.921126f
C4807 a_n7636_8799.n71 gnd 0.053239f
C4808 a_n7636_8799.t54 gnd 0.612465f
C4809 a_n7636_8799.n72 gnd 0.273539f
C4810 a_n7636_8799.n73 gnd 0.053239f
C4811 a_n7636_8799.n74 gnd 0.012081f
C4812 a_n7636_8799.t62 gnd 0.612465f
C4813 a_n7636_8799.n75 gnd 0.169503f
C4814 a_n7636_8799.t68 gnd 0.612465f
C4815 a_n7636_8799.t75 gnd 0.624057f
C4816 a_n7636_8799.n76 gnd 0.256755f
C4817 a_n7636_8799.n77 gnd 0.27042f
C4818 a_n7636_8799.n78 gnd 0.012081f
C4819 a_n7636_8799.t82 gnd 0.612465f
C4820 a_n7636_8799.n79 gnd 0.273539f
C4821 a_n7636_8799.n80 gnd 0.053239f
C4822 a_n7636_8799.n81 gnd 0.053239f
C4823 a_n7636_8799.n82 gnd 0.053239f
C4824 a_n7636_8799.n83 gnd 0.270749f
C4825 a_n7636_8799.t89 gnd 0.612465f
C4826 a_n7636_8799.n84 gnd 0.270749f
C4827 a_n7636_8799.n85 gnd 0.012081f
C4828 a_n7636_8799.n86 gnd 0.053239f
C4829 a_n7636_8799.n87 gnd 0.053239f
C4830 a_n7636_8799.n88 gnd 0.053239f
C4831 a_n7636_8799.n89 gnd 0.012081f
C4832 a_n7636_8799.t48 gnd 0.612465f
C4833 a_n7636_8799.n90 gnd 0.27042f
C4834 a_n7636_8799.t72 gnd 0.612465f
C4835 a_n7636_8799.n91 gnd 0.267958f
C4836 a_n7636_8799.n92 gnd 0.133864f
C4837 a_n7636_8799.n93 gnd 1.946f
C4838 a_n7636_8799.n94 gnd 0.053239f
C4839 a_n7636_8799.t50 gnd 0.612465f
C4840 a_n7636_8799.t49 gnd 0.612465f
C4841 a_n7636_8799.t80 gnd 0.612465f
C4842 a_n7636_8799.n95 gnd 0.273539f
C4843 a_n7636_8799.n96 gnd 0.053239f
C4844 a_n7636_8799.t57 gnd 0.612465f
C4845 a_n7636_8799.t51 gnd 0.612465f
C4846 a_n7636_8799.n97 gnd 0.053239f
C4847 a_n7636_8799.t84 gnd 0.612465f
C4848 a_n7636_8799.n98 gnd 0.273539f
C4849 a_n7636_8799.t58 gnd 0.624057f
C4850 a_n7636_8799.n99 gnd 0.256755f
C4851 a_n7636_8799.t67 gnd 0.612465f
C4852 a_n7636_8799.n100 gnd 0.27042f
C4853 a_n7636_8799.n101 gnd 0.012081f
C4854 a_n7636_8799.n102 gnd 0.169503f
C4855 a_n7636_8799.n103 gnd 0.053239f
C4856 a_n7636_8799.n104 gnd 0.053239f
C4857 a_n7636_8799.n105 gnd 0.012081f
C4858 a_n7636_8799.n106 gnd 0.270749f
C4859 a_n7636_8799.n107 gnd 0.270749f
C4860 a_n7636_8799.n108 gnd 0.012081f
C4861 a_n7636_8799.n109 gnd 0.053239f
C4862 a_n7636_8799.n110 gnd 0.053239f
C4863 a_n7636_8799.n111 gnd 0.053239f
C4864 a_n7636_8799.n112 gnd 0.012081f
C4865 a_n7636_8799.n113 gnd 0.27042f
C4866 a_n7636_8799.n114 gnd 0.267958f
C4867 a_n7636_8799.n115 gnd 0.30294f
C4868 a_n7636_8799.n116 gnd 0.053239f
C4869 a_n7636_8799.t53 gnd 0.612465f
C4870 a_n7636_8799.t52 gnd 0.612465f
C4871 a_n7636_8799.t91 gnd 0.612465f
C4872 a_n7636_8799.n117 gnd 0.273539f
C4873 a_n7636_8799.n118 gnd 0.053239f
C4874 a_n7636_8799.t60 gnd 0.612465f
C4875 a_n7636_8799.t56 gnd 0.612465f
C4876 a_n7636_8799.n119 gnd 0.053239f
C4877 a_n7636_8799.t92 gnd 0.612465f
C4878 a_n7636_8799.n120 gnd 0.273539f
C4879 a_n7636_8799.t61 gnd 0.624057f
C4880 a_n7636_8799.n121 gnd 0.256755f
C4881 a_n7636_8799.t74 gnd 0.612465f
C4882 a_n7636_8799.n122 gnd 0.27042f
C4883 a_n7636_8799.n123 gnd 0.012081f
C4884 a_n7636_8799.n124 gnd 0.169503f
C4885 a_n7636_8799.n125 gnd 0.053239f
C4886 a_n7636_8799.n126 gnd 0.053239f
C4887 a_n7636_8799.n127 gnd 0.012081f
C4888 a_n7636_8799.n128 gnd 0.270749f
C4889 a_n7636_8799.n129 gnd 0.270749f
C4890 a_n7636_8799.n130 gnd 0.012081f
C4891 a_n7636_8799.n131 gnd 0.053239f
C4892 a_n7636_8799.n132 gnd 0.053239f
C4893 a_n7636_8799.n133 gnd 0.053239f
C4894 a_n7636_8799.n134 gnd 0.012081f
C4895 a_n7636_8799.n135 gnd 0.27042f
C4896 a_n7636_8799.n136 gnd 0.267958f
C4897 a_n7636_8799.n137 gnd 0.133864f
C4898 a_n7636_8799.n138 gnd 0.921126f
C4899 a_n7636_8799.n139 gnd 0.053239f
C4900 a_n7636_8799.t73 gnd 0.612465f
C4901 a_n7636_8799.t79 gnd 0.612465f
C4902 a_n7636_8799.t55 gnd 0.612465f
C4903 a_n7636_8799.n140 gnd 0.273539f
C4904 a_n7636_8799.n141 gnd 0.053239f
C4905 a_n7636_8799.t90 gnd 0.612465f
C4906 a_n7636_8799.t63 gnd 0.612465f
C4907 a_n7636_8799.n142 gnd 0.053239f
C4908 a_n7636_8799.t85 gnd 0.612465f
C4909 a_n7636_8799.n143 gnd 0.273539f
C4910 a_n7636_8799.t76 gnd 0.624057f
C4911 a_n7636_8799.n144 gnd 0.256755f
C4912 a_n7636_8799.t59 gnd 0.612465f
C4913 a_n7636_8799.n145 gnd 0.27042f
C4914 a_n7636_8799.n146 gnd 0.012081f
C4915 a_n7636_8799.n147 gnd 0.169503f
C4916 a_n7636_8799.n148 gnd 0.053239f
C4917 a_n7636_8799.n149 gnd 0.053239f
C4918 a_n7636_8799.n150 gnd 0.012081f
C4919 a_n7636_8799.n151 gnd 0.270749f
C4920 a_n7636_8799.n152 gnd 0.270749f
C4921 a_n7636_8799.n153 gnd 0.012081f
C4922 a_n7636_8799.n154 gnd 0.053239f
C4923 a_n7636_8799.n155 gnd 0.053239f
C4924 a_n7636_8799.n156 gnd 0.053239f
C4925 a_n7636_8799.n157 gnd 0.012081f
C4926 a_n7636_8799.n158 gnd 0.27042f
C4927 a_n7636_8799.n159 gnd 0.267958f
C4928 a_n7636_8799.n160 gnd 0.133864f
C4929 a_n7636_8799.n161 gnd 1.41081f
C4930 a_n7636_8799.n162 gnd 17.7867f
C4931 a_n7636_8799.n163 gnd 4.48235f
C4932 a_n7636_8799.t14 gnd 0.114884f
C4933 a_n7636_8799.t15 gnd 0.114884f
C4934 a_n7636_8799.n164 gnd 1.01741f
C4935 a_n7636_8799.t8 gnd 0.114884f
C4936 a_n7636_8799.t9 gnd 0.114884f
C4937 a_n7636_8799.n165 gnd 1.01515f
C4938 a_n7636_8799.n166 gnd 0.808616f
C4939 a_n7636_8799.t7 gnd 0.114884f
C4940 a_n7636_8799.t25 gnd 0.114884f
C4941 a_n7636_8799.n167 gnd 1.01515f
C4942 a_n7636_8799.n168 gnd 0.33765f
C4943 a_n7636_8799.n169 gnd 0.482056f
C4944 a_n7636_8799.t27 gnd 0.114884f
C4945 a_n7636_8799.t20 gnd 0.114884f
C4946 a_n7636_8799.n170 gnd 1.01515f
C4947 a_n7636_8799.n171 gnd 0.33765f
C4948 a_n7636_8799.t22 gnd 0.114884f
C4949 a_n7636_8799.t6 gnd 0.114884f
C4950 a_n7636_8799.n172 gnd 1.01515f
C4951 a_n7636_8799.n173 gnd 0.397072f
C4952 a_n7636_8799.t24 gnd 0.114884f
C4953 a_n7636_8799.t26 gnd 0.114884f
C4954 a_n7636_8799.n174 gnd 1.01515f
C4955 a_n7636_8799.n175 gnd 2.92329f
C4956 a_n7636_8799.t21 gnd 0.114884f
C4957 a_n7636_8799.t19 gnd 0.114884f
C4958 a_n7636_8799.n176 gnd 1.01741f
C4959 a_n7636_8799.t10 gnd 0.114884f
C4960 a_n7636_8799.t16 gnd 0.114884f
C4961 a_n7636_8799.n177 gnd 1.01515f
C4962 a_n7636_8799.n178 gnd 0.808618f
C4963 a_n7636_8799.t28 gnd 0.114884f
C4964 a_n7636_8799.t11 gnd 0.114884f
C4965 a_n7636_8799.n179 gnd 1.01515f
C4966 a_n7636_8799.n180 gnd 0.337651f
C4967 a_n7636_8799.n181 gnd 2.46037f
C4968 a_n7636_8799.n182 gnd 0.337654f
C4969 a_n7636_8799.n183 gnd 1.01515f
C4970 a_n7636_8799.t29 gnd 0.114884f
C4971 a_n3827_n3924.n0 gnd 1.99733f
C4972 a_n3827_n3924.n1 gnd 2.17486f
C4973 a_n3827_n3924.n2 gnd 1.44807f
C4974 a_n3827_n3924.n3 gnd 1.31657f
C4975 a_n3827_n3924.n4 gnd 1.81285f
C4976 a_n3827_n3924.n5 gnd 3.90473f
C4977 a_n3827_n3924.n6 gnd 0.724032f
C4978 a_n3827_n3924.n7 gnd 1.77302f
C4979 a_n3827_n3924.n8 gnd 0.886511f
C4980 a_n3827_n3924.n9 gnd 2.49022f
C4981 a_n3827_n3924.n10 gnd 0.954549f
C4982 a_n3827_n3924.n11 gnd 1.2733f
C4983 a_n3827_n3924.t32 gnd 0.097472f
C4984 a_n3827_n3924.t31 gnd 0.097472f
C4985 a_n3827_n3924.t43 gnd 0.097472f
C4986 a_n3827_n3924.n12 gnd 0.796069f
C4987 a_n3827_n3924.t52 gnd 1.26084f
C4988 a_n3827_n3924.t56 gnd 0.097472f
C4989 a_n3827_n3924.t38 gnd 0.097472f
C4990 a_n3827_n3924.n13 gnd 0.796069f
C4991 a_n3827_n3924.t36 gnd 0.097472f
C4992 a_n3827_n3924.t2 gnd 0.097472f
C4993 a_n3827_n3924.n14 gnd 0.796069f
C4994 a_n3827_n3924.t34 gnd 1.01304f
C4995 a_n3827_n3924.t45 gnd 1.26048f
C4996 a_n3827_n3924.t54 gnd 1.25868f
C4997 a_n3827_n3924.t57 gnd 1.25868f
C4998 a_n3827_n3924.t4 gnd 1.25868f
C4999 a_n3827_n3924.t53 gnd 1.25868f
C5000 a_n3827_n3924.t41 gnd 1.25868f
C5001 a_n3827_n3924.t49 gnd 1.25868f
C5002 a_n3827_n3924.t48 gnd 1.25868f
C5003 a_n3827_n3924.t42 gnd 1.25868f
C5004 a_n3827_n3924.n15 gnd 0.914318f
C5005 a_n3827_n3924.t12 gnd 1.01304f
C5006 a_n3827_n3924.t24 gnd 0.097472f
C5007 a_n3827_n3924.t27 gnd 0.097472f
C5008 a_n3827_n3924.n16 gnd 0.796068f
C5009 a_n3827_n3924.t18 gnd 0.097472f
C5010 a_n3827_n3924.t17 gnd 0.097472f
C5011 a_n3827_n3924.n17 gnd 0.796068f
C5012 a_n3827_n3924.t8 gnd 0.097472f
C5013 a_n3827_n3924.t14 gnd 0.097472f
C5014 a_n3827_n3924.n18 gnd 0.796068f
C5015 a_n3827_n3924.t22 gnd 0.097472f
C5016 a_n3827_n3924.t19 gnd 0.097472f
C5017 a_n3827_n3924.n19 gnd 0.796068f
C5018 a_n3827_n3924.t26 gnd 0.097472f
C5019 a_n3827_n3924.t28 gnd 0.097472f
C5020 a_n3827_n3924.n20 gnd 0.796068f
C5021 a_n3827_n3924.t15 gnd 1.01304f
C5022 a_n3827_n3924.t3 gnd 1.01304f
C5023 a_n3827_n3924.t47 gnd 0.097472f
C5024 a_n3827_n3924.t50 gnd 0.097472f
C5025 a_n3827_n3924.n21 gnd 0.796068f
C5026 a_n3827_n3924.t51 gnd 0.097472f
C5027 a_n3827_n3924.t40 gnd 0.097472f
C5028 a_n3827_n3924.n22 gnd 0.796068f
C5029 a_n3827_n3924.t35 gnd 0.097472f
C5030 a_n3827_n3924.t30 gnd 0.097472f
C5031 a_n3827_n3924.n23 gnd 0.796068f
C5032 a_n3827_n3924.t33 gnd 0.097472f
C5033 a_n3827_n3924.t39 gnd 0.097472f
C5034 a_n3827_n3924.n24 gnd 0.796068f
C5035 a_n3827_n3924.t29 gnd 0.097472f
C5036 a_n3827_n3924.t37 gnd 0.097472f
C5037 a_n3827_n3924.n25 gnd 0.796068f
C5038 a_n3827_n3924.t46 gnd 1.01304f
C5039 a_n3827_n3924.n26 gnd 0.914318f
C5040 a_n3827_n3924.t11 gnd 1.01304f
C5041 a_n3827_n3924.t6 gnd 0.097472f
C5042 a_n3827_n3924.t20 gnd 0.097472f
C5043 a_n3827_n3924.n27 gnd 0.796069f
C5044 a_n3827_n3924.t25 gnd 0.097472f
C5045 a_n3827_n3924.t10 gnd 0.097472f
C5046 a_n3827_n3924.n28 gnd 0.796069f
C5047 a_n3827_n3924.t23 gnd 0.097472f
C5048 a_n3827_n3924.t16 gnd 0.097472f
C5049 a_n3827_n3924.n29 gnd 0.796069f
C5050 a_n3827_n3924.t9 gnd 0.097472f
C5051 a_n3827_n3924.t13 gnd 0.097472f
C5052 a_n3827_n3924.n30 gnd 0.796069f
C5053 a_n3827_n3924.t7 gnd 0.097472f
C5054 a_n3827_n3924.t5 gnd 0.097472f
C5055 a_n3827_n3924.n31 gnd 0.796069f
C5056 a_n3827_n3924.t21 gnd 1.01304f
C5057 a_n3827_n3924.t55 gnd 1.01304f
C5058 a_n3827_n3924.t44 gnd 0.097472f
C5059 a_n3827_n3924.t1 gnd 0.097472f
C5060 a_n3827_n3924.n32 gnd 0.796069f
C5061 a_n3827_n3924.n33 gnd 0.79607f
C5062 a_n3827_n3924.t0 gnd 0.097472f
C5063 plus.n0 gnd 0.023071f
C5064 plus.t21 gnd 0.326322f
C5065 plus.n1 gnd 0.023071f
C5066 plus.t22 gnd 0.326322f
C5067 plus.t16 gnd 0.326322f
C5068 plus.n2 gnd 0.144963f
C5069 plus.n3 gnd 0.023071f
C5070 plus.t17 gnd 0.326322f
C5071 plus.t11 gnd 0.326322f
C5072 plus.n4 gnd 0.144963f
C5073 plus.n5 gnd 0.023071f
C5074 plus.t5 gnd 0.326322f
C5075 plus.t6 gnd 0.326322f
C5076 plus.n6 gnd 0.144963f
C5077 plus.n7 gnd 0.023071f
C5078 plus.t23 gnd 0.326322f
C5079 plus.t24 gnd 0.326322f
C5080 plus.n8 gnd 0.144963f
C5081 plus.n9 gnd 0.023071f
C5082 plus.t18 gnd 0.326322f
C5083 plus.t13 gnd 0.326322f
C5084 plus.n10 gnd 0.149684f
C5085 plus.t15 gnd 0.338168f
C5086 plus.n11 gnd 0.134346f
C5087 plus.n12 gnd 0.099323f
C5088 plus.n13 gnd 0.005235f
C5089 plus.n14 gnd 0.144963f
C5090 plus.n15 gnd 0.005235f
C5091 plus.n16 gnd 0.023071f
C5092 plus.n17 gnd 0.023071f
C5093 plus.n18 gnd 0.023071f
C5094 plus.n19 gnd 0.005235f
C5095 plus.n20 gnd 0.144963f
C5096 plus.n21 gnd 0.005235f
C5097 plus.n22 gnd 0.023071f
C5098 plus.n23 gnd 0.023071f
C5099 plus.n24 gnd 0.023071f
C5100 plus.n25 gnd 0.005235f
C5101 plus.n26 gnd 0.144963f
C5102 plus.n27 gnd 0.005235f
C5103 plus.n28 gnd 0.023071f
C5104 plus.n29 gnd 0.023071f
C5105 plus.n30 gnd 0.023071f
C5106 plus.n31 gnd 0.005235f
C5107 plus.n32 gnd 0.144963f
C5108 plus.n33 gnd 0.005235f
C5109 plus.n34 gnd 0.023071f
C5110 plus.n35 gnd 0.023071f
C5111 plus.n36 gnd 0.023071f
C5112 plus.n37 gnd 0.005235f
C5113 plus.n38 gnd 0.144963f
C5114 plus.n39 gnd 0.005235f
C5115 plus.n40 gnd 0.145176f
C5116 plus.n41 gnd 0.261247f
C5117 plus.n42 gnd 0.023071f
C5118 plus.n43 gnd 0.005235f
C5119 plus.t10 gnd 0.326322f
C5120 plus.n44 gnd 0.023071f
C5121 plus.n45 gnd 0.005235f
C5122 plus.t12 gnd 0.326322f
C5123 plus.n46 gnd 0.023071f
C5124 plus.n47 gnd 0.005235f
C5125 plus.t7 gnd 0.326322f
C5126 plus.n48 gnd 0.023071f
C5127 plus.n49 gnd 0.005235f
C5128 plus.t27 gnd 0.326322f
C5129 plus.n50 gnd 0.023071f
C5130 plus.n51 gnd 0.005235f
C5131 plus.t26 gnd 0.326322f
C5132 plus.t20 gnd 0.338168f
C5133 plus.t19 gnd 0.326322f
C5134 plus.n52 gnd 0.149684f
C5135 plus.n53 gnd 0.134346f
C5136 plus.n54 gnd 0.099323f
C5137 plus.n55 gnd 0.023071f
C5138 plus.n56 gnd 0.144963f
C5139 plus.n57 gnd 0.005235f
C5140 plus.t25 gnd 0.326322f
C5141 plus.n58 gnd 0.144963f
C5142 plus.n59 gnd 0.023071f
C5143 plus.n60 gnd 0.023071f
C5144 plus.n61 gnd 0.023071f
C5145 plus.n62 gnd 0.144963f
C5146 plus.n63 gnd 0.005235f
C5147 plus.t9 gnd 0.326322f
C5148 plus.n64 gnd 0.144963f
C5149 plus.n65 gnd 0.023071f
C5150 plus.n66 gnd 0.023071f
C5151 plus.n67 gnd 0.023071f
C5152 plus.n68 gnd 0.144963f
C5153 plus.n69 gnd 0.005235f
C5154 plus.t14 gnd 0.326322f
C5155 plus.n70 gnd 0.144963f
C5156 plus.n71 gnd 0.023071f
C5157 plus.n72 gnd 0.023071f
C5158 plus.n73 gnd 0.023071f
C5159 plus.n74 gnd 0.144963f
C5160 plus.n75 gnd 0.005235f
C5161 plus.t28 gnd 0.326322f
C5162 plus.n76 gnd 0.144963f
C5163 plus.n77 gnd 0.023071f
C5164 plus.n78 gnd 0.023071f
C5165 plus.n79 gnd 0.023071f
C5166 plus.n80 gnd 0.144963f
C5167 plus.n81 gnd 0.005235f
C5168 plus.t8 gnd 0.326322f
C5169 plus.n82 gnd 0.145176f
C5170 plus.n83 gnd 0.763663f
C5171 plus.n84 gnd 1.14249f
C5172 plus.t2 gnd 0.039828f
C5173 plus.t3 gnd 0.007112f
C5174 plus.t1 gnd 0.007112f
C5175 plus.n85 gnd 0.023066f
C5176 plus.n86 gnd 0.179065f
C5177 plus.t4 gnd 0.007112f
C5178 plus.t0 gnd 0.007112f
C5179 plus.n87 gnd 0.023066f
C5180 plus.n88 gnd 0.13441f
C5181 plus.n89 gnd 3.15838f
C5182 commonsourceibias.n0 gnd 0.012818f
C5183 commonsourceibias.t104 gnd 0.19409f
C5184 commonsourceibias.t181 gnd 0.179464f
C5185 commonsourceibias.n1 gnd 0.00935f
C5186 commonsourceibias.n2 gnd 0.009606f
C5187 commonsourceibias.t124 gnd 0.179464f
C5188 commonsourceibias.n3 gnd 0.012358f
C5189 commonsourceibias.n4 gnd 0.009606f
C5190 commonsourceibias.t197 gnd 0.179464f
C5191 commonsourceibias.n5 gnd 0.071606f
C5192 commonsourceibias.t142 gnd 0.179464f
C5193 commonsourceibias.n6 gnd 0.009057f
C5194 commonsourceibias.n7 gnd 0.009606f
C5195 commonsourceibias.t101 gnd 0.179464f
C5196 commonsourceibias.n8 gnd 0.012175f
C5197 commonsourceibias.n9 gnd 0.009606f
C5198 commonsourceibias.t156 gnd 0.179464f
C5199 commonsourceibias.n10 gnd 0.071606f
C5200 commonsourceibias.t143 gnd 0.179464f
C5201 commonsourceibias.n11 gnd 0.008798f
C5202 commonsourceibias.n12 gnd 0.009606f
C5203 commonsourceibias.t193 gnd 0.179464f
C5204 commonsourceibias.n13 gnd 0.01197f
C5205 commonsourceibias.n14 gnd 0.012818f
C5206 commonsourceibias.t72 gnd 0.19409f
C5207 commonsourceibias.t54 gnd 0.179464f
C5208 commonsourceibias.n15 gnd 0.00935f
C5209 commonsourceibias.n16 gnd 0.009606f
C5210 commonsourceibias.t14 gnd 0.179464f
C5211 commonsourceibias.n17 gnd 0.012358f
C5212 commonsourceibias.n18 gnd 0.009606f
C5213 commonsourceibias.t64 gnd 0.179464f
C5214 commonsourceibias.n19 gnd 0.071606f
C5215 commonsourceibias.t48 gnd 0.179464f
C5216 commonsourceibias.n20 gnd 0.009057f
C5217 commonsourceibias.n21 gnd 0.009606f
C5218 commonsourceibias.t74 gnd 0.179464f
C5219 commonsourceibias.n22 gnd 0.012175f
C5220 commonsourceibias.n23 gnd 0.009606f
C5221 commonsourceibias.t36 gnd 0.179464f
C5222 commonsourceibias.n24 gnd 0.071606f
C5223 commonsourceibias.t46 gnd 0.179464f
C5224 commonsourceibias.n25 gnd 0.008798f
C5225 commonsourceibias.n26 gnd 0.009606f
C5226 commonsourceibias.t66 gnd 0.179464f
C5227 commonsourceibias.n27 gnd 0.01197f
C5228 commonsourceibias.n28 gnd 0.009606f
C5229 commonsourceibias.t2 gnd 0.179464f
C5230 commonsourceibias.n29 gnd 0.071606f
C5231 commonsourceibias.t20 gnd 0.179464f
C5232 commonsourceibias.n30 gnd 0.008572f
C5233 commonsourceibias.n31 gnd 0.009606f
C5234 commonsourceibias.t38 gnd 0.179464f
C5235 commonsourceibias.n32 gnd 0.011742f
C5236 commonsourceibias.n33 gnd 0.009606f
C5237 commonsourceibias.t0 gnd 0.179464f
C5238 commonsourceibias.n34 gnd 0.071606f
C5239 commonsourceibias.t10 gnd 0.179464f
C5240 commonsourceibias.n35 gnd 0.008375f
C5241 commonsourceibias.n36 gnd 0.009606f
C5242 commonsourceibias.t52 gnd 0.179464f
C5243 commonsourceibias.n37 gnd 0.011489f
C5244 commonsourceibias.n38 gnd 0.009606f
C5245 commonsourceibias.t56 gnd 0.179464f
C5246 commonsourceibias.n39 gnd 0.071606f
C5247 commonsourceibias.t16 gnd 0.179464f
C5248 commonsourceibias.n40 gnd 0.008208f
C5249 commonsourceibias.n41 gnd 0.009606f
C5250 commonsourceibias.t60 gnd 0.179464f
C5251 commonsourceibias.n42 gnd 0.011208f
C5252 commonsourceibias.t76 gnd 0.199531f
C5253 commonsourceibias.t24 gnd 0.179464f
C5254 commonsourceibias.n43 gnd 0.078223f
C5255 commonsourceibias.n44 gnd 0.08584f
C5256 commonsourceibias.n45 gnd 0.039831f
C5257 commonsourceibias.n46 gnd 0.009606f
C5258 commonsourceibias.n47 gnd 0.00935f
C5259 commonsourceibias.n48 gnd 0.013398f
C5260 commonsourceibias.n49 gnd 0.071606f
C5261 commonsourceibias.n50 gnd 0.013389f
C5262 commonsourceibias.n51 gnd 0.009606f
C5263 commonsourceibias.n52 gnd 0.009606f
C5264 commonsourceibias.n53 gnd 0.009606f
C5265 commonsourceibias.n54 gnd 0.012358f
C5266 commonsourceibias.n55 gnd 0.071606f
C5267 commonsourceibias.n56 gnd 0.012648f
C5268 commonsourceibias.n57 gnd 0.012289f
C5269 commonsourceibias.n58 gnd 0.009606f
C5270 commonsourceibias.n59 gnd 0.009606f
C5271 commonsourceibias.n60 gnd 0.009606f
C5272 commonsourceibias.n61 gnd 0.009057f
C5273 commonsourceibias.n62 gnd 0.01341f
C5274 commonsourceibias.n63 gnd 0.071606f
C5275 commonsourceibias.n64 gnd 0.013406f
C5276 commonsourceibias.n65 gnd 0.009606f
C5277 commonsourceibias.n66 gnd 0.009606f
C5278 commonsourceibias.n67 gnd 0.009606f
C5279 commonsourceibias.n68 gnd 0.012175f
C5280 commonsourceibias.n69 gnd 0.071606f
C5281 commonsourceibias.n70 gnd 0.012558f
C5282 commonsourceibias.n71 gnd 0.012378f
C5283 commonsourceibias.n72 gnd 0.009606f
C5284 commonsourceibias.n73 gnd 0.009606f
C5285 commonsourceibias.n74 gnd 0.009606f
C5286 commonsourceibias.n75 gnd 0.008798f
C5287 commonsourceibias.n76 gnd 0.013416f
C5288 commonsourceibias.n77 gnd 0.071606f
C5289 commonsourceibias.n78 gnd 0.013414f
C5290 commonsourceibias.n79 gnd 0.009606f
C5291 commonsourceibias.n80 gnd 0.009606f
C5292 commonsourceibias.n81 gnd 0.009606f
C5293 commonsourceibias.n82 gnd 0.01197f
C5294 commonsourceibias.n83 gnd 0.071606f
C5295 commonsourceibias.n84 gnd 0.012468f
C5296 commonsourceibias.n85 gnd 0.012468f
C5297 commonsourceibias.n86 gnd 0.009606f
C5298 commonsourceibias.n87 gnd 0.009606f
C5299 commonsourceibias.n88 gnd 0.009606f
C5300 commonsourceibias.n89 gnd 0.008572f
C5301 commonsourceibias.n90 gnd 0.013414f
C5302 commonsourceibias.n91 gnd 0.071606f
C5303 commonsourceibias.n92 gnd 0.013416f
C5304 commonsourceibias.n93 gnd 0.009606f
C5305 commonsourceibias.n94 gnd 0.009606f
C5306 commonsourceibias.n95 gnd 0.009606f
C5307 commonsourceibias.n96 gnd 0.011742f
C5308 commonsourceibias.n97 gnd 0.071606f
C5309 commonsourceibias.n98 gnd 0.012378f
C5310 commonsourceibias.n99 gnd 0.012558f
C5311 commonsourceibias.n100 gnd 0.009606f
C5312 commonsourceibias.n101 gnd 0.009606f
C5313 commonsourceibias.n102 gnd 0.009606f
C5314 commonsourceibias.n103 gnd 0.008375f
C5315 commonsourceibias.n104 gnd 0.013406f
C5316 commonsourceibias.n105 gnd 0.071606f
C5317 commonsourceibias.n106 gnd 0.01341f
C5318 commonsourceibias.n107 gnd 0.009606f
C5319 commonsourceibias.n108 gnd 0.009606f
C5320 commonsourceibias.n109 gnd 0.009606f
C5321 commonsourceibias.n110 gnd 0.011489f
C5322 commonsourceibias.n111 gnd 0.071606f
C5323 commonsourceibias.n112 gnd 0.012289f
C5324 commonsourceibias.n113 gnd 0.012648f
C5325 commonsourceibias.n114 gnd 0.009606f
C5326 commonsourceibias.n115 gnd 0.009606f
C5327 commonsourceibias.n116 gnd 0.009606f
C5328 commonsourceibias.n117 gnd 0.008208f
C5329 commonsourceibias.n118 gnd 0.013389f
C5330 commonsourceibias.n119 gnd 0.071606f
C5331 commonsourceibias.n120 gnd 0.013398f
C5332 commonsourceibias.n121 gnd 0.009606f
C5333 commonsourceibias.n122 gnd 0.009606f
C5334 commonsourceibias.n123 gnd 0.009606f
C5335 commonsourceibias.n124 gnd 0.011208f
C5336 commonsourceibias.n125 gnd 0.071606f
C5337 commonsourceibias.n126 gnd 0.011785f
C5338 commonsourceibias.n127 gnd 0.085921f
C5339 commonsourceibias.n128 gnd 0.095704f
C5340 commonsourceibias.t73 gnd 0.020728f
C5341 commonsourceibias.t55 gnd 0.020728f
C5342 commonsourceibias.n129 gnd 0.183161f
C5343 commonsourceibias.n130 gnd 0.158435f
C5344 commonsourceibias.t15 gnd 0.020728f
C5345 commonsourceibias.t65 gnd 0.020728f
C5346 commonsourceibias.n131 gnd 0.183161f
C5347 commonsourceibias.n132 gnd 0.084133f
C5348 commonsourceibias.t49 gnd 0.020728f
C5349 commonsourceibias.t75 gnd 0.020728f
C5350 commonsourceibias.n133 gnd 0.183161f
C5351 commonsourceibias.n134 gnd 0.084133f
C5352 commonsourceibias.t37 gnd 0.020728f
C5353 commonsourceibias.t47 gnd 0.020728f
C5354 commonsourceibias.n135 gnd 0.183161f
C5355 commonsourceibias.n136 gnd 0.084133f
C5356 commonsourceibias.t67 gnd 0.020728f
C5357 commonsourceibias.t3 gnd 0.020728f
C5358 commonsourceibias.n137 gnd 0.183161f
C5359 commonsourceibias.n138 gnd 0.070289f
C5360 commonsourceibias.t25 gnd 0.020728f
C5361 commonsourceibias.t77 gnd 0.020728f
C5362 commonsourceibias.n139 gnd 0.183774f
C5363 commonsourceibias.t17 gnd 0.020728f
C5364 commonsourceibias.t61 gnd 0.020728f
C5365 commonsourceibias.n140 gnd 0.183161f
C5366 commonsourceibias.n141 gnd 0.170671f
C5367 commonsourceibias.t53 gnd 0.020728f
C5368 commonsourceibias.t57 gnd 0.020728f
C5369 commonsourceibias.n142 gnd 0.183161f
C5370 commonsourceibias.n143 gnd 0.084133f
C5371 commonsourceibias.t1 gnd 0.020728f
C5372 commonsourceibias.t11 gnd 0.020728f
C5373 commonsourceibias.n144 gnd 0.183161f
C5374 commonsourceibias.n145 gnd 0.084133f
C5375 commonsourceibias.t21 gnd 0.020728f
C5376 commonsourceibias.t39 gnd 0.020728f
C5377 commonsourceibias.n146 gnd 0.183161f
C5378 commonsourceibias.n147 gnd 0.070289f
C5379 commonsourceibias.n148 gnd 0.085113f
C5380 commonsourceibias.n149 gnd 0.062168f
C5381 commonsourceibias.t136 gnd 0.179464f
C5382 commonsourceibias.n150 gnd 0.071606f
C5383 commonsourceibias.t119 gnd 0.179464f
C5384 commonsourceibias.n151 gnd 0.071606f
C5385 commonsourceibias.n152 gnd 0.009606f
C5386 commonsourceibias.t155 gnd 0.179464f
C5387 commonsourceibias.n153 gnd 0.071606f
C5388 commonsourceibias.n154 gnd 0.009606f
C5389 commonsourceibias.t140 gnd 0.179464f
C5390 commonsourceibias.n155 gnd 0.071606f
C5391 commonsourceibias.n156 gnd 0.009606f
C5392 commonsourceibias.t109 gnd 0.179464f
C5393 commonsourceibias.n157 gnd 0.008375f
C5394 commonsourceibias.n158 gnd 0.009606f
C5395 commonsourceibias.t182 gnd 0.179464f
C5396 commonsourceibias.n159 gnd 0.011489f
C5397 commonsourceibias.n160 gnd 0.009606f
C5398 commonsourceibias.t166 gnd 0.179464f
C5399 commonsourceibias.n161 gnd 0.071606f
C5400 commonsourceibias.t123 gnd 0.179464f
C5401 commonsourceibias.n162 gnd 0.008208f
C5402 commonsourceibias.n163 gnd 0.009606f
C5403 commonsourceibias.t84 gnd 0.179464f
C5404 commonsourceibias.n164 gnd 0.011208f
C5405 commonsourceibias.t100 gnd 0.199531f
C5406 commonsourceibias.t131 gnd 0.179464f
C5407 commonsourceibias.n165 gnd 0.078223f
C5408 commonsourceibias.n166 gnd 0.08584f
C5409 commonsourceibias.n167 gnd 0.039831f
C5410 commonsourceibias.n168 gnd 0.009606f
C5411 commonsourceibias.n169 gnd 0.00935f
C5412 commonsourceibias.n170 gnd 0.013398f
C5413 commonsourceibias.n171 gnd 0.071606f
C5414 commonsourceibias.n172 gnd 0.013389f
C5415 commonsourceibias.n173 gnd 0.009606f
C5416 commonsourceibias.n174 gnd 0.009606f
C5417 commonsourceibias.n175 gnd 0.009606f
C5418 commonsourceibias.n176 gnd 0.012358f
C5419 commonsourceibias.n177 gnd 0.071606f
C5420 commonsourceibias.n178 gnd 0.012648f
C5421 commonsourceibias.n179 gnd 0.012289f
C5422 commonsourceibias.n180 gnd 0.009606f
C5423 commonsourceibias.n181 gnd 0.009606f
C5424 commonsourceibias.n182 gnd 0.009606f
C5425 commonsourceibias.n183 gnd 0.009057f
C5426 commonsourceibias.n184 gnd 0.01341f
C5427 commonsourceibias.n185 gnd 0.071606f
C5428 commonsourceibias.n186 gnd 0.013406f
C5429 commonsourceibias.n187 gnd 0.009606f
C5430 commonsourceibias.n188 gnd 0.009606f
C5431 commonsourceibias.n189 gnd 0.009606f
C5432 commonsourceibias.n190 gnd 0.012175f
C5433 commonsourceibias.n191 gnd 0.071606f
C5434 commonsourceibias.n192 gnd 0.012558f
C5435 commonsourceibias.n193 gnd 0.012378f
C5436 commonsourceibias.n194 gnd 0.009606f
C5437 commonsourceibias.n195 gnd 0.009606f
C5438 commonsourceibias.n196 gnd 0.011742f
C5439 commonsourceibias.n197 gnd 0.008798f
C5440 commonsourceibias.n198 gnd 0.013416f
C5441 commonsourceibias.n199 gnd 0.009606f
C5442 commonsourceibias.n200 gnd 0.009606f
C5443 commonsourceibias.n201 gnd 0.013414f
C5444 commonsourceibias.n202 gnd 0.008572f
C5445 commonsourceibias.n203 gnd 0.01197f
C5446 commonsourceibias.n204 gnd 0.009606f
C5447 commonsourceibias.n205 gnd 0.008392f
C5448 commonsourceibias.n206 gnd 0.012468f
C5449 commonsourceibias.n207 gnd 0.012468f
C5450 commonsourceibias.n208 gnd 0.008392f
C5451 commonsourceibias.n209 gnd 0.009606f
C5452 commonsourceibias.n210 gnd 0.009606f
C5453 commonsourceibias.n211 gnd 0.008572f
C5454 commonsourceibias.n212 gnd 0.013414f
C5455 commonsourceibias.n213 gnd 0.071606f
C5456 commonsourceibias.n214 gnd 0.013416f
C5457 commonsourceibias.n215 gnd 0.009606f
C5458 commonsourceibias.n216 gnd 0.009606f
C5459 commonsourceibias.n217 gnd 0.009606f
C5460 commonsourceibias.n218 gnd 0.011742f
C5461 commonsourceibias.n219 gnd 0.071606f
C5462 commonsourceibias.n220 gnd 0.012378f
C5463 commonsourceibias.n221 gnd 0.012558f
C5464 commonsourceibias.n222 gnd 0.009606f
C5465 commonsourceibias.n223 gnd 0.009606f
C5466 commonsourceibias.n224 gnd 0.009606f
C5467 commonsourceibias.n225 gnd 0.008375f
C5468 commonsourceibias.n226 gnd 0.013406f
C5469 commonsourceibias.n227 gnd 0.071606f
C5470 commonsourceibias.n228 gnd 0.01341f
C5471 commonsourceibias.n229 gnd 0.009606f
C5472 commonsourceibias.n230 gnd 0.009606f
C5473 commonsourceibias.n231 gnd 0.009606f
C5474 commonsourceibias.n232 gnd 0.011489f
C5475 commonsourceibias.n233 gnd 0.071606f
C5476 commonsourceibias.n234 gnd 0.012289f
C5477 commonsourceibias.n235 gnd 0.012648f
C5478 commonsourceibias.n236 gnd 0.009606f
C5479 commonsourceibias.n237 gnd 0.009606f
C5480 commonsourceibias.n238 gnd 0.009606f
C5481 commonsourceibias.n239 gnd 0.008208f
C5482 commonsourceibias.n240 gnd 0.013389f
C5483 commonsourceibias.n241 gnd 0.071606f
C5484 commonsourceibias.n242 gnd 0.013398f
C5485 commonsourceibias.n243 gnd 0.009606f
C5486 commonsourceibias.n244 gnd 0.009606f
C5487 commonsourceibias.n245 gnd 0.009606f
C5488 commonsourceibias.n246 gnd 0.011208f
C5489 commonsourceibias.n247 gnd 0.071606f
C5490 commonsourceibias.n248 gnd 0.011785f
C5491 commonsourceibias.n249 gnd 0.085921f
C5492 commonsourceibias.n250 gnd 0.056157f
C5493 commonsourceibias.n251 gnd 0.012818f
C5494 commonsourceibias.t145 gnd 0.19409f
C5495 commonsourceibias.t172 gnd 0.179464f
C5496 commonsourceibias.n252 gnd 0.00935f
C5497 commonsourceibias.n253 gnd 0.009606f
C5498 commonsourceibias.t160 gnd 0.179464f
C5499 commonsourceibias.n254 gnd 0.012358f
C5500 commonsourceibias.n255 gnd 0.009606f
C5501 commonsourceibias.t146 gnd 0.179464f
C5502 commonsourceibias.n256 gnd 0.071606f
C5503 commonsourceibias.t173 gnd 0.179464f
C5504 commonsourceibias.n257 gnd 0.009057f
C5505 commonsourceibias.n258 gnd 0.009606f
C5506 commonsourceibias.t158 gnd 0.179464f
C5507 commonsourceibias.n259 gnd 0.012175f
C5508 commonsourceibias.n260 gnd 0.009606f
C5509 commonsourceibias.t144 gnd 0.179464f
C5510 commonsourceibias.n261 gnd 0.071606f
C5511 commonsourceibias.t174 gnd 0.179464f
C5512 commonsourceibias.n262 gnd 0.008798f
C5513 commonsourceibias.n263 gnd 0.009606f
C5514 commonsourceibias.t159 gnd 0.179464f
C5515 commonsourceibias.n264 gnd 0.01197f
C5516 commonsourceibias.n265 gnd 0.009606f
C5517 commonsourceibias.t185 gnd 0.179464f
C5518 commonsourceibias.n266 gnd 0.071606f
C5519 commonsourceibias.t175 gnd 0.179464f
C5520 commonsourceibias.n267 gnd 0.008572f
C5521 commonsourceibias.n268 gnd 0.009606f
C5522 commonsourceibias.t157 gnd 0.179464f
C5523 commonsourceibias.n269 gnd 0.011742f
C5524 commonsourceibias.n270 gnd 0.009606f
C5525 commonsourceibias.t190 gnd 0.179464f
C5526 commonsourceibias.n271 gnd 0.071606f
C5527 commonsourceibias.t91 gnd 0.179464f
C5528 commonsourceibias.n272 gnd 0.008375f
C5529 commonsourceibias.n273 gnd 0.009606f
C5530 commonsourceibias.t169 gnd 0.179464f
C5531 commonsourceibias.n274 gnd 0.011489f
C5532 commonsourceibias.n275 gnd 0.009606f
C5533 commonsourceibias.t82 gnd 0.179464f
C5534 commonsourceibias.n276 gnd 0.071606f
C5535 commonsourceibias.t95 gnd 0.179464f
C5536 commonsourceibias.n277 gnd 0.008208f
C5537 commonsourceibias.n278 gnd 0.009606f
C5538 commonsourceibias.t90 gnd 0.179464f
C5539 commonsourceibias.n279 gnd 0.011208f
C5540 commonsourceibias.t94 gnd 0.199531f
C5541 commonsourceibias.t80 gnd 0.179464f
C5542 commonsourceibias.n280 gnd 0.078223f
C5543 commonsourceibias.n281 gnd 0.08584f
C5544 commonsourceibias.n282 gnd 0.039831f
C5545 commonsourceibias.n283 gnd 0.009606f
C5546 commonsourceibias.n284 gnd 0.00935f
C5547 commonsourceibias.n285 gnd 0.013398f
C5548 commonsourceibias.n286 gnd 0.071606f
C5549 commonsourceibias.n287 gnd 0.013389f
C5550 commonsourceibias.n288 gnd 0.009606f
C5551 commonsourceibias.n289 gnd 0.009606f
C5552 commonsourceibias.n290 gnd 0.009606f
C5553 commonsourceibias.n291 gnd 0.012358f
C5554 commonsourceibias.n292 gnd 0.071606f
C5555 commonsourceibias.n293 gnd 0.012648f
C5556 commonsourceibias.n294 gnd 0.012289f
C5557 commonsourceibias.n295 gnd 0.009606f
C5558 commonsourceibias.n296 gnd 0.009606f
C5559 commonsourceibias.n297 gnd 0.009606f
C5560 commonsourceibias.n298 gnd 0.009057f
C5561 commonsourceibias.n299 gnd 0.01341f
C5562 commonsourceibias.n300 gnd 0.071606f
C5563 commonsourceibias.n301 gnd 0.013406f
C5564 commonsourceibias.n302 gnd 0.009606f
C5565 commonsourceibias.n303 gnd 0.009606f
C5566 commonsourceibias.n304 gnd 0.009606f
C5567 commonsourceibias.n305 gnd 0.012175f
C5568 commonsourceibias.n306 gnd 0.071606f
C5569 commonsourceibias.n307 gnd 0.012558f
C5570 commonsourceibias.n308 gnd 0.012378f
C5571 commonsourceibias.n309 gnd 0.009606f
C5572 commonsourceibias.n310 gnd 0.009606f
C5573 commonsourceibias.n311 gnd 0.009606f
C5574 commonsourceibias.n312 gnd 0.008798f
C5575 commonsourceibias.n313 gnd 0.013416f
C5576 commonsourceibias.n314 gnd 0.071606f
C5577 commonsourceibias.n315 gnd 0.013414f
C5578 commonsourceibias.n316 gnd 0.009606f
C5579 commonsourceibias.n317 gnd 0.009606f
C5580 commonsourceibias.n318 gnd 0.009606f
C5581 commonsourceibias.n319 gnd 0.01197f
C5582 commonsourceibias.n320 gnd 0.071606f
C5583 commonsourceibias.n321 gnd 0.012468f
C5584 commonsourceibias.n322 gnd 0.012468f
C5585 commonsourceibias.n323 gnd 0.009606f
C5586 commonsourceibias.n324 gnd 0.009606f
C5587 commonsourceibias.n325 gnd 0.009606f
C5588 commonsourceibias.n326 gnd 0.008572f
C5589 commonsourceibias.n327 gnd 0.013414f
C5590 commonsourceibias.n328 gnd 0.071606f
C5591 commonsourceibias.n329 gnd 0.013416f
C5592 commonsourceibias.n330 gnd 0.009606f
C5593 commonsourceibias.n331 gnd 0.009606f
C5594 commonsourceibias.n332 gnd 0.009606f
C5595 commonsourceibias.n333 gnd 0.011742f
C5596 commonsourceibias.n334 gnd 0.071606f
C5597 commonsourceibias.n335 gnd 0.012378f
C5598 commonsourceibias.n336 gnd 0.012558f
C5599 commonsourceibias.n337 gnd 0.009606f
C5600 commonsourceibias.n338 gnd 0.009606f
C5601 commonsourceibias.n339 gnd 0.009606f
C5602 commonsourceibias.n340 gnd 0.008375f
C5603 commonsourceibias.n341 gnd 0.013406f
C5604 commonsourceibias.n342 gnd 0.071606f
C5605 commonsourceibias.n343 gnd 0.01341f
C5606 commonsourceibias.n344 gnd 0.009606f
C5607 commonsourceibias.n345 gnd 0.009606f
C5608 commonsourceibias.n346 gnd 0.009606f
C5609 commonsourceibias.n347 gnd 0.011489f
C5610 commonsourceibias.n348 gnd 0.071606f
C5611 commonsourceibias.n349 gnd 0.012289f
C5612 commonsourceibias.n350 gnd 0.012648f
C5613 commonsourceibias.n351 gnd 0.009606f
C5614 commonsourceibias.n352 gnd 0.009606f
C5615 commonsourceibias.n353 gnd 0.009606f
C5616 commonsourceibias.n354 gnd 0.008208f
C5617 commonsourceibias.n355 gnd 0.013389f
C5618 commonsourceibias.n356 gnd 0.071606f
C5619 commonsourceibias.n357 gnd 0.013398f
C5620 commonsourceibias.n358 gnd 0.009606f
C5621 commonsourceibias.n359 gnd 0.009606f
C5622 commonsourceibias.n360 gnd 0.009606f
C5623 commonsourceibias.n361 gnd 0.011208f
C5624 commonsourceibias.n362 gnd 0.071606f
C5625 commonsourceibias.n363 gnd 0.011785f
C5626 commonsourceibias.n364 gnd 0.085921f
C5627 commonsourceibias.n365 gnd 0.029883f
C5628 commonsourceibias.n366 gnd 0.153513f
C5629 commonsourceibias.n367 gnd 0.012818f
C5630 commonsourceibias.t89 gnd 0.179464f
C5631 commonsourceibias.n368 gnd 0.00935f
C5632 commonsourceibias.n369 gnd 0.009606f
C5633 commonsourceibias.t107 gnd 0.179464f
C5634 commonsourceibias.n370 gnd 0.012358f
C5635 commonsourceibias.n371 gnd 0.009606f
C5636 commonsourceibias.t168 gnd 0.179464f
C5637 commonsourceibias.n372 gnd 0.071606f
C5638 commonsourceibias.t199 gnd 0.179464f
C5639 commonsourceibias.n373 gnd 0.009057f
C5640 commonsourceibias.n374 gnd 0.009606f
C5641 commonsourceibias.t98 gnd 0.179464f
C5642 commonsourceibias.n375 gnd 0.012175f
C5643 commonsourceibias.n376 gnd 0.009606f
C5644 commonsourceibias.t150 gnd 0.179464f
C5645 commonsourceibias.n377 gnd 0.071606f
C5646 commonsourceibias.t141 gnd 0.179464f
C5647 commonsourceibias.n378 gnd 0.008798f
C5648 commonsourceibias.n379 gnd 0.009606f
C5649 commonsourceibias.t88 gnd 0.179464f
C5650 commonsourceibias.n380 gnd 0.01197f
C5651 commonsourceibias.n381 gnd 0.009606f
C5652 commonsourceibias.t108 gnd 0.179464f
C5653 commonsourceibias.n382 gnd 0.071606f
C5654 commonsourceibias.t130 gnd 0.179464f
C5655 commonsourceibias.n383 gnd 0.008572f
C5656 commonsourceibias.n384 gnd 0.009606f
C5657 commonsourceibias.t198 gnd 0.179464f
C5658 commonsourceibias.n385 gnd 0.011742f
C5659 commonsourceibias.n386 gnd 0.009606f
C5660 commonsourceibias.t186 gnd 0.179464f
C5661 commonsourceibias.n387 gnd 0.071606f
C5662 commonsourceibias.t92 gnd 0.179464f
C5663 commonsourceibias.n388 gnd 0.008375f
C5664 commonsourceibias.n389 gnd 0.009606f
C5665 commonsourceibias.t177 gnd 0.179464f
C5666 commonsourceibias.n390 gnd 0.011489f
C5667 commonsourceibias.n391 gnd 0.009606f
C5668 commonsourceibias.t170 gnd 0.179464f
C5669 commonsourceibias.n392 gnd 0.071606f
C5670 commonsourceibias.t81 gnd 0.179464f
C5671 commonsourceibias.n393 gnd 0.008208f
C5672 commonsourceibias.n394 gnd 0.009606f
C5673 commonsourceibias.t99 gnd 0.179464f
C5674 commonsourceibias.n395 gnd 0.011208f
C5675 commonsourceibias.t184 gnd 0.199531f
C5676 commonsourceibias.t151 gnd 0.179464f
C5677 commonsourceibias.n396 gnd 0.078223f
C5678 commonsourceibias.n397 gnd 0.08584f
C5679 commonsourceibias.n398 gnd 0.039831f
C5680 commonsourceibias.n399 gnd 0.009606f
C5681 commonsourceibias.n400 gnd 0.00935f
C5682 commonsourceibias.n401 gnd 0.013398f
C5683 commonsourceibias.n402 gnd 0.071606f
C5684 commonsourceibias.n403 gnd 0.013389f
C5685 commonsourceibias.n404 gnd 0.009606f
C5686 commonsourceibias.n405 gnd 0.009606f
C5687 commonsourceibias.n406 gnd 0.009606f
C5688 commonsourceibias.n407 gnd 0.012358f
C5689 commonsourceibias.n408 gnd 0.071606f
C5690 commonsourceibias.n409 gnd 0.012648f
C5691 commonsourceibias.n410 gnd 0.012289f
C5692 commonsourceibias.n411 gnd 0.009606f
C5693 commonsourceibias.n412 gnd 0.009606f
C5694 commonsourceibias.n413 gnd 0.009606f
C5695 commonsourceibias.n414 gnd 0.009057f
C5696 commonsourceibias.n415 gnd 0.01341f
C5697 commonsourceibias.n416 gnd 0.071606f
C5698 commonsourceibias.n417 gnd 0.013406f
C5699 commonsourceibias.n418 gnd 0.009606f
C5700 commonsourceibias.n419 gnd 0.009606f
C5701 commonsourceibias.n420 gnd 0.009606f
C5702 commonsourceibias.n421 gnd 0.012175f
C5703 commonsourceibias.n422 gnd 0.071606f
C5704 commonsourceibias.n423 gnd 0.012558f
C5705 commonsourceibias.n424 gnd 0.012378f
C5706 commonsourceibias.n425 gnd 0.009606f
C5707 commonsourceibias.n426 gnd 0.009606f
C5708 commonsourceibias.n427 gnd 0.009606f
C5709 commonsourceibias.n428 gnd 0.008798f
C5710 commonsourceibias.n429 gnd 0.013416f
C5711 commonsourceibias.n430 gnd 0.071606f
C5712 commonsourceibias.n431 gnd 0.013414f
C5713 commonsourceibias.n432 gnd 0.009606f
C5714 commonsourceibias.n433 gnd 0.009606f
C5715 commonsourceibias.n434 gnd 0.009606f
C5716 commonsourceibias.n435 gnd 0.01197f
C5717 commonsourceibias.n436 gnd 0.071606f
C5718 commonsourceibias.n437 gnd 0.012468f
C5719 commonsourceibias.n438 gnd 0.012468f
C5720 commonsourceibias.n439 gnd 0.009606f
C5721 commonsourceibias.n440 gnd 0.009606f
C5722 commonsourceibias.n441 gnd 0.009606f
C5723 commonsourceibias.n442 gnd 0.008572f
C5724 commonsourceibias.n443 gnd 0.013414f
C5725 commonsourceibias.n444 gnd 0.071606f
C5726 commonsourceibias.n445 gnd 0.013416f
C5727 commonsourceibias.n446 gnd 0.009606f
C5728 commonsourceibias.n447 gnd 0.009606f
C5729 commonsourceibias.n448 gnd 0.009606f
C5730 commonsourceibias.n449 gnd 0.011742f
C5731 commonsourceibias.n450 gnd 0.071606f
C5732 commonsourceibias.n451 gnd 0.012378f
C5733 commonsourceibias.n452 gnd 0.012558f
C5734 commonsourceibias.n453 gnd 0.009606f
C5735 commonsourceibias.n454 gnd 0.009606f
C5736 commonsourceibias.n455 gnd 0.009606f
C5737 commonsourceibias.n456 gnd 0.008375f
C5738 commonsourceibias.n457 gnd 0.013406f
C5739 commonsourceibias.n458 gnd 0.071606f
C5740 commonsourceibias.n459 gnd 0.01341f
C5741 commonsourceibias.n460 gnd 0.009606f
C5742 commonsourceibias.n461 gnd 0.009606f
C5743 commonsourceibias.n462 gnd 0.009606f
C5744 commonsourceibias.n463 gnd 0.011489f
C5745 commonsourceibias.n464 gnd 0.071606f
C5746 commonsourceibias.n465 gnd 0.012289f
C5747 commonsourceibias.n466 gnd 0.012648f
C5748 commonsourceibias.n467 gnd 0.009606f
C5749 commonsourceibias.n468 gnd 0.009606f
C5750 commonsourceibias.n469 gnd 0.009606f
C5751 commonsourceibias.n470 gnd 0.008208f
C5752 commonsourceibias.n471 gnd 0.013389f
C5753 commonsourceibias.n472 gnd 0.071606f
C5754 commonsourceibias.n473 gnd 0.013398f
C5755 commonsourceibias.n474 gnd 0.009606f
C5756 commonsourceibias.n475 gnd 0.009606f
C5757 commonsourceibias.n476 gnd 0.009606f
C5758 commonsourceibias.n477 gnd 0.011208f
C5759 commonsourceibias.n478 gnd 0.071606f
C5760 commonsourceibias.n479 gnd 0.011785f
C5761 commonsourceibias.t183 gnd 0.19409f
C5762 commonsourceibias.n480 gnd 0.085921f
C5763 commonsourceibias.n481 gnd 0.029883f
C5764 commonsourceibias.n482 gnd 0.5392f
C5765 commonsourceibias.n483 gnd 0.012818f
C5766 commonsourceibias.t191 gnd 0.19409f
C5767 commonsourceibias.t134 gnd 0.179464f
C5768 commonsourceibias.n484 gnd 0.00935f
C5769 commonsourceibias.n485 gnd 0.009606f
C5770 commonsourceibias.t97 gnd 0.179464f
C5771 commonsourceibias.n486 gnd 0.012358f
C5772 commonsourceibias.n487 gnd 0.009606f
C5773 commonsourceibias.t117 gnd 0.179464f
C5774 commonsourceibias.n488 gnd 0.009057f
C5775 commonsourceibias.n489 gnd 0.009606f
C5776 commonsourceibias.t187 gnd 0.179464f
C5777 commonsourceibias.n490 gnd 0.012175f
C5778 commonsourceibias.n491 gnd 0.009606f
C5779 commonsourceibias.t118 gnd 0.179464f
C5780 commonsourceibias.n492 gnd 0.008798f
C5781 commonsourceibias.n493 gnd 0.009606f
C5782 commonsourceibias.t149 gnd 0.179464f
C5783 commonsourceibias.n494 gnd 0.01197f
C5784 commonsourceibias.t41 gnd 0.020728f
C5785 commonsourceibias.t59 gnd 0.020728f
C5786 commonsourceibias.n495 gnd 0.183774f
C5787 commonsourceibias.t35 gnd 0.020728f
C5788 commonsourceibias.t69 gnd 0.020728f
C5789 commonsourceibias.n496 gnd 0.183161f
C5790 commonsourceibias.n497 gnd 0.170671f
C5791 commonsourceibias.t9 gnd 0.020728f
C5792 commonsourceibias.t7 gnd 0.020728f
C5793 commonsourceibias.n498 gnd 0.183161f
C5794 commonsourceibias.n499 gnd 0.084133f
C5795 commonsourceibias.t63 gnd 0.020728f
C5796 commonsourceibias.t31 gnd 0.020728f
C5797 commonsourceibias.n500 gnd 0.183161f
C5798 commonsourceibias.n501 gnd 0.084133f
C5799 commonsourceibias.t19 gnd 0.020728f
C5800 commonsourceibias.t13 gnd 0.020728f
C5801 commonsourceibias.n502 gnd 0.183161f
C5802 commonsourceibias.n503 gnd 0.070289f
C5803 commonsourceibias.n504 gnd 0.012818f
C5804 commonsourceibias.t4 gnd 0.179464f
C5805 commonsourceibias.n505 gnd 0.00935f
C5806 commonsourceibias.n506 gnd 0.009606f
C5807 commonsourceibias.t78 gnd 0.179464f
C5808 commonsourceibias.n507 gnd 0.012358f
C5809 commonsourceibias.n508 gnd 0.009606f
C5810 commonsourceibias.t28 gnd 0.179464f
C5811 commonsourceibias.n509 gnd 0.009057f
C5812 commonsourceibias.n510 gnd 0.009606f
C5813 commonsourceibias.t50 gnd 0.179464f
C5814 commonsourceibias.n511 gnd 0.012175f
C5815 commonsourceibias.n512 gnd 0.009606f
C5816 commonsourceibias.t26 gnd 0.179464f
C5817 commonsourceibias.n513 gnd 0.008798f
C5818 commonsourceibias.n514 gnd 0.009606f
C5819 commonsourceibias.t44 gnd 0.179464f
C5820 commonsourceibias.n515 gnd 0.01197f
C5821 commonsourceibias.n516 gnd 0.009606f
C5822 commonsourceibias.t12 gnd 0.179464f
C5823 commonsourceibias.n517 gnd 0.008572f
C5824 commonsourceibias.n518 gnd 0.009606f
C5825 commonsourceibias.t18 gnd 0.179464f
C5826 commonsourceibias.n519 gnd 0.011742f
C5827 commonsourceibias.n520 gnd 0.009606f
C5828 commonsourceibias.t62 gnd 0.179464f
C5829 commonsourceibias.n521 gnd 0.008375f
C5830 commonsourceibias.n522 gnd 0.009606f
C5831 commonsourceibias.t6 gnd 0.179464f
C5832 commonsourceibias.n523 gnd 0.011489f
C5833 commonsourceibias.n524 gnd 0.009606f
C5834 commonsourceibias.t68 gnd 0.179464f
C5835 commonsourceibias.n525 gnd 0.008208f
C5836 commonsourceibias.n526 gnd 0.009606f
C5837 commonsourceibias.t34 gnd 0.179464f
C5838 commonsourceibias.n527 gnd 0.011208f
C5839 commonsourceibias.t40 gnd 0.199531f
C5840 commonsourceibias.t58 gnd 0.179464f
C5841 commonsourceibias.n528 gnd 0.078223f
C5842 commonsourceibias.n529 gnd 0.08584f
C5843 commonsourceibias.n530 gnd 0.039831f
C5844 commonsourceibias.n531 gnd 0.009606f
C5845 commonsourceibias.n532 gnd 0.00935f
C5846 commonsourceibias.n533 gnd 0.013398f
C5847 commonsourceibias.n534 gnd 0.071606f
C5848 commonsourceibias.n535 gnd 0.013389f
C5849 commonsourceibias.n536 gnd 0.009606f
C5850 commonsourceibias.n537 gnd 0.009606f
C5851 commonsourceibias.n538 gnd 0.009606f
C5852 commonsourceibias.n539 gnd 0.012358f
C5853 commonsourceibias.n540 gnd 0.071606f
C5854 commonsourceibias.n541 gnd 0.012648f
C5855 commonsourceibias.t8 gnd 0.179464f
C5856 commonsourceibias.n542 gnd 0.071606f
C5857 commonsourceibias.n543 gnd 0.012289f
C5858 commonsourceibias.n544 gnd 0.009606f
C5859 commonsourceibias.n545 gnd 0.009606f
C5860 commonsourceibias.n546 gnd 0.009606f
C5861 commonsourceibias.n547 gnd 0.009057f
C5862 commonsourceibias.n548 gnd 0.01341f
C5863 commonsourceibias.n549 gnd 0.071606f
C5864 commonsourceibias.n550 gnd 0.013406f
C5865 commonsourceibias.n551 gnd 0.009606f
C5866 commonsourceibias.n552 gnd 0.009606f
C5867 commonsourceibias.n553 gnd 0.009606f
C5868 commonsourceibias.n554 gnd 0.012175f
C5869 commonsourceibias.n555 gnd 0.071606f
C5870 commonsourceibias.n556 gnd 0.012558f
C5871 commonsourceibias.t30 gnd 0.179464f
C5872 commonsourceibias.n557 gnd 0.071606f
C5873 commonsourceibias.n558 gnd 0.012378f
C5874 commonsourceibias.n559 gnd 0.009606f
C5875 commonsourceibias.n560 gnd 0.009606f
C5876 commonsourceibias.n561 gnd 0.009606f
C5877 commonsourceibias.n562 gnd 0.008798f
C5878 commonsourceibias.n563 gnd 0.013416f
C5879 commonsourceibias.n564 gnd 0.071606f
C5880 commonsourceibias.n565 gnd 0.013414f
C5881 commonsourceibias.n566 gnd 0.009606f
C5882 commonsourceibias.n567 gnd 0.009606f
C5883 commonsourceibias.n568 gnd 0.009606f
C5884 commonsourceibias.n569 gnd 0.01197f
C5885 commonsourceibias.n570 gnd 0.071606f
C5886 commonsourceibias.n571 gnd 0.012468f
C5887 commonsourceibias.t32 gnd 0.179464f
C5888 commonsourceibias.n572 gnd 0.071606f
C5889 commonsourceibias.n573 gnd 0.012468f
C5890 commonsourceibias.n574 gnd 0.009606f
C5891 commonsourceibias.n575 gnd 0.009606f
C5892 commonsourceibias.n576 gnd 0.009606f
C5893 commonsourceibias.n577 gnd 0.008572f
C5894 commonsourceibias.n578 gnd 0.013414f
C5895 commonsourceibias.n579 gnd 0.071606f
C5896 commonsourceibias.n580 gnd 0.013416f
C5897 commonsourceibias.n581 gnd 0.009606f
C5898 commonsourceibias.n582 gnd 0.009606f
C5899 commonsourceibias.n583 gnd 0.009606f
C5900 commonsourceibias.n584 gnd 0.011742f
C5901 commonsourceibias.n585 gnd 0.071606f
C5902 commonsourceibias.n586 gnd 0.012378f
C5903 commonsourceibias.t22 gnd 0.179464f
C5904 commonsourceibias.n587 gnd 0.071606f
C5905 commonsourceibias.n588 gnd 0.012558f
C5906 commonsourceibias.n589 gnd 0.009606f
C5907 commonsourceibias.n590 gnd 0.009606f
C5908 commonsourceibias.n591 gnd 0.009606f
C5909 commonsourceibias.n592 gnd 0.008375f
C5910 commonsourceibias.n593 gnd 0.013406f
C5911 commonsourceibias.n594 gnd 0.071606f
C5912 commonsourceibias.n595 gnd 0.01341f
C5913 commonsourceibias.n596 gnd 0.009606f
C5914 commonsourceibias.n597 gnd 0.009606f
C5915 commonsourceibias.n598 gnd 0.009606f
C5916 commonsourceibias.n599 gnd 0.011489f
C5917 commonsourceibias.n600 gnd 0.071606f
C5918 commonsourceibias.n601 gnd 0.012289f
C5919 commonsourceibias.t42 gnd 0.179464f
C5920 commonsourceibias.n602 gnd 0.071606f
C5921 commonsourceibias.n603 gnd 0.012648f
C5922 commonsourceibias.n604 gnd 0.009606f
C5923 commonsourceibias.n605 gnd 0.009606f
C5924 commonsourceibias.n606 gnd 0.009606f
C5925 commonsourceibias.n607 gnd 0.008208f
C5926 commonsourceibias.n608 gnd 0.013389f
C5927 commonsourceibias.n609 gnd 0.071606f
C5928 commonsourceibias.n610 gnd 0.013398f
C5929 commonsourceibias.n611 gnd 0.009606f
C5930 commonsourceibias.n612 gnd 0.009606f
C5931 commonsourceibias.n613 gnd 0.009606f
C5932 commonsourceibias.n614 gnd 0.011208f
C5933 commonsourceibias.n615 gnd 0.071606f
C5934 commonsourceibias.n616 gnd 0.011785f
C5935 commonsourceibias.t70 gnd 0.19409f
C5936 commonsourceibias.n617 gnd 0.085921f
C5937 commonsourceibias.n618 gnd 0.095704f
C5938 commonsourceibias.t5 gnd 0.020728f
C5939 commonsourceibias.t71 gnd 0.020728f
C5940 commonsourceibias.n619 gnd 0.183161f
C5941 commonsourceibias.n620 gnd 0.158435f
C5942 commonsourceibias.t43 gnd 0.020728f
C5943 commonsourceibias.t79 gnd 0.020728f
C5944 commonsourceibias.n621 gnd 0.183161f
C5945 commonsourceibias.n622 gnd 0.084133f
C5946 commonsourceibias.t51 gnd 0.020728f
C5947 commonsourceibias.t29 gnd 0.020728f
C5948 commonsourceibias.n623 gnd 0.183161f
C5949 commonsourceibias.n624 gnd 0.084133f
C5950 commonsourceibias.t27 gnd 0.020728f
C5951 commonsourceibias.t23 gnd 0.020728f
C5952 commonsourceibias.n625 gnd 0.183161f
C5953 commonsourceibias.n626 gnd 0.084133f
C5954 commonsourceibias.t33 gnd 0.020728f
C5955 commonsourceibias.t45 gnd 0.020728f
C5956 commonsourceibias.n627 gnd 0.183161f
C5957 commonsourceibias.n628 gnd 0.070289f
C5958 commonsourceibias.n629 gnd 0.085113f
C5959 commonsourceibias.n630 gnd 0.062168f
C5960 commonsourceibias.t105 gnd 0.179464f
C5961 commonsourceibias.n631 gnd 0.071606f
C5962 commonsourceibias.n632 gnd 0.009606f
C5963 commonsourceibias.t122 gnd 0.179464f
C5964 commonsourceibias.n633 gnd 0.071606f
C5965 commonsourceibias.n634 gnd 0.009606f
C5966 commonsourceibias.t115 gnd 0.179464f
C5967 commonsourceibias.n635 gnd 0.071606f
C5968 commonsourceibias.n636 gnd 0.009606f
C5969 commonsourceibias.t83 gnd 0.179464f
C5970 commonsourceibias.n637 gnd 0.008375f
C5971 commonsourceibias.n638 gnd 0.009606f
C5972 commonsourceibias.t111 gnd 0.179464f
C5973 commonsourceibias.n639 gnd 0.011489f
C5974 commonsourceibias.n640 gnd 0.009606f
C5975 commonsourceibias.t192 gnd 0.179464f
C5976 commonsourceibias.n641 gnd 0.008208f
C5977 commonsourceibias.n642 gnd 0.009606f
C5978 commonsourceibias.t127 gnd 0.179464f
C5979 commonsourceibias.n643 gnd 0.011208f
C5980 commonsourceibias.t153 gnd 0.199531f
C5981 commonsourceibias.t86 gnd 0.179464f
C5982 commonsourceibias.n644 gnd 0.078223f
C5983 commonsourceibias.n645 gnd 0.08584f
C5984 commonsourceibias.n646 gnd 0.039831f
C5985 commonsourceibias.n647 gnd 0.009606f
C5986 commonsourceibias.n648 gnd 0.00935f
C5987 commonsourceibias.n649 gnd 0.013398f
C5988 commonsourceibias.n650 gnd 0.071606f
C5989 commonsourceibias.n651 gnd 0.013389f
C5990 commonsourceibias.n652 gnd 0.009606f
C5991 commonsourceibias.n653 gnd 0.009606f
C5992 commonsourceibias.n654 gnd 0.009606f
C5993 commonsourceibias.n655 gnd 0.012358f
C5994 commonsourceibias.n656 gnd 0.071606f
C5995 commonsourceibias.n657 gnd 0.012648f
C5996 commonsourceibias.t110 gnd 0.179464f
C5997 commonsourceibias.n658 gnd 0.071606f
C5998 commonsourceibias.n659 gnd 0.012289f
C5999 commonsourceibias.n660 gnd 0.009606f
C6000 commonsourceibias.n661 gnd 0.009606f
C6001 commonsourceibias.n662 gnd 0.009606f
C6002 commonsourceibias.n663 gnd 0.009057f
C6003 commonsourceibias.n664 gnd 0.01341f
C6004 commonsourceibias.n665 gnd 0.071606f
C6005 commonsourceibias.n666 gnd 0.013406f
C6006 commonsourceibias.n667 gnd 0.009606f
C6007 commonsourceibias.n668 gnd 0.009606f
C6008 commonsourceibias.n669 gnd 0.009606f
C6009 commonsourceibias.n670 gnd 0.012175f
C6010 commonsourceibias.n671 gnd 0.071606f
C6011 commonsourceibias.n672 gnd 0.012558f
C6012 commonsourceibias.n673 gnd 0.012378f
C6013 commonsourceibias.n674 gnd 0.009606f
C6014 commonsourceibias.n675 gnd 0.009606f
C6015 commonsourceibias.n676 gnd 0.011742f
C6016 commonsourceibias.n677 gnd 0.008798f
C6017 commonsourceibias.n678 gnd 0.013416f
C6018 commonsourceibias.n679 gnd 0.009606f
C6019 commonsourceibias.n680 gnd 0.009606f
C6020 commonsourceibias.n681 gnd 0.013414f
C6021 commonsourceibias.n682 gnd 0.008572f
C6022 commonsourceibias.n683 gnd 0.01197f
C6023 commonsourceibias.n684 gnd 0.009606f
C6024 commonsourceibias.n685 gnd 0.008392f
C6025 commonsourceibias.n686 gnd 0.012468f
C6026 commonsourceibias.t114 gnd 0.179464f
C6027 commonsourceibias.n687 gnd 0.071606f
C6028 commonsourceibias.n688 gnd 0.012468f
C6029 commonsourceibias.n689 gnd 0.008392f
C6030 commonsourceibias.n690 gnd 0.009606f
C6031 commonsourceibias.n691 gnd 0.009606f
C6032 commonsourceibias.n692 gnd 0.008572f
C6033 commonsourceibias.n693 gnd 0.013414f
C6034 commonsourceibias.n694 gnd 0.071606f
C6035 commonsourceibias.n695 gnd 0.013416f
C6036 commonsourceibias.n696 gnd 0.009606f
C6037 commonsourceibias.n697 gnd 0.009606f
C6038 commonsourceibias.n698 gnd 0.009606f
C6039 commonsourceibias.n699 gnd 0.011742f
C6040 commonsourceibias.n700 gnd 0.071606f
C6041 commonsourceibias.n701 gnd 0.012378f
C6042 commonsourceibias.t132 gnd 0.179464f
C6043 commonsourceibias.n702 gnd 0.071606f
C6044 commonsourceibias.n703 gnd 0.012558f
C6045 commonsourceibias.n704 gnd 0.009606f
C6046 commonsourceibias.n705 gnd 0.009606f
C6047 commonsourceibias.n706 gnd 0.009606f
C6048 commonsourceibias.n707 gnd 0.008375f
C6049 commonsourceibias.n708 gnd 0.013406f
C6050 commonsourceibias.n709 gnd 0.071606f
C6051 commonsourceibias.n710 gnd 0.01341f
C6052 commonsourceibias.n711 gnd 0.009606f
C6053 commonsourceibias.n712 gnd 0.009606f
C6054 commonsourceibias.n713 gnd 0.009606f
C6055 commonsourceibias.n714 gnd 0.011489f
C6056 commonsourceibias.n715 gnd 0.071606f
C6057 commonsourceibias.n716 gnd 0.012289f
C6058 commonsourceibias.t152 gnd 0.179464f
C6059 commonsourceibias.n717 gnd 0.071606f
C6060 commonsourceibias.n718 gnd 0.012648f
C6061 commonsourceibias.n719 gnd 0.009606f
C6062 commonsourceibias.n720 gnd 0.009606f
C6063 commonsourceibias.n721 gnd 0.009606f
C6064 commonsourceibias.n722 gnd 0.008208f
C6065 commonsourceibias.n723 gnd 0.013389f
C6066 commonsourceibias.n724 gnd 0.071606f
C6067 commonsourceibias.n725 gnd 0.013398f
C6068 commonsourceibias.n726 gnd 0.009606f
C6069 commonsourceibias.n727 gnd 0.009606f
C6070 commonsourceibias.n728 gnd 0.009606f
C6071 commonsourceibias.n729 gnd 0.011208f
C6072 commonsourceibias.n730 gnd 0.071606f
C6073 commonsourceibias.n731 gnd 0.011785f
C6074 commonsourceibias.n732 gnd 0.085921f
C6075 commonsourceibias.n733 gnd 0.056157f
C6076 commonsourceibias.n734 gnd 0.012818f
C6077 commonsourceibias.t148 gnd 0.179464f
C6078 commonsourceibias.n735 gnd 0.00935f
C6079 commonsourceibias.n736 gnd 0.009606f
C6080 commonsourceibias.t139 gnd 0.179464f
C6081 commonsourceibias.n737 gnd 0.012358f
C6082 commonsourceibias.n738 gnd 0.009606f
C6083 commonsourceibias.t147 gnd 0.179464f
C6084 commonsourceibias.n739 gnd 0.009057f
C6085 commonsourceibias.n740 gnd 0.009606f
C6086 commonsourceibias.t138 gnd 0.179464f
C6087 commonsourceibias.n741 gnd 0.012175f
C6088 commonsourceibias.n742 gnd 0.009606f
C6089 commonsourceibias.t154 gnd 0.179464f
C6090 commonsourceibias.n743 gnd 0.008798f
C6091 commonsourceibias.n744 gnd 0.009606f
C6092 commonsourceibias.t137 gnd 0.179464f
C6093 commonsourceibias.n745 gnd 0.01197f
C6094 commonsourceibias.n746 gnd 0.009606f
C6095 commonsourceibias.t195 gnd 0.179464f
C6096 commonsourceibias.n747 gnd 0.008572f
C6097 commonsourceibias.n748 gnd 0.009606f
C6098 commonsourceibias.t135 gnd 0.179464f
C6099 commonsourceibias.n749 gnd 0.011742f
C6100 commonsourceibias.n750 gnd 0.009606f
C6101 commonsourceibias.t194 gnd 0.179464f
C6102 commonsourceibias.n751 gnd 0.008375f
C6103 commonsourceibias.n752 gnd 0.009606f
C6104 commonsourceibias.t176 gnd 0.179464f
C6105 commonsourceibias.n753 gnd 0.011489f
C6106 commonsourceibias.n754 gnd 0.009606f
C6107 commonsourceibias.t189 gnd 0.179464f
C6108 commonsourceibias.n755 gnd 0.008208f
C6109 commonsourceibias.n756 gnd 0.009606f
C6110 commonsourceibias.t180 gnd 0.179464f
C6111 commonsourceibias.n757 gnd 0.011208f
C6112 commonsourceibias.t188 gnd 0.199531f
C6113 commonsourceibias.t163 gnd 0.179464f
C6114 commonsourceibias.n758 gnd 0.078223f
C6115 commonsourceibias.n759 gnd 0.08584f
C6116 commonsourceibias.n760 gnd 0.039831f
C6117 commonsourceibias.n761 gnd 0.009606f
C6118 commonsourceibias.n762 gnd 0.00935f
C6119 commonsourceibias.n763 gnd 0.013398f
C6120 commonsourceibias.n764 gnd 0.071606f
C6121 commonsourceibias.n765 gnd 0.013389f
C6122 commonsourceibias.n766 gnd 0.009606f
C6123 commonsourceibias.n767 gnd 0.009606f
C6124 commonsourceibias.n768 gnd 0.009606f
C6125 commonsourceibias.n769 gnd 0.012358f
C6126 commonsourceibias.n770 gnd 0.071606f
C6127 commonsourceibias.n771 gnd 0.012648f
C6128 commonsourceibias.t164 gnd 0.179464f
C6129 commonsourceibias.n772 gnd 0.071606f
C6130 commonsourceibias.n773 gnd 0.012289f
C6131 commonsourceibias.n774 gnd 0.009606f
C6132 commonsourceibias.n775 gnd 0.009606f
C6133 commonsourceibias.n776 gnd 0.009606f
C6134 commonsourceibias.n777 gnd 0.009057f
C6135 commonsourceibias.n778 gnd 0.01341f
C6136 commonsourceibias.n779 gnd 0.071606f
C6137 commonsourceibias.n780 gnd 0.013406f
C6138 commonsourceibias.n781 gnd 0.009606f
C6139 commonsourceibias.n782 gnd 0.009606f
C6140 commonsourceibias.n783 gnd 0.009606f
C6141 commonsourceibias.n784 gnd 0.012175f
C6142 commonsourceibias.n785 gnd 0.071606f
C6143 commonsourceibias.n786 gnd 0.012558f
C6144 commonsourceibias.t171 gnd 0.179464f
C6145 commonsourceibias.n787 gnd 0.071606f
C6146 commonsourceibias.n788 gnd 0.012378f
C6147 commonsourceibias.n789 gnd 0.009606f
C6148 commonsourceibias.n790 gnd 0.009606f
C6149 commonsourceibias.n791 gnd 0.009606f
C6150 commonsourceibias.n792 gnd 0.008798f
C6151 commonsourceibias.n793 gnd 0.013416f
C6152 commonsourceibias.n794 gnd 0.071606f
C6153 commonsourceibias.n795 gnd 0.013414f
C6154 commonsourceibias.n796 gnd 0.009606f
C6155 commonsourceibias.n797 gnd 0.009606f
C6156 commonsourceibias.n798 gnd 0.009606f
C6157 commonsourceibias.n799 gnd 0.01197f
C6158 commonsourceibias.n800 gnd 0.071606f
C6159 commonsourceibias.n801 gnd 0.012468f
C6160 commonsourceibias.t161 gnd 0.179464f
C6161 commonsourceibias.n802 gnd 0.071606f
C6162 commonsourceibias.n803 gnd 0.012468f
C6163 commonsourceibias.n804 gnd 0.009606f
C6164 commonsourceibias.n805 gnd 0.009606f
C6165 commonsourceibias.n806 gnd 0.009606f
C6166 commonsourceibias.n807 gnd 0.008572f
C6167 commonsourceibias.n808 gnd 0.013414f
C6168 commonsourceibias.n809 gnd 0.071606f
C6169 commonsourceibias.n810 gnd 0.013416f
C6170 commonsourceibias.n811 gnd 0.009606f
C6171 commonsourceibias.n812 gnd 0.009606f
C6172 commonsourceibias.n813 gnd 0.009606f
C6173 commonsourceibias.n814 gnd 0.011742f
C6174 commonsourceibias.n815 gnd 0.071606f
C6175 commonsourceibias.n816 gnd 0.012378f
C6176 commonsourceibias.t162 gnd 0.179464f
C6177 commonsourceibias.n817 gnd 0.071606f
C6178 commonsourceibias.n818 gnd 0.012558f
C6179 commonsourceibias.n819 gnd 0.009606f
C6180 commonsourceibias.n820 gnd 0.009606f
C6181 commonsourceibias.n821 gnd 0.009606f
C6182 commonsourceibias.n822 gnd 0.008375f
C6183 commonsourceibias.n823 gnd 0.013406f
C6184 commonsourceibias.n824 gnd 0.071606f
C6185 commonsourceibias.n825 gnd 0.01341f
C6186 commonsourceibias.n826 gnd 0.009606f
C6187 commonsourceibias.n827 gnd 0.009606f
C6188 commonsourceibias.n828 gnd 0.009606f
C6189 commonsourceibias.n829 gnd 0.011489f
C6190 commonsourceibias.n830 gnd 0.071606f
C6191 commonsourceibias.n831 gnd 0.012289f
C6192 commonsourceibias.t128 gnd 0.179464f
C6193 commonsourceibias.n832 gnd 0.071606f
C6194 commonsourceibias.n833 gnd 0.012648f
C6195 commonsourceibias.n834 gnd 0.009606f
C6196 commonsourceibias.n835 gnd 0.009606f
C6197 commonsourceibias.n836 gnd 0.009606f
C6198 commonsourceibias.n837 gnd 0.008208f
C6199 commonsourceibias.n838 gnd 0.013389f
C6200 commonsourceibias.n839 gnd 0.071606f
C6201 commonsourceibias.n840 gnd 0.013398f
C6202 commonsourceibias.n841 gnd 0.009606f
C6203 commonsourceibias.n842 gnd 0.009606f
C6204 commonsourceibias.n843 gnd 0.009606f
C6205 commonsourceibias.n844 gnd 0.011208f
C6206 commonsourceibias.n845 gnd 0.071606f
C6207 commonsourceibias.n846 gnd 0.011785f
C6208 commonsourceibias.t129 gnd 0.19409f
C6209 commonsourceibias.n847 gnd 0.085921f
C6210 commonsourceibias.n848 gnd 0.029883f
C6211 commonsourceibias.n849 gnd 0.153513f
C6212 commonsourceibias.n850 gnd 0.012818f
C6213 commonsourceibias.t113 gnd 0.179464f
C6214 commonsourceibias.n851 gnd 0.00935f
C6215 commonsourceibias.n852 gnd 0.009606f
C6216 commonsourceibias.t125 gnd 0.179464f
C6217 commonsourceibias.n853 gnd 0.012358f
C6218 commonsourceibias.n854 gnd 0.009606f
C6219 commonsourceibias.t103 gnd 0.179464f
C6220 commonsourceibias.n855 gnd 0.009057f
C6221 commonsourceibias.n856 gnd 0.009606f
C6222 commonsourceibias.t120 gnd 0.179464f
C6223 commonsourceibias.n857 gnd 0.012175f
C6224 commonsourceibias.n858 gnd 0.009606f
C6225 commonsourceibias.t179 gnd 0.179464f
C6226 commonsourceibias.n859 gnd 0.008798f
C6227 commonsourceibias.n860 gnd 0.009606f
C6228 commonsourceibias.t112 gnd 0.179464f
C6229 commonsourceibias.n861 gnd 0.01197f
C6230 commonsourceibias.n862 gnd 0.009606f
C6231 commonsourceibias.t121 gnd 0.179464f
C6232 commonsourceibias.n863 gnd 0.008572f
C6233 commonsourceibias.n864 gnd 0.009606f
C6234 commonsourceibias.t102 gnd 0.179464f
C6235 commonsourceibias.n865 gnd 0.011742f
C6236 commonsourceibias.n866 gnd 0.009606f
C6237 commonsourceibias.t116 gnd 0.179464f
C6238 commonsourceibias.n867 gnd 0.008375f
C6239 commonsourceibias.n868 gnd 0.009606f
C6240 commonsourceibias.t167 gnd 0.179464f
C6241 commonsourceibias.n869 gnd 0.011489f
C6242 commonsourceibias.n870 gnd 0.009606f
C6243 commonsourceibias.t87 gnd 0.179464f
C6244 commonsourceibias.n871 gnd 0.008208f
C6245 commonsourceibias.n872 gnd 0.009606f
C6246 commonsourceibias.t106 gnd 0.179464f
C6247 commonsourceibias.n873 gnd 0.011208f
C6248 commonsourceibias.t196 gnd 0.199531f
C6249 commonsourceibias.t165 gnd 0.179464f
C6250 commonsourceibias.n874 gnd 0.078223f
C6251 commonsourceibias.n875 gnd 0.08584f
C6252 commonsourceibias.n876 gnd 0.039831f
C6253 commonsourceibias.n877 gnd 0.009606f
C6254 commonsourceibias.n878 gnd 0.00935f
C6255 commonsourceibias.n879 gnd 0.013398f
C6256 commonsourceibias.n880 gnd 0.071606f
C6257 commonsourceibias.n881 gnd 0.013389f
C6258 commonsourceibias.n882 gnd 0.009606f
C6259 commonsourceibias.n883 gnd 0.009606f
C6260 commonsourceibias.n884 gnd 0.009606f
C6261 commonsourceibias.n885 gnd 0.012358f
C6262 commonsourceibias.n886 gnd 0.071606f
C6263 commonsourceibias.n887 gnd 0.012648f
C6264 commonsourceibias.t178 gnd 0.179464f
C6265 commonsourceibias.n888 gnd 0.071606f
C6266 commonsourceibias.n889 gnd 0.012289f
C6267 commonsourceibias.n890 gnd 0.009606f
C6268 commonsourceibias.n891 gnd 0.009606f
C6269 commonsourceibias.n892 gnd 0.009606f
C6270 commonsourceibias.n893 gnd 0.009057f
C6271 commonsourceibias.n894 gnd 0.01341f
C6272 commonsourceibias.n895 gnd 0.071606f
C6273 commonsourceibias.n896 gnd 0.013406f
C6274 commonsourceibias.n897 gnd 0.009606f
C6275 commonsourceibias.n898 gnd 0.009606f
C6276 commonsourceibias.n899 gnd 0.009606f
C6277 commonsourceibias.n900 gnd 0.012175f
C6278 commonsourceibias.n901 gnd 0.071606f
C6279 commonsourceibias.n902 gnd 0.012558f
C6280 commonsourceibias.t96 gnd 0.179464f
C6281 commonsourceibias.n903 gnd 0.071606f
C6282 commonsourceibias.n904 gnd 0.012378f
C6283 commonsourceibias.n905 gnd 0.009606f
C6284 commonsourceibias.n906 gnd 0.009606f
C6285 commonsourceibias.n907 gnd 0.009606f
C6286 commonsourceibias.n908 gnd 0.008798f
C6287 commonsourceibias.n909 gnd 0.013416f
C6288 commonsourceibias.n910 gnd 0.071606f
C6289 commonsourceibias.n911 gnd 0.013414f
C6290 commonsourceibias.n912 gnd 0.009606f
C6291 commonsourceibias.n913 gnd 0.009606f
C6292 commonsourceibias.n914 gnd 0.009606f
C6293 commonsourceibias.n915 gnd 0.01197f
C6294 commonsourceibias.n916 gnd 0.071606f
C6295 commonsourceibias.n917 gnd 0.012468f
C6296 commonsourceibias.t126 gnd 0.179464f
C6297 commonsourceibias.n918 gnd 0.071606f
C6298 commonsourceibias.n919 gnd 0.012468f
C6299 commonsourceibias.n920 gnd 0.009606f
C6300 commonsourceibias.n921 gnd 0.009606f
C6301 commonsourceibias.n922 gnd 0.009606f
C6302 commonsourceibias.n923 gnd 0.008572f
C6303 commonsourceibias.n924 gnd 0.013414f
C6304 commonsourceibias.n925 gnd 0.071606f
C6305 commonsourceibias.n926 gnd 0.013416f
C6306 commonsourceibias.n927 gnd 0.009606f
C6307 commonsourceibias.n928 gnd 0.009606f
C6308 commonsourceibias.n929 gnd 0.009606f
C6309 commonsourceibias.n930 gnd 0.011742f
C6310 commonsourceibias.n931 gnd 0.071606f
C6311 commonsourceibias.n932 gnd 0.012378f
C6312 commonsourceibias.t133 gnd 0.179464f
C6313 commonsourceibias.n933 gnd 0.071606f
C6314 commonsourceibias.n934 gnd 0.012558f
C6315 commonsourceibias.n935 gnd 0.009606f
C6316 commonsourceibias.n936 gnd 0.009606f
C6317 commonsourceibias.n937 gnd 0.009606f
C6318 commonsourceibias.n938 gnd 0.008375f
C6319 commonsourceibias.n939 gnd 0.013406f
C6320 commonsourceibias.n940 gnd 0.071606f
C6321 commonsourceibias.n941 gnd 0.01341f
C6322 commonsourceibias.n942 gnd 0.009606f
C6323 commonsourceibias.n943 gnd 0.009606f
C6324 commonsourceibias.n944 gnd 0.009606f
C6325 commonsourceibias.n945 gnd 0.011489f
C6326 commonsourceibias.n946 gnd 0.071606f
C6327 commonsourceibias.n947 gnd 0.012289f
C6328 commonsourceibias.t85 gnd 0.179464f
C6329 commonsourceibias.n948 gnd 0.071606f
C6330 commonsourceibias.n949 gnd 0.012648f
C6331 commonsourceibias.n950 gnd 0.009606f
C6332 commonsourceibias.n951 gnd 0.009606f
C6333 commonsourceibias.n952 gnd 0.009606f
C6334 commonsourceibias.n953 gnd 0.008208f
C6335 commonsourceibias.n954 gnd 0.013389f
C6336 commonsourceibias.n955 gnd 0.071606f
C6337 commonsourceibias.n956 gnd 0.013398f
C6338 commonsourceibias.n957 gnd 0.009606f
C6339 commonsourceibias.n958 gnd 0.009606f
C6340 commonsourceibias.n959 gnd 0.009606f
C6341 commonsourceibias.n960 gnd 0.011208f
C6342 commonsourceibias.n961 gnd 0.071606f
C6343 commonsourceibias.n962 gnd 0.011785f
C6344 commonsourceibias.t93 gnd 0.19409f
C6345 commonsourceibias.n963 gnd 0.085921f
C6346 commonsourceibias.n964 gnd 0.029883f
C6347 commonsourceibias.n965 gnd 0.202576f
C6348 commonsourceibias.n966 gnd 5.69738f
.ends

