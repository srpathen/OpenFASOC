* NGSPICE file created from opamp474.ext - technology: sky130A

.subckt opamp474 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 a_n8964_8799.t37 plus.t5 a_n2903_n3924.t35 gnd.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X1 a_n2804_13878.t25 a_n2982_13878.t44 a_n2982_13878.t45 vdd.t44 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X2 CSoutput.t215 commonsourceibias.t80 gnd.t160 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X3 a_n2804_13878.t30 a_n2982_13878.t64 vdd.t57 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 vdd.t191 a_n8964_8799.t40 CSoutput.t95 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X5 gnd.t92 commonsourceibias.t81 CSoutput.t214 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X6 CSoutput.t213 commonsourceibias.t82 gnd.t104 gnd.t103 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 CSoutput.t212 commonsourceibias.t83 gnd.t119 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 CSoutput.t94 a_n8964_8799.t41 vdd.t190 vdd.t82 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X9 a_n2903_n3924.t31 plus.t6 a_n8964_8799.t36 gnd.t345 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X10 gnd.t43 commonsourceibias.t84 CSoutput.t211 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X11 CSoutput.t216 a_n2982_8322.t37 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X12 plus.t3 gnd.t284 gnd.t286 gnd.t285 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X13 vdd.t189 a_n8964_8799.t42 CSoutput.t93 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X14 a_n2982_8322.t23 a_n2982_13878.t65 a_n8964_8799.t0 vdd.t54 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X15 CSoutput.t92 a_n8964_8799.t43 vdd.t188 vdd.t101 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X16 vdd.t187 a_n8964_8799.t44 CSoutput.t91 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X17 vdd.t60 CSoutput.t217 output.t18 gnd.t118 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X18 CSoutput.t90 a_n8964_8799.t45 vdd.t186 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X19 CSoutput.t210 commonsourceibias.t85 gnd.t61 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X20 gnd.t124 commonsourceibias.t86 CSoutput.t209 gnd.t123 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X21 CSoutput.t208 commonsourceibias.t87 gnd.t294 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X22 gnd.t394 commonsourceibias.t88 CSoutput.t207 gnd.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X23 vdd.t184 a_n8964_8799.t46 CSoutput.t89 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X24 vdd.t185 a_n8964_8799.t47 CSoutput.t88 vdd.t129 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X25 CSoutput.t206 commonsourceibias.t89 gnd.t370 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X26 CSoutput.t205 commonsourceibias.t90 gnd.t346 gnd.t108 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X27 gnd.t399 commonsourceibias.t91 CSoutput.t204 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X28 gnd.t283 gnd.t280 gnd.t282 gnd.t281 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X29 gnd.t279 gnd.t277 gnd.t278 gnd.t183 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X30 commonsourceibias.t79 commonsourceibias.t78 gnd.t379 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X31 CSoutput.t203 commonsourceibias.t92 gnd.t31 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 gnd.t276 gnd.t274 gnd.t275 gnd.t179 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X33 a_n8964_8799.t18 a_n2982_13878.t66 a_n2982_8322.t22 vdd.t40 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X34 vdd.t183 a_n8964_8799.t48 CSoutput.t87 vdd.t76 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X35 a_n2982_13878.t63 minus.t5 a_n2903_n3924.t39 gnd.t344 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X36 vdd.t182 a_n8964_8799.t49 CSoutput.t86 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X37 a_n8964_8799.t19 a_n2982_13878.t67 a_n2982_8322.t21 vdd.t3 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X38 CSoutput.t202 commonsourceibias.t93 gnd.t354 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X39 gnd.t153 commonsourceibias.t94 CSoutput.t201 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X40 gnd.t273 gnd.t271 gnd.t272 gnd.t197 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X41 CSoutput.t200 commonsourceibias.t95 gnd.t143 gnd.t130 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X42 CSoutput.t199 commonsourceibias.t96 gnd.t139 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X43 a_n2903_n3924.t7 minus.t6 a_n2982_13878.t5 gnd.t94 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X44 gnd.t270 gnd.t268 minus.t4 gnd.t269 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X45 CSoutput.t198 commonsourceibias.t97 gnd.t161 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X46 a_n2903_n3924.t21 diffpairibias.t16 gnd.t341 gnd.t340 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X47 gnd.t45 commonsourceibias.t98 CSoutput.t197 gnd.t44 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X48 CSoutput.t85 a_n8964_8799.t50 vdd.t181 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X49 gnd.t32 commonsourceibias.t99 CSoutput.t196 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X50 gnd.t267 gnd.t265 gnd.t266 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X51 CSoutput.t195 commonsourceibias.t100 gnd.t317 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 vdd.t180 a_n8964_8799.t51 CSoutput.t84 vdd.t76 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X53 CSoutput.t194 commonsourceibias.t101 gnd.t318 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X54 gnd.t353 commonsourceibias.t76 commonsourceibias.t77 gnd.t49 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X55 CSoutput.t193 commonsourceibias.t102 gnd.t309 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X56 gnd.t295 commonsourceibias.t103 CSoutput.t192 gnd.t111 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X57 a_n2903_n3924.t26 plus.t7 a_n8964_8799.t35 gnd.t107 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X58 vdd.t179 a_n8964_8799.t52 CSoutput.t83 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X59 a_n2804_13878.t24 a_n2982_13878.t32 a_n2982_13878.t33 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X60 CSoutput.t191 commonsourceibias.t104 gnd.t63 gnd.t62 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X61 CSoutput.t190 commonsourceibias.t105 gnd.t154 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X62 gnd.t380 commonsourceibias.t106 CSoutput.t189 gnd.t111 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X63 vdd.t58 CSoutput.t218 output.t17 gnd.t101 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X64 a_n2982_13878.t21 a_n2982_13878.t20 a_n2804_13878.t23 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X65 CSoutput.t188 commonsourceibias.t107 gnd.t371 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X66 gnd.t125 commonsourceibias.t108 CSoutput.t187 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X67 CSoutput.t219 a_n2982_8322.t36 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X68 a_n8964_8799.t34 plus.t8 a_n2903_n3924.t27 gnd.t314 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X69 CSoutput.t82 a_n8964_8799.t53 vdd.t178 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X70 vdd.t268 vdd.t266 vdd.t267 vdd.t243 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X71 gnd.t60 commonsourceibias.t74 commonsourceibias.t75 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X72 vdd.t177 a_n8964_8799.t54 CSoutput.t81 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X73 CSoutput.t186 commonsourceibias.t109 gnd.t93 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X74 vdd.t175 a_n8964_8799.t55 CSoutput.t80 vdd.t129 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X75 gnd.t264 gnd.t262 gnd.t263 gnd.t197 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X76 CSoutput.t185 commonsourceibias.t110 gnd.t106 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X77 diffpairibias.t15 diffpairibias.t14 gnd.t397 gnd.t396 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X78 gnd.t120 commonsourceibias.t111 CSoutput.t184 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X79 a_n2982_13878.t0 minus.t7 a_n2903_n3924.t0 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X80 a_n2982_13878.t17 a_n2982_13878.t16 a_n2804_13878.t22 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X81 CSoutput.t183 commonsourceibias.t112 gnd.t46 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X82 CSoutput.t79 a_n8964_8799.t56 vdd.t174 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X83 CSoutput.t182 commonsourceibias.t113 gnd.t64 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X84 gnd.t126 commonsourceibias.t114 CSoutput.t181 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 a_n8964_8799.t9 a_n2982_13878.t68 a_n2982_8322.t20 vdd.t34 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X86 gnd.t296 commonsourceibias.t115 CSoutput.t180 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X87 vdd.t173 a_n8964_8799.t57 CSoutput.t78 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X88 CSoutput.t77 a_n8964_8799.t58 vdd.t172 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X89 gnd.t395 commonsourceibias.t116 CSoutput.t179 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 a_n2982_13878.t31 a_n2982_13878.t30 a_n2804_13878.t21 vdd.t55 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X91 vdd.t171 a_n8964_8799.t59 CSoutput.t76 vdd.t84 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X92 vdd.t170 a_n8964_8799.t60 CSoutput.t75 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X93 a_n8964_8799.t1 a_n2982_13878.t69 a_n2982_8322.t19 vdd.t32 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X94 CSoutput.t178 commonsourceibias.t117 gnd.t372 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X95 diffpairibias.t13 diffpairibias.t12 gnd.t89 gnd.t88 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X96 CSoutput.t74 a_n8964_8799.t61 vdd.t169 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X97 gnd.t316 commonsourceibias.t72 commonsourceibias.t73 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X98 gnd.t157 commonsourceibias.t118 CSoutput.t177 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X99 a_n8964_8799.t16 a_n2982_13878.t70 a_n2982_8322.t18 vdd.t47 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X100 CSoutput.t176 commonsourceibias.t119 gnd.t48 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X101 gnd.t95 commonsourceibias.t120 CSoutput.t175 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X102 CSoutput.t174 commonsourceibias.t121 gnd.t109 gnd.t108 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X103 CSoutput.t173 commonsourceibias.t122 gnd.t17 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X104 a_n2982_8322.t17 a_n2982_13878.t71 a_n8964_8799.t14 vdd.t55 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X105 CSoutput.t172 commonsourceibias.t123 gnd.t121 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X106 gnd.t381 commonsourceibias.t124 CSoutput.t171 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X107 CSoutput.t73 a_n8964_8799.t62 vdd.t168 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X108 gnd.t315 commonsourceibias.t70 commonsourceibias.t71 gnd.t72 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X109 gnd.t398 commonsourceibias.t68 commonsourceibias.t69 gnd.t44 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X110 CSoutput.t170 commonsourceibias.t125 gnd.t55 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X111 vdd.t59 CSoutput.t220 output.t16 gnd.t102 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X112 output.t15 CSoutput.t221 vdd.t0 gnd.t90 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X113 CSoutput.t169 commonsourceibias.t126 gnd.t158 gnd.t62 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X114 a_n2903_n3924.t24 plus.t9 a_n8964_8799.t33 gnd.t313 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X115 gnd.t248 gnd.t246 minus.t3 gnd.t247 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X116 gnd.t382 commonsourceibias.t127 CSoutput.t168 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X117 vdd.t265 vdd.t263 vdd.t264 vdd.t239 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X118 a_n2903_n3924.t9 diffpairibias.t17 gnd.t116 gnd.t115 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X119 CSoutput.t222 a_n2982_8322.t35 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X120 vdd.t167 a_n8964_8799.t63 CSoutput.t72 vdd.t127 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X121 gnd.t261 gnd.t259 gnd.t260 gnd.t175 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X122 vdd.t166 a_n8964_8799.t64 CSoutput.t71 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X123 a_n2982_13878.t23 a_n2982_13878.t22 a_n2804_13878.t20 vdd.t54 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X124 vdd.t165 a_n8964_8799.t65 CSoutput.t70 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X125 gnd.t4 commonsourceibias.t128 CSoutput.t167 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X126 gnd.t258 gnd.t255 gnd.t257 gnd.t256 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X127 a_n8964_8799.t39 a_n2982_13878.t72 a_n2982_8322.t16 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X128 a_n2982_13878.t9 a_n2982_13878.t8 a_n2804_13878.t19 vdd.t6 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X129 gnd.t254 gnd.t252 gnd.t253 gnd.t175 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X130 gnd.t97 commonsourceibias.t129 CSoutput.t166 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X131 CSoutput.t165 commonsourceibias.t130 gnd.t110 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X132 commonsourceibias.t67 commonsourceibias.t66 gnd.t393 gnd.t62 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X133 CSoutput.t69 a_n8964_8799.t66 vdd.t164 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X134 gnd.t383 commonsourceibias.t131 CSoutput.t164 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X135 a_n2982_13878.t58 minus.t8 a_n2903_n3924.t15 gnd.t312 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X136 gnd.t19 commonsourceibias.t132 CSoutput.t163 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X137 vdd.t262 vdd.t260 vdd.t261 vdd.t250 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X138 gnd.t308 commonsourceibias.t64 commonsourceibias.t65 gnd.t123 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X139 gnd.t50 commonsourceibias.t133 CSoutput.t162 gnd.t49 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X140 CSoutput.t68 a_n8964_8799.t67 vdd.t163 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X141 vdd.t259 vdd.t256 vdd.t258 vdd.t257 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X142 gnd.t251 gnd.t249 gnd.t250 gnd.t193 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X143 a_n2804_13878.t18 a_n2982_13878.t18 a_n2982_13878.t19 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X144 a_n2903_n3924.t5 minus.t9 a_n2982_13878.t4 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X145 CSoutput.t67 a_n8964_8799.t68 vdd.t162 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X146 gnd.t245 gnd.t243 gnd.t244 gnd.t179 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X147 vdd.t161 a_n8964_8799.t69 CSoutput.t66 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X148 vdd.t53 a_n2982_13878.t73 a_n2982_8322.t31 vdd.t52 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X149 a_n2982_13878.t49 a_n2982_13878.t48 a_n2804_13878.t17 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X150 CSoutput.t161 commonsourceibias.t134 gnd.t57 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X151 a_n2982_8322.t30 a_n2982_13878.t74 vdd.t51 vdd.t50 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X152 gnd.t99 commonsourceibias.t135 CSoutput.t160 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X153 a_n2903_n3924.t18 diffpairibias.t18 gnd.t333 gnd.t332 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X154 output.t14 CSoutput.t223 vdd.t1 gnd.t91 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X155 CSoutput.t65 a_n8964_8799.t70 vdd.t160 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X156 vdd.t269 CSoutput.t224 output.t13 gnd.t361 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X157 gnd.t112 commonsourceibias.t136 CSoutput.t159 gnd.t111 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X158 gnd.t79 commonsourceibias.t62 commonsourceibias.t63 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X159 CSoutput.t158 commonsourceibias.t137 gnd.t122 gnd.t108 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X160 gnd.t100 commonsourceibias.t138 CSoutput.t157 gnd.t72 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X161 CSoutput.t156 commonsourceibias.t139 gnd.t6 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X162 CSoutput.t155 commonsourceibias.t140 gnd.t297 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X163 CSoutput.t154 commonsourceibias.t141 gnd.t21 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X164 a_n2903_n3924.t19 minus.t10 a_n2982_13878.t61 gnd.t334 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X165 gnd.t242 gnd.t240 plus.t4 gnd.t241 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X166 vdd.t49 a_n2982_13878.t75 a_n2804_13878.t29 vdd.t48 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X167 vdd.t255 vdd.t253 vdd.t254 vdd.t239 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X168 a_n2903_n3924.t37 plus.t10 a_n8964_8799.t32 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X169 vdd.t252 vdd.t249 vdd.t251 vdd.t250 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X170 vdd.t159 a_n8964_8799.t71 CSoutput.t64 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X171 vdd.t270 CSoutput.t225 output.t12 gnd.t362 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X172 gnd.t239 gnd.t237 gnd.t238 gnd.t175 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X173 a_n2804_13878.t16 a_n2982_13878.t10 a_n2982_13878.t11 vdd.t47 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X174 vdd.t157 a_n8964_8799.t72 CSoutput.t63 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X175 a_n2982_8322.t15 a_n2982_13878.t76 a_n8964_8799.t12 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X176 a_n8964_8799.t31 plus.t11 a_n2903_n3924.t22 gnd.t155 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X177 a_n8964_8799.t30 plus.t12 a_n2903_n3924.t36 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X178 vdd.t248 vdd.t246 vdd.t247 vdd.t216 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X179 vdd.t245 vdd.t242 vdd.t244 vdd.t243 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X180 a_n2982_8322.t29 a_n2982_13878.t77 vdd.t46 vdd.t45 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X181 a_n8964_8799.t15 a_n2982_13878.t78 a_n2982_8322.t14 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X182 CSoutput.t62 a_n8964_8799.t73 vdd.t156 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X183 diffpairibias.t11 diffpairibias.t10 gnd.t147 gnd.t146 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X184 vdd.t155 a_n8964_8799.t74 CSoutput.t61 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X185 a_n2982_13878.t57 minus.t11 a_n2903_n3924.t13 gnd.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X186 a_n2982_13878.t43 a_n2982_13878.t42 a_n2804_13878.t15 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X187 CSoutput.t153 commonsourceibias.t142 gnd.t373 gnd.t103 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X188 a_n8964_8799.t38 a_n2982_13878.t79 a_n2982_8322.t13 vdd.t44 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X189 CSoutput.t60 a_n8964_8799.t75 vdd.t153 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X190 CSoutput.t59 a_n8964_8799.t76 vdd.t151 vdd.t122 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X191 commonsourceibias.t61 commonsourceibias.t60 gnd.t159 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X192 output.t11 CSoutput.t226 vdd.t271 gnd.t363 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X193 gnd.t51 commonsourceibias.t143 CSoutput.t152 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X194 a_n2804_13878.t14 a_n2982_13878.t46 a_n2982_13878.t47 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X195 gnd.t369 commonsourceibias.t58 commonsourceibias.t59 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 a_n2903_n3924.t3 minus.t12 a_n2982_13878.t3 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X197 CSoutput.t151 commonsourceibias.t144 gnd.t81 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X198 minus.t2 gnd.t234 gnd.t236 gnd.t235 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X199 vdd.t241 vdd.t238 vdd.t240 vdd.t239 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X200 vdd.t237 vdd.t235 vdd.t236 vdd.t212 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X201 vdd.t234 vdd.t232 vdd.t233 vdd.t198 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X202 CSoutput.t58 a_n8964_8799.t77 vdd.t150 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X203 output.t10 CSoutput.t227 vdd.t273 gnd.t384 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X204 CSoutput.t150 commonsourceibias.t145 gnd.t127 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X205 vdd.t42 a_n2982_13878.t80 a_n2982_8322.t28 vdd.t41 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X206 a_n2804_13878.t13 a_n2982_13878.t36 a_n2982_13878.t37 vdd.t40 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X207 vdd.t149 a_n8964_8799.t78 CSoutput.t57 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X208 vdd.t148 a_n8964_8799.t79 CSoutput.t56 vdd.t138 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X209 gnd.t82 commonsourceibias.t146 CSoutput.t149 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X210 gnd.t128 commonsourceibias.t147 CSoutput.t148 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X211 a_n2982_13878.t15 a_n2982_13878.t14 a_n2804_13878.t12 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X212 gnd.t319 commonsourceibias.t148 CSoutput.t147 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X213 gnd.t320 commonsourceibias.t149 CSoutput.t146 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X214 commonsourceibias.t57 commonsourceibias.t56 gnd.t378 gnd.t108 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X215 gnd.t83 commonsourceibias.t150 CSoutput.t145 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X216 gnd.t233 gnd.t231 gnd.t232 gnd.t183 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X217 gnd.t53 commonsourceibias.t151 CSoutput.t144 gnd.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X218 vdd.t143 a_n8964_8799.t80 CSoutput.t55 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X219 CSoutput.t143 commonsourceibias.t152 gnd.t359 gnd.t130 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X220 a_n2903_n3924.t4 diffpairibias.t19 gnd.t37 gnd.t36 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X221 gnd.t230 gnd.t227 gnd.t229 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X222 a_n2903_n3924.t20 diffpairibias.t20 gnd.t339 gnd.t338 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X223 commonsourceibias.t55 commonsourceibias.t54 gnd.t138 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X224 vdd.t147 a_n8964_8799.t81 CSoutput.t54 vdd.t138 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X225 vdd.t146 a_n8964_8799.t82 CSoutput.t53 vdd.t127 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X226 CSoutput.t52 a_n8964_8799.t83 vdd.t145 vdd.t80 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X227 gnd.t226 gnd.t224 gnd.t225 gnd.t197 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X228 vdd.t231 vdd.t229 vdd.t230 vdd.t216 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X229 CSoutput.t142 commonsourceibias.t153 gnd.t355 gnd.t103 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X230 CSoutput.t141 commonsourceibias.t154 gnd.t321 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X231 a_n2804_13878.t11 a_n2982_13878.t26 a_n2982_13878.t27 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X232 CSoutput.t51 a_n8964_8799.t84 vdd.t144 vdd.t122 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X233 commonsourceibias.t53 commonsourceibias.t52 gnd.t142 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X234 gnd.t223 gnd.t220 gnd.t222 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X235 a_n2982_8322.t12 a_n2982_13878.t81 a_n8964_8799.t5 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X236 output.t1 outputibias.t8 gnd.t141 gnd.t140 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X237 CSoutput.t50 a_n8964_8799.t85 vdd.t142 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X238 CSoutput.t140 commonsourceibias.t155 gnd.t84 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X239 commonsourceibias.t51 commonsourceibias.t50 gnd.t152 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X240 CSoutput.t139 commonsourceibias.t156 gnd.t129 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X241 outputibias.t7 outputibias.t6 gnd.t390 gnd.t389 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X242 gnd.t350 commonsourceibias.t48 commonsourceibias.t49 gnd.t111 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X243 vdd.t274 CSoutput.t228 output.t9 gnd.t385 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X244 diffpairibias.t9 diffpairibias.t8 gnd.t375 gnd.t374 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X245 a_n2804_13878.t31 a_n2982_13878.t82 vdd.t38 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X246 output.t2 outputibias.t9 gnd.t150 gnd.t149 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X247 vdd.t36 a_n2982_13878.t83 a_n2804_13878.t28 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X248 CSoutput.t138 commonsourceibias.t157 gnd.t131 gnd.t130 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X249 CSoutput.t137 commonsourceibias.t158 gnd.t328 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X250 CSoutput.t49 a_n8964_8799.t86 vdd.t141 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X251 CSoutput.t136 commonsourceibias.t159 gnd.t300 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X252 gnd.t29 commonsourceibias.t46 commonsourceibias.t47 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X253 vdd.t139 a_n8964_8799.t87 CSoutput.t48 vdd.t138 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X254 vdd.t137 a_n8964_8799.t88 CSoutput.t47 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X255 gnd.t219 gnd.t216 gnd.t218 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X256 gnd.t215 gnd.t213 plus.t2 gnd.t214 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X257 outputibias.t5 outputibias.t4 gnd.t368 gnd.t367 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X258 vdd.t135 a_n8964_8799.t89 CSoutput.t46 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X259 commonsourceibias.t45 commonsourceibias.t44 gnd.t78 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X260 gnd.t66 commonsourceibias.t160 CSoutput.t135 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X261 CSoutput.t45 a_n8964_8799.t90 vdd.t133 vdd.t112 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X262 a_n2804_13878.t10 a_n2982_13878.t6 a_n2982_13878.t7 vdd.t34 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X263 gnd.t299 commonsourceibias.t42 commonsourceibias.t43 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X264 a_n2903_n3924.t8 minus.t13 a_n2982_13878.t54 gnd.t107 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X265 gnd.t329 commonsourceibias.t161 CSoutput.t134 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X266 commonsourceibias.t41 commonsourceibias.t40 gnd.t293 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X267 vdd.t132 a_n8964_8799.t91 CSoutput.t44 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X268 gnd.t307 commonsourceibias.t38 commonsourceibias.t39 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X269 a_n2982_8322.t11 a_n2982_13878.t84 a_n8964_8799.t6 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X270 a_n2982_13878.t29 a_n2982_13878.t28 a_n2804_13878.t9 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X271 CSoutput.t133 commonsourceibias.t162 gnd.t301 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X272 CSoutput.t43 a_n8964_8799.t92 vdd.t131 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X273 diffpairibias.t7 diffpairibias.t6 gnd.t114 gnd.t113 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X274 vdd.t130 a_n8964_8799.t93 CSoutput.t42 vdd.t129 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X275 a_n2804_13878.t8 a_n2982_13878.t24 a_n2982_13878.t25 vdd.t32 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X276 commonsourceibias.t37 commonsourceibias.t36 gnd.t27 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X277 a_n2982_13878.t60 minus.t14 a_n2903_n3924.t17 gnd.t314 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X278 a_n2982_13878.t55 minus.t15 a_n2903_n3924.t10 gnd.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X279 gnd.t212 gnd.t210 gnd.t211 gnd.t183 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X280 vdd.t31 a_n2982_13878.t85 a_n2982_8322.t27 vdd.t30 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X281 vdd.t128 a_n8964_8799.t94 CSoutput.t41 vdd.t127 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X282 a_n8964_8799.t29 plus.t13 a_n2903_n3924.t23 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X283 gnd.t68 commonsourceibias.t163 CSoutput.t132 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X284 CSoutput.t40 a_n8964_8799.t95 vdd.t126 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X285 a_n2903_n3924.t38 minus.t16 a_n2982_13878.t62 gnd.t345 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X286 gnd.t1 commonsourceibias.t34 commonsourceibias.t35 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X287 CSoutput.t131 commonsourceibias.t164 gnd.t330 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X288 a_n2804_13878.t0 a_n2982_13878.t86 vdd.t29 vdd.t28 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X289 vdd.t228 vdd.t226 vdd.t227 vdd.t212 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X290 vdd.t125 a_n8964_8799.t96 CSoutput.t39 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X291 output.t8 CSoutput.t229 vdd.t275 gnd.t386 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X292 CSoutput.t38 a_n8964_8799.t97 vdd.t123 vdd.t122 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X293 CSoutput.t37 a_n8964_8799.t98 vdd.t121 vdd.t112 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X294 gnd.t70 commonsourceibias.t165 CSoutput.t130 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X295 vdd.t120 a_n8964_8799.t99 CSoutput.t36 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X296 gnd.t209 gnd.t206 gnd.t208 gnd.t207 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X297 vdd.t225 vdd.t223 vdd.t224 vdd.t202 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X298 a_n2903_n3924.t14 diffpairibias.t21 gnd.t311 gnd.t310 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X299 a_n2982_8322.t10 a_n2982_13878.t87 a_n8964_8799.t17 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X300 vdd.t26 a_n2982_13878.t88 a_n2982_8322.t26 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X301 CSoutput.t230 a_n2982_8322.t34 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X302 gnd.t306 commonsourceibias.t32 commonsourceibias.t33 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X303 outputibias.t3 outputibias.t2 gnd.t392 gnd.t391 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X304 vdd.t119 a_n8964_8799.t100 CSoutput.t35 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X305 a_n8964_8799.t28 plus.t14 a_n2903_n3924.t30 gnd.t344 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X306 output.t19 outputibias.t10 gnd.t349 gnd.t348 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X307 gnd.t205 gnd.t203 plus.t1 gnd.t204 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X308 gnd.t366 commonsourceibias.t30 commonsourceibias.t31 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X309 vdd.t222 vdd.t219 vdd.t221 vdd.t220 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X310 CSoutput.t129 commonsourceibias.t166 gnd.t357 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X311 a_n2903_n3924.t28 plus.t15 a_n8964_8799.t27 gnd.t94 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X312 vdd.t118 a_n8964_8799.t101 CSoutput.t34 vdd.t74 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X313 gnd.t202 gnd.t200 gnd.t201 gnd.t179 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X314 vdd.t192 CSoutput.t231 output.t7 gnd.t289 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X315 CSoutput.t33 a_n8964_8799.t102 vdd.t117 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X316 CSoutput.t128 commonsourceibias.t167 gnd.t351 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X317 CSoutput.t32 a_n8964_8799.t103 vdd.t69 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X318 CSoutput.t31 a_n8964_8799.t104 vdd.t115 vdd.t101 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X319 a_n2804_13878.t7 a_n2982_13878.t34 a_n2982_13878.t35 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X320 a_n2982_8322.t9 a_n2982_13878.t89 a_n8964_8799.t4 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X321 diffpairibias.t5 diffpairibias.t4 gnd.t23 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X322 CSoutput.t232 a_n2982_8322.t33 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X323 gnd.t199 gnd.t196 gnd.t198 gnd.t197 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X324 CSoutput.t30 a_n8964_8799.t105 vdd.t110 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X325 CSoutput.t29 a_n8964_8799.t106 vdd.t114 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X326 gnd.t388 commonsourceibias.t28 commonsourceibias.t29 gnd.t98 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X327 output.t6 CSoutput.t233 vdd.t61 gnd.t135 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X328 vdd.t218 vdd.t215 vdd.t217 vdd.t216 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X329 vdd.t214 vdd.t211 vdd.t213 vdd.t212 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X330 CSoutput.t127 commonsourceibias.t168 gnd.t33 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X331 commonsourceibias.t27 commonsourceibias.t26 gnd.t292 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X332 a_n2982_8322.t25 a_n2982_13878.t90 vdd.t23 vdd.t22 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X333 CSoutput.t28 a_n8964_8799.t107 vdd.t113 vdd.t112 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X334 gnd.t195 gnd.t192 gnd.t194 gnd.t193 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X335 vdd.t111 a_n8964_8799.t108 CSoutput.t27 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X336 gnd.t85 commonsourceibias.t169 CSoutput.t126 gnd.t49 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X337 CSoutput.t26 a_n8964_8799.t109 vdd.t108 vdd.t82 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X338 vdd.t21 a_n2982_13878.t91 a_n2804_13878.t26 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X339 vdd.t73 a_n8964_8799.t110 CSoutput.t25 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X340 CSoutput.t24 a_n8964_8799.t111 vdd.t107 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X341 vdd.t105 a_n8964_8799.t112 CSoutput.t23 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X342 gnd.t132 commonsourceibias.t170 CSoutput.t125 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X343 gnd.t322 commonsourceibias.t171 CSoutput.t124 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X344 output.t5 CSoutput.t234 vdd.t62 gnd.t136 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X345 a_n2982_8322.t8 a_n2982_13878.t92 a_n8964_8799.t7 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X346 commonsourceibias.t25 commonsourceibias.t24 gnd.t305 gnd.t103 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X347 gnd.t191 gnd.t189 minus.t1 gnd.t190 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X348 a_n8964_8799.t2 a_n2982_13878.t93 a_n2982_8322.t7 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X349 a_n2804_13878.t27 a_n2982_13878.t94 vdd.t18 vdd.t17 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X350 gnd.t323 commonsourceibias.t172 CSoutput.t123 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X351 vdd.t210 vdd.t208 vdd.t209 vdd.t194 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X352 vdd.t103 a_n8964_8799.t113 CSoutput.t22 vdd.t84 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X353 a_n2982_13878.t56 minus.t17 a_n2903_n3924.t12 gnd.t155 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X354 CSoutput.t21 a_n8964_8799.t114 vdd.t102 vdd.t101 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X355 CSoutput.t20 a_n8964_8799.t115 vdd.t100 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X356 CSoutput.t19 a_n8964_8799.t116 vdd.t99 vdd.t80 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X357 commonsourceibias.t23 commonsourceibias.t22 gnd.t365 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X358 a_n2982_13878.t13 a_n2982_13878.t12 a_n2804_13878.t6 vdd.t7 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X359 a_n8964_8799.t13 a_n2982_13878.t95 a_n2982_8322.t6 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X360 output.t4 CSoutput.t235 vdd.t63 gnd.t137 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X361 minus.t0 gnd.t186 gnd.t188 gnd.t187 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X362 a_n8964_8799.t20 a_n2982_13878.t96 a_n2982_8322.t5 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X363 gnd.t185 gnd.t182 gnd.t184 gnd.t183 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X364 gnd.t87 commonsourceibias.t173 CSoutput.t122 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X365 a_n2982_8322.t4 a_n2982_13878.t97 a_n8964_8799.t21 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X366 commonsourceibias.t21 commonsourceibias.t20 gnd.t387 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X367 a_n8964_8799.t26 plus.t16 a_n2903_n3924.t32 gnd.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X368 gnd.t59 commonsourceibias.t174 CSoutput.t121 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X369 CSoutput.t120 commonsourceibias.t175 gnd.t360 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X370 a_n2903_n3924.t16 minus.t18 a_n2982_13878.t59 gnd.t313 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X371 vdd.t98 a_n8964_8799.t117 CSoutput.t18 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X372 gnd.t291 commonsourceibias.t18 commonsourceibias.t19 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X373 CSoutput.t17 a_n8964_8799.t118 vdd.t95 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X374 CSoutput.t16 a_n8964_8799.t119 vdd.t96 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X375 CSoutput.t15 a_n8964_8799.t120 vdd.t93 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X376 a_n2804_13878.t5 a_n2982_13878.t38 a_n2982_13878.t39 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X377 outputibias.t1 outputibias.t0 gnd.t327 gnd.t326 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X378 vdd.t92 a_n8964_8799.t121 CSoutput.t14 vdd.t78 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X379 a_n2903_n3924.t29 plus.t17 a_n8964_8799.t25 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X380 gnd.t364 commonsourceibias.t16 commonsourceibias.t17 gnd.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X381 commonsourceibias.t15 commonsourceibias.t14 gnd.t377 gnd.t130 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X382 gnd.t181 gnd.t178 gnd.t180 gnd.t179 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X383 gnd.t356 commonsourceibias.t176 CSoutput.t119 gnd.t72 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X384 gnd.t133 commonsourceibias.t177 CSoutput.t118 gnd.t44 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X385 a_n2903_n3924.t11 diffpairibias.t22 gnd.t145 gnd.t144 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X386 gnd.t324 commonsourceibias.t178 CSoutput.t117 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X387 vdd.t91 a_n8964_8799.t122 CSoutput.t13 vdd.t74 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X388 CSoutput.t116 commonsourceibias.t179 gnd.t134 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X389 gnd.t337 commonsourceibias.t180 CSoutput.t115 gnd.t49 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X390 CSoutput.t12 a_n8964_8799.t123 vdd.t90 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X391 CSoutput.t114 commonsourceibias.t181 gnd.t9 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X392 a_n2982_13878.t51 a_n2982_13878.t50 a_n2804_13878.t4 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X393 gnd.t177 gnd.t174 gnd.t176 gnd.t175 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X394 a_n8964_8799.t11 a_n2982_13878.t98 a_n2982_8322.t3 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X395 vdd.t272 CSoutput.t236 output.t3 gnd.t376 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X396 vdd.t89 a_n8964_8799.t124 CSoutput.t11 vdd.t78 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X397 CSoutput.t10 a_n8964_8799.t125 vdd.t88 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X398 vdd.t207 vdd.t205 vdd.t206 vdd.t202 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X399 a_n8964_8799.t24 plus.t18 a_n2903_n3924.t25 gnd.t312 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X400 CSoutput.t113 commonsourceibias.t182 gnd.t35 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X401 gnd.t71 commonsourceibias.t183 CSoutput.t112 gnd.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X402 commonsourceibias.t13 commonsourceibias.t12 gnd.t148 gnd.t16 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X403 CSoutput.t111 commonsourceibias.t184 gnd.t331 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X404 CSoutput.t9 a_n8964_8799.t126 vdd.t86 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X405 gnd.t173 gnd.t170 gnd.t172 gnd.t171 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X406 diffpairibias.t3 diffpairibias.t2 gnd.t336 gnd.t335 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X407 a_n2982_8322.t2 a_n2982_13878.t99 a_n8964_8799.t3 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X408 CSoutput.t110 commonsourceibias.t185 gnd.t302 gnd.t62 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X409 gnd.t303 commonsourceibias.t186 CSoutput.t109 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X410 a_n2903_n3924.t34 plus.t19 a_n8964_8799.t23 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X411 vdd.t85 a_n8964_8799.t127 CSoutput.t8 vdd.t84 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X412 CSoutput.t7 a_n8964_8799.t128 vdd.t81 vdd.t80 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X413 CSoutput.t6 a_n8964_8799.t129 vdd.t83 vdd.t82 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X414 diffpairibias.t1 diffpairibias.t0 gnd.t288 gnd.t287 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X415 gnd.t73 commonsourceibias.t187 CSoutput.t108 gnd.t72 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X416 CSoutput.t237 a_n2982_8322.t32 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X417 commonsourceibias.t11 commonsourceibias.t10 gnd.t347 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X418 gnd.t342 commonsourceibias.t188 CSoutput.t107 gnd.t123 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X419 a_n2903_n3924.t33 plus.t20 a_n8964_8799.t22 gnd.t334 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X420 commonsourceibias.t9 commonsourceibias.t8 gnd.t25 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X421 CSoutput.t106 commonsourceibias.t189 gnd.t39 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X422 vdd.t9 a_n2982_13878.t100 a_n2804_13878.t1 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X423 CSoutput.t5 a_n8964_8799.t130 vdd.t71 vdd.t70 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X424 gnd.t76 commonsourceibias.t6 commonsourceibias.t7 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X425 a_n2903_n3924.t1 minus.t19 a_n2982_13878.t1 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X426 vdd.t79 a_n8964_8799.t131 CSoutput.t4 vdd.t78 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X427 gnd.t298 commonsourceibias.t4 commonsourceibias.t5 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X428 a_n2982_8322.t1 a_n2982_13878.t101 a_n8964_8799.t10 vdd.t7 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X429 gnd.t343 commonsourceibias.t190 CSoutput.t105 gnd.t69 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X430 a_n2982_13878.t2 minus.t20 a_n2903_n3924.t2 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X431 commonsourceibias.t3 commonsourceibias.t2 gnd.t290 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X432 gnd.t358 commonsourceibias.t191 CSoutput.t104 gnd.t44 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X433 gnd.t352 commonsourceibias.t192 CSoutput.t103 gnd.t123 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X434 gnd.t41 commonsourceibias.t193 CSoutput.t102 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X435 a_n2982_8322.t0 a_n2982_13878.t102 a_n8964_8799.t8 vdd.t6 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X436 vdd.t75 a_n8964_8799.t132 CSoutput.t3 vdd.t74 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X437 vdd.t77 a_n8964_8799.t133 CSoutput.t2 vdd.t76 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X438 output.t0 outputibias.t11 gnd.t13 gnd.t12 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X439 CSoutput.t1 a_n8964_8799.t134 vdd.t67 vdd.t66 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X440 gnd.t11 commonsourceibias.t194 CSoutput.t101 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X441 plus.t0 gnd.t167 gnd.t169 gnd.t168 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X442 vdd.t204 vdd.t201 vdd.t203 vdd.t202 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X443 a_n2982_8322.t24 a_n2982_13878.t103 vdd.t5 vdd.t4 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X444 gnd.t163 commonsourceibias.t195 CSoutput.t100 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X445 a_n2804_13878.t3 a_n2982_13878.t40 a_n2982_13878.t41 vdd.t3 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X446 gnd.t164 commonsourceibias.t196 CSoutput.t99 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X447 CSoutput.t98 commonsourceibias.t197 gnd.t165 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X448 commonsourceibias.t1 commonsourceibias.t0 gnd.t325 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X449 CSoutput.t97 commonsourceibias.t198 gnd.t166 gnd.t30 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X450 vdd.t200 vdd.t197 vdd.t199 vdd.t198 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X451 a_n2903_n3924.t6 diffpairibias.t23 gnd.t75 gnd.t74 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X452 vdd.t196 vdd.t193 vdd.t195 vdd.t194 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X453 CSoutput.t0 a_n8964_8799.t135 vdd.t65 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X454 a_n2982_13878.t53 a_n2982_13878.t52 a_n2804_13878.t2 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X455 gnd.t304 commonsourceibias.t199 CSoutput.t96 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
R0 plus.n33 plus.t15 321.495
R1 plus.n7 plus.t12 321.495
R2 plus.n32 plus.t14 297.12
R3 plus.n36 plus.t19 297.12
R4 plus.n38 plus.t18 297.12
R5 plus.n42 plus.t20 297.12
R6 plus.n44 plus.t8 297.12
R7 plus.n48 plus.t7 297.12
R8 plus.n50 plus.t11 297.12
R9 plus.n24 plus.t9 297.12
R10 plus.n22 plus.t5 297.12
R11 plus.n2 plus.t6 297.12
R12 plus.n16 plus.t16 297.12
R13 plus.n4 plus.t17 297.12
R14 plus.n10 plus.t13 297.12
R15 plus.n6 plus.t10 297.12
R16 plus.n54 plus.t4 243.97
R17 plus.n54 plus.n53 223.454
R18 plus.n56 plus.n55 223.454
R19 plus.n51 plus.n50 161.3
R20 plus.n49 plus.n26 161.3
R21 plus.n48 plus.n47 161.3
R22 plus.n46 plus.n27 161.3
R23 plus.n45 plus.n44 161.3
R24 plus.n43 plus.n28 161.3
R25 plus.n42 plus.n41 161.3
R26 plus.n40 plus.n29 161.3
R27 plus.n39 plus.n38 161.3
R28 plus.n37 plus.n30 161.3
R29 plus.n36 plus.n35 161.3
R30 plus.n34 plus.n31 161.3
R31 plus.n9 plus.n8 161.3
R32 plus.n10 plus.n5 161.3
R33 plus.n12 plus.n11 161.3
R34 plus.n13 plus.n4 161.3
R35 plus.n15 plus.n14 161.3
R36 plus.n16 plus.n3 161.3
R37 plus.n18 plus.n17 161.3
R38 plus.n19 plus.n2 161.3
R39 plus.n21 plus.n20 161.3
R40 plus.n22 plus.n1 161.3
R41 plus.n23 plus.n0 161.3
R42 plus.n25 plus.n24 161.3
R43 plus.n34 plus.n33 44.9377
R44 plus.n8 plus.n7 44.9377
R45 plus.n50 plus.n49 37.246
R46 plus.n24 plus.n23 37.246
R47 plus.n32 plus.n31 32.8641
R48 plus.n48 plus.n27 32.8641
R49 plus.n22 plus.n21 32.8641
R50 plus.n9 plus.n6 32.8641
R51 plus.n52 plus.n51 30.0327
R52 plus.n37 plus.n36 28.4823
R53 plus.n44 plus.n43 28.4823
R54 plus.n17 plus.n2 28.4823
R55 plus.n11 plus.n10 28.4823
R56 plus.n38 plus.n29 24.1005
R57 plus.n42 plus.n29 24.1005
R58 plus.n16 plus.n15 24.1005
R59 plus.n15 plus.n4 24.1005
R60 plus.n53 plus.t2 19.8005
R61 plus.n53 plus.t3 19.8005
R62 plus.n55 plus.t1 19.8005
R63 plus.n55 plus.t0 19.8005
R64 plus.n38 plus.n37 19.7187
R65 plus.n43 plus.n42 19.7187
R66 plus.n17 plus.n16 19.7187
R67 plus.n11 plus.n4 19.7187
R68 plus.n33 plus.n32 17.0522
R69 plus.n7 plus.n6 17.0522
R70 plus.n36 plus.n31 15.3369
R71 plus.n44 plus.n27 15.3369
R72 plus.n21 plus.n2 15.3369
R73 plus.n10 plus.n9 15.3369
R74 plus plus.n57 14.6484
R75 plus.n52 plus.n25 11.8547
R76 plus.n49 plus.n48 10.955
R77 plus.n23 plus.n22 10.955
R78 plus.n57 plus.n56 5.40567
R79 plus.n57 plus.n52 1.188
R80 plus.n56 plus.n54 0.716017
R81 plus.n35 plus.n34 0.189894
R82 plus.n35 plus.n30 0.189894
R83 plus.n39 plus.n30 0.189894
R84 plus.n40 plus.n39 0.189894
R85 plus.n41 plus.n40 0.189894
R86 plus.n41 plus.n28 0.189894
R87 plus.n45 plus.n28 0.189894
R88 plus.n46 plus.n45 0.189894
R89 plus.n47 plus.n46 0.189894
R90 plus.n47 plus.n26 0.189894
R91 plus.n51 plus.n26 0.189894
R92 plus.n25 plus.n0 0.189894
R93 plus.n1 plus.n0 0.189894
R94 plus.n20 plus.n1 0.189894
R95 plus.n20 plus.n19 0.189894
R96 plus.n19 plus.n18 0.189894
R97 plus.n18 plus.n3 0.189894
R98 plus.n14 plus.n3 0.189894
R99 plus.n14 plus.n13 0.189894
R100 plus.n13 plus.n12 0.189894
R101 plus.n12 plus.n5 0.189894
R102 plus.n8 plus.n5 0.189894
R103 a_n2903_n3924.n7 a_n2903_n3924.t14 214.994
R104 a_n2903_n3924.n4 a_n2903_n3924.t18 214.714
R105 a_n2903_n3924.n4 a_n2903_n3924.t11 214.321
R106 a_n2903_n3924.n5 a_n2903_n3924.t20 214.321
R107 a_n2903_n3924.n5 a_n2903_n3924.t6 214.321
R108 a_n2903_n3924.n6 a_n2903_n3924.t4 214.321
R109 a_n2903_n3924.n7 a_n2903_n3924.t21 214.321
R110 a_n2903_n3924.n7 a_n2903_n3924.t9 214.321
R111 a_n2903_n3924.n3 a_n2903_n3924.t28 55.8337
R112 a_n2903_n3924.n3 a_n2903_n3924.t2 55.8337
R113 a_n2903_n3924.n9 a_n2903_n3924.t16 55.8337
R114 a_n2903_n3924.n0 a_n2903_n3924.t22 55.8335
R115 a_n2903_n3924.n1 a_n2903_n3924.t12 55.8335
R116 a_n2903_n3924.n8 a_n2903_n3924.t7 55.8335
R117 a_n2903_n3924.n8 a_n2903_n3924.t36 55.8335
R118 a_n2903_n3924.n2 a_n2903_n3924.t24 55.8335
R119 a_n2903_n3924.n0 a_n2903_n3924.n20 53.0052
R120 a_n2903_n3924.n0 a_n2903_n3924.n21 53.0052
R121 a_n2903_n3924.n0 a_n2903_n3924.n22 53.0052
R122 a_n2903_n3924.n3 a_n2903_n3924.n10 53.0052
R123 a_n2903_n3924.n9 a_n2903_n3924.n11 53.0052
R124 a_n2903_n3924.n1 a_n2903_n3924.n18 53.0051
R125 a_n2903_n3924.n1 a_n2903_n3924.n17 53.0051
R126 a_n2903_n3924.n1 a_n2903_n3924.n16 53.0051
R127 a_n2903_n3924.n8 a_n2903_n3924.n15 53.0051
R128 a_n2903_n3924.n2 a_n2903_n3924.n14 53.0051
R129 a_n2903_n3924.n2 a_n2903_n3924.n13 53.0051
R130 a_n2903_n3924.n23 a_n2903_n3924.n3 53.0051
R131 a_n2903_n3924.n12 a_n2903_n3924.n9 12.1986
R132 a_n2903_n3924.n0 a_n2903_n3924.n19 12.1986
R133 a_n2903_n3924.n2 a_n2903_n3924.n12 5.11903
R134 a_n2903_n3924.n19 a_n2903_n3924.n1 5.11903
R135 a_n2903_n3924.n20 a_n2903_n3924.t27 2.82907
R136 a_n2903_n3924.n20 a_n2903_n3924.t26 2.82907
R137 a_n2903_n3924.n21 a_n2903_n3924.t25 2.82907
R138 a_n2903_n3924.n21 a_n2903_n3924.t33 2.82907
R139 a_n2903_n3924.n22 a_n2903_n3924.t30 2.82907
R140 a_n2903_n3924.n22 a_n2903_n3924.t34 2.82907
R141 a_n2903_n3924.n10 a_n2903_n3924.t13 2.82907
R142 a_n2903_n3924.n10 a_n2903_n3924.t3 2.82907
R143 a_n2903_n3924.n11 a_n2903_n3924.t10 2.82907
R144 a_n2903_n3924.n11 a_n2903_n3924.t38 2.82907
R145 a_n2903_n3924.n18 a_n2903_n3924.t17 2.82907
R146 a_n2903_n3924.n18 a_n2903_n3924.t8 2.82907
R147 a_n2903_n3924.n17 a_n2903_n3924.t15 2.82907
R148 a_n2903_n3924.n17 a_n2903_n3924.t19 2.82907
R149 a_n2903_n3924.n16 a_n2903_n3924.t39 2.82907
R150 a_n2903_n3924.n16 a_n2903_n3924.t5 2.82907
R151 a_n2903_n3924.n15 a_n2903_n3924.t23 2.82907
R152 a_n2903_n3924.n15 a_n2903_n3924.t37 2.82907
R153 a_n2903_n3924.n14 a_n2903_n3924.t32 2.82907
R154 a_n2903_n3924.n14 a_n2903_n3924.t29 2.82907
R155 a_n2903_n3924.n13 a_n2903_n3924.t35 2.82907
R156 a_n2903_n3924.n13 a_n2903_n3924.t31 2.82907
R157 a_n2903_n3924.t0 a_n2903_n3924.n23 2.82907
R158 a_n2903_n3924.n23 a_n2903_n3924.t1 2.82907
R159 a_n2903_n3924.n3 a_n2903_n3924.n0 2.45524
R160 a_n2903_n3924.n1 a_n2903_n3924.n8 2.01128
R161 a_n2903_n3924.n19 a_n2903_n3924.n4 1.95694
R162 a_n2903_n3924.n12 a_n2903_n3924.n7 1.95694
R163 a_n2903_n3924.n8 a_n2903_n3924.n2 1.77636
R164 a_n2903_n3924.n6 a_n2903_n3924.n5 1.34352
R165 a_n2903_n3924.n7 a_n2903_n3924.n6 1.34352
R166 a_n2903_n3924.n9 a_n2903_n3924.n3 1.3324
R167 a_n2903_n3924.n5 a_n2903_n3924.n4 0.951808
R168 a_n8964_8799.n183 a_n8964_8799.t116 485.149
R169 a_n8964_8799.n231 a_n8964_8799.t128 485.149
R170 a_n8964_8799.n280 a_n8964_8799.t83 485.149
R171 a_n8964_8799.n35 a_n8964_8799.t79 485.149
R172 a_n8964_8799.n83 a_n8964_8799.t87 485.149
R173 a_n8964_8799.n132 a_n8964_8799.t81 485.149
R174 a_n8964_8799.n215 a_n8964_8799.t47 464.166
R175 a_n8964_8799.n214 a_n8964_8799.t45 464.166
R176 a_n8964_8799.n170 a_n8964_8799.t113 464.166
R177 a_n8964_8799.n208 a_n8964_8799.t61 464.166
R178 a_n8964_8799.n207 a_n8964_8799.t49 464.166
R179 a_n8964_8799.n173 a_n8964_8799.t119 464.166
R180 a_n8964_8799.n201 a_n8964_8799.t82 464.166
R181 a_n8964_8799.n200 a_n8964_8799.t62 464.166
R182 a_n8964_8799.n176 a_n8964_8799.t133 464.166
R183 a_n8964_8799.n195 a_n8964_8799.t98 464.166
R184 a_n8964_8799.n193 a_n8964_8799.t64 464.166
R185 a_n8964_8799.n179 a_n8964_8799.t129 464.166
R186 a_n8964_8799.n188 a_n8964_8799.t100 464.166
R187 a_n8964_8799.n186 a_n8964_8799.t76 464.166
R188 a_n8964_8799.n182 a_n8964_8799.t46 464.166
R189 a_n8964_8799.n263 a_n8964_8799.t55 464.166
R190 a_n8964_8799.n262 a_n8964_8799.t53 464.166
R191 a_n8964_8799.n218 a_n8964_8799.t127 464.166
R192 a_n8964_8799.n256 a_n8964_8799.t67 464.166
R193 a_n8964_8799.n255 a_n8964_8799.t60 464.166
R194 a_n8964_8799.n221 a_n8964_8799.t130 464.166
R195 a_n8964_8799.n249 a_n8964_8799.t94 464.166
R196 a_n8964_8799.n248 a_n8964_8799.t70 464.166
R197 a_n8964_8799.n224 a_n8964_8799.t48 464.166
R198 a_n8964_8799.n243 a_n8964_8799.t107 464.166
R199 a_n8964_8799.n241 a_n8964_8799.t71 464.166
R200 a_n8964_8799.n227 a_n8964_8799.t41 464.166
R201 a_n8964_8799.n236 a_n8964_8799.t112 464.166
R202 a_n8964_8799.n234 a_n8964_8799.t84 464.166
R203 a_n8964_8799.n230 a_n8964_8799.t54 464.166
R204 a_n8964_8799.n312 a_n8964_8799.t93 464.166
R205 a_n8964_8799.n311 a_n8964_8799.t111 464.166
R206 a_n8964_8799.n267 a_n8964_8799.t59 464.166
R207 a_n8964_8799.n305 a_n8964_8799.t125 464.166
R208 a_n8964_8799.n304 a_n8964_8799.t74 464.166
R209 a_n8964_8799.n270 a_n8964_8799.t120 464.166
R210 a_n8964_8799.n298 a_n8964_8799.t63 464.166
R211 a_n8964_8799.n297 a_n8964_8799.t102 464.166
R212 a_n8964_8799.n273 a_n8964_8799.t51 464.166
R213 a_n8964_8799.n292 a_n8964_8799.t90 464.166
R214 a_n8964_8799.n290 a_n8964_8799.t69 464.166
R215 a_n8964_8799.n276 a_n8964_8799.t109 464.166
R216 a_n8964_8799.n285 a_n8964_8799.t57 464.166
R217 a_n8964_8799.n283 a_n8964_8799.t97 464.166
R218 a_n8964_8799.n279 a_n8964_8799.t44 464.166
R219 a_n8964_8799.n34 a_n8964_8799.t104 464.166
R220 a_n8964_8799.n38 a_n8964_8799.t42 464.166
R221 a_n8964_8799.n32 a_n8964_8799.t66 464.166
R222 a_n8964_8799.n43 a_n8964_8799.t99 464.166
R223 a_n8964_8799.n45 a_n8964_8799.t126 464.166
R224 a_n8964_8799.n49 a_n8964_8799.t65 464.166
R225 a_n8964_8799.n50 a_n8964_8799.t95 464.166
R226 a_n8964_8799.n28 a_n8964_8799.t122 464.166
R227 a_n8964_8799.n55 a_n8964_8799.t123 464.166
R228 a_n8964_8799.n57 a_n8964_8799.t80 464.166
R229 a_n8964_8799.n61 a_n8964_8799.t106 464.166
R230 a_n8964_8799.n62 a_n8964_8799.t121 464.166
R231 a_n8964_8799.n24 a_n8964_8799.t77 464.166
R232 a_n8964_8799.n68 a_n8964_8799.t78 464.166
R233 a_n8964_8799.n69 a_n8964_8799.t103 464.166
R234 a_n8964_8799.n82 a_n8964_8799.t114 464.166
R235 a_n8964_8799.n86 a_n8964_8799.t52 464.166
R236 a_n8964_8799.n80 a_n8964_8799.t75 464.166
R237 a_n8964_8799.n91 a_n8964_8799.t108 464.166
R238 a_n8964_8799.n93 a_n8964_8799.t135 464.166
R239 a_n8964_8799.n97 a_n8964_8799.t72 464.166
R240 a_n8964_8799.n98 a_n8964_8799.t105 464.166
R241 a_n8964_8799.n76 a_n8964_8799.t132 464.166
R242 a_n8964_8799.n103 a_n8964_8799.t134 464.166
R243 a_n8964_8799.n105 a_n8964_8799.t91 464.166
R244 a_n8964_8799.n109 a_n8964_8799.t118 464.166
R245 a_n8964_8799.n110 a_n8964_8799.t131 464.166
R246 a_n8964_8799.n72 a_n8964_8799.t86 464.166
R247 a_n8964_8799.n116 a_n8964_8799.t88 464.166
R248 a_n8964_8799.n117 a_n8964_8799.t115 464.166
R249 a_n8964_8799.n131 a_n8964_8799.t43 464.166
R250 a_n8964_8799.n135 a_n8964_8799.t96 464.166
R251 a_n8964_8799.n129 a_n8964_8799.t56 464.166
R252 a_n8964_8799.n140 a_n8964_8799.t110 464.166
R253 a_n8964_8799.n142 a_n8964_8799.t68 464.166
R254 a_n8964_8799.n146 a_n8964_8799.t89 464.166
R255 a_n8964_8799.n147 a_n8964_8799.t50 464.166
R256 a_n8964_8799.n125 a_n8964_8799.t101 464.166
R257 a_n8964_8799.n152 a_n8964_8799.t85 464.166
R258 a_n8964_8799.n154 a_n8964_8799.t117 464.166
R259 a_n8964_8799.n158 a_n8964_8799.t73 464.166
R260 a_n8964_8799.n159 a_n8964_8799.t124 464.166
R261 a_n8964_8799.n121 a_n8964_8799.t58 464.166
R262 a_n8964_8799.n165 a_n8964_8799.t40 464.166
R263 a_n8964_8799.n166 a_n8964_8799.t92 464.166
R264 a_n8964_8799.n185 a_n8964_8799.n184 161.3
R265 a_n8964_8799.n186 a_n8964_8799.n181 161.3
R266 a_n8964_8799.n187 a_n8964_8799.n180 161.3
R267 a_n8964_8799.n189 a_n8964_8799.n188 161.3
R268 a_n8964_8799.n190 a_n8964_8799.n179 161.3
R269 a_n8964_8799.n192 a_n8964_8799.n191 161.3
R270 a_n8964_8799.n193 a_n8964_8799.n178 161.3
R271 a_n8964_8799.n194 a_n8964_8799.n177 161.3
R272 a_n8964_8799.n196 a_n8964_8799.n195 161.3
R273 a_n8964_8799.n197 a_n8964_8799.n176 161.3
R274 a_n8964_8799.n199 a_n8964_8799.n198 161.3
R275 a_n8964_8799.n200 a_n8964_8799.n175 161.3
R276 a_n8964_8799.n201 a_n8964_8799.n174 161.3
R277 a_n8964_8799.n203 a_n8964_8799.n202 161.3
R278 a_n8964_8799.n204 a_n8964_8799.n173 161.3
R279 a_n8964_8799.n206 a_n8964_8799.n205 161.3
R280 a_n8964_8799.n207 a_n8964_8799.n172 161.3
R281 a_n8964_8799.n208 a_n8964_8799.n171 161.3
R282 a_n8964_8799.n210 a_n8964_8799.n209 161.3
R283 a_n8964_8799.n211 a_n8964_8799.n170 161.3
R284 a_n8964_8799.n213 a_n8964_8799.n212 161.3
R285 a_n8964_8799.n214 a_n8964_8799.n169 161.3
R286 a_n8964_8799.n216 a_n8964_8799.n215 161.3
R287 a_n8964_8799.n233 a_n8964_8799.n232 161.3
R288 a_n8964_8799.n234 a_n8964_8799.n229 161.3
R289 a_n8964_8799.n235 a_n8964_8799.n228 161.3
R290 a_n8964_8799.n237 a_n8964_8799.n236 161.3
R291 a_n8964_8799.n238 a_n8964_8799.n227 161.3
R292 a_n8964_8799.n240 a_n8964_8799.n239 161.3
R293 a_n8964_8799.n241 a_n8964_8799.n226 161.3
R294 a_n8964_8799.n242 a_n8964_8799.n225 161.3
R295 a_n8964_8799.n244 a_n8964_8799.n243 161.3
R296 a_n8964_8799.n245 a_n8964_8799.n224 161.3
R297 a_n8964_8799.n247 a_n8964_8799.n246 161.3
R298 a_n8964_8799.n248 a_n8964_8799.n223 161.3
R299 a_n8964_8799.n249 a_n8964_8799.n222 161.3
R300 a_n8964_8799.n251 a_n8964_8799.n250 161.3
R301 a_n8964_8799.n252 a_n8964_8799.n221 161.3
R302 a_n8964_8799.n254 a_n8964_8799.n253 161.3
R303 a_n8964_8799.n255 a_n8964_8799.n220 161.3
R304 a_n8964_8799.n256 a_n8964_8799.n219 161.3
R305 a_n8964_8799.n258 a_n8964_8799.n257 161.3
R306 a_n8964_8799.n259 a_n8964_8799.n218 161.3
R307 a_n8964_8799.n261 a_n8964_8799.n260 161.3
R308 a_n8964_8799.n262 a_n8964_8799.n217 161.3
R309 a_n8964_8799.n264 a_n8964_8799.n263 161.3
R310 a_n8964_8799.n282 a_n8964_8799.n281 161.3
R311 a_n8964_8799.n283 a_n8964_8799.n278 161.3
R312 a_n8964_8799.n284 a_n8964_8799.n277 161.3
R313 a_n8964_8799.n286 a_n8964_8799.n285 161.3
R314 a_n8964_8799.n287 a_n8964_8799.n276 161.3
R315 a_n8964_8799.n289 a_n8964_8799.n288 161.3
R316 a_n8964_8799.n290 a_n8964_8799.n275 161.3
R317 a_n8964_8799.n291 a_n8964_8799.n274 161.3
R318 a_n8964_8799.n293 a_n8964_8799.n292 161.3
R319 a_n8964_8799.n294 a_n8964_8799.n273 161.3
R320 a_n8964_8799.n296 a_n8964_8799.n295 161.3
R321 a_n8964_8799.n297 a_n8964_8799.n272 161.3
R322 a_n8964_8799.n298 a_n8964_8799.n271 161.3
R323 a_n8964_8799.n300 a_n8964_8799.n299 161.3
R324 a_n8964_8799.n301 a_n8964_8799.n270 161.3
R325 a_n8964_8799.n303 a_n8964_8799.n302 161.3
R326 a_n8964_8799.n304 a_n8964_8799.n269 161.3
R327 a_n8964_8799.n305 a_n8964_8799.n268 161.3
R328 a_n8964_8799.n307 a_n8964_8799.n306 161.3
R329 a_n8964_8799.n308 a_n8964_8799.n267 161.3
R330 a_n8964_8799.n310 a_n8964_8799.n309 161.3
R331 a_n8964_8799.n311 a_n8964_8799.n266 161.3
R332 a_n8964_8799.n313 a_n8964_8799.n312 161.3
R333 a_n8964_8799.n70 a_n8964_8799.n69 161.3
R334 a_n8964_8799.n68 a_n8964_8799.n23 161.3
R335 a_n8964_8799.n67 a_n8964_8799.n66 161.3
R336 a_n8964_8799.n65 a_n8964_8799.n24 161.3
R337 a_n8964_8799.n64 a_n8964_8799.n63 161.3
R338 a_n8964_8799.n62 a_n8964_8799.n25 161.3
R339 a_n8964_8799.n61 a_n8964_8799.n60 161.3
R340 a_n8964_8799.n59 a_n8964_8799.n26 161.3
R341 a_n8964_8799.n58 a_n8964_8799.n57 161.3
R342 a_n8964_8799.n56 a_n8964_8799.n27 161.3
R343 a_n8964_8799.n55 a_n8964_8799.n54 161.3
R344 a_n8964_8799.n53 a_n8964_8799.n28 161.3
R345 a_n8964_8799.n52 a_n8964_8799.n51 161.3
R346 a_n8964_8799.n50 a_n8964_8799.n29 161.3
R347 a_n8964_8799.n49 a_n8964_8799.n48 161.3
R348 a_n8964_8799.n47 a_n8964_8799.n30 161.3
R349 a_n8964_8799.n46 a_n8964_8799.n45 161.3
R350 a_n8964_8799.n44 a_n8964_8799.n31 161.3
R351 a_n8964_8799.n43 a_n8964_8799.n42 161.3
R352 a_n8964_8799.n41 a_n8964_8799.n32 161.3
R353 a_n8964_8799.n40 a_n8964_8799.n39 161.3
R354 a_n8964_8799.n38 a_n8964_8799.n33 161.3
R355 a_n8964_8799.n37 a_n8964_8799.n36 161.3
R356 a_n8964_8799.n118 a_n8964_8799.n117 161.3
R357 a_n8964_8799.n116 a_n8964_8799.n71 161.3
R358 a_n8964_8799.n115 a_n8964_8799.n114 161.3
R359 a_n8964_8799.n113 a_n8964_8799.n72 161.3
R360 a_n8964_8799.n112 a_n8964_8799.n111 161.3
R361 a_n8964_8799.n110 a_n8964_8799.n73 161.3
R362 a_n8964_8799.n109 a_n8964_8799.n108 161.3
R363 a_n8964_8799.n107 a_n8964_8799.n74 161.3
R364 a_n8964_8799.n106 a_n8964_8799.n105 161.3
R365 a_n8964_8799.n104 a_n8964_8799.n75 161.3
R366 a_n8964_8799.n103 a_n8964_8799.n102 161.3
R367 a_n8964_8799.n101 a_n8964_8799.n76 161.3
R368 a_n8964_8799.n100 a_n8964_8799.n99 161.3
R369 a_n8964_8799.n98 a_n8964_8799.n77 161.3
R370 a_n8964_8799.n97 a_n8964_8799.n96 161.3
R371 a_n8964_8799.n95 a_n8964_8799.n78 161.3
R372 a_n8964_8799.n94 a_n8964_8799.n93 161.3
R373 a_n8964_8799.n92 a_n8964_8799.n79 161.3
R374 a_n8964_8799.n91 a_n8964_8799.n90 161.3
R375 a_n8964_8799.n89 a_n8964_8799.n80 161.3
R376 a_n8964_8799.n88 a_n8964_8799.n87 161.3
R377 a_n8964_8799.n86 a_n8964_8799.n81 161.3
R378 a_n8964_8799.n85 a_n8964_8799.n84 161.3
R379 a_n8964_8799.n167 a_n8964_8799.n166 161.3
R380 a_n8964_8799.n165 a_n8964_8799.n120 161.3
R381 a_n8964_8799.n164 a_n8964_8799.n163 161.3
R382 a_n8964_8799.n162 a_n8964_8799.n121 161.3
R383 a_n8964_8799.n161 a_n8964_8799.n160 161.3
R384 a_n8964_8799.n159 a_n8964_8799.n122 161.3
R385 a_n8964_8799.n158 a_n8964_8799.n157 161.3
R386 a_n8964_8799.n156 a_n8964_8799.n123 161.3
R387 a_n8964_8799.n155 a_n8964_8799.n154 161.3
R388 a_n8964_8799.n153 a_n8964_8799.n124 161.3
R389 a_n8964_8799.n152 a_n8964_8799.n151 161.3
R390 a_n8964_8799.n150 a_n8964_8799.n125 161.3
R391 a_n8964_8799.n149 a_n8964_8799.n148 161.3
R392 a_n8964_8799.n147 a_n8964_8799.n126 161.3
R393 a_n8964_8799.n146 a_n8964_8799.n145 161.3
R394 a_n8964_8799.n144 a_n8964_8799.n127 161.3
R395 a_n8964_8799.n143 a_n8964_8799.n142 161.3
R396 a_n8964_8799.n141 a_n8964_8799.n128 161.3
R397 a_n8964_8799.n140 a_n8964_8799.n139 161.3
R398 a_n8964_8799.n138 a_n8964_8799.n129 161.3
R399 a_n8964_8799.n137 a_n8964_8799.n136 161.3
R400 a_n8964_8799.n135 a_n8964_8799.n130 161.3
R401 a_n8964_8799.n134 a_n8964_8799.n133 161.3
R402 a_n8964_8799.n13 a_n8964_8799.n11 98.9633
R403 a_n8964_8799.n2 a_n8964_8799.n0 98.9631
R404 a_n8964_8799.n21 a_n8964_8799.n20 98.6055
R405 a_n8964_8799.n19 a_n8964_8799.n18 98.6055
R406 a_n8964_8799.n17 a_n8964_8799.n16 98.6055
R407 a_n8964_8799.n15 a_n8964_8799.n14 98.6055
R408 a_n8964_8799.n13 a_n8964_8799.n12 98.6055
R409 a_n8964_8799.n2 a_n8964_8799.n1 98.6055
R410 a_n8964_8799.n4 a_n8964_8799.n3 98.6055
R411 a_n8964_8799.n6 a_n8964_8799.n5 98.6055
R412 a_n8964_8799.n8 a_n8964_8799.n7 98.6055
R413 a_n8964_8799.n10 a_n8964_8799.n9 98.6055
R414 a_n8964_8799.n331 a_n8964_8799.n330 81.3766
R415 a_n8964_8799.n319 a_n8964_8799.n317 81.3764
R416 a_n8964_8799.n327 a_n8964_8799.n325 81.3764
R417 a_n8964_8799.n324 a_n8964_8799.n323 80.9324
R418 a_n8964_8799.n322 a_n8964_8799.n321 80.9324
R419 a_n8964_8799.n319 a_n8964_8799.n318 80.9324
R420 a_n8964_8799.n327 a_n8964_8799.n326 80.9324
R421 a_n8964_8799.n330 a_n8964_8799.n329 80.9324
R422 a_n8964_8799.n184 a_n8964_8799.n183 70.4033
R423 a_n8964_8799.n232 a_n8964_8799.n231 70.4033
R424 a_n8964_8799.n281 a_n8964_8799.n280 70.4033
R425 a_n8964_8799.n36 a_n8964_8799.n35 70.4033
R426 a_n8964_8799.n84 a_n8964_8799.n83 70.4033
R427 a_n8964_8799.n133 a_n8964_8799.n132 70.4033
R428 a_n8964_8799.n215 a_n8964_8799.n214 48.2005
R429 a_n8964_8799.n208 a_n8964_8799.n207 48.2005
R430 a_n8964_8799.n201 a_n8964_8799.n200 48.2005
R431 a_n8964_8799.n195 a_n8964_8799.n176 48.2005
R432 a_n8964_8799.n188 a_n8964_8799.n179 48.2005
R433 a_n8964_8799.n263 a_n8964_8799.n262 48.2005
R434 a_n8964_8799.n256 a_n8964_8799.n255 48.2005
R435 a_n8964_8799.n249 a_n8964_8799.n248 48.2005
R436 a_n8964_8799.n243 a_n8964_8799.n224 48.2005
R437 a_n8964_8799.n236 a_n8964_8799.n227 48.2005
R438 a_n8964_8799.n312 a_n8964_8799.n311 48.2005
R439 a_n8964_8799.n305 a_n8964_8799.n304 48.2005
R440 a_n8964_8799.n298 a_n8964_8799.n297 48.2005
R441 a_n8964_8799.n292 a_n8964_8799.n273 48.2005
R442 a_n8964_8799.n285 a_n8964_8799.n276 48.2005
R443 a_n8964_8799.n43 a_n8964_8799.n32 48.2005
R444 a_n8964_8799.n50 a_n8964_8799.n49 48.2005
R445 a_n8964_8799.n55 a_n8964_8799.n28 48.2005
R446 a_n8964_8799.n62 a_n8964_8799.n61 48.2005
R447 a_n8964_8799.n69 a_n8964_8799.n68 48.2005
R448 a_n8964_8799.n91 a_n8964_8799.n80 48.2005
R449 a_n8964_8799.n98 a_n8964_8799.n97 48.2005
R450 a_n8964_8799.n103 a_n8964_8799.n76 48.2005
R451 a_n8964_8799.n110 a_n8964_8799.n109 48.2005
R452 a_n8964_8799.n117 a_n8964_8799.n116 48.2005
R453 a_n8964_8799.n140 a_n8964_8799.n129 48.2005
R454 a_n8964_8799.n147 a_n8964_8799.n146 48.2005
R455 a_n8964_8799.n152 a_n8964_8799.n125 48.2005
R456 a_n8964_8799.n159 a_n8964_8799.n158 48.2005
R457 a_n8964_8799.n166 a_n8964_8799.n165 48.2005
R458 a_n8964_8799.n202 a_n8964_8799.n173 47.4702
R459 a_n8964_8799.n194 a_n8964_8799.n193 47.4702
R460 a_n8964_8799.n250 a_n8964_8799.n221 47.4702
R461 a_n8964_8799.n242 a_n8964_8799.n241 47.4702
R462 a_n8964_8799.n299 a_n8964_8799.n270 47.4702
R463 a_n8964_8799.n291 a_n8964_8799.n290 47.4702
R464 a_n8964_8799.n45 a_n8964_8799.n30 47.4702
R465 a_n8964_8799.n57 a_n8964_8799.n56 47.4702
R466 a_n8964_8799.n93 a_n8964_8799.n78 47.4702
R467 a_n8964_8799.n105 a_n8964_8799.n104 47.4702
R468 a_n8964_8799.n142 a_n8964_8799.n127 47.4702
R469 a_n8964_8799.n154 a_n8964_8799.n153 47.4702
R470 a_n8964_8799.n209 a_n8964_8799.n170 46.0096
R471 a_n8964_8799.n187 a_n8964_8799.n186 46.0096
R472 a_n8964_8799.n257 a_n8964_8799.n218 46.0096
R473 a_n8964_8799.n235 a_n8964_8799.n234 46.0096
R474 a_n8964_8799.n306 a_n8964_8799.n267 46.0096
R475 a_n8964_8799.n284 a_n8964_8799.n283 46.0096
R476 a_n8964_8799.n39 a_n8964_8799.n38 46.0096
R477 a_n8964_8799.n63 a_n8964_8799.n24 46.0096
R478 a_n8964_8799.n87 a_n8964_8799.n86 46.0096
R479 a_n8964_8799.n111 a_n8964_8799.n72 46.0096
R480 a_n8964_8799.n136 a_n8964_8799.n135 46.0096
R481 a_n8964_8799.n160 a_n8964_8799.n121 46.0096
R482 a_n8964_8799.n22 a_n8964_8799.n10 33.7114
R483 a_n8964_8799.n328 a_n8964_8799.n324 32.0866
R484 a_n8964_8799.n213 a_n8964_8799.n170 27.0217
R485 a_n8964_8799.n186 a_n8964_8799.n185 27.0217
R486 a_n8964_8799.n261 a_n8964_8799.n218 27.0217
R487 a_n8964_8799.n234 a_n8964_8799.n233 27.0217
R488 a_n8964_8799.n310 a_n8964_8799.n267 27.0217
R489 a_n8964_8799.n283 a_n8964_8799.n282 27.0217
R490 a_n8964_8799.n38 a_n8964_8799.n37 27.0217
R491 a_n8964_8799.n67 a_n8964_8799.n24 27.0217
R492 a_n8964_8799.n86 a_n8964_8799.n85 27.0217
R493 a_n8964_8799.n115 a_n8964_8799.n72 27.0217
R494 a_n8964_8799.n135 a_n8964_8799.n134 27.0217
R495 a_n8964_8799.n164 a_n8964_8799.n121 27.0217
R496 a_n8964_8799.n206 a_n8964_8799.n173 25.5611
R497 a_n8964_8799.n193 a_n8964_8799.n192 25.5611
R498 a_n8964_8799.n254 a_n8964_8799.n221 25.5611
R499 a_n8964_8799.n241 a_n8964_8799.n240 25.5611
R500 a_n8964_8799.n303 a_n8964_8799.n270 25.5611
R501 a_n8964_8799.n290 a_n8964_8799.n289 25.5611
R502 a_n8964_8799.n45 a_n8964_8799.n44 25.5611
R503 a_n8964_8799.n57 a_n8964_8799.n26 25.5611
R504 a_n8964_8799.n93 a_n8964_8799.n92 25.5611
R505 a_n8964_8799.n105 a_n8964_8799.n74 25.5611
R506 a_n8964_8799.n142 a_n8964_8799.n141 25.5611
R507 a_n8964_8799.n154 a_n8964_8799.n123 25.5611
R508 a_n8964_8799.n200 a_n8964_8799.n199 24.1005
R509 a_n8964_8799.n199 a_n8964_8799.n176 24.1005
R510 a_n8964_8799.n248 a_n8964_8799.n247 24.1005
R511 a_n8964_8799.n247 a_n8964_8799.n224 24.1005
R512 a_n8964_8799.n297 a_n8964_8799.n296 24.1005
R513 a_n8964_8799.n296 a_n8964_8799.n273 24.1005
R514 a_n8964_8799.n51 a_n8964_8799.n50 24.1005
R515 a_n8964_8799.n51 a_n8964_8799.n28 24.1005
R516 a_n8964_8799.n99 a_n8964_8799.n98 24.1005
R517 a_n8964_8799.n99 a_n8964_8799.n76 24.1005
R518 a_n8964_8799.n148 a_n8964_8799.n147 24.1005
R519 a_n8964_8799.n148 a_n8964_8799.n125 24.1005
R520 a_n8964_8799.n207 a_n8964_8799.n206 22.6399
R521 a_n8964_8799.n192 a_n8964_8799.n179 22.6399
R522 a_n8964_8799.n255 a_n8964_8799.n254 22.6399
R523 a_n8964_8799.n240 a_n8964_8799.n227 22.6399
R524 a_n8964_8799.n304 a_n8964_8799.n303 22.6399
R525 a_n8964_8799.n289 a_n8964_8799.n276 22.6399
R526 a_n8964_8799.n44 a_n8964_8799.n43 22.6399
R527 a_n8964_8799.n61 a_n8964_8799.n26 22.6399
R528 a_n8964_8799.n92 a_n8964_8799.n91 22.6399
R529 a_n8964_8799.n109 a_n8964_8799.n74 22.6399
R530 a_n8964_8799.n141 a_n8964_8799.n140 22.6399
R531 a_n8964_8799.n158 a_n8964_8799.n123 22.6399
R532 a_n8964_8799.n214 a_n8964_8799.n213 21.1793
R533 a_n8964_8799.n185 a_n8964_8799.n182 21.1793
R534 a_n8964_8799.n262 a_n8964_8799.n261 21.1793
R535 a_n8964_8799.n233 a_n8964_8799.n230 21.1793
R536 a_n8964_8799.n311 a_n8964_8799.n310 21.1793
R537 a_n8964_8799.n282 a_n8964_8799.n279 21.1793
R538 a_n8964_8799.n37 a_n8964_8799.n34 21.1793
R539 a_n8964_8799.n68 a_n8964_8799.n67 21.1793
R540 a_n8964_8799.n85 a_n8964_8799.n82 21.1793
R541 a_n8964_8799.n116 a_n8964_8799.n115 21.1793
R542 a_n8964_8799.n134 a_n8964_8799.n131 21.1793
R543 a_n8964_8799.n165 a_n8964_8799.n164 21.1793
R544 a_n8964_8799.n22 a_n8964_8799.n21 21.1779
R545 a_n8964_8799.n183 a_n8964_8799.n182 20.9576
R546 a_n8964_8799.n231 a_n8964_8799.n230 20.9576
R547 a_n8964_8799.n280 a_n8964_8799.n279 20.9576
R548 a_n8964_8799.n35 a_n8964_8799.n34 20.9576
R549 a_n8964_8799.n83 a_n8964_8799.n82 20.9576
R550 a_n8964_8799.n132 a_n8964_8799.n131 20.9576
R551 a_n8964_8799.n320 a_n8964_8799.n316 12.3339
R552 a_n8964_8799.n316 a_n8964_8799.n22 11.4887
R553 a_n8964_8799.n265 a_n8964_8799.n216 9.07815
R554 a_n8964_8799.n119 a_n8964_8799.n70 9.07815
R555 a_n8964_8799.n315 a_n8964_8799.n168 7.14965
R556 a_n8964_8799.n315 a_n8964_8799.n314 6.85731
R557 a_n8964_8799.n265 a_n8964_8799.n264 4.9702
R558 a_n8964_8799.n314 a_n8964_8799.n313 4.9702
R559 a_n8964_8799.n119 a_n8964_8799.n118 4.9702
R560 a_n8964_8799.n168 a_n8964_8799.n167 4.9702
R561 a_n8964_8799.n314 a_n8964_8799.n265 4.10845
R562 a_n8964_8799.n168 a_n8964_8799.n119 4.10845
R563 a_n8964_8799.n20 a_n8964_8799.t12 3.61217
R564 a_n8964_8799.n20 a_n8964_8799.t13 3.61217
R565 a_n8964_8799.n18 a_n8964_8799.t5 3.61217
R566 a_n8964_8799.n18 a_n8964_8799.t1 3.61217
R567 a_n8964_8799.n16 a_n8964_8799.t3 3.61217
R568 a_n8964_8799.n16 a_n8964_8799.t18 3.61217
R569 a_n8964_8799.n14 a_n8964_8799.t4 3.61217
R570 a_n8964_8799.n14 a_n8964_8799.t11 3.61217
R571 a_n8964_8799.n12 a_n8964_8799.t6 3.61217
R572 a_n8964_8799.n12 a_n8964_8799.t39 3.61217
R573 a_n8964_8799.n11 a_n8964_8799.t8 3.61217
R574 a_n8964_8799.n11 a_n8964_8799.t38 3.61217
R575 a_n8964_8799.n0 a_n8964_8799.t17 3.61217
R576 a_n8964_8799.n0 a_n8964_8799.t19 3.61217
R577 a_n8964_8799.n1 a_n8964_8799.t0 3.61217
R578 a_n8964_8799.n1 a_n8964_8799.t15 3.61217
R579 a_n8964_8799.n3 a_n8964_8799.t7 3.61217
R580 a_n8964_8799.n3 a_n8964_8799.t2 3.61217
R581 a_n8964_8799.n5 a_n8964_8799.t21 3.61217
R582 a_n8964_8799.n5 a_n8964_8799.t9 3.61217
R583 a_n8964_8799.n7 a_n8964_8799.t14 3.61217
R584 a_n8964_8799.n7 a_n8964_8799.t20 3.61217
R585 a_n8964_8799.n9 a_n8964_8799.t10 3.61217
R586 a_n8964_8799.n9 a_n8964_8799.t16 3.61217
R587 a_n8964_8799.n316 a_n8964_8799.n315 3.4105
R588 a_n8964_8799.n325 a_n8964_8799.t32 2.82907
R589 a_n8964_8799.n325 a_n8964_8799.t30 2.82907
R590 a_n8964_8799.n326 a_n8964_8799.t25 2.82907
R591 a_n8964_8799.n326 a_n8964_8799.t29 2.82907
R592 a_n8964_8799.n329 a_n8964_8799.t36 2.82907
R593 a_n8964_8799.n329 a_n8964_8799.t26 2.82907
R594 a_n8964_8799.n323 a_n8964_8799.t35 2.82907
R595 a_n8964_8799.n323 a_n8964_8799.t31 2.82907
R596 a_n8964_8799.n321 a_n8964_8799.t22 2.82907
R597 a_n8964_8799.n321 a_n8964_8799.t34 2.82907
R598 a_n8964_8799.n318 a_n8964_8799.t23 2.82907
R599 a_n8964_8799.n318 a_n8964_8799.t24 2.82907
R600 a_n8964_8799.n317 a_n8964_8799.t27 2.82907
R601 a_n8964_8799.n317 a_n8964_8799.t28 2.82907
R602 a_n8964_8799.n331 a_n8964_8799.t33 2.82907
R603 a_n8964_8799.t37 a_n8964_8799.n331 2.82907
R604 a_n8964_8799.n209 a_n8964_8799.n208 2.19141
R605 a_n8964_8799.n188 a_n8964_8799.n187 2.19141
R606 a_n8964_8799.n257 a_n8964_8799.n256 2.19141
R607 a_n8964_8799.n236 a_n8964_8799.n235 2.19141
R608 a_n8964_8799.n306 a_n8964_8799.n305 2.19141
R609 a_n8964_8799.n285 a_n8964_8799.n284 2.19141
R610 a_n8964_8799.n39 a_n8964_8799.n32 2.19141
R611 a_n8964_8799.n63 a_n8964_8799.n62 2.19141
R612 a_n8964_8799.n87 a_n8964_8799.n80 2.19141
R613 a_n8964_8799.n111 a_n8964_8799.n110 2.19141
R614 a_n8964_8799.n136 a_n8964_8799.n129 2.19141
R615 a_n8964_8799.n160 a_n8964_8799.n159 2.19141
R616 a_n8964_8799.n202 a_n8964_8799.n201 0.730803
R617 a_n8964_8799.n195 a_n8964_8799.n194 0.730803
R618 a_n8964_8799.n250 a_n8964_8799.n249 0.730803
R619 a_n8964_8799.n243 a_n8964_8799.n242 0.730803
R620 a_n8964_8799.n299 a_n8964_8799.n298 0.730803
R621 a_n8964_8799.n292 a_n8964_8799.n291 0.730803
R622 a_n8964_8799.n49 a_n8964_8799.n30 0.730803
R623 a_n8964_8799.n56 a_n8964_8799.n55 0.730803
R624 a_n8964_8799.n97 a_n8964_8799.n78 0.730803
R625 a_n8964_8799.n104 a_n8964_8799.n103 0.730803
R626 a_n8964_8799.n146 a_n8964_8799.n127 0.730803
R627 a_n8964_8799.n153 a_n8964_8799.n152 0.730803
R628 a_n8964_8799.n324 a_n8964_8799.n322 0.444466
R629 a_n8964_8799.n15 a_n8964_8799.n13 0.358259
R630 a_n8964_8799.n17 a_n8964_8799.n15 0.358259
R631 a_n8964_8799.n19 a_n8964_8799.n17 0.358259
R632 a_n8964_8799.n21 a_n8964_8799.n19 0.358259
R633 a_n8964_8799.n10 a_n8964_8799.n8 0.358259
R634 a_n8964_8799.n8 a_n8964_8799.n6 0.358259
R635 a_n8964_8799.n6 a_n8964_8799.n4 0.358259
R636 a_n8964_8799.n4 a_n8964_8799.n2 0.358259
R637 a_n8964_8799.n320 a_n8964_8799.n319 0.222483
R638 a_n8964_8799.n322 a_n8964_8799.n320 0.222483
R639 a_n8964_8799.n330 a_n8964_8799.n328 0.222483
R640 a_n8964_8799.n328 a_n8964_8799.n327 0.222483
R641 a_n8964_8799.n216 a_n8964_8799.n169 0.189894
R642 a_n8964_8799.n212 a_n8964_8799.n169 0.189894
R643 a_n8964_8799.n212 a_n8964_8799.n211 0.189894
R644 a_n8964_8799.n211 a_n8964_8799.n210 0.189894
R645 a_n8964_8799.n210 a_n8964_8799.n171 0.189894
R646 a_n8964_8799.n172 a_n8964_8799.n171 0.189894
R647 a_n8964_8799.n205 a_n8964_8799.n172 0.189894
R648 a_n8964_8799.n205 a_n8964_8799.n204 0.189894
R649 a_n8964_8799.n204 a_n8964_8799.n203 0.189894
R650 a_n8964_8799.n203 a_n8964_8799.n174 0.189894
R651 a_n8964_8799.n175 a_n8964_8799.n174 0.189894
R652 a_n8964_8799.n198 a_n8964_8799.n175 0.189894
R653 a_n8964_8799.n198 a_n8964_8799.n197 0.189894
R654 a_n8964_8799.n197 a_n8964_8799.n196 0.189894
R655 a_n8964_8799.n196 a_n8964_8799.n177 0.189894
R656 a_n8964_8799.n178 a_n8964_8799.n177 0.189894
R657 a_n8964_8799.n191 a_n8964_8799.n178 0.189894
R658 a_n8964_8799.n191 a_n8964_8799.n190 0.189894
R659 a_n8964_8799.n190 a_n8964_8799.n189 0.189894
R660 a_n8964_8799.n189 a_n8964_8799.n180 0.189894
R661 a_n8964_8799.n181 a_n8964_8799.n180 0.189894
R662 a_n8964_8799.n184 a_n8964_8799.n181 0.189894
R663 a_n8964_8799.n264 a_n8964_8799.n217 0.189894
R664 a_n8964_8799.n260 a_n8964_8799.n217 0.189894
R665 a_n8964_8799.n260 a_n8964_8799.n259 0.189894
R666 a_n8964_8799.n259 a_n8964_8799.n258 0.189894
R667 a_n8964_8799.n258 a_n8964_8799.n219 0.189894
R668 a_n8964_8799.n220 a_n8964_8799.n219 0.189894
R669 a_n8964_8799.n253 a_n8964_8799.n220 0.189894
R670 a_n8964_8799.n253 a_n8964_8799.n252 0.189894
R671 a_n8964_8799.n252 a_n8964_8799.n251 0.189894
R672 a_n8964_8799.n251 a_n8964_8799.n222 0.189894
R673 a_n8964_8799.n223 a_n8964_8799.n222 0.189894
R674 a_n8964_8799.n246 a_n8964_8799.n223 0.189894
R675 a_n8964_8799.n246 a_n8964_8799.n245 0.189894
R676 a_n8964_8799.n245 a_n8964_8799.n244 0.189894
R677 a_n8964_8799.n244 a_n8964_8799.n225 0.189894
R678 a_n8964_8799.n226 a_n8964_8799.n225 0.189894
R679 a_n8964_8799.n239 a_n8964_8799.n226 0.189894
R680 a_n8964_8799.n239 a_n8964_8799.n238 0.189894
R681 a_n8964_8799.n238 a_n8964_8799.n237 0.189894
R682 a_n8964_8799.n237 a_n8964_8799.n228 0.189894
R683 a_n8964_8799.n229 a_n8964_8799.n228 0.189894
R684 a_n8964_8799.n232 a_n8964_8799.n229 0.189894
R685 a_n8964_8799.n313 a_n8964_8799.n266 0.189894
R686 a_n8964_8799.n309 a_n8964_8799.n266 0.189894
R687 a_n8964_8799.n309 a_n8964_8799.n308 0.189894
R688 a_n8964_8799.n308 a_n8964_8799.n307 0.189894
R689 a_n8964_8799.n307 a_n8964_8799.n268 0.189894
R690 a_n8964_8799.n269 a_n8964_8799.n268 0.189894
R691 a_n8964_8799.n302 a_n8964_8799.n269 0.189894
R692 a_n8964_8799.n302 a_n8964_8799.n301 0.189894
R693 a_n8964_8799.n301 a_n8964_8799.n300 0.189894
R694 a_n8964_8799.n300 a_n8964_8799.n271 0.189894
R695 a_n8964_8799.n272 a_n8964_8799.n271 0.189894
R696 a_n8964_8799.n295 a_n8964_8799.n272 0.189894
R697 a_n8964_8799.n295 a_n8964_8799.n294 0.189894
R698 a_n8964_8799.n294 a_n8964_8799.n293 0.189894
R699 a_n8964_8799.n293 a_n8964_8799.n274 0.189894
R700 a_n8964_8799.n275 a_n8964_8799.n274 0.189894
R701 a_n8964_8799.n288 a_n8964_8799.n275 0.189894
R702 a_n8964_8799.n288 a_n8964_8799.n287 0.189894
R703 a_n8964_8799.n287 a_n8964_8799.n286 0.189894
R704 a_n8964_8799.n286 a_n8964_8799.n277 0.189894
R705 a_n8964_8799.n278 a_n8964_8799.n277 0.189894
R706 a_n8964_8799.n281 a_n8964_8799.n278 0.189894
R707 a_n8964_8799.n36 a_n8964_8799.n33 0.189894
R708 a_n8964_8799.n40 a_n8964_8799.n33 0.189894
R709 a_n8964_8799.n41 a_n8964_8799.n40 0.189894
R710 a_n8964_8799.n42 a_n8964_8799.n41 0.189894
R711 a_n8964_8799.n42 a_n8964_8799.n31 0.189894
R712 a_n8964_8799.n46 a_n8964_8799.n31 0.189894
R713 a_n8964_8799.n47 a_n8964_8799.n46 0.189894
R714 a_n8964_8799.n48 a_n8964_8799.n47 0.189894
R715 a_n8964_8799.n48 a_n8964_8799.n29 0.189894
R716 a_n8964_8799.n52 a_n8964_8799.n29 0.189894
R717 a_n8964_8799.n53 a_n8964_8799.n52 0.189894
R718 a_n8964_8799.n54 a_n8964_8799.n53 0.189894
R719 a_n8964_8799.n54 a_n8964_8799.n27 0.189894
R720 a_n8964_8799.n58 a_n8964_8799.n27 0.189894
R721 a_n8964_8799.n59 a_n8964_8799.n58 0.189894
R722 a_n8964_8799.n60 a_n8964_8799.n59 0.189894
R723 a_n8964_8799.n60 a_n8964_8799.n25 0.189894
R724 a_n8964_8799.n64 a_n8964_8799.n25 0.189894
R725 a_n8964_8799.n65 a_n8964_8799.n64 0.189894
R726 a_n8964_8799.n66 a_n8964_8799.n65 0.189894
R727 a_n8964_8799.n66 a_n8964_8799.n23 0.189894
R728 a_n8964_8799.n70 a_n8964_8799.n23 0.189894
R729 a_n8964_8799.n84 a_n8964_8799.n81 0.189894
R730 a_n8964_8799.n88 a_n8964_8799.n81 0.189894
R731 a_n8964_8799.n89 a_n8964_8799.n88 0.189894
R732 a_n8964_8799.n90 a_n8964_8799.n89 0.189894
R733 a_n8964_8799.n90 a_n8964_8799.n79 0.189894
R734 a_n8964_8799.n94 a_n8964_8799.n79 0.189894
R735 a_n8964_8799.n95 a_n8964_8799.n94 0.189894
R736 a_n8964_8799.n96 a_n8964_8799.n95 0.189894
R737 a_n8964_8799.n96 a_n8964_8799.n77 0.189894
R738 a_n8964_8799.n100 a_n8964_8799.n77 0.189894
R739 a_n8964_8799.n101 a_n8964_8799.n100 0.189894
R740 a_n8964_8799.n102 a_n8964_8799.n101 0.189894
R741 a_n8964_8799.n102 a_n8964_8799.n75 0.189894
R742 a_n8964_8799.n106 a_n8964_8799.n75 0.189894
R743 a_n8964_8799.n107 a_n8964_8799.n106 0.189894
R744 a_n8964_8799.n108 a_n8964_8799.n107 0.189894
R745 a_n8964_8799.n108 a_n8964_8799.n73 0.189894
R746 a_n8964_8799.n112 a_n8964_8799.n73 0.189894
R747 a_n8964_8799.n113 a_n8964_8799.n112 0.189894
R748 a_n8964_8799.n114 a_n8964_8799.n113 0.189894
R749 a_n8964_8799.n114 a_n8964_8799.n71 0.189894
R750 a_n8964_8799.n118 a_n8964_8799.n71 0.189894
R751 a_n8964_8799.n133 a_n8964_8799.n130 0.189894
R752 a_n8964_8799.n137 a_n8964_8799.n130 0.189894
R753 a_n8964_8799.n138 a_n8964_8799.n137 0.189894
R754 a_n8964_8799.n139 a_n8964_8799.n138 0.189894
R755 a_n8964_8799.n139 a_n8964_8799.n128 0.189894
R756 a_n8964_8799.n143 a_n8964_8799.n128 0.189894
R757 a_n8964_8799.n144 a_n8964_8799.n143 0.189894
R758 a_n8964_8799.n145 a_n8964_8799.n144 0.189894
R759 a_n8964_8799.n145 a_n8964_8799.n126 0.189894
R760 a_n8964_8799.n149 a_n8964_8799.n126 0.189894
R761 a_n8964_8799.n150 a_n8964_8799.n149 0.189894
R762 a_n8964_8799.n151 a_n8964_8799.n150 0.189894
R763 a_n8964_8799.n151 a_n8964_8799.n124 0.189894
R764 a_n8964_8799.n155 a_n8964_8799.n124 0.189894
R765 a_n8964_8799.n156 a_n8964_8799.n155 0.189894
R766 a_n8964_8799.n157 a_n8964_8799.n156 0.189894
R767 a_n8964_8799.n157 a_n8964_8799.n122 0.189894
R768 a_n8964_8799.n161 a_n8964_8799.n122 0.189894
R769 a_n8964_8799.n162 a_n8964_8799.n161 0.189894
R770 a_n8964_8799.n163 a_n8964_8799.n162 0.189894
R771 a_n8964_8799.n163 a_n8964_8799.n120 0.189894
R772 a_n8964_8799.n167 a_n8964_8799.n120 0.189894
R773 gnd.n7376 gnd.n493 1564.47
R774 gnd.n6672 gnd.n6625 939.716
R775 gnd.n4522 gnd.n4521 771.183
R776 gnd.n6094 gnd.n2998 771.183
R777 gnd.n4782 gnd.n3907 771.183
R778 gnd.n6096 gnd.n2993 771.183
R779 gnd.n6687 gnd.n1006 766.379
R780 gnd.n2354 gnd.n1003 766.379
R781 gnd.n1625 gnd.n1528 766.379
R782 gnd.n1621 gnd.n1526 766.379
R783 gnd.n6671 gnd.n1000 756.769
R784 gnd.n6682 gnd.n6681 756.769
R785 gnd.n1718 gnd.n1435 756.769
R786 gnd.n1716 gnd.n1438 756.769
R787 gnd.n257 gnd.n246 751.963
R788 gnd.n7675 gnd.n7674 751.963
R789 gnd.n3174 gnd.n3062 751.963
R790 gnd.n5905 gnd.n3176 751.963
R791 gnd.n2766 gnd.n2754 751.963
R792 gnd.n4767 gnd.n3936 751.963
R793 gnd.n4136 gnd.n2393 751.963
R794 gnd.n4092 gnd.n4091 751.963
R795 gnd.n6884 gnd.n785 703.915
R796 gnd.n7375 gnd.n494 703.915
R797 gnd.n7589 gnd.n7587 703.915
R798 gnd.n4202 gnd.n4195 703.915
R799 gnd.n7854 gnd.n250 696.707
R800 gnd.n7730 gnd.n7729 696.707
R801 gnd.n5908 gnd.n5907 696.707
R802 gnd.n6025 gnd.n3108 696.707
R803 gnd.n6325 gnd.n2759 696.707
R804 gnd.n4751 gnd.n3935 696.707
R805 gnd.n6503 gnd.n2466 696.707
R806 gnd.n6623 gnd.n2397 696.707
R807 gnd.n6884 gnd.n6883 585
R808 gnd.n6885 gnd.n6884 585
R809 gnd.n6882 gnd.n787 585
R810 gnd.n787 gnd.n786 585
R811 gnd.n6881 gnd.n6880 585
R812 gnd.n6880 gnd.n6879 585
R813 gnd.n792 gnd.n791 585
R814 gnd.n6878 gnd.n792 585
R815 gnd.n6876 gnd.n6875 585
R816 gnd.n6877 gnd.n6876 585
R817 gnd.n6874 gnd.n794 585
R818 gnd.n794 gnd.n793 585
R819 gnd.n6873 gnd.n6872 585
R820 gnd.n6872 gnd.n6871 585
R821 gnd.n800 gnd.n799 585
R822 gnd.n6870 gnd.n800 585
R823 gnd.n6868 gnd.n6867 585
R824 gnd.n6869 gnd.n6868 585
R825 gnd.n6866 gnd.n802 585
R826 gnd.n802 gnd.n801 585
R827 gnd.n6865 gnd.n6864 585
R828 gnd.n6864 gnd.n6863 585
R829 gnd.n808 gnd.n807 585
R830 gnd.n6862 gnd.n808 585
R831 gnd.n6860 gnd.n6859 585
R832 gnd.n6861 gnd.n6860 585
R833 gnd.n6858 gnd.n810 585
R834 gnd.n810 gnd.n809 585
R835 gnd.n6857 gnd.n6856 585
R836 gnd.n6856 gnd.n6855 585
R837 gnd.n816 gnd.n815 585
R838 gnd.n6854 gnd.n816 585
R839 gnd.n6852 gnd.n6851 585
R840 gnd.n6853 gnd.n6852 585
R841 gnd.n6850 gnd.n818 585
R842 gnd.n818 gnd.n817 585
R843 gnd.n6849 gnd.n6848 585
R844 gnd.n6848 gnd.n6847 585
R845 gnd.n824 gnd.n823 585
R846 gnd.n6846 gnd.n824 585
R847 gnd.n6844 gnd.n6843 585
R848 gnd.n6845 gnd.n6844 585
R849 gnd.n6842 gnd.n826 585
R850 gnd.n826 gnd.n825 585
R851 gnd.n6841 gnd.n6840 585
R852 gnd.n6840 gnd.n6839 585
R853 gnd.n832 gnd.n831 585
R854 gnd.n6838 gnd.n832 585
R855 gnd.n6836 gnd.n6835 585
R856 gnd.n6837 gnd.n6836 585
R857 gnd.n6834 gnd.n834 585
R858 gnd.n834 gnd.n833 585
R859 gnd.n6833 gnd.n6832 585
R860 gnd.n6832 gnd.n6831 585
R861 gnd.n840 gnd.n839 585
R862 gnd.n6830 gnd.n840 585
R863 gnd.n6828 gnd.n6827 585
R864 gnd.n6829 gnd.n6828 585
R865 gnd.n6826 gnd.n842 585
R866 gnd.n842 gnd.n841 585
R867 gnd.n6825 gnd.n6824 585
R868 gnd.n6824 gnd.n6823 585
R869 gnd.n848 gnd.n847 585
R870 gnd.n6822 gnd.n848 585
R871 gnd.n6820 gnd.n6819 585
R872 gnd.n6821 gnd.n6820 585
R873 gnd.n6818 gnd.n850 585
R874 gnd.n850 gnd.n849 585
R875 gnd.n6817 gnd.n6816 585
R876 gnd.n6816 gnd.n6815 585
R877 gnd.n856 gnd.n855 585
R878 gnd.n6814 gnd.n856 585
R879 gnd.n6812 gnd.n6811 585
R880 gnd.n6813 gnd.n6812 585
R881 gnd.n6810 gnd.n858 585
R882 gnd.n858 gnd.n857 585
R883 gnd.n6809 gnd.n6808 585
R884 gnd.n6808 gnd.n6807 585
R885 gnd.n864 gnd.n863 585
R886 gnd.n6806 gnd.n864 585
R887 gnd.n6804 gnd.n6803 585
R888 gnd.n6805 gnd.n6804 585
R889 gnd.n6802 gnd.n866 585
R890 gnd.n866 gnd.n865 585
R891 gnd.n6801 gnd.n6800 585
R892 gnd.n6800 gnd.n6799 585
R893 gnd.n872 gnd.n871 585
R894 gnd.n6798 gnd.n872 585
R895 gnd.n6796 gnd.n6795 585
R896 gnd.n6797 gnd.n6796 585
R897 gnd.n6794 gnd.n874 585
R898 gnd.n874 gnd.n873 585
R899 gnd.n6793 gnd.n6792 585
R900 gnd.n6792 gnd.n6791 585
R901 gnd.n880 gnd.n879 585
R902 gnd.n6790 gnd.n880 585
R903 gnd.n6788 gnd.n6787 585
R904 gnd.n6789 gnd.n6788 585
R905 gnd.n6786 gnd.n882 585
R906 gnd.n882 gnd.n881 585
R907 gnd.n6785 gnd.n6784 585
R908 gnd.n6784 gnd.n6783 585
R909 gnd.n888 gnd.n887 585
R910 gnd.n6782 gnd.n888 585
R911 gnd.n6780 gnd.n6779 585
R912 gnd.n6781 gnd.n6780 585
R913 gnd.n6778 gnd.n890 585
R914 gnd.n890 gnd.n889 585
R915 gnd.n6777 gnd.n6776 585
R916 gnd.n6776 gnd.n6775 585
R917 gnd.n896 gnd.n895 585
R918 gnd.n6774 gnd.n896 585
R919 gnd.n6772 gnd.n6771 585
R920 gnd.n6773 gnd.n6772 585
R921 gnd.n6770 gnd.n898 585
R922 gnd.n898 gnd.n897 585
R923 gnd.n6769 gnd.n6768 585
R924 gnd.n6768 gnd.n6767 585
R925 gnd.n904 gnd.n903 585
R926 gnd.n6766 gnd.n904 585
R927 gnd.n6764 gnd.n6763 585
R928 gnd.n6765 gnd.n6764 585
R929 gnd.n6762 gnd.n906 585
R930 gnd.n906 gnd.n905 585
R931 gnd.n6761 gnd.n6760 585
R932 gnd.n6760 gnd.n6759 585
R933 gnd.n912 gnd.n911 585
R934 gnd.n6758 gnd.n912 585
R935 gnd.n6756 gnd.n6755 585
R936 gnd.n6757 gnd.n6756 585
R937 gnd.n6754 gnd.n914 585
R938 gnd.n914 gnd.n913 585
R939 gnd.n6753 gnd.n6752 585
R940 gnd.n6752 gnd.n6751 585
R941 gnd.n920 gnd.n919 585
R942 gnd.n6750 gnd.n920 585
R943 gnd.n6748 gnd.n6747 585
R944 gnd.n6749 gnd.n6748 585
R945 gnd.n6746 gnd.n922 585
R946 gnd.n922 gnd.n921 585
R947 gnd.n6745 gnd.n6744 585
R948 gnd.n6744 gnd.n6743 585
R949 gnd.n928 gnd.n927 585
R950 gnd.n6742 gnd.n928 585
R951 gnd.n6740 gnd.n6739 585
R952 gnd.n6741 gnd.n6740 585
R953 gnd.n6738 gnd.n930 585
R954 gnd.n930 gnd.n929 585
R955 gnd.n6737 gnd.n6736 585
R956 gnd.n6736 gnd.n6735 585
R957 gnd.n936 gnd.n935 585
R958 gnd.n6734 gnd.n936 585
R959 gnd.n6732 gnd.n6731 585
R960 gnd.n6733 gnd.n6732 585
R961 gnd.n6730 gnd.n938 585
R962 gnd.n938 gnd.n937 585
R963 gnd.n6729 gnd.n6728 585
R964 gnd.n6728 gnd.n6727 585
R965 gnd.n944 gnd.n943 585
R966 gnd.n6726 gnd.n944 585
R967 gnd.n6724 gnd.n6723 585
R968 gnd.n6725 gnd.n6724 585
R969 gnd.n6722 gnd.n946 585
R970 gnd.n946 gnd.n945 585
R971 gnd.n6721 gnd.n6720 585
R972 gnd.n6720 gnd.n6719 585
R973 gnd.n952 gnd.n951 585
R974 gnd.n6718 gnd.n952 585
R975 gnd.n785 gnd.n784 585
R976 gnd.n6886 gnd.n785 585
R977 gnd.n6889 gnd.n6888 585
R978 gnd.n6888 gnd.n6887 585
R979 gnd.n782 gnd.n781 585
R980 gnd.n781 gnd.n780 585
R981 gnd.n6894 gnd.n6893 585
R982 gnd.n6895 gnd.n6894 585
R983 gnd.n779 gnd.n778 585
R984 gnd.n6896 gnd.n779 585
R985 gnd.n6899 gnd.n6898 585
R986 gnd.n6898 gnd.n6897 585
R987 gnd.n776 gnd.n775 585
R988 gnd.n775 gnd.n774 585
R989 gnd.n6904 gnd.n6903 585
R990 gnd.n6905 gnd.n6904 585
R991 gnd.n773 gnd.n772 585
R992 gnd.n6906 gnd.n773 585
R993 gnd.n6909 gnd.n6908 585
R994 gnd.n6908 gnd.n6907 585
R995 gnd.n770 gnd.n769 585
R996 gnd.n769 gnd.n768 585
R997 gnd.n6914 gnd.n6913 585
R998 gnd.n6915 gnd.n6914 585
R999 gnd.n767 gnd.n766 585
R1000 gnd.n6916 gnd.n767 585
R1001 gnd.n6919 gnd.n6918 585
R1002 gnd.n6918 gnd.n6917 585
R1003 gnd.n764 gnd.n763 585
R1004 gnd.n763 gnd.n762 585
R1005 gnd.n6924 gnd.n6923 585
R1006 gnd.n6925 gnd.n6924 585
R1007 gnd.n761 gnd.n760 585
R1008 gnd.n6926 gnd.n761 585
R1009 gnd.n6929 gnd.n6928 585
R1010 gnd.n6928 gnd.n6927 585
R1011 gnd.n758 gnd.n757 585
R1012 gnd.n757 gnd.n756 585
R1013 gnd.n6934 gnd.n6933 585
R1014 gnd.n6935 gnd.n6934 585
R1015 gnd.n755 gnd.n754 585
R1016 gnd.n6936 gnd.n755 585
R1017 gnd.n6939 gnd.n6938 585
R1018 gnd.n6938 gnd.n6937 585
R1019 gnd.n752 gnd.n751 585
R1020 gnd.n751 gnd.n750 585
R1021 gnd.n6944 gnd.n6943 585
R1022 gnd.n6945 gnd.n6944 585
R1023 gnd.n749 gnd.n748 585
R1024 gnd.n6946 gnd.n749 585
R1025 gnd.n6949 gnd.n6948 585
R1026 gnd.n6948 gnd.n6947 585
R1027 gnd.n746 gnd.n745 585
R1028 gnd.n745 gnd.n744 585
R1029 gnd.n6954 gnd.n6953 585
R1030 gnd.n6955 gnd.n6954 585
R1031 gnd.n743 gnd.n742 585
R1032 gnd.n6956 gnd.n743 585
R1033 gnd.n6959 gnd.n6958 585
R1034 gnd.n6958 gnd.n6957 585
R1035 gnd.n740 gnd.n739 585
R1036 gnd.n739 gnd.n738 585
R1037 gnd.n6964 gnd.n6963 585
R1038 gnd.n6965 gnd.n6964 585
R1039 gnd.n737 gnd.n736 585
R1040 gnd.n6966 gnd.n737 585
R1041 gnd.n6969 gnd.n6968 585
R1042 gnd.n6968 gnd.n6967 585
R1043 gnd.n734 gnd.n733 585
R1044 gnd.n733 gnd.n732 585
R1045 gnd.n6974 gnd.n6973 585
R1046 gnd.n6975 gnd.n6974 585
R1047 gnd.n731 gnd.n730 585
R1048 gnd.n6976 gnd.n731 585
R1049 gnd.n6979 gnd.n6978 585
R1050 gnd.n6978 gnd.n6977 585
R1051 gnd.n728 gnd.n727 585
R1052 gnd.n727 gnd.n726 585
R1053 gnd.n6984 gnd.n6983 585
R1054 gnd.n6985 gnd.n6984 585
R1055 gnd.n725 gnd.n724 585
R1056 gnd.n6986 gnd.n725 585
R1057 gnd.n6989 gnd.n6988 585
R1058 gnd.n6988 gnd.n6987 585
R1059 gnd.n722 gnd.n721 585
R1060 gnd.n721 gnd.n720 585
R1061 gnd.n6994 gnd.n6993 585
R1062 gnd.n6995 gnd.n6994 585
R1063 gnd.n719 gnd.n718 585
R1064 gnd.n6996 gnd.n719 585
R1065 gnd.n6999 gnd.n6998 585
R1066 gnd.n6998 gnd.n6997 585
R1067 gnd.n716 gnd.n715 585
R1068 gnd.n715 gnd.n714 585
R1069 gnd.n7004 gnd.n7003 585
R1070 gnd.n7005 gnd.n7004 585
R1071 gnd.n713 gnd.n712 585
R1072 gnd.n7006 gnd.n713 585
R1073 gnd.n7009 gnd.n7008 585
R1074 gnd.n7008 gnd.n7007 585
R1075 gnd.n710 gnd.n709 585
R1076 gnd.n709 gnd.n708 585
R1077 gnd.n7014 gnd.n7013 585
R1078 gnd.n7015 gnd.n7014 585
R1079 gnd.n707 gnd.n706 585
R1080 gnd.n7016 gnd.n707 585
R1081 gnd.n7019 gnd.n7018 585
R1082 gnd.n7018 gnd.n7017 585
R1083 gnd.n704 gnd.n703 585
R1084 gnd.n703 gnd.n702 585
R1085 gnd.n7024 gnd.n7023 585
R1086 gnd.n7025 gnd.n7024 585
R1087 gnd.n701 gnd.n700 585
R1088 gnd.n7026 gnd.n701 585
R1089 gnd.n7029 gnd.n7028 585
R1090 gnd.n7028 gnd.n7027 585
R1091 gnd.n698 gnd.n697 585
R1092 gnd.n697 gnd.n696 585
R1093 gnd.n7034 gnd.n7033 585
R1094 gnd.n7035 gnd.n7034 585
R1095 gnd.n695 gnd.n694 585
R1096 gnd.n7036 gnd.n695 585
R1097 gnd.n7039 gnd.n7038 585
R1098 gnd.n7038 gnd.n7037 585
R1099 gnd.n692 gnd.n691 585
R1100 gnd.n691 gnd.n690 585
R1101 gnd.n7044 gnd.n7043 585
R1102 gnd.n7045 gnd.n7044 585
R1103 gnd.n689 gnd.n688 585
R1104 gnd.n7046 gnd.n689 585
R1105 gnd.n7049 gnd.n7048 585
R1106 gnd.n7048 gnd.n7047 585
R1107 gnd.n686 gnd.n685 585
R1108 gnd.n685 gnd.n684 585
R1109 gnd.n7054 gnd.n7053 585
R1110 gnd.n7055 gnd.n7054 585
R1111 gnd.n683 gnd.n682 585
R1112 gnd.n7056 gnd.n683 585
R1113 gnd.n7059 gnd.n7058 585
R1114 gnd.n7058 gnd.n7057 585
R1115 gnd.n680 gnd.n679 585
R1116 gnd.n679 gnd.n678 585
R1117 gnd.n7064 gnd.n7063 585
R1118 gnd.n7065 gnd.n7064 585
R1119 gnd.n677 gnd.n676 585
R1120 gnd.n7066 gnd.n677 585
R1121 gnd.n7069 gnd.n7068 585
R1122 gnd.n7068 gnd.n7067 585
R1123 gnd.n674 gnd.n673 585
R1124 gnd.n673 gnd.n672 585
R1125 gnd.n7074 gnd.n7073 585
R1126 gnd.n7075 gnd.n7074 585
R1127 gnd.n671 gnd.n670 585
R1128 gnd.n7076 gnd.n671 585
R1129 gnd.n7079 gnd.n7078 585
R1130 gnd.n7078 gnd.n7077 585
R1131 gnd.n668 gnd.n667 585
R1132 gnd.n667 gnd.n666 585
R1133 gnd.n7084 gnd.n7083 585
R1134 gnd.n7085 gnd.n7084 585
R1135 gnd.n665 gnd.n664 585
R1136 gnd.n7086 gnd.n665 585
R1137 gnd.n7089 gnd.n7088 585
R1138 gnd.n7088 gnd.n7087 585
R1139 gnd.n662 gnd.n661 585
R1140 gnd.n661 gnd.n660 585
R1141 gnd.n7094 gnd.n7093 585
R1142 gnd.n7095 gnd.n7094 585
R1143 gnd.n659 gnd.n658 585
R1144 gnd.n7096 gnd.n659 585
R1145 gnd.n7099 gnd.n7098 585
R1146 gnd.n7098 gnd.n7097 585
R1147 gnd.n656 gnd.n655 585
R1148 gnd.n655 gnd.n654 585
R1149 gnd.n7104 gnd.n7103 585
R1150 gnd.n7105 gnd.n7104 585
R1151 gnd.n653 gnd.n652 585
R1152 gnd.n7106 gnd.n653 585
R1153 gnd.n7109 gnd.n7108 585
R1154 gnd.n7108 gnd.n7107 585
R1155 gnd.n650 gnd.n649 585
R1156 gnd.n649 gnd.n648 585
R1157 gnd.n7114 gnd.n7113 585
R1158 gnd.n7115 gnd.n7114 585
R1159 gnd.n647 gnd.n646 585
R1160 gnd.n7116 gnd.n647 585
R1161 gnd.n7119 gnd.n7118 585
R1162 gnd.n7118 gnd.n7117 585
R1163 gnd.n644 gnd.n643 585
R1164 gnd.n643 gnd.n642 585
R1165 gnd.n7124 gnd.n7123 585
R1166 gnd.n7125 gnd.n7124 585
R1167 gnd.n641 gnd.n640 585
R1168 gnd.n7126 gnd.n641 585
R1169 gnd.n7129 gnd.n7128 585
R1170 gnd.n7128 gnd.n7127 585
R1171 gnd.n638 gnd.n637 585
R1172 gnd.n637 gnd.n636 585
R1173 gnd.n7134 gnd.n7133 585
R1174 gnd.n7135 gnd.n7134 585
R1175 gnd.n635 gnd.n634 585
R1176 gnd.n7136 gnd.n635 585
R1177 gnd.n7139 gnd.n7138 585
R1178 gnd.n7138 gnd.n7137 585
R1179 gnd.n632 gnd.n631 585
R1180 gnd.n631 gnd.n630 585
R1181 gnd.n7144 gnd.n7143 585
R1182 gnd.n7145 gnd.n7144 585
R1183 gnd.n629 gnd.n628 585
R1184 gnd.n7146 gnd.n629 585
R1185 gnd.n7149 gnd.n7148 585
R1186 gnd.n7148 gnd.n7147 585
R1187 gnd.n626 gnd.n625 585
R1188 gnd.n625 gnd.n624 585
R1189 gnd.n7154 gnd.n7153 585
R1190 gnd.n7155 gnd.n7154 585
R1191 gnd.n623 gnd.n622 585
R1192 gnd.n7156 gnd.n623 585
R1193 gnd.n7159 gnd.n7158 585
R1194 gnd.n7158 gnd.n7157 585
R1195 gnd.n620 gnd.n619 585
R1196 gnd.n619 gnd.n618 585
R1197 gnd.n7164 gnd.n7163 585
R1198 gnd.n7165 gnd.n7164 585
R1199 gnd.n617 gnd.n616 585
R1200 gnd.n7166 gnd.n617 585
R1201 gnd.n7169 gnd.n7168 585
R1202 gnd.n7168 gnd.n7167 585
R1203 gnd.n614 gnd.n613 585
R1204 gnd.n613 gnd.n612 585
R1205 gnd.n7174 gnd.n7173 585
R1206 gnd.n7175 gnd.n7174 585
R1207 gnd.n611 gnd.n610 585
R1208 gnd.n7176 gnd.n611 585
R1209 gnd.n7179 gnd.n7178 585
R1210 gnd.n7178 gnd.n7177 585
R1211 gnd.n608 gnd.n607 585
R1212 gnd.n607 gnd.n606 585
R1213 gnd.n7184 gnd.n7183 585
R1214 gnd.n7185 gnd.n7184 585
R1215 gnd.n605 gnd.n604 585
R1216 gnd.n7186 gnd.n605 585
R1217 gnd.n7189 gnd.n7188 585
R1218 gnd.n7188 gnd.n7187 585
R1219 gnd.n602 gnd.n601 585
R1220 gnd.n601 gnd.n600 585
R1221 gnd.n7194 gnd.n7193 585
R1222 gnd.n7195 gnd.n7194 585
R1223 gnd.n599 gnd.n598 585
R1224 gnd.n7196 gnd.n599 585
R1225 gnd.n7199 gnd.n7198 585
R1226 gnd.n7198 gnd.n7197 585
R1227 gnd.n596 gnd.n595 585
R1228 gnd.n595 gnd.n594 585
R1229 gnd.n7204 gnd.n7203 585
R1230 gnd.n7205 gnd.n7204 585
R1231 gnd.n593 gnd.n592 585
R1232 gnd.n7206 gnd.n593 585
R1233 gnd.n7209 gnd.n7208 585
R1234 gnd.n7208 gnd.n7207 585
R1235 gnd.n590 gnd.n589 585
R1236 gnd.n589 gnd.n588 585
R1237 gnd.n7214 gnd.n7213 585
R1238 gnd.n7215 gnd.n7214 585
R1239 gnd.n587 gnd.n586 585
R1240 gnd.n7216 gnd.n587 585
R1241 gnd.n7219 gnd.n7218 585
R1242 gnd.n7218 gnd.n7217 585
R1243 gnd.n584 gnd.n583 585
R1244 gnd.n583 gnd.n582 585
R1245 gnd.n7224 gnd.n7223 585
R1246 gnd.n7225 gnd.n7224 585
R1247 gnd.n581 gnd.n580 585
R1248 gnd.n7226 gnd.n581 585
R1249 gnd.n7229 gnd.n7228 585
R1250 gnd.n7228 gnd.n7227 585
R1251 gnd.n578 gnd.n577 585
R1252 gnd.n577 gnd.n576 585
R1253 gnd.n7234 gnd.n7233 585
R1254 gnd.n7235 gnd.n7234 585
R1255 gnd.n575 gnd.n574 585
R1256 gnd.n7236 gnd.n575 585
R1257 gnd.n7239 gnd.n7238 585
R1258 gnd.n7238 gnd.n7237 585
R1259 gnd.n572 gnd.n571 585
R1260 gnd.n571 gnd.n570 585
R1261 gnd.n7244 gnd.n7243 585
R1262 gnd.n7245 gnd.n7244 585
R1263 gnd.n569 gnd.n568 585
R1264 gnd.n7246 gnd.n569 585
R1265 gnd.n7249 gnd.n7248 585
R1266 gnd.n7248 gnd.n7247 585
R1267 gnd.n566 gnd.n565 585
R1268 gnd.n565 gnd.n564 585
R1269 gnd.n7254 gnd.n7253 585
R1270 gnd.n7255 gnd.n7254 585
R1271 gnd.n563 gnd.n562 585
R1272 gnd.n7256 gnd.n563 585
R1273 gnd.n7259 gnd.n7258 585
R1274 gnd.n7258 gnd.n7257 585
R1275 gnd.n560 gnd.n559 585
R1276 gnd.n559 gnd.n558 585
R1277 gnd.n7264 gnd.n7263 585
R1278 gnd.n7265 gnd.n7264 585
R1279 gnd.n557 gnd.n556 585
R1280 gnd.n7266 gnd.n557 585
R1281 gnd.n7269 gnd.n7268 585
R1282 gnd.n7268 gnd.n7267 585
R1283 gnd.n554 gnd.n553 585
R1284 gnd.n553 gnd.n552 585
R1285 gnd.n7274 gnd.n7273 585
R1286 gnd.n7275 gnd.n7274 585
R1287 gnd.n551 gnd.n550 585
R1288 gnd.n7276 gnd.n551 585
R1289 gnd.n7279 gnd.n7278 585
R1290 gnd.n7278 gnd.n7277 585
R1291 gnd.n548 gnd.n547 585
R1292 gnd.n547 gnd.n546 585
R1293 gnd.n7284 gnd.n7283 585
R1294 gnd.n7285 gnd.n7284 585
R1295 gnd.n545 gnd.n544 585
R1296 gnd.n7286 gnd.n545 585
R1297 gnd.n7289 gnd.n7288 585
R1298 gnd.n7288 gnd.n7287 585
R1299 gnd.n542 gnd.n541 585
R1300 gnd.n541 gnd.n540 585
R1301 gnd.n7294 gnd.n7293 585
R1302 gnd.n7295 gnd.n7294 585
R1303 gnd.n539 gnd.n538 585
R1304 gnd.n7296 gnd.n539 585
R1305 gnd.n7299 gnd.n7298 585
R1306 gnd.n7298 gnd.n7297 585
R1307 gnd.n536 gnd.n535 585
R1308 gnd.n535 gnd.n534 585
R1309 gnd.n7304 gnd.n7303 585
R1310 gnd.n7305 gnd.n7304 585
R1311 gnd.n533 gnd.n532 585
R1312 gnd.n7306 gnd.n533 585
R1313 gnd.n7309 gnd.n7308 585
R1314 gnd.n7308 gnd.n7307 585
R1315 gnd.n530 gnd.n529 585
R1316 gnd.n529 gnd.n528 585
R1317 gnd.n7314 gnd.n7313 585
R1318 gnd.n7315 gnd.n7314 585
R1319 gnd.n527 gnd.n526 585
R1320 gnd.n7316 gnd.n527 585
R1321 gnd.n7319 gnd.n7318 585
R1322 gnd.n7318 gnd.n7317 585
R1323 gnd.n524 gnd.n523 585
R1324 gnd.n523 gnd.n522 585
R1325 gnd.n7324 gnd.n7323 585
R1326 gnd.n7325 gnd.n7324 585
R1327 gnd.n521 gnd.n520 585
R1328 gnd.n7326 gnd.n521 585
R1329 gnd.n7329 gnd.n7328 585
R1330 gnd.n7328 gnd.n7327 585
R1331 gnd.n518 gnd.n517 585
R1332 gnd.n517 gnd.n516 585
R1333 gnd.n7334 gnd.n7333 585
R1334 gnd.n7335 gnd.n7334 585
R1335 gnd.n515 gnd.n514 585
R1336 gnd.n7336 gnd.n515 585
R1337 gnd.n7339 gnd.n7338 585
R1338 gnd.n7338 gnd.n7337 585
R1339 gnd.n512 gnd.n511 585
R1340 gnd.n511 gnd.n510 585
R1341 gnd.n7344 gnd.n7343 585
R1342 gnd.n7345 gnd.n7344 585
R1343 gnd.n509 gnd.n508 585
R1344 gnd.n7346 gnd.n509 585
R1345 gnd.n7349 gnd.n7348 585
R1346 gnd.n7348 gnd.n7347 585
R1347 gnd.n506 gnd.n505 585
R1348 gnd.n505 gnd.n504 585
R1349 gnd.n7354 gnd.n7353 585
R1350 gnd.n7355 gnd.n7354 585
R1351 gnd.n503 gnd.n502 585
R1352 gnd.n7356 gnd.n503 585
R1353 gnd.n7359 gnd.n7358 585
R1354 gnd.n7358 gnd.n7357 585
R1355 gnd.n500 gnd.n499 585
R1356 gnd.n499 gnd.n498 585
R1357 gnd.n7365 gnd.n7364 585
R1358 gnd.n7366 gnd.n7365 585
R1359 gnd.n497 gnd.n496 585
R1360 gnd.n7367 gnd.n497 585
R1361 gnd.n7370 gnd.n7369 585
R1362 gnd.n7369 gnd.n7368 585
R1363 gnd.n7371 gnd.n494 585
R1364 gnd.n494 gnd.n493 585
R1365 gnd.n369 gnd.n368 585
R1366 gnd.n7578 gnd.n368 585
R1367 gnd.n7581 gnd.n7580 585
R1368 gnd.n7580 gnd.n7579 585
R1369 gnd.n372 gnd.n371 585
R1370 gnd.n7577 gnd.n372 585
R1371 gnd.n7575 gnd.n7574 585
R1372 gnd.n7576 gnd.n7575 585
R1373 gnd.n375 gnd.n374 585
R1374 gnd.n374 gnd.n373 585
R1375 gnd.n7570 gnd.n7569 585
R1376 gnd.n7569 gnd.n7568 585
R1377 gnd.n378 gnd.n377 585
R1378 gnd.n7567 gnd.n378 585
R1379 gnd.n7565 gnd.n7564 585
R1380 gnd.n7566 gnd.n7565 585
R1381 gnd.n381 gnd.n380 585
R1382 gnd.n380 gnd.n379 585
R1383 gnd.n7560 gnd.n7559 585
R1384 gnd.n7559 gnd.n7558 585
R1385 gnd.n384 gnd.n383 585
R1386 gnd.n7557 gnd.n384 585
R1387 gnd.n7555 gnd.n7554 585
R1388 gnd.n7556 gnd.n7555 585
R1389 gnd.n387 gnd.n386 585
R1390 gnd.n386 gnd.n385 585
R1391 gnd.n7550 gnd.n7549 585
R1392 gnd.n7549 gnd.n7548 585
R1393 gnd.n390 gnd.n389 585
R1394 gnd.n7547 gnd.n390 585
R1395 gnd.n7545 gnd.n7544 585
R1396 gnd.n7546 gnd.n7545 585
R1397 gnd.n393 gnd.n392 585
R1398 gnd.n392 gnd.n391 585
R1399 gnd.n7540 gnd.n7539 585
R1400 gnd.n7539 gnd.n7538 585
R1401 gnd.n396 gnd.n395 585
R1402 gnd.n7537 gnd.n396 585
R1403 gnd.n7535 gnd.n7534 585
R1404 gnd.n7536 gnd.n7535 585
R1405 gnd.n399 gnd.n398 585
R1406 gnd.n398 gnd.n397 585
R1407 gnd.n7530 gnd.n7529 585
R1408 gnd.n7529 gnd.n7528 585
R1409 gnd.n402 gnd.n401 585
R1410 gnd.n7527 gnd.n402 585
R1411 gnd.n7525 gnd.n7524 585
R1412 gnd.n7526 gnd.n7525 585
R1413 gnd.n405 gnd.n404 585
R1414 gnd.n404 gnd.n403 585
R1415 gnd.n7520 gnd.n7519 585
R1416 gnd.n7519 gnd.n7518 585
R1417 gnd.n408 gnd.n407 585
R1418 gnd.n7517 gnd.n408 585
R1419 gnd.n7515 gnd.n7514 585
R1420 gnd.n7516 gnd.n7515 585
R1421 gnd.n411 gnd.n410 585
R1422 gnd.n410 gnd.n409 585
R1423 gnd.n7510 gnd.n7509 585
R1424 gnd.n7509 gnd.n7508 585
R1425 gnd.n414 gnd.n413 585
R1426 gnd.n7507 gnd.n414 585
R1427 gnd.n7505 gnd.n7504 585
R1428 gnd.n7506 gnd.n7505 585
R1429 gnd.n417 gnd.n416 585
R1430 gnd.n416 gnd.n415 585
R1431 gnd.n7500 gnd.n7499 585
R1432 gnd.n7499 gnd.n7498 585
R1433 gnd.n420 gnd.n419 585
R1434 gnd.n7497 gnd.n420 585
R1435 gnd.n7495 gnd.n7494 585
R1436 gnd.n7496 gnd.n7495 585
R1437 gnd.n423 gnd.n422 585
R1438 gnd.n422 gnd.n421 585
R1439 gnd.n7490 gnd.n7489 585
R1440 gnd.n7489 gnd.n7488 585
R1441 gnd.n426 gnd.n425 585
R1442 gnd.n7487 gnd.n426 585
R1443 gnd.n7485 gnd.n7484 585
R1444 gnd.n7486 gnd.n7485 585
R1445 gnd.n429 gnd.n428 585
R1446 gnd.n428 gnd.n427 585
R1447 gnd.n7480 gnd.n7479 585
R1448 gnd.n7479 gnd.n7478 585
R1449 gnd.n432 gnd.n431 585
R1450 gnd.n7477 gnd.n432 585
R1451 gnd.n7475 gnd.n7474 585
R1452 gnd.n7476 gnd.n7475 585
R1453 gnd.n435 gnd.n434 585
R1454 gnd.n434 gnd.n433 585
R1455 gnd.n7470 gnd.n7469 585
R1456 gnd.n7469 gnd.n7468 585
R1457 gnd.n438 gnd.n437 585
R1458 gnd.n7467 gnd.n438 585
R1459 gnd.n7465 gnd.n7464 585
R1460 gnd.n7466 gnd.n7465 585
R1461 gnd.n441 gnd.n440 585
R1462 gnd.n440 gnd.n439 585
R1463 gnd.n7460 gnd.n7459 585
R1464 gnd.n7459 gnd.n7458 585
R1465 gnd.n444 gnd.n443 585
R1466 gnd.n7457 gnd.n444 585
R1467 gnd.n7455 gnd.n7454 585
R1468 gnd.n7456 gnd.n7455 585
R1469 gnd.n447 gnd.n446 585
R1470 gnd.n446 gnd.n445 585
R1471 gnd.n7450 gnd.n7449 585
R1472 gnd.n7449 gnd.n7448 585
R1473 gnd.n450 gnd.n449 585
R1474 gnd.n7447 gnd.n450 585
R1475 gnd.n7445 gnd.n7444 585
R1476 gnd.n7446 gnd.n7445 585
R1477 gnd.n453 gnd.n452 585
R1478 gnd.n452 gnd.n451 585
R1479 gnd.n7440 gnd.n7439 585
R1480 gnd.n7439 gnd.n7438 585
R1481 gnd.n456 gnd.n455 585
R1482 gnd.n7437 gnd.n456 585
R1483 gnd.n7435 gnd.n7434 585
R1484 gnd.n7436 gnd.n7435 585
R1485 gnd.n459 gnd.n458 585
R1486 gnd.n458 gnd.n457 585
R1487 gnd.n7430 gnd.n7429 585
R1488 gnd.n7429 gnd.n7428 585
R1489 gnd.n462 gnd.n461 585
R1490 gnd.n7427 gnd.n462 585
R1491 gnd.n7425 gnd.n7424 585
R1492 gnd.n7426 gnd.n7425 585
R1493 gnd.n465 gnd.n464 585
R1494 gnd.n464 gnd.n463 585
R1495 gnd.n7420 gnd.n7419 585
R1496 gnd.n7419 gnd.n7418 585
R1497 gnd.n468 gnd.n467 585
R1498 gnd.n7417 gnd.n468 585
R1499 gnd.n7415 gnd.n7414 585
R1500 gnd.n7416 gnd.n7415 585
R1501 gnd.n471 gnd.n470 585
R1502 gnd.n470 gnd.n469 585
R1503 gnd.n7410 gnd.n7409 585
R1504 gnd.n7409 gnd.n7408 585
R1505 gnd.n474 gnd.n473 585
R1506 gnd.n7407 gnd.n474 585
R1507 gnd.n7405 gnd.n7404 585
R1508 gnd.n7406 gnd.n7405 585
R1509 gnd.n477 gnd.n476 585
R1510 gnd.n476 gnd.n475 585
R1511 gnd.n7400 gnd.n7399 585
R1512 gnd.n7399 gnd.n7398 585
R1513 gnd.n480 gnd.n479 585
R1514 gnd.n7397 gnd.n480 585
R1515 gnd.n7395 gnd.n7394 585
R1516 gnd.n7396 gnd.n7395 585
R1517 gnd.n483 gnd.n482 585
R1518 gnd.n482 gnd.n481 585
R1519 gnd.n7390 gnd.n7389 585
R1520 gnd.n7389 gnd.n7388 585
R1521 gnd.n486 gnd.n485 585
R1522 gnd.n7387 gnd.n486 585
R1523 gnd.n7385 gnd.n7384 585
R1524 gnd.n7386 gnd.n7385 585
R1525 gnd.n489 gnd.n488 585
R1526 gnd.n488 gnd.n487 585
R1527 gnd.n7380 gnd.n7379 585
R1528 gnd.n7379 gnd.n7378 585
R1529 gnd.n492 gnd.n491 585
R1530 gnd.n7377 gnd.n492 585
R1531 gnd.n7375 gnd.n7374 585
R1532 gnd.n7376 gnd.n7375 585
R1533 gnd.n2754 gnd.n2753 585
R1534 gnd.n4768 gnd.n2754 585
R1535 gnd.n6334 gnd.n6333 585
R1536 gnd.n6333 gnd.n6332 585
R1537 gnd.n6335 gnd.n2749 585
R1538 gnd.n4760 gnd.n2749 585
R1539 gnd.n6337 gnd.n6336 585
R1540 gnd.n6338 gnd.n6337 585
R1541 gnd.n2733 gnd.n2732 585
R1542 gnd.n4473 gnd.n2733 585
R1543 gnd.n6346 gnd.n6345 585
R1544 gnd.n6345 gnd.n6344 585
R1545 gnd.n6347 gnd.n2728 585
R1546 gnd.n4465 gnd.n2728 585
R1547 gnd.n6349 gnd.n6348 585
R1548 gnd.n6350 gnd.n6349 585
R1549 gnd.n2714 gnd.n2713 585
R1550 gnd.n4459 gnd.n2714 585
R1551 gnd.n6358 gnd.n6357 585
R1552 gnd.n6357 gnd.n6356 585
R1553 gnd.n6359 gnd.n2709 585
R1554 gnd.n4451 gnd.n2709 585
R1555 gnd.n6361 gnd.n6360 585
R1556 gnd.n6362 gnd.n6361 585
R1557 gnd.n2693 gnd.n2692 585
R1558 gnd.n4391 gnd.n2693 585
R1559 gnd.n6370 gnd.n6369 585
R1560 gnd.n6369 gnd.n6368 585
R1561 gnd.n6371 gnd.n2688 585
R1562 gnd.n4382 gnd.n2688 585
R1563 gnd.n6373 gnd.n6372 585
R1564 gnd.n6374 gnd.n6373 585
R1565 gnd.n2674 gnd.n2673 585
R1566 gnd.n4377 gnd.n2674 585
R1567 gnd.n6382 gnd.n6381 585
R1568 gnd.n6381 gnd.n6380 585
R1569 gnd.n6383 gnd.n2669 585
R1570 gnd.n4405 gnd.n2669 585
R1571 gnd.n6385 gnd.n6384 585
R1572 gnd.n6386 gnd.n6385 585
R1573 gnd.n2653 gnd.n2652 585
R1574 gnd.n4370 gnd.n2653 585
R1575 gnd.n6394 gnd.n6393 585
R1576 gnd.n6393 gnd.n6392 585
R1577 gnd.n6395 gnd.n2648 585
R1578 gnd.n4362 gnd.n2648 585
R1579 gnd.n6397 gnd.n6396 585
R1580 gnd.n6398 gnd.n6397 585
R1581 gnd.n2635 gnd.n2634 585
R1582 gnd.n4356 gnd.n2635 585
R1583 gnd.n6406 gnd.n6405 585
R1584 gnd.n6405 gnd.n6404 585
R1585 gnd.n6407 gnd.n2629 585
R1586 gnd.n4348 gnd.n2629 585
R1587 gnd.n6409 gnd.n6408 585
R1588 gnd.n6410 gnd.n6409 585
R1589 gnd.n2630 gnd.n2628 585
R1590 gnd.n4317 gnd.n2628 585
R1591 gnd.n4299 gnd.n4298 585
R1592 gnd.n4298 gnd.n3988 585
R1593 gnd.n4300 gnd.n3998 585
R1594 gnd.n4309 gnd.n3998 585
R1595 gnd.n4302 gnd.n4301 585
R1596 gnd.n4303 gnd.n4302 585
R1597 gnd.n4005 gnd.n4004 585
R1598 gnd.n4287 gnd.n4004 585
R1599 gnd.n4240 gnd.n4239 585
R1600 gnd.n4239 gnd.n4238 585
R1601 gnd.n2607 gnd.n2606 585
R1602 gnd.n4279 gnd.n2607 585
R1603 gnd.n6419 gnd.n6418 585
R1604 gnd.n6418 gnd.n6417 585
R1605 gnd.n6420 gnd.n2602 585
R1606 gnd.n4247 gnd.n2602 585
R1607 gnd.n6422 gnd.n6421 585
R1608 gnd.n6423 gnd.n6422 585
R1609 gnd.n2588 gnd.n2587 585
R1610 gnd.n4253 gnd.n2588 585
R1611 gnd.n6431 gnd.n6430 585
R1612 gnd.n6430 gnd.n6429 585
R1613 gnd.n6432 gnd.n2583 585
R1614 gnd.n4229 gnd.n2583 585
R1615 gnd.n6434 gnd.n6433 585
R1616 gnd.n6435 gnd.n6434 585
R1617 gnd.n2568 gnd.n2567 585
R1618 gnd.n4220 gnd.n2568 585
R1619 gnd.n6443 gnd.n6442 585
R1620 gnd.n6442 gnd.n6441 585
R1621 gnd.n6444 gnd.n2563 585
R1622 gnd.n4183 gnd.n2563 585
R1623 gnd.n6446 gnd.n6445 585
R1624 gnd.n6447 gnd.n6446 585
R1625 gnd.n2548 gnd.n2547 585
R1626 gnd.n4189 gnd.n2548 585
R1627 gnd.n6455 gnd.n6454 585
R1628 gnd.n6454 gnd.n6453 585
R1629 gnd.n6456 gnd.n2543 585
R1630 gnd.n4171 gnd.n2543 585
R1631 gnd.n6458 gnd.n6457 585
R1632 gnd.n6459 gnd.n6458 585
R1633 gnd.n2528 gnd.n2527 585
R1634 gnd.n2532 gnd.n2528 585
R1635 gnd.n6467 gnd.n6466 585
R1636 gnd.n6466 gnd.n6465 585
R1637 gnd.n6468 gnd.n2523 585
R1638 gnd.n2523 gnd.n2522 585
R1639 gnd.n6470 gnd.n6469 585
R1640 gnd.n6471 gnd.n6470 585
R1641 gnd.n2509 gnd.n2508 585
R1642 gnd.n2519 gnd.n2509 585
R1643 gnd.n6479 gnd.n6478 585
R1644 gnd.n6478 gnd.n6477 585
R1645 gnd.n6480 gnd.n2504 585
R1646 gnd.n2504 gnd.n2503 585
R1647 gnd.n6482 gnd.n6481 585
R1648 gnd.n6483 gnd.n6482 585
R1649 gnd.n2490 gnd.n2489 585
R1650 gnd.n2493 gnd.n2490 585
R1651 gnd.n6491 gnd.n6490 585
R1652 gnd.n6490 gnd.n6489 585
R1653 gnd.n6492 gnd.n2483 585
R1654 gnd.n2483 gnd.n2481 585
R1655 gnd.n6494 gnd.n6493 585
R1656 gnd.n6495 gnd.n6494 585
R1657 gnd.n2485 gnd.n2482 585
R1658 gnd.n2482 gnd.n2478 585
R1659 gnd.n2484 gnd.n2469 585
R1660 gnd.n6501 gnd.n2469 585
R1661 gnd.n4091 gnd.n2463 585
R1662 gnd.n4091 gnd.n2394 585
R1663 gnd.n4093 gnd.n4092 585
R1664 gnd.n4095 gnd.n4094 585
R1665 gnd.n4097 gnd.n4096 585
R1666 gnd.n4101 gnd.n4089 585
R1667 gnd.n4103 gnd.n4102 585
R1668 gnd.n4105 gnd.n4104 585
R1669 gnd.n4107 gnd.n4106 585
R1670 gnd.n4111 gnd.n4087 585
R1671 gnd.n4113 gnd.n4112 585
R1672 gnd.n4115 gnd.n4114 585
R1673 gnd.n4117 gnd.n4116 585
R1674 gnd.n4121 gnd.n4085 585
R1675 gnd.n4123 gnd.n4122 585
R1676 gnd.n4125 gnd.n4124 585
R1677 gnd.n4127 gnd.n4126 585
R1678 gnd.n4082 gnd.n4081 585
R1679 gnd.n4131 gnd.n4083 585
R1680 gnd.n4132 gnd.n4078 585
R1681 gnd.n4133 gnd.n2393 585
R1682 gnd.n6625 gnd.n2393 585
R1683 gnd.n4602 gnd.n3936 585
R1684 gnd.n4594 gnd.n4593 585
R1685 gnd.n4609 gnd.n4590 585
R1686 gnd.n4610 gnd.n4589 585
R1687 gnd.n4588 gnd.n4580 585
R1688 gnd.n4617 gnd.n4579 585
R1689 gnd.n4618 gnd.n4578 585
R1690 gnd.n4572 gnd.n4571 585
R1691 gnd.n4625 gnd.n4570 585
R1692 gnd.n4626 gnd.n4569 585
R1693 gnd.n4568 gnd.n4560 585
R1694 gnd.n4633 gnd.n4559 585
R1695 gnd.n4634 gnd.n4558 585
R1696 gnd.n4552 gnd.n4551 585
R1697 gnd.n4641 gnd.n4550 585
R1698 gnd.n4642 gnd.n4549 585
R1699 gnd.n4548 gnd.n4540 585
R1700 gnd.n4649 gnd.n4539 585
R1701 gnd.n4650 gnd.n2766 585
R1702 gnd.n6324 gnd.n2766 585
R1703 gnd.n4767 gnd.n4766 585
R1704 gnd.n4768 gnd.n4767 585
R1705 gnd.n3937 gnd.n2757 585
R1706 gnd.n6332 gnd.n2757 585
R1707 gnd.n4762 gnd.n4761 585
R1708 gnd.n4761 gnd.n4760 585
R1709 gnd.n3939 gnd.n2747 585
R1710 gnd.n6338 gnd.n2747 585
R1711 gnd.n4472 gnd.n4471 585
R1712 gnd.n4473 gnd.n4472 585
R1713 gnd.n3942 gnd.n2736 585
R1714 gnd.n6344 gnd.n2736 585
R1715 gnd.n4467 gnd.n4466 585
R1716 gnd.n4466 gnd.n4465 585
R1717 gnd.n3944 gnd.n2727 585
R1718 gnd.n6350 gnd.n2727 585
R1719 gnd.n4458 gnd.n4457 585
R1720 gnd.n4459 gnd.n4458 585
R1721 gnd.n3948 gnd.n2716 585
R1722 gnd.n6356 gnd.n2716 585
R1723 gnd.n4453 gnd.n4452 585
R1724 gnd.n4452 gnd.n4451 585
R1725 gnd.n3950 gnd.n2707 585
R1726 gnd.n6362 gnd.n2707 585
R1727 gnd.n4393 gnd.n4392 585
R1728 gnd.n4392 gnd.n4391 585
R1729 gnd.n3970 gnd.n2696 585
R1730 gnd.n6368 gnd.n2696 585
R1731 gnd.n4397 gnd.n3969 585
R1732 gnd.n4382 gnd.n3969 585
R1733 gnd.n4398 gnd.n2687 585
R1734 gnd.n6374 gnd.n2687 585
R1735 gnd.n4399 gnd.n3968 585
R1736 gnd.n4377 gnd.n3968 585
R1737 gnd.n3965 gnd.n2676 585
R1738 gnd.n6380 gnd.n2676 585
R1739 gnd.n4404 gnd.n4403 585
R1740 gnd.n4405 gnd.n4404 585
R1741 gnd.n3964 gnd.n2667 585
R1742 gnd.n6386 gnd.n2667 585
R1743 gnd.n4369 gnd.n4368 585
R1744 gnd.n4370 gnd.n4369 585
R1745 gnd.n3973 gnd.n2656 585
R1746 gnd.n6392 gnd.n2656 585
R1747 gnd.n4364 gnd.n4363 585
R1748 gnd.n4363 gnd.n4362 585
R1749 gnd.n3975 gnd.n2647 585
R1750 gnd.n6398 gnd.n2647 585
R1751 gnd.n4355 gnd.n4354 585
R1752 gnd.n4356 gnd.n4355 585
R1753 gnd.n3979 gnd.n2637 585
R1754 gnd.n6404 gnd.n2637 585
R1755 gnd.n4350 gnd.n4349 585
R1756 gnd.n4349 gnd.n4348 585
R1757 gnd.n3981 gnd.n2626 585
R1758 gnd.n6410 gnd.n2626 585
R1759 gnd.n4316 gnd.n4315 585
R1760 gnd.n4317 gnd.n4316 585
R1761 gnd.n3991 gnd.n3990 585
R1762 gnd.n3990 gnd.n3988 585
R1763 gnd.n4311 gnd.n4310 585
R1764 gnd.n4310 gnd.n4309 585
R1765 gnd.n3994 gnd.n3993 585
R1766 gnd.n4303 gnd.n3994 585
R1767 gnd.n4286 gnd.n4285 585
R1768 gnd.n4287 gnd.n4286 585
R1769 gnd.n4014 gnd.n4013 585
R1770 gnd.n4238 gnd.n4013 585
R1771 gnd.n4281 gnd.n4280 585
R1772 gnd.n4280 gnd.n4279 585
R1773 gnd.n4016 gnd.n2610 585
R1774 gnd.n6417 gnd.n2610 585
R1775 gnd.n4249 gnd.n4248 585
R1776 gnd.n4248 gnd.n4247 585
R1777 gnd.n4250 gnd.n2600 585
R1778 gnd.n6423 gnd.n2600 585
R1779 gnd.n4252 gnd.n4251 585
R1780 gnd.n4253 gnd.n4252 585
R1781 gnd.n4027 gnd.n2591 585
R1782 gnd.n6429 gnd.n2591 585
R1783 gnd.n4228 gnd.n4227 585
R1784 gnd.n4229 gnd.n4228 585
R1785 gnd.n4032 gnd.n2581 585
R1786 gnd.n6435 gnd.n2581 585
R1787 gnd.n4222 gnd.n4221 585
R1788 gnd.n4221 gnd.n4220 585
R1789 gnd.n4034 gnd.n2571 585
R1790 gnd.n6441 gnd.n2571 585
R1791 gnd.n4185 gnd.n4184 585
R1792 gnd.n4184 gnd.n4183 585
R1793 gnd.n4186 gnd.n2561 585
R1794 gnd.n6447 gnd.n2561 585
R1795 gnd.n4188 gnd.n4187 585
R1796 gnd.n4189 gnd.n4188 585
R1797 gnd.n4041 gnd.n2551 585
R1798 gnd.n6453 gnd.n2551 585
R1799 gnd.n4170 gnd.n4169 585
R1800 gnd.n4171 gnd.n4170 585
R1801 gnd.n4069 gnd.n2541 585
R1802 gnd.n6459 gnd.n2541 585
R1803 gnd.n4164 gnd.n4163 585
R1804 gnd.n4163 gnd.n2532 585
R1805 gnd.n4162 gnd.n2531 585
R1806 gnd.n6465 gnd.n2531 585
R1807 gnd.n4161 gnd.n4160 585
R1808 gnd.n4160 gnd.n2522 585
R1809 gnd.n4071 gnd.n2521 585
R1810 gnd.n6471 gnd.n2521 585
R1811 gnd.n4156 gnd.n4155 585
R1812 gnd.n4155 gnd.n2519 585
R1813 gnd.n4154 gnd.n2511 585
R1814 gnd.n6477 gnd.n2511 585
R1815 gnd.n4153 gnd.n4152 585
R1816 gnd.n4152 gnd.n2503 585
R1817 gnd.n4073 gnd.n2502 585
R1818 gnd.n6483 gnd.n2502 585
R1819 gnd.n4148 gnd.n4147 585
R1820 gnd.n4147 gnd.n2493 585
R1821 gnd.n4146 gnd.n2492 585
R1822 gnd.n6489 gnd.n2492 585
R1823 gnd.n4145 gnd.n4144 585
R1824 gnd.n4144 gnd.n2481 585
R1825 gnd.n4075 gnd.n2480 585
R1826 gnd.n6495 gnd.n2480 585
R1827 gnd.n4140 gnd.n4139 585
R1828 gnd.n4139 gnd.n2478 585
R1829 gnd.n4138 gnd.n2468 585
R1830 gnd.n6501 gnd.n2468 585
R1831 gnd.n4137 gnd.n4136 585
R1832 gnd.n4136 gnd.n2394 585
R1833 gnd.n6687 gnd.n6686 585
R1834 gnd.n6688 gnd.n6687 585
R1835 gnd.n1007 gnd.n1005 585
R1836 gnd.n1005 gnd.n1001 585
R1837 gnd.n987 gnd.n986 585
R1838 gnd.n2346 gnd.n987 585
R1839 gnd.n6698 gnd.n6697 585
R1840 gnd.n6697 gnd.n6696 585
R1841 gnd.n6699 gnd.n981 585
R1842 gnd.n2022 gnd.n981 585
R1843 gnd.n6701 gnd.n6700 585
R1844 gnd.n6702 gnd.n6701 585
R1845 gnd.n982 gnd.n980 585
R1846 gnd.n980 gnd.n976 585
R1847 gnd.n963 gnd.n962 585
R1848 gnd.n967 gnd.n963 585
R1849 gnd.n6712 gnd.n6711 585
R1850 gnd.n6711 gnd.n6710 585
R1851 gnd.n6713 gnd.n957 585
R1852 gnd.n2031 gnd.n957 585
R1853 gnd.n6715 gnd.n6714 585
R1854 gnd.n6716 gnd.n6715 585
R1855 gnd.n958 gnd.n956 585
R1856 gnd.n2035 gnd.n956 585
R1857 gnd.n2059 gnd.n2058 585
R1858 gnd.n2058 gnd.n2057 585
R1859 gnd.n1122 gnd.n1121 585
R1860 gnd.n2041 gnd.n1122 585
R1861 gnd.n2001 gnd.n1141 585
R1862 gnd.n1141 gnd.n1131 585
R1863 gnd.n2003 gnd.n2002 585
R1864 gnd.n2004 gnd.n2003 585
R1865 gnd.n1142 gnd.n1140 585
R1866 gnd.n1149 gnd.n1140 585
R1867 gnd.n1977 gnd.n1161 585
R1868 gnd.n1926 gnd.n1161 585
R1869 gnd.n1979 gnd.n1978 585
R1870 gnd.n1980 gnd.n1979 585
R1871 gnd.n1162 gnd.n1160 585
R1872 gnd.n1160 gnd.n1156 585
R1873 gnd.n1965 gnd.n1964 585
R1874 gnd.n1964 gnd.n1963 585
R1875 gnd.n1167 gnd.n1166 585
R1876 gnd.n1176 gnd.n1167 585
R1877 gnd.n1954 gnd.n1953 585
R1878 gnd.n1953 gnd.n1952 585
R1879 gnd.n1174 gnd.n1173 585
R1880 gnd.n1940 gnd.n1174 585
R1881 gnd.n1911 gnd.n1192 585
R1882 gnd.n1192 gnd.n1183 585
R1883 gnd.n1913 gnd.n1912 585
R1884 gnd.n1914 gnd.n1913 585
R1885 gnd.n1193 gnd.n1191 585
R1886 gnd.n1201 gnd.n1191 585
R1887 gnd.n1888 gnd.n1213 585
R1888 gnd.n1213 gnd.n1200 585
R1889 gnd.n1890 gnd.n1889 585
R1890 gnd.n1891 gnd.n1890 585
R1891 gnd.n1214 gnd.n1212 585
R1892 gnd.n1212 gnd.n1208 585
R1893 gnd.n1876 gnd.n1875 585
R1894 gnd.n1875 gnd.n1874 585
R1895 gnd.n1219 gnd.n1218 585
R1896 gnd.n1223 gnd.n1219 585
R1897 gnd.n1860 gnd.n1859 585
R1898 gnd.n1861 gnd.n1860 585
R1899 gnd.n1233 gnd.n1232 585
R1900 gnd.n1851 gnd.n1232 585
R1901 gnd.n1351 gnd.n1350 585
R1902 gnd.n1351 gnd.n1240 585
R1903 gnd.n1838 gnd.n1837 585
R1904 gnd.n1837 gnd.n1836 585
R1905 gnd.n1839 gnd.n1343 585
R1906 gnd.n1816 gnd.n1343 585
R1907 gnd.n1841 gnd.n1840 585
R1908 gnd.n1842 gnd.n1841 585
R1909 gnd.n1344 gnd.n1342 585
R1910 gnd.n1824 gnd.n1342 585
R1911 gnd.n1808 gnd.n1807 585
R1912 gnd.n1807 gnd.n1361 585
R1913 gnd.n1806 gnd.n1366 585
R1914 gnd.n1806 gnd.n1805 585
R1915 gnd.n1791 gnd.n1367 585
R1916 gnd.n1375 gnd.n1367 585
R1917 gnd.n1793 gnd.n1792 585
R1918 gnd.n1794 gnd.n1793 585
R1919 gnd.n1378 gnd.n1377 585
R1920 gnd.n1385 gnd.n1377 585
R1921 gnd.n1766 gnd.n1765 585
R1922 gnd.n1767 gnd.n1766 585
R1923 gnd.n1397 gnd.n1396 585
R1924 gnd.n1396 gnd.n1392 585
R1925 gnd.n1756 gnd.n1755 585
R1926 gnd.n1757 gnd.n1756 585
R1927 gnd.n1407 gnd.n1406 585
R1928 gnd.n1412 gnd.n1406 585
R1929 gnd.n1734 gnd.n1425 585
R1930 gnd.n1425 gnd.n1411 585
R1931 gnd.n1736 gnd.n1735 585
R1932 gnd.n1737 gnd.n1736 585
R1933 gnd.n1426 gnd.n1424 585
R1934 gnd.n1424 gnd.n1420 585
R1935 gnd.n1725 gnd.n1724 585
R1936 gnd.n1726 gnd.n1725 585
R1937 gnd.n1433 gnd.n1432 585
R1938 gnd.n1437 gnd.n1432 585
R1939 gnd.n1702 gnd.n1454 585
R1940 gnd.n1454 gnd.n1436 585
R1941 gnd.n1704 gnd.n1703 585
R1942 gnd.n1705 gnd.n1704 585
R1943 gnd.n1455 gnd.n1453 585
R1944 gnd.n1453 gnd.n1444 585
R1945 gnd.n1697 gnd.n1696 585
R1946 gnd.n1696 gnd.n1695 585
R1947 gnd.n1502 gnd.n1501 585
R1948 gnd.n1503 gnd.n1502 585
R1949 gnd.n1656 gnd.n1655 585
R1950 gnd.n1657 gnd.n1656 585
R1951 gnd.n1512 gnd.n1511 585
R1952 gnd.n1511 gnd.n1510 585
R1953 gnd.n1651 gnd.n1650 585
R1954 gnd.n1650 gnd.n1649 585
R1955 gnd.n1515 gnd.n1514 585
R1956 gnd.n1516 gnd.n1515 585
R1957 gnd.n1640 gnd.n1639 585
R1958 gnd.n1641 gnd.n1640 585
R1959 gnd.n1523 gnd.n1522 585
R1960 gnd.n1632 gnd.n1522 585
R1961 gnd.n1635 gnd.n1634 585
R1962 gnd.n1634 gnd.n1633 585
R1963 gnd.n1526 gnd.n1525 585
R1964 gnd.n1527 gnd.n1526 585
R1965 gnd.n1621 gnd.n1620 585
R1966 gnd.n1619 gnd.n1545 585
R1967 gnd.n1618 gnd.n1544 585
R1968 gnd.n1623 gnd.n1544 585
R1969 gnd.n1617 gnd.n1616 585
R1970 gnd.n1615 gnd.n1614 585
R1971 gnd.n1613 gnd.n1612 585
R1972 gnd.n1611 gnd.n1610 585
R1973 gnd.n1609 gnd.n1608 585
R1974 gnd.n1607 gnd.n1606 585
R1975 gnd.n1605 gnd.n1604 585
R1976 gnd.n1603 gnd.n1602 585
R1977 gnd.n1601 gnd.n1600 585
R1978 gnd.n1599 gnd.n1598 585
R1979 gnd.n1597 gnd.n1596 585
R1980 gnd.n1595 gnd.n1594 585
R1981 gnd.n1593 gnd.n1592 585
R1982 gnd.n1591 gnd.n1590 585
R1983 gnd.n1589 gnd.n1588 585
R1984 gnd.n1587 gnd.n1586 585
R1985 gnd.n1585 gnd.n1584 585
R1986 gnd.n1583 gnd.n1582 585
R1987 gnd.n1581 gnd.n1580 585
R1988 gnd.n1579 gnd.n1578 585
R1989 gnd.n1577 gnd.n1576 585
R1990 gnd.n1575 gnd.n1574 585
R1991 gnd.n1532 gnd.n1531 585
R1992 gnd.n1626 gnd.n1625 585
R1993 gnd.n2354 gnd.n2353 585
R1994 gnd.n1031 gnd.n1030 585
R1995 gnd.n1107 gnd.n1106 585
R1996 gnd.n1105 gnd.n1104 585
R1997 gnd.n1103 gnd.n1102 585
R1998 gnd.n1096 gnd.n1036 585
R1999 gnd.n1098 gnd.n1097 585
R2000 gnd.n1095 gnd.n1094 585
R2001 gnd.n1093 gnd.n1092 585
R2002 gnd.n1086 gnd.n1038 585
R2003 gnd.n1088 gnd.n1087 585
R2004 gnd.n1085 gnd.n1084 585
R2005 gnd.n1083 gnd.n1082 585
R2006 gnd.n1076 gnd.n1040 585
R2007 gnd.n1078 gnd.n1077 585
R2008 gnd.n1075 gnd.n1074 585
R2009 gnd.n1073 gnd.n1072 585
R2010 gnd.n1066 gnd.n1042 585
R2011 gnd.n1068 gnd.n1067 585
R2012 gnd.n1065 gnd.n1064 585
R2013 gnd.n1063 gnd.n1062 585
R2014 gnd.n1056 gnd.n1044 585
R2015 gnd.n1058 gnd.n1057 585
R2016 gnd.n1055 gnd.n1054 585
R2017 gnd.n1053 gnd.n1052 585
R2018 gnd.n1047 gnd.n1046 585
R2019 gnd.n1048 gnd.n1006 585
R2020 gnd.n6672 gnd.n1006 585
R2021 gnd.n2350 gnd.n1003 585
R2022 gnd.n6688 gnd.n1003 585
R2023 gnd.n2349 gnd.n2348 585
R2024 gnd.n2348 gnd.n1001 585
R2025 gnd.n2347 gnd.n1111 585
R2026 gnd.n2347 gnd.n2346 585
R2027 gnd.n2021 gnd.n989 585
R2028 gnd.n6696 gnd.n989 585
R2029 gnd.n2024 gnd.n2023 585
R2030 gnd.n2023 gnd.n2022 585
R2031 gnd.n2025 gnd.n978 585
R2032 gnd.n6702 gnd.n978 585
R2033 gnd.n2027 gnd.n2026 585
R2034 gnd.n2027 gnd.n976 585
R2035 gnd.n2029 gnd.n2028 585
R2036 gnd.n2028 gnd.n967 585
R2037 gnd.n2030 gnd.n965 585
R2038 gnd.n6710 gnd.n965 585
R2039 gnd.n2033 gnd.n2032 585
R2040 gnd.n2032 gnd.n2031 585
R2041 gnd.n2034 gnd.n954 585
R2042 gnd.n6716 gnd.n954 585
R2043 gnd.n2037 gnd.n2036 585
R2044 gnd.n2036 gnd.n2035 585
R2045 gnd.n2038 gnd.n1124 585
R2046 gnd.n2057 gnd.n1124 585
R2047 gnd.n2040 gnd.n2039 585
R2048 gnd.n2041 gnd.n2040 585
R2049 gnd.n1134 gnd.n1133 585
R2050 gnd.n1133 gnd.n1131 585
R2051 gnd.n2006 gnd.n2005 585
R2052 gnd.n2005 gnd.n2004 585
R2053 gnd.n1137 gnd.n1136 585
R2054 gnd.n1149 gnd.n1137 585
R2055 gnd.n1928 gnd.n1927 585
R2056 gnd.n1927 gnd.n1926 585
R2057 gnd.n1929 gnd.n1158 585
R2058 gnd.n1980 gnd.n1158 585
R2059 gnd.n1931 gnd.n1930 585
R2060 gnd.n1930 gnd.n1156 585
R2061 gnd.n1932 gnd.n1169 585
R2062 gnd.n1963 gnd.n1169 585
R2063 gnd.n1934 gnd.n1933 585
R2064 gnd.n1933 gnd.n1176 585
R2065 gnd.n1935 gnd.n1175 585
R2066 gnd.n1952 gnd.n1175 585
R2067 gnd.n1937 gnd.n1936 585
R2068 gnd.n1940 gnd.n1937 585
R2069 gnd.n1186 gnd.n1185 585
R2070 gnd.n1185 gnd.n1183 585
R2071 gnd.n1916 gnd.n1915 585
R2072 gnd.n1915 gnd.n1914 585
R2073 gnd.n1189 gnd.n1188 585
R2074 gnd.n1201 gnd.n1189 585
R2075 gnd.n1248 gnd.n1247 585
R2076 gnd.n1247 gnd.n1200 585
R2077 gnd.n1249 gnd.n1210 585
R2078 gnd.n1891 gnd.n1210 585
R2079 gnd.n1251 gnd.n1250 585
R2080 gnd.n1250 gnd.n1208 585
R2081 gnd.n1252 gnd.n1220 585
R2082 gnd.n1874 gnd.n1220 585
R2083 gnd.n1244 gnd.n1243 585
R2084 gnd.n1243 gnd.n1223 585
R2085 gnd.n1848 gnd.n1230 585
R2086 gnd.n1861 gnd.n1230 585
R2087 gnd.n1850 gnd.n1849 585
R2088 gnd.n1851 gnd.n1850 585
R2089 gnd.n1352 gnd.n1241 585
R2090 gnd.n1241 gnd.n1240 585
R2091 gnd.n1354 gnd.n1353 585
R2092 gnd.n1836 gnd.n1354 585
R2093 gnd.n1339 gnd.n1337 585
R2094 gnd.n1816 gnd.n1339 585
R2095 gnd.n1844 gnd.n1843 585
R2096 gnd.n1843 gnd.n1842 585
R2097 gnd.n1338 gnd.n1336 585
R2098 gnd.n1824 gnd.n1338 585
R2099 gnd.n1801 gnd.n1370 585
R2100 gnd.n1370 gnd.n1361 585
R2101 gnd.n1803 gnd.n1802 585
R2102 gnd.n1805 gnd.n1803 585
R2103 gnd.n1371 gnd.n1369 585
R2104 gnd.n1375 gnd.n1369 585
R2105 gnd.n1796 gnd.n1795 585
R2106 gnd.n1795 gnd.n1794 585
R2107 gnd.n1374 gnd.n1373 585
R2108 gnd.n1385 gnd.n1374 585
R2109 gnd.n1675 gnd.n1394 585
R2110 gnd.n1767 gnd.n1394 585
R2111 gnd.n1677 gnd.n1676 585
R2112 gnd.n1676 gnd.n1392 585
R2113 gnd.n1678 gnd.n1405 585
R2114 gnd.n1757 gnd.n1405 585
R2115 gnd.n1680 gnd.n1679 585
R2116 gnd.n1680 gnd.n1412 585
R2117 gnd.n1682 gnd.n1681 585
R2118 gnd.n1681 gnd.n1411 585
R2119 gnd.n1683 gnd.n1422 585
R2120 gnd.n1737 gnd.n1422 585
R2121 gnd.n1685 gnd.n1684 585
R2122 gnd.n1684 gnd.n1420 585
R2123 gnd.n1686 gnd.n1431 585
R2124 gnd.n1726 gnd.n1431 585
R2125 gnd.n1688 gnd.n1687 585
R2126 gnd.n1688 gnd.n1437 585
R2127 gnd.n1690 gnd.n1689 585
R2128 gnd.n1689 gnd.n1436 585
R2129 gnd.n1691 gnd.n1452 585
R2130 gnd.n1705 gnd.n1452 585
R2131 gnd.n1692 gnd.n1505 585
R2132 gnd.n1505 gnd.n1444 585
R2133 gnd.n1694 gnd.n1693 585
R2134 gnd.n1695 gnd.n1694 585
R2135 gnd.n1506 gnd.n1504 585
R2136 gnd.n1504 gnd.n1503 585
R2137 gnd.n1659 gnd.n1658 585
R2138 gnd.n1658 gnd.n1657 585
R2139 gnd.n1509 gnd.n1508 585
R2140 gnd.n1510 gnd.n1509 585
R2141 gnd.n1648 gnd.n1647 585
R2142 gnd.n1649 gnd.n1648 585
R2143 gnd.n1518 gnd.n1517 585
R2144 gnd.n1517 gnd.n1516 585
R2145 gnd.n1643 gnd.n1642 585
R2146 gnd.n1642 gnd.n1641 585
R2147 gnd.n1521 gnd.n1520 585
R2148 gnd.n1632 gnd.n1521 585
R2149 gnd.n1631 gnd.n1630 585
R2150 gnd.n1633 gnd.n1631 585
R2151 gnd.n1529 gnd.n1528 585
R2152 gnd.n1528 gnd.n1527 585
R2153 gnd.n246 gnd.n245 585
R2154 gnd.n249 gnd.n246 585
R2155 gnd.n7863 gnd.n7862 585
R2156 gnd.n7862 gnd.n7861 585
R2157 gnd.n7864 gnd.n241 585
R2158 gnd.n241 gnd.n240 585
R2159 gnd.n7866 gnd.n7865 585
R2160 gnd.n7867 gnd.n7866 585
R2161 gnd.n226 gnd.n225 585
R2162 gnd.n230 gnd.n226 585
R2163 gnd.n7875 gnd.n7874 585
R2164 gnd.n7874 gnd.n7873 585
R2165 gnd.n7876 gnd.n221 585
R2166 gnd.n227 gnd.n221 585
R2167 gnd.n7878 gnd.n7877 585
R2168 gnd.n7879 gnd.n7878 585
R2169 gnd.n208 gnd.n207 585
R2170 gnd.n211 gnd.n208 585
R2171 gnd.n7887 gnd.n7886 585
R2172 gnd.n7886 gnd.n7885 585
R2173 gnd.n7888 gnd.n203 585
R2174 gnd.n203 gnd.n202 585
R2175 gnd.n7890 gnd.n7889 585
R2176 gnd.n7891 gnd.n7890 585
R2177 gnd.n187 gnd.n186 585
R2178 gnd.n199 gnd.n187 585
R2179 gnd.n7899 gnd.n7898 585
R2180 gnd.n7898 gnd.n7897 585
R2181 gnd.n7900 gnd.n182 585
R2182 gnd.n188 gnd.n182 585
R2183 gnd.n7902 gnd.n7901 585
R2184 gnd.n7903 gnd.n7902 585
R2185 gnd.n168 gnd.n167 585
R2186 gnd.n7701 gnd.n168 585
R2187 gnd.n7911 gnd.n7910 585
R2188 gnd.n7910 gnd.n7909 585
R2189 gnd.n7912 gnd.n163 585
R2190 gnd.n7596 gnd.n163 585
R2191 gnd.n7914 gnd.n7913 585
R2192 gnd.n7915 gnd.n7914 585
R2193 gnd.n147 gnd.n146 585
R2194 gnd.n5765 gnd.n147 585
R2195 gnd.n7923 gnd.n7922 585
R2196 gnd.n7922 gnd.n7921 585
R2197 gnd.n7924 gnd.n142 585
R2198 gnd.n5771 gnd.n142 585
R2199 gnd.n7926 gnd.n7925 585
R2200 gnd.n7927 gnd.n7926 585
R2201 gnd.n129 gnd.n128 585
R2202 gnd.n5777 gnd.n129 585
R2203 gnd.n7935 gnd.n7934 585
R2204 gnd.n7934 gnd.n7933 585
R2205 gnd.n7936 gnd.n123 585
R2206 gnd.n5783 gnd.n123 585
R2207 gnd.n7938 gnd.n7937 585
R2208 gnd.n7939 gnd.n7938 585
R2209 gnd.n124 gnd.n122 585
R2210 gnd.n5722 gnd.n122 585
R2211 gnd.n5794 gnd.n5793 585
R2212 gnd.n5795 gnd.n5794 585
R2213 gnd.n3347 gnd.n104 585
R2214 gnd.n7947 gnd.n104 585
R2215 gnd.n5803 gnd.n5802 585
R2216 gnd.n5802 gnd.n5801 585
R2217 gnd.n5804 gnd.n3342 585
R2218 gnd.n3350 gnd.n3342 585
R2219 gnd.n5806 gnd.n5805 585
R2220 gnd.n5807 gnd.n5806 585
R2221 gnd.n3343 gnd.n3332 585
R2222 gnd.n5812 gnd.n3332 585
R2223 gnd.n5693 gnd.n5692 585
R2224 gnd.n5692 gnd.n3328 585
R2225 gnd.n5691 gnd.n5690 585
R2226 gnd.n5691 gnd.n3321 585
R2227 gnd.n3313 gnd.n3312 585
R2228 gnd.n5821 gnd.n3313 585
R2229 gnd.n5828 gnd.n5827 585
R2230 gnd.n5827 gnd.n5826 585
R2231 gnd.n5829 gnd.n3308 585
R2232 gnd.n5681 gnd.n3308 585
R2233 gnd.n5831 gnd.n5830 585
R2234 gnd.n5832 gnd.n5831 585
R2235 gnd.n3291 gnd.n3290 585
R2236 gnd.n5661 gnd.n3291 585
R2237 gnd.n5840 gnd.n5839 585
R2238 gnd.n5839 gnd.n5838 585
R2239 gnd.n5841 gnd.n3286 585
R2240 gnd.n5654 gnd.n3286 585
R2241 gnd.n5843 gnd.n5842 585
R2242 gnd.n5844 gnd.n5843 585
R2243 gnd.n3271 gnd.n3270 585
R2244 gnd.n5646 gnd.n3271 585
R2245 gnd.n5852 gnd.n5851 585
R2246 gnd.n5851 gnd.n5850 585
R2247 gnd.n5853 gnd.n3266 585
R2248 gnd.n5639 gnd.n3266 585
R2249 gnd.n5855 gnd.n5854 585
R2250 gnd.n5856 gnd.n5855 585
R2251 gnd.n3250 gnd.n3249 585
R2252 gnd.n5631 gnd.n3250 585
R2253 gnd.n5864 gnd.n5863 585
R2254 gnd.n5863 gnd.n5862 585
R2255 gnd.n5865 gnd.n3245 585
R2256 gnd.n5624 gnd.n3245 585
R2257 gnd.n5867 gnd.n5866 585
R2258 gnd.n5868 gnd.n5867 585
R2259 gnd.n3230 gnd.n3229 585
R2260 gnd.n5616 gnd.n3230 585
R2261 gnd.n5876 gnd.n5875 585
R2262 gnd.n5875 gnd.n5874 585
R2263 gnd.n5877 gnd.n3225 585
R2264 gnd.n5609 gnd.n3225 585
R2265 gnd.n5879 gnd.n5878 585
R2266 gnd.n5880 gnd.n5879 585
R2267 gnd.n3209 gnd.n3208 585
R2268 gnd.n5601 gnd.n3209 585
R2269 gnd.n5888 gnd.n5887 585
R2270 gnd.n5887 gnd.n5886 585
R2271 gnd.n5889 gnd.n3202 585
R2272 gnd.n5594 gnd.n3202 585
R2273 gnd.n5891 gnd.n5890 585
R2274 gnd.n5892 gnd.n5891 585
R2275 gnd.n3203 gnd.n3201 585
R2276 gnd.n5586 gnd.n3201 585
R2277 gnd.n3185 gnd.n3179 585
R2278 gnd.n5898 gnd.n3185 585
R2279 gnd.n5903 gnd.n3177 585
R2280 gnd.n5562 gnd.n3177 585
R2281 gnd.n5905 gnd.n5904 585
R2282 gnd.n5906 gnd.n5905 585
R2283 gnd.n3176 gnd.n3016 585
R2284 gnd.n6073 gnd.n3017 585
R2285 gnd.n6072 gnd.n3018 585
R2286 gnd.n3093 gnd.n3019 585
R2287 gnd.n6065 gnd.n3025 585
R2288 gnd.n6064 gnd.n3026 585
R2289 gnd.n3096 gnd.n3027 585
R2290 gnd.n6057 gnd.n3033 585
R2291 gnd.n6056 gnd.n3034 585
R2292 gnd.n3098 gnd.n3035 585
R2293 gnd.n6049 gnd.n3041 585
R2294 gnd.n6048 gnd.n3042 585
R2295 gnd.n3101 gnd.n3043 585
R2296 gnd.n6041 gnd.n3049 585
R2297 gnd.n6040 gnd.n3050 585
R2298 gnd.n3103 gnd.n3051 585
R2299 gnd.n6033 gnd.n3059 585
R2300 gnd.n6032 gnd.n6029 585
R2301 gnd.n3062 gnd.n3060 585
R2302 gnd.n6027 gnd.n3062 585
R2303 gnd.n7674 gnd.n7673 585
R2304 gnd.n7667 gnd.n7620 585
R2305 gnd.n7669 gnd.n7668 585
R2306 gnd.n7666 gnd.n7665 585
R2307 gnd.n7664 gnd.n7663 585
R2308 gnd.n7657 gnd.n7622 585
R2309 gnd.n7659 gnd.n7658 585
R2310 gnd.n7656 gnd.n7655 585
R2311 gnd.n7654 gnd.n7653 585
R2312 gnd.n7647 gnd.n7624 585
R2313 gnd.n7649 gnd.n7648 585
R2314 gnd.n7646 gnd.n7645 585
R2315 gnd.n7644 gnd.n7643 585
R2316 gnd.n7637 gnd.n7626 585
R2317 gnd.n7639 gnd.n7638 585
R2318 gnd.n7636 gnd.n7635 585
R2319 gnd.n7634 gnd.n7633 585
R2320 gnd.n7630 gnd.n7629 585
R2321 gnd.n7628 gnd.n257 585
R2322 gnd.n7853 gnd.n257 585
R2323 gnd.n7676 gnd.n7675 585
R2324 gnd.n7675 gnd.n249 585
R2325 gnd.n7677 gnd.n248 585
R2326 gnd.n7861 gnd.n248 585
R2327 gnd.n7679 gnd.n7678 585
R2328 gnd.n7678 gnd.n240 585
R2329 gnd.n7680 gnd.n239 585
R2330 gnd.n7867 gnd.n239 585
R2331 gnd.n7682 gnd.n7681 585
R2332 gnd.n7681 gnd.n230 585
R2333 gnd.n7683 gnd.n229 585
R2334 gnd.n7873 gnd.n229 585
R2335 gnd.n7685 gnd.n7684 585
R2336 gnd.n7684 gnd.n227 585
R2337 gnd.n7686 gnd.n220 585
R2338 gnd.n7879 gnd.n220 585
R2339 gnd.n7688 gnd.n7687 585
R2340 gnd.n7687 gnd.n211 585
R2341 gnd.n7689 gnd.n210 585
R2342 gnd.n7885 gnd.n210 585
R2343 gnd.n7691 gnd.n7690 585
R2344 gnd.n7690 gnd.n202 585
R2345 gnd.n7692 gnd.n201 585
R2346 gnd.n7891 gnd.n201 585
R2347 gnd.n7694 gnd.n7693 585
R2348 gnd.n7693 gnd.n199 585
R2349 gnd.n7695 gnd.n190 585
R2350 gnd.n7897 gnd.n190 585
R2351 gnd.n7697 gnd.n7696 585
R2352 gnd.n7696 gnd.n188 585
R2353 gnd.n7698 gnd.n181 585
R2354 gnd.n7903 gnd.n181 585
R2355 gnd.n7700 gnd.n7699 585
R2356 gnd.n7701 gnd.n7700 585
R2357 gnd.n357 gnd.n170 585
R2358 gnd.n7909 gnd.n170 585
R2359 gnd.n7598 gnd.n7597 585
R2360 gnd.n7597 gnd.n7596 585
R2361 gnd.n359 gnd.n161 585
R2362 gnd.n7915 gnd.n161 585
R2363 gnd.n5767 gnd.n5766 585
R2364 gnd.n5766 gnd.n5765 585
R2365 gnd.n5768 gnd.n150 585
R2366 gnd.n7921 gnd.n150 585
R2367 gnd.n5770 gnd.n5769 585
R2368 gnd.n5771 gnd.n5770 585
R2369 gnd.n5730 gnd.n141 585
R2370 gnd.n7927 gnd.n141 585
R2371 gnd.n5779 gnd.n5778 585
R2372 gnd.n5778 gnd.n5777 585
R2373 gnd.n5780 gnd.n131 585
R2374 gnd.n7933 gnd.n131 585
R2375 gnd.n5782 gnd.n5781 585
R2376 gnd.n5783 gnd.n5782 585
R2377 gnd.n5720 gnd.n120 585
R2378 gnd.n7939 gnd.n120 585
R2379 gnd.n5724 gnd.n5723 585
R2380 gnd.n5723 gnd.n5722 585
R2381 gnd.n100 gnd.n99 585
R2382 gnd.n5795 gnd.n100 585
R2383 gnd.n7949 gnd.n7948 585
R2384 gnd.n7948 gnd.n7947 585
R2385 gnd.n7950 gnd.n98 585
R2386 gnd.n5801 gnd.n98 585
R2387 gnd.n3349 gnd.n96 585
R2388 gnd.n3350 gnd.n3349 585
R2389 gnd.n5669 gnd.n3340 585
R2390 gnd.n5807 gnd.n3340 585
R2391 gnd.n5670 gnd.n3330 585
R2392 gnd.n5812 gnd.n3330 585
R2393 gnd.n5673 gnd.n5668 585
R2394 gnd.n5668 gnd.n3328 585
R2395 gnd.n5674 gnd.n5667 585
R2396 gnd.n5667 gnd.n3321 585
R2397 gnd.n5675 gnd.n3320 585
R2398 gnd.n5821 gnd.n3320 585
R2399 gnd.n3356 gnd.n3316 585
R2400 gnd.n5826 gnd.n3316 585
R2401 gnd.n5680 gnd.n5679 585
R2402 gnd.n5681 gnd.n5680 585
R2403 gnd.n3355 gnd.n3306 585
R2404 gnd.n5832 gnd.n3306 585
R2405 gnd.n5663 gnd.n5662 585
R2406 gnd.n5662 gnd.n5661 585
R2407 gnd.n3358 gnd.n3294 585
R2408 gnd.n5838 gnd.n3294 585
R2409 gnd.n5653 gnd.n5652 585
R2410 gnd.n5654 gnd.n5653 585
R2411 gnd.n3361 gnd.n3285 585
R2412 gnd.n5844 gnd.n3285 585
R2413 gnd.n5648 gnd.n5647 585
R2414 gnd.n5647 gnd.n5646 585
R2415 gnd.n3363 gnd.n3274 585
R2416 gnd.n5850 gnd.n3274 585
R2417 gnd.n5638 gnd.n5637 585
R2418 gnd.n5639 gnd.n5638 585
R2419 gnd.n3365 gnd.n3264 585
R2420 gnd.n5856 gnd.n3264 585
R2421 gnd.n5633 gnd.n5632 585
R2422 gnd.n5632 gnd.n5631 585
R2423 gnd.n3367 gnd.n3253 585
R2424 gnd.n5862 gnd.n3253 585
R2425 gnd.n5623 gnd.n5622 585
R2426 gnd.n5624 gnd.n5623 585
R2427 gnd.n3370 gnd.n3244 585
R2428 gnd.n5868 gnd.n3244 585
R2429 gnd.n5618 gnd.n5617 585
R2430 gnd.n5617 gnd.n5616 585
R2431 gnd.n3372 gnd.n3233 585
R2432 gnd.n5874 gnd.n3233 585
R2433 gnd.n5608 gnd.n5607 585
R2434 gnd.n5609 gnd.n5608 585
R2435 gnd.n3374 gnd.n3223 585
R2436 gnd.n5880 gnd.n3223 585
R2437 gnd.n5603 gnd.n5602 585
R2438 gnd.n5602 gnd.n5601 585
R2439 gnd.n3376 gnd.n3212 585
R2440 gnd.n5886 gnd.n3212 585
R2441 gnd.n5593 gnd.n5592 585
R2442 gnd.n5594 gnd.n5593 585
R2443 gnd.n3378 gnd.n3199 585
R2444 gnd.n5892 gnd.n3199 585
R2445 gnd.n5588 gnd.n5587 585
R2446 gnd.n5587 gnd.n5586 585
R2447 gnd.n5585 gnd.n3183 585
R2448 gnd.n5898 gnd.n3183 585
R2449 gnd.n5584 gnd.n3381 585
R2450 gnd.n5562 gnd.n3381 585
R2451 gnd.n3380 gnd.n3174 585
R2452 gnd.n5906 gnd.n3174 585
R2453 gnd.n1000 gnd.n999 585
R2454 gnd.n1004 gnd.n1000 585
R2455 gnd.n6691 gnd.n6690 585
R2456 gnd.n6690 gnd.n6689 585
R2457 gnd.n6692 gnd.n992 585
R2458 gnd.n2345 gnd.n992 585
R2459 gnd.n6694 gnd.n6693 585
R2460 gnd.n6695 gnd.n6694 585
R2461 gnd.n993 gnd.n991 585
R2462 gnd.n991 gnd.n988 585
R2463 gnd.n975 gnd.n974 585
R2464 gnd.n979 gnd.n975 585
R2465 gnd.n6705 gnd.n6704 585
R2466 gnd.n6704 gnd.n6703 585
R2467 gnd.n6706 gnd.n969 585
R2468 gnd.n1112 gnd.n969 585
R2469 gnd.n6708 gnd.n6707 585
R2470 gnd.n6709 gnd.n6708 585
R2471 gnd.n970 gnd.n968 585
R2472 gnd.n968 gnd.n964 585
R2473 gnd.n2052 gnd.n2051 585
R2474 gnd.n2051 gnd.n955 585
R2475 gnd.n2053 gnd.n1126 585
R2476 gnd.n1126 gnd.n953 585
R2477 gnd.n2055 gnd.n2054 585
R2478 gnd.n2056 gnd.n2055 585
R2479 gnd.n1127 gnd.n1125 585
R2480 gnd.n1125 gnd.n1123 585
R2481 gnd.n2044 gnd.n2043 585
R2482 gnd.n2043 gnd.n2042 585
R2483 gnd.n1130 gnd.n1129 585
R2484 gnd.n1139 gnd.n1130 585
R2485 gnd.n1988 gnd.n1151 585
R2486 gnd.n1151 gnd.n1138 585
R2487 gnd.n1990 gnd.n1989 585
R2488 gnd.n1991 gnd.n1990 585
R2489 gnd.n1152 gnd.n1150 585
R2490 gnd.n1159 gnd.n1150 585
R2491 gnd.n1983 gnd.n1982 585
R2492 gnd.n1982 gnd.n1981 585
R2493 gnd.n1155 gnd.n1154 585
R2494 gnd.n1962 gnd.n1155 585
R2495 gnd.n1948 gnd.n1178 585
R2496 gnd.n1178 gnd.n1168 585
R2497 gnd.n1950 gnd.n1949 585
R2498 gnd.n1951 gnd.n1950 585
R2499 gnd.n1179 gnd.n1177 585
R2500 gnd.n1939 gnd.n1177 585
R2501 gnd.n1943 gnd.n1942 585
R2502 gnd.n1942 gnd.n1941 585
R2503 gnd.n1182 gnd.n1181 585
R2504 gnd.n1905 gnd.n1182 585
R2505 gnd.n1899 gnd.n1203 585
R2506 gnd.n1203 gnd.n1190 585
R2507 gnd.n1901 gnd.n1900 585
R2508 gnd.n1902 gnd.n1901 585
R2509 gnd.n1204 gnd.n1202 585
R2510 gnd.n1211 gnd.n1202 585
R2511 gnd.n1894 gnd.n1893 585
R2512 gnd.n1893 gnd.n1892 585
R2513 gnd.n1207 gnd.n1206 585
R2514 gnd.n1873 gnd.n1207 585
R2515 gnd.n1869 gnd.n1868 585
R2516 gnd.n1870 gnd.n1869 585
R2517 gnd.n1225 gnd.n1224 585
R2518 gnd.n1231 gnd.n1224 585
R2519 gnd.n1864 gnd.n1863 585
R2520 gnd.n1863 gnd.n1862 585
R2521 gnd.n1228 gnd.n1227 585
R2522 gnd.n1852 gnd.n1228 585
R2523 gnd.n1834 gnd.n1833 585
R2524 gnd.n1835 gnd.n1834 585
R2525 gnd.n1356 gnd.n1355 585
R2526 gnd.n1817 gnd.n1355 585
R2527 gnd.n1829 gnd.n1828 585
R2528 gnd.n1828 gnd.n1341 585
R2529 gnd.n1827 gnd.n1358 585
R2530 gnd.n1827 gnd.n1340 585
R2531 gnd.n1826 gnd.n1360 585
R2532 gnd.n1826 gnd.n1825 585
R2533 gnd.n1778 gnd.n1359 585
R2534 gnd.n1804 gnd.n1359 585
R2535 gnd.n1780 gnd.n1779 585
R2536 gnd.n1779 gnd.n1368 585
R2537 gnd.n1781 gnd.n1387 585
R2538 gnd.n1387 gnd.n1376 585
R2539 gnd.n1783 gnd.n1782 585
R2540 gnd.n1784 gnd.n1783 585
R2541 gnd.n1388 gnd.n1386 585
R2542 gnd.n1395 gnd.n1386 585
R2543 gnd.n1770 gnd.n1769 585
R2544 gnd.n1769 gnd.n1768 585
R2545 gnd.n1391 gnd.n1390 585
R2546 gnd.n1758 gnd.n1391 585
R2547 gnd.n1745 gnd.n1415 585
R2548 gnd.n1415 gnd.n1414 585
R2549 gnd.n1747 gnd.n1746 585
R2550 gnd.n1748 gnd.n1747 585
R2551 gnd.n1416 gnd.n1413 585
R2552 gnd.n1423 gnd.n1413 585
R2553 gnd.n1740 gnd.n1739 585
R2554 gnd.n1739 gnd.n1738 585
R2555 gnd.n1419 gnd.n1418 585
R2556 gnd.n1727 gnd.n1419 585
R2557 gnd.n1714 gnd.n1440 585
R2558 gnd.n1440 gnd.n1439 585
R2559 gnd.n1716 gnd.n1715 585
R2560 gnd.n1717 gnd.n1716 585
R2561 gnd.n1710 gnd.n1438 585
R2562 gnd.n1709 gnd.n1708 585
R2563 gnd.n1443 gnd.n1442 585
R2564 gnd.n1706 gnd.n1443 585
R2565 gnd.n1465 gnd.n1464 585
R2566 gnd.n1468 gnd.n1467 585
R2567 gnd.n1466 gnd.n1461 585
R2568 gnd.n1473 gnd.n1472 585
R2569 gnd.n1475 gnd.n1474 585
R2570 gnd.n1478 gnd.n1477 585
R2571 gnd.n1476 gnd.n1459 585
R2572 gnd.n1483 gnd.n1482 585
R2573 gnd.n1485 gnd.n1484 585
R2574 gnd.n1488 gnd.n1487 585
R2575 gnd.n1486 gnd.n1457 585
R2576 gnd.n1493 gnd.n1492 585
R2577 gnd.n1497 gnd.n1494 585
R2578 gnd.n1498 gnd.n1435 585
R2579 gnd.n6681 gnd.n6680 585
R2580 gnd.n6674 gnd.n1014 585
R2581 gnd.n6676 gnd.n6675 585
R2582 gnd.n1017 gnd.n1016 585
R2583 gnd.n6646 gnd.n6645 585
R2584 gnd.n6648 gnd.n6647 585
R2585 gnd.n6650 gnd.n6649 585
R2586 gnd.n6652 gnd.n6651 585
R2587 gnd.n6654 gnd.n6653 585
R2588 gnd.n6656 gnd.n6655 585
R2589 gnd.n6658 gnd.n6657 585
R2590 gnd.n6660 gnd.n6659 585
R2591 gnd.n6662 gnd.n6661 585
R2592 gnd.n6665 gnd.n6664 585
R2593 gnd.n6663 gnd.n6635 585
R2594 gnd.n6669 gnd.n6632 585
R2595 gnd.n6671 gnd.n6670 585
R2596 gnd.n6672 gnd.n6671 585
R2597 gnd.n6683 gnd.n6682 585
R2598 gnd.n6682 gnd.n1004 585
R2599 gnd.n1010 gnd.n1002 585
R2600 gnd.n6689 gnd.n1002 585
R2601 gnd.n2344 gnd.n2343 585
R2602 gnd.n2345 gnd.n2344 585
R2603 gnd.n2338 gnd.n990 585
R2604 gnd.n6695 gnd.n990 585
R2605 gnd.n2337 gnd.n2336 585
R2606 gnd.n2336 gnd.n988 585
R2607 gnd.n2335 gnd.n2333 585
R2608 gnd.n2335 gnd.n979 585
R2609 gnd.n2075 gnd.n977 585
R2610 gnd.n6703 gnd.n977 585
R2611 gnd.n1114 gnd.n1113 585
R2612 gnd.n1113 gnd.n1112 585
R2613 gnd.n2069 gnd.n966 585
R2614 gnd.n6709 gnd.n966 585
R2615 gnd.n2068 gnd.n2067 585
R2616 gnd.n2067 gnd.n964 585
R2617 gnd.n2066 gnd.n1116 585
R2618 gnd.n2066 gnd.n955 585
R2619 gnd.n2065 gnd.n2064 585
R2620 gnd.n2065 gnd.n953 585
R2621 gnd.n1119 gnd.n1118 585
R2622 gnd.n2056 gnd.n1118 585
R2623 gnd.n1997 gnd.n1996 585
R2624 gnd.n1996 gnd.n1123 585
R2625 gnd.n1998 gnd.n1132 585
R2626 gnd.n2042 gnd.n1132 585
R2627 gnd.n1995 gnd.n1994 585
R2628 gnd.n1994 gnd.n1139 585
R2629 gnd.n1993 gnd.n1146 585
R2630 gnd.n1993 gnd.n1138 585
R2631 gnd.n1992 gnd.n1148 585
R2632 gnd.n1992 gnd.n1991 585
R2633 gnd.n1971 gnd.n1147 585
R2634 gnd.n1159 gnd.n1147 585
R2635 gnd.n1970 gnd.n1157 585
R2636 gnd.n1981 gnd.n1157 585
R2637 gnd.n1961 gnd.n1164 585
R2638 gnd.n1962 gnd.n1961 585
R2639 gnd.n1960 gnd.n1959 585
R2640 gnd.n1960 gnd.n1168 585
R2641 gnd.n1958 gnd.n1170 585
R2642 gnd.n1951 gnd.n1170 585
R2643 gnd.n1938 gnd.n1171 585
R2644 gnd.n1939 gnd.n1938 585
R2645 gnd.n1908 gnd.n1184 585
R2646 gnd.n1941 gnd.n1184 585
R2647 gnd.n1907 gnd.n1906 585
R2648 gnd.n1906 gnd.n1905 585
R2649 gnd.n1904 gnd.n1197 585
R2650 gnd.n1904 gnd.n1190 585
R2651 gnd.n1903 gnd.n1199 585
R2652 gnd.n1903 gnd.n1902 585
R2653 gnd.n1882 gnd.n1198 585
R2654 gnd.n1211 gnd.n1198 585
R2655 gnd.n1881 gnd.n1209 585
R2656 gnd.n1892 gnd.n1209 585
R2657 gnd.n1872 gnd.n1216 585
R2658 gnd.n1873 gnd.n1872 585
R2659 gnd.n1871 gnd.n1222 585
R2660 gnd.n1871 gnd.n1870 585
R2661 gnd.n1856 gnd.n1221 585
R2662 gnd.n1231 gnd.n1221 585
R2663 gnd.n1855 gnd.n1229 585
R2664 gnd.n1862 gnd.n1229 585
R2665 gnd.n1854 gnd.n1853 585
R2666 gnd.n1853 gnd.n1852 585
R2667 gnd.n1239 gnd.n1236 585
R2668 gnd.n1835 gnd.n1239 585
R2669 gnd.n1818 gnd.n1815 585
R2670 gnd.n1818 gnd.n1817 585
R2671 gnd.n1820 gnd.n1819 585
R2672 gnd.n1819 gnd.n1341 585
R2673 gnd.n1821 gnd.n1363 585
R2674 gnd.n1363 gnd.n1340 585
R2675 gnd.n1823 gnd.n1822 585
R2676 gnd.n1825 gnd.n1823 585
R2677 gnd.n1364 gnd.n1362 585
R2678 gnd.n1804 gnd.n1362 585
R2679 gnd.n1788 gnd.n1787 585
R2680 gnd.n1787 gnd.n1368 585
R2681 gnd.n1786 gnd.n1382 585
R2682 gnd.n1786 gnd.n1376 585
R2683 gnd.n1785 gnd.n1384 585
R2684 gnd.n1785 gnd.n1784 585
R2685 gnd.n1762 gnd.n1383 585
R2686 gnd.n1395 gnd.n1383 585
R2687 gnd.n1761 gnd.n1393 585
R2688 gnd.n1768 gnd.n1393 585
R2689 gnd.n1760 gnd.n1759 585
R2690 gnd.n1759 gnd.n1758 585
R2691 gnd.n1404 gnd.n1401 585
R2692 gnd.n1414 gnd.n1404 585
R2693 gnd.n1750 gnd.n1749 585
R2694 gnd.n1749 gnd.n1748 585
R2695 gnd.n1410 gnd.n1409 585
R2696 gnd.n1423 gnd.n1410 585
R2697 gnd.n1730 gnd.n1421 585
R2698 gnd.n1738 gnd.n1421 585
R2699 gnd.n1729 gnd.n1728 585
R2700 gnd.n1728 gnd.n1727 585
R2701 gnd.n1430 gnd.n1428 585
R2702 gnd.n1439 gnd.n1430 585
R2703 gnd.n1719 gnd.n1718 585
R2704 gnd.n1718 gnd.n1717 585
R2705 gnd.n5402 gnd.n3473 585
R2706 gnd.n3473 gnd.n3460 585
R2707 gnd.n5404 gnd.n5403 585
R2708 gnd.n5405 gnd.n5404 585
R2709 gnd.n3474 gnd.n3472 585
R2710 gnd.n3472 gnd.n3467 585
R2711 gnd.n5273 gnd.n5272 585
R2712 gnd.n5274 gnd.n5273 585
R2713 gnd.n5271 gnd.n3547 585
R2714 gnd.n3552 gnd.n3547 585
R2715 gnd.n5270 gnd.n5269 585
R2716 gnd.n5269 gnd.n5268 585
R2717 gnd.n3549 gnd.n3548 585
R2718 gnd.n5245 gnd.n3549 585
R2719 gnd.n5257 gnd.n5256 585
R2720 gnd.n5258 gnd.n5257 585
R2721 gnd.n5255 gnd.n3562 585
R2722 gnd.n5251 gnd.n3562 585
R2723 gnd.n5254 gnd.n5253 585
R2724 gnd.n5253 gnd.n5252 585
R2725 gnd.n3564 gnd.n3563 585
R2726 gnd.n5239 gnd.n3564 585
R2727 gnd.n5225 gnd.n5224 585
R2728 gnd.n5224 gnd.n3569 585
R2729 gnd.n5226 gnd.n3581 585
R2730 gnd.n3581 gnd.n3579 585
R2731 gnd.n5228 gnd.n5227 585
R2732 gnd.n5229 gnd.n5228 585
R2733 gnd.n5223 gnd.n3580 585
R2734 gnd.n3580 gnd.n3576 585
R2735 gnd.n5222 gnd.n5221 585
R2736 gnd.n5221 gnd.n5220 585
R2737 gnd.n3583 gnd.n3582 585
R2738 gnd.n3584 gnd.n3583 585
R2739 gnd.n5171 gnd.n3607 585
R2740 gnd.n5171 gnd.n5170 585
R2741 gnd.n5173 gnd.n5172 585
R2742 gnd.n5172 gnd.n3592 585
R2743 gnd.n5174 gnd.n3605 585
R2744 gnd.n5156 gnd.n3605 585
R2745 gnd.n5176 gnd.n5175 585
R2746 gnd.n5177 gnd.n5176 585
R2747 gnd.n3606 gnd.n3604 585
R2748 gnd.n3604 gnd.n3600 585
R2749 gnd.n5150 gnd.n5149 585
R2750 gnd.n5151 gnd.n5150 585
R2751 gnd.n5148 gnd.n3613 585
R2752 gnd.n3619 gnd.n3613 585
R2753 gnd.n5147 gnd.n5146 585
R2754 gnd.n5146 gnd.n5145 585
R2755 gnd.n3615 gnd.n3614 585
R2756 gnd.n3616 gnd.n3615 585
R2757 gnd.n5134 gnd.n5133 585
R2758 gnd.n5135 gnd.n5134 585
R2759 gnd.n5132 gnd.n3629 585
R2760 gnd.n3629 gnd.n3626 585
R2761 gnd.n5131 gnd.n5130 585
R2762 gnd.n5130 gnd.n5129 585
R2763 gnd.n3631 gnd.n3630 585
R2764 gnd.n3638 gnd.n3631 585
R2765 gnd.n5116 gnd.n5115 585
R2766 gnd.n5117 gnd.n5116 585
R2767 gnd.n5114 gnd.n3641 585
R2768 gnd.n3641 gnd.n3637 585
R2769 gnd.n5113 gnd.n5112 585
R2770 gnd.n5112 gnd.n5111 585
R2771 gnd.n3643 gnd.n3642 585
R2772 gnd.n3655 gnd.n3643 585
R2773 gnd.n5098 gnd.n5097 585
R2774 gnd.n5099 gnd.n5098 585
R2775 gnd.n5096 gnd.n3656 585
R2776 gnd.n3656 gnd.n3652 585
R2777 gnd.n5095 gnd.n5094 585
R2778 gnd.n5094 gnd.n5093 585
R2779 gnd.n3658 gnd.n3657 585
R2780 gnd.n5033 gnd.n3658 585
R2781 gnd.n3681 gnd.n3680 585
R2782 gnd.n3681 gnd.n3667 585
R2783 gnd.n5041 gnd.n5040 585
R2784 gnd.n5040 gnd.n5039 585
R2785 gnd.n5042 gnd.n3678 585
R2786 gnd.n3678 gnd.n3676 585
R2787 gnd.n5044 gnd.n5043 585
R2788 gnd.n5045 gnd.n5044 585
R2789 gnd.n3679 gnd.n3677 585
R2790 gnd.n5021 gnd.n3677 585
R2791 gnd.n3709 gnd.n3708 585
R2792 gnd.n3708 gnd.n3687 585
R2793 gnd.n3711 gnd.n3710 585
R2794 gnd.n4991 gnd.n3711 585
R2795 gnd.n4994 gnd.n3707 585
R2796 gnd.n4994 gnd.n4993 585
R2797 gnd.n4996 gnd.n4995 585
R2798 gnd.n4995 gnd.n3694 585
R2799 gnd.n4997 gnd.n3705 585
R2800 gnd.n4984 gnd.n3705 585
R2801 gnd.n4999 gnd.n4998 585
R2802 gnd.n5000 gnd.n4999 585
R2803 gnd.n3706 gnd.n3704 585
R2804 gnd.n3704 gnd.n3701 585
R2805 gnd.n4975 gnd.n4974 585
R2806 gnd.n4976 gnd.n4975 585
R2807 gnd.n4973 gnd.n3716 585
R2808 gnd.n3721 gnd.n3716 585
R2809 gnd.n4972 gnd.n4971 585
R2810 gnd.n4971 gnd.n4970 585
R2811 gnd.n3718 gnd.n3717 585
R2812 gnd.n4947 gnd.n3718 585
R2813 gnd.n4959 gnd.n4958 585
R2814 gnd.n4960 gnd.n4959 585
R2815 gnd.n4957 gnd.n3730 585
R2816 gnd.n3730 gnd.n3727 585
R2817 gnd.n4956 gnd.n4955 585
R2818 gnd.n4955 gnd.n4954 585
R2819 gnd.n3732 gnd.n3731 585
R2820 gnd.n3745 gnd.n3732 585
R2821 gnd.n4917 gnd.n4916 585
R2822 gnd.n4916 gnd.n3744 585
R2823 gnd.n4918 gnd.n3755 585
R2824 gnd.n4880 gnd.n3755 585
R2825 gnd.n4920 gnd.n4919 585
R2826 gnd.n4921 gnd.n4920 585
R2827 gnd.n4915 gnd.n3754 585
R2828 gnd.n3754 gnd.n3751 585
R2829 gnd.n4914 gnd.n4913 585
R2830 gnd.n4913 gnd.n4912 585
R2831 gnd.n3757 gnd.n3756 585
R2832 gnd.n3758 gnd.n3757 585
R2833 gnd.n4898 gnd.n4897 585
R2834 gnd.n4899 gnd.n4898 585
R2835 gnd.n4896 gnd.n3772 585
R2836 gnd.n3772 gnd.n3765 585
R2837 gnd.n4895 gnd.n4894 585
R2838 gnd.n4894 gnd.n4893 585
R2839 gnd.n3774 gnd.n3773 585
R2840 gnd.n3774 gnd.n2909 585
R2841 gnd.n4871 gnd.n4870 585
R2842 gnd.n4872 gnd.n4871 585
R2843 gnd.n2895 gnd.n2894 585
R2844 gnd.n2899 gnd.n2895 585
R2845 gnd.n6202 gnd.n6201 585
R2846 gnd.n6201 gnd.n6200 585
R2847 gnd.n6203 gnd.n2873 585
R2848 gnd.n3842 gnd.n2873 585
R2849 gnd.n6268 gnd.n6267 585
R2850 gnd.n6266 gnd.n2872 585
R2851 gnd.n6265 gnd.n2871 585
R2852 gnd.n6270 gnd.n2871 585
R2853 gnd.n6264 gnd.n6263 585
R2854 gnd.n6262 gnd.n6261 585
R2855 gnd.n6260 gnd.n6259 585
R2856 gnd.n6258 gnd.n6257 585
R2857 gnd.n6256 gnd.n6255 585
R2858 gnd.n6254 gnd.n6253 585
R2859 gnd.n6252 gnd.n6251 585
R2860 gnd.n6250 gnd.n6249 585
R2861 gnd.n6248 gnd.n6247 585
R2862 gnd.n6246 gnd.n6245 585
R2863 gnd.n6244 gnd.n6243 585
R2864 gnd.n6242 gnd.n6241 585
R2865 gnd.n6240 gnd.n6239 585
R2866 gnd.n6238 gnd.n6237 585
R2867 gnd.n6236 gnd.n6235 585
R2868 gnd.n6234 gnd.n6233 585
R2869 gnd.n6232 gnd.n6231 585
R2870 gnd.n6230 gnd.n6229 585
R2871 gnd.n6228 gnd.n6227 585
R2872 gnd.n6226 gnd.n6225 585
R2873 gnd.n6224 gnd.n6223 585
R2874 gnd.n6222 gnd.n6221 585
R2875 gnd.n6220 gnd.n6219 585
R2876 gnd.n6218 gnd.n6217 585
R2877 gnd.n6216 gnd.n6215 585
R2878 gnd.n6214 gnd.n6213 585
R2879 gnd.n6212 gnd.n6211 585
R2880 gnd.n6210 gnd.n6209 585
R2881 gnd.n6208 gnd.n2836 585
R2882 gnd.n6273 gnd.n6272 585
R2883 gnd.n2838 gnd.n2835 585
R2884 gnd.n3780 gnd.n3779 585
R2885 gnd.n3782 gnd.n3781 585
R2886 gnd.n3785 gnd.n3784 585
R2887 gnd.n3787 gnd.n3786 585
R2888 gnd.n3789 gnd.n3788 585
R2889 gnd.n3791 gnd.n3790 585
R2890 gnd.n3793 gnd.n3792 585
R2891 gnd.n3795 gnd.n3794 585
R2892 gnd.n3797 gnd.n3796 585
R2893 gnd.n3799 gnd.n3798 585
R2894 gnd.n3801 gnd.n3800 585
R2895 gnd.n3803 gnd.n3802 585
R2896 gnd.n3805 gnd.n3804 585
R2897 gnd.n3807 gnd.n3806 585
R2898 gnd.n3809 gnd.n3808 585
R2899 gnd.n3811 gnd.n3810 585
R2900 gnd.n3813 gnd.n3812 585
R2901 gnd.n3815 gnd.n3814 585
R2902 gnd.n3817 gnd.n3816 585
R2903 gnd.n3819 gnd.n3818 585
R2904 gnd.n3821 gnd.n3820 585
R2905 gnd.n3823 gnd.n3822 585
R2906 gnd.n3825 gnd.n3824 585
R2907 gnd.n3827 gnd.n3826 585
R2908 gnd.n3829 gnd.n3828 585
R2909 gnd.n3831 gnd.n3830 585
R2910 gnd.n3833 gnd.n3832 585
R2911 gnd.n3835 gnd.n3834 585
R2912 gnd.n3837 gnd.n3836 585
R2913 gnd.n3839 gnd.n3838 585
R2914 gnd.n3841 gnd.n3840 585
R2915 gnd.n5283 gnd.n5282 585
R2916 gnd.n5284 gnd.n3543 585
R2917 gnd.n5286 gnd.n5285 585
R2918 gnd.n5288 gnd.n3541 585
R2919 gnd.n5290 gnd.n5289 585
R2920 gnd.n5291 gnd.n3540 585
R2921 gnd.n5293 gnd.n5292 585
R2922 gnd.n5295 gnd.n3538 585
R2923 gnd.n5297 gnd.n5296 585
R2924 gnd.n5298 gnd.n3537 585
R2925 gnd.n5300 gnd.n5299 585
R2926 gnd.n5302 gnd.n3535 585
R2927 gnd.n5304 gnd.n5303 585
R2928 gnd.n5305 gnd.n3534 585
R2929 gnd.n5307 gnd.n5306 585
R2930 gnd.n5309 gnd.n3532 585
R2931 gnd.n5311 gnd.n5310 585
R2932 gnd.n5312 gnd.n3531 585
R2933 gnd.n5314 gnd.n5313 585
R2934 gnd.n5316 gnd.n3529 585
R2935 gnd.n5318 gnd.n5317 585
R2936 gnd.n5319 gnd.n3528 585
R2937 gnd.n5321 gnd.n5320 585
R2938 gnd.n5323 gnd.n3526 585
R2939 gnd.n5325 gnd.n5324 585
R2940 gnd.n5326 gnd.n3525 585
R2941 gnd.n5328 gnd.n5327 585
R2942 gnd.n5330 gnd.n3523 585
R2943 gnd.n5332 gnd.n5331 585
R2944 gnd.n5334 gnd.n3520 585
R2945 gnd.n5336 gnd.n5335 585
R2946 gnd.n5338 gnd.n3519 585
R2947 gnd.n5339 gnd.n3461 585
R2948 gnd.n5342 gnd.n3137 585
R2949 gnd.n5344 gnd.n5343 585
R2950 gnd.n5346 gnd.n3517 585
R2951 gnd.n5348 gnd.n5347 585
R2952 gnd.n5350 gnd.n3514 585
R2953 gnd.n5352 gnd.n5351 585
R2954 gnd.n5354 gnd.n3512 585
R2955 gnd.n5356 gnd.n5355 585
R2956 gnd.n5357 gnd.n3511 585
R2957 gnd.n5359 gnd.n5358 585
R2958 gnd.n5361 gnd.n3509 585
R2959 gnd.n5363 gnd.n5362 585
R2960 gnd.n5364 gnd.n3508 585
R2961 gnd.n5366 gnd.n5365 585
R2962 gnd.n5368 gnd.n3506 585
R2963 gnd.n5370 gnd.n5369 585
R2964 gnd.n5371 gnd.n3505 585
R2965 gnd.n5373 gnd.n5372 585
R2966 gnd.n5375 gnd.n3503 585
R2967 gnd.n5377 gnd.n5376 585
R2968 gnd.n5378 gnd.n3502 585
R2969 gnd.n5380 gnd.n5379 585
R2970 gnd.n5382 gnd.n3500 585
R2971 gnd.n5384 gnd.n5383 585
R2972 gnd.n5385 gnd.n3499 585
R2973 gnd.n5387 gnd.n5386 585
R2974 gnd.n5389 gnd.n3497 585
R2975 gnd.n5391 gnd.n5390 585
R2976 gnd.n5392 gnd.n3496 585
R2977 gnd.n5394 gnd.n5393 585
R2978 gnd.n5396 gnd.n3495 585
R2979 gnd.n5397 gnd.n3494 585
R2980 gnd.n5400 gnd.n5399 585
R2981 gnd.n5281 gnd.n5279 585
R2982 gnd.n5281 gnd.n3460 585
R2983 gnd.n5278 gnd.n3469 585
R2984 gnd.n5405 gnd.n3469 585
R2985 gnd.n5277 gnd.n5276 585
R2986 gnd.n5276 gnd.n3467 585
R2987 gnd.n5275 gnd.n3544 585
R2988 gnd.n5275 gnd.n5274 585
R2989 gnd.n5243 gnd.n3545 585
R2990 gnd.n3552 gnd.n3545 585
R2991 gnd.n5244 gnd.n3550 585
R2992 gnd.n5268 gnd.n3550 585
R2993 gnd.n5247 gnd.n5246 585
R2994 gnd.n5246 gnd.n5245 585
R2995 gnd.n5248 gnd.n3559 585
R2996 gnd.n5258 gnd.n3559 585
R2997 gnd.n5250 gnd.n5249 585
R2998 gnd.n5251 gnd.n5250 585
R2999 gnd.n5242 gnd.n3566 585
R3000 gnd.n5252 gnd.n3566 585
R3001 gnd.n5241 gnd.n5240 585
R3002 gnd.n5240 gnd.n5239 585
R3003 gnd.n3568 gnd.n3567 585
R3004 gnd.n3569 gnd.n3568 585
R3005 gnd.n5161 gnd.n5160 585
R3006 gnd.n5160 gnd.n3579 585
R3007 gnd.n5162 gnd.n3578 585
R3008 gnd.n5229 gnd.n3578 585
R3009 gnd.n5164 gnd.n5163 585
R3010 gnd.n5163 gnd.n3576 585
R3011 gnd.n5165 gnd.n3585 585
R3012 gnd.n5220 gnd.n3585 585
R3013 gnd.n5166 gnd.n3609 585
R3014 gnd.n3609 gnd.n3584 585
R3015 gnd.n5168 gnd.n5167 585
R3016 gnd.n5170 gnd.n5168 585
R3017 gnd.n5159 gnd.n3608 585
R3018 gnd.n3608 gnd.n3592 585
R3019 gnd.n5158 gnd.n5157 585
R3020 gnd.n5157 gnd.n5156 585
R3021 gnd.n5155 gnd.n3602 585
R3022 gnd.n5177 gnd.n3602 585
R3023 gnd.n5154 gnd.n5153 585
R3024 gnd.n5153 gnd.n3600 585
R3025 gnd.n5152 gnd.n3610 585
R3026 gnd.n5152 gnd.n5151 585
R3027 gnd.n5121 gnd.n3611 585
R3028 gnd.n3619 gnd.n3611 585
R3029 gnd.n5122 gnd.n3617 585
R3030 gnd.n5145 gnd.n3617 585
R3031 gnd.n5124 gnd.n5123 585
R3032 gnd.n5123 gnd.n3616 585
R3033 gnd.n5125 gnd.n3628 585
R3034 gnd.n5135 gnd.n3628 585
R3035 gnd.n5126 gnd.n3634 585
R3036 gnd.n3634 gnd.n3626 585
R3037 gnd.n5128 gnd.n5127 585
R3038 gnd.n5129 gnd.n5128 585
R3039 gnd.n5120 gnd.n3633 585
R3040 gnd.n3638 gnd.n3633 585
R3041 gnd.n5119 gnd.n5118 585
R3042 gnd.n5118 gnd.n5117 585
R3043 gnd.n3636 gnd.n3635 585
R3044 gnd.n3637 gnd.n3636 585
R3045 gnd.n5026 gnd.n3644 585
R3046 gnd.n5111 gnd.n3644 585
R3047 gnd.n5028 gnd.n5027 585
R3048 gnd.n5027 gnd.n3655 585
R3049 gnd.n5029 gnd.n3654 585
R3050 gnd.n5099 gnd.n3654 585
R3051 gnd.n5031 gnd.n5030 585
R3052 gnd.n5030 gnd.n3652 585
R3053 gnd.n5032 gnd.n3660 585
R3054 gnd.n5093 gnd.n3660 585
R3055 gnd.n5035 gnd.n5034 585
R3056 gnd.n5034 gnd.n5033 585
R3057 gnd.n5036 gnd.n3684 585
R3058 gnd.n3684 gnd.n3667 585
R3059 gnd.n5038 gnd.n5037 585
R3060 gnd.n5039 gnd.n5038 585
R3061 gnd.n5025 gnd.n3683 585
R3062 gnd.n3683 gnd.n3676 585
R3063 gnd.n5024 gnd.n3675 585
R3064 gnd.n5045 gnd.n3675 585
R3065 gnd.n5023 gnd.n5022 585
R3066 gnd.n5022 gnd.n5021 585
R3067 gnd.n3686 gnd.n3685 585
R3068 gnd.n3687 gnd.n3686 585
R3069 gnd.n4990 gnd.n4989 585
R3070 gnd.n4991 gnd.n4990 585
R3071 gnd.n4988 gnd.n3712 585
R3072 gnd.n4993 gnd.n3712 585
R3073 gnd.n4987 gnd.n4986 585
R3074 gnd.n4986 gnd.n3694 585
R3075 gnd.n4985 gnd.n4981 585
R3076 gnd.n4985 gnd.n4984 585
R3077 gnd.n4980 gnd.n3703 585
R3078 gnd.n5000 gnd.n3703 585
R3079 gnd.n4979 gnd.n4978 585
R3080 gnd.n4978 gnd.n3701 585
R3081 gnd.n4977 gnd.n3713 585
R3082 gnd.n4977 gnd.n4976 585
R3083 gnd.n3737 gnd.n3714 585
R3084 gnd.n3721 gnd.n3714 585
R3085 gnd.n3738 gnd.n3719 585
R3086 gnd.n4970 gnd.n3719 585
R3087 gnd.n4949 gnd.n4948 585
R3088 gnd.n4948 gnd.n4947 585
R3089 gnd.n4950 gnd.n3729 585
R3090 gnd.n4960 gnd.n3729 585
R3091 gnd.n4951 gnd.n3735 585
R3092 gnd.n3735 gnd.n3727 585
R3093 gnd.n4953 gnd.n4952 585
R3094 gnd.n4954 gnd.n4953 585
R3095 gnd.n3736 gnd.n3734 585
R3096 gnd.n3745 gnd.n3734 585
R3097 gnd.n4877 gnd.n4876 585
R3098 gnd.n4877 gnd.n3744 585
R3099 gnd.n4882 gnd.n4881 585
R3100 gnd.n4881 gnd.n4880 585
R3101 gnd.n4883 gnd.n3753 585
R3102 gnd.n4921 gnd.n3753 585
R3103 gnd.n4885 gnd.n4884 585
R3104 gnd.n4884 gnd.n3751 585
R3105 gnd.n4886 gnd.n3759 585
R3106 gnd.n4912 gnd.n3759 585
R3107 gnd.n4888 gnd.n4887 585
R3108 gnd.n4887 gnd.n3758 585
R3109 gnd.n4889 gnd.n3766 585
R3110 gnd.n4899 gnd.n3766 585
R3111 gnd.n4890 gnd.n3776 585
R3112 gnd.n3776 gnd.n3765 585
R3113 gnd.n4892 gnd.n4891 585
R3114 gnd.n4893 gnd.n4892 585
R3115 gnd.n4875 gnd.n3775 585
R3116 gnd.n3775 gnd.n2909 585
R3117 gnd.n4874 gnd.n4873 585
R3118 gnd.n4873 gnd.n4872 585
R3119 gnd.n3847 gnd.n3846 585
R3120 gnd.n3847 gnd.n2899 585
R3121 gnd.n3845 gnd.n2897 585
R3122 gnd.n6200 gnd.n2897 585
R3123 gnd.n3844 gnd.n3843 585
R3124 gnd.n3843 gnd.n3842 585
R3125 gnd.n6329 gnd.n2759 585
R3126 gnd.n4768 gnd.n2759 585
R3127 gnd.n6331 gnd.n6330 585
R3128 gnd.n6332 gnd.n6331 585
R3129 gnd.n2744 gnd.n2743 585
R3130 gnd.n4760 gnd.n2744 585
R3131 gnd.n6340 gnd.n6339 585
R3132 gnd.n6339 gnd.n6338 585
R3133 gnd.n6341 gnd.n2738 585
R3134 gnd.n4473 gnd.n2738 585
R3135 gnd.n6343 gnd.n6342 585
R3136 gnd.n6344 gnd.n6343 585
R3137 gnd.n2724 gnd.n2723 585
R3138 gnd.n4465 gnd.n2724 585
R3139 gnd.n6352 gnd.n6351 585
R3140 gnd.n6351 gnd.n6350 585
R3141 gnd.n6353 gnd.n2718 585
R3142 gnd.n4459 gnd.n2718 585
R3143 gnd.n6355 gnd.n6354 585
R3144 gnd.n6356 gnd.n6355 585
R3145 gnd.n2704 gnd.n2703 585
R3146 gnd.n4451 gnd.n2704 585
R3147 gnd.n6364 gnd.n6363 585
R3148 gnd.n6363 gnd.n6362 585
R3149 gnd.n6365 gnd.n2698 585
R3150 gnd.n4391 gnd.n2698 585
R3151 gnd.n6367 gnd.n6366 585
R3152 gnd.n6368 gnd.n6367 585
R3153 gnd.n2684 gnd.n2683 585
R3154 gnd.n4382 gnd.n2684 585
R3155 gnd.n6376 gnd.n6375 585
R3156 gnd.n6375 gnd.n6374 585
R3157 gnd.n6377 gnd.n2678 585
R3158 gnd.n4377 gnd.n2678 585
R3159 gnd.n6379 gnd.n6378 585
R3160 gnd.n6380 gnd.n6379 585
R3161 gnd.n2664 gnd.n2663 585
R3162 gnd.n4405 gnd.n2664 585
R3163 gnd.n6388 gnd.n6387 585
R3164 gnd.n6387 gnd.n6386 585
R3165 gnd.n6389 gnd.n2658 585
R3166 gnd.n4370 gnd.n2658 585
R3167 gnd.n6391 gnd.n6390 585
R3168 gnd.n6392 gnd.n6391 585
R3169 gnd.n2644 gnd.n2643 585
R3170 gnd.n4362 gnd.n2644 585
R3171 gnd.n6400 gnd.n6399 585
R3172 gnd.n6399 gnd.n6398 585
R3173 gnd.n6401 gnd.n2639 585
R3174 gnd.n4356 gnd.n2639 585
R3175 gnd.n6403 gnd.n6402 585
R3176 gnd.n6404 gnd.n6403 585
R3177 gnd.n2623 gnd.n2621 585
R3178 gnd.n4348 gnd.n2623 585
R3179 gnd.n6412 gnd.n6411 585
R3180 gnd.n6411 gnd.n6410 585
R3181 gnd.n2622 gnd.n2620 585
R3182 gnd.n4317 gnd.n2622 585
R3183 gnd.n4306 gnd.n4305 585
R3184 gnd.n4305 gnd.n3988 585
R3185 gnd.n4308 gnd.n4307 585
R3186 gnd.n4309 gnd.n4308 585
R3187 gnd.n4304 gnd.n4001 585
R3188 gnd.n4304 gnd.n4303 585
R3189 gnd.n4000 gnd.n3999 585
R3190 gnd.n4287 gnd.n3999 585
R3191 gnd.n4237 gnd.n4236 585
R3192 gnd.n4238 gnd.n4237 585
R3193 gnd.n2614 gnd.n2612 585
R3194 gnd.n4279 gnd.n2612 585
R3195 gnd.n6416 gnd.n6415 585
R3196 gnd.n6417 gnd.n6416 585
R3197 gnd.n2613 gnd.n2597 585
R3198 gnd.n4247 gnd.n2597 585
R3199 gnd.n6425 gnd.n6424 585
R3200 gnd.n6424 gnd.n6423 585
R3201 gnd.n6426 gnd.n2592 585
R3202 gnd.n4253 gnd.n2592 585
R3203 gnd.n6428 gnd.n6427 585
R3204 gnd.n6429 gnd.n6428 585
R3205 gnd.n2579 gnd.n2578 585
R3206 gnd.n4229 gnd.n2579 585
R3207 gnd.n6437 gnd.n6436 585
R3208 gnd.n6436 gnd.n6435 585
R3209 gnd.n6438 gnd.n2573 585
R3210 gnd.n4220 gnd.n2573 585
R3211 gnd.n6440 gnd.n6439 585
R3212 gnd.n6441 gnd.n6440 585
R3213 gnd.n2558 gnd.n2557 585
R3214 gnd.n4183 gnd.n2558 585
R3215 gnd.n6449 gnd.n6448 585
R3216 gnd.n6448 gnd.n6447 585
R3217 gnd.n6450 gnd.n2552 585
R3218 gnd.n4189 gnd.n2552 585
R3219 gnd.n6452 gnd.n6451 585
R3220 gnd.n6453 gnd.n6452 585
R3221 gnd.n2539 gnd.n2538 585
R3222 gnd.n4171 gnd.n2539 585
R3223 gnd.n6461 gnd.n6460 585
R3224 gnd.n6460 gnd.n6459 585
R3225 gnd.n6462 gnd.n2533 585
R3226 gnd.n2533 gnd.n2532 585
R3227 gnd.n6464 gnd.n6463 585
R3228 gnd.n6465 gnd.n6464 585
R3229 gnd.n2518 gnd.n2517 585
R3230 gnd.n2522 gnd.n2518 585
R3231 gnd.n6473 gnd.n6472 585
R3232 gnd.n6472 gnd.n6471 585
R3233 gnd.n6474 gnd.n2512 585
R3234 gnd.n2519 gnd.n2512 585
R3235 gnd.n6476 gnd.n6475 585
R3236 gnd.n6477 gnd.n6476 585
R3237 gnd.n2500 gnd.n2499 585
R3238 gnd.n2503 gnd.n2500 585
R3239 gnd.n6485 gnd.n6484 585
R3240 gnd.n6484 gnd.n6483 585
R3241 gnd.n6486 gnd.n2494 585
R3242 gnd.n2494 gnd.n2493 585
R3243 gnd.n6488 gnd.n6487 585
R3244 gnd.n6489 gnd.n6488 585
R3245 gnd.n2477 gnd.n2476 585
R3246 gnd.n2481 gnd.n2477 585
R3247 gnd.n6497 gnd.n6496 585
R3248 gnd.n6496 gnd.n6495 585
R3249 gnd.n6498 gnd.n2470 585
R3250 gnd.n2478 gnd.n2470 585
R3251 gnd.n6500 gnd.n6499 585
R3252 gnd.n6501 gnd.n6500 585
R3253 gnd.n2471 gnd.n2397 585
R3254 gnd.n2397 gnd.n2394 585
R3255 gnd.n6623 gnd.n6622 585
R3256 gnd.n6621 gnd.n2396 585
R3257 gnd.n6620 gnd.n2395 585
R3258 gnd.n6625 gnd.n2395 585
R3259 gnd.n6619 gnd.n6618 585
R3260 gnd.n6617 gnd.n6616 585
R3261 gnd.n6615 gnd.n6614 585
R3262 gnd.n6613 gnd.n6612 585
R3263 gnd.n6611 gnd.n6610 585
R3264 gnd.n6609 gnd.n6608 585
R3265 gnd.n6607 gnd.n6606 585
R3266 gnd.n6605 gnd.n6604 585
R3267 gnd.n6603 gnd.n6602 585
R3268 gnd.n6601 gnd.n6600 585
R3269 gnd.n6599 gnd.n6598 585
R3270 gnd.n6597 gnd.n6596 585
R3271 gnd.n6595 gnd.n6594 585
R3272 gnd.n6593 gnd.n6592 585
R3273 gnd.n6591 gnd.n6590 585
R3274 gnd.n6588 gnd.n6587 585
R3275 gnd.n6586 gnd.n6585 585
R3276 gnd.n6584 gnd.n6583 585
R3277 gnd.n6582 gnd.n6581 585
R3278 gnd.n6580 gnd.n6579 585
R3279 gnd.n6578 gnd.n6577 585
R3280 gnd.n6576 gnd.n6575 585
R3281 gnd.n6574 gnd.n6573 585
R3282 gnd.n6572 gnd.n6571 585
R3283 gnd.n6570 gnd.n6569 585
R3284 gnd.n6568 gnd.n6567 585
R3285 gnd.n6566 gnd.n6565 585
R3286 gnd.n6564 gnd.n6563 585
R3287 gnd.n6562 gnd.n6561 585
R3288 gnd.n6560 gnd.n6559 585
R3289 gnd.n6558 gnd.n6557 585
R3290 gnd.n6556 gnd.n6555 585
R3291 gnd.n6554 gnd.n6553 585
R3292 gnd.n6552 gnd.n6551 585
R3293 gnd.n6550 gnd.n6549 585
R3294 gnd.n6548 gnd.n6547 585
R3295 gnd.n6546 gnd.n6545 585
R3296 gnd.n6544 gnd.n6543 585
R3297 gnd.n6542 gnd.n6541 585
R3298 gnd.n6540 gnd.n6539 585
R3299 gnd.n6538 gnd.n6537 585
R3300 gnd.n6536 gnd.n6535 585
R3301 gnd.n6534 gnd.n6533 585
R3302 gnd.n6532 gnd.n6531 585
R3303 gnd.n6530 gnd.n6529 585
R3304 gnd.n6528 gnd.n6527 585
R3305 gnd.n6526 gnd.n6525 585
R3306 gnd.n6524 gnd.n6523 585
R3307 gnd.n6522 gnd.n6521 585
R3308 gnd.n6520 gnd.n6519 585
R3309 gnd.n6518 gnd.n6517 585
R3310 gnd.n6516 gnd.n6515 585
R3311 gnd.n6514 gnd.n6513 585
R3312 gnd.n6512 gnd.n6511 585
R3313 gnd.n6510 gnd.n6509 585
R3314 gnd.n2466 gnd.n2459 585
R3315 gnd.n4752 gnd.n4751 585
R3316 gnd.n4750 gnd.n4661 585
R3317 gnd.n4749 gnd.n4748 585
R3318 gnd.n4742 gnd.n4662 585
R3319 gnd.n4744 gnd.n4743 585
R3320 gnd.n4741 gnd.n4740 585
R3321 gnd.n4739 gnd.n4738 585
R3322 gnd.n4732 gnd.n4664 585
R3323 gnd.n4734 gnd.n4733 585
R3324 gnd.n4731 gnd.n4730 585
R3325 gnd.n4729 gnd.n4728 585
R3326 gnd.n4722 gnd.n4666 585
R3327 gnd.n4724 gnd.n4723 585
R3328 gnd.n4721 gnd.n4720 585
R3329 gnd.n4719 gnd.n4718 585
R3330 gnd.n4712 gnd.n4668 585
R3331 gnd.n4714 gnd.n4713 585
R3332 gnd.n4711 gnd.n4710 585
R3333 gnd.n4709 gnd.n4708 585
R3334 gnd.n4702 gnd.n4670 585
R3335 gnd.n4704 gnd.n4703 585
R3336 gnd.n4701 gnd.n4674 585
R3337 gnd.n4700 gnd.n4699 585
R3338 gnd.n4693 gnd.n4675 585
R3339 gnd.n4695 gnd.n4694 585
R3340 gnd.n4692 gnd.n4691 585
R3341 gnd.n4690 gnd.n4689 585
R3342 gnd.n4683 gnd.n4677 585
R3343 gnd.n4685 gnd.n4684 585
R3344 gnd.n4682 gnd.n4681 585
R3345 gnd.n4680 gnd.n2832 585
R3346 gnd.n6276 gnd.n6275 585
R3347 gnd.n6278 gnd.n6277 585
R3348 gnd.n6280 gnd.n6279 585
R3349 gnd.n6282 gnd.n6281 585
R3350 gnd.n6284 gnd.n6283 585
R3351 gnd.n6286 gnd.n6285 585
R3352 gnd.n6288 gnd.n6287 585
R3353 gnd.n6290 gnd.n6289 585
R3354 gnd.n6293 gnd.n6292 585
R3355 gnd.n6295 gnd.n6294 585
R3356 gnd.n6297 gnd.n6296 585
R3357 gnd.n6299 gnd.n6298 585
R3358 gnd.n6301 gnd.n6300 585
R3359 gnd.n6303 gnd.n6302 585
R3360 gnd.n6305 gnd.n6304 585
R3361 gnd.n6307 gnd.n6306 585
R3362 gnd.n6309 gnd.n6308 585
R3363 gnd.n6311 gnd.n6310 585
R3364 gnd.n6313 gnd.n6312 585
R3365 gnd.n6315 gnd.n6314 585
R3366 gnd.n6317 gnd.n6316 585
R3367 gnd.n6319 gnd.n6318 585
R3368 gnd.n6320 gnd.n2805 585
R3369 gnd.n6322 gnd.n6321 585
R3370 gnd.n2764 gnd.n2763 585
R3371 gnd.n6326 gnd.n6325 585
R3372 gnd.n6325 gnd.n6324 585
R3373 gnd.n4756 gnd.n3935 585
R3374 gnd.n4768 gnd.n3935 585
R3375 gnd.n4757 gnd.n2756 585
R3376 gnd.n6332 gnd.n2756 585
R3377 gnd.n4759 gnd.n4758 585
R3378 gnd.n4760 gnd.n4759 585
R3379 gnd.n4476 gnd.n2746 585
R3380 gnd.n6338 gnd.n2746 585
R3381 gnd.n4475 gnd.n4474 585
R3382 gnd.n4474 gnd.n4473 585
R3383 gnd.n3940 gnd.n2735 585
R3384 gnd.n6344 gnd.n2735 585
R3385 gnd.n4464 gnd.n4463 585
R3386 gnd.n4465 gnd.n4464 585
R3387 gnd.n4462 gnd.n2726 585
R3388 gnd.n6350 gnd.n2726 585
R3389 gnd.n4461 gnd.n4460 585
R3390 gnd.n4460 gnd.n4459 585
R3391 gnd.n3946 gnd.n2715 585
R3392 gnd.n6356 gnd.n2715 585
R3393 gnd.n4387 gnd.n3951 585
R3394 gnd.n4451 gnd.n3951 585
R3395 gnd.n4388 gnd.n2706 585
R3396 gnd.n6362 gnd.n2706 585
R3397 gnd.n4390 gnd.n4389 585
R3398 gnd.n4391 gnd.n4390 585
R3399 gnd.n4385 gnd.n2695 585
R3400 gnd.n6368 gnd.n2695 585
R3401 gnd.n4384 gnd.n4383 585
R3402 gnd.n4383 gnd.n4382 585
R3403 gnd.n4380 gnd.n2686 585
R3404 gnd.n6374 gnd.n2686 585
R3405 gnd.n4379 gnd.n4378 585
R3406 gnd.n4378 gnd.n4377 585
R3407 gnd.n4375 gnd.n2675 585
R3408 gnd.n6380 gnd.n2675 585
R3409 gnd.n4374 gnd.n3963 585
R3410 gnd.n4405 gnd.n3963 585
R3411 gnd.n4373 gnd.n2666 585
R3412 gnd.n6386 gnd.n2666 585
R3413 gnd.n4372 gnd.n4371 585
R3414 gnd.n4371 gnd.n4370 585
R3415 gnd.n3971 gnd.n2655 585
R3416 gnd.n6392 gnd.n2655 585
R3417 gnd.n4361 gnd.n4360 585
R3418 gnd.n4362 gnd.n4361 585
R3419 gnd.n4359 gnd.n2646 585
R3420 gnd.n6398 gnd.n2646 585
R3421 gnd.n4358 gnd.n4357 585
R3422 gnd.n4357 gnd.n4356 585
R3423 gnd.n3977 gnd.n2636 585
R3424 gnd.n6404 gnd.n2636 585
R3425 gnd.n4292 gnd.n3982 585
R3426 gnd.n4348 gnd.n3982 585
R3427 gnd.n4293 gnd.n2625 585
R3428 gnd.n6410 gnd.n2625 585
R3429 gnd.n4294 gnd.n3989 585
R3430 gnd.n4317 gnd.n3989 585
R3431 gnd.n4296 gnd.n4295 585
R3432 gnd.n4295 gnd.n3988 585
R3433 gnd.n4291 gnd.n3996 585
R3434 gnd.n4309 gnd.n3996 585
R3435 gnd.n4290 gnd.n4003 585
R3436 gnd.n4303 gnd.n4003 585
R3437 gnd.n4289 gnd.n4288 585
R3438 gnd.n4288 gnd.n4287 585
R3439 gnd.n4011 gnd.n4009 585
R3440 gnd.n4238 gnd.n4011 585
R3441 gnd.n4243 gnd.n4017 585
R3442 gnd.n4279 gnd.n4017 585
R3443 gnd.n4244 gnd.n2609 585
R3444 gnd.n6417 gnd.n2609 585
R3445 gnd.n4246 gnd.n4245 585
R3446 gnd.n4247 gnd.n4246 585
R3447 gnd.n4235 gnd.n2599 585
R3448 gnd.n6423 gnd.n2599 585
R3449 gnd.n4234 gnd.n4026 585
R3450 gnd.n4253 gnd.n4026 585
R3451 gnd.n4232 gnd.n2590 585
R3452 gnd.n6429 gnd.n2590 585
R3453 gnd.n4231 gnd.n4230 585
R3454 gnd.n4230 gnd.n4229 585
R3455 gnd.n4031 gnd.n2580 585
R3456 gnd.n6435 gnd.n2580 585
R3457 gnd.n4179 gnd.n4035 585
R3458 gnd.n4220 gnd.n4035 585
R3459 gnd.n4180 gnd.n2570 585
R3460 gnd.n6441 gnd.n2570 585
R3461 gnd.n4182 gnd.n4181 585
R3462 gnd.n4183 gnd.n4182 585
R3463 gnd.n4177 gnd.n2560 585
R3464 gnd.n6447 gnd.n2560 585
R3465 gnd.n4176 gnd.n4040 585
R3466 gnd.n4189 gnd.n4040 585
R3467 gnd.n4174 gnd.n2550 585
R3468 gnd.n6453 gnd.n2550 585
R3469 gnd.n4173 gnd.n4172 585
R3470 gnd.n4172 gnd.n4171 585
R3471 gnd.n4068 gnd.n2540 585
R3472 gnd.n6459 gnd.n2540 585
R3473 gnd.n4067 gnd.n4066 585
R3474 gnd.n4066 gnd.n2532 585
R3475 gnd.n4064 gnd.n2530 585
R3476 gnd.n6465 gnd.n2530 585
R3477 gnd.n4063 gnd.n4062 585
R3478 gnd.n4062 gnd.n2522 585
R3479 gnd.n4061 gnd.n2520 585
R3480 gnd.n6471 gnd.n2520 585
R3481 gnd.n4060 gnd.n4059 585
R3482 gnd.n4059 gnd.n2519 585
R3483 gnd.n4057 gnd.n2510 585
R3484 gnd.n6477 gnd.n2510 585
R3485 gnd.n4056 gnd.n4055 585
R3486 gnd.n4055 gnd.n2503 585
R3487 gnd.n4054 gnd.n2501 585
R3488 gnd.n6483 gnd.n2501 585
R3489 gnd.n4053 gnd.n4052 585
R3490 gnd.n4052 gnd.n2493 585
R3491 gnd.n4050 gnd.n2491 585
R3492 gnd.n6489 gnd.n2491 585
R3493 gnd.n4049 gnd.n4048 585
R3494 gnd.n4048 gnd.n2481 585
R3495 gnd.n4047 gnd.n2479 585
R3496 gnd.n6495 gnd.n2479 585
R3497 gnd.n4046 gnd.n2467 585
R3498 gnd.n2478 gnd.n2467 585
R3499 gnd.n6502 gnd.n2465 585
R3500 gnd.n6502 gnd.n6501 585
R3501 gnd.n6504 gnd.n6503 585
R3502 gnd.n6503 gnd.n2394 585
R3503 gnd.n7858 gnd.n250 585
R3504 gnd.n250 gnd.n249 585
R3505 gnd.n7860 gnd.n7859 585
R3506 gnd.n7861 gnd.n7860 585
R3507 gnd.n237 gnd.n236 585
R3508 gnd.n240 gnd.n237 585
R3509 gnd.n7869 gnd.n7868 585
R3510 gnd.n7868 gnd.n7867 585
R3511 gnd.n7870 gnd.n231 585
R3512 gnd.n231 gnd.n230 585
R3513 gnd.n7872 gnd.n7871 585
R3514 gnd.n7873 gnd.n7872 585
R3515 gnd.n218 gnd.n217 585
R3516 gnd.n227 gnd.n218 585
R3517 gnd.n7881 gnd.n7880 585
R3518 gnd.n7880 gnd.n7879 585
R3519 gnd.n7882 gnd.n212 585
R3520 gnd.n212 gnd.n211 585
R3521 gnd.n7884 gnd.n7883 585
R3522 gnd.n7885 gnd.n7884 585
R3523 gnd.n198 gnd.n197 585
R3524 gnd.n202 gnd.n198 585
R3525 gnd.n7893 gnd.n7892 585
R3526 gnd.n7892 gnd.n7891 585
R3527 gnd.n7894 gnd.n192 585
R3528 gnd.n199 gnd.n192 585
R3529 gnd.n7896 gnd.n7895 585
R3530 gnd.n7897 gnd.n7896 585
R3531 gnd.n178 gnd.n177 585
R3532 gnd.n188 gnd.n178 585
R3533 gnd.n7905 gnd.n7904 585
R3534 gnd.n7904 gnd.n7903 585
R3535 gnd.n7906 gnd.n172 585
R3536 gnd.n7701 gnd.n172 585
R3537 gnd.n7908 gnd.n7907 585
R3538 gnd.n7909 gnd.n7908 585
R3539 gnd.n158 gnd.n157 585
R3540 gnd.n7596 gnd.n158 585
R3541 gnd.n7917 gnd.n7916 585
R3542 gnd.n7916 gnd.n7915 585
R3543 gnd.n7918 gnd.n152 585
R3544 gnd.n5765 gnd.n152 585
R3545 gnd.n7920 gnd.n7919 585
R3546 gnd.n7921 gnd.n7920 585
R3547 gnd.n138 gnd.n137 585
R3548 gnd.n5771 gnd.n138 585
R3549 gnd.n7929 gnd.n7928 585
R3550 gnd.n7928 gnd.n7927 585
R3551 gnd.n7930 gnd.n133 585
R3552 gnd.n5777 gnd.n133 585
R3553 gnd.n7932 gnd.n7931 585
R3554 gnd.n7933 gnd.n7932 585
R3555 gnd.n117 gnd.n115 585
R3556 gnd.n5783 gnd.n117 585
R3557 gnd.n7941 gnd.n7940 585
R3558 gnd.n7940 gnd.n7939 585
R3559 gnd.n116 gnd.n108 585
R3560 gnd.n5722 gnd.n116 585
R3561 gnd.n7944 gnd.n106 585
R3562 gnd.n5795 gnd.n106 585
R3563 gnd.n7946 gnd.n7945 585
R3564 gnd.n7947 gnd.n7946 585
R3565 gnd.n3336 gnd.n105 585
R3566 gnd.n5801 gnd.n105 585
R3567 gnd.n3338 gnd.n3337 585
R3568 gnd.n3350 gnd.n3338 585
R3569 gnd.n5809 gnd.n5808 585
R3570 gnd.n5808 gnd.n5807 585
R3571 gnd.n5811 gnd.n5810 585
R3572 gnd.n5812 gnd.n5811 585
R3573 gnd.n3335 gnd.n3334 585
R3574 gnd.n3335 gnd.n3328 585
R3575 gnd.n3333 gnd.n3318 585
R3576 gnd.n3321 gnd.n3318 585
R3577 gnd.n5823 gnd.n5822 585
R3578 gnd.n5822 gnd.n5821 585
R3579 gnd.n5825 gnd.n5824 585
R3580 gnd.n5826 gnd.n5825 585
R3581 gnd.n3303 gnd.n3302 585
R3582 gnd.n5681 gnd.n3303 585
R3583 gnd.n5834 gnd.n5833 585
R3584 gnd.n5833 gnd.n5832 585
R3585 gnd.n5835 gnd.n3296 585
R3586 gnd.n5661 gnd.n3296 585
R3587 gnd.n5837 gnd.n5836 585
R3588 gnd.n5838 gnd.n5837 585
R3589 gnd.n3282 gnd.n3281 585
R3590 gnd.n5654 gnd.n3282 585
R3591 gnd.n5846 gnd.n5845 585
R3592 gnd.n5845 gnd.n5844 585
R3593 gnd.n5847 gnd.n3276 585
R3594 gnd.n5646 gnd.n3276 585
R3595 gnd.n5849 gnd.n5848 585
R3596 gnd.n5850 gnd.n5849 585
R3597 gnd.n3261 gnd.n3260 585
R3598 gnd.n5639 gnd.n3261 585
R3599 gnd.n5858 gnd.n5857 585
R3600 gnd.n5857 gnd.n5856 585
R3601 gnd.n5859 gnd.n3255 585
R3602 gnd.n5631 gnd.n3255 585
R3603 gnd.n5861 gnd.n5860 585
R3604 gnd.n5862 gnd.n5861 585
R3605 gnd.n3241 gnd.n3240 585
R3606 gnd.n5624 gnd.n3241 585
R3607 gnd.n5870 gnd.n5869 585
R3608 gnd.n5869 gnd.n5868 585
R3609 gnd.n5871 gnd.n3235 585
R3610 gnd.n5616 gnd.n3235 585
R3611 gnd.n5873 gnd.n5872 585
R3612 gnd.n5874 gnd.n5873 585
R3613 gnd.n3220 gnd.n3219 585
R3614 gnd.n5609 gnd.n3220 585
R3615 gnd.n5882 gnd.n5881 585
R3616 gnd.n5881 gnd.n5880 585
R3617 gnd.n5883 gnd.n3214 585
R3618 gnd.n5601 gnd.n3214 585
R3619 gnd.n5885 gnd.n5884 585
R3620 gnd.n5886 gnd.n5885 585
R3621 gnd.n3196 gnd.n3195 585
R3622 gnd.n5594 gnd.n3196 585
R3623 gnd.n5894 gnd.n5893 585
R3624 gnd.n5893 gnd.n5892 585
R3625 gnd.n5895 gnd.n3187 585
R3626 gnd.n5586 gnd.n3187 585
R3627 gnd.n5897 gnd.n5896 585
R3628 gnd.n5898 gnd.n5897 585
R3629 gnd.n3188 gnd.n3186 585
R3630 gnd.n5562 gnd.n3186 585
R3631 gnd.n3189 gnd.n3108 585
R3632 gnd.n5906 gnd.n3108 585
R3633 gnd.n6025 gnd.n6024 585
R3634 gnd.n6023 gnd.n3107 585
R3635 gnd.n6022 gnd.n3106 585
R3636 gnd.n6027 gnd.n3106 585
R3637 gnd.n6021 gnd.n6020 585
R3638 gnd.n6019 gnd.n6018 585
R3639 gnd.n6017 gnd.n6016 585
R3640 gnd.n6015 gnd.n6014 585
R3641 gnd.n6013 gnd.n6012 585
R3642 gnd.n6011 gnd.n6010 585
R3643 gnd.n6009 gnd.n6008 585
R3644 gnd.n6007 gnd.n6006 585
R3645 gnd.n6005 gnd.n6004 585
R3646 gnd.n6003 gnd.n6002 585
R3647 gnd.n6001 gnd.n6000 585
R3648 gnd.n5999 gnd.n5998 585
R3649 gnd.n5997 gnd.n5996 585
R3650 gnd.n5995 gnd.n5994 585
R3651 gnd.n5993 gnd.n5992 585
R3652 gnd.n5990 gnd.n5989 585
R3653 gnd.n5988 gnd.n5987 585
R3654 gnd.n5986 gnd.n5985 585
R3655 gnd.n5984 gnd.n5983 585
R3656 gnd.n5982 gnd.n5981 585
R3657 gnd.n5980 gnd.n5979 585
R3658 gnd.n5978 gnd.n5977 585
R3659 gnd.n5976 gnd.n5975 585
R3660 gnd.n5973 gnd.n5972 585
R3661 gnd.n5971 gnd.n5970 585
R3662 gnd.n5969 gnd.n5968 585
R3663 gnd.n5967 gnd.n5966 585
R3664 gnd.n5965 gnd.n5964 585
R3665 gnd.n5963 gnd.n5962 585
R3666 gnd.n5961 gnd.n5960 585
R3667 gnd.n5959 gnd.n5958 585
R3668 gnd.n5957 gnd.n5956 585
R3669 gnd.n5955 gnd.n5954 585
R3670 gnd.n5953 gnd.n5952 585
R3671 gnd.n5951 gnd.n5950 585
R3672 gnd.n5949 gnd.n5948 585
R3673 gnd.n5947 gnd.n5946 585
R3674 gnd.n5945 gnd.n5944 585
R3675 gnd.n5943 gnd.n5942 585
R3676 gnd.n5941 gnd.n5940 585
R3677 gnd.n5939 gnd.n5938 585
R3678 gnd.n5937 gnd.n5936 585
R3679 gnd.n5935 gnd.n5934 585
R3680 gnd.n5933 gnd.n5932 585
R3681 gnd.n5931 gnd.n5930 585
R3682 gnd.n5929 gnd.n5928 585
R3683 gnd.n5927 gnd.n5926 585
R3684 gnd.n5925 gnd.n5924 585
R3685 gnd.n5923 gnd.n5922 585
R3686 gnd.n5921 gnd.n5920 585
R3687 gnd.n5919 gnd.n5918 585
R3688 gnd.n5917 gnd.n5916 585
R3689 gnd.n5915 gnd.n5914 585
R3690 gnd.n5909 gnd.n5908 585
R3691 gnd.n7729 gnd.n351 585
R3692 gnd.n7737 gnd.n7736 585
R3693 gnd.n7739 gnd.n7738 585
R3694 gnd.n7741 gnd.n7740 585
R3695 gnd.n7743 gnd.n7742 585
R3696 gnd.n7745 gnd.n7744 585
R3697 gnd.n7747 gnd.n7746 585
R3698 gnd.n7749 gnd.n7748 585
R3699 gnd.n7751 gnd.n7750 585
R3700 gnd.n7753 gnd.n7752 585
R3701 gnd.n7755 gnd.n7754 585
R3702 gnd.n7757 gnd.n7756 585
R3703 gnd.n7759 gnd.n7758 585
R3704 gnd.n7761 gnd.n7760 585
R3705 gnd.n7763 gnd.n7762 585
R3706 gnd.n7765 gnd.n7764 585
R3707 gnd.n7767 gnd.n7766 585
R3708 gnd.n7769 gnd.n7768 585
R3709 gnd.n7771 gnd.n7770 585
R3710 gnd.n7774 gnd.n7773 585
R3711 gnd.n7772 gnd.n331 585
R3712 gnd.n7779 gnd.n7778 585
R3713 gnd.n7781 gnd.n7780 585
R3714 gnd.n7783 gnd.n7782 585
R3715 gnd.n7785 gnd.n7784 585
R3716 gnd.n7787 gnd.n7786 585
R3717 gnd.n7789 gnd.n7788 585
R3718 gnd.n7791 gnd.n7790 585
R3719 gnd.n7793 gnd.n7792 585
R3720 gnd.n7795 gnd.n7794 585
R3721 gnd.n7797 gnd.n7796 585
R3722 gnd.n7799 gnd.n7798 585
R3723 gnd.n7801 gnd.n7800 585
R3724 gnd.n7803 gnd.n7802 585
R3725 gnd.n7805 gnd.n7804 585
R3726 gnd.n7807 gnd.n7806 585
R3727 gnd.n7809 gnd.n7808 585
R3728 gnd.n7811 gnd.n7810 585
R3729 gnd.n7813 gnd.n7812 585
R3730 gnd.n7815 gnd.n7814 585
R3731 gnd.n7817 gnd.n7816 585
R3732 gnd.n7822 gnd.n7821 585
R3733 gnd.n7824 gnd.n7823 585
R3734 gnd.n7826 gnd.n7825 585
R3735 gnd.n7828 gnd.n7827 585
R3736 gnd.n7830 gnd.n7829 585
R3737 gnd.n7832 gnd.n7831 585
R3738 gnd.n7834 gnd.n7833 585
R3739 gnd.n7836 gnd.n7835 585
R3740 gnd.n7838 gnd.n7837 585
R3741 gnd.n7840 gnd.n7839 585
R3742 gnd.n7842 gnd.n7841 585
R3743 gnd.n7844 gnd.n7843 585
R3744 gnd.n7846 gnd.n7845 585
R3745 gnd.n7848 gnd.n7847 585
R3746 gnd.n7849 gnd.n295 585
R3747 gnd.n7851 gnd.n7850 585
R3748 gnd.n255 gnd.n254 585
R3749 gnd.n7855 gnd.n7854 585
R3750 gnd.n7854 gnd.n7853 585
R3751 gnd.n7731 gnd.n7730 585
R3752 gnd.n7730 gnd.n249 585
R3753 gnd.n7728 gnd.n247 585
R3754 gnd.n7861 gnd.n247 585
R3755 gnd.n7727 gnd.n7726 585
R3756 gnd.n7726 gnd.n240 585
R3757 gnd.n7725 gnd.n238 585
R3758 gnd.n7867 gnd.n238 585
R3759 gnd.n7724 gnd.n7723 585
R3760 gnd.n7723 gnd.n230 585
R3761 gnd.n7721 gnd.n228 585
R3762 gnd.n7873 gnd.n228 585
R3763 gnd.n7720 gnd.n7719 585
R3764 gnd.n7719 gnd.n227 585
R3765 gnd.n7718 gnd.n219 585
R3766 gnd.n7879 gnd.n219 585
R3767 gnd.n7717 gnd.n7716 585
R3768 gnd.n7716 gnd.n211 585
R3769 gnd.n7714 gnd.n209 585
R3770 gnd.n7885 gnd.n209 585
R3771 gnd.n7713 gnd.n7712 585
R3772 gnd.n7712 gnd.n202 585
R3773 gnd.n7711 gnd.n200 585
R3774 gnd.n7891 gnd.n200 585
R3775 gnd.n7710 gnd.n7709 585
R3776 gnd.n7709 gnd.n199 585
R3777 gnd.n7707 gnd.n189 585
R3778 gnd.n7897 gnd.n189 585
R3779 gnd.n7706 gnd.n7705 585
R3780 gnd.n7705 gnd.n188 585
R3781 gnd.n7704 gnd.n180 585
R3782 gnd.n7903 gnd.n180 585
R3783 gnd.n7703 gnd.n7702 585
R3784 gnd.n7702 gnd.n7701 585
R3785 gnd.n355 gnd.n169 585
R3786 gnd.n7909 gnd.n169 585
R3787 gnd.n5761 gnd.n360 585
R3788 gnd.n7596 gnd.n360 585
R3789 gnd.n5762 gnd.n160 585
R3790 gnd.n7915 gnd.n160 585
R3791 gnd.n5764 gnd.n5763 585
R3792 gnd.n5765 gnd.n5764 585
R3793 gnd.n5735 gnd.n149 585
R3794 gnd.n7921 gnd.n149 585
R3795 gnd.n5773 gnd.n5772 585
R3796 gnd.n5772 gnd.n5771 585
R3797 gnd.n5774 gnd.n140 585
R3798 gnd.n7927 gnd.n140 585
R3799 gnd.n5776 gnd.n5775 585
R3800 gnd.n5777 gnd.n5776 585
R3801 gnd.n5733 gnd.n130 585
R3802 gnd.n7933 gnd.n130 585
R3803 gnd.n5732 gnd.n5719 585
R3804 gnd.n5783 gnd.n5719 585
R3805 gnd.n5731 gnd.n119 585
R3806 gnd.n7939 gnd.n119 585
R3807 gnd.n5703 gnd.n5702 585
R3808 gnd.n5722 gnd.n5703 585
R3809 gnd.n5797 gnd.n5796 585
R3810 gnd.n5796 gnd.n5795 585
R3811 gnd.n5798 gnd.n102 585
R3812 gnd.n7947 gnd.n102 585
R3813 gnd.n5800 gnd.n5799 585
R3814 gnd.n5801 gnd.n5800 585
R3815 gnd.n5698 gnd.n3351 585
R3816 gnd.n3351 gnd.n3350 585
R3817 gnd.n5697 gnd.n3339 585
R3818 gnd.n5807 gnd.n3339 585
R3819 gnd.n5696 gnd.n3329 585
R3820 gnd.n5812 gnd.n3329 585
R3821 gnd.n5686 gnd.n3352 585
R3822 gnd.n5686 gnd.n3328 585
R3823 gnd.n5688 gnd.n5687 585
R3824 gnd.n5687 gnd.n3321 585
R3825 gnd.n5685 gnd.n3319 585
R3826 gnd.n5821 gnd.n3319 585
R3827 gnd.n5684 gnd.n3315 585
R3828 gnd.n5826 gnd.n3315 585
R3829 gnd.n5683 gnd.n5682 585
R3830 gnd.n5682 gnd.n5681 585
R3831 gnd.n3354 gnd.n3305 585
R3832 gnd.n5832 gnd.n3305 585
R3833 gnd.n5660 gnd.n5659 585
R3834 gnd.n5661 gnd.n5660 585
R3835 gnd.n5657 gnd.n3293 585
R3836 gnd.n5838 gnd.n3293 585
R3837 gnd.n5656 gnd.n5655 585
R3838 gnd.n5655 gnd.n5654 585
R3839 gnd.n3359 gnd.n3284 585
R3840 gnd.n5844 gnd.n3284 585
R3841 gnd.n5645 gnd.n5644 585
R3842 gnd.n5646 gnd.n5645 585
R3843 gnd.n5642 gnd.n3273 585
R3844 gnd.n5850 gnd.n3273 585
R3845 gnd.n5641 gnd.n5640 585
R3846 gnd.n5640 gnd.n5639 585
R3847 gnd.n3364 gnd.n3263 585
R3848 gnd.n5856 gnd.n3263 585
R3849 gnd.n5630 gnd.n5629 585
R3850 gnd.n5631 gnd.n5630 585
R3851 gnd.n5627 gnd.n3252 585
R3852 gnd.n5862 gnd.n3252 585
R3853 gnd.n5626 gnd.n5625 585
R3854 gnd.n5625 gnd.n5624 585
R3855 gnd.n3368 gnd.n3243 585
R3856 gnd.n5868 gnd.n3243 585
R3857 gnd.n5615 gnd.n5614 585
R3858 gnd.n5616 gnd.n5615 585
R3859 gnd.n5612 gnd.n3232 585
R3860 gnd.n5874 gnd.n3232 585
R3861 gnd.n5611 gnd.n5610 585
R3862 gnd.n5610 gnd.n5609 585
R3863 gnd.n3373 gnd.n3222 585
R3864 gnd.n5880 gnd.n3222 585
R3865 gnd.n5600 gnd.n5599 585
R3866 gnd.n5601 gnd.n5600 585
R3867 gnd.n5597 gnd.n3211 585
R3868 gnd.n5886 gnd.n3211 585
R3869 gnd.n5596 gnd.n5595 585
R3870 gnd.n5595 gnd.n5594 585
R3871 gnd.n3377 gnd.n3198 585
R3872 gnd.n5892 gnd.n3198 585
R3873 gnd.n3182 gnd.n3181 585
R3874 gnd.n5586 gnd.n3182 585
R3875 gnd.n5900 gnd.n5899 585
R3876 gnd.n5899 gnd.n5898 585
R3877 gnd.n5901 gnd.n3171 585
R3878 gnd.n5562 gnd.n3171 585
R3879 gnd.n5907 gnd.n3172 585
R3880 gnd.n5907 gnd.n5906 585
R3881 gnd.n4197 gnd.n4195 585
R3882 gnd.n4195 gnd.n2529 585
R3883 gnd.n7587 gnd.n7586 585
R3884 gnd.n7587 gnd.n191 585
R3885 gnd.n7589 gnd.n367 585
R3886 gnd.n7589 gnd.n7588 585
R3887 gnd.n7591 gnd.n7590 585
R3888 gnd.n7590 gnd.n179 585
R3889 gnd.n7592 gnd.n362 585
R3890 gnd.n362 gnd.n171 585
R3891 gnd.n7594 gnd.n7593 585
R3892 gnd.n7595 gnd.n7594 585
R3893 gnd.n363 gnd.n361 585
R3894 gnd.n361 gnd.n162 585
R3895 gnd.n5749 gnd.n5748 585
R3896 gnd.n5749 gnd.n159 585
R3897 gnd.n5751 gnd.n5750 585
R3898 gnd.n5750 gnd.n151 585
R3899 gnd.n5752 gnd.n5737 585
R3900 gnd.n5737 gnd.n148 585
R3901 gnd.n5754 gnd.n5753 585
R3902 gnd.n5755 gnd.n5754 585
R3903 gnd.n5738 gnd.n5736 585
R3904 gnd.n5736 gnd.n139 585
R3905 gnd.n5740 gnd.n5718 585
R3906 gnd.n5718 gnd.n132 585
R3907 gnd.n5785 gnd.n5717 585
R3908 gnd.n5785 gnd.n5784 585
R3909 gnd.n5787 gnd.n5786 585
R3910 gnd.n5786 gnd.n121 585
R3911 gnd.n5788 gnd.n5705 585
R3912 gnd.n5705 gnd.n118 585
R3913 gnd.n5791 gnd.n5790 585
R3914 gnd.n5792 gnd.n5791 585
R3915 gnd.n5715 gnd.n5704 585
R3916 gnd.n5704 gnd.n103 585
R3917 gnd.n5713 gnd.n5712 585
R3918 gnd.n5712 gnd.n101 585
R3919 gnd.n5711 gnd.n5706 585
R3920 gnd.n5711 gnd.n3348 585
R3921 gnd.n5710 gnd.n5709 585
R3922 gnd.n5710 gnd.n3341 585
R3923 gnd.n5707 gnd.n3326 585
R3924 gnd.n3331 gnd.n3326 585
R3925 gnd.n5815 gnd.n5814 585
R3926 gnd.n5814 gnd.n5813 585
R3927 gnd.n5816 gnd.n3323 585
R3928 gnd.n3327 gnd.n3323 585
R3929 gnd.n5819 gnd.n5818 585
R3930 gnd.n5820 gnd.n5819 585
R3931 gnd.n3324 gnd.n3322 585
R3932 gnd.n3322 gnd.n3317 585
R3933 gnd.n5527 gnd.n5526 585
R3934 gnd.n5526 gnd.n3314 585
R3935 gnd.n5528 gnd.n5520 585
R3936 gnd.n5520 gnd.n3307 585
R3937 gnd.n5530 gnd.n5529 585
R3938 gnd.n5530 gnd.n3304 585
R3939 gnd.n5531 gnd.n5519 585
R3940 gnd.n5531 gnd.n3295 585
R3941 gnd.n5533 gnd.n5532 585
R3942 gnd.n5532 gnd.n3292 585
R3943 gnd.n5534 gnd.n5514 585
R3944 gnd.n5514 gnd.n3360 585
R3945 gnd.n5536 gnd.n5535 585
R3946 gnd.n5536 gnd.n3283 585
R3947 gnd.n5537 gnd.n5513 585
R3948 gnd.n5537 gnd.n3275 585
R3949 gnd.n5539 gnd.n5538 585
R3950 gnd.n5538 gnd.n3272 585
R3951 gnd.n5540 gnd.n5508 585
R3952 gnd.n5508 gnd.n3265 585
R3953 gnd.n5542 gnd.n5541 585
R3954 gnd.n5542 gnd.n3262 585
R3955 gnd.n5543 gnd.n5507 585
R3956 gnd.n5543 gnd.n3254 585
R3957 gnd.n5545 gnd.n5544 585
R3958 gnd.n5544 gnd.n3251 585
R3959 gnd.n5546 gnd.n5502 585
R3960 gnd.n5502 gnd.n3369 585
R3961 gnd.n5548 gnd.n5547 585
R3962 gnd.n5548 gnd.n3242 585
R3963 gnd.n5549 gnd.n5501 585
R3964 gnd.n5549 gnd.n3234 585
R3965 gnd.n5551 gnd.n5550 585
R3966 gnd.n5550 gnd.n3231 585
R3967 gnd.n5552 gnd.n5496 585
R3968 gnd.n5496 gnd.n3224 585
R3969 gnd.n5554 gnd.n5553 585
R3970 gnd.n5554 gnd.n3221 585
R3971 gnd.n5555 gnd.n5495 585
R3972 gnd.n5555 gnd.n3213 585
R3973 gnd.n5557 gnd.n5556 585
R3974 gnd.n5556 gnd.n3210 585
R3975 gnd.n5558 gnd.n5490 585
R3976 gnd.n5490 gnd.n3200 585
R3977 gnd.n5560 gnd.n5559 585
R3978 gnd.n5560 gnd.n3197 585
R3979 gnd.n5561 gnd.n5489 585
R3980 gnd.n5561 gnd.n3184 585
R3981 gnd.n5565 gnd.n5564 585
R3982 gnd.n5564 gnd.n5563 585
R3983 gnd.n5566 gnd.n5484 585
R3984 gnd.n5484 gnd.n3175 585
R3985 gnd.n5568 gnd.n5567 585
R3986 gnd.n5568 gnd.n3173 585
R3987 gnd.n5569 gnd.n5483 585
R3988 gnd.n5569 gnd.n3105 585
R3989 gnd.n5571 gnd.n5570 585
R3990 gnd.n5570 gnd.n3063 585
R3991 gnd.n5572 gnd.n3410 585
R3992 gnd.n3410 gnd.n3408 585
R3993 gnd.n5574 gnd.n5573 585
R3994 gnd.n5575 gnd.n5574 585
R3995 gnd.n3411 gnd.n3409 585
R3996 gnd.n3409 gnd.n2996 585
R3997 gnd.n5477 gnd.n2995 585
R3998 gnd.n6095 gnd.n2995 585
R3999 gnd.n5476 gnd.n5475 585
R4000 gnd.n5475 gnd.n2994 585
R4001 gnd.n5474 gnd.n3413 585
R4002 gnd.n5474 gnd.n5473 585
R4003 gnd.n5462 gnd.n3414 585
R4004 gnd.n3415 gnd.n3414 585
R4005 gnd.n5464 gnd.n5463 585
R4006 gnd.n5465 gnd.n5464 585
R4007 gnd.n3424 gnd.n3423 585
R4008 gnd.n3423 gnd.n3422 585
R4009 gnd.n5456 gnd.n5455 585
R4010 gnd.n5455 gnd.n5454 585
R4011 gnd.n3427 gnd.n3426 585
R4012 gnd.n3435 gnd.n3427 585
R4013 gnd.n5445 gnd.n5444 585
R4014 gnd.n5446 gnd.n5445 585
R4015 gnd.n3437 gnd.n3436 585
R4016 gnd.n3436 gnd.n3434 585
R4017 gnd.n5440 gnd.n5439 585
R4018 gnd.n5439 gnd.n5438 585
R4019 gnd.n3440 gnd.n3439 585
R4020 gnd.n3448 gnd.n3440 585
R4021 gnd.n5429 gnd.n5428 585
R4022 gnd.n5430 gnd.n5429 585
R4023 gnd.n3450 gnd.n3449 585
R4024 gnd.n3449 gnd.n3447 585
R4025 gnd.n5424 gnd.n5423 585
R4026 gnd.n5423 gnd.n5422 585
R4027 gnd.n3453 gnd.n3452 585
R4028 gnd.n3454 gnd.n3453 585
R4029 gnd.n5413 gnd.n5412 585
R4030 gnd.n5414 gnd.n5413 585
R4031 gnd.n3463 gnd.n3462 585
R4032 gnd.n3471 gnd.n3462 585
R4033 gnd.n5408 gnd.n5407 585
R4034 gnd.n5407 gnd.n5406 585
R4035 gnd.n3466 gnd.n3465 585
R4036 gnd.n3546 gnd.n3466 585
R4037 gnd.n5266 gnd.n5265 585
R4038 gnd.n5267 gnd.n5266 585
R4039 gnd.n3554 gnd.n3553 585
R4040 gnd.n3561 gnd.n3553 585
R4041 gnd.n5261 gnd.n5260 585
R4042 gnd.n5260 gnd.n5259 585
R4043 gnd.n3557 gnd.n3556 585
R4044 gnd.n3565 gnd.n3557 585
R4045 gnd.n5237 gnd.n5236 585
R4046 gnd.n5238 gnd.n5237 585
R4047 gnd.n3572 gnd.n3571 585
R4048 gnd.n5195 gnd.n3571 585
R4049 gnd.n5232 gnd.n5231 585
R4050 gnd.n5231 gnd.n5230 585
R4051 gnd.n3575 gnd.n3574 585
R4052 gnd.n5219 gnd.n3575 585
R4053 gnd.n5185 gnd.n3595 585
R4054 gnd.n5169 gnd.n3595 585
R4055 gnd.n5187 gnd.n5186 585
R4056 gnd.n5188 gnd.n5187 585
R4057 gnd.n3596 gnd.n3594 585
R4058 gnd.n3603 gnd.n3594 585
R4059 gnd.n5180 gnd.n5179 585
R4060 gnd.n5179 gnd.n5178 585
R4061 gnd.n3599 gnd.n3598 585
R4062 gnd.n3612 gnd.n3599 585
R4063 gnd.n5143 gnd.n5142 585
R4064 gnd.n5144 gnd.n5143 585
R4065 gnd.n3622 gnd.n3621 585
R4066 gnd.n5069 gnd.n3621 585
R4067 gnd.n5138 gnd.n5137 585
R4068 gnd.n5137 gnd.n5136 585
R4069 gnd.n3625 gnd.n3624 585
R4070 gnd.n3632 gnd.n3625 585
R4071 gnd.n5107 gnd.n3647 585
R4072 gnd.n3647 gnd.n3640 585
R4073 gnd.n5109 gnd.n5108 585
R4074 gnd.n5110 gnd.n5109 585
R4075 gnd.n3648 gnd.n3646 585
R4076 gnd.n5063 gnd.n3646 585
R4077 gnd.n5102 gnd.n5101 585
R4078 gnd.n5101 gnd.n5100 585
R4079 gnd.n3651 gnd.n3650 585
R4080 gnd.n5092 gnd.n3651 585
R4081 gnd.n5054 gnd.n3669 585
R4082 gnd.n3669 gnd.n3659 585
R4083 gnd.n5056 gnd.n5055 585
R4084 gnd.n5057 gnd.n5056 585
R4085 gnd.n3670 gnd.n3668 585
R4086 gnd.n3682 gnd.n3668 585
R4087 gnd.n5049 gnd.n5048 585
R4088 gnd.n5048 gnd.n5047 585
R4089 gnd.n3673 gnd.n3672 585
R4090 gnd.n5020 gnd.n3673 585
R4091 gnd.n5008 gnd.n3696 585
R4092 gnd.n4992 gnd.n3696 585
R4093 gnd.n5010 gnd.n5009 585
R4094 gnd.n5011 gnd.n5010 585
R4095 gnd.n3697 gnd.n3695 585
R4096 gnd.n4983 gnd.n3695 585
R4097 gnd.n5003 gnd.n5002 585
R4098 gnd.n5002 gnd.n5001 585
R4099 gnd.n3700 gnd.n3699 585
R4100 gnd.n3715 gnd.n3700 585
R4101 gnd.n4968 gnd.n4967 585
R4102 gnd.n4969 gnd.n4968 585
R4103 gnd.n3723 gnd.n3722 585
R4104 gnd.n4946 gnd.n3722 585
R4105 gnd.n4963 gnd.n4962 585
R4106 gnd.n4962 gnd.n4961 585
R4107 gnd.n3726 gnd.n3725 585
R4108 gnd.n3733 gnd.n3726 585
R4109 gnd.n4929 gnd.n4928 585
R4110 gnd.n4930 gnd.n4929 585
R4111 gnd.n3747 gnd.n3746 585
R4112 gnd.n4879 gnd.n3746 585
R4113 gnd.n4924 gnd.n4923 585
R4114 gnd.n4923 gnd.n4922 585
R4115 gnd.n3750 gnd.n3749 585
R4116 gnd.n4911 gnd.n3750 585
R4117 gnd.n3770 gnd.n3769 585
R4118 gnd.n3771 gnd.n3770 585
R4119 gnd.n2908 gnd.n2907 585
R4120 gnd.n4900 gnd.n2908 585
R4121 gnd.n6195 gnd.n6194 585
R4122 gnd.n6194 gnd.n6193 585
R4123 gnd.n6196 gnd.n2902 585
R4124 gnd.n4869 gnd.n2902 585
R4125 gnd.n6198 gnd.n6197 585
R4126 gnd.n6199 gnd.n6198 585
R4127 gnd.n2903 gnd.n2901 585
R4128 gnd.n2901 gnd.n2896 585
R4129 gnd.n4856 gnd.n3856 585
R4130 gnd.n3856 gnd.n2870 585
R4131 gnd.n4858 gnd.n4857 585
R4132 gnd.n4859 gnd.n4858 585
R4133 gnd.n3857 gnd.n3855 585
R4134 gnd.n3855 gnd.n3853 585
R4135 gnd.n4850 gnd.n4849 585
R4136 gnd.n4849 gnd.n4848 585
R4137 gnd.n3860 gnd.n3859 585
R4138 gnd.n3861 gnd.n3860 585
R4139 gnd.n4828 gnd.n4827 585
R4140 gnd.n4829 gnd.n4828 585
R4141 gnd.n3872 gnd.n3871 585
R4142 gnd.n3878 gnd.n3871 585
R4143 gnd.n4823 gnd.n4822 585
R4144 gnd.n4822 gnd.n4821 585
R4145 gnd.n3875 gnd.n3874 585
R4146 gnd.n3876 gnd.n3875 585
R4147 gnd.n4812 gnd.n4811 585
R4148 gnd.n4813 gnd.n4812 585
R4149 gnd.n3886 gnd.n3885 585
R4150 gnd.n3892 gnd.n3885 585
R4151 gnd.n4807 gnd.n4806 585
R4152 gnd.n4806 gnd.n4805 585
R4153 gnd.n3889 gnd.n3888 585
R4154 gnd.n3890 gnd.n3889 585
R4155 gnd.n4796 gnd.n4795 585
R4156 gnd.n4797 gnd.n4796 585
R4157 gnd.n3901 gnd.n3900 585
R4158 gnd.n3900 gnd.n3898 585
R4159 gnd.n4791 gnd.n4790 585
R4160 gnd.n4790 gnd.n4789 585
R4161 gnd.n3904 gnd.n3903 585
R4162 gnd.n3905 gnd.n3904 585
R4163 gnd.n4778 gnd.n3929 585
R4164 gnd.n3929 gnd.n3927 585
R4165 gnd.n4780 gnd.n4779 585
R4166 gnd.n4781 gnd.n4780 585
R4167 gnd.n3930 gnd.n3928 585
R4168 gnd.n3928 gnd.n3912 585
R4169 gnd.n4773 gnd.n4772 585
R4170 gnd.n4772 gnd.n2776 585
R4171 gnd.n4771 gnd.n3932 585
R4172 gnd.n4771 gnd.n2765 585
R4173 gnd.n4770 gnd.n3934 585
R4174 gnd.n4770 gnd.n4769 585
R4175 gnd.n4435 gnd.n3933 585
R4176 gnd.n3933 gnd.n2758 585
R4177 gnd.n4437 gnd.n4436 585
R4178 gnd.n4437 gnd.n2755 585
R4179 gnd.n4438 gnd.n4430 585
R4180 gnd.n4438 gnd.n2748 585
R4181 gnd.n4440 gnd.n4439 585
R4182 gnd.n4439 gnd.n2745 585
R4183 gnd.n4441 gnd.n4425 585
R4184 gnd.n4425 gnd.n2737 585
R4185 gnd.n4443 gnd.n4442 585
R4186 gnd.n4443 gnd.n2734 585
R4187 gnd.n4444 gnd.n4424 585
R4188 gnd.n4444 gnd.n3945 585
R4189 gnd.n4446 gnd.n4445 585
R4190 gnd.n4445 gnd.n2725 585
R4191 gnd.n4447 gnd.n3953 585
R4192 gnd.n3953 gnd.n2717 585
R4193 gnd.n4449 gnd.n4448 585
R4194 gnd.n4450 gnd.n4449 585
R4195 gnd.n3954 gnd.n3952 585
R4196 gnd.n3952 gnd.n2708 585
R4197 gnd.n4418 gnd.n4417 585
R4198 gnd.n4417 gnd.n2705 585
R4199 gnd.n4416 gnd.n3956 585
R4200 gnd.n4416 gnd.n2697 585
R4201 gnd.n4415 gnd.n4414 585
R4202 gnd.n4415 gnd.n2694 585
R4203 gnd.n3958 gnd.n3957 585
R4204 gnd.n4381 gnd.n3957 585
R4205 gnd.n4410 gnd.n4409 585
R4206 gnd.n4409 gnd.n2685 585
R4207 gnd.n4408 gnd.n3960 585
R4208 gnd.n4408 gnd.n2677 585
R4209 gnd.n4407 gnd.n3962 585
R4210 gnd.n4407 gnd.n4406 585
R4211 gnd.n4335 gnd.n3961 585
R4212 gnd.n3961 gnd.n2668 585
R4213 gnd.n4337 gnd.n4336 585
R4214 gnd.n4336 gnd.n2665 585
R4215 gnd.n4338 gnd.n4328 585
R4216 gnd.n4328 gnd.n2657 585
R4217 gnd.n4340 gnd.n4339 585
R4218 gnd.n4340 gnd.n2654 585
R4219 gnd.n4341 gnd.n4327 585
R4220 gnd.n4341 gnd.n3976 585
R4221 gnd.n4343 gnd.n4342 585
R4222 gnd.n4342 gnd.n2645 585
R4223 gnd.n4344 gnd.n3984 585
R4224 gnd.n3984 gnd.n2638 585
R4225 gnd.n4346 gnd.n4345 585
R4226 gnd.n4347 gnd.n4346 585
R4227 gnd.n4322 gnd.n3983 585
R4228 gnd.n3983 gnd.n2627 585
R4229 gnd.n4321 gnd.n4320 585
R4230 gnd.n4320 gnd.n2624 585
R4231 gnd.n4319 gnd.n3987 585
R4232 gnd.n4319 gnd.n4318 585
R4233 gnd.n4268 gnd.n3986 585
R4234 gnd.n3997 gnd.n3986 585
R4235 gnd.n4271 gnd.n4270 585
R4236 gnd.n4271 gnd.n3995 585
R4237 gnd.n4273 gnd.n4272 585
R4238 gnd.n4272 gnd.n4002 585
R4239 gnd.n4275 gnd.n4019 585
R4240 gnd.n4019 gnd.n4012 585
R4241 gnd.n4277 gnd.n4276 585
R4242 gnd.n4278 gnd.n4277 585
R4243 gnd.n4266 gnd.n4018 585
R4244 gnd.n4018 gnd.n2611 585
R4245 gnd.n4265 gnd.n4264 585
R4246 gnd.n4264 gnd.n2608 585
R4247 gnd.n4263 gnd.n4262 585
R4248 gnd.n4263 gnd.n2601 585
R4249 gnd.n4261 gnd.n4021 585
R4250 gnd.n4021 gnd.n2598 585
R4251 gnd.n4255 gnd.n4022 585
R4252 gnd.n4255 gnd.n4254 585
R4253 gnd.n4257 gnd.n4256 585
R4254 gnd.n4256 gnd.n2589 585
R4255 gnd.n4025 gnd.n4024 585
R4256 gnd.n4025 gnd.n2582 585
R4257 gnd.n4218 gnd.n4217 585
R4258 gnd.n4219 gnd.n4218 585
R4259 gnd.n4037 gnd.n4036 585
R4260 gnd.n4036 gnd.n2572 585
R4261 gnd.n4213 gnd.n4212 585
R4262 gnd.n4212 gnd.n2569 585
R4263 gnd.n4211 gnd.n4039 585
R4264 gnd.n4211 gnd.n2562 585
R4265 gnd.n4210 gnd.n4209 585
R4266 gnd.n4210 gnd.n2559 585
R4267 gnd.n4192 gnd.n4191 585
R4268 gnd.n4191 gnd.n4190 585
R4269 gnd.n4205 gnd.n4204 585
R4270 gnd.n4204 gnd.n2549 585
R4271 gnd.n4203 gnd.n4194 585
R4272 gnd.n4203 gnd.n2542 585
R4273 gnd.n4202 gnd.n4200 585
R4274 gnd.n4202 gnd.n4201 585
R4275 gnd.n6094 gnd.n6093 585
R4276 gnd.n6095 gnd.n6094 585
R4277 gnd.n2999 gnd.n2997 585
R4278 gnd.n2997 gnd.n2994 585
R4279 gnd.n5472 gnd.n5471 585
R4280 gnd.n5473 gnd.n5472 585
R4281 gnd.n3417 gnd.n3416 585
R4282 gnd.n3416 gnd.n3415 585
R4283 gnd.n5467 gnd.n5466 585
R4284 gnd.n5466 gnd.n5465 585
R4285 gnd.n3420 gnd.n3419 585
R4286 gnd.n3422 gnd.n3420 585
R4287 gnd.n5453 gnd.n5452 585
R4288 gnd.n5454 gnd.n5453 585
R4289 gnd.n3429 gnd.n3428 585
R4290 gnd.n3435 gnd.n3428 585
R4291 gnd.n5448 gnd.n5447 585
R4292 gnd.n5447 gnd.n5446 585
R4293 gnd.n3432 gnd.n3431 585
R4294 gnd.n3434 gnd.n3432 585
R4295 gnd.n5437 gnd.n5436 585
R4296 gnd.n5438 gnd.n5437 585
R4297 gnd.n3442 gnd.n3441 585
R4298 gnd.n3448 gnd.n3441 585
R4299 gnd.n5432 gnd.n5431 585
R4300 gnd.n5431 gnd.n5430 585
R4301 gnd.n3445 gnd.n3444 585
R4302 gnd.n3447 gnd.n3445 585
R4303 gnd.n5421 gnd.n5420 585
R4304 gnd.n5422 gnd.n5421 585
R4305 gnd.n3456 gnd.n3455 585
R4306 gnd.n3455 gnd.n3454 585
R4307 gnd.n5416 gnd.n5415 585
R4308 gnd.n5415 gnd.n5414 585
R4309 gnd.n3459 gnd.n3458 585
R4310 gnd.n3471 gnd.n3459 585
R4311 gnd.n5202 gnd.n3468 585
R4312 gnd.n5406 gnd.n3468 585
R4313 gnd.n5205 gnd.n5201 585
R4314 gnd.n5201 gnd.n3546 585
R4315 gnd.n5206 gnd.n3551 585
R4316 gnd.n5267 gnd.n3551 585
R4317 gnd.n5207 gnd.n5200 585
R4318 gnd.n5200 gnd.n3561 585
R4319 gnd.n5198 gnd.n3558 585
R4320 gnd.n5259 gnd.n3558 585
R4321 gnd.n5211 gnd.n5197 585
R4322 gnd.n5197 gnd.n3565 585
R4323 gnd.n5212 gnd.n3570 585
R4324 gnd.n5238 gnd.n3570 585
R4325 gnd.n5213 gnd.n5196 585
R4326 gnd.n5196 gnd.n5195 585
R4327 gnd.n3588 gnd.n3577 585
R4328 gnd.n5230 gnd.n3577 585
R4329 gnd.n5218 gnd.n5217 585
R4330 gnd.n5219 gnd.n5218 585
R4331 gnd.n3587 gnd.n3586 585
R4332 gnd.n5169 gnd.n3586 585
R4333 gnd.n5190 gnd.n5189 585
R4334 gnd.n5189 gnd.n5188 585
R4335 gnd.n3591 gnd.n3590 585
R4336 gnd.n3603 gnd.n3591 585
R4337 gnd.n5073 gnd.n3601 585
R4338 gnd.n5178 gnd.n3601 585
R4339 gnd.n5072 gnd.n5071 585
R4340 gnd.n5071 gnd.n3612 585
R4341 gnd.n5077 gnd.n3618 585
R4342 gnd.n5144 gnd.n3618 585
R4343 gnd.n5078 gnd.n5070 585
R4344 gnd.n5070 gnd.n5069 585
R4345 gnd.n5079 gnd.n3627 585
R4346 gnd.n5136 gnd.n3627 585
R4347 gnd.n5067 gnd.n5066 585
R4348 gnd.n5066 gnd.n3632 585
R4349 gnd.n5083 gnd.n5065 585
R4350 gnd.n5065 gnd.n3640 585
R4351 gnd.n5084 gnd.n3645 585
R4352 gnd.n5110 gnd.n3645 585
R4353 gnd.n5085 gnd.n5064 585
R4354 gnd.n5064 gnd.n5063 585
R4355 gnd.n3663 gnd.n3653 585
R4356 gnd.n5100 gnd.n3653 585
R4357 gnd.n5090 gnd.n5089 585
R4358 gnd.n5092 gnd.n5090 585
R4359 gnd.n3662 gnd.n3661 585
R4360 gnd.n3661 gnd.n3659 585
R4361 gnd.n5059 gnd.n5058 585
R4362 gnd.n5058 gnd.n5057 585
R4363 gnd.n3666 gnd.n3665 585
R4364 gnd.n3682 gnd.n3666 585
R4365 gnd.n3690 gnd.n3674 585
R4366 gnd.n5047 gnd.n3674 585
R4367 gnd.n5019 gnd.n5018 585
R4368 gnd.n5020 gnd.n5019 585
R4369 gnd.n3689 gnd.n3688 585
R4370 gnd.n4992 gnd.n3688 585
R4371 gnd.n5013 gnd.n5012 585
R4372 gnd.n5012 gnd.n5011 585
R4373 gnd.n3693 gnd.n3692 585
R4374 gnd.n4983 gnd.n3693 585
R4375 gnd.n4938 gnd.n3702 585
R4376 gnd.n5001 gnd.n3702 585
R4377 gnd.n4939 gnd.n4937 585
R4378 gnd.n4937 gnd.n3715 585
R4379 gnd.n3740 gnd.n3720 585
R4380 gnd.n4969 gnd.n3720 585
R4381 gnd.n4944 gnd.n4943 585
R4382 gnd.n4946 gnd.n4944 585
R4383 gnd.n3739 gnd.n3728 585
R4384 gnd.n4961 gnd.n3728 585
R4385 gnd.n4933 gnd.n4932 585
R4386 gnd.n4932 gnd.n3733 585
R4387 gnd.n4931 gnd.n3742 585
R4388 gnd.n4931 gnd.n4930 585
R4389 gnd.n4905 gnd.n3743 585
R4390 gnd.n4879 gnd.n3743 585
R4391 gnd.n3762 gnd.n3752 585
R4392 gnd.n4922 gnd.n3752 585
R4393 gnd.n4910 gnd.n4909 585
R4394 gnd.n4911 gnd.n4910 585
R4395 gnd.n3761 gnd.n3760 585
R4396 gnd.n3771 gnd.n3760 585
R4397 gnd.n4902 gnd.n4901 585
R4398 gnd.n4901 gnd.n4900 585
R4399 gnd.n3764 gnd.n2910 585
R4400 gnd.n6193 gnd.n2910 585
R4401 gnd.n4868 gnd.n4867 585
R4402 gnd.n4869 gnd.n4868 585
R4403 gnd.n3848 gnd.n2898 585
R4404 gnd.n6199 gnd.n2898 585
R4405 gnd.n4863 gnd.n4862 585
R4406 gnd.n4862 gnd.n2896 585
R4407 gnd.n4861 gnd.n3850 585
R4408 gnd.n4861 gnd.n2870 585
R4409 gnd.n4860 gnd.n3852 585
R4410 gnd.n4860 gnd.n4859 585
R4411 gnd.n4498 gnd.n3851 585
R4412 gnd.n3853 gnd.n3851 585
R4413 gnd.n4496 gnd.n3862 585
R4414 gnd.n4848 gnd.n3862 585
R4415 gnd.n4502 gnd.n4495 585
R4416 gnd.n4495 gnd.n3861 585
R4417 gnd.n4503 gnd.n3870 585
R4418 gnd.n4829 gnd.n3870 585
R4419 gnd.n4504 gnd.n4494 585
R4420 gnd.n4494 gnd.n3878 585
R4421 gnd.n4492 gnd.n3877 585
R4422 gnd.n4821 gnd.n3877 585
R4423 gnd.n4508 gnd.n4491 585
R4424 gnd.n4491 gnd.n3876 585
R4425 gnd.n4509 gnd.n3884 585
R4426 gnd.n4813 gnd.n3884 585
R4427 gnd.n4510 gnd.n4490 585
R4428 gnd.n4490 gnd.n3892 585
R4429 gnd.n4488 gnd.n3891 585
R4430 gnd.n4805 gnd.n3891 585
R4431 gnd.n4514 gnd.n4487 585
R4432 gnd.n4487 gnd.n3890 585
R4433 gnd.n4515 gnd.n3899 585
R4434 gnd.n4797 gnd.n3899 585
R4435 gnd.n4516 gnd.n4486 585
R4436 gnd.n4486 gnd.n3898 585
R4437 gnd.n4484 gnd.n3906 585
R4438 gnd.n4789 gnd.n3906 585
R4439 gnd.n4521 gnd.n4520 585
R4440 gnd.n4521 gnd.n3905 585
R4441 gnd.n4523 gnd.n4522 585
R4442 gnd.n4525 gnd.n4524 585
R4443 gnd.n4527 gnd.n4526 585
R4444 gnd.n4480 gnd.n4479 585
R4445 gnd.n4531 gnd.n4481 585
R4446 gnd.n4533 gnd.n4532 585
R4447 gnd.n4655 gnd.n4534 585
R4448 gnd.n4654 gnd.n4535 585
R4449 gnd.n4653 gnd.n4536 585
R4450 gnd.n4542 gnd.n4537 585
R4451 gnd.n4646 gnd.n4543 585
R4452 gnd.n4645 gnd.n4544 585
R4453 gnd.n4546 gnd.n4545 585
R4454 gnd.n4638 gnd.n4554 585
R4455 gnd.n4637 gnd.n4555 585
R4456 gnd.n4562 gnd.n4556 585
R4457 gnd.n4630 gnd.n4563 585
R4458 gnd.n4629 gnd.n4564 585
R4459 gnd.n4566 gnd.n4565 585
R4460 gnd.n4622 gnd.n4574 585
R4461 gnd.n4621 gnd.n4575 585
R4462 gnd.n4582 gnd.n4576 585
R4463 gnd.n4614 gnd.n4583 585
R4464 gnd.n4613 gnd.n4584 585
R4465 gnd.n4586 gnd.n4585 585
R4466 gnd.n4606 gnd.n4599 585
R4467 gnd.n4605 gnd.n4600 585
R4468 gnd.n3911 gnd.n3910 585
R4469 gnd.n4783 gnd.n4782 585
R4470 gnd.n4782 gnd.n4781 585
R4471 gnd.n6097 gnd.n6096 585
R4472 gnd.n6096 gnd.n6095 585
R4473 gnd.n2992 gnd.n2990 585
R4474 gnd.n2994 gnd.n2992 585
R4475 gnd.n6101 gnd.n2989 585
R4476 gnd.n5473 gnd.n2989 585
R4477 gnd.n6102 gnd.n2988 585
R4478 gnd.n3415 gnd.n2988 585
R4479 gnd.n6103 gnd.n2987 585
R4480 gnd.n5465 gnd.n2987 585
R4481 gnd.n3421 gnd.n2985 585
R4482 gnd.n3422 gnd.n3421 585
R4483 gnd.n6107 gnd.n2984 585
R4484 gnd.n5454 gnd.n2984 585
R4485 gnd.n6108 gnd.n2983 585
R4486 gnd.n3435 gnd.n2983 585
R4487 gnd.n6109 gnd.n2982 585
R4488 gnd.n5446 gnd.n2982 585
R4489 gnd.n3433 gnd.n2980 585
R4490 gnd.n3434 gnd.n3433 585
R4491 gnd.n6113 gnd.n2979 585
R4492 gnd.n5438 gnd.n2979 585
R4493 gnd.n6114 gnd.n2978 585
R4494 gnd.n3448 gnd.n2978 585
R4495 gnd.n6115 gnd.n2977 585
R4496 gnd.n5430 gnd.n2977 585
R4497 gnd.n3446 gnd.n2975 585
R4498 gnd.n3447 gnd.n3446 585
R4499 gnd.n6119 gnd.n2974 585
R4500 gnd.n5422 gnd.n2974 585
R4501 gnd.n6120 gnd.n2973 585
R4502 gnd.n3454 gnd.n2973 585
R4503 gnd.n6121 gnd.n2972 585
R4504 gnd.n5414 gnd.n2972 585
R4505 gnd.n3470 gnd.n2970 585
R4506 gnd.n3471 gnd.n3470 585
R4507 gnd.n6125 gnd.n2969 585
R4508 gnd.n5406 gnd.n2969 585
R4509 gnd.n6126 gnd.n2968 585
R4510 gnd.n3546 gnd.n2968 585
R4511 gnd.n6127 gnd.n2967 585
R4512 gnd.n5267 gnd.n2967 585
R4513 gnd.n3560 gnd.n2965 585
R4514 gnd.n3561 gnd.n3560 585
R4515 gnd.n6131 gnd.n2964 585
R4516 gnd.n5259 gnd.n2964 585
R4517 gnd.n6132 gnd.n2963 585
R4518 gnd.n3565 gnd.n2963 585
R4519 gnd.n6133 gnd.n2962 585
R4520 gnd.n5238 gnd.n2962 585
R4521 gnd.n5194 gnd.n2960 585
R4522 gnd.n5195 gnd.n5194 585
R4523 gnd.n6137 gnd.n2959 585
R4524 gnd.n5230 gnd.n2959 585
R4525 gnd.n6138 gnd.n2958 585
R4526 gnd.n5219 gnd.n2958 585
R4527 gnd.n6139 gnd.n2957 585
R4528 gnd.n5169 gnd.n2957 585
R4529 gnd.n3593 gnd.n2955 585
R4530 gnd.n5188 gnd.n3593 585
R4531 gnd.n6143 gnd.n2954 585
R4532 gnd.n3603 gnd.n2954 585
R4533 gnd.n6144 gnd.n2953 585
R4534 gnd.n5178 gnd.n2953 585
R4535 gnd.n6145 gnd.n2952 585
R4536 gnd.n3612 gnd.n2952 585
R4537 gnd.n3620 gnd.n2950 585
R4538 gnd.n5144 gnd.n3620 585
R4539 gnd.n6149 gnd.n2949 585
R4540 gnd.n5069 gnd.n2949 585
R4541 gnd.n6150 gnd.n2948 585
R4542 gnd.n5136 gnd.n2948 585
R4543 gnd.n6151 gnd.n2947 585
R4544 gnd.n3632 gnd.n2947 585
R4545 gnd.n3639 gnd.n2945 585
R4546 gnd.n3640 gnd.n3639 585
R4547 gnd.n6155 gnd.n2944 585
R4548 gnd.n5110 gnd.n2944 585
R4549 gnd.n6156 gnd.n2943 585
R4550 gnd.n5063 gnd.n2943 585
R4551 gnd.n6157 gnd.n2942 585
R4552 gnd.n5100 gnd.n2942 585
R4553 gnd.n5091 gnd.n2940 585
R4554 gnd.n5092 gnd.n5091 585
R4555 gnd.n6161 gnd.n2939 585
R4556 gnd.n3659 gnd.n2939 585
R4557 gnd.n6162 gnd.n2938 585
R4558 gnd.n5057 gnd.n2938 585
R4559 gnd.n6163 gnd.n2937 585
R4560 gnd.n3682 gnd.n2937 585
R4561 gnd.n5046 gnd.n2935 585
R4562 gnd.n5047 gnd.n5046 585
R4563 gnd.n6167 gnd.n2934 585
R4564 gnd.n5020 gnd.n2934 585
R4565 gnd.n6168 gnd.n2933 585
R4566 gnd.n4992 gnd.n2933 585
R4567 gnd.n6169 gnd.n2932 585
R4568 gnd.n5011 gnd.n2932 585
R4569 gnd.n4982 gnd.n2930 585
R4570 gnd.n4983 gnd.n4982 585
R4571 gnd.n6173 gnd.n2929 585
R4572 gnd.n5001 gnd.n2929 585
R4573 gnd.n6174 gnd.n2928 585
R4574 gnd.n3715 gnd.n2928 585
R4575 gnd.n6175 gnd.n2927 585
R4576 gnd.n4969 gnd.n2927 585
R4577 gnd.n4945 gnd.n2925 585
R4578 gnd.n4946 gnd.n4945 585
R4579 gnd.n6179 gnd.n2924 585
R4580 gnd.n4961 gnd.n2924 585
R4581 gnd.n6180 gnd.n2923 585
R4582 gnd.n3733 gnd.n2923 585
R4583 gnd.n6181 gnd.n2922 585
R4584 gnd.n4930 gnd.n2922 585
R4585 gnd.n4878 gnd.n2920 585
R4586 gnd.n4879 gnd.n4878 585
R4587 gnd.n6185 gnd.n2919 585
R4588 gnd.n4922 gnd.n2919 585
R4589 gnd.n6186 gnd.n2918 585
R4590 gnd.n4911 gnd.n2918 585
R4591 gnd.n6187 gnd.n2917 585
R4592 gnd.n3771 gnd.n2917 585
R4593 gnd.n2914 gnd.n2912 585
R4594 gnd.n4900 gnd.n2912 585
R4595 gnd.n6192 gnd.n6191 585
R4596 gnd.n6193 gnd.n6192 585
R4597 gnd.n2913 gnd.n2911 585
R4598 gnd.n4869 gnd.n2911 585
R4599 gnd.n4837 gnd.n2900 585
R4600 gnd.n6199 gnd.n2900 585
R4601 gnd.n4840 gnd.n4836 585
R4602 gnd.n4836 gnd.n2896 585
R4603 gnd.n4841 gnd.n4835 585
R4604 gnd.n4835 gnd.n2870 585
R4605 gnd.n4842 gnd.n3854 585
R4606 gnd.n4859 gnd.n3854 585
R4607 gnd.n3866 gnd.n3864 585
R4608 gnd.n3864 gnd.n3853 585
R4609 gnd.n4847 gnd.n4846 585
R4610 gnd.n4848 gnd.n4847 585
R4611 gnd.n3865 gnd.n3863 585
R4612 gnd.n3863 gnd.n3861 585
R4613 gnd.n4831 gnd.n4830 585
R4614 gnd.n4830 gnd.n4829 585
R4615 gnd.n3869 gnd.n3868 585
R4616 gnd.n3878 gnd.n3869 585
R4617 gnd.n4820 gnd.n4819 585
R4618 gnd.n4821 gnd.n4820 585
R4619 gnd.n3880 gnd.n3879 585
R4620 gnd.n3879 gnd.n3876 585
R4621 gnd.n4815 gnd.n4814 585
R4622 gnd.n4814 gnd.n4813 585
R4623 gnd.n3883 gnd.n3882 585
R4624 gnd.n3892 gnd.n3883 585
R4625 gnd.n4804 gnd.n4803 585
R4626 gnd.n4805 gnd.n4804 585
R4627 gnd.n3894 gnd.n3893 585
R4628 gnd.n3893 gnd.n3890 585
R4629 gnd.n4799 gnd.n4798 585
R4630 gnd.n4798 gnd.n4797 585
R4631 gnd.n3897 gnd.n3896 585
R4632 gnd.n3898 gnd.n3897 585
R4633 gnd.n4788 gnd.n4787 585
R4634 gnd.n4789 gnd.n4788 585
R4635 gnd.n3908 gnd.n3907 585
R4636 gnd.n3907 gnd.n3905 585
R4637 gnd.n6036 gnd.n3054 585
R4638 gnd.n6037 gnd.n3053 585
R4639 gnd.n3403 gnd.n3047 585
R4640 gnd.n6044 gnd.n3046 585
R4641 gnd.n6045 gnd.n3045 585
R4642 gnd.n3400 gnd.n3039 585
R4643 gnd.n6052 gnd.n3038 585
R4644 gnd.n6053 gnd.n3037 585
R4645 gnd.n3398 gnd.n3031 585
R4646 gnd.n6060 gnd.n3030 585
R4647 gnd.n6061 gnd.n3029 585
R4648 gnd.n3395 gnd.n3023 585
R4649 gnd.n6068 gnd.n3022 585
R4650 gnd.n6069 gnd.n3021 585
R4651 gnd.n3393 gnd.n3014 585
R4652 gnd.n6076 gnd.n3013 585
R4653 gnd.n6077 gnd.n3012 585
R4654 gnd.n3390 gnd.n3009 585
R4655 gnd.n6082 gnd.n3008 585
R4656 gnd.n6083 gnd.n3007 585
R4657 gnd.n6084 gnd.n3006 585
R4658 gnd.n3387 gnd.n3004 585
R4659 gnd.n6088 gnd.n3003 585
R4660 gnd.n6089 gnd.n3002 585
R4661 gnd.n6090 gnd.n2998 585
R4662 gnd.n5578 gnd.n2993 585
R4663 gnd.n5575 gnd.n2993 585
R4664 gnd.n5579 gnd.n5577 585
R4665 gnd.n3385 gnd.n3384 585
R4666 gnd.n3406 gnd.n3405 585
R4667 gnd.n5399 gnd.n3473 463.671
R4668 gnd.n5282 gnd.n5281 463.671
R4669 gnd.n3843 gnd.n3841 463.671
R4670 gnd.n6268 gnd.n2873 463.671
R4671 gnd.n6886 gnd.n6885 452.659
R4672 gnd.n3777 gnd.t192 443.966
R4673 gnd.n3521 gnd.t216 443.966
R4674 gnd.n6205 gnd.t249 443.966
R4675 gnd.n3515 gnd.t265 443.966
R4676 gnd.n4596 gnd.t227 371.625
R4677 gnd.n6030 gnd.t259 371.625
R4678 gnd.n4591 gnd.t271 371.625
R4679 gnd.n3127 gnd.t252 371.625
R4680 gnd.n3150 gnd.t237 371.625
R4681 gnd.n5910 gnd.t174 371.625
R4682 gnd.n352 gnd.t277 371.625
R4683 gnd.n332 gnd.t182 371.625
R4684 gnd.n7818 gnd.t210 371.625
R4685 gnd.n7618 gnd.t231 371.625
R4686 gnd.n2416 gnd.t243 371.625
R4687 gnd.n2438 gnd.t178 371.625
R4688 gnd.n2460 gnd.t200 371.625
R4689 gnd.n4079 gnd.t274 371.625
R4690 gnd.n2822 gnd.t262 371.625
R4691 gnd.n4659 gnd.t196 371.625
R4692 gnd.n4672 gnd.t224 371.625
R4693 gnd.n3055 gnd.t206 371.625
R4694 gnd.n1495 gnd.t220 323.425
R4695 gnd.n1012 gnd.t255 323.425
R4696 gnd.n2324 gnd.n2298 289.615
R4697 gnd.n2292 gnd.n2266 289.615
R4698 gnd.n2260 gnd.n2234 289.615
R4699 gnd.n2229 gnd.n2203 289.615
R4700 gnd.n2197 gnd.n2171 289.615
R4701 gnd.n2165 gnd.n2139 289.615
R4702 gnd.n2133 gnd.n2107 289.615
R4703 gnd.n2102 gnd.n2076 289.615
R4704 gnd.n1569 gnd.t170 279.217
R4705 gnd.n1033 gnd.t280 279.217
R4706 gnd.n2880 gnd.t205 260.649
R4707 gnd.n3486 gnd.t191 260.649
R4708 gnd.n6270 gnd.n6269 256.663
R4709 gnd.n6270 gnd.n2839 256.663
R4710 gnd.n6270 gnd.n2840 256.663
R4711 gnd.n6270 gnd.n2841 256.663
R4712 gnd.n6270 gnd.n2842 256.663
R4713 gnd.n6270 gnd.n2843 256.663
R4714 gnd.n6270 gnd.n2844 256.663
R4715 gnd.n6270 gnd.n2845 256.663
R4716 gnd.n6270 gnd.n2846 256.663
R4717 gnd.n6270 gnd.n2847 256.663
R4718 gnd.n6270 gnd.n2848 256.663
R4719 gnd.n6270 gnd.n2849 256.663
R4720 gnd.n6270 gnd.n2850 256.663
R4721 gnd.n6270 gnd.n2851 256.663
R4722 gnd.n6270 gnd.n2852 256.663
R4723 gnd.n6270 gnd.n2853 256.663
R4724 gnd.n6273 gnd.n2837 256.663
R4725 gnd.n6271 gnd.n6270 256.663
R4726 gnd.n6270 gnd.n2854 256.663
R4727 gnd.n6270 gnd.n2855 256.663
R4728 gnd.n6270 gnd.n2856 256.663
R4729 gnd.n6270 gnd.n2857 256.663
R4730 gnd.n6270 gnd.n2858 256.663
R4731 gnd.n6270 gnd.n2859 256.663
R4732 gnd.n6270 gnd.n2860 256.663
R4733 gnd.n6270 gnd.n2861 256.663
R4734 gnd.n6270 gnd.n2862 256.663
R4735 gnd.n6270 gnd.n2863 256.663
R4736 gnd.n6270 gnd.n2864 256.663
R4737 gnd.n6270 gnd.n2865 256.663
R4738 gnd.n6270 gnd.n2866 256.663
R4739 gnd.n6270 gnd.n2867 256.663
R4740 gnd.n6270 gnd.n2868 256.663
R4741 gnd.n6270 gnd.n2869 256.663
R4742 gnd.n5280 gnd.n3461 256.663
R4743 gnd.n5287 gnd.n3461 256.663
R4744 gnd.n3542 gnd.n3461 256.663
R4745 gnd.n5294 gnd.n3461 256.663
R4746 gnd.n3539 gnd.n3461 256.663
R4747 gnd.n5301 gnd.n3461 256.663
R4748 gnd.n3536 gnd.n3461 256.663
R4749 gnd.n5308 gnd.n3461 256.663
R4750 gnd.n3533 gnd.n3461 256.663
R4751 gnd.n5315 gnd.n3461 256.663
R4752 gnd.n3530 gnd.n3461 256.663
R4753 gnd.n5322 gnd.n3461 256.663
R4754 gnd.n3527 gnd.n3461 256.663
R4755 gnd.n5329 gnd.n3461 256.663
R4756 gnd.n3524 gnd.n3461 256.663
R4757 gnd.n5337 gnd.n3461 256.663
R4758 gnd.n5340 gnd.n3137 256.663
R4759 gnd.n5341 gnd.n3461 256.663
R4760 gnd.n5345 gnd.n3461 256.663
R4761 gnd.n3518 gnd.n3461 256.663
R4762 gnd.n5353 gnd.n3461 256.663
R4763 gnd.n3513 gnd.n3461 256.663
R4764 gnd.n5360 gnd.n3461 256.663
R4765 gnd.n3510 gnd.n3461 256.663
R4766 gnd.n5367 gnd.n3461 256.663
R4767 gnd.n3507 gnd.n3461 256.663
R4768 gnd.n5374 gnd.n3461 256.663
R4769 gnd.n3504 gnd.n3461 256.663
R4770 gnd.n5381 gnd.n3461 256.663
R4771 gnd.n3501 gnd.n3461 256.663
R4772 gnd.n5388 gnd.n3461 256.663
R4773 gnd.n3498 gnd.n3461 256.663
R4774 gnd.n5395 gnd.n3461 256.663
R4775 gnd.n5398 gnd.n3461 256.663
R4776 gnd.n6625 gnd.n2384 242.672
R4777 gnd.n6625 gnd.n2385 242.672
R4778 gnd.n6625 gnd.n2386 242.672
R4779 gnd.n6625 gnd.n2387 242.672
R4780 gnd.n6625 gnd.n2388 242.672
R4781 gnd.n6625 gnd.n2389 242.672
R4782 gnd.n6625 gnd.n2390 242.672
R4783 gnd.n6625 gnd.n2391 242.672
R4784 gnd.n6625 gnd.n2392 242.672
R4785 gnd.n6324 gnd.n2775 242.672
R4786 gnd.n6324 gnd.n2774 242.672
R4787 gnd.n6324 gnd.n2773 242.672
R4788 gnd.n6324 gnd.n2772 242.672
R4789 gnd.n6324 gnd.n2771 242.672
R4790 gnd.n6324 gnd.n2770 242.672
R4791 gnd.n6324 gnd.n2769 242.672
R4792 gnd.n6324 gnd.n2768 242.672
R4793 gnd.n6324 gnd.n2767 242.672
R4794 gnd.n1623 gnd.n1622 242.672
R4795 gnd.n1623 gnd.n1533 242.672
R4796 gnd.n1623 gnd.n1534 242.672
R4797 gnd.n1623 gnd.n1535 242.672
R4798 gnd.n1623 gnd.n1536 242.672
R4799 gnd.n1623 gnd.n1537 242.672
R4800 gnd.n1623 gnd.n1538 242.672
R4801 gnd.n1623 gnd.n1539 242.672
R4802 gnd.n1623 gnd.n1540 242.672
R4803 gnd.n1623 gnd.n1541 242.672
R4804 gnd.n1623 gnd.n1542 242.672
R4805 gnd.n1623 gnd.n1543 242.672
R4806 gnd.n1624 gnd.n1623 242.672
R4807 gnd.n6672 gnd.n2355 242.672
R4808 gnd.n6672 gnd.n1029 242.672
R4809 gnd.n6672 gnd.n1028 242.672
R4810 gnd.n6672 gnd.n1027 242.672
R4811 gnd.n6672 gnd.n1026 242.672
R4812 gnd.n6672 gnd.n1025 242.672
R4813 gnd.n6672 gnd.n1024 242.672
R4814 gnd.n6672 gnd.n1023 242.672
R4815 gnd.n6672 gnd.n1022 242.672
R4816 gnd.n6672 gnd.n1021 242.672
R4817 gnd.n6672 gnd.n1020 242.672
R4818 gnd.n6672 gnd.n1019 242.672
R4819 gnd.n6672 gnd.n1018 242.672
R4820 gnd.n6027 gnd.n3092 242.672
R4821 gnd.n6027 gnd.n3094 242.672
R4822 gnd.n6027 gnd.n3095 242.672
R4823 gnd.n6027 gnd.n3097 242.672
R4824 gnd.n6027 gnd.n3099 242.672
R4825 gnd.n6027 gnd.n3100 242.672
R4826 gnd.n6027 gnd.n3102 242.672
R4827 gnd.n6027 gnd.n3104 242.672
R4828 gnd.n6028 gnd.n6027 242.672
R4829 gnd.n7853 gnd.n266 242.672
R4830 gnd.n7853 gnd.n265 242.672
R4831 gnd.n7853 gnd.n264 242.672
R4832 gnd.n7853 gnd.n263 242.672
R4833 gnd.n7853 gnd.n262 242.672
R4834 gnd.n7853 gnd.n261 242.672
R4835 gnd.n7853 gnd.n260 242.672
R4836 gnd.n7853 gnd.n259 242.672
R4837 gnd.n7853 gnd.n258 242.672
R4838 gnd.n1707 gnd.n1706 242.672
R4839 gnd.n1706 gnd.n1445 242.672
R4840 gnd.n1706 gnd.n1446 242.672
R4841 gnd.n1706 gnd.n1447 242.672
R4842 gnd.n1706 gnd.n1448 242.672
R4843 gnd.n1706 gnd.n1449 242.672
R4844 gnd.n1706 gnd.n1450 242.672
R4845 gnd.n1706 gnd.n1451 242.672
R4846 gnd.n6672 gnd.n1011 242.672
R4847 gnd.n6673 gnd.n6672 242.672
R4848 gnd.n6672 gnd.n6626 242.672
R4849 gnd.n6672 gnd.n6627 242.672
R4850 gnd.n6672 gnd.n6628 242.672
R4851 gnd.n6672 gnd.n6629 242.672
R4852 gnd.n6672 gnd.n6630 242.672
R4853 gnd.n6672 gnd.n6631 242.672
R4854 gnd.n6625 gnd.n6624 242.672
R4855 gnd.n6625 gnd.n2356 242.672
R4856 gnd.n6625 gnd.n2357 242.672
R4857 gnd.n6625 gnd.n2358 242.672
R4858 gnd.n6625 gnd.n2359 242.672
R4859 gnd.n6625 gnd.n2360 242.672
R4860 gnd.n6625 gnd.n2361 242.672
R4861 gnd.n6625 gnd.n2362 242.672
R4862 gnd.n6625 gnd.n2363 242.672
R4863 gnd.n6625 gnd.n2364 242.672
R4864 gnd.n6625 gnd.n2365 242.672
R4865 gnd.n6625 gnd.n2366 242.672
R4866 gnd.n6625 gnd.n2367 242.672
R4867 gnd.n6625 gnd.n2368 242.672
R4868 gnd.n6625 gnd.n2369 242.672
R4869 gnd.n6625 gnd.n2370 242.672
R4870 gnd.n6625 gnd.n2371 242.672
R4871 gnd.n6625 gnd.n2372 242.672
R4872 gnd.n6625 gnd.n2373 242.672
R4873 gnd.n6625 gnd.n2374 242.672
R4874 gnd.n6625 gnd.n2375 242.672
R4875 gnd.n6625 gnd.n2376 242.672
R4876 gnd.n6625 gnd.n2377 242.672
R4877 gnd.n6625 gnd.n2378 242.672
R4878 gnd.n6625 gnd.n2379 242.672
R4879 gnd.n6625 gnd.n2380 242.672
R4880 gnd.n6625 gnd.n2381 242.672
R4881 gnd.n6625 gnd.n2382 242.672
R4882 gnd.n6625 gnd.n2383 242.672
R4883 gnd.n6324 gnd.n2777 242.672
R4884 gnd.n6324 gnd.n2778 242.672
R4885 gnd.n6324 gnd.n2779 242.672
R4886 gnd.n6324 gnd.n2780 242.672
R4887 gnd.n6324 gnd.n2781 242.672
R4888 gnd.n6324 gnd.n2782 242.672
R4889 gnd.n6324 gnd.n2783 242.672
R4890 gnd.n6324 gnd.n2784 242.672
R4891 gnd.n6324 gnd.n2785 242.672
R4892 gnd.n6324 gnd.n2786 242.672
R4893 gnd.n6324 gnd.n2787 242.672
R4894 gnd.n6324 gnd.n2788 242.672
R4895 gnd.n6324 gnd.n2789 242.672
R4896 gnd.n6324 gnd.n2790 242.672
R4897 gnd.n6324 gnd.n2791 242.672
R4898 gnd.n6324 gnd.n2792 242.672
R4899 gnd.n6274 gnd.n2833 242.672
R4900 gnd.n6324 gnd.n2793 242.672
R4901 gnd.n6324 gnd.n2794 242.672
R4902 gnd.n6324 gnd.n2795 242.672
R4903 gnd.n6324 gnd.n2796 242.672
R4904 gnd.n6324 gnd.n2797 242.672
R4905 gnd.n6324 gnd.n2798 242.672
R4906 gnd.n6324 gnd.n2799 242.672
R4907 gnd.n6324 gnd.n2800 242.672
R4908 gnd.n6324 gnd.n2801 242.672
R4909 gnd.n6324 gnd.n2802 242.672
R4910 gnd.n6324 gnd.n2803 242.672
R4911 gnd.n6324 gnd.n2804 242.672
R4912 gnd.n6324 gnd.n6323 242.672
R4913 gnd.n6027 gnd.n6026 242.672
R4914 gnd.n6027 gnd.n3064 242.672
R4915 gnd.n6027 gnd.n3065 242.672
R4916 gnd.n6027 gnd.n3066 242.672
R4917 gnd.n6027 gnd.n3067 242.672
R4918 gnd.n6027 gnd.n3068 242.672
R4919 gnd.n6027 gnd.n3069 242.672
R4920 gnd.n6027 gnd.n3070 242.672
R4921 gnd.n6027 gnd.n3071 242.672
R4922 gnd.n6027 gnd.n3072 242.672
R4923 gnd.n6027 gnd.n3073 242.672
R4924 gnd.n6027 gnd.n3074 242.672
R4925 gnd.n6027 gnd.n3075 242.672
R4926 gnd.n5974 gnd.n3138 242.672
R4927 gnd.n6027 gnd.n3076 242.672
R4928 gnd.n6027 gnd.n3077 242.672
R4929 gnd.n6027 gnd.n3078 242.672
R4930 gnd.n6027 gnd.n3079 242.672
R4931 gnd.n6027 gnd.n3080 242.672
R4932 gnd.n6027 gnd.n3081 242.672
R4933 gnd.n6027 gnd.n3082 242.672
R4934 gnd.n6027 gnd.n3083 242.672
R4935 gnd.n6027 gnd.n3084 242.672
R4936 gnd.n6027 gnd.n3085 242.672
R4937 gnd.n6027 gnd.n3086 242.672
R4938 gnd.n6027 gnd.n3087 242.672
R4939 gnd.n6027 gnd.n3088 242.672
R4940 gnd.n6027 gnd.n3089 242.672
R4941 gnd.n6027 gnd.n3090 242.672
R4942 gnd.n6027 gnd.n3091 242.672
R4943 gnd.n7853 gnd.n267 242.672
R4944 gnd.n7853 gnd.n268 242.672
R4945 gnd.n7853 gnd.n269 242.672
R4946 gnd.n7853 gnd.n270 242.672
R4947 gnd.n7853 gnd.n271 242.672
R4948 gnd.n7853 gnd.n272 242.672
R4949 gnd.n7853 gnd.n273 242.672
R4950 gnd.n7853 gnd.n274 242.672
R4951 gnd.n7853 gnd.n275 242.672
R4952 gnd.n7853 gnd.n276 242.672
R4953 gnd.n7853 gnd.n277 242.672
R4954 gnd.n7853 gnd.n278 242.672
R4955 gnd.n7853 gnd.n279 242.672
R4956 gnd.n7853 gnd.n280 242.672
R4957 gnd.n7853 gnd.n281 242.672
R4958 gnd.n7853 gnd.n282 242.672
R4959 gnd.n7853 gnd.n283 242.672
R4960 gnd.n7853 gnd.n284 242.672
R4961 gnd.n7853 gnd.n285 242.672
R4962 gnd.n7853 gnd.n286 242.672
R4963 gnd.n7853 gnd.n287 242.672
R4964 gnd.n7853 gnd.n288 242.672
R4965 gnd.n7853 gnd.n289 242.672
R4966 gnd.n7853 gnd.n290 242.672
R4967 gnd.n7853 gnd.n291 242.672
R4968 gnd.n7853 gnd.n292 242.672
R4969 gnd.n7853 gnd.n293 242.672
R4970 gnd.n7853 gnd.n294 242.672
R4971 gnd.n7853 gnd.n7852 242.672
R4972 gnd.n4781 gnd.n3913 242.672
R4973 gnd.n4781 gnd.n3914 242.672
R4974 gnd.n4781 gnd.n3915 242.672
R4975 gnd.n4781 gnd.n3916 242.672
R4976 gnd.n4781 gnd.n3917 242.672
R4977 gnd.n4781 gnd.n3918 242.672
R4978 gnd.n4781 gnd.n3919 242.672
R4979 gnd.n4781 gnd.n3920 242.672
R4980 gnd.n4781 gnd.n3921 242.672
R4981 gnd.n4781 gnd.n3922 242.672
R4982 gnd.n4781 gnd.n3923 242.672
R4983 gnd.n4781 gnd.n3924 242.672
R4984 gnd.n4781 gnd.n3925 242.672
R4985 gnd.n4781 gnd.n3926 242.672
R4986 gnd.n5575 gnd.n3407 242.672
R4987 gnd.n5575 gnd.n3404 242.672
R4988 gnd.n5575 gnd.n3402 242.672
R4989 gnd.n5575 gnd.n3401 242.672
R4990 gnd.n5575 gnd.n3399 242.672
R4991 gnd.n5575 gnd.n3397 242.672
R4992 gnd.n5575 gnd.n3396 242.672
R4993 gnd.n5575 gnd.n3394 242.672
R4994 gnd.n5575 gnd.n3392 242.672
R4995 gnd.n5575 gnd.n3391 242.672
R4996 gnd.n5575 gnd.n3389 242.672
R4997 gnd.n5575 gnd.n3388 242.672
R4998 gnd.n5575 gnd.n3386 242.672
R4999 gnd.n5576 gnd.n5575 242.672
R5000 gnd.n7854 gnd.n255 240.244
R5001 gnd.n7851 gnd.n295 240.244
R5002 gnd.n7847 gnd.n7846 240.244
R5003 gnd.n7843 gnd.n7842 240.244
R5004 gnd.n7839 gnd.n7838 240.244
R5005 gnd.n7835 gnd.n7834 240.244
R5006 gnd.n7831 gnd.n7830 240.244
R5007 gnd.n7827 gnd.n7826 240.244
R5008 gnd.n7823 gnd.n7822 240.244
R5009 gnd.n7816 gnd.n7815 240.244
R5010 gnd.n7812 gnd.n7811 240.244
R5011 gnd.n7808 gnd.n7807 240.244
R5012 gnd.n7804 gnd.n7803 240.244
R5013 gnd.n7800 gnd.n7799 240.244
R5014 gnd.n7796 gnd.n7795 240.244
R5015 gnd.n7792 gnd.n7791 240.244
R5016 gnd.n7788 gnd.n7787 240.244
R5017 gnd.n7784 gnd.n7783 240.244
R5018 gnd.n7780 gnd.n7779 240.244
R5019 gnd.n7773 gnd.n7772 240.244
R5020 gnd.n7770 gnd.n7769 240.244
R5021 gnd.n7766 gnd.n7765 240.244
R5022 gnd.n7762 gnd.n7761 240.244
R5023 gnd.n7758 gnd.n7757 240.244
R5024 gnd.n7754 gnd.n7753 240.244
R5025 gnd.n7750 gnd.n7749 240.244
R5026 gnd.n7746 gnd.n7745 240.244
R5027 gnd.n7742 gnd.n7741 240.244
R5028 gnd.n7738 gnd.n7737 240.244
R5029 gnd.n5907 gnd.n3171 240.244
R5030 gnd.n5899 gnd.n3171 240.244
R5031 gnd.n5899 gnd.n3182 240.244
R5032 gnd.n3198 gnd.n3182 240.244
R5033 gnd.n5595 gnd.n3198 240.244
R5034 gnd.n5595 gnd.n3211 240.244
R5035 gnd.n5600 gnd.n3211 240.244
R5036 gnd.n5600 gnd.n3222 240.244
R5037 gnd.n5610 gnd.n3222 240.244
R5038 gnd.n5610 gnd.n3232 240.244
R5039 gnd.n5615 gnd.n3232 240.244
R5040 gnd.n5615 gnd.n3243 240.244
R5041 gnd.n5625 gnd.n3243 240.244
R5042 gnd.n5625 gnd.n3252 240.244
R5043 gnd.n5630 gnd.n3252 240.244
R5044 gnd.n5630 gnd.n3263 240.244
R5045 gnd.n5640 gnd.n3263 240.244
R5046 gnd.n5640 gnd.n3273 240.244
R5047 gnd.n5645 gnd.n3273 240.244
R5048 gnd.n5645 gnd.n3284 240.244
R5049 gnd.n5655 gnd.n3284 240.244
R5050 gnd.n5655 gnd.n3293 240.244
R5051 gnd.n5660 gnd.n3293 240.244
R5052 gnd.n5660 gnd.n3305 240.244
R5053 gnd.n5682 gnd.n3305 240.244
R5054 gnd.n5682 gnd.n3315 240.244
R5055 gnd.n3319 gnd.n3315 240.244
R5056 gnd.n5687 gnd.n3319 240.244
R5057 gnd.n5687 gnd.n5686 240.244
R5058 gnd.n5686 gnd.n3329 240.244
R5059 gnd.n3339 gnd.n3329 240.244
R5060 gnd.n3351 gnd.n3339 240.244
R5061 gnd.n5800 gnd.n3351 240.244
R5062 gnd.n5800 gnd.n102 240.244
R5063 gnd.n5796 gnd.n102 240.244
R5064 gnd.n5796 gnd.n5703 240.244
R5065 gnd.n5703 gnd.n119 240.244
R5066 gnd.n5719 gnd.n119 240.244
R5067 gnd.n5719 gnd.n130 240.244
R5068 gnd.n5776 gnd.n130 240.244
R5069 gnd.n5776 gnd.n140 240.244
R5070 gnd.n5772 gnd.n140 240.244
R5071 gnd.n5772 gnd.n149 240.244
R5072 gnd.n5764 gnd.n149 240.244
R5073 gnd.n5764 gnd.n160 240.244
R5074 gnd.n360 gnd.n160 240.244
R5075 gnd.n360 gnd.n169 240.244
R5076 gnd.n7702 gnd.n169 240.244
R5077 gnd.n7702 gnd.n180 240.244
R5078 gnd.n7705 gnd.n180 240.244
R5079 gnd.n7705 gnd.n189 240.244
R5080 gnd.n7709 gnd.n189 240.244
R5081 gnd.n7709 gnd.n200 240.244
R5082 gnd.n7712 gnd.n200 240.244
R5083 gnd.n7712 gnd.n209 240.244
R5084 gnd.n7716 gnd.n209 240.244
R5085 gnd.n7716 gnd.n219 240.244
R5086 gnd.n7719 gnd.n219 240.244
R5087 gnd.n7719 gnd.n228 240.244
R5088 gnd.n7723 gnd.n228 240.244
R5089 gnd.n7723 gnd.n238 240.244
R5090 gnd.n7726 gnd.n238 240.244
R5091 gnd.n7726 gnd.n247 240.244
R5092 gnd.n7730 gnd.n247 240.244
R5093 gnd.n3107 gnd.n3106 240.244
R5094 gnd.n6020 gnd.n3106 240.244
R5095 gnd.n6018 gnd.n6017 240.244
R5096 gnd.n6014 gnd.n6013 240.244
R5097 gnd.n6010 gnd.n6009 240.244
R5098 gnd.n6006 gnd.n6005 240.244
R5099 gnd.n6002 gnd.n6001 240.244
R5100 gnd.n5998 gnd.n5997 240.244
R5101 gnd.n5994 gnd.n5993 240.244
R5102 gnd.n5989 gnd.n5988 240.244
R5103 gnd.n5985 gnd.n5984 240.244
R5104 gnd.n5981 gnd.n5980 240.244
R5105 gnd.n5977 gnd.n5976 240.244
R5106 gnd.n5972 gnd.n5971 240.244
R5107 gnd.n5968 gnd.n5967 240.244
R5108 gnd.n5964 gnd.n5963 240.244
R5109 gnd.n5960 gnd.n5959 240.244
R5110 gnd.n5956 gnd.n5955 240.244
R5111 gnd.n5952 gnd.n5951 240.244
R5112 gnd.n5948 gnd.n5947 240.244
R5113 gnd.n5944 gnd.n5943 240.244
R5114 gnd.n5940 gnd.n5939 240.244
R5115 gnd.n5936 gnd.n5935 240.244
R5116 gnd.n5932 gnd.n5931 240.244
R5117 gnd.n5928 gnd.n5927 240.244
R5118 gnd.n5924 gnd.n5923 240.244
R5119 gnd.n5920 gnd.n5919 240.244
R5120 gnd.n5916 gnd.n5915 240.244
R5121 gnd.n3186 gnd.n3108 240.244
R5122 gnd.n5897 gnd.n3186 240.244
R5123 gnd.n5897 gnd.n3187 240.244
R5124 gnd.n5893 gnd.n3187 240.244
R5125 gnd.n5893 gnd.n3196 240.244
R5126 gnd.n5885 gnd.n3196 240.244
R5127 gnd.n5885 gnd.n3214 240.244
R5128 gnd.n5881 gnd.n3214 240.244
R5129 gnd.n5881 gnd.n3220 240.244
R5130 gnd.n5873 gnd.n3220 240.244
R5131 gnd.n5873 gnd.n3235 240.244
R5132 gnd.n5869 gnd.n3235 240.244
R5133 gnd.n5869 gnd.n3241 240.244
R5134 gnd.n5861 gnd.n3241 240.244
R5135 gnd.n5861 gnd.n3255 240.244
R5136 gnd.n5857 gnd.n3255 240.244
R5137 gnd.n5857 gnd.n3261 240.244
R5138 gnd.n5849 gnd.n3261 240.244
R5139 gnd.n5849 gnd.n3276 240.244
R5140 gnd.n5845 gnd.n3276 240.244
R5141 gnd.n5845 gnd.n3282 240.244
R5142 gnd.n5837 gnd.n3282 240.244
R5143 gnd.n5837 gnd.n3296 240.244
R5144 gnd.n5833 gnd.n3296 240.244
R5145 gnd.n5833 gnd.n3303 240.244
R5146 gnd.n5825 gnd.n3303 240.244
R5147 gnd.n5825 gnd.n5822 240.244
R5148 gnd.n5822 gnd.n3318 240.244
R5149 gnd.n3335 gnd.n3318 240.244
R5150 gnd.n5811 gnd.n3335 240.244
R5151 gnd.n5811 gnd.n5808 240.244
R5152 gnd.n5808 gnd.n3338 240.244
R5153 gnd.n3338 gnd.n105 240.244
R5154 gnd.n7946 gnd.n105 240.244
R5155 gnd.n7946 gnd.n106 240.244
R5156 gnd.n116 gnd.n106 240.244
R5157 gnd.n7940 gnd.n116 240.244
R5158 gnd.n7940 gnd.n117 240.244
R5159 gnd.n7932 gnd.n117 240.244
R5160 gnd.n7932 gnd.n133 240.244
R5161 gnd.n7928 gnd.n133 240.244
R5162 gnd.n7928 gnd.n138 240.244
R5163 gnd.n7920 gnd.n138 240.244
R5164 gnd.n7920 gnd.n152 240.244
R5165 gnd.n7916 gnd.n152 240.244
R5166 gnd.n7916 gnd.n158 240.244
R5167 gnd.n7908 gnd.n158 240.244
R5168 gnd.n7908 gnd.n172 240.244
R5169 gnd.n7904 gnd.n172 240.244
R5170 gnd.n7904 gnd.n178 240.244
R5171 gnd.n7896 gnd.n178 240.244
R5172 gnd.n7896 gnd.n192 240.244
R5173 gnd.n7892 gnd.n192 240.244
R5174 gnd.n7892 gnd.n198 240.244
R5175 gnd.n7884 gnd.n198 240.244
R5176 gnd.n7884 gnd.n212 240.244
R5177 gnd.n7880 gnd.n212 240.244
R5178 gnd.n7880 gnd.n218 240.244
R5179 gnd.n7872 gnd.n218 240.244
R5180 gnd.n7872 gnd.n231 240.244
R5181 gnd.n7868 gnd.n231 240.244
R5182 gnd.n7868 gnd.n237 240.244
R5183 gnd.n7860 gnd.n237 240.244
R5184 gnd.n7860 gnd.n250 240.244
R5185 gnd.n6325 gnd.n2764 240.244
R5186 gnd.n6322 gnd.n2805 240.244
R5187 gnd.n6318 gnd.n6317 240.244
R5188 gnd.n6314 gnd.n6313 240.244
R5189 gnd.n6310 gnd.n6309 240.244
R5190 gnd.n6306 gnd.n6305 240.244
R5191 gnd.n6302 gnd.n6301 240.244
R5192 gnd.n6298 gnd.n6297 240.244
R5193 gnd.n6294 gnd.n6293 240.244
R5194 gnd.n6289 gnd.n6288 240.244
R5195 gnd.n6285 gnd.n6284 240.244
R5196 gnd.n6281 gnd.n6280 240.244
R5197 gnd.n6277 gnd.n6276 240.244
R5198 gnd.n4681 gnd.n4680 240.244
R5199 gnd.n4684 gnd.n4683 240.244
R5200 gnd.n4691 gnd.n4690 240.244
R5201 gnd.n4694 gnd.n4693 240.244
R5202 gnd.n4699 gnd.n4674 240.244
R5203 gnd.n4703 gnd.n4702 240.244
R5204 gnd.n4710 gnd.n4709 240.244
R5205 gnd.n4713 gnd.n4712 240.244
R5206 gnd.n4720 gnd.n4719 240.244
R5207 gnd.n4723 gnd.n4722 240.244
R5208 gnd.n4730 gnd.n4729 240.244
R5209 gnd.n4733 gnd.n4732 240.244
R5210 gnd.n4740 gnd.n4739 240.244
R5211 gnd.n4743 gnd.n4742 240.244
R5212 gnd.n4748 gnd.n4661 240.244
R5213 gnd.n6503 gnd.n6502 240.244
R5214 gnd.n6502 gnd.n2467 240.244
R5215 gnd.n2479 gnd.n2467 240.244
R5216 gnd.n4048 gnd.n2479 240.244
R5217 gnd.n4048 gnd.n2491 240.244
R5218 gnd.n4052 gnd.n2491 240.244
R5219 gnd.n4052 gnd.n2501 240.244
R5220 gnd.n4055 gnd.n2501 240.244
R5221 gnd.n4055 gnd.n2510 240.244
R5222 gnd.n4059 gnd.n2510 240.244
R5223 gnd.n4059 gnd.n2520 240.244
R5224 gnd.n4062 gnd.n2520 240.244
R5225 gnd.n4062 gnd.n2530 240.244
R5226 gnd.n4066 gnd.n2530 240.244
R5227 gnd.n4066 gnd.n2540 240.244
R5228 gnd.n4172 gnd.n2540 240.244
R5229 gnd.n4172 gnd.n2550 240.244
R5230 gnd.n4040 gnd.n2550 240.244
R5231 gnd.n4040 gnd.n2560 240.244
R5232 gnd.n4182 gnd.n2560 240.244
R5233 gnd.n4182 gnd.n2570 240.244
R5234 gnd.n4035 gnd.n2570 240.244
R5235 gnd.n4035 gnd.n2580 240.244
R5236 gnd.n4230 gnd.n2580 240.244
R5237 gnd.n4230 gnd.n2590 240.244
R5238 gnd.n4026 gnd.n2590 240.244
R5239 gnd.n4026 gnd.n2599 240.244
R5240 gnd.n4246 gnd.n2599 240.244
R5241 gnd.n4246 gnd.n2609 240.244
R5242 gnd.n4017 gnd.n2609 240.244
R5243 gnd.n4017 gnd.n4011 240.244
R5244 gnd.n4288 gnd.n4011 240.244
R5245 gnd.n4288 gnd.n4003 240.244
R5246 gnd.n4003 gnd.n3996 240.244
R5247 gnd.n4295 gnd.n3996 240.244
R5248 gnd.n4295 gnd.n3989 240.244
R5249 gnd.n3989 gnd.n2625 240.244
R5250 gnd.n3982 gnd.n2625 240.244
R5251 gnd.n3982 gnd.n2636 240.244
R5252 gnd.n4357 gnd.n2636 240.244
R5253 gnd.n4357 gnd.n2646 240.244
R5254 gnd.n4361 gnd.n2646 240.244
R5255 gnd.n4361 gnd.n2655 240.244
R5256 gnd.n4371 gnd.n2655 240.244
R5257 gnd.n4371 gnd.n2666 240.244
R5258 gnd.n3963 gnd.n2666 240.244
R5259 gnd.n3963 gnd.n2675 240.244
R5260 gnd.n4378 gnd.n2675 240.244
R5261 gnd.n4378 gnd.n2686 240.244
R5262 gnd.n4383 gnd.n2686 240.244
R5263 gnd.n4383 gnd.n2695 240.244
R5264 gnd.n4390 gnd.n2695 240.244
R5265 gnd.n4390 gnd.n2706 240.244
R5266 gnd.n3951 gnd.n2706 240.244
R5267 gnd.n3951 gnd.n2715 240.244
R5268 gnd.n4460 gnd.n2715 240.244
R5269 gnd.n4460 gnd.n2726 240.244
R5270 gnd.n4464 gnd.n2726 240.244
R5271 gnd.n4464 gnd.n2735 240.244
R5272 gnd.n4474 gnd.n2735 240.244
R5273 gnd.n4474 gnd.n2746 240.244
R5274 gnd.n4759 gnd.n2746 240.244
R5275 gnd.n4759 gnd.n2756 240.244
R5276 gnd.n3935 gnd.n2756 240.244
R5277 gnd.n2396 gnd.n2395 240.244
R5278 gnd.n6618 gnd.n2395 240.244
R5279 gnd.n6616 gnd.n6615 240.244
R5280 gnd.n6612 gnd.n6611 240.244
R5281 gnd.n6608 gnd.n6607 240.244
R5282 gnd.n6604 gnd.n6603 240.244
R5283 gnd.n6600 gnd.n6599 240.244
R5284 gnd.n6596 gnd.n6595 240.244
R5285 gnd.n6592 gnd.n6591 240.244
R5286 gnd.n6587 gnd.n6586 240.244
R5287 gnd.n6583 gnd.n6582 240.244
R5288 gnd.n6579 gnd.n6578 240.244
R5289 gnd.n6575 gnd.n6574 240.244
R5290 gnd.n6571 gnd.n6570 240.244
R5291 gnd.n6567 gnd.n6566 240.244
R5292 gnd.n6563 gnd.n6562 240.244
R5293 gnd.n6559 gnd.n6558 240.244
R5294 gnd.n6555 gnd.n6554 240.244
R5295 gnd.n6551 gnd.n6550 240.244
R5296 gnd.n6547 gnd.n6546 240.244
R5297 gnd.n6543 gnd.n6542 240.244
R5298 gnd.n6539 gnd.n6538 240.244
R5299 gnd.n6535 gnd.n6534 240.244
R5300 gnd.n6531 gnd.n6530 240.244
R5301 gnd.n6527 gnd.n6526 240.244
R5302 gnd.n6523 gnd.n6522 240.244
R5303 gnd.n6519 gnd.n6518 240.244
R5304 gnd.n6515 gnd.n6514 240.244
R5305 gnd.n6511 gnd.n6510 240.244
R5306 gnd.n6500 gnd.n2397 240.244
R5307 gnd.n6500 gnd.n2470 240.244
R5308 gnd.n6496 gnd.n2470 240.244
R5309 gnd.n6496 gnd.n2477 240.244
R5310 gnd.n6488 gnd.n2477 240.244
R5311 gnd.n6488 gnd.n2494 240.244
R5312 gnd.n6484 gnd.n2494 240.244
R5313 gnd.n6484 gnd.n2500 240.244
R5314 gnd.n6476 gnd.n2500 240.244
R5315 gnd.n6476 gnd.n2512 240.244
R5316 gnd.n6472 gnd.n2512 240.244
R5317 gnd.n6472 gnd.n2518 240.244
R5318 gnd.n6464 gnd.n2518 240.244
R5319 gnd.n6464 gnd.n2533 240.244
R5320 gnd.n6460 gnd.n2533 240.244
R5321 gnd.n6460 gnd.n2539 240.244
R5322 gnd.n6452 gnd.n2539 240.244
R5323 gnd.n6452 gnd.n2552 240.244
R5324 gnd.n6448 gnd.n2552 240.244
R5325 gnd.n6448 gnd.n2558 240.244
R5326 gnd.n6440 gnd.n2558 240.244
R5327 gnd.n6440 gnd.n2573 240.244
R5328 gnd.n6436 gnd.n2573 240.244
R5329 gnd.n6436 gnd.n2579 240.244
R5330 gnd.n6428 gnd.n2579 240.244
R5331 gnd.n6428 gnd.n2592 240.244
R5332 gnd.n6424 gnd.n2592 240.244
R5333 gnd.n6424 gnd.n2597 240.244
R5334 gnd.n6416 gnd.n2597 240.244
R5335 gnd.n6416 gnd.n2612 240.244
R5336 gnd.n4237 gnd.n2612 240.244
R5337 gnd.n4237 gnd.n3999 240.244
R5338 gnd.n4304 gnd.n3999 240.244
R5339 gnd.n4308 gnd.n4304 240.244
R5340 gnd.n4308 gnd.n4305 240.244
R5341 gnd.n4305 gnd.n2622 240.244
R5342 gnd.n6411 gnd.n2622 240.244
R5343 gnd.n6411 gnd.n2623 240.244
R5344 gnd.n6403 gnd.n2623 240.244
R5345 gnd.n6403 gnd.n2639 240.244
R5346 gnd.n6399 gnd.n2639 240.244
R5347 gnd.n6399 gnd.n2644 240.244
R5348 gnd.n6391 gnd.n2644 240.244
R5349 gnd.n6391 gnd.n2658 240.244
R5350 gnd.n6387 gnd.n2658 240.244
R5351 gnd.n6387 gnd.n2664 240.244
R5352 gnd.n6379 gnd.n2664 240.244
R5353 gnd.n6379 gnd.n2678 240.244
R5354 gnd.n6375 gnd.n2678 240.244
R5355 gnd.n6375 gnd.n2684 240.244
R5356 gnd.n6367 gnd.n2684 240.244
R5357 gnd.n6367 gnd.n2698 240.244
R5358 gnd.n6363 gnd.n2698 240.244
R5359 gnd.n6363 gnd.n2704 240.244
R5360 gnd.n6355 gnd.n2704 240.244
R5361 gnd.n6355 gnd.n2718 240.244
R5362 gnd.n6351 gnd.n2718 240.244
R5363 gnd.n6351 gnd.n2724 240.244
R5364 gnd.n6343 gnd.n2724 240.244
R5365 gnd.n6343 gnd.n2738 240.244
R5366 gnd.n6339 gnd.n2738 240.244
R5367 gnd.n6339 gnd.n2744 240.244
R5368 gnd.n6331 gnd.n2744 240.244
R5369 gnd.n6331 gnd.n2759 240.244
R5370 gnd.n6671 gnd.n6632 240.244
R5371 gnd.n6664 gnd.n6663 240.244
R5372 gnd.n6661 gnd.n6660 240.244
R5373 gnd.n6657 gnd.n6656 240.244
R5374 gnd.n6653 gnd.n6652 240.244
R5375 gnd.n6649 gnd.n6648 240.244
R5376 gnd.n6645 gnd.n1017 240.244
R5377 gnd.n6675 gnd.n6674 240.244
R5378 gnd.n1718 gnd.n1430 240.244
R5379 gnd.n1728 gnd.n1430 240.244
R5380 gnd.n1728 gnd.n1421 240.244
R5381 gnd.n1421 gnd.n1410 240.244
R5382 gnd.n1749 gnd.n1410 240.244
R5383 gnd.n1749 gnd.n1404 240.244
R5384 gnd.n1759 gnd.n1404 240.244
R5385 gnd.n1759 gnd.n1393 240.244
R5386 gnd.n1393 gnd.n1383 240.244
R5387 gnd.n1785 gnd.n1383 240.244
R5388 gnd.n1786 gnd.n1785 240.244
R5389 gnd.n1787 gnd.n1786 240.244
R5390 gnd.n1787 gnd.n1362 240.244
R5391 gnd.n1823 gnd.n1362 240.244
R5392 gnd.n1823 gnd.n1363 240.244
R5393 gnd.n1819 gnd.n1363 240.244
R5394 gnd.n1819 gnd.n1818 240.244
R5395 gnd.n1818 gnd.n1239 240.244
R5396 gnd.n1853 gnd.n1239 240.244
R5397 gnd.n1853 gnd.n1229 240.244
R5398 gnd.n1229 gnd.n1221 240.244
R5399 gnd.n1871 gnd.n1221 240.244
R5400 gnd.n1872 gnd.n1871 240.244
R5401 gnd.n1872 gnd.n1209 240.244
R5402 gnd.n1209 gnd.n1198 240.244
R5403 gnd.n1903 gnd.n1198 240.244
R5404 gnd.n1904 gnd.n1903 240.244
R5405 gnd.n1906 gnd.n1904 240.244
R5406 gnd.n1906 gnd.n1184 240.244
R5407 gnd.n1938 gnd.n1184 240.244
R5408 gnd.n1938 gnd.n1170 240.244
R5409 gnd.n1960 gnd.n1170 240.244
R5410 gnd.n1961 gnd.n1960 240.244
R5411 gnd.n1961 gnd.n1157 240.244
R5412 gnd.n1157 gnd.n1147 240.244
R5413 gnd.n1992 gnd.n1147 240.244
R5414 gnd.n1993 gnd.n1992 240.244
R5415 gnd.n1994 gnd.n1993 240.244
R5416 gnd.n1994 gnd.n1132 240.244
R5417 gnd.n1996 gnd.n1132 240.244
R5418 gnd.n1996 gnd.n1118 240.244
R5419 gnd.n2065 gnd.n1118 240.244
R5420 gnd.n2066 gnd.n2065 240.244
R5421 gnd.n2067 gnd.n2066 240.244
R5422 gnd.n2067 gnd.n966 240.244
R5423 gnd.n1113 gnd.n966 240.244
R5424 gnd.n1113 gnd.n977 240.244
R5425 gnd.n2335 gnd.n977 240.244
R5426 gnd.n2336 gnd.n2335 240.244
R5427 gnd.n2336 gnd.n990 240.244
R5428 gnd.n2344 gnd.n990 240.244
R5429 gnd.n2344 gnd.n1002 240.244
R5430 gnd.n6682 gnd.n1002 240.244
R5431 gnd.n1708 gnd.n1443 240.244
R5432 gnd.n1464 gnd.n1443 240.244
R5433 gnd.n1467 gnd.n1466 240.244
R5434 gnd.n1474 gnd.n1473 240.244
R5435 gnd.n1477 gnd.n1476 240.244
R5436 gnd.n1484 gnd.n1483 240.244
R5437 gnd.n1487 gnd.n1486 240.244
R5438 gnd.n1494 gnd.n1493 240.244
R5439 gnd.n1716 gnd.n1440 240.244
R5440 gnd.n1440 gnd.n1419 240.244
R5441 gnd.n1739 gnd.n1419 240.244
R5442 gnd.n1739 gnd.n1413 240.244
R5443 gnd.n1747 gnd.n1413 240.244
R5444 gnd.n1747 gnd.n1415 240.244
R5445 gnd.n1415 gnd.n1391 240.244
R5446 gnd.n1769 gnd.n1391 240.244
R5447 gnd.n1769 gnd.n1386 240.244
R5448 gnd.n1783 gnd.n1386 240.244
R5449 gnd.n1783 gnd.n1387 240.244
R5450 gnd.n1779 gnd.n1387 240.244
R5451 gnd.n1779 gnd.n1359 240.244
R5452 gnd.n1826 gnd.n1359 240.244
R5453 gnd.n1827 gnd.n1826 240.244
R5454 gnd.n1828 gnd.n1827 240.244
R5455 gnd.n1828 gnd.n1355 240.244
R5456 gnd.n1834 gnd.n1355 240.244
R5457 gnd.n1834 gnd.n1228 240.244
R5458 gnd.n1863 gnd.n1228 240.244
R5459 gnd.n1863 gnd.n1224 240.244
R5460 gnd.n1869 gnd.n1224 240.244
R5461 gnd.n1869 gnd.n1207 240.244
R5462 gnd.n1893 gnd.n1207 240.244
R5463 gnd.n1893 gnd.n1202 240.244
R5464 gnd.n1901 gnd.n1202 240.244
R5465 gnd.n1901 gnd.n1203 240.244
R5466 gnd.n1203 gnd.n1182 240.244
R5467 gnd.n1942 gnd.n1182 240.244
R5468 gnd.n1942 gnd.n1177 240.244
R5469 gnd.n1950 gnd.n1177 240.244
R5470 gnd.n1950 gnd.n1178 240.244
R5471 gnd.n1178 gnd.n1155 240.244
R5472 gnd.n1982 gnd.n1155 240.244
R5473 gnd.n1982 gnd.n1150 240.244
R5474 gnd.n1990 gnd.n1150 240.244
R5475 gnd.n1990 gnd.n1151 240.244
R5476 gnd.n1151 gnd.n1130 240.244
R5477 gnd.n2043 gnd.n1130 240.244
R5478 gnd.n2043 gnd.n1125 240.244
R5479 gnd.n2055 gnd.n1125 240.244
R5480 gnd.n2055 gnd.n1126 240.244
R5481 gnd.n2051 gnd.n1126 240.244
R5482 gnd.n2051 gnd.n968 240.244
R5483 gnd.n6708 gnd.n968 240.244
R5484 gnd.n6708 gnd.n969 240.244
R5485 gnd.n6704 gnd.n969 240.244
R5486 gnd.n6704 gnd.n975 240.244
R5487 gnd.n991 gnd.n975 240.244
R5488 gnd.n6694 gnd.n991 240.244
R5489 gnd.n6694 gnd.n992 240.244
R5490 gnd.n6690 gnd.n992 240.244
R5491 gnd.n6690 gnd.n1000 240.244
R5492 gnd.n7629 gnd.n257 240.244
R5493 gnd.n7635 gnd.n7634 240.244
R5494 gnd.n7638 gnd.n7637 240.244
R5495 gnd.n7645 gnd.n7644 240.244
R5496 gnd.n7648 gnd.n7647 240.244
R5497 gnd.n7655 gnd.n7654 240.244
R5498 gnd.n7658 gnd.n7657 240.244
R5499 gnd.n7665 gnd.n7664 240.244
R5500 gnd.n7668 gnd.n7667 240.244
R5501 gnd.n3381 gnd.n3174 240.244
R5502 gnd.n3381 gnd.n3183 240.244
R5503 gnd.n5587 gnd.n3183 240.244
R5504 gnd.n5587 gnd.n3199 240.244
R5505 gnd.n5593 gnd.n3199 240.244
R5506 gnd.n5593 gnd.n3212 240.244
R5507 gnd.n5602 gnd.n3212 240.244
R5508 gnd.n5602 gnd.n3223 240.244
R5509 gnd.n5608 gnd.n3223 240.244
R5510 gnd.n5608 gnd.n3233 240.244
R5511 gnd.n5617 gnd.n3233 240.244
R5512 gnd.n5617 gnd.n3244 240.244
R5513 gnd.n5623 gnd.n3244 240.244
R5514 gnd.n5623 gnd.n3253 240.244
R5515 gnd.n5632 gnd.n3253 240.244
R5516 gnd.n5632 gnd.n3264 240.244
R5517 gnd.n5638 gnd.n3264 240.244
R5518 gnd.n5638 gnd.n3274 240.244
R5519 gnd.n5647 gnd.n3274 240.244
R5520 gnd.n5647 gnd.n3285 240.244
R5521 gnd.n5653 gnd.n3285 240.244
R5522 gnd.n5653 gnd.n3294 240.244
R5523 gnd.n5662 gnd.n3294 240.244
R5524 gnd.n5662 gnd.n3306 240.244
R5525 gnd.n5680 gnd.n3306 240.244
R5526 gnd.n5680 gnd.n3316 240.244
R5527 gnd.n3320 gnd.n3316 240.244
R5528 gnd.n5667 gnd.n3320 240.244
R5529 gnd.n5668 gnd.n5667 240.244
R5530 gnd.n5668 gnd.n3330 240.244
R5531 gnd.n3340 gnd.n3330 240.244
R5532 gnd.n3349 gnd.n3340 240.244
R5533 gnd.n3349 gnd.n98 240.244
R5534 gnd.n7948 gnd.n98 240.244
R5535 gnd.n7948 gnd.n100 240.244
R5536 gnd.n5723 gnd.n100 240.244
R5537 gnd.n5723 gnd.n120 240.244
R5538 gnd.n5782 gnd.n120 240.244
R5539 gnd.n5782 gnd.n131 240.244
R5540 gnd.n5778 gnd.n131 240.244
R5541 gnd.n5778 gnd.n141 240.244
R5542 gnd.n5770 gnd.n141 240.244
R5543 gnd.n5770 gnd.n150 240.244
R5544 gnd.n5766 gnd.n150 240.244
R5545 gnd.n5766 gnd.n161 240.244
R5546 gnd.n7597 gnd.n161 240.244
R5547 gnd.n7597 gnd.n170 240.244
R5548 gnd.n7700 gnd.n170 240.244
R5549 gnd.n7700 gnd.n181 240.244
R5550 gnd.n7696 gnd.n181 240.244
R5551 gnd.n7696 gnd.n190 240.244
R5552 gnd.n7693 gnd.n190 240.244
R5553 gnd.n7693 gnd.n201 240.244
R5554 gnd.n7690 gnd.n201 240.244
R5555 gnd.n7690 gnd.n210 240.244
R5556 gnd.n7687 gnd.n210 240.244
R5557 gnd.n7687 gnd.n220 240.244
R5558 gnd.n7684 gnd.n220 240.244
R5559 gnd.n7684 gnd.n229 240.244
R5560 gnd.n7681 gnd.n229 240.244
R5561 gnd.n7681 gnd.n239 240.244
R5562 gnd.n7678 gnd.n239 240.244
R5563 gnd.n7678 gnd.n248 240.244
R5564 gnd.n7675 gnd.n248 240.244
R5565 gnd.n3018 gnd.n3017 240.244
R5566 gnd.n3093 gnd.n3025 240.244
R5567 gnd.n3096 gnd.n3026 240.244
R5568 gnd.n3034 gnd.n3033 240.244
R5569 gnd.n3098 gnd.n3041 240.244
R5570 gnd.n3101 gnd.n3042 240.244
R5571 gnd.n3050 gnd.n3049 240.244
R5572 gnd.n3103 gnd.n3059 240.244
R5573 gnd.n6029 gnd.n3062 240.244
R5574 gnd.n5905 gnd.n3177 240.244
R5575 gnd.n3185 gnd.n3177 240.244
R5576 gnd.n3201 gnd.n3185 240.244
R5577 gnd.n5891 gnd.n3201 240.244
R5578 gnd.n5891 gnd.n3202 240.244
R5579 gnd.n5887 gnd.n3202 240.244
R5580 gnd.n5887 gnd.n3209 240.244
R5581 gnd.n5879 gnd.n3209 240.244
R5582 gnd.n5879 gnd.n3225 240.244
R5583 gnd.n5875 gnd.n3225 240.244
R5584 gnd.n5875 gnd.n3230 240.244
R5585 gnd.n5867 gnd.n3230 240.244
R5586 gnd.n5867 gnd.n3245 240.244
R5587 gnd.n5863 gnd.n3245 240.244
R5588 gnd.n5863 gnd.n3250 240.244
R5589 gnd.n5855 gnd.n3250 240.244
R5590 gnd.n5855 gnd.n3266 240.244
R5591 gnd.n5851 gnd.n3266 240.244
R5592 gnd.n5851 gnd.n3271 240.244
R5593 gnd.n5843 gnd.n3271 240.244
R5594 gnd.n5843 gnd.n3286 240.244
R5595 gnd.n5839 gnd.n3286 240.244
R5596 gnd.n5839 gnd.n3291 240.244
R5597 gnd.n5831 gnd.n3291 240.244
R5598 gnd.n5831 gnd.n3308 240.244
R5599 gnd.n5827 gnd.n3308 240.244
R5600 gnd.n5827 gnd.n3313 240.244
R5601 gnd.n5691 gnd.n3313 240.244
R5602 gnd.n5692 gnd.n5691 240.244
R5603 gnd.n5692 gnd.n3332 240.244
R5604 gnd.n5806 gnd.n3332 240.244
R5605 gnd.n5806 gnd.n3342 240.244
R5606 gnd.n5802 gnd.n3342 240.244
R5607 gnd.n5802 gnd.n104 240.244
R5608 gnd.n5794 gnd.n104 240.244
R5609 gnd.n5794 gnd.n122 240.244
R5610 gnd.n7938 gnd.n122 240.244
R5611 gnd.n7938 gnd.n123 240.244
R5612 gnd.n7934 gnd.n123 240.244
R5613 gnd.n7934 gnd.n129 240.244
R5614 gnd.n7926 gnd.n129 240.244
R5615 gnd.n7926 gnd.n142 240.244
R5616 gnd.n7922 gnd.n142 240.244
R5617 gnd.n7922 gnd.n147 240.244
R5618 gnd.n7914 gnd.n147 240.244
R5619 gnd.n7914 gnd.n163 240.244
R5620 gnd.n7910 gnd.n163 240.244
R5621 gnd.n7910 gnd.n168 240.244
R5622 gnd.n7902 gnd.n168 240.244
R5623 gnd.n7902 gnd.n182 240.244
R5624 gnd.n7898 gnd.n182 240.244
R5625 gnd.n7898 gnd.n187 240.244
R5626 gnd.n7890 gnd.n187 240.244
R5627 gnd.n7890 gnd.n203 240.244
R5628 gnd.n7886 gnd.n203 240.244
R5629 gnd.n7886 gnd.n208 240.244
R5630 gnd.n7878 gnd.n208 240.244
R5631 gnd.n7878 gnd.n221 240.244
R5632 gnd.n7874 gnd.n221 240.244
R5633 gnd.n7874 gnd.n226 240.244
R5634 gnd.n7866 gnd.n226 240.244
R5635 gnd.n7866 gnd.n241 240.244
R5636 gnd.n7862 gnd.n241 240.244
R5637 gnd.n7862 gnd.n246 240.244
R5638 gnd.n1046 gnd.n1006 240.244
R5639 gnd.n1054 gnd.n1053 240.244
R5640 gnd.n1057 gnd.n1056 240.244
R5641 gnd.n1064 gnd.n1063 240.244
R5642 gnd.n1067 gnd.n1066 240.244
R5643 gnd.n1074 gnd.n1073 240.244
R5644 gnd.n1077 gnd.n1076 240.244
R5645 gnd.n1084 gnd.n1083 240.244
R5646 gnd.n1087 gnd.n1086 240.244
R5647 gnd.n1094 gnd.n1093 240.244
R5648 gnd.n1097 gnd.n1096 240.244
R5649 gnd.n1104 gnd.n1103 240.244
R5650 gnd.n1106 gnd.n1030 240.244
R5651 gnd.n1631 gnd.n1528 240.244
R5652 gnd.n1631 gnd.n1521 240.244
R5653 gnd.n1642 gnd.n1521 240.244
R5654 gnd.n1642 gnd.n1517 240.244
R5655 gnd.n1648 gnd.n1517 240.244
R5656 gnd.n1648 gnd.n1509 240.244
R5657 gnd.n1658 gnd.n1509 240.244
R5658 gnd.n1658 gnd.n1504 240.244
R5659 gnd.n1694 gnd.n1504 240.244
R5660 gnd.n1694 gnd.n1505 240.244
R5661 gnd.n1505 gnd.n1452 240.244
R5662 gnd.n1689 gnd.n1452 240.244
R5663 gnd.n1689 gnd.n1688 240.244
R5664 gnd.n1688 gnd.n1431 240.244
R5665 gnd.n1684 gnd.n1431 240.244
R5666 gnd.n1684 gnd.n1422 240.244
R5667 gnd.n1681 gnd.n1422 240.244
R5668 gnd.n1681 gnd.n1680 240.244
R5669 gnd.n1680 gnd.n1405 240.244
R5670 gnd.n1676 gnd.n1405 240.244
R5671 gnd.n1676 gnd.n1394 240.244
R5672 gnd.n1394 gnd.n1374 240.244
R5673 gnd.n1795 gnd.n1374 240.244
R5674 gnd.n1795 gnd.n1369 240.244
R5675 gnd.n1803 gnd.n1369 240.244
R5676 gnd.n1803 gnd.n1370 240.244
R5677 gnd.n1370 gnd.n1338 240.244
R5678 gnd.n1843 gnd.n1338 240.244
R5679 gnd.n1843 gnd.n1339 240.244
R5680 gnd.n1354 gnd.n1339 240.244
R5681 gnd.n1354 gnd.n1241 240.244
R5682 gnd.n1850 gnd.n1241 240.244
R5683 gnd.n1850 gnd.n1230 240.244
R5684 gnd.n1243 gnd.n1230 240.244
R5685 gnd.n1243 gnd.n1220 240.244
R5686 gnd.n1250 gnd.n1220 240.244
R5687 gnd.n1250 gnd.n1210 240.244
R5688 gnd.n1247 gnd.n1210 240.244
R5689 gnd.n1247 gnd.n1189 240.244
R5690 gnd.n1915 gnd.n1189 240.244
R5691 gnd.n1915 gnd.n1185 240.244
R5692 gnd.n1937 gnd.n1185 240.244
R5693 gnd.n1937 gnd.n1175 240.244
R5694 gnd.n1933 gnd.n1175 240.244
R5695 gnd.n1933 gnd.n1169 240.244
R5696 gnd.n1930 gnd.n1169 240.244
R5697 gnd.n1930 gnd.n1158 240.244
R5698 gnd.n1927 gnd.n1158 240.244
R5699 gnd.n1927 gnd.n1137 240.244
R5700 gnd.n2005 gnd.n1137 240.244
R5701 gnd.n2005 gnd.n1133 240.244
R5702 gnd.n2040 gnd.n1133 240.244
R5703 gnd.n2040 gnd.n1124 240.244
R5704 gnd.n2036 gnd.n1124 240.244
R5705 gnd.n2036 gnd.n954 240.244
R5706 gnd.n2032 gnd.n954 240.244
R5707 gnd.n2032 gnd.n965 240.244
R5708 gnd.n2028 gnd.n965 240.244
R5709 gnd.n2028 gnd.n2027 240.244
R5710 gnd.n2027 gnd.n978 240.244
R5711 gnd.n2023 gnd.n978 240.244
R5712 gnd.n2023 gnd.n989 240.244
R5713 gnd.n2347 gnd.n989 240.244
R5714 gnd.n2348 gnd.n2347 240.244
R5715 gnd.n2348 gnd.n1003 240.244
R5716 gnd.n1545 gnd.n1544 240.244
R5717 gnd.n1616 gnd.n1544 240.244
R5718 gnd.n1614 gnd.n1613 240.244
R5719 gnd.n1610 gnd.n1609 240.244
R5720 gnd.n1606 gnd.n1605 240.244
R5721 gnd.n1602 gnd.n1601 240.244
R5722 gnd.n1598 gnd.n1597 240.244
R5723 gnd.n1594 gnd.n1593 240.244
R5724 gnd.n1590 gnd.n1589 240.244
R5725 gnd.n1586 gnd.n1585 240.244
R5726 gnd.n1582 gnd.n1581 240.244
R5727 gnd.n1578 gnd.n1577 240.244
R5728 gnd.n1574 gnd.n1532 240.244
R5729 gnd.n1634 gnd.n1526 240.244
R5730 gnd.n1634 gnd.n1522 240.244
R5731 gnd.n1640 gnd.n1522 240.244
R5732 gnd.n1640 gnd.n1515 240.244
R5733 gnd.n1650 gnd.n1515 240.244
R5734 gnd.n1650 gnd.n1511 240.244
R5735 gnd.n1656 gnd.n1511 240.244
R5736 gnd.n1656 gnd.n1502 240.244
R5737 gnd.n1696 gnd.n1502 240.244
R5738 gnd.n1696 gnd.n1453 240.244
R5739 gnd.n1704 gnd.n1453 240.244
R5740 gnd.n1704 gnd.n1454 240.244
R5741 gnd.n1454 gnd.n1432 240.244
R5742 gnd.n1725 gnd.n1432 240.244
R5743 gnd.n1725 gnd.n1424 240.244
R5744 gnd.n1736 gnd.n1424 240.244
R5745 gnd.n1736 gnd.n1425 240.244
R5746 gnd.n1425 gnd.n1406 240.244
R5747 gnd.n1756 gnd.n1406 240.244
R5748 gnd.n1756 gnd.n1396 240.244
R5749 gnd.n1766 gnd.n1396 240.244
R5750 gnd.n1766 gnd.n1377 240.244
R5751 gnd.n1793 gnd.n1377 240.244
R5752 gnd.n1793 gnd.n1367 240.244
R5753 gnd.n1806 gnd.n1367 240.244
R5754 gnd.n1807 gnd.n1806 240.244
R5755 gnd.n1807 gnd.n1342 240.244
R5756 gnd.n1841 gnd.n1342 240.244
R5757 gnd.n1841 gnd.n1343 240.244
R5758 gnd.n1837 gnd.n1343 240.244
R5759 gnd.n1837 gnd.n1351 240.244
R5760 gnd.n1351 gnd.n1232 240.244
R5761 gnd.n1860 gnd.n1232 240.244
R5762 gnd.n1860 gnd.n1219 240.244
R5763 gnd.n1875 gnd.n1219 240.244
R5764 gnd.n1875 gnd.n1212 240.244
R5765 gnd.n1890 gnd.n1212 240.244
R5766 gnd.n1890 gnd.n1213 240.244
R5767 gnd.n1213 gnd.n1191 240.244
R5768 gnd.n1913 gnd.n1191 240.244
R5769 gnd.n1913 gnd.n1192 240.244
R5770 gnd.n1192 gnd.n1174 240.244
R5771 gnd.n1953 gnd.n1174 240.244
R5772 gnd.n1953 gnd.n1167 240.244
R5773 gnd.n1964 gnd.n1167 240.244
R5774 gnd.n1964 gnd.n1160 240.244
R5775 gnd.n1979 gnd.n1160 240.244
R5776 gnd.n1979 gnd.n1161 240.244
R5777 gnd.n1161 gnd.n1140 240.244
R5778 gnd.n2003 gnd.n1140 240.244
R5779 gnd.n2003 gnd.n1141 240.244
R5780 gnd.n1141 gnd.n1122 240.244
R5781 gnd.n2058 gnd.n1122 240.244
R5782 gnd.n2058 gnd.n956 240.244
R5783 gnd.n6715 gnd.n956 240.244
R5784 gnd.n6715 gnd.n957 240.244
R5785 gnd.n6711 gnd.n957 240.244
R5786 gnd.n6711 gnd.n963 240.244
R5787 gnd.n980 gnd.n963 240.244
R5788 gnd.n6701 gnd.n980 240.244
R5789 gnd.n6701 gnd.n981 240.244
R5790 gnd.n6697 gnd.n981 240.244
R5791 gnd.n6697 gnd.n987 240.244
R5792 gnd.n1005 gnd.n987 240.244
R5793 gnd.n6687 gnd.n1005 240.244
R5794 gnd.n4539 gnd.n2766 240.244
R5795 gnd.n4549 gnd.n4548 240.244
R5796 gnd.n4551 gnd.n4550 240.244
R5797 gnd.n4559 gnd.n4558 240.244
R5798 gnd.n4569 gnd.n4568 240.244
R5799 gnd.n4571 gnd.n4570 240.244
R5800 gnd.n4579 gnd.n4578 240.244
R5801 gnd.n4589 gnd.n4588 240.244
R5802 gnd.n4593 gnd.n4590 240.244
R5803 gnd.n4136 gnd.n2468 240.244
R5804 gnd.n4139 gnd.n2468 240.244
R5805 gnd.n4139 gnd.n2480 240.244
R5806 gnd.n4144 gnd.n2480 240.244
R5807 gnd.n4144 gnd.n2492 240.244
R5808 gnd.n4147 gnd.n2492 240.244
R5809 gnd.n4147 gnd.n2502 240.244
R5810 gnd.n4152 gnd.n2502 240.244
R5811 gnd.n4152 gnd.n2511 240.244
R5812 gnd.n4155 gnd.n2511 240.244
R5813 gnd.n4155 gnd.n2521 240.244
R5814 gnd.n4160 gnd.n2521 240.244
R5815 gnd.n4160 gnd.n2531 240.244
R5816 gnd.n4163 gnd.n2531 240.244
R5817 gnd.n4163 gnd.n2541 240.244
R5818 gnd.n4170 gnd.n2541 240.244
R5819 gnd.n4170 gnd.n2551 240.244
R5820 gnd.n4188 gnd.n2551 240.244
R5821 gnd.n4188 gnd.n2561 240.244
R5822 gnd.n4184 gnd.n2561 240.244
R5823 gnd.n4184 gnd.n2571 240.244
R5824 gnd.n4221 gnd.n2571 240.244
R5825 gnd.n4221 gnd.n2581 240.244
R5826 gnd.n4228 gnd.n2581 240.244
R5827 gnd.n4228 gnd.n2591 240.244
R5828 gnd.n4252 gnd.n2591 240.244
R5829 gnd.n4252 gnd.n2600 240.244
R5830 gnd.n4248 gnd.n2600 240.244
R5831 gnd.n4248 gnd.n2610 240.244
R5832 gnd.n4280 gnd.n2610 240.244
R5833 gnd.n4280 gnd.n4013 240.244
R5834 gnd.n4286 gnd.n4013 240.244
R5835 gnd.n4286 gnd.n3994 240.244
R5836 gnd.n4310 gnd.n3994 240.244
R5837 gnd.n4310 gnd.n3990 240.244
R5838 gnd.n4316 gnd.n3990 240.244
R5839 gnd.n4316 gnd.n2626 240.244
R5840 gnd.n4349 gnd.n2626 240.244
R5841 gnd.n4349 gnd.n2637 240.244
R5842 gnd.n4355 gnd.n2637 240.244
R5843 gnd.n4355 gnd.n2647 240.244
R5844 gnd.n4363 gnd.n2647 240.244
R5845 gnd.n4363 gnd.n2656 240.244
R5846 gnd.n4369 gnd.n2656 240.244
R5847 gnd.n4369 gnd.n2667 240.244
R5848 gnd.n4404 gnd.n2667 240.244
R5849 gnd.n4404 gnd.n2676 240.244
R5850 gnd.n3968 gnd.n2676 240.244
R5851 gnd.n3968 gnd.n2687 240.244
R5852 gnd.n3969 gnd.n2687 240.244
R5853 gnd.n3969 gnd.n2696 240.244
R5854 gnd.n4392 gnd.n2696 240.244
R5855 gnd.n4392 gnd.n2707 240.244
R5856 gnd.n4452 gnd.n2707 240.244
R5857 gnd.n4452 gnd.n2716 240.244
R5858 gnd.n4458 gnd.n2716 240.244
R5859 gnd.n4458 gnd.n2727 240.244
R5860 gnd.n4466 gnd.n2727 240.244
R5861 gnd.n4466 gnd.n2736 240.244
R5862 gnd.n4472 gnd.n2736 240.244
R5863 gnd.n4472 gnd.n2747 240.244
R5864 gnd.n4761 gnd.n2747 240.244
R5865 gnd.n4761 gnd.n2757 240.244
R5866 gnd.n4767 gnd.n2757 240.244
R5867 gnd.n4096 gnd.n4095 240.244
R5868 gnd.n4102 gnd.n4101 240.244
R5869 gnd.n4106 gnd.n4105 240.244
R5870 gnd.n4112 gnd.n4111 240.244
R5871 gnd.n4116 gnd.n4115 240.244
R5872 gnd.n4122 gnd.n4121 240.244
R5873 gnd.n4126 gnd.n4125 240.244
R5874 gnd.n4083 gnd.n4082 240.244
R5875 gnd.n4078 gnd.n2393 240.244
R5876 gnd.n4091 gnd.n2469 240.244
R5877 gnd.n2482 gnd.n2469 240.244
R5878 gnd.n6494 gnd.n2482 240.244
R5879 gnd.n6494 gnd.n2483 240.244
R5880 gnd.n6490 gnd.n2483 240.244
R5881 gnd.n6490 gnd.n2490 240.244
R5882 gnd.n6482 gnd.n2490 240.244
R5883 gnd.n6482 gnd.n2504 240.244
R5884 gnd.n6478 gnd.n2504 240.244
R5885 gnd.n6478 gnd.n2509 240.244
R5886 gnd.n6470 gnd.n2509 240.244
R5887 gnd.n6470 gnd.n2523 240.244
R5888 gnd.n6466 gnd.n2523 240.244
R5889 gnd.n6466 gnd.n2528 240.244
R5890 gnd.n6458 gnd.n2528 240.244
R5891 gnd.n6458 gnd.n2543 240.244
R5892 gnd.n6454 gnd.n2543 240.244
R5893 gnd.n6454 gnd.n2548 240.244
R5894 gnd.n6446 gnd.n2548 240.244
R5895 gnd.n6446 gnd.n2563 240.244
R5896 gnd.n6442 gnd.n2563 240.244
R5897 gnd.n6442 gnd.n2568 240.244
R5898 gnd.n6434 gnd.n2568 240.244
R5899 gnd.n6434 gnd.n2583 240.244
R5900 gnd.n6430 gnd.n2583 240.244
R5901 gnd.n6430 gnd.n2588 240.244
R5902 gnd.n6422 gnd.n2588 240.244
R5903 gnd.n6422 gnd.n2602 240.244
R5904 gnd.n6418 gnd.n2602 240.244
R5905 gnd.n6418 gnd.n2607 240.244
R5906 gnd.n4239 gnd.n2607 240.244
R5907 gnd.n4239 gnd.n4004 240.244
R5908 gnd.n4302 gnd.n4004 240.244
R5909 gnd.n4302 gnd.n3998 240.244
R5910 gnd.n4298 gnd.n3998 240.244
R5911 gnd.n4298 gnd.n2628 240.244
R5912 gnd.n6409 gnd.n2628 240.244
R5913 gnd.n6409 gnd.n2629 240.244
R5914 gnd.n6405 gnd.n2629 240.244
R5915 gnd.n6405 gnd.n2635 240.244
R5916 gnd.n6397 gnd.n2635 240.244
R5917 gnd.n6397 gnd.n2648 240.244
R5918 gnd.n6393 gnd.n2648 240.244
R5919 gnd.n6393 gnd.n2653 240.244
R5920 gnd.n6385 gnd.n2653 240.244
R5921 gnd.n6385 gnd.n2669 240.244
R5922 gnd.n6381 gnd.n2669 240.244
R5923 gnd.n6381 gnd.n2674 240.244
R5924 gnd.n6373 gnd.n2674 240.244
R5925 gnd.n6373 gnd.n2688 240.244
R5926 gnd.n6369 gnd.n2688 240.244
R5927 gnd.n6369 gnd.n2693 240.244
R5928 gnd.n6361 gnd.n2693 240.244
R5929 gnd.n6361 gnd.n2709 240.244
R5930 gnd.n6357 gnd.n2709 240.244
R5931 gnd.n6357 gnd.n2714 240.244
R5932 gnd.n6349 gnd.n2714 240.244
R5933 gnd.n6349 gnd.n2728 240.244
R5934 gnd.n6345 gnd.n2728 240.244
R5935 gnd.n6345 gnd.n2733 240.244
R5936 gnd.n6337 gnd.n2733 240.244
R5937 gnd.n6337 gnd.n2749 240.244
R5938 gnd.n6333 gnd.n2749 240.244
R5939 gnd.n6333 gnd.n2754 240.244
R5940 gnd.n6888 gnd.n785 240.244
R5941 gnd.n6888 gnd.n781 240.244
R5942 gnd.n6894 gnd.n781 240.244
R5943 gnd.n6894 gnd.n779 240.244
R5944 gnd.n6898 gnd.n779 240.244
R5945 gnd.n6898 gnd.n775 240.244
R5946 gnd.n6904 gnd.n775 240.244
R5947 gnd.n6904 gnd.n773 240.244
R5948 gnd.n6908 gnd.n773 240.244
R5949 gnd.n6908 gnd.n769 240.244
R5950 gnd.n6914 gnd.n769 240.244
R5951 gnd.n6914 gnd.n767 240.244
R5952 gnd.n6918 gnd.n767 240.244
R5953 gnd.n6918 gnd.n763 240.244
R5954 gnd.n6924 gnd.n763 240.244
R5955 gnd.n6924 gnd.n761 240.244
R5956 gnd.n6928 gnd.n761 240.244
R5957 gnd.n6928 gnd.n757 240.244
R5958 gnd.n6934 gnd.n757 240.244
R5959 gnd.n6934 gnd.n755 240.244
R5960 gnd.n6938 gnd.n755 240.244
R5961 gnd.n6938 gnd.n751 240.244
R5962 gnd.n6944 gnd.n751 240.244
R5963 gnd.n6944 gnd.n749 240.244
R5964 gnd.n6948 gnd.n749 240.244
R5965 gnd.n6948 gnd.n745 240.244
R5966 gnd.n6954 gnd.n745 240.244
R5967 gnd.n6954 gnd.n743 240.244
R5968 gnd.n6958 gnd.n743 240.244
R5969 gnd.n6958 gnd.n739 240.244
R5970 gnd.n6964 gnd.n739 240.244
R5971 gnd.n6964 gnd.n737 240.244
R5972 gnd.n6968 gnd.n737 240.244
R5973 gnd.n6968 gnd.n733 240.244
R5974 gnd.n6974 gnd.n733 240.244
R5975 gnd.n6974 gnd.n731 240.244
R5976 gnd.n6978 gnd.n731 240.244
R5977 gnd.n6978 gnd.n727 240.244
R5978 gnd.n6984 gnd.n727 240.244
R5979 gnd.n6984 gnd.n725 240.244
R5980 gnd.n6988 gnd.n725 240.244
R5981 gnd.n6988 gnd.n721 240.244
R5982 gnd.n6994 gnd.n721 240.244
R5983 gnd.n6994 gnd.n719 240.244
R5984 gnd.n6998 gnd.n719 240.244
R5985 gnd.n6998 gnd.n715 240.244
R5986 gnd.n7004 gnd.n715 240.244
R5987 gnd.n7004 gnd.n713 240.244
R5988 gnd.n7008 gnd.n713 240.244
R5989 gnd.n7008 gnd.n709 240.244
R5990 gnd.n7014 gnd.n709 240.244
R5991 gnd.n7014 gnd.n707 240.244
R5992 gnd.n7018 gnd.n707 240.244
R5993 gnd.n7018 gnd.n703 240.244
R5994 gnd.n7024 gnd.n703 240.244
R5995 gnd.n7024 gnd.n701 240.244
R5996 gnd.n7028 gnd.n701 240.244
R5997 gnd.n7028 gnd.n697 240.244
R5998 gnd.n7034 gnd.n697 240.244
R5999 gnd.n7034 gnd.n695 240.244
R6000 gnd.n7038 gnd.n695 240.244
R6001 gnd.n7038 gnd.n691 240.244
R6002 gnd.n7044 gnd.n691 240.244
R6003 gnd.n7044 gnd.n689 240.244
R6004 gnd.n7048 gnd.n689 240.244
R6005 gnd.n7048 gnd.n685 240.244
R6006 gnd.n7054 gnd.n685 240.244
R6007 gnd.n7054 gnd.n683 240.244
R6008 gnd.n7058 gnd.n683 240.244
R6009 gnd.n7058 gnd.n679 240.244
R6010 gnd.n7064 gnd.n679 240.244
R6011 gnd.n7064 gnd.n677 240.244
R6012 gnd.n7068 gnd.n677 240.244
R6013 gnd.n7068 gnd.n673 240.244
R6014 gnd.n7074 gnd.n673 240.244
R6015 gnd.n7074 gnd.n671 240.244
R6016 gnd.n7078 gnd.n671 240.244
R6017 gnd.n7078 gnd.n667 240.244
R6018 gnd.n7084 gnd.n667 240.244
R6019 gnd.n7084 gnd.n665 240.244
R6020 gnd.n7088 gnd.n665 240.244
R6021 gnd.n7088 gnd.n661 240.244
R6022 gnd.n7094 gnd.n661 240.244
R6023 gnd.n7094 gnd.n659 240.244
R6024 gnd.n7098 gnd.n659 240.244
R6025 gnd.n7098 gnd.n655 240.244
R6026 gnd.n7104 gnd.n655 240.244
R6027 gnd.n7104 gnd.n653 240.244
R6028 gnd.n7108 gnd.n653 240.244
R6029 gnd.n7108 gnd.n649 240.244
R6030 gnd.n7114 gnd.n649 240.244
R6031 gnd.n7114 gnd.n647 240.244
R6032 gnd.n7118 gnd.n647 240.244
R6033 gnd.n7118 gnd.n643 240.244
R6034 gnd.n7124 gnd.n643 240.244
R6035 gnd.n7124 gnd.n641 240.244
R6036 gnd.n7128 gnd.n641 240.244
R6037 gnd.n7128 gnd.n637 240.244
R6038 gnd.n7134 gnd.n637 240.244
R6039 gnd.n7134 gnd.n635 240.244
R6040 gnd.n7138 gnd.n635 240.244
R6041 gnd.n7138 gnd.n631 240.244
R6042 gnd.n7144 gnd.n631 240.244
R6043 gnd.n7144 gnd.n629 240.244
R6044 gnd.n7148 gnd.n629 240.244
R6045 gnd.n7148 gnd.n625 240.244
R6046 gnd.n7154 gnd.n625 240.244
R6047 gnd.n7154 gnd.n623 240.244
R6048 gnd.n7158 gnd.n623 240.244
R6049 gnd.n7158 gnd.n619 240.244
R6050 gnd.n7164 gnd.n619 240.244
R6051 gnd.n7164 gnd.n617 240.244
R6052 gnd.n7168 gnd.n617 240.244
R6053 gnd.n7168 gnd.n613 240.244
R6054 gnd.n7174 gnd.n613 240.244
R6055 gnd.n7174 gnd.n611 240.244
R6056 gnd.n7178 gnd.n611 240.244
R6057 gnd.n7178 gnd.n607 240.244
R6058 gnd.n7184 gnd.n607 240.244
R6059 gnd.n7184 gnd.n605 240.244
R6060 gnd.n7188 gnd.n605 240.244
R6061 gnd.n7188 gnd.n601 240.244
R6062 gnd.n7194 gnd.n601 240.244
R6063 gnd.n7194 gnd.n599 240.244
R6064 gnd.n7198 gnd.n599 240.244
R6065 gnd.n7198 gnd.n595 240.244
R6066 gnd.n7204 gnd.n595 240.244
R6067 gnd.n7204 gnd.n593 240.244
R6068 gnd.n7208 gnd.n593 240.244
R6069 gnd.n7208 gnd.n589 240.244
R6070 gnd.n7214 gnd.n589 240.244
R6071 gnd.n7214 gnd.n587 240.244
R6072 gnd.n7218 gnd.n587 240.244
R6073 gnd.n7218 gnd.n583 240.244
R6074 gnd.n7224 gnd.n583 240.244
R6075 gnd.n7224 gnd.n581 240.244
R6076 gnd.n7228 gnd.n581 240.244
R6077 gnd.n7228 gnd.n577 240.244
R6078 gnd.n7234 gnd.n577 240.244
R6079 gnd.n7234 gnd.n575 240.244
R6080 gnd.n7238 gnd.n575 240.244
R6081 gnd.n7238 gnd.n571 240.244
R6082 gnd.n7244 gnd.n571 240.244
R6083 gnd.n7244 gnd.n569 240.244
R6084 gnd.n7248 gnd.n569 240.244
R6085 gnd.n7248 gnd.n565 240.244
R6086 gnd.n7254 gnd.n565 240.244
R6087 gnd.n7254 gnd.n563 240.244
R6088 gnd.n7258 gnd.n563 240.244
R6089 gnd.n7258 gnd.n559 240.244
R6090 gnd.n7264 gnd.n559 240.244
R6091 gnd.n7264 gnd.n557 240.244
R6092 gnd.n7268 gnd.n557 240.244
R6093 gnd.n7268 gnd.n553 240.244
R6094 gnd.n7274 gnd.n553 240.244
R6095 gnd.n7274 gnd.n551 240.244
R6096 gnd.n7278 gnd.n551 240.244
R6097 gnd.n7278 gnd.n547 240.244
R6098 gnd.n7284 gnd.n547 240.244
R6099 gnd.n7284 gnd.n545 240.244
R6100 gnd.n7288 gnd.n545 240.244
R6101 gnd.n7288 gnd.n541 240.244
R6102 gnd.n7294 gnd.n541 240.244
R6103 gnd.n7294 gnd.n539 240.244
R6104 gnd.n7298 gnd.n539 240.244
R6105 gnd.n7298 gnd.n535 240.244
R6106 gnd.n7304 gnd.n535 240.244
R6107 gnd.n7304 gnd.n533 240.244
R6108 gnd.n7308 gnd.n533 240.244
R6109 gnd.n7308 gnd.n529 240.244
R6110 gnd.n7314 gnd.n529 240.244
R6111 gnd.n7314 gnd.n527 240.244
R6112 gnd.n7318 gnd.n527 240.244
R6113 gnd.n7318 gnd.n523 240.244
R6114 gnd.n7324 gnd.n523 240.244
R6115 gnd.n7324 gnd.n521 240.244
R6116 gnd.n7328 gnd.n521 240.244
R6117 gnd.n7328 gnd.n517 240.244
R6118 gnd.n7334 gnd.n517 240.244
R6119 gnd.n7334 gnd.n515 240.244
R6120 gnd.n7338 gnd.n515 240.244
R6121 gnd.n7338 gnd.n511 240.244
R6122 gnd.n7344 gnd.n511 240.244
R6123 gnd.n7344 gnd.n509 240.244
R6124 gnd.n7348 gnd.n509 240.244
R6125 gnd.n7348 gnd.n505 240.244
R6126 gnd.n7354 gnd.n505 240.244
R6127 gnd.n7354 gnd.n503 240.244
R6128 gnd.n7358 gnd.n503 240.244
R6129 gnd.n7358 gnd.n499 240.244
R6130 gnd.n7365 gnd.n499 240.244
R6131 gnd.n7365 gnd.n497 240.244
R6132 gnd.n7369 gnd.n497 240.244
R6133 gnd.n7369 gnd.n494 240.244
R6134 gnd.n7375 gnd.n492 240.244
R6135 gnd.n7379 gnd.n492 240.244
R6136 gnd.n7379 gnd.n488 240.244
R6137 gnd.n7385 gnd.n488 240.244
R6138 gnd.n7385 gnd.n486 240.244
R6139 gnd.n7389 gnd.n486 240.244
R6140 gnd.n7389 gnd.n482 240.244
R6141 gnd.n7395 gnd.n482 240.244
R6142 gnd.n7395 gnd.n480 240.244
R6143 gnd.n7399 gnd.n480 240.244
R6144 gnd.n7399 gnd.n476 240.244
R6145 gnd.n7405 gnd.n476 240.244
R6146 gnd.n7405 gnd.n474 240.244
R6147 gnd.n7409 gnd.n474 240.244
R6148 gnd.n7409 gnd.n470 240.244
R6149 gnd.n7415 gnd.n470 240.244
R6150 gnd.n7415 gnd.n468 240.244
R6151 gnd.n7419 gnd.n468 240.244
R6152 gnd.n7419 gnd.n464 240.244
R6153 gnd.n7425 gnd.n464 240.244
R6154 gnd.n7425 gnd.n462 240.244
R6155 gnd.n7429 gnd.n462 240.244
R6156 gnd.n7429 gnd.n458 240.244
R6157 gnd.n7435 gnd.n458 240.244
R6158 gnd.n7435 gnd.n456 240.244
R6159 gnd.n7439 gnd.n456 240.244
R6160 gnd.n7439 gnd.n452 240.244
R6161 gnd.n7445 gnd.n452 240.244
R6162 gnd.n7445 gnd.n450 240.244
R6163 gnd.n7449 gnd.n450 240.244
R6164 gnd.n7449 gnd.n446 240.244
R6165 gnd.n7455 gnd.n446 240.244
R6166 gnd.n7455 gnd.n444 240.244
R6167 gnd.n7459 gnd.n444 240.244
R6168 gnd.n7459 gnd.n440 240.244
R6169 gnd.n7465 gnd.n440 240.244
R6170 gnd.n7465 gnd.n438 240.244
R6171 gnd.n7469 gnd.n438 240.244
R6172 gnd.n7469 gnd.n434 240.244
R6173 gnd.n7475 gnd.n434 240.244
R6174 gnd.n7475 gnd.n432 240.244
R6175 gnd.n7479 gnd.n432 240.244
R6176 gnd.n7479 gnd.n428 240.244
R6177 gnd.n7485 gnd.n428 240.244
R6178 gnd.n7485 gnd.n426 240.244
R6179 gnd.n7489 gnd.n426 240.244
R6180 gnd.n7489 gnd.n422 240.244
R6181 gnd.n7495 gnd.n422 240.244
R6182 gnd.n7495 gnd.n420 240.244
R6183 gnd.n7499 gnd.n420 240.244
R6184 gnd.n7499 gnd.n416 240.244
R6185 gnd.n7505 gnd.n416 240.244
R6186 gnd.n7505 gnd.n414 240.244
R6187 gnd.n7509 gnd.n414 240.244
R6188 gnd.n7509 gnd.n410 240.244
R6189 gnd.n7515 gnd.n410 240.244
R6190 gnd.n7515 gnd.n408 240.244
R6191 gnd.n7519 gnd.n408 240.244
R6192 gnd.n7519 gnd.n404 240.244
R6193 gnd.n7525 gnd.n404 240.244
R6194 gnd.n7525 gnd.n402 240.244
R6195 gnd.n7529 gnd.n402 240.244
R6196 gnd.n7529 gnd.n398 240.244
R6197 gnd.n7535 gnd.n398 240.244
R6198 gnd.n7535 gnd.n396 240.244
R6199 gnd.n7539 gnd.n396 240.244
R6200 gnd.n7539 gnd.n392 240.244
R6201 gnd.n7545 gnd.n392 240.244
R6202 gnd.n7545 gnd.n390 240.244
R6203 gnd.n7549 gnd.n390 240.244
R6204 gnd.n7549 gnd.n386 240.244
R6205 gnd.n7555 gnd.n386 240.244
R6206 gnd.n7555 gnd.n384 240.244
R6207 gnd.n7559 gnd.n384 240.244
R6208 gnd.n7559 gnd.n380 240.244
R6209 gnd.n7565 gnd.n380 240.244
R6210 gnd.n7565 gnd.n378 240.244
R6211 gnd.n7569 gnd.n378 240.244
R6212 gnd.n7569 gnd.n374 240.244
R6213 gnd.n7575 gnd.n374 240.244
R6214 gnd.n7575 gnd.n372 240.244
R6215 gnd.n7580 gnd.n372 240.244
R6216 gnd.n7580 gnd.n368 240.244
R6217 gnd.n7587 gnd.n368 240.244
R6218 gnd.n4203 gnd.n4202 240.244
R6219 gnd.n4204 gnd.n4203 240.244
R6220 gnd.n4204 gnd.n4191 240.244
R6221 gnd.n4210 gnd.n4191 240.244
R6222 gnd.n4211 gnd.n4210 240.244
R6223 gnd.n4212 gnd.n4211 240.244
R6224 gnd.n4212 gnd.n4036 240.244
R6225 gnd.n4218 gnd.n4036 240.244
R6226 gnd.n4218 gnd.n4025 240.244
R6227 gnd.n4256 gnd.n4025 240.244
R6228 gnd.n4256 gnd.n4255 240.244
R6229 gnd.n4255 gnd.n4021 240.244
R6230 gnd.n4263 gnd.n4021 240.244
R6231 gnd.n4264 gnd.n4263 240.244
R6232 gnd.n4264 gnd.n4018 240.244
R6233 gnd.n4277 gnd.n4018 240.244
R6234 gnd.n4277 gnd.n4019 240.244
R6235 gnd.n4272 gnd.n4019 240.244
R6236 gnd.n4272 gnd.n4271 240.244
R6237 gnd.n4271 gnd.n3986 240.244
R6238 gnd.n4319 gnd.n3986 240.244
R6239 gnd.n4320 gnd.n4319 240.244
R6240 gnd.n4320 gnd.n3983 240.244
R6241 gnd.n4346 gnd.n3983 240.244
R6242 gnd.n4346 gnd.n3984 240.244
R6243 gnd.n4342 gnd.n3984 240.244
R6244 gnd.n4342 gnd.n4341 240.244
R6245 gnd.n4341 gnd.n4340 240.244
R6246 gnd.n4340 gnd.n4328 240.244
R6247 gnd.n4336 gnd.n4328 240.244
R6248 gnd.n4336 gnd.n3961 240.244
R6249 gnd.n4407 gnd.n3961 240.244
R6250 gnd.n4408 gnd.n4407 240.244
R6251 gnd.n4409 gnd.n4408 240.244
R6252 gnd.n4409 gnd.n3957 240.244
R6253 gnd.n4415 gnd.n3957 240.244
R6254 gnd.n4416 gnd.n4415 240.244
R6255 gnd.n4417 gnd.n4416 240.244
R6256 gnd.n4417 gnd.n3952 240.244
R6257 gnd.n4449 gnd.n3952 240.244
R6258 gnd.n4449 gnd.n3953 240.244
R6259 gnd.n4445 gnd.n3953 240.244
R6260 gnd.n4445 gnd.n4444 240.244
R6261 gnd.n4444 gnd.n4443 240.244
R6262 gnd.n4443 gnd.n4425 240.244
R6263 gnd.n4439 gnd.n4425 240.244
R6264 gnd.n4439 gnd.n4438 240.244
R6265 gnd.n4438 gnd.n4437 240.244
R6266 gnd.n4437 gnd.n3933 240.244
R6267 gnd.n4770 gnd.n3933 240.244
R6268 gnd.n4771 gnd.n4770 240.244
R6269 gnd.n4772 gnd.n4771 240.244
R6270 gnd.n4772 gnd.n3928 240.244
R6271 gnd.n4780 gnd.n3928 240.244
R6272 gnd.n4780 gnd.n3929 240.244
R6273 gnd.n3929 gnd.n3904 240.244
R6274 gnd.n4790 gnd.n3904 240.244
R6275 gnd.n4790 gnd.n3900 240.244
R6276 gnd.n4796 gnd.n3900 240.244
R6277 gnd.n4796 gnd.n3889 240.244
R6278 gnd.n4806 gnd.n3889 240.244
R6279 gnd.n4806 gnd.n3885 240.244
R6280 gnd.n4812 gnd.n3885 240.244
R6281 gnd.n4812 gnd.n3875 240.244
R6282 gnd.n4822 gnd.n3875 240.244
R6283 gnd.n4822 gnd.n3871 240.244
R6284 gnd.n4828 gnd.n3871 240.244
R6285 gnd.n4828 gnd.n3860 240.244
R6286 gnd.n4849 gnd.n3860 240.244
R6287 gnd.n4849 gnd.n3855 240.244
R6288 gnd.n4858 gnd.n3855 240.244
R6289 gnd.n4858 gnd.n3856 240.244
R6290 gnd.n3856 gnd.n2901 240.244
R6291 gnd.n6198 gnd.n2901 240.244
R6292 gnd.n6198 gnd.n2902 240.244
R6293 gnd.n6194 gnd.n2902 240.244
R6294 gnd.n6194 gnd.n2908 240.244
R6295 gnd.n3770 gnd.n2908 240.244
R6296 gnd.n3770 gnd.n3750 240.244
R6297 gnd.n4923 gnd.n3750 240.244
R6298 gnd.n4923 gnd.n3746 240.244
R6299 gnd.n4929 gnd.n3746 240.244
R6300 gnd.n4929 gnd.n3726 240.244
R6301 gnd.n4962 gnd.n3726 240.244
R6302 gnd.n4962 gnd.n3722 240.244
R6303 gnd.n4968 gnd.n3722 240.244
R6304 gnd.n4968 gnd.n3700 240.244
R6305 gnd.n5002 gnd.n3700 240.244
R6306 gnd.n5002 gnd.n3695 240.244
R6307 gnd.n5010 gnd.n3695 240.244
R6308 gnd.n5010 gnd.n3696 240.244
R6309 gnd.n3696 gnd.n3673 240.244
R6310 gnd.n5048 gnd.n3673 240.244
R6311 gnd.n5048 gnd.n3668 240.244
R6312 gnd.n5056 gnd.n3668 240.244
R6313 gnd.n5056 gnd.n3669 240.244
R6314 gnd.n3669 gnd.n3651 240.244
R6315 gnd.n5101 gnd.n3651 240.244
R6316 gnd.n5101 gnd.n3646 240.244
R6317 gnd.n5109 gnd.n3646 240.244
R6318 gnd.n5109 gnd.n3647 240.244
R6319 gnd.n3647 gnd.n3625 240.244
R6320 gnd.n5137 gnd.n3625 240.244
R6321 gnd.n5137 gnd.n3621 240.244
R6322 gnd.n5143 gnd.n3621 240.244
R6323 gnd.n5143 gnd.n3599 240.244
R6324 gnd.n5179 gnd.n3599 240.244
R6325 gnd.n5179 gnd.n3594 240.244
R6326 gnd.n5187 gnd.n3594 240.244
R6327 gnd.n5187 gnd.n3595 240.244
R6328 gnd.n3595 gnd.n3575 240.244
R6329 gnd.n5231 gnd.n3575 240.244
R6330 gnd.n5231 gnd.n3571 240.244
R6331 gnd.n5237 gnd.n3571 240.244
R6332 gnd.n5237 gnd.n3557 240.244
R6333 gnd.n5260 gnd.n3557 240.244
R6334 gnd.n5260 gnd.n3553 240.244
R6335 gnd.n5266 gnd.n3553 240.244
R6336 gnd.n5266 gnd.n3466 240.244
R6337 gnd.n5407 gnd.n3466 240.244
R6338 gnd.n5407 gnd.n3462 240.244
R6339 gnd.n5413 gnd.n3462 240.244
R6340 gnd.n5413 gnd.n3453 240.244
R6341 gnd.n5423 gnd.n3453 240.244
R6342 gnd.n5423 gnd.n3449 240.244
R6343 gnd.n5429 gnd.n3449 240.244
R6344 gnd.n5429 gnd.n3440 240.244
R6345 gnd.n5439 gnd.n3440 240.244
R6346 gnd.n5439 gnd.n3436 240.244
R6347 gnd.n5445 gnd.n3436 240.244
R6348 gnd.n5445 gnd.n3427 240.244
R6349 gnd.n5455 gnd.n3427 240.244
R6350 gnd.n5455 gnd.n3423 240.244
R6351 gnd.n5464 gnd.n3423 240.244
R6352 gnd.n5464 gnd.n3414 240.244
R6353 gnd.n5474 gnd.n3414 240.244
R6354 gnd.n5475 gnd.n5474 240.244
R6355 gnd.n5475 gnd.n2995 240.244
R6356 gnd.n3409 gnd.n2995 240.244
R6357 gnd.n5574 gnd.n3409 240.244
R6358 gnd.n5574 gnd.n3410 240.244
R6359 gnd.n5570 gnd.n3410 240.244
R6360 gnd.n5570 gnd.n5569 240.244
R6361 gnd.n5569 gnd.n5568 240.244
R6362 gnd.n5568 gnd.n5484 240.244
R6363 gnd.n5564 gnd.n5484 240.244
R6364 gnd.n5564 gnd.n5561 240.244
R6365 gnd.n5561 gnd.n5560 240.244
R6366 gnd.n5560 gnd.n5490 240.244
R6367 gnd.n5556 gnd.n5490 240.244
R6368 gnd.n5556 gnd.n5555 240.244
R6369 gnd.n5555 gnd.n5554 240.244
R6370 gnd.n5554 gnd.n5496 240.244
R6371 gnd.n5550 gnd.n5496 240.244
R6372 gnd.n5550 gnd.n5549 240.244
R6373 gnd.n5549 gnd.n5548 240.244
R6374 gnd.n5548 gnd.n5502 240.244
R6375 gnd.n5544 gnd.n5502 240.244
R6376 gnd.n5544 gnd.n5543 240.244
R6377 gnd.n5543 gnd.n5542 240.244
R6378 gnd.n5542 gnd.n5508 240.244
R6379 gnd.n5538 gnd.n5508 240.244
R6380 gnd.n5538 gnd.n5537 240.244
R6381 gnd.n5537 gnd.n5536 240.244
R6382 gnd.n5536 gnd.n5514 240.244
R6383 gnd.n5532 gnd.n5514 240.244
R6384 gnd.n5532 gnd.n5531 240.244
R6385 gnd.n5531 gnd.n5530 240.244
R6386 gnd.n5530 gnd.n5520 240.244
R6387 gnd.n5526 gnd.n5520 240.244
R6388 gnd.n5526 gnd.n3322 240.244
R6389 gnd.n5819 gnd.n3322 240.244
R6390 gnd.n5819 gnd.n3323 240.244
R6391 gnd.n5814 gnd.n3323 240.244
R6392 gnd.n5814 gnd.n3326 240.244
R6393 gnd.n5710 gnd.n3326 240.244
R6394 gnd.n5711 gnd.n5710 240.244
R6395 gnd.n5712 gnd.n5711 240.244
R6396 gnd.n5712 gnd.n5704 240.244
R6397 gnd.n5791 gnd.n5704 240.244
R6398 gnd.n5791 gnd.n5705 240.244
R6399 gnd.n5786 gnd.n5705 240.244
R6400 gnd.n5786 gnd.n5785 240.244
R6401 gnd.n5785 gnd.n5718 240.244
R6402 gnd.n5736 gnd.n5718 240.244
R6403 gnd.n5754 gnd.n5736 240.244
R6404 gnd.n5754 gnd.n5737 240.244
R6405 gnd.n5750 gnd.n5737 240.244
R6406 gnd.n5750 gnd.n5749 240.244
R6407 gnd.n5749 gnd.n361 240.244
R6408 gnd.n7594 gnd.n361 240.244
R6409 gnd.n7594 gnd.n362 240.244
R6410 gnd.n7590 gnd.n362 240.244
R6411 gnd.n7590 gnd.n7589 240.244
R6412 gnd.n6884 gnd.n787 240.244
R6413 gnd.n6880 gnd.n787 240.244
R6414 gnd.n6880 gnd.n792 240.244
R6415 gnd.n6876 gnd.n792 240.244
R6416 gnd.n6876 gnd.n794 240.244
R6417 gnd.n6872 gnd.n794 240.244
R6418 gnd.n6872 gnd.n800 240.244
R6419 gnd.n6868 gnd.n800 240.244
R6420 gnd.n6868 gnd.n802 240.244
R6421 gnd.n6864 gnd.n802 240.244
R6422 gnd.n6864 gnd.n808 240.244
R6423 gnd.n6860 gnd.n808 240.244
R6424 gnd.n6860 gnd.n810 240.244
R6425 gnd.n6856 gnd.n810 240.244
R6426 gnd.n6856 gnd.n816 240.244
R6427 gnd.n6852 gnd.n816 240.244
R6428 gnd.n6852 gnd.n818 240.244
R6429 gnd.n6848 gnd.n818 240.244
R6430 gnd.n6848 gnd.n824 240.244
R6431 gnd.n6844 gnd.n824 240.244
R6432 gnd.n6844 gnd.n826 240.244
R6433 gnd.n6840 gnd.n826 240.244
R6434 gnd.n6840 gnd.n832 240.244
R6435 gnd.n6836 gnd.n832 240.244
R6436 gnd.n6836 gnd.n834 240.244
R6437 gnd.n6832 gnd.n834 240.244
R6438 gnd.n6832 gnd.n840 240.244
R6439 gnd.n6828 gnd.n840 240.244
R6440 gnd.n6828 gnd.n842 240.244
R6441 gnd.n6824 gnd.n842 240.244
R6442 gnd.n6824 gnd.n848 240.244
R6443 gnd.n6820 gnd.n848 240.244
R6444 gnd.n6820 gnd.n850 240.244
R6445 gnd.n6816 gnd.n850 240.244
R6446 gnd.n6816 gnd.n856 240.244
R6447 gnd.n6812 gnd.n856 240.244
R6448 gnd.n6812 gnd.n858 240.244
R6449 gnd.n6808 gnd.n858 240.244
R6450 gnd.n6808 gnd.n864 240.244
R6451 gnd.n6804 gnd.n864 240.244
R6452 gnd.n6804 gnd.n866 240.244
R6453 gnd.n6800 gnd.n866 240.244
R6454 gnd.n6800 gnd.n872 240.244
R6455 gnd.n6796 gnd.n872 240.244
R6456 gnd.n6796 gnd.n874 240.244
R6457 gnd.n6792 gnd.n874 240.244
R6458 gnd.n6792 gnd.n880 240.244
R6459 gnd.n6788 gnd.n880 240.244
R6460 gnd.n6788 gnd.n882 240.244
R6461 gnd.n6784 gnd.n882 240.244
R6462 gnd.n6784 gnd.n888 240.244
R6463 gnd.n6780 gnd.n888 240.244
R6464 gnd.n6780 gnd.n890 240.244
R6465 gnd.n6776 gnd.n890 240.244
R6466 gnd.n6776 gnd.n896 240.244
R6467 gnd.n6772 gnd.n896 240.244
R6468 gnd.n6772 gnd.n898 240.244
R6469 gnd.n6768 gnd.n898 240.244
R6470 gnd.n6768 gnd.n904 240.244
R6471 gnd.n6764 gnd.n904 240.244
R6472 gnd.n6764 gnd.n906 240.244
R6473 gnd.n6760 gnd.n906 240.244
R6474 gnd.n6760 gnd.n912 240.244
R6475 gnd.n6756 gnd.n912 240.244
R6476 gnd.n6756 gnd.n914 240.244
R6477 gnd.n6752 gnd.n914 240.244
R6478 gnd.n6752 gnd.n920 240.244
R6479 gnd.n6748 gnd.n920 240.244
R6480 gnd.n6748 gnd.n922 240.244
R6481 gnd.n6744 gnd.n922 240.244
R6482 gnd.n6744 gnd.n928 240.244
R6483 gnd.n6740 gnd.n928 240.244
R6484 gnd.n6740 gnd.n930 240.244
R6485 gnd.n6736 gnd.n930 240.244
R6486 gnd.n6736 gnd.n936 240.244
R6487 gnd.n6732 gnd.n936 240.244
R6488 gnd.n6732 gnd.n938 240.244
R6489 gnd.n6728 gnd.n938 240.244
R6490 gnd.n6728 gnd.n944 240.244
R6491 gnd.n6724 gnd.n944 240.244
R6492 gnd.n6724 gnd.n946 240.244
R6493 gnd.n6720 gnd.n946 240.244
R6494 gnd.n6720 gnd.n952 240.244
R6495 gnd.n4195 gnd.n952 240.244
R6496 gnd.n4521 gnd.n3906 240.244
R6497 gnd.n4486 gnd.n3906 240.244
R6498 gnd.n4486 gnd.n3899 240.244
R6499 gnd.n4487 gnd.n3899 240.244
R6500 gnd.n4487 gnd.n3891 240.244
R6501 gnd.n4490 gnd.n3891 240.244
R6502 gnd.n4490 gnd.n3884 240.244
R6503 gnd.n4491 gnd.n3884 240.244
R6504 gnd.n4491 gnd.n3877 240.244
R6505 gnd.n4494 gnd.n3877 240.244
R6506 gnd.n4494 gnd.n3870 240.244
R6507 gnd.n4495 gnd.n3870 240.244
R6508 gnd.n4495 gnd.n3862 240.244
R6509 gnd.n3862 gnd.n3851 240.244
R6510 gnd.n4860 gnd.n3851 240.244
R6511 gnd.n4861 gnd.n4860 240.244
R6512 gnd.n4862 gnd.n4861 240.244
R6513 gnd.n4862 gnd.n2898 240.244
R6514 gnd.n4868 gnd.n2898 240.244
R6515 gnd.n4868 gnd.n2910 240.244
R6516 gnd.n4901 gnd.n2910 240.244
R6517 gnd.n4901 gnd.n3760 240.244
R6518 gnd.n4910 gnd.n3760 240.244
R6519 gnd.n4910 gnd.n3752 240.244
R6520 gnd.n3752 gnd.n3743 240.244
R6521 gnd.n4931 gnd.n3743 240.244
R6522 gnd.n4932 gnd.n4931 240.244
R6523 gnd.n4932 gnd.n3728 240.244
R6524 gnd.n4944 gnd.n3728 240.244
R6525 gnd.n4944 gnd.n3720 240.244
R6526 gnd.n4937 gnd.n3720 240.244
R6527 gnd.n4937 gnd.n3702 240.244
R6528 gnd.n3702 gnd.n3693 240.244
R6529 gnd.n5012 gnd.n3693 240.244
R6530 gnd.n5012 gnd.n3688 240.244
R6531 gnd.n5019 gnd.n3688 240.244
R6532 gnd.n5019 gnd.n3674 240.244
R6533 gnd.n3674 gnd.n3666 240.244
R6534 gnd.n5058 gnd.n3666 240.244
R6535 gnd.n5058 gnd.n3661 240.244
R6536 gnd.n5090 gnd.n3661 240.244
R6537 gnd.n5090 gnd.n3653 240.244
R6538 gnd.n5064 gnd.n3653 240.244
R6539 gnd.n5064 gnd.n3645 240.244
R6540 gnd.n5065 gnd.n3645 240.244
R6541 gnd.n5066 gnd.n5065 240.244
R6542 gnd.n5066 gnd.n3627 240.244
R6543 gnd.n5070 gnd.n3627 240.244
R6544 gnd.n5070 gnd.n3618 240.244
R6545 gnd.n5071 gnd.n3618 240.244
R6546 gnd.n5071 gnd.n3601 240.244
R6547 gnd.n3601 gnd.n3591 240.244
R6548 gnd.n5189 gnd.n3591 240.244
R6549 gnd.n5189 gnd.n3586 240.244
R6550 gnd.n5218 gnd.n3586 240.244
R6551 gnd.n5218 gnd.n3577 240.244
R6552 gnd.n5196 gnd.n3577 240.244
R6553 gnd.n5196 gnd.n3570 240.244
R6554 gnd.n5197 gnd.n3570 240.244
R6555 gnd.n5197 gnd.n3558 240.244
R6556 gnd.n5200 gnd.n3558 240.244
R6557 gnd.n5200 gnd.n3551 240.244
R6558 gnd.n5201 gnd.n3551 240.244
R6559 gnd.n5201 gnd.n3468 240.244
R6560 gnd.n3468 gnd.n3459 240.244
R6561 gnd.n5415 gnd.n3459 240.244
R6562 gnd.n5415 gnd.n3455 240.244
R6563 gnd.n5421 gnd.n3455 240.244
R6564 gnd.n5421 gnd.n3445 240.244
R6565 gnd.n5431 gnd.n3445 240.244
R6566 gnd.n5431 gnd.n3441 240.244
R6567 gnd.n5437 gnd.n3441 240.244
R6568 gnd.n5437 gnd.n3432 240.244
R6569 gnd.n5447 gnd.n3432 240.244
R6570 gnd.n5447 gnd.n3428 240.244
R6571 gnd.n5453 gnd.n3428 240.244
R6572 gnd.n5453 gnd.n3420 240.244
R6573 gnd.n5466 gnd.n3420 240.244
R6574 gnd.n5466 gnd.n3416 240.244
R6575 gnd.n5472 gnd.n3416 240.244
R6576 gnd.n5472 gnd.n2997 240.244
R6577 gnd.n6094 gnd.n2997 240.244
R6578 gnd.n4526 gnd.n4525 240.244
R6579 gnd.n4481 gnd.n4480 240.244
R6580 gnd.n4534 gnd.n4533 240.244
R6581 gnd.n4536 gnd.n4535 240.244
R6582 gnd.n4543 gnd.n4542 240.244
R6583 gnd.n4545 gnd.n4544 240.244
R6584 gnd.n4555 gnd.n4554 240.244
R6585 gnd.n4563 gnd.n4562 240.244
R6586 gnd.n4565 gnd.n4564 240.244
R6587 gnd.n4575 gnd.n4574 240.244
R6588 gnd.n4583 gnd.n4582 240.244
R6589 gnd.n4585 gnd.n4584 240.244
R6590 gnd.n4600 gnd.n4599 240.244
R6591 gnd.n4782 gnd.n3911 240.244
R6592 gnd.n4788 gnd.n3907 240.244
R6593 gnd.n4788 gnd.n3897 240.244
R6594 gnd.n4798 gnd.n3897 240.244
R6595 gnd.n4798 gnd.n3893 240.244
R6596 gnd.n4804 gnd.n3893 240.244
R6597 gnd.n4804 gnd.n3883 240.244
R6598 gnd.n4814 gnd.n3883 240.244
R6599 gnd.n4814 gnd.n3879 240.244
R6600 gnd.n4820 gnd.n3879 240.244
R6601 gnd.n4820 gnd.n3869 240.244
R6602 gnd.n4830 gnd.n3869 240.244
R6603 gnd.n4830 gnd.n3863 240.244
R6604 gnd.n4847 gnd.n3863 240.244
R6605 gnd.n4847 gnd.n3864 240.244
R6606 gnd.n3864 gnd.n3854 240.244
R6607 gnd.n4835 gnd.n3854 240.244
R6608 gnd.n4836 gnd.n4835 240.244
R6609 gnd.n4836 gnd.n2900 240.244
R6610 gnd.n2911 gnd.n2900 240.244
R6611 gnd.n6192 gnd.n2911 240.244
R6612 gnd.n6192 gnd.n2912 240.244
R6613 gnd.n2917 gnd.n2912 240.244
R6614 gnd.n2918 gnd.n2917 240.244
R6615 gnd.n2919 gnd.n2918 240.244
R6616 gnd.n4878 gnd.n2919 240.244
R6617 gnd.n4878 gnd.n2922 240.244
R6618 gnd.n2923 gnd.n2922 240.244
R6619 gnd.n2924 gnd.n2923 240.244
R6620 gnd.n4945 gnd.n2924 240.244
R6621 gnd.n4945 gnd.n2927 240.244
R6622 gnd.n2928 gnd.n2927 240.244
R6623 gnd.n2929 gnd.n2928 240.244
R6624 gnd.n4982 gnd.n2929 240.244
R6625 gnd.n4982 gnd.n2932 240.244
R6626 gnd.n2933 gnd.n2932 240.244
R6627 gnd.n2934 gnd.n2933 240.244
R6628 gnd.n5046 gnd.n2934 240.244
R6629 gnd.n5046 gnd.n2937 240.244
R6630 gnd.n2938 gnd.n2937 240.244
R6631 gnd.n2939 gnd.n2938 240.244
R6632 gnd.n5091 gnd.n2939 240.244
R6633 gnd.n5091 gnd.n2942 240.244
R6634 gnd.n2943 gnd.n2942 240.244
R6635 gnd.n2944 gnd.n2943 240.244
R6636 gnd.n3639 gnd.n2944 240.244
R6637 gnd.n3639 gnd.n2947 240.244
R6638 gnd.n2948 gnd.n2947 240.244
R6639 gnd.n2949 gnd.n2948 240.244
R6640 gnd.n3620 gnd.n2949 240.244
R6641 gnd.n3620 gnd.n2952 240.244
R6642 gnd.n2953 gnd.n2952 240.244
R6643 gnd.n2954 gnd.n2953 240.244
R6644 gnd.n3593 gnd.n2954 240.244
R6645 gnd.n3593 gnd.n2957 240.244
R6646 gnd.n2958 gnd.n2957 240.244
R6647 gnd.n2959 gnd.n2958 240.244
R6648 gnd.n5194 gnd.n2959 240.244
R6649 gnd.n5194 gnd.n2962 240.244
R6650 gnd.n2963 gnd.n2962 240.244
R6651 gnd.n2964 gnd.n2963 240.244
R6652 gnd.n3560 gnd.n2964 240.244
R6653 gnd.n3560 gnd.n2967 240.244
R6654 gnd.n2968 gnd.n2967 240.244
R6655 gnd.n2969 gnd.n2968 240.244
R6656 gnd.n3470 gnd.n2969 240.244
R6657 gnd.n3470 gnd.n2972 240.244
R6658 gnd.n2973 gnd.n2972 240.244
R6659 gnd.n2974 gnd.n2973 240.244
R6660 gnd.n3446 gnd.n2974 240.244
R6661 gnd.n3446 gnd.n2977 240.244
R6662 gnd.n2978 gnd.n2977 240.244
R6663 gnd.n2979 gnd.n2978 240.244
R6664 gnd.n3433 gnd.n2979 240.244
R6665 gnd.n3433 gnd.n2982 240.244
R6666 gnd.n2983 gnd.n2982 240.244
R6667 gnd.n2984 gnd.n2983 240.244
R6668 gnd.n3421 gnd.n2984 240.244
R6669 gnd.n3421 gnd.n2987 240.244
R6670 gnd.n2988 gnd.n2987 240.244
R6671 gnd.n2989 gnd.n2988 240.244
R6672 gnd.n2992 gnd.n2989 240.244
R6673 gnd.n6096 gnd.n2992 240.244
R6674 gnd.n3003 gnd.n3002 240.244
R6675 gnd.n3387 gnd.n3006 240.244
R6676 gnd.n3008 gnd.n3007 240.244
R6677 gnd.n3390 gnd.n3012 240.244
R6678 gnd.n3393 gnd.n3013 240.244
R6679 gnd.n3022 gnd.n3021 240.244
R6680 gnd.n3395 gnd.n3029 240.244
R6681 gnd.n3398 gnd.n3030 240.244
R6682 gnd.n3038 gnd.n3037 240.244
R6683 gnd.n3400 gnd.n3045 240.244
R6684 gnd.n3403 gnd.n3046 240.244
R6685 gnd.n3054 gnd.n3053 240.244
R6686 gnd.n3406 gnd.n3385 240.244
R6687 gnd.n5577 gnd.n2993 240.244
R6688 gnd.n2880 gnd.n2879 240.132
R6689 gnd.n3486 gnd.n3485 240.132
R6690 gnd.n6887 gnd.n6886 225.874
R6691 gnd.n6887 gnd.n780 225.874
R6692 gnd.n6895 gnd.n780 225.874
R6693 gnd.n6896 gnd.n6895 225.874
R6694 gnd.n6897 gnd.n6896 225.874
R6695 gnd.n6897 gnd.n774 225.874
R6696 gnd.n6905 gnd.n774 225.874
R6697 gnd.n6906 gnd.n6905 225.874
R6698 gnd.n6907 gnd.n6906 225.874
R6699 gnd.n6907 gnd.n768 225.874
R6700 gnd.n6915 gnd.n768 225.874
R6701 gnd.n6916 gnd.n6915 225.874
R6702 gnd.n6917 gnd.n6916 225.874
R6703 gnd.n6917 gnd.n762 225.874
R6704 gnd.n6925 gnd.n762 225.874
R6705 gnd.n6926 gnd.n6925 225.874
R6706 gnd.n6927 gnd.n6926 225.874
R6707 gnd.n6927 gnd.n756 225.874
R6708 gnd.n6935 gnd.n756 225.874
R6709 gnd.n6936 gnd.n6935 225.874
R6710 gnd.n6937 gnd.n6936 225.874
R6711 gnd.n6937 gnd.n750 225.874
R6712 gnd.n6945 gnd.n750 225.874
R6713 gnd.n6946 gnd.n6945 225.874
R6714 gnd.n6947 gnd.n6946 225.874
R6715 gnd.n6947 gnd.n744 225.874
R6716 gnd.n6955 gnd.n744 225.874
R6717 gnd.n6956 gnd.n6955 225.874
R6718 gnd.n6957 gnd.n6956 225.874
R6719 gnd.n6957 gnd.n738 225.874
R6720 gnd.n6965 gnd.n738 225.874
R6721 gnd.n6966 gnd.n6965 225.874
R6722 gnd.n6967 gnd.n6966 225.874
R6723 gnd.n6967 gnd.n732 225.874
R6724 gnd.n6975 gnd.n732 225.874
R6725 gnd.n6976 gnd.n6975 225.874
R6726 gnd.n6977 gnd.n6976 225.874
R6727 gnd.n6977 gnd.n726 225.874
R6728 gnd.n6985 gnd.n726 225.874
R6729 gnd.n6986 gnd.n6985 225.874
R6730 gnd.n6987 gnd.n6986 225.874
R6731 gnd.n6987 gnd.n720 225.874
R6732 gnd.n6995 gnd.n720 225.874
R6733 gnd.n6996 gnd.n6995 225.874
R6734 gnd.n6997 gnd.n6996 225.874
R6735 gnd.n6997 gnd.n714 225.874
R6736 gnd.n7005 gnd.n714 225.874
R6737 gnd.n7006 gnd.n7005 225.874
R6738 gnd.n7007 gnd.n7006 225.874
R6739 gnd.n7007 gnd.n708 225.874
R6740 gnd.n7015 gnd.n708 225.874
R6741 gnd.n7016 gnd.n7015 225.874
R6742 gnd.n7017 gnd.n7016 225.874
R6743 gnd.n7017 gnd.n702 225.874
R6744 gnd.n7025 gnd.n702 225.874
R6745 gnd.n7026 gnd.n7025 225.874
R6746 gnd.n7027 gnd.n7026 225.874
R6747 gnd.n7027 gnd.n696 225.874
R6748 gnd.n7035 gnd.n696 225.874
R6749 gnd.n7036 gnd.n7035 225.874
R6750 gnd.n7037 gnd.n7036 225.874
R6751 gnd.n7037 gnd.n690 225.874
R6752 gnd.n7045 gnd.n690 225.874
R6753 gnd.n7046 gnd.n7045 225.874
R6754 gnd.n7047 gnd.n7046 225.874
R6755 gnd.n7047 gnd.n684 225.874
R6756 gnd.n7055 gnd.n684 225.874
R6757 gnd.n7056 gnd.n7055 225.874
R6758 gnd.n7057 gnd.n7056 225.874
R6759 gnd.n7057 gnd.n678 225.874
R6760 gnd.n7065 gnd.n678 225.874
R6761 gnd.n7066 gnd.n7065 225.874
R6762 gnd.n7067 gnd.n7066 225.874
R6763 gnd.n7067 gnd.n672 225.874
R6764 gnd.n7075 gnd.n672 225.874
R6765 gnd.n7076 gnd.n7075 225.874
R6766 gnd.n7077 gnd.n7076 225.874
R6767 gnd.n7077 gnd.n666 225.874
R6768 gnd.n7085 gnd.n666 225.874
R6769 gnd.n7086 gnd.n7085 225.874
R6770 gnd.n7087 gnd.n7086 225.874
R6771 gnd.n7087 gnd.n660 225.874
R6772 gnd.n7095 gnd.n660 225.874
R6773 gnd.n7096 gnd.n7095 225.874
R6774 gnd.n7097 gnd.n7096 225.874
R6775 gnd.n7097 gnd.n654 225.874
R6776 gnd.n7105 gnd.n654 225.874
R6777 gnd.n7106 gnd.n7105 225.874
R6778 gnd.n7107 gnd.n7106 225.874
R6779 gnd.n7107 gnd.n648 225.874
R6780 gnd.n7115 gnd.n648 225.874
R6781 gnd.n7116 gnd.n7115 225.874
R6782 gnd.n7117 gnd.n7116 225.874
R6783 gnd.n7117 gnd.n642 225.874
R6784 gnd.n7125 gnd.n642 225.874
R6785 gnd.n7126 gnd.n7125 225.874
R6786 gnd.n7127 gnd.n7126 225.874
R6787 gnd.n7127 gnd.n636 225.874
R6788 gnd.n7135 gnd.n636 225.874
R6789 gnd.n7136 gnd.n7135 225.874
R6790 gnd.n7137 gnd.n7136 225.874
R6791 gnd.n7137 gnd.n630 225.874
R6792 gnd.n7145 gnd.n630 225.874
R6793 gnd.n7146 gnd.n7145 225.874
R6794 gnd.n7147 gnd.n7146 225.874
R6795 gnd.n7147 gnd.n624 225.874
R6796 gnd.n7155 gnd.n624 225.874
R6797 gnd.n7156 gnd.n7155 225.874
R6798 gnd.n7157 gnd.n7156 225.874
R6799 gnd.n7157 gnd.n618 225.874
R6800 gnd.n7165 gnd.n618 225.874
R6801 gnd.n7166 gnd.n7165 225.874
R6802 gnd.n7167 gnd.n7166 225.874
R6803 gnd.n7167 gnd.n612 225.874
R6804 gnd.n7175 gnd.n612 225.874
R6805 gnd.n7176 gnd.n7175 225.874
R6806 gnd.n7177 gnd.n7176 225.874
R6807 gnd.n7177 gnd.n606 225.874
R6808 gnd.n7185 gnd.n606 225.874
R6809 gnd.n7186 gnd.n7185 225.874
R6810 gnd.n7187 gnd.n7186 225.874
R6811 gnd.n7187 gnd.n600 225.874
R6812 gnd.n7195 gnd.n600 225.874
R6813 gnd.n7196 gnd.n7195 225.874
R6814 gnd.n7197 gnd.n7196 225.874
R6815 gnd.n7197 gnd.n594 225.874
R6816 gnd.n7205 gnd.n594 225.874
R6817 gnd.n7206 gnd.n7205 225.874
R6818 gnd.n7207 gnd.n7206 225.874
R6819 gnd.n7207 gnd.n588 225.874
R6820 gnd.n7215 gnd.n588 225.874
R6821 gnd.n7216 gnd.n7215 225.874
R6822 gnd.n7217 gnd.n7216 225.874
R6823 gnd.n7217 gnd.n582 225.874
R6824 gnd.n7225 gnd.n582 225.874
R6825 gnd.n7226 gnd.n7225 225.874
R6826 gnd.n7227 gnd.n7226 225.874
R6827 gnd.n7227 gnd.n576 225.874
R6828 gnd.n7235 gnd.n576 225.874
R6829 gnd.n7236 gnd.n7235 225.874
R6830 gnd.n7237 gnd.n7236 225.874
R6831 gnd.n7237 gnd.n570 225.874
R6832 gnd.n7245 gnd.n570 225.874
R6833 gnd.n7246 gnd.n7245 225.874
R6834 gnd.n7247 gnd.n7246 225.874
R6835 gnd.n7247 gnd.n564 225.874
R6836 gnd.n7255 gnd.n564 225.874
R6837 gnd.n7256 gnd.n7255 225.874
R6838 gnd.n7257 gnd.n7256 225.874
R6839 gnd.n7257 gnd.n558 225.874
R6840 gnd.n7265 gnd.n558 225.874
R6841 gnd.n7266 gnd.n7265 225.874
R6842 gnd.n7267 gnd.n7266 225.874
R6843 gnd.n7267 gnd.n552 225.874
R6844 gnd.n7275 gnd.n552 225.874
R6845 gnd.n7276 gnd.n7275 225.874
R6846 gnd.n7277 gnd.n7276 225.874
R6847 gnd.n7277 gnd.n546 225.874
R6848 gnd.n7285 gnd.n546 225.874
R6849 gnd.n7286 gnd.n7285 225.874
R6850 gnd.n7287 gnd.n7286 225.874
R6851 gnd.n7287 gnd.n540 225.874
R6852 gnd.n7295 gnd.n540 225.874
R6853 gnd.n7296 gnd.n7295 225.874
R6854 gnd.n7297 gnd.n7296 225.874
R6855 gnd.n7297 gnd.n534 225.874
R6856 gnd.n7305 gnd.n534 225.874
R6857 gnd.n7306 gnd.n7305 225.874
R6858 gnd.n7307 gnd.n7306 225.874
R6859 gnd.n7307 gnd.n528 225.874
R6860 gnd.n7315 gnd.n528 225.874
R6861 gnd.n7316 gnd.n7315 225.874
R6862 gnd.n7317 gnd.n7316 225.874
R6863 gnd.n7317 gnd.n522 225.874
R6864 gnd.n7325 gnd.n522 225.874
R6865 gnd.n7326 gnd.n7325 225.874
R6866 gnd.n7327 gnd.n7326 225.874
R6867 gnd.n7327 gnd.n516 225.874
R6868 gnd.n7335 gnd.n516 225.874
R6869 gnd.n7336 gnd.n7335 225.874
R6870 gnd.n7337 gnd.n7336 225.874
R6871 gnd.n7337 gnd.n510 225.874
R6872 gnd.n7345 gnd.n510 225.874
R6873 gnd.n7346 gnd.n7345 225.874
R6874 gnd.n7347 gnd.n7346 225.874
R6875 gnd.n7347 gnd.n504 225.874
R6876 gnd.n7355 gnd.n504 225.874
R6877 gnd.n7356 gnd.n7355 225.874
R6878 gnd.n7357 gnd.n7356 225.874
R6879 gnd.n7357 gnd.n498 225.874
R6880 gnd.n7366 gnd.n498 225.874
R6881 gnd.n7367 gnd.n7366 225.874
R6882 gnd.n7368 gnd.n7367 225.874
R6883 gnd.n7368 gnd.n493 225.874
R6884 gnd.n1569 gnd.t173 224.174
R6885 gnd.n1033 gnd.t282 224.174
R6886 gnd.n3138 gnd.n3075 199.319
R6887 gnd.n3138 gnd.n3076 199.319
R6888 gnd.n2833 gnd.n2793 199.319
R6889 gnd.n2833 gnd.n2792 199.319
R6890 gnd.n2881 gnd.n2878 186.49
R6891 gnd.n3487 gnd.n3484 186.49
R6892 gnd.n2325 gnd.n2324 185
R6893 gnd.n2323 gnd.n2322 185
R6894 gnd.n2302 gnd.n2301 185
R6895 gnd.n2317 gnd.n2316 185
R6896 gnd.n2315 gnd.n2314 185
R6897 gnd.n2306 gnd.n2305 185
R6898 gnd.n2309 gnd.n2308 185
R6899 gnd.n2293 gnd.n2292 185
R6900 gnd.n2291 gnd.n2290 185
R6901 gnd.n2270 gnd.n2269 185
R6902 gnd.n2285 gnd.n2284 185
R6903 gnd.n2283 gnd.n2282 185
R6904 gnd.n2274 gnd.n2273 185
R6905 gnd.n2277 gnd.n2276 185
R6906 gnd.n2261 gnd.n2260 185
R6907 gnd.n2259 gnd.n2258 185
R6908 gnd.n2238 gnd.n2237 185
R6909 gnd.n2253 gnd.n2252 185
R6910 gnd.n2251 gnd.n2250 185
R6911 gnd.n2242 gnd.n2241 185
R6912 gnd.n2245 gnd.n2244 185
R6913 gnd.n2230 gnd.n2229 185
R6914 gnd.n2228 gnd.n2227 185
R6915 gnd.n2207 gnd.n2206 185
R6916 gnd.n2222 gnd.n2221 185
R6917 gnd.n2220 gnd.n2219 185
R6918 gnd.n2211 gnd.n2210 185
R6919 gnd.n2214 gnd.n2213 185
R6920 gnd.n2198 gnd.n2197 185
R6921 gnd.n2196 gnd.n2195 185
R6922 gnd.n2175 gnd.n2174 185
R6923 gnd.n2190 gnd.n2189 185
R6924 gnd.n2188 gnd.n2187 185
R6925 gnd.n2179 gnd.n2178 185
R6926 gnd.n2182 gnd.n2181 185
R6927 gnd.n2166 gnd.n2165 185
R6928 gnd.n2164 gnd.n2163 185
R6929 gnd.n2143 gnd.n2142 185
R6930 gnd.n2158 gnd.n2157 185
R6931 gnd.n2156 gnd.n2155 185
R6932 gnd.n2147 gnd.n2146 185
R6933 gnd.n2150 gnd.n2149 185
R6934 gnd.n2134 gnd.n2133 185
R6935 gnd.n2132 gnd.n2131 185
R6936 gnd.n2111 gnd.n2110 185
R6937 gnd.n2126 gnd.n2125 185
R6938 gnd.n2124 gnd.n2123 185
R6939 gnd.n2115 gnd.n2114 185
R6940 gnd.n2118 gnd.n2117 185
R6941 gnd.n2103 gnd.n2102 185
R6942 gnd.n2101 gnd.n2100 185
R6943 gnd.n2080 gnd.n2079 185
R6944 gnd.n2095 gnd.n2094 185
R6945 gnd.n2093 gnd.n2092 185
R6946 gnd.n2084 gnd.n2083 185
R6947 gnd.n2087 gnd.n2086 185
R6948 gnd.n1570 gnd.t172 178.987
R6949 gnd.n1034 gnd.t283 178.987
R6950 gnd.n1 gnd.t311 170.774
R6951 gnd.n7 gnd.t333 170.103
R6952 gnd.n6 gnd.t145 170.103
R6953 gnd.n5 gnd.t339 170.103
R6954 gnd.n4 gnd.t75 170.103
R6955 gnd.n3 gnd.t37 170.103
R6956 gnd.n2 gnd.t341 170.103
R6957 gnd.n1 gnd.t116 170.103
R6958 gnd.n5397 gnd.n5396 163.367
R6959 gnd.n5394 gnd.n3496 163.367
R6960 gnd.n5390 gnd.n5389 163.367
R6961 gnd.n5387 gnd.n3499 163.367
R6962 gnd.n5383 gnd.n5382 163.367
R6963 gnd.n5380 gnd.n3502 163.367
R6964 gnd.n5376 gnd.n5375 163.367
R6965 gnd.n5373 gnd.n3505 163.367
R6966 gnd.n5369 gnd.n5368 163.367
R6967 gnd.n5366 gnd.n3508 163.367
R6968 gnd.n5362 gnd.n5361 163.367
R6969 gnd.n5359 gnd.n3511 163.367
R6970 gnd.n5355 gnd.n5354 163.367
R6971 gnd.n5352 gnd.n3514 163.367
R6972 gnd.n5347 gnd.n5346 163.367
R6973 gnd.n5344 gnd.n5342 163.367
R6974 gnd.n5339 gnd.n5338 163.367
R6975 gnd.n5336 gnd.n3520 163.367
R6976 gnd.n5331 gnd.n5330 163.367
R6977 gnd.n5328 gnd.n3525 163.367
R6978 gnd.n5324 gnd.n5323 163.367
R6979 gnd.n5321 gnd.n3528 163.367
R6980 gnd.n5317 gnd.n5316 163.367
R6981 gnd.n5314 gnd.n3531 163.367
R6982 gnd.n5310 gnd.n5309 163.367
R6983 gnd.n5307 gnd.n3534 163.367
R6984 gnd.n5303 gnd.n5302 163.367
R6985 gnd.n5300 gnd.n3537 163.367
R6986 gnd.n5296 gnd.n5295 163.367
R6987 gnd.n5293 gnd.n3540 163.367
R6988 gnd.n5289 gnd.n5288 163.367
R6989 gnd.n5286 gnd.n3543 163.367
R6990 gnd.n3843 gnd.n2897 163.367
R6991 gnd.n3847 gnd.n2897 163.367
R6992 gnd.n4873 gnd.n3847 163.367
R6993 gnd.n4873 gnd.n3775 163.367
R6994 gnd.n4892 gnd.n3775 163.367
R6995 gnd.n4892 gnd.n3776 163.367
R6996 gnd.n3776 gnd.n3766 163.367
R6997 gnd.n4887 gnd.n3766 163.367
R6998 gnd.n4887 gnd.n3759 163.367
R6999 gnd.n4884 gnd.n3759 163.367
R7000 gnd.n4884 gnd.n3753 163.367
R7001 gnd.n4881 gnd.n3753 163.367
R7002 gnd.n4881 gnd.n4877 163.367
R7003 gnd.n4877 gnd.n3734 163.367
R7004 gnd.n4953 gnd.n3734 163.367
R7005 gnd.n4953 gnd.n3735 163.367
R7006 gnd.n3735 gnd.n3729 163.367
R7007 gnd.n4948 gnd.n3729 163.367
R7008 gnd.n4948 gnd.n3719 163.367
R7009 gnd.n3719 gnd.n3714 163.367
R7010 gnd.n4977 gnd.n3714 163.367
R7011 gnd.n4978 gnd.n4977 163.367
R7012 gnd.n4978 gnd.n3703 163.367
R7013 gnd.n4985 gnd.n3703 163.367
R7014 gnd.n4986 gnd.n4985 163.367
R7015 gnd.n4986 gnd.n3712 163.367
R7016 gnd.n4990 gnd.n3712 163.367
R7017 gnd.n4990 gnd.n3686 163.367
R7018 gnd.n5022 gnd.n3686 163.367
R7019 gnd.n5022 gnd.n3675 163.367
R7020 gnd.n3683 gnd.n3675 163.367
R7021 gnd.n5038 gnd.n3683 163.367
R7022 gnd.n5038 gnd.n3684 163.367
R7023 gnd.n5034 gnd.n3684 163.367
R7024 gnd.n5034 gnd.n3660 163.367
R7025 gnd.n5030 gnd.n3660 163.367
R7026 gnd.n5030 gnd.n3654 163.367
R7027 gnd.n5027 gnd.n3654 163.367
R7028 gnd.n5027 gnd.n3644 163.367
R7029 gnd.n3644 gnd.n3636 163.367
R7030 gnd.n5118 gnd.n3636 163.367
R7031 gnd.n5118 gnd.n3633 163.367
R7032 gnd.n5128 gnd.n3633 163.367
R7033 gnd.n5128 gnd.n3634 163.367
R7034 gnd.n3634 gnd.n3628 163.367
R7035 gnd.n5123 gnd.n3628 163.367
R7036 gnd.n5123 gnd.n3617 163.367
R7037 gnd.n3617 gnd.n3611 163.367
R7038 gnd.n5152 gnd.n3611 163.367
R7039 gnd.n5153 gnd.n5152 163.367
R7040 gnd.n5153 gnd.n3602 163.367
R7041 gnd.n5157 gnd.n3602 163.367
R7042 gnd.n5157 gnd.n3608 163.367
R7043 gnd.n5168 gnd.n3608 163.367
R7044 gnd.n5168 gnd.n3609 163.367
R7045 gnd.n3609 gnd.n3585 163.367
R7046 gnd.n5163 gnd.n3585 163.367
R7047 gnd.n5163 gnd.n3578 163.367
R7048 gnd.n5160 gnd.n3578 163.367
R7049 gnd.n5160 gnd.n3568 163.367
R7050 gnd.n5240 gnd.n3568 163.367
R7051 gnd.n5240 gnd.n3566 163.367
R7052 gnd.n5250 gnd.n3566 163.367
R7053 gnd.n5250 gnd.n3559 163.367
R7054 gnd.n5246 gnd.n3559 163.367
R7055 gnd.n5246 gnd.n3550 163.367
R7056 gnd.n3550 gnd.n3545 163.367
R7057 gnd.n5275 gnd.n3545 163.367
R7058 gnd.n5276 gnd.n5275 163.367
R7059 gnd.n5276 gnd.n3469 163.367
R7060 gnd.n5281 gnd.n3469 163.367
R7061 gnd.n2872 gnd.n2871 163.367
R7062 gnd.n6263 gnd.n2871 163.367
R7063 gnd.n6261 gnd.n6260 163.367
R7064 gnd.n6257 gnd.n6256 163.367
R7065 gnd.n6253 gnd.n6252 163.367
R7066 gnd.n6249 gnd.n6248 163.367
R7067 gnd.n6245 gnd.n6244 163.367
R7068 gnd.n6241 gnd.n6240 163.367
R7069 gnd.n6237 gnd.n6236 163.367
R7070 gnd.n6233 gnd.n6232 163.367
R7071 gnd.n6229 gnd.n6228 163.367
R7072 gnd.n6225 gnd.n6224 163.367
R7073 gnd.n6221 gnd.n6220 163.367
R7074 gnd.n6217 gnd.n6216 163.367
R7075 gnd.n6213 gnd.n6212 163.367
R7076 gnd.n6209 gnd.n6208 163.367
R7077 gnd.n6272 gnd.n2838 163.367
R7078 gnd.n3781 gnd.n3780 163.367
R7079 gnd.n3786 gnd.n3785 163.367
R7080 gnd.n3790 gnd.n3789 163.367
R7081 gnd.n3794 gnd.n3793 163.367
R7082 gnd.n3798 gnd.n3797 163.367
R7083 gnd.n3802 gnd.n3801 163.367
R7084 gnd.n3806 gnd.n3805 163.367
R7085 gnd.n3810 gnd.n3809 163.367
R7086 gnd.n3814 gnd.n3813 163.367
R7087 gnd.n3818 gnd.n3817 163.367
R7088 gnd.n3822 gnd.n3821 163.367
R7089 gnd.n3826 gnd.n3825 163.367
R7090 gnd.n3830 gnd.n3829 163.367
R7091 gnd.n3834 gnd.n3833 163.367
R7092 gnd.n3838 gnd.n3837 163.367
R7093 gnd.n6201 gnd.n2873 163.367
R7094 gnd.n6201 gnd.n2895 163.367
R7095 gnd.n4871 gnd.n2895 163.367
R7096 gnd.n4871 gnd.n3774 163.367
R7097 gnd.n4894 gnd.n3774 163.367
R7098 gnd.n4894 gnd.n3772 163.367
R7099 gnd.n4898 gnd.n3772 163.367
R7100 gnd.n4898 gnd.n3757 163.367
R7101 gnd.n4913 gnd.n3757 163.367
R7102 gnd.n4913 gnd.n3754 163.367
R7103 gnd.n4920 gnd.n3754 163.367
R7104 gnd.n4920 gnd.n3755 163.367
R7105 gnd.n4916 gnd.n3755 163.367
R7106 gnd.n4916 gnd.n3732 163.367
R7107 gnd.n4955 gnd.n3732 163.367
R7108 gnd.n4955 gnd.n3730 163.367
R7109 gnd.n4959 gnd.n3730 163.367
R7110 gnd.n4959 gnd.n3718 163.367
R7111 gnd.n4971 gnd.n3718 163.367
R7112 gnd.n4971 gnd.n3716 163.367
R7113 gnd.n4975 gnd.n3716 163.367
R7114 gnd.n4975 gnd.n3704 163.367
R7115 gnd.n4999 gnd.n3704 163.367
R7116 gnd.n4999 gnd.n3705 163.367
R7117 gnd.n4995 gnd.n3705 163.367
R7118 gnd.n4995 gnd.n4994 163.367
R7119 gnd.n4994 gnd.n3711 163.367
R7120 gnd.n3711 gnd.n3708 163.367
R7121 gnd.n3708 gnd.n3677 163.367
R7122 gnd.n5044 gnd.n3677 163.367
R7123 gnd.n5044 gnd.n3678 163.367
R7124 gnd.n5040 gnd.n3678 163.367
R7125 gnd.n5040 gnd.n3681 163.367
R7126 gnd.n3681 gnd.n3658 163.367
R7127 gnd.n5094 gnd.n3658 163.367
R7128 gnd.n5094 gnd.n3656 163.367
R7129 gnd.n5098 gnd.n3656 163.367
R7130 gnd.n5098 gnd.n3643 163.367
R7131 gnd.n5112 gnd.n3643 163.367
R7132 gnd.n5112 gnd.n3641 163.367
R7133 gnd.n5116 gnd.n3641 163.367
R7134 gnd.n5116 gnd.n3631 163.367
R7135 gnd.n5130 gnd.n3631 163.367
R7136 gnd.n5130 gnd.n3629 163.367
R7137 gnd.n5134 gnd.n3629 163.367
R7138 gnd.n5134 gnd.n3615 163.367
R7139 gnd.n5146 gnd.n3615 163.367
R7140 gnd.n5146 gnd.n3613 163.367
R7141 gnd.n5150 gnd.n3613 163.367
R7142 gnd.n5150 gnd.n3604 163.367
R7143 gnd.n5176 gnd.n3604 163.367
R7144 gnd.n5176 gnd.n3605 163.367
R7145 gnd.n5172 gnd.n3605 163.367
R7146 gnd.n5172 gnd.n5171 163.367
R7147 gnd.n5171 gnd.n3583 163.367
R7148 gnd.n5221 gnd.n3583 163.367
R7149 gnd.n5221 gnd.n3580 163.367
R7150 gnd.n5228 gnd.n3580 163.367
R7151 gnd.n5228 gnd.n3581 163.367
R7152 gnd.n5224 gnd.n3581 163.367
R7153 gnd.n5224 gnd.n3564 163.367
R7154 gnd.n5253 gnd.n3564 163.367
R7155 gnd.n5253 gnd.n3562 163.367
R7156 gnd.n5257 gnd.n3562 163.367
R7157 gnd.n5257 gnd.n3549 163.367
R7158 gnd.n5269 gnd.n3549 163.367
R7159 gnd.n5269 gnd.n3547 163.367
R7160 gnd.n5273 gnd.n3547 163.367
R7161 gnd.n5273 gnd.n3472 163.367
R7162 gnd.n5404 gnd.n3472 163.367
R7163 gnd.n5404 gnd.n3473 163.367
R7164 gnd.n3493 gnd.n3492 156.462
R7165 gnd.n2265 gnd.n2233 153.042
R7166 gnd.n2329 gnd.n2328 152.079
R7167 gnd.n2297 gnd.n2296 152.079
R7168 gnd.n2265 gnd.n2264 152.079
R7169 gnd.n2886 gnd.n2885 152
R7170 gnd.n2887 gnd.n2876 152
R7171 gnd.n2889 gnd.n2888 152
R7172 gnd.n2891 gnd.n2874 152
R7173 gnd.n2893 gnd.n2892 152
R7174 gnd.n3491 gnd.n3475 152
R7175 gnd.n3483 gnd.n3476 152
R7176 gnd.n3482 gnd.n3481 152
R7177 gnd.n3480 gnd.n3477 152
R7178 gnd.n3478 gnd.t189 150.546
R7179 gnd.n7377 gnd.n7376 150.119
R7180 gnd.n7378 gnd.n7377 150.119
R7181 gnd.n7378 gnd.n487 150.119
R7182 gnd.n7386 gnd.n487 150.119
R7183 gnd.n7387 gnd.n7386 150.119
R7184 gnd.n7388 gnd.n7387 150.119
R7185 gnd.n7388 gnd.n481 150.119
R7186 gnd.n7396 gnd.n481 150.119
R7187 gnd.n7397 gnd.n7396 150.119
R7188 gnd.n7398 gnd.n7397 150.119
R7189 gnd.n7398 gnd.n475 150.119
R7190 gnd.n7406 gnd.n475 150.119
R7191 gnd.n7407 gnd.n7406 150.119
R7192 gnd.n7408 gnd.n7407 150.119
R7193 gnd.n7408 gnd.n469 150.119
R7194 gnd.n7416 gnd.n469 150.119
R7195 gnd.n7417 gnd.n7416 150.119
R7196 gnd.n7418 gnd.n7417 150.119
R7197 gnd.n7418 gnd.n463 150.119
R7198 gnd.n7426 gnd.n463 150.119
R7199 gnd.n7427 gnd.n7426 150.119
R7200 gnd.n7428 gnd.n7427 150.119
R7201 gnd.n7428 gnd.n457 150.119
R7202 gnd.n7436 gnd.n457 150.119
R7203 gnd.n7437 gnd.n7436 150.119
R7204 gnd.n7438 gnd.n7437 150.119
R7205 gnd.n7438 gnd.n451 150.119
R7206 gnd.n7446 gnd.n451 150.119
R7207 gnd.n7447 gnd.n7446 150.119
R7208 gnd.n7448 gnd.n7447 150.119
R7209 gnd.n7448 gnd.n445 150.119
R7210 gnd.n7456 gnd.n445 150.119
R7211 gnd.n7457 gnd.n7456 150.119
R7212 gnd.n7458 gnd.n7457 150.119
R7213 gnd.n7458 gnd.n439 150.119
R7214 gnd.n7466 gnd.n439 150.119
R7215 gnd.n7467 gnd.n7466 150.119
R7216 gnd.n7468 gnd.n7467 150.119
R7217 gnd.n7468 gnd.n433 150.119
R7218 gnd.n7476 gnd.n433 150.119
R7219 gnd.n7477 gnd.n7476 150.119
R7220 gnd.n7478 gnd.n7477 150.119
R7221 gnd.n7478 gnd.n427 150.119
R7222 gnd.n7486 gnd.n427 150.119
R7223 gnd.n7487 gnd.n7486 150.119
R7224 gnd.n7488 gnd.n7487 150.119
R7225 gnd.n7488 gnd.n421 150.119
R7226 gnd.n7496 gnd.n421 150.119
R7227 gnd.n7497 gnd.n7496 150.119
R7228 gnd.n7498 gnd.n7497 150.119
R7229 gnd.n7498 gnd.n415 150.119
R7230 gnd.n7506 gnd.n415 150.119
R7231 gnd.n7507 gnd.n7506 150.119
R7232 gnd.n7508 gnd.n7507 150.119
R7233 gnd.n7508 gnd.n409 150.119
R7234 gnd.n7516 gnd.n409 150.119
R7235 gnd.n7517 gnd.n7516 150.119
R7236 gnd.n7518 gnd.n7517 150.119
R7237 gnd.n7518 gnd.n403 150.119
R7238 gnd.n7526 gnd.n403 150.119
R7239 gnd.n7527 gnd.n7526 150.119
R7240 gnd.n7528 gnd.n7527 150.119
R7241 gnd.n7528 gnd.n397 150.119
R7242 gnd.n7536 gnd.n397 150.119
R7243 gnd.n7537 gnd.n7536 150.119
R7244 gnd.n7538 gnd.n7537 150.119
R7245 gnd.n7538 gnd.n391 150.119
R7246 gnd.n7546 gnd.n391 150.119
R7247 gnd.n7547 gnd.n7546 150.119
R7248 gnd.n7548 gnd.n7547 150.119
R7249 gnd.n7548 gnd.n385 150.119
R7250 gnd.n7556 gnd.n385 150.119
R7251 gnd.n7557 gnd.n7556 150.119
R7252 gnd.n7558 gnd.n7557 150.119
R7253 gnd.n7558 gnd.n379 150.119
R7254 gnd.n7566 gnd.n379 150.119
R7255 gnd.n7567 gnd.n7566 150.119
R7256 gnd.n7568 gnd.n7567 150.119
R7257 gnd.n7568 gnd.n373 150.119
R7258 gnd.n7576 gnd.n373 150.119
R7259 gnd.n7577 gnd.n7576 150.119
R7260 gnd.n7579 gnd.n7577 150.119
R7261 gnd.n7579 gnd.n7578 150.119
R7262 gnd.t141 gnd.n2307 147.661
R7263 gnd.t349 gnd.n2275 147.661
R7264 gnd.t13 gnd.n2243 147.661
R7265 gnd.t150 gnd.n2212 147.661
R7266 gnd.t390 gnd.n2180 147.661
R7267 gnd.t327 gnd.n2148 147.661
R7268 gnd.t392 gnd.n2116 147.661
R7269 gnd.t368 gnd.n2085 147.661
R7270 gnd.n5341 gnd.n5340 143.351
R7271 gnd.n2853 gnd.n2837 143.351
R7272 gnd.n6271 gnd.n2837 143.351
R7273 gnd.n5974 gnd.n3137 131.649
R7274 gnd.n6274 gnd.n6273 131.649
R7275 gnd.n2883 gnd.t240 130.484
R7276 gnd.n2892 gnd.t203 126.766
R7277 gnd.n2890 gnd.t167 126.766
R7278 gnd.n2876 gnd.t213 126.766
R7279 gnd.n2884 gnd.t284 126.766
R7280 gnd.n3479 gnd.t186 126.766
R7281 gnd.n3481 gnd.t246 126.766
R7282 gnd.n3490 gnd.t234 126.766
R7283 gnd.n3492 gnd.t268 126.766
R7284 gnd.n2324 gnd.n2323 104.615
R7285 gnd.n2323 gnd.n2301 104.615
R7286 gnd.n2316 gnd.n2301 104.615
R7287 gnd.n2316 gnd.n2315 104.615
R7288 gnd.n2315 gnd.n2305 104.615
R7289 gnd.n2308 gnd.n2305 104.615
R7290 gnd.n2292 gnd.n2291 104.615
R7291 gnd.n2291 gnd.n2269 104.615
R7292 gnd.n2284 gnd.n2269 104.615
R7293 gnd.n2284 gnd.n2283 104.615
R7294 gnd.n2283 gnd.n2273 104.615
R7295 gnd.n2276 gnd.n2273 104.615
R7296 gnd.n2260 gnd.n2259 104.615
R7297 gnd.n2259 gnd.n2237 104.615
R7298 gnd.n2252 gnd.n2237 104.615
R7299 gnd.n2252 gnd.n2251 104.615
R7300 gnd.n2251 gnd.n2241 104.615
R7301 gnd.n2244 gnd.n2241 104.615
R7302 gnd.n2229 gnd.n2228 104.615
R7303 gnd.n2228 gnd.n2206 104.615
R7304 gnd.n2221 gnd.n2206 104.615
R7305 gnd.n2221 gnd.n2220 104.615
R7306 gnd.n2220 gnd.n2210 104.615
R7307 gnd.n2213 gnd.n2210 104.615
R7308 gnd.n2197 gnd.n2196 104.615
R7309 gnd.n2196 gnd.n2174 104.615
R7310 gnd.n2189 gnd.n2174 104.615
R7311 gnd.n2189 gnd.n2188 104.615
R7312 gnd.n2188 gnd.n2178 104.615
R7313 gnd.n2181 gnd.n2178 104.615
R7314 gnd.n2165 gnd.n2164 104.615
R7315 gnd.n2164 gnd.n2142 104.615
R7316 gnd.n2157 gnd.n2142 104.615
R7317 gnd.n2157 gnd.n2156 104.615
R7318 gnd.n2156 gnd.n2146 104.615
R7319 gnd.n2149 gnd.n2146 104.615
R7320 gnd.n2133 gnd.n2132 104.615
R7321 gnd.n2132 gnd.n2110 104.615
R7322 gnd.n2125 gnd.n2110 104.615
R7323 gnd.n2125 gnd.n2124 104.615
R7324 gnd.n2124 gnd.n2114 104.615
R7325 gnd.n2117 gnd.n2114 104.615
R7326 gnd.n2102 gnd.n2101 104.615
R7327 gnd.n2101 gnd.n2079 104.615
R7328 gnd.n2094 gnd.n2079 104.615
R7329 gnd.n2094 gnd.n2093 104.615
R7330 gnd.n2093 gnd.n2083 104.615
R7331 gnd.n2086 gnd.n2083 104.615
R7332 gnd.n1495 gnd.t223 100.632
R7333 gnd.n1012 gnd.t257 100.632
R7334 gnd.n7852 gnd.n7851 99.6594
R7335 gnd.n7847 gnd.n294 99.6594
R7336 gnd.n7843 gnd.n293 99.6594
R7337 gnd.n7839 gnd.n292 99.6594
R7338 gnd.n7835 gnd.n291 99.6594
R7339 gnd.n7831 gnd.n290 99.6594
R7340 gnd.n7827 gnd.n289 99.6594
R7341 gnd.n7823 gnd.n288 99.6594
R7342 gnd.n7816 gnd.n287 99.6594
R7343 gnd.n7812 gnd.n286 99.6594
R7344 gnd.n7808 gnd.n285 99.6594
R7345 gnd.n7804 gnd.n284 99.6594
R7346 gnd.n7800 gnd.n283 99.6594
R7347 gnd.n7796 gnd.n282 99.6594
R7348 gnd.n7792 gnd.n281 99.6594
R7349 gnd.n7788 gnd.n280 99.6594
R7350 gnd.n7784 gnd.n279 99.6594
R7351 gnd.n7780 gnd.n278 99.6594
R7352 gnd.n7772 gnd.n277 99.6594
R7353 gnd.n7770 gnd.n276 99.6594
R7354 gnd.n7766 gnd.n275 99.6594
R7355 gnd.n7762 gnd.n274 99.6594
R7356 gnd.n7758 gnd.n273 99.6594
R7357 gnd.n7754 gnd.n272 99.6594
R7358 gnd.n7750 gnd.n271 99.6594
R7359 gnd.n7746 gnd.n270 99.6594
R7360 gnd.n7742 gnd.n269 99.6594
R7361 gnd.n7738 gnd.n268 99.6594
R7362 gnd.n7729 gnd.n267 99.6594
R7363 gnd.n6026 gnd.n6025 99.6594
R7364 gnd.n6020 gnd.n3064 99.6594
R7365 gnd.n6017 gnd.n3065 99.6594
R7366 gnd.n6013 gnd.n3066 99.6594
R7367 gnd.n6009 gnd.n3067 99.6594
R7368 gnd.n6005 gnd.n3068 99.6594
R7369 gnd.n6001 gnd.n3069 99.6594
R7370 gnd.n5997 gnd.n3070 99.6594
R7371 gnd.n5993 gnd.n3071 99.6594
R7372 gnd.n5988 gnd.n3072 99.6594
R7373 gnd.n5984 gnd.n3073 99.6594
R7374 gnd.n5980 gnd.n3074 99.6594
R7375 gnd.n5976 gnd.n3075 99.6594
R7376 gnd.n5971 gnd.n3077 99.6594
R7377 gnd.n5967 gnd.n3078 99.6594
R7378 gnd.n5963 gnd.n3079 99.6594
R7379 gnd.n5959 gnd.n3080 99.6594
R7380 gnd.n5955 gnd.n3081 99.6594
R7381 gnd.n5951 gnd.n3082 99.6594
R7382 gnd.n5947 gnd.n3083 99.6594
R7383 gnd.n5943 gnd.n3084 99.6594
R7384 gnd.n5939 gnd.n3085 99.6594
R7385 gnd.n5935 gnd.n3086 99.6594
R7386 gnd.n5931 gnd.n3087 99.6594
R7387 gnd.n5927 gnd.n3088 99.6594
R7388 gnd.n5923 gnd.n3089 99.6594
R7389 gnd.n5919 gnd.n3090 99.6594
R7390 gnd.n5915 gnd.n3091 99.6594
R7391 gnd.n6323 gnd.n6322 99.6594
R7392 gnd.n6318 gnd.n2804 99.6594
R7393 gnd.n6314 gnd.n2803 99.6594
R7394 gnd.n6310 gnd.n2802 99.6594
R7395 gnd.n6306 gnd.n2801 99.6594
R7396 gnd.n6302 gnd.n2800 99.6594
R7397 gnd.n6298 gnd.n2799 99.6594
R7398 gnd.n6294 gnd.n2798 99.6594
R7399 gnd.n6289 gnd.n2797 99.6594
R7400 gnd.n6285 gnd.n2796 99.6594
R7401 gnd.n6281 gnd.n2795 99.6594
R7402 gnd.n6277 gnd.n2794 99.6594
R7403 gnd.n4680 gnd.n2792 99.6594
R7404 gnd.n4684 gnd.n2791 99.6594
R7405 gnd.n4690 gnd.n2790 99.6594
R7406 gnd.n4694 gnd.n2789 99.6594
R7407 gnd.n4699 gnd.n2788 99.6594
R7408 gnd.n4703 gnd.n2787 99.6594
R7409 gnd.n4709 gnd.n2786 99.6594
R7410 gnd.n4713 gnd.n2785 99.6594
R7411 gnd.n4719 gnd.n2784 99.6594
R7412 gnd.n4723 gnd.n2783 99.6594
R7413 gnd.n4729 gnd.n2782 99.6594
R7414 gnd.n4733 gnd.n2781 99.6594
R7415 gnd.n4739 gnd.n2780 99.6594
R7416 gnd.n4743 gnd.n2779 99.6594
R7417 gnd.n4748 gnd.n2778 99.6594
R7418 gnd.n4751 gnd.n2777 99.6594
R7419 gnd.n6624 gnd.n6623 99.6594
R7420 gnd.n6618 gnd.n2356 99.6594
R7421 gnd.n6615 gnd.n2357 99.6594
R7422 gnd.n6611 gnd.n2358 99.6594
R7423 gnd.n6607 gnd.n2359 99.6594
R7424 gnd.n6603 gnd.n2360 99.6594
R7425 gnd.n6599 gnd.n2361 99.6594
R7426 gnd.n6595 gnd.n2362 99.6594
R7427 gnd.n6591 gnd.n2363 99.6594
R7428 gnd.n6586 gnd.n2364 99.6594
R7429 gnd.n6582 gnd.n2365 99.6594
R7430 gnd.n6578 gnd.n2366 99.6594
R7431 gnd.n6574 gnd.n2367 99.6594
R7432 gnd.n6570 gnd.n2368 99.6594
R7433 gnd.n6566 gnd.n2369 99.6594
R7434 gnd.n6562 gnd.n2370 99.6594
R7435 gnd.n6558 gnd.n2371 99.6594
R7436 gnd.n6554 gnd.n2372 99.6594
R7437 gnd.n6550 gnd.n2373 99.6594
R7438 gnd.n6546 gnd.n2374 99.6594
R7439 gnd.n6542 gnd.n2375 99.6594
R7440 gnd.n6538 gnd.n2376 99.6594
R7441 gnd.n6534 gnd.n2377 99.6594
R7442 gnd.n6530 gnd.n2378 99.6594
R7443 gnd.n6526 gnd.n2379 99.6594
R7444 gnd.n6522 gnd.n2380 99.6594
R7445 gnd.n6518 gnd.n2381 99.6594
R7446 gnd.n6514 gnd.n2382 99.6594
R7447 gnd.n6510 gnd.n2383 99.6594
R7448 gnd.n6663 gnd.n6631 99.6594
R7449 gnd.n6661 gnd.n6630 99.6594
R7450 gnd.n6657 gnd.n6629 99.6594
R7451 gnd.n6653 gnd.n6628 99.6594
R7452 gnd.n6649 gnd.n6627 99.6594
R7453 gnd.n6645 gnd.n6626 99.6594
R7454 gnd.n6675 gnd.n6673 99.6594
R7455 gnd.n6681 gnd.n1011 99.6594
R7456 gnd.n1707 gnd.n1438 99.6594
R7457 gnd.n1464 gnd.n1445 99.6594
R7458 gnd.n1466 gnd.n1446 99.6594
R7459 gnd.n1474 gnd.n1447 99.6594
R7460 gnd.n1476 gnd.n1448 99.6594
R7461 gnd.n1484 gnd.n1449 99.6594
R7462 gnd.n1486 gnd.n1450 99.6594
R7463 gnd.n1494 gnd.n1451 99.6594
R7464 gnd.n7634 gnd.n258 99.6594
R7465 gnd.n7638 gnd.n259 99.6594
R7466 gnd.n7644 gnd.n260 99.6594
R7467 gnd.n7648 gnd.n261 99.6594
R7468 gnd.n7654 gnd.n262 99.6594
R7469 gnd.n7658 gnd.n263 99.6594
R7470 gnd.n7664 gnd.n264 99.6594
R7471 gnd.n7668 gnd.n265 99.6594
R7472 gnd.n7674 gnd.n266 99.6594
R7473 gnd.n3176 gnd.n3092 99.6594
R7474 gnd.n3094 gnd.n3018 99.6594
R7475 gnd.n3095 gnd.n3025 99.6594
R7476 gnd.n3097 gnd.n3096 99.6594
R7477 gnd.n3099 gnd.n3034 99.6594
R7478 gnd.n3100 gnd.n3041 99.6594
R7479 gnd.n3102 gnd.n3101 99.6594
R7480 gnd.n3104 gnd.n3050 99.6594
R7481 gnd.n6028 gnd.n3059 99.6594
R7482 gnd.n1053 gnd.n1018 99.6594
R7483 gnd.n1057 gnd.n1019 99.6594
R7484 gnd.n1063 gnd.n1020 99.6594
R7485 gnd.n1067 gnd.n1021 99.6594
R7486 gnd.n1073 gnd.n1022 99.6594
R7487 gnd.n1077 gnd.n1023 99.6594
R7488 gnd.n1083 gnd.n1024 99.6594
R7489 gnd.n1087 gnd.n1025 99.6594
R7490 gnd.n1093 gnd.n1026 99.6594
R7491 gnd.n1097 gnd.n1027 99.6594
R7492 gnd.n1103 gnd.n1028 99.6594
R7493 gnd.n1106 gnd.n1029 99.6594
R7494 gnd.n2355 gnd.n2354 99.6594
R7495 gnd.n1622 gnd.n1621 99.6594
R7496 gnd.n1616 gnd.n1533 99.6594
R7497 gnd.n1613 gnd.n1534 99.6594
R7498 gnd.n1609 gnd.n1535 99.6594
R7499 gnd.n1605 gnd.n1536 99.6594
R7500 gnd.n1601 gnd.n1537 99.6594
R7501 gnd.n1597 gnd.n1538 99.6594
R7502 gnd.n1593 gnd.n1539 99.6594
R7503 gnd.n1589 gnd.n1540 99.6594
R7504 gnd.n1585 gnd.n1541 99.6594
R7505 gnd.n1581 gnd.n1542 99.6594
R7506 gnd.n1577 gnd.n1543 99.6594
R7507 gnd.n1624 gnd.n1532 99.6594
R7508 gnd.n4548 gnd.n2767 99.6594
R7509 gnd.n4550 gnd.n2768 99.6594
R7510 gnd.n4558 gnd.n2769 99.6594
R7511 gnd.n4568 gnd.n2770 99.6594
R7512 gnd.n4570 gnd.n2771 99.6594
R7513 gnd.n4578 gnd.n2772 99.6594
R7514 gnd.n4588 gnd.n2773 99.6594
R7515 gnd.n4590 gnd.n2774 99.6594
R7516 gnd.n3936 gnd.n2775 99.6594
R7517 gnd.n4092 gnd.n2384 99.6594
R7518 gnd.n4096 gnd.n2385 99.6594
R7519 gnd.n4102 gnd.n2386 99.6594
R7520 gnd.n4106 gnd.n2387 99.6594
R7521 gnd.n4112 gnd.n2388 99.6594
R7522 gnd.n4116 gnd.n2389 99.6594
R7523 gnd.n4122 gnd.n2390 99.6594
R7524 gnd.n4126 gnd.n2391 99.6594
R7525 gnd.n4083 gnd.n2392 99.6594
R7526 gnd.n4095 gnd.n2384 99.6594
R7527 gnd.n4101 gnd.n2385 99.6594
R7528 gnd.n4105 gnd.n2386 99.6594
R7529 gnd.n4111 gnd.n2387 99.6594
R7530 gnd.n4115 gnd.n2388 99.6594
R7531 gnd.n4121 gnd.n2389 99.6594
R7532 gnd.n4125 gnd.n2390 99.6594
R7533 gnd.n4082 gnd.n2391 99.6594
R7534 gnd.n4078 gnd.n2392 99.6594
R7535 gnd.n4593 gnd.n2775 99.6594
R7536 gnd.n4589 gnd.n2774 99.6594
R7537 gnd.n4579 gnd.n2773 99.6594
R7538 gnd.n4571 gnd.n2772 99.6594
R7539 gnd.n4569 gnd.n2771 99.6594
R7540 gnd.n4559 gnd.n2770 99.6594
R7541 gnd.n4551 gnd.n2769 99.6594
R7542 gnd.n4549 gnd.n2768 99.6594
R7543 gnd.n4539 gnd.n2767 99.6594
R7544 gnd.n1622 gnd.n1545 99.6594
R7545 gnd.n1614 gnd.n1533 99.6594
R7546 gnd.n1610 gnd.n1534 99.6594
R7547 gnd.n1606 gnd.n1535 99.6594
R7548 gnd.n1602 gnd.n1536 99.6594
R7549 gnd.n1598 gnd.n1537 99.6594
R7550 gnd.n1594 gnd.n1538 99.6594
R7551 gnd.n1590 gnd.n1539 99.6594
R7552 gnd.n1586 gnd.n1540 99.6594
R7553 gnd.n1582 gnd.n1541 99.6594
R7554 gnd.n1578 gnd.n1542 99.6594
R7555 gnd.n1574 gnd.n1543 99.6594
R7556 gnd.n1625 gnd.n1624 99.6594
R7557 gnd.n2355 gnd.n1030 99.6594
R7558 gnd.n1104 gnd.n1029 99.6594
R7559 gnd.n1096 gnd.n1028 99.6594
R7560 gnd.n1094 gnd.n1027 99.6594
R7561 gnd.n1086 gnd.n1026 99.6594
R7562 gnd.n1084 gnd.n1025 99.6594
R7563 gnd.n1076 gnd.n1024 99.6594
R7564 gnd.n1074 gnd.n1023 99.6594
R7565 gnd.n1066 gnd.n1022 99.6594
R7566 gnd.n1064 gnd.n1021 99.6594
R7567 gnd.n1056 gnd.n1020 99.6594
R7568 gnd.n1054 gnd.n1019 99.6594
R7569 gnd.n1046 gnd.n1018 99.6594
R7570 gnd.n3092 gnd.n3017 99.6594
R7571 gnd.n3094 gnd.n3093 99.6594
R7572 gnd.n3095 gnd.n3026 99.6594
R7573 gnd.n3097 gnd.n3033 99.6594
R7574 gnd.n3099 gnd.n3098 99.6594
R7575 gnd.n3100 gnd.n3042 99.6594
R7576 gnd.n3102 gnd.n3049 99.6594
R7577 gnd.n3104 gnd.n3103 99.6594
R7578 gnd.n6029 gnd.n6028 99.6594
R7579 gnd.n7667 gnd.n266 99.6594
R7580 gnd.n7665 gnd.n265 99.6594
R7581 gnd.n7657 gnd.n264 99.6594
R7582 gnd.n7655 gnd.n263 99.6594
R7583 gnd.n7647 gnd.n262 99.6594
R7584 gnd.n7645 gnd.n261 99.6594
R7585 gnd.n7637 gnd.n260 99.6594
R7586 gnd.n7635 gnd.n259 99.6594
R7587 gnd.n7629 gnd.n258 99.6594
R7588 gnd.n1708 gnd.n1707 99.6594
R7589 gnd.n1467 gnd.n1445 99.6594
R7590 gnd.n1473 gnd.n1446 99.6594
R7591 gnd.n1477 gnd.n1447 99.6594
R7592 gnd.n1483 gnd.n1448 99.6594
R7593 gnd.n1487 gnd.n1449 99.6594
R7594 gnd.n1493 gnd.n1450 99.6594
R7595 gnd.n1451 gnd.n1435 99.6594
R7596 gnd.n6674 gnd.n1011 99.6594
R7597 gnd.n6673 gnd.n1017 99.6594
R7598 gnd.n6648 gnd.n6626 99.6594
R7599 gnd.n6652 gnd.n6627 99.6594
R7600 gnd.n6656 gnd.n6628 99.6594
R7601 gnd.n6660 gnd.n6629 99.6594
R7602 gnd.n6664 gnd.n6630 99.6594
R7603 gnd.n6632 gnd.n6631 99.6594
R7604 gnd.n6624 gnd.n2396 99.6594
R7605 gnd.n6616 gnd.n2356 99.6594
R7606 gnd.n6612 gnd.n2357 99.6594
R7607 gnd.n6608 gnd.n2358 99.6594
R7608 gnd.n6604 gnd.n2359 99.6594
R7609 gnd.n6600 gnd.n2360 99.6594
R7610 gnd.n6596 gnd.n2361 99.6594
R7611 gnd.n6592 gnd.n2362 99.6594
R7612 gnd.n6587 gnd.n2363 99.6594
R7613 gnd.n6583 gnd.n2364 99.6594
R7614 gnd.n6579 gnd.n2365 99.6594
R7615 gnd.n6575 gnd.n2366 99.6594
R7616 gnd.n6571 gnd.n2367 99.6594
R7617 gnd.n6567 gnd.n2368 99.6594
R7618 gnd.n6563 gnd.n2369 99.6594
R7619 gnd.n6559 gnd.n2370 99.6594
R7620 gnd.n6555 gnd.n2371 99.6594
R7621 gnd.n6551 gnd.n2372 99.6594
R7622 gnd.n6547 gnd.n2373 99.6594
R7623 gnd.n6543 gnd.n2374 99.6594
R7624 gnd.n6539 gnd.n2375 99.6594
R7625 gnd.n6535 gnd.n2376 99.6594
R7626 gnd.n6531 gnd.n2377 99.6594
R7627 gnd.n6527 gnd.n2378 99.6594
R7628 gnd.n6523 gnd.n2379 99.6594
R7629 gnd.n6519 gnd.n2380 99.6594
R7630 gnd.n6515 gnd.n2381 99.6594
R7631 gnd.n6511 gnd.n2382 99.6594
R7632 gnd.n2466 gnd.n2383 99.6594
R7633 gnd.n4661 gnd.n2777 99.6594
R7634 gnd.n4742 gnd.n2778 99.6594
R7635 gnd.n4740 gnd.n2779 99.6594
R7636 gnd.n4732 gnd.n2780 99.6594
R7637 gnd.n4730 gnd.n2781 99.6594
R7638 gnd.n4722 gnd.n2782 99.6594
R7639 gnd.n4720 gnd.n2783 99.6594
R7640 gnd.n4712 gnd.n2784 99.6594
R7641 gnd.n4710 gnd.n2785 99.6594
R7642 gnd.n4702 gnd.n2786 99.6594
R7643 gnd.n4674 gnd.n2787 99.6594
R7644 gnd.n4693 gnd.n2788 99.6594
R7645 gnd.n4691 gnd.n2789 99.6594
R7646 gnd.n4683 gnd.n2790 99.6594
R7647 gnd.n4681 gnd.n2791 99.6594
R7648 gnd.n6276 gnd.n2793 99.6594
R7649 gnd.n6280 gnd.n2794 99.6594
R7650 gnd.n6284 gnd.n2795 99.6594
R7651 gnd.n6288 gnd.n2796 99.6594
R7652 gnd.n6293 gnd.n2797 99.6594
R7653 gnd.n6297 gnd.n2798 99.6594
R7654 gnd.n6301 gnd.n2799 99.6594
R7655 gnd.n6305 gnd.n2800 99.6594
R7656 gnd.n6309 gnd.n2801 99.6594
R7657 gnd.n6313 gnd.n2802 99.6594
R7658 gnd.n6317 gnd.n2803 99.6594
R7659 gnd.n2805 gnd.n2804 99.6594
R7660 gnd.n6323 gnd.n2764 99.6594
R7661 gnd.n6026 gnd.n3107 99.6594
R7662 gnd.n6018 gnd.n3064 99.6594
R7663 gnd.n6014 gnd.n3065 99.6594
R7664 gnd.n6010 gnd.n3066 99.6594
R7665 gnd.n6006 gnd.n3067 99.6594
R7666 gnd.n6002 gnd.n3068 99.6594
R7667 gnd.n5998 gnd.n3069 99.6594
R7668 gnd.n5994 gnd.n3070 99.6594
R7669 gnd.n5989 gnd.n3071 99.6594
R7670 gnd.n5985 gnd.n3072 99.6594
R7671 gnd.n5981 gnd.n3073 99.6594
R7672 gnd.n5977 gnd.n3074 99.6594
R7673 gnd.n5972 gnd.n3076 99.6594
R7674 gnd.n5968 gnd.n3077 99.6594
R7675 gnd.n5964 gnd.n3078 99.6594
R7676 gnd.n5960 gnd.n3079 99.6594
R7677 gnd.n5956 gnd.n3080 99.6594
R7678 gnd.n5952 gnd.n3081 99.6594
R7679 gnd.n5948 gnd.n3082 99.6594
R7680 gnd.n5944 gnd.n3083 99.6594
R7681 gnd.n5940 gnd.n3084 99.6594
R7682 gnd.n5936 gnd.n3085 99.6594
R7683 gnd.n5932 gnd.n3086 99.6594
R7684 gnd.n5928 gnd.n3087 99.6594
R7685 gnd.n5924 gnd.n3088 99.6594
R7686 gnd.n5920 gnd.n3089 99.6594
R7687 gnd.n5916 gnd.n3090 99.6594
R7688 gnd.n5908 gnd.n3091 99.6594
R7689 gnd.n7737 gnd.n267 99.6594
R7690 gnd.n7741 gnd.n268 99.6594
R7691 gnd.n7745 gnd.n269 99.6594
R7692 gnd.n7749 gnd.n270 99.6594
R7693 gnd.n7753 gnd.n271 99.6594
R7694 gnd.n7757 gnd.n272 99.6594
R7695 gnd.n7761 gnd.n273 99.6594
R7696 gnd.n7765 gnd.n274 99.6594
R7697 gnd.n7769 gnd.n275 99.6594
R7698 gnd.n7773 gnd.n276 99.6594
R7699 gnd.n7779 gnd.n277 99.6594
R7700 gnd.n7783 gnd.n278 99.6594
R7701 gnd.n7787 gnd.n279 99.6594
R7702 gnd.n7791 gnd.n280 99.6594
R7703 gnd.n7795 gnd.n281 99.6594
R7704 gnd.n7799 gnd.n282 99.6594
R7705 gnd.n7803 gnd.n283 99.6594
R7706 gnd.n7807 gnd.n284 99.6594
R7707 gnd.n7811 gnd.n285 99.6594
R7708 gnd.n7815 gnd.n286 99.6594
R7709 gnd.n7822 gnd.n287 99.6594
R7710 gnd.n7826 gnd.n288 99.6594
R7711 gnd.n7830 gnd.n289 99.6594
R7712 gnd.n7834 gnd.n290 99.6594
R7713 gnd.n7838 gnd.n291 99.6594
R7714 gnd.n7842 gnd.n292 99.6594
R7715 gnd.n7846 gnd.n293 99.6594
R7716 gnd.n295 gnd.n294 99.6594
R7717 gnd.n7852 gnd.n255 99.6594
R7718 gnd.n4522 gnd.n3913 99.6594
R7719 gnd.n4526 gnd.n3914 99.6594
R7720 gnd.n4481 gnd.n3915 99.6594
R7721 gnd.n4534 gnd.n3916 99.6594
R7722 gnd.n4536 gnd.n3917 99.6594
R7723 gnd.n4543 gnd.n3918 99.6594
R7724 gnd.n4545 gnd.n3919 99.6594
R7725 gnd.n4555 gnd.n3920 99.6594
R7726 gnd.n4563 gnd.n3921 99.6594
R7727 gnd.n4565 gnd.n3922 99.6594
R7728 gnd.n4575 gnd.n3923 99.6594
R7729 gnd.n4583 gnd.n3924 99.6594
R7730 gnd.n4585 gnd.n3925 99.6594
R7731 gnd.n4600 gnd.n3926 99.6594
R7732 gnd.n4525 gnd.n3913 99.6594
R7733 gnd.n4480 gnd.n3914 99.6594
R7734 gnd.n4533 gnd.n3915 99.6594
R7735 gnd.n4535 gnd.n3916 99.6594
R7736 gnd.n4542 gnd.n3917 99.6594
R7737 gnd.n4544 gnd.n3918 99.6594
R7738 gnd.n4554 gnd.n3919 99.6594
R7739 gnd.n4562 gnd.n3920 99.6594
R7740 gnd.n4564 gnd.n3921 99.6594
R7741 gnd.n4574 gnd.n3922 99.6594
R7742 gnd.n4582 gnd.n3923 99.6594
R7743 gnd.n4584 gnd.n3924 99.6594
R7744 gnd.n4599 gnd.n3925 99.6594
R7745 gnd.n3926 gnd.n3911 99.6594
R7746 gnd.n3386 gnd.n2998 99.6594
R7747 gnd.n3388 gnd.n3003 99.6594
R7748 gnd.n3389 gnd.n3006 99.6594
R7749 gnd.n3391 gnd.n3008 99.6594
R7750 gnd.n3392 gnd.n3012 99.6594
R7751 gnd.n3394 gnd.n3393 99.6594
R7752 gnd.n3396 gnd.n3022 99.6594
R7753 gnd.n3397 gnd.n3029 99.6594
R7754 gnd.n3399 gnd.n3398 99.6594
R7755 gnd.n3401 gnd.n3038 99.6594
R7756 gnd.n3402 gnd.n3045 99.6594
R7757 gnd.n3404 gnd.n3403 99.6594
R7758 gnd.n3407 gnd.n3054 99.6594
R7759 gnd.n5576 gnd.n3385 99.6594
R7760 gnd.n3404 gnd.n3053 99.6594
R7761 gnd.n3402 gnd.n3046 99.6594
R7762 gnd.n3401 gnd.n3400 99.6594
R7763 gnd.n3399 gnd.n3037 99.6594
R7764 gnd.n3397 gnd.n3030 99.6594
R7765 gnd.n3396 gnd.n3395 99.6594
R7766 gnd.n3394 gnd.n3021 99.6594
R7767 gnd.n3392 gnd.n3013 99.6594
R7768 gnd.n3391 gnd.n3390 99.6594
R7769 gnd.n3389 gnd.n3007 99.6594
R7770 gnd.n3388 gnd.n3387 99.6594
R7771 gnd.n3386 gnd.n3002 99.6594
R7772 gnd.n5577 gnd.n5576 99.6594
R7773 gnd.n3407 gnd.n3406 99.6594
R7774 gnd.n4596 gnd.t230 98.63
R7775 gnd.n6030 gnd.t261 98.63
R7776 gnd.n4591 gnd.t272 98.63
R7777 gnd.n3127 gnd.t254 98.63
R7778 gnd.n3150 gnd.t239 98.63
R7779 gnd.n5910 gnd.t177 98.63
R7780 gnd.n352 gnd.t278 98.63
R7781 gnd.n332 gnd.t184 98.63
R7782 gnd.n7818 gnd.t211 98.63
R7783 gnd.n7618 gnd.t232 98.63
R7784 gnd.n2416 gnd.t245 98.63
R7785 gnd.n2438 gnd.t181 98.63
R7786 gnd.n2460 gnd.t202 98.63
R7787 gnd.n4079 gnd.t276 98.63
R7788 gnd.n2822 gnd.t263 98.63
R7789 gnd.n4659 gnd.t198 98.63
R7790 gnd.n4672 gnd.t225 98.63
R7791 gnd.n3055 gnd.t208 98.63
R7792 gnd.n3777 gnd.t195 92.8196
R7793 gnd.n3521 gnd.t218 92.8196
R7794 gnd.n6205 gnd.t251 92.8118
R7795 gnd.n3515 gnd.t266 92.8118
R7796 gnd.n7578 gnd.n256 90.0721
R7797 gnd.n2883 gnd.n2882 81.8399
R7798 gnd.n1496 gnd.t222 74.8376
R7799 gnd.n1013 gnd.t258 74.8376
R7800 gnd.n3778 gnd.t194 72.8438
R7801 gnd.n3522 gnd.t219 72.8438
R7802 gnd.n2884 gnd.n2877 72.8411
R7803 gnd.n2890 gnd.n2875 72.8411
R7804 gnd.n3490 gnd.n3489 72.8411
R7805 gnd.n4597 gnd.t229 72.836
R7806 gnd.n6206 gnd.t250 72.836
R7807 gnd.n3516 gnd.t267 72.836
R7808 gnd.n6031 gnd.t260 72.836
R7809 gnd.n4592 gnd.t273 72.836
R7810 gnd.n3128 gnd.t253 72.836
R7811 gnd.n3151 gnd.t238 72.836
R7812 gnd.n5911 gnd.t176 72.836
R7813 gnd.n353 gnd.t279 72.836
R7814 gnd.n333 gnd.t185 72.836
R7815 gnd.n7819 gnd.t212 72.836
R7816 gnd.n7619 gnd.t233 72.836
R7817 gnd.n2417 gnd.t244 72.836
R7818 gnd.n2439 gnd.t180 72.836
R7819 gnd.n2461 gnd.t201 72.836
R7820 gnd.n4080 gnd.t275 72.836
R7821 gnd.n2823 gnd.t264 72.836
R7822 gnd.n4660 gnd.t199 72.836
R7823 gnd.n4673 gnd.t226 72.836
R7824 gnd.n3056 gnd.t209 72.836
R7825 gnd.n5398 gnd.n5397 71.676
R7826 gnd.n5395 gnd.n5394 71.676
R7827 gnd.n5390 gnd.n3498 71.676
R7828 gnd.n5388 gnd.n5387 71.676
R7829 gnd.n5383 gnd.n3501 71.676
R7830 gnd.n5381 gnd.n5380 71.676
R7831 gnd.n5376 gnd.n3504 71.676
R7832 gnd.n5374 gnd.n5373 71.676
R7833 gnd.n5369 gnd.n3507 71.676
R7834 gnd.n5367 gnd.n5366 71.676
R7835 gnd.n5362 gnd.n3510 71.676
R7836 gnd.n5360 gnd.n5359 71.676
R7837 gnd.n5355 gnd.n3513 71.676
R7838 gnd.n5353 gnd.n5352 71.676
R7839 gnd.n5347 gnd.n3518 71.676
R7840 gnd.n5345 gnd.n5344 71.676
R7841 gnd.n5340 gnd.n5339 71.676
R7842 gnd.n5337 gnd.n5336 71.676
R7843 gnd.n5331 gnd.n3524 71.676
R7844 gnd.n5329 gnd.n5328 71.676
R7845 gnd.n5324 gnd.n3527 71.676
R7846 gnd.n5322 gnd.n5321 71.676
R7847 gnd.n5317 gnd.n3530 71.676
R7848 gnd.n5315 gnd.n5314 71.676
R7849 gnd.n5310 gnd.n3533 71.676
R7850 gnd.n5308 gnd.n5307 71.676
R7851 gnd.n5303 gnd.n3536 71.676
R7852 gnd.n5301 gnd.n5300 71.676
R7853 gnd.n5296 gnd.n3539 71.676
R7854 gnd.n5294 gnd.n5293 71.676
R7855 gnd.n5289 gnd.n3542 71.676
R7856 gnd.n5287 gnd.n5286 71.676
R7857 gnd.n5282 gnd.n5280 71.676
R7858 gnd.n6269 gnd.n6268 71.676
R7859 gnd.n6263 gnd.n2839 71.676
R7860 gnd.n6260 gnd.n2840 71.676
R7861 gnd.n6256 gnd.n2841 71.676
R7862 gnd.n6252 gnd.n2842 71.676
R7863 gnd.n6248 gnd.n2843 71.676
R7864 gnd.n6244 gnd.n2844 71.676
R7865 gnd.n6240 gnd.n2845 71.676
R7866 gnd.n6236 gnd.n2846 71.676
R7867 gnd.n6232 gnd.n2847 71.676
R7868 gnd.n6228 gnd.n2848 71.676
R7869 gnd.n6224 gnd.n2849 71.676
R7870 gnd.n6220 gnd.n2850 71.676
R7871 gnd.n6216 gnd.n2851 71.676
R7872 gnd.n6212 gnd.n2852 71.676
R7873 gnd.n6208 gnd.n2853 71.676
R7874 gnd.n2854 gnd.n2838 71.676
R7875 gnd.n3781 gnd.n2855 71.676
R7876 gnd.n3786 gnd.n2856 71.676
R7877 gnd.n3790 gnd.n2857 71.676
R7878 gnd.n3794 gnd.n2858 71.676
R7879 gnd.n3798 gnd.n2859 71.676
R7880 gnd.n3802 gnd.n2860 71.676
R7881 gnd.n3806 gnd.n2861 71.676
R7882 gnd.n3810 gnd.n2862 71.676
R7883 gnd.n3814 gnd.n2863 71.676
R7884 gnd.n3818 gnd.n2864 71.676
R7885 gnd.n3822 gnd.n2865 71.676
R7886 gnd.n3826 gnd.n2866 71.676
R7887 gnd.n3830 gnd.n2867 71.676
R7888 gnd.n3834 gnd.n2868 71.676
R7889 gnd.n3838 gnd.n2869 71.676
R7890 gnd.n6269 gnd.n2872 71.676
R7891 gnd.n6261 gnd.n2839 71.676
R7892 gnd.n6257 gnd.n2840 71.676
R7893 gnd.n6253 gnd.n2841 71.676
R7894 gnd.n6249 gnd.n2842 71.676
R7895 gnd.n6245 gnd.n2843 71.676
R7896 gnd.n6241 gnd.n2844 71.676
R7897 gnd.n6237 gnd.n2845 71.676
R7898 gnd.n6233 gnd.n2846 71.676
R7899 gnd.n6229 gnd.n2847 71.676
R7900 gnd.n6225 gnd.n2848 71.676
R7901 gnd.n6221 gnd.n2849 71.676
R7902 gnd.n6217 gnd.n2850 71.676
R7903 gnd.n6213 gnd.n2851 71.676
R7904 gnd.n6209 gnd.n2852 71.676
R7905 gnd.n6272 gnd.n6271 71.676
R7906 gnd.n3780 gnd.n2854 71.676
R7907 gnd.n3785 gnd.n2855 71.676
R7908 gnd.n3789 gnd.n2856 71.676
R7909 gnd.n3793 gnd.n2857 71.676
R7910 gnd.n3797 gnd.n2858 71.676
R7911 gnd.n3801 gnd.n2859 71.676
R7912 gnd.n3805 gnd.n2860 71.676
R7913 gnd.n3809 gnd.n2861 71.676
R7914 gnd.n3813 gnd.n2862 71.676
R7915 gnd.n3817 gnd.n2863 71.676
R7916 gnd.n3821 gnd.n2864 71.676
R7917 gnd.n3825 gnd.n2865 71.676
R7918 gnd.n3829 gnd.n2866 71.676
R7919 gnd.n3833 gnd.n2867 71.676
R7920 gnd.n3837 gnd.n2868 71.676
R7921 gnd.n3841 gnd.n2869 71.676
R7922 gnd.n5280 gnd.n3543 71.676
R7923 gnd.n5288 gnd.n5287 71.676
R7924 gnd.n3542 gnd.n3540 71.676
R7925 gnd.n5295 gnd.n5294 71.676
R7926 gnd.n3539 gnd.n3537 71.676
R7927 gnd.n5302 gnd.n5301 71.676
R7928 gnd.n3536 gnd.n3534 71.676
R7929 gnd.n5309 gnd.n5308 71.676
R7930 gnd.n3533 gnd.n3531 71.676
R7931 gnd.n5316 gnd.n5315 71.676
R7932 gnd.n3530 gnd.n3528 71.676
R7933 gnd.n5323 gnd.n5322 71.676
R7934 gnd.n3527 gnd.n3525 71.676
R7935 gnd.n5330 gnd.n5329 71.676
R7936 gnd.n3524 gnd.n3520 71.676
R7937 gnd.n5338 gnd.n5337 71.676
R7938 gnd.n5342 gnd.n5341 71.676
R7939 gnd.n5346 gnd.n5345 71.676
R7940 gnd.n3518 gnd.n3514 71.676
R7941 gnd.n5354 gnd.n5353 71.676
R7942 gnd.n3513 gnd.n3511 71.676
R7943 gnd.n5361 gnd.n5360 71.676
R7944 gnd.n3510 gnd.n3508 71.676
R7945 gnd.n5368 gnd.n5367 71.676
R7946 gnd.n3507 gnd.n3505 71.676
R7947 gnd.n5375 gnd.n5374 71.676
R7948 gnd.n3504 gnd.n3502 71.676
R7949 gnd.n5382 gnd.n5381 71.676
R7950 gnd.n3501 gnd.n3499 71.676
R7951 gnd.n5389 gnd.n5388 71.676
R7952 gnd.n3498 gnd.n3496 71.676
R7953 gnd.n5396 gnd.n5395 71.676
R7954 gnd.n5399 gnd.n5398 71.676
R7955 gnd.n8 gnd.t397 69.1507
R7956 gnd.n14 gnd.t288 68.4792
R7957 gnd.n13 gnd.t375 68.4792
R7958 gnd.n12 gnd.t147 68.4792
R7959 gnd.n11 gnd.t114 68.4792
R7960 gnd.n10 gnd.t336 68.4792
R7961 gnd.n9 gnd.t89 68.4792
R7962 gnd.n8 gnd.t23 68.4792
R7963 gnd.n1623 gnd.n1527 64.369
R7964 gnd.n3783 gnd.n3778 59.5399
R7965 gnd.n5333 gnd.n3522 59.5399
R7966 gnd.n6207 gnd.n6206 59.5399
R7967 gnd.n5349 gnd.n3516 59.5399
R7968 gnd.n6204 gnd.n2893 59.1804
R7969 gnd.n6672 gnd.n1004 57.3586
R7970 gnd.n1314 gnd.t293 56.407
R7971 gnd.n1255 gnd.t318 56.407
R7972 gnd.n1274 gnd.t39 56.407
R7973 gnd.n1294 gnd.t46 56.407
R7974 gnd.n76 gnd.t364 56.407
R7975 gnd.n17 gnd.t71 56.407
R7976 gnd.n36 gnd.t394 56.407
R7977 gnd.n56 gnd.t53 56.407
R7978 gnd.n1331 gnd.t398 55.8337
R7979 gnd.n1272 gnd.t358 55.8337
R7980 gnd.n1291 gnd.t45 55.8337
R7981 gnd.n1311 gnd.t133 55.8337
R7982 gnd.n93 gnd.t292 55.8337
R7983 gnd.n34 gnd.t331 55.8337
R7984 gnd.n53 gnd.t57 55.8337
R7985 gnd.n73 gnd.t297 55.8337
R7986 gnd.n2881 gnd.n2880 54.358
R7987 gnd.n3487 gnd.n3486 54.358
R7988 gnd.n1314 gnd.n1313 53.0052
R7989 gnd.n1316 gnd.n1315 53.0052
R7990 gnd.n1318 gnd.n1317 53.0052
R7991 gnd.n1320 gnd.n1319 53.0052
R7992 gnd.n1322 gnd.n1321 53.0052
R7993 gnd.n1324 gnd.n1323 53.0052
R7994 gnd.n1326 gnd.n1325 53.0052
R7995 gnd.n1328 gnd.n1327 53.0052
R7996 gnd.n1330 gnd.n1329 53.0052
R7997 gnd.n1255 gnd.n1254 53.0052
R7998 gnd.n1257 gnd.n1256 53.0052
R7999 gnd.n1259 gnd.n1258 53.0052
R8000 gnd.n1261 gnd.n1260 53.0052
R8001 gnd.n1263 gnd.n1262 53.0052
R8002 gnd.n1265 gnd.n1264 53.0052
R8003 gnd.n1267 gnd.n1266 53.0052
R8004 gnd.n1269 gnd.n1268 53.0052
R8005 gnd.n1271 gnd.n1270 53.0052
R8006 gnd.n1274 gnd.n1273 53.0052
R8007 gnd.n1276 gnd.n1275 53.0052
R8008 gnd.n1278 gnd.n1277 53.0052
R8009 gnd.n1280 gnd.n1279 53.0052
R8010 gnd.n1282 gnd.n1281 53.0052
R8011 gnd.n1284 gnd.n1283 53.0052
R8012 gnd.n1286 gnd.n1285 53.0052
R8013 gnd.n1288 gnd.n1287 53.0052
R8014 gnd.n1290 gnd.n1289 53.0052
R8015 gnd.n1294 gnd.n1293 53.0052
R8016 gnd.n1296 gnd.n1295 53.0052
R8017 gnd.n1298 gnd.n1297 53.0052
R8018 gnd.n1300 gnd.n1299 53.0052
R8019 gnd.n1302 gnd.n1301 53.0052
R8020 gnd.n1304 gnd.n1303 53.0052
R8021 gnd.n1306 gnd.n1305 53.0052
R8022 gnd.n1308 gnd.n1307 53.0052
R8023 gnd.n1310 gnd.n1309 53.0052
R8024 gnd.n92 gnd.n91 53.0052
R8025 gnd.n90 gnd.n89 53.0052
R8026 gnd.n88 gnd.n87 53.0052
R8027 gnd.n86 gnd.n85 53.0052
R8028 gnd.n84 gnd.n83 53.0052
R8029 gnd.n82 gnd.n81 53.0052
R8030 gnd.n80 gnd.n79 53.0052
R8031 gnd.n78 gnd.n77 53.0052
R8032 gnd.n76 gnd.n75 53.0052
R8033 gnd.n33 gnd.n32 53.0052
R8034 gnd.n31 gnd.n30 53.0052
R8035 gnd.n29 gnd.n28 53.0052
R8036 gnd.n27 gnd.n26 53.0052
R8037 gnd.n25 gnd.n24 53.0052
R8038 gnd.n23 gnd.n22 53.0052
R8039 gnd.n21 gnd.n20 53.0052
R8040 gnd.n19 gnd.n18 53.0052
R8041 gnd.n17 gnd.n16 53.0052
R8042 gnd.n52 gnd.n51 53.0052
R8043 gnd.n50 gnd.n49 53.0052
R8044 gnd.n48 gnd.n47 53.0052
R8045 gnd.n46 gnd.n45 53.0052
R8046 gnd.n44 gnd.n43 53.0052
R8047 gnd.n42 gnd.n41 53.0052
R8048 gnd.n40 gnd.n39 53.0052
R8049 gnd.n38 gnd.n37 53.0052
R8050 gnd.n36 gnd.n35 53.0052
R8051 gnd.n72 gnd.n71 53.0052
R8052 gnd.n70 gnd.n69 53.0052
R8053 gnd.n68 gnd.n67 53.0052
R8054 gnd.n66 gnd.n65 53.0052
R8055 gnd.n64 gnd.n63 53.0052
R8056 gnd.n62 gnd.n61 53.0052
R8057 gnd.n60 gnd.n59 53.0052
R8058 gnd.n58 gnd.n57 53.0052
R8059 gnd.n56 gnd.n55 53.0052
R8060 gnd.n3478 gnd.n3477 52.4801
R8061 gnd.n2308 gnd.t141 52.3082
R8062 gnd.n2276 gnd.t349 52.3082
R8063 gnd.n2244 gnd.t13 52.3082
R8064 gnd.n2213 gnd.t150 52.3082
R8065 gnd.n2181 gnd.t390 52.3082
R8066 gnd.n2149 gnd.t327 52.3082
R8067 gnd.n2117 gnd.t392 52.3082
R8068 gnd.n2086 gnd.t368 52.3082
R8069 gnd.n6625 gnd.n2394 51.6227
R8070 gnd.n2138 gnd.n2106 51.4173
R8071 gnd.n2202 gnd.n2201 50.455
R8072 gnd.n2170 gnd.n2169 50.455
R8073 gnd.n2138 gnd.n2137 50.455
R8074 gnd.n1570 gnd.n1569 45.1884
R8075 gnd.n1034 gnd.n1033 45.1884
R8076 gnd.n5401 gnd.n3493 44.3322
R8077 gnd.n2884 gnd.n2883 44.3189
R8078 gnd.n4598 gnd.n4597 42.2793
R8079 gnd.n6032 gnd.n6031 42.2793
R8080 gnd.n1571 gnd.n1570 42.2793
R8081 gnd.n1035 gnd.n1034 42.2793
R8082 gnd.n1497 gnd.n1496 42.2793
R8083 gnd.n1014 gnd.n1013 42.2793
R8084 gnd.n4594 gnd.n4592 42.2793
R8085 gnd.n5991 gnd.n3128 42.2793
R8086 gnd.n5954 gnd.n3151 42.2793
R8087 gnd.n5914 gnd.n5911 42.2793
R8088 gnd.n7736 gnd.n353 42.2793
R8089 gnd.n7778 gnd.n333 42.2793
R8090 gnd.n7820 gnd.n7819 42.2793
R8091 gnd.n7620 gnd.n7619 42.2793
R8092 gnd.n6589 gnd.n2417 42.2793
R8093 gnd.n6549 gnd.n2439 42.2793
R8094 gnd.n6509 gnd.n2461 42.2793
R8095 gnd.n4132 gnd.n4080 42.2793
R8096 gnd.n6291 gnd.n2823 42.2793
R8097 gnd.n4750 gnd.n4660 42.2793
R8098 gnd.n4701 gnd.n4673 42.2793
R8099 gnd.n3057 gnd.n3056 42.2793
R8100 gnd.n2882 gnd.n2881 41.6274
R8101 gnd.n3488 gnd.n3487 41.6274
R8102 gnd.n2891 gnd.n2890 40.8975
R8103 gnd.n3491 gnd.n3490 40.8975
R8104 gnd.n6885 gnd.n786 38.268
R8105 gnd.n6879 gnd.n786 38.268
R8106 gnd.n6879 gnd.n6878 38.268
R8107 gnd.n6878 gnd.n6877 38.268
R8108 gnd.n6877 gnd.n793 38.268
R8109 gnd.n6871 gnd.n793 38.268
R8110 gnd.n6871 gnd.n6870 38.268
R8111 gnd.n6870 gnd.n6869 38.268
R8112 gnd.n6869 gnd.n801 38.268
R8113 gnd.n6863 gnd.n801 38.268
R8114 gnd.n6863 gnd.n6862 38.268
R8115 gnd.n6862 gnd.n6861 38.268
R8116 gnd.n6861 gnd.n809 38.268
R8117 gnd.n6855 gnd.n809 38.268
R8118 gnd.n6855 gnd.n6854 38.268
R8119 gnd.n6854 gnd.n6853 38.268
R8120 gnd.n6853 gnd.n817 38.268
R8121 gnd.n6847 gnd.n817 38.268
R8122 gnd.n6847 gnd.n6846 38.268
R8123 gnd.n6846 gnd.n6845 38.268
R8124 gnd.n6845 gnd.n825 38.268
R8125 gnd.n6839 gnd.n825 38.268
R8126 gnd.n6839 gnd.n6838 38.268
R8127 gnd.n6838 gnd.n6837 38.268
R8128 gnd.n6837 gnd.n833 38.268
R8129 gnd.n6831 gnd.n833 38.268
R8130 gnd.n6831 gnd.n6830 38.268
R8131 gnd.n6830 gnd.n6829 38.268
R8132 gnd.n6829 gnd.n841 38.268
R8133 gnd.n6823 gnd.n841 38.268
R8134 gnd.n6823 gnd.n6822 38.268
R8135 gnd.n6822 gnd.n6821 38.268
R8136 gnd.n6821 gnd.n849 38.268
R8137 gnd.n6815 gnd.n849 38.268
R8138 gnd.n6815 gnd.n6814 38.268
R8139 gnd.n6814 gnd.n6813 38.268
R8140 gnd.n6813 gnd.n857 38.268
R8141 gnd.n6807 gnd.n857 38.268
R8142 gnd.n6807 gnd.n6806 38.268
R8143 gnd.n6806 gnd.n6805 38.268
R8144 gnd.n6805 gnd.n865 38.268
R8145 gnd.n6799 gnd.n865 38.268
R8146 gnd.n6799 gnd.n6798 38.268
R8147 gnd.n6798 gnd.n6797 38.268
R8148 gnd.n6797 gnd.n873 38.268
R8149 gnd.n6791 gnd.n873 38.268
R8150 gnd.n6791 gnd.n6790 38.268
R8151 gnd.n6790 gnd.n6789 38.268
R8152 gnd.n6789 gnd.n881 38.268
R8153 gnd.n6783 gnd.n881 38.268
R8154 gnd.n6783 gnd.n6782 38.268
R8155 gnd.n6782 gnd.n6781 38.268
R8156 gnd.n6781 gnd.n889 38.268
R8157 gnd.n6775 gnd.n889 38.268
R8158 gnd.n6775 gnd.n6774 38.268
R8159 gnd.n6774 gnd.n6773 38.268
R8160 gnd.n6773 gnd.n897 38.268
R8161 gnd.n6767 gnd.n897 38.268
R8162 gnd.n6767 gnd.n6766 38.268
R8163 gnd.n6766 gnd.n6765 38.268
R8164 gnd.n6765 gnd.n905 38.268
R8165 gnd.n6759 gnd.n905 38.268
R8166 gnd.n6759 gnd.n6758 38.268
R8167 gnd.n6758 gnd.n6757 38.268
R8168 gnd.n6757 gnd.n913 38.268
R8169 gnd.n6751 gnd.n913 38.268
R8170 gnd.n6751 gnd.n6750 38.268
R8171 gnd.n6750 gnd.n6749 38.268
R8172 gnd.n6749 gnd.n921 38.268
R8173 gnd.n6743 gnd.n921 38.268
R8174 gnd.n6743 gnd.n6742 38.268
R8175 gnd.n6742 gnd.n6741 38.268
R8176 gnd.n6741 gnd.n929 38.268
R8177 gnd.n6735 gnd.n929 38.268
R8178 gnd.n6735 gnd.n6734 38.268
R8179 gnd.n6734 gnd.n6733 38.268
R8180 gnd.n6733 gnd.n937 38.268
R8181 gnd.n6727 gnd.n937 38.268
R8182 gnd.n6727 gnd.n6726 38.268
R8183 gnd.n6726 gnd.n6725 38.268
R8184 gnd.n6725 gnd.n945 38.268
R8185 gnd.n6719 gnd.n945 38.268
R8186 gnd.n6719 gnd.n6718 38.268
R8187 gnd.n7853 gnd.n256 35.69
R8188 gnd.n2890 gnd.n2889 35.055
R8189 gnd.n2885 gnd.n2884 35.055
R8190 gnd.n3480 gnd.n3479 35.055
R8191 gnd.n3490 gnd.n3476 35.055
R8192 gnd.n1633 gnd.n1527 31.8661
R8193 gnd.n1633 gnd.n1632 31.8661
R8194 gnd.n1641 gnd.n1516 31.8661
R8195 gnd.n1649 gnd.n1516 31.8661
R8196 gnd.n1649 gnd.n1510 31.8661
R8197 gnd.n1657 gnd.n1510 31.8661
R8198 gnd.n1657 gnd.n1503 31.8661
R8199 gnd.n1695 gnd.n1503 31.8661
R8200 gnd.n1705 gnd.n1436 31.8661
R8201 gnd.n6501 gnd.n2394 31.8661
R8202 gnd.n6495 gnd.n2478 31.8661
R8203 gnd.n6495 gnd.n2481 31.8661
R8204 gnd.n6489 gnd.n2481 31.8661
R8205 gnd.n6489 gnd.n2493 31.8661
R8206 gnd.n6483 gnd.n2503 31.8661
R8207 gnd.n6477 gnd.n2503 31.8661
R8208 gnd.n6471 gnd.n2519 31.8661
R8209 gnd.n6471 gnd.n2522 31.8661
R8210 gnd.n6465 gnd.n2532 31.8661
R8211 gnd.n4769 gnd.n2765 31.8661
R8212 gnd.n3912 gnd.n2776 31.8661
R8213 gnd.n4781 gnd.n3912 31.8661
R8214 gnd.n4781 gnd.n3927 31.8661
R8215 gnd.n3927 gnd.n3905 31.8661
R8216 gnd.n4789 gnd.n3905 31.8661
R8217 gnd.n4797 gnd.n3898 31.8661
R8218 gnd.n4797 gnd.n3890 31.8661
R8219 gnd.n4805 gnd.n3890 31.8661
R8220 gnd.n4805 gnd.n3892 31.8661
R8221 gnd.n4813 gnd.n3876 31.8661
R8222 gnd.n4821 gnd.n3876 31.8661
R8223 gnd.n4821 gnd.n3878 31.8661
R8224 gnd.n4829 gnd.n3861 31.8661
R8225 gnd.n4848 gnd.n3861 31.8661
R8226 gnd.n4848 gnd.n3853 31.8661
R8227 gnd.n4859 gnd.n3853 31.8661
R8228 gnd.n5422 gnd.n3454 31.8661
R8229 gnd.n5422 gnd.n3447 31.8661
R8230 gnd.n5430 gnd.n3447 31.8661
R8231 gnd.n5430 gnd.n3448 31.8661
R8232 gnd.n5438 gnd.n3434 31.8661
R8233 gnd.n5446 gnd.n3434 31.8661
R8234 gnd.n5446 gnd.n3435 31.8661
R8235 gnd.n5454 gnd.n3422 31.8661
R8236 gnd.n5465 gnd.n3422 31.8661
R8237 gnd.n5465 gnd.n3415 31.8661
R8238 gnd.n5473 gnd.n3415 31.8661
R8239 gnd.n6095 gnd.n2994 31.8661
R8240 gnd.n6095 gnd.n2996 31.8661
R8241 gnd.n5575 gnd.n2996 31.8661
R8242 gnd.n5575 gnd.n3408 31.8661
R8243 gnd.n3408 gnd.n3063 31.8661
R8244 gnd.n3173 gnd.n3105 31.8661
R8245 gnd.n7897 gnd.n188 31.8661
R8246 gnd.n7891 gnd.n199 31.8661
R8247 gnd.n7891 gnd.n202 31.8661
R8248 gnd.n7885 gnd.n211 31.8661
R8249 gnd.n7879 gnd.n211 31.8661
R8250 gnd.n7873 gnd.n227 31.8661
R8251 gnd.n7873 gnd.n230 31.8661
R8252 gnd.n7867 gnd.n230 31.8661
R8253 gnd.n7867 gnd.n240 31.8661
R8254 gnd.n7861 gnd.n249 31.8661
R8255 gnd.n3878 gnd.t396 30.9101
R8256 gnd.n5438 gnd.t332 30.9101
R8257 gnd.n5283 gnd.n5279 30.1273
R8258 gnd.n3844 gnd.n3840 30.1273
R8259 gnd.n6501 gnd.t179 28.3609
R8260 gnd.n7861 gnd.t183 28.3609
R8261 gnd.n6324 gnd.n2776 27.4049
R8262 gnd.n5414 gnd.n3460 27.4049
R8263 gnd.n6027 gnd.n3063 27.4049
R8264 gnd.n4597 gnd.n4596 25.7944
R8265 gnd.n6031 gnd.n6030 25.7944
R8266 gnd.n1496 gnd.n1495 25.7944
R8267 gnd.n1013 gnd.n1012 25.7944
R8268 gnd.n4592 gnd.n4591 25.7944
R8269 gnd.n3128 gnd.n3127 25.7944
R8270 gnd.n3151 gnd.n3150 25.7944
R8271 gnd.n5911 gnd.n5910 25.7944
R8272 gnd.n353 gnd.n352 25.7944
R8273 gnd.n333 gnd.n332 25.7944
R8274 gnd.n7819 gnd.n7818 25.7944
R8275 gnd.n7619 gnd.n7618 25.7944
R8276 gnd.n2417 gnd.n2416 25.7944
R8277 gnd.n2439 gnd.n2438 25.7944
R8278 gnd.n2461 gnd.n2460 25.7944
R8279 gnd.n4080 gnd.n4079 25.7944
R8280 gnd.n2823 gnd.n2822 25.7944
R8281 gnd.n4660 gnd.n4659 25.7944
R8282 gnd.n4673 gnd.n4672 25.7944
R8283 gnd.n3056 gnd.n3055 25.7944
R8284 gnd.n1717 gnd.n1437 24.8557
R8285 gnd.n1727 gnd.n1420 24.8557
R8286 gnd.n1423 gnd.n1411 24.8557
R8287 gnd.n1748 gnd.n1412 24.8557
R8288 gnd.n1758 gnd.n1392 24.8557
R8289 gnd.n1768 gnd.n1767 24.8557
R8290 gnd.n1376 gnd.n1375 24.8557
R8291 gnd.n1805 gnd.n1368 24.8557
R8292 gnd.n1804 gnd.n1361 24.8557
R8293 gnd.n1842 gnd.n1340 24.8557
R8294 gnd.n1816 gnd.n1341 24.8557
R8295 gnd.n1835 gnd.n1240 24.8557
R8296 gnd.n1852 gnd.n1851 24.8557
R8297 gnd.n1862 gnd.n1861 24.8557
R8298 gnd.n1231 gnd.n1223 24.8557
R8299 gnd.n1892 gnd.n1891 24.8557
R8300 gnd.n1902 gnd.n1201 24.8557
R8301 gnd.n1914 gnd.n1190 24.8557
R8302 gnd.n1905 gnd.n1183 24.8557
R8303 gnd.n1941 gnd.n1940 24.8557
R8304 gnd.n1951 gnd.n1176 24.8557
R8305 gnd.n1963 gnd.n1168 24.8557
R8306 gnd.n1981 gnd.n1980 24.8557
R8307 gnd.n1926 gnd.n1159 24.8557
R8308 gnd.n1991 gnd.n1149 24.8557
R8309 gnd.n2004 gnd.n1138 24.8557
R8310 gnd.n2042 gnd.n2041 24.8557
R8311 gnd.n2057 gnd.n1123 24.8557
R8312 gnd.n6710 gnd.n964 24.8557
R8313 gnd.n6709 gnd.n967 24.8557
R8314 gnd.n6703 gnd.n6702 24.8557
R8315 gnd.n2022 gnd.n979 24.8557
R8316 gnd.n6696 gnd.n988 24.8557
R8317 gnd.n6689 gnd.n6688 24.8557
R8318 gnd.n1738 gnd.t367 23.2624
R8319 gnd.t44 gnd.n2493 23.2624
R8320 gnd.n227 gnd.t56 23.2624
R8321 gnd.n6718 gnd.n6717 22.961
R8322 gnd.n1439 gnd.t221 22.6251
R8323 gnd.n2529 gnd.t18 22.3064
R8324 gnd.t204 gnd.n2870 22.3064
R8325 gnd.t54 gnd.n191 22.3064
R8326 gnd.n4893 gnd.n3765 21.6691
R8327 gnd.n4912 gnd.n3758 21.6691
R8328 gnd.n4880 gnd.n3744 21.6691
R8329 gnd.n4954 gnd.n3727 21.6691
R8330 gnd.n4976 gnd.n3701 21.6691
R8331 gnd.n4984 gnd.n3694 21.6691
R8332 gnd.n4991 gnd.n3687 21.6691
R8333 gnd.n5045 gnd.n3676 21.6691
R8334 gnd.n5033 gnd.n3667 21.6691
R8335 gnd.n5099 gnd.n3655 21.6691
R8336 gnd.n5117 gnd.n3637 21.6691
R8337 gnd.n5129 gnd.n3626 21.6691
R8338 gnd.n5145 gnd.n3616 21.6691
R8339 gnd.n5151 gnd.n3600 21.6691
R8340 gnd.n5220 gnd.n3584 21.6691
R8341 gnd.n5229 gnd.n3579 21.6691
R8342 gnd.n5252 gnd.n5251 21.6691
R8343 gnd.t149 gnd.n1444 21.3504
R8344 gnd.n5093 gnd.n3659 21.0318
R8345 gnd.n5100 gnd.n3652 21.0318
R8346 gnd.n5239 gnd.n3565 21.0318
R8347 gnd.t247 gnd.n3467 21.0318
R8348 gnd.n2035 gnd.t361 20.7131
R8349 gnd.n4813 gnd.t310 20.7131
R8350 gnd.n3435 gnd.t287 20.7131
R8351 gnd.t90 gnd.n1156 20.0758
R8352 gnd.n3778 gnd.n3777 19.9763
R8353 gnd.n3522 gnd.n3521 19.9763
R8354 gnd.n6206 gnd.n6205 19.9763
R8355 gnd.n3516 gnd.n3515 19.9763
R8356 gnd.n2879 gnd.t169 19.8005
R8357 gnd.n2879 gnd.t215 19.8005
R8358 gnd.n2878 gnd.t286 19.8005
R8359 gnd.n2878 gnd.t242 19.8005
R8360 gnd.n3485 gnd.t188 19.8005
R8361 gnd.n3485 gnd.t248 19.8005
R8362 gnd.n3484 gnd.t236 19.8005
R8363 gnd.n3484 gnd.t270 19.8005
R8364 gnd.n4900 gnd.n4899 19.7572
R8365 gnd.n5039 gnd.n3682 19.7572
R8366 gnd.n5111 gnd.n5110 19.7572
R8367 gnd.n5258 gnd.n3561 19.7572
R8368 gnd.n2875 gnd.n2874 19.5087
R8369 gnd.n2888 gnd.n2875 19.5087
R8370 gnd.n2886 gnd.n2877 19.5087
R8371 gnd.n3489 gnd.n3483 19.5087
R8372 gnd.t101 gnd.n1200 19.4385
R8373 gnd.n2519 gnd.t24 19.4385
R8374 gnd.t42 gnd.n202 19.4385
R8375 gnd.n4787 gnd.n3908 19.3944
R8376 gnd.n4787 gnd.n3896 19.3944
R8377 gnd.n4799 gnd.n3896 19.3944
R8378 gnd.n4799 gnd.n3894 19.3944
R8379 gnd.n4803 gnd.n3894 19.3944
R8380 gnd.n4803 gnd.n3882 19.3944
R8381 gnd.n4815 gnd.n3882 19.3944
R8382 gnd.n4815 gnd.n3880 19.3944
R8383 gnd.n4819 gnd.n3880 19.3944
R8384 gnd.n4819 gnd.n3868 19.3944
R8385 gnd.n4831 gnd.n3868 19.3944
R8386 gnd.n4831 gnd.n3865 19.3944
R8387 gnd.n4846 gnd.n3865 19.3944
R8388 gnd.n4846 gnd.n3866 19.3944
R8389 gnd.n4842 gnd.n3866 19.3944
R8390 gnd.n4842 gnd.n4841 19.3944
R8391 gnd.n4841 gnd.n4840 19.3944
R8392 gnd.n4840 gnd.n4837 19.3944
R8393 gnd.n4837 gnd.n2913 19.3944
R8394 gnd.n6191 gnd.n2913 19.3944
R8395 gnd.n6191 gnd.n2914 19.3944
R8396 gnd.n6187 gnd.n2914 19.3944
R8397 gnd.n6187 gnd.n6186 19.3944
R8398 gnd.n6186 gnd.n6185 19.3944
R8399 gnd.n6185 gnd.n2920 19.3944
R8400 gnd.n6181 gnd.n2920 19.3944
R8401 gnd.n6181 gnd.n6180 19.3944
R8402 gnd.n6180 gnd.n6179 19.3944
R8403 gnd.n6179 gnd.n2925 19.3944
R8404 gnd.n6175 gnd.n2925 19.3944
R8405 gnd.n6175 gnd.n6174 19.3944
R8406 gnd.n6174 gnd.n6173 19.3944
R8407 gnd.n6173 gnd.n2930 19.3944
R8408 gnd.n6169 gnd.n2930 19.3944
R8409 gnd.n6169 gnd.n6168 19.3944
R8410 gnd.n6168 gnd.n6167 19.3944
R8411 gnd.n6167 gnd.n2935 19.3944
R8412 gnd.n6163 gnd.n2935 19.3944
R8413 gnd.n6163 gnd.n6162 19.3944
R8414 gnd.n6162 gnd.n6161 19.3944
R8415 gnd.n6161 gnd.n2940 19.3944
R8416 gnd.n6157 gnd.n2940 19.3944
R8417 gnd.n6157 gnd.n6156 19.3944
R8418 gnd.n6156 gnd.n6155 19.3944
R8419 gnd.n6155 gnd.n2945 19.3944
R8420 gnd.n6151 gnd.n2945 19.3944
R8421 gnd.n6151 gnd.n6150 19.3944
R8422 gnd.n6150 gnd.n6149 19.3944
R8423 gnd.n6149 gnd.n2950 19.3944
R8424 gnd.n6145 gnd.n2950 19.3944
R8425 gnd.n6145 gnd.n6144 19.3944
R8426 gnd.n6144 gnd.n6143 19.3944
R8427 gnd.n6143 gnd.n2955 19.3944
R8428 gnd.n6139 gnd.n2955 19.3944
R8429 gnd.n6139 gnd.n6138 19.3944
R8430 gnd.n6138 gnd.n6137 19.3944
R8431 gnd.n6137 gnd.n2960 19.3944
R8432 gnd.n6133 gnd.n2960 19.3944
R8433 gnd.n6133 gnd.n6132 19.3944
R8434 gnd.n6132 gnd.n6131 19.3944
R8435 gnd.n6131 gnd.n2965 19.3944
R8436 gnd.n6127 gnd.n2965 19.3944
R8437 gnd.n6127 gnd.n6126 19.3944
R8438 gnd.n6126 gnd.n6125 19.3944
R8439 gnd.n6125 gnd.n2970 19.3944
R8440 gnd.n6121 gnd.n2970 19.3944
R8441 gnd.n6121 gnd.n6120 19.3944
R8442 gnd.n6120 gnd.n6119 19.3944
R8443 gnd.n6119 gnd.n2975 19.3944
R8444 gnd.n6115 gnd.n2975 19.3944
R8445 gnd.n6115 gnd.n6114 19.3944
R8446 gnd.n6114 gnd.n6113 19.3944
R8447 gnd.n6113 gnd.n2980 19.3944
R8448 gnd.n6109 gnd.n2980 19.3944
R8449 gnd.n6109 gnd.n6108 19.3944
R8450 gnd.n6108 gnd.n6107 19.3944
R8451 gnd.n6107 gnd.n2985 19.3944
R8452 gnd.n6103 gnd.n2985 19.3944
R8453 gnd.n6103 gnd.n6102 19.3944
R8454 gnd.n6102 gnd.n6101 19.3944
R8455 gnd.n6101 gnd.n2990 19.3944
R8456 gnd.n6097 gnd.n2990 19.3944
R8457 gnd.n4606 gnd.n4605 19.3944
R8458 gnd.n4605 gnd.n3910 19.3944
R8459 gnd.n4783 gnd.n3910 19.3944
R8460 gnd.n4524 gnd.n4523 19.3944
R8461 gnd.n4527 gnd.n4524 19.3944
R8462 gnd.n4527 gnd.n4479 19.3944
R8463 gnd.n4531 gnd.n4479 19.3944
R8464 gnd.n4532 gnd.n4531 19.3944
R8465 gnd.n4655 gnd.n4532 19.3944
R8466 gnd.n4655 gnd.n4654 19.3944
R8467 gnd.n4654 gnd.n4653 19.3944
R8468 gnd.n4653 gnd.n4537 19.3944
R8469 gnd.n4646 gnd.n4537 19.3944
R8470 gnd.n4646 gnd.n4645 19.3944
R8471 gnd.n4645 gnd.n4546 19.3944
R8472 gnd.n4638 gnd.n4546 19.3944
R8473 gnd.n4638 gnd.n4637 19.3944
R8474 gnd.n4637 gnd.n4556 19.3944
R8475 gnd.n4630 gnd.n4556 19.3944
R8476 gnd.n4630 gnd.n4629 19.3944
R8477 gnd.n4629 gnd.n4566 19.3944
R8478 gnd.n4622 gnd.n4566 19.3944
R8479 gnd.n4622 gnd.n4621 19.3944
R8480 gnd.n4621 gnd.n4576 19.3944
R8481 gnd.n4614 gnd.n4576 19.3944
R8482 gnd.n4614 gnd.n4613 19.3944
R8483 gnd.n4613 gnd.n4586 19.3944
R8484 gnd.n6073 gnd.n3016 19.3944
R8485 gnd.n6073 gnd.n6072 19.3944
R8486 gnd.n6072 gnd.n3019 19.3944
R8487 gnd.n6065 gnd.n3019 19.3944
R8488 gnd.n6065 gnd.n6064 19.3944
R8489 gnd.n6064 gnd.n3027 19.3944
R8490 gnd.n6057 gnd.n3027 19.3944
R8491 gnd.n6057 gnd.n6056 19.3944
R8492 gnd.n6056 gnd.n3035 19.3944
R8493 gnd.n6049 gnd.n3035 19.3944
R8494 gnd.n6049 gnd.n6048 19.3944
R8495 gnd.n6048 gnd.n3043 19.3944
R8496 gnd.n6041 gnd.n3043 19.3944
R8497 gnd.n6041 gnd.n6040 19.3944
R8498 gnd.n6040 gnd.n3051 19.3944
R8499 gnd.n6033 gnd.n3051 19.3944
R8500 gnd.n1620 gnd.n1619 19.3944
R8501 gnd.n1619 gnd.n1618 19.3944
R8502 gnd.n1618 gnd.n1617 19.3944
R8503 gnd.n1617 gnd.n1615 19.3944
R8504 gnd.n1615 gnd.n1612 19.3944
R8505 gnd.n1612 gnd.n1611 19.3944
R8506 gnd.n1611 gnd.n1608 19.3944
R8507 gnd.n1608 gnd.n1607 19.3944
R8508 gnd.n1607 gnd.n1604 19.3944
R8509 gnd.n1604 gnd.n1603 19.3944
R8510 gnd.n1603 gnd.n1600 19.3944
R8511 gnd.n1600 gnd.n1599 19.3944
R8512 gnd.n1599 gnd.n1596 19.3944
R8513 gnd.n1596 gnd.n1595 19.3944
R8514 gnd.n1595 gnd.n1592 19.3944
R8515 gnd.n1592 gnd.n1591 19.3944
R8516 gnd.n1591 gnd.n1588 19.3944
R8517 gnd.n1588 gnd.n1587 19.3944
R8518 gnd.n1587 gnd.n1584 19.3944
R8519 gnd.n1584 gnd.n1583 19.3944
R8520 gnd.n1583 gnd.n1580 19.3944
R8521 gnd.n1580 gnd.n1579 19.3944
R8522 gnd.n1576 gnd.n1575 19.3944
R8523 gnd.n1575 gnd.n1531 19.3944
R8524 gnd.n1626 gnd.n1531 19.3944
R8525 gnd.n1107 gnd.n1105 19.3944
R8526 gnd.n1107 gnd.n1031 19.3944
R8527 gnd.n2353 gnd.n1031 19.3944
R8528 gnd.n1048 gnd.n1047 19.3944
R8529 gnd.n1052 gnd.n1047 19.3944
R8530 gnd.n1055 gnd.n1052 19.3944
R8531 gnd.n1058 gnd.n1055 19.3944
R8532 gnd.n1058 gnd.n1044 19.3944
R8533 gnd.n1062 gnd.n1044 19.3944
R8534 gnd.n1065 gnd.n1062 19.3944
R8535 gnd.n1068 gnd.n1065 19.3944
R8536 gnd.n1068 gnd.n1042 19.3944
R8537 gnd.n1072 gnd.n1042 19.3944
R8538 gnd.n1075 gnd.n1072 19.3944
R8539 gnd.n1078 gnd.n1075 19.3944
R8540 gnd.n1078 gnd.n1040 19.3944
R8541 gnd.n1082 gnd.n1040 19.3944
R8542 gnd.n1085 gnd.n1082 19.3944
R8543 gnd.n1088 gnd.n1085 19.3944
R8544 gnd.n1088 gnd.n1038 19.3944
R8545 gnd.n1092 gnd.n1038 19.3944
R8546 gnd.n1095 gnd.n1092 19.3944
R8547 gnd.n1098 gnd.n1095 19.3944
R8548 gnd.n1098 gnd.n1036 19.3944
R8549 gnd.n1102 gnd.n1036 19.3944
R8550 gnd.n1719 gnd.n1428 19.3944
R8551 gnd.n1729 gnd.n1428 19.3944
R8552 gnd.n1730 gnd.n1729 19.3944
R8553 gnd.n1730 gnd.n1409 19.3944
R8554 gnd.n1750 gnd.n1409 19.3944
R8555 gnd.n1750 gnd.n1401 19.3944
R8556 gnd.n1760 gnd.n1401 19.3944
R8557 gnd.n1761 gnd.n1760 19.3944
R8558 gnd.n1762 gnd.n1761 19.3944
R8559 gnd.n1762 gnd.n1384 19.3944
R8560 gnd.n1384 gnd.n1382 19.3944
R8561 gnd.n1788 gnd.n1382 19.3944
R8562 gnd.n1788 gnd.n1364 19.3944
R8563 gnd.n1822 gnd.n1364 19.3944
R8564 gnd.n1822 gnd.n1821 19.3944
R8565 gnd.n1821 gnd.n1820 19.3944
R8566 gnd.n1820 gnd.n1815 19.3944
R8567 gnd.n1815 gnd.n1236 19.3944
R8568 gnd.n1854 gnd.n1236 19.3944
R8569 gnd.n1855 gnd.n1854 19.3944
R8570 gnd.n1856 gnd.n1855 19.3944
R8571 gnd.n1856 gnd.n1222 19.3944
R8572 gnd.n1222 gnd.n1216 19.3944
R8573 gnd.n1881 gnd.n1216 19.3944
R8574 gnd.n1882 gnd.n1881 19.3944
R8575 gnd.n1882 gnd.n1199 19.3944
R8576 gnd.n1199 gnd.n1197 19.3944
R8577 gnd.n1907 gnd.n1197 19.3944
R8578 gnd.n1908 gnd.n1907 19.3944
R8579 gnd.n1908 gnd.n1171 19.3944
R8580 gnd.n1958 gnd.n1171 19.3944
R8581 gnd.n1959 gnd.n1958 19.3944
R8582 gnd.n1959 gnd.n1164 19.3944
R8583 gnd.n1970 gnd.n1164 19.3944
R8584 gnd.n1971 gnd.n1970 19.3944
R8585 gnd.n1971 gnd.n1148 19.3944
R8586 gnd.n1148 gnd.n1146 19.3944
R8587 gnd.n1995 gnd.n1146 19.3944
R8588 gnd.n1998 gnd.n1995 19.3944
R8589 gnd.n1998 gnd.n1997 19.3944
R8590 gnd.n1997 gnd.n1119 19.3944
R8591 gnd.n2064 gnd.n1119 19.3944
R8592 gnd.n2064 gnd.n1116 19.3944
R8593 gnd.n2068 gnd.n1116 19.3944
R8594 gnd.n2069 gnd.n2068 19.3944
R8595 gnd.n2069 gnd.n1114 19.3944
R8596 gnd.n2075 gnd.n1114 19.3944
R8597 gnd.n2333 gnd.n2075 19.3944
R8598 gnd.n2337 gnd.n2333 19.3944
R8599 gnd.n2338 gnd.n2337 19.3944
R8600 gnd.n2343 gnd.n2338 19.3944
R8601 gnd.n2343 gnd.n1010 19.3944
R8602 gnd.n6683 gnd.n1010 19.3944
R8603 gnd.n1710 gnd.n1709 19.3944
R8604 gnd.n1709 gnd.n1442 19.3944
R8605 gnd.n1465 gnd.n1442 19.3944
R8606 gnd.n1468 gnd.n1465 19.3944
R8607 gnd.n1468 gnd.n1461 19.3944
R8608 gnd.n1472 gnd.n1461 19.3944
R8609 gnd.n1475 gnd.n1472 19.3944
R8610 gnd.n1478 gnd.n1475 19.3944
R8611 gnd.n1478 gnd.n1459 19.3944
R8612 gnd.n1482 gnd.n1459 19.3944
R8613 gnd.n1485 gnd.n1482 19.3944
R8614 gnd.n1488 gnd.n1485 19.3944
R8615 gnd.n1488 gnd.n1457 19.3944
R8616 gnd.n1492 gnd.n1457 19.3944
R8617 gnd.n1715 gnd.n1714 19.3944
R8618 gnd.n1714 gnd.n1418 19.3944
R8619 gnd.n1740 gnd.n1418 19.3944
R8620 gnd.n1740 gnd.n1416 19.3944
R8621 gnd.n1746 gnd.n1416 19.3944
R8622 gnd.n1746 gnd.n1745 19.3944
R8623 gnd.n1745 gnd.n1390 19.3944
R8624 gnd.n1770 gnd.n1390 19.3944
R8625 gnd.n1770 gnd.n1388 19.3944
R8626 gnd.n1782 gnd.n1388 19.3944
R8627 gnd.n1782 gnd.n1781 19.3944
R8628 gnd.n1781 gnd.n1780 19.3944
R8629 gnd.n1780 gnd.n1778 19.3944
R8630 gnd.n1778 gnd.n1360 19.3944
R8631 gnd.n1360 gnd.n1358 19.3944
R8632 gnd.n1829 gnd.n1358 19.3944
R8633 gnd.n1829 gnd.n1356 19.3944
R8634 gnd.n1833 gnd.n1356 19.3944
R8635 gnd.n1833 gnd.n1227 19.3944
R8636 gnd.n1864 gnd.n1227 19.3944
R8637 gnd.n1864 gnd.n1225 19.3944
R8638 gnd.n1868 gnd.n1225 19.3944
R8639 gnd.n1868 gnd.n1206 19.3944
R8640 gnd.n1894 gnd.n1206 19.3944
R8641 gnd.n1894 gnd.n1204 19.3944
R8642 gnd.n1900 gnd.n1204 19.3944
R8643 gnd.n1900 gnd.n1899 19.3944
R8644 gnd.n1899 gnd.n1181 19.3944
R8645 gnd.n1943 gnd.n1181 19.3944
R8646 gnd.n1943 gnd.n1179 19.3944
R8647 gnd.n1949 gnd.n1179 19.3944
R8648 gnd.n1949 gnd.n1948 19.3944
R8649 gnd.n1948 gnd.n1154 19.3944
R8650 gnd.n1983 gnd.n1154 19.3944
R8651 gnd.n1983 gnd.n1152 19.3944
R8652 gnd.n1989 gnd.n1152 19.3944
R8653 gnd.n1989 gnd.n1988 19.3944
R8654 gnd.n1988 gnd.n1129 19.3944
R8655 gnd.n2044 gnd.n1129 19.3944
R8656 gnd.n2044 gnd.n1127 19.3944
R8657 gnd.n2054 gnd.n1127 19.3944
R8658 gnd.n2054 gnd.n2053 19.3944
R8659 gnd.n2053 gnd.n2052 19.3944
R8660 gnd.n2052 gnd.n970 19.3944
R8661 gnd.n6707 gnd.n970 19.3944
R8662 gnd.n6707 gnd.n6706 19.3944
R8663 gnd.n6706 gnd.n6705 19.3944
R8664 gnd.n6705 gnd.n974 19.3944
R8665 gnd.n993 gnd.n974 19.3944
R8666 gnd.n6693 gnd.n993 19.3944
R8667 gnd.n6693 gnd.n6692 19.3944
R8668 gnd.n6692 gnd.n6691 19.3944
R8669 gnd.n6691 gnd.n999 19.3944
R8670 gnd.n6670 gnd.n6669 19.3944
R8671 gnd.n6669 gnd.n6635 19.3944
R8672 gnd.n6665 gnd.n6635 19.3944
R8673 gnd.n6665 gnd.n6662 19.3944
R8674 gnd.n6662 gnd.n6659 19.3944
R8675 gnd.n6659 gnd.n6658 19.3944
R8676 gnd.n6658 gnd.n6655 19.3944
R8677 gnd.n6655 gnd.n6654 19.3944
R8678 gnd.n6654 gnd.n6651 19.3944
R8679 gnd.n6651 gnd.n6650 19.3944
R8680 gnd.n6650 gnd.n6647 19.3944
R8681 gnd.n6647 gnd.n6646 19.3944
R8682 gnd.n6646 gnd.n1016 19.3944
R8683 gnd.n6676 gnd.n1016 19.3944
R8684 gnd.n1630 gnd.n1529 19.3944
R8685 gnd.n1630 gnd.n1520 19.3944
R8686 gnd.n1643 gnd.n1520 19.3944
R8687 gnd.n1643 gnd.n1518 19.3944
R8688 gnd.n1647 gnd.n1518 19.3944
R8689 gnd.n1647 gnd.n1508 19.3944
R8690 gnd.n1659 gnd.n1508 19.3944
R8691 gnd.n1659 gnd.n1506 19.3944
R8692 gnd.n1693 gnd.n1506 19.3944
R8693 gnd.n1693 gnd.n1692 19.3944
R8694 gnd.n1692 gnd.n1691 19.3944
R8695 gnd.n1691 gnd.n1690 19.3944
R8696 gnd.n1690 gnd.n1687 19.3944
R8697 gnd.n1687 gnd.n1686 19.3944
R8698 gnd.n1686 gnd.n1685 19.3944
R8699 gnd.n1685 gnd.n1683 19.3944
R8700 gnd.n1683 gnd.n1682 19.3944
R8701 gnd.n1682 gnd.n1679 19.3944
R8702 gnd.n1679 gnd.n1678 19.3944
R8703 gnd.n1678 gnd.n1677 19.3944
R8704 gnd.n1677 gnd.n1675 19.3944
R8705 gnd.n1675 gnd.n1373 19.3944
R8706 gnd.n1796 gnd.n1373 19.3944
R8707 gnd.n1796 gnd.n1371 19.3944
R8708 gnd.n1802 gnd.n1371 19.3944
R8709 gnd.n1802 gnd.n1801 19.3944
R8710 gnd.n1801 gnd.n1336 19.3944
R8711 gnd.n1844 gnd.n1336 19.3944
R8712 gnd.n1844 gnd.n1337 19.3944
R8713 gnd.n1353 gnd.n1352 19.3944
R8714 gnd.n1849 gnd.n1848 19.3944
R8715 gnd.n1252 gnd.n1244 19.3944
R8716 gnd.n1251 gnd.n1249 19.3944
R8717 gnd.n1249 gnd.n1248 19.3944
R8718 gnd.n1248 gnd.n1188 19.3944
R8719 gnd.n1916 gnd.n1188 19.3944
R8720 gnd.n1916 gnd.n1186 19.3944
R8721 gnd.n1936 gnd.n1186 19.3944
R8722 gnd.n1936 gnd.n1935 19.3944
R8723 gnd.n1935 gnd.n1934 19.3944
R8724 gnd.n1934 gnd.n1932 19.3944
R8725 gnd.n1932 gnd.n1931 19.3944
R8726 gnd.n1931 gnd.n1929 19.3944
R8727 gnd.n1929 gnd.n1928 19.3944
R8728 gnd.n1928 gnd.n1136 19.3944
R8729 gnd.n2006 gnd.n1136 19.3944
R8730 gnd.n2006 gnd.n1134 19.3944
R8731 gnd.n2039 gnd.n1134 19.3944
R8732 gnd.n2039 gnd.n2038 19.3944
R8733 gnd.n2038 gnd.n2037 19.3944
R8734 gnd.n2037 gnd.n2034 19.3944
R8735 gnd.n2034 gnd.n2033 19.3944
R8736 gnd.n2033 gnd.n2030 19.3944
R8737 gnd.n2030 gnd.n2029 19.3944
R8738 gnd.n2029 gnd.n2026 19.3944
R8739 gnd.n2026 gnd.n2025 19.3944
R8740 gnd.n2025 gnd.n2024 19.3944
R8741 gnd.n2024 gnd.n2021 19.3944
R8742 gnd.n2021 gnd.n1111 19.3944
R8743 gnd.n2349 gnd.n1111 19.3944
R8744 gnd.n2350 gnd.n2349 19.3944
R8745 gnd.n1635 gnd.n1525 19.3944
R8746 gnd.n1635 gnd.n1523 19.3944
R8747 gnd.n1639 gnd.n1523 19.3944
R8748 gnd.n1639 gnd.n1514 19.3944
R8749 gnd.n1651 gnd.n1514 19.3944
R8750 gnd.n1651 gnd.n1512 19.3944
R8751 gnd.n1655 gnd.n1512 19.3944
R8752 gnd.n1655 gnd.n1501 19.3944
R8753 gnd.n1697 gnd.n1501 19.3944
R8754 gnd.n1697 gnd.n1455 19.3944
R8755 gnd.n1703 gnd.n1455 19.3944
R8756 gnd.n1703 gnd.n1702 19.3944
R8757 gnd.n1702 gnd.n1433 19.3944
R8758 gnd.n1724 gnd.n1433 19.3944
R8759 gnd.n1724 gnd.n1426 19.3944
R8760 gnd.n1735 gnd.n1426 19.3944
R8761 gnd.n1735 gnd.n1734 19.3944
R8762 gnd.n1734 gnd.n1407 19.3944
R8763 gnd.n1755 gnd.n1407 19.3944
R8764 gnd.n1755 gnd.n1397 19.3944
R8765 gnd.n1765 gnd.n1397 19.3944
R8766 gnd.n1765 gnd.n1378 19.3944
R8767 gnd.n1792 gnd.n1378 19.3944
R8768 gnd.n1792 gnd.n1791 19.3944
R8769 gnd.n1791 gnd.n1366 19.3944
R8770 gnd.n1808 gnd.n1366 19.3944
R8771 gnd.n1808 gnd.n1344 19.3944
R8772 gnd.n1840 gnd.n1344 19.3944
R8773 gnd.n1840 gnd.n1839 19.3944
R8774 gnd.n1839 gnd.n1838 19.3944
R8775 gnd.n1838 gnd.n1350 19.3944
R8776 gnd.n1350 gnd.n1233 19.3944
R8777 gnd.n1859 gnd.n1233 19.3944
R8778 gnd.n1859 gnd.n1218 19.3944
R8779 gnd.n1876 gnd.n1218 19.3944
R8780 gnd.n1876 gnd.n1214 19.3944
R8781 gnd.n1889 gnd.n1214 19.3944
R8782 gnd.n1889 gnd.n1888 19.3944
R8783 gnd.n1888 gnd.n1193 19.3944
R8784 gnd.n1912 gnd.n1193 19.3944
R8785 gnd.n1912 gnd.n1911 19.3944
R8786 gnd.n1911 gnd.n1173 19.3944
R8787 gnd.n1954 gnd.n1173 19.3944
R8788 gnd.n1954 gnd.n1166 19.3944
R8789 gnd.n1965 gnd.n1166 19.3944
R8790 gnd.n1965 gnd.n1162 19.3944
R8791 gnd.n1978 gnd.n1162 19.3944
R8792 gnd.n1978 gnd.n1977 19.3944
R8793 gnd.n1977 gnd.n1142 19.3944
R8794 gnd.n2002 gnd.n1142 19.3944
R8795 gnd.n2002 gnd.n2001 19.3944
R8796 gnd.n2001 gnd.n1121 19.3944
R8797 gnd.n2059 gnd.n1121 19.3944
R8798 gnd.n2059 gnd.n958 19.3944
R8799 gnd.n6714 gnd.n958 19.3944
R8800 gnd.n6714 gnd.n6713 19.3944
R8801 gnd.n6713 gnd.n6712 19.3944
R8802 gnd.n6712 gnd.n962 19.3944
R8803 gnd.n982 gnd.n962 19.3944
R8804 gnd.n6700 gnd.n982 19.3944
R8805 gnd.n6700 gnd.n6699 19.3944
R8806 gnd.n6699 gnd.n6698 19.3944
R8807 gnd.n6698 gnd.n986 19.3944
R8808 gnd.n1007 gnd.n986 19.3944
R8809 gnd.n6686 gnd.n1007 19.3944
R8810 gnd.n4650 gnd.n4649 19.3944
R8811 gnd.n4649 gnd.n4540 19.3944
R8812 gnd.n4642 gnd.n4540 19.3944
R8813 gnd.n4642 gnd.n4641 19.3944
R8814 gnd.n4641 gnd.n4552 19.3944
R8815 gnd.n4634 gnd.n4552 19.3944
R8816 gnd.n4634 gnd.n4633 19.3944
R8817 gnd.n4633 gnd.n4560 19.3944
R8818 gnd.n4626 gnd.n4560 19.3944
R8819 gnd.n4626 gnd.n4625 19.3944
R8820 gnd.n4625 gnd.n4572 19.3944
R8821 gnd.n4618 gnd.n4572 19.3944
R8822 gnd.n4618 gnd.n4617 19.3944
R8823 gnd.n4617 gnd.n4580 19.3944
R8824 gnd.n4610 gnd.n4580 19.3944
R8825 gnd.n4610 gnd.n4609 19.3944
R8826 gnd.n7374 gnd.n491 19.3944
R8827 gnd.n7380 gnd.n491 19.3944
R8828 gnd.n7380 gnd.n489 19.3944
R8829 gnd.n7384 gnd.n489 19.3944
R8830 gnd.n7384 gnd.n485 19.3944
R8831 gnd.n7390 gnd.n485 19.3944
R8832 gnd.n7390 gnd.n483 19.3944
R8833 gnd.n7394 gnd.n483 19.3944
R8834 gnd.n7394 gnd.n479 19.3944
R8835 gnd.n7400 gnd.n479 19.3944
R8836 gnd.n7400 gnd.n477 19.3944
R8837 gnd.n7404 gnd.n477 19.3944
R8838 gnd.n7404 gnd.n473 19.3944
R8839 gnd.n7410 gnd.n473 19.3944
R8840 gnd.n7410 gnd.n471 19.3944
R8841 gnd.n7414 gnd.n471 19.3944
R8842 gnd.n7414 gnd.n467 19.3944
R8843 gnd.n7420 gnd.n467 19.3944
R8844 gnd.n7420 gnd.n465 19.3944
R8845 gnd.n7424 gnd.n465 19.3944
R8846 gnd.n7424 gnd.n461 19.3944
R8847 gnd.n7430 gnd.n461 19.3944
R8848 gnd.n7430 gnd.n459 19.3944
R8849 gnd.n7434 gnd.n459 19.3944
R8850 gnd.n7434 gnd.n455 19.3944
R8851 gnd.n7440 gnd.n455 19.3944
R8852 gnd.n7440 gnd.n453 19.3944
R8853 gnd.n7444 gnd.n453 19.3944
R8854 gnd.n7444 gnd.n449 19.3944
R8855 gnd.n7450 gnd.n449 19.3944
R8856 gnd.n7450 gnd.n447 19.3944
R8857 gnd.n7454 gnd.n447 19.3944
R8858 gnd.n7454 gnd.n443 19.3944
R8859 gnd.n7460 gnd.n443 19.3944
R8860 gnd.n7460 gnd.n441 19.3944
R8861 gnd.n7464 gnd.n441 19.3944
R8862 gnd.n7464 gnd.n437 19.3944
R8863 gnd.n7470 gnd.n437 19.3944
R8864 gnd.n7470 gnd.n435 19.3944
R8865 gnd.n7474 gnd.n435 19.3944
R8866 gnd.n7474 gnd.n431 19.3944
R8867 gnd.n7480 gnd.n431 19.3944
R8868 gnd.n7480 gnd.n429 19.3944
R8869 gnd.n7484 gnd.n429 19.3944
R8870 gnd.n7484 gnd.n425 19.3944
R8871 gnd.n7490 gnd.n425 19.3944
R8872 gnd.n7490 gnd.n423 19.3944
R8873 gnd.n7494 gnd.n423 19.3944
R8874 gnd.n7494 gnd.n419 19.3944
R8875 gnd.n7500 gnd.n419 19.3944
R8876 gnd.n7500 gnd.n417 19.3944
R8877 gnd.n7504 gnd.n417 19.3944
R8878 gnd.n7504 gnd.n413 19.3944
R8879 gnd.n7510 gnd.n413 19.3944
R8880 gnd.n7510 gnd.n411 19.3944
R8881 gnd.n7514 gnd.n411 19.3944
R8882 gnd.n7514 gnd.n407 19.3944
R8883 gnd.n7520 gnd.n407 19.3944
R8884 gnd.n7520 gnd.n405 19.3944
R8885 gnd.n7524 gnd.n405 19.3944
R8886 gnd.n7524 gnd.n401 19.3944
R8887 gnd.n7530 gnd.n401 19.3944
R8888 gnd.n7530 gnd.n399 19.3944
R8889 gnd.n7534 gnd.n399 19.3944
R8890 gnd.n7534 gnd.n395 19.3944
R8891 gnd.n7540 gnd.n395 19.3944
R8892 gnd.n7540 gnd.n393 19.3944
R8893 gnd.n7544 gnd.n393 19.3944
R8894 gnd.n7544 gnd.n389 19.3944
R8895 gnd.n7550 gnd.n389 19.3944
R8896 gnd.n7550 gnd.n387 19.3944
R8897 gnd.n7554 gnd.n387 19.3944
R8898 gnd.n7554 gnd.n383 19.3944
R8899 gnd.n7560 gnd.n383 19.3944
R8900 gnd.n7560 gnd.n381 19.3944
R8901 gnd.n7564 gnd.n381 19.3944
R8902 gnd.n7564 gnd.n377 19.3944
R8903 gnd.n7570 gnd.n377 19.3944
R8904 gnd.n7570 gnd.n375 19.3944
R8905 gnd.n7574 gnd.n375 19.3944
R8906 gnd.n7574 gnd.n371 19.3944
R8907 gnd.n7581 gnd.n371 19.3944
R8908 gnd.n7581 gnd.n369 19.3944
R8909 gnd.n7586 gnd.n369 19.3944
R8910 gnd.n6889 gnd.n784 19.3944
R8911 gnd.n6889 gnd.n782 19.3944
R8912 gnd.n6893 gnd.n782 19.3944
R8913 gnd.n6893 gnd.n778 19.3944
R8914 gnd.n6899 gnd.n778 19.3944
R8915 gnd.n6899 gnd.n776 19.3944
R8916 gnd.n6903 gnd.n776 19.3944
R8917 gnd.n6903 gnd.n772 19.3944
R8918 gnd.n6909 gnd.n772 19.3944
R8919 gnd.n6909 gnd.n770 19.3944
R8920 gnd.n6913 gnd.n770 19.3944
R8921 gnd.n6913 gnd.n766 19.3944
R8922 gnd.n6919 gnd.n766 19.3944
R8923 gnd.n6919 gnd.n764 19.3944
R8924 gnd.n6923 gnd.n764 19.3944
R8925 gnd.n6923 gnd.n760 19.3944
R8926 gnd.n6929 gnd.n760 19.3944
R8927 gnd.n6929 gnd.n758 19.3944
R8928 gnd.n6933 gnd.n758 19.3944
R8929 gnd.n6933 gnd.n754 19.3944
R8930 gnd.n6939 gnd.n754 19.3944
R8931 gnd.n6939 gnd.n752 19.3944
R8932 gnd.n6943 gnd.n752 19.3944
R8933 gnd.n6943 gnd.n748 19.3944
R8934 gnd.n6949 gnd.n748 19.3944
R8935 gnd.n6949 gnd.n746 19.3944
R8936 gnd.n6953 gnd.n746 19.3944
R8937 gnd.n6953 gnd.n742 19.3944
R8938 gnd.n6959 gnd.n742 19.3944
R8939 gnd.n6959 gnd.n740 19.3944
R8940 gnd.n6963 gnd.n740 19.3944
R8941 gnd.n6963 gnd.n736 19.3944
R8942 gnd.n6969 gnd.n736 19.3944
R8943 gnd.n6969 gnd.n734 19.3944
R8944 gnd.n6973 gnd.n734 19.3944
R8945 gnd.n6973 gnd.n730 19.3944
R8946 gnd.n6979 gnd.n730 19.3944
R8947 gnd.n6979 gnd.n728 19.3944
R8948 gnd.n6983 gnd.n728 19.3944
R8949 gnd.n6983 gnd.n724 19.3944
R8950 gnd.n6989 gnd.n724 19.3944
R8951 gnd.n6989 gnd.n722 19.3944
R8952 gnd.n6993 gnd.n722 19.3944
R8953 gnd.n6993 gnd.n718 19.3944
R8954 gnd.n6999 gnd.n718 19.3944
R8955 gnd.n6999 gnd.n716 19.3944
R8956 gnd.n7003 gnd.n716 19.3944
R8957 gnd.n7003 gnd.n712 19.3944
R8958 gnd.n7009 gnd.n712 19.3944
R8959 gnd.n7009 gnd.n710 19.3944
R8960 gnd.n7013 gnd.n710 19.3944
R8961 gnd.n7013 gnd.n706 19.3944
R8962 gnd.n7019 gnd.n706 19.3944
R8963 gnd.n7019 gnd.n704 19.3944
R8964 gnd.n7023 gnd.n704 19.3944
R8965 gnd.n7023 gnd.n700 19.3944
R8966 gnd.n7029 gnd.n700 19.3944
R8967 gnd.n7029 gnd.n698 19.3944
R8968 gnd.n7033 gnd.n698 19.3944
R8969 gnd.n7033 gnd.n694 19.3944
R8970 gnd.n7039 gnd.n694 19.3944
R8971 gnd.n7039 gnd.n692 19.3944
R8972 gnd.n7043 gnd.n692 19.3944
R8973 gnd.n7043 gnd.n688 19.3944
R8974 gnd.n7049 gnd.n688 19.3944
R8975 gnd.n7049 gnd.n686 19.3944
R8976 gnd.n7053 gnd.n686 19.3944
R8977 gnd.n7053 gnd.n682 19.3944
R8978 gnd.n7059 gnd.n682 19.3944
R8979 gnd.n7059 gnd.n680 19.3944
R8980 gnd.n7063 gnd.n680 19.3944
R8981 gnd.n7063 gnd.n676 19.3944
R8982 gnd.n7069 gnd.n676 19.3944
R8983 gnd.n7069 gnd.n674 19.3944
R8984 gnd.n7073 gnd.n674 19.3944
R8985 gnd.n7073 gnd.n670 19.3944
R8986 gnd.n7079 gnd.n670 19.3944
R8987 gnd.n7079 gnd.n668 19.3944
R8988 gnd.n7083 gnd.n668 19.3944
R8989 gnd.n7083 gnd.n664 19.3944
R8990 gnd.n7089 gnd.n664 19.3944
R8991 gnd.n7089 gnd.n662 19.3944
R8992 gnd.n7093 gnd.n662 19.3944
R8993 gnd.n7093 gnd.n658 19.3944
R8994 gnd.n7099 gnd.n658 19.3944
R8995 gnd.n7099 gnd.n656 19.3944
R8996 gnd.n7103 gnd.n656 19.3944
R8997 gnd.n7103 gnd.n652 19.3944
R8998 gnd.n7109 gnd.n652 19.3944
R8999 gnd.n7109 gnd.n650 19.3944
R9000 gnd.n7113 gnd.n650 19.3944
R9001 gnd.n7113 gnd.n646 19.3944
R9002 gnd.n7119 gnd.n646 19.3944
R9003 gnd.n7119 gnd.n644 19.3944
R9004 gnd.n7123 gnd.n644 19.3944
R9005 gnd.n7123 gnd.n640 19.3944
R9006 gnd.n7129 gnd.n640 19.3944
R9007 gnd.n7129 gnd.n638 19.3944
R9008 gnd.n7133 gnd.n638 19.3944
R9009 gnd.n7133 gnd.n634 19.3944
R9010 gnd.n7139 gnd.n634 19.3944
R9011 gnd.n7139 gnd.n632 19.3944
R9012 gnd.n7143 gnd.n632 19.3944
R9013 gnd.n7143 gnd.n628 19.3944
R9014 gnd.n7149 gnd.n628 19.3944
R9015 gnd.n7149 gnd.n626 19.3944
R9016 gnd.n7153 gnd.n626 19.3944
R9017 gnd.n7153 gnd.n622 19.3944
R9018 gnd.n7159 gnd.n622 19.3944
R9019 gnd.n7159 gnd.n620 19.3944
R9020 gnd.n7163 gnd.n620 19.3944
R9021 gnd.n7163 gnd.n616 19.3944
R9022 gnd.n7169 gnd.n616 19.3944
R9023 gnd.n7169 gnd.n614 19.3944
R9024 gnd.n7173 gnd.n614 19.3944
R9025 gnd.n7173 gnd.n610 19.3944
R9026 gnd.n7179 gnd.n610 19.3944
R9027 gnd.n7179 gnd.n608 19.3944
R9028 gnd.n7183 gnd.n608 19.3944
R9029 gnd.n7183 gnd.n604 19.3944
R9030 gnd.n7189 gnd.n604 19.3944
R9031 gnd.n7189 gnd.n602 19.3944
R9032 gnd.n7193 gnd.n602 19.3944
R9033 gnd.n7193 gnd.n598 19.3944
R9034 gnd.n7199 gnd.n598 19.3944
R9035 gnd.n7199 gnd.n596 19.3944
R9036 gnd.n7203 gnd.n596 19.3944
R9037 gnd.n7203 gnd.n592 19.3944
R9038 gnd.n7209 gnd.n592 19.3944
R9039 gnd.n7209 gnd.n590 19.3944
R9040 gnd.n7213 gnd.n590 19.3944
R9041 gnd.n7213 gnd.n586 19.3944
R9042 gnd.n7219 gnd.n586 19.3944
R9043 gnd.n7219 gnd.n584 19.3944
R9044 gnd.n7223 gnd.n584 19.3944
R9045 gnd.n7223 gnd.n580 19.3944
R9046 gnd.n7229 gnd.n580 19.3944
R9047 gnd.n7229 gnd.n578 19.3944
R9048 gnd.n7233 gnd.n578 19.3944
R9049 gnd.n7233 gnd.n574 19.3944
R9050 gnd.n7239 gnd.n574 19.3944
R9051 gnd.n7239 gnd.n572 19.3944
R9052 gnd.n7243 gnd.n572 19.3944
R9053 gnd.n7243 gnd.n568 19.3944
R9054 gnd.n7249 gnd.n568 19.3944
R9055 gnd.n7249 gnd.n566 19.3944
R9056 gnd.n7253 gnd.n566 19.3944
R9057 gnd.n7253 gnd.n562 19.3944
R9058 gnd.n7259 gnd.n562 19.3944
R9059 gnd.n7259 gnd.n560 19.3944
R9060 gnd.n7263 gnd.n560 19.3944
R9061 gnd.n7263 gnd.n556 19.3944
R9062 gnd.n7269 gnd.n556 19.3944
R9063 gnd.n7269 gnd.n554 19.3944
R9064 gnd.n7273 gnd.n554 19.3944
R9065 gnd.n7273 gnd.n550 19.3944
R9066 gnd.n7279 gnd.n550 19.3944
R9067 gnd.n7279 gnd.n548 19.3944
R9068 gnd.n7283 gnd.n548 19.3944
R9069 gnd.n7283 gnd.n544 19.3944
R9070 gnd.n7289 gnd.n544 19.3944
R9071 gnd.n7289 gnd.n542 19.3944
R9072 gnd.n7293 gnd.n542 19.3944
R9073 gnd.n7293 gnd.n538 19.3944
R9074 gnd.n7299 gnd.n538 19.3944
R9075 gnd.n7299 gnd.n536 19.3944
R9076 gnd.n7303 gnd.n536 19.3944
R9077 gnd.n7303 gnd.n532 19.3944
R9078 gnd.n7309 gnd.n532 19.3944
R9079 gnd.n7309 gnd.n530 19.3944
R9080 gnd.n7313 gnd.n530 19.3944
R9081 gnd.n7313 gnd.n526 19.3944
R9082 gnd.n7319 gnd.n526 19.3944
R9083 gnd.n7319 gnd.n524 19.3944
R9084 gnd.n7323 gnd.n524 19.3944
R9085 gnd.n7323 gnd.n520 19.3944
R9086 gnd.n7329 gnd.n520 19.3944
R9087 gnd.n7329 gnd.n518 19.3944
R9088 gnd.n7333 gnd.n518 19.3944
R9089 gnd.n7333 gnd.n514 19.3944
R9090 gnd.n7339 gnd.n514 19.3944
R9091 gnd.n7339 gnd.n512 19.3944
R9092 gnd.n7343 gnd.n512 19.3944
R9093 gnd.n7343 gnd.n508 19.3944
R9094 gnd.n7349 gnd.n508 19.3944
R9095 gnd.n7349 gnd.n506 19.3944
R9096 gnd.n7353 gnd.n506 19.3944
R9097 gnd.n7353 gnd.n502 19.3944
R9098 gnd.n7359 gnd.n502 19.3944
R9099 gnd.n7359 gnd.n500 19.3944
R9100 gnd.n7364 gnd.n500 19.3944
R9101 gnd.n7364 gnd.n496 19.3944
R9102 gnd.n7370 gnd.n496 19.3944
R9103 gnd.n7371 gnd.n7370 19.3944
R9104 gnd.n6024 gnd.n6023 19.3944
R9105 gnd.n6023 gnd.n6022 19.3944
R9106 gnd.n6022 gnd.n6021 19.3944
R9107 gnd.n6021 gnd.n6019 19.3944
R9108 gnd.n6019 gnd.n6016 19.3944
R9109 gnd.n6016 gnd.n6015 19.3944
R9110 gnd.n6015 gnd.n6012 19.3944
R9111 gnd.n6012 gnd.n6011 19.3944
R9112 gnd.n6011 gnd.n6008 19.3944
R9113 gnd.n6008 gnd.n6007 19.3944
R9114 gnd.n6007 gnd.n6004 19.3944
R9115 gnd.n6004 gnd.n6003 19.3944
R9116 gnd.n6003 gnd.n6000 19.3944
R9117 gnd.n6000 gnd.n5999 19.3944
R9118 gnd.n5999 gnd.n5996 19.3944
R9119 gnd.n5996 gnd.n5995 19.3944
R9120 gnd.n5995 gnd.n5992 19.3944
R9121 gnd.n5990 gnd.n5987 19.3944
R9122 gnd.n5987 gnd.n5986 19.3944
R9123 gnd.n5986 gnd.n5983 19.3944
R9124 gnd.n5983 gnd.n5982 19.3944
R9125 gnd.n5982 gnd.n5979 19.3944
R9126 gnd.n5979 gnd.n5978 19.3944
R9127 gnd.n5978 gnd.n5975 19.3944
R9128 gnd.n5973 gnd.n5970 19.3944
R9129 gnd.n5970 gnd.n5969 19.3944
R9130 gnd.n5969 gnd.n5966 19.3944
R9131 gnd.n5966 gnd.n5965 19.3944
R9132 gnd.n5965 gnd.n5962 19.3944
R9133 gnd.n5962 gnd.n5961 19.3944
R9134 gnd.n5961 gnd.n5958 19.3944
R9135 gnd.n5958 gnd.n5957 19.3944
R9136 gnd.n5953 gnd.n5950 19.3944
R9137 gnd.n5950 gnd.n5949 19.3944
R9138 gnd.n5949 gnd.n5946 19.3944
R9139 gnd.n5946 gnd.n5945 19.3944
R9140 gnd.n5945 gnd.n5942 19.3944
R9141 gnd.n5942 gnd.n5941 19.3944
R9142 gnd.n5941 gnd.n5938 19.3944
R9143 gnd.n5938 gnd.n5937 19.3944
R9144 gnd.n5937 gnd.n5934 19.3944
R9145 gnd.n5934 gnd.n5933 19.3944
R9146 gnd.n5933 gnd.n5930 19.3944
R9147 gnd.n5930 gnd.n5929 19.3944
R9148 gnd.n5929 gnd.n5926 19.3944
R9149 gnd.n5926 gnd.n5925 19.3944
R9150 gnd.n5925 gnd.n5922 19.3944
R9151 gnd.n5922 gnd.n5921 19.3944
R9152 gnd.n5921 gnd.n5918 19.3944
R9153 gnd.n5918 gnd.n5917 19.3944
R9154 gnd.n5901 gnd.n3172 19.3944
R9155 gnd.n5901 gnd.n5900 19.3944
R9156 gnd.n5900 gnd.n3181 19.3944
R9157 gnd.n3377 gnd.n3181 19.3944
R9158 gnd.n5596 gnd.n3377 19.3944
R9159 gnd.n5597 gnd.n5596 19.3944
R9160 gnd.n5599 gnd.n5597 19.3944
R9161 gnd.n5599 gnd.n3373 19.3944
R9162 gnd.n5611 gnd.n3373 19.3944
R9163 gnd.n5612 gnd.n5611 19.3944
R9164 gnd.n5614 gnd.n5612 19.3944
R9165 gnd.n5614 gnd.n3368 19.3944
R9166 gnd.n5626 gnd.n3368 19.3944
R9167 gnd.n5627 gnd.n5626 19.3944
R9168 gnd.n5629 gnd.n5627 19.3944
R9169 gnd.n5629 gnd.n3364 19.3944
R9170 gnd.n5641 gnd.n3364 19.3944
R9171 gnd.n5642 gnd.n5641 19.3944
R9172 gnd.n5644 gnd.n5642 19.3944
R9173 gnd.n5644 gnd.n3359 19.3944
R9174 gnd.n5656 gnd.n3359 19.3944
R9175 gnd.n5657 gnd.n5656 19.3944
R9176 gnd.n5659 gnd.n5657 19.3944
R9177 gnd.n5659 gnd.n3354 19.3944
R9178 gnd.n5683 gnd.n3354 19.3944
R9179 gnd.n5684 gnd.n5683 19.3944
R9180 gnd.n5685 gnd.n5684 19.3944
R9181 gnd.n5688 gnd.n5685 19.3944
R9182 gnd.n5688 gnd.n3352 19.3944
R9183 gnd.n5696 gnd.n3352 19.3944
R9184 gnd.n5697 gnd.n5696 19.3944
R9185 gnd.n5698 gnd.n5697 19.3944
R9186 gnd.n5799 gnd.n5698 19.3944
R9187 gnd.n5799 gnd.n5798 19.3944
R9188 gnd.n5798 gnd.n5797 19.3944
R9189 gnd.n5797 gnd.n5702 19.3944
R9190 gnd.n5731 gnd.n5702 19.3944
R9191 gnd.n5732 gnd.n5731 19.3944
R9192 gnd.n5733 gnd.n5732 19.3944
R9193 gnd.n5775 gnd.n5733 19.3944
R9194 gnd.n5775 gnd.n5774 19.3944
R9195 gnd.n5774 gnd.n5773 19.3944
R9196 gnd.n5773 gnd.n5735 19.3944
R9197 gnd.n5763 gnd.n5735 19.3944
R9198 gnd.n5763 gnd.n5762 19.3944
R9199 gnd.n5762 gnd.n5761 19.3944
R9200 gnd.n5761 gnd.n355 19.3944
R9201 gnd.n7703 gnd.n355 19.3944
R9202 gnd.n7704 gnd.n7703 19.3944
R9203 gnd.n7706 gnd.n7704 19.3944
R9204 gnd.n7707 gnd.n7706 19.3944
R9205 gnd.n7710 gnd.n7707 19.3944
R9206 gnd.n7711 gnd.n7710 19.3944
R9207 gnd.n7713 gnd.n7711 19.3944
R9208 gnd.n7714 gnd.n7713 19.3944
R9209 gnd.n7717 gnd.n7714 19.3944
R9210 gnd.n7718 gnd.n7717 19.3944
R9211 gnd.n7720 gnd.n7718 19.3944
R9212 gnd.n7721 gnd.n7720 19.3944
R9213 gnd.n7724 gnd.n7721 19.3944
R9214 gnd.n7725 gnd.n7724 19.3944
R9215 gnd.n7727 gnd.n7725 19.3944
R9216 gnd.n7728 gnd.n7727 19.3944
R9217 gnd.n7731 gnd.n7728 19.3944
R9218 gnd.n5904 gnd.n5903 19.3944
R9219 gnd.n5903 gnd.n3179 19.3944
R9220 gnd.n3203 gnd.n3179 19.3944
R9221 gnd.n5890 gnd.n3203 19.3944
R9222 gnd.n5890 gnd.n5889 19.3944
R9223 gnd.n5889 gnd.n5888 19.3944
R9224 gnd.n5888 gnd.n3208 19.3944
R9225 gnd.n5878 gnd.n3208 19.3944
R9226 gnd.n5878 gnd.n5877 19.3944
R9227 gnd.n5877 gnd.n5876 19.3944
R9228 gnd.n5876 gnd.n3229 19.3944
R9229 gnd.n5866 gnd.n3229 19.3944
R9230 gnd.n5866 gnd.n5865 19.3944
R9231 gnd.n5865 gnd.n5864 19.3944
R9232 gnd.n5864 gnd.n3249 19.3944
R9233 gnd.n5854 gnd.n3249 19.3944
R9234 gnd.n5854 gnd.n5853 19.3944
R9235 gnd.n5853 gnd.n5852 19.3944
R9236 gnd.n5852 gnd.n3270 19.3944
R9237 gnd.n5842 gnd.n3270 19.3944
R9238 gnd.n5842 gnd.n5841 19.3944
R9239 gnd.n5841 gnd.n5840 19.3944
R9240 gnd.n5840 gnd.n3290 19.3944
R9241 gnd.n5830 gnd.n3290 19.3944
R9242 gnd.n5830 gnd.n5829 19.3944
R9243 gnd.n5829 gnd.n5828 19.3944
R9244 gnd.n5828 gnd.n3312 19.3944
R9245 gnd.n5690 gnd.n3312 19.3944
R9246 gnd.n5693 gnd.n5690 19.3944
R9247 gnd.n5693 gnd.n3343 19.3944
R9248 gnd.n5805 gnd.n3343 19.3944
R9249 gnd.n5805 gnd.n5804 19.3944
R9250 gnd.n5804 gnd.n5803 19.3944
R9251 gnd.n5803 gnd.n3347 19.3944
R9252 gnd.n5793 gnd.n3347 19.3944
R9253 gnd.n5793 gnd.n124 19.3944
R9254 gnd.n7937 gnd.n124 19.3944
R9255 gnd.n7937 gnd.n7936 19.3944
R9256 gnd.n7936 gnd.n7935 19.3944
R9257 gnd.n7935 gnd.n128 19.3944
R9258 gnd.n7925 gnd.n128 19.3944
R9259 gnd.n7925 gnd.n7924 19.3944
R9260 gnd.n7924 gnd.n7923 19.3944
R9261 gnd.n7923 gnd.n146 19.3944
R9262 gnd.n7913 gnd.n146 19.3944
R9263 gnd.n7913 gnd.n7912 19.3944
R9264 gnd.n7912 gnd.n7911 19.3944
R9265 gnd.n7911 gnd.n167 19.3944
R9266 gnd.n7901 gnd.n167 19.3944
R9267 gnd.n7901 gnd.n7900 19.3944
R9268 gnd.n7900 gnd.n7899 19.3944
R9269 gnd.n7899 gnd.n186 19.3944
R9270 gnd.n7889 gnd.n186 19.3944
R9271 gnd.n7889 gnd.n7888 19.3944
R9272 gnd.n7888 gnd.n7887 19.3944
R9273 gnd.n7887 gnd.n207 19.3944
R9274 gnd.n7877 gnd.n207 19.3944
R9275 gnd.n7877 gnd.n7876 19.3944
R9276 gnd.n7876 gnd.n7875 19.3944
R9277 gnd.n7875 gnd.n225 19.3944
R9278 gnd.n7865 gnd.n225 19.3944
R9279 gnd.n7865 gnd.n7864 19.3944
R9280 gnd.n7864 gnd.n7863 19.3944
R9281 gnd.n7863 gnd.n245 19.3944
R9282 gnd.n7774 gnd.n331 19.3944
R9283 gnd.n7774 gnd.n7771 19.3944
R9284 gnd.n7771 gnd.n7768 19.3944
R9285 gnd.n7768 gnd.n7767 19.3944
R9286 gnd.n7767 gnd.n7764 19.3944
R9287 gnd.n7764 gnd.n7763 19.3944
R9288 gnd.n7763 gnd.n7760 19.3944
R9289 gnd.n7760 gnd.n7759 19.3944
R9290 gnd.n7759 gnd.n7756 19.3944
R9291 gnd.n7756 gnd.n7755 19.3944
R9292 gnd.n7755 gnd.n7752 19.3944
R9293 gnd.n7752 gnd.n7751 19.3944
R9294 gnd.n7751 gnd.n7748 19.3944
R9295 gnd.n7748 gnd.n7747 19.3944
R9296 gnd.n7747 gnd.n7744 19.3944
R9297 gnd.n7744 gnd.n7743 19.3944
R9298 gnd.n7743 gnd.n7740 19.3944
R9299 gnd.n7740 gnd.n7739 19.3944
R9300 gnd.n7817 gnd.n7814 19.3944
R9301 gnd.n7814 gnd.n7813 19.3944
R9302 gnd.n7813 gnd.n7810 19.3944
R9303 gnd.n7810 gnd.n7809 19.3944
R9304 gnd.n7809 gnd.n7806 19.3944
R9305 gnd.n7806 gnd.n7805 19.3944
R9306 gnd.n7805 gnd.n7802 19.3944
R9307 gnd.n7802 gnd.n7801 19.3944
R9308 gnd.n7801 gnd.n7798 19.3944
R9309 gnd.n7798 gnd.n7797 19.3944
R9310 gnd.n7797 gnd.n7794 19.3944
R9311 gnd.n7794 gnd.n7793 19.3944
R9312 gnd.n7793 gnd.n7790 19.3944
R9313 gnd.n7790 gnd.n7789 19.3944
R9314 gnd.n7789 gnd.n7786 19.3944
R9315 gnd.n7786 gnd.n7785 19.3944
R9316 gnd.n7785 gnd.n7782 19.3944
R9317 gnd.n7782 gnd.n7781 19.3944
R9318 gnd.n7855 gnd.n254 19.3944
R9319 gnd.n7850 gnd.n254 19.3944
R9320 gnd.n7850 gnd.n7849 19.3944
R9321 gnd.n7849 gnd.n7848 19.3944
R9322 gnd.n7848 gnd.n7845 19.3944
R9323 gnd.n7845 gnd.n7844 19.3944
R9324 gnd.n7844 gnd.n7841 19.3944
R9325 gnd.n7841 gnd.n7840 19.3944
R9326 gnd.n7840 gnd.n7837 19.3944
R9327 gnd.n7837 gnd.n7836 19.3944
R9328 gnd.n7836 gnd.n7833 19.3944
R9329 gnd.n7833 gnd.n7832 19.3944
R9330 gnd.n7832 gnd.n7829 19.3944
R9331 gnd.n7829 gnd.n7828 19.3944
R9332 gnd.n7828 gnd.n7825 19.3944
R9333 gnd.n7825 gnd.n7824 19.3944
R9334 gnd.n7824 gnd.n7821 19.3944
R9335 gnd.n7630 gnd.n7628 19.3944
R9336 gnd.n7633 gnd.n7630 19.3944
R9337 gnd.n7636 gnd.n7633 19.3944
R9338 gnd.n7639 gnd.n7636 19.3944
R9339 gnd.n7639 gnd.n7626 19.3944
R9340 gnd.n7643 gnd.n7626 19.3944
R9341 gnd.n7646 gnd.n7643 19.3944
R9342 gnd.n7649 gnd.n7646 19.3944
R9343 gnd.n7649 gnd.n7624 19.3944
R9344 gnd.n7653 gnd.n7624 19.3944
R9345 gnd.n7656 gnd.n7653 19.3944
R9346 gnd.n7659 gnd.n7656 19.3944
R9347 gnd.n7659 gnd.n7622 19.3944
R9348 gnd.n7663 gnd.n7622 19.3944
R9349 gnd.n7666 gnd.n7663 19.3944
R9350 gnd.n7669 gnd.n7666 19.3944
R9351 gnd.n5584 gnd.n3380 19.3944
R9352 gnd.n5585 gnd.n5584 19.3944
R9353 gnd.n5588 gnd.n5585 19.3944
R9354 gnd.n5588 gnd.n3378 19.3944
R9355 gnd.n5592 gnd.n3378 19.3944
R9356 gnd.n5592 gnd.n3376 19.3944
R9357 gnd.n5603 gnd.n3376 19.3944
R9358 gnd.n5603 gnd.n3374 19.3944
R9359 gnd.n5607 gnd.n3374 19.3944
R9360 gnd.n5607 gnd.n3372 19.3944
R9361 gnd.n5618 gnd.n3372 19.3944
R9362 gnd.n5618 gnd.n3370 19.3944
R9363 gnd.n5622 gnd.n3370 19.3944
R9364 gnd.n5622 gnd.n3367 19.3944
R9365 gnd.n5633 gnd.n3367 19.3944
R9366 gnd.n5633 gnd.n3365 19.3944
R9367 gnd.n5637 gnd.n3365 19.3944
R9368 gnd.n5637 gnd.n3363 19.3944
R9369 gnd.n5648 gnd.n3363 19.3944
R9370 gnd.n5648 gnd.n3361 19.3944
R9371 gnd.n5652 gnd.n3361 19.3944
R9372 gnd.n5652 gnd.n3358 19.3944
R9373 gnd.n5663 gnd.n3358 19.3944
R9374 gnd.n5663 gnd.n3355 19.3944
R9375 gnd.n5679 gnd.n3355 19.3944
R9376 gnd.n5679 gnd.n3356 19.3944
R9377 gnd.n5675 gnd.n3356 19.3944
R9378 gnd.n5675 gnd.n5674 19.3944
R9379 gnd.n5674 gnd.n5673 19.3944
R9380 gnd.n5673 gnd.n5670 19.3944
R9381 gnd.n5670 gnd.n5669 19.3944
R9382 gnd.n5669 gnd.n96 19.3944
R9383 gnd.n7950 gnd.n96 19.3944
R9384 gnd.n7950 gnd.n7949 19.3944
R9385 gnd.n7949 gnd.n99 19.3944
R9386 gnd.n5724 gnd.n99 19.3944
R9387 gnd.n5724 gnd.n5720 19.3944
R9388 gnd.n5781 gnd.n5720 19.3944
R9389 gnd.n5781 gnd.n5780 19.3944
R9390 gnd.n5780 gnd.n5779 19.3944
R9391 gnd.n5779 gnd.n5730 19.3944
R9392 gnd.n5769 gnd.n5730 19.3944
R9393 gnd.n5769 gnd.n5768 19.3944
R9394 gnd.n5768 gnd.n5767 19.3944
R9395 gnd.n5767 gnd.n359 19.3944
R9396 gnd.n7598 gnd.n359 19.3944
R9397 gnd.n7598 gnd.n357 19.3944
R9398 gnd.n7699 gnd.n357 19.3944
R9399 gnd.n7699 gnd.n7698 19.3944
R9400 gnd.n7698 gnd.n7697 19.3944
R9401 gnd.n7697 gnd.n7695 19.3944
R9402 gnd.n7695 gnd.n7694 19.3944
R9403 gnd.n7694 gnd.n7692 19.3944
R9404 gnd.n7692 gnd.n7691 19.3944
R9405 gnd.n7691 gnd.n7689 19.3944
R9406 gnd.n7689 gnd.n7688 19.3944
R9407 gnd.n7688 gnd.n7686 19.3944
R9408 gnd.n7686 gnd.n7685 19.3944
R9409 gnd.n7685 gnd.n7683 19.3944
R9410 gnd.n7683 gnd.n7682 19.3944
R9411 gnd.n7682 gnd.n7680 19.3944
R9412 gnd.n7680 gnd.n7679 19.3944
R9413 gnd.n7679 gnd.n7677 19.3944
R9414 gnd.n7677 gnd.n7676 19.3944
R9415 gnd.n3189 gnd.n3188 19.3944
R9416 gnd.n5896 gnd.n3188 19.3944
R9417 gnd.n5896 gnd.n5895 19.3944
R9418 gnd.n5895 gnd.n5894 19.3944
R9419 gnd.n5894 gnd.n3195 19.3944
R9420 gnd.n5884 gnd.n3195 19.3944
R9421 gnd.n5884 gnd.n5883 19.3944
R9422 gnd.n5883 gnd.n5882 19.3944
R9423 gnd.n5882 gnd.n3219 19.3944
R9424 gnd.n5872 gnd.n3219 19.3944
R9425 gnd.n5872 gnd.n5871 19.3944
R9426 gnd.n5871 gnd.n5870 19.3944
R9427 gnd.n5870 gnd.n3240 19.3944
R9428 gnd.n5860 gnd.n3240 19.3944
R9429 gnd.n5860 gnd.n5859 19.3944
R9430 gnd.n5859 gnd.n5858 19.3944
R9431 gnd.n5858 gnd.n3260 19.3944
R9432 gnd.n5848 gnd.n3260 19.3944
R9433 gnd.n5848 gnd.n5847 19.3944
R9434 gnd.n5847 gnd.n5846 19.3944
R9435 gnd.n5846 gnd.n3281 19.3944
R9436 gnd.n5836 gnd.n3281 19.3944
R9437 gnd.n5836 gnd.n5835 19.3944
R9438 gnd.n5835 gnd.n5834 19.3944
R9439 gnd.n5834 gnd.n3302 19.3944
R9440 gnd.n5824 gnd.n3302 19.3944
R9441 gnd.n5824 gnd.n5823 19.3944
R9442 gnd.n3334 gnd.n3333 19.3944
R9443 gnd.n5810 gnd.n5809 19.3944
R9444 gnd.n3337 gnd.n3336 19.3944
R9445 gnd.n7945 gnd.n7944 19.3944
R9446 gnd.n7941 gnd.n108 19.3944
R9447 gnd.n7941 gnd.n115 19.3944
R9448 gnd.n7931 gnd.n115 19.3944
R9449 gnd.n7931 gnd.n7930 19.3944
R9450 gnd.n7930 gnd.n7929 19.3944
R9451 gnd.n7929 gnd.n137 19.3944
R9452 gnd.n7919 gnd.n137 19.3944
R9453 gnd.n7919 gnd.n7918 19.3944
R9454 gnd.n7918 gnd.n7917 19.3944
R9455 gnd.n7917 gnd.n157 19.3944
R9456 gnd.n7907 gnd.n157 19.3944
R9457 gnd.n7907 gnd.n7906 19.3944
R9458 gnd.n7906 gnd.n7905 19.3944
R9459 gnd.n7905 gnd.n177 19.3944
R9460 gnd.n7895 gnd.n177 19.3944
R9461 gnd.n7895 gnd.n7894 19.3944
R9462 gnd.n7894 gnd.n7893 19.3944
R9463 gnd.n7893 gnd.n197 19.3944
R9464 gnd.n7883 gnd.n197 19.3944
R9465 gnd.n7883 gnd.n7882 19.3944
R9466 gnd.n7882 gnd.n7881 19.3944
R9467 gnd.n7881 gnd.n217 19.3944
R9468 gnd.n7871 gnd.n217 19.3944
R9469 gnd.n7871 gnd.n7870 19.3944
R9470 gnd.n7870 gnd.n7869 19.3944
R9471 gnd.n7869 gnd.n236 19.3944
R9472 gnd.n7859 gnd.n236 19.3944
R9473 gnd.n7859 gnd.n7858 19.3944
R9474 gnd.n4200 gnd.n4194 19.3944
R9475 gnd.n4205 gnd.n4194 19.3944
R9476 gnd.n4205 gnd.n4192 19.3944
R9477 gnd.n4209 gnd.n4192 19.3944
R9478 gnd.n4209 gnd.n4039 19.3944
R9479 gnd.n4213 gnd.n4039 19.3944
R9480 gnd.n4213 gnd.n4037 19.3944
R9481 gnd.n4217 gnd.n4037 19.3944
R9482 gnd.n4217 gnd.n4024 19.3944
R9483 gnd.n4257 gnd.n4024 19.3944
R9484 gnd.n4257 gnd.n4022 19.3944
R9485 gnd.n4261 gnd.n4022 19.3944
R9486 gnd.n4262 gnd.n4261 19.3944
R9487 gnd.n4266 gnd.n4265 19.3944
R9488 gnd.n4276 gnd.n4275 19.3944
R9489 gnd.n4273 gnd.n4270 19.3944
R9490 gnd.n4268 gnd.n3987 19.3944
R9491 gnd.n4322 gnd.n4321 19.3944
R9492 gnd.n4345 gnd.n4322 19.3944
R9493 gnd.n4345 gnd.n4344 19.3944
R9494 gnd.n4344 gnd.n4343 19.3944
R9495 gnd.n4343 gnd.n4327 19.3944
R9496 gnd.n4339 gnd.n4327 19.3944
R9497 gnd.n4339 gnd.n4338 19.3944
R9498 gnd.n4338 gnd.n4337 19.3944
R9499 gnd.n4337 gnd.n4335 19.3944
R9500 gnd.n4335 gnd.n3962 19.3944
R9501 gnd.n3962 gnd.n3960 19.3944
R9502 gnd.n4410 gnd.n3960 19.3944
R9503 gnd.n4410 gnd.n3958 19.3944
R9504 gnd.n4414 gnd.n3958 19.3944
R9505 gnd.n4414 gnd.n3956 19.3944
R9506 gnd.n4418 gnd.n3956 19.3944
R9507 gnd.n4418 gnd.n3954 19.3944
R9508 gnd.n4448 gnd.n3954 19.3944
R9509 gnd.n4448 gnd.n4447 19.3944
R9510 gnd.n4447 gnd.n4446 19.3944
R9511 gnd.n4446 gnd.n4424 19.3944
R9512 gnd.n4442 gnd.n4424 19.3944
R9513 gnd.n4442 gnd.n4441 19.3944
R9514 gnd.n4441 gnd.n4440 19.3944
R9515 gnd.n4440 gnd.n4430 19.3944
R9516 gnd.n4436 gnd.n4430 19.3944
R9517 gnd.n4436 gnd.n4435 19.3944
R9518 gnd.n4435 gnd.n3934 19.3944
R9519 gnd.n3934 gnd.n3932 19.3944
R9520 gnd.n4773 gnd.n3932 19.3944
R9521 gnd.n4773 gnd.n3930 19.3944
R9522 gnd.n4779 gnd.n3930 19.3944
R9523 gnd.n4779 gnd.n4778 19.3944
R9524 gnd.n4778 gnd.n3903 19.3944
R9525 gnd.n4791 gnd.n3903 19.3944
R9526 gnd.n4791 gnd.n3901 19.3944
R9527 gnd.n4795 gnd.n3901 19.3944
R9528 gnd.n4795 gnd.n3888 19.3944
R9529 gnd.n4807 gnd.n3888 19.3944
R9530 gnd.n4807 gnd.n3886 19.3944
R9531 gnd.n4811 gnd.n3886 19.3944
R9532 gnd.n4811 gnd.n3874 19.3944
R9533 gnd.n4823 gnd.n3874 19.3944
R9534 gnd.n4823 gnd.n3872 19.3944
R9535 gnd.n4827 gnd.n3872 19.3944
R9536 gnd.n4827 gnd.n3859 19.3944
R9537 gnd.n4850 gnd.n3859 19.3944
R9538 gnd.n4850 gnd.n3857 19.3944
R9539 gnd.n4857 gnd.n3857 19.3944
R9540 gnd.n4857 gnd.n4856 19.3944
R9541 gnd.n4856 gnd.n2903 19.3944
R9542 gnd.n6197 gnd.n2903 19.3944
R9543 gnd.n6197 gnd.n6196 19.3944
R9544 gnd.n6196 gnd.n6195 19.3944
R9545 gnd.n6195 gnd.n2907 19.3944
R9546 gnd.n3769 gnd.n2907 19.3944
R9547 gnd.n3769 gnd.n3749 19.3944
R9548 gnd.n4924 gnd.n3749 19.3944
R9549 gnd.n4924 gnd.n3747 19.3944
R9550 gnd.n4928 gnd.n3747 19.3944
R9551 gnd.n4928 gnd.n3725 19.3944
R9552 gnd.n4963 gnd.n3725 19.3944
R9553 gnd.n4963 gnd.n3723 19.3944
R9554 gnd.n4967 gnd.n3723 19.3944
R9555 gnd.n4967 gnd.n3699 19.3944
R9556 gnd.n5003 gnd.n3699 19.3944
R9557 gnd.n5003 gnd.n3697 19.3944
R9558 gnd.n5009 gnd.n3697 19.3944
R9559 gnd.n5009 gnd.n5008 19.3944
R9560 gnd.n5008 gnd.n3672 19.3944
R9561 gnd.n5049 gnd.n3672 19.3944
R9562 gnd.n5049 gnd.n3670 19.3944
R9563 gnd.n5055 gnd.n3670 19.3944
R9564 gnd.n5055 gnd.n5054 19.3944
R9565 gnd.n5054 gnd.n3650 19.3944
R9566 gnd.n5102 gnd.n3650 19.3944
R9567 gnd.n5102 gnd.n3648 19.3944
R9568 gnd.n5108 gnd.n3648 19.3944
R9569 gnd.n5108 gnd.n5107 19.3944
R9570 gnd.n5107 gnd.n3624 19.3944
R9571 gnd.n5138 gnd.n3624 19.3944
R9572 gnd.n5138 gnd.n3622 19.3944
R9573 gnd.n5142 gnd.n3622 19.3944
R9574 gnd.n5142 gnd.n3598 19.3944
R9575 gnd.n5180 gnd.n3598 19.3944
R9576 gnd.n5180 gnd.n3596 19.3944
R9577 gnd.n5186 gnd.n3596 19.3944
R9578 gnd.n5186 gnd.n5185 19.3944
R9579 gnd.n5185 gnd.n3574 19.3944
R9580 gnd.n5232 gnd.n3574 19.3944
R9581 gnd.n5232 gnd.n3572 19.3944
R9582 gnd.n5236 gnd.n3572 19.3944
R9583 gnd.n5236 gnd.n3556 19.3944
R9584 gnd.n5261 gnd.n3556 19.3944
R9585 gnd.n5261 gnd.n3554 19.3944
R9586 gnd.n5265 gnd.n3554 19.3944
R9587 gnd.n5265 gnd.n3465 19.3944
R9588 gnd.n5408 gnd.n3465 19.3944
R9589 gnd.n5408 gnd.n3463 19.3944
R9590 gnd.n5412 gnd.n3463 19.3944
R9591 gnd.n5412 gnd.n3452 19.3944
R9592 gnd.n5424 gnd.n3452 19.3944
R9593 gnd.n5424 gnd.n3450 19.3944
R9594 gnd.n5428 gnd.n3450 19.3944
R9595 gnd.n5428 gnd.n3439 19.3944
R9596 gnd.n5440 gnd.n3439 19.3944
R9597 gnd.n5440 gnd.n3437 19.3944
R9598 gnd.n5444 gnd.n3437 19.3944
R9599 gnd.n5444 gnd.n3426 19.3944
R9600 gnd.n5456 gnd.n3426 19.3944
R9601 gnd.n5456 gnd.n3424 19.3944
R9602 gnd.n5463 gnd.n3424 19.3944
R9603 gnd.n5463 gnd.n5462 19.3944
R9604 gnd.n5462 gnd.n3413 19.3944
R9605 gnd.n5476 gnd.n3413 19.3944
R9606 gnd.n5477 gnd.n5476 19.3944
R9607 gnd.n5477 gnd.n3411 19.3944
R9608 gnd.n5573 gnd.n3411 19.3944
R9609 gnd.n5573 gnd.n5572 19.3944
R9610 gnd.n5572 gnd.n5571 19.3944
R9611 gnd.n5571 gnd.n5483 19.3944
R9612 gnd.n5567 gnd.n5483 19.3944
R9613 gnd.n5567 gnd.n5566 19.3944
R9614 gnd.n5566 gnd.n5565 19.3944
R9615 gnd.n5565 gnd.n5489 19.3944
R9616 gnd.n5559 gnd.n5489 19.3944
R9617 gnd.n5559 gnd.n5558 19.3944
R9618 gnd.n5558 gnd.n5557 19.3944
R9619 gnd.n5557 gnd.n5495 19.3944
R9620 gnd.n5553 gnd.n5495 19.3944
R9621 gnd.n5553 gnd.n5552 19.3944
R9622 gnd.n5552 gnd.n5551 19.3944
R9623 gnd.n5551 gnd.n5501 19.3944
R9624 gnd.n5547 gnd.n5501 19.3944
R9625 gnd.n5547 gnd.n5546 19.3944
R9626 gnd.n5546 gnd.n5545 19.3944
R9627 gnd.n5545 gnd.n5507 19.3944
R9628 gnd.n5541 gnd.n5507 19.3944
R9629 gnd.n5541 gnd.n5540 19.3944
R9630 gnd.n5540 gnd.n5539 19.3944
R9631 gnd.n5539 gnd.n5513 19.3944
R9632 gnd.n5535 gnd.n5513 19.3944
R9633 gnd.n5535 gnd.n5534 19.3944
R9634 gnd.n5534 gnd.n5533 19.3944
R9635 gnd.n5533 gnd.n5519 19.3944
R9636 gnd.n5529 gnd.n5519 19.3944
R9637 gnd.n5529 gnd.n5528 19.3944
R9638 gnd.n5528 gnd.n5527 19.3944
R9639 gnd.n5527 gnd.n3324 19.3944
R9640 gnd.n5818 gnd.n3324 19.3944
R9641 gnd.n5816 gnd.n5815 19.3944
R9642 gnd.n5709 gnd.n5707 19.3944
R9643 gnd.n5713 gnd.n5706 19.3944
R9644 gnd.n5790 gnd.n5715 19.3944
R9645 gnd.n5788 gnd.n5787 19.3944
R9646 gnd.n5787 gnd.n5717 19.3944
R9647 gnd.n5740 gnd.n5717 19.3944
R9648 gnd.n5740 gnd.n5738 19.3944
R9649 gnd.n5753 gnd.n5738 19.3944
R9650 gnd.n5753 gnd.n5752 19.3944
R9651 gnd.n5752 gnd.n5751 19.3944
R9652 gnd.n5751 gnd.n5748 19.3944
R9653 gnd.n5748 gnd.n363 19.3944
R9654 gnd.n7593 gnd.n363 19.3944
R9655 gnd.n7593 gnd.n7592 19.3944
R9656 gnd.n7592 gnd.n7591 19.3944
R9657 gnd.n7591 gnd.n367 19.3944
R9658 gnd.n6622 gnd.n6621 19.3944
R9659 gnd.n6621 gnd.n6620 19.3944
R9660 gnd.n6620 gnd.n6619 19.3944
R9661 gnd.n6619 gnd.n6617 19.3944
R9662 gnd.n6617 gnd.n6614 19.3944
R9663 gnd.n6614 gnd.n6613 19.3944
R9664 gnd.n6613 gnd.n6610 19.3944
R9665 gnd.n6610 gnd.n6609 19.3944
R9666 gnd.n6609 gnd.n6606 19.3944
R9667 gnd.n6606 gnd.n6605 19.3944
R9668 gnd.n6605 gnd.n6602 19.3944
R9669 gnd.n6602 gnd.n6601 19.3944
R9670 gnd.n6601 gnd.n6598 19.3944
R9671 gnd.n6598 gnd.n6597 19.3944
R9672 gnd.n6597 gnd.n6594 19.3944
R9673 gnd.n6594 gnd.n6593 19.3944
R9674 gnd.n6593 gnd.n6590 19.3944
R9675 gnd.n6588 gnd.n6585 19.3944
R9676 gnd.n6585 gnd.n6584 19.3944
R9677 gnd.n6584 gnd.n6581 19.3944
R9678 gnd.n6581 gnd.n6580 19.3944
R9679 gnd.n6580 gnd.n6577 19.3944
R9680 gnd.n6577 gnd.n6576 19.3944
R9681 gnd.n6576 gnd.n6573 19.3944
R9682 gnd.n6573 gnd.n6572 19.3944
R9683 gnd.n6572 gnd.n6569 19.3944
R9684 gnd.n6569 gnd.n6568 19.3944
R9685 gnd.n6568 gnd.n6565 19.3944
R9686 gnd.n6565 gnd.n6564 19.3944
R9687 gnd.n6564 gnd.n6561 19.3944
R9688 gnd.n6561 gnd.n6560 19.3944
R9689 gnd.n6560 gnd.n6557 19.3944
R9690 gnd.n6557 gnd.n6556 19.3944
R9691 gnd.n6556 gnd.n6553 19.3944
R9692 gnd.n6553 gnd.n6552 19.3944
R9693 gnd.n6548 gnd.n6545 19.3944
R9694 gnd.n6545 gnd.n6544 19.3944
R9695 gnd.n6544 gnd.n6541 19.3944
R9696 gnd.n6541 gnd.n6540 19.3944
R9697 gnd.n6540 gnd.n6537 19.3944
R9698 gnd.n6537 gnd.n6536 19.3944
R9699 gnd.n6536 gnd.n6533 19.3944
R9700 gnd.n6533 gnd.n6532 19.3944
R9701 gnd.n6532 gnd.n6529 19.3944
R9702 gnd.n6529 gnd.n6528 19.3944
R9703 gnd.n6528 gnd.n6525 19.3944
R9704 gnd.n6525 gnd.n6524 19.3944
R9705 gnd.n6524 gnd.n6521 19.3944
R9706 gnd.n6521 gnd.n6520 19.3944
R9707 gnd.n6520 gnd.n6517 19.3944
R9708 gnd.n6517 gnd.n6516 19.3944
R9709 gnd.n6516 gnd.n6513 19.3944
R9710 gnd.n6513 gnd.n6512 19.3944
R9711 gnd.n4094 gnd.n4093 19.3944
R9712 gnd.n4097 gnd.n4094 19.3944
R9713 gnd.n4097 gnd.n4089 19.3944
R9714 gnd.n4103 gnd.n4089 19.3944
R9715 gnd.n4104 gnd.n4103 19.3944
R9716 gnd.n4107 gnd.n4104 19.3944
R9717 gnd.n4107 gnd.n4087 19.3944
R9718 gnd.n4113 gnd.n4087 19.3944
R9719 gnd.n4114 gnd.n4113 19.3944
R9720 gnd.n4117 gnd.n4114 19.3944
R9721 gnd.n4117 gnd.n4085 19.3944
R9722 gnd.n4123 gnd.n4085 19.3944
R9723 gnd.n4124 gnd.n4123 19.3944
R9724 gnd.n4127 gnd.n4124 19.3944
R9725 gnd.n4127 gnd.n4081 19.3944
R9726 gnd.n4131 gnd.n4081 19.3944
R9727 gnd.n4138 gnd.n4137 19.3944
R9728 gnd.n4140 gnd.n4138 19.3944
R9729 gnd.n4140 gnd.n4075 19.3944
R9730 gnd.n4145 gnd.n4075 19.3944
R9731 gnd.n4146 gnd.n4145 19.3944
R9732 gnd.n4148 gnd.n4146 19.3944
R9733 gnd.n4148 gnd.n4073 19.3944
R9734 gnd.n4153 gnd.n4073 19.3944
R9735 gnd.n4154 gnd.n4153 19.3944
R9736 gnd.n4156 gnd.n4154 19.3944
R9737 gnd.n4156 gnd.n4071 19.3944
R9738 gnd.n4161 gnd.n4071 19.3944
R9739 gnd.n4162 gnd.n4161 19.3944
R9740 gnd.n4164 gnd.n4162 19.3944
R9741 gnd.n4164 gnd.n4069 19.3944
R9742 gnd.n4169 gnd.n4069 19.3944
R9743 gnd.n4169 gnd.n4041 19.3944
R9744 gnd.n4187 gnd.n4041 19.3944
R9745 gnd.n4187 gnd.n4186 19.3944
R9746 gnd.n4186 gnd.n4185 19.3944
R9747 gnd.n4185 gnd.n4034 19.3944
R9748 gnd.n4222 gnd.n4034 19.3944
R9749 gnd.n4222 gnd.n4032 19.3944
R9750 gnd.n4227 gnd.n4032 19.3944
R9751 gnd.n4227 gnd.n4027 19.3944
R9752 gnd.n4251 gnd.n4027 19.3944
R9753 gnd.n4251 gnd.n4250 19.3944
R9754 gnd.n4250 gnd.n4249 19.3944
R9755 gnd.n4249 gnd.n4016 19.3944
R9756 gnd.n4281 gnd.n4016 19.3944
R9757 gnd.n4281 gnd.n4014 19.3944
R9758 gnd.n4285 gnd.n4014 19.3944
R9759 gnd.n4285 gnd.n3993 19.3944
R9760 gnd.n4311 gnd.n3993 19.3944
R9761 gnd.n4311 gnd.n3991 19.3944
R9762 gnd.n4315 gnd.n3991 19.3944
R9763 gnd.n4315 gnd.n3981 19.3944
R9764 gnd.n4350 gnd.n3981 19.3944
R9765 gnd.n4350 gnd.n3979 19.3944
R9766 gnd.n4354 gnd.n3979 19.3944
R9767 gnd.n4354 gnd.n3975 19.3944
R9768 gnd.n4364 gnd.n3975 19.3944
R9769 gnd.n4364 gnd.n3973 19.3944
R9770 gnd.n4368 gnd.n3973 19.3944
R9771 gnd.n4368 gnd.n3964 19.3944
R9772 gnd.n4403 gnd.n3964 19.3944
R9773 gnd.n4403 gnd.n3965 19.3944
R9774 gnd.n4399 gnd.n3965 19.3944
R9775 gnd.n4399 gnd.n4398 19.3944
R9776 gnd.n4398 gnd.n4397 19.3944
R9777 gnd.n4397 gnd.n3970 19.3944
R9778 gnd.n4393 gnd.n3970 19.3944
R9779 gnd.n4393 gnd.n3950 19.3944
R9780 gnd.n4453 gnd.n3950 19.3944
R9781 gnd.n4453 gnd.n3948 19.3944
R9782 gnd.n4457 gnd.n3948 19.3944
R9783 gnd.n4457 gnd.n3944 19.3944
R9784 gnd.n4467 gnd.n3944 19.3944
R9785 gnd.n4467 gnd.n3942 19.3944
R9786 gnd.n4471 gnd.n3942 19.3944
R9787 gnd.n4471 gnd.n3939 19.3944
R9788 gnd.n4762 gnd.n3939 19.3944
R9789 gnd.n4762 gnd.n3937 19.3944
R9790 gnd.n4766 gnd.n3937 19.3944
R9791 gnd.n6504 gnd.n2465 19.3944
R9792 gnd.n4046 gnd.n2465 19.3944
R9793 gnd.n4047 gnd.n4046 19.3944
R9794 gnd.n4049 gnd.n4047 19.3944
R9795 gnd.n4050 gnd.n4049 19.3944
R9796 gnd.n4053 gnd.n4050 19.3944
R9797 gnd.n4054 gnd.n4053 19.3944
R9798 gnd.n4056 gnd.n4054 19.3944
R9799 gnd.n4057 gnd.n4056 19.3944
R9800 gnd.n4060 gnd.n4057 19.3944
R9801 gnd.n4061 gnd.n4060 19.3944
R9802 gnd.n4063 gnd.n4061 19.3944
R9803 gnd.n4064 gnd.n4063 19.3944
R9804 gnd.n4067 gnd.n4064 19.3944
R9805 gnd.n4068 gnd.n4067 19.3944
R9806 gnd.n4173 gnd.n4068 19.3944
R9807 gnd.n4174 gnd.n4173 19.3944
R9808 gnd.n4176 gnd.n4174 19.3944
R9809 gnd.n4177 gnd.n4176 19.3944
R9810 gnd.n4181 gnd.n4177 19.3944
R9811 gnd.n4181 gnd.n4180 19.3944
R9812 gnd.n4180 gnd.n4179 19.3944
R9813 gnd.n4179 gnd.n4031 19.3944
R9814 gnd.n4231 gnd.n4031 19.3944
R9815 gnd.n4232 gnd.n4231 19.3944
R9816 gnd.n4234 gnd.n4232 19.3944
R9817 gnd.n4235 gnd.n4234 19.3944
R9818 gnd.n4245 gnd.n4235 19.3944
R9819 gnd.n4245 gnd.n4244 19.3944
R9820 gnd.n4244 gnd.n4243 19.3944
R9821 gnd.n4243 gnd.n4009 19.3944
R9822 gnd.n4289 gnd.n4009 19.3944
R9823 gnd.n4290 gnd.n4289 19.3944
R9824 gnd.n4291 gnd.n4290 19.3944
R9825 gnd.n4296 gnd.n4291 19.3944
R9826 gnd.n4296 gnd.n4294 19.3944
R9827 gnd.n4294 gnd.n4293 19.3944
R9828 gnd.n4293 gnd.n4292 19.3944
R9829 gnd.n4292 gnd.n3977 19.3944
R9830 gnd.n4358 gnd.n3977 19.3944
R9831 gnd.n4359 gnd.n4358 19.3944
R9832 gnd.n4360 gnd.n4359 19.3944
R9833 gnd.n4360 gnd.n3971 19.3944
R9834 gnd.n4372 gnd.n3971 19.3944
R9835 gnd.n4373 gnd.n4372 19.3944
R9836 gnd.n4374 gnd.n4373 19.3944
R9837 gnd.n4375 gnd.n4374 19.3944
R9838 gnd.n4379 gnd.n4375 19.3944
R9839 gnd.n4380 gnd.n4379 19.3944
R9840 gnd.n4384 gnd.n4380 19.3944
R9841 gnd.n4385 gnd.n4384 19.3944
R9842 gnd.n4389 gnd.n4385 19.3944
R9843 gnd.n4389 gnd.n4388 19.3944
R9844 gnd.n4388 gnd.n4387 19.3944
R9845 gnd.n4387 gnd.n3946 19.3944
R9846 gnd.n4461 gnd.n3946 19.3944
R9847 gnd.n4462 gnd.n4461 19.3944
R9848 gnd.n4463 gnd.n4462 19.3944
R9849 gnd.n4463 gnd.n3940 19.3944
R9850 gnd.n4475 gnd.n3940 19.3944
R9851 gnd.n4476 gnd.n4475 19.3944
R9852 gnd.n4758 gnd.n4476 19.3944
R9853 gnd.n4758 gnd.n4757 19.3944
R9854 gnd.n4757 gnd.n4756 19.3944
R9855 gnd.n2484 gnd.n2463 19.3944
R9856 gnd.n2485 gnd.n2484 19.3944
R9857 gnd.n6493 gnd.n2485 19.3944
R9858 gnd.n6493 gnd.n6492 19.3944
R9859 gnd.n6492 gnd.n6491 19.3944
R9860 gnd.n6491 gnd.n2489 19.3944
R9861 gnd.n6481 gnd.n2489 19.3944
R9862 gnd.n6481 gnd.n6480 19.3944
R9863 gnd.n6480 gnd.n6479 19.3944
R9864 gnd.n6479 gnd.n2508 19.3944
R9865 gnd.n6469 gnd.n2508 19.3944
R9866 gnd.n6469 gnd.n6468 19.3944
R9867 gnd.n6468 gnd.n6467 19.3944
R9868 gnd.n6467 gnd.n2527 19.3944
R9869 gnd.n6457 gnd.n2527 19.3944
R9870 gnd.n6457 gnd.n6456 19.3944
R9871 gnd.n6456 gnd.n6455 19.3944
R9872 gnd.n6455 gnd.n2547 19.3944
R9873 gnd.n6445 gnd.n2547 19.3944
R9874 gnd.n6445 gnd.n6444 19.3944
R9875 gnd.n6444 gnd.n6443 19.3944
R9876 gnd.n6443 gnd.n2567 19.3944
R9877 gnd.n6433 gnd.n2567 19.3944
R9878 gnd.n6433 gnd.n6432 19.3944
R9879 gnd.n6432 gnd.n6431 19.3944
R9880 gnd.n6431 gnd.n2587 19.3944
R9881 gnd.n6421 gnd.n2587 19.3944
R9882 gnd.n6421 gnd.n6420 19.3944
R9883 gnd.n6420 gnd.n6419 19.3944
R9884 gnd.n6419 gnd.n2606 19.3944
R9885 gnd.n4240 gnd.n2606 19.3944
R9886 gnd.n4240 gnd.n4005 19.3944
R9887 gnd.n4301 gnd.n4005 19.3944
R9888 gnd.n4301 gnd.n4300 19.3944
R9889 gnd.n4300 gnd.n4299 19.3944
R9890 gnd.n4299 gnd.n2630 19.3944
R9891 gnd.n6408 gnd.n2630 19.3944
R9892 gnd.n6408 gnd.n6407 19.3944
R9893 gnd.n6407 gnd.n6406 19.3944
R9894 gnd.n6406 gnd.n2634 19.3944
R9895 gnd.n6396 gnd.n2634 19.3944
R9896 gnd.n6396 gnd.n6395 19.3944
R9897 gnd.n6395 gnd.n6394 19.3944
R9898 gnd.n6394 gnd.n2652 19.3944
R9899 gnd.n6384 gnd.n2652 19.3944
R9900 gnd.n6384 gnd.n6383 19.3944
R9901 gnd.n6383 gnd.n6382 19.3944
R9902 gnd.n6382 gnd.n2673 19.3944
R9903 gnd.n6372 gnd.n2673 19.3944
R9904 gnd.n6372 gnd.n6371 19.3944
R9905 gnd.n6371 gnd.n6370 19.3944
R9906 gnd.n6370 gnd.n2692 19.3944
R9907 gnd.n6360 gnd.n2692 19.3944
R9908 gnd.n6360 gnd.n6359 19.3944
R9909 gnd.n6359 gnd.n6358 19.3944
R9910 gnd.n6358 gnd.n2713 19.3944
R9911 gnd.n6348 gnd.n2713 19.3944
R9912 gnd.n6348 gnd.n6347 19.3944
R9913 gnd.n6347 gnd.n6346 19.3944
R9914 gnd.n6346 gnd.n2732 19.3944
R9915 gnd.n6336 gnd.n2732 19.3944
R9916 gnd.n6336 gnd.n6335 19.3944
R9917 gnd.n6335 gnd.n6334 19.3944
R9918 gnd.n6334 gnd.n2753 19.3944
R9919 gnd.n6326 gnd.n2763 19.3944
R9920 gnd.n6321 gnd.n2763 19.3944
R9921 gnd.n6321 gnd.n6320 19.3944
R9922 gnd.n6320 gnd.n6319 19.3944
R9923 gnd.n6319 gnd.n6316 19.3944
R9924 gnd.n6316 gnd.n6315 19.3944
R9925 gnd.n6315 gnd.n6312 19.3944
R9926 gnd.n6312 gnd.n6311 19.3944
R9927 gnd.n6311 gnd.n6308 19.3944
R9928 gnd.n6308 gnd.n6307 19.3944
R9929 gnd.n6307 gnd.n6304 19.3944
R9930 gnd.n6304 gnd.n6303 19.3944
R9931 gnd.n6303 gnd.n6300 19.3944
R9932 gnd.n6300 gnd.n6299 19.3944
R9933 gnd.n6299 gnd.n6296 19.3944
R9934 gnd.n6296 gnd.n6295 19.3944
R9935 gnd.n6295 gnd.n6292 19.3944
R9936 gnd.n4704 gnd.n4670 19.3944
R9937 gnd.n4708 gnd.n4670 19.3944
R9938 gnd.n4711 gnd.n4708 19.3944
R9939 gnd.n4714 gnd.n4711 19.3944
R9940 gnd.n4714 gnd.n4668 19.3944
R9941 gnd.n4718 gnd.n4668 19.3944
R9942 gnd.n4721 gnd.n4718 19.3944
R9943 gnd.n4724 gnd.n4721 19.3944
R9944 gnd.n4724 gnd.n4666 19.3944
R9945 gnd.n4728 gnd.n4666 19.3944
R9946 gnd.n4731 gnd.n4728 19.3944
R9947 gnd.n4734 gnd.n4731 19.3944
R9948 gnd.n4734 gnd.n4664 19.3944
R9949 gnd.n4738 gnd.n4664 19.3944
R9950 gnd.n4741 gnd.n4738 19.3944
R9951 gnd.n4744 gnd.n4741 19.3944
R9952 gnd.n4744 gnd.n4662 19.3944
R9953 gnd.n4749 gnd.n4662 19.3944
R9954 gnd.n4682 gnd.n2832 19.3944
R9955 gnd.n4685 gnd.n4682 19.3944
R9956 gnd.n4685 gnd.n4677 19.3944
R9957 gnd.n4689 gnd.n4677 19.3944
R9958 gnd.n4692 gnd.n4689 19.3944
R9959 gnd.n4695 gnd.n4692 19.3944
R9960 gnd.n4695 gnd.n4675 19.3944
R9961 gnd.n4700 gnd.n4675 19.3944
R9962 gnd.n6290 gnd.n6287 19.3944
R9963 gnd.n6287 gnd.n6286 19.3944
R9964 gnd.n6286 gnd.n6283 19.3944
R9965 gnd.n6283 gnd.n6282 19.3944
R9966 gnd.n6282 gnd.n6279 19.3944
R9967 gnd.n6279 gnd.n6278 19.3944
R9968 gnd.n6278 gnd.n6275 19.3944
R9969 gnd.n6499 gnd.n2471 19.3944
R9970 gnd.n6499 gnd.n6498 19.3944
R9971 gnd.n6498 gnd.n6497 19.3944
R9972 gnd.n6497 gnd.n2476 19.3944
R9973 gnd.n6487 gnd.n2476 19.3944
R9974 gnd.n6487 gnd.n6486 19.3944
R9975 gnd.n6486 gnd.n6485 19.3944
R9976 gnd.n6485 gnd.n2499 19.3944
R9977 gnd.n6475 gnd.n2499 19.3944
R9978 gnd.n6475 gnd.n6474 19.3944
R9979 gnd.n6474 gnd.n6473 19.3944
R9980 gnd.n6473 gnd.n2517 19.3944
R9981 gnd.n6463 gnd.n2517 19.3944
R9982 gnd.n6463 gnd.n6462 19.3944
R9983 gnd.n6462 gnd.n6461 19.3944
R9984 gnd.n6461 gnd.n2538 19.3944
R9985 gnd.n6451 gnd.n2538 19.3944
R9986 gnd.n6451 gnd.n6450 19.3944
R9987 gnd.n6450 gnd.n6449 19.3944
R9988 gnd.n6449 gnd.n2557 19.3944
R9989 gnd.n6439 gnd.n2557 19.3944
R9990 gnd.n6439 gnd.n6438 19.3944
R9991 gnd.n6438 gnd.n6437 19.3944
R9992 gnd.n6437 gnd.n2578 19.3944
R9993 gnd.n6427 gnd.n2578 19.3944
R9994 gnd.n6427 gnd.n6426 19.3944
R9995 gnd.n6426 gnd.n6425 19.3944
R9996 gnd.n6415 gnd.n2613 19.3944
R9997 gnd.n4236 gnd.n2614 19.3944
R9998 gnd.n4001 gnd.n4000 19.3944
R9999 gnd.n4307 gnd.n4306 19.3944
R10000 gnd.n6412 gnd.n2620 19.3944
R10001 gnd.n6412 gnd.n2621 19.3944
R10002 gnd.n6402 gnd.n2621 19.3944
R10003 gnd.n6402 gnd.n6401 19.3944
R10004 gnd.n6401 gnd.n6400 19.3944
R10005 gnd.n6400 gnd.n2643 19.3944
R10006 gnd.n6390 gnd.n2643 19.3944
R10007 gnd.n6390 gnd.n6389 19.3944
R10008 gnd.n6389 gnd.n6388 19.3944
R10009 gnd.n6388 gnd.n2663 19.3944
R10010 gnd.n6378 gnd.n2663 19.3944
R10011 gnd.n6378 gnd.n6377 19.3944
R10012 gnd.n6377 gnd.n6376 19.3944
R10013 gnd.n6376 gnd.n2683 19.3944
R10014 gnd.n6366 gnd.n2683 19.3944
R10015 gnd.n6366 gnd.n6365 19.3944
R10016 gnd.n6365 gnd.n6364 19.3944
R10017 gnd.n6364 gnd.n2703 19.3944
R10018 gnd.n6354 gnd.n2703 19.3944
R10019 gnd.n6354 gnd.n6353 19.3944
R10020 gnd.n6353 gnd.n6352 19.3944
R10021 gnd.n6352 gnd.n2723 19.3944
R10022 gnd.n6342 gnd.n2723 19.3944
R10023 gnd.n6342 gnd.n6341 19.3944
R10024 gnd.n6341 gnd.n6340 19.3944
R10025 gnd.n6340 gnd.n2743 19.3944
R10026 gnd.n6330 gnd.n2743 19.3944
R10027 gnd.n6330 gnd.n6329 19.3944
R10028 gnd.n6883 gnd.n6882 19.3944
R10029 gnd.n6882 gnd.n6881 19.3944
R10030 gnd.n6881 gnd.n791 19.3944
R10031 gnd.n6875 gnd.n791 19.3944
R10032 gnd.n6875 gnd.n6874 19.3944
R10033 gnd.n6874 gnd.n6873 19.3944
R10034 gnd.n6873 gnd.n799 19.3944
R10035 gnd.n6867 gnd.n799 19.3944
R10036 gnd.n6867 gnd.n6866 19.3944
R10037 gnd.n6866 gnd.n6865 19.3944
R10038 gnd.n6865 gnd.n807 19.3944
R10039 gnd.n6859 gnd.n807 19.3944
R10040 gnd.n6859 gnd.n6858 19.3944
R10041 gnd.n6858 gnd.n6857 19.3944
R10042 gnd.n6857 gnd.n815 19.3944
R10043 gnd.n6851 gnd.n815 19.3944
R10044 gnd.n6851 gnd.n6850 19.3944
R10045 gnd.n6850 gnd.n6849 19.3944
R10046 gnd.n6849 gnd.n823 19.3944
R10047 gnd.n6843 gnd.n823 19.3944
R10048 gnd.n6843 gnd.n6842 19.3944
R10049 gnd.n6842 gnd.n6841 19.3944
R10050 gnd.n6841 gnd.n831 19.3944
R10051 gnd.n6835 gnd.n831 19.3944
R10052 gnd.n6835 gnd.n6834 19.3944
R10053 gnd.n6834 gnd.n6833 19.3944
R10054 gnd.n6833 gnd.n839 19.3944
R10055 gnd.n6827 gnd.n839 19.3944
R10056 gnd.n6827 gnd.n6826 19.3944
R10057 gnd.n6826 gnd.n6825 19.3944
R10058 gnd.n6825 gnd.n847 19.3944
R10059 gnd.n6819 gnd.n847 19.3944
R10060 gnd.n6819 gnd.n6818 19.3944
R10061 gnd.n6818 gnd.n6817 19.3944
R10062 gnd.n6817 gnd.n855 19.3944
R10063 gnd.n6811 gnd.n855 19.3944
R10064 gnd.n6811 gnd.n6810 19.3944
R10065 gnd.n6810 gnd.n6809 19.3944
R10066 gnd.n6809 gnd.n863 19.3944
R10067 gnd.n6803 gnd.n863 19.3944
R10068 gnd.n6803 gnd.n6802 19.3944
R10069 gnd.n6802 gnd.n6801 19.3944
R10070 gnd.n6801 gnd.n871 19.3944
R10071 gnd.n6795 gnd.n871 19.3944
R10072 gnd.n6795 gnd.n6794 19.3944
R10073 gnd.n6794 gnd.n6793 19.3944
R10074 gnd.n6793 gnd.n879 19.3944
R10075 gnd.n6787 gnd.n879 19.3944
R10076 gnd.n6787 gnd.n6786 19.3944
R10077 gnd.n6786 gnd.n6785 19.3944
R10078 gnd.n6785 gnd.n887 19.3944
R10079 gnd.n6779 gnd.n887 19.3944
R10080 gnd.n6779 gnd.n6778 19.3944
R10081 gnd.n6778 gnd.n6777 19.3944
R10082 gnd.n6777 gnd.n895 19.3944
R10083 gnd.n6771 gnd.n895 19.3944
R10084 gnd.n6771 gnd.n6770 19.3944
R10085 gnd.n6770 gnd.n6769 19.3944
R10086 gnd.n6769 gnd.n903 19.3944
R10087 gnd.n6763 gnd.n903 19.3944
R10088 gnd.n6763 gnd.n6762 19.3944
R10089 gnd.n6762 gnd.n6761 19.3944
R10090 gnd.n6761 gnd.n911 19.3944
R10091 gnd.n6755 gnd.n911 19.3944
R10092 gnd.n6755 gnd.n6754 19.3944
R10093 gnd.n6754 gnd.n6753 19.3944
R10094 gnd.n6753 gnd.n919 19.3944
R10095 gnd.n6747 gnd.n919 19.3944
R10096 gnd.n6747 gnd.n6746 19.3944
R10097 gnd.n6746 gnd.n6745 19.3944
R10098 gnd.n6745 gnd.n927 19.3944
R10099 gnd.n6739 gnd.n927 19.3944
R10100 gnd.n6739 gnd.n6738 19.3944
R10101 gnd.n6738 gnd.n6737 19.3944
R10102 gnd.n6737 gnd.n935 19.3944
R10103 gnd.n6731 gnd.n935 19.3944
R10104 gnd.n6731 gnd.n6730 19.3944
R10105 gnd.n6730 gnd.n6729 19.3944
R10106 gnd.n6729 gnd.n943 19.3944
R10107 gnd.n6723 gnd.n943 19.3944
R10108 gnd.n6723 gnd.n6722 19.3944
R10109 gnd.n6722 gnd.n6721 19.3944
R10110 gnd.n6721 gnd.n951 19.3944
R10111 gnd.n4197 gnd.n951 19.3944
R10112 gnd.n4520 gnd.n4484 19.3944
R10113 gnd.n4516 gnd.n4484 19.3944
R10114 gnd.n4516 gnd.n4515 19.3944
R10115 gnd.n4515 gnd.n4514 19.3944
R10116 gnd.n4514 gnd.n4488 19.3944
R10117 gnd.n4510 gnd.n4488 19.3944
R10118 gnd.n4510 gnd.n4509 19.3944
R10119 gnd.n4509 gnd.n4508 19.3944
R10120 gnd.n4508 gnd.n4492 19.3944
R10121 gnd.n4504 gnd.n4492 19.3944
R10122 gnd.n4504 gnd.n4503 19.3944
R10123 gnd.n4503 gnd.n4502 19.3944
R10124 gnd.n4502 gnd.n4496 19.3944
R10125 gnd.n4498 gnd.n4496 19.3944
R10126 gnd.n4498 gnd.n3852 19.3944
R10127 gnd.n3852 gnd.n3850 19.3944
R10128 gnd.n4863 gnd.n3850 19.3944
R10129 gnd.n4863 gnd.n3848 19.3944
R10130 gnd.n4867 gnd.n3848 19.3944
R10131 gnd.n4867 gnd.n3764 19.3944
R10132 gnd.n4902 gnd.n3764 19.3944
R10133 gnd.n4902 gnd.n3761 19.3944
R10134 gnd.n4909 gnd.n3761 19.3944
R10135 gnd.n4909 gnd.n3762 19.3944
R10136 gnd.n4905 gnd.n3762 19.3944
R10137 gnd.n4905 gnd.n3742 19.3944
R10138 gnd.n4933 gnd.n3742 19.3944
R10139 gnd.n4933 gnd.n3739 19.3944
R10140 gnd.n4943 gnd.n3739 19.3944
R10141 gnd.n4943 gnd.n3740 19.3944
R10142 gnd.n4939 gnd.n3740 19.3944
R10143 gnd.n4939 gnd.n4938 19.3944
R10144 gnd.n4938 gnd.n3692 19.3944
R10145 gnd.n5013 gnd.n3692 19.3944
R10146 gnd.n5013 gnd.n3689 19.3944
R10147 gnd.n5018 gnd.n3689 19.3944
R10148 gnd.n5018 gnd.n3690 19.3944
R10149 gnd.n3690 gnd.n3665 19.3944
R10150 gnd.n5059 gnd.n3665 19.3944
R10151 gnd.n5059 gnd.n3662 19.3944
R10152 gnd.n5089 gnd.n3662 19.3944
R10153 gnd.n5089 gnd.n3663 19.3944
R10154 gnd.n5085 gnd.n3663 19.3944
R10155 gnd.n5085 gnd.n5084 19.3944
R10156 gnd.n5084 gnd.n5083 19.3944
R10157 gnd.n5083 gnd.n5067 19.3944
R10158 gnd.n5079 gnd.n5067 19.3944
R10159 gnd.n5079 gnd.n5078 19.3944
R10160 gnd.n5078 gnd.n5077 19.3944
R10161 gnd.n5077 gnd.n5072 19.3944
R10162 gnd.n5073 gnd.n5072 19.3944
R10163 gnd.n5073 gnd.n3590 19.3944
R10164 gnd.n5190 gnd.n3590 19.3944
R10165 gnd.n5190 gnd.n3587 19.3944
R10166 gnd.n5217 gnd.n3587 19.3944
R10167 gnd.n5217 gnd.n3588 19.3944
R10168 gnd.n5213 gnd.n3588 19.3944
R10169 gnd.n5213 gnd.n5212 19.3944
R10170 gnd.n5212 gnd.n5211 19.3944
R10171 gnd.n5211 gnd.n5198 19.3944
R10172 gnd.n5207 gnd.n5198 19.3944
R10173 gnd.n5207 gnd.n5206 19.3944
R10174 gnd.n5206 gnd.n5205 19.3944
R10175 gnd.n5205 gnd.n5202 19.3944
R10176 gnd.n5202 gnd.n3458 19.3944
R10177 gnd.n5416 gnd.n3458 19.3944
R10178 gnd.n5416 gnd.n3456 19.3944
R10179 gnd.n5420 gnd.n3456 19.3944
R10180 gnd.n5420 gnd.n3444 19.3944
R10181 gnd.n5432 gnd.n3444 19.3944
R10182 gnd.n5432 gnd.n3442 19.3944
R10183 gnd.n5436 gnd.n3442 19.3944
R10184 gnd.n5436 gnd.n3431 19.3944
R10185 gnd.n5448 gnd.n3431 19.3944
R10186 gnd.n5448 gnd.n3429 19.3944
R10187 gnd.n5452 gnd.n3429 19.3944
R10188 gnd.n5452 gnd.n3419 19.3944
R10189 gnd.n5467 gnd.n3419 19.3944
R10190 gnd.n5467 gnd.n3417 19.3944
R10191 gnd.n5471 gnd.n3417 19.3944
R10192 gnd.n5471 gnd.n2999 19.3944
R10193 gnd.n6093 gnd.n2999 19.3944
R10194 gnd.n6090 gnd.n6089 19.3944
R10195 gnd.n6089 gnd.n6088 19.3944
R10196 gnd.n6088 gnd.n3004 19.3944
R10197 gnd.n6084 gnd.n3004 19.3944
R10198 gnd.n6084 gnd.n6083 19.3944
R10199 gnd.n6083 gnd.n6082 19.3944
R10200 gnd.n6082 gnd.n3009 19.3944
R10201 gnd.n6077 gnd.n3009 19.3944
R10202 gnd.n6077 gnd.n6076 19.3944
R10203 gnd.n6076 gnd.n3014 19.3944
R10204 gnd.n6069 gnd.n3014 19.3944
R10205 gnd.n6069 gnd.n6068 19.3944
R10206 gnd.n6068 gnd.n3023 19.3944
R10207 gnd.n6061 gnd.n3023 19.3944
R10208 gnd.n6061 gnd.n6060 19.3944
R10209 gnd.n6060 gnd.n3031 19.3944
R10210 gnd.n6053 gnd.n3031 19.3944
R10211 gnd.n6053 gnd.n6052 19.3944
R10212 gnd.n6052 gnd.n3039 19.3944
R10213 gnd.n6045 gnd.n3039 19.3944
R10214 gnd.n6045 gnd.n6044 19.3944
R10215 gnd.n6044 gnd.n3047 19.3944
R10216 gnd.n6037 gnd.n3047 19.3944
R10217 gnd.n6037 gnd.n6036 19.3944
R10218 gnd.n3405 gnd.n3384 19.3944
R10219 gnd.n5579 gnd.n3384 19.3944
R10220 gnd.n5579 gnd.n5578 19.3944
R10221 gnd.n1836 gnd.t135 18.8012
R10222 gnd.n1873 gnd.t348 18.8012
R10223 gnd.n4859 gnd.t115 18.8012
R10224 gnd.n1706 gnd.n1705 18.4825
R10225 gnd.n6717 gnd.n953 18.4825
R10226 gnd.n4869 gnd.n2909 18.4825
R10227 gnd.n5021 gnd.n5020 18.4825
R10228 gnd.n3638 gnd.n3632 18.4825
R10229 gnd.n3552 gnd.n3546 18.4825
R10230 gnd.n5975 gnd.n5974 18.4247
R10231 gnd.n6275 gnd.n6274 18.4247
R10232 gnd.n6033 gnd.n6032 18.2308
R10233 gnd.n4609 gnd.n4594 18.2308
R10234 gnd.n7669 gnd.n7620 18.2308
R10235 gnd.n4132 gnd.n4131 18.2308
R10236 gnd.t362 gnd.n1385 18.1639
R10237 gnd.n6204 gnd.n6203 17.9517
R10238 gnd.n5402 gnd.n5401 17.9517
R10239 gnd.t269 gnd.n3454 17.8452
R10240 gnd.n1414 gnd.t137 17.5266
R10241 gnd.n6200 gnd.n2896 17.2079
R10242 gnd.n4872 gnd.t168 17.2079
R10243 gnd.n1825 gnd.t102 16.8893
R10244 gnd.n5957 gnd.n5954 16.6793
R10245 gnd.n7781 gnd.n7778 16.6793
R10246 gnd.n6552 gnd.n6549 16.6793
R10247 gnd.n4701 gnd.n4700 16.6793
R10248 gnd.n4171 gnd.n2542 16.5706
R10249 gnd.n6453 gnd.n2549 16.5706
R10250 gnd.n4190 gnd.n4189 16.5706
R10251 gnd.n6447 gnd.n2559 16.5706
R10252 gnd.n4183 gnd.n2562 16.5706
R10253 gnd.n6441 gnd.n2569 16.5706
R10254 gnd.n4220 gnd.n2572 16.5706
R10255 gnd.n4229 gnd.n2582 16.5706
R10256 gnd.n6429 gnd.n2589 16.5706
R10257 gnd.n4254 gnd.n4253 16.5706
R10258 gnd.n6423 gnd.n2598 16.5706
R10259 gnd.n4247 gnd.n2601 16.5706
R10260 gnd.n6417 gnd.n2608 16.5706
R10261 gnd.n4279 gnd.n2611 16.5706
R10262 gnd.n4287 gnd.n4012 16.5706
R10263 gnd.n4303 gnd.n4002 16.5706
R10264 gnd.n4309 gnd.n3995 16.5706
R10265 gnd.n3997 gnd.n3988 16.5706
R10266 gnd.n6410 gnd.n2624 16.5706
R10267 gnd.n4348 gnd.n2627 16.5706
R10268 gnd.n4356 gnd.n2638 16.5706
R10269 gnd.n6398 gnd.n2645 16.5706
R10270 gnd.n4362 gnd.n3976 16.5706
R10271 gnd.n6392 gnd.n2654 16.5706
R10272 gnd.n6386 gnd.n2665 16.5706
R10273 gnd.n4405 gnd.n2668 16.5706
R10274 gnd.n4377 gnd.n2677 16.5706
R10275 gnd.n6374 gnd.n2685 16.5706
R10276 gnd.n4382 gnd.n4381 16.5706
R10277 gnd.n6368 gnd.n2694 16.5706
R10278 gnd.n6362 gnd.n2705 16.5706
R10279 gnd.n4451 gnd.n2708 16.5706
R10280 gnd.n4459 gnd.n2717 16.5706
R10281 gnd.n6350 gnd.n2725 16.5706
R10282 gnd.n4465 gnd.n3945 16.5706
R10283 gnd.n6344 gnd.n2734 16.5706
R10284 gnd.n4473 gnd.n2737 16.5706
R10285 gnd.n6338 gnd.n2745 16.5706
R10286 gnd.n4760 gnd.n2748 16.5706
R10287 gnd.n6332 gnd.n2755 16.5706
R10288 gnd.n4768 gnd.n2758 16.5706
R10289 gnd.n5906 gnd.n3175 16.5706
R10290 gnd.n5563 gnd.n5562 16.5706
R10291 gnd.n5898 gnd.n3184 16.5706
R10292 gnd.n5586 gnd.n3197 16.5706
R10293 gnd.n5892 gnd.n3200 16.5706
R10294 gnd.n5594 gnd.n3210 16.5706
R10295 gnd.n5886 gnd.n3213 16.5706
R10296 gnd.n5601 gnd.n3221 16.5706
R10297 gnd.n5880 gnd.n3224 16.5706
R10298 gnd.n5874 gnd.n3234 16.5706
R10299 gnd.n5616 gnd.n3242 16.5706
R10300 gnd.n5624 gnd.n3251 16.5706
R10301 gnd.n5862 gnd.n3254 16.5706
R10302 gnd.n5631 gnd.n3262 16.5706
R10303 gnd.n5856 gnd.n3265 16.5706
R10304 gnd.n5850 gnd.n3275 16.5706
R10305 gnd.n5646 gnd.n3283 16.5706
R10306 gnd.n5654 gnd.n3292 16.5706
R10307 gnd.n5838 gnd.n3295 16.5706
R10308 gnd.n5661 gnd.n3304 16.5706
R10309 gnd.n5832 gnd.n3307 16.5706
R10310 gnd.n5826 gnd.n3317 16.5706
R10311 gnd.n5821 gnd.n5820 16.5706
R10312 gnd.n5813 gnd.n3328 16.5706
R10313 gnd.n5812 gnd.n3331 16.5706
R10314 gnd.n5807 gnd.n3341 16.5706
R10315 gnd.n3350 gnd.n3348 16.5706
R10316 gnd.n7947 gnd.n103 16.5706
R10317 gnd.n5795 gnd.n5792 16.5706
R10318 gnd.n5722 gnd.n118 16.5706
R10319 gnd.n7939 gnd.n121 16.5706
R10320 gnd.n5784 gnd.n5783 16.5706
R10321 gnd.n7933 gnd.n132 16.5706
R10322 gnd.n5777 gnd.n139 16.5706
R10323 gnd.n5771 gnd.n148 16.5706
R10324 gnd.n7921 gnd.n151 16.5706
R10325 gnd.n5765 gnd.n159 16.5706
R10326 gnd.n7915 gnd.n162 16.5706
R10327 gnd.n7596 gnd.n7595 16.5706
R10328 gnd.n7909 gnd.n171 16.5706
R10329 gnd.n7701 gnd.n179 16.5706
R10330 gnd.n1641 gnd.t171 16.2519
R10331 gnd.n1870 gnd.t91 16.2519
R10332 gnd.n4318 gnd.t77 16.2519
R10333 gnd.n4789 gnd.t228 16.2519
R10334 gnd.t207 gnd.n2994 16.2519
R10335 gnd.n3327 gnd.t86 16.2519
R10336 gnd.n5001 gnd.n5000 15.9333
R10337 gnd.n3619 gnd.n3612 15.9333
R10338 gnd.n256 gnd.n249 15.9333
R10339 gnd.n2309 gnd.n2307 15.6674
R10340 gnd.n2277 gnd.n2275 15.6674
R10341 gnd.n2245 gnd.n2243 15.6674
R10342 gnd.n2214 gnd.n2212 15.6674
R10343 gnd.n2182 gnd.n2180 15.6674
R10344 gnd.n2150 gnd.n2148 15.6674
R10345 gnd.n2118 gnd.n2116 15.6674
R10346 gnd.n2087 gnd.n2085 15.6674
R10347 gnd.n1632 gnd.t171 15.6146
R10348 gnd.n2346 gnd.t281 15.6146
R10349 gnd.t256 gnd.n1001 15.6146
R10350 gnd.t28 gnd.n2657 15.6146
R10351 gnd.t228 gnd.n3898 15.6146
R10352 gnd.n5473 gnd.t207 15.6146
R10353 gnd.n3360 gnd.t105 15.6146
R10354 gnd.n5914 gnd.n5909 15.3217
R10355 gnd.n7736 gnd.n351 15.3217
R10356 gnd.n6509 gnd.n2459 15.3217
R10357 gnd.n4752 gnd.n4750 15.3217
R10358 gnd.n4201 gnd.n2532 15.296
R10359 gnd.n6459 gnd.n2542 15.296
R10360 gnd.n4171 gnd.n2549 15.296
R10361 gnd.n4189 gnd.n2559 15.296
R10362 gnd.n6447 gnd.n2562 15.296
R10363 gnd.n6441 gnd.n2572 15.296
R10364 gnd.n4220 gnd.n4219 15.296
R10365 gnd.n6435 gnd.n2582 15.296
R10366 gnd.n4229 gnd.n2589 15.296
R10367 gnd.n4253 gnd.n2598 15.296
R10368 gnd.n6423 gnd.n2601 15.296
R10369 gnd.n6417 gnd.n2611 15.296
R10370 gnd.n4279 gnd.n4278 15.296
R10371 gnd.n4238 gnd.n4012 15.296
R10372 gnd.n4287 gnd.n4002 15.296
R10373 gnd.n4309 gnd.n3997 15.296
R10374 gnd.n4318 gnd.n3988 15.296
R10375 gnd.n4317 gnd.n2624 15.296
R10376 gnd.n6410 gnd.n2627 15.296
R10377 gnd.n4348 gnd.n4347 15.296
R10378 gnd.n6404 gnd.n2638 15.296
R10379 gnd.n4356 gnd.n2645 15.296
R10380 gnd.n4362 gnd.n2654 15.296
R10381 gnd.n6392 gnd.n2657 15.296
R10382 gnd.n4370 gnd.n2665 15.296
R10383 gnd.n6386 gnd.n2668 15.296
R10384 gnd.n4406 gnd.n4405 15.296
R10385 gnd.n6380 gnd.n2677 15.296
R10386 gnd.n4377 gnd.n2685 15.296
R10387 gnd.n4382 gnd.n2694 15.296
R10388 gnd.n6368 gnd.n2697 15.296
R10389 gnd.n4391 gnd.n2705 15.296
R10390 gnd.n6362 gnd.n2708 15.296
R10391 gnd.n4451 gnd.n4450 15.296
R10392 gnd.n6356 gnd.n2717 15.296
R10393 gnd.n4459 gnd.n2725 15.296
R10394 gnd.n4465 gnd.n2734 15.296
R10395 gnd.n6344 gnd.n2737 15.296
R10396 gnd.n4473 gnd.n2745 15.296
R10397 gnd.n6338 gnd.n2748 15.296
R10398 gnd.n6332 gnd.n2758 15.296
R10399 gnd.n4769 gnd.n4768 15.296
R10400 gnd.t117 gnd.n3733 15.296
R10401 gnd.n5219 gnd.t107 15.296
R10402 gnd.n5906 gnd.n3173 15.296
R10403 gnd.n5562 gnd.n3175 15.296
R10404 gnd.n5586 gnd.n3184 15.296
R10405 gnd.n5892 gnd.n3197 15.296
R10406 gnd.n5594 gnd.n3200 15.296
R10407 gnd.n5886 gnd.n3210 15.296
R10408 gnd.n5880 gnd.n3221 15.296
R10409 gnd.n5609 gnd.n3224 15.296
R10410 gnd.n5874 gnd.n3231 15.296
R10411 gnd.n5616 gnd.n3234 15.296
R10412 gnd.n5868 gnd.n3242 15.296
R10413 gnd.n5624 gnd.n3369 15.296
R10414 gnd.n5862 gnd.n3251 15.296
R10415 gnd.n5856 gnd.n3262 15.296
R10416 gnd.n5639 gnd.n3265 15.296
R10417 gnd.n5850 gnd.n3272 15.296
R10418 gnd.n5646 gnd.n3275 15.296
R10419 gnd.n5844 gnd.n3283 15.296
R10420 gnd.n5654 gnd.n3360 15.296
R10421 gnd.n5838 gnd.n3292 15.296
R10422 gnd.n5832 gnd.n3304 15.296
R10423 gnd.n5681 gnd.n3307 15.296
R10424 gnd.n5826 gnd.n3314 15.296
R10425 gnd.n5821 gnd.n3317 15.296
R10426 gnd.n5820 gnd.n3321 15.296
R10427 gnd.n3328 gnd.n3327 15.296
R10428 gnd.n5813 gnd.n5812 15.296
R10429 gnd.n3350 gnd.n3341 15.296
R10430 gnd.n5801 gnd.n3348 15.296
R10431 gnd.n7947 gnd.n101 15.296
R10432 gnd.n5795 gnd.n103 15.296
R10433 gnd.n7939 gnd.n118 15.296
R10434 gnd.n5783 gnd.n121 15.296
R10435 gnd.n5777 gnd.n132 15.296
R10436 gnd.n7927 gnd.n139 15.296
R10437 gnd.n5771 gnd.n5755 15.296
R10438 gnd.n7921 gnd.n148 15.296
R10439 gnd.n7915 gnd.n159 15.296
R10440 gnd.n7596 gnd.n162 15.296
R10441 gnd.n7701 gnd.n171 15.296
R10442 gnd.n7903 gnd.n179 15.296
R10443 gnd.n7588 gnd.n188 15.296
R10444 gnd.n3479 gnd.n3478 15.0827
R10445 gnd.n2882 gnd.n2877 15.0481
R10446 gnd.n3489 gnd.n3488 15.0481
R10447 gnd.n1139 gnd.t136 14.9773
R10448 gnd.t123 gnd.n2608 14.9773
R10449 gnd.t103 gnd.n2697 14.9773
R10450 gnd.n4993 gnd.t36 14.9773
R10451 gnd.n5135 gnd.t113 14.9773
R10452 gnd.n3369 gnd.t67 14.9773
R10453 gnd.n5792 gnd.t26 14.9773
R10454 gnd.n6200 gnd.n6199 14.6587
R10455 gnd.n4969 gnd.n3721 14.6587
R10456 gnd.n5177 gnd.n3603 14.6587
R10457 gnd.n5406 gnd.n5405 14.6587
R10458 gnd.t389 gnd.n955 14.34
R10459 gnd.n1112 gnd.t376 14.34
R10460 gnd.t8 gnd.n2569 14.34
R10461 gnd.t69 gnd.n151 14.34
R10462 gnd.n1794 gnd.t12 13.7027
R10463 gnd.n1498 gnd.n1497 13.5763
R10464 gnd.n6680 gnd.n1014 13.5763
R10465 gnd.n1706 gnd.n1444 13.384
R10466 gnd.n6193 gnd.n2909 13.384
R10467 gnd.n4961 gnd.n4960 13.384
R10468 gnd.n4946 gnd.t345 13.384
R10469 gnd.n5188 gnd.t314 13.384
R10470 gnd.n5170 gnd.n5169 13.384
R10471 gnd.n5267 gnd.n3552 13.384
R10472 gnd.n2893 gnd.n2874 13.1884
R10473 gnd.n2888 gnd.n2887 13.1884
R10474 gnd.n2887 gnd.n2886 13.1884
R10475 gnd.n3482 gnd.n3477 13.1884
R10476 gnd.n3483 gnd.n3482 13.1884
R10477 gnd.n2889 gnd.n2876 13.146
R10478 gnd.n2885 gnd.n2876 13.146
R10479 gnd.n3481 gnd.n3480 13.146
R10480 gnd.n3481 gnd.n3476 13.146
R10481 gnd.n2310 gnd.n2306 12.8005
R10482 gnd.n2278 gnd.n2274 12.8005
R10483 gnd.n2246 gnd.n2242 12.8005
R10484 gnd.n2215 gnd.n2211 12.8005
R10485 gnd.n2183 gnd.n2179 12.8005
R10486 gnd.n2151 gnd.n2147 12.8005
R10487 gnd.n2119 gnd.n2115 12.8005
R10488 gnd.n2088 gnd.n2084 12.8005
R10489 gnd.n5245 gnd.t187 12.7467
R10490 gnd.n6477 gnd.t24 12.4281
R10491 gnd.n6356 gnd.t49 12.4281
R10492 gnd.n5609 gnd.t30 12.4281
R10493 gnd.n7885 gnd.t42 12.4281
R10494 gnd.n1497 gnd.n1492 12.4126
R10495 gnd.n6676 gnd.n1014 12.4126
R10496 gnd.n6267 gnd.n6204 12.1761
R10497 gnd.n5401 gnd.n5400 12.1761
R10498 gnd.n4930 gnd.n3745 12.1094
R10499 gnd.n5230 gnd.n3576 12.1094
R10500 gnd.n5259 gnd.n5258 12.1094
R10501 gnd.n2314 gnd.n2313 12.0247
R10502 gnd.n2282 gnd.n2281 12.0247
R10503 gnd.n2250 gnd.n2249 12.0247
R10504 gnd.n2219 gnd.n2218 12.0247
R10505 gnd.n2187 gnd.n2186 12.0247
R10506 gnd.n2155 gnd.n2154 12.0247
R10507 gnd.n2123 gnd.n2122 12.0247
R10508 gnd.n2092 gnd.n2091 12.0247
R10509 gnd.n6453 gnd.t98 11.7908
R10510 gnd.n6380 gnd.t16 11.7908
R10511 gnd.t197 gnd.n2755 11.7908
R10512 gnd.t340 gnd.t313 11.7908
R10513 gnd.t146 gnd.t155 11.7908
R10514 gnd.n5563 gnd.t175 11.7908
R10515 gnd.n5639 gnd.t10 11.7908
R10516 gnd.n7909 gnd.t5 11.7908
R10517 gnd.t156 gnd.n3715 11.4721
R10518 gnd.n5178 gnd.t334 11.4721
R10519 gnd.n2317 gnd.n2304 11.249
R10520 gnd.n2285 gnd.n2272 11.249
R10521 gnd.n2253 gnd.n2240 11.249
R10522 gnd.n2222 gnd.n2209 11.249
R10523 gnd.n2190 gnd.n2177 11.249
R10524 gnd.n2158 gnd.n2145 11.249
R10525 gnd.n2126 gnd.n2113 11.249
R10526 gnd.n2095 gnd.n2082 11.249
R10527 gnd.n1784 gnd.t12 11.1535
R10528 gnd.n6429 gnd.t47 11.1535
R10529 gnd.n6404 gnd.t3 11.1535
R10530 gnd.n3892 gnd.t310 11.1535
R10531 gnd.n4947 gnd.t88 11.1535
R10532 gnd.t338 gnd.n3592 11.1535
R10533 gnd.n5454 gnd.t287 11.1535
R10534 gnd.n5681 gnd.t34 11.1535
R10535 gnd.n7933 gnd.t72 11.1535
R10536 gnd.n4911 gnd.t241 10.8348
R10537 gnd.n4922 gnd.n3751 10.8348
R10538 gnd.n4922 gnd.n4921 10.8348
R10539 gnd.n5093 gnd.n5092 10.8348
R10540 gnd.n5092 gnd.n3652 10.8348
R10541 gnd.n5238 gnd.n3569 10.8348
R10542 gnd.n5239 gnd.n5238 10.8348
R10543 gnd.n5917 gnd.n5914 10.6672
R10544 gnd.n7739 gnd.n7736 10.6672
R10545 gnd.n6512 gnd.n6509 10.6672
R10546 gnd.n4750 gnd.n4749 10.6672
R10547 gnd.n5335 gnd.n3519 10.6151
R10548 gnd.n5335 gnd.n5334 10.6151
R10549 gnd.n5332 gnd.n3523 10.6151
R10550 gnd.n5327 gnd.n3523 10.6151
R10551 gnd.n5327 gnd.n5326 10.6151
R10552 gnd.n5326 gnd.n5325 10.6151
R10553 gnd.n5325 gnd.n3526 10.6151
R10554 gnd.n5320 gnd.n3526 10.6151
R10555 gnd.n5320 gnd.n5319 10.6151
R10556 gnd.n5319 gnd.n5318 10.6151
R10557 gnd.n5318 gnd.n3529 10.6151
R10558 gnd.n5313 gnd.n3529 10.6151
R10559 gnd.n5313 gnd.n5312 10.6151
R10560 gnd.n5312 gnd.n5311 10.6151
R10561 gnd.n5311 gnd.n3532 10.6151
R10562 gnd.n5306 gnd.n3532 10.6151
R10563 gnd.n5306 gnd.n5305 10.6151
R10564 gnd.n5305 gnd.n5304 10.6151
R10565 gnd.n5304 gnd.n3535 10.6151
R10566 gnd.n5299 gnd.n3535 10.6151
R10567 gnd.n5299 gnd.n5298 10.6151
R10568 gnd.n5298 gnd.n5297 10.6151
R10569 gnd.n5297 gnd.n3538 10.6151
R10570 gnd.n5292 gnd.n3538 10.6151
R10571 gnd.n5292 gnd.n5291 10.6151
R10572 gnd.n5291 gnd.n5290 10.6151
R10573 gnd.n5290 gnd.n3541 10.6151
R10574 gnd.n5285 gnd.n3541 10.6151
R10575 gnd.n5285 gnd.n5284 10.6151
R10576 gnd.n5284 gnd.n5283 10.6151
R10577 gnd.n3845 gnd.n3844 10.6151
R10578 gnd.n3846 gnd.n3845 10.6151
R10579 gnd.n4874 gnd.n3846 10.6151
R10580 gnd.n4875 gnd.n4874 10.6151
R10581 gnd.n4891 gnd.n4875 10.6151
R10582 gnd.n4891 gnd.n4890 10.6151
R10583 gnd.n4890 gnd.n4889 10.6151
R10584 gnd.n4889 gnd.n4888 10.6151
R10585 gnd.n4888 gnd.n4886 10.6151
R10586 gnd.n4886 gnd.n4885 10.6151
R10587 gnd.n4885 gnd.n4883 10.6151
R10588 gnd.n4883 gnd.n4882 10.6151
R10589 gnd.n4882 gnd.n4876 10.6151
R10590 gnd.n4876 gnd.n3736 10.6151
R10591 gnd.n4952 gnd.n3736 10.6151
R10592 gnd.n4952 gnd.n4951 10.6151
R10593 gnd.n4951 gnd.n4950 10.6151
R10594 gnd.n4950 gnd.n4949 10.6151
R10595 gnd.n4949 gnd.n3738 10.6151
R10596 gnd.n3738 gnd.n3737 10.6151
R10597 gnd.n3737 gnd.n3713 10.6151
R10598 gnd.n4979 gnd.n3713 10.6151
R10599 gnd.n4980 gnd.n4979 10.6151
R10600 gnd.n4981 gnd.n4980 10.6151
R10601 gnd.n4987 gnd.n4981 10.6151
R10602 gnd.n4988 gnd.n4987 10.6151
R10603 gnd.n4989 gnd.n4988 10.6151
R10604 gnd.n4989 gnd.n3685 10.6151
R10605 gnd.n5023 gnd.n3685 10.6151
R10606 gnd.n5024 gnd.n5023 10.6151
R10607 gnd.n5025 gnd.n5024 10.6151
R10608 gnd.n5037 gnd.n5025 10.6151
R10609 gnd.n5037 gnd.n5036 10.6151
R10610 gnd.n5036 gnd.n5035 10.6151
R10611 gnd.n5035 gnd.n5032 10.6151
R10612 gnd.n5032 gnd.n5031 10.6151
R10613 gnd.n5031 gnd.n5029 10.6151
R10614 gnd.n5029 gnd.n5028 10.6151
R10615 gnd.n5028 gnd.n5026 10.6151
R10616 gnd.n5026 gnd.n3635 10.6151
R10617 gnd.n5119 gnd.n3635 10.6151
R10618 gnd.n5120 gnd.n5119 10.6151
R10619 gnd.n5127 gnd.n5120 10.6151
R10620 gnd.n5127 gnd.n5126 10.6151
R10621 gnd.n5126 gnd.n5125 10.6151
R10622 gnd.n5125 gnd.n5124 10.6151
R10623 gnd.n5124 gnd.n5122 10.6151
R10624 gnd.n5122 gnd.n5121 10.6151
R10625 gnd.n5121 gnd.n3610 10.6151
R10626 gnd.n5154 gnd.n3610 10.6151
R10627 gnd.n5155 gnd.n5154 10.6151
R10628 gnd.n5158 gnd.n5155 10.6151
R10629 gnd.n5159 gnd.n5158 10.6151
R10630 gnd.n5167 gnd.n5159 10.6151
R10631 gnd.n5167 gnd.n5166 10.6151
R10632 gnd.n5166 gnd.n5165 10.6151
R10633 gnd.n5165 gnd.n5164 10.6151
R10634 gnd.n5164 gnd.n5162 10.6151
R10635 gnd.n5162 gnd.n5161 10.6151
R10636 gnd.n5161 gnd.n3567 10.6151
R10637 gnd.n5241 gnd.n3567 10.6151
R10638 gnd.n5242 gnd.n5241 10.6151
R10639 gnd.n5249 gnd.n5242 10.6151
R10640 gnd.n5249 gnd.n5248 10.6151
R10641 gnd.n5248 gnd.n5247 10.6151
R10642 gnd.n5247 gnd.n5244 10.6151
R10643 gnd.n5244 gnd.n5243 10.6151
R10644 gnd.n5243 gnd.n3544 10.6151
R10645 gnd.n5277 gnd.n3544 10.6151
R10646 gnd.n5278 gnd.n5277 10.6151
R10647 gnd.n5279 gnd.n5278 10.6151
R10648 gnd.n3779 gnd.n2835 10.6151
R10649 gnd.n3782 gnd.n3779 10.6151
R10650 gnd.n3787 gnd.n3784 10.6151
R10651 gnd.n3788 gnd.n3787 10.6151
R10652 gnd.n3791 gnd.n3788 10.6151
R10653 gnd.n3792 gnd.n3791 10.6151
R10654 gnd.n3795 gnd.n3792 10.6151
R10655 gnd.n3796 gnd.n3795 10.6151
R10656 gnd.n3799 gnd.n3796 10.6151
R10657 gnd.n3800 gnd.n3799 10.6151
R10658 gnd.n3803 gnd.n3800 10.6151
R10659 gnd.n3804 gnd.n3803 10.6151
R10660 gnd.n3807 gnd.n3804 10.6151
R10661 gnd.n3808 gnd.n3807 10.6151
R10662 gnd.n3811 gnd.n3808 10.6151
R10663 gnd.n3812 gnd.n3811 10.6151
R10664 gnd.n3815 gnd.n3812 10.6151
R10665 gnd.n3816 gnd.n3815 10.6151
R10666 gnd.n3819 gnd.n3816 10.6151
R10667 gnd.n3820 gnd.n3819 10.6151
R10668 gnd.n3823 gnd.n3820 10.6151
R10669 gnd.n3824 gnd.n3823 10.6151
R10670 gnd.n3827 gnd.n3824 10.6151
R10671 gnd.n3828 gnd.n3827 10.6151
R10672 gnd.n3831 gnd.n3828 10.6151
R10673 gnd.n3832 gnd.n3831 10.6151
R10674 gnd.n3835 gnd.n3832 10.6151
R10675 gnd.n3836 gnd.n3835 10.6151
R10676 gnd.n3839 gnd.n3836 10.6151
R10677 gnd.n3840 gnd.n3839 10.6151
R10678 gnd.n6267 gnd.n6266 10.6151
R10679 gnd.n6266 gnd.n6265 10.6151
R10680 gnd.n6265 gnd.n6264 10.6151
R10681 gnd.n6264 gnd.n6262 10.6151
R10682 gnd.n6262 gnd.n6259 10.6151
R10683 gnd.n6259 gnd.n6258 10.6151
R10684 gnd.n6258 gnd.n6255 10.6151
R10685 gnd.n6255 gnd.n6254 10.6151
R10686 gnd.n6254 gnd.n6251 10.6151
R10687 gnd.n6251 gnd.n6250 10.6151
R10688 gnd.n6250 gnd.n6247 10.6151
R10689 gnd.n6247 gnd.n6246 10.6151
R10690 gnd.n6246 gnd.n6243 10.6151
R10691 gnd.n6243 gnd.n6242 10.6151
R10692 gnd.n6242 gnd.n6239 10.6151
R10693 gnd.n6239 gnd.n6238 10.6151
R10694 gnd.n6238 gnd.n6235 10.6151
R10695 gnd.n6235 gnd.n6234 10.6151
R10696 gnd.n6234 gnd.n6231 10.6151
R10697 gnd.n6231 gnd.n6230 10.6151
R10698 gnd.n6230 gnd.n6227 10.6151
R10699 gnd.n6227 gnd.n6226 10.6151
R10700 gnd.n6226 gnd.n6223 10.6151
R10701 gnd.n6223 gnd.n6222 10.6151
R10702 gnd.n6222 gnd.n6219 10.6151
R10703 gnd.n6219 gnd.n6218 10.6151
R10704 gnd.n6218 gnd.n6215 10.6151
R10705 gnd.n6215 gnd.n6214 10.6151
R10706 gnd.n6211 gnd.n6210 10.6151
R10707 gnd.n6210 gnd.n2836 10.6151
R10708 gnd.n5400 gnd.n3494 10.6151
R10709 gnd.n3495 gnd.n3494 10.6151
R10710 gnd.n5393 gnd.n3495 10.6151
R10711 gnd.n5393 gnd.n5392 10.6151
R10712 gnd.n5392 gnd.n5391 10.6151
R10713 gnd.n5391 gnd.n3497 10.6151
R10714 gnd.n5386 gnd.n3497 10.6151
R10715 gnd.n5386 gnd.n5385 10.6151
R10716 gnd.n5385 gnd.n5384 10.6151
R10717 gnd.n5384 gnd.n3500 10.6151
R10718 gnd.n5379 gnd.n3500 10.6151
R10719 gnd.n5379 gnd.n5378 10.6151
R10720 gnd.n5378 gnd.n5377 10.6151
R10721 gnd.n5377 gnd.n3503 10.6151
R10722 gnd.n5372 gnd.n3503 10.6151
R10723 gnd.n5372 gnd.n5371 10.6151
R10724 gnd.n5371 gnd.n5370 10.6151
R10725 gnd.n5370 gnd.n3506 10.6151
R10726 gnd.n5365 gnd.n3506 10.6151
R10727 gnd.n5365 gnd.n5364 10.6151
R10728 gnd.n5364 gnd.n5363 10.6151
R10729 gnd.n5363 gnd.n3509 10.6151
R10730 gnd.n5358 gnd.n3509 10.6151
R10731 gnd.n5358 gnd.n5357 10.6151
R10732 gnd.n5357 gnd.n5356 10.6151
R10733 gnd.n5356 gnd.n3512 10.6151
R10734 gnd.n5351 gnd.n3512 10.6151
R10735 gnd.n5351 gnd.n5350 10.6151
R10736 gnd.n5348 gnd.n3517 10.6151
R10737 gnd.n5343 gnd.n3517 10.6151
R10738 gnd.n6203 gnd.n6202 10.6151
R10739 gnd.n6202 gnd.n2894 10.6151
R10740 gnd.n4870 gnd.n2894 10.6151
R10741 gnd.n4870 gnd.n3773 10.6151
R10742 gnd.n4895 gnd.n3773 10.6151
R10743 gnd.n4896 gnd.n4895 10.6151
R10744 gnd.n4897 gnd.n4896 10.6151
R10745 gnd.n4897 gnd.n3756 10.6151
R10746 gnd.n4914 gnd.n3756 10.6151
R10747 gnd.n4915 gnd.n4914 10.6151
R10748 gnd.n4919 gnd.n4915 10.6151
R10749 gnd.n4919 gnd.n4918 10.6151
R10750 gnd.n4918 gnd.n4917 10.6151
R10751 gnd.n4917 gnd.n3731 10.6151
R10752 gnd.n4956 gnd.n3731 10.6151
R10753 gnd.n4957 gnd.n4956 10.6151
R10754 gnd.n4958 gnd.n4957 10.6151
R10755 gnd.n4958 gnd.n3717 10.6151
R10756 gnd.n4972 gnd.n3717 10.6151
R10757 gnd.n4973 gnd.n4972 10.6151
R10758 gnd.n4974 gnd.n4973 10.6151
R10759 gnd.n4974 gnd.n3706 10.6151
R10760 gnd.n4998 gnd.n3706 10.6151
R10761 gnd.n4998 gnd.n4997 10.6151
R10762 gnd.n4997 gnd.n4996 10.6151
R10763 gnd.n4996 gnd.n3707 10.6151
R10764 gnd.n3710 gnd.n3707 10.6151
R10765 gnd.n3710 gnd.n3709 10.6151
R10766 gnd.n3709 gnd.n3679 10.6151
R10767 gnd.n5043 gnd.n3679 10.6151
R10768 gnd.n5043 gnd.n5042 10.6151
R10769 gnd.n5042 gnd.n5041 10.6151
R10770 gnd.n5041 gnd.n3680 10.6151
R10771 gnd.n3680 gnd.n3657 10.6151
R10772 gnd.n5095 gnd.n3657 10.6151
R10773 gnd.n5096 gnd.n5095 10.6151
R10774 gnd.n5097 gnd.n5096 10.6151
R10775 gnd.n5097 gnd.n3642 10.6151
R10776 gnd.n5113 gnd.n3642 10.6151
R10777 gnd.n5114 gnd.n5113 10.6151
R10778 gnd.n5115 gnd.n5114 10.6151
R10779 gnd.n5115 gnd.n3630 10.6151
R10780 gnd.n5131 gnd.n3630 10.6151
R10781 gnd.n5132 gnd.n5131 10.6151
R10782 gnd.n5133 gnd.n5132 10.6151
R10783 gnd.n5133 gnd.n3614 10.6151
R10784 gnd.n5147 gnd.n3614 10.6151
R10785 gnd.n5148 gnd.n5147 10.6151
R10786 gnd.n5149 gnd.n5148 10.6151
R10787 gnd.n5149 gnd.n3606 10.6151
R10788 gnd.n5175 gnd.n3606 10.6151
R10789 gnd.n5175 gnd.n5174 10.6151
R10790 gnd.n5174 gnd.n5173 10.6151
R10791 gnd.n5173 gnd.n3607 10.6151
R10792 gnd.n3607 gnd.n3582 10.6151
R10793 gnd.n5222 gnd.n3582 10.6151
R10794 gnd.n5223 gnd.n5222 10.6151
R10795 gnd.n5227 gnd.n5223 10.6151
R10796 gnd.n5227 gnd.n5226 10.6151
R10797 gnd.n5226 gnd.n5225 10.6151
R10798 gnd.n5225 gnd.n3563 10.6151
R10799 gnd.n5254 gnd.n3563 10.6151
R10800 gnd.n5255 gnd.n5254 10.6151
R10801 gnd.n5256 gnd.n5255 10.6151
R10802 gnd.n5256 gnd.n3548 10.6151
R10803 gnd.n5270 gnd.n3548 10.6151
R10804 gnd.n5271 gnd.n5270 10.6151
R10805 gnd.n5272 gnd.n5271 10.6151
R10806 gnd.n5272 gnd.n3474 10.6151
R10807 gnd.n5403 gnd.n3474 10.6151
R10808 gnd.n5403 gnd.n5402 10.6151
R10809 gnd.n1695 gnd.t149 10.5161
R10810 gnd.n2031 gnd.t389 10.5161
R10811 gnd.t376 gnd.n976 10.5161
R10812 gnd.n4238 gnd.t151 10.5161
R10813 gnd.n4303 gnd.t58 10.5161
R10814 gnd.n4970 gnd.t88 10.5161
R10815 gnd.n5156 gnd.t338 10.5161
R10816 gnd.n5807 gnd.t20 10.5161
R10817 gnd.n5801 gnd.t162 10.5161
R10818 gnd.n2318 gnd.n2302 10.4732
R10819 gnd.n2286 gnd.n2270 10.4732
R10820 gnd.n2254 gnd.n2238 10.4732
R10821 gnd.n2223 gnd.n2207 10.4732
R10822 gnd.n2191 gnd.n2175 10.4732
R10823 gnd.n2159 gnd.n2143 10.4732
R10824 gnd.n2127 gnd.n2111 10.4732
R10825 gnd.n2096 gnd.n2080 10.4732
R10826 gnd.t285 gnd.n3771 10.1975
R10827 gnd.t241 gnd.n3751 10.1975
R10828 gnd.n5405 gnd.t235 10.1975
R10829 gnd.t136 gnd.n1131 9.87883
R10830 gnd.n6435 gnd.t111 9.87883
R10831 gnd.n6398 gnd.t108 9.87883
R10832 gnd.n5661 gnd.t0 9.87883
R10833 gnd.n7927 gnd.t80 9.87883
R10834 gnd.n2322 gnd.n2321 9.69747
R10835 gnd.n2290 gnd.n2289 9.69747
R10836 gnd.n2258 gnd.n2257 9.69747
R10837 gnd.n2227 gnd.n2226 9.69747
R10838 gnd.n2195 gnd.n2194 9.69747
R10839 gnd.n2163 gnd.n2162 9.69747
R10840 gnd.n2131 gnd.n2130 9.69747
R10841 gnd.n2100 gnd.n2099 9.69747
R10842 gnd.n3771 gnd.n3758 9.56018
R10843 gnd.n4930 gnd.n3744 9.56018
R10844 gnd.n4983 gnd.t15 9.56018
R10845 gnd.n5057 gnd.n3667 9.56018
R10846 gnd.n5063 gnd.n3655 9.56018
R10847 gnd.n5144 gnd.t312 9.56018
R10848 gnd.n5230 gnd.n5229 9.56018
R10849 gnd.n2328 gnd.n2327 9.45567
R10850 gnd.n2296 gnd.n2295 9.45567
R10851 gnd.n2264 gnd.n2263 9.45567
R10852 gnd.n2233 gnd.n2232 9.45567
R10853 gnd.n2201 gnd.n2200 9.45567
R10854 gnd.n2169 gnd.n2168 9.45567
R10855 gnd.n2137 gnd.n2136 9.45567
R10856 gnd.n2106 gnd.n2105 9.45567
R10857 gnd.n5954 gnd.n5953 9.30959
R10858 gnd.n7778 gnd.n331 9.30959
R10859 gnd.n6549 gnd.n6548 9.30959
R10860 gnd.n4704 gnd.n4701 9.30959
R10861 gnd.n2327 gnd.n2326 9.3005
R10862 gnd.n2300 gnd.n2299 9.3005
R10863 gnd.n2321 gnd.n2320 9.3005
R10864 gnd.n2319 gnd.n2318 9.3005
R10865 gnd.n2304 gnd.n2303 9.3005
R10866 gnd.n2313 gnd.n2312 9.3005
R10867 gnd.n2311 gnd.n2310 9.3005
R10868 gnd.n2295 gnd.n2294 9.3005
R10869 gnd.n2268 gnd.n2267 9.3005
R10870 gnd.n2289 gnd.n2288 9.3005
R10871 gnd.n2287 gnd.n2286 9.3005
R10872 gnd.n2272 gnd.n2271 9.3005
R10873 gnd.n2281 gnd.n2280 9.3005
R10874 gnd.n2279 gnd.n2278 9.3005
R10875 gnd.n2263 gnd.n2262 9.3005
R10876 gnd.n2236 gnd.n2235 9.3005
R10877 gnd.n2257 gnd.n2256 9.3005
R10878 gnd.n2255 gnd.n2254 9.3005
R10879 gnd.n2240 gnd.n2239 9.3005
R10880 gnd.n2249 gnd.n2248 9.3005
R10881 gnd.n2247 gnd.n2246 9.3005
R10882 gnd.n2232 gnd.n2231 9.3005
R10883 gnd.n2205 gnd.n2204 9.3005
R10884 gnd.n2226 gnd.n2225 9.3005
R10885 gnd.n2224 gnd.n2223 9.3005
R10886 gnd.n2209 gnd.n2208 9.3005
R10887 gnd.n2218 gnd.n2217 9.3005
R10888 gnd.n2216 gnd.n2215 9.3005
R10889 gnd.n2200 gnd.n2199 9.3005
R10890 gnd.n2173 gnd.n2172 9.3005
R10891 gnd.n2194 gnd.n2193 9.3005
R10892 gnd.n2192 gnd.n2191 9.3005
R10893 gnd.n2177 gnd.n2176 9.3005
R10894 gnd.n2186 gnd.n2185 9.3005
R10895 gnd.n2184 gnd.n2183 9.3005
R10896 gnd.n2168 gnd.n2167 9.3005
R10897 gnd.n2141 gnd.n2140 9.3005
R10898 gnd.n2162 gnd.n2161 9.3005
R10899 gnd.n2160 gnd.n2159 9.3005
R10900 gnd.n2145 gnd.n2144 9.3005
R10901 gnd.n2154 gnd.n2153 9.3005
R10902 gnd.n2152 gnd.n2151 9.3005
R10903 gnd.n2136 gnd.n2135 9.3005
R10904 gnd.n2109 gnd.n2108 9.3005
R10905 gnd.n2130 gnd.n2129 9.3005
R10906 gnd.n2128 gnd.n2127 9.3005
R10907 gnd.n2113 gnd.n2112 9.3005
R10908 gnd.n2122 gnd.n2121 9.3005
R10909 gnd.n2120 gnd.n2119 9.3005
R10910 gnd.n2105 gnd.n2104 9.3005
R10911 gnd.n2078 gnd.n2077 9.3005
R10912 gnd.n2099 gnd.n2098 9.3005
R10913 gnd.n2097 gnd.n2096 9.3005
R10914 gnd.n2082 gnd.n2081 9.3005
R10915 gnd.n2091 gnd.n2090 9.3005
R10916 gnd.n2089 gnd.n2088 9.3005
R10917 gnd.n6669 gnd.n6668 9.3005
R10918 gnd.n6667 gnd.n6635 9.3005
R10919 gnd.n6666 gnd.n6665 9.3005
R10920 gnd.n6662 gnd.n6636 9.3005
R10921 gnd.n6659 gnd.n6637 9.3005
R10922 gnd.n6658 gnd.n6638 9.3005
R10923 gnd.n6655 gnd.n6639 9.3005
R10924 gnd.n6654 gnd.n6640 9.3005
R10925 gnd.n6651 gnd.n6641 9.3005
R10926 gnd.n6650 gnd.n6642 9.3005
R10927 gnd.n6647 gnd.n6643 9.3005
R10928 gnd.n6646 gnd.n6644 9.3005
R10929 gnd.n1016 gnd.n1015 9.3005
R10930 gnd.n6677 gnd.n6676 9.3005
R10931 gnd.n6678 gnd.n1014 9.3005
R10932 gnd.n6680 gnd.n6679 9.3005
R10933 gnd.n6670 gnd.n6634 9.3005
R10934 gnd.n1714 gnd.n1713 9.3005
R10935 gnd.n1418 gnd.n1417 9.3005
R10936 gnd.n1741 gnd.n1740 9.3005
R10937 gnd.n1742 gnd.n1416 9.3005
R10938 gnd.n1746 gnd.n1743 9.3005
R10939 gnd.n1745 gnd.n1744 9.3005
R10940 gnd.n1390 gnd.n1389 9.3005
R10941 gnd.n1771 gnd.n1770 9.3005
R10942 gnd.n1772 gnd.n1388 9.3005
R10943 gnd.n1782 gnd.n1773 9.3005
R10944 gnd.n1781 gnd.n1774 9.3005
R10945 gnd.n1780 gnd.n1775 9.3005
R10946 gnd.n1778 gnd.n1777 9.3005
R10947 gnd.n1776 gnd.n1360 9.3005
R10948 gnd.n1358 gnd.n1357 9.3005
R10949 gnd.n1830 gnd.n1829 9.3005
R10950 gnd.n1831 gnd.n1356 9.3005
R10951 gnd.n1833 gnd.n1832 9.3005
R10952 gnd.n1227 gnd.n1226 9.3005
R10953 gnd.n1865 gnd.n1864 9.3005
R10954 gnd.n1866 gnd.n1225 9.3005
R10955 gnd.n1868 gnd.n1867 9.3005
R10956 gnd.n1206 gnd.n1205 9.3005
R10957 gnd.n1895 gnd.n1894 9.3005
R10958 gnd.n1896 gnd.n1204 9.3005
R10959 gnd.n1900 gnd.n1897 9.3005
R10960 gnd.n1899 gnd.n1898 9.3005
R10961 gnd.n1181 gnd.n1180 9.3005
R10962 gnd.n1944 gnd.n1943 9.3005
R10963 gnd.n1945 gnd.n1179 9.3005
R10964 gnd.n1949 gnd.n1946 9.3005
R10965 gnd.n1948 gnd.n1947 9.3005
R10966 gnd.n1154 gnd.n1153 9.3005
R10967 gnd.n1984 gnd.n1983 9.3005
R10968 gnd.n1985 gnd.n1152 9.3005
R10969 gnd.n1989 gnd.n1986 9.3005
R10970 gnd.n1988 gnd.n1987 9.3005
R10971 gnd.n1129 gnd.n1128 9.3005
R10972 gnd.n2045 gnd.n2044 9.3005
R10973 gnd.n2046 gnd.n1127 9.3005
R10974 gnd.n2054 gnd.n2047 9.3005
R10975 gnd.n2053 gnd.n2048 9.3005
R10976 gnd.n2052 gnd.n2050 9.3005
R10977 gnd.n2049 gnd.n970 9.3005
R10978 gnd.n6707 gnd.n971 9.3005
R10979 gnd.n6706 gnd.n972 9.3005
R10980 gnd.n6705 gnd.n973 9.3005
R10981 gnd.n994 gnd.n974 9.3005
R10982 gnd.n995 gnd.n993 9.3005
R10983 gnd.n6693 gnd.n996 9.3005
R10984 gnd.n6692 gnd.n997 9.3005
R10985 gnd.n6691 gnd.n998 9.3005
R10986 gnd.n6633 gnd.n999 9.3005
R10987 gnd.n1715 gnd.n1712 9.3005
R10988 gnd.n1497 gnd.n1456 9.3005
R10989 gnd.n1492 gnd.n1491 9.3005
R10990 gnd.n1490 gnd.n1457 9.3005
R10991 gnd.n1489 gnd.n1488 9.3005
R10992 gnd.n1485 gnd.n1458 9.3005
R10993 gnd.n1482 gnd.n1481 9.3005
R10994 gnd.n1480 gnd.n1459 9.3005
R10995 gnd.n1479 gnd.n1478 9.3005
R10996 gnd.n1475 gnd.n1460 9.3005
R10997 gnd.n1472 gnd.n1471 9.3005
R10998 gnd.n1470 gnd.n1461 9.3005
R10999 gnd.n1469 gnd.n1468 9.3005
R11000 gnd.n1465 gnd.n1463 9.3005
R11001 gnd.n1462 gnd.n1442 9.3005
R11002 gnd.n1709 gnd.n1441 9.3005
R11003 gnd.n1711 gnd.n1710 9.3005
R11004 gnd.n1499 gnd.n1498 9.3005
R11005 gnd.n1722 gnd.n1428 9.3005
R11006 gnd.n1729 gnd.n1429 9.3005
R11007 gnd.n1731 gnd.n1730 9.3005
R11008 gnd.n1732 gnd.n1409 9.3005
R11009 gnd.n1751 gnd.n1750 9.3005
R11010 gnd.n1753 gnd.n1401 9.3005
R11011 gnd.n1760 gnd.n1403 9.3005
R11012 gnd.n1761 gnd.n1398 9.3005
R11013 gnd.n1763 gnd.n1762 9.3005
R11014 gnd.n1399 gnd.n1384 9.3005
R11015 gnd.n1382 gnd.n1380 9.3005
R11016 gnd.n1789 gnd.n1788 9.3005
R11017 gnd.n1365 gnd.n1364 9.3005
R11018 gnd.n1822 gnd.n1810 9.3005
R11019 gnd.n1821 gnd.n1812 9.3005
R11020 gnd.n1820 gnd.n1813 9.3005
R11021 gnd.n1815 gnd.n1814 9.3005
R11022 gnd.n1348 gnd.n1236 9.3005
R11023 gnd.n1854 gnd.n1238 9.3005
R11024 gnd.n1855 gnd.n1234 9.3005
R11025 gnd.n1857 gnd.n1856 9.3005
R11026 gnd.n1222 gnd.n1217 9.3005
R11027 gnd.n1878 gnd.n1216 9.3005
R11028 gnd.n1881 gnd.n1880 9.3005
R11029 gnd.n1883 gnd.n1882 9.3005
R11030 gnd.n1886 gnd.n1199 9.3005
R11031 gnd.n1884 gnd.n1197 9.3005
R11032 gnd.n1907 gnd.n1195 9.3005
R11033 gnd.n1909 gnd.n1908 9.3005
R11034 gnd.n1172 gnd.n1171 9.3005
R11035 gnd.n1958 gnd.n1957 9.3005
R11036 gnd.n1959 gnd.n1165 9.3005
R11037 gnd.n1967 gnd.n1164 9.3005
R11038 gnd.n1970 gnd.n1969 9.3005
R11039 gnd.n1972 gnd.n1971 9.3005
R11040 gnd.n1975 gnd.n1148 9.3005
R11041 gnd.n1973 gnd.n1146 9.3005
R11042 gnd.n1995 gnd.n1144 9.3005
R11043 gnd.n1999 gnd.n1998 9.3005
R11044 gnd.n1997 gnd.n1120 9.3005
R11045 gnd.n2061 gnd.n1119 9.3005
R11046 gnd.n2064 gnd.n2063 9.3005
R11047 gnd.n1116 gnd.n1115 9.3005
R11048 gnd.n2068 gnd.n1117 9.3005
R11049 gnd.n2070 gnd.n2069 9.3005
R11050 gnd.n2072 gnd.n1114 9.3005
R11051 gnd.n2075 gnd.n2074 9.3005
R11052 gnd.n2333 gnd.n2332 9.3005
R11053 gnd.n2337 gnd.n2334 9.3005
R11054 gnd.n2339 gnd.n2338 9.3005
R11055 gnd.n2343 gnd.n2342 9.3005
R11056 gnd.n1010 gnd.n1008 9.3005
R11057 gnd.n6684 gnd.n6683 9.3005
R11058 gnd.n1720 gnd.n1719 9.3005
R11059 gnd.n1050 gnd.n1047 9.3005
R11060 gnd.n1052 gnd.n1051 9.3005
R11061 gnd.n1055 gnd.n1045 9.3005
R11062 gnd.n1059 gnd.n1058 9.3005
R11063 gnd.n1060 gnd.n1044 9.3005
R11064 gnd.n1062 gnd.n1061 9.3005
R11065 gnd.n1065 gnd.n1043 9.3005
R11066 gnd.n1069 gnd.n1068 9.3005
R11067 gnd.n1070 gnd.n1042 9.3005
R11068 gnd.n1072 gnd.n1071 9.3005
R11069 gnd.n1075 gnd.n1041 9.3005
R11070 gnd.n1079 gnd.n1078 9.3005
R11071 gnd.n1080 gnd.n1040 9.3005
R11072 gnd.n1082 gnd.n1081 9.3005
R11073 gnd.n1085 gnd.n1039 9.3005
R11074 gnd.n1089 gnd.n1088 9.3005
R11075 gnd.n1090 gnd.n1038 9.3005
R11076 gnd.n1092 gnd.n1091 9.3005
R11077 gnd.n1095 gnd.n1037 9.3005
R11078 gnd.n1099 gnd.n1098 9.3005
R11079 gnd.n1100 gnd.n1036 9.3005
R11080 gnd.n1102 gnd.n1101 9.3005
R11081 gnd.n1105 gnd.n1032 9.3005
R11082 gnd.n1108 gnd.n1107 9.3005
R11083 gnd.n1109 gnd.n1031 9.3005
R11084 gnd.n2353 gnd.n2352 9.3005
R11085 gnd.n1049 gnd.n1048 9.3005
R11086 gnd.n1249 gnd.n1245 9.3005
R11087 gnd.n1248 gnd.n1246 9.3005
R11088 gnd.n1188 gnd.n1187 9.3005
R11089 gnd.n1917 gnd.n1916 9.3005
R11090 gnd.n1918 gnd.n1186 9.3005
R11091 gnd.n1936 gnd.n1919 9.3005
R11092 gnd.n1935 gnd.n1920 9.3005
R11093 gnd.n1934 gnd.n1921 9.3005
R11094 gnd.n1932 gnd.n1922 9.3005
R11095 gnd.n1931 gnd.n1923 9.3005
R11096 gnd.n1929 gnd.n1924 9.3005
R11097 gnd.n1928 gnd.n1925 9.3005
R11098 gnd.n1136 gnd.n1135 9.3005
R11099 gnd.n2007 gnd.n2006 9.3005
R11100 gnd.n2008 gnd.n1134 9.3005
R11101 gnd.n2039 gnd.n2009 9.3005
R11102 gnd.n2038 gnd.n2010 9.3005
R11103 gnd.n2037 gnd.n2011 9.3005
R11104 gnd.n2034 gnd.n2012 9.3005
R11105 gnd.n2033 gnd.n2013 9.3005
R11106 gnd.n2030 gnd.n2014 9.3005
R11107 gnd.n2029 gnd.n2015 9.3005
R11108 gnd.n2026 gnd.n2016 9.3005
R11109 gnd.n2025 gnd.n2017 9.3005
R11110 gnd.n2024 gnd.n2018 9.3005
R11111 gnd.n2021 gnd.n2020 9.3005
R11112 gnd.n2019 gnd.n1111 9.3005
R11113 gnd.n2349 gnd.n1110 9.3005
R11114 gnd.n2351 gnd.n2350 9.3005
R11115 gnd.n1630 gnd.n1629 9.3005
R11116 gnd.n1520 gnd.n1519 9.3005
R11117 gnd.n1644 gnd.n1643 9.3005
R11118 gnd.n1645 gnd.n1518 9.3005
R11119 gnd.n1647 gnd.n1646 9.3005
R11120 gnd.n1508 gnd.n1507 9.3005
R11121 gnd.n1660 gnd.n1659 9.3005
R11122 gnd.n1661 gnd.n1506 9.3005
R11123 gnd.n1693 gnd.n1662 9.3005
R11124 gnd.n1692 gnd.n1663 9.3005
R11125 gnd.n1691 gnd.n1664 9.3005
R11126 gnd.n1690 gnd.n1665 9.3005
R11127 gnd.n1687 gnd.n1666 9.3005
R11128 gnd.n1686 gnd.n1667 9.3005
R11129 gnd.n1685 gnd.n1668 9.3005
R11130 gnd.n1683 gnd.n1669 9.3005
R11131 gnd.n1682 gnd.n1670 9.3005
R11132 gnd.n1679 gnd.n1671 9.3005
R11133 gnd.n1678 gnd.n1672 9.3005
R11134 gnd.n1677 gnd.n1673 9.3005
R11135 gnd.n1675 gnd.n1674 9.3005
R11136 gnd.n1373 gnd.n1372 9.3005
R11137 gnd.n1797 gnd.n1796 9.3005
R11138 gnd.n1798 gnd.n1371 9.3005
R11139 gnd.n1802 gnd.n1799 9.3005
R11140 gnd.n1801 gnd.n1800 9.3005
R11141 gnd.n1336 gnd.n1335 9.3005
R11142 gnd.n1845 gnd.n1844 9.3005
R11143 gnd.n1628 gnd.n1529 9.3005
R11144 gnd.n1531 gnd.n1530 9.3005
R11145 gnd.n1575 gnd.n1573 9.3005
R11146 gnd.n1576 gnd.n1572 9.3005
R11147 gnd.n1579 gnd.n1568 9.3005
R11148 gnd.n1580 gnd.n1567 9.3005
R11149 gnd.n1583 gnd.n1566 9.3005
R11150 gnd.n1584 gnd.n1565 9.3005
R11151 gnd.n1587 gnd.n1564 9.3005
R11152 gnd.n1588 gnd.n1563 9.3005
R11153 gnd.n1591 gnd.n1562 9.3005
R11154 gnd.n1592 gnd.n1561 9.3005
R11155 gnd.n1595 gnd.n1560 9.3005
R11156 gnd.n1596 gnd.n1559 9.3005
R11157 gnd.n1599 gnd.n1558 9.3005
R11158 gnd.n1600 gnd.n1557 9.3005
R11159 gnd.n1603 gnd.n1556 9.3005
R11160 gnd.n1604 gnd.n1555 9.3005
R11161 gnd.n1607 gnd.n1554 9.3005
R11162 gnd.n1608 gnd.n1553 9.3005
R11163 gnd.n1611 gnd.n1552 9.3005
R11164 gnd.n1612 gnd.n1551 9.3005
R11165 gnd.n1615 gnd.n1550 9.3005
R11166 gnd.n1617 gnd.n1549 9.3005
R11167 gnd.n1618 gnd.n1548 9.3005
R11168 gnd.n1619 gnd.n1547 9.3005
R11169 gnd.n1620 gnd.n1546 9.3005
R11170 gnd.n1627 gnd.n1626 9.3005
R11171 gnd.n1636 gnd.n1635 9.3005
R11172 gnd.n1637 gnd.n1523 9.3005
R11173 gnd.n1639 gnd.n1638 9.3005
R11174 gnd.n1514 gnd.n1513 9.3005
R11175 gnd.n1652 gnd.n1651 9.3005
R11176 gnd.n1653 gnd.n1512 9.3005
R11177 gnd.n1655 gnd.n1654 9.3005
R11178 gnd.n1501 gnd.n1500 9.3005
R11179 gnd.n1698 gnd.n1697 9.3005
R11180 gnd.n1699 gnd.n1455 9.3005
R11181 gnd.n1703 gnd.n1701 9.3005
R11182 gnd.n1702 gnd.n1434 9.3005
R11183 gnd.n1721 gnd.n1433 9.3005
R11184 gnd.n1724 gnd.n1723 9.3005
R11185 gnd.n1427 gnd.n1426 9.3005
R11186 gnd.n1735 gnd.n1733 9.3005
R11187 gnd.n1734 gnd.n1408 9.3005
R11188 gnd.n1752 gnd.n1407 9.3005
R11189 gnd.n1755 gnd.n1754 9.3005
R11190 gnd.n1402 gnd.n1397 9.3005
R11191 gnd.n1765 gnd.n1764 9.3005
R11192 gnd.n1400 gnd.n1378 9.3005
R11193 gnd.n1792 gnd.n1379 9.3005
R11194 gnd.n1791 gnd.n1790 9.3005
R11195 gnd.n1381 gnd.n1366 9.3005
R11196 gnd.n1809 gnd.n1808 9.3005
R11197 gnd.n1811 gnd.n1344 9.3005
R11198 gnd.n1840 gnd.n1345 9.3005
R11199 gnd.n1839 gnd.n1346 9.3005
R11200 gnd.n1838 gnd.n1347 9.3005
R11201 gnd.n1350 gnd.n1349 9.3005
R11202 gnd.n1237 gnd.n1233 9.3005
R11203 gnd.n1859 gnd.n1858 9.3005
R11204 gnd.n1235 gnd.n1218 9.3005
R11205 gnd.n1877 gnd.n1876 9.3005
R11206 gnd.n1879 gnd.n1214 9.3005
R11207 gnd.n1889 gnd.n1215 9.3005
R11208 gnd.n1888 gnd.n1887 9.3005
R11209 gnd.n1885 gnd.n1193 9.3005
R11210 gnd.n1912 gnd.n1194 9.3005
R11211 gnd.n1911 gnd.n1910 9.3005
R11212 gnd.n1196 gnd.n1173 9.3005
R11213 gnd.n1955 gnd.n1954 9.3005
R11214 gnd.n1956 gnd.n1166 9.3005
R11215 gnd.n1966 gnd.n1965 9.3005
R11216 gnd.n1968 gnd.n1162 9.3005
R11217 gnd.n1978 gnd.n1163 9.3005
R11218 gnd.n1977 gnd.n1976 9.3005
R11219 gnd.n1974 gnd.n1142 9.3005
R11220 gnd.n2002 gnd.n1143 9.3005
R11221 gnd.n2001 gnd.n2000 9.3005
R11222 gnd.n1145 gnd.n1121 9.3005
R11223 gnd.n2060 gnd.n2059 9.3005
R11224 gnd.n2062 gnd.n958 9.3005
R11225 gnd.n6714 gnd.n959 9.3005
R11226 gnd.n6713 gnd.n960 9.3005
R11227 gnd.n6712 gnd.n961 9.3005
R11228 gnd.n2071 gnd.n962 9.3005
R11229 gnd.n2073 gnd.n982 9.3005
R11230 gnd.n6700 gnd.n983 9.3005
R11231 gnd.n6699 gnd.n984 9.3005
R11232 gnd.n6698 gnd.n985 9.3005
R11233 gnd.n2340 gnd.n986 9.3005
R11234 gnd.n2341 gnd.n1007 9.3005
R11235 gnd.n6686 gnd.n6685 9.3005
R11236 gnd.n1525 gnd.n1524 9.3005
R11237 gnd.n784 gnd.n783 9.3005
R11238 gnd.n6890 gnd.n6889 9.3005
R11239 gnd.n6891 gnd.n782 9.3005
R11240 gnd.n6893 gnd.n6892 9.3005
R11241 gnd.n778 gnd.n777 9.3005
R11242 gnd.n6900 gnd.n6899 9.3005
R11243 gnd.n6901 gnd.n776 9.3005
R11244 gnd.n6903 gnd.n6902 9.3005
R11245 gnd.n772 gnd.n771 9.3005
R11246 gnd.n6910 gnd.n6909 9.3005
R11247 gnd.n6911 gnd.n770 9.3005
R11248 gnd.n6913 gnd.n6912 9.3005
R11249 gnd.n766 gnd.n765 9.3005
R11250 gnd.n6920 gnd.n6919 9.3005
R11251 gnd.n6921 gnd.n764 9.3005
R11252 gnd.n6923 gnd.n6922 9.3005
R11253 gnd.n760 gnd.n759 9.3005
R11254 gnd.n6930 gnd.n6929 9.3005
R11255 gnd.n6931 gnd.n758 9.3005
R11256 gnd.n6933 gnd.n6932 9.3005
R11257 gnd.n754 gnd.n753 9.3005
R11258 gnd.n6940 gnd.n6939 9.3005
R11259 gnd.n6941 gnd.n752 9.3005
R11260 gnd.n6943 gnd.n6942 9.3005
R11261 gnd.n748 gnd.n747 9.3005
R11262 gnd.n6950 gnd.n6949 9.3005
R11263 gnd.n6951 gnd.n746 9.3005
R11264 gnd.n6953 gnd.n6952 9.3005
R11265 gnd.n742 gnd.n741 9.3005
R11266 gnd.n6960 gnd.n6959 9.3005
R11267 gnd.n6961 gnd.n740 9.3005
R11268 gnd.n6963 gnd.n6962 9.3005
R11269 gnd.n736 gnd.n735 9.3005
R11270 gnd.n6970 gnd.n6969 9.3005
R11271 gnd.n6971 gnd.n734 9.3005
R11272 gnd.n6973 gnd.n6972 9.3005
R11273 gnd.n730 gnd.n729 9.3005
R11274 gnd.n6980 gnd.n6979 9.3005
R11275 gnd.n6981 gnd.n728 9.3005
R11276 gnd.n6983 gnd.n6982 9.3005
R11277 gnd.n724 gnd.n723 9.3005
R11278 gnd.n6990 gnd.n6989 9.3005
R11279 gnd.n6991 gnd.n722 9.3005
R11280 gnd.n6993 gnd.n6992 9.3005
R11281 gnd.n718 gnd.n717 9.3005
R11282 gnd.n7000 gnd.n6999 9.3005
R11283 gnd.n7001 gnd.n716 9.3005
R11284 gnd.n7003 gnd.n7002 9.3005
R11285 gnd.n712 gnd.n711 9.3005
R11286 gnd.n7010 gnd.n7009 9.3005
R11287 gnd.n7011 gnd.n710 9.3005
R11288 gnd.n7013 gnd.n7012 9.3005
R11289 gnd.n706 gnd.n705 9.3005
R11290 gnd.n7020 gnd.n7019 9.3005
R11291 gnd.n7021 gnd.n704 9.3005
R11292 gnd.n7023 gnd.n7022 9.3005
R11293 gnd.n700 gnd.n699 9.3005
R11294 gnd.n7030 gnd.n7029 9.3005
R11295 gnd.n7031 gnd.n698 9.3005
R11296 gnd.n7033 gnd.n7032 9.3005
R11297 gnd.n694 gnd.n693 9.3005
R11298 gnd.n7040 gnd.n7039 9.3005
R11299 gnd.n7041 gnd.n692 9.3005
R11300 gnd.n7043 gnd.n7042 9.3005
R11301 gnd.n688 gnd.n687 9.3005
R11302 gnd.n7050 gnd.n7049 9.3005
R11303 gnd.n7051 gnd.n686 9.3005
R11304 gnd.n7053 gnd.n7052 9.3005
R11305 gnd.n682 gnd.n681 9.3005
R11306 gnd.n7060 gnd.n7059 9.3005
R11307 gnd.n7061 gnd.n680 9.3005
R11308 gnd.n7063 gnd.n7062 9.3005
R11309 gnd.n676 gnd.n675 9.3005
R11310 gnd.n7070 gnd.n7069 9.3005
R11311 gnd.n7071 gnd.n674 9.3005
R11312 gnd.n7073 gnd.n7072 9.3005
R11313 gnd.n670 gnd.n669 9.3005
R11314 gnd.n7080 gnd.n7079 9.3005
R11315 gnd.n7081 gnd.n668 9.3005
R11316 gnd.n7083 gnd.n7082 9.3005
R11317 gnd.n664 gnd.n663 9.3005
R11318 gnd.n7090 gnd.n7089 9.3005
R11319 gnd.n7091 gnd.n662 9.3005
R11320 gnd.n7093 gnd.n7092 9.3005
R11321 gnd.n658 gnd.n657 9.3005
R11322 gnd.n7100 gnd.n7099 9.3005
R11323 gnd.n7101 gnd.n656 9.3005
R11324 gnd.n7103 gnd.n7102 9.3005
R11325 gnd.n652 gnd.n651 9.3005
R11326 gnd.n7110 gnd.n7109 9.3005
R11327 gnd.n7111 gnd.n650 9.3005
R11328 gnd.n7113 gnd.n7112 9.3005
R11329 gnd.n646 gnd.n645 9.3005
R11330 gnd.n7120 gnd.n7119 9.3005
R11331 gnd.n7121 gnd.n644 9.3005
R11332 gnd.n7123 gnd.n7122 9.3005
R11333 gnd.n640 gnd.n639 9.3005
R11334 gnd.n7130 gnd.n7129 9.3005
R11335 gnd.n7131 gnd.n638 9.3005
R11336 gnd.n7133 gnd.n7132 9.3005
R11337 gnd.n634 gnd.n633 9.3005
R11338 gnd.n7140 gnd.n7139 9.3005
R11339 gnd.n7141 gnd.n632 9.3005
R11340 gnd.n7143 gnd.n7142 9.3005
R11341 gnd.n628 gnd.n627 9.3005
R11342 gnd.n7150 gnd.n7149 9.3005
R11343 gnd.n7151 gnd.n626 9.3005
R11344 gnd.n7153 gnd.n7152 9.3005
R11345 gnd.n622 gnd.n621 9.3005
R11346 gnd.n7160 gnd.n7159 9.3005
R11347 gnd.n7161 gnd.n620 9.3005
R11348 gnd.n7163 gnd.n7162 9.3005
R11349 gnd.n616 gnd.n615 9.3005
R11350 gnd.n7170 gnd.n7169 9.3005
R11351 gnd.n7171 gnd.n614 9.3005
R11352 gnd.n7173 gnd.n7172 9.3005
R11353 gnd.n610 gnd.n609 9.3005
R11354 gnd.n7180 gnd.n7179 9.3005
R11355 gnd.n7181 gnd.n608 9.3005
R11356 gnd.n7183 gnd.n7182 9.3005
R11357 gnd.n604 gnd.n603 9.3005
R11358 gnd.n7190 gnd.n7189 9.3005
R11359 gnd.n7191 gnd.n602 9.3005
R11360 gnd.n7193 gnd.n7192 9.3005
R11361 gnd.n598 gnd.n597 9.3005
R11362 gnd.n7200 gnd.n7199 9.3005
R11363 gnd.n7201 gnd.n596 9.3005
R11364 gnd.n7203 gnd.n7202 9.3005
R11365 gnd.n592 gnd.n591 9.3005
R11366 gnd.n7210 gnd.n7209 9.3005
R11367 gnd.n7211 gnd.n590 9.3005
R11368 gnd.n7213 gnd.n7212 9.3005
R11369 gnd.n586 gnd.n585 9.3005
R11370 gnd.n7220 gnd.n7219 9.3005
R11371 gnd.n7221 gnd.n584 9.3005
R11372 gnd.n7223 gnd.n7222 9.3005
R11373 gnd.n580 gnd.n579 9.3005
R11374 gnd.n7230 gnd.n7229 9.3005
R11375 gnd.n7231 gnd.n578 9.3005
R11376 gnd.n7233 gnd.n7232 9.3005
R11377 gnd.n574 gnd.n573 9.3005
R11378 gnd.n7240 gnd.n7239 9.3005
R11379 gnd.n7241 gnd.n572 9.3005
R11380 gnd.n7243 gnd.n7242 9.3005
R11381 gnd.n568 gnd.n567 9.3005
R11382 gnd.n7250 gnd.n7249 9.3005
R11383 gnd.n7251 gnd.n566 9.3005
R11384 gnd.n7253 gnd.n7252 9.3005
R11385 gnd.n562 gnd.n561 9.3005
R11386 gnd.n7260 gnd.n7259 9.3005
R11387 gnd.n7261 gnd.n560 9.3005
R11388 gnd.n7263 gnd.n7262 9.3005
R11389 gnd.n556 gnd.n555 9.3005
R11390 gnd.n7270 gnd.n7269 9.3005
R11391 gnd.n7271 gnd.n554 9.3005
R11392 gnd.n7273 gnd.n7272 9.3005
R11393 gnd.n550 gnd.n549 9.3005
R11394 gnd.n7280 gnd.n7279 9.3005
R11395 gnd.n7281 gnd.n548 9.3005
R11396 gnd.n7283 gnd.n7282 9.3005
R11397 gnd.n544 gnd.n543 9.3005
R11398 gnd.n7290 gnd.n7289 9.3005
R11399 gnd.n7291 gnd.n542 9.3005
R11400 gnd.n7293 gnd.n7292 9.3005
R11401 gnd.n538 gnd.n537 9.3005
R11402 gnd.n7300 gnd.n7299 9.3005
R11403 gnd.n7301 gnd.n536 9.3005
R11404 gnd.n7303 gnd.n7302 9.3005
R11405 gnd.n532 gnd.n531 9.3005
R11406 gnd.n7310 gnd.n7309 9.3005
R11407 gnd.n7311 gnd.n530 9.3005
R11408 gnd.n7313 gnd.n7312 9.3005
R11409 gnd.n526 gnd.n525 9.3005
R11410 gnd.n7320 gnd.n7319 9.3005
R11411 gnd.n7321 gnd.n524 9.3005
R11412 gnd.n7323 gnd.n7322 9.3005
R11413 gnd.n520 gnd.n519 9.3005
R11414 gnd.n7330 gnd.n7329 9.3005
R11415 gnd.n7331 gnd.n518 9.3005
R11416 gnd.n7333 gnd.n7332 9.3005
R11417 gnd.n514 gnd.n513 9.3005
R11418 gnd.n7340 gnd.n7339 9.3005
R11419 gnd.n7341 gnd.n512 9.3005
R11420 gnd.n7343 gnd.n7342 9.3005
R11421 gnd.n508 gnd.n507 9.3005
R11422 gnd.n7350 gnd.n7349 9.3005
R11423 gnd.n7351 gnd.n506 9.3005
R11424 gnd.n7353 gnd.n7352 9.3005
R11425 gnd.n502 gnd.n501 9.3005
R11426 gnd.n7360 gnd.n7359 9.3005
R11427 gnd.n7361 gnd.n500 9.3005
R11428 gnd.n7364 gnd.n7363 9.3005
R11429 gnd.n7362 gnd.n496 9.3005
R11430 gnd.n7370 gnd.n495 9.3005
R11431 gnd.n7372 gnd.n7371 9.3005
R11432 gnd.n491 gnd.n490 9.3005
R11433 gnd.n7381 gnd.n7380 9.3005
R11434 gnd.n7382 gnd.n489 9.3005
R11435 gnd.n7384 gnd.n7383 9.3005
R11436 gnd.n485 gnd.n484 9.3005
R11437 gnd.n7391 gnd.n7390 9.3005
R11438 gnd.n7392 gnd.n483 9.3005
R11439 gnd.n7394 gnd.n7393 9.3005
R11440 gnd.n479 gnd.n478 9.3005
R11441 gnd.n7401 gnd.n7400 9.3005
R11442 gnd.n7402 gnd.n477 9.3005
R11443 gnd.n7404 gnd.n7403 9.3005
R11444 gnd.n473 gnd.n472 9.3005
R11445 gnd.n7411 gnd.n7410 9.3005
R11446 gnd.n7412 gnd.n471 9.3005
R11447 gnd.n7414 gnd.n7413 9.3005
R11448 gnd.n467 gnd.n466 9.3005
R11449 gnd.n7421 gnd.n7420 9.3005
R11450 gnd.n7422 gnd.n465 9.3005
R11451 gnd.n7424 gnd.n7423 9.3005
R11452 gnd.n461 gnd.n460 9.3005
R11453 gnd.n7431 gnd.n7430 9.3005
R11454 gnd.n7432 gnd.n459 9.3005
R11455 gnd.n7434 gnd.n7433 9.3005
R11456 gnd.n455 gnd.n454 9.3005
R11457 gnd.n7441 gnd.n7440 9.3005
R11458 gnd.n7442 gnd.n453 9.3005
R11459 gnd.n7444 gnd.n7443 9.3005
R11460 gnd.n449 gnd.n448 9.3005
R11461 gnd.n7451 gnd.n7450 9.3005
R11462 gnd.n7452 gnd.n447 9.3005
R11463 gnd.n7454 gnd.n7453 9.3005
R11464 gnd.n443 gnd.n442 9.3005
R11465 gnd.n7461 gnd.n7460 9.3005
R11466 gnd.n7462 gnd.n441 9.3005
R11467 gnd.n7464 gnd.n7463 9.3005
R11468 gnd.n437 gnd.n436 9.3005
R11469 gnd.n7471 gnd.n7470 9.3005
R11470 gnd.n7472 gnd.n435 9.3005
R11471 gnd.n7474 gnd.n7473 9.3005
R11472 gnd.n431 gnd.n430 9.3005
R11473 gnd.n7481 gnd.n7480 9.3005
R11474 gnd.n7482 gnd.n429 9.3005
R11475 gnd.n7484 gnd.n7483 9.3005
R11476 gnd.n425 gnd.n424 9.3005
R11477 gnd.n7491 gnd.n7490 9.3005
R11478 gnd.n7492 gnd.n423 9.3005
R11479 gnd.n7494 gnd.n7493 9.3005
R11480 gnd.n419 gnd.n418 9.3005
R11481 gnd.n7501 gnd.n7500 9.3005
R11482 gnd.n7502 gnd.n417 9.3005
R11483 gnd.n7504 gnd.n7503 9.3005
R11484 gnd.n413 gnd.n412 9.3005
R11485 gnd.n7511 gnd.n7510 9.3005
R11486 gnd.n7512 gnd.n411 9.3005
R11487 gnd.n7514 gnd.n7513 9.3005
R11488 gnd.n407 gnd.n406 9.3005
R11489 gnd.n7521 gnd.n7520 9.3005
R11490 gnd.n7522 gnd.n405 9.3005
R11491 gnd.n7524 gnd.n7523 9.3005
R11492 gnd.n401 gnd.n400 9.3005
R11493 gnd.n7531 gnd.n7530 9.3005
R11494 gnd.n7532 gnd.n399 9.3005
R11495 gnd.n7534 gnd.n7533 9.3005
R11496 gnd.n395 gnd.n394 9.3005
R11497 gnd.n7541 gnd.n7540 9.3005
R11498 gnd.n7542 gnd.n393 9.3005
R11499 gnd.n7544 gnd.n7543 9.3005
R11500 gnd.n389 gnd.n388 9.3005
R11501 gnd.n7551 gnd.n7550 9.3005
R11502 gnd.n7552 gnd.n387 9.3005
R11503 gnd.n7554 gnd.n7553 9.3005
R11504 gnd.n383 gnd.n382 9.3005
R11505 gnd.n7561 gnd.n7560 9.3005
R11506 gnd.n7562 gnd.n381 9.3005
R11507 gnd.n7564 gnd.n7563 9.3005
R11508 gnd.n377 gnd.n376 9.3005
R11509 gnd.n7571 gnd.n7570 9.3005
R11510 gnd.n7572 gnd.n375 9.3005
R11511 gnd.n7574 gnd.n7573 9.3005
R11512 gnd.n371 gnd.n370 9.3005
R11513 gnd.n7582 gnd.n7581 9.3005
R11514 gnd.n7583 gnd.n369 9.3005
R11515 gnd.n7586 gnd.n7585 9.3005
R11516 gnd.n7374 gnd.n7373 9.3005
R11517 gnd.n7951 gnd.n7950 9.3005
R11518 gnd.n7949 gnd.n97 9.3005
R11519 gnd.n5721 gnd.n99 9.3005
R11520 gnd.n5725 gnd.n5724 9.3005
R11521 gnd.n5726 gnd.n5720 9.3005
R11522 gnd.n5781 gnd.n5727 9.3005
R11523 gnd.n5780 gnd.n5728 9.3005
R11524 gnd.n5779 gnd.n5729 9.3005
R11525 gnd.n5756 gnd.n5730 9.3005
R11526 gnd.n5769 gnd.n5757 9.3005
R11527 gnd.n5768 gnd.n5758 9.3005
R11528 gnd.n5767 gnd.n5759 9.3005
R11529 gnd.n359 gnd.n358 9.3005
R11530 gnd.n7599 gnd.n7598 9.3005
R11531 gnd.n7600 gnd.n357 9.3005
R11532 gnd.n7699 gnd.n7601 9.3005
R11533 gnd.n7698 gnd.n7602 9.3005
R11534 gnd.n7697 gnd.n7603 9.3005
R11535 gnd.n7695 gnd.n7604 9.3005
R11536 gnd.n7694 gnd.n7605 9.3005
R11537 gnd.n7692 gnd.n7606 9.3005
R11538 gnd.n7691 gnd.n7607 9.3005
R11539 gnd.n7689 gnd.n7608 9.3005
R11540 gnd.n7688 gnd.n7609 9.3005
R11541 gnd.n7686 gnd.n7610 9.3005
R11542 gnd.n7685 gnd.n7611 9.3005
R11543 gnd.n7683 gnd.n7612 9.3005
R11544 gnd.n7682 gnd.n7613 9.3005
R11545 gnd.n7680 gnd.n7614 9.3005
R11546 gnd.n7679 gnd.n7615 9.3005
R11547 gnd.n7677 gnd.n7616 9.3005
R11548 gnd.n7676 gnd.n7617 9.3005
R11549 gnd.n7631 gnd.n7630 9.3005
R11550 gnd.n7633 gnd.n7632 9.3005
R11551 gnd.n7636 gnd.n7627 9.3005
R11552 gnd.n7640 gnd.n7639 9.3005
R11553 gnd.n7641 gnd.n7626 9.3005
R11554 gnd.n7643 gnd.n7642 9.3005
R11555 gnd.n7646 gnd.n7625 9.3005
R11556 gnd.n7650 gnd.n7649 9.3005
R11557 gnd.n7651 gnd.n7624 9.3005
R11558 gnd.n7653 gnd.n7652 9.3005
R11559 gnd.n7656 gnd.n7623 9.3005
R11560 gnd.n7660 gnd.n7659 9.3005
R11561 gnd.n7661 gnd.n7622 9.3005
R11562 gnd.n7663 gnd.n7662 9.3005
R11563 gnd.n7666 gnd.n7621 9.3005
R11564 gnd.n7670 gnd.n7669 9.3005
R11565 gnd.n7671 gnd.n7620 9.3005
R11566 gnd.n7673 gnd.n7672 9.3005
R11567 gnd.n7628 gnd.n354 9.3005
R11568 gnd.n254 gnd.n253 9.3005
R11569 gnd.n7850 gnd.n296 9.3005
R11570 gnd.n7849 gnd.n297 9.3005
R11571 gnd.n7848 gnd.n298 9.3005
R11572 gnd.n7845 gnd.n299 9.3005
R11573 gnd.n7844 gnd.n300 9.3005
R11574 gnd.n7841 gnd.n301 9.3005
R11575 gnd.n7840 gnd.n302 9.3005
R11576 gnd.n7837 gnd.n303 9.3005
R11577 gnd.n7836 gnd.n304 9.3005
R11578 gnd.n7833 gnd.n305 9.3005
R11579 gnd.n7832 gnd.n306 9.3005
R11580 gnd.n7829 gnd.n307 9.3005
R11581 gnd.n7828 gnd.n308 9.3005
R11582 gnd.n7825 gnd.n309 9.3005
R11583 gnd.n7824 gnd.n310 9.3005
R11584 gnd.n7821 gnd.n311 9.3005
R11585 gnd.n7817 gnd.n312 9.3005
R11586 gnd.n7814 gnd.n313 9.3005
R11587 gnd.n7813 gnd.n314 9.3005
R11588 gnd.n7810 gnd.n315 9.3005
R11589 gnd.n7809 gnd.n316 9.3005
R11590 gnd.n7806 gnd.n317 9.3005
R11591 gnd.n7805 gnd.n318 9.3005
R11592 gnd.n7802 gnd.n319 9.3005
R11593 gnd.n7801 gnd.n320 9.3005
R11594 gnd.n7798 gnd.n321 9.3005
R11595 gnd.n7797 gnd.n322 9.3005
R11596 gnd.n7794 gnd.n323 9.3005
R11597 gnd.n7793 gnd.n324 9.3005
R11598 gnd.n7790 gnd.n325 9.3005
R11599 gnd.n7789 gnd.n326 9.3005
R11600 gnd.n7786 gnd.n327 9.3005
R11601 gnd.n7785 gnd.n328 9.3005
R11602 gnd.n7782 gnd.n329 9.3005
R11603 gnd.n7781 gnd.n330 9.3005
R11604 gnd.n7778 gnd.n7777 9.3005
R11605 gnd.n7776 gnd.n331 9.3005
R11606 gnd.n7775 gnd.n7774 9.3005
R11607 gnd.n7771 gnd.n334 9.3005
R11608 gnd.n7768 gnd.n335 9.3005
R11609 gnd.n7767 gnd.n336 9.3005
R11610 gnd.n7764 gnd.n337 9.3005
R11611 gnd.n7763 gnd.n338 9.3005
R11612 gnd.n7760 gnd.n339 9.3005
R11613 gnd.n7759 gnd.n340 9.3005
R11614 gnd.n7756 gnd.n341 9.3005
R11615 gnd.n7755 gnd.n342 9.3005
R11616 gnd.n7752 gnd.n343 9.3005
R11617 gnd.n7751 gnd.n344 9.3005
R11618 gnd.n7748 gnd.n345 9.3005
R11619 gnd.n7747 gnd.n346 9.3005
R11620 gnd.n7744 gnd.n347 9.3005
R11621 gnd.n7743 gnd.n348 9.3005
R11622 gnd.n7740 gnd.n349 9.3005
R11623 gnd.n7739 gnd.n350 9.3005
R11624 gnd.n7736 gnd.n7735 9.3005
R11625 gnd.n7734 gnd.n351 9.3005
R11626 gnd.n7856 gnd.n7855 9.3005
R11627 gnd.n5903 gnd.n5902 9.3005
R11628 gnd.n3180 gnd.n3179 9.3005
R11629 gnd.n3204 gnd.n3203 9.3005
R11630 gnd.n5890 gnd.n3205 9.3005
R11631 gnd.n5889 gnd.n3206 9.3005
R11632 gnd.n5888 gnd.n3207 9.3005
R11633 gnd.n5598 gnd.n3208 9.3005
R11634 gnd.n5878 gnd.n3226 9.3005
R11635 gnd.n5877 gnd.n3227 9.3005
R11636 gnd.n5876 gnd.n3228 9.3005
R11637 gnd.n5613 gnd.n3229 9.3005
R11638 gnd.n5866 gnd.n3246 9.3005
R11639 gnd.n5865 gnd.n3247 9.3005
R11640 gnd.n5864 gnd.n3248 9.3005
R11641 gnd.n5628 gnd.n3249 9.3005
R11642 gnd.n5854 gnd.n3267 9.3005
R11643 gnd.n5853 gnd.n3268 9.3005
R11644 gnd.n5852 gnd.n3269 9.3005
R11645 gnd.n5643 gnd.n3270 9.3005
R11646 gnd.n5842 gnd.n3287 9.3005
R11647 gnd.n5841 gnd.n3288 9.3005
R11648 gnd.n5840 gnd.n3289 9.3005
R11649 gnd.n5658 gnd.n3290 9.3005
R11650 gnd.n5830 gnd.n3309 9.3005
R11651 gnd.n5829 gnd.n3310 9.3005
R11652 gnd.n5828 gnd.n3311 9.3005
R11653 gnd.n3353 gnd.n3312 9.3005
R11654 gnd.n5690 gnd.n5689 9.3005
R11655 gnd.n5694 gnd.n5693 9.3005
R11656 gnd.n5695 gnd.n3343 9.3005
R11657 gnd.n5805 gnd.n3344 9.3005
R11658 gnd.n5804 gnd.n3345 9.3005
R11659 gnd.n5803 gnd.n3346 9.3005
R11660 gnd.n5699 gnd.n3347 9.3005
R11661 gnd.n5793 gnd.n5700 9.3005
R11662 gnd.n5701 gnd.n124 9.3005
R11663 gnd.n7937 gnd.n125 9.3005
R11664 gnd.n7936 gnd.n126 9.3005
R11665 gnd.n7935 gnd.n127 9.3005
R11666 gnd.n5734 gnd.n128 9.3005
R11667 gnd.n7925 gnd.n143 9.3005
R11668 gnd.n7924 gnd.n144 9.3005
R11669 gnd.n7923 gnd.n145 9.3005
R11670 gnd.n5760 gnd.n146 9.3005
R11671 gnd.n7913 gnd.n164 9.3005
R11672 gnd.n7912 gnd.n165 9.3005
R11673 gnd.n7911 gnd.n166 9.3005
R11674 gnd.n356 gnd.n167 9.3005
R11675 gnd.n7901 gnd.n183 9.3005
R11676 gnd.n7900 gnd.n184 9.3005
R11677 gnd.n7899 gnd.n185 9.3005
R11678 gnd.n7708 gnd.n186 9.3005
R11679 gnd.n7889 gnd.n204 9.3005
R11680 gnd.n7888 gnd.n205 9.3005
R11681 gnd.n7887 gnd.n206 9.3005
R11682 gnd.n7715 gnd.n207 9.3005
R11683 gnd.n7877 gnd.n222 9.3005
R11684 gnd.n7876 gnd.n223 9.3005
R11685 gnd.n7875 gnd.n224 9.3005
R11686 gnd.n7722 gnd.n225 9.3005
R11687 gnd.n7865 gnd.n242 9.3005
R11688 gnd.n7864 gnd.n243 9.3005
R11689 gnd.n7863 gnd.n244 9.3005
R11690 gnd.n7732 gnd.n245 9.3005
R11691 gnd.n5904 gnd.n3178 9.3005
R11692 gnd.n5902 gnd.n5901 9.3005
R11693 gnd.n5900 gnd.n3180 9.3005
R11694 gnd.n3204 gnd.n3181 9.3005
R11695 gnd.n3377 gnd.n3205 9.3005
R11696 gnd.n5596 gnd.n3206 9.3005
R11697 gnd.n5597 gnd.n3207 9.3005
R11698 gnd.n5599 gnd.n5598 9.3005
R11699 gnd.n3373 gnd.n3226 9.3005
R11700 gnd.n5611 gnd.n3227 9.3005
R11701 gnd.n5612 gnd.n3228 9.3005
R11702 gnd.n5614 gnd.n5613 9.3005
R11703 gnd.n3368 gnd.n3246 9.3005
R11704 gnd.n5626 gnd.n3247 9.3005
R11705 gnd.n5627 gnd.n3248 9.3005
R11706 gnd.n5629 gnd.n5628 9.3005
R11707 gnd.n3364 gnd.n3267 9.3005
R11708 gnd.n5641 gnd.n3268 9.3005
R11709 gnd.n5642 gnd.n3269 9.3005
R11710 gnd.n5644 gnd.n5643 9.3005
R11711 gnd.n3359 gnd.n3287 9.3005
R11712 gnd.n5656 gnd.n3288 9.3005
R11713 gnd.n5657 gnd.n3289 9.3005
R11714 gnd.n5659 gnd.n5658 9.3005
R11715 gnd.n3354 gnd.n3309 9.3005
R11716 gnd.n5683 gnd.n3310 9.3005
R11717 gnd.n5684 gnd.n3311 9.3005
R11718 gnd.n5685 gnd.n3353 9.3005
R11719 gnd.n5689 gnd.n5688 9.3005
R11720 gnd.n5694 gnd.n3352 9.3005
R11721 gnd.n5696 gnd.n5695 9.3005
R11722 gnd.n5697 gnd.n3344 9.3005
R11723 gnd.n5698 gnd.n3345 9.3005
R11724 gnd.n5799 gnd.n3346 9.3005
R11725 gnd.n5798 gnd.n5699 9.3005
R11726 gnd.n5797 gnd.n5700 9.3005
R11727 gnd.n5702 gnd.n5701 9.3005
R11728 gnd.n5731 gnd.n125 9.3005
R11729 gnd.n5732 gnd.n126 9.3005
R11730 gnd.n5733 gnd.n127 9.3005
R11731 gnd.n5775 gnd.n5734 9.3005
R11732 gnd.n5774 gnd.n143 9.3005
R11733 gnd.n5773 gnd.n144 9.3005
R11734 gnd.n5735 gnd.n145 9.3005
R11735 gnd.n5763 gnd.n5760 9.3005
R11736 gnd.n5762 gnd.n164 9.3005
R11737 gnd.n5761 gnd.n165 9.3005
R11738 gnd.n355 gnd.n166 9.3005
R11739 gnd.n7703 gnd.n356 9.3005
R11740 gnd.n7704 gnd.n183 9.3005
R11741 gnd.n7706 gnd.n184 9.3005
R11742 gnd.n7707 gnd.n185 9.3005
R11743 gnd.n7710 gnd.n7708 9.3005
R11744 gnd.n7711 gnd.n204 9.3005
R11745 gnd.n7713 gnd.n205 9.3005
R11746 gnd.n7714 gnd.n206 9.3005
R11747 gnd.n7717 gnd.n7715 9.3005
R11748 gnd.n7718 gnd.n222 9.3005
R11749 gnd.n7720 gnd.n223 9.3005
R11750 gnd.n7721 gnd.n224 9.3005
R11751 gnd.n7724 gnd.n7722 9.3005
R11752 gnd.n7725 gnd.n242 9.3005
R11753 gnd.n7727 gnd.n243 9.3005
R11754 gnd.n7728 gnd.n244 9.3005
R11755 gnd.n7732 gnd.n7731 9.3005
R11756 gnd.n3178 gnd.n3172 9.3005
R11757 gnd.n5914 gnd.n5913 9.3005
R11758 gnd.n5917 gnd.n3170 9.3005
R11759 gnd.n5918 gnd.n3169 9.3005
R11760 gnd.n5921 gnd.n3168 9.3005
R11761 gnd.n5922 gnd.n3167 9.3005
R11762 gnd.n5925 gnd.n3166 9.3005
R11763 gnd.n5926 gnd.n3165 9.3005
R11764 gnd.n5929 gnd.n3164 9.3005
R11765 gnd.n5930 gnd.n3163 9.3005
R11766 gnd.n5933 gnd.n3162 9.3005
R11767 gnd.n5934 gnd.n3161 9.3005
R11768 gnd.n5937 gnd.n3160 9.3005
R11769 gnd.n5938 gnd.n3159 9.3005
R11770 gnd.n5941 gnd.n3158 9.3005
R11771 gnd.n5942 gnd.n3157 9.3005
R11772 gnd.n5945 gnd.n3156 9.3005
R11773 gnd.n5946 gnd.n3155 9.3005
R11774 gnd.n5949 gnd.n3154 9.3005
R11775 gnd.n5950 gnd.n3153 9.3005
R11776 gnd.n5953 gnd.n3152 9.3005
R11777 gnd.n5957 gnd.n3148 9.3005
R11778 gnd.n5958 gnd.n3147 9.3005
R11779 gnd.n5961 gnd.n3146 9.3005
R11780 gnd.n5962 gnd.n3145 9.3005
R11781 gnd.n5965 gnd.n3144 9.3005
R11782 gnd.n5966 gnd.n3143 9.3005
R11783 gnd.n5969 gnd.n3142 9.3005
R11784 gnd.n5970 gnd.n3141 9.3005
R11785 gnd.n5973 gnd.n3140 9.3005
R11786 gnd.n5975 gnd.n3136 9.3005
R11787 gnd.n5978 gnd.n3135 9.3005
R11788 gnd.n5979 gnd.n3134 9.3005
R11789 gnd.n5982 gnd.n3133 9.3005
R11790 gnd.n5983 gnd.n3132 9.3005
R11791 gnd.n5986 gnd.n3131 9.3005
R11792 gnd.n5987 gnd.n3130 9.3005
R11793 gnd.n5990 gnd.n3129 9.3005
R11794 gnd.n5992 gnd.n3126 9.3005
R11795 gnd.n5995 gnd.n3125 9.3005
R11796 gnd.n5996 gnd.n3124 9.3005
R11797 gnd.n5999 gnd.n3123 9.3005
R11798 gnd.n6000 gnd.n3122 9.3005
R11799 gnd.n6003 gnd.n3121 9.3005
R11800 gnd.n6004 gnd.n3120 9.3005
R11801 gnd.n6007 gnd.n3119 9.3005
R11802 gnd.n6008 gnd.n3118 9.3005
R11803 gnd.n6011 gnd.n3117 9.3005
R11804 gnd.n6012 gnd.n3116 9.3005
R11805 gnd.n6015 gnd.n3115 9.3005
R11806 gnd.n6016 gnd.n3114 9.3005
R11807 gnd.n6019 gnd.n3113 9.3005
R11808 gnd.n6021 gnd.n3112 9.3005
R11809 gnd.n6022 gnd.n3111 9.3005
R11810 gnd.n6023 gnd.n3110 9.3005
R11811 gnd.n6024 gnd.n3109 9.3005
R11812 gnd.n5954 gnd.n3149 9.3005
R11813 gnd.n5912 gnd.n5909 9.3005
R11814 gnd.n3191 gnd.n3188 9.3005
R11815 gnd.n5896 gnd.n3192 9.3005
R11816 gnd.n5895 gnd.n3193 9.3005
R11817 gnd.n5894 gnd.n3194 9.3005
R11818 gnd.n3215 gnd.n3195 9.3005
R11819 gnd.n5884 gnd.n3216 9.3005
R11820 gnd.n5883 gnd.n3217 9.3005
R11821 gnd.n5882 gnd.n3218 9.3005
R11822 gnd.n3236 gnd.n3219 9.3005
R11823 gnd.n5872 gnd.n3237 9.3005
R11824 gnd.n5871 gnd.n3238 9.3005
R11825 gnd.n5870 gnd.n3239 9.3005
R11826 gnd.n3256 gnd.n3240 9.3005
R11827 gnd.n5860 gnd.n3257 9.3005
R11828 gnd.n5859 gnd.n3258 9.3005
R11829 gnd.n5858 gnd.n3259 9.3005
R11830 gnd.n3277 gnd.n3260 9.3005
R11831 gnd.n5848 gnd.n3278 9.3005
R11832 gnd.n5847 gnd.n3279 9.3005
R11833 gnd.n5846 gnd.n3280 9.3005
R11834 gnd.n3297 gnd.n3281 9.3005
R11835 gnd.n5836 gnd.n3298 9.3005
R11836 gnd.n5835 gnd.n3299 9.3005
R11837 gnd.n5834 gnd.n3300 9.3005
R11838 gnd.n3302 gnd.n3301 9.3005
R11839 gnd.n5824 gnd.n110 9.3005
R11840 gnd.n115 gnd.n109 9.3005
R11841 gnd.n7931 gnd.n134 9.3005
R11842 gnd.n7930 gnd.n135 9.3005
R11843 gnd.n7929 gnd.n136 9.3005
R11844 gnd.n153 gnd.n137 9.3005
R11845 gnd.n7919 gnd.n154 9.3005
R11846 gnd.n7918 gnd.n155 9.3005
R11847 gnd.n7917 gnd.n156 9.3005
R11848 gnd.n173 gnd.n157 9.3005
R11849 gnd.n7907 gnd.n174 9.3005
R11850 gnd.n7906 gnd.n175 9.3005
R11851 gnd.n7905 gnd.n176 9.3005
R11852 gnd.n193 gnd.n177 9.3005
R11853 gnd.n7895 gnd.n194 9.3005
R11854 gnd.n7894 gnd.n195 9.3005
R11855 gnd.n7893 gnd.n196 9.3005
R11856 gnd.n213 gnd.n197 9.3005
R11857 gnd.n7883 gnd.n214 9.3005
R11858 gnd.n7882 gnd.n215 9.3005
R11859 gnd.n7881 gnd.n216 9.3005
R11860 gnd.n232 gnd.n217 9.3005
R11861 gnd.n7871 gnd.n233 9.3005
R11862 gnd.n7870 gnd.n234 9.3005
R11863 gnd.n7869 gnd.n235 9.3005
R11864 gnd.n251 gnd.n236 9.3005
R11865 gnd.n7859 gnd.n252 9.3005
R11866 gnd.n7858 gnd.n7857 9.3005
R11867 gnd.n3190 gnd.n3189 9.3005
R11868 gnd.n7942 gnd.n7941 9.3005
R11869 gnd.n4323 gnd.n4322 9.3005
R11870 gnd.n4345 gnd.n4324 9.3005
R11871 gnd.n4344 gnd.n4325 9.3005
R11872 gnd.n4343 gnd.n4326 9.3005
R11873 gnd.n4329 gnd.n4327 9.3005
R11874 gnd.n4339 gnd.n4330 9.3005
R11875 gnd.n4338 gnd.n4331 9.3005
R11876 gnd.n4337 gnd.n4332 9.3005
R11877 gnd.n4335 gnd.n4334 9.3005
R11878 gnd.n4333 gnd.n3962 9.3005
R11879 gnd.n3960 gnd.n3959 9.3005
R11880 gnd.n4411 gnd.n4410 9.3005
R11881 gnd.n4412 gnd.n3958 9.3005
R11882 gnd.n4414 gnd.n4413 9.3005
R11883 gnd.n3956 gnd.n3955 9.3005
R11884 gnd.n4419 gnd.n4418 9.3005
R11885 gnd.n4420 gnd.n3954 9.3005
R11886 gnd.n4448 gnd.n4421 9.3005
R11887 gnd.n4447 gnd.n4422 9.3005
R11888 gnd.n4446 gnd.n4423 9.3005
R11889 gnd.n4426 gnd.n4424 9.3005
R11890 gnd.n4442 gnd.n4427 9.3005
R11891 gnd.n4441 gnd.n4428 9.3005
R11892 gnd.n4440 gnd.n4429 9.3005
R11893 gnd.n4431 gnd.n4430 9.3005
R11894 gnd.n4436 gnd.n4432 9.3005
R11895 gnd.n4435 gnd.n4434 9.3005
R11896 gnd.n4433 gnd.n3934 9.3005
R11897 gnd.n3932 gnd.n3931 9.3005
R11898 gnd.n4774 gnd.n4773 9.3005
R11899 gnd.n4775 gnd.n3930 9.3005
R11900 gnd.n4779 gnd.n4776 9.3005
R11901 gnd.n4778 gnd.n4777 9.3005
R11902 gnd.n3903 gnd.n3902 9.3005
R11903 gnd.n4792 gnd.n4791 9.3005
R11904 gnd.n4793 gnd.n3901 9.3005
R11905 gnd.n4795 gnd.n4794 9.3005
R11906 gnd.n3888 gnd.n3887 9.3005
R11907 gnd.n4808 gnd.n4807 9.3005
R11908 gnd.n4809 gnd.n3886 9.3005
R11909 gnd.n4811 gnd.n4810 9.3005
R11910 gnd.n3874 gnd.n3873 9.3005
R11911 gnd.n4824 gnd.n4823 9.3005
R11912 gnd.n4825 gnd.n3872 9.3005
R11913 gnd.n4827 gnd.n4826 9.3005
R11914 gnd.n3859 gnd.n3858 9.3005
R11915 gnd.n4851 gnd.n4850 9.3005
R11916 gnd.n4852 gnd.n3857 9.3005
R11917 gnd.n4857 gnd.n4853 9.3005
R11918 gnd.n4856 gnd.n4855 9.3005
R11919 gnd.n4854 gnd.n2903 9.3005
R11920 gnd.n6197 gnd.n2904 9.3005
R11921 gnd.n6196 gnd.n2905 9.3005
R11922 gnd.n6195 gnd.n2906 9.3005
R11923 gnd.n3767 gnd.n2907 9.3005
R11924 gnd.n3769 gnd.n3768 9.3005
R11925 gnd.n3749 gnd.n3748 9.3005
R11926 gnd.n4925 gnd.n4924 9.3005
R11927 gnd.n4926 gnd.n3747 9.3005
R11928 gnd.n4928 gnd.n4927 9.3005
R11929 gnd.n3725 gnd.n3724 9.3005
R11930 gnd.n4964 gnd.n4963 9.3005
R11931 gnd.n4965 gnd.n3723 9.3005
R11932 gnd.n4967 gnd.n4966 9.3005
R11933 gnd.n3699 gnd.n3698 9.3005
R11934 gnd.n5004 gnd.n5003 9.3005
R11935 gnd.n5005 gnd.n3697 9.3005
R11936 gnd.n5009 gnd.n5006 9.3005
R11937 gnd.n5008 gnd.n5007 9.3005
R11938 gnd.n3672 gnd.n3671 9.3005
R11939 gnd.n5050 gnd.n5049 9.3005
R11940 gnd.n5051 gnd.n3670 9.3005
R11941 gnd.n5055 gnd.n5052 9.3005
R11942 gnd.n5054 gnd.n5053 9.3005
R11943 gnd.n3650 gnd.n3649 9.3005
R11944 gnd.n5103 gnd.n5102 9.3005
R11945 gnd.n5104 gnd.n3648 9.3005
R11946 gnd.n5108 gnd.n5105 9.3005
R11947 gnd.n5107 gnd.n5106 9.3005
R11948 gnd.n3624 gnd.n3623 9.3005
R11949 gnd.n5139 gnd.n5138 9.3005
R11950 gnd.n5140 gnd.n3622 9.3005
R11951 gnd.n5142 gnd.n5141 9.3005
R11952 gnd.n3598 gnd.n3597 9.3005
R11953 gnd.n5181 gnd.n5180 9.3005
R11954 gnd.n5182 gnd.n3596 9.3005
R11955 gnd.n5186 gnd.n5183 9.3005
R11956 gnd.n5185 gnd.n5184 9.3005
R11957 gnd.n3574 gnd.n3573 9.3005
R11958 gnd.n5233 gnd.n5232 9.3005
R11959 gnd.n5234 gnd.n3572 9.3005
R11960 gnd.n5236 gnd.n5235 9.3005
R11961 gnd.n3556 gnd.n3555 9.3005
R11962 gnd.n5262 gnd.n5261 9.3005
R11963 gnd.n5263 gnd.n3554 9.3005
R11964 gnd.n5265 gnd.n5264 9.3005
R11965 gnd.n3465 gnd.n3464 9.3005
R11966 gnd.n5409 gnd.n5408 9.3005
R11967 gnd.n5410 gnd.n3463 9.3005
R11968 gnd.n5412 gnd.n5411 9.3005
R11969 gnd.n3452 gnd.n3451 9.3005
R11970 gnd.n5425 gnd.n5424 9.3005
R11971 gnd.n5426 gnd.n3450 9.3005
R11972 gnd.n5428 gnd.n5427 9.3005
R11973 gnd.n3439 gnd.n3438 9.3005
R11974 gnd.n5441 gnd.n5440 9.3005
R11975 gnd.n5442 gnd.n3437 9.3005
R11976 gnd.n5444 gnd.n5443 9.3005
R11977 gnd.n3426 gnd.n3425 9.3005
R11978 gnd.n5457 gnd.n5456 9.3005
R11979 gnd.n5458 gnd.n3424 9.3005
R11980 gnd.n5463 gnd.n5459 9.3005
R11981 gnd.n5462 gnd.n5461 9.3005
R11982 gnd.n5460 gnd.n3413 9.3005
R11983 gnd.n5476 gnd.n3412 9.3005
R11984 gnd.n5478 gnd.n5477 9.3005
R11985 gnd.n5479 gnd.n3411 9.3005
R11986 gnd.n5573 gnd.n5480 9.3005
R11987 gnd.n5572 gnd.n5481 9.3005
R11988 gnd.n5571 gnd.n5482 9.3005
R11989 gnd.n5485 gnd.n5483 9.3005
R11990 gnd.n5567 gnd.n5486 9.3005
R11991 gnd.n5566 gnd.n5487 9.3005
R11992 gnd.n5565 gnd.n5488 9.3005
R11993 gnd.n5491 gnd.n5489 9.3005
R11994 gnd.n5559 gnd.n5492 9.3005
R11995 gnd.n5558 gnd.n5493 9.3005
R11996 gnd.n5557 gnd.n5494 9.3005
R11997 gnd.n5497 gnd.n5495 9.3005
R11998 gnd.n5553 gnd.n5498 9.3005
R11999 gnd.n5552 gnd.n5499 9.3005
R12000 gnd.n5551 gnd.n5500 9.3005
R12001 gnd.n5503 gnd.n5501 9.3005
R12002 gnd.n5547 gnd.n5504 9.3005
R12003 gnd.n5546 gnd.n5505 9.3005
R12004 gnd.n5545 gnd.n5506 9.3005
R12005 gnd.n5509 gnd.n5507 9.3005
R12006 gnd.n5541 gnd.n5510 9.3005
R12007 gnd.n5540 gnd.n5511 9.3005
R12008 gnd.n5539 gnd.n5512 9.3005
R12009 gnd.n5515 gnd.n5513 9.3005
R12010 gnd.n5535 gnd.n5516 9.3005
R12011 gnd.n5534 gnd.n5517 9.3005
R12012 gnd.n5533 gnd.n5518 9.3005
R12013 gnd.n5521 gnd.n5519 9.3005
R12014 gnd.n5529 gnd.n5522 9.3005
R12015 gnd.n5528 gnd.n5523 9.3005
R12016 gnd.n5527 gnd.n5525 9.3005
R12017 gnd.n5524 gnd.n3324 9.3005
R12018 gnd.n5787 gnd.n5716 9.3005
R12019 gnd.n5739 gnd.n5717 9.3005
R12020 gnd.n5741 gnd.n5740 9.3005
R12021 gnd.n5742 gnd.n5738 9.3005
R12022 gnd.n5753 gnd.n5743 9.3005
R12023 gnd.n5752 gnd.n5744 9.3005
R12024 gnd.n5751 gnd.n5745 9.3005
R12025 gnd.n5748 gnd.n5747 9.3005
R12026 gnd.n5746 gnd.n363 9.3005
R12027 gnd.n7593 gnd.n364 9.3005
R12028 gnd.n7592 gnd.n365 9.3005
R12029 gnd.n7591 gnd.n366 9.3005
R12030 gnd.n7584 gnd.n367 9.3005
R12031 gnd.n4285 gnd.n4284 9.3005
R12032 gnd.n4138 gnd.n4076 9.3005
R12033 gnd.n4141 gnd.n4140 9.3005
R12034 gnd.n4142 gnd.n4075 9.3005
R12035 gnd.n4145 gnd.n4143 9.3005
R12036 gnd.n4146 gnd.n4074 9.3005
R12037 gnd.n4149 gnd.n4148 9.3005
R12038 gnd.n4150 gnd.n4073 9.3005
R12039 gnd.n4153 gnd.n4151 9.3005
R12040 gnd.n4154 gnd.n4072 9.3005
R12041 gnd.n4157 gnd.n4156 9.3005
R12042 gnd.n4158 gnd.n4071 9.3005
R12043 gnd.n4161 gnd.n4159 9.3005
R12044 gnd.n4162 gnd.n4070 9.3005
R12045 gnd.n4165 gnd.n4164 9.3005
R12046 gnd.n4166 gnd.n4069 9.3005
R12047 gnd.n4169 gnd.n4168 9.3005
R12048 gnd.n4167 gnd.n4041 9.3005
R12049 gnd.n4187 gnd.n4042 9.3005
R12050 gnd.n4186 gnd.n4043 9.3005
R12051 gnd.n4185 gnd.n4044 9.3005
R12052 gnd.n4034 gnd.n4033 9.3005
R12053 gnd.n4223 gnd.n4222 9.3005
R12054 gnd.n4224 gnd.n4032 9.3005
R12055 gnd.n4227 gnd.n4226 9.3005
R12056 gnd.n4225 gnd.n4027 9.3005
R12057 gnd.n4251 gnd.n4028 9.3005
R12058 gnd.n4250 gnd.n4029 9.3005
R12059 gnd.n4249 gnd.n4030 9.3005
R12060 gnd.n4016 gnd.n4015 9.3005
R12061 gnd.n4282 gnd.n4281 9.3005
R12062 gnd.n4283 gnd.n4014 9.3005
R12063 gnd.n4137 gnd.n4135 9.3005
R12064 gnd.n4131 gnd.n4130 9.3005
R12065 gnd.n4129 gnd.n4081 9.3005
R12066 gnd.n4128 gnd.n4127 9.3005
R12067 gnd.n4124 gnd.n4084 9.3005
R12068 gnd.n4123 gnd.n4120 9.3005
R12069 gnd.n4119 gnd.n4085 9.3005
R12070 gnd.n4118 gnd.n4117 9.3005
R12071 gnd.n4114 gnd.n4086 9.3005
R12072 gnd.n4113 gnd.n4110 9.3005
R12073 gnd.n4109 gnd.n4087 9.3005
R12074 gnd.n4108 gnd.n4107 9.3005
R12075 gnd.n4104 gnd.n4088 9.3005
R12076 gnd.n4103 gnd.n4100 9.3005
R12077 gnd.n4099 gnd.n4089 9.3005
R12078 gnd.n4098 gnd.n4097 9.3005
R12079 gnd.n4094 gnd.n4090 9.3005
R12080 gnd.n4093 gnd.n2462 9.3005
R12081 gnd.n4132 gnd.n4077 9.3005
R12082 gnd.n4134 gnd.n4133 9.3005
R12083 gnd.n6275 gnd.n2831 9.3005
R12084 gnd.n6278 gnd.n2830 9.3005
R12085 gnd.n6279 gnd.n2829 9.3005
R12086 gnd.n6282 gnd.n2828 9.3005
R12087 gnd.n6283 gnd.n2827 9.3005
R12088 gnd.n6286 gnd.n2826 9.3005
R12089 gnd.n6287 gnd.n2825 9.3005
R12090 gnd.n6290 gnd.n2824 9.3005
R12091 gnd.n6292 gnd.n2821 9.3005
R12092 gnd.n6295 gnd.n2820 9.3005
R12093 gnd.n6296 gnd.n2819 9.3005
R12094 gnd.n6299 gnd.n2818 9.3005
R12095 gnd.n6300 gnd.n2817 9.3005
R12096 gnd.n6303 gnd.n2816 9.3005
R12097 gnd.n6304 gnd.n2815 9.3005
R12098 gnd.n6307 gnd.n2814 9.3005
R12099 gnd.n6308 gnd.n2813 9.3005
R12100 gnd.n6311 gnd.n2812 9.3005
R12101 gnd.n6312 gnd.n2811 9.3005
R12102 gnd.n6315 gnd.n2810 9.3005
R12103 gnd.n6316 gnd.n2809 9.3005
R12104 gnd.n6319 gnd.n2808 9.3005
R12105 gnd.n6320 gnd.n2807 9.3005
R12106 gnd.n6321 gnd.n2806 9.3005
R12107 gnd.n2763 gnd.n2762 9.3005
R12108 gnd.n6327 gnd.n6326 9.3005
R12109 gnd.n4682 gnd.n4679 9.3005
R12110 gnd.n4686 gnd.n4685 9.3005
R12111 gnd.n4687 gnd.n4677 9.3005
R12112 gnd.n4689 gnd.n4688 9.3005
R12113 gnd.n4692 gnd.n4676 9.3005
R12114 gnd.n4696 gnd.n4695 9.3005
R12115 gnd.n4697 gnd.n4675 9.3005
R12116 gnd.n4700 gnd.n4698 9.3005
R12117 gnd.n4701 gnd.n4671 9.3005
R12118 gnd.n4705 gnd.n4704 9.3005
R12119 gnd.n4706 gnd.n4670 9.3005
R12120 gnd.n4708 gnd.n4707 9.3005
R12121 gnd.n4711 gnd.n4669 9.3005
R12122 gnd.n4715 gnd.n4714 9.3005
R12123 gnd.n4716 gnd.n4668 9.3005
R12124 gnd.n4718 gnd.n4717 9.3005
R12125 gnd.n4721 gnd.n4667 9.3005
R12126 gnd.n4725 gnd.n4724 9.3005
R12127 gnd.n4726 gnd.n4666 9.3005
R12128 gnd.n4728 gnd.n4727 9.3005
R12129 gnd.n4731 gnd.n4665 9.3005
R12130 gnd.n4735 gnd.n4734 9.3005
R12131 gnd.n4736 gnd.n4664 9.3005
R12132 gnd.n4738 gnd.n4737 9.3005
R12133 gnd.n4741 gnd.n4663 9.3005
R12134 gnd.n4745 gnd.n4744 9.3005
R12135 gnd.n4746 gnd.n4662 9.3005
R12136 gnd.n4749 gnd.n4747 9.3005
R12137 gnd.n4750 gnd.n4658 9.3005
R12138 gnd.n4753 gnd.n4752 9.3005
R12139 gnd.n4678 gnd.n2832 9.3005
R12140 gnd.n2484 gnd.n2464 9.3005
R12141 gnd.n4045 gnd.n2485 9.3005
R12142 gnd.n6493 gnd.n2486 9.3005
R12143 gnd.n6492 gnd.n2487 9.3005
R12144 gnd.n6491 gnd.n2488 9.3005
R12145 gnd.n4051 gnd.n2489 9.3005
R12146 gnd.n6481 gnd.n2505 9.3005
R12147 gnd.n6480 gnd.n2506 9.3005
R12148 gnd.n6479 gnd.n2507 9.3005
R12149 gnd.n4058 gnd.n2508 9.3005
R12150 gnd.n6469 gnd.n2524 9.3005
R12151 gnd.n6468 gnd.n2525 9.3005
R12152 gnd.n6467 gnd.n2526 9.3005
R12153 gnd.n4065 gnd.n2527 9.3005
R12154 gnd.n6457 gnd.n2544 9.3005
R12155 gnd.n6456 gnd.n2545 9.3005
R12156 gnd.n6455 gnd.n2546 9.3005
R12157 gnd.n4175 gnd.n2547 9.3005
R12158 gnd.n6445 gnd.n2564 9.3005
R12159 gnd.n6444 gnd.n2565 9.3005
R12160 gnd.n6443 gnd.n2566 9.3005
R12161 gnd.n4178 gnd.n2567 9.3005
R12162 gnd.n6433 gnd.n2584 9.3005
R12163 gnd.n6432 gnd.n2585 9.3005
R12164 gnd.n6431 gnd.n2586 9.3005
R12165 gnd.n4233 gnd.n2587 9.3005
R12166 gnd.n6421 gnd.n2603 9.3005
R12167 gnd.n6420 gnd.n2604 9.3005
R12168 gnd.n6419 gnd.n2605 9.3005
R12169 gnd.n4242 gnd.n2606 9.3005
R12170 gnd.n4241 gnd.n4240 9.3005
R12171 gnd.n4010 gnd.n4005 9.3005
R12172 gnd.n4301 gnd.n4006 9.3005
R12173 gnd.n4300 gnd.n4007 9.3005
R12174 gnd.n4299 gnd.n4297 9.3005
R12175 gnd.n4008 gnd.n2630 9.3005
R12176 gnd.n6408 gnd.n2631 9.3005
R12177 gnd.n6407 gnd.n2632 9.3005
R12178 gnd.n6406 gnd.n2633 9.3005
R12179 gnd.n3978 gnd.n2634 9.3005
R12180 gnd.n6396 gnd.n2649 9.3005
R12181 gnd.n6395 gnd.n2650 9.3005
R12182 gnd.n6394 gnd.n2651 9.3005
R12183 gnd.n3972 gnd.n2652 9.3005
R12184 gnd.n6384 gnd.n2670 9.3005
R12185 gnd.n6383 gnd.n2671 9.3005
R12186 gnd.n6382 gnd.n2672 9.3005
R12187 gnd.n4376 gnd.n2673 9.3005
R12188 gnd.n6372 gnd.n2689 9.3005
R12189 gnd.n6371 gnd.n2690 9.3005
R12190 gnd.n6370 gnd.n2691 9.3005
R12191 gnd.n4386 gnd.n2692 9.3005
R12192 gnd.n6360 gnd.n2710 9.3005
R12193 gnd.n6359 gnd.n2711 9.3005
R12194 gnd.n6358 gnd.n2712 9.3005
R12195 gnd.n3947 gnd.n2713 9.3005
R12196 gnd.n6348 gnd.n2729 9.3005
R12197 gnd.n6347 gnd.n2730 9.3005
R12198 gnd.n6346 gnd.n2731 9.3005
R12199 gnd.n3941 gnd.n2732 9.3005
R12200 gnd.n6336 gnd.n2750 9.3005
R12201 gnd.n6335 gnd.n2751 9.3005
R12202 gnd.n6334 gnd.n2752 9.3005
R12203 gnd.n4755 gnd.n2753 9.3005
R12204 gnd.n6505 gnd.n2463 9.3005
R12205 gnd.n2465 gnd.n2464 9.3005
R12206 gnd.n4046 gnd.n4045 9.3005
R12207 gnd.n4047 gnd.n2486 9.3005
R12208 gnd.n4049 gnd.n2487 9.3005
R12209 gnd.n4050 gnd.n2488 9.3005
R12210 gnd.n4053 gnd.n4051 9.3005
R12211 gnd.n4054 gnd.n2505 9.3005
R12212 gnd.n4056 gnd.n2506 9.3005
R12213 gnd.n4057 gnd.n2507 9.3005
R12214 gnd.n4060 gnd.n4058 9.3005
R12215 gnd.n4061 gnd.n2524 9.3005
R12216 gnd.n4063 gnd.n2525 9.3005
R12217 gnd.n4064 gnd.n2526 9.3005
R12218 gnd.n4067 gnd.n4065 9.3005
R12219 gnd.n4068 gnd.n2544 9.3005
R12220 gnd.n4173 gnd.n2545 9.3005
R12221 gnd.n4174 gnd.n2546 9.3005
R12222 gnd.n4176 gnd.n4175 9.3005
R12223 gnd.n4177 gnd.n2564 9.3005
R12224 gnd.n4181 gnd.n2565 9.3005
R12225 gnd.n4180 gnd.n2566 9.3005
R12226 gnd.n4179 gnd.n4178 9.3005
R12227 gnd.n4031 gnd.n2584 9.3005
R12228 gnd.n4231 gnd.n2585 9.3005
R12229 gnd.n4232 gnd.n2586 9.3005
R12230 gnd.n4234 gnd.n4233 9.3005
R12231 gnd.n4235 gnd.n2603 9.3005
R12232 gnd.n4245 gnd.n2604 9.3005
R12233 gnd.n4244 gnd.n2605 9.3005
R12234 gnd.n4243 gnd.n4242 9.3005
R12235 gnd.n4241 gnd.n4009 9.3005
R12236 gnd.n4289 gnd.n4010 9.3005
R12237 gnd.n4290 gnd.n4006 9.3005
R12238 gnd.n4291 gnd.n4007 9.3005
R12239 gnd.n4297 gnd.n4296 9.3005
R12240 gnd.n4294 gnd.n4008 9.3005
R12241 gnd.n4293 gnd.n2631 9.3005
R12242 gnd.n4292 gnd.n2632 9.3005
R12243 gnd.n3977 gnd.n2633 9.3005
R12244 gnd.n4358 gnd.n3978 9.3005
R12245 gnd.n4359 gnd.n2649 9.3005
R12246 gnd.n4360 gnd.n2650 9.3005
R12247 gnd.n3971 gnd.n2651 9.3005
R12248 gnd.n4372 gnd.n3972 9.3005
R12249 gnd.n4373 gnd.n2670 9.3005
R12250 gnd.n4374 gnd.n2671 9.3005
R12251 gnd.n4375 gnd.n2672 9.3005
R12252 gnd.n4379 gnd.n4376 9.3005
R12253 gnd.n4380 gnd.n2689 9.3005
R12254 gnd.n4384 gnd.n2690 9.3005
R12255 gnd.n4385 gnd.n2691 9.3005
R12256 gnd.n4389 gnd.n4386 9.3005
R12257 gnd.n4388 gnd.n2710 9.3005
R12258 gnd.n4387 gnd.n2711 9.3005
R12259 gnd.n3946 gnd.n2712 9.3005
R12260 gnd.n4461 gnd.n3947 9.3005
R12261 gnd.n4462 gnd.n2729 9.3005
R12262 gnd.n4463 gnd.n2730 9.3005
R12263 gnd.n3940 gnd.n2731 9.3005
R12264 gnd.n4475 gnd.n3941 9.3005
R12265 gnd.n4476 gnd.n2750 9.3005
R12266 gnd.n4758 gnd.n2751 9.3005
R12267 gnd.n4757 gnd.n2752 9.3005
R12268 gnd.n4756 gnd.n4755 9.3005
R12269 gnd.n6505 gnd.n6504 9.3005
R12270 gnd.n6509 gnd.n6508 9.3005
R12271 gnd.n6512 gnd.n2458 9.3005
R12272 gnd.n6513 gnd.n2457 9.3005
R12273 gnd.n6516 gnd.n2456 9.3005
R12274 gnd.n6517 gnd.n2455 9.3005
R12275 gnd.n6520 gnd.n2454 9.3005
R12276 gnd.n6521 gnd.n2453 9.3005
R12277 gnd.n6524 gnd.n2452 9.3005
R12278 gnd.n6525 gnd.n2451 9.3005
R12279 gnd.n6528 gnd.n2450 9.3005
R12280 gnd.n6529 gnd.n2449 9.3005
R12281 gnd.n6532 gnd.n2448 9.3005
R12282 gnd.n6533 gnd.n2447 9.3005
R12283 gnd.n6536 gnd.n2446 9.3005
R12284 gnd.n6537 gnd.n2445 9.3005
R12285 gnd.n6540 gnd.n2444 9.3005
R12286 gnd.n6541 gnd.n2443 9.3005
R12287 gnd.n6544 gnd.n2442 9.3005
R12288 gnd.n6545 gnd.n2441 9.3005
R12289 gnd.n6548 gnd.n2440 9.3005
R12290 gnd.n6552 gnd.n2436 9.3005
R12291 gnd.n6553 gnd.n2435 9.3005
R12292 gnd.n6556 gnd.n2434 9.3005
R12293 gnd.n6557 gnd.n2433 9.3005
R12294 gnd.n6560 gnd.n2432 9.3005
R12295 gnd.n6561 gnd.n2431 9.3005
R12296 gnd.n6564 gnd.n2430 9.3005
R12297 gnd.n6565 gnd.n2429 9.3005
R12298 gnd.n6568 gnd.n2428 9.3005
R12299 gnd.n6569 gnd.n2427 9.3005
R12300 gnd.n6572 gnd.n2426 9.3005
R12301 gnd.n6573 gnd.n2425 9.3005
R12302 gnd.n6576 gnd.n2424 9.3005
R12303 gnd.n6577 gnd.n2423 9.3005
R12304 gnd.n6580 gnd.n2422 9.3005
R12305 gnd.n6581 gnd.n2421 9.3005
R12306 gnd.n6584 gnd.n2420 9.3005
R12307 gnd.n6585 gnd.n2419 9.3005
R12308 gnd.n6588 gnd.n2418 9.3005
R12309 gnd.n6590 gnd.n2415 9.3005
R12310 gnd.n6593 gnd.n2414 9.3005
R12311 gnd.n6594 gnd.n2413 9.3005
R12312 gnd.n6597 gnd.n2412 9.3005
R12313 gnd.n6598 gnd.n2411 9.3005
R12314 gnd.n6601 gnd.n2410 9.3005
R12315 gnd.n6602 gnd.n2409 9.3005
R12316 gnd.n6605 gnd.n2408 9.3005
R12317 gnd.n6606 gnd.n2407 9.3005
R12318 gnd.n6609 gnd.n2406 9.3005
R12319 gnd.n6610 gnd.n2405 9.3005
R12320 gnd.n6613 gnd.n2404 9.3005
R12321 gnd.n6614 gnd.n2403 9.3005
R12322 gnd.n6617 gnd.n2402 9.3005
R12323 gnd.n6619 gnd.n2401 9.3005
R12324 gnd.n6620 gnd.n2400 9.3005
R12325 gnd.n6621 gnd.n2399 9.3005
R12326 gnd.n6622 gnd.n2398 9.3005
R12327 gnd.n6549 gnd.n2437 9.3005
R12328 gnd.n6507 gnd.n2459 9.3005
R12329 gnd.n6499 gnd.n2473 9.3005
R12330 gnd.n6498 gnd.n2474 9.3005
R12331 gnd.n6497 gnd.n2475 9.3005
R12332 gnd.n2495 gnd.n2476 9.3005
R12333 gnd.n6487 gnd.n2496 9.3005
R12334 gnd.n6486 gnd.n2497 9.3005
R12335 gnd.n6485 gnd.n2498 9.3005
R12336 gnd.n2513 gnd.n2499 9.3005
R12337 gnd.n6475 gnd.n2514 9.3005
R12338 gnd.n6474 gnd.n2515 9.3005
R12339 gnd.n6473 gnd.n2516 9.3005
R12340 gnd.n2534 gnd.n2517 9.3005
R12341 gnd.n6463 gnd.n2535 9.3005
R12342 gnd.n6462 gnd.n2536 9.3005
R12343 gnd.n6461 gnd.n2537 9.3005
R12344 gnd.n2553 gnd.n2538 9.3005
R12345 gnd.n6451 gnd.n2554 9.3005
R12346 gnd.n6450 gnd.n2555 9.3005
R12347 gnd.n6449 gnd.n2556 9.3005
R12348 gnd.n2574 gnd.n2557 9.3005
R12349 gnd.n6439 gnd.n2575 9.3005
R12350 gnd.n6438 gnd.n2576 9.3005
R12351 gnd.n6437 gnd.n2577 9.3005
R12352 gnd.n2593 gnd.n2578 9.3005
R12353 gnd.n6427 gnd.n2594 9.3005
R12354 gnd.n6426 gnd.n2595 9.3005
R12355 gnd.n2621 gnd.n2615 9.3005
R12356 gnd.n6402 gnd.n2640 9.3005
R12357 gnd.n6401 gnd.n2641 9.3005
R12358 gnd.n6400 gnd.n2642 9.3005
R12359 gnd.n2659 gnd.n2643 9.3005
R12360 gnd.n6390 gnd.n2660 9.3005
R12361 gnd.n6389 gnd.n2661 9.3005
R12362 gnd.n6388 gnd.n2662 9.3005
R12363 gnd.n2679 gnd.n2663 9.3005
R12364 gnd.n6378 gnd.n2680 9.3005
R12365 gnd.n6377 gnd.n2681 9.3005
R12366 gnd.n6376 gnd.n2682 9.3005
R12367 gnd.n2699 gnd.n2683 9.3005
R12368 gnd.n6366 gnd.n2700 9.3005
R12369 gnd.n6365 gnd.n2701 9.3005
R12370 gnd.n6364 gnd.n2702 9.3005
R12371 gnd.n2719 gnd.n2703 9.3005
R12372 gnd.n6354 gnd.n2720 9.3005
R12373 gnd.n6353 gnd.n2721 9.3005
R12374 gnd.n6352 gnd.n2722 9.3005
R12375 gnd.n2739 gnd.n2723 9.3005
R12376 gnd.n6342 gnd.n2740 9.3005
R12377 gnd.n6341 gnd.n2741 9.3005
R12378 gnd.n6340 gnd.n2742 9.3005
R12379 gnd.n2760 gnd.n2743 9.3005
R12380 gnd.n6330 gnd.n2761 9.3005
R12381 gnd.n6329 gnd.n6328 9.3005
R12382 gnd.n2472 gnd.n2471 9.3005
R12383 gnd.n6413 gnd.n6412 9.3005
R12384 gnd.n4194 gnd.n4193 9.3005
R12385 gnd.n4206 gnd.n4205 9.3005
R12386 gnd.n4207 gnd.n4192 9.3005
R12387 gnd.n4209 gnd.n4208 9.3005
R12388 gnd.n4039 gnd.n4038 9.3005
R12389 gnd.n4214 gnd.n4213 9.3005
R12390 gnd.n4215 gnd.n4037 9.3005
R12391 gnd.n4217 gnd.n4216 9.3005
R12392 gnd.n4024 gnd.n4023 9.3005
R12393 gnd.n4258 gnd.n4257 9.3005
R12394 gnd.n4259 gnd.n4022 9.3005
R12395 gnd.n4261 gnd.n4260 9.3005
R12396 gnd.n4200 gnd.n4199 9.3005
R12397 gnd.n4196 gnd.n951 9.3005
R12398 gnd.n6721 gnd.n950 9.3005
R12399 gnd.n6722 gnd.n949 9.3005
R12400 gnd.n6723 gnd.n948 9.3005
R12401 gnd.n947 gnd.n943 9.3005
R12402 gnd.n6729 gnd.n942 9.3005
R12403 gnd.n6730 gnd.n941 9.3005
R12404 gnd.n6731 gnd.n940 9.3005
R12405 gnd.n939 gnd.n935 9.3005
R12406 gnd.n6737 gnd.n934 9.3005
R12407 gnd.n6738 gnd.n933 9.3005
R12408 gnd.n6739 gnd.n932 9.3005
R12409 gnd.n931 gnd.n927 9.3005
R12410 gnd.n6745 gnd.n926 9.3005
R12411 gnd.n6746 gnd.n925 9.3005
R12412 gnd.n6747 gnd.n924 9.3005
R12413 gnd.n923 gnd.n919 9.3005
R12414 gnd.n6753 gnd.n918 9.3005
R12415 gnd.n6754 gnd.n917 9.3005
R12416 gnd.n6755 gnd.n916 9.3005
R12417 gnd.n915 gnd.n911 9.3005
R12418 gnd.n6761 gnd.n910 9.3005
R12419 gnd.n6762 gnd.n909 9.3005
R12420 gnd.n6763 gnd.n908 9.3005
R12421 gnd.n907 gnd.n903 9.3005
R12422 gnd.n6769 gnd.n902 9.3005
R12423 gnd.n6770 gnd.n901 9.3005
R12424 gnd.n6771 gnd.n900 9.3005
R12425 gnd.n899 gnd.n895 9.3005
R12426 gnd.n6777 gnd.n894 9.3005
R12427 gnd.n6778 gnd.n893 9.3005
R12428 gnd.n6779 gnd.n892 9.3005
R12429 gnd.n891 gnd.n887 9.3005
R12430 gnd.n6785 gnd.n886 9.3005
R12431 gnd.n6786 gnd.n885 9.3005
R12432 gnd.n6787 gnd.n884 9.3005
R12433 gnd.n883 gnd.n879 9.3005
R12434 gnd.n6793 gnd.n878 9.3005
R12435 gnd.n6794 gnd.n877 9.3005
R12436 gnd.n6795 gnd.n876 9.3005
R12437 gnd.n875 gnd.n871 9.3005
R12438 gnd.n6801 gnd.n870 9.3005
R12439 gnd.n6802 gnd.n869 9.3005
R12440 gnd.n6803 gnd.n868 9.3005
R12441 gnd.n867 gnd.n863 9.3005
R12442 gnd.n6809 gnd.n862 9.3005
R12443 gnd.n6810 gnd.n861 9.3005
R12444 gnd.n6811 gnd.n860 9.3005
R12445 gnd.n859 gnd.n855 9.3005
R12446 gnd.n6817 gnd.n854 9.3005
R12447 gnd.n6818 gnd.n853 9.3005
R12448 gnd.n6819 gnd.n852 9.3005
R12449 gnd.n851 gnd.n847 9.3005
R12450 gnd.n6825 gnd.n846 9.3005
R12451 gnd.n6826 gnd.n845 9.3005
R12452 gnd.n6827 gnd.n844 9.3005
R12453 gnd.n843 gnd.n839 9.3005
R12454 gnd.n6833 gnd.n838 9.3005
R12455 gnd.n6834 gnd.n837 9.3005
R12456 gnd.n6835 gnd.n836 9.3005
R12457 gnd.n835 gnd.n831 9.3005
R12458 gnd.n6841 gnd.n830 9.3005
R12459 gnd.n6842 gnd.n829 9.3005
R12460 gnd.n6843 gnd.n828 9.3005
R12461 gnd.n827 gnd.n823 9.3005
R12462 gnd.n6849 gnd.n822 9.3005
R12463 gnd.n6850 gnd.n821 9.3005
R12464 gnd.n6851 gnd.n820 9.3005
R12465 gnd.n819 gnd.n815 9.3005
R12466 gnd.n6857 gnd.n814 9.3005
R12467 gnd.n6858 gnd.n813 9.3005
R12468 gnd.n6859 gnd.n812 9.3005
R12469 gnd.n811 gnd.n807 9.3005
R12470 gnd.n6865 gnd.n806 9.3005
R12471 gnd.n6866 gnd.n805 9.3005
R12472 gnd.n6867 gnd.n804 9.3005
R12473 gnd.n803 gnd.n799 9.3005
R12474 gnd.n6873 gnd.n798 9.3005
R12475 gnd.n6874 gnd.n797 9.3005
R12476 gnd.n6875 gnd.n796 9.3005
R12477 gnd.n795 gnd.n791 9.3005
R12478 gnd.n6881 gnd.n790 9.3005
R12479 gnd.n6882 gnd.n789 9.3005
R12480 gnd.n6883 gnd.n788 9.3005
R12481 gnd.n4198 gnd.n4197 9.3005
R12482 gnd.n5578 gnd.n2991 9.3005
R12483 gnd.n4787 gnd.n4786 9.3005
R12484 gnd.n3896 gnd.n3895 9.3005
R12485 gnd.n4800 gnd.n4799 9.3005
R12486 gnd.n4801 gnd.n3894 9.3005
R12487 gnd.n4803 gnd.n4802 9.3005
R12488 gnd.n3882 gnd.n3881 9.3005
R12489 gnd.n4816 gnd.n4815 9.3005
R12490 gnd.n4817 gnd.n3880 9.3005
R12491 gnd.n4819 gnd.n4818 9.3005
R12492 gnd.n3868 gnd.n3867 9.3005
R12493 gnd.n4832 gnd.n4831 9.3005
R12494 gnd.n4833 gnd.n3865 9.3005
R12495 gnd.n4846 gnd.n4845 9.3005
R12496 gnd.n4844 gnd.n3866 9.3005
R12497 gnd.n4843 gnd.n4842 9.3005
R12498 gnd.n4841 gnd.n4834 9.3005
R12499 gnd.n4840 gnd.n4839 9.3005
R12500 gnd.n4838 gnd.n4837 9.3005
R12501 gnd.n2915 gnd.n2913 9.3005
R12502 gnd.n6191 gnd.n6190 9.3005
R12503 gnd.n6189 gnd.n2914 9.3005
R12504 gnd.n6188 gnd.n6187 9.3005
R12505 gnd.n6186 gnd.n2916 9.3005
R12506 gnd.n6185 gnd.n6184 9.3005
R12507 gnd.n6183 gnd.n2920 9.3005
R12508 gnd.n6182 gnd.n6181 9.3005
R12509 gnd.n6180 gnd.n2921 9.3005
R12510 gnd.n6179 gnd.n6178 9.3005
R12511 gnd.n6177 gnd.n2925 9.3005
R12512 gnd.n6176 gnd.n6175 9.3005
R12513 gnd.n6174 gnd.n2926 9.3005
R12514 gnd.n6173 gnd.n6172 9.3005
R12515 gnd.n6171 gnd.n2930 9.3005
R12516 gnd.n6170 gnd.n6169 9.3005
R12517 gnd.n6168 gnd.n2931 9.3005
R12518 gnd.n6167 gnd.n6166 9.3005
R12519 gnd.n6165 gnd.n2935 9.3005
R12520 gnd.n6164 gnd.n6163 9.3005
R12521 gnd.n6162 gnd.n2936 9.3005
R12522 gnd.n6161 gnd.n6160 9.3005
R12523 gnd.n6159 gnd.n2940 9.3005
R12524 gnd.n6158 gnd.n6157 9.3005
R12525 gnd.n6156 gnd.n2941 9.3005
R12526 gnd.n6155 gnd.n6154 9.3005
R12527 gnd.n6153 gnd.n2945 9.3005
R12528 gnd.n6152 gnd.n6151 9.3005
R12529 gnd.n6150 gnd.n2946 9.3005
R12530 gnd.n6149 gnd.n6148 9.3005
R12531 gnd.n6147 gnd.n2950 9.3005
R12532 gnd.n6146 gnd.n6145 9.3005
R12533 gnd.n6144 gnd.n2951 9.3005
R12534 gnd.n6143 gnd.n6142 9.3005
R12535 gnd.n6141 gnd.n2955 9.3005
R12536 gnd.n6140 gnd.n6139 9.3005
R12537 gnd.n6138 gnd.n2956 9.3005
R12538 gnd.n6137 gnd.n6136 9.3005
R12539 gnd.n6135 gnd.n2960 9.3005
R12540 gnd.n6134 gnd.n6133 9.3005
R12541 gnd.n6132 gnd.n2961 9.3005
R12542 gnd.n6131 gnd.n6130 9.3005
R12543 gnd.n6129 gnd.n2965 9.3005
R12544 gnd.n6128 gnd.n6127 9.3005
R12545 gnd.n6126 gnd.n2966 9.3005
R12546 gnd.n6125 gnd.n6124 9.3005
R12547 gnd.n6123 gnd.n2970 9.3005
R12548 gnd.n6122 gnd.n6121 9.3005
R12549 gnd.n6120 gnd.n2971 9.3005
R12550 gnd.n6119 gnd.n6118 9.3005
R12551 gnd.n6117 gnd.n2975 9.3005
R12552 gnd.n6116 gnd.n6115 9.3005
R12553 gnd.n6114 gnd.n2976 9.3005
R12554 gnd.n6113 gnd.n6112 9.3005
R12555 gnd.n6111 gnd.n2980 9.3005
R12556 gnd.n6110 gnd.n6109 9.3005
R12557 gnd.n6108 gnd.n2981 9.3005
R12558 gnd.n6107 gnd.n6106 9.3005
R12559 gnd.n6105 gnd.n2985 9.3005
R12560 gnd.n6104 gnd.n6103 9.3005
R12561 gnd.n6102 gnd.n2986 9.3005
R12562 gnd.n6101 gnd.n6100 9.3005
R12563 gnd.n6099 gnd.n2990 9.3005
R12564 gnd.n6098 gnd.n6097 9.3005
R12565 gnd.n4785 gnd.n3908 9.3005
R12566 gnd.n4784 gnd.n4783 9.3005
R12567 gnd.n3993 gnd.n3992 9.3005
R12568 gnd.n4312 gnd.n4311 9.3005
R12569 gnd.n4313 gnd.n3991 9.3005
R12570 gnd.n4315 gnd.n4314 9.3005
R12571 gnd.n3981 gnd.n3980 9.3005
R12572 gnd.n4351 gnd.n4350 9.3005
R12573 gnd.n4352 gnd.n3979 9.3005
R12574 gnd.n4354 gnd.n4353 9.3005
R12575 gnd.n3975 gnd.n3974 9.3005
R12576 gnd.n4365 gnd.n4364 9.3005
R12577 gnd.n4366 gnd.n3973 9.3005
R12578 gnd.n4368 gnd.n4367 9.3005
R12579 gnd.n3966 gnd.n3964 9.3005
R12580 gnd.n4403 gnd.n4402 9.3005
R12581 gnd.n4401 gnd.n3965 9.3005
R12582 gnd.n4400 gnd.n4399 9.3005
R12583 gnd.n4398 gnd.n3967 9.3005
R12584 gnd.n4397 gnd.n4396 9.3005
R12585 gnd.n4395 gnd.n3970 9.3005
R12586 gnd.n4394 gnd.n4393 9.3005
R12587 gnd.n3950 gnd.n3949 9.3005
R12588 gnd.n4454 gnd.n4453 9.3005
R12589 gnd.n4455 gnd.n3948 9.3005
R12590 gnd.n4457 gnd.n4456 9.3005
R12591 gnd.n3944 gnd.n3943 9.3005
R12592 gnd.n4468 gnd.n4467 9.3005
R12593 gnd.n4469 gnd.n3942 9.3005
R12594 gnd.n4471 gnd.n4470 9.3005
R12595 gnd.n3939 gnd.n3938 9.3005
R12596 gnd.n4763 gnd.n4762 9.3005
R12597 gnd.n4764 gnd.n3937 9.3005
R12598 gnd.n4766 gnd.n4765 9.3005
R12599 gnd.n4649 gnd.n4648 9.3005
R12600 gnd.n4541 gnd.n4540 9.3005
R12601 gnd.n4643 gnd.n4642 9.3005
R12602 gnd.n4641 gnd.n4640 9.3005
R12603 gnd.n4553 gnd.n4552 9.3005
R12604 gnd.n4635 gnd.n4634 9.3005
R12605 gnd.n4633 gnd.n4632 9.3005
R12606 gnd.n4561 gnd.n4560 9.3005
R12607 gnd.n4627 gnd.n4626 9.3005
R12608 gnd.n4625 gnd.n4624 9.3005
R12609 gnd.n4573 gnd.n4572 9.3005
R12610 gnd.n4619 gnd.n4618 9.3005
R12611 gnd.n4617 gnd.n4616 9.3005
R12612 gnd.n4581 gnd.n4580 9.3005
R12613 gnd.n4611 gnd.n4610 9.3005
R12614 gnd.n4609 gnd.n4608 9.3005
R12615 gnd.n4595 gnd.n4594 9.3005
R12616 gnd.n4603 gnd.n4602 9.3005
R12617 gnd.n4651 gnd.n4650 9.3005
R12618 gnd.n4601 gnd.n3910 9.3005
R12619 gnd.n4605 gnd.n4604 9.3005
R12620 gnd.n4607 gnd.n4606 9.3005
R12621 gnd.n4587 gnd.n4586 9.3005
R12622 gnd.n4613 gnd.n4612 9.3005
R12623 gnd.n4615 gnd.n4614 9.3005
R12624 gnd.n4577 gnd.n4576 9.3005
R12625 gnd.n4621 gnd.n4620 9.3005
R12626 gnd.n4623 gnd.n4622 9.3005
R12627 gnd.n4567 gnd.n4566 9.3005
R12628 gnd.n4629 gnd.n4628 9.3005
R12629 gnd.n4631 gnd.n4630 9.3005
R12630 gnd.n4557 gnd.n4556 9.3005
R12631 gnd.n4637 gnd.n4636 9.3005
R12632 gnd.n4639 gnd.n4638 9.3005
R12633 gnd.n4547 gnd.n4546 9.3005
R12634 gnd.n4645 gnd.n4644 9.3005
R12635 gnd.n4647 gnd.n4646 9.3005
R12636 gnd.n4538 gnd.n4537 9.3005
R12637 gnd.n4653 gnd.n4652 9.3005
R12638 gnd.n4654 gnd.n4477 9.3005
R12639 gnd.n4656 gnd.n4655 9.3005
R12640 gnd.n4532 gnd.n4478 9.3005
R12641 gnd.n4531 gnd.n4530 9.3005
R12642 gnd.n4529 gnd.n4479 9.3005
R12643 gnd.n4528 gnd.n4527 9.3005
R12644 gnd.n4524 gnd.n4482 9.3005
R12645 gnd.n4523 gnd.n4483 9.3005
R12646 gnd.n4518 gnd.n4484 9.3005
R12647 gnd.n4517 gnd.n4516 9.3005
R12648 gnd.n4515 gnd.n4485 9.3005
R12649 gnd.n4514 gnd.n4513 9.3005
R12650 gnd.n4512 gnd.n4488 9.3005
R12651 gnd.n4511 gnd.n4510 9.3005
R12652 gnd.n4509 gnd.n4489 9.3005
R12653 gnd.n4508 gnd.n4507 9.3005
R12654 gnd.n4506 gnd.n4492 9.3005
R12655 gnd.n4505 gnd.n4504 9.3005
R12656 gnd.n4503 gnd.n4493 9.3005
R12657 gnd.n4502 gnd.n4501 9.3005
R12658 gnd.n4500 gnd.n4496 9.3005
R12659 gnd.n4499 gnd.n4498 9.3005
R12660 gnd.n4497 gnd.n3852 9.3005
R12661 gnd.n3850 gnd.n3849 9.3005
R12662 gnd.n4864 gnd.n4863 9.3005
R12663 gnd.n4865 gnd.n3848 9.3005
R12664 gnd.n4867 gnd.n4866 9.3005
R12665 gnd.n3764 gnd.n3763 9.3005
R12666 gnd.n4903 gnd.n4902 9.3005
R12667 gnd.n4904 gnd.n3761 9.3005
R12668 gnd.n4909 gnd.n4908 9.3005
R12669 gnd.n4907 gnd.n3762 9.3005
R12670 gnd.n4906 gnd.n4905 9.3005
R12671 gnd.n3742 gnd.n3741 9.3005
R12672 gnd.n4934 gnd.n4933 9.3005
R12673 gnd.n4935 gnd.n3739 9.3005
R12674 gnd.n4943 gnd.n4942 9.3005
R12675 gnd.n4941 gnd.n3740 9.3005
R12676 gnd.n4940 gnd.n4939 9.3005
R12677 gnd.n4938 gnd.n4936 9.3005
R12678 gnd.n3692 gnd.n3691 9.3005
R12679 gnd.n5014 gnd.n5013 9.3005
R12680 gnd.n5015 gnd.n3689 9.3005
R12681 gnd.n5018 gnd.n5017 9.3005
R12682 gnd.n5016 gnd.n3690 9.3005
R12683 gnd.n3665 gnd.n3664 9.3005
R12684 gnd.n5060 gnd.n5059 9.3005
R12685 gnd.n5061 gnd.n3662 9.3005
R12686 gnd.n5089 gnd.n5088 9.3005
R12687 gnd.n5087 gnd.n3663 9.3005
R12688 gnd.n5086 gnd.n5085 9.3005
R12689 gnd.n5084 gnd.n5062 9.3005
R12690 gnd.n5083 gnd.n5082 9.3005
R12691 gnd.n5081 gnd.n5067 9.3005
R12692 gnd.n5080 gnd.n5079 9.3005
R12693 gnd.n5078 gnd.n5068 9.3005
R12694 gnd.n5077 gnd.n5076 9.3005
R12695 gnd.n5075 gnd.n5072 9.3005
R12696 gnd.n5074 gnd.n5073 9.3005
R12697 gnd.n3590 gnd.n3589 9.3005
R12698 gnd.n5191 gnd.n5190 9.3005
R12699 gnd.n5192 gnd.n3587 9.3005
R12700 gnd.n5217 gnd.n5216 9.3005
R12701 gnd.n5215 gnd.n3588 9.3005
R12702 gnd.n5214 gnd.n5213 9.3005
R12703 gnd.n5212 gnd.n5193 9.3005
R12704 gnd.n5211 gnd.n5210 9.3005
R12705 gnd.n5209 gnd.n5198 9.3005
R12706 gnd.n5208 gnd.n5207 9.3005
R12707 gnd.n5206 gnd.n5199 9.3005
R12708 gnd.n5205 gnd.n5204 9.3005
R12709 gnd.n5203 gnd.n5202 9.3005
R12710 gnd.n3458 gnd.n3457 9.3005
R12711 gnd.n5417 gnd.n5416 9.3005
R12712 gnd.n5418 gnd.n3456 9.3005
R12713 gnd.n5420 gnd.n5419 9.3005
R12714 gnd.n3444 gnd.n3443 9.3005
R12715 gnd.n5433 gnd.n5432 9.3005
R12716 gnd.n5434 gnd.n3442 9.3005
R12717 gnd.n5436 gnd.n5435 9.3005
R12718 gnd.n3431 gnd.n3430 9.3005
R12719 gnd.n5449 gnd.n5448 9.3005
R12720 gnd.n5450 gnd.n3429 9.3005
R12721 gnd.n5452 gnd.n5451 9.3005
R12722 gnd.n3419 gnd.n3418 9.3005
R12723 gnd.n5468 gnd.n5467 9.3005
R12724 gnd.n5469 gnd.n3417 9.3005
R12725 gnd.n5471 gnd.n5470 9.3005
R12726 gnd.n3000 gnd.n2999 9.3005
R12727 gnd.n6093 gnd.n6092 9.3005
R12728 gnd.n4520 gnd.n4519 9.3005
R12729 gnd.n6089 gnd.n3001 9.3005
R12730 gnd.n6088 gnd.n6087 9.3005
R12731 gnd.n6086 gnd.n3004 9.3005
R12732 gnd.n6085 gnd.n6084 9.3005
R12733 gnd.n6083 gnd.n3005 9.3005
R12734 gnd.n6082 gnd.n6081 9.3005
R12735 gnd.n6091 gnd.n6090 9.3005
R12736 gnd.n6034 gnd.n6033 9.3005
R12737 gnd.n3052 gnd.n3051 9.3005
R12738 gnd.n6040 gnd.n6039 9.3005
R12739 gnd.n6042 gnd.n6041 9.3005
R12740 gnd.n3044 gnd.n3043 9.3005
R12741 gnd.n6048 gnd.n6047 9.3005
R12742 gnd.n6050 gnd.n6049 9.3005
R12743 gnd.n3036 gnd.n3035 9.3005
R12744 gnd.n6056 gnd.n6055 9.3005
R12745 gnd.n6058 gnd.n6057 9.3005
R12746 gnd.n3028 gnd.n3027 9.3005
R12747 gnd.n6064 gnd.n6063 9.3005
R12748 gnd.n6066 gnd.n6065 9.3005
R12749 gnd.n3020 gnd.n3019 9.3005
R12750 gnd.n6072 gnd.n6071 9.3005
R12751 gnd.n6074 gnd.n6073 9.3005
R12752 gnd.n3016 gnd.n3011 9.3005
R12753 gnd.n6032 gnd.n3061 9.3005
R12754 gnd.n3382 gnd.n3060 9.3005
R12755 gnd.n6079 gnd.n3009 9.3005
R12756 gnd.n6078 gnd.n6077 9.3005
R12757 gnd.n6076 gnd.n6075 9.3005
R12758 gnd.n3015 gnd.n3014 9.3005
R12759 gnd.n6070 gnd.n6069 9.3005
R12760 gnd.n6068 gnd.n6067 9.3005
R12761 gnd.n3024 gnd.n3023 9.3005
R12762 gnd.n6062 gnd.n6061 9.3005
R12763 gnd.n6060 gnd.n6059 9.3005
R12764 gnd.n3032 gnd.n3031 9.3005
R12765 gnd.n6054 gnd.n6053 9.3005
R12766 gnd.n6052 gnd.n6051 9.3005
R12767 gnd.n3040 gnd.n3039 9.3005
R12768 gnd.n6046 gnd.n6045 9.3005
R12769 gnd.n6044 gnd.n6043 9.3005
R12770 gnd.n3048 gnd.n3047 9.3005
R12771 gnd.n6038 gnd.n6037 9.3005
R12772 gnd.n6036 gnd.n6035 9.3005
R12773 gnd.n3405 gnd.n3058 9.3005
R12774 gnd.n3384 gnd.n3383 9.3005
R12775 gnd.n5580 gnd.n5579 9.3005
R12776 gnd.n5584 gnd.n5583 9.3005
R12777 gnd.n5585 gnd.n3379 9.3005
R12778 gnd.n5589 gnd.n5588 9.3005
R12779 gnd.n5590 gnd.n3378 9.3005
R12780 gnd.n5592 gnd.n5591 9.3005
R12781 gnd.n3376 gnd.n3375 9.3005
R12782 gnd.n5604 gnd.n5603 9.3005
R12783 gnd.n5605 gnd.n3374 9.3005
R12784 gnd.n5607 gnd.n5606 9.3005
R12785 gnd.n3372 gnd.n3371 9.3005
R12786 gnd.n5619 gnd.n5618 9.3005
R12787 gnd.n5620 gnd.n3370 9.3005
R12788 gnd.n5622 gnd.n5621 9.3005
R12789 gnd.n3367 gnd.n3366 9.3005
R12790 gnd.n5634 gnd.n5633 9.3005
R12791 gnd.n5635 gnd.n3365 9.3005
R12792 gnd.n5637 gnd.n5636 9.3005
R12793 gnd.n3363 gnd.n3362 9.3005
R12794 gnd.n5649 gnd.n5648 9.3005
R12795 gnd.n5650 gnd.n3361 9.3005
R12796 gnd.n5652 gnd.n5651 9.3005
R12797 gnd.n3358 gnd.n3357 9.3005
R12798 gnd.n5664 gnd.n5663 9.3005
R12799 gnd.n5665 gnd.n3355 9.3005
R12800 gnd.n5679 gnd.n5678 9.3005
R12801 gnd.n5677 gnd.n3356 9.3005
R12802 gnd.n5676 gnd.n5675 9.3005
R12803 gnd.n5674 gnd.n5666 9.3005
R12804 gnd.n5673 gnd.n5672 9.3005
R12805 gnd.n5671 gnd.n5670 9.3005
R12806 gnd.n5669 gnd.n95 9.3005
R12807 gnd.n5582 gnd.n3380 9.3005
R12808 gnd.n7952 gnd.n96 9.3005
R12809 gnd.n1952 gnd.t289 9.24152
R12810 gnd.n6695 gnd.t281 9.24152
R12811 gnd.n2345 gnd.t256 9.24152
R12812 gnd.n6459 gnd.t62 9.24152
R12813 gnd.n6374 gnd.t40 9.24152
R12814 gnd.n6270 gnd.n2870 9.24152
R12815 gnd.n5414 gnd.n3461 9.24152
R12816 gnd.n5631 gnd.t130 9.24152
R12817 gnd.n7903 gnd.t96 9.24152
R12818 gnd.t326 gnd.t289 8.92286
R12819 gnd.n5268 gnd.t187 8.92286
R12820 gnd.n2325 gnd.n2300 8.92171
R12821 gnd.n2293 gnd.n2268 8.92171
R12822 gnd.n2261 gnd.n2236 8.92171
R12823 gnd.n2230 gnd.n2205 8.92171
R12824 gnd.n2198 gnd.n2173 8.92171
R12825 gnd.n2166 gnd.n2141 8.92171
R12826 gnd.n2134 gnd.n2109 8.92171
R12827 gnd.n2103 gnd.n2078 8.92171
R12828 gnd.n3493 gnd.n3475 8.72777
R12829 gnd.n1874 gnd.t91 8.60421
R12830 gnd.n6483 gnd.t44 8.60421
R12831 gnd.n6350 gnd.t38 8.60421
R12832 gnd.n5601 gnd.t52 8.60421
R12833 gnd.n7879 gnd.t56 8.60421
R12834 gnd.n1292 gnd.n1272 8.43656
R12835 gnd.n54 gnd.n34 8.43656
R12836 gnd.n4961 gnd.n3727 8.28555
R12837 gnd.n5047 gnd.n5045 8.28555
R12838 gnd.n5117 gnd.n3640 8.28555
R12839 gnd.n5169 gnd.n3584 8.28555
R12840 gnd.n2326 gnd.n2298 8.14595
R12841 gnd.n2294 gnd.n2266 8.14595
R12842 gnd.n2262 gnd.n2234 8.14595
R12843 gnd.n2231 gnd.n2203 8.14595
R12844 gnd.n2199 gnd.n2171 8.14595
R12845 gnd.n2167 gnd.n2139 8.14595
R12846 gnd.n2135 gnd.n2107 8.14595
R12847 gnd.n2104 gnd.n2076 8.14595
R12848 gnd.n4284 gnd.n0 8.10675
R12849 gnd.n7953 gnd.n7952 8.10675
R12850 gnd.n2331 gnd.n2330 7.97301
R12851 gnd.t102 gnd.n1824 7.9669
R12852 gnd.n6465 gnd.n2529 7.9669
R12853 gnd.n7897 gnd.n191 7.9669
R12854 gnd.n7953 gnd.n94 7.95236
R12855 gnd.n6032 gnd.n3060 7.75808
R12856 gnd.n4602 gnd.n4594 7.75808
R12857 gnd.n7673 gnd.n7620 7.75808
R12858 gnd.n4133 gnd.n4132 7.75808
R12859 gnd.t2 gnd.n4992 7.64824
R12860 gnd.n5021 gnd.t7 7.64824
R12861 gnd.t344 gnd.n3638 7.64824
R12862 gnd.n5136 gnd.t65 7.64824
R12863 gnd.n1333 gnd.n1332 7.53171
R12864 gnd.n1757 gnd.t137 7.32958
R12865 gnd.n4201 gnd.t62 7.32958
R12866 gnd.n7588 gnd.t96 7.32958
R12867 gnd.n2892 gnd.n2891 7.30353
R12868 gnd.n3492 gnd.n3491 7.30353
R12869 gnd.n1717 gnd.n1436 7.01093
R12870 gnd.n1439 gnd.n1437 7.01093
R12871 gnd.n1727 gnd.n1726 7.01093
R12872 gnd.n1738 gnd.n1420 7.01093
R12873 gnd.n1737 gnd.n1423 7.01093
R12874 gnd.n1748 gnd.n1411 7.01093
R12875 gnd.n1414 gnd.n1412 7.01093
R12876 gnd.n1758 gnd.n1757 7.01093
R12877 gnd.n1768 gnd.n1392 7.01093
R12878 gnd.n1767 gnd.n1395 7.01093
R12879 gnd.n1784 gnd.n1385 7.01093
R12880 gnd.n1794 gnd.n1376 7.01093
R12881 gnd.n1805 gnd.n1804 7.01093
R12882 gnd.n1825 gnd.n1361 7.01093
R12883 gnd.n1824 gnd.n1340 7.01093
R12884 gnd.n1842 gnd.n1341 7.01093
R12885 gnd.n1836 gnd.n1835 7.01093
R12886 gnd.n1852 gnd.n1240 7.01093
R12887 gnd.n1861 gnd.n1231 7.01093
R12888 gnd.n1870 gnd.n1223 7.01093
R12889 gnd.n1874 gnd.n1873 7.01093
R12890 gnd.n1892 gnd.n1208 7.01093
R12891 gnd.n1891 gnd.n1211 7.01093
R12892 gnd.n1902 gnd.n1200 7.01093
R12893 gnd.n1201 gnd.n1190 7.01093
R12894 gnd.n1941 gnd.n1183 7.01093
R12895 gnd.n1940 gnd.n1939 7.01093
R12896 gnd.n1952 gnd.n1951 7.01093
R12897 gnd.n1176 gnd.n1168 7.01093
R12898 gnd.n1963 gnd.n1962 7.01093
R12899 gnd.n1981 gnd.n1156 7.01093
R12900 gnd.n1980 gnd.n1159 7.01093
R12901 gnd.n2004 gnd.n1139 7.01093
R12902 gnd.n2042 gnd.n1131 7.01093
R12903 gnd.n2041 gnd.n1123 7.01093
R12904 gnd.n2057 gnd.n2056 7.01093
R12905 gnd.n2035 gnd.n953 7.01093
R12906 gnd.n6716 gnd.n955 7.01093
R12907 gnd.n6710 gnd.n6709 7.01093
R12908 gnd.n1112 gnd.n967 7.01093
R12909 gnd.n6703 gnd.n976 7.01093
R12910 gnd.n6702 gnd.n979 7.01093
R12911 gnd.n2022 gnd.n988 7.01093
R12912 gnd.n6696 gnd.n6695 7.01093
R12913 gnd.n2346 gnd.n2345 7.01093
R12914 gnd.n6689 gnd.n1001 7.01093
R12915 gnd.n6688 gnd.n1004 7.01093
R12916 gnd.n6199 gnd.n2899 7.01093
R12917 gnd.n4970 gnd.n4969 7.01093
R12918 gnd.n4993 gnd.t2 7.01093
R12919 gnd.n4992 gnd.n4991 7.01093
R12920 gnd.n5136 gnd.n3626 7.01093
R12921 gnd.t65 gnd.n5135 7.01093
R12922 gnd.n5156 gnd.n3603 7.01093
R12923 gnd.n5406 gnd.n3467 7.01093
R12924 gnd.t235 gnd.n3471 7.01093
R12925 gnd.n1395 gnd.t362 6.69227
R12926 gnd.n1939 gnd.t326 6.69227
R12927 gnd.t363 gnd.n964 6.69227
R12928 gnd.n4219 gnd.t111 6.69227
R12929 gnd.n3945 gnd.t38 6.69227
R12930 gnd.t144 gnd.n5267 6.69227
R12931 gnd.t52 gnd.n3213 6.69227
R12932 gnd.n5755 gnd.t80 6.69227
R12933 gnd.n5334 gnd.n5333 6.5566
R12934 gnd.n3783 gnd.n3782 6.5566
R12935 gnd.n6211 gnd.n6207 6.5566
R12936 gnd.n5349 gnd.n5348 6.5566
R12937 gnd.n6717 gnd.n6716 6.37362
R12938 gnd.n5000 gnd.t15 6.37362
R12939 gnd.t312 gnd.n3619 6.37362
R12940 gnd.n5259 gnd.t190 6.37362
R12941 gnd.n4606 gnd.n4598 6.20656
R12942 gnd.n3405 gnd.n3057 6.20656
R12943 gnd.t391 gnd.n1816 6.05496
R12944 gnd.n1817 gnd.t135 6.05496
R12945 gnd.t348 gnd.n1208 6.05496
R12946 gnd.n1991 gnd.t118 6.05496
R12947 gnd.n4278 gnd.t151 6.05496
R12948 gnd.n4381 gnd.t40 6.05496
R12949 gnd.t22 gnd.t214 6.05496
R12950 gnd.t335 gnd.t14 6.05496
R12951 gnd.t94 gnd.t74 6.05496
R12952 gnd.t130 gnd.n3254 6.05496
R12953 gnd.t162 gnd.n101 6.05496
R12954 gnd.n2328 gnd.n2298 5.81868
R12955 gnd.n2296 gnd.n2266 5.81868
R12956 gnd.n2264 gnd.n2234 5.81868
R12957 gnd.n2233 gnd.n2203 5.81868
R12958 gnd.n2201 gnd.n2171 5.81868
R12959 gnd.n2169 gnd.n2139 5.81868
R12960 gnd.n2137 gnd.n2107 5.81868
R12961 gnd.n2106 gnd.n2076 5.81868
R12962 gnd.n3721 gnd.t156 5.73631
R12963 gnd.n5001 gnd.n3701 5.73631
R12964 gnd.n4984 gnd.n4983 5.73631
R12965 gnd.n5047 gnd.t7 5.73631
R12966 gnd.n3640 gnd.t344 5.73631
R12967 gnd.n5145 gnd.n5144 5.73631
R12968 gnd.n5151 gnd.n3612 5.73631
R12969 gnd.t334 gnd.n5177 5.73631
R12970 gnd.n3519 gnd.n3137 5.62001
R12971 gnd.n6273 gnd.n2835 5.62001
R12972 gnd.n6273 gnd.n2836 5.62001
R12973 gnd.n5343 gnd.n3137 5.62001
R12974 gnd.n1576 gnd.n1571 5.4308
R12975 gnd.n1105 gnd.n1035 5.4308
R12976 gnd.n1211 gnd.t101 5.41765
R12977 gnd.n1905 gnd.t386 5.41765
R12978 gnd.t140 gnd.n1138 5.41765
R12979 gnd.n4347 gnd.t3 5.41765
R12980 gnd.n3976 gnd.t108 5.41765
R12981 gnd.n4879 gnd.t340 5.41765
R12982 gnd.n5195 gnd.t146 5.41765
R12983 gnd.t0 gnd.n3295 5.41765
R12984 gnd.t34 gnd.n3314 5.41765
R12985 gnd.n3842 gnd.t204 5.09899
R12986 gnd.n4960 gnd.t345 5.09899
R12987 gnd.n5170 gnd.t314 5.09899
R12988 gnd.n2326 gnd.n2325 5.04292
R12989 gnd.n2294 gnd.n2293 5.04292
R12990 gnd.n2262 gnd.n2261 5.04292
R12991 gnd.n2231 gnd.n2230 5.04292
R12992 gnd.n2199 gnd.n2198 5.04292
R12993 gnd.n2167 gnd.n2166 5.04292
R12994 gnd.n2135 gnd.n2134 5.04292
R12995 gnd.n2104 gnd.n2103 5.04292
R12996 gnd.n1862 gnd.t385 4.78034
R12997 gnd.n1962 gnd.t90 4.78034
R12998 gnd.t58 gnd.n3995 4.78034
R12999 gnd.n4406 gnd.t16 4.78034
R13000 gnd.t10 gnd.n3272 4.78034
R13001 gnd.t20 gnd.n3331 4.78034
R13002 gnd.n1337 gnd.n1334 4.74817
R13003 gnd.n1849 gnd.n1242 4.74817
R13004 gnd.n1847 gnd.n1244 4.74817
R13005 gnd.n1253 gnd.n1251 4.74817
R13006 gnd.n1353 gnd.n1334 4.74817
R13007 gnd.n1352 gnd.n1242 4.74817
R13008 gnd.n1848 gnd.n1847 4.74817
R13009 gnd.n1253 gnd.n1252 4.74817
R13010 gnd.n3333 gnd.n114 4.74817
R13011 gnd.n5810 gnd.n113 4.74817
R13012 gnd.n3337 gnd.n112 4.74817
R13013 gnd.n7945 gnd.n107 4.74817
R13014 gnd.n7943 gnd.n108 4.74817
R13015 gnd.n5823 gnd.n114 4.74817
R13016 gnd.n3334 gnd.n113 4.74817
R13017 gnd.n5809 gnd.n112 4.74817
R13018 gnd.n3336 gnd.n107 4.74817
R13019 gnd.n7944 gnd.n7943 4.74817
R13020 gnd.n4262 gnd.n4020 4.74817
R13021 gnd.n4276 gnd.n4267 4.74817
R13022 gnd.n4274 gnd.n4273 4.74817
R13023 gnd.n4269 gnd.n4268 4.74817
R13024 gnd.n4321 gnd.n3985 4.74817
R13025 gnd.n5817 gnd.n5816 4.74817
R13026 gnd.n5707 gnd.n3325 4.74817
R13027 gnd.n5708 gnd.n5706 4.74817
R13028 gnd.n5715 gnd.n5714 4.74817
R13029 gnd.n5789 gnd.n5788 4.74817
R13030 gnd.n5818 gnd.n5817 4.74817
R13031 gnd.n5815 gnd.n3325 4.74817
R13032 gnd.n5709 gnd.n5708 4.74817
R13033 gnd.n5714 gnd.n5713 4.74817
R13034 gnd.n5790 gnd.n5789 4.74817
R13035 gnd.n2613 gnd.n2596 4.74817
R13036 gnd.n6414 gnd.n2614 4.74817
R13037 gnd.n4000 gnd.n2619 4.74817
R13038 gnd.n4307 gnd.n2618 4.74817
R13039 gnd.n2620 gnd.n2617 4.74817
R13040 gnd.n6425 gnd.n2596 4.74817
R13041 gnd.n6415 gnd.n6414 4.74817
R13042 gnd.n4236 gnd.n2619 4.74817
R13043 gnd.n4001 gnd.n2618 4.74817
R13044 gnd.n4306 gnd.n2617 4.74817
R13045 gnd.n4265 gnd.n4020 4.74817
R13046 gnd.n4267 gnd.n4266 4.74817
R13047 gnd.n4275 gnd.n4274 4.74817
R13048 gnd.n4270 gnd.n4269 4.74817
R13049 gnd.n3987 gnd.n3985 4.74817
R13050 gnd.n1332 gnd.n1331 4.74296
R13051 gnd.n94 gnd.n93 4.74296
R13052 gnd.n1292 gnd.n1291 4.7074
R13053 gnd.n1312 gnd.n1311 4.7074
R13054 gnd.n54 gnd.n53 4.7074
R13055 gnd.n74 gnd.n73 4.7074
R13056 gnd.n1332 gnd.n1312 4.65959
R13057 gnd.n94 gnd.n74 4.65959
R13058 gnd.n5974 gnd.n3139 4.6132
R13059 gnd.n6274 gnd.n2834 4.6132
R13060 gnd.n6324 gnd.n2765 4.46168
R13061 gnd.n3842 gnd.n2896 4.46168
R13062 gnd.t168 gnd.n2899 4.46168
R13063 gnd.n3745 gnd.t117 4.46168
R13064 gnd.n4976 gnd.n3715 4.46168
R13065 gnd.n5011 gnd.n3694 4.46168
R13066 gnd.n5069 gnd.n3616 4.46168
R13067 gnd.n5178 gnd.n3600 4.46168
R13068 gnd.t107 gnd.n3576 4.46168
R13069 gnd.n3471 gnd.n3460 4.46168
R13070 gnd.n6027 gnd.n3105 4.46168
R13071 gnd.n3488 gnd.n3475 4.46111
R13072 gnd.n2311 gnd.n2307 4.38594
R13073 gnd.n2279 gnd.n2275 4.38594
R13074 gnd.n2247 gnd.n2243 4.38594
R13075 gnd.n2216 gnd.n2212 4.38594
R13076 gnd.n2184 gnd.n2180 4.38594
R13077 gnd.n2152 gnd.n2148 4.38594
R13078 gnd.n2120 gnd.n2116 4.38594
R13079 gnd.n2089 gnd.n2085 4.38594
R13080 gnd.n2322 gnd.n2300 4.26717
R13081 gnd.n2290 gnd.n2268 4.26717
R13082 gnd.n2258 gnd.n2236 4.26717
R13083 gnd.n2227 gnd.n2205 4.26717
R13084 gnd.n2195 gnd.n2173 4.26717
R13085 gnd.n2163 gnd.n2141 4.26717
R13086 gnd.n2131 gnd.n2109 4.26717
R13087 gnd.n2100 gnd.n2078 4.26717
R13088 gnd.t384 gnd.n1368 4.14303
R13089 gnd.n2056 gnd.t361 4.14303
R13090 gnd.n4254 gnd.t47 4.14303
R13091 gnd.n4450 gnd.t49 4.14303
R13092 gnd.t30 gnd.n3231 4.14303
R13093 gnd.n5784 gnd.t72 4.14303
R13094 gnd.n2330 gnd.n2329 4.08274
R13095 gnd.n5333 gnd.n5332 4.05904
R13096 gnd.n3784 gnd.n3783 4.05904
R13097 gnd.n6214 gnd.n6207 4.05904
R13098 gnd.n5350 gnd.n5349 4.05904
R13099 gnd.n15 gnd.n7 3.99943
R13100 gnd.n6270 gnd.t115 3.82437
R13101 gnd.n4921 gnd.t313 3.82437
R13102 gnd.n5057 gnd.t14 3.82437
R13103 gnd.n5063 gnd.t94 3.82437
R13104 gnd.t155 gnd.n3569 3.82437
R13105 gnd.n3461 gnd.t374 3.82437
R13106 gnd.n1846 gnd.n1333 3.81325
R13107 gnd.n1312 gnd.n1292 3.72967
R13108 gnd.n74 gnd.n54 3.72967
R13109 gnd.n2330 gnd.n2202 3.70378
R13110 gnd.n15 gnd.n14 3.60163
R13111 gnd.n2478 gnd.t179 3.50571
R13112 gnd.n4190 gnd.t98 3.50571
R13113 gnd.n4760 gnd.t197 3.50571
R13114 gnd.n5898 gnd.t175 3.50571
R13115 gnd.n7595 gnd.t5 3.50571
R13116 gnd.t183 gnd.n240 3.50571
R13117 gnd.n2321 gnd.n2302 3.49141
R13118 gnd.n2289 gnd.n2270 3.49141
R13119 gnd.n2257 gnd.n2238 3.49141
R13120 gnd.n2226 gnd.n2207 3.49141
R13121 gnd.n2194 gnd.n2175 3.49141
R13122 gnd.n2162 gnd.n2143 3.49141
R13123 gnd.n2130 gnd.n2111 3.49141
R13124 gnd.n2099 gnd.n2080 3.49141
R13125 gnd.n5992 gnd.n5991 3.29747
R13126 gnd.n5991 gnd.n5990 3.29747
R13127 gnd.n7820 gnd.n7817 3.29747
R13128 gnd.n7821 gnd.n7820 3.29747
R13129 gnd.n6590 gnd.n6589 3.29747
R13130 gnd.n6589 gnd.n6588 3.29747
R13131 gnd.n6292 gnd.n6291 3.29747
R13132 gnd.n6291 gnd.n6290 3.29747
R13133 gnd.n4872 gnd.n4869 3.18706
R13134 gnd.n4947 gnd.n4946 3.18706
R13135 gnd.n5020 gnd.n3687 3.18706
R13136 gnd.n5129 gnd.n3632 3.18706
R13137 gnd.n5188 gnd.n3592 3.18706
R13138 gnd.n5251 gnd.t190 3.18706
R13139 gnd.n5274 gnd.n3546 3.18706
R13140 gnd.n1375 gnd.t384 2.8684
R13141 gnd.n1313 gnd.t305 2.82907
R13142 gnd.n1313 gnd.t353 2.82907
R13143 gnd.n1315 gnd.t148 2.82907
R13144 gnd.n1315 gnd.t307 2.82907
R13145 gnd.n1317 gnd.t378 2.82907
R13146 gnd.n1317 gnd.t29 2.82907
R13147 gnd.n1319 gnd.t78 2.82907
R13148 gnd.n1319 gnd.t306 2.82907
R13149 gnd.n1321 gnd.t152 2.82907
R13150 gnd.n1321 gnd.t316 2.82907
R13151 gnd.n1323 gnd.t290 2.82907
R13152 gnd.n1323 gnd.t308 2.82907
R13153 gnd.n1325 gnd.t379 2.82907
R13154 gnd.n1325 gnd.t350 2.82907
R13155 gnd.n1327 gnd.t393 2.82907
R13156 gnd.n1327 gnd.t388 2.82907
R13157 gnd.n1329 gnd.t25 2.82907
R13158 gnd.n1329 gnd.t76 2.82907
R13159 gnd.n1254 gnd.t355 2.82907
R13160 gnd.n1254 gnd.t50 2.82907
R13161 gnd.n1256 gnd.t17 2.82907
R13162 gnd.n1256 gnd.t132 2.82907
R13163 gnd.n1258 gnd.t122 2.82907
R13164 gnd.n1258 gnd.t51 2.82907
R13165 gnd.n1260 gnd.t294 2.82907
R13166 gnd.n1260 gnd.t32 2.82907
R13167 gnd.n1262 gnd.t351 2.82907
R13168 gnd.n1262 gnd.t382 2.82907
R13169 gnd.n1264 gnd.t371 2.82907
R13170 gnd.n1264 gnd.t352 2.82907
R13171 gnd.n1266 gnd.t9 2.82907
R13172 gnd.n1266 gnd.t112 2.82907
R13173 gnd.n1268 gnd.t158 2.82907
R13174 gnd.n1268 gnd.t399 2.82907
R13175 gnd.n1270 gnd.t129 2.82907
R13176 gnd.n1270 gnd.t82 2.82907
R13177 gnd.n1273 gnd.t104 2.82907
R13178 gnd.n1273 gnd.t337 2.82907
R13179 gnd.n1275 gnd.t134 2.82907
R13180 gnd.n1275 gnd.t41 2.82907
R13181 gnd.n1277 gnd.t109 2.82907
R13182 gnd.n1277 gnd.t92 2.82907
R13183 gnd.n1279 gnd.t370 2.82907
R13184 gnd.n1279 gnd.t324 2.82907
R13185 gnd.n1281 gnd.t161 2.82907
R13186 gnd.n1281 gnd.t95 2.82907
R13187 gnd.n1283 gnd.t48 2.82907
R13188 gnd.n1283 gnd.t124 2.82907
R13189 gnd.n1285 gnd.t61 2.82907
R13190 gnd.n1285 gnd.t380 2.82907
R13191 gnd.n1287 gnd.t63 2.82907
R13192 gnd.n1287 gnd.t157 2.82907
R13193 gnd.n1289 gnd.t121 2.82907
R13194 gnd.n1289 gnd.t19 2.82907
R13195 gnd.n1293 gnd.t373 2.82907
R13196 gnd.n1293 gnd.t85 2.82907
R13197 gnd.n1295 gnd.t321 2.82907
R13198 gnd.n1295 gnd.t395 2.82907
R13199 gnd.n1297 gnd.t346 2.82907
R13200 gnd.n1297 gnd.t125 2.82907
R13201 gnd.n1299 gnd.t93 2.82907
R13202 gnd.n1299 gnd.t4 2.82907
R13203 gnd.n1301 gnd.t309 2.82907
R13204 gnd.n1301 gnd.t59 2.82907
R13205 gnd.n1303 gnd.t301 2.82907
R13206 gnd.n1303 gnd.t342 2.82907
R13207 gnd.n1305 gnd.t357 2.82907
R13208 gnd.n1305 gnd.t295 2.82907
R13209 gnd.n1307 gnd.t302 2.82907
R13210 gnd.n1307 gnd.t99 2.82907
R13211 gnd.n1309 gnd.t300 2.82907
R13212 gnd.n1309 gnd.t66 2.82907
R13213 gnd.n91 gnd.t142 2.82907
R13214 gnd.n91 gnd.t369 2.82907
R13215 gnd.n89 gnd.t325 2.82907
R13216 gnd.n89 gnd.t299 2.82907
R13217 gnd.n87 gnd.t365 2.82907
R13218 gnd.n87 gnd.t79 2.82907
R13219 gnd.n85 gnd.t27 2.82907
R13220 gnd.n85 gnd.t315 2.82907
R13221 gnd.n83 gnd.t138 2.82907
R13222 gnd.n83 gnd.t366 2.82907
R13223 gnd.n81 gnd.t347 2.82907
R13224 gnd.n81 gnd.t291 2.82907
R13225 gnd.n79 gnd.t387 2.82907
R13226 gnd.n79 gnd.t1 2.82907
R13227 gnd.n77 gnd.t377 2.82907
R13228 gnd.n77 gnd.t60 2.82907
R13229 gnd.n75 gnd.t159 2.82907
R13230 gnd.n75 gnd.t298 2.82907
R13231 gnd.n32 gnd.t84 2.82907
R13232 gnd.n32 gnd.t83 2.82907
R13233 gnd.n30 gnd.t360 2.82907
R13234 gnd.n30 gnd.t304 2.82907
R13235 gnd.n28 gnd.t139 2.82907
R13236 gnd.n28 gnd.t70 2.82907
R13237 gnd.n26 gnd.t33 2.82907
R13238 gnd.n26 gnd.t73 2.82907
R13239 gnd.n24 gnd.t160 2.82907
R13240 gnd.n24 gnd.t323 2.82907
R13241 gnd.n22 gnd.t35 2.82907
R13242 gnd.n22 gnd.t87 2.82907
R13243 gnd.n20 gnd.t106 2.82907
R13244 gnd.n20 gnd.t320 2.82907
R13245 gnd.n18 gnd.t131 2.82907
R13246 gnd.n18 gnd.t11 2.82907
R13247 gnd.n16 gnd.t31 2.82907
R13248 gnd.n16 gnd.t68 2.82907
R13249 gnd.n51 gnd.t55 2.82907
R13250 gnd.n51 gnd.t128 2.82907
R13251 gnd.n49 gnd.t6 2.82907
R13252 gnd.n49 gnd.t97 2.82907
R13253 gnd.n47 gnd.t110 2.82907
R13254 gnd.n47 gnd.t126 2.82907
R13255 gnd.n45 gnd.t64 2.82907
R13256 gnd.n45 gnd.t100 2.82907
R13257 gnd.n43 gnd.t21 2.82907
R13258 gnd.n43 gnd.t163 2.82907
R13259 gnd.n41 gnd.t165 2.82907
R13260 gnd.n41 gnd.t296 2.82907
R13261 gnd.n39 gnd.t154 2.82907
R13262 gnd.n39 gnd.t153 2.82907
R13263 gnd.n37 gnd.t143 2.82907
R13264 gnd.n37 gnd.t164 2.82907
R13265 gnd.n35 gnd.t166 2.82907
R13266 gnd.n35 gnd.t303 2.82907
R13267 gnd.n71 gnd.t317 2.82907
R13268 gnd.n71 gnd.t43 2.82907
R13269 gnd.n69 gnd.t330 2.82907
R13270 gnd.n69 gnd.t120 2.82907
R13271 gnd.n67 gnd.t81 2.82907
R13272 gnd.n67 gnd.t343 2.82907
R13273 gnd.n65 gnd.t372 2.82907
R13274 gnd.n65 gnd.t356 2.82907
R13275 gnd.n63 gnd.t354 2.82907
R13276 gnd.n63 gnd.t383 2.82907
R13277 gnd.n61 gnd.t328 2.82907
R13278 gnd.n61 gnd.t319 2.82907
R13279 gnd.n59 gnd.t127 2.82907
R13280 gnd.n59 gnd.t381 2.82907
R13281 gnd.n57 gnd.t359 2.82907
R13282 gnd.n57 gnd.t322 2.82907
R13283 gnd.n55 gnd.t119 2.82907
R13284 gnd.n55 gnd.t329 2.82907
R13285 gnd.n2318 gnd.n2317 2.71565
R13286 gnd.n2286 gnd.n2285 2.71565
R13287 gnd.n2254 gnd.n2253 2.71565
R13288 gnd.n2223 gnd.n2222 2.71565
R13289 gnd.n2191 gnd.n2190 2.71565
R13290 gnd.n2159 gnd.n2158 2.71565
R13291 gnd.n2127 gnd.n2126 2.71565
R13292 gnd.n2096 gnd.n2095 2.71565
R13293 gnd.n1846 gnd.n1334 2.27742
R13294 gnd.n1846 gnd.n1242 2.27742
R13295 gnd.n1847 gnd.n1846 2.27742
R13296 gnd.n1846 gnd.n1253 2.27742
R13297 gnd.n7942 gnd.n114 2.27742
R13298 gnd.n7942 gnd.n113 2.27742
R13299 gnd.n7942 gnd.n112 2.27742
R13300 gnd.n7942 gnd.n107 2.27742
R13301 gnd.n7943 gnd.n7942 2.27742
R13302 gnd.n5817 gnd.n111 2.27742
R13303 gnd.n3325 gnd.n111 2.27742
R13304 gnd.n5708 gnd.n111 2.27742
R13305 gnd.n5714 gnd.n111 2.27742
R13306 gnd.n5789 gnd.n111 2.27742
R13307 gnd.n6413 gnd.n2596 2.27742
R13308 gnd.n6414 gnd.n6413 2.27742
R13309 gnd.n6413 gnd.n2619 2.27742
R13310 gnd.n6413 gnd.n2618 2.27742
R13311 gnd.n6413 gnd.n2617 2.27742
R13312 gnd.n4020 gnd.n2616 2.27742
R13313 gnd.n4267 gnd.n2616 2.27742
R13314 gnd.n4274 gnd.n2616 2.27742
R13315 gnd.n4269 gnd.n2616 2.27742
R13316 gnd.n3985 gnd.n2616 2.27742
R13317 gnd.n1726 gnd.t221 2.23109
R13318 gnd.n1851 gnd.t385 2.23109
R13319 gnd.n5011 gnd.t36 2.23109
R13320 gnd.n5039 gnd.t335 2.23109
R13321 gnd.n5111 gnd.t74 2.23109
R13322 gnd.n5069 gnd.t113 2.23109
R13323 gnd.n2314 gnd.n2304 1.93989
R13324 gnd.n2282 gnd.n2272 1.93989
R13325 gnd.n2250 gnd.n2240 1.93989
R13326 gnd.n2219 gnd.n2209 1.93989
R13327 gnd.n2187 gnd.n2177 1.93989
R13328 gnd.n2155 gnd.n2145 1.93989
R13329 gnd.n2123 gnd.n2113 1.93989
R13330 gnd.n2092 gnd.n2082 1.93989
R13331 gnd.n4900 gnd.n3765 1.91244
R13332 gnd.n4899 gnd.t285 1.91244
R13333 gnd.n4954 gnd.n3733 1.91244
R13334 gnd.n3682 gnd.n3676 1.91244
R13335 gnd.n5110 gnd.n3637 1.91244
R13336 gnd.n5220 gnd.n5219 1.91244
R13337 gnd.n5245 gnd.n3561 1.91244
R13338 gnd.t367 gnd.n1737 1.59378
R13339 gnd.n1914 gnd.t386 1.59378
R13340 gnd.n1149 gnd.t140 1.59378
R13341 gnd.t18 gnd.n2522 1.59378
R13342 gnd.n4391 gnd.t103 1.59378
R13343 gnd.n5868 gnd.t67 1.59378
R13344 gnd.n199 gnd.t54 1.59378
R13345 gnd.n4893 gnd.t193 1.27512
R13346 gnd.n5268 gnd.t217 1.27512
R13347 gnd.n1579 gnd.n1571 1.16414
R13348 gnd.n1102 gnd.n1035 1.16414
R13349 gnd.n2313 gnd.n2306 1.16414
R13350 gnd.n2281 gnd.n2274 1.16414
R13351 gnd.n2249 gnd.n2242 1.16414
R13352 gnd.n2218 gnd.n2211 1.16414
R13353 gnd.n2186 gnd.n2179 1.16414
R13354 gnd.n2154 gnd.n2147 1.16414
R13355 gnd.n2122 gnd.n2115 1.16414
R13356 gnd.n2091 gnd.n2084 1.16414
R13357 gnd.n5974 gnd.n5973 0.970197
R13358 gnd.n6274 gnd.n2832 0.970197
R13359 gnd.n2297 gnd.n2265 0.962709
R13360 gnd.n2329 gnd.n2297 0.962709
R13361 gnd.n2170 gnd.n2138 0.962709
R13362 gnd.n2202 gnd.n2170 0.962709
R13363 gnd.n1817 gnd.t391 0.956468
R13364 gnd.n1926 gnd.t118 0.956468
R13365 gnd.n4183 gnd.t8 0.956468
R13366 gnd.n4370 gnd.t28 0.956468
R13367 gnd.n4829 gnd.t396 0.956468
R13368 gnd.t374 gnd.t269 0.956468
R13369 gnd.n3448 gnd.t332 0.956468
R13370 gnd.n5844 gnd.t105 0.956468
R13371 gnd.n5765 gnd.t69 0.956468
R13372 gnd.n2 gnd.n1 0.672012
R13373 gnd.n3 gnd.n2 0.672012
R13374 gnd.n4 gnd.n3 0.672012
R13375 gnd.n5 gnd.n4 0.672012
R13376 gnd.n6 gnd.n5 0.672012
R13377 gnd.n7 gnd.n6 0.672012
R13378 gnd.n9 gnd.n8 0.672012
R13379 gnd.n10 gnd.n9 0.672012
R13380 gnd.n11 gnd.n10 0.672012
R13381 gnd.n12 gnd.n11 0.672012
R13382 gnd.n13 gnd.n12 0.672012
R13383 gnd.n14 gnd.n13 0.672012
R13384 gnd.n6193 gnd.t214 0.637812
R13385 gnd.n4912 gnd.n4911 0.637812
R13386 gnd.n4880 gnd.n4879 0.637812
R13387 gnd.n5033 gnd.n3659 0.637812
R13388 gnd.n5100 gnd.n5099 0.637812
R13389 gnd.n5195 gnd.n3579 0.637812
R13390 gnd.n5252 gnd.n3565 0.637812
R13391 gnd.n5274 gnd.t247 0.637812
R13392 gnd.n7954 gnd.n7953 0.63688
R13393 gnd gnd.n0 0.634843
R13394 gnd.n1331 gnd.n1330 0.573776
R13395 gnd.n1330 gnd.n1328 0.573776
R13396 gnd.n1328 gnd.n1326 0.573776
R13397 gnd.n1326 gnd.n1324 0.573776
R13398 gnd.n1324 gnd.n1322 0.573776
R13399 gnd.n1322 gnd.n1320 0.573776
R13400 gnd.n1320 gnd.n1318 0.573776
R13401 gnd.n1318 gnd.n1316 0.573776
R13402 gnd.n1316 gnd.n1314 0.573776
R13403 gnd.n1272 gnd.n1271 0.573776
R13404 gnd.n1271 gnd.n1269 0.573776
R13405 gnd.n1269 gnd.n1267 0.573776
R13406 gnd.n1267 gnd.n1265 0.573776
R13407 gnd.n1265 gnd.n1263 0.573776
R13408 gnd.n1263 gnd.n1261 0.573776
R13409 gnd.n1261 gnd.n1259 0.573776
R13410 gnd.n1259 gnd.n1257 0.573776
R13411 gnd.n1257 gnd.n1255 0.573776
R13412 gnd.n1291 gnd.n1290 0.573776
R13413 gnd.n1290 gnd.n1288 0.573776
R13414 gnd.n1288 gnd.n1286 0.573776
R13415 gnd.n1286 gnd.n1284 0.573776
R13416 gnd.n1284 gnd.n1282 0.573776
R13417 gnd.n1282 gnd.n1280 0.573776
R13418 gnd.n1280 gnd.n1278 0.573776
R13419 gnd.n1278 gnd.n1276 0.573776
R13420 gnd.n1276 gnd.n1274 0.573776
R13421 gnd.n1311 gnd.n1310 0.573776
R13422 gnd.n1310 gnd.n1308 0.573776
R13423 gnd.n1308 gnd.n1306 0.573776
R13424 gnd.n1306 gnd.n1304 0.573776
R13425 gnd.n1304 gnd.n1302 0.573776
R13426 gnd.n1302 gnd.n1300 0.573776
R13427 gnd.n1300 gnd.n1298 0.573776
R13428 gnd.n1298 gnd.n1296 0.573776
R13429 gnd.n1296 gnd.n1294 0.573776
R13430 gnd.n78 gnd.n76 0.573776
R13431 gnd.n80 gnd.n78 0.573776
R13432 gnd.n82 gnd.n80 0.573776
R13433 gnd.n84 gnd.n82 0.573776
R13434 gnd.n86 gnd.n84 0.573776
R13435 gnd.n88 gnd.n86 0.573776
R13436 gnd.n90 gnd.n88 0.573776
R13437 gnd.n92 gnd.n90 0.573776
R13438 gnd.n93 gnd.n92 0.573776
R13439 gnd.n19 gnd.n17 0.573776
R13440 gnd.n21 gnd.n19 0.573776
R13441 gnd.n23 gnd.n21 0.573776
R13442 gnd.n25 gnd.n23 0.573776
R13443 gnd.n27 gnd.n25 0.573776
R13444 gnd.n29 gnd.n27 0.573776
R13445 gnd.n31 gnd.n29 0.573776
R13446 gnd.n33 gnd.n31 0.573776
R13447 gnd.n34 gnd.n33 0.573776
R13448 gnd.n38 gnd.n36 0.573776
R13449 gnd.n40 gnd.n38 0.573776
R13450 gnd.n42 gnd.n40 0.573776
R13451 gnd.n44 gnd.n42 0.573776
R13452 gnd.n46 gnd.n44 0.573776
R13453 gnd.n48 gnd.n46 0.573776
R13454 gnd.n50 gnd.n48 0.573776
R13455 gnd.n52 gnd.n50 0.573776
R13456 gnd.n53 gnd.n52 0.573776
R13457 gnd.n58 gnd.n56 0.573776
R13458 gnd.n60 gnd.n58 0.573776
R13459 gnd.n62 gnd.n60 0.573776
R13460 gnd.n64 gnd.n62 0.573776
R13461 gnd.n66 gnd.n64 0.573776
R13462 gnd.n68 gnd.n66 0.573776
R13463 gnd.n70 gnd.n68 0.573776
R13464 gnd.n72 gnd.n70 0.573776
R13465 gnd.n73 gnd.n72 0.573776
R13466 gnd.n6098 gnd.n2991 0.489829
R13467 gnd.n4785 gnd.n4784 0.489829
R13468 gnd.n4519 gnd.n4483 0.489829
R13469 gnd.n6092 gnd.n6091 0.489829
R13470 gnd.n2352 gnd.n2351 0.486781
R13471 gnd.n1628 gnd.n1627 0.48678
R13472 gnd.n6634 gnd.n6633 0.480683
R13473 gnd.n1712 gnd.n1711 0.480683
R13474 gnd.n7672 gnd.n7617 0.477634
R13475 gnd.n4135 gnd.n4134 0.477634
R13476 gnd.n788 gnd.n783 0.447146
R13477 gnd.n7373 gnd.n7372 0.447146
R13478 gnd.n7585 gnd.n7584 0.447146
R13479 gnd.n4199 gnd.n4198 0.447146
R13480 gnd.n7857 gnd.n7856 0.442573
R13481 gnd.n3190 gnd.n3109 0.442573
R13482 gnd.n6328 gnd.n6327 0.442573
R13483 gnd.n2472 gnd.n2398 0.442573
R13484 gnd.n7942 gnd.n111 0.4255
R13485 gnd.n6413 gnd.n2616 0.4255
R13486 gnd.n4598 gnd.n4586 0.388379
R13487 gnd.n2310 gnd.n2309 0.388379
R13488 gnd.n2278 gnd.n2277 0.388379
R13489 gnd.n2246 gnd.n2245 0.388379
R13490 gnd.n2215 gnd.n2214 0.388379
R13491 gnd.n2183 gnd.n2182 0.388379
R13492 gnd.n2151 gnd.n2150 0.388379
R13493 gnd.n2119 gnd.n2118 0.388379
R13494 gnd.n2088 gnd.n2087 0.388379
R13495 gnd.n6036 gnd.n3057 0.388379
R13496 gnd.n7954 gnd.n15 0.374463
R13497 gnd.n2031 gnd.t363 0.319156
R13498 gnd.n4247 gnd.t123 0.319156
R13499 gnd.t77 gnd.n4317 0.319156
R13500 gnd.t193 gnd.t22 0.319156
R13501 gnd.t217 gnd.t144 0.319156
R13502 gnd.t86 gnd.n3321 0.319156
R13503 gnd.n5722 gnd.t26 0.319156
R13504 gnd.n1546 gnd.n1524 0.311721
R13505 gnd gnd.n7954 0.295112
R13506 gnd.n7733 gnd.n354 0.293183
R13507 gnd.n6506 gnd.n2462 0.293183
R13508 gnd.n6679 gnd.n1009 0.268793
R13509 gnd.n7734 gnd.n7733 0.258122
R13510 gnd.n5912 gnd.n3010 0.258122
R13511 gnd.n4754 gnd.n4753 0.258122
R13512 gnd.n6507 gnd.n6506 0.258122
R13513 gnd.n4765 gnd.n3909 0.247451
R13514 gnd.n5582 gnd.n5581 0.247451
R13515 gnd.n1049 gnd.n1009 0.241354
R13516 gnd.n3139 gnd.n3136 0.229039
R13517 gnd.n3140 gnd.n3139 0.229039
R13518 gnd.n2834 gnd.n2831 0.229039
R13519 gnd.n4678 gnd.n2834 0.229039
R13520 gnd.n1333 gnd.n0 0.210825
R13521 gnd.n1700 gnd.n1499 0.206293
R13522 gnd.n2327 gnd.n2299 0.155672
R13523 gnd.n2320 gnd.n2299 0.155672
R13524 gnd.n2320 gnd.n2319 0.155672
R13525 gnd.n2319 gnd.n2303 0.155672
R13526 gnd.n2312 gnd.n2303 0.155672
R13527 gnd.n2312 gnd.n2311 0.155672
R13528 gnd.n2295 gnd.n2267 0.155672
R13529 gnd.n2288 gnd.n2267 0.155672
R13530 gnd.n2288 gnd.n2287 0.155672
R13531 gnd.n2287 gnd.n2271 0.155672
R13532 gnd.n2280 gnd.n2271 0.155672
R13533 gnd.n2280 gnd.n2279 0.155672
R13534 gnd.n2263 gnd.n2235 0.155672
R13535 gnd.n2256 gnd.n2235 0.155672
R13536 gnd.n2256 gnd.n2255 0.155672
R13537 gnd.n2255 gnd.n2239 0.155672
R13538 gnd.n2248 gnd.n2239 0.155672
R13539 gnd.n2248 gnd.n2247 0.155672
R13540 gnd.n2232 gnd.n2204 0.155672
R13541 gnd.n2225 gnd.n2204 0.155672
R13542 gnd.n2225 gnd.n2224 0.155672
R13543 gnd.n2224 gnd.n2208 0.155672
R13544 gnd.n2217 gnd.n2208 0.155672
R13545 gnd.n2217 gnd.n2216 0.155672
R13546 gnd.n2200 gnd.n2172 0.155672
R13547 gnd.n2193 gnd.n2172 0.155672
R13548 gnd.n2193 gnd.n2192 0.155672
R13549 gnd.n2192 gnd.n2176 0.155672
R13550 gnd.n2185 gnd.n2176 0.155672
R13551 gnd.n2185 gnd.n2184 0.155672
R13552 gnd.n2168 gnd.n2140 0.155672
R13553 gnd.n2161 gnd.n2140 0.155672
R13554 gnd.n2161 gnd.n2160 0.155672
R13555 gnd.n2160 gnd.n2144 0.155672
R13556 gnd.n2153 gnd.n2144 0.155672
R13557 gnd.n2153 gnd.n2152 0.155672
R13558 gnd.n2136 gnd.n2108 0.155672
R13559 gnd.n2129 gnd.n2108 0.155672
R13560 gnd.n2129 gnd.n2128 0.155672
R13561 gnd.n2128 gnd.n2112 0.155672
R13562 gnd.n2121 gnd.n2112 0.155672
R13563 gnd.n2121 gnd.n2120 0.155672
R13564 gnd.n2105 gnd.n2077 0.155672
R13565 gnd.n2098 gnd.n2077 0.155672
R13566 gnd.n2098 gnd.n2097 0.155672
R13567 gnd.n2097 gnd.n2081 0.155672
R13568 gnd.n2090 gnd.n2081 0.155672
R13569 gnd.n2090 gnd.n2089 0.155672
R13570 gnd.n6668 gnd.n6634 0.152939
R13571 gnd.n6668 gnd.n6667 0.152939
R13572 gnd.n6667 gnd.n6666 0.152939
R13573 gnd.n6666 gnd.n6636 0.152939
R13574 gnd.n6637 gnd.n6636 0.152939
R13575 gnd.n6638 gnd.n6637 0.152939
R13576 gnd.n6639 gnd.n6638 0.152939
R13577 gnd.n6640 gnd.n6639 0.152939
R13578 gnd.n6641 gnd.n6640 0.152939
R13579 gnd.n6642 gnd.n6641 0.152939
R13580 gnd.n6643 gnd.n6642 0.152939
R13581 gnd.n6644 gnd.n6643 0.152939
R13582 gnd.n6644 gnd.n1015 0.152939
R13583 gnd.n6677 gnd.n1015 0.152939
R13584 gnd.n6678 gnd.n6677 0.152939
R13585 gnd.n6679 gnd.n6678 0.152939
R13586 gnd.n1713 gnd.n1712 0.152939
R13587 gnd.n1713 gnd.n1417 0.152939
R13588 gnd.n1741 gnd.n1417 0.152939
R13589 gnd.n1742 gnd.n1741 0.152939
R13590 gnd.n1743 gnd.n1742 0.152939
R13591 gnd.n1744 gnd.n1743 0.152939
R13592 gnd.n1744 gnd.n1389 0.152939
R13593 gnd.n1771 gnd.n1389 0.152939
R13594 gnd.n1772 gnd.n1771 0.152939
R13595 gnd.n1773 gnd.n1772 0.152939
R13596 gnd.n1774 gnd.n1773 0.152939
R13597 gnd.n1775 gnd.n1774 0.152939
R13598 gnd.n1777 gnd.n1775 0.152939
R13599 gnd.n1777 gnd.n1776 0.152939
R13600 gnd.n1776 gnd.n1357 0.152939
R13601 gnd.n1830 gnd.n1357 0.152939
R13602 gnd.n1831 gnd.n1830 0.152939
R13603 gnd.n1832 gnd.n1831 0.152939
R13604 gnd.n1832 gnd.n1226 0.152939
R13605 gnd.n1865 gnd.n1226 0.152939
R13606 gnd.n1866 gnd.n1865 0.152939
R13607 gnd.n1867 gnd.n1866 0.152939
R13608 gnd.n1867 gnd.n1205 0.152939
R13609 gnd.n1895 gnd.n1205 0.152939
R13610 gnd.n1896 gnd.n1895 0.152939
R13611 gnd.n1897 gnd.n1896 0.152939
R13612 gnd.n1898 gnd.n1897 0.152939
R13613 gnd.n1898 gnd.n1180 0.152939
R13614 gnd.n1944 gnd.n1180 0.152939
R13615 gnd.n1945 gnd.n1944 0.152939
R13616 gnd.n1946 gnd.n1945 0.152939
R13617 gnd.n1947 gnd.n1946 0.152939
R13618 gnd.n1947 gnd.n1153 0.152939
R13619 gnd.n1984 gnd.n1153 0.152939
R13620 gnd.n1985 gnd.n1984 0.152939
R13621 gnd.n1986 gnd.n1985 0.152939
R13622 gnd.n1987 gnd.n1986 0.152939
R13623 gnd.n1987 gnd.n1128 0.152939
R13624 gnd.n2045 gnd.n1128 0.152939
R13625 gnd.n2046 gnd.n2045 0.152939
R13626 gnd.n2047 gnd.n2046 0.152939
R13627 gnd.n2048 gnd.n2047 0.152939
R13628 gnd.n2050 gnd.n2048 0.152939
R13629 gnd.n2050 gnd.n2049 0.152939
R13630 gnd.n2049 gnd.n971 0.152939
R13631 gnd.n972 gnd.n971 0.152939
R13632 gnd.n973 gnd.n972 0.152939
R13633 gnd.n994 gnd.n973 0.152939
R13634 gnd.n995 gnd.n994 0.152939
R13635 gnd.n996 gnd.n995 0.152939
R13636 gnd.n997 gnd.n996 0.152939
R13637 gnd.n998 gnd.n997 0.152939
R13638 gnd.n6633 gnd.n998 0.152939
R13639 gnd.n1711 gnd.n1441 0.152939
R13640 gnd.n1462 gnd.n1441 0.152939
R13641 gnd.n1463 gnd.n1462 0.152939
R13642 gnd.n1469 gnd.n1463 0.152939
R13643 gnd.n1470 gnd.n1469 0.152939
R13644 gnd.n1471 gnd.n1470 0.152939
R13645 gnd.n1471 gnd.n1460 0.152939
R13646 gnd.n1479 gnd.n1460 0.152939
R13647 gnd.n1480 gnd.n1479 0.152939
R13648 gnd.n1481 gnd.n1480 0.152939
R13649 gnd.n1481 gnd.n1458 0.152939
R13650 gnd.n1489 gnd.n1458 0.152939
R13651 gnd.n1490 gnd.n1489 0.152939
R13652 gnd.n1491 gnd.n1490 0.152939
R13653 gnd.n1491 gnd.n1456 0.152939
R13654 gnd.n1499 gnd.n1456 0.152939
R13655 gnd.n1050 gnd.n1049 0.152939
R13656 gnd.n1051 gnd.n1050 0.152939
R13657 gnd.n1051 gnd.n1045 0.152939
R13658 gnd.n1059 gnd.n1045 0.152939
R13659 gnd.n1060 gnd.n1059 0.152939
R13660 gnd.n1061 gnd.n1060 0.152939
R13661 gnd.n1061 gnd.n1043 0.152939
R13662 gnd.n1069 gnd.n1043 0.152939
R13663 gnd.n1070 gnd.n1069 0.152939
R13664 gnd.n1071 gnd.n1070 0.152939
R13665 gnd.n1071 gnd.n1041 0.152939
R13666 gnd.n1079 gnd.n1041 0.152939
R13667 gnd.n1080 gnd.n1079 0.152939
R13668 gnd.n1081 gnd.n1080 0.152939
R13669 gnd.n1081 gnd.n1039 0.152939
R13670 gnd.n1089 gnd.n1039 0.152939
R13671 gnd.n1090 gnd.n1089 0.152939
R13672 gnd.n1091 gnd.n1090 0.152939
R13673 gnd.n1091 gnd.n1037 0.152939
R13674 gnd.n1099 gnd.n1037 0.152939
R13675 gnd.n1100 gnd.n1099 0.152939
R13676 gnd.n1101 gnd.n1100 0.152939
R13677 gnd.n1101 gnd.n1032 0.152939
R13678 gnd.n1108 gnd.n1032 0.152939
R13679 gnd.n1109 gnd.n1108 0.152939
R13680 gnd.n2352 gnd.n1109 0.152939
R13681 gnd.n1246 gnd.n1245 0.152939
R13682 gnd.n1246 gnd.n1187 0.152939
R13683 gnd.n1917 gnd.n1187 0.152939
R13684 gnd.n1918 gnd.n1917 0.152939
R13685 gnd.n1919 gnd.n1918 0.152939
R13686 gnd.n1920 gnd.n1919 0.152939
R13687 gnd.n1921 gnd.n1920 0.152939
R13688 gnd.n1922 gnd.n1921 0.152939
R13689 gnd.n1923 gnd.n1922 0.152939
R13690 gnd.n1924 gnd.n1923 0.152939
R13691 gnd.n1925 gnd.n1924 0.152939
R13692 gnd.n1925 gnd.n1135 0.152939
R13693 gnd.n2007 gnd.n1135 0.152939
R13694 gnd.n2008 gnd.n2007 0.152939
R13695 gnd.n2009 gnd.n2008 0.152939
R13696 gnd.n2010 gnd.n2009 0.152939
R13697 gnd.n2011 gnd.n2010 0.152939
R13698 gnd.n2012 gnd.n2011 0.152939
R13699 gnd.n2013 gnd.n2012 0.152939
R13700 gnd.n2014 gnd.n2013 0.152939
R13701 gnd.n2015 gnd.n2014 0.152939
R13702 gnd.n2016 gnd.n2015 0.152939
R13703 gnd.n2017 gnd.n2016 0.152939
R13704 gnd.n2018 gnd.n2017 0.152939
R13705 gnd.n2020 gnd.n2018 0.152939
R13706 gnd.n2020 gnd.n2019 0.152939
R13707 gnd.n2019 gnd.n1110 0.152939
R13708 gnd.n2351 gnd.n1110 0.152939
R13709 gnd.n1629 gnd.n1628 0.152939
R13710 gnd.n1629 gnd.n1519 0.152939
R13711 gnd.n1644 gnd.n1519 0.152939
R13712 gnd.n1645 gnd.n1644 0.152939
R13713 gnd.n1646 gnd.n1645 0.152939
R13714 gnd.n1646 gnd.n1507 0.152939
R13715 gnd.n1660 gnd.n1507 0.152939
R13716 gnd.n1661 gnd.n1660 0.152939
R13717 gnd.n1662 gnd.n1661 0.152939
R13718 gnd.n1663 gnd.n1662 0.152939
R13719 gnd.n1664 gnd.n1663 0.152939
R13720 gnd.n1665 gnd.n1664 0.152939
R13721 gnd.n1666 gnd.n1665 0.152939
R13722 gnd.n1667 gnd.n1666 0.152939
R13723 gnd.n1668 gnd.n1667 0.152939
R13724 gnd.n1669 gnd.n1668 0.152939
R13725 gnd.n1670 gnd.n1669 0.152939
R13726 gnd.n1671 gnd.n1670 0.152939
R13727 gnd.n1672 gnd.n1671 0.152939
R13728 gnd.n1673 gnd.n1672 0.152939
R13729 gnd.n1674 gnd.n1673 0.152939
R13730 gnd.n1674 gnd.n1372 0.152939
R13731 gnd.n1797 gnd.n1372 0.152939
R13732 gnd.n1798 gnd.n1797 0.152939
R13733 gnd.n1799 gnd.n1798 0.152939
R13734 gnd.n1800 gnd.n1799 0.152939
R13735 gnd.n1800 gnd.n1335 0.152939
R13736 gnd.n1845 gnd.n1335 0.152939
R13737 gnd.n1547 gnd.n1546 0.152939
R13738 gnd.n1548 gnd.n1547 0.152939
R13739 gnd.n1549 gnd.n1548 0.152939
R13740 gnd.n1550 gnd.n1549 0.152939
R13741 gnd.n1551 gnd.n1550 0.152939
R13742 gnd.n1552 gnd.n1551 0.152939
R13743 gnd.n1553 gnd.n1552 0.152939
R13744 gnd.n1554 gnd.n1553 0.152939
R13745 gnd.n1555 gnd.n1554 0.152939
R13746 gnd.n1556 gnd.n1555 0.152939
R13747 gnd.n1557 gnd.n1556 0.152939
R13748 gnd.n1558 gnd.n1557 0.152939
R13749 gnd.n1559 gnd.n1558 0.152939
R13750 gnd.n1560 gnd.n1559 0.152939
R13751 gnd.n1561 gnd.n1560 0.152939
R13752 gnd.n1562 gnd.n1561 0.152939
R13753 gnd.n1563 gnd.n1562 0.152939
R13754 gnd.n1564 gnd.n1563 0.152939
R13755 gnd.n1565 gnd.n1564 0.152939
R13756 gnd.n1566 gnd.n1565 0.152939
R13757 gnd.n1567 gnd.n1566 0.152939
R13758 gnd.n1568 gnd.n1567 0.152939
R13759 gnd.n1572 gnd.n1568 0.152939
R13760 gnd.n1573 gnd.n1572 0.152939
R13761 gnd.n1573 gnd.n1530 0.152939
R13762 gnd.n1627 gnd.n1530 0.152939
R13763 gnd.n6890 gnd.n783 0.152939
R13764 gnd.n6891 gnd.n6890 0.152939
R13765 gnd.n6892 gnd.n6891 0.152939
R13766 gnd.n6892 gnd.n777 0.152939
R13767 gnd.n6900 gnd.n777 0.152939
R13768 gnd.n6901 gnd.n6900 0.152939
R13769 gnd.n6902 gnd.n6901 0.152939
R13770 gnd.n6902 gnd.n771 0.152939
R13771 gnd.n6910 gnd.n771 0.152939
R13772 gnd.n6911 gnd.n6910 0.152939
R13773 gnd.n6912 gnd.n6911 0.152939
R13774 gnd.n6912 gnd.n765 0.152939
R13775 gnd.n6920 gnd.n765 0.152939
R13776 gnd.n6921 gnd.n6920 0.152939
R13777 gnd.n6922 gnd.n6921 0.152939
R13778 gnd.n6922 gnd.n759 0.152939
R13779 gnd.n6930 gnd.n759 0.152939
R13780 gnd.n6931 gnd.n6930 0.152939
R13781 gnd.n6932 gnd.n6931 0.152939
R13782 gnd.n6932 gnd.n753 0.152939
R13783 gnd.n6940 gnd.n753 0.152939
R13784 gnd.n6941 gnd.n6940 0.152939
R13785 gnd.n6942 gnd.n6941 0.152939
R13786 gnd.n6942 gnd.n747 0.152939
R13787 gnd.n6950 gnd.n747 0.152939
R13788 gnd.n6951 gnd.n6950 0.152939
R13789 gnd.n6952 gnd.n6951 0.152939
R13790 gnd.n6952 gnd.n741 0.152939
R13791 gnd.n6960 gnd.n741 0.152939
R13792 gnd.n6961 gnd.n6960 0.152939
R13793 gnd.n6962 gnd.n6961 0.152939
R13794 gnd.n6962 gnd.n735 0.152939
R13795 gnd.n6970 gnd.n735 0.152939
R13796 gnd.n6971 gnd.n6970 0.152939
R13797 gnd.n6972 gnd.n6971 0.152939
R13798 gnd.n6972 gnd.n729 0.152939
R13799 gnd.n6980 gnd.n729 0.152939
R13800 gnd.n6981 gnd.n6980 0.152939
R13801 gnd.n6982 gnd.n6981 0.152939
R13802 gnd.n6982 gnd.n723 0.152939
R13803 gnd.n6990 gnd.n723 0.152939
R13804 gnd.n6991 gnd.n6990 0.152939
R13805 gnd.n6992 gnd.n6991 0.152939
R13806 gnd.n6992 gnd.n717 0.152939
R13807 gnd.n7000 gnd.n717 0.152939
R13808 gnd.n7001 gnd.n7000 0.152939
R13809 gnd.n7002 gnd.n7001 0.152939
R13810 gnd.n7002 gnd.n711 0.152939
R13811 gnd.n7010 gnd.n711 0.152939
R13812 gnd.n7011 gnd.n7010 0.152939
R13813 gnd.n7012 gnd.n7011 0.152939
R13814 gnd.n7012 gnd.n705 0.152939
R13815 gnd.n7020 gnd.n705 0.152939
R13816 gnd.n7021 gnd.n7020 0.152939
R13817 gnd.n7022 gnd.n7021 0.152939
R13818 gnd.n7022 gnd.n699 0.152939
R13819 gnd.n7030 gnd.n699 0.152939
R13820 gnd.n7031 gnd.n7030 0.152939
R13821 gnd.n7032 gnd.n7031 0.152939
R13822 gnd.n7032 gnd.n693 0.152939
R13823 gnd.n7040 gnd.n693 0.152939
R13824 gnd.n7041 gnd.n7040 0.152939
R13825 gnd.n7042 gnd.n7041 0.152939
R13826 gnd.n7042 gnd.n687 0.152939
R13827 gnd.n7050 gnd.n687 0.152939
R13828 gnd.n7051 gnd.n7050 0.152939
R13829 gnd.n7052 gnd.n7051 0.152939
R13830 gnd.n7052 gnd.n681 0.152939
R13831 gnd.n7060 gnd.n681 0.152939
R13832 gnd.n7061 gnd.n7060 0.152939
R13833 gnd.n7062 gnd.n7061 0.152939
R13834 gnd.n7062 gnd.n675 0.152939
R13835 gnd.n7070 gnd.n675 0.152939
R13836 gnd.n7071 gnd.n7070 0.152939
R13837 gnd.n7072 gnd.n7071 0.152939
R13838 gnd.n7072 gnd.n669 0.152939
R13839 gnd.n7080 gnd.n669 0.152939
R13840 gnd.n7081 gnd.n7080 0.152939
R13841 gnd.n7082 gnd.n7081 0.152939
R13842 gnd.n7082 gnd.n663 0.152939
R13843 gnd.n7090 gnd.n663 0.152939
R13844 gnd.n7091 gnd.n7090 0.152939
R13845 gnd.n7092 gnd.n7091 0.152939
R13846 gnd.n7092 gnd.n657 0.152939
R13847 gnd.n7100 gnd.n657 0.152939
R13848 gnd.n7101 gnd.n7100 0.152939
R13849 gnd.n7102 gnd.n7101 0.152939
R13850 gnd.n7102 gnd.n651 0.152939
R13851 gnd.n7110 gnd.n651 0.152939
R13852 gnd.n7111 gnd.n7110 0.152939
R13853 gnd.n7112 gnd.n7111 0.152939
R13854 gnd.n7112 gnd.n645 0.152939
R13855 gnd.n7120 gnd.n645 0.152939
R13856 gnd.n7121 gnd.n7120 0.152939
R13857 gnd.n7122 gnd.n7121 0.152939
R13858 gnd.n7122 gnd.n639 0.152939
R13859 gnd.n7130 gnd.n639 0.152939
R13860 gnd.n7131 gnd.n7130 0.152939
R13861 gnd.n7132 gnd.n7131 0.152939
R13862 gnd.n7132 gnd.n633 0.152939
R13863 gnd.n7140 gnd.n633 0.152939
R13864 gnd.n7141 gnd.n7140 0.152939
R13865 gnd.n7142 gnd.n7141 0.152939
R13866 gnd.n7142 gnd.n627 0.152939
R13867 gnd.n7150 gnd.n627 0.152939
R13868 gnd.n7151 gnd.n7150 0.152939
R13869 gnd.n7152 gnd.n7151 0.152939
R13870 gnd.n7152 gnd.n621 0.152939
R13871 gnd.n7160 gnd.n621 0.152939
R13872 gnd.n7161 gnd.n7160 0.152939
R13873 gnd.n7162 gnd.n7161 0.152939
R13874 gnd.n7162 gnd.n615 0.152939
R13875 gnd.n7170 gnd.n615 0.152939
R13876 gnd.n7171 gnd.n7170 0.152939
R13877 gnd.n7172 gnd.n7171 0.152939
R13878 gnd.n7172 gnd.n609 0.152939
R13879 gnd.n7180 gnd.n609 0.152939
R13880 gnd.n7181 gnd.n7180 0.152939
R13881 gnd.n7182 gnd.n7181 0.152939
R13882 gnd.n7182 gnd.n603 0.152939
R13883 gnd.n7190 gnd.n603 0.152939
R13884 gnd.n7191 gnd.n7190 0.152939
R13885 gnd.n7192 gnd.n7191 0.152939
R13886 gnd.n7192 gnd.n597 0.152939
R13887 gnd.n7200 gnd.n597 0.152939
R13888 gnd.n7201 gnd.n7200 0.152939
R13889 gnd.n7202 gnd.n7201 0.152939
R13890 gnd.n7202 gnd.n591 0.152939
R13891 gnd.n7210 gnd.n591 0.152939
R13892 gnd.n7211 gnd.n7210 0.152939
R13893 gnd.n7212 gnd.n7211 0.152939
R13894 gnd.n7212 gnd.n585 0.152939
R13895 gnd.n7220 gnd.n585 0.152939
R13896 gnd.n7221 gnd.n7220 0.152939
R13897 gnd.n7222 gnd.n7221 0.152939
R13898 gnd.n7222 gnd.n579 0.152939
R13899 gnd.n7230 gnd.n579 0.152939
R13900 gnd.n7231 gnd.n7230 0.152939
R13901 gnd.n7232 gnd.n7231 0.152939
R13902 gnd.n7232 gnd.n573 0.152939
R13903 gnd.n7240 gnd.n573 0.152939
R13904 gnd.n7241 gnd.n7240 0.152939
R13905 gnd.n7242 gnd.n7241 0.152939
R13906 gnd.n7242 gnd.n567 0.152939
R13907 gnd.n7250 gnd.n567 0.152939
R13908 gnd.n7251 gnd.n7250 0.152939
R13909 gnd.n7252 gnd.n7251 0.152939
R13910 gnd.n7252 gnd.n561 0.152939
R13911 gnd.n7260 gnd.n561 0.152939
R13912 gnd.n7261 gnd.n7260 0.152939
R13913 gnd.n7262 gnd.n7261 0.152939
R13914 gnd.n7262 gnd.n555 0.152939
R13915 gnd.n7270 gnd.n555 0.152939
R13916 gnd.n7271 gnd.n7270 0.152939
R13917 gnd.n7272 gnd.n7271 0.152939
R13918 gnd.n7272 gnd.n549 0.152939
R13919 gnd.n7280 gnd.n549 0.152939
R13920 gnd.n7281 gnd.n7280 0.152939
R13921 gnd.n7282 gnd.n7281 0.152939
R13922 gnd.n7282 gnd.n543 0.152939
R13923 gnd.n7290 gnd.n543 0.152939
R13924 gnd.n7291 gnd.n7290 0.152939
R13925 gnd.n7292 gnd.n7291 0.152939
R13926 gnd.n7292 gnd.n537 0.152939
R13927 gnd.n7300 gnd.n537 0.152939
R13928 gnd.n7301 gnd.n7300 0.152939
R13929 gnd.n7302 gnd.n7301 0.152939
R13930 gnd.n7302 gnd.n531 0.152939
R13931 gnd.n7310 gnd.n531 0.152939
R13932 gnd.n7311 gnd.n7310 0.152939
R13933 gnd.n7312 gnd.n7311 0.152939
R13934 gnd.n7312 gnd.n525 0.152939
R13935 gnd.n7320 gnd.n525 0.152939
R13936 gnd.n7321 gnd.n7320 0.152939
R13937 gnd.n7322 gnd.n7321 0.152939
R13938 gnd.n7322 gnd.n519 0.152939
R13939 gnd.n7330 gnd.n519 0.152939
R13940 gnd.n7331 gnd.n7330 0.152939
R13941 gnd.n7332 gnd.n7331 0.152939
R13942 gnd.n7332 gnd.n513 0.152939
R13943 gnd.n7340 gnd.n513 0.152939
R13944 gnd.n7341 gnd.n7340 0.152939
R13945 gnd.n7342 gnd.n7341 0.152939
R13946 gnd.n7342 gnd.n507 0.152939
R13947 gnd.n7350 gnd.n507 0.152939
R13948 gnd.n7351 gnd.n7350 0.152939
R13949 gnd.n7352 gnd.n7351 0.152939
R13950 gnd.n7352 gnd.n501 0.152939
R13951 gnd.n7360 gnd.n501 0.152939
R13952 gnd.n7361 gnd.n7360 0.152939
R13953 gnd.n7363 gnd.n7361 0.152939
R13954 gnd.n7363 gnd.n7362 0.152939
R13955 gnd.n7362 gnd.n495 0.152939
R13956 gnd.n7372 gnd.n495 0.152939
R13957 gnd.n7373 gnd.n490 0.152939
R13958 gnd.n7381 gnd.n490 0.152939
R13959 gnd.n7382 gnd.n7381 0.152939
R13960 gnd.n7383 gnd.n7382 0.152939
R13961 gnd.n7383 gnd.n484 0.152939
R13962 gnd.n7391 gnd.n484 0.152939
R13963 gnd.n7392 gnd.n7391 0.152939
R13964 gnd.n7393 gnd.n7392 0.152939
R13965 gnd.n7393 gnd.n478 0.152939
R13966 gnd.n7401 gnd.n478 0.152939
R13967 gnd.n7402 gnd.n7401 0.152939
R13968 gnd.n7403 gnd.n7402 0.152939
R13969 gnd.n7403 gnd.n472 0.152939
R13970 gnd.n7411 gnd.n472 0.152939
R13971 gnd.n7412 gnd.n7411 0.152939
R13972 gnd.n7413 gnd.n7412 0.152939
R13973 gnd.n7413 gnd.n466 0.152939
R13974 gnd.n7421 gnd.n466 0.152939
R13975 gnd.n7422 gnd.n7421 0.152939
R13976 gnd.n7423 gnd.n7422 0.152939
R13977 gnd.n7423 gnd.n460 0.152939
R13978 gnd.n7431 gnd.n460 0.152939
R13979 gnd.n7432 gnd.n7431 0.152939
R13980 gnd.n7433 gnd.n7432 0.152939
R13981 gnd.n7433 gnd.n454 0.152939
R13982 gnd.n7441 gnd.n454 0.152939
R13983 gnd.n7442 gnd.n7441 0.152939
R13984 gnd.n7443 gnd.n7442 0.152939
R13985 gnd.n7443 gnd.n448 0.152939
R13986 gnd.n7451 gnd.n448 0.152939
R13987 gnd.n7452 gnd.n7451 0.152939
R13988 gnd.n7453 gnd.n7452 0.152939
R13989 gnd.n7453 gnd.n442 0.152939
R13990 gnd.n7461 gnd.n442 0.152939
R13991 gnd.n7462 gnd.n7461 0.152939
R13992 gnd.n7463 gnd.n7462 0.152939
R13993 gnd.n7463 gnd.n436 0.152939
R13994 gnd.n7471 gnd.n436 0.152939
R13995 gnd.n7472 gnd.n7471 0.152939
R13996 gnd.n7473 gnd.n7472 0.152939
R13997 gnd.n7473 gnd.n430 0.152939
R13998 gnd.n7481 gnd.n430 0.152939
R13999 gnd.n7482 gnd.n7481 0.152939
R14000 gnd.n7483 gnd.n7482 0.152939
R14001 gnd.n7483 gnd.n424 0.152939
R14002 gnd.n7491 gnd.n424 0.152939
R14003 gnd.n7492 gnd.n7491 0.152939
R14004 gnd.n7493 gnd.n7492 0.152939
R14005 gnd.n7493 gnd.n418 0.152939
R14006 gnd.n7501 gnd.n418 0.152939
R14007 gnd.n7502 gnd.n7501 0.152939
R14008 gnd.n7503 gnd.n7502 0.152939
R14009 gnd.n7503 gnd.n412 0.152939
R14010 gnd.n7511 gnd.n412 0.152939
R14011 gnd.n7512 gnd.n7511 0.152939
R14012 gnd.n7513 gnd.n7512 0.152939
R14013 gnd.n7513 gnd.n406 0.152939
R14014 gnd.n7521 gnd.n406 0.152939
R14015 gnd.n7522 gnd.n7521 0.152939
R14016 gnd.n7523 gnd.n7522 0.152939
R14017 gnd.n7523 gnd.n400 0.152939
R14018 gnd.n7531 gnd.n400 0.152939
R14019 gnd.n7532 gnd.n7531 0.152939
R14020 gnd.n7533 gnd.n7532 0.152939
R14021 gnd.n7533 gnd.n394 0.152939
R14022 gnd.n7541 gnd.n394 0.152939
R14023 gnd.n7542 gnd.n7541 0.152939
R14024 gnd.n7543 gnd.n7542 0.152939
R14025 gnd.n7543 gnd.n388 0.152939
R14026 gnd.n7551 gnd.n388 0.152939
R14027 gnd.n7552 gnd.n7551 0.152939
R14028 gnd.n7553 gnd.n7552 0.152939
R14029 gnd.n7553 gnd.n382 0.152939
R14030 gnd.n7561 gnd.n382 0.152939
R14031 gnd.n7562 gnd.n7561 0.152939
R14032 gnd.n7563 gnd.n7562 0.152939
R14033 gnd.n7563 gnd.n376 0.152939
R14034 gnd.n7571 gnd.n376 0.152939
R14035 gnd.n7572 gnd.n7571 0.152939
R14036 gnd.n7573 gnd.n7572 0.152939
R14037 gnd.n7573 gnd.n370 0.152939
R14038 gnd.n7582 gnd.n370 0.152939
R14039 gnd.n7583 gnd.n7582 0.152939
R14040 gnd.n7585 gnd.n7583 0.152939
R14041 gnd.n5739 gnd.n5716 0.152939
R14042 gnd.n5741 gnd.n5739 0.152939
R14043 gnd.n5742 gnd.n5741 0.152939
R14044 gnd.n5743 gnd.n5742 0.152939
R14045 gnd.n5744 gnd.n5743 0.152939
R14046 gnd.n5745 gnd.n5744 0.152939
R14047 gnd.n5747 gnd.n5745 0.152939
R14048 gnd.n5747 gnd.n5746 0.152939
R14049 gnd.n5746 gnd.n364 0.152939
R14050 gnd.n365 gnd.n364 0.152939
R14051 gnd.n366 gnd.n365 0.152939
R14052 gnd.n7584 gnd.n366 0.152939
R14053 gnd.n7942 gnd.n109 0.152939
R14054 gnd.n134 gnd.n109 0.152939
R14055 gnd.n135 gnd.n134 0.152939
R14056 gnd.n136 gnd.n135 0.152939
R14057 gnd.n153 gnd.n136 0.152939
R14058 gnd.n154 gnd.n153 0.152939
R14059 gnd.n155 gnd.n154 0.152939
R14060 gnd.n156 gnd.n155 0.152939
R14061 gnd.n173 gnd.n156 0.152939
R14062 gnd.n174 gnd.n173 0.152939
R14063 gnd.n175 gnd.n174 0.152939
R14064 gnd.n176 gnd.n175 0.152939
R14065 gnd.n193 gnd.n176 0.152939
R14066 gnd.n194 gnd.n193 0.152939
R14067 gnd.n195 gnd.n194 0.152939
R14068 gnd.n196 gnd.n195 0.152939
R14069 gnd.n213 gnd.n196 0.152939
R14070 gnd.n214 gnd.n213 0.152939
R14071 gnd.n215 gnd.n214 0.152939
R14072 gnd.n216 gnd.n215 0.152939
R14073 gnd.n232 gnd.n216 0.152939
R14074 gnd.n233 gnd.n232 0.152939
R14075 gnd.n234 gnd.n233 0.152939
R14076 gnd.n235 gnd.n234 0.152939
R14077 gnd.n251 gnd.n235 0.152939
R14078 gnd.n252 gnd.n251 0.152939
R14079 gnd.n7857 gnd.n252 0.152939
R14080 gnd.n7951 gnd.n97 0.152939
R14081 gnd.n5721 gnd.n97 0.152939
R14082 gnd.n5725 gnd.n5721 0.152939
R14083 gnd.n5726 gnd.n5725 0.152939
R14084 gnd.n5727 gnd.n5726 0.152939
R14085 gnd.n5728 gnd.n5727 0.152939
R14086 gnd.n5729 gnd.n5728 0.152939
R14087 gnd.n5756 gnd.n5729 0.152939
R14088 gnd.n5757 gnd.n5756 0.152939
R14089 gnd.n5758 gnd.n5757 0.152939
R14090 gnd.n5759 gnd.n5758 0.152939
R14091 gnd.n5759 gnd.n358 0.152939
R14092 gnd.n7599 gnd.n358 0.152939
R14093 gnd.n7600 gnd.n7599 0.152939
R14094 gnd.n7601 gnd.n7600 0.152939
R14095 gnd.n7602 gnd.n7601 0.152939
R14096 gnd.n7603 gnd.n7602 0.152939
R14097 gnd.n7604 gnd.n7603 0.152939
R14098 gnd.n7605 gnd.n7604 0.152939
R14099 gnd.n7606 gnd.n7605 0.152939
R14100 gnd.n7607 gnd.n7606 0.152939
R14101 gnd.n7608 gnd.n7607 0.152939
R14102 gnd.n7609 gnd.n7608 0.152939
R14103 gnd.n7610 gnd.n7609 0.152939
R14104 gnd.n7611 gnd.n7610 0.152939
R14105 gnd.n7612 gnd.n7611 0.152939
R14106 gnd.n7613 gnd.n7612 0.152939
R14107 gnd.n7614 gnd.n7613 0.152939
R14108 gnd.n7615 gnd.n7614 0.152939
R14109 gnd.n7616 gnd.n7615 0.152939
R14110 gnd.n7617 gnd.n7616 0.152939
R14111 gnd.n7631 gnd.n354 0.152939
R14112 gnd.n7632 gnd.n7631 0.152939
R14113 gnd.n7632 gnd.n7627 0.152939
R14114 gnd.n7640 gnd.n7627 0.152939
R14115 gnd.n7641 gnd.n7640 0.152939
R14116 gnd.n7642 gnd.n7641 0.152939
R14117 gnd.n7642 gnd.n7625 0.152939
R14118 gnd.n7650 gnd.n7625 0.152939
R14119 gnd.n7651 gnd.n7650 0.152939
R14120 gnd.n7652 gnd.n7651 0.152939
R14121 gnd.n7652 gnd.n7623 0.152939
R14122 gnd.n7660 gnd.n7623 0.152939
R14123 gnd.n7661 gnd.n7660 0.152939
R14124 gnd.n7662 gnd.n7661 0.152939
R14125 gnd.n7662 gnd.n7621 0.152939
R14126 gnd.n7670 gnd.n7621 0.152939
R14127 gnd.n7671 gnd.n7670 0.152939
R14128 gnd.n7672 gnd.n7671 0.152939
R14129 gnd.n7856 gnd.n253 0.152939
R14130 gnd.n296 gnd.n253 0.152939
R14131 gnd.n297 gnd.n296 0.152939
R14132 gnd.n298 gnd.n297 0.152939
R14133 gnd.n299 gnd.n298 0.152939
R14134 gnd.n300 gnd.n299 0.152939
R14135 gnd.n301 gnd.n300 0.152939
R14136 gnd.n302 gnd.n301 0.152939
R14137 gnd.n303 gnd.n302 0.152939
R14138 gnd.n304 gnd.n303 0.152939
R14139 gnd.n305 gnd.n304 0.152939
R14140 gnd.n306 gnd.n305 0.152939
R14141 gnd.n307 gnd.n306 0.152939
R14142 gnd.n308 gnd.n307 0.152939
R14143 gnd.n309 gnd.n308 0.152939
R14144 gnd.n310 gnd.n309 0.152939
R14145 gnd.n311 gnd.n310 0.152939
R14146 gnd.n312 gnd.n311 0.152939
R14147 gnd.n313 gnd.n312 0.152939
R14148 gnd.n314 gnd.n313 0.152939
R14149 gnd.n315 gnd.n314 0.152939
R14150 gnd.n316 gnd.n315 0.152939
R14151 gnd.n317 gnd.n316 0.152939
R14152 gnd.n318 gnd.n317 0.152939
R14153 gnd.n319 gnd.n318 0.152939
R14154 gnd.n320 gnd.n319 0.152939
R14155 gnd.n321 gnd.n320 0.152939
R14156 gnd.n322 gnd.n321 0.152939
R14157 gnd.n323 gnd.n322 0.152939
R14158 gnd.n324 gnd.n323 0.152939
R14159 gnd.n325 gnd.n324 0.152939
R14160 gnd.n326 gnd.n325 0.152939
R14161 gnd.n327 gnd.n326 0.152939
R14162 gnd.n328 gnd.n327 0.152939
R14163 gnd.n329 gnd.n328 0.152939
R14164 gnd.n330 gnd.n329 0.152939
R14165 gnd.n7777 gnd.n330 0.152939
R14166 gnd.n7777 gnd.n7776 0.152939
R14167 gnd.n7776 gnd.n7775 0.152939
R14168 gnd.n7775 gnd.n334 0.152939
R14169 gnd.n335 gnd.n334 0.152939
R14170 gnd.n336 gnd.n335 0.152939
R14171 gnd.n337 gnd.n336 0.152939
R14172 gnd.n338 gnd.n337 0.152939
R14173 gnd.n339 gnd.n338 0.152939
R14174 gnd.n340 gnd.n339 0.152939
R14175 gnd.n341 gnd.n340 0.152939
R14176 gnd.n342 gnd.n341 0.152939
R14177 gnd.n343 gnd.n342 0.152939
R14178 gnd.n344 gnd.n343 0.152939
R14179 gnd.n345 gnd.n344 0.152939
R14180 gnd.n346 gnd.n345 0.152939
R14181 gnd.n347 gnd.n346 0.152939
R14182 gnd.n348 gnd.n347 0.152939
R14183 gnd.n349 gnd.n348 0.152939
R14184 gnd.n350 gnd.n349 0.152939
R14185 gnd.n7735 gnd.n350 0.152939
R14186 gnd.n7735 gnd.n7734 0.152939
R14187 gnd.n3110 gnd.n3109 0.152939
R14188 gnd.n3111 gnd.n3110 0.152939
R14189 gnd.n3112 gnd.n3111 0.152939
R14190 gnd.n3113 gnd.n3112 0.152939
R14191 gnd.n3114 gnd.n3113 0.152939
R14192 gnd.n3115 gnd.n3114 0.152939
R14193 gnd.n3116 gnd.n3115 0.152939
R14194 gnd.n3117 gnd.n3116 0.152939
R14195 gnd.n3118 gnd.n3117 0.152939
R14196 gnd.n3119 gnd.n3118 0.152939
R14197 gnd.n3120 gnd.n3119 0.152939
R14198 gnd.n3121 gnd.n3120 0.152939
R14199 gnd.n3122 gnd.n3121 0.152939
R14200 gnd.n3123 gnd.n3122 0.152939
R14201 gnd.n3124 gnd.n3123 0.152939
R14202 gnd.n3125 gnd.n3124 0.152939
R14203 gnd.n3126 gnd.n3125 0.152939
R14204 gnd.n3129 gnd.n3126 0.152939
R14205 gnd.n3130 gnd.n3129 0.152939
R14206 gnd.n3131 gnd.n3130 0.152939
R14207 gnd.n3132 gnd.n3131 0.152939
R14208 gnd.n3133 gnd.n3132 0.152939
R14209 gnd.n3134 gnd.n3133 0.152939
R14210 gnd.n3135 gnd.n3134 0.152939
R14211 gnd.n3136 gnd.n3135 0.152939
R14212 gnd.n3141 gnd.n3140 0.152939
R14213 gnd.n3142 gnd.n3141 0.152939
R14214 gnd.n3143 gnd.n3142 0.152939
R14215 gnd.n3144 gnd.n3143 0.152939
R14216 gnd.n3145 gnd.n3144 0.152939
R14217 gnd.n3146 gnd.n3145 0.152939
R14218 gnd.n3147 gnd.n3146 0.152939
R14219 gnd.n3148 gnd.n3147 0.152939
R14220 gnd.n3149 gnd.n3148 0.152939
R14221 gnd.n3152 gnd.n3149 0.152939
R14222 gnd.n3153 gnd.n3152 0.152939
R14223 gnd.n3154 gnd.n3153 0.152939
R14224 gnd.n3155 gnd.n3154 0.152939
R14225 gnd.n3156 gnd.n3155 0.152939
R14226 gnd.n3157 gnd.n3156 0.152939
R14227 gnd.n3158 gnd.n3157 0.152939
R14228 gnd.n3159 gnd.n3158 0.152939
R14229 gnd.n3160 gnd.n3159 0.152939
R14230 gnd.n3161 gnd.n3160 0.152939
R14231 gnd.n3162 gnd.n3161 0.152939
R14232 gnd.n3163 gnd.n3162 0.152939
R14233 gnd.n3164 gnd.n3163 0.152939
R14234 gnd.n3165 gnd.n3164 0.152939
R14235 gnd.n3166 gnd.n3165 0.152939
R14236 gnd.n3167 gnd.n3166 0.152939
R14237 gnd.n3168 gnd.n3167 0.152939
R14238 gnd.n3169 gnd.n3168 0.152939
R14239 gnd.n3170 gnd.n3169 0.152939
R14240 gnd.n5913 gnd.n3170 0.152939
R14241 gnd.n5913 gnd.n5912 0.152939
R14242 gnd.n3191 gnd.n3190 0.152939
R14243 gnd.n3192 gnd.n3191 0.152939
R14244 gnd.n3193 gnd.n3192 0.152939
R14245 gnd.n3194 gnd.n3193 0.152939
R14246 gnd.n3215 gnd.n3194 0.152939
R14247 gnd.n3216 gnd.n3215 0.152939
R14248 gnd.n3217 gnd.n3216 0.152939
R14249 gnd.n3218 gnd.n3217 0.152939
R14250 gnd.n3236 gnd.n3218 0.152939
R14251 gnd.n3237 gnd.n3236 0.152939
R14252 gnd.n3238 gnd.n3237 0.152939
R14253 gnd.n3239 gnd.n3238 0.152939
R14254 gnd.n3256 gnd.n3239 0.152939
R14255 gnd.n3257 gnd.n3256 0.152939
R14256 gnd.n3258 gnd.n3257 0.152939
R14257 gnd.n3259 gnd.n3258 0.152939
R14258 gnd.n3277 gnd.n3259 0.152939
R14259 gnd.n3278 gnd.n3277 0.152939
R14260 gnd.n3279 gnd.n3278 0.152939
R14261 gnd.n3280 gnd.n3279 0.152939
R14262 gnd.n3297 gnd.n3280 0.152939
R14263 gnd.n3298 gnd.n3297 0.152939
R14264 gnd.n3299 gnd.n3298 0.152939
R14265 gnd.n3300 gnd.n3299 0.152939
R14266 gnd.n3301 gnd.n3300 0.152939
R14267 gnd.n3301 gnd.n110 0.152939
R14268 gnd.n7942 gnd.n110 0.152939
R14269 gnd.n4324 gnd.n4323 0.152939
R14270 gnd.n4325 gnd.n4324 0.152939
R14271 gnd.n4326 gnd.n4325 0.152939
R14272 gnd.n4329 gnd.n4326 0.152939
R14273 gnd.n4330 gnd.n4329 0.152939
R14274 gnd.n4331 gnd.n4330 0.152939
R14275 gnd.n4332 gnd.n4331 0.152939
R14276 gnd.n4334 gnd.n4332 0.152939
R14277 gnd.n4334 gnd.n4333 0.152939
R14278 gnd.n4333 gnd.n3959 0.152939
R14279 gnd.n4411 gnd.n3959 0.152939
R14280 gnd.n4412 gnd.n4411 0.152939
R14281 gnd.n4413 gnd.n4412 0.152939
R14282 gnd.n4413 gnd.n3955 0.152939
R14283 gnd.n4419 gnd.n3955 0.152939
R14284 gnd.n4420 gnd.n4419 0.152939
R14285 gnd.n4421 gnd.n4420 0.152939
R14286 gnd.n4422 gnd.n4421 0.152939
R14287 gnd.n4423 gnd.n4422 0.152939
R14288 gnd.n4426 gnd.n4423 0.152939
R14289 gnd.n4427 gnd.n4426 0.152939
R14290 gnd.n4428 gnd.n4427 0.152939
R14291 gnd.n4429 gnd.n4428 0.152939
R14292 gnd.n4431 gnd.n4429 0.152939
R14293 gnd.n4432 gnd.n4431 0.152939
R14294 gnd.n4434 gnd.n4432 0.152939
R14295 gnd.n4434 gnd.n4433 0.152939
R14296 gnd.n4433 gnd.n3931 0.152939
R14297 gnd.n4774 gnd.n3931 0.152939
R14298 gnd.n4775 gnd.n4774 0.152939
R14299 gnd.n4776 gnd.n4775 0.152939
R14300 gnd.n4777 gnd.n4776 0.152939
R14301 gnd.n4777 gnd.n3902 0.152939
R14302 gnd.n4792 gnd.n3902 0.152939
R14303 gnd.n4793 gnd.n4792 0.152939
R14304 gnd.n4794 gnd.n4793 0.152939
R14305 gnd.n4794 gnd.n3887 0.152939
R14306 gnd.n4808 gnd.n3887 0.152939
R14307 gnd.n4809 gnd.n4808 0.152939
R14308 gnd.n4810 gnd.n4809 0.152939
R14309 gnd.n4810 gnd.n3873 0.152939
R14310 gnd.n4824 gnd.n3873 0.152939
R14311 gnd.n4825 gnd.n4824 0.152939
R14312 gnd.n4826 gnd.n4825 0.152939
R14313 gnd.n4826 gnd.n3858 0.152939
R14314 gnd.n4851 gnd.n3858 0.152939
R14315 gnd.n4852 gnd.n4851 0.152939
R14316 gnd.n4853 gnd.n4852 0.152939
R14317 gnd.n4855 gnd.n4853 0.152939
R14318 gnd.n4855 gnd.n4854 0.152939
R14319 gnd.n4854 gnd.n2904 0.152939
R14320 gnd.n2905 gnd.n2904 0.152939
R14321 gnd.n2906 gnd.n2905 0.152939
R14322 gnd.n3767 gnd.n2906 0.152939
R14323 gnd.n3768 gnd.n3767 0.152939
R14324 gnd.n3768 gnd.n3748 0.152939
R14325 gnd.n4925 gnd.n3748 0.152939
R14326 gnd.n4926 gnd.n4925 0.152939
R14327 gnd.n4927 gnd.n4926 0.152939
R14328 gnd.n4927 gnd.n3724 0.152939
R14329 gnd.n4964 gnd.n3724 0.152939
R14330 gnd.n4965 gnd.n4964 0.152939
R14331 gnd.n4966 gnd.n4965 0.152939
R14332 gnd.n4966 gnd.n3698 0.152939
R14333 gnd.n5004 gnd.n3698 0.152939
R14334 gnd.n5005 gnd.n5004 0.152939
R14335 gnd.n5006 gnd.n5005 0.152939
R14336 gnd.n5007 gnd.n5006 0.152939
R14337 gnd.n5007 gnd.n3671 0.152939
R14338 gnd.n5050 gnd.n3671 0.152939
R14339 gnd.n5051 gnd.n5050 0.152939
R14340 gnd.n5052 gnd.n5051 0.152939
R14341 gnd.n5053 gnd.n5052 0.152939
R14342 gnd.n5053 gnd.n3649 0.152939
R14343 gnd.n5103 gnd.n3649 0.152939
R14344 gnd.n5104 gnd.n5103 0.152939
R14345 gnd.n5105 gnd.n5104 0.152939
R14346 gnd.n5106 gnd.n5105 0.152939
R14347 gnd.n5106 gnd.n3623 0.152939
R14348 gnd.n5139 gnd.n3623 0.152939
R14349 gnd.n5140 gnd.n5139 0.152939
R14350 gnd.n5141 gnd.n5140 0.152939
R14351 gnd.n5141 gnd.n3597 0.152939
R14352 gnd.n5181 gnd.n3597 0.152939
R14353 gnd.n5182 gnd.n5181 0.152939
R14354 gnd.n5183 gnd.n5182 0.152939
R14355 gnd.n5184 gnd.n5183 0.152939
R14356 gnd.n5184 gnd.n3573 0.152939
R14357 gnd.n5233 gnd.n3573 0.152939
R14358 gnd.n5234 gnd.n5233 0.152939
R14359 gnd.n5235 gnd.n5234 0.152939
R14360 gnd.n5235 gnd.n3555 0.152939
R14361 gnd.n5262 gnd.n3555 0.152939
R14362 gnd.n5263 gnd.n5262 0.152939
R14363 gnd.n5264 gnd.n5263 0.152939
R14364 gnd.n5264 gnd.n3464 0.152939
R14365 gnd.n5409 gnd.n3464 0.152939
R14366 gnd.n5410 gnd.n5409 0.152939
R14367 gnd.n5411 gnd.n5410 0.152939
R14368 gnd.n5411 gnd.n3451 0.152939
R14369 gnd.n5425 gnd.n3451 0.152939
R14370 gnd.n5426 gnd.n5425 0.152939
R14371 gnd.n5427 gnd.n5426 0.152939
R14372 gnd.n5427 gnd.n3438 0.152939
R14373 gnd.n5441 gnd.n3438 0.152939
R14374 gnd.n5442 gnd.n5441 0.152939
R14375 gnd.n5443 gnd.n5442 0.152939
R14376 gnd.n5443 gnd.n3425 0.152939
R14377 gnd.n5457 gnd.n3425 0.152939
R14378 gnd.n5458 gnd.n5457 0.152939
R14379 gnd.n5459 gnd.n5458 0.152939
R14380 gnd.n5461 gnd.n5459 0.152939
R14381 gnd.n5461 gnd.n5460 0.152939
R14382 gnd.n5460 gnd.n3412 0.152939
R14383 gnd.n5478 gnd.n3412 0.152939
R14384 gnd.n5479 gnd.n5478 0.152939
R14385 gnd.n5480 gnd.n5479 0.152939
R14386 gnd.n5481 gnd.n5480 0.152939
R14387 gnd.n5482 gnd.n5481 0.152939
R14388 gnd.n5485 gnd.n5482 0.152939
R14389 gnd.n5486 gnd.n5485 0.152939
R14390 gnd.n5487 gnd.n5486 0.152939
R14391 gnd.n5488 gnd.n5487 0.152939
R14392 gnd.n5491 gnd.n5488 0.152939
R14393 gnd.n5492 gnd.n5491 0.152939
R14394 gnd.n5493 gnd.n5492 0.152939
R14395 gnd.n5494 gnd.n5493 0.152939
R14396 gnd.n5497 gnd.n5494 0.152939
R14397 gnd.n5498 gnd.n5497 0.152939
R14398 gnd.n5499 gnd.n5498 0.152939
R14399 gnd.n5500 gnd.n5499 0.152939
R14400 gnd.n5503 gnd.n5500 0.152939
R14401 gnd.n5504 gnd.n5503 0.152939
R14402 gnd.n5505 gnd.n5504 0.152939
R14403 gnd.n5506 gnd.n5505 0.152939
R14404 gnd.n5509 gnd.n5506 0.152939
R14405 gnd.n5510 gnd.n5509 0.152939
R14406 gnd.n5511 gnd.n5510 0.152939
R14407 gnd.n5512 gnd.n5511 0.152939
R14408 gnd.n5515 gnd.n5512 0.152939
R14409 gnd.n5516 gnd.n5515 0.152939
R14410 gnd.n5517 gnd.n5516 0.152939
R14411 gnd.n5518 gnd.n5517 0.152939
R14412 gnd.n5521 gnd.n5518 0.152939
R14413 gnd.n5522 gnd.n5521 0.152939
R14414 gnd.n5523 gnd.n5522 0.152939
R14415 gnd.n5525 gnd.n5523 0.152939
R14416 gnd.n5525 gnd.n5524 0.152939
R14417 gnd.n4135 gnd.n4076 0.152939
R14418 gnd.n4141 gnd.n4076 0.152939
R14419 gnd.n4142 gnd.n4141 0.152939
R14420 gnd.n4143 gnd.n4142 0.152939
R14421 gnd.n4143 gnd.n4074 0.152939
R14422 gnd.n4149 gnd.n4074 0.152939
R14423 gnd.n4150 gnd.n4149 0.152939
R14424 gnd.n4151 gnd.n4150 0.152939
R14425 gnd.n4151 gnd.n4072 0.152939
R14426 gnd.n4157 gnd.n4072 0.152939
R14427 gnd.n4158 gnd.n4157 0.152939
R14428 gnd.n4159 gnd.n4158 0.152939
R14429 gnd.n4159 gnd.n4070 0.152939
R14430 gnd.n4165 gnd.n4070 0.152939
R14431 gnd.n4166 gnd.n4165 0.152939
R14432 gnd.n4168 gnd.n4166 0.152939
R14433 gnd.n4168 gnd.n4167 0.152939
R14434 gnd.n4167 gnd.n4042 0.152939
R14435 gnd.n4043 gnd.n4042 0.152939
R14436 gnd.n4044 gnd.n4043 0.152939
R14437 gnd.n4044 gnd.n4033 0.152939
R14438 gnd.n4223 gnd.n4033 0.152939
R14439 gnd.n4224 gnd.n4223 0.152939
R14440 gnd.n4226 gnd.n4224 0.152939
R14441 gnd.n4226 gnd.n4225 0.152939
R14442 gnd.n4225 gnd.n4028 0.152939
R14443 gnd.n4029 gnd.n4028 0.152939
R14444 gnd.n4030 gnd.n4029 0.152939
R14445 gnd.n4030 gnd.n4015 0.152939
R14446 gnd.n4282 gnd.n4015 0.152939
R14447 gnd.n4283 gnd.n4282 0.152939
R14448 gnd.n4090 gnd.n2462 0.152939
R14449 gnd.n4098 gnd.n4090 0.152939
R14450 gnd.n4099 gnd.n4098 0.152939
R14451 gnd.n4100 gnd.n4099 0.152939
R14452 gnd.n4100 gnd.n4088 0.152939
R14453 gnd.n4108 gnd.n4088 0.152939
R14454 gnd.n4109 gnd.n4108 0.152939
R14455 gnd.n4110 gnd.n4109 0.152939
R14456 gnd.n4110 gnd.n4086 0.152939
R14457 gnd.n4118 gnd.n4086 0.152939
R14458 gnd.n4119 gnd.n4118 0.152939
R14459 gnd.n4120 gnd.n4119 0.152939
R14460 gnd.n4120 gnd.n4084 0.152939
R14461 gnd.n4128 gnd.n4084 0.152939
R14462 gnd.n4129 gnd.n4128 0.152939
R14463 gnd.n4130 gnd.n4129 0.152939
R14464 gnd.n4130 gnd.n4077 0.152939
R14465 gnd.n4134 gnd.n4077 0.152939
R14466 gnd.n6413 gnd.n2615 0.152939
R14467 gnd.n2640 gnd.n2615 0.152939
R14468 gnd.n2641 gnd.n2640 0.152939
R14469 gnd.n2642 gnd.n2641 0.152939
R14470 gnd.n2659 gnd.n2642 0.152939
R14471 gnd.n2660 gnd.n2659 0.152939
R14472 gnd.n2661 gnd.n2660 0.152939
R14473 gnd.n2662 gnd.n2661 0.152939
R14474 gnd.n2679 gnd.n2662 0.152939
R14475 gnd.n2680 gnd.n2679 0.152939
R14476 gnd.n2681 gnd.n2680 0.152939
R14477 gnd.n2682 gnd.n2681 0.152939
R14478 gnd.n2699 gnd.n2682 0.152939
R14479 gnd.n2700 gnd.n2699 0.152939
R14480 gnd.n2701 gnd.n2700 0.152939
R14481 gnd.n2702 gnd.n2701 0.152939
R14482 gnd.n2719 gnd.n2702 0.152939
R14483 gnd.n2720 gnd.n2719 0.152939
R14484 gnd.n2721 gnd.n2720 0.152939
R14485 gnd.n2722 gnd.n2721 0.152939
R14486 gnd.n2739 gnd.n2722 0.152939
R14487 gnd.n2740 gnd.n2739 0.152939
R14488 gnd.n2741 gnd.n2740 0.152939
R14489 gnd.n2742 gnd.n2741 0.152939
R14490 gnd.n2760 gnd.n2742 0.152939
R14491 gnd.n2761 gnd.n2760 0.152939
R14492 gnd.n6328 gnd.n2761 0.152939
R14493 gnd.n6327 gnd.n2762 0.152939
R14494 gnd.n2806 gnd.n2762 0.152939
R14495 gnd.n2807 gnd.n2806 0.152939
R14496 gnd.n2808 gnd.n2807 0.152939
R14497 gnd.n2809 gnd.n2808 0.152939
R14498 gnd.n2810 gnd.n2809 0.152939
R14499 gnd.n2811 gnd.n2810 0.152939
R14500 gnd.n2812 gnd.n2811 0.152939
R14501 gnd.n2813 gnd.n2812 0.152939
R14502 gnd.n2814 gnd.n2813 0.152939
R14503 gnd.n2815 gnd.n2814 0.152939
R14504 gnd.n2816 gnd.n2815 0.152939
R14505 gnd.n2817 gnd.n2816 0.152939
R14506 gnd.n2818 gnd.n2817 0.152939
R14507 gnd.n2819 gnd.n2818 0.152939
R14508 gnd.n2820 gnd.n2819 0.152939
R14509 gnd.n2821 gnd.n2820 0.152939
R14510 gnd.n2824 gnd.n2821 0.152939
R14511 gnd.n2825 gnd.n2824 0.152939
R14512 gnd.n2826 gnd.n2825 0.152939
R14513 gnd.n2827 gnd.n2826 0.152939
R14514 gnd.n2828 gnd.n2827 0.152939
R14515 gnd.n2829 gnd.n2828 0.152939
R14516 gnd.n2830 gnd.n2829 0.152939
R14517 gnd.n2831 gnd.n2830 0.152939
R14518 gnd.n4679 gnd.n4678 0.152939
R14519 gnd.n4686 gnd.n4679 0.152939
R14520 gnd.n4687 gnd.n4686 0.152939
R14521 gnd.n4688 gnd.n4687 0.152939
R14522 gnd.n4688 gnd.n4676 0.152939
R14523 gnd.n4696 gnd.n4676 0.152939
R14524 gnd.n4697 gnd.n4696 0.152939
R14525 gnd.n4698 gnd.n4697 0.152939
R14526 gnd.n4698 gnd.n4671 0.152939
R14527 gnd.n4705 gnd.n4671 0.152939
R14528 gnd.n4706 gnd.n4705 0.152939
R14529 gnd.n4707 gnd.n4706 0.152939
R14530 gnd.n4707 gnd.n4669 0.152939
R14531 gnd.n4715 gnd.n4669 0.152939
R14532 gnd.n4716 gnd.n4715 0.152939
R14533 gnd.n4717 gnd.n4716 0.152939
R14534 gnd.n4717 gnd.n4667 0.152939
R14535 gnd.n4725 gnd.n4667 0.152939
R14536 gnd.n4726 gnd.n4725 0.152939
R14537 gnd.n4727 gnd.n4726 0.152939
R14538 gnd.n4727 gnd.n4665 0.152939
R14539 gnd.n4735 gnd.n4665 0.152939
R14540 gnd.n4736 gnd.n4735 0.152939
R14541 gnd.n4737 gnd.n4736 0.152939
R14542 gnd.n4737 gnd.n4663 0.152939
R14543 gnd.n4745 gnd.n4663 0.152939
R14544 gnd.n4746 gnd.n4745 0.152939
R14545 gnd.n4747 gnd.n4746 0.152939
R14546 gnd.n4747 gnd.n4658 0.152939
R14547 gnd.n4753 gnd.n4658 0.152939
R14548 gnd.n2399 gnd.n2398 0.152939
R14549 gnd.n2400 gnd.n2399 0.152939
R14550 gnd.n2401 gnd.n2400 0.152939
R14551 gnd.n2402 gnd.n2401 0.152939
R14552 gnd.n2403 gnd.n2402 0.152939
R14553 gnd.n2404 gnd.n2403 0.152939
R14554 gnd.n2405 gnd.n2404 0.152939
R14555 gnd.n2406 gnd.n2405 0.152939
R14556 gnd.n2407 gnd.n2406 0.152939
R14557 gnd.n2408 gnd.n2407 0.152939
R14558 gnd.n2409 gnd.n2408 0.152939
R14559 gnd.n2410 gnd.n2409 0.152939
R14560 gnd.n2411 gnd.n2410 0.152939
R14561 gnd.n2412 gnd.n2411 0.152939
R14562 gnd.n2413 gnd.n2412 0.152939
R14563 gnd.n2414 gnd.n2413 0.152939
R14564 gnd.n2415 gnd.n2414 0.152939
R14565 gnd.n2418 gnd.n2415 0.152939
R14566 gnd.n2419 gnd.n2418 0.152939
R14567 gnd.n2420 gnd.n2419 0.152939
R14568 gnd.n2421 gnd.n2420 0.152939
R14569 gnd.n2422 gnd.n2421 0.152939
R14570 gnd.n2423 gnd.n2422 0.152939
R14571 gnd.n2424 gnd.n2423 0.152939
R14572 gnd.n2425 gnd.n2424 0.152939
R14573 gnd.n2426 gnd.n2425 0.152939
R14574 gnd.n2427 gnd.n2426 0.152939
R14575 gnd.n2428 gnd.n2427 0.152939
R14576 gnd.n2429 gnd.n2428 0.152939
R14577 gnd.n2430 gnd.n2429 0.152939
R14578 gnd.n2431 gnd.n2430 0.152939
R14579 gnd.n2432 gnd.n2431 0.152939
R14580 gnd.n2433 gnd.n2432 0.152939
R14581 gnd.n2434 gnd.n2433 0.152939
R14582 gnd.n2435 gnd.n2434 0.152939
R14583 gnd.n2436 gnd.n2435 0.152939
R14584 gnd.n2437 gnd.n2436 0.152939
R14585 gnd.n2440 gnd.n2437 0.152939
R14586 gnd.n2441 gnd.n2440 0.152939
R14587 gnd.n2442 gnd.n2441 0.152939
R14588 gnd.n2443 gnd.n2442 0.152939
R14589 gnd.n2444 gnd.n2443 0.152939
R14590 gnd.n2445 gnd.n2444 0.152939
R14591 gnd.n2446 gnd.n2445 0.152939
R14592 gnd.n2447 gnd.n2446 0.152939
R14593 gnd.n2448 gnd.n2447 0.152939
R14594 gnd.n2449 gnd.n2448 0.152939
R14595 gnd.n2450 gnd.n2449 0.152939
R14596 gnd.n2451 gnd.n2450 0.152939
R14597 gnd.n2452 gnd.n2451 0.152939
R14598 gnd.n2453 gnd.n2452 0.152939
R14599 gnd.n2454 gnd.n2453 0.152939
R14600 gnd.n2455 gnd.n2454 0.152939
R14601 gnd.n2456 gnd.n2455 0.152939
R14602 gnd.n2457 gnd.n2456 0.152939
R14603 gnd.n2458 gnd.n2457 0.152939
R14604 gnd.n6508 gnd.n2458 0.152939
R14605 gnd.n6508 gnd.n6507 0.152939
R14606 gnd.n2473 gnd.n2472 0.152939
R14607 gnd.n2474 gnd.n2473 0.152939
R14608 gnd.n2475 gnd.n2474 0.152939
R14609 gnd.n2495 gnd.n2475 0.152939
R14610 gnd.n2496 gnd.n2495 0.152939
R14611 gnd.n2497 gnd.n2496 0.152939
R14612 gnd.n2498 gnd.n2497 0.152939
R14613 gnd.n2513 gnd.n2498 0.152939
R14614 gnd.n2514 gnd.n2513 0.152939
R14615 gnd.n2515 gnd.n2514 0.152939
R14616 gnd.n2516 gnd.n2515 0.152939
R14617 gnd.n2534 gnd.n2516 0.152939
R14618 gnd.n2535 gnd.n2534 0.152939
R14619 gnd.n2536 gnd.n2535 0.152939
R14620 gnd.n2537 gnd.n2536 0.152939
R14621 gnd.n2553 gnd.n2537 0.152939
R14622 gnd.n2554 gnd.n2553 0.152939
R14623 gnd.n2555 gnd.n2554 0.152939
R14624 gnd.n2556 gnd.n2555 0.152939
R14625 gnd.n2574 gnd.n2556 0.152939
R14626 gnd.n2575 gnd.n2574 0.152939
R14627 gnd.n2576 gnd.n2575 0.152939
R14628 gnd.n2577 gnd.n2576 0.152939
R14629 gnd.n2593 gnd.n2577 0.152939
R14630 gnd.n2594 gnd.n2593 0.152939
R14631 gnd.n2595 gnd.n2594 0.152939
R14632 gnd.n6413 gnd.n2595 0.152939
R14633 gnd.n4199 gnd.n4193 0.152939
R14634 gnd.n4206 gnd.n4193 0.152939
R14635 gnd.n4207 gnd.n4206 0.152939
R14636 gnd.n4208 gnd.n4207 0.152939
R14637 gnd.n4208 gnd.n4038 0.152939
R14638 gnd.n4214 gnd.n4038 0.152939
R14639 gnd.n4215 gnd.n4214 0.152939
R14640 gnd.n4216 gnd.n4215 0.152939
R14641 gnd.n4216 gnd.n4023 0.152939
R14642 gnd.n4258 gnd.n4023 0.152939
R14643 gnd.n4259 gnd.n4258 0.152939
R14644 gnd.n4260 gnd.n4259 0.152939
R14645 gnd.n789 gnd.n788 0.152939
R14646 gnd.n790 gnd.n789 0.152939
R14647 gnd.n795 gnd.n790 0.152939
R14648 gnd.n796 gnd.n795 0.152939
R14649 gnd.n797 gnd.n796 0.152939
R14650 gnd.n798 gnd.n797 0.152939
R14651 gnd.n803 gnd.n798 0.152939
R14652 gnd.n804 gnd.n803 0.152939
R14653 gnd.n805 gnd.n804 0.152939
R14654 gnd.n806 gnd.n805 0.152939
R14655 gnd.n811 gnd.n806 0.152939
R14656 gnd.n812 gnd.n811 0.152939
R14657 gnd.n813 gnd.n812 0.152939
R14658 gnd.n814 gnd.n813 0.152939
R14659 gnd.n819 gnd.n814 0.152939
R14660 gnd.n820 gnd.n819 0.152939
R14661 gnd.n821 gnd.n820 0.152939
R14662 gnd.n822 gnd.n821 0.152939
R14663 gnd.n827 gnd.n822 0.152939
R14664 gnd.n828 gnd.n827 0.152939
R14665 gnd.n829 gnd.n828 0.152939
R14666 gnd.n830 gnd.n829 0.152939
R14667 gnd.n835 gnd.n830 0.152939
R14668 gnd.n836 gnd.n835 0.152939
R14669 gnd.n837 gnd.n836 0.152939
R14670 gnd.n838 gnd.n837 0.152939
R14671 gnd.n843 gnd.n838 0.152939
R14672 gnd.n844 gnd.n843 0.152939
R14673 gnd.n845 gnd.n844 0.152939
R14674 gnd.n846 gnd.n845 0.152939
R14675 gnd.n851 gnd.n846 0.152939
R14676 gnd.n852 gnd.n851 0.152939
R14677 gnd.n853 gnd.n852 0.152939
R14678 gnd.n854 gnd.n853 0.152939
R14679 gnd.n859 gnd.n854 0.152939
R14680 gnd.n860 gnd.n859 0.152939
R14681 gnd.n861 gnd.n860 0.152939
R14682 gnd.n862 gnd.n861 0.152939
R14683 gnd.n867 gnd.n862 0.152939
R14684 gnd.n868 gnd.n867 0.152939
R14685 gnd.n869 gnd.n868 0.152939
R14686 gnd.n870 gnd.n869 0.152939
R14687 gnd.n875 gnd.n870 0.152939
R14688 gnd.n876 gnd.n875 0.152939
R14689 gnd.n877 gnd.n876 0.152939
R14690 gnd.n878 gnd.n877 0.152939
R14691 gnd.n883 gnd.n878 0.152939
R14692 gnd.n884 gnd.n883 0.152939
R14693 gnd.n885 gnd.n884 0.152939
R14694 gnd.n886 gnd.n885 0.152939
R14695 gnd.n891 gnd.n886 0.152939
R14696 gnd.n892 gnd.n891 0.152939
R14697 gnd.n893 gnd.n892 0.152939
R14698 gnd.n894 gnd.n893 0.152939
R14699 gnd.n899 gnd.n894 0.152939
R14700 gnd.n900 gnd.n899 0.152939
R14701 gnd.n901 gnd.n900 0.152939
R14702 gnd.n902 gnd.n901 0.152939
R14703 gnd.n907 gnd.n902 0.152939
R14704 gnd.n908 gnd.n907 0.152939
R14705 gnd.n909 gnd.n908 0.152939
R14706 gnd.n910 gnd.n909 0.152939
R14707 gnd.n915 gnd.n910 0.152939
R14708 gnd.n916 gnd.n915 0.152939
R14709 gnd.n917 gnd.n916 0.152939
R14710 gnd.n918 gnd.n917 0.152939
R14711 gnd.n923 gnd.n918 0.152939
R14712 gnd.n924 gnd.n923 0.152939
R14713 gnd.n925 gnd.n924 0.152939
R14714 gnd.n926 gnd.n925 0.152939
R14715 gnd.n931 gnd.n926 0.152939
R14716 gnd.n932 gnd.n931 0.152939
R14717 gnd.n933 gnd.n932 0.152939
R14718 gnd.n934 gnd.n933 0.152939
R14719 gnd.n939 gnd.n934 0.152939
R14720 gnd.n940 gnd.n939 0.152939
R14721 gnd.n941 gnd.n940 0.152939
R14722 gnd.n942 gnd.n941 0.152939
R14723 gnd.n947 gnd.n942 0.152939
R14724 gnd.n948 gnd.n947 0.152939
R14725 gnd.n949 gnd.n948 0.152939
R14726 gnd.n950 gnd.n949 0.152939
R14727 gnd.n4196 gnd.n950 0.152939
R14728 gnd.n4198 gnd.n4196 0.152939
R14729 gnd.n4786 gnd.n4785 0.152939
R14730 gnd.n4786 gnd.n3895 0.152939
R14731 gnd.n4800 gnd.n3895 0.152939
R14732 gnd.n4801 gnd.n4800 0.152939
R14733 gnd.n4802 gnd.n4801 0.152939
R14734 gnd.n4802 gnd.n3881 0.152939
R14735 gnd.n4816 gnd.n3881 0.152939
R14736 gnd.n4817 gnd.n4816 0.152939
R14737 gnd.n4818 gnd.n4817 0.152939
R14738 gnd.n4818 gnd.n3867 0.152939
R14739 gnd.n4832 gnd.n3867 0.152939
R14740 gnd.n4833 gnd.n4832 0.152939
R14741 gnd.n4845 gnd.n4833 0.152939
R14742 gnd.n4845 gnd.n4844 0.152939
R14743 gnd.n4844 gnd.n4843 0.152939
R14744 gnd.n4843 gnd.n4834 0.152939
R14745 gnd.n4839 gnd.n4834 0.152939
R14746 gnd.n4839 gnd.n4838 0.152939
R14747 gnd.n4838 gnd.n2915 0.152939
R14748 gnd.n6190 gnd.n2915 0.152939
R14749 gnd.n6190 gnd.n6189 0.152939
R14750 gnd.n6189 gnd.n6188 0.152939
R14751 gnd.n6188 gnd.n2916 0.152939
R14752 gnd.n6184 gnd.n2916 0.152939
R14753 gnd.n6184 gnd.n6183 0.152939
R14754 gnd.n6183 gnd.n6182 0.152939
R14755 gnd.n6182 gnd.n2921 0.152939
R14756 gnd.n6178 gnd.n2921 0.152939
R14757 gnd.n6178 gnd.n6177 0.152939
R14758 gnd.n6177 gnd.n6176 0.152939
R14759 gnd.n6176 gnd.n2926 0.152939
R14760 gnd.n6172 gnd.n2926 0.152939
R14761 gnd.n6172 gnd.n6171 0.152939
R14762 gnd.n6171 gnd.n6170 0.152939
R14763 gnd.n6170 gnd.n2931 0.152939
R14764 gnd.n6166 gnd.n2931 0.152939
R14765 gnd.n6166 gnd.n6165 0.152939
R14766 gnd.n6165 gnd.n6164 0.152939
R14767 gnd.n6164 gnd.n2936 0.152939
R14768 gnd.n6160 gnd.n2936 0.152939
R14769 gnd.n6160 gnd.n6159 0.152939
R14770 gnd.n6159 gnd.n6158 0.152939
R14771 gnd.n6158 gnd.n2941 0.152939
R14772 gnd.n6154 gnd.n2941 0.152939
R14773 gnd.n6154 gnd.n6153 0.152939
R14774 gnd.n6153 gnd.n6152 0.152939
R14775 gnd.n6152 gnd.n2946 0.152939
R14776 gnd.n6148 gnd.n2946 0.152939
R14777 gnd.n6148 gnd.n6147 0.152939
R14778 gnd.n6147 gnd.n6146 0.152939
R14779 gnd.n6146 gnd.n2951 0.152939
R14780 gnd.n6142 gnd.n2951 0.152939
R14781 gnd.n6142 gnd.n6141 0.152939
R14782 gnd.n6141 gnd.n6140 0.152939
R14783 gnd.n6140 gnd.n2956 0.152939
R14784 gnd.n6136 gnd.n2956 0.152939
R14785 gnd.n6136 gnd.n6135 0.152939
R14786 gnd.n6135 gnd.n6134 0.152939
R14787 gnd.n6134 gnd.n2961 0.152939
R14788 gnd.n6130 gnd.n2961 0.152939
R14789 gnd.n6130 gnd.n6129 0.152939
R14790 gnd.n6129 gnd.n6128 0.152939
R14791 gnd.n6128 gnd.n2966 0.152939
R14792 gnd.n6124 gnd.n2966 0.152939
R14793 gnd.n6124 gnd.n6123 0.152939
R14794 gnd.n6123 gnd.n6122 0.152939
R14795 gnd.n6122 gnd.n2971 0.152939
R14796 gnd.n6118 gnd.n2971 0.152939
R14797 gnd.n6118 gnd.n6117 0.152939
R14798 gnd.n6117 gnd.n6116 0.152939
R14799 gnd.n6116 gnd.n2976 0.152939
R14800 gnd.n6112 gnd.n2976 0.152939
R14801 gnd.n6112 gnd.n6111 0.152939
R14802 gnd.n6111 gnd.n6110 0.152939
R14803 gnd.n6110 gnd.n2981 0.152939
R14804 gnd.n6106 gnd.n2981 0.152939
R14805 gnd.n6106 gnd.n6105 0.152939
R14806 gnd.n6105 gnd.n6104 0.152939
R14807 gnd.n6104 gnd.n2986 0.152939
R14808 gnd.n6100 gnd.n2986 0.152939
R14809 gnd.n6100 gnd.n6099 0.152939
R14810 gnd.n6099 gnd.n6098 0.152939
R14811 gnd.n4312 gnd.n3992 0.152939
R14812 gnd.n4313 gnd.n4312 0.152939
R14813 gnd.n4314 gnd.n4313 0.152939
R14814 gnd.n4314 gnd.n3980 0.152939
R14815 gnd.n4351 gnd.n3980 0.152939
R14816 gnd.n4352 gnd.n4351 0.152939
R14817 gnd.n4353 gnd.n4352 0.152939
R14818 gnd.n4353 gnd.n3974 0.152939
R14819 gnd.n4365 gnd.n3974 0.152939
R14820 gnd.n4366 gnd.n4365 0.152939
R14821 gnd.n4367 gnd.n4366 0.152939
R14822 gnd.n4367 gnd.n3966 0.152939
R14823 gnd.n4402 gnd.n3966 0.152939
R14824 gnd.n4402 gnd.n4401 0.152939
R14825 gnd.n4401 gnd.n4400 0.152939
R14826 gnd.n4400 gnd.n3967 0.152939
R14827 gnd.n4396 gnd.n3967 0.152939
R14828 gnd.n4396 gnd.n4395 0.152939
R14829 gnd.n4395 gnd.n4394 0.152939
R14830 gnd.n4394 gnd.n3949 0.152939
R14831 gnd.n4454 gnd.n3949 0.152939
R14832 gnd.n4455 gnd.n4454 0.152939
R14833 gnd.n4456 gnd.n4455 0.152939
R14834 gnd.n4456 gnd.n3943 0.152939
R14835 gnd.n4468 gnd.n3943 0.152939
R14836 gnd.n4469 gnd.n4468 0.152939
R14837 gnd.n4470 gnd.n4469 0.152939
R14838 gnd.n4470 gnd.n3938 0.152939
R14839 gnd.n4763 gnd.n3938 0.152939
R14840 gnd.n4764 gnd.n4763 0.152939
R14841 gnd.n4765 gnd.n4764 0.152939
R14842 gnd.n4483 gnd.n4482 0.152939
R14843 gnd.n4528 gnd.n4482 0.152939
R14844 gnd.n4529 gnd.n4528 0.152939
R14845 gnd.n4530 gnd.n4529 0.152939
R14846 gnd.n4530 gnd.n4478 0.152939
R14847 gnd.n4656 gnd.n4478 0.152939
R14848 gnd.n4519 gnd.n4518 0.152939
R14849 gnd.n4518 gnd.n4517 0.152939
R14850 gnd.n4517 gnd.n4485 0.152939
R14851 gnd.n4513 gnd.n4485 0.152939
R14852 gnd.n4513 gnd.n4512 0.152939
R14853 gnd.n4512 gnd.n4511 0.152939
R14854 gnd.n4511 gnd.n4489 0.152939
R14855 gnd.n4507 gnd.n4489 0.152939
R14856 gnd.n4507 gnd.n4506 0.152939
R14857 gnd.n4506 gnd.n4505 0.152939
R14858 gnd.n4505 gnd.n4493 0.152939
R14859 gnd.n4501 gnd.n4493 0.152939
R14860 gnd.n4501 gnd.n4500 0.152939
R14861 gnd.n4500 gnd.n4499 0.152939
R14862 gnd.n4499 gnd.n4497 0.152939
R14863 gnd.n4497 gnd.n3849 0.152939
R14864 gnd.n4864 gnd.n3849 0.152939
R14865 gnd.n4865 gnd.n4864 0.152939
R14866 gnd.n4866 gnd.n4865 0.152939
R14867 gnd.n4866 gnd.n3763 0.152939
R14868 gnd.n4903 gnd.n3763 0.152939
R14869 gnd.n4904 gnd.n4903 0.152939
R14870 gnd.n4908 gnd.n4904 0.152939
R14871 gnd.n4908 gnd.n4907 0.152939
R14872 gnd.n4907 gnd.n4906 0.152939
R14873 gnd.n4906 gnd.n3741 0.152939
R14874 gnd.n4934 gnd.n3741 0.152939
R14875 gnd.n4935 gnd.n4934 0.152939
R14876 gnd.n4942 gnd.n4935 0.152939
R14877 gnd.n4942 gnd.n4941 0.152939
R14878 gnd.n4941 gnd.n4940 0.152939
R14879 gnd.n4940 gnd.n4936 0.152939
R14880 gnd.n4936 gnd.n3691 0.152939
R14881 gnd.n5014 gnd.n3691 0.152939
R14882 gnd.n5015 gnd.n5014 0.152939
R14883 gnd.n5017 gnd.n5015 0.152939
R14884 gnd.n5017 gnd.n5016 0.152939
R14885 gnd.n5016 gnd.n3664 0.152939
R14886 gnd.n5060 gnd.n3664 0.152939
R14887 gnd.n5061 gnd.n5060 0.152939
R14888 gnd.n5088 gnd.n5061 0.152939
R14889 gnd.n5088 gnd.n5087 0.152939
R14890 gnd.n5087 gnd.n5086 0.152939
R14891 gnd.n5086 gnd.n5062 0.152939
R14892 gnd.n5082 gnd.n5062 0.152939
R14893 gnd.n5082 gnd.n5081 0.152939
R14894 gnd.n5081 gnd.n5080 0.152939
R14895 gnd.n5080 gnd.n5068 0.152939
R14896 gnd.n5076 gnd.n5068 0.152939
R14897 gnd.n5076 gnd.n5075 0.152939
R14898 gnd.n5075 gnd.n5074 0.152939
R14899 gnd.n5074 gnd.n3589 0.152939
R14900 gnd.n5191 gnd.n3589 0.152939
R14901 gnd.n5192 gnd.n5191 0.152939
R14902 gnd.n5216 gnd.n5192 0.152939
R14903 gnd.n5216 gnd.n5215 0.152939
R14904 gnd.n5215 gnd.n5214 0.152939
R14905 gnd.n5214 gnd.n5193 0.152939
R14906 gnd.n5210 gnd.n5193 0.152939
R14907 gnd.n5210 gnd.n5209 0.152939
R14908 gnd.n5209 gnd.n5208 0.152939
R14909 gnd.n5208 gnd.n5199 0.152939
R14910 gnd.n5204 gnd.n5199 0.152939
R14911 gnd.n5204 gnd.n5203 0.152939
R14912 gnd.n5203 gnd.n3457 0.152939
R14913 gnd.n5417 gnd.n3457 0.152939
R14914 gnd.n5418 gnd.n5417 0.152939
R14915 gnd.n5419 gnd.n5418 0.152939
R14916 gnd.n5419 gnd.n3443 0.152939
R14917 gnd.n5433 gnd.n3443 0.152939
R14918 gnd.n5434 gnd.n5433 0.152939
R14919 gnd.n5435 gnd.n5434 0.152939
R14920 gnd.n5435 gnd.n3430 0.152939
R14921 gnd.n5449 gnd.n3430 0.152939
R14922 gnd.n5450 gnd.n5449 0.152939
R14923 gnd.n5451 gnd.n5450 0.152939
R14924 gnd.n5451 gnd.n3418 0.152939
R14925 gnd.n5468 gnd.n3418 0.152939
R14926 gnd.n5469 gnd.n5468 0.152939
R14927 gnd.n5470 gnd.n5469 0.152939
R14928 gnd.n5470 gnd.n3000 0.152939
R14929 gnd.n6092 gnd.n3000 0.152939
R14930 gnd.n6091 gnd.n3001 0.152939
R14931 gnd.n6087 gnd.n3001 0.152939
R14932 gnd.n6087 gnd.n6086 0.152939
R14933 gnd.n6086 gnd.n6085 0.152939
R14934 gnd.n6085 gnd.n3005 0.152939
R14935 gnd.n6081 gnd.n3005 0.152939
R14936 gnd.n5583 gnd.n5582 0.152939
R14937 gnd.n5583 gnd.n3379 0.152939
R14938 gnd.n5589 gnd.n3379 0.152939
R14939 gnd.n5590 gnd.n5589 0.152939
R14940 gnd.n5591 gnd.n5590 0.152939
R14941 gnd.n5591 gnd.n3375 0.152939
R14942 gnd.n5604 gnd.n3375 0.152939
R14943 gnd.n5605 gnd.n5604 0.152939
R14944 gnd.n5606 gnd.n5605 0.152939
R14945 gnd.n5606 gnd.n3371 0.152939
R14946 gnd.n5619 gnd.n3371 0.152939
R14947 gnd.n5620 gnd.n5619 0.152939
R14948 gnd.n5621 gnd.n5620 0.152939
R14949 gnd.n5621 gnd.n3366 0.152939
R14950 gnd.n5634 gnd.n3366 0.152939
R14951 gnd.n5635 gnd.n5634 0.152939
R14952 gnd.n5636 gnd.n5635 0.152939
R14953 gnd.n5636 gnd.n3362 0.152939
R14954 gnd.n5649 gnd.n3362 0.152939
R14955 gnd.n5650 gnd.n5649 0.152939
R14956 gnd.n5651 gnd.n5650 0.152939
R14957 gnd.n5651 gnd.n3357 0.152939
R14958 gnd.n5664 gnd.n3357 0.152939
R14959 gnd.n5665 gnd.n5664 0.152939
R14960 gnd.n5678 gnd.n5665 0.152939
R14961 gnd.n5678 gnd.n5677 0.152939
R14962 gnd.n5677 gnd.n5676 0.152939
R14963 gnd.n5676 gnd.n5666 0.152939
R14964 gnd.n5672 gnd.n5666 0.152939
R14965 gnd.n5672 gnd.n5671 0.152939
R14966 gnd.n5671 gnd.n95 0.152939
R14967 gnd.n7952 gnd.n7951 0.145814
R14968 gnd.n4284 gnd.n4283 0.145814
R14969 gnd.n4284 gnd.n3992 0.145814
R14970 gnd.n7952 gnd.n95 0.145814
R14971 gnd.n4657 gnd.n4656 0.128549
R14972 gnd.n6081 gnd.n6080 0.128549
R14973 gnd.n5716 gnd.n111 0.0797683
R14974 gnd.n4260 gnd.n2616 0.0797683
R14975 gnd.n1846 gnd.n1245 0.0767195
R14976 gnd.n1846 gnd.n1845 0.0767195
R14977 gnd.n4323 gnd.n2616 0.0736707
R14978 gnd.n5524 gnd.n111 0.0736707
R14979 gnd.n4754 gnd.n4657 0.063
R14980 gnd.n6080 gnd.n3010 0.063
R14981 gnd.n6684 gnd.n1009 0.0477147
R14982 gnd.n1636 gnd.n1524 0.0442063
R14983 gnd.n1637 gnd.n1636 0.0442063
R14984 gnd.n1638 gnd.n1637 0.0442063
R14985 gnd.n1638 gnd.n1513 0.0442063
R14986 gnd.n1652 gnd.n1513 0.0442063
R14987 gnd.n1653 gnd.n1652 0.0442063
R14988 gnd.n1654 gnd.n1653 0.0442063
R14989 gnd.n1654 gnd.n1500 0.0442063
R14990 gnd.n1698 gnd.n1500 0.0442063
R14991 gnd.n1699 gnd.n1698 0.0442063
R14992 gnd.n3178 gnd.n3010 0.0416005
R14993 gnd.n7733 gnd.n7732 0.0416005
R14994 gnd.n6506 gnd.n6505 0.0416005
R14995 gnd.n4755 gnd.n4754 0.0416005
R14996 gnd.n1701 gnd.n1434 0.0344674
R14997 gnd.n5902 gnd.n3178 0.0344674
R14998 gnd.n5902 gnd.n3180 0.0344674
R14999 gnd.n3204 gnd.n3180 0.0344674
R15000 gnd.n3205 gnd.n3204 0.0344674
R15001 gnd.n3206 gnd.n3205 0.0344674
R15002 gnd.n3207 gnd.n3206 0.0344674
R15003 gnd.n5598 gnd.n3207 0.0344674
R15004 gnd.n5598 gnd.n3226 0.0344674
R15005 gnd.n3227 gnd.n3226 0.0344674
R15006 gnd.n3228 gnd.n3227 0.0344674
R15007 gnd.n5613 gnd.n3228 0.0344674
R15008 gnd.n5613 gnd.n3246 0.0344674
R15009 gnd.n3247 gnd.n3246 0.0344674
R15010 gnd.n3248 gnd.n3247 0.0344674
R15011 gnd.n5628 gnd.n3248 0.0344674
R15012 gnd.n5628 gnd.n3267 0.0344674
R15013 gnd.n3268 gnd.n3267 0.0344674
R15014 gnd.n3269 gnd.n3268 0.0344674
R15015 gnd.n5643 gnd.n3269 0.0344674
R15016 gnd.n5643 gnd.n3287 0.0344674
R15017 gnd.n3288 gnd.n3287 0.0344674
R15018 gnd.n3289 gnd.n3288 0.0344674
R15019 gnd.n5658 gnd.n3289 0.0344674
R15020 gnd.n5658 gnd.n3309 0.0344674
R15021 gnd.n3310 gnd.n3309 0.0344674
R15022 gnd.n3311 gnd.n3310 0.0344674
R15023 gnd.n3353 gnd.n3311 0.0344674
R15024 gnd.n5689 gnd.n3353 0.0344674
R15025 gnd.n5694 gnd.n5689 0.0344674
R15026 gnd.n5695 gnd.n5694 0.0344674
R15027 gnd.n5695 gnd.n3344 0.0344674
R15028 gnd.n3345 gnd.n3344 0.0344674
R15029 gnd.n3346 gnd.n3345 0.0344674
R15030 gnd.n5699 gnd.n3346 0.0344674
R15031 gnd.n5700 gnd.n5699 0.0344674
R15032 gnd.n5701 gnd.n5700 0.0344674
R15033 gnd.n5701 gnd.n125 0.0344674
R15034 gnd.n126 gnd.n125 0.0344674
R15035 gnd.n127 gnd.n126 0.0344674
R15036 gnd.n5734 gnd.n127 0.0344674
R15037 gnd.n5734 gnd.n143 0.0344674
R15038 gnd.n144 gnd.n143 0.0344674
R15039 gnd.n145 gnd.n144 0.0344674
R15040 gnd.n5760 gnd.n145 0.0344674
R15041 gnd.n5760 gnd.n164 0.0344674
R15042 gnd.n165 gnd.n164 0.0344674
R15043 gnd.n166 gnd.n165 0.0344674
R15044 gnd.n356 gnd.n166 0.0344674
R15045 gnd.n356 gnd.n183 0.0344674
R15046 gnd.n184 gnd.n183 0.0344674
R15047 gnd.n185 gnd.n184 0.0344674
R15048 gnd.n7708 gnd.n185 0.0344674
R15049 gnd.n7708 gnd.n204 0.0344674
R15050 gnd.n205 gnd.n204 0.0344674
R15051 gnd.n206 gnd.n205 0.0344674
R15052 gnd.n7715 gnd.n206 0.0344674
R15053 gnd.n7715 gnd.n222 0.0344674
R15054 gnd.n223 gnd.n222 0.0344674
R15055 gnd.n224 gnd.n223 0.0344674
R15056 gnd.n7722 gnd.n224 0.0344674
R15057 gnd.n7722 gnd.n242 0.0344674
R15058 gnd.n243 gnd.n242 0.0344674
R15059 gnd.n244 gnd.n243 0.0344674
R15060 gnd.n7732 gnd.n244 0.0344674
R15061 gnd.n6505 gnd.n2464 0.0344674
R15062 gnd.n4045 gnd.n2464 0.0344674
R15063 gnd.n4045 gnd.n2486 0.0344674
R15064 gnd.n2487 gnd.n2486 0.0344674
R15065 gnd.n2488 gnd.n2487 0.0344674
R15066 gnd.n4051 gnd.n2488 0.0344674
R15067 gnd.n4051 gnd.n2505 0.0344674
R15068 gnd.n2506 gnd.n2505 0.0344674
R15069 gnd.n2507 gnd.n2506 0.0344674
R15070 gnd.n4058 gnd.n2507 0.0344674
R15071 gnd.n4058 gnd.n2524 0.0344674
R15072 gnd.n2525 gnd.n2524 0.0344674
R15073 gnd.n2526 gnd.n2525 0.0344674
R15074 gnd.n4065 gnd.n2526 0.0344674
R15075 gnd.n4065 gnd.n2544 0.0344674
R15076 gnd.n2545 gnd.n2544 0.0344674
R15077 gnd.n2546 gnd.n2545 0.0344674
R15078 gnd.n4175 gnd.n2546 0.0344674
R15079 gnd.n4175 gnd.n2564 0.0344674
R15080 gnd.n2565 gnd.n2564 0.0344674
R15081 gnd.n2566 gnd.n2565 0.0344674
R15082 gnd.n4178 gnd.n2566 0.0344674
R15083 gnd.n4178 gnd.n2584 0.0344674
R15084 gnd.n2585 gnd.n2584 0.0344674
R15085 gnd.n2586 gnd.n2585 0.0344674
R15086 gnd.n4233 gnd.n2586 0.0344674
R15087 gnd.n4233 gnd.n2603 0.0344674
R15088 gnd.n2604 gnd.n2603 0.0344674
R15089 gnd.n2605 gnd.n2604 0.0344674
R15090 gnd.n4242 gnd.n2605 0.0344674
R15091 gnd.n4242 gnd.n4241 0.0344674
R15092 gnd.n4241 gnd.n4010 0.0344674
R15093 gnd.n4010 gnd.n4006 0.0344674
R15094 gnd.n4007 gnd.n4006 0.0344674
R15095 gnd.n4297 gnd.n4007 0.0344674
R15096 gnd.n4297 gnd.n4008 0.0344674
R15097 gnd.n4008 gnd.n2631 0.0344674
R15098 gnd.n2632 gnd.n2631 0.0344674
R15099 gnd.n2633 gnd.n2632 0.0344674
R15100 gnd.n3978 gnd.n2633 0.0344674
R15101 gnd.n3978 gnd.n2649 0.0344674
R15102 gnd.n2650 gnd.n2649 0.0344674
R15103 gnd.n2651 gnd.n2650 0.0344674
R15104 gnd.n3972 gnd.n2651 0.0344674
R15105 gnd.n3972 gnd.n2670 0.0344674
R15106 gnd.n2671 gnd.n2670 0.0344674
R15107 gnd.n2672 gnd.n2671 0.0344674
R15108 gnd.n4376 gnd.n2672 0.0344674
R15109 gnd.n4376 gnd.n2689 0.0344674
R15110 gnd.n2690 gnd.n2689 0.0344674
R15111 gnd.n2691 gnd.n2690 0.0344674
R15112 gnd.n4386 gnd.n2691 0.0344674
R15113 gnd.n4386 gnd.n2710 0.0344674
R15114 gnd.n2711 gnd.n2710 0.0344674
R15115 gnd.n2712 gnd.n2711 0.0344674
R15116 gnd.n3947 gnd.n2712 0.0344674
R15117 gnd.n3947 gnd.n2729 0.0344674
R15118 gnd.n2730 gnd.n2729 0.0344674
R15119 gnd.n2731 gnd.n2730 0.0344674
R15120 gnd.n3941 gnd.n2731 0.0344674
R15121 gnd.n3941 gnd.n2750 0.0344674
R15122 gnd.n2751 gnd.n2750 0.0344674
R15123 gnd.n2752 gnd.n2751 0.0344674
R15124 gnd.n4755 gnd.n2752 0.0344674
R15125 gnd.n4652 gnd.n4477 0.0344674
R15126 gnd.n6079 gnd.n6078 0.0344674
R15127 gnd.n4601 gnd.n3909 0.029712
R15128 gnd.n5581 gnd.n5580 0.029712
R15129 gnd.n1721 gnd.n1720 0.0269946
R15130 gnd.n1723 gnd.n1722 0.0269946
R15131 gnd.n1429 gnd.n1427 0.0269946
R15132 gnd.n1733 gnd.n1731 0.0269946
R15133 gnd.n1732 gnd.n1408 0.0269946
R15134 gnd.n1752 gnd.n1751 0.0269946
R15135 gnd.n1754 gnd.n1753 0.0269946
R15136 gnd.n1403 gnd.n1402 0.0269946
R15137 gnd.n1764 gnd.n1398 0.0269946
R15138 gnd.n1763 gnd.n1400 0.0269946
R15139 gnd.n1399 gnd.n1379 0.0269946
R15140 gnd.n1790 gnd.n1380 0.0269946
R15141 gnd.n1789 gnd.n1381 0.0269946
R15142 gnd.n1809 gnd.n1365 0.0269946
R15143 gnd.n1811 gnd.n1810 0.0269946
R15144 gnd.n1812 gnd.n1345 0.0269946
R15145 gnd.n1813 gnd.n1346 0.0269946
R15146 gnd.n1814 gnd.n1347 0.0269946
R15147 gnd.n1349 gnd.n1348 0.0269946
R15148 gnd.n1238 gnd.n1237 0.0269946
R15149 gnd.n1858 gnd.n1234 0.0269946
R15150 gnd.n1857 gnd.n1235 0.0269946
R15151 gnd.n1877 gnd.n1217 0.0269946
R15152 gnd.n1879 gnd.n1878 0.0269946
R15153 gnd.n1880 gnd.n1215 0.0269946
R15154 gnd.n1887 gnd.n1883 0.0269946
R15155 gnd.n1886 gnd.n1885 0.0269946
R15156 gnd.n1884 gnd.n1194 0.0269946
R15157 gnd.n1910 gnd.n1195 0.0269946
R15158 gnd.n1909 gnd.n1196 0.0269946
R15159 gnd.n1955 gnd.n1172 0.0269946
R15160 gnd.n1957 gnd.n1956 0.0269946
R15161 gnd.n1966 gnd.n1165 0.0269946
R15162 gnd.n1968 gnd.n1967 0.0269946
R15163 gnd.n1969 gnd.n1163 0.0269946
R15164 gnd.n1976 gnd.n1972 0.0269946
R15165 gnd.n1975 gnd.n1974 0.0269946
R15166 gnd.n1973 gnd.n1143 0.0269946
R15167 gnd.n2000 gnd.n1144 0.0269946
R15168 gnd.n1999 gnd.n1145 0.0269946
R15169 gnd.n2060 gnd.n1120 0.0269946
R15170 gnd.n2062 gnd.n2061 0.0269946
R15171 gnd.n2063 gnd.n959 0.0269946
R15172 gnd.n1115 gnd.n960 0.0269946
R15173 gnd.n1117 gnd.n961 0.0269946
R15174 gnd.n2071 gnd.n2070 0.0269946
R15175 gnd.n2073 gnd.n2072 0.0269946
R15176 gnd.n2074 gnd.n983 0.0269946
R15177 gnd.n2334 gnd.n985 0.0269946
R15178 gnd.n2340 gnd.n2339 0.0269946
R15179 gnd.n2342 gnd.n2341 0.0269946
R15180 gnd.n6685 gnd.n1008 0.0269946
R15181 gnd.n4651 gnd.n4538 0.0225788
R15182 gnd.n4648 gnd.n4647 0.0225788
R15183 gnd.n4644 gnd.n4541 0.0225788
R15184 gnd.n4643 gnd.n4547 0.0225788
R15185 gnd.n4640 gnd.n4639 0.0225788
R15186 gnd.n4636 gnd.n4553 0.0225788
R15187 gnd.n4635 gnd.n4557 0.0225788
R15188 gnd.n4632 gnd.n4631 0.0225788
R15189 gnd.n4628 gnd.n4561 0.0225788
R15190 gnd.n4627 gnd.n4567 0.0225788
R15191 gnd.n4624 gnd.n4623 0.0225788
R15192 gnd.n4620 gnd.n4573 0.0225788
R15193 gnd.n4619 gnd.n4577 0.0225788
R15194 gnd.n4616 gnd.n4615 0.0225788
R15195 gnd.n4612 gnd.n4581 0.0225788
R15196 gnd.n4611 gnd.n4587 0.0225788
R15197 gnd.n4608 gnd.n4607 0.0225788
R15198 gnd.n4604 gnd.n4595 0.0225788
R15199 gnd.n4603 gnd.n4601 0.0225788
R15200 gnd.n6075 gnd.n3011 0.0225788
R15201 gnd.n6074 gnd.n3015 0.0225788
R15202 gnd.n6071 gnd.n6070 0.0225788
R15203 gnd.n6067 gnd.n3020 0.0225788
R15204 gnd.n6066 gnd.n3024 0.0225788
R15205 gnd.n6063 gnd.n6062 0.0225788
R15206 gnd.n6059 gnd.n3028 0.0225788
R15207 gnd.n6058 gnd.n3032 0.0225788
R15208 gnd.n6055 gnd.n6054 0.0225788
R15209 gnd.n6051 gnd.n3036 0.0225788
R15210 gnd.n6050 gnd.n3040 0.0225788
R15211 gnd.n6047 gnd.n6046 0.0225788
R15212 gnd.n6043 gnd.n3044 0.0225788
R15213 gnd.n6042 gnd.n3048 0.0225788
R15214 gnd.n6039 gnd.n6038 0.0225788
R15215 gnd.n6035 gnd.n3052 0.0225788
R15216 gnd.n6034 gnd.n3058 0.0225788
R15217 gnd.n3383 gnd.n3061 0.0225788
R15218 gnd.n5580 gnd.n3382 0.0225788
R15219 gnd.n5581 gnd.n2991 0.0218415
R15220 gnd.n4784 gnd.n3909 0.0218415
R15221 gnd.n1701 gnd.n1700 0.0202011
R15222 gnd.n1700 gnd.n1699 0.0148637
R15223 gnd.n2332 gnd.n2331 0.0144266
R15224 gnd.n2331 gnd.n984 0.0130679
R15225 gnd.n4652 gnd.n4651 0.0123886
R15226 gnd.n4648 gnd.n4538 0.0123886
R15227 gnd.n4647 gnd.n4541 0.0123886
R15228 gnd.n4644 gnd.n4643 0.0123886
R15229 gnd.n4640 gnd.n4547 0.0123886
R15230 gnd.n4639 gnd.n4553 0.0123886
R15231 gnd.n4636 gnd.n4635 0.0123886
R15232 gnd.n4632 gnd.n4557 0.0123886
R15233 gnd.n4631 gnd.n4561 0.0123886
R15234 gnd.n4628 gnd.n4627 0.0123886
R15235 gnd.n4624 gnd.n4567 0.0123886
R15236 gnd.n4623 gnd.n4573 0.0123886
R15237 gnd.n4620 gnd.n4619 0.0123886
R15238 gnd.n4616 gnd.n4577 0.0123886
R15239 gnd.n4615 gnd.n4581 0.0123886
R15240 gnd.n4612 gnd.n4611 0.0123886
R15241 gnd.n4608 gnd.n4587 0.0123886
R15242 gnd.n4607 gnd.n4595 0.0123886
R15243 gnd.n4604 gnd.n4603 0.0123886
R15244 gnd.n6078 gnd.n3011 0.0123886
R15245 gnd.n6075 gnd.n6074 0.0123886
R15246 gnd.n6071 gnd.n3015 0.0123886
R15247 gnd.n6070 gnd.n3020 0.0123886
R15248 gnd.n6067 gnd.n6066 0.0123886
R15249 gnd.n6063 gnd.n3024 0.0123886
R15250 gnd.n6062 gnd.n3028 0.0123886
R15251 gnd.n6059 gnd.n6058 0.0123886
R15252 gnd.n6055 gnd.n3032 0.0123886
R15253 gnd.n6054 gnd.n3036 0.0123886
R15254 gnd.n6051 gnd.n6050 0.0123886
R15255 gnd.n6047 gnd.n3040 0.0123886
R15256 gnd.n6046 gnd.n3044 0.0123886
R15257 gnd.n6043 gnd.n6042 0.0123886
R15258 gnd.n6039 gnd.n3048 0.0123886
R15259 gnd.n6038 gnd.n3052 0.0123886
R15260 gnd.n6035 gnd.n6034 0.0123886
R15261 gnd.n3061 gnd.n3058 0.0123886
R15262 gnd.n3383 gnd.n3382 0.0123886
R15263 gnd.n1720 gnd.n1434 0.00797283
R15264 gnd.n1722 gnd.n1721 0.00797283
R15265 gnd.n1723 gnd.n1429 0.00797283
R15266 gnd.n1731 gnd.n1427 0.00797283
R15267 gnd.n1733 gnd.n1732 0.00797283
R15268 gnd.n1751 gnd.n1408 0.00797283
R15269 gnd.n1753 gnd.n1752 0.00797283
R15270 gnd.n1754 gnd.n1403 0.00797283
R15271 gnd.n1402 gnd.n1398 0.00797283
R15272 gnd.n1764 gnd.n1763 0.00797283
R15273 gnd.n1400 gnd.n1399 0.00797283
R15274 gnd.n1380 gnd.n1379 0.00797283
R15275 gnd.n1790 gnd.n1789 0.00797283
R15276 gnd.n1381 gnd.n1365 0.00797283
R15277 gnd.n1810 gnd.n1809 0.00797283
R15278 gnd.n1812 gnd.n1811 0.00797283
R15279 gnd.n1813 gnd.n1345 0.00797283
R15280 gnd.n1814 gnd.n1346 0.00797283
R15281 gnd.n1348 gnd.n1347 0.00797283
R15282 gnd.n1349 gnd.n1238 0.00797283
R15283 gnd.n1237 gnd.n1234 0.00797283
R15284 gnd.n1858 gnd.n1857 0.00797283
R15285 gnd.n1235 gnd.n1217 0.00797283
R15286 gnd.n1878 gnd.n1877 0.00797283
R15287 gnd.n1880 gnd.n1879 0.00797283
R15288 gnd.n1883 gnd.n1215 0.00797283
R15289 gnd.n1887 gnd.n1886 0.00797283
R15290 gnd.n1885 gnd.n1884 0.00797283
R15291 gnd.n1195 gnd.n1194 0.00797283
R15292 gnd.n1910 gnd.n1909 0.00797283
R15293 gnd.n1196 gnd.n1172 0.00797283
R15294 gnd.n1957 gnd.n1955 0.00797283
R15295 gnd.n1956 gnd.n1165 0.00797283
R15296 gnd.n1967 gnd.n1966 0.00797283
R15297 gnd.n1969 gnd.n1968 0.00797283
R15298 gnd.n1972 gnd.n1163 0.00797283
R15299 gnd.n1976 gnd.n1975 0.00797283
R15300 gnd.n1974 gnd.n1973 0.00797283
R15301 gnd.n1144 gnd.n1143 0.00797283
R15302 gnd.n2000 gnd.n1999 0.00797283
R15303 gnd.n1145 gnd.n1120 0.00797283
R15304 gnd.n2061 gnd.n2060 0.00797283
R15305 gnd.n2063 gnd.n2062 0.00797283
R15306 gnd.n1115 gnd.n959 0.00797283
R15307 gnd.n1117 gnd.n960 0.00797283
R15308 gnd.n2070 gnd.n961 0.00797283
R15309 gnd.n2072 gnd.n2071 0.00797283
R15310 gnd.n2074 gnd.n2073 0.00797283
R15311 gnd.n2332 gnd.n983 0.00797283
R15312 gnd.n2334 gnd.n984 0.00797283
R15313 gnd.n2339 gnd.n985 0.00797283
R15314 gnd.n2342 gnd.n2340 0.00797283
R15315 gnd.n2341 gnd.n1008 0.00797283
R15316 gnd.n6685 gnd.n6684 0.00797283
R15317 gnd.n4657 gnd.n4477 0.00593478
R15318 gnd.n6080 gnd.n6079 0.00593478
R15319 a_n2982_13878.n74 a_n2982_13878.t12 532.5
R15320 a_n2982_13878.n149 a_n2982_13878.t10 512.366
R15321 a_n2982_13878.n148 a_n2982_13878.t30 512.366
R15322 a_n2982_13878.n83 a_n2982_13878.t26 512.366
R15323 a_n2982_13878.n147 a_n2982_13878.t48 512.366
R15324 a_n2982_13878.n146 a_n2982_13878.t6 512.366
R15325 a_n2982_13878.n84 a_n2982_13878.t50 512.366
R15326 a_n2982_13878.n145 a_n2982_13878.t34 512.366
R15327 a_n2982_13878.n144 a_n2982_13878.t22 512.366
R15328 a_n2982_13878.n85 a_n2982_13878.t38 512.366
R15329 a_n2982_13878.n143 a_n2982_13878.t42 512.366
R15330 a_n2982_13878.n12 a_n2982_13878.t102 538.698
R15331 a_n2982_13878.n134 a_n2982_13878.t79 512.366
R15332 a_n2982_13878.n133 a_n2982_13878.t84 512.366
R15333 a_n2982_13878.n86 a_n2982_13878.t72 512.366
R15334 a_n2982_13878.n132 a_n2982_13878.t89 512.366
R15335 a_n2982_13878.n131 a_n2982_13878.t98 512.366
R15336 a_n2982_13878.n87 a_n2982_13878.t99 512.366
R15337 a_n2982_13878.n130 a_n2982_13878.t66 512.366
R15338 a_n2982_13878.n129 a_n2982_13878.t81 512.366
R15339 a_n2982_13878.n88 a_n2982_13878.t69 512.366
R15340 a_n2982_13878.n128 a_n2982_13878.t76 512.366
R15341 a_n2982_13878.n27 a_n2982_13878.t8 538.698
R15342 a_n2982_13878.n108 a_n2982_13878.t44 512.366
R15343 a_n2982_13878.n97 a_n2982_13878.t52 512.366
R15344 a_n2982_13878.n109 a_n2982_13878.t46 512.366
R15345 a_n2982_13878.n96 a_n2982_13878.t20 512.366
R15346 a_n2982_13878.n110 a_n2982_13878.t32 512.366
R15347 a_n2982_13878.n111 a_n2982_13878.t14 512.366
R15348 a_n2982_13878.n95 a_n2982_13878.t36 512.366
R15349 a_n2982_13878.n112 a_n2982_13878.t16 512.366
R15350 a_n2982_13878.n94 a_n2982_13878.t24 512.366
R15351 a_n2982_13878.n113 a_n2982_13878.t28 512.366
R15352 a_n2982_13878.n33 a_n2982_13878.t101 538.698
R15353 a_n2982_13878.n102 a_n2982_13878.t70 512.366
R15354 a_n2982_13878.n101 a_n2982_13878.t71 512.366
R15355 a_n2982_13878.n103 a_n2982_13878.t96 512.366
R15356 a_n2982_13878.n100 a_n2982_13878.t97 512.366
R15357 a_n2982_13878.n104 a_n2982_13878.t68 512.366
R15358 a_n2982_13878.n105 a_n2982_13878.t92 512.366
R15359 a_n2982_13878.n99 a_n2982_13878.t93 512.366
R15360 a_n2982_13878.n106 a_n2982_13878.t65 512.366
R15361 a_n2982_13878.n98 a_n2982_13878.t78 512.366
R15362 a_n2982_13878.n107 a_n2982_13878.t87 512.366
R15363 a_n2982_13878.n125 a_n2982_13878.t86 512.366
R15364 a_n2982_13878.n115 a_n2982_13878.t75 512.366
R15365 a_n2982_13878.n126 a_n2982_13878.t64 512.366
R15366 a_n2982_13878.n123 a_n2982_13878.t94 512.366
R15367 a_n2982_13878.n116 a_n2982_13878.t83 512.366
R15368 a_n2982_13878.n124 a_n2982_13878.t82 512.366
R15369 a_n2982_13878.n121 a_n2982_13878.t90 512.366
R15370 a_n2982_13878.n117 a_n2982_13878.t73 512.366
R15371 a_n2982_13878.n122 a_n2982_13878.t74 512.366
R15372 a_n2982_13878.n119 a_n2982_13878.t77 512.366
R15373 a_n2982_13878.n118 a_n2982_13878.t88 512.366
R15374 a_n2982_13878.n120 a_n2982_13878.t103 512.366
R15375 a_n2982_13878.n35 a_n2982_13878.n34 44.7878
R15376 a_n2982_13878.n73 a_n2982_13878.n7 70.5844
R15377 a_n2982_13878.n23 a_n2982_13878.n57 70.5844
R15378 a_n2982_13878.n29 a_n2982_13878.n49 70.5844
R15379 a_n2982_13878.n48 a_n2982_13878.n29 70.1674
R15380 a_n2982_13878.n48 a_n2982_13878.n98 20.9683
R15381 a_n2982_13878.n28 a_n2982_13878.n47 74.73
R15382 a_n2982_13878.n106 a_n2982_13878.n47 11.843
R15383 a_n2982_13878.n46 a_n2982_13878.n28 80.4688
R15384 a_n2982_13878.n46 a_n2982_13878.n99 0.365327
R15385 a_n2982_13878.n30 a_n2982_13878.n45 75.0448
R15386 a_n2982_13878.n44 a_n2982_13878.n30 70.1674
R15387 a_n2982_13878.n44 a_n2982_13878.n100 20.9683
R15388 a_n2982_13878.n31 a_n2982_13878.n43 70.3058
R15389 a_n2982_13878.n103 a_n2982_13878.n43 20.6913
R15390 a_n2982_13878.n42 a_n2982_13878.n31 75.3623
R15391 a_n2982_13878.n42 a_n2982_13878.n101 10.5784
R15392 a_n2982_13878.n33 a_n2982_13878.n32 44.7878
R15393 a_n2982_13878.n56 a_n2982_13878.n23 70.1674
R15394 a_n2982_13878.n56 a_n2982_13878.n94 20.9683
R15395 a_n2982_13878.n22 a_n2982_13878.n55 74.73
R15396 a_n2982_13878.n112 a_n2982_13878.n55 11.843
R15397 a_n2982_13878.n54 a_n2982_13878.n22 80.4688
R15398 a_n2982_13878.n54 a_n2982_13878.n95 0.365327
R15399 a_n2982_13878.n24 a_n2982_13878.n53 75.0448
R15400 a_n2982_13878.n52 a_n2982_13878.n24 70.1674
R15401 a_n2982_13878.n52 a_n2982_13878.n96 20.9683
R15402 a_n2982_13878.n25 a_n2982_13878.n51 70.3058
R15403 a_n2982_13878.n109 a_n2982_13878.n51 20.6913
R15404 a_n2982_13878.n50 a_n2982_13878.n25 75.3623
R15405 a_n2982_13878.n50 a_n2982_13878.n97 10.5784
R15406 a_n2982_13878.n27 a_n2982_13878.n26 44.7878
R15407 a_n2982_13878.n13 a_n2982_13878.n65 70.1674
R15408 a_n2982_13878.n15 a_n2982_13878.n63 70.1674
R15409 a_n2982_13878.n17 a_n2982_13878.n61 70.1674
R15410 a_n2982_13878.n20 a_n2982_13878.n59 70.1674
R15411 a_n2982_13878.n120 a_n2982_13878.n59 20.9683
R15412 a_n2982_13878.n58 a_n2982_13878.n21 75.0448
R15413 a_n2982_13878.n58 a_n2982_13878.n118 11.2134
R15414 a_n2982_13878.n21 a_n2982_13878.n119 161.3
R15415 a_n2982_13878.n122 a_n2982_13878.n61 20.9683
R15416 a_n2982_13878.n60 a_n2982_13878.n18 75.0448
R15417 a_n2982_13878.n60 a_n2982_13878.n117 11.2134
R15418 a_n2982_13878.n18 a_n2982_13878.n121 161.3
R15419 a_n2982_13878.n124 a_n2982_13878.n63 20.9683
R15420 a_n2982_13878.n62 a_n2982_13878.n16 75.0448
R15421 a_n2982_13878.n62 a_n2982_13878.n116 11.2134
R15422 a_n2982_13878.n16 a_n2982_13878.n123 161.3
R15423 a_n2982_13878.n126 a_n2982_13878.n65 20.9683
R15424 a_n2982_13878.n64 a_n2982_13878.n14 75.0448
R15425 a_n2982_13878.n64 a_n2982_13878.n115 11.2134
R15426 a_n2982_13878.n14 a_n2982_13878.n125 161.3
R15427 a_n2982_13878.n7 a_n2982_13878.n72 70.1674
R15428 a_n2982_13878.n72 a_n2982_13878.n88 20.9683
R15429 a_n2982_13878.n71 a_n2982_13878.n8 74.73
R15430 a_n2982_13878.n129 a_n2982_13878.n71 11.843
R15431 a_n2982_13878.n70 a_n2982_13878.n8 80.4688
R15432 a_n2982_13878.n70 a_n2982_13878.n130 0.365327
R15433 a_n2982_13878.n9 a_n2982_13878.n69 75.0448
R15434 a_n2982_13878.n68 a_n2982_13878.n9 70.1674
R15435 a_n2982_13878.n132 a_n2982_13878.n68 20.9683
R15436 a_n2982_13878.n11 a_n2982_13878.n67 70.3058
R15437 a_n2982_13878.n67 a_n2982_13878.n86 20.6913
R15438 a_n2982_13878.n66 a_n2982_13878.n11 75.3623
R15439 a_n2982_13878.n133 a_n2982_13878.n66 10.5784
R15440 a_n2982_13878.n10 a_n2982_13878.n12 44.7878
R15441 a_n2982_13878.n35 a_n2982_13878.n143 14.1668
R15442 a_n2982_13878.n82 a_n2982_13878.n81 75.3623
R15443 a_n2982_13878.n80 a_n2982_13878.n3 70.3058
R15444 a_n2982_13878.n3 a_n2982_13878.n79 70.1674
R15445 a_n2982_13878.n79 a_n2982_13878.n84 20.9683
R15446 a_n2982_13878.n78 a_n2982_13878.n4 75.0448
R15447 a_n2982_13878.n146 a_n2982_13878.n78 11.2134
R15448 a_n2982_13878.n77 a_n2982_13878.n4 80.4688
R15449 a_n2982_13878.n6 a_n2982_13878.n76 74.73
R15450 a_n2982_13878.n75 a_n2982_13878.n6 70.1674
R15451 a_n2982_13878.n149 a_n2982_13878.n75 20.9683
R15452 a_n2982_13878.n5 a_n2982_13878.n74 70.5844
R15453 a_n2982_13878.n1 a_n2982_13878.n141 81.3764
R15454 a_n2982_13878.n2 a_n2982_13878.n137 81.3764
R15455 a_n2982_13878.n2 a_n2982_13878.n135 81.3764
R15456 a_n2982_13878.n1 a_n2982_13878.n142 80.9324
R15457 a_n2982_13878.n1 a_n2982_13878.n140 80.9324
R15458 a_n2982_13878.n0 a_n2982_13878.n139 80.9324
R15459 a_n2982_13878.n2 a_n2982_13878.n138 80.9324
R15460 a_n2982_13878.n2 a_n2982_13878.n136 80.9324
R15461 a_n2982_13878.n40 a_n2982_13878.t41 74.6477
R15462 a_n2982_13878.n36 a_n2982_13878.t9 74.6477
R15463 a_n2982_13878.n39 a_n2982_13878.t13 74.2899
R15464 a_n2982_13878.n38 a_n2982_13878.t19 74.2897
R15465 a_n2982_13878.n40 a_n2982_13878.n153 70.6783
R15466 a_n2982_13878.n40 a_n2982_13878.n154 70.6783
R15467 a_n2982_13878.n41 a_n2982_13878.n152 70.6783
R15468 a_n2982_13878.n39 a_n2982_13878.n151 70.6783
R15469 a_n2982_13878.n38 a_n2982_13878.n93 70.6783
R15470 a_n2982_13878.n37 a_n2982_13878.n92 70.6783
R15471 a_n2982_13878.n37 a_n2982_13878.n91 70.6783
R15472 a_n2982_13878.n36 a_n2982_13878.n90 70.6783
R15473 a_n2982_13878.n36 a_n2982_13878.n89 70.6783
R15474 a_n2982_13878.n155 a_n2982_13878.n41 70.6782
R15475 a_n2982_13878.n75 a_n2982_13878.n148 20.9683
R15476 a_n2982_13878.n147 a_n2982_13878.n146 48.2005
R15477 a_n2982_13878.n145 a_n2982_13878.n79 20.9683
R15478 a_n2982_13878.n143 a_n2982_13878.n85 48.2005
R15479 a_n2982_13878.n134 a_n2982_13878.n133 48.2005
R15480 a_n2982_13878.n68 a_n2982_13878.n131 20.9683
R15481 a_n2982_13878.n130 a_n2982_13878.n87 48.2005
R15482 a_n2982_13878.n128 a_n2982_13878.n72 20.9683
R15483 a_n2982_13878.n108 a_n2982_13878.n97 48.2005
R15484 a_n2982_13878.n110 a_n2982_13878.n52 20.9683
R15485 a_n2982_13878.n111 a_n2982_13878.n95 48.2005
R15486 a_n2982_13878.n113 a_n2982_13878.n56 20.9683
R15487 a_n2982_13878.n102 a_n2982_13878.n101 48.2005
R15488 a_n2982_13878.n104 a_n2982_13878.n44 20.9683
R15489 a_n2982_13878.n105 a_n2982_13878.n99 48.2005
R15490 a_n2982_13878.n107 a_n2982_13878.n48 20.9683
R15491 a_n2982_13878.n125 a_n2982_13878.n115 48.2005
R15492 a_n2982_13878.t91 a_n2982_13878.n65 533.335
R15493 a_n2982_13878.n123 a_n2982_13878.n116 48.2005
R15494 a_n2982_13878.t100 a_n2982_13878.n63 533.335
R15495 a_n2982_13878.n121 a_n2982_13878.n117 48.2005
R15496 a_n2982_13878.t85 a_n2982_13878.n61 533.335
R15497 a_n2982_13878.n119 a_n2982_13878.n118 48.2005
R15498 a_n2982_13878.t80 a_n2982_13878.n59 533.335
R15499 a_n2982_13878.n77 a_n2982_13878.n83 47.835
R15500 a_n2982_13878.n80 a_n2982_13878.n144 20.6913
R15501 a_n2982_13878.n132 a_n2982_13878.n67 21.4216
R15502 a_n2982_13878.n96 a_n2982_13878.n51 21.4216
R15503 a_n2982_13878.n100 a_n2982_13878.n43 21.4216
R15504 a_n2982_13878.n73 a_n2982_13878.t95 532.5
R15505 a_n2982_13878.t18 a_n2982_13878.n57 532.5
R15506 a_n2982_13878.t67 a_n2982_13878.n49 532.5
R15507 a_n2982_13878.n76 a_n2982_13878.n83 11.843
R15508 a_n2982_13878.n144 a_n2982_13878.n81 36.139
R15509 a_n2982_13878.n71 a_n2982_13878.n88 34.4824
R15510 a_n2982_13878.n94 a_n2982_13878.n55 34.4824
R15511 a_n2982_13878.n98 a_n2982_13878.n47 34.4824
R15512 a_n2982_13878.n78 a_n2982_13878.n84 35.3134
R15513 a_n2982_13878.n131 a_n2982_13878.n69 35.3134
R15514 a_n2982_13878.n69 a_n2982_13878.n87 11.2134
R15515 a_n2982_13878.n53 a_n2982_13878.n110 35.3134
R15516 a_n2982_13878.n111 a_n2982_13878.n53 11.2134
R15517 a_n2982_13878.n45 a_n2982_13878.n104 35.3134
R15518 a_n2982_13878.n105 a_n2982_13878.n45 11.2134
R15519 a_n2982_13878.n126 a_n2982_13878.n64 35.3134
R15520 a_n2982_13878.n124 a_n2982_13878.n62 35.3134
R15521 a_n2982_13878.n122 a_n2982_13878.n60 35.3134
R15522 a_n2982_13878.n120 a_n2982_13878.n58 35.3134
R15523 a_n2982_13878.n34 a_n2982_13878.n1 23.891
R15524 a_n2982_13878.n148 a_n2982_13878.n76 34.4824
R15525 a_n2982_13878.n81 a_n2982_13878.n85 10.5784
R15526 a_n2982_13878.n66 a_n2982_13878.n86 36.139
R15527 a_n2982_13878.n109 a_n2982_13878.n50 36.139
R15528 a_n2982_13878.n103 a_n2982_13878.n42 36.139
R15529 a_n2982_13878.n32 a_n2982_13878.n19 13.9285
R15530 a_n2982_13878.n7 a_n2982_13878.n127 13.724
R15531 a_n2982_13878.n150 a_n2982_13878.n5 12.4191
R15532 a_n2982_13878.n21 a_n2982_13878.n19 11.2486
R15533 a_n2982_13878.n127 a_n2982_13878.n13 11.2486
R15534 a_n2982_13878.n114 a_n2982_13878.n38 10.5745
R15535 a_n2982_13878.n114 a_n2982_13878.n23 8.58383
R15536 a_n2982_13878.n39 a_n2982_13878.n150 6.7311
R15537 a_n2982_13878.n127 a_n2982_13878.n114 5.3452
R15538 a_n2982_13878.n26 a_n2982_13878.n29 3.94368
R15539 a_n2982_13878.n34 a_n2982_13878.n10 3.7202
R15540 a_n2982_13878.n153 a_n2982_13878.t39 3.61217
R15541 a_n2982_13878.n153 a_n2982_13878.t43 3.61217
R15542 a_n2982_13878.n154 a_n2982_13878.t35 3.61217
R15543 a_n2982_13878.n154 a_n2982_13878.t23 3.61217
R15544 a_n2982_13878.n152 a_n2982_13878.t27 3.61217
R15545 a_n2982_13878.n152 a_n2982_13878.t49 3.61217
R15546 a_n2982_13878.n151 a_n2982_13878.t11 3.61217
R15547 a_n2982_13878.n151 a_n2982_13878.t31 3.61217
R15548 a_n2982_13878.n93 a_n2982_13878.t25 3.61217
R15549 a_n2982_13878.n93 a_n2982_13878.t29 3.61217
R15550 a_n2982_13878.n92 a_n2982_13878.t37 3.61217
R15551 a_n2982_13878.n92 a_n2982_13878.t17 3.61217
R15552 a_n2982_13878.n91 a_n2982_13878.t33 3.61217
R15553 a_n2982_13878.n91 a_n2982_13878.t15 3.61217
R15554 a_n2982_13878.n90 a_n2982_13878.t47 3.61217
R15555 a_n2982_13878.n90 a_n2982_13878.t21 3.61217
R15556 a_n2982_13878.n89 a_n2982_13878.t45 3.61217
R15557 a_n2982_13878.n89 a_n2982_13878.t53 3.61217
R15558 a_n2982_13878.t7 a_n2982_13878.n155 3.61217
R15559 a_n2982_13878.n155 a_n2982_13878.t51 3.61217
R15560 a_n2982_13878.n141 a_n2982_13878.t1 2.82907
R15561 a_n2982_13878.n141 a_n2982_13878.t2 2.82907
R15562 a_n2982_13878.n142 a_n2982_13878.t3 2.82907
R15563 a_n2982_13878.n142 a_n2982_13878.t0 2.82907
R15564 a_n2982_13878.n140 a_n2982_13878.t62 2.82907
R15565 a_n2982_13878.n140 a_n2982_13878.t57 2.82907
R15566 a_n2982_13878.n139 a_n2982_13878.t59 2.82907
R15567 a_n2982_13878.n139 a_n2982_13878.t55 2.82907
R15568 a_n2982_13878.n137 a_n2982_13878.t54 2.82907
R15569 a_n2982_13878.n137 a_n2982_13878.t56 2.82907
R15570 a_n2982_13878.n138 a_n2982_13878.t61 2.82907
R15571 a_n2982_13878.n138 a_n2982_13878.t60 2.82907
R15572 a_n2982_13878.n136 a_n2982_13878.t4 2.82907
R15573 a_n2982_13878.n136 a_n2982_13878.t58 2.82907
R15574 a_n2982_13878.n135 a_n2982_13878.t5 2.82907
R15575 a_n2982_13878.n135 a_n2982_13878.t63 2.82907
R15576 a_n2982_13878.n74 a_n2982_13878.n149 22.3251
R15577 a_n2982_13878.n35 a_n2982_13878.t40 538.698
R15578 a_n2982_13878.n12 a_n2982_13878.n134 14.1668
R15579 a_n2982_13878.n128 a_n2982_13878.n73 22.3251
R15580 a_n2982_13878.n108 a_n2982_13878.n27 14.1668
R15581 a_n2982_13878.n57 a_n2982_13878.n113 22.3251
R15582 a_n2982_13878.n102 a_n2982_13878.n33 14.1668
R15583 a_n2982_13878.n49 a_n2982_13878.n107 22.3251
R15584 a_n2982_13878.n150 a_n2982_13878.n19 1.30542
R15585 a_n2982_13878.n16 a_n2982_13878.n17 1.04595
R15586 a_n2982_13878.n77 a_n2982_13878.n147 0.365327
R15587 a_n2982_13878.n145 a_n2982_13878.n80 21.4216
R15588 a_n2982_13878.n70 a_n2982_13878.n129 47.835
R15589 a_n2982_13878.n112 a_n2982_13878.n54 47.835
R15590 a_n2982_13878.n106 a_n2982_13878.n46 47.835
R15591 a_n2982_13878.n0 a_n2982_13878.n2 31.7919
R15592 a_n2982_13878.n29 a_n2982_13878.n28 1.13686
R15593 a_n2982_13878.n23 a_n2982_13878.n22 1.13686
R15594 a_n2982_13878.n8 a_n2982_13878.n7 1.13686
R15595 a_n2982_13878.n41 a_n2982_13878.n39 1.07378
R15596 a_n2982_13878.n37 a_n2982_13878.n36 1.07378
R15597 a_n2982_13878.n1 a_n2982_13878.n0 0.888431
R15598 a_n2982_13878.n31 a_n2982_13878.n32 0.758076
R15599 a_n2982_13878.n30 a_n2982_13878.n31 0.758076
R15600 a_n2982_13878.n28 a_n2982_13878.n30 0.758076
R15601 a_n2982_13878.n25 a_n2982_13878.n26 0.758076
R15602 a_n2982_13878.n24 a_n2982_13878.n25 0.758076
R15603 a_n2982_13878.n22 a_n2982_13878.n24 0.758076
R15604 a_n2982_13878.n21 a_n2982_13878.n20 0.758076
R15605 a_n2982_13878.n18 a_n2982_13878.n17 0.758076
R15606 a_n2982_13878.n16 a_n2982_13878.n15 0.758076
R15607 a_n2982_13878.n14 a_n2982_13878.n13 0.758076
R15608 a_n2982_13878.n11 a_n2982_13878.n10 0.758076
R15609 a_n2982_13878.n11 a_n2982_13878.n9 0.758076
R15610 a_n2982_13878.n9 a_n2982_13878.n8 0.758076
R15611 a_n2982_13878.n6 a_n2982_13878.n4 0.758076
R15612 a_n2982_13878.n4 a_n2982_13878.n3 0.758076
R15613 a_n2982_13878.n82 a_n2982_13878.n3 0.758076
R15614 a_n2982_13878.n82 a_n2982_13878.n34 0.754288
R15615 a_n2982_13878.n41 a_n2982_13878.n40 0.716017
R15616 a_n2982_13878.n38 a_n2982_13878.n37 0.716017
R15617 a_n2982_13878.n18 a_n2982_13878.n20 0.67853
R15618 a_n2982_13878.n14 a_n2982_13878.n15 0.67853
R15619 a_n2982_13878.n6 a_n2982_13878.n5 0.568682
R15620 a_n2804_13878.n29 a_n2804_13878.n28 98.9632
R15621 a_n2804_13878.n2 a_n2804_13878.n0 98.7517
R15622 a_n2804_13878.n22 a_n2804_13878.n21 98.6055
R15623 a_n2804_13878.n24 a_n2804_13878.n23 98.6055
R15624 a_n2804_13878.n26 a_n2804_13878.n25 98.6055
R15625 a_n2804_13878.n28 a_n2804_13878.n27 98.6055
R15626 a_n2804_13878.n10 a_n2804_13878.n9 98.6055
R15627 a_n2804_13878.n8 a_n2804_13878.n7 98.6055
R15628 a_n2804_13878.n6 a_n2804_13878.n5 98.6055
R15629 a_n2804_13878.n4 a_n2804_13878.n3 98.6055
R15630 a_n2804_13878.n2 a_n2804_13878.n1 98.6055
R15631 a_n2804_13878.n20 a_n2804_13878.n19 98.6054
R15632 a_n2804_13878.n12 a_n2804_13878.t27 74.6477
R15633 a_n2804_13878.n17 a_n2804_13878.t26 74.2899
R15634 a_n2804_13878.n14 a_n2804_13878.t0 74.2899
R15635 a_n2804_13878.n13 a_n2804_13878.t1 74.2899
R15636 a_n2804_13878.n16 a_n2804_13878.n15 70.6783
R15637 a_n2804_13878.n12 a_n2804_13878.n11 70.6783
R15638 a_n2804_13878.n18 a_n2804_13878.n10 15.7159
R15639 a_n2804_13878.n20 a_n2804_13878.n18 12.6495
R15640 a_n2804_13878.n18 a_n2804_13878.n17 8.38735
R15641 a_n2804_13878.n19 a_n2804_13878.t9 3.61217
R15642 a_n2804_13878.n19 a_n2804_13878.t18 3.61217
R15643 a_n2804_13878.n21 a_n2804_13878.t22 3.61217
R15644 a_n2804_13878.n21 a_n2804_13878.t8 3.61217
R15645 a_n2804_13878.n23 a_n2804_13878.t12 3.61217
R15646 a_n2804_13878.n23 a_n2804_13878.t13 3.61217
R15647 a_n2804_13878.n25 a_n2804_13878.t23 3.61217
R15648 a_n2804_13878.n25 a_n2804_13878.t24 3.61217
R15649 a_n2804_13878.n27 a_n2804_13878.t2 3.61217
R15650 a_n2804_13878.n27 a_n2804_13878.t14 3.61217
R15651 a_n2804_13878.n15 a_n2804_13878.t29 3.61217
R15652 a_n2804_13878.n15 a_n2804_13878.t30 3.61217
R15653 a_n2804_13878.n11 a_n2804_13878.t28 3.61217
R15654 a_n2804_13878.n11 a_n2804_13878.t31 3.61217
R15655 a_n2804_13878.n9 a_n2804_13878.t15 3.61217
R15656 a_n2804_13878.n9 a_n2804_13878.t3 3.61217
R15657 a_n2804_13878.n7 a_n2804_13878.t20 3.61217
R15658 a_n2804_13878.n7 a_n2804_13878.t5 3.61217
R15659 a_n2804_13878.n5 a_n2804_13878.t4 3.61217
R15660 a_n2804_13878.n5 a_n2804_13878.t7 3.61217
R15661 a_n2804_13878.n3 a_n2804_13878.t17 3.61217
R15662 a_n2804_13878.n3 a_n2804_13878.t10 3.61217
R15663 a_n2804_13878.n1 a_n2804_13878.t21 3.61217
R15664 a_n2804_13878.n1 a_n2804_13878.t11 3.61217
R15665 a_n2804_13878.n0 a_n2804_13878.t6 3.61217
R15666 a_n2804_13878.n0 a_n2804_13878.t16 3.61217
R15667 a_n2804_13878.n29 a_n2804_13878.t19 3.61217
R15668 a_n2804_13878.t25 a_n2804_13878.n29 3.61217
R15669 a_n2804_13878.n13 a_n2804_13878.n12 0.358259
R15670 a_n2804_13878.n16 a_n2804_13878.n14 0.358259
R15671 a_n2804_13878.n17 a_n2804_13878.n16 0.358259
R15672 a_n2804_13878.n28 a_n2804_13878.n26 0.358259
R15673 a_n2804_13878.n26 a_n2804_13878.n24 0.358259
R15674 a_n2804_13878.n24 a_n2804_13878.n22 0.358259
R15675 a_n2804_13878.n22 a_n2804_13878.n20 0.358259
R15676 a_n2804_13878.n4 a_n2804_13878.n2 0.146627
R15677 a_n2804_13878.n6 a_n2804_13878.n4 0.146627
R15678 a_n2804_13878.n8 a_n2804_13878.n6 0.146627
R15679 a_n2804_13878.n10 a_n2804_13878.n8 0.146627
R15680 a_n2804_13878.n14 a_n2804_13878.n13 0.101793
R15681 vdd.n315 vdd.n279 756.745
R15682 vdd.n260 vdd.n224 756.745
R15683 vdd.n217 vdd.n181 756.745
R15684 vdd.n162 vdd.n126 756.745
R15685 vdd.n120 vdd.n84 756.745
R15686 vdd.n65 vdd.n29 756.745
R15687 vdd.n2139 vdd.n2103 756.745
R15688 vdd.n2194 vdd.n2158 756.745
R15689 vdd.n2041 vdd.n2005 756.745
R15690 vdd.n2096 vdd.n2060 756.745
R15691 vdd.n1944 vdd.n1908 756.745
R15692 vdd.n1999 vdd.n1963 756.745
R15693 vdd.n1286 vdd.t197 640.208
R15694 vdd.n981 vdd.t242 640.208
R15695 vdd.n1290 vdd.t232 640.208
R15696 vdd.n972 vdd.t266 640.208
R15697 vdd.n867 vdd.t219 640.208
R15698 vdd.n2740 vdd.t260 640.208
R15699 vdd.n804 vdd.t208 640.208
R15700 vdd.n2737 vdd.t249 640.208
R15701 vdd.n768 vdd.t193 640.208
R15702 vdd.n1042 vdd.t256 640.208
R15703 vdd.n1603 vdd.t238 592.009
R15704 vdd.n1759 vdd.t253 592.009
R15705 vdd.n1795 vdd.t263 592.009
R15706 vdd.n2279 vdd.t223 592.009
R15707 vdd.n1219 vdd.t201 592.009
R15708 vdd.n1179 vdd.t205 592.009
R15709 vdd.n405 vdd.t235 592.009
R15710 vdd.n419 vdd.t211 592.009
R15711 vdd.n431 vdd.t226 592.009
R15712 vdd.n723 vdd.t229 592.009
R15713 vdd.n686 vdd.t246 592.009
R15714 vdd.n3285 vdd.t215 592.009
R15715 vdd.n316 vdd.n315 585
R15716 vdd.n314 vdd.n281 585
R15717 vdd.n313 vdd.n312 585
R15718 vdd.n284 vdd.n282 585
R15719 vdd.n307 vdd.n306 585
R15720 vdd.n305 vdd.n304 585
R15721 vdd.n288 vdd.n287 585
R15722 vdd.n299 vdd.n298 585
R15723 vdd.n297 vdd.n296 585
R15724 vdd.n292 vdd.n291 585
R15725 vdd.n261 vdd.n260 585
R15726 vdd.n259 vdd.n226 585
R15727 vdd.n258 vdd.n257 585
R15728 vdd.n229 vdd.n227 585
R15729 vdd.n252 vdd.n251 585
R15730 vdd.n250 vdd.n249 585
R15731 vdd.n233 vdd.n232 585
R15732 vdd.n244 vdd.n243 585
R15733 vdd.n242 vdd.n241 585
R15734 vdd.n237 vdd.n236 585
R15735 vdd.n218 vdd.n217 585
R15736 vdd.n216 vdd.n183 585
R15737 vdd.n215 vdd.n214 585
R15738 vdd.n186 vdd.n184 585
R15739 vdd.n209 vdd.n208 585
R15740 vdd.n207 vdd.n206 585
R15741 vdd.n190 vdd.n189 585
R15742 vdd.n201 vdd.n200 585
R15743 vdd.n199 vdd.n198 585
R15744 vdd.n194 vdd.n193 585
R15745 vdd.n163 vdd.n162 585
R15746 vdd.n161 vdd.n128 585
R15747 vdd.n160 vdd.n159 585
R15748 vdd.n131 vdd.n129 585
R15749 vdd.n154 vdd.n153 585
R15750 vdd.n152 vdd.n151 585
R15751 vdd.n135 vdd.n134 585
R15752 vdd.n146 vdd.n145 585
R15753 vdd.n144 vdd.n143 585
R15754 vdd.n139 vdd.n138 585
R15755 vdd.n121 vdd.n120 585
R15756 vdd.n119 vdd.n86 585
R15757 vdd.n118 vdd.n117 585
R15758 vdd.n89 vdd.n87 585
R15759 vdd.n112 vdd.n111 585
R15760 vdd.n110 vdd.n109 585
R15761 vdd.n93 vdd.n92 585
R15762 vdd.n104 vdd.n103 585
R15763 vdd.n102 vdd.n101 585
R15764 vdd.n97 vdd.n96 585
R15765 vdd.n66 vdd.n65 585
R15766 vdd.n64 vdd.n31 585
R15767 vdd.n63 vdd.n62 585
R15768 vdd.n34 vdd.n32 585
R15769 vdd.n57 vdd.n56 585
R15770 vdd.n55 vdd.n54 585
R15771 vdd.n38 vdd.n37 585
R15772 vdd.n49 vdd.n48 585
R15773 vdd.n47 vdd.n46 585
R15774 vdd.n42 vdd.n41 585
R15775 vdd.n2140 vdd.n2139 585
R15776 vdd.n2138 vdd.n2105 585
R15777 vdd.n2137 vdd.n2136 585
R15778 vdd.n2108 vdd.n2106 585
R15779 vdd.n2131 vdd.n2130 585
R15780 vdd.n2129 vdd.n2128 585
R15781 vdd.n2112 vdd.n2111 585
R15782 vdd.n2123 vdd.n2122 585
R15783 vdd.n2121 vdd.n2120 585
R15784 vdd.n2116 vdd.n2115 585
R15785 vdd.n2195 vdd.n2194 585
R15786 vdd.n2193 vdd.n2160 585
R15787 vdd.n2192 vdd.n2191 585
R15788 vdd.n2163 vdd.n2161 585
R15789 vdd.n2186 vdd.n2185 585
R15790 vdd.n2184 vdd.n2183 585
R15791 vdd.n2167 vdd.n2166 585
R15792 vdd.n2178 vdd.n2177 585
R15793 vdd.n2176 vdd.n2175 585
R15794 vdd.n2171 vdd.n2170 585
R15795 vdd.n2042 vdd.n2041 585
R15796 vdd.n2040 vdd.n2007 585
R15797 vdd.n2039 vdd.n2038 585
R15798 vdd.n2010 vdd.n2008 585
R15799 vdd.n2033 vdd.n2032 585
R15800 vdd.n2031 vdd.n2030 585
R15801 vdd.n2014 vdd.n2013 585
R15802 vdd.n2025 vdd.n2024 585
R15803 vdd.n2023 vdd.n2022 585
R15804 vdd.n2018 vdd.n2017 585
R15805 vdd.n2097 vdd.n2096 585
R15806 vdd.n2095 vdd.n2062 585
R15807 vdd.n2094 vdd.n2093 585
R15808 vdd.n2065 vdd.n2063 585
R15809 vdd.n2088 vdd.n2087 585
R15810 vdd.n2086 vdd.n2085 585
R15811 vdd.n2069 vdd.n2068 585
R15812 vdd.n2080 vdd.n2079 585
R15813 vdd.n2078 vdd.n2077 585
R15814 vdd.n2073 vdd.n2072 585
R15815 vdd.n1945 vdd.n1944 585
R15816 vdd.n1943 vdd.n1910 585
R15817 vdd.n1942 vdd.n1941 585
R15818 vdd.n1913 vdd.n1911 585
R15819 vdd.n1936 vdd.n1935 585
R15820 vdd.n1934 vdd.n1933 585
R15821 vdd.n1917 vdd.n1916 585
R15822 vdd.n1928 vdd.n1927 585
R15823 vdd.n1926 vdd.n1925 585
R15824 vdd.n1921 vdd.n1920 585
R15825 vdd.n2000 vdd.n1999 585
R15826 vdd.n1998 vdd.n1965 585
R15827 vdd.n1997 vdd.n1996 585
R15828 vdd.n1968 vdd.n1966 585
R15829 vdd.n1991 vdd.n1990 585
R15830 vdd.n1989 vdd.n1988 585
R15831 vdd.n1972 vdd.n1971 585
R15832 vdd.n1983 vdd.n1982 585
R15833 vdd.n1981 vdd.n1980 585
R15834 vdd.n1976 vdd.n1975 585
R15835 vdd.n445 vdd.n370 462.44
R15836 vdd.n3523 vdd.n372 462.44
R15837 vdd.n3418 vdd.n657 462.44
R15838 vdd.n3416 vdd.n660 462.44
R15839 vdd.n2274 vdd.n1502 462.44
R15840 vdd.n2277 vdd.n2276 462.44
R15841 vdd.n1830 vdd.n1600 462.44
R15842 vdd.n1827 vdd.n1598 462.44
R15843 vdd.n293 vdd.t99 329.043
R15844 vdd.n238 vdd.t185 329.043
R15845 vdd.n195 vdd.t81 329.043
R15846 vdd.n140 vdd.t175 329.043
R15847 vdd.n98 vdd.t145 329.043
R15848 vdd.n43 vdd.t130 329.043
R15849 vdd.n2117 vdd.t69 329.043
R15850 vdd.n2172 vdd.t148 329.043
R15851 vdd.n2019 vdd.t100 329.043
R15852 vdd.n2074 vdd.t139 329.043
R15853 vdd.n1922 vdd.t131 329.043
R15854 vdd.n1977 vdd.t147 329.043
R15855 vdd.n1603 vdd.t241 319.788
R15856 vdd.n1759 vdd.t255 319.788
R15857 vdd.n1795 vdd.t265 319.788
R15858 vdd.n2279 vdd.t224 319.788
R15859 vdd.n1219 vdd.t203 319.788
R15860 vdd.n1179 vdd.t206 319.788
R15861 vdd.n405 vdd.t236 319.788
R15862 vdd.n419 vdd.t213 319.788
R15863 vdd.n431 vdd.t227 319.788
R15864 vdd.n723 vdd.t231 319.788
R15865 vdd.n686 vdd.t248 319.788
R15866 vdd.n3285 vdd.t218 319.788
R15867 vdd.n1604 vdd.t240 303.69
R15868 vdd.n1760 vdd.t254 303.69
R15869 vdd.n1796 vdd.t264 303.69
R15870 vdd.n2280 vdd.t225 303.69
R15871 vdd.n1220 vdd.t204 303.69
R15872 vdd.n1180 vdd.t207 303.69
R15873 vdd.n406 vdd.t237 303.69
R15874 vdd.n420 vdd.t214 303.69
R15875 vdd.n432 vdd.t228 303.69
R15876 vdd.n724 vdd.t230 303.69
R15877 vdd.n687 vdd.t247 303.69
R15878 vdd.n3286 vdd.t217 303.69
R15879 vdd.n3007 vdd.n931 279.512
R15880 vdd.n3247 vdd.n778 279.512
R15881 vdd.n3184 vdd.n775 279.512
R15882 vdd.n2939 vdd.n2938 279.512
R15883 vdd.n2700 vdd.n969 279.512
R15884 vdd.n2631 vdd.n2630 279.512
R15885 vdd.n1326 vdd.n1325 279.512
R15886 vdd.n2425 vdd.n1109 279.512
R15887 vdd.n3163 vdd.n776 279.512
R15888 vdd.n3250 vdd.n3249 279.512
R15889 vdd.n2812 vdd.n2735 279.512
R15890 vdd.n2743 vdd.n927 279.512
R15891 vdd.n2628 vdd.n979 279.512
R15892 vdd.n977 vdd.n951 279.512
R15893 vdd.n1451 vdd.n1146 279.512
R15894 vdd.n1251 vdd.n1104 279.512
R15895 vdd.n2423 vdd.n1112 254.619
R15896 vdd.n756 vdd.n658 254.619
R15897 vdd.n3165 vdd.n776 185
R15898 vdd.n3248 vdd.n776 185
R15899 vdd.n3167 vdd.n3166 185
R15900 vdd.n3166 vdd.n774 185
R15901 vdd.n3168 vdd.n810 185
R15902 vdd.n3178 vdd.n810 185
R15903 vdd.n3169 vdd.n819 185
R15904 vdd.n819 vdd.n817 185
R15905 vdd.n3171 vdd.n3170 185
R15906 vdd.n3172 vdd.n3171 185
R15907 vdd.n3124 vdd.n818 185
R15908 vdd.n818 vdd.n814 185
R15909 vdd.n3123 vdd.n3122 185
R15910 vdd.n3122 vdd.n3121 185
R15911 vdd.n821 vdd.n820 185
R15912 vdd.n822 vdd.n821 185
R15913 vdd.n3114 vdd.n3113 185
R15914 vdd.n3115 vdd.n3114 185
R15915 vdd.n3112 vdd.n830 185
R15916 vdd.n835 vdd.n830 185
R15917 vdd.n3111 vdd.n3110 185
R15918 vdd.n3110 vdd.n3109 185
R15919 vdd.n832 vdd.n831 185
R15920 vdd.n841 vdd.n832 185
R15921 vdd.n3102 vdd.n3101 185
R15922 vdd.n3103 vdd.n3102 185
R15923 vdd.n3100 vdd.n842 185
R15924 vdd.n848 vdd.n842 185
R15925 vdd.n3099 vdd.n3098 185
R15926 vdd.n3098 vdd.n3097 185
R15927 vdd.n844 vdd.n843 185
R15928 vdd.n845 vdd.n844 185
R15929 vdd.n3090 vdd.n3089 185
R15930 vdd.n3091 vdd.n3090 185
R15931 vdd.n3088 vdd.n855 185
R15932 vdd.n855 vdd.n852 185
R15933 vdd.n3087 vdd.n3086 185
R15934 vdd.n3086 vdd.n3085 185
R15935 vdd.n857 vdd.n856 185
R15936 vdd.n858 vdd.n857 185
R15937 vdd.n3078 vdd.n3077 185
R15938 vdd.n3079 vdd.n3078 185
R15939 vdd.n3076 vdd.n866 185
R15940 vdd.n872 vdd.n866 185
R15941 vdd.n3075 vdd.n3074 185
R15942 vdd.n3074 vdd.n3073 185
R15943 vdd.n3064 vdd.n869 185
R15944 vdd.n879 vdd.n869 185
R15945 vdd.n3066 vdd.n3065 185
R15946 vdd.n3067 vdd.n3066 185
R15947 vdd.n3063 vdd.n880 185
R15948 vdd.n880 vdd.n876 185
R15949 vdd.n3062 vdd.n3061 185
R15950 vdd.n3061 vdd.n3060 185
R15951 vdd.n882 vdd.n881 185
R15952 vdd.n883 vdd.n882 185
R15953 vdd.n3053 vdd.n3052 185
R15954 vdd.n3054 vdd.n3053 185
R15955 vdd.n3051 vdd.n891 185
R15956 vdd.n896 vdd.n891 185
R15957 vdd.n3050 vdd.n3049 185
R15958 vdd.n3049 vdd.n3048 185
R15959 vdd.n893 vdd.n892 185
R15960 vdd.n902 vdd.n893 185
R15961 vdd.n3041 vdd.n3040 185
R15962 vdd.n3042 vdd.n3041 185
R15963 vdd.n3039 vdd.n903 185
R15964 vdd.n2915 vdd.n903 185
R15965 vdd.n3038 vdd.n3037 185
R15966 vdd.n3037 vdd.n3036 185
R15967 vdd.n905 vdd.n904 185
R15968 vdd.n2921 vdd.n905 185
R15969 vdd.n3029 vdd.n3028 185
R15970 vdd.n3030 vdd.n3029 185
R15971 vdd.n3027 vdd.n914 185
R15972 vdd.n914 vdd.n911 185
R15973 vdd.n3026 vdd.n3025 185
R15974 vdd.n3025 vdd.n3024 185
R15975 vdd.n916 vdd.n915 185
R15976 vdd.n917 vdd.n916 185
R15977 vdd.n3017 vdd.n3016 185
R15978 vdd.n3018 vdd.n3017 185
R15979 vdd.n3015 vdd.n925 185
R15980 vdd.n2933 vdd.n925 185
R15981 vdd.n3014 vdd.n3013 185
R15982 vdd.n3013 vdd.n3012 185
R15983 vdd.n927 vdd.n926 185
R15984 vdd.n928 vdd.n927 185
R15985 vdd.n2744 vdd.n2743 185
R15986 vdd.n2746 vdd.n2745 185
R15987 vdd.n2748 vdd.n2747 185
R15988 vdd.n2750 vdd.n2749 185
R15989 vdd.n2752 vdd.n2751 185
R15990 vdd.n2754 vdd.n2753 185
R15991 vdd.n2756 vdd.n2755 185
R15992 vdd.n2758 vdd.n2757 185
R15993 vdd.n2760 vdd.n2759 185
R15994 vdd.n2762 vdd.n2761 185
R15995 vdd.n2764 vdd.n2763 185
R15996 vdd.n2766 vdd.n2765 185
R15997 vdd.n2768 vdd.n2767 185
R15998 vdd.n2770 vdd.n2769 185
R15999 vdd.n2772 vdd.n2771 185
R16000 vdd.n2774 vdd.n2773 185
R16001 vdd.n2776 vdd.n2775 185
R16002 vdd.n2778 vdd.n2777 185
R16003 vdd.n2780 vdd.n2779 185
R16004 vdd.n2782 vdd.n2781 185
R16005 vdd.n2784 vdd.n2783 185
R16006 vdd.n2786 vdd.n2785 185
R16007 vdd.n2788 vdd.n2787 185
R16008 vdd.n2790 vdd.n2789 185
R16009 vdd.n2792 vdd.n2791 185
R16010 vdd.n2794 vdd.n2793 185
R16011 vdd.n2796 vdd.n2795 185
R16012 vdd.n2798 vdd.n2797 185
R16013 vdd.n2800 vdd.n2799 185
R16014 vdd.n2802 vdd.n2801 185
R16015 vdd.n2804 vdd.n2803 185
R16016 vdd.n2806 vdd.n2805 185
R16017 vdd.n2808 vdd.n2807 185
R16018 vdd.n2810 vdd.n2809 185
R16019 vdd.n2811 vdd.n2735 185
R16020 vdd.n3005 vdd.n2735 185
R16021 vdd.n3251 vdd.n3250 185
R16022 vdd.n3252 vdd.n767 185
R16023 vdd.n3254 vdd.n3253 185
R16024 vdd.n3256 vdd.n765 185
R16025 vdd.n3258 vdd.n3257 185
R16026 vdd.n3259 vdd.n764 185
R16027 vdd.n3261 vdd.n3260 185
R16028 vdd.n3263 vdd.n762 185
R16029 vdd.n3265 vdd.n3264 185
R16030 vdd.n3266 vdd.n761 185
R16031 vdd.n3268 vdd.n3267 185
R16032 vdd.n3270 vdd.n759 185
R16033 vdd.n3272 vdd.n3271 185
R16034 vdd.n3273 vdd.n758 185
R16035 vdd.n3275 vdd.n3274 185
R16036 vdd.n3277 vdd.n757 185
R16037 vdd.n3278 vdd.n754 185
R16038 vdd.n3281 vdd.n3280 185
R16039 vdd.n755 vdd.n753 185
R16040 vdd.n3137 vdd.n3136 185
R16041 vdd.n3139 vdd.n3138 185
R16042 vdd.n3141 vdd.n3133 185
R16043 vdd.n3143 vdd.n3142 185
R16044 vdd.n3144 vdd.n3132 185
R16045 vdd.n3146 vdd.n3145 185
R16046 vdd.n3148 vdd.n3130 185
R16047 vdd.n3150 vdd.n3149 185
R16048 vdd.n3151 vdd.n3129 185
R16049 vdd.n3153 vdd.n3152 185
R16050 vdd.n3155 vdd.n3127 185
R16051 vdd.n3157 vdd.n3156 185
R16052 vdd.n3158 vdd.n3126 185
R16053 vdd.n3160 vdd.n3159 185
R16054 vdd.n3162 vdd.n3125 185
R16055 vdd.n3164 vdd.n3163 185
R16056 vdd.n3163 vdd.n756 185
R16057 vdd.n3249 vdd.n771 185
R16058 vdd.n3249 vdd.n3248 185
R16059 vdd.n2866 vdd.n773 185
R16060 vdd.n774 vdd.n773 185
R16061 vdd.n2867 vdd.n809 185
R16062 vdd.n3178 vdd.n809 185
R16063 vdd.n2869 vdd.n2868 185
R16064 vdd.n2868 vdd.n817 185
R16065 vdd.n2870 vdd.n816 185
R16066 vdd.n3172 vdd.n816 185
R16067 vdd.n2872 vdd.n2871 185
R16068 vdd.n2871 vdd.n814 185
R16069 vdd.n2873 vdd.n824 185
R16070 vdd.n3121 vdd.n824 185
R16071 vdd.n2875 vdd.n2874 185
R16072 vdd.n2874 vdd.n822 185
R16073 vdd.n2876 vdd.n829 185
R16074 vdd.n3115 vdd.n829 185
R16075 vdd.n2878 vdd.n2877 185
R16076 vdd.n2877 vdd.n835 185
R16077 vdd.n2879 vdd.n834 185
R16078 vdd.n3109 vdd.n834 185
R16079 vdd.n2881 vdd.n2880 185
R16080 vdd.n2880 vdd.n841 185
R16081 vdd.n2882 vdd.n840 185
R16082 vdd.n3103 vdd.n840 185
R16083 vdd.n2884 vdd.n2883 185
R16084 vdd.n2883 vdd.n848 185
R16085 vdd.n2885 vdd.n847 185
R16086 vdd.n3097 vdd.n847 185
R16087 vdd.n2887 vdd.n2886 185
R16088 vdd.n2886 vdd.n845 185
R16089 vdd.n2888 vdd.n854 185
R16090 vdd.n3091 vdd.n854 185
R16091 vdd.n2890 vdd.n2889 185
R16092 vdd.n2889 vdd.n852 185
R16093 vdd.n2891 vdd.n860 185
R16094 vdd.n3085 vdd.n860 185
R16095 vdd.n2893 vdd.n2892 185
R16096 vdd.n2892 vdd.n858 185
R16097 vdd.n2894 vdd.n865 185
R16098 vdd.n3079 vdd.n865 185
R16099 vdd.n2896 vdd.n2895 185
R16100 vdd.n2895 vdd.n872 185
R16101 vdd.n2897 vdd.n871 185
R16102 vdd.n3073 vdd.n871 185
R16103 vdd.n2899 vdd.n2898 185
R16104 vdd.n2898 vdd.n879 185
R16105 vdd.n2900 vdd.n878 185
R16106 vdd.n3067 vdd.n878 185
R16107 vdd.n2902 vdd.n2901 185
R16108 vdd.n2901 vdd.n876 185
R16109 vdd.n2903 vdd.n885 185
R16110 vdd.n3060 vdd.n885 185
R16111 vdd.n2905 vdd.n2904 185
R16112 vdd.n2904 vdd.n883 185
R16113 vdd.n2906 vdd.n890 185
R16114 vdd.n3054 vdd.n890 185
R16115 vdd.n2908 vdd.n2907 185
R16116 vdd.n2907 vdd.n896 185
R16117 vdd.n2909 vdd.n895 185
R16118 vdd.n3048 vdd.n895 185
R16119 vdd.n2911 vdd.n2910 185
R16120 vdd.n2910 vdd.n902 185
R16121 vdd.n2912 vdd.n901 185
R16122 vdd.n3042 vdd.n901 185
R16123 vdd.n2914 vdd.n2913 185
R16124 vdd.n2915 vdd.n2914 185
R16125 vdd.n2815 vdd.n907 185
R16126 vdd.n3036 vdd.n907 185
R16127 vdd.n2923 vdd.n2922 185
R16128 vdd.n2922 vdd.n2921 185
R16129 vdd.n2924 vdd.n913 185
R16130 vdd.n3030 vdd.n913 185
R16131 vdd.n2926 vdd.n2925 185
R16132 vdd.n2925 vdd.n911 185
R16133 vdd.n2927 vdd.n919 185
R16134 vdd.n3024 vdd.n919 185
R16135 vdd.n2929 vdd.n2928 185
R16136 vdd.n2928 vdd.n917 185
R16137 vdd.n2930 vdd.n924 185
R16138 vdd.n3018 vdd.n924 185
R16139 vdd.n2932 vdd.n2931 185
R16140 vdd.n2933 vdd.n2932 185
R16141 vdd.n2814 vdd.n930 185
R16142 vdd.n3012 vdd.n930 185
R16143 vdd.n2813 vdd.n2812 185
R16144 vdd.n2812 vdd.n928 185
R16145 vdd.n2274 vdd.n2273 185
R16146 vdd.n2275 vdd.n2274 185
R16147 vdd.n1503 vdd.n1501 185
R16148 vdd.n1501 vdd.n1500 185
R16149 vdd.n2269 vdd.n2268 185
R16150 vdd.n2268 vdd.n2267 185
R16151 vdd.n1506 vdd.n1505 185
R16152 vdd.n1507 vdd.n1506 185
R16153 vdd.n2256 vdd.n2255 185
R16154 vdd.n2257 vdd.n2256 185
R16155 vdd.n1515 vdd.n1514 185
R16156 vdd.n2248 vdd.n1514 185
R16157 vdd.n2251 vdd.n2250 185
R16158 vdd.n2250 vdd.n2249 185
R16159 vdd.n1518 vdd.n1517 185
R16160 vdd.n1524 vdd.n1518 185
R16161 vdd.n2239 vdd.n2238 185
R16162 vdd.n2240 vdd.n2239 185
R16163 vdd.n1526 vdd.n1525 185
R16164 vdd.n2231 vdd.n1525 185
R16165 vdd.n2234 vdd.n2233 185
R16166 vdd.n2233 vdd.n2232 185
R16167 vdd.n1529 vdd.n1528 185
R16168 vdd.n1530 vdd.n1529 185
R16169 vdd.n2222 vdd.n2221 185
R16170 vdd.n2223 vdd.n2222 185
R16171 vdd.n1538 vdd.n1537 185
R16172 vdd.n1537 vdd.n1536 185
R16173 vdd.n2217 vdd.n2216 185
R16174 vdd.n2216 vdd.n2215 185
R16175 vdd.n1541 vdd.n1540 185
R16176 vdd.n1547 vdd.n1541 185
R16177 vdd.n2206 vdd.n2205 185
R16178 vdd.n2207 vdd.n2206 185
R16179 vdd.n1549 vdd.n1548 185
R16180 vdd.n1903 vdd.n1548 185
R16181 vdd.n1906 vdd.n1905 185
R16182 vdd.n1905 vdd.n1904 185
R16183 vdd.n1552 vdd.n1551 185
R16184 vdd.n1559 vdd.n1552 185
R16185 vdd.n1894 vdd.n1893 185
R16186 vdd.n1895 vdd.n1894 185
R16187 vdd.n1561 vdd.n1560 185
R16188 vdd.n1560 vdd.n1558 185
R16189 vdd.n1889 vdd.n1888 185
R16190 vdd.n1888 vdd.n1887 185
R16191 vdd.n1564 vdd.n1563 185
R16192 vdd.n1565 vdd.n1564 185
R16193 vdd.n1878 vdd.n1877 185
R16194 vdd.n1879 vdd.n1878 185
R16195 vdd.n1572 vdd.n1571 185
R16196 vdd.n1870 vdd.n1571 185
R16197 vdd.n1873 vdd.n1872 185
R16198 vdd.n1872 vdd.n1871 185
R16199 vdd.n1575 vdd.n1574 185
R16200 vdd.n1581 vdd.n1575 185
R16201 vdd.n1861 vdd.n1860 185
R16202 vdd.n1862 vdd.n1861 185
R16203 vdd.n1583 vdd.n1582 185
R16204 vdd.n1853 vdd.n1582 185
R16205 vdd.n1856 vdd.n1855 185
R16206 vdd.n1855 vdd.n1854 185
R16207 vdd.n1586 vdd.n1585 185
R16208 vdd.n1587 vdd.n1586 185
R16209 vdd.n1844 vdd.n1843 185
R16210 vdd.n1845 vdd.n1844 185
R16211 vdd.n1595 vdd.n1594 185
R16212 vdd.n1594 vdd.n1593 185
R16213 vdd.n1839 vdd.n1838 185
R16214 vdd.n1838 vdd.n1837 185
R16215 vdd.n1598 vdd.n1597 185
R16216 vdd.n1599 vdd.n1598 185
R16217 vdd.n1827 vdd.n1826 185
R16218 vdd.n1825 vdd.n1638 185
R16219 vdd.n1640 vdd.n1637 185
R16220 vdd.n1829 vdd.n1637 185
R16221 vdd.n1821 vdd.n1642 185
R16222 vdd.n1820 vdd.n1643 185
R16223 vdd.n1819 vdd.n1644 185
R16224 vdd.n1647 vdd.n1645 185
R16225 vdd.n1815 vdd.n1648 185
R16226 vdd.n1814 vdd.n1649 185
R16227 vdd.n1813 vdd.n1650 185
R16228 vdd.n1653 vdd.n1651 185
R16229 vdd.n1809 vdd.n1654 185
R16230 vdd.n1808 vdd.n1655 185
R16231 vdd.n1807 vdd.n1656 185
R16232 vdd.n1659 vdd.n1657 185
R16233 vdd.n1803 vdd.n1660 185
R16234 vdd.n1802 vdd.n1661 185
R16235 vdd.n1801 vdd.n1662 185
R16236 vdd.n1793 vdd.n1663 185
R16237 vdd.n1797 vdd.n1794 185
R16238 vdd.n1792 vdd.n1665 185
R16239 vdd.n1791 vdd.n1666 185
R16240 vdd.n1669 vdd.n1667 185
R16241 vdd.n1787 vdd.n1670 185
R16242 vdd.n1786 vdd.n1671 185
R16243 vdd.n1785 vdd.n1672 185
R16244 vdd.n1675 vdd.n1673 185
R16245 vdd.n1781 vdd.n1676 185
R16246 vdd.n1780 vdd.n1677 185
R16247 vdd.n1779 vdd.n1678 185
R16248 vdd.n1681 vdd.n1679 185
R16249 vdd.n1775 vdd.n1682 185
R16250 vdd.n1774 vdd.n1683 185
R16251 vdd.n1773 vdd.n1684 185
R16252 vdd.n1687 vdd.n1685 185
R16253 vdd.n1769 vdd.n1688 185
R16254 vdd.n1768 vdd.n1689 185
R16255 vdd.n1767 vdd.n1690 185
R16256 vdd.n1693 vdd.n1691 185
R16257 vdd.n1763 vdd.n1694 185
R16258 vdd.n1762 vdd.n1695 185
R16259 vdd.n1761 vdd.n1758 185
R16260 vdd.n1698 vdd.n1696 185
R16261 vdd.n1754 vdd.n1699 185
R16262 vdd.n1753 vdd.n1700 185
R16263 vdd.n1752 vdd.n1701 185
R16264 vdd.n1704 vdd.n1702 185
R16265 vdd.n1748 vdd.n1705 185
R16266 vdd.n1747 vdd.n1706 185
R16267 vdd.n1746 vdd.n1707 185
R16268 vdd.n1710 vdd.n1708 185
R16269 vdd.n1742 vdd.n1711 185
R16270 vdd.n1741 vdd.n1712 185
R16271 vdd.n1740 vdd.n1713 185
R16272 vdd.n1716 vdd.n1714 185
R16273 vdd.n1736 vdd.n1717 185
R16274 vdd.n1735 vdd.n1718 185
R16275 vdd.n1734 vdd.n1719 185
R16276 vdd.n1722 vdd.n1720 185
R16277 vdd.n1730 vdd.n1723 185
R16278 vdd.n1729 vdd.n1724 185
R16279 vdd.n1728 vdd.n1725 185
R16280 vdd.n1726 vdd.n1606 185
R16281 vdd.n1831 vdd.n1830 185
R16282 vdd.n1830 vdd.n1829 185
R16283 vdd.n2278 vdd.n2277 185
R16284 vdd.n2282 vdd.n1496 185
R16285 vdd.n1495 vdd.n1489 185
R16286 vdd.n1493 vdd.n1492 185
R16287 vdd.n1491 vdd.n1250 185
R16288 vdd.n2286 vdd.n1247 185
R16289 vdd.n2288 vdd.n2287 185
R16290 vdd.n2290 vdd.n1245 185
R16291 vdd.n2292 vdd.n2291 185
R16292 vdd.n2293 vdd.n1240 185
R16293 vdd.n2295 vdd.n2294 185
R16294 vdd.n2297 vdd.n1238 185
R16295 vdd.n2299 vdd.n2298 185
R16296 vdd.n2300 vdd.n1233 185
R16297 vdd.n2302 vdd.n2301 185
R16298 vdd.n2304 vdd.n1231 185
R16299 vdd.n2306 vdd.n2305 185
R16300 vdd.n2307 vdd.n1227 185
R16301 vdd.n2309 vdd.n2308 185
R16302 vdd.n2311 vdd.n1224 185
R16303 vdd.n2313 vdd.n2312 185
R16304 vdd.n1225 vdd.n1218 185
R16305 vdd.n2317 vdd.n1222 185
R16306 vdd.n2318 vdd.n1214 185
R16307 vdd.n2320 vdd.n2319 185
R16308 vdd.n2322 vdd.n1212 185
R16309 vdd.n2324 vdd.n2323 185
R16310 vdd.n2325 vdd.n1207 185
R16311 vdd.n2327 vdd.n2326 185
R16312 vdd.n2329 vdd.n1205 185
R16313 vdd.n2331 vdd.n2330 185
R16314 vdd.n2332 vdd.n1200 185
R16315 vdd.n2334 vdd.n2333 185
R16316 vdd.n2336 vdd.n1198 185
R16317 vdd.n2338 vdd.n2337 185
R16318 vdd.n2339 vdd.n1193 185
R16319 vdd.n2341 vdd.n2340 185
R16320 vdd.n2343 vdd.n1191 185
R16321 vdd.n2345 vdd.n2344 185
R16322 vdd.n2346 vdd.n1187 185
R16323 vdd.n2348 vdd.n2347 185
R16324 vdd.n2350 vdd.n1184 185
R16325 vdd.n2352 vdd.n2351 185
R16326 vdd.n1185 vdd.n1178 185
R16327 vdd.n2356 vdd.n1182 185
R16328 vdd.n2357 vdd.n1174 185
R16329 vdd.n2359 vdd.n2358 185
R16330 vdd.n2361 vdd.n1172 185
R16331 vdd.n2363 vdd.n2362 185
R16332 vdd.n2364 vdd.n1167 185
R16333 vdd.n2366 vdd.n2365 185
R16334 vdd.n2368 vdd.n1165 185
R16335 vdd.n2370 vdd.n2369 185
R16336 vdd.n2371 vdd.n1160 185
R16337 vdd.n2373 vdd.n2372 185
R16338 vdd.n2375 vdd.n1158 185
R16339 vdd.n2377 vdd.n2376 185
R16340 vdd.n2378 vdd.n1156 185
R16341 vdd.n2380 vdd.n2379 185
R16342 vdd.n2383 vdd.n2382 185
R16343 vdd.n2385 vdd.n2384 185
R16344 vdd.n2387 vdd.n1154 185
R16345 vdd.n2389 vdd.n2388 185
R16346 vdd.n1502 vdd.n1153 185
R16347 vdd.n2276 vdd.n1499 185
R16348 vdd.n2276 vdd.n2275 185
R16349 vdd.n1510 vdd.n1498 185
R16350 vdd.n1500 vdd.n1498 185
R16351 vdd.n2266 vdd.n2265 185
R16352 vdd.n2267 vdd.n2266 185
R16353 vdd.n1509 vdd.n1508 185
R16354 vdd.n1508 vdd.n1507 185
R16355 vdd.n2259 vdd.n2258 185
R16356 vdd.n2258 vdd.n2257 185
R16357 vdd.n1513 vdd.n1512 185
R16358 vdd.n2248 vdd.n1513 185
R16359 vdd.n2247 vdd.n2246 185
R16360 vdd.n2249 vdd.n2247 185
R16361 vdd.n1520 vdd.n1519 185
R16362 vdd.n1524 vdd.n1519 185
R16363 vdd.n2242 vdd.n2241 185
R16364 vdd.n2241 vdd.n2240 185
R16365 vdd.n1523 vdd.n1522 185
R16366 vdd.n2231 vdd.n1523 185
R16367 vdd.n2230 vdd.n2229 185
R16368 vdd.n2232 vdd.n2230 185
R16369 vdd.n1532 vdd.n1531 185
R16370 vdd.n1531 vdd.n1530 185
R16371 vdd.n2225 vdd.n2224 185
R16372 vdd.n2224 vdd.n2223 185
R16373 vdd.n1535 vdd.n1534 185
R16374 vdd.n1536 vdd.n1535 185
R16375 vdd.n2214 vdd.n2213 185
R16376 vdd.n2215 vdd.n2214 185
R16377 vdd.n1543 vdd.n1542 185
R16378 vdd.n1547 vdd.n1542 185
R16379 vdd.n2209 vdd.n2208 185
R16380 vdd.n2208 vdd.n2207 185
R16381 vdd.n1546 vdd.n1545 185
R16382 vdd.n1903 vdd.n1546 185
R16383 vdd.n1902 vdd.n1901 185
R16384 vdd.n1904 vdd.n1902 185
R16385 vdd.n1554 vdd.n1553 185
R16386 vdd.n1559 vdd.n1553 185
R16387 vdd.n1897 vdd.n1896 185
R16388 vdd.n1896 vdd.n1895 185
R16389 vdd.n1557 vdd.n1556 185
R16390 vdd.n1558 vdd.n1557 185
R16391 vdd.n1886 vdd.n1885 185
R16392 vdd.n1887 vdd.n1886 185
R16393 vdd.n1567 vdd.n1566 185
R16394 vdd.n1566 vdd.n1565 185
R16395 vdd.n1881 vdd.n1880 185
R16396 vdd.n1880 vdd.n1879 185
R16397 vdd.n1570 vdd.n1569 185
R16398 vdd.n1870 vdd.n1570 185
R16399 vdd.n1869 vdd.n1868 185
R16400 vdd.n1871 vdd.n1869 185
R16401 vdd.n1577 vdd.n1576 185
R16402 vdd.n1581 vdd.n1576 185
R16403 vdd.n1864 vdd.n1863 185
R16404 vdd.n1863 vdd.n1862 185
R16405 vdd.n1580 vdd.n1579 185
R16406 vdd.n1853 vdd.n1580 185
R16407 vdd.n1852 vdd.n1851 185
R16408 vdd.n1854 vdd.n1852 185
R16409 vdd.n1589 vdd.n1588 185
R16410 vdd.n1588 vdd.n1587 185
R16411 vdd.n1847 vdd.n1846 185
R16412 vdd.n1846 vdd.n1845 185
R16413 vdd.n1592 vdd.n1591 185
R16414 vdd.n1593 vdd.n1592 185
R16415 vdd.n1836 vdd.n1835 185
R16416 vdd.n1837 vdd.n1836 185
R16417 vdd.n1601 vdd.n1600 185
R16418 vdd.n1600 vdd.n1599 185
R16419 vdd.n971 vdd.n969 185
R16420 vdd.n2629 vdd.n969 185
R16421 vdd.n2551 vdd.n989 185
R16422 vdd.n989 vdd.n976 185
R16423 vdd.n2553 vdd.n2552 185
R16424 vdd.n2554 vdd.n2553 185
R16425 vdd.n2550 vdd.n988 185
R16426 vdd.n1370 vdd.n988 185
R16427 vdd.n2549 vdd.n2548 185
R16428 vdd.n2548 vdd.n2547 185
R16429 vdd.n991 vdd.n990 185
R16430 vdd.n992 vdd.n991 185
R16431 vdd.n2538 vdd.n2537 185
R16432 vdd.n2539 vdd.n2538 185
R16433 vdd.n2536 vdd.n1002 185
R16434 vdd.n1002 vdd.n999 185
R16435 vdd.n2535 vdd.n2534 185
R16436 vdd.n2534 vdd.n2533 185
R16437 vdd.n1004 vdd.n1003 185
R16438 vdd.n1396 vdd.n1004 185
R16439 vdd.n2526 vdd.n2525 185
R16440 vdd.n2527 vdd.n2526 185
R16441 vdd.n2524 vdd.n1012 185
R16442 vdd.n1017 vdd.n1012 185
R16443 vdd.n2523 vdd.n2522 185
R16444 vdd.n2522 vdd.n2521 185
R16445 vdd.n1014 vdd.n1013 185
R16446 vdd.n1023 vdd.n1014 185
R16447 vdd.n2514 vdd.n2513 185
R16448 vdd.n2515 vdd.n2514 185
R16449 vdd.n2512 vdd.n1024 185
R16450 vdd.n1408 vdd.n1024 185
R16451 vdd.n2511 vdd.n2510 185
R16452 vdd.n2510 vdd.n2509 185
R16453 vdd.n1026 vdd.n1025 185
R16454 vdd.n1027 vdd.n1026 185
R16455 vdd.n2502 vdd.n2501 185
R16456 vdd.n2503 vdd.n2502 185
R16457 vdd.n2500 vdd.n1036 185
R16458 vdd.n1036 vdd.n1033 185
R16459 vdd.n2499 vdd.n2498 185
R16460 vdd.n2498 vdd.n2497 185
R16461 vdd.n1038 vdd.n1037 185
R16462 vdd.n1047 vdd.n1038 185
R16463 vdd.n2489 vdd.n2488 185
R16464 vdd.n2490 vdd.n2489 185
R16465 vdd.n2487 vdd.n1048 185
R16466 vdd.n1054 vdd.n1048 185
R16467 vdd.n2486 vdd.n2485 185
R16468 vdd.n2485 vdd.n2484 185
R16469 vdd.n1050 vdd.n1049 185
R16470 vdd.n1051 vdd.n1050 185
R16471 vdd.n2477 vdd.n2476 185
R16472 vdd.n2478 vdd.n2477 185
R16473 vdd.n2475 vdd.n1061 185
R16474 vdd.n1061 vdd.n1058 185
R16475 vdd.n2474 vdd.n2473 185
R16476 vdd.n2473 vdd.n2472 185
R16477 vdd.n1063 vdd.n1062 185
R16478 vdd.n1064 vdd.n1063 185
R16479 vdd.n2465 vdd.n2464 185
R16480 vdd.n2466 vdd.n2465 185
R16481 vdd.n2463 vdd.n1072 185
R16482 vdd.n1077 vdd.n1072 185
R16483 vdd.n2462 vdd.n2461 185
R16484 vdd.n2461 vdd.n2460 185
R16485 vdd.n1074 vdd.n1073 185
R16486 vdd.n1083 vdd.n1074 185
R16487 vdd.n2453 vdd.n2452 185
R16488 vdd.n2454 vdd.n2453 185
R16489 vdd.n2451 vdd.n1084 185
R16490 vdd.n1090 vdd.n1084 185
R16491 vdd.n2450 vdd.n2449 185
R16492 vdd.n2449 vdd.n2448 185
R16493 vdd.n1086 vdd.n1085 185
R16494 vdd.n1087 vdd.n1086 185
R16495 vdd.n2441 vdd.n2440 185
R16496 vdd.n2442 vdd.n2441 185
R16497 vdd.n2439 vdd.n1097 185
R16498 vdd.n1097 vdd.n1094 185
R16499 vdd.n2438 vdd.n2437 185
R16500 vdd.n2437 vdd.n2436 185
R16501 vdd.n1099 vdd.n1098 185
R16502 vdd.n1108 vdd.n1099 185
R16503 vdd.n2429 vdd.n2428 185
R16504 vdd.n2430 vdd.n2429 185
R16505 vdd.n2427 vdd.n1109 185
R16506 vdd.n1109 vdd.n1105 185
R16507 vdd.n2426 vdd.n2425 185
R16508 vdd.n1111 vdd.n1110 185
R16509 vdd.n2422 vdd.n2421 185
R16510 vdd.n2423 vdd.n2422 185
R16511 vdd.n2420 vdd.n1147 185
R16512 vdd.n2419 vdd.n2418 185
R16513 vdd.n2417 vdd.n2416 185
R16514 vdd.n2415 vdd.n2414 185
R16515 vdd.n2413 vdd.n2412 185
R16516 vdd.n2411 vdd.n2410 185
R16517 vdd.n2409 vdd.n2408 185
R16518 vdd.n2407 vdd.n2406 185
R16519 vdd.n2405 vdd.n2404 185
R16520 vdd.n2403 vdd.n2402 185
R16521 vdd.n2401 vdd.n2400 185
R16522 vdd.n2399 vdd.n2398 185
R16523 vdd.n2397 vdd.n2396 185
R16524 vdd.n2395 vdd.n2394 185
R16525 vdd.n2393 vdd.n2392 185
R16526 vdd.n1292 vdd.n1148 185
R16527 vdd.n1294 vdd.n1293 185
R16528 vdd.n1296 vdd.n1295 185
R16529 vdd.n1298 vdd.n1297 185
R16530 vdd.n1300 vdd.n1299 185
R16531 vdd.n1302 vdd.n1301 185
R16532 vdd.n1304 vdd.n1303 185
R16533 vdd.n1306 vdd.n1305 185
R16534 vdd.n1308 vdd.n1307 185
R16535 vdd.n1310 vdd.n1309 185
R16536 vdd.n1312 vdd.n1311 185
R16537 vdd.n1314 vdd.n1313 185
R16538 vdd.n1316 vdd.n1315 185
R16539 vdd.n1318 vdd.n1317 185
R16540 vdd.n1321 vdd.n1320 185
R16541 vdd.n1323 vdd.n1322 185
R16542 vdd.n1325 vdd.n1324 185
R16543 vdd.n2632 vdd.n2631 185
R16544 vdd.n2634 vdd.n2633 185
R16545 vdd.n2636 vdd.n2635 185
R16546 vdd.n2639 vdd.n2638 185
R16547 vdd.n2641 vdd.n2640 185
R16548 vdd.n2643 vdd.n2642 185
R16549 vdd.n2645 vdd.n2644 185
R16550 vdd.n2647 vdd.n2646 185
R16551 vdd.n2649 vdd.n2648 185
R16552 vdd.n2651 vdd.n2650 185
R16553 vdd.n2653 vdd.n2652 185
R16554 vdd.n2655 vdd.n2654 185
R16555 vdd.n2657 vdd.n2656 185
R16556 vdd.n2659 vdd.n2658 185
R16557 vdd.n2661 vdd.n2660 185
R16558 vdd.n2663 vdd.n2662 185
R16559 vdd.n2665 vdd.n2664 185
R16560 vdd.n2667 vdd.n2666 185
R16561 vdd.n2669 vdd.n2668 185
R16562 vdd.n2671 vdd.n2670 185
R16563 vdd.n2673 vdd.n2672 185
R16564 vdd.n2675 vdd.n2674 185
R16565 vdd.n2677 vdd.n2676 185
R16566 vdd.n2679 vdd.n2678 185
R16567 vdd.n2681 vdd.n2680 185
R16568 vdd.n2683 vdd.n2682 185
R16569 vdd.n2685 vdd.n2684 185
R16570 vdd.n2687 vdd.n2686 185
R16571 vdd.n2689 vdd.n2688 185
R16572 vdd.n2691 vdd.n2690 185
R16573 vdd.n2693 vdd.n2692 185
R16574 vdd.n2695 vdd.n2694 185
R16575 vdd.n2697 vdd.n2696 185
R16576 vdd.n2698 vdd.n970 185
R16577 vdd.n2700 vdd.n2699 185
R16578 vdd.n2701 vdd.n2700 185
R16579 vdd.n2630 vdd.n974 185
R16580 vdd.n2630 vdd.n2629 185
R16581 vdd.n1368 vdd.n975 185
R16582 vdd.n976 vdd.n975 185
R16583 vdd.n1369 vdd.n986 185
R16584 vdd.n2554 vdd.n986 185
R16585 vdd.n1372 vdd.n1371 185
R16586 vdd.n1371 vdd.n1370 185
R16587 vdd.n1373 vdd.n993 185
R16588 vdd.n2547 vdd.n993 185
R16589 vdd.n1375 vdd.n1374 185
R16590 vdd.n1374 vdd.n992 185
R16591 vdd.n1376 vdd.n1000 185
R16592 vdd.n2539 vdd.n1000 185
R16593 vdd.n1378 vdd.n1377 185
R16594 vdd.n1377 vdd.n999 185
R16595 vdd.n1379 vdd.n1005 185
R16596 vdd.n2533 vdd.n1005 185
R16597 vdd.n1398 vdd.n1397 185
R16598 vdd.n1397 vdd.n1396 185
R16599 vdd.n1399 vdd.n1010 185
R16600 vdd.n2527 vdd.n1010 185
R16601 vdd.n1401 vdd.n1400 185
R16602 vdd.n1400 vdd.n1017 185
R16603 vdd.n1402 vdd.n1015 185
R16604 vdd.n2521 vdd.n1015 185
R16605 vdd.n1404 vdd.n1403 185
R16606 vdd.n1403 vdd.n1023 185
R16607 vdd.n1405 vdd.n1021 185
R16608 vdd.n2515 vdd.n1021 185
R16609 vdd.n1407 vdd.n1406 185
R16610 vdd.n1408 vdd.n1407 185
R16611 vdd.n1367 vdd.n1028 185
R16612 vdd.n2509 vdd.n1028 185
R16613 vdd.n1366 vdd.n1365 185
R16614 vdd.n1365 vdd.n1027 185
R16615 vdd.n1364 vdd.n1034 185
R16616 vdd.n2503 vdd.n1034 185
R16617 vdd.n1363 vdd.n1362 185
R16618 vdd.n1362 vdd.n1033 185
R16619 vdd.n1361 vdd.n1039 185
R16620 vdd.n2497 vdd.n1039 185
R16621 vdd.n1360 vdd.n1359 185
R16622 vdd.n1359 vdd.n1047 185
R16623 vdd.n1358 vdd.n1045 185
R16624 vdd.n2490 vdd.n1045 185
R16625 vdd.n1357 vdd.n1356 185
R16626 vdd.n1356 vdd.n1054 185
R16627 vdd.n1355 vdd.n1052 185
R16628 vdd.n2484 vdd.n1052 185
R16629 vdd.n1354 vdd.n1353 185
R16630 vdd.n1353 vdd.n1051 185
R16631 vdd.n1352 vdd.n1059 185
R16632 vdd.n2478 vdd.n1059 185
R16633 vdd.n1351 vdd.n1350 185
R16634 vdd.n1350 vdd.n1058 185
R16635 vdd.n1349 vdd.n1065 185
R16636 vdd.n2472 vdd.n1065 185
R16637 vdd.n1348 vdd.n1347 185
R16638 vdd.n1347 vdd.n1064 185
R16639 vdd.n1346 vdd.n1070 185
R16640 vdd.n2466 vdd.n1070 185
R16641 vdd.n1345 vdd.n1344 185
R16642 vdd.n1344 vdd.n1077 185
R16643 vdd.n1343 vdd.n1075 185
R16644 vdd.n2460 vdd.n1075 185
R16645 vdd.n1342 vdd.n1341 185
R16646 vdd.n1341 vdd.n1083 185
R16647 vdd.n1340 vdd.n1081 185
R16648 vdd.n2454 vdd.n1081 185
R16649 vdd.n1339 vdd.n1338 185
R16650 vdd.n1338 vdd.n1090 185
R16651 vdd.n1337 vdd.n1088 185
R16652 vdd.n2448 vdd.n1088 185
R16653 vdd.n1336 vdd.n1335 185
R16654 vdd.n1335 vdd.n1087 185
R16655 vdd.n1334 vdd.n1095 185
R16656 vdd.n2442 vdd.n1095 185
R16657 vdd.n1333 vdd.n1332 185
R16658 vdd.n1332 vdd.n1094 185
R16659 vdd.n1331 vdd.n1100 185
R16660 vdd.n2436 vdd.n1100 185
R16661 vdd.n1330 vdd.n1329 185
R16662 vdd.n1329 vdd.n1108 185
R16663 vdd.n1328 vdd.n1106 185
R16664 vdd.n2430 vdd.n1106 185
R16665 vdd.n1327 vdd.n1326 185
R16666 vdd.n1326 vdd.n1105 185
R16667 vdd.n370 vdd.n369 185
R16668 vdd.n3526 vdd.n370 185
R16669 vdd.n3529 vdd.n3528 185
R16670 vdd.n3528 vdd.n3527 185
R16671 vdd.n3530 vdd.n364 185
R16672 vdd.n364 vdd.n363 185
R16673 vdd.n3532 vdd.n3531 185
R16674 vdd.n3533 vdd.n3532 185
R16675 vdd.n359 vdd.n358 185
R16676 vdd.n3534 vdd.n359 185
R16677 vdd.n3537 vdd.n3536 185
R16678 vdd.n3536 vdd.n3535 185
R16679 vdd.n3538 vdd.n353 185
R16680 vdd.n3508 vdd.n353 185
R16681 vdd.n3540 vdd.n3539 185
R16682 vdd.n3541 vdd.n3540 185
R16683 vdd.n348 vdd.n347 185
R16684 vdd.n3542 vdd.n348 185
R16685 vdd.n3545 vdd.n3544 185
R16686 vdd.n3544 vdd.n3543 185
R16687 vdd.n3546 vdd.n342 185
R16688 vdd.n349 vdd.n342 185
R16689 vdd.n3548 vdd.n3547 185
R16690 vdd.n3549 vdd.n3548 185
R16691 vdd.n338 vdd.n337 185
R16692 vdd.n3550 vdd.n338 185
R16693 vdd.n3553 vdd.n3552 185
R16694 vdd.n3552 vdd.n3551 185
R16695 vdd.n3554 vdd.n333 185
R16696 vdd.n333 vdd.n332 185
R16697 vdd.n3556 vdd.n3555 185
R16698 vdd.n3557 vdd.n3556 185
R16699 vdd.n327 vdd.n325 185
R16700 vdd.n3558 vdd.n327 185
R16701 vdd.n3561 vdd.n3560 185
R16702 vdd.n3560 vdd.n3559 185
R16703 vdd.n326 vdd.n324 185
R16704 vdd.n328 vdd.n326 185
R16705 vdd.n3484 vdd.n3483 185
R16706 vdd.n3485 vdd.n3484 185
R16707 vdd.n615 vdd.n614 185
R16708 vdd.n614 vdd.n613 185
R16709 vdd.n3479 vdd.n3478 185
R16710 vdd.n3478 vdd.n3477 185
R16711 vdd.n618 vdd.n617 185
R16712 vdd.n624 vdd.n618 185
R16713 vdd.n3465 vdd.n3464 185
R16714 vdd.n3466 vdd.n3465 185
R16715 vdd.n626 vdd.n625 185
R16716 vdd.n3457 vdd.n625 185
R16717 vdd.n3460 vdd.n3459 185
R16718 vdd.n3459 vdd.n3458 185
R16719 vdd.n629 vdd.n628 185
R16720 vdd.n636 vdd.n629 185
R16721 vdd.n3448 vdd.n3447 185
R16722 vdd.n3449 vdd.n3448 185
R16723 vdd.n638 vdd.n637 185
R16724 vdd.n637 vdd.n635 185
R16725 vdd.n3443 vdd.n3442 185
R16726 vdd.n3442 vdd.n3441 185
R16727 vdd.n641 vdd.n640 185
R16728 vdd.n642 vdd.n641 185
R16729 vdd.n3432 vdd.n3431 185
R16730 vdd.n3433 vdd.n3432 185
R16731 vdd.n650 vdd.n649 185
R16732 vdd.n649 vdd.n648 185
R16733 vdd.n3427 vdd.n3426 185
R16734 vdd.n3426 vdd.n3425 185
R16735 vdd.n653 vdd.n652 185
R16736 vdd.n659 vdd.n653 185
R16737 vdd.n3416 vdd.n3415 185
R16738 vdd.n3417 vdd.n3416 185
R16739 vdd.n3412 vdd.n660 185
R16740 vdd.n3411 vdd.n3410 185
R16741 vdd.n3408 vdd.n662 185
R16742 vdd.n3408 vdd.n658 185
R16743 vdd.n3407 vdd.n3406 185
R16744 vdd.n3405 vdd.n3404 185
R16745 vdd.n3403 vdd.n3402 185
R16746 vdd.n3401 vdd.n3400 185
R16747 vdd.n3399 vdd.n668 185
R16748 vdd.n3397 vdd.n3396 185
R16749 vdd.n3395 vdd.n669 185
R16750 vdd.n3394 vdd.n3393 185
R16751 vdd.n3391 vdd.n674 185
R16752 vdd.n3389 vdd.n3388 185
R16753 vdd.n3387 vdd.n675 185
R16754 vdd.n3386 vdd.n3385 185
R16755 vdd.n3383 vdd.n680 185
R16756 vdd.n3381 vdd.n3380 185
R16757 vdd.n3379 vdd.n681 185
R16758 vdd.n3378 vdd.n3377 185
R16759 vdd.n3375 vdd.n688 185
R16760 vdd.n3373 vdd.n3372 185
R16761 vdd.n3371 vdd.n689 185
R16762 vdd.n3370 vdd.n3369 185
R16763 vdd.n3367 vdd.n694 185
R16764 vdd.n3365 vdd.n3364 185
R16765 vdd.n3363 vdd.n695 185
R16766 vdd.n3362 vdd.n3361 185
R16767 vdd.n3359 vdd.n700 185
R16768 vdd.n3357 vdd.n3356 185
R16769 vdd.n3355 vdd.n701 185
R16770 vdd.n3354 vdd.n3353 185
R16771 vdd.n3351 vdd.n706 185
R16772 vdd.n3349 vdd.n3348 185
R16773 vdd.n3347 vdd.n707 185
R16774 vdd.n3346 vdd.n3345 185
R16775 vdd.n3343 vdd.n712 185
R16776 vdd.n3341 vdd.n3340 185
R16777 vdd.n3339 vdd.n713 185
R16778 vdd.n3338 vdd.n3337 185
R16779 vdd.n3335 vdd.n718 185
R16780 vdd.n3333 vdd.n3332 185
R16781 vdd.n3331 vdd.n719 185
R16782 vdd.n728 vdd.n722 185
R16783 vdd.n3327 vdd.n3326 185
R16784 vdd.n3324 vdd.n726 185
R16785 vdd.n3323 vdd.n3322 185
R16786 vdd.n3321 vdd.n3320 185
R16787 vdd.n3319 vdd.n732 185
R16788 vdd.n3317 vdd.n3316 185
R16789 vdd.n3315 vdd.n733 185
R16790 vdd.n3314 vdd.n3313 185
R16791 vdd.n3311 vdd.n738 185
R16792 vdd.n3309 vdd.n3308 185
R16793 vdd.n3307 vdd.n739 185
R16794 vdd.n3306 vdd.n3305 185
R16795 vdd.n3303 vdd.n744 185
R16796 vdd.n3301 vdd.n3300 185
R16797 vdd.n3299 vdd.n745 185
R16798 vdd.n3298 vdd.n3297 185
R16799 vdd.n3295 vdd.n3294 185
R16800 vdd.n3293 vdd.n3292 185
R16801 vdd.n3291 vdd.n3290 185
R16802 vdd.n3289 vdd.n3288 185
R16803 vdd.n3284 vdd.n657 185
R16804 vdd.n658 vdd.n657 185
R16805 vdd.n3523 vdd.n3522 185
R16806 vdd.n599 vdd.n404 185
R16807 vdd.n598 vdd.n597 185
R16808 vdd.n596 vdd.n595 185
R16809 vdd.n594 vdd.n409 185
R16810 vdd.n590 vdd.n589 185
R16811 vdd.n588 vdd.n587 185
R16812 vdd.n586 vdd.n585 185
R16813 vdd.n584 vdd.n411 185
R16814 vdd.n580 vdd.n579 185
R16815 vdd.n578 vdd.n577 185
R16816 vdd.n576 vdd.n575 185
R16817 vdd.n574 vdd.n413 185
R16818 vdd.n570 vdd.n569 185
R16819 vdd.n568 vdd.n567 185
R16820 vdd.n566 vdd.n565 185
R16821 vdd.n564 vdd.n415 185
R16822 vdd.n560 vdd.n559 185
R16823 vdd.n558 vdd.n557 185
R16824 vdd.n556 vdd.n555 185
R16825 vdd.n554 vdd.n417 185
R16826 vdd.n550 vdd.n549 185
R16827 vdd.n548 vdd.n547 185
R16828 vdd.n546 vdd.n545 185
R16829 vdd.n544 vdd.n421 185
R16830 vdd.n540 vdd.n539 185
R16831 vdd.n538 vdd.n537 185
R16832 vdd.n536 vdd.n535 185
R16833 vdd.n534 vdd.n423 185
R16834 vdd.n530 vdd.n529 185
R16835 vdd.n528 vdd.n527 185
R16836 vdd.n526 vdd.n525 185
R16837 vdd.n524 vdd.n425 185
R16838 vdd.n520 vdd.n519 185
R16839 vdd.n518 vdd.n517 185
R16840 vdd.n516 vdd.n515 185
R16841 vdd.n514 vdd.n427 185
R16842 vdd.n510 vdd.n509 185
R16843 vdd.n508 vdd.n507 185
R16844 vdd.n506 vdd.n505 185
R16845 vdd.n504 vdd.n429 185
R16846 vdd.n500 vdd.n499 185
R16847 vdd.n498 vdd.n497 185
R16848 vdd.n496 vdd.n495 185
R16849 vdd.n494 vdd.n433 185
R16850 vdd.n490 vdd.n489 185
R16851 vdd.n488 vdd.n487 185
R16852 vdd.n486 vdd.n485 185
R16853 vdd.n484 vdd.n435 185
R16854 vdd.n480 vdd.n479 185
R16855 vdd.n478 vdd.n477 185
R16856 vdd.n476 vdd.n475 185
R16857 vdd.n474 vdd.n437 185
R16858 vdd.n470 vdd.n469 185
R16859 vdd.n468 vdd.n467 185
R16860 vdd.n466 vdd.n465 185
R16861 vdd.n464 vdd.n439 185
R16862 vdd.n460 vdd.n459 185
R16863 vdd.n458 vdd.n457 185
R16864 vdd.n456 vdd.n455 185
R16865 vdd.n454 vdd.n441 185
R16866 vdd.n450 vdd.n449 185
R16867 vdd.n448 vdd.n447 185
R16868 vdd.n446 vdd.n445 185
R16869 vdd.n3519 vdd.n372 185
R16870 vdd.n3526 vdd.n372 185
R16871 vdd.n3518 vdd.n371 185
R16872 vdd.n3527 vdd.n371 185
R16873 vdd.n3517 vdd.n3516 185
R16874 vdd.n3516 vdd.n363 185
R16875 vdd.n602 vdd.n362 185
R16876 vdd.n3533 vdd.n362 185
R16877 vdd.n3512 vdd.n361 185
R16878 vdd.n3534 vdd.n361 185
R16879 vdd.n3511 vdd.n360 185
R16880 vdd.n3535 vdd.n360 185
R16881 vdd.n3510 vdd.n3509 185
R16882 vdd.n3509 vdd.n3508 185
R16883 vdd.n604 vdd.n352 185
R16884 vdd.n3541 vdd.n352 185
R16885 vdd.n3504 vdd.n351 185
R16886 vdd.n3542 vdd.n351 185
R16887 vdd.n3503 vdd.n350 185
R16888 vdd.n3543 vdd.n350 185
R16889 vdd.n3502 vdd.n3501 185
R16890 vdd.n3501 vdd.n349 185
R16891 vdd.n606 vdd.n341 185
R16892 vdd.n3549 vdd.n341 185
R16893 vdd.n3497 vdd.n340 185
R16894 vdd.n3550 vdd.n340 185
R16895 vdd.n3496 vdd.n339 185
R16896 vdd.n3551 vdd.n339 185
R16897 vdd.n3495 vdd.n3494 185
R16898 vdd.n3494 vdd.n332 185
R16899 vdd.n608 vdd.n331 185
R16900 vdd.n3557 vdd.n331 185
R16901 vdd.n3490 vdd.n330 185
R16902 vdd.n3558 vdd.n330 185
R16903 vdd.n3489 vdd.n329 185
R16904 vdd.n3559 vdd.n329 185
R16905 vdd.n3488 vdd.n3487 185
R16906 vdd.n3487 vdd.n328 185
R16907 vdd.n3486 vdd.n610 185
R16908 vdd.n3486 vdd.n3485 185
R16909 vdd.n3474 vdd.n612 185
R16910 vdd.n613 vdd.n612 185
R16911 vdd.n3476 vdd.n3475 185
R16912 vdd.n3477 vdd.n3476 185
R16913 vdd.n620 vdd.n619 185
R16914 vdd.n624 vdd.n619 185
R16915 vdd.n3468 vdd.n3467 185
R16916 vdd.n3467 vdd.n3466 185
R16917 vdd.n623 vdd.n622 185
R16918 vdd.n3457 vdd.n623 185
R16919 vdd.n3456 vdd.n3455 185
R16920 vdd.n3458 vdd.n3456 185
R16921 vdd.n631 vdd.n630 185
R16922 vdd.n636 vdd.n630 185
R16923 vdd.n3451 vdd.n3450 185
R16924 vdd.n3450 vdd.n3449 185
R16925 vdd.n634 vdd.n633 185
R16926 vdd.n635 vdd.n634 185
R16927 vdd.n3440 vdd.n3439 185
R16928 vdd.n3441 vdd.n3440 185
R16929 vdd.n644 vdd.n643 185
R16930 vdd.n643 vdd.n642 185
R16931 vdd.n3435 vdd.n3434 185
R16932 vdd.n3434 vdd.n3433 185
R16933 vdd.n647 vdd.n646 185
R16934 vdd.n648 vdd.n647 185
R16935 vdd.n3424 vdd.n3423 185
R16936 vdd.n3425 vdd.n3424 185
R16937 vdd.n655 vdd.n654 185
R16938 vdd.n659 vdd.n654 185
R16939 vdd.n3419 vdd.n3418 185
R16940 vdd.n3418 vdd.n3417 185
R16941 vdd.n3008 vdd.n3007 185
R16942 vdd.n933 vdd.n932 185
R16943 vdd.n3004 vdd.n3003 185
R16944 vdd.n3005 vdd.n3004 185
R16945 vdd.n3002 vdd.n2736 185
R16946 vdd.n3001 vdd.n3000 185
R16947 vdd.n2999 vdd.n2998 185
R16948 vdd.n2997 vdd.n2996 185
R16949 vdd.n2995 vdd.n2994 185
R16950 vdd.n2993 vdd.n2992 185
R16951 vdd.n2991 vdd.n2990 185
R16952 vdd.n2989 vdd.n2988 185
R16953 vdd.n2987 vdd.n2986 185
R16954 vdd.n2985 vdd.n2984 185
R16955 vdd.n2983 vdd.n2982 185
R16956 vdd.n2981 vdd.n2980 185
R16957 vdd.n2979 vdd.n2978 185
R16958 vdd.n2977 vdd.n2976 185
R16959 vdd.n2975 vdd.n2974 185
R16960 vdd.n2973 vdd.n2972 185
R16961 vdd.n2971 vdd.n2970 185
R16962 vdd.n2969 vdd.n2968 185
R16963 vdd.n2967 vdd.n2966 185
R16964 vdd.n2965 vdd.n2964 185
R16965 vdd.n2963 vdd.n2962 185
R16966 vdd.n2961 vdd.n2960 185
R16967 vdd.n2959 vdd.n2958 185
R16968 vdd.n2957 vdd.n2956 185
R16969 vdd.n2955 vdd.n2954 185
R16970 vdd.n2953 vdd.n2952 185
R16971 vdd.n2951 vdd.n2950 185
R16972 vdd.n2949 vdd.n2948 185
R16973 vdd.n2947 vdd.n2946 185
R16974 vdd.n2944 vdd.n2943 185
R16975 vdd.n2942 vdd.n2941 185
R16976 vdd.n2940 vdd.n2939 185
R16977 vdd.n3185 vdd.n3184 185
R16978 vdd.n3186 vdd.n803 185
R16979 vdd.n3188 vdd.n3187 185
R16980 vdd.n3190 vdd.n801 185
R16981 vdd.n3192 vdd.n3191 185
R16982 vdd.n3193 vdd.n800 185
R16983 vdd.n3195 vdd.n3194 185
R16984 vdd.n3197 vdd.n798 185
R16985 vdd.n3199 vdd.n3198 185
R16986 vdd.n3200 vdd.n797 185
R16987 vdd.n3202 vdd.n3201 185
R16988 vdd.n3204 vdd.n795 185
R16989 vdd.n3206 vdd.n3205 185
R16990 vdd.n3207 vdd.n794 185
R16991 vdd.n3209 vdd.n3208 185
R16992 vdd.n3211 vdd.n792 185
R16993 vdd.n3213 vdd.n3212 185
R16994 vdd.n3215 vdd.n791 185
R16995 vdd.n3217 vdd.n3216 185
R16996 vdd.n3219 vdd.n789 185
R16997 vdd.n3221 vdd.n3220 185
R16998 vdd.n3222 vdd.n788 185
R16999 vdd.n3224 vdd.n3223 185
R17000 vdd.n3226 vdd.n786 185
R17001 vdd.n3228 vdd.n3227 185
R17002 vdd.n3229 vdd.n785 185
R17003 vdd.n3231 vdd.n3230 185
R17004 vdd.n3233 vdd.n783 185
R17005 vdd.n3235 vdd.n3234 185
R17006 vdd.n3236 vdd.n782 185
R17007 vdd.n3238 vdd.n3237 185
R17008 vdd.n3240 vdd.n781 185
R17009 vdd.n3241 vdd.n780 185
R17010 vdd.n3244 vdd.n3243 185
R17011 vdd.n3245 vdd.n778 185
R17012 vdd.n778 vdd.n756 185
R17013 vdd.n3182 vdd.n775 185
R17014 vdd.n3248 vdd.n775 185
R17015 vdd.n3181 vdd.n3180 185
R17016 vdd.n3180 vdd.n774 185
R17017 vdd.n3179 vdd.n807 185
R17018 vdd.n3179 vdd.n3178 185
R17019 vdd.n2822 vdd.n808 185
R17020 vdd.n817 vdd.n808 185
R17021 vdd.n2823 vdd.n815 185
R17022 vdd.n3172 vdd.n815 185
R17023 vdd.n2825 vdd.n2824 185
R17024 vdd.n2824 vdd.n814 185
R17025 vdd.n2826 vdd.n823 185
R17026 vdd.n3121 vdd.n823 185
R17027 vdd.n2828 vdd.n2827 185
R17028 vdd.n2827 vdd.n822 185
R17029 vdd.n2829 vdd.n828 185
R17030 vdd.n3115 vdd.n828 185
R17031 vdd.n2831 vdd.n2830 185
R17032 vdd.n2830 vdd.n835 185
R17033 vdd.n2832 vdd.n833 185
R17034 vdd.n3109 vdd.n833 185
R17035 vdd.n2834 vdd.n2833 185
R17036 vdd.n2833 vdd.n841 185
R17037 vdd.n2835 vdd.n839 185
R17038 vdd.n3103 vdd.n839 185
R17039 vdd.n2837 vdd.n2836 185
R17040 vdd.n2836 vdd.n848 185
R17041 vdd.n2838 vdd.n846 185
R17042 vdd.n3097 vdd.n846 185
R17043 vdd.n2840 vdd.n2839 185
R17044 vdd.n2839 vdd.n845 185
R17045 vdd.n2841 vdd.n853 185
R17046 vdd.n3091 vdd.n853 185
R17047 vdd.n2843 vdd.n2842 185
R17048 vdd.n2842 vdd.n852 185
R17049 vdd.n2844 vdd.n859 185
R17050 vdd.n3085 vdd.n859 185
R17051 vdd.n2846 vdd.n2845 185
R17052 vdd.n2845 vdd.n858 185
R17053 vdd.n2847 vdd.n864 185
R17054 vdd.n3079 vdd.n864 185
R17055 vdd.n2849 vdd.n2848 185
R17056 vdd.n2848 vdd.n872 185
R17057 vdd.n2850 vdd.n870 185
R17058 vdd.n3073 vdd.n870 185
R17059 vdd.n2852 vdd.n2851 185
R17060 vdd.n2851 vdd.n879 185
R17061 vdd.n2853 vdd.n877 185
R17062 vdd.n3067 vdd.n877 185
R17063 vdd.n2855 vdd.n2854 185
R17064 vdd.n2854 vdd.n876 185
R17065 vdd.n2856 vdd.n884 185
R17066 vdd.n3060 vdd.n884 185
R17067 vdd.n2858 vdd.n2857 185
R17068 vdd.n2857 vdd.n883 185
R17069 vdd.n2859 vdd.n889 185
R17070 vdd.n3054 vdd.n889 185
R17071 vdd.n2861 vdd.n2860 185
R17072 vdd.n2860 vdd.n896 185
R17073 vdd.n2862 vdd.n894 185
R17074 vdd.n3048 vdd.n894 185
R17075 vdd.n2864 vdd.n2863 185
R17076 vdd.n2863 vdd.n902 185
R17077 vdd.n2865 vdd.n900 185
R17078 vdd.n3042 vdd.n900 185
R17079 vdd.n2917 vdd.n2916 185
R17080 vdd.n2916 vdd.n2915 185
R17081 vdd.n2918 vdd.n906 185
R17082 vdd.n3036 vdd.n906 185
R17083 vdd.n2920 vdd.n2919 185
R17084 vdd.n2921 vdd.n2920 185
R17085 vdd.n2821 vdd.n912 185
R17086 vdd.n3030 vdd.n912 185
R17087 vdd.n2820 vdd.n2819 185
R17088 vdd.n2819 vdd.n911 185
R17089 vdd.n2818 vdd.n918 185
R17090 vdd.n3024 vdd.n918 185
R17091 vdd.n2817 vdd.n2816 185
R17092 vdd.n2816 vdd.n917 185
R17093 vdd.n2739 vdd.n923 185
R17094 vdd.n3018 vdd.n923 185
R17095 vdd.n2935 vdd.n2934 185
R17096 vdd.n2934 vdd.n2933 185
R17097 vdd.n2936 vdd.n929 185
R17098 vdd.n3012 vdd.n929 185
R17099 vdd.n2938 vdd.n2937 185
R17100 vdd.n2938 vdd.n928 185
R17101 vdd.n3009 vdd.n931 185
R17102 vdd.n931 vdd.n928 185
R17103 vdd.n3011 vdd.n3010 185
R17104 vdd.n3012 vdd.n3011 185
R17105 vdd.n922 vdd.n921 185
R17106 vdd.n2933 vdd.n922 185
R17107 vdd.n3020 vdd.n3019 185
R17108 vdd.n3019 vdd.n3018 185
R17109 vdd.n3021 vdd.n920 185
R17110 vdd.n920 vdd.n917 185
R17111 vdd.n3023 vdd.n3022 185
R17112 vdd.n3024 vdd.n3023 185
R17113 vdd.n910 vdd.n909 185
R17114 vdd.n911 vdd.n910 185
R17115 vdd.n3032 vdd.n3031 185
R17116 vdd.n3031 vdd.n3030 185
R17117 vdd.n3033 vdd.n908 185
R17118 vdd.n2921 vdd.n908 185
R17119 vdd.n3035 vdd.n3034 185
R17120 vdd.n3036 vdd.n3035 185
R17121 vdd.n899 vdd.n898 185
R17122 vdd.n2915 vdd.n899 185
R17123 vdd.n3044 vdd.n3043 185
R17124 vdd.n3043 vdd.n3042 185
R17125 vdd.n3045 vdd.n897 185
R17126 vdd.n902 vdd.n897 185
R17127 vdd.n3047 vdd.n3046 185
R17128 vdd.n3048 vdd.n3047 185
R17129 vdd.n888 vdd.n887 185
R17130 vdd.n896 vdd.n888 185
R17131 vdd.n3056 vdd.n3055 185
R17132 vdd.n3055 vdd.n3054 185
R17133 vdd.n3057 vdd.n886 185
R17134 vdd.n886 vdd.n883 185
R17135 vdd.n3059 vdd.n3058 185
R17136 vdd.n3060 vdd.n3059 185
R17137 vdd.n875 vdd.n874 185
R17138 vdd.n876 vdd.n875 185
R17139 vdd.n3069 vdd.n3068 185
R17140 vdd.n3068 vdd.n3067 185
R17141 vdd.n3070 vdd.n873 185
R17142 vdd.n879 vdd.n873 185
R17143 vdd.n3072 vdd.n3071 185
R17144 vdd.n3073 vdd.n3072 185
R17145 vdd.n863 vdd.n862 185
R17146 vdd.n872 vdd.n863 185
R17147 vdd.n3081 vdd.n3080 185
R17148 vdd.n3080 vdd.n3079 185
R17149 vdd.n3082 vdd.n861 185
R17150 vdd.n861 vdd.n858 185
R17151 vdd.n3084 vdd.n3083 185
R17152 vdd.n3085 vdd.n3084 185
R17153 vdd.n851 vdd.n850 185
R17154 vdd.n852 vdd.n851 185
R17155 vdd.n3093 vdd.n3092 185
R17156 vdd.n3092 vdd.n3091 185
R17157 vdd.n3094 vdd.n849 185
R17158 vdd.n849 vdd.n845 185
R17159 vdd.n3096 vdd.n3095 185
R17160 vdd.n3097 vdd.n3096 185
R17161 vdd.n838 vdd.n837 185
R17162 vdd.n848 vdd.n838 185
R17163 vdd.n3105 vdd.n3104 185
R17164 vdd.n3104 vdd.n3103 185
R17165 vdd.n3106 vdd.n836 185
R17166 vdd.n841 vdd.n836 185
R17167 vdd.n3108 vdd.n3107 185
R17168 vdd.n3109 vdd.n3108 185
R17169 vdd.n827 vdd.n826 185
R17170 vdd.n835 vdd.n827 185
R17171 vdd.n3117 vdd.n3116 185
R17172 vdd.n3116 vdd.n3115 185
R17173 vdd.n3118 vdd.n825 185
R17174 vdd.n825 vdd.n822 185
R17175 vdd.n3120 vdd.n3119 185
R17176 vdd.n3121 vdd.n3120 185
R17177 vdd.n813 vdd.n812 185
R17178 vdd.n814 vdd.n813 185
R17179 vdd.n3174 vdd.n3173 185
R17180 vdd.n3173 vdd.n3172 185
R17181 vdd.n3175 vdd.n811 185
R17182 vdd.n817 vdd.n811 185
R17183 vdd.n3177 vdd.n3176 185
R17184 vdd.n3178 vdd.n3177 185
R17185 vdd.n779 vdd.n777 185
R17186 vdd.n777 vdd.n774 185
R17187 vdd.n3247 vdd.n3246 185
R17188 vdd.n3248 vdd.n3247 185
R17189 vdd.n2628 vdd.n2627 185
R17190 vdd.n2629 vdd.n2628 185
R17191 vdd.n980 vdd.n978 185
R17192 vdd.n978 vdd.n976 185
R17193 vdd.n2543 vdd.n987 185
R17194 vdd.n2554 vdd.n987 185
R17195 vdd.n2544 vdd.n996 185
R17196 vdd.n1370 vdd.n996 185
R17197 vdd.n2546 vdd.n2545 185
R17198 vdd.n2547 vdd.n2546 185
R17199 vdd.n2542 vdd.n995 185
R17200 vdd.n995 vdd.n992 185
R17201 vdd.n2541 vdd.n2540 185
R17202 vdd.n2540 vdd.n2539 185
R17203 vdd.n998 vdd.n997 185
R17204 vdd.n999 vdd.n998 185
R17205 vdd.n2532 vdd.n2531 185
R17206 vdd.n2533 vdd.n2532 185
R17207 vdd.n2530 vdd.n1007 185
R17208 vdd.n1396 vdd.n1007 185
R17209 vdd.n2529 vdd.n2528 185
R17210 vdd.n2528 vdd.n2527 185
R17211 vdd.n1009 vdd.n1008 185
R17212 vdd.n1017 vdd.n1009 185
R17213 vdd.n2520 vdd.n2519 185
R17214 vdd.n2521 vdd.n2520 185
R17215 vdd.n2518 vdd.n1018 185
R17216 vdd.n1023 vdd.n1018 185
R17217 vdd.n2517 vdd.n2516 185
R17218 vdd.n2516 vdd.n2515 185
R17219 vdd.n1020 vdd.n1019 185
R17220 vdd.n1408 vdd.n1020 185
R17221 vdd.n2508 vdd.n2507 185
R17222 vdd.n2509 vdd.n2508 185
R17223 vdd.n2506 vdd.n1030 185
R17224 vdd.n1030 vdd.n1027 185
R17225 vdd.n2505 vdd.n2504 185
R17226 vdd.n2504 vdd.n2503 185
R17227 vdd.n1032 vdd.n1031 185
R17228 vdd.n1033 vdd.n1032 185
R17229 vdd.n2496 vdd.n2495 185
R17230 vdd.n2497 vdd.n2496 185
R17231 vdd.n2493 vdd.n1041 185
R17232 vdd.n1047 vdd.n1041 185
R17233 vdd.n2492 vdd.n2491 185
R17234 vdd.n2491 vdd.n2490 185
R17235 vdd.n1044 vdd.n1043 185
R17236 vdd.n1054 vdd.n1044 185
R17237 vdd.n2483 vdd.n2482 185
R17238 vdd.n2484 vdd.n2483 185
R17239 vdd.n2481 vdd.n1055 185
R17240 vdd.n1055 vdd.n1051 185
R17241 vdd.n2480 vdd.n2479 185
R17242 vdd.n2479 vdd.n2478 185
R17243 vdd.n1057 vdd.n1056 185
R17244 vdd.n1058 vdd.n1057 185
R17245 vdd.n2471 vdd.n2470 185
R17246 vdd.n2472 vdd.n2471 185
R17247 vdd.n2469 vdd.n1067 185
R17248 vdd.n1067 vdd.n1064 185
R17249 vdd.n2468 vdd.n2467 185
R17250 vdd.n2467 vdd.n2466 185
R17251 vdd.n1069 vdd.n1068 185
R17252 vdd.n1077 vdd.n1069 185
R17253 vdd.n2459 vdd.n2458 185
R17254 vdd.n2460 vdd.n2459 185
R17255 vdd.n2457 vdd.n1078 185
R17256 vdd.n1083 vdd.n1078 185
R17257 vdd.n2456 vdd.n2455 185
R17258 vdd.n2455 vdd.n2454 185
R17259 vdd.n1080 vdd.n1079 185
R17260 vdd.n1090 vdd.n1080 185
R17261 vdd.n2447 vdd.n2446 185
R17262 vdd.n2448 vdd.n2447 185
R17263 vdd.n2445 vdd.n1091 185
R17264 vdd.n1091 vdd.n1087 185
R17265 vdd.n2444 vdd.n2443 185
R17266 vdd.n2443 vdd.n2442 185
R17267 vdd.n1093 vdd.n1092 185
R17268 vdd.n1094 vdd.n1093 185
R17269 vdd.n2435 vdd.n2434 185
R17270 vdd.n2436 vdd.n2435 185
R17271 vdd.n2433 vdd.n1102 185
R17272 vdd.n1108 vdd.n1102 185
R17273 vdd.n2432 vdd.n2431 185
R17274 vdd.n2431 vdd.n2430 185
R17275 vdd.n1104 vdd.n1103 185
R17276 vdd.n1105 vdd.n1104 185
R17277 vdd.n2559 vdd.n951 185
R17278 vdd.n2701 vdd.n951 185
R17279 vdd.n2561 vdd.n2560 185
R17280 vdd.n2563 vdd.n2562 185
R17281 vdd.n2565 vdd.n2564 185
R17282 vdd.n2567 vdd.n2566 185
R17283 vdd.n2569 vdd.n2568 185
R17284 vdd.n2571 vdd.n2570 185
R17285 vdd.n2573 vdd.n2572 185
R17286 vdd.n2575 vdd.n2574 185
R17287 vdd.n2577 vdd.n2576 185
R17288 vdd.n2579 vdd.n2578 185
R17289 vdd.n2581 vdd.n2580 185
R17290 vdd.n2583 vdd.n2582 185
R17291 vdd.n2585 vdd.n2584 185
R17292 vdd.n2587 vdd.n2586 185
R17293 vdd.n2589 vdd.n2588 185
R17294 vdd.n2591 vdd.n2590 185
R17295 vdd.n2593 vdd.n2592 185
R17296 vdd.n2595 vdd.n2594 185
R17297 vdd.n2597 vdd.n2596 185
R17298 vdd.n2599 vdd.n2598 185
R17299 vdd.n2601 vdd.n2600 185
R17300 vdd.n2603 vdd.n2602 185
R17301 vdd.n2605 vdd.n2604 185
R17302 vdd.n2607 vdd.n2606 185
R17303 vdd.n2609 vdd.n2608 185
R17304 vdd.n2611 vdd.n2610 185
R17305 vdd.n2613 vdd.n2612 185
R17306 vdd.n2615 vdd.n2614 185
R17307 vdd.n2617 vdd.n2616 185
R17308 vdd.n2619 vdd.n2618 185
R17309 vdd.n2621 vdd.n2620 185
R17310 vdd.n2623 vdd.n2622 185
R17311 vdd.n2625 vdd.n2624 185
R17312 vdd.n2626 vdd.n979 185
R17313 vdd.n2558 vdd.n977 185
R17314 vdd.n2629 vdd.n977 185
R17315 vdd.n2557 vdd.n2556 185
R17316 vdd.n2556 vdd.n976 185
R17317 vdd.n2555 vdd.n984 185
R17318 vdd.n2555 vdd.n2554 185
R17319 vdd.n1386 vdd.n985 185
R17320 vdd.n1370 vdd.n985 185
R17321 vdd.n1387 vdd.n994 185
R17322 vdd.n2547 vdd.n994 185
R17323 vdd.n1389 vdd.n1388 185
R17324 vdd.n1388 vdd.n992 185
R17325 vdd.n1390 vdd.n1001 185
R17326 vdd.n2539 vdd.n1001 185
R17327 vdd.n1392 vdd.n1391 185
R17328 vdd.n1391 vdd.n999 185
R17329 vdd.n1393 vdd.n1006 185
R17330 vdd.n2533 vdd.n1006 185
R17331 vdd.n1395 vdd.n1394 185
R17332 vdd.n1396 vdd.n1395 185
R17333 vdd.n1385 vdd.n1011 185
R17334 vdd.n2527 vdd.n1011 185
R17335 vdd.n1384 vdd.n1383 185
R17336 vdd.n1383 vdd.n1017 185
R17337 vdd.n1382 vdd.n1016 185
R17338 vdd.n2521 vdd.n1016 185
R17339 vdd.n1381 vdd.n1380 185
R17340 vdd.n1380 vdd.n1023 185
R17341 vdd.n1289 vdd.n1022 185
R17342 vdd.n2515 vdd.n1022 185
R17343 vdd.n1410 vdd.n1409 185
R17344 vdd.n1409 vdd.n1408 185
R17345 vdd.n1411 vdd.n1029 185
R17346 vdd.n2509 vdd.n1029 185
R17347 vdd.n1413 vdd.n1412 185
R17348 vdd.n1412 vdd.n1027 185
R17349 vdd.n1414 vdd.n1035 185
R17350 vdd.n2503 vdd.n1035 185
R17351 vdd.n1416 vdd.n1415 185
R17352 vdd.n1415 vdd.n1033 185
R17353 vdd.n1417 vdd.n1040 185
R17354 vdd.n2497 vdd.n1040 185
R17355 vdd.n1419 vdd.n1418 185
R17356 vdd.n1418 vdd.n1047 185
R17357 vdd.n1420 vdd.n1046 185
R17358 vdd.n2490 vdd.n1046 185
R17359 vdd.n1422 vdd.n1421 185
R17360 vdd.n1421 vdd.n1054 185
R17361 vdd.n1423 vdd.n1053 185
R17362 vdd.n2484 vdd.n1053 185
R17363 vdd.n1425 vdd.n1424 185
R17364 vdd.n1424 vdd.n1051 185
R17365 vdd.n1426 vdd.n1060 185
R17366 vdd.n2478 vdd.n1060 185
R17367 vdd.n1428 vdd.n1427 185
R17368 vdd.n1427 vdd.n1058 185
R17369 vdd.n1429 vdd.n1066 185
R17370 vdd.n2472 vdd.n1066 185
R17371 vdd.n1431 vdd.n1430 185
R17372 vdd.n1430 vdd.n1064 185
R17373 vdd.n1432 vdd.n1071 185
R17374 vdd.n2466 vdd.n1071 185
R17375 vdd.n1434 vdd.n1433 185
R17376 vdd.n1433 vdd.n1077 185
R17377 vdd.n1435 vdd.n1076 185
R17378 vdd.n2460 vdd.n1076 185
R17379 vdd.n1437 vdd.n1436 185
R17380 vdd.n1436 vdd.n1083 185
R17381 vdd.n1438 vdd.n1082 185
R17382 vdd.n2454 vdd.n1082 185
R17383 vdd.n1440 vdd.n1439 185
R17384 vdd.n1439 vdd.n1090 185
R17385 vdd.n1441 vdd.n1089 185
R17386 vdd.n2448 vdd.n1089 185
R17387 vdd.n1443 vdd.n1442 185
R17388 vdd.n1442 vdd.n1087 185
R17389 vdd.n1444 vdd.n1096 185
R17390 vdd.n2442 vdd.n1096 185
R17391 vdd.n1446 vdd.n1445 185
R17392 vdd.n1445 vdd.n1094 185
R17393 vdd.n1447 vdd.n1101 185
R17394 vdd.n2436 vdd.n1101 185
R17395 vdd.n1449 vdd.n1448 185
R17396 vdd.n1448 vdd.n1108 185
R17397 vdd.n1450 vdd.n1107 185
R17398 vdd.n2430 vdd.n1107 185
R17399 vdd.n1452 vdd.n1451 185
R17400 vdd.n1451 vdd.n1105 185
R17401 vdd.n1252 vdd.n1251 185
R17402 vdd.n1254 vdd.n1253 185
R17403 vdd.n1256 vdd.n1255 185
R17404 vdd.n1258 vdd.n1257 185
R17405 vdd.n1260 vdd.n1259 185
R17406 vdd.n1262 vdd.n1261 185
R17407 vdd.n1264 vdd.n1263 185
R17408 vdd.n1266 vdd.n1265 185
R17409 vdd.n1268 vdd.n1267 185
R17410 vdd.n1270 vdd.n1269 185
R17411 vdd.n1272 vdd.n1271 185
R17412 vdd.n1274 vdd.n1273 185
R17413 vdd.n1276 vdd.n1275 185
R17414 vdd.n1278 vdd.n1277 185
R17415 vdd.n1280 vdd.n1279 185
R17416 vdd.n1282 vdd.n1281 185
R17417 vdd.n1284 vdd.n1283 185
R17418 vdd.n1486 vdd.n1285 185
R17419 vdd.n1485 vdd.n1484 185
R17420 vdd.n1483 vdd.n1482 185
R17421 vdd.n1481 vdd.n1480 185
R17422 vdd.n1479 vdd.n1478 185
R17423 vdd.n1477 vdd.n1476 185
R17424 vdd.n1475 vdd.n1474 185
R17425 vdd.n1473 vdd.n1472 185
R17426 vdd.n1471 vdd.n1470 185
R17427 vdd.n1469 vdd.n1468 185
R17428 vdd.n1467 vdd.n1466 185
R17429 vdd.n1465 vdd.n1464 185
R17430 vdd.n1463 vdd.n1462 185
R17431 vdd.n1461 vdd.n1460 185
R17432 vdd.n1459 vdd.n1458 185
R17433 vdd.n1457 vdd.n1456 185
R17434 vdd.n1455 vdd.n1454 185
R17435 vdd.n1453 vdd.n1146 185
R17436 vdd.n2423 vdd.n1146 185
R17437 vdd.n315 vdd.n314 171.744
R17438 vdd.n314 vdd.n313 171.744
R17439 vdd.n313 vdd.n282 171.744
R17440 vdd.n306 vdd.n282 171.744
R17441 vdd.n306 vdd.n305 171.744
R17442 vdd.n305 vdd.n287 171.744
R17443 vdd.n298 vdd.n287 171.744
R17444 vdd.n298 vdd.n297 171.744
R17445 vdd.n297 vdd.n291 171.744
R17446 vdd.n260 vdd.n259 171.744
R17447 vdd.n259 vdd.n258 171.744
R17448 vdd.n258 vdd.n227 171.744
R17449 vdd.n251 vdd.n227 171.744
R17450 vdd.n251 vdd.n250 171.744
R17451 vdd.n250 vdd.n232 171.744
R17452 vdd.n243 vdd.n232 171.744
R17453 vdd.n243 vdd.n242 171.744
R17454 vdd.n242 vdd.n236 171.744
R17455 vdd.n217 vdd.n216 171.744
R17456 vdd.n216 vdd.n215 171.744
R17457 vdd.n215 vdd.n184 171.744
R17458 vdd.n208 vdd.n184 171.744
R17459 vdd.n208 vdd.n207 171.744
R17460 vdd.n207 vdd.n189 171.744
R17461 vdd.n200 vdd.n189 171.744
R17462 vdd.n200 vdd.n199 171.744
R17463 vdd.n199 vdd.n193 171.744
R17464 vdd.n162 vdd.n161 171.744
R17465 vdd.n161 vdd.n160 171.744
R17466 vdd.n160 vdd.n129 171.744
R17467 vdd.n153 vdd.n129 171.744
R17468 vdd.n153 vdd.n152 171.744
R17469 vdd.n152 vdd.n134 171.744
R17470 vdd.n145 vdd.n134 171.744
R17471 vdd.n145 vdd.n144 171.744
R17472 vdd.n144 vdd.n138 171.744
R17473 vdd.n120 vdd.n119 171.744
R17474 vdd.n119 vdd.n118 171.744
R17475 vdd.n118 vdd.n87 171.744
R17476 vdd.n111 vdd.n87 171.744
R17477 vdd.n111 vdd.n110 171.744
R17478 vdd.n110 vdd.n92 171.744
R17479 vdd.n103 vdd.n92 171.744
R17480 vdd.n103 vdd.n102 171.744
R17481 vdd.n102 vdd.n96 171.744
R17482 vdd.n65 vdd.n64 171.744
R17483 vdd.n64 vdd.n63 171.744
R17484 vdd.n63 vdd.n32 171.744
R17485 vdd.n56 vdd.n32 171.744
R17486 vdd.n56 vdd.n55 171.744
R17487 vdd.n55 vdd.n37 171.744
R17488 vdd.n48 vdd.n37 171.744
R17489 vdd.n48 vdd.n47 171.744
R17490 vdd.n47 vdd.n41 171.744
R17491 vdd.n2139 vdd.n2138 171.744
R17492 vdd.n2138 vdd.n2137 171.744
R17493 vdd.n2137 vdd.n2106 171.744
R17494 vdd.n2130 vdd.n2106 171.744
R17495 vdd.n2130 vdd.n2129 171.744
R17496 vdd.n2129 vdd.n2111 171.744
R17497 vdd.n2122 vdd.n2111 171.744
R17498 vdd.n2122 vdd.n2121 171.744
R17499 vdd.n2121 vdd.n2115 171.744
R17500 vdd.n2194 vdd.n2193 171.744
R17501 vdd.n2193 vdd.n2192 171.744
R17502 vdd.n2192 vdd.n2161 171.744
R17503 vdd.n2185 vdd.n2161 171.744
R17504 vdd.n2185 vdd.n2184 171.744
R17505 vdd.n2184 vdd.n2166 171.744
R17506 vdd.n2177 vdd.n2166 171.744
R17507 vdd.n2177 vdd.n2176 171.744
R17508 vdd.n2176 vdd.n2170 171.744
R17509 vdd.n2041 vdd.n2040 171.744
R17510 vdd.n2040 vdd.n2039 171.744
R17511 vdd.n2039 vdd.n2008 171.744
R17512 vdd.n2032 vdd.n2008 171.744
R17513 vdd.n2032 vdd.n2031 171.744
R17514 vdd.n2031 vdd.n2013 171.744
R17515 vdd.n2024 vdd.n2013 171.744
R17516 vdd.n2024 vdd.n2023 171.744
R17517 vdd.n2023 vdd.n2017 171.744
R17518 vdd.n2096 vdd.n2095 171.744
R17519 vdd.n2095 vdd.n2094 171.744
R17520 vdd.n2094 vdd.n2063 171.744
R17521 vdd.n2087 vdd.n2063 171.744
R17522 vdd.n2087 vdd.n2086 171.744
R17523 vdd.n2086 vdd.n2068 171.744
R17524 vdd.n2079 vdd.n2068 171.744
R17525 vdd.n2079 vdd.n2078 171.744
R17526 vdd.n2078 vdd.n2072 171.744
R17527 vdd.n1944 vdd.n1943 171.744
R17528 vdd.n1943 vdd.n1942 171.744
R17529 vdd.n1942 vdd.n1911 171.744
R17530 vdd.n1935 vdd.n1911 171.744
R17531 vdd.n1935 vdd.n1934 171.744
R17532 vdd.n1934 vdd.n1916 171.744
R17533 vdd.n1927 vdd.n1916 171.744
R17534 vdd.n1927 vdd.n1926 171.744
R17535 vdd.n1926 vdd.n1920 171.744
R17536 vdd.n1999 vdd.n1998 171.744
R17537 vdd.n1998 vdd.n1997 171.744
R17538 vdd.n1997 vdd.n1966 171.744
R17539 vdd.n1990 vdd.n1966 171.744
R17540 vdd.n1990 vdd.n1989 171.744
R17541 vdd.n1989 vdd.n1971 171.744
R17542 vdd.n1982 vdd.n1971 171.744
R17543 vdd.n1982 vdd.n1981 171.744
R17544 vdd.n1981 vdd.n1975 171.744
R17545 vdd.n449 vdd.n448 146.341
R17546 vdd.n455 vdd.n454 146.341
R17547 vdd.n459 vdd.n458 146.341
R17548 vdd.n465 vdd.n464 146.341
R17549 vdd.n469 vdd.n468 146.341
R17550 vdd.n475 vdd.n474 146.341
R17551 vdd.n479 vdd.n478 146.341
R17552 vdd.n485 vdd.n484 146.341
R17553 vdd.n489 vdd.n488 146.341
R17554 vdd.n495 vdd.n494 146.341
R17555 vdd.n499 vdd.n498 146.341
R17556 vdd.n505 vdd.n504 146.341
R17557 vdd.n509 vdd.n508 146.341
R17558 vdd.n515 vdd.n514 146.341
R17559 vdd.n519 vdd.n518 146.341
R17560 vdd.n525 vdd.n524 146.341
R17561 vdd.n529 vdd.n528 146.341
R17562 vdd.n535 vdd.n534 146.341
R17563 vdd.n539 vdd.n538 146.341
R17564 vdd.n545 vdd.n544 146.341
R17565 vdd.n549 vdd.n548 146.341
R17566 vdd.n555 vdd.n554 146.341
R17567 vdd.n559 vdd.n558 146.341
R17568 vdd.n565 vdd.n564 146.341
R17569 vdd.n569 vdd.n568 146.341
R17570 vdd.n575 vdd.n574 146.341
R17571 vdd.n579 vdd.n578 146.341
R17572 vdd.n585 vdd.n584 146.341
R17573 vdd.n589 vdd.n588 146.341
R17574 vdd.n595 vdd.n594 146.341
R17575 vdd.n597 vdd.n404 146.341
R17576 vdd.n3418 vdd.n654 146.341
R17577 vdd.n3424 vdd.n654 146.341
R17578 vdd.n3424 vdd.n647 146.341
R17579 vdd.n3434 vdd.n647 146.341
R17580 vdd.n3434 vdd.n643 146.341
R17581 vdd.n3440 vdd.n643 146.341
R17582 vdd.n3440 vdd.n634 146.341
R17583 vdd.n3450 vdd.n634 146.341
R17584 vdd.n3450 vdd.n630 146.341
R17585 vdd.n3456 vdd.n630 146.341
R17586 vdd.n3456 vdd.n623 146.341
R17587 vdd.n3467 vdd.n623 146.341
R17588 vdd.n3467 vdd.n619 146.341
R17589 vdd.n3476 vdd.n619 146.341
R17590 vdd.n3476 vdd.n612 146.341
R17591 vdd.n3486 vdd.n612 146.341
R17592 vdd.n3487 vdd.n3486 146.341
R17593 vdd.n3487 vdd.n329 146.341
R17594 vdd.n330 vdd.n329 146.341
R17595 vdd.n331 vdd.n330 146.341
R17596 vdd.n3494 vdd.n331 146.341
R17597 vdd.n3494 vdd.n339 146.341
R17598 vdd.n340 vdd.n339 146.341
R17599 vdd.n341 vdd.n340 146.341
R17600 vdd.n3501 vdd.n341 146.341
R17601 vdd.n3501 vdd.n350 146.341
R17602 vdd.n351 vdd.n350 146.341
R17603 vdd.n352 vdd.n351 146.341
R17604 vdd.n3509 vdd.n352 146.341
R17605 vdd.n3509 vdd.n360 146.341
R17606 vdd.n361 vdd.n360 146.341
R17607 vdd.n362 vdd.n361 146.341
R17608 vdd.n3516 vdd.n362 146.341
R17609 vdd.n3516 vdd.n371 146.341
R17610 vdd.n372 vdd.n371 146.341
R17611 vdd.n3410 vdd.n3408 146.341
R17612 vdd.n3408 vdd.n3407 146.341
R17613 vdd.n3404 vdd.n3403 146.341
R17614 vdd.n3400 vdd.n3399 146.341
R17615 vdd.n3397 vdd.n669 146.341
R17616 vdd.n3393 vdd.n3391 146.341
R17617 vdd.n3389 vdd.n675 146.341
R17618 vdd.n3385 vdd.n3383 146.341
R17619 vdd.n3381 vdd.n681 146.341
R17620 vdd.n3377 vdd.n3375 146.341
R17621 vdd.n3373 vdd.n689 146.341
R17622 vdd.n3369 vdd.n3367 146.341
R17623 vdd.n3365 vdd.n695 146.341
R17624 vdd.n3361 vdd.n3359 146.341
R17625 vdd.n3357 vdd.n701 146.341
R17626 vdd.n3353 vdd.n3351 146.341
R17627 vdd.n3349 vdd.n707 146.341
R17628 vdd.n3345 vdd.n3343 146.341
R17629 vdd.n3341 vdd.n713 146.341
R17630 vdd.n3337 vdd.n3335 146.341
R17631 vdd.n3333 vdd.n719 146.341
R17632 vdd.n3326 vdd.n728 146.341
R17633 vdd.n3324 vdd.n3323 146.341
R17634 vdd.n3320 vdd.n3319 146.341
R17635 vdd.n3317 vdd.n733 146.341
R17636 vdd.n3313 vdd.n3311 146.341
R17637 vdd.n3309 vdd.n739 146.341
R17638 vdd.n3305 vdd.n3303 146.341
R17639 vdd.n3301 vdd.n745 146.341
R17640 vdd.n3297 vdd.n3295 146.341
R17641 vdd.n3292 vdd.n3291 146.341
R17642 vdd.n3288 vdd.n657 146.341
R17643 vdd.n3416 vdd.n653 146.341
R17644 vdd.n3426 vdd.n653 146.341
R17645 vdd.n3426 vdd.n649 146.341
R17646 vdd.n3432 vdd.n649 146.341
R17647 vdd.n3432 vdd.n641 146.341
R17648 vdd.n3442 vdd.n641 146.341
R17649 vdd.n3442 vdd.n637 146.341
R17650 vdd.n3448 vdd.n637 146.341
R17651 vdd.n3448 vdd.n629 146.341
R17652 vdd.n3459 vdd.n629 146.341
R17653 vdd.n3459 vdd.n625 146.341
R17654 vdd.n3465 vdd.n625 146.341
R17655 vdd.n3465 vdd.n618 146.341
R17656 vdd.n3478 vdd.n618 146.341
R17657 vdd.n3478 vdd.n614 146.341
R17658 vdd.n3484 vdd.n614 146.341
R17659 vdd.n3484 vdd.n326 146.341
R17660 vdd.n3560 vdd.n326 146.341
R17661 vdd.n3560 vdd.n327 146.341
R17662 vdd.n3556 vdd.n327 146.341
R17663 vdd.n3556 vdd.n333 146.341
R17664 vdd.n3552 vdd.n333 146.341
R17665 vdd.n3552 vdd.n338 146.341
R17666 vdd.n3548 vdd.n338 146.341
R17667 vdd.n3548 vdd.n342 146.341
R17668 vdd.n3544 vdd.n342 146.341
R17669 vdd.n3544 vdd.n348 146.341
R17670 vdd.n3540 vdd.n348 146.341
R17671 vdd.n3540 vdd.n353 146.341
R17672 vdd.n3536 vdd.n353 146.341
R17673 vdd.n3536 vdd.n359 146.341
R17674 vdd.n3532 vdd.n359 146.341
R17675 vdd.n3532 vdd.n364 146.341
R17676 vdd.n3528 vdd.n364 146.341
R17677 vdd.n3528 vdd.n370 146.341
R17678 vdd.n2388 vdd.n2387 146.341
R17679 vdd.n2385 vdd.n2382 146.341
R17680 vdd.n2380 vdd.n1156 146.341
R17681 vdd.n2376 vdd.n2375 146.341
R17682 vdd.n2373 vdd.n1160 146.341
R17683 vdd.n2369 vdd.n2368 146.341
R17684 vdd.n2366 vdd.n1167 146.341
R17685 vdd.n2362 vdd.n2361 146.341
R17686 vdd.n2359 vdd.n1174 146.341
R17687 vdd.n1185 vdd.n1182 146.341
R17688 vdd.n2351 vdd.n2350 146.341
R17689 vdd.n2348 vdd.n1187 146.341
R17690 vdd.n2344 vdd.n2343 146.341
R17691 vdd.n2341 vdd.n1193 146.341
R17692 vdd.n2337 vdd.n2336 146.341
R17693 vdd.n2334 vdd.n1200 146.341
R17694 vdd.n2330 vdd.n2329 146.341
R17695 vdd.n2327 vdd.n1207 146.341
R17696 vdd.n2323 vdd.n2322 146.341
R17697 vdd.n2320 vdd.n1214 146.341
R17698 vdd.n1225 vdd.n1222 146.341
R17699 vdd.n2312 vdd.n2311 146.341
R17700 vdd.n2309 vdd.n1227 146.341
R17701 vdd.n2305 vdd.n2304 146.341
R17702 vdd.n2302 vdd.n1233 146.341
R17703 vdd.n2298 vdd.n2297 146.341
R17704 vdd.n2295 vdd.n1240 146.341
R17705 vdd.n2291 vdd.n2290 146.341
R17706 vdd.n2288 vdd.n1247 146.341
R17707 vdd.n1493 vdd.n1491 146.341
R17708 vdd.n1496 vdd.n1495 146.341
R17709 vdd.n1836 vdd.n1600 146.341
R17710 vdd.n1836 vdd.n1592 146.341
R17711 vdd.n1846 vdd.n1592 146.341
R17712 vdd.n1846 vdd.n1588 146.341
R17713 vdd.n1852 vdd.n1588 146.341
R17714 vdd.n1852 vdd.n1580 146.341
R17715 vdd.n1863 vdd.n1580 146.341
R17716 vdd.n1863 vdd.n1576 146.341
R17717 vdd.n1869 vdd.n1576 146.341
R17718 vdd.n1869 vdd.n1570 146.341
R17719 vdd.n1880 vdd.n1570 146.341
R17720 vdd.n1880 vdd.n1566 146.341
R17721 vdd.n1886 vdd.n1566 146.341
R17722 vdd.n1886 vdd.n1557 146.341
R17723 vdd.n1896 vdd.n1557 146.341
R17724 vdd.n1896 vdd.n1553 146.341
R17725 vdd.n1902 vdd.n1553 146.341
R17726 vdd.n1902 vdd.n1546 146.341
R17727 vdd.n2208 vdd.n1546 146.341
R17728 vdd.n2208 vdd.n1542 146.341
R17729 vdd.n2214 vdd.n1542 146.341
R17730 vdd.n2214 vdd.n1535 146.341
R17731 vdd.n2224 vdd.n1535 146.341
R17732 vdd.n2224 vdd.n1531 146.341
R17733 vdd.n2230 vdd.n1531 146.341
R17734 vdd.n2230 vdd.n1523 146.341
R17735 vdd.n2241 vdd.n1523 146.341
R17736 vdd.n2241 vdd.n1519 146.341
R17737 vdd.n2247 vdd.n1519 146.341
R17738 vdd.n2247 vdd.n1513 146.341
R17739 vdd.n2258 vdd.n1513 146.341
R17740 vdd.n2258 vdd.n1508 146.341
R17741 vdd.n2266 vdd.n1508 146.341
R17742 vdd.n2266 vdd.n1498 146.341
R17743 vdd.n2276 vdd.n1498 146.341
R17744 vdd.n1638 vdd.n1637 146.341
R17745 vdd.n1642 vdd.n1637 146.341
R17746 vdd.n1644 vdd.n1643 146.341
R17747 vdd.n1648 vdd.n1647 146.341
R17748 vdd.n1650 vdd.n1649 146.341
R17749 vdd.n1654 vdd.n1653 146.341
R17750 vdd.n1656 vdd.n1655 146.341
R17751 vdd.n1660 vdd.n1659 146.341
R17752 vdd.n1662 vdd.n1661 146.341
R17753 vdd.n1794 vdd.n1793 146.341
R17754 vdd.n1666 vdd.n1665 146.341
R17755 vdd.n1670 vdd.n1669 146.341
R17756 vdd.n1672 vdd.n1671 146.341
R17757 vdd.n1676 vdd.n1675 146.341
R17758 vdd.n1678 vdd.n1677 146.341
R17759 vdd.n1682 vdd.n1681 146.341
R17760 vdd.n1684 vdd.n1683 146.341
R17761 vdd.n1688 vdd.n1687 146.341
R17762 vdd.n1690 vdd.n1689 146.341
R17763 vdd.n1694 vdd.n1693 146.341
R17764 vdd.n1758 vdd.n1695 146.341
R17765 vdd.n1699 vdd.n1698 146.341
R17766 vdd.n1701 vdd.n1700 146.341
R17767 vdd.n1705 vdd.n1704 146.341
R17768 vdd.n1707 vdd.n1706 146.341
R17769 vdd.n1711 vdd.n1710 146.341
R17770 vdd.n1713 vdd.n1712 146.341
R17771 vdd.n1717 vdd.n1716 146.341
R17772 vdd.n1719 vdd.n1718 146.341
R17773 vdd.n1723 vdd.n1722 146.341
R17774 vdd.n1725 vdd.n1724 146.341
R17775 vdd.n1830 vdd.n1606 146.341
R17776 vdd.n1838 vdd.n1598 146.341
R17777 vdd.n1838 vdd.n1594 146.341
R17778 vdd.n1844 vdd.n1594 146.341
R17779 vdd.n1844 vdd.n1586 146.341
R17780 vdd.n1855 vdd.n1586 146.341
R17781 vdd.n1855 vdd.n1582 146.341
R17782 vdd.n1861 vdd.n1582 146.341
R17783 vdd.n1861 vdd.n1575 146.341
R17784 vdd.n1872 vdd.n1575 146.341
R17785 vdd.n1872 vdd.n1571 146.341
R17786 vdd.n1878 vdd.n1571 146.341
R17787 vdd.n1878 vdd.n1564 146.341
R17788 vdd.n1888 vdd.n1564 146.341
R17789 vdd.n1888 vdd.n1560 146.341
R17790 vdd.n1894 vdd.n1560 146.341
R17791 vdd.n1894 vdd.n1552 146.341
R17792 vdd.n1905 vdd.n1552 146.341
R17793 vdd.n1905 vdd.n1548 146.341
R17794 vdd.n2206 vdd.n1548 146.341
R17795 vdd.n2206 vdd.n1541 146.341
R17796 vdd.n2216 vdd.n1541 146.341
R17797 vdd.n2216 vdd.n1537 146.341
R17798 vdd.n2222 vdd.n1537 146.341
R17799 vdd.n2222 vdd.n1529 146.341
R17800 vdd.n2233 vdd.n1529 146.341
R17801 vdd.n2233 vdd.n1525 146.341
R17802 vdd.n2239 vdd.n1525 146.341
R17803 vdd.n2239 vdd.n1518 146.341
R17804 vdd.n2250 vdd.n1518 146.341
R17805 vdd.n2250 vdd.n1514 146.341
R17806 vdd.n2256 vdd.n1514 146.341
R17807 vdd.n2256 vdd.n1506 146.341
R17808 vdd.n2268 vdd.n1506 146.341
R17809 vdd.n2268 vdd.n1501 146.341
R17810 vdd.n2274 vdd.n1501 146.341
R17811 vdd.n1286 vdd.t200 127.284
R17812 vdd.n981 vdd.t244 127.284
R17813 vdd.n1290 vdd.t234 127.284
R17814 vdd.n972 vdd.t267 127.284
R17815 vdd.n867 vdd.t221 127.284
R17816 vdd.n867 vdd.t222 127.284
R17817 vdd.n2740 vdd.t262 127.284
R17818 vdd.n804 vdd.t209 127.284
R17819 vdd.n2737 vdd.t252 127.284
R17820 vdd.n768 vdd.t195 127.284
R17821 vdd.n1042 vdd.t258 127.284
R17822 vdd.n1042 vdd.t259 127.284
R17823 vdd.n22 vdd.n20 117.314
R17824 vdd.n17 vdd.n15 117.314
R17825 vdd.n27 vdd.n26 116.927
R17826 vdd.n24 vdd.n23 116.927
R17827 vdd.n22 vdd.n21 116.927
R17828 vdd.n17 vdd.n16 116.927
R17829 vdd.n19 vdd.n18 116.927
R17830 vdd.n27 vdd.n25 116.927
R17831 vdd.n1287 vdd.t199 111.188
R17832 vdd.n982 vdd.t245 111.188
R17833 vdd.n1291 vdd.t233 111.188
R17834 vdd.n973 vdd.t268 111.188
R17835 vdd.n2741 vdd.t261 111.188
R17836 vdd.n805 vdd.t210 111.188
R17837 vdd.n2738 vdd.t251 111.188
R17838 vdd.n769 vdd.t196 111.188
R17839 vdd.n3011 vdd.n931 99.5127
R17840 vdd.n3011 vdd.n922 99.5127
R17841 vdd.n3019 vdd.n922 99.5127
R17842 vdd.n3019 vdd.n920 99.5127
R17843 vdd.n3023 vdd.n920 99.5127
R17844 vdd.n3023 vdd.n910 99.5127
R17845 vdd.n3031 vdd.n910 99.5127
R17846 vdd.n3031 vdd.n908 99.5127
R17847 vdd.n3035 vdd.n908 99.5127
R17848 vdd.n3035 vdd.n899 99.5127
R17849 vdd.n3043 vdd.n899 99.5127
R17850 vdd.n3043 vdd.n897 99.5127
R17851 vdd.n3047 vdd.n897 99.5127
R17852 vdd.n3047 vdd.n888 99.5127
R17853 vdd.n3055 vdd.n888 99.5127
R17854 vdd.n3055 vdd.n886 99.5127
R17855 vdd.n3059 vdd.n886 99.5127
R17856 vdd.n3059 vdd.n875 99.5127
R17857 vdd.n3068 vdd.n875 99.5127
R17858 vdd.n3068 vdd.n873 99.5127
R17859 vdd.n3072 vdd.n873 99.5127
R17860 vdd.n3072 vdd.n863 99.5127
R17861 vdd.n3080 vdd.n863 99.5127
R17862 vdd.n3080 vdd.n861 99.5127
R17863 vdd.n3084 vdd.n861 99.5127
R17864 vdd.n3084 vdd.n851 99.5127
R17865 vdd.n3092 vdd.n851 99.5127
R17866 vdd.n3092 vdd.n849 99.5127
R17867 vdd.n3096 vdd.n849 99.5127
R17868 vdd.n3096 vdd.n838 99.5127
R17869 vdd.n3104 vdd.n838 99.5127
R17870 vdd.n3104 vdd.n836 99.5127
R17871 vdd.n3108 vdd.n836 99.5127
R17872 vdd.n3108 vdd.n827 99.5127
R17873 vdd.n3116 vdd.n827 99.5127
R17874 vdd.n3116 vdd.n825 99.5127
R17875 vdd.n3120 vdd.n825 99.5127
R17876 vdd.n3120 vdd.n813 99.5127
R17877 vdd.n3173 vdd.n813 99.5127
R17878 vdd.n3173 vdd.n811 99.5127
R17879 vdd.n3177 vdd.n811 99.5127
R17880 vdd.n3177 vdd.n777 99.5127
R17881 vdd.n3247 vdd.n777 99.5127
R17882 vdd.n3243 vdd.n778 99.5127
R17883 vdd.n3241 vdd.n3240 99.5127
R17884 vdd.n3238 vdd.n782 99.5127
R17885 vdd.n3234 vdd.n3233 99.5127
R17886 vdd.n3231 vdd.n785 99.5127
R17887 vdd.n3227 vdd.n3226 99.5127
R17888 vdd.n3224 vdd.n788 99.5127
R17889 vdd.n3220 vdd.n3219 99.5127
R17890 vdd.n3217 vdd.n791 99.5127
R17891 vdd.n3212 vdd.n3211 99.5127
R17892 vdd.n3209 vdd.n794 99.5127
R17893 vdd.n3205 vdd.n3204 99.5127
R17894 vdd.n3202 vdd.n797 99.5127
R17895 vdd.n3198 vdd.n3197 99.5127
R17896 vdd.n3195 vdd.n800 99.5127
R17897 vdd.n3191 vdd.n3190 99.5127
R17898 vdd.n3188 vdd.n803 99.5127
R17899 vdd.n2938 vdd.n929 99.5127
R17900 vdd.n2934 vdd.n929 99.5127
R17901 vdd.n2934 vdd.n923 99.5127
R17902 vdd.n2816 vdd.n923 99.5127
R17903 vdd.n2816 vdd.n918 99.5127
R17904 vdd.n2819 vdd.n918 99.5127
R17905 vdd.n2819 vdd.n912 99.5127
R17906 vdd.n2920 vdd.n912 99.5127
R17907 vdd.n2920 vdd.n906 99.5127
R17908 vdd.n2916 vdd.n906 99.5127
R17909 vdd.n2916 vdd.n900 99.5127
R17910 vdd.n2863 vdd.n900 99.5127
R17911 vdd.n2863 vdd.n894 99.5127
R17912 vdd.n2860 vdd.n894 99.5127
R17913 vdd.n2860 vdd.n889 99.5127
R17914 vdd.n2857 vdd.n889 99.5127
R17915 vdd.n2857 vdd.n884 99.5127
R17916 vdd.n2854 vdd.n884 99.5127
R17917 vdd.n2854 vdd.n877 99.5127
R17918 vdd.n2851 vdd.n877 99.5127
R17919 vdd.n2851 vdd.n870 99.5127
R17920 vdd.n2848 vdd.n870 99.5127
R17921 vdd.n2848 vdd.n864 99.5127
R17922 vdd.n2845 vdd.n864 99.5127
R17923 vdd.n2845 vdd.n859 99.5127
R17924 vdd.n2842 vdd.n859 99.5127
R17925 vdd.n2842 vdd.n853 99.5127
R17926 vdd.n2839 vdd.n853 99.5127
R17927 vdd.n2839 vdd.n846 99.5127
R17928 vdd.n2836 vdd.n846 99.5127
R17929 vdd.n2836 vdd.n839 99.5127
R17930 vdd.n2833 vdd.n839 99.5127
R17931 vdd.n2833 vdd.n833 99.5127
R17932 vdd.n2830 vdd.n833 99.5127
R17933 vdd.n2830 vdd.n828 99.5127
R17934 vdd.n2827 vdd.n828 99.5127
R17935 vdd.n2827 vdd.n823 99.5127
R17936 vdd.n2824 vdd.n823 99.5127
R17937 vdd.n2824 vdd.n815 99.5127
R17938 vdd.n815 vdd.n808 99.5127
R17939 vdd.n3179 vdd.n808 99.5127
R17940 vdd.n3180 vdd.n3179 99.5127
R17941 vdd.n3180 vdd.n775 99.5127
R17942 vdd.n3004 vdd.n933 99.5127
R17943 vdd.n3004 vdd.n2736 99.5127
R17944 vdd.n3000 vdd.n2999 99.5127
R17945 vdd.n2996 vdd.n2995 99.5127
R17946 vdd.n2992 vdd.n2991 99.5127
R17947 vdd.n2988 vdd.n2987 99.5127
R17948 vdd.n2984 vdd.n2983 99.5127
R17949 vdd.n2980 vdd.n2979 99.5127
R17950 vdd.n2976 vdd.n2975 99.5127
R17951 vdd.n2972 vdd.n2971 99.5127
R17952 vdd.n2968 vdd.n2967 99.5127
R17953 vdd.n2964 vdd.n2963 99.5127
R17954 vdd.n2960 vdd.n2959 99.5127
R17955 vdd.n2956 vdd.n2955 99.5127
R17956 vdd.n2952 vdd.n2951 99.5127
R17957 vdd.n2948 vdd.n2947 99.5127
R17958 vdd.n2943 vdd.n2942 99.5127
R17959 vdd.n2700 vdd.n970 99.5127
R17960 vdd.n2696 vdd.n2695 99.5127
R17961 vdd.n2692 vdd.n2691 99.5127
R17962 vdd.n2688 vdd.n2687 99.5127
R17963 vdd.n2684 vdd.n2683 99.5127
R17964 vdd.n2680 vdd.n2679 99.5127
R17965 vdd.n2676 vdd.n2675 99.5127
R17966 vdd.n2672 vdd.n2671 99.5127
R17967 vdd.n2668 vdd.n2667 99.5127
R17968 vdd.n2664 vdd.n2663 99.5127
R17969 vdd.n2660 vdd.n2659 99.5127
R17970 vdd.n2656 vdd.n2655 99.5127
R17971 vdd.n2652 vdd.n2651 99.5127
R17972 vdd.n2648 vdd.n2647 99.5127
R17973 vdd.n2644 vdd.n2643 99.5127
R17974 vdd.n2640 vdd.n2639 99.5127
R17975 vdd.n2635 vdd.n2634 99.5127
R17976 vdd.n1326 vdd.n1106 99.5127
R17977 vdd.n1329 vdd.n1106 99.5127
R17978 vdd.n1329 vdd.n1100 99.5127
R17979 vdd.n1332 vdd.n1100 99.5127
R17980 vdd.n1332 vdd.n1095 99.5127
R17981 vdd.n1335 vdd.n1095 99.5127
R17982 vdd.n1335 vdd.n1088 99.5127
R17983 vdd.n1338 vdd.n1088 99.5127
R17984 vdd.n1338 vdd.n1081 99.5127
R17985 vdd.n1341 vdd.n1081 99.5127
R17986 vdd.n1341 vdd.n1075 99.5127
R17987 vdd.n1344 vdd.n1075 99.5127
R17988 vdd.n1344 vdd.n1070 99.5127
R17989 vdd.n1347 vdd.n1070 99.5127
R17990 vdd.n1347 vdd.n1065 99.5127
R17991 vdd.n1350 vdd.n1065 99.5127
R17992 vdd.n1350 vdd.n1059 99.5127
R17993 vdd.n1353 vdd.n1059 99.5127
R17994 vdd.n1353 vdd.n1052 99.5127
R17995 vdd.n1356 vdd.n1052 99.5127
R17996 vdd.n1356 vdd.n1045 99.5127
R17997 vdd.n1359 vdd.n1045 99.5127
R17998 vdd.n1359 vdd.n1039 99.5127
R17999 vdd.n1362 vdd.n1039 99.5127
R18000 vdd.n1362 vdd.n1034 99.5127
R18001 vdd.n1365 vdd.n1034 99.5127
R18002 vdd.n1365 vdd.n1028 99.5127
R18003 vdd.n1407 vdd.n1028 99.5127
R18004 vdd.n1407 vdd.n1021 99.5127
R18005 vdd.n1403 vdd.n1021 99.5127
R18006 vdd.n1403 vdd.n1015 99.5127
R18007 vdd.n1400 vdd.n1015 99.5127
R18008 vdd.n1400 vdd.n1010 99.5127
R18009 vdd.n1397 vdd.n1010 99.5127
R18010 vdd.n1397 vdd.n1005 99.5127
R18011 vdd.n1377 vdd.n1005 99.5127
R18012 vdd.n1377 vdd.n1000 99.5127
R18013 vdd.n1374 vdd.n1000 99.5127
R18014 vdd.n1374 vdd.n993 99.5127
R18015 vdd.n1371 vdd.n993 99.5127
R18016 vdd.n1371 vdd.n986 99.5127
R18017 vdd.n986 vdd.n975 99.5127
R18018 vdd.n2630 vdd.n975 99.5127
R18019 vdd.n2422 vdd.n1111 99.5127
R18020 vdd.n2422 vdd.n1147 99.5127
R18021 vdd.n2418 vdd.n2417 99.5127
R18022 vdd.n2414 vdd.n2413 99.5127
R18023 vdd.n2410 vdd.n2409 99.5127
R18024 vdd.n2406 vdd.n2405 99.5127
R18025 vdd.n2402 vdd.n2401 99.5127
R18026 vdd.n2398 vdd.n2397 99.5127
R18027 vdd.n2394 vdd.n2393 99.5127
R18028 vdd.n1293 vdd.n1292 99.5127
R18029 vdd.n1297 vdd.n1296 99.5127
R18030 vdd.n1301 vdd.n1300 99.5127
R18031 vdd.n1305 vdd.n1304 99.5127
R18032 vdd.n1309 vdd.n1308 99.5127
R18033 vdd.n1313 vdd.n1312 99.5127
R18034 vdd.n1317 vdd.n1316 99.5127
R18035 vdd.n1322 vdd.n1321 99.5127
R18036 vdd.n2429 vdd.n1109 99.5127
R18037 vdd.n2429 vdd.n1099 99.5127
R18038 vdd.n2437 vdd.n1099 99.5127
R18039 vdd.n2437 vdd.n1097 99.5127
R18040 vdd.n2441 vdd.n1097 99.5127
R18041 vdd.n2441 vdd.n1086 99.5127
R18042 vdd.n2449 vdd.n1086 99.5127
R18043 vdd.n2449 vdd.n1084 99.5127
R18044 vdd.n2453 vdd.n1084 99.5127
R18045 vdd.n2453 vdd.n1074 99.5127
R18046 vdd.n2461 vdd.n1074 99.5127
R18047 vdd.n2461 vdd.n1072 99.5127
R18048 vdd.n2465 vdd.n1072 99.5127
R18049 vdd.n2465 vdd.n1063 99.5127
R18050 vdd.n2473 vdd.n1063 99.5127
R18051 vdd.n2473 vdd.n1061 99.5127
R18052 vdd.n2477 vdd.n1061 99.5127
R18053 vdd.n2477 vdd.n1050 99.5127
R18054 vdd.n2485 vdd.n1050 99.5127
R18055 vdd.n2485 vdd.n1048 99.5127
R18056 vdd.n2489 vdd.n1048 99.5127
R18057 vdd.n2489 vdd.n1038 99.5127
R18058 vdd.n2498 vdd.n1038 99.5127
R18059 vdd.n2498 vdd.n1036 99.5127
R18060 vdd.n2502 vdd.n1036 99.5127
R18061 vdd.n2502 vdd.n1026 99.5127
R18062 vdd.n2510 vdd.n1026 99.5127
R18063 vdd.n2510 vdd.n1024 99.5127
R18064 vdd.n2514 vdd.n1024 99.5127
R18065 vdd.n2514 vdd.n1014 99.5127
R18066 vdd.n2522 vdd.n1014 99.5127
R18067 vdd.n2522 vdd.n1012 99.5127
R18068 vdd.n2526 vdd.n1012 99.5127
R18069 vdd.n2526 vdd.n1004 99.5127
R18070 vdd.n2534 vdd.n1004 99.5127
R18071 vdd.n2534 vdd.n1002 99.5127
R18072 vdd.n2538 vdd.n1002 99.5127
R18073 vdd.n2538 vdd.n991 99.5127
R18074 vdd.n2548 vdd.n991 99.5127
R18075 vdd.n2548 vdd.n988 99.5127
R18076 vdd.n2553 vdd.n988 99.5127
R18077 vdd.n2553 vdd.n989 99.5127
R18078 vdd.n989 vdd.n969 99.5127
R18079 vdd.n3163 vdd.n3162 99.5127
R18080 vdd.n3160 vdd.n3126 99.5127
R18081 vdd.n3156 vdd.n3155 99.5127
R18082 vdd.n3153 vdd.n3129 99.5127
R18083 vdd.n3149 vdd.n3148 99.5127
R18084 vdd.n3146 vdd.n3132 99.5127
R18085 vdd.n3142 vdd.n3141 99.5127
R18086 vdd.n3139 vdd.n3136 99.5127
R18087 vdd.n3280 vdd.n755 99.5127
R18088 vdd.n3278 vdd.n3277 99.5127
R18089 vdd.n3275 vdd.n758 99.5127
R18090 vdd.n3271 vdd.n3270 99.5127
R18091 vdd.n3268 vdd.n761 99.5127
R18092 vdd.n3264 vdd.n3263 99.5127
R18093 vdd.n3261 vdd.n764 99.5127
R18094 vdd.n3257 vdd.n3256 99.5127
R18095 vdd.n3254 vdd.n767 99.5127
R18096 vdd.n2812 vdd.n930 99.5127
R18097 vdd.n2932 vdd.n930 99.5127
R18098 vdd.n2932 vdd.n924 99.5127
R18099 vdd.n2928 vdd.n924 99.5127
R18100 vdd.n2928 vdd.n919 99.5127
R18101 vdd.n2925 vdd.n919 99.5127
R18102 vdd.n2925 vdd.n913 99.5127
R18103 vdd.n2922 vdd.n913 99.5127
R18104 vdd.n2922 vdd.n907 99.5127
R18105 vdd.n2914 vdd.n907 99.5127
R18106 vdd.n2914 vdd.n901 99.5127
R18107 vdd.n2910 vdd.n901 99.5127
R18108 vdd.n2910 vdd.n895 99.5127
R18109 vdd.n2907 vdd.n895 99.5127
R18110 vdd.n2907 vdd.n890 99.5127
R18111 vdd.n2904 vdd.n890 99.5127
R18112 vdd.n2904 vdd.n885 99.5127
R18113 vdd.n2901 vdd.n885 99.5127
R18114 vdd.n2901 vdd.n878 99.5127
R18115 vdd.n2898 vdd.n878 99.5127
R18116 vdd.n2898 vdd.n871 99.5127
R18117 vdd.n2895 vdd.n871 99.5127
R18118 vdd.n2895 vdd.n865 99.5127
R18119 vdd.n2892 vdd.n865 99.5127
R18120 vdd.n2892 vdd.n860 99.5127
R18121 vdd.n2889 vdd.n860 99.5127
R18122 vdd.n2889 vdd.n854 99.5127
R18123 vdd.n2886 vdd.n854 99.5127
R18124 vdd.n2886 vdd.n847 99.5127
R18125 vdd.n2883 vdd.n847 99.5127
R18126 vdd.n2883 vdd.n840 99.5127
R18127 vdd.n2880 vdd.n840 99.5127
R18128 vdd.n2880 vdd.n834 99.5127
R18129 vdd.n2877 vdd.n834 99.5127
R18130 vdd.n2877 vdd.n829 99.5127
R18131 vdd.n2874 vdd.n829 99.5127
R18132 vdd.n2874 vdd.n824 99.5127
R18133 vdd.n2871 vdd.n824 99.5127
R18134 vdd.n2871 vdd.n816 99.5127
R18135 vdd.n2868 vdd.n816 99.5127
R18136 vdd.n2868 vdd.n809 99.5127
R18137 vdd.n809 vdd.n773 99.5127
R18138 vdd.n3249 vdd.n773 99.5127
R18139 vdd.n2747 vdd.n2746 99.5127
R18140 vdd.n2751 vdd.n2750 99.5127
R18141 vdd.n2755 vdd.n2754 99.5127
R18142 vdd.n2759 vdd.n2758 99.5127
R18143 vdd.n2763 vdd.n2762 99.5127
R18144 vdd.n2767 vdd.n2766 99.5127
R18145 vdd.n2771 vdd.n2770 99.5127
R18146 vdd.n2775 vdd.n2774 99.5127
R18147 vdd.n2779 vdd.n2778 99.5127
R18148 vdd.n2783 vdd.n2782 99.5127
R18149 vdd.n2787 vdd.n2786 99.5127
R18150 vdd.n2791 vdd.n2790 99.5127
R18151 vdd.n2795 vdd.n2794 99.5127
R18152 vdd.n2799 vdd.n2798 99.5127
R18153 vdd.n2803 vdd.n2802 99.5127
R18154 vdd.n2807 vdd.n2806 99.5127
R18155 vdd.n2809 vdd.n2735 99.5127
R18156 vdd.n3013 vdd.n927 99.5127
R18157 vdd.n3013 vdd.n925 99.5127
R18158 vdd.n3017 vdd.n925 99.5127
R18159 vdd.n3017 vdd.n916 99.5127
R18160 vdd.n3025 vdd.n916 99.5127
R18161 vdd.n3025 vdd.n914 99.5127
R18162 vdd.n3029 vdd.n914 99.5127
R18163 vdd.n3029 vdd.n905 99.5127
R18164 vdd.n3037 vdd.n905 99.5127
R18165 vdd.n3037 vdd.n903 99.5127
R18166 vdd.n3041 vdd.n903 99.5127
R18167 vdd.n3041 vdd.n893 99.5127
R18168 vdd.n3049 vdd.n893 99.5127
R18169 vdd.n3049 vdd.n891 99.5127
R18170 vdd.n3053 vdd.n891 99.5127
R18171 vdd.n3053 vdd.n882 99.5127
R18172 vdd.n3061 vdd.n882 99.5127
R18173 vdd.n3061 vdd.n880 99.5127
R18174 vdd.n3066 vdd.n880 99.5127
R18175 vdd.n3066 vdd.n869 99.5127
R18176 vdd.n3074 vdd.n869 99.5127
R18177 vdd.n3074 vdd.n866 99.5127
R18178 vdd.n3078 vdd.n866 99.5127
R18179 vdd.n3078 vdd.n857 99.5127
R18180 vdd.n3086 vdd.n857 99.5127
R18181 vdd.n3086 vdd.n855 99.5127
R18182 vdd.n3090 vdd.n855 99.5127
R18183 vdd.n3090 vdd.n844 99.5127
R18184 vdd.n3098 vdd.n844 99.5127
R18185 vdd.n3098 vdd.n842 99.5127
R18186 vdd.n3102 vdd.n842 99.5127
R18187 vdd.n3102 vdd.n832 99.5127
R18188 vdd.n3110 vdd.n832 99.5127
R18189 vdd.n3110 vdd.n830 99.5127
R18190 vdd.n3114 vdd.n830 99.5127
R18191 vdd.n3114 vdd.n821 99.5127
R18192 vdd.n3122 vdd.n821 99.5127
R18193 vdd.n3122 vdd.n818 99.5127
R18194 vdd.n3171 vdd.n818 99.5127
R18195 vdd.n3171 vdd.n819 99.5127
R18196 vdd.n819 vdd.n810 99.5127
R18197 vdd.n3166 vdd.n810 99.5127
R18198 vdd.n3166 vdd.n776 99.5127
R18199 vdd.n2624 vdd.n2623 99.5127
R18200 vdd.n2620 vdd.n2619 99.5127
R18201 vdd.n2616 vdd.n2615 99.5127
R18202 vdd.n2612 vdd.n2611 99.5127
R18203 vdd.n2608 vdd.n2607 99.5127
R18204 vdd.n2604 vdd.n2603 99.5127
R18205 vdd.n2600 vdd.n2599 99.5127
R18206 vdd.n2596 vdd.n2595 99.5127
R18207 vdd.n2592 vdd.n2591 99.5127
R18208 vdd.n2588 vdd.n2587 99.5127
R18209 vdd.n2584 vdd.n2583 99.5127
R18210 vdd.n2580 vdd.n2579 99.5127
R18211 vdd.n2576 vdd.n2575 99.5127
R18212 vdd.n2572 vdd.n2571 99.5127
R18213 vdd.n2568 vdd.n2567 99.5127
R18214 vdd.n2564 vdd.n2563 99.5127
R18215 vdd.n2560 vdd.n951 99.5127
R18216 vdd.n1451 vdd.n1107 99.5127
R18217 vdd.n1448 vdd.n1107 99.5127
R18218 vdd.n1448 vdd.n1101 99.5127
R18219 vdd.n1445 vdd.n1101 99.5127
R18220 vdd.n1445 vdd.n1096 99.5127
R18221 vdd.n1442 vdd.n1096 99.5127
R18222 vdd.n1442 vdd.n1089 99.5127
R18223 vdd.n1439 vdd.n1089 99.5127
R18224 vdd.n1439 vdd.n1082 99.5127
R18225 vdd.n1436 vdd.n1082 99.5127
R18226 vdd.n1436 vdd.n1076 99.5127
R18227 vdd.n1433 vdd.n1076 99.5127
R18228 vdd.n1433 vdd.n1071 99.5127
R18229 vdd.n1430 vdd.n1071 99.5127
R18230 vdd.n1430 vdd.n1066 99.5127
R18231 vdd.n1427 vdd.n1066 99.5127
R18232 vdd.n1427 vdd.n1060 99.5127
R18233 vdd.n1424 vdd.n1060 99.5127
R18234 vdd.n1424 vdd.n1053 99.5127
R18235 vdd.n1421 vdd.n1053 99.5127
R18236 vdd.n1421 vdd.n1046 99.5127
R18237 vdd.n1418 vdd.n1046 99.5127
R18238 vdd.n1418 vdd.n1040 99.5127
R18239 vdd.n1415 vdd.n1040 99.5127
R18240 vdd.n1415 vdd.n1035 99.5127
R18241 vdd.n1412 vdd.n1035 99.5127
R18242 vdd.n1412 vdd.n1029 99.5127
R18243 vdd.n1409 vdd.n1029 99.5127
R18244 vdd.n1409 vdd.n1022 99.5127
R18245 vdd.n1380 vdd.n1022 99.5127
R18246 vdd.n1380 vdd.n1016 99.5127
R18247 vdd.n1383 vdd.n1016 99.5127
R18248 vdd.n1383 vdd.n1011 99.5127
R18249 vdd.n1395 vdd.n1011 99.5127
R18250 vdd.n1395 vdd.n1006 99.5127
R18251 vdd.n1391 vdd.n1006 99.5127
R18252 vdd.n1391 vdd.n1001 99.5127
R18253 vdd.n1388 vdd.n1001 99.5127
R18254 vdd.n1388 vdd.n994 99.5127
R18255 vdd.n994 vdd.n985 99.5127
R18256 vdd.n2555 vdd.n985 99.5127
R18257 vdd.n2556 vdd.n2555 99.5127
R18258 vdd.n2556 vdd.n977 99.5127
R18259 vdd.n1255 vdd.n1254 99.5127
R18260 vdd.n1259 vdd.n1258 99.5127
R18261 vdd.n1263 vdd.n1262 99.5127
R18262 vdd.n1267 vdd.n1266 99.5127
R18263 vdd.n1271 vdd.n1270 99.5127
R18264 vdd.n1275 vdd.n1274 99.5127
R18265 vdd.n1279 vdd.n1278 99.5127
R18266 vdd.n1283 vdd.n1282 99.5127
R18267 vdd.n1484 vdd.n1285 99.5127
R18268 vdd.n1482 vdd.n1481 99.5127
R18269 vdd.n1478 vdd.n1477 99.5127
R18270 vdd.n1474 vdd.n1473 99.5127
R18271 vdd.n1470 vdd.n1469 99.5127
R18272 vdd.n1466 vdd.n1465 99.5127
R18273 vdd.n1462 vdd.n1461 99.5127
R18274 vdd.n1458 vdd.n1457 99.5127
R18275 vdd.n1454 vdd.n1146 99.5127
R18276 vdd.n2431 vdd.n1104 99.5127
R18277 vdd.n2431 vdd.n1102 99.5127
R18278 vdd.n2435 vdd.n1102 99.5127
R18279 vdd.n2435 vdd.n1093 99.5127
R18280 vdd.n2443 vdd.n1093 99.5127
R18281 vdd.n2443 vdd.n1091 99.5127
R18282 vdd.n2447 vdd.n1091 99.5127
R18283 vdd.n2447 vdd.n1080 99.5127
R18284 vdd.n2455 vdd.n1080 99.5127
R18285 vdd.n2455 vdd.n1078 99.5127
R18286 vdd.n2459 vdd.n1078 99.5127
R18287 vdd.n2459 vdd.n1069 99.5127
R18288 vdd.n2467 vdd.n1069 99.5127
R18289 vdd.n2467 vdd.n1067 99.5127
R18290 vdd.n2471 vdd.n1067 99.5127
R18291 vdd.n2471 vdd.n1057 99.5127
R18292 vdd.n2479 vdd.n1057 99.5127
R18293 vdd.n2479 vdd.n1055 99.5127
R18294 vdd.n2483 vdd.n1055 99.5127
R18295 vdd.n2483 vdd.n1044 99.5127
R18296 vdd.n2491 vdd.n1044 99.5127
R18297 vdd.n2491 vdd.n1041 99.5127
R18298 vdd.n2496 vdd.n1041 99.5127
R18299 vdd.n2496 vdd.n1032 99.5127
R18300 vdd.n2504 vdd.n1032 99.5127
R18301 vdd.n2504 vdd.n1030 99.5127
R18302 vdd.n2508 vdd.n1030 99.5127
R18303 vdd.n2508 vdd.n1020 99.5127
R18304 vdd.n2516 vdd.n1020 99.5127
R18305 vdd.n2516 vdd.n1018 99.5127
R18306 vdd.n2520 vdd.n1018 99.5127
R18307 vdd.n2520 vdd.n1009 99.5127
R18308 vdd.n2528 vdd.n1009 99.5127
R18309 vdd.n2528 vdd.n1007 99.5127
R18310 vdd.n2532 vdd.n1007 99.5127
R18311 vdd.n2532 vdd.n998 99.5127
R18312 vdd.n2540 vdd.n998 99.5127
R18313 vdd.n2540 vdd.n995 99.5127
R18314 vdd.n2546 vdd.n995 99.5127
R18315 vdd.n2546 vdd.n996 99.5127
R18316 vdd.n996 vdd.n987 99.5127
R18317 vdd.n987 vdd.n978 99.5127
R18318 vdd.n2628 vdd.n978 99.5127
R18319 vdd.n9 vdd.n7 98.9633
R18320 vdd.n2 vdd.n0 98.9633
R18321 vdd.n9 vdd.n8 98.6055
R18322 vdd.n11 vdd.n10 98.6055
R18323 vdd.n13 vdd.n12 98.6055
R18324 vdd.n6 vdd.n5 98.6055
R18325 vdd.n4 vdd.n3 98.6055
R18326 vdd.n2 vdd.n1 98.6055
R18327 vdd.t99 vdd.n291 85.8723
R18328 vdd.t185 vdd.n236 85.8723
R18329 vdd.t81 vdd.n193 85.8723
R18330 vdd.t175 vdd.n138 85.8723
R18331 vdd.t145 vdd.n96 85.8723
R18332 vdd.t130 vdd.n41 85.8723
R18333 vdd.t69 vdd.n2115 85.8723
R18334 vdd.t148 vdd.n2170 85.8723
R18335 vdd.t100 vdd.n2017 85.8723
R18336 vdd.t139 vdd.n2072 85.8723
R18337 vdd.t131 vdd.n1920 85.8723
R18338 vdd.t147 vdd.n1975 85.8723
R18339 vdd.n868 vdd.n867 78.546
R18340 vdd.n2494 vdd.n1042 78.546
R18341 vdd.n278 vdd.n277 75.1835
R18342 vdd.n276 vdd.n275 75.1835
R18343 vdd.n274 vdd.n273 75.1835
R18344 vdd.n272 vdd.n271 75.1835
R18345 vdd.n270 vdd.n269 75.1835
R18346 vdd.n268 vdd.n267 75.1835
R18347 vdd.n266 vdd.n265 75.1835
R18348 vdd.n180 vdd.n179 75.1835
R18349 vdd.n178 vdd.n177 75.1835
R18350 vdd.n176 vdd.n175 75.1835
R18351 vdd.n174 vdd.n173 75.1835
R18352 vdd.n172 vdd.n171 75.1835
R18353 vdd.n170 vdd.n169 75.1835
R18354 vdd.n168 vdd.n167 75.1835
R18355 vdd.n83 vdd.n82 75.1835
R18356 vdd.n81 vdd.n80 75.1835
R18357 vdd.n79 vdd.n78 75.1835
R18358 vdd.n77 vdd.n76 75.1835
R18359 vdd.n75 vdd.n74 75.1835
R18360 vdd.n73 vdd.n72 75.1835
R18361 vdd.n71 vdd.n70 75.1835
R18362 vdd.n2145 vdd.n2144 75.1835
R18363 vdd.n2147 vdd.n2146 75.1835
R18364 vdd.n2149 vdd.n2148 75.1835
R18365 vdd.n2151 vdd.n2150 75.1835
R18366 vdd.n2153 vdd.n2152 75.1835
R18367 vdd.n2155 vdd.n2154 75.1835
R18368 vdd.n2157 vdd.n2156 75.1835
R18369 vdd.n2047 vdd.n2046 75.1835
R18370 vdd.n2049 vdd.n2048 75.1835
R18371 vdd.n2051 vdd.n2050 75.1835
R18372 vdd.n2053 vdd.n2052 75.1835
R18373 vdd.n2055 vdd.n2054 75.1835
R18374 vdd.n2057 vdd.n2056 75.1835
R18375 vdd.n2059 vdd.n2058 75.1835
R18376 vdd.n1950 vdd.n1949 75.1835
R18377 vdd.n1952 vdd.n1951 75.1835
R18378 vdd.n1954 vdd.n1953 75.1835
R18379 vdd.n1956 vdd.n1955 75.1835
R18380 vdd.n1958 vdd.n1957 75.1835
R18381 vdd.n1960 vdd.n1959 75.1835
R18382 vdd.n1962 vdd.n1961 75.1835
R18383 vdd.n3005 vdd.n2718 72.8958
R18384 vdd.n3005 vdd.n2719 72.8958
R18385 vdd.n3005 vdd.n2720 72.8958
R18386 vdd.n3005 vdd.n2721 72.8958
R18387 vdd.n3005 vdd.n2722 72.8958
R18388 vdd.n3005 vdd.n2723 72.8958
R18389 vdd.n3005 vdd.n2724 72.8958
R18390 vdd.n3005 vdd.n2725 72.8958
R18391 vdd.n3005 vdd.n2726 72.8958
R18392 vdd.n3005 vdd.n2727 72.8958
R18393 vdd.n3005 vdd.n2728 72.8958
R18394 vdd.n3005 vdd.n2729 72.8958
R18395 vdd.n3005 vdd.n2730 72.8958
R18396 vdd.n3005 vdd.n2731 72.8958
R18397 vdd.n3005 vdd.n2732 72.8958
R18398 vdd.n3005 vdd.n2733 72.8958
R18399 vdd.n3005 vdd.n2734 72.8958
R18400 vdd.n772 vdd.n756 72.8958
R18401 vdd.n3255 vdd.n756 72.8958
R18402 vdd.n766 vdd.n756 72.8958
R18403 vdd.n3262 vdd.n756 72.8958
R18404 vdd.n763 vdd.n756 72.8958
R18405 vdd.n3269 vdd.n756 72.8958
R18406 vdd.n760 vdd.n756 72.8958
R18407 vdd.n3276 vdd.n756 72.8958
R18408 vdd.n3279 vdd.n756 72.8958
R18409 vdd.n3135 vdd.n756 72.8958
R18410 vdd.n3140 vdd.n756 72.8958
R18411 vdd.n3134 vdd.n756 72.8958
R18412 vdd.n3147 vdd.n756 72.8958
R18413 vdd.n3131 vdd.n756 72.8958
R18414 vdd.n3154 vdd.n756 72.8958
R18415 vdd.n3128 vdd.n756 72.8958
R18416 vdd.n3161 vdd.n756 72.8958
R18417 vdd.n2424 vdd.n2423 72.8958
R18418 vdd.n2423 vdd.n1113 72.8958
R18419 vdd.n2423 vdd.n1114 72.8958
R18420 vdd.n2423 vdd.n1115 72.8958
R18421 vdd.n2423 vdd.n1116 72.8958
R18422 vdd.n2423 vdd.n1117 72.8958
R18423 vdd.n2423 vdd.n1118 72.8958
R18424 vdd.n2423 vdd.n1119 72.8958
R18425 vdd.n2423 vdd.n1120 72.8958
R18426 vdd.n2423 vdd.n1121 72.8958
R18427 vdd.n2423 vdd.n1122 72.8958
R18428 vdd.n2423 vdd.n1123 72.8958
R18429 vdd.n2423 vdd.n1124 72.8958
R18430 vdd.n2423 vdd.n1125 72.8958
R18431 vdd.n2423 vdd.n1126 72.8958
R18432 vdd.n2423 vdd.n1127 72.8958
R18433 vdd.n2423 vdd.n1128 72.8958
R18434 vdd.n2701 vdd.n952 72.8958
R18435 vdd.n2701 vdd.n953 72.8958
R18436 vdd.n2701 vdd.n954 72.8958
R18437 vdd.n2701 vdd.n955 72.8958
R18438 vdd.n2701 vdd.n956 72.8958
R18439 vdd.n2701 vdd.n957 72.8958
R18440 vdd.n2701 vdd.n958 72.8958
R18441 vdd.n2701 vdd.n959 72.8958
R18442 vdd.n2701 vdd.n960 72.8958
R18443 vdd.n2701 vdd.n961 72.8958
R18444 vdd.n2701 vdd.n962 72.8958
R18445 vdd.n2701 vdd.n963 72.8958
R18446 vdd.n2701 vdd.n964 72.8958
R18447 vdd.n2701 vdd.n965 72.8958
R18448 vdd.n2701 vdd.n966 72.8958
R18449 vdd.n2701 vdd.n967 72.8958
R18450 vdd.n2701 vdd.n968 72.8958
R18451 vdd.n3006 vdd.n3005 72.8958
R18452 vdd.n3005 vdd.n2702 72.8958
R18453 vdd.n3005 vdd.n2703 72.8958
R18454 vdd.n3005 vdd.n2704 72.8958
R18455 vdd.n3005 vdd.n2705 72.8958
R18456 vdd.n3005 vdd.n2706 72.8958
R18457 vdd.n3005 vdd.n2707 72.8958
R18458 vdd.n3005 vdd.n2708 72.8958
R18459 vdd.n3005 vdd.n2709 72.8958
R18460 vdd.n3005 vdd.n2710 72.8958
R18461 vdd.n3005 vdd.n2711 72.8958
R18462 vdd.n3005 vdd.n2712 72.8958
R18463 vdd.n3005 vdd.n2713 72.8958
R18464 vdd.n3005 vdd.n2714 72.8958
R18465 vdd.n3005 vdd.n2715 72.8958
R18466 vdd.n3005 vdd.n2716 72.8958
R18467 vdd.n3005 vdd.n2717 72.8958
R18468 vdd.n3183 vdd.n756 72.8958
R18469 vdd.n3189 vdd.n756 72.8958
R18470 vdd.n802 vdd.n756 72.8958
R18471 vdd.n3196 vdd.n756 72.8958
R18472 vdd.n799 vdd.n756 72.8958
R18473 vdd.n3203 vdd.n756 72.8958
R18474 vdd.n796 vdd.n756 72.8958
R18475 vdd.n3210 vdd.n756 72.8958
R18476 vdd.n793 vdd.n756 72.8958
R18477 vdd.n3218 vdd.n756 72.8958
R18478 vdd.n790 vdd.n756 72.8958
R18479 vdd.n3225 vdd.n756 72.8958
R18480 vdd.n787 vdd.n756 72.8958
R18481 vdd.n3232 vdd.n756 72.8958
R18482 vdd.n784 vdd.n756 72.8958
R18483 vdd.n3239 vdd.n756 72.8958
R18484 vdd.n3242 vdd.n756 72.8958
R18485 vdd.n2701 vdd.n950 72.8958
R18486 vdd.n2701 vdd.n949 72.8958
R18487 vdd.n2701 vdd.n948 72.8958
R18488 vdd.n2701 vdd.n947 72.8958
R18489 vdd.n2701 vdd.n946 72.8958
R18490 vdd.n2701 vdd.n945 72.8958
R18491 vdd.n2701 vdd.n944 72.8958
R18492 vdd.n2701 vdd.n943 72.8958
R18493 vdd.n2701 vdd.n942 72.8958
R18494 vdd.n2701 vdd.n941 72.8958
R18495 vdd.n2701 vdd.n940 72.8958
R18496 vdd.n2701 vdd.n939 72.8958
R18497 vdd.n2701 vdd.n938 72.8958
R18498 vdd.n2701 vdd.n937 72.8958
R18499 vdd.n2701 vdd.n936 72.8958
R18500 vdd.n2701 vdd.n935 72.8958
R18501 vdd.n2701 vdd.n934 72.8958
R18502 vdd.n2423 vdd.n1129 72.8958
R18503 vdd.n2423 vdd.n1130 72.8958
R18504 vdd.n2423 vdd.n1131 72.8958
R18505 vdd.n2423 vdd.n1132 72.8958
R18506 vdd.n2423 vdd.n1133 72.8958
R18507 vdd.n2423 vdd.n1134 72.8958
R18508 vdd.n2423 vdd.n1135 72.8958
R18509 vdd.n2423 vdd.n1136 72.8958
R18510 vdd.n2423 vdd.n1137 72.8958
R18511 vdd.n2423 vdd.n1138 72.8958
R18512 vdd.n2423 vdd.n1139 72.8958
R18513 vdd.n2423 vdd.n1140 72.8958
R18514 vdd.n2423 vdd.n1141 72.8958
R18515 vdd.n2423 vdd.n1142 72.8958
R18516 vdd.n2423 vdd.n1143 72.8958
R18517 vdd.n2423 vdd.n1144 72.8958
R18518 vdd.n2423 vdd.n1145 72.8958
R18519 vdd.n1829 vdd.n1828 66.2847
R18520 vdd.n1829 vdd.n1607 66.2847
R18521 vdd.n1829 vdd.n1608 66.2847
R18522 vdd.n1829 vdd.n1609 66.2847
R18523 vdd.n1829 vdd.n1610 66.2847
R18524 vdd.n1829 vdd.n1611 66.2847
R18525 vdd.n1829 vdd.n1612 66.2847
R18526 vdd.n1829 vdd.n1613 66.2847
R18527 vdd.n1829 vdd.n1614 66.2847
R18528 vdd.n1829 vdd.n1615 66.2847
R18529 vdd.n1829 vdd.n1616 66.2847
R18530 vdd.n1829 vdd.n1617 66.2847
R18531 vdd.n1829 vdd.n1618 66.2847
R18532 vdd.n1829 vdd.n1619 66.2847
R18533 vdd.n1829 vdd.n1620 66.2847
R18534 vdd.n1829 vdd.n1621 66.2847
R18535 vdd.n1829 vdd.n1622 66.2847
R18536 vdd.n1829 vdd.n1623 66.2847
R18537 vdd.n1829 vdd.n1624 66.2847
R18538 vdd.n1829 vdd.n1625 66.2847
R18539 vdd.n1829 vdd.n1626 66.2847
R18540 vdd.n1829 vdd.n1627 66.2847
R18541 vdd.n1829 vdd.n1628 66.2847
R18542 vdd.n1829 vdd.n1629 66.2847
R18543 vdd.n1829 vdd.n1630 66.2847
R18544 vdd.n1829 vdd.n1631 66.2847
R18545 vdd.n1829 vdd.n1632 66.2847
R18546 vdd.n1829 vdd.n1633 66.2847
R18547 vdd.n1829 vdd.n1634 66.2847
R18548 vdd.n1829 vdd.n1635 66.2847
R18549 vdd.n1829 vdd.n1636 66.2847
R18550 vdd.n1497 vdd.n1112 66.2847
R18551 vdd.n1494 vdd.n1112 66.2847
R18552 vdd.n1490 vdd.n1112 66.2847
R18553 vdd.n2289 vdd.n1112 66.2847
R18554 vdd.n1246 vdd.n1112 66.2847
R18555 vdd.n2296 vdd.n1112 66.2847
R18556 vdd.n1239 vdd.n1112 66.2847
R18557 vdd.n2303 vdd.n1112 66.2847
R18558 vdd.n1232 vdd.n1112 66.2847
R18559 vdd.n2310 vdd.n1112 66.2847
R18560 vdd.n1226 vdd.n1112 66.2847
R18561 vdd.n1221 vdd.n1112 66.2847
R18562 vdd.n2321 vdd.n1112 66.2847
R18563 vdd.n1213 vdd.n1112 66.2847
R18564 vdd.n2328 vdd.n1112 66.2847
R18565 vdd.n1206 vdd.n1112 66.2847
R18566 vdd.n2335 vdd.n1112 66.2847
R18567 vdd.n1199 vdd.n1112 66.2847
R18568 vdd.n2342 vdd.n1112 66.2847
R18569 vdd.n1192 vdd.n1112 66.2847
R18570 vdd.n2349 vdd.n1112 66.2847
R18571 vdd.n1186 vdd.n1112 66.2847
R18572 vdd.n1181 vdd.n1112 66.2847
R18573 vdd.n2360 vdd.n1112 66.2847
R18574 vdd.n1173 vdd.n1112 66.2847
R18575 vdd.n2367 vdd.n1112 66.2847
R18576 vdd.n1166 vdd.n1112 66.2847
R18577 vdd.n2374 vdd.n1112 66.2847
R18578 vdd.n1159 vdd.n1112 66.2847
R18579 vdd.n2381 vdd.n1112 66.2847
R18580 vdd.n2386 vdd.n1112 66.2847
R18581 vdd.n1155 vdd.n1112 66.2847
R18582 vdd.n3409 vdd.n658 66.2847
R18583 vdd.n663 vdd.n658 66.2847
R18584 vdd.n666 vdd.n658 66.2847
R18585 vdd.n3398 vdd.n658 66.2847
R18586 vdd.n3392 vdd.n658 66.2847
R18587 vdd.n3390 vdd.n658 66.2847
R18588 vdd.n3384 vdd.n658 66.2847
R18589 vdd.n3382 vdd.n658 66.2847
R18590 vdd.n3376 vdd.n658 66.2847
R18591 vdd.n3374 vdd.n658 66.2847
R18592 vdd.n3368 vdd.n658 66.2847
R18593 vdd.n3366 vdd.n658 66.2847
R18594 vdd.n3360 vdd.n658 66.2847
R18595 vdd.n3358 vdd.n658 66.2847
R18596 vdd.n3352 vdd.n658 66.2847
R18597 vdd.n3350 vdd.n658 66.2847
R18598 vdd.n3344 vdd.n658 66.2847
R18599 vdd.n3342 vdd.n658 66.2847
R18600 vdd.n3336 vdd.n658 66.2847
R18601 vdd.n3334 vdd.n658 66.2847
R18602 vdd.n727 vdd.n658 66.2847
R18603 vdd.n3325 vdd.n658 66.2847
R18604 vdd.n729 vdd.n658 66.2847
R18605 vdd.n3318 vdd.n658 66.2847
R18606 vdd.n3312 vdd.n658 66.2847
R18607 vdd.n3310 vdd.n658 66.2847
R18608 vdd.n3304 vdd.n658 66.2847
R18609 vdd.n3302 vdd.n658 66.2847
R18610 vdd.n3296 vdd.n658 66.2847
R18611 vdd.n750 vdd.n658 66.2847
R18612 vdd.n752 vdd.n658 66.2847
R18613 vdd.n3525 vdd.n3524 66.2847
R18614 vdd.n3525 vdd.n403 66.2847
R18615 vdd.n3525 vdd.n402 66.2847
R18616 vdd.n3525 vdd.n401 66.2847
R18617 vdd.n3525 vdd.n400 66.2847
R18618 vdd.n3525 vdd.n399 66.2847
R18619 vdd.n3525 vdd.n398 66.2847
R18620 vdd.n3525 vdd.n397 66.2847
R18621 vdd.n3525 vdd.n396 66.2847
R18622 vdd.n3525 vdd.n395 66.2847
R18623 vdd.n3525 vdd.n394 66.2847
R18624 vdd.n3525 vdd.n393 66.2847
R18625 vdd.n3525 vdd.n392 66.2847
R18626 vdd.n3525 vdd.n391 66.2847
R18627 vdd.n3525 vdd.n390 66.2847
R18628 vdd.n3525 vdd.n389 66.2847
R18629 vdd.n3525 vdd.n388 66.2847
R18630 vdd.n3525 vdd.n387 66.2847
R18631 vdd.n3525 vdd.n386 66.2847
R18632 vdd.n3525 vdd.n385 66.2847
R18633 vdd.n3525 vdd.n384 66.2847
R18634 vdd.n3525 vdd.n383 66.2847
R18635 vdd.n3525 vdd.n382 66.2847
R18636 vdd.n3525 vdd.n381 66.2847
R18637 vdd.n3525 vdd.n380 66.2847
R18638 vdd.n3525 vdd.n379 66.2847
R18639 vdd.n3525 vdd.n378 66.2847
R18640 vdd.n3525 vdd.n377 66.2847
R18641 vdd.n3525 vdd.n376 66.2847
R18642 vdd.n3525 vdd.n375 66.2847
R18643 vdd.n3525 vdd.n374 66.2847
R18644 vdd.n3525 vdd.n373 66.2847
R18645 vdd.n448 vdd.n373 52.4337
R18646 vdd.n454 vdd.n374 52.4337
R18647 vdd.n458 vdd.n375 52.4337
R18648 vdd.n464 vdd.n376 52.4337
R18649 vdd.n468 vdd.n377 52.4337
R18650 vdd.n474 vdd.n378 52.4337
R18651 vdd.n478 vdd.n379 52.4337
R18652 vdd.n484 vdd.n380 52.4337
R18653 vdd.n488 vdd.n381 52.4337
R18654 vdd.n494 vdd.n382 52.4337
R18655 vdd.n498 vdd.n383 52.4337
R18656 vdd.n504 vdd.n384 52.4337
R18657 vdd.n508 vdd.n385 52.4337
R18658 vdd.n514 vdd.n386 52.4337
R18659 vdd.n518 vdd.n387 52.4337
R18660 vdd.n524 vdd.n388 52.4337
R18661 vdd.n528 vdd.n389 52.4337
R18662 vdd.n534 vdd.n390 52.4337
R18663 vdd.n538 vdd.n391 52.4337
R18664 vdd.n544 vdd.n392 52.4337
R18665 vdd.n548 vdd.n393 52.4337
R18666 vdd.n554 vdd.n394 52.4337
R18667 vdd.n558 vdd.n395 52.4337
R18668 vdd.n564 vdd.n396 52.4337
R18669 vdd.n568 vdd.n397 52.4337
R18670 vdd.n574 vdd.n398 52.4337
R18671 vdd.n578 vdd.n399 52.4337
R18672 vdd.n584 vdd.n400 52.4337
R18673 vdd.n588 vdd.n401 52.4337
R18674 vdd.n594 vdd.n402 52.4337
R18675 vdd.n597 vdd.n403 52.4337
R18676 vdd.n3524 vdd.n3523 52.4337
R18677 vdd.n3409 vdd.n660 52.4337
R18678 vdd.n3407 vdd.n663 52.4337
R18679 vdd.n3403 vdd.n666 52.4337
R18680 vdd.n3399 vdd.n3398 52.4337
R18681 vdd.n3392 vdd.n669 52.4337
R18682 vdd.n3391 vdd.n3390 52.4337
R18683 vdd.n3384 vdd.n675 52.4337
R18684 vdd.n3383 vdd.n3382 52.4337
R18685 vdd.n3376 vdd.n681 52.4337
R18686 vdd.n3375 vdd.n3374 52.4337
R18687 vdd.n3368 vdd.n689 52.4337
R18688 vdd.n3367 vdd.n3366 52.4337
R18689 vdd.n3360 vdd.n695 52.4337
R18690 vdd.n3359 vdd.n3358 52.4337
R18691 vdd.n3352 vdd.n701 52.4337
R18692 vdd.n3351 vdd.n3350 52.4337
R18693 vdd.n3344 vdd.n707 52.4337
R18694 vdd.n3343 vdd.n3342 52.4337
R18695 vdd.n3336 vdd.n713 52.4337
R18696 vdd.n3335 vdd.n3334 52.4337
R18697 vdd.n727 vdd.n719 52.4337
R18698 vdd.n3326 vdd.n3325 52.4337
R18699 vdd.n3323 vdd.n729 52.4337
R18700 vdd.n3319 vdd.n3318 52.4337
R18701 vdd.n3312 vdd.n733 52.4337
R18702 vdd.n3311 vdd.n3310 52.4337
R18703 vdd.n3304 vdd.n739 52.4337
R18704 vdd.n3303 vdd.n3302 52.4337
R18705 vdd.n3296 vdd.n745 52.4337
R18706 vdd.n3295 vdd.n750 52.4337
R18707 vdd.n3291 vdd.n752 52.4337
R18708 vdd.n2388 vdd.n1155 52.4337
R18709 vdd.n2386 vdd.n2385 52.4337
R18710 vdd.n2381 vdd.n2380 52.4337
R18711 vdd.n2376 vdd.n1159 52.4337
R18712 vdd.n2374 vdd.n2373 52.4337
R18713 vdd.n2369 vdd.n1166 52.4337
R18714 vdd.n2367 vdd.n2366 52.4337
R18715 vdd.n2362 vdd.n1173 52.4337
R18716 vdd.n2360 vdd.n2359 52.4337
R18717 vdd.n1182 vdd.n1181 52.4337
R18718 vdd.n2351 vdd.n1186 52.4337
R18719 vdd.n2349 vdd.n2348 52.4337
R18720 vdd.n2344 vdd.n1192 52.4337
R18721 vdd.n2342 vdd.n2341 52.4337
R18722 vdd.n2337 vdd.n1199 52.4337
R18723 vdd.n2335 vdd.n2334 52.4337
R18724 vdd.n2330 vdd.n1206 52.4337
R18725 vdd.n2328 vdd.n2327 52.4337
R18726 vdd.n2323 vdd.n1213 52.4337
R18727 vdd.n2321 vdd.n2320 52.4337
R18728 vdd.n1222 vdd.n1221 52.4337
R18729 vdd.n2312 vdd.n1226 52.4337
R18730 vdd.n2310 vdd.n2309 52.4337
R18731 vdd.n2305 vdd.n1232 52.4337
R18732 vdd.n2303 vdd.n2302 52.4337
R18733 vdd.n2298 vdd.n1239 52.4337
R18734 vdd.n2296 vdd.n2295 52.4337
R18735 vdd.n2291 vdd.n1246 52.4337
R18736 vdd.n2289 vdd.n2288 52.4337
R18737 vdd.n1491 vdd.n1490 52.4337
R18738 vdd.n1495 vdd.n1494 52.4337
R18739 vdd.n2277 vdd.n1497 52.4337
R18740 vdd.n1828 vdd.n1827 52.4337
R18741 vdd.n1642 vdd.n1607 52.4337
R18742 vdd.n1644 vdd.n1608 52.4337
R18743 vdd.n1648 vdd.n1609 52.4337
R18744 vdd.n1650 vdd.n1610 52.4337
R18745 vdd.n1654 vdd.n1611 52.4337
R18746 vdd.n1656 vdd.n1612 52.4337
R18747 vdd.n1660 vdd.n1613 52.4337
R18748 vdd.n1662 vdd.n1614 52.4337
R18749 vdd.n1794 vdd.n1615 52.4337
R18750 vdd.n1666 vdd.n1616 52.4337
R18751 vdd.n1670 vdd.n1617 52.4337
R18752 vdd.n1672 vdd.n1618 52.4337
R18753 vdd.n1676 vdd.n1619 52.4337
R18754 vdd.n1678 vdd.n1620 52.4337
R18755 vdd.n1682 vdd.n1621 52.4337
R18756 vdd.n1684 vdd.n1622 52.4337
R18757 vdd.n1688 vdd.n1623 52.4337
R18758 vdd.n1690 vdd.n1624 52.4337
R18759 vdd.n1694 vdd.n1625 52.4337
R18760 vdd.n1758 vdd.n1626 52.4337
R18761 vdd.n1699 vdd.n1627 52.4337
R18762 vdd.n1701 vdd.n1628 52.4337
R18763 vdd.n1705 vdd.n1629 52.4337
R18764 vdd.n1707 vdd.n1630 52.4337
R18765 vdd.n1711 vdd.n1631 52.4337
R18766 vdd.n1713 vdd.n1632 52.4337
R18767 vdd.n1717 vdd.n1633 52.4337
R18768 vdd.n1719 vdd.n1634 52.4337
R18769 vdd.n1723 vdd.n1635 52.4337
R18770 vdd.n1725 vdd.n1636 52.4337
R18771 vdd.n1828 vdd.n1638 52.4337
R18772 vdd.n1643 vdd.n1607 52.4337
R18773 vdd.n1647 vdd.n1608 52.4337
R18774 vdd.n1649 vdd.n1609 52.4337
R18775 vdd.n1653 vdd.n1610 52.4337
R18776 vdd.n1655 vdd.n1611 52.4337
R18777 vdd.n1659 vdd.n1612 52.4337
R18778 vdd.n1661 vdd.n1613 52.4337
R18779 vdd.n1793 vdd.n1614 52.4337
R18780 vdd.n1665 vdd.n1615 52.4337
R18781 vdd.n1669 vdd.n1616 52.4337
R18782 vdd.n1671 vdd.n1617 52.4337
R18783 vdd.n1675 vdd.n1618 52.4337
R18784 vdd.n1677 vdd.n1619 52.4337
R18785 vdd.n1681 vdd.n1620 52.4337
R18786 vdd.n1683 vdd.n1621 52.4337
R18787 vdd.n1687 vdd.n1622 52.4337
R18788 vdd.n1689 vdd.n1623 52.4337
R18789 vdd.n1693 vdd.n1624 52.4337
R18790 vdd.n1695 vdd.n1625 52.4337
R18791 vdd.n1698 vdd.n1626 52.4337
R18792 vdd.n1700 vdd.n1627 52.4337
R18793 vdd.n1704 vdd.n1628 52.4337
R18794 vdd.n1706 vdd.n1629 52.4337
R18795 vdd.n1710 vdd.n1630 52.4337
R18796 vdd.n1712 vdd.n1631 52.4337
R18797 vdd.n1716 vdd.n1632 52.4337
R18798 vdd.n1718 vdd.n1633 52.4337
R18799 vdd.n1722 vdd.n1634 52.4337
R18800 vdd.n1724 vdd.n1635 52.4337
R18801 vdd.n1636 vdd.n1606 52.4337
R18802 vdd.n1497 vdd.n1496 52.4337
R18803 vdd.n1494 vdd.n1493 52.4337
R18804 vdd.n1490 vdd.n1247 52.4337
R18805 vdd.n2290 vdd.n2289 52.4337
R18806 vdd.n1246 vdd.n1240 52.4337
R18807 vdd.n2297 vdd.n2296 52.4337
R18808 vdd.n1239 vdd.n1233 52.4337
R18809 vdd.n2304 vdd.n2303 52.4337
R18810 vdd.n1232 vdd.n1227 52.4337
R18811 vdd.n2311 vdd.n2310 52.4337
R18812 vdd.n1226 vdd.n1225 52.4337
R18813 vdd.n1221 vdd.n1214 52.4337
R18814 vdd.n2322 vdd.n2321 52.4337
R18815 vdd.n1213 vdd.n1207 52.4337
R18816 vdd.n2329 vdd.n2328 52.4337
R18817 vdd.n1206 vdd.n1200 52.4337
R18818 vdd.n2336 vdd.n2335 52.4337
R18819 vdd.n1199 vdd.n1193 52.4337
R18820 vdd.n2343 vdd.n2342 52.4337
R18821 vdd.n1192 vdd.n1187 52.4337
R18822 vdd.n2350 vdd.n2349 52.4337
R18823 vdd.n1186 vdd.n1185 52.4337
R18824 vdd.n1181 vdd.n1174 52.4337
R18825 vdd.n2361 vdd.n2360 52.4337
R18826 vdd.n1173 vdd.n1167 52.4337
R18827 vdd.n2368 vdd.n2367 52.4337
R18828 vdd.n1166 vdd.n1160 52.4337
R18829 vdd.n2375 vdd.n2374 52.4337
R18830 vdd.n1159 vdd.n1156 52.4337
R18831 vdd.n2382 vdd.n2381 52.4337
R18832 vdd.n2387 vdd.n2386 52.4337
R18833 vdd.n1502 vdd.n1155 52.4337
R18834 vdd.n3410 vdd.n3409 52.4337
R18835 vdd.n3404 vdd.n663 52.4337
R18836 vdd.n3400 vdd.n666 52.4337
R18837 vdd.n3398 vdd.n3397 52.4337
R18838 vdd.n3393 vdd.n3392 52.4337
R18839 vdd.n3390 vdd.n3389 52.4337
R18840 vdd.n3385 vdd.n3384 52.4337
R18841 vdd.n3382 vdd.n3381 52.4337
R18842 vdd.n3377 vdd.n3376 52.4337
R18843 vdd.n3374 vdd.n3373 52.4337
R18844 vdd.n3369 vdd.n3368 52.4337
R18845 vdd.n3366 vdd.n3365 52.4337
R18846 vdd.n3361 vdd.n3360 52.4337
R18847 vdd.n3358 vdd.n3357 52.4337
R18848 vdd.n3353 vdd.n3352 52.4337
R18849 vdd.n3350 vdd.n3349 52.4337
R18850 vdd.n3345 vdd.n3344 52.4337
R18851 vdd.n3342 vdd.n3341 52.4337
R18852 vdd.n3337 vdd.n3336 52.4337
R18853 vdd.n3334 vdd.n3333 52.4337
R18854 vdd.n728 vdd.n727 52.4337
R18855 vdd.n3325 vdd.n3324 52.4337
R18856 vdd.n3320 vdd.n729 52.4337
R18857 vdd.n3318 vdd.n3317 52.4337
R18858 vdd.n3313 vdd.n3312 52.4337
R18859 vdd.n3310 vdd.n3309 52.4337
R18860 vdd.n3305 vdd.n3304 52.4337
R18861 vdd.n3302 vdd.n3301 52.4337
R18862 vdd.n3297 vdd.n3296 52.4337
R18863 vdd.n3292 vdd.n750 52.4337
R18864 vdd.n3288 vdd.n752 52.4337
R18865 vdd.n3524 vdd.n404 52.4337
R18866 vdd.n595 vdd.n403 52.4337
R18867 vdd.n589 vdd.n402 52.4337
R18868 vdd.n585 vdd.n401 52.4337
R18869 vdd.n579 vdd.n400 52.4337
R18870 vdd.n575 vdd.n399 52.4337
R18871 vdd.n569 vdd.n398 52.4337
R18872 vdd.n565 vdd.n397 52.4337
R18873 vdd.n559 vdd.n396 52.4337
R18874 vdd.n555 vdd.n395 52.4337
R18875 vdd.n549 vdd.n394 52.4337
R18876 vdd.n545 vdd.n393 52.4337
R18877 vdd.n539 vdd.n392 52.4337
R18878 vdd.n535 vdd.n391 52.4337
R18879 vdd.n529 vdd.n390 52.4337
R18880 vdd.n525 vdd.n389 52.4337
R18881 vdd.n519 vdd.n388 52.4337
R18882 vdd.n515 vdd.n387 52.4337
R18883 vdd.n509 vdd.n386 52.4337
R18884 vdd.n505 vdd.n385 52.4337
R18885 vdd.n499 vdd.n384 52.4337
R18886 vdd.n495 vdd.n383 52.4337
R18887 vdd.n489 vdd.n382 52.4337
R18888 vdd.n485 vdd.n381 52.4337
R18889 vdd.n479 vdd.n380 52.4337
R18890 vdd.n475 vdd.n379 52.4337
R18891 vdd.n469 vdd.n378 52.4337
R18892 vdd.n465 vdd.n377 52.4337
R18893 vdd.n459 vdd.n376 52.4337
R18894 vdd.n455 vdd.n375 52.4337
R18895 vdd.n449 vdd.n374 52.4337
R18896 vdd.n445 vdd.n373 52.4337
R18897 vdd.t17 vdd.t30 51.4683
R18898 vdd.n266 vdd.n264 42.0461
R18899 vdd.n168 vdd.n166 42.0461
R18900 vdd.n71 vdd.n69 42.0461
R18901 vdd.n2145 vdd.n2143 42.0461
R18902 vdd.n2047 vdd.n2045 42.0461
R18903 vdd.n1950 vdd.n1948 42.0461
R18904 vdd.n320 vdd.n319 41.6884
R18905 vdd.n222 vdd.n221 41.6884
R18906 vdd.n125 vdd.n124 41.6884
R18907 vdd.n2199 vdd.n2198 41.6884
R18908 vdd.n2101 vdd.n2100 41.6884
R18909 vdd.n2004 vdd.n2003 41.6884
R18910 vdd.n1605 vdd.n1604 41.1157
R18911 vdd.n1761 vdd.n1760 41.1157
R18912 vdd.n1797 vdd.n1796 41.1157
R18913 vdd.n407 vdd.n406 41.1157
R18914 vdd.n547 vdd.n420 41.1157
R18915 vdd.n433 vdd.n432 41.1157
R18916 vdd.n3242 vdd.n3241 39.2114
R18917 vdd.n3239 vdd.n3238 39.2114
R18918 vdd.n3234 vdd.n784 39.2114
R18919 vdd.n3232 vdd.n3231 39.2114
R18920 vdd.n3227 vdd.n787 39.2114
R18921 vdd.n3225 vdd.n3224 39.2114
R18922 vdd.n3220 vdd.n790 39.2114
R18923 vdd.n3218 vdd.n3217 39.2114
R18924 vdd.n3212 vdd.n793 39.2114
R18925 vdd.n3210 vdd.n3209 39.2114
R18926 vdd.n3205 vdd.n796 39.2114
R18927 vdd.n3203 vdd.n3202 39.2114
R18928 vdd.n3198 vdd.n799 39.2114
R18929 vdd.n3196 vdd.n3195 39.2114
R18930 vdd.n3191 vdd.n802 39.2114
R18931 vdd.n3189 vdd.n3188 39.2114
R18932 vdd.n3184 vdd.n3183 39.2114
R18933 vdd.n3007 vdd.n3006 39.2114
R18934 vdd.n2736 vdd.n2702 39.2114
R18935 vdd.n2999 vdd.n2703 39.2114
R18936 vdd.n2995 vdd.n2704 39.2114
R18937 vdd.n2991 vdd.n2705 39.2114
R18938 vdd.n2987 vdd.n2706 39.2114
R18939 vdd.n2983 vdd.n2707 39.2114
R18940 vdd.n2979 vdd.n2708 39.2114
R18941 vdd.n2975 vdd.n2709 39.2114
R18942 vdd.n2971 vdd.n2710 39.2114
R18943 vdd.n2967 vdd.n2711 39.2114
R18944 vdd.n2963 vdd.n2712 39.2114
R18945 vdd.n2959 vdd.n2713 39.2114
R18946 vdd.n2955 vdd.n2714 39.2114
R18947 vdd.n2951 vdd.n2715 39.2114
R18948 vdd.n2947 vdd.n2716 39.2114
R18949 vdd.n2942 vdd.n2717 39.2114
R18950 vdd.n2696 vdd.n968 39.2114
R18951 vdd.n2692 vdd.n967 39.2114
R18952 vdd.n2688 vdd.n966 39.2114
R18953 vdd.n2684 vdd.n965 39.2114
R18954 vdd.n2680 vdd.n964 39.2114
R18955 vdd.n2676 vdd.n963 39.2114
R18956 vdd.n2672 vdd.n962 39.2114
R18957 vdd.n2668 vdd.n961 39.2114
R18958 vdd.n2664 vdd.n960 39.2114
R18959 vdd.n2660 vdd.n959 39.2114
R18960 vdd.n2656 vdd.n958 39.2114
R18961 vdd.n2652 vdd.n957 39.2114
R18962 vdd.n2648 vdd.n956 39.2114
R18963 vdd.n2644 vdd.n955 39.2114
R18964 vdd.n2640 vdd.n954 39.2114
R18965 vdd.n2635 vdd.n953 39.2114
R18966 vdd.n2631 vdd.n952 39.2114
R18967 vdd.n2425 vdd.n2424 39.2114
R18968 vdd.n1147 vdd.n1113 39.2114
R18969 vdd.n2417 vdd.n1114 39.2114
R18970 vdd.n2413 vdd.n1115 39.2114
R18971 vdd.n2409 vdd.n1116 39.2114
R18972 vdd.n2405 vdd.n1117 39.2114
R18973 vdd.n2401 vdd.n1118 39.2114
R18974 vdd.n2397 vdd.n1119 39.2114
R18975 vdd.n2393 vdd.n1120 39.2114
R18976 vdd.n1293 vdd.n1121 39.2114
R18977 vdd.n1297 vdd.n1122 39.2114
R18978 vdd.n1301 vdd.n1123 39.2114
R18979 vdd.n1305 vdd.n1124 39.2114
R18980 vdd.n1309 vdd.n1125 39.2114
R18981 vdd.n1313 vdd.n1126 39.2114
R18982 vdd.n1317 vdd.n1127 39.2114
R18983 vdd.n1322 vdd.n1128 39.2114
R18984 vdd.n3161 vdd.n3160 39.2114
R18985 vdd.n3156 vdd.n3128 39.2114
R18986 vdd.n3154 vdd.n3153 39.2114
R18987 vdd.n3149 vdd.n3131 39.2114
R18988 vdd.n3147 vdd.n3146 39.2114
R18989 vdd.n3142 vdd.n3134 39.2114
R18990 vdd.n3140 vdd.n3139 39.2114
R18991 vdd.n3135 vdd.n755 39.2114
R18992 vdd.n3279 vdd.n3278 39.2114
R18993 vdd.n3276 vdd.n3275 39.2114
R18994 vdd.n3271 vdd.n760 39.2114
R18995 vdd.n3269 vdd.n3268 39.2114
R18996 vdd.n3264 vdd.n763 39.2114
R18997 vdd.n3262 vdd.n3261 39.2114
R18998 vdd.n3257 vdd.n766 39.2114
R18999 vdd.n3255 vdd.n3254 39.2114
R19000 vdd.n3250 vdd.n772 39.2114
R19001 vdd.n2743 vdd.n2718 39.2114
R19002 vdd.n2747 vdd.n2719 39.2114
R19003 vdd.n2751 vdd.n2720 39.2114
R19004 vdd.n2755 vdd.n2721 39.2114
R19005 vdd.n2759 vdd.n2722 39.2114
R19006 vdd.n2763 vdd.n2723 39.2114
R19007 vdd.n2767 vdd.n2724 39.2114
R19008 vdd.n2771 vdd.n2725 39.2114
R19009 vdd.n2775 vdd.n2726 39.2114
R19010 vdd.n2779 vdd.n2727 39.2114
R19011 vdd.n2783 vdd.n2728 39.2114
R19012 vdd.n2787 vdd.n2729 39.2114
R19013 vdd.n2791 vdd.n2730 39.2114
R19014 vdd.n2795 vdd.n2731 39.2114
R19015 vdd.n2799 vdd.n2732 39.2114
R19016 vdd.n2803 vdd.n2733 39.2114
R19017 vdd.n2807 vdd.n2734 39.2114
R19018 vdd.n2746 vdd.n2718 39.2114
R19019 vdd.n2750 vdd.n2719 39.2114
R19020 vdd.n2754 vdd.n2720 39.2114
R19021 vdd.n2758 vdd.n2721 39.2114
R19022 vdd.n2762 vdd.n2722 39.2114
R19023 vdd.n2766 vdd.n2723 39.2114
R19024 vdd.n2770 vdd.n2724 39.2114
R19025 vdd.n2774 vdd.n2725 39.2114
R19026 vdd.n2778 vdd.n2726 39.2114
R19027 vdd.n2782 vdd.n2727 39.2114
R19028 vdd.n2786 vdd.n2728 39.2114
R19029 vdd.n2790 vdd.n2729 39.2114
R19030 vdd.n2794 vdd.n2730 39.2114
R19031 vdd.n2798 vdd.n2731 39.2114
R19032 vdd.n2802 vdd.n2732 39.2114
R19033 vdd.n2806 vdd.n2733 39.2114
R19034 vdd.n2809 vdd.n2734 39.2114
R19035 vdd.n772 vdd.n767 39.2114
R19036 vdd.n3256 vdd.n3255 39.2114
R19037 vdd.n766 vdd.n764 39.2114
R19038 vdd.n3263 vdd.n3262 39.2114
R19039 vdd.n763 vdd.n761 39.2114
R19040 vdd.n3270 vdd.n3269 39.2114
R19041 vdd.n760 vdd.n758 39.2114
R19042 vdd.n3277 vdd.n3276 39.2114
R19043 vdd.n3280 vdd.n3279 39.2114
R19044 vdd.n3136 vdd.n3135 39.2114
R19045 vdd.n3141 vdd.n3140 39.2114
R19046 vdd.n3134 vdd.n3132 39.2114
R19047 vdd.n3148 vdd.n3147 39.2114
R19048 vdd.n3131 vdd.n3129 39.2114
R19049 vdd.n3155 vdd.n3154 39.2114
R19050 vdd.n3128 vdd.n3126 39.2114
R19051 vdd.n3162 vdd.n3161 39.2114
R19052 vdd.n2424 vdd.n1111 39.2114
R19053 vdd.n2418 vdd.n1113 39.2114
R19054 vdd.n2414 vdd.n1114 39.2114
R19055 vdd.n2410 vdd.n1115 39.2114
R19056 vdd.n2406 vdd.n1116 39.2114
R19057 vdd.n2402 vdd.n1117 39.2114
R19058 vdd.n2398 vdd.n1118 39.2114
R19059 vdd.n2394 vdd.n1119 39.2114
R19060 vdd.n1292 vdd.n1120 39.2114
R19061 vdd.n1296 vdd.n1121 39.2114
R19062 vdd.n1300 vdd.n1122 39.2114
R19063 vdd.n1304 vdd.n1123 39.2114
R19064 vdd.n1308 vdd.n1124 39.2114
R19065 vdd.n1312 vdd.n1125 39.2114
R19066 vdd.n1316 vdd.n1126 39.2114
R19067 vdd.n1321 vdd.n1127 39.2114
R19068 vdd.n1325 vdd.n1128 39.2114
R19069 vdd.n2634 vdd.n952 39.2114
R19070 vdd.n2639 vdd.n953 39.2114
R19071 vdd.n2643 vdd.n954 39.2114
R19072 vdd.n2647 vdd.n955 39.2114
R19073 vdd.n2651 vdd.n956 39.2114
R19074 vdd.n2655 vdd.n957 39.2114
R19075 vdd.n2659 vdd.n958 39.2114
R19076 vdd.n2663 vdd.n959 39.2114
R19077 vdd.n2667 vdd.n960 39.2114
R19078 vdd.n2671 vdd.n961 39.2114
R19079 vdd.n2675 vdd.n962 39.2114
R19080 vdd.n2679 vdd.n963 39.2114
R19081 vdd.n2683 vdd.n964 39.2114
R19082 vdd.n2687 vdd.n965 39.2114
R19083 vdd.n2691 vdd.n966 39.2114
R19084 vdd.n2695 vdd.n967 39.2114
R19085 vdd.n970 vdd.n968 39.2114
R19086 vdd.n3006 vdd.n933 39.2114
R19087 vdd.n3000 vdd.n2702 39.2114
R19088 vdd.n2996 vdd.n2703 39.2114
R19089 vdd.n2992 vdd.n2704 39.2114
R19090 vdd.n2988 vdd.n2705 39.2114
R19091 vdd.n2984 vdd.n2706 39.2114
R19092 vdd.n2980 vdd.n2707 39.2114
R19093 vdd.n2976 vdd.n2708 39.2114
R19094 vdd.n2972 vdd.n2709 39.2114
R19095 vdd.n2968 vdd.n2710 39.2114
R19096 vdd.n2964 vdd.n2711 39.2114
R19097 vdd.n2960 vdd.n2712 39.2114
R19098 vdd.n2956 vdd.n2713 39.2114
R19099 vdd.n2952 vdd.n2714 39.2114
R19100 vdd.n2948 vdd.n2715 39.2114
R19101 vdd.n2943 vdd.n2716 39.2114
R19102 vdd.n2939 vdd.n2717 39.2114
R19103 vdd.n3183 vdd.n803 39.2114
R19104 vdd.n3190 vdd.n3189 39.2114
R19105 vdd.n802 vdd.n800 39.2114
R19106 vdd.n3197 vdd.n3196 39.2114
R19107 vdd.n799 vdd.n797 39.2114
R19108 vdd.n3204 vdd.n3203 39.2114
R19109 vdd.n796 vdd.n794 39.2114
R19110 vdd.n3211 vdd.n3210 39.2114
R19111 vdd.n793 vdd.n791 39.2114
R19112 vdd.n3219 vdd.n3218 39.2114
R19113 vdd.n790 vdd.n788 39.2114
R19114 vdd.n3226 vdd.n3225 39.2114
R19115 vdd.n787 vdd.n785 39.2114
R19116 vdd.n3233 vdd.n3232 39.2114
R19117 vdd.n784 vdd.n782 39.2114
R19118 vdd.n3240 vdd.n3239 39.2114
R19119 vdd.n3243 vdd.n3242 39.2114
R19120 vdd.n979 vdd.n934 39.2114
R19121 vdd.n2623 vdd.n935 39.2114
R19122 vdd.n2619 vdd.n936 39.2114
R19123 vdd.n2615 vdd.n937 39.2114
R19124 vdd.n2611 vdd.n938 39.2114
R19125 vdd.n2607 vdd.n939 39.2114
R19126 vdd.n2603 vdd.n940 39.2114
R19127 vdd.n2599 vdd.n941 39.2114
R19128 vdd.n2595 vdd.n942 39.2114
R19129 vdd.n2591 vdd.n943 39.2114
R19130 vdd.n2587 vdd.n944 39.2114
R19131 vdd.n2583 vdd.n945 39.2114
R19132 vdd.n2579 vdd.n946 39.2114
R19133 vdd.n2575 vdd.n947 39.2114
R19134 vdd.n2571 vdd.n948 39.2114
R19135 vdd.n2567 vdd.n949 39.2114
R19136 vdd.n2563 vdd.n950 39.2114
R19137 vdd.n1251 vdd.n1129 39.2114
R19138 vdd.n1255 vdd.n1130 39.2114
R19139 vdd.n1259 vdd.n1131 39.2114
R19140 vdd.n1263 vdd.n1132 39.2114
R19141 vdd.n1267 vdd.n1133 39.2114
R19142 vdd.n1271 vdd.n1134 39.2114
R19143 vdd.n1275 vdd.n1135 39.2114
R19144 vdd.n1279 vdd.n1136 39.2114
R19145 vdd.n1283 vdd.n1137 39.2114
R19146 vdd.n1484 vdd.n1138 39.2114
R19147 vdd.n1481 vdd.n1139 39.2114
R19148 vdd.n1477 vdd.n1140 39.2114
R19149 vdd.n1473 vdd.n1141 39.2114
R19150 vdd.n1469 vdd.n1142 39.2114
R19151 vdd.n1465 vdd.n1143 39.2114
R19152 vdd.n1461 vdd.n1144 39.2114
R19153 vdd.n1457 vdd.n1145 39.2114
R19154 vdd.n2560 vdd.n950 39.2114
R19155 vdd.n2564 vdd.n949 39.2114
R19156 vdd.n2568 vdd.n948 39.2114
R19157 vdd.n2572 vdd.n947 39.2114
R19158 vdd.n2576 vdd.n946 39.2114
R19159 vdd.n2580 vdd.n945 39.2114
R19160 vdd.n2584 vdd.n944 39.2114
R19161 vdd.n2588 vdd.n943 39.2114
R19162 vdd.n2592 vdd.n942 39.2114
R19163 vdd.n2596 vdd.n941 39.2114
R19164 vdd.n2600 vdd.n940 39.2114
R19165 vdd.n2604 vdd.n939 39.2114
R19166 vdd.n2608 vdd.n938 39.2114
R19167 vdd.n2612 vdd.n937 39.2114
R19168 vdd.n2616 vdd.n936 39.2114
R19169 vdd.n2620 vdd.n935 39.2114
R19170 vdd.n2624 vdd.n934 39.2114
R19171 vdd.n1254 vdd.n1129 39.2114
R19172 vdd.n1258 vdd.n1130 39.2114
R19173 vdd.n1262 vdd.n1131 39.2114
R19174 vdd.n1266 vdd.n1132 39.2114
R19175 vdd.n1270 vdd.n1133 39.2114
R19176 vdd.n1274 vdd.n1134 39.2114
R19177 vdd.n1278 vdd.n1135 39.2114
R19178 vdd.n1282 vdd.n1136 39.2114
R19179 vdd.n1285 vdd.n1137 39.2114
R19180 vdd.n1482 vdd.n1138 39.2114
R19181 vdd.n1478 vdd.n1139 39.2114
R19182 vdd.n1474 vdd.n1140 39.2114
R19183 vdd.n1470 vdd.n1141 39.2114
R19184 vdd.n1466 vdd.n1142 39.2114
R19185 vdd.n1462 vdd.n1143 39.2114
R19186 vdd.n1458 vdd.n1144 39.2114
R19187 vdd.n1454 vdd.n1145 39.2114
R19188 vdd.n2281 vdd.n2280 37.2369
R19189 vdd.n2317 vdd.n1220 37.2369
R19190 vdd.n2356 vdd.n1180 37.2369
R19191 vdd.n3331 vdd.n724 37.2369
R19192 vdd.n688 vdd.n687 37.2369
R19193 vdd.n3287 vdd.n3286 37.2369
R19194 vdd.n1288 vdd.n1287 30.449
R19195 vdd.n983 vdd.n982 30.449
R19196 vdd.n1319 vdd.n1291 30.449
R19197 vdd.n2637 vdd.n973 30.449
R19198 vdd.n2742 vdd.n2741 30.449
R19199 vdd.n806 vdd.n805 30.449
R19200 vdd.n2945 vdd.n2738 30.449
R19201 vdd.n770 vdd.n769 30.449
R19202 vdd.n2427 vdd.n2426 29.8151
R19203 vdd.n2699 vdd.n971 29.8151
R19204 vdd.n2632 vdd.n974 29.8151
R19205 vdd.n1327 vdd.n1324 29.8151
R19206 vdd.n2940 vdd.n2937 29.8151
R19207 vdd.n3185 vdd.n3182 29.8151
R19208 vdd.n3009 vdd.n3008 29.8151
R19209 vdd.n3246 vdd.n3245 29.8151
R19210 vdd.n3165 vdd.n3164 29.8151
R19211 vdd.n3251 vdd.n771 29.8151
R19212 vdd.n2813 vdd.n2811 29.8151
R19213 vdd.n2744 vdd.n926 29.8151
R19214 vdd.n1252 vdd.n1103 29.8151
R19215 vdd.n2627 vdd.n2626 29.8151
R19216 vdd.n2559 vdd.n2558 29.8151
R19217 vdd.n1453 vdd.n1452 29.8151
R19218 vdd.n1835 vdd.n1601 19.3944
R19219 vdd.n1835 vdd.n1591 19.3944
R19220 vdd.n1847 vdd.n1591 19.3944
R19221 vdd.n1847 vdd.n1589 19.3944
R19222 vdd.n1851 vdd.n1589 19.3944
R19223 vdd.n1851 vdd.n1579 19.3944
R19224 vdd.n1864 vdd.n1579 19.3944
R19225 vdd.n1864 vdd.n1577 19.3944
R19226 vdd.n1868 vdd.n1577 19.3944
R19227 vdd.n1868 vdd.n1569 19.3944
R19228 vdd.n1881 vdd.n1569 19.3944
R19229 vdd.n1881 vdd.n1567 19.3944
R19230 vdd.n1885 vdd.n1567 19.3944
R19231 vdd.n1885 vdd.n1556 19.3944
R19232 vdd.n1897 vdd.n1556 19.3944
R19233 vdd.n1897 vdd.n1554 19.3944
R19234 vdd.n1901 vdd.n1554 19.3944
R19235 vdd.n1901 vdd.n1545 19.3944
R19236 vdd.n2209 vdd.n1545 19.3944
R19237 vdd.n2209 vdd.n1543 19.3944
R19238 vdd.n2213 vdd.n1543 19.3944
R19239 vdd.n2213 vdd.n1534 19.3944
R19240 vdd.n2225 vdd.n1534 19.3944
R19241 vdd.n2225 vdd.n1532 19.3944
R19242 vdd.n2229 vdd.n1532 19.3944
R19243 vdd.n2229 vdd.n1522 19.3944
R19244 vdd.n2242 vdd.n1522 19.3944
R19245 vdd.n2242 vdd.n1520 19.3944
R19246 vdd.n2246 vdd.n1520 19.3944
R19247 vdd.n2246 vdd.n1512 19.3944
R19248 vdd.n2259 vdd.n1512 19.3944
R19249 vdd.n2259 vdd.n1509 19.3944
R19250 vdd.n2265 vdd.n1509 19.3944
R19251 vdd.n2265 vdd.n1510 19.3944
R19252 vdd.n1510 vdd.n1499 19.3944
R19253 vdd.n1754 vdd.n1696 19.3944
R19254 vdd.n1754 vdd.n1753 19.3944
R19255 vdd.n1753 vdd.n1752 19.3944
R19256 vdd.n1752 vdd.n1702 19.3944
R19257 vdd.n1748 vdd.n1702 19.3944
R19258 vdd.n1748 vdd.n1747 19.3944
R19259 vdd.n1747 vdd.n1746 19.3944
R19260 vdd.n1746 vdd.n1708 19.3944
R19261 vdd.n1742 vdd.n1708 19.3944
R19262 vdd.n1742 vdd.n1741 19.3944
R19263 vdd.n1741 vdd.n1740 19.3944
R19264 vdd.n1740 vdd.n1714 19.3944
R19265 vdd.n1736 vdd.n1714 19.3944
R19266 vdd.n1736 vdd.n1735 19.3944
R19267 vdd.n1735 vdd.n1734 19.3944
R19268 vdd.n1734 vdd.n1720 19.3944
R19269 vdd.n1730 vdd.n1720 19.3944
R19270 vdd.n1730 vdd.n1729 19.3944
R19271 vdd.n1729 vdd.n1728 19.3944
R19272 vdd.n1728 vdd.n1726 19.3944
R19273 vdd.n1792 vdd.n1791 19.3944
R19274 vdd.n1791 vdd.n1667 19.3944
R19275 vdd.n1787 vdd.n1667 19.3944
R19276 vdd.n1787 vdd.n1786 19.3944
R19277 vdd.n1786 vdd.n1785 19.3944
R19278 vdd.n1785 vdd.n1673 19.3944
R19279 vdd.n1781 vdd.n1673 19.3944
R19280 vdd.n1781 vdd.n1780 19.3944
R19281 vdd.n1780 vdd.n1779 19.3944
R19282 vdd.n1779 vdd.n1679 19.3944
R19283 vdd.n1775 vdd.n1679 19.3944
R19284 vdd.n1775 vdd.n1774 19.3944
R19285 vdd.n1774 vdd.n1773 19.3944
R19286 vdd.n1773 vdd.n1685 19.3944
R19287 vdd.n1769 vdd.n1685 19.3944
R19288 vdd.n1769 vdd.n1768 19.3944
R19289 vdd.n1768 vdd.n1767 19.3944
R19290 vdd.n1767 vdd.n1691 19.3944
R19291 vdd.n1763 vdd.n1691 19.3944
R19292 vdd.n1763 vdd.n1762 19.3944
R19293 vdd.n1826 vdd.n1825 19.3944
R19294 vdd.n1825 vdd.n1640 19.3944
R19295 vdd.n1821 vdd.n1640 19.3944
R19296 vdd.n1821 vdd.n1820 19.3944
R19297 vdd.n1820 vdd.n1819 19.3944
R19298 vdd.n1819 vdd.n1645 19.3944
R19299 vdd.n1815 vdd.n1645 19.3944
R19300 vdd.n1815 vdd.n1814 19.3944
R19301 vdd.n1814 vdd.n1813 19.3944
R19302 vdd.n1813 vdd.n1651 19.3944
R19303 vdd.n1809 vdd.n1651 19.3944
R19304 vdd.n1809 vdd.n1808 19.3944
R19305 vdd.n1808 vdd.n1807 19.3944
R19306 vdd.n1807 vdd.n1657 19.3944
R19307 vdd.n1803 vdd.n1657 19.3944
R19308 vdd.n1803 vdd.n1802 19.3944
R19309 vdd.n1802 vdd.n1801 19.3944
R19310 vdd.n1801 vdd.n1663 19.3944
R19311 vdd.n2313 vdd.n1218 19.3944
R19312 vdd.n2313 vdd.n1224 19.3944
R19313 vdd.n2308 vdd.n1224 19.3944
R19314 vdd.n2308 vdd.n2307 19.3944
R19315 vdd.n2307 vdd.n2306 19.3944
R19316 vdd.n2306 vdd.n1231 19.3944
R19317 vdd.n2301 vdd.n1231 19.3944
R19318 vdd.n2301 vdd.n2300 19.3944
R19319 vdd.n2300 vdd.n2299 19.3944
R19320 vdd.n2299 vdd.n1238 19.3944
R19321 vdd.n2294 vdd.n1238 19.3944
R19322 vdd.n2294 vdd.n2293 19.3944
R19323 vdd.n2293 vdd.n2292 19.3944
R19324 vdd.n2292 vdd.n1245 19.3944
R19325 vdd.n2287 vdd.n1245 19.3944
R19326 vdd.n2287 vdd.n2286 19.3944
R19327 vdd.n1492 vdd.n1250 19.3944
R19328 vdd.n2282 vdd.n1489 19.3944
R19329 vdd.n2352 vdd.n1178 19.3944
R19330 vdd.n2352 vdd.n1184 19.3944
R19331 vdd.n2347 vdd.n1184 19.3944
R19332 vdd.n2347 vdd.n2346 19.3944
R19333 vdd.n2346 vdd.n2345 19.3944
R19334 vdd.n2345 vdd.n1191 19.3944
R19335 vdd.n2340 vdd.n1191 19.3944
R19336 vdd.n2340 vdd.n2339 19.3944
R19337 vdd.n2339 vdd.n2338 19.3944
R19338 vdd.n2338 vdd.n1198 19.3944
R19339 vdd.n2333 vdd.n1198 19.3944
R19340 vdd.n2333 vdd.n2332 19.3944
R19341 vdd.n2332 vdd.n2331 19.3944
R19342 vdd.n2331 vdd.n1205 19.3944
R19343 vdd.n2326 vdd.n1205 19.3944
R19344 vdd.n2326 vdd.n2325 19.3944
R19345 vdd.n2325 vdd.n2324 19.3944
R19346 vdd.n2324 vdd.n1212 19.3944
R19347 vdd.n2319 vdd.n1212 19.3944
R19348 vdd.n2319 vdd.n2318 19.3944
R19349 vdd.n2389 vdd.n1153 19.3944
R19350 vdd.n2389 vdd.n1154 19.3944
R19351 vdd.n2384 vdd.n2383 19.3944
R19352 vdd.n2379 vdd.n2378 19.3944
R19353 vdd.n2378 vdd.n2377 19.3944
R19354 vdd.n2377 vdd.n1158 19.3944
R19355 vdd.n2372 vdd.n1158 19.3944
R19356 vdd.n2372 vdd.n2371 19.3944
R19357 vdd.n2371 vdd.n2370 19.3944
R19358 vdd.n2370 vdd.n1165 19.3944
R19359 vdd.n2365 vdd.n1165 19.3944
R19360 vdd.n2365 vdd.n2364 19.3944
R19361 vdd.n2364 vdd.n2363 19.3944
R19362 vdd.n2363 vdd.n1172 19.3944
R19363 vdd.n2358 vdd.n1172 19.3944
R19364 vdd.n2358 vdd.n2357 19.3944
R19365 vdd.n1839 vdd.n1597 19.3944
R19366 vdd.n1839 vdd.n1595 19.3944
R19367 vdd.n1843 vdd.n1595 19.3944
R19368 vdd.n1843 vdd.n1585 19.3944
R19369 vdd.n1856 vdd.n1585 19.3944
R19370 vdd.n1856 vdd.n1583 19.3944
R19371 vdd.n1860 vdd.n1583 19.3944
R19372 vdd.n1860 vdd.n1574 19.3944
R19373 vdd.n1873 vdd.n1574 19.3944
R19374 vdd.n1873 vdd.n1572 19.3944
R19375 vdd.n1877 vdd.n1572 19.3944
R19376 vdd.n1877 vdd.n1563 19.3944
R19377 vdd.n1889 vdd.n1563 19.3944
R19378 vdd.n1889 vdd.n1561 19.3944
R19379 vdd.n1893 vdd.n1561 19.3944
R19380 vdd.n1893 vdd.n1551 19.3944
R19381 vdd.n1906 vdd.n1551 19.3944
R19382 vdd.n1906 vdd.n1549 19.3944
R19383 vdd.n2205 vdd.n1549 19.3944
R19384 vdd.n2205 vdd.n1540 19.3944
R19385 vdd.n2217 vdd.n1540 19.3944
R19386 vdd.n2217 vdd.n1538 19.3944
R19387 vdd.n2221 vdd.n1538 19.3944
R19388 vdd.n2221 vdd.n1528 19.3944
R19389 vdd.n2234 vdd.n1528 19.3944
R19390 vdd.n2234 vdd.n1526 19.3944
R19391 vdd.n2238 vdd.n1526 19.3944
R19392 vdd.n2238 vdd.n1517 19.3944
R19393 vdd.n2251 vdd.n1517 19.3944
R19394 vdd.n2251 vdd.n1515 19.3944
R19395 vdd.n2255 vdd.n1515 19.3944
R19396 vdd.n2255 vdd.n1505 19.3944
R19397 vdd.n2269 vdd.n1505 19.3944
R19398 vdd.n2269 vdd.n1503 19.3944
R19399 vdd.n2273 vdd.n1503 19.3944
R19400 vdd.n3419 vdd.n655 19.3944
R19401 vdd.n3423 vdd.n655 19.3944
R19402 vdd.n3423 vdd.n646 19.3944
R19403 vdd.n3435 vdd.n646 19.3944
R19404 vdd.n3435 vdd.n644 19.3944
R19405 vdd.n3439 vdd.n644 19.3944
R19406 vdd.n3439 vdd.n633 19.3944
R19407 vdd.n3451 vdd.n633 19.3944
R19408 vdd.n3451 vdd.n631 19.3944
R19409 vdd.n3455 vdd.n631 19.3944
R19410 vdd.n3455 vdd.n622 19.3944
R19411 vdd.n3468 vdd.n622 19.3944
R19412 vdd.n3468 vdd.n620 19.3944
R19413 vdd.n3475 vdd.n620 19.3944
R19414 vdd.n3475 vdd.n3474 19.3944
R19415 vdd.n3474 vdd.n610 19.3944
R19416 vdd.n3488 vdd.n610 19.3944
R19417 vdd.n3489 vdd.n3488 19.3944
R19418 vdd.n3490 vdd.n3489 19.3944
R19419 vdd.n3490 vdd.n608 19.3944
R19420 vdd.n3495 vdd.n608 19.3944
R19421 vdd.n3496 vdd.n3495 19.3944
R19422 vdd.n3497 vdd.n3496 19.3944
R19423 vdd.n3497 vdd.n606 19.3944
R19424 vdd.n3502 vdd.n606 19.3944
R19425 vdd.n3503 vdd.n3502 19.3944
R19426 vdd.n3504 vdd.n3503 19.3944
R19427 vdd.n3504 vdd.n604 19.3944
R19428 vdd.n3510 vdd.n604 19.3944
R19429 vdd.n3511 vdd.n3510 19.3944
R19430 vdd.n3512 vdd.n3511 19.3944
R19431 vdd.n3512 vdd.n602 19.3944
R19432 vdd.n3517 vdd.n602 19.3944
R19433 vdd.n3518 vdd.n3517 19.3944
R19434 vdd.n3519 vdd.n3518 19.3944
R19435 vdd.n550 vdd.n417 19.3944
R19436 vdd.n556 vdd.n417 19.3944
R19437 vdd.n557 vdd.n556 19.3944
R19438 vdd.n560 vdd.n557 19.3944
R19439 vdd.n560 vdd.n415 19.3944
R19440 vdd.n566 vdd.n415 19.3944
R19441 vdd.n567 vdd.n566 19.3944
R19442 vdd.n570 vdd.n567 19.3944
R19443 vdd.n570 vdd.n413 19.3944
R19444 vdd.n576 vdd.n413 19.3944
R19445 vdd.n577 vdd.n576 19.3944
R19446 vdd.n580 vdd.n577 19.3944
R19447 vdd.n580 vdd.n411 19.3944
R19448 vdd.n586 vdd.n411 19.3944
R19449 vdd.n587 vdd.n586 19.3944
R19450 vdd.n590 vdd.n587 19.3944
R19451 vdd.n590 vdd.n409 19.3944
R19452 vdd.n596 vdd.n409 19.3944
R19453 vdd.n598 vdd.n596 19.3944
R19454 vdd.n599 vdd.n598 19.3944
R19455 vdd.n497 vdd.n496 19.3944
R19456 vdd.n500 vdd.n497 19.3944
R19457 vdd.n500 vdd.n429 19.3944
R19458 vdd.n506 vdd.n429 19.3944
R19459 vdd.n507 vdd.n506 19.3944
R19460 vdd.n510 vdd.n507 19.3944
R19461 vdd.n510 vdd.n427 19.3944
R19462 vdd.n516 vdd.n427 19.3944
R19463 vdd.n517 vdd.n516 19.3944
R19464 vdd.n520 vdd.n517 19.3944
R19465 vdd.n520 vdd.n425 19.3944
R19466 vdd.n526 vdd.n425 19.3944
R19467 vdd.n527 vdd.n526 19.3944
R19468 vdd.n530 vdd.n527 19.3944
R19469 vdd.n530 vdd.n423 19.3944
R19470 vdd.n536 vdd.n423 19.3944
R19471 vdd.n537 vdd.n536 19.3944
R19472 vdd.n540 vdd.n537 19.3944
R19473 vdd.n540 vdd.n421 19.3944
R19474 vdd.n546 vdd.n421 19.3944
R19475 vdd.n447 vdd.n446 19.3944
R19476 vdd.n450 vdd.n447 19.3944
R19477 vdd.n450 vdd.n441 19.3944
R19478 vdd.n456 vdd.n441 19.3944
R19479 vdd.n457 vdd.n456 19.3944
R19480 vdd.n460 vdd.n457 19.3944
R19481 vdd.n460 vdd.n439 19.3944
R19482 vdd.n466 vdd.n439 19.3944
R19483 vdd.n467 vdd.n466 19.3944
R19484 vdd.n470 vdd.n467 19.3944
R19485 vdd.n470 vdd.n437 19.3944
R19486 vdd.n476 vdd.n437 19.3944
R19487 vdd.n477 vdd.n476 19.3944
R19488 vdd.n480 vdd.n477 19.3944
R19489 vdd.n480 vdd.n435 19.3944
R19490 vdd.n486 vdd.n435 19.3944
R19491 vdd.n487 vdd.n486 19.3944
R19492 vdd.n490 vdd.n487 19.3944
R19493 vdd.n3415 vdd.n652 19.3944
R19494 vdd.n3427 vdd.n652 19.3944
R19495 vdd.n3427 vdd.n650 19.3944
R19496 vdd.n3431 vdd.n650 19.3944
R19497 vdd.n3431 vdd.n640 19.3944
R19498 vdd.n3443 vdd.n640 19.3944
R19499 vdd.n3443 vdd.n638 19.3944
R19500 vdd.n3447 vdd.n638 19.3944
R19501 vdd.n3447 vdd.n628 19.3944
R19502 vdd.n3460 vdd.n628 19.3944
R19503 vdd.n3460 vdd.n626 19.3944
R19504 vdd.n3464 vdd.n626 19.3944
R19505 vdd.n3464 vdd.n617 19.3944
R19506 vdd.n3479 vdd.n617 19.3944
R19507 vdd.n3479 vdd.n615 19.3944
R19508 vdd.n3483 vdd.n615 19.3944
R19509 vdd.n3483 vdd.n324 19.3944
R19510 vdd.n3561 vdd.n324 19.3944
R19511 vdd.n3561 vdd.n325 19.3944
R19512 vdd.n3555 vdd.n325 19.3944
R19513 vdd.n3555 vdd.n3554 19.3944
R19514 vdd.n3554 vdd.n3553 19.3944
R19515 vdd.n3553 vdd.n337 19.3944
R19516 vdd.n3547 vdd.n337 19.3944
R19517 vdd.n3547 vdd.n3546 19.3944
R19518 vdd.n3546 vdd.n3545 19.3944
R19519 vdd.n3545 vdd.n347 19.3944
R19520 vdd.n3539 vdd.n347 19.3944
R19521 vdd.n3539 vdd.n3538 19.3944
R19522 vdd.n3538 vdd.n3537 19.3944
R19523 vdd.n3537 vdd.n358 19.3944
R19524 vdd.n3531 vdd.n358 19.3944
R19525 vdd.n3531 vdd.n3530 19.3944
R19526 vdd.n3530 vdd.n3529 19.3944
R19527 vdd.n3529 vdd.n369 19.3944
R19528 vdd.n3372 vdd.n3371 19.3944
R19529 vdd.n3371 vdd.n3370 19.3944
R19530 vdd.n3370 vdd.n694 19.3944
R19531 vdd.n3364 vdd.n694 19.3944
R19532 vdd.n3364 vdd.n3363 19.3944
R19533 vdd.n3363 vdd.n3362 19.3944
R19534 vdd.n3362 vdd.n700 19.3944
R19535 vdd.n3356 vdd.n700 19.3944
R19536 vdd.n3356 vdd.n3355 19.3944
R19537 vdd.n3355 vdd.n3354 19.3944
R19538 vdd.n3354 vdd.n706 19.3944
R19539 vdd.n3348 vdd.n706 19.3944
R19540 vdd.n3348 vdd.n3347 19.3944
R19541 vdd.n3347 vdd.n3346 19.3944
R19542 vdd.n3346 vdd.n712 19.3944
R19543 vdd.n3340 vdd.n712 19.3944
R19544 vdd.n3340 vdd.n3339 19.3944
R19545 vdd.n3339 vdd.n3338 19.3944
R19546 vdd.n3338 vdd.n718 19.3944
R19547 vdd.n3332 vdd.n718 19.3944
R19548 vdd.n3412 vdd.n3411 19.3944
R19549 vdd.n3411 vdd.n662 19.3944
R19550 vdd.n3406 vdd.n3405 19.3944
R19551 vdd.n3402 vdd.n3401 19.3944
R19552 vdd.n3401 vdd.n668 19.3944
R19553 vdd.n3396 vdd.n668 19.3944
R19554 vdd.n3396 vdd.n3395 19.3944
R19555 vdd.n3395 vdd.n3394 19.3944
R19556 vdd.n3394 vdd.n674 19.3944
R19557 vdd.n3388 vdd.n674 19.3944
R19558 vdd.n3388 vdd.n3387 19.3944
R19559 vdd.n3387 vdd.n3386 19.3944
R19560 vdd.n3386 vdd.n680 19.3944
R19561 vdd.n3380 vdd.n680 19.3944
R19562 vdd.n3380 vdd.n3379 19.3944
R19563 vdd.n3379 vdd.n3378 19.3944
R19564 vdd.n3327 vdd.n722 19.3944
R19565 vdd.n3327 vdd.n726 19.3944
R19566 vdd.n3322 vdd.n726 19.3944
R19567 vdd.n3322 vdd.n3321 19.3944
R19568 vdd.n3321 vdd.n732 19.3944
R19569 vdd.n3316 vdd.n732 19.3944
R19570 vdd.n3316 vdd.n3315 19.3944
R19571 vdd.n3315 vdd.n3314 19.3944
R19572 vdd.n3314 vdd.n738 19.3944
R19573 vdd.n3308 vdd.n738 19.3944
R19574 vdd.n3308 vdd.n3307 19.3944
R19575 vdd.n3307 vdd.n3306 19.3944
R19576 vdd.n3306 vdd.n744 19.3944
R19577 vdd.n3300 vdd.n744 19.3944
R19578 vdd.n3300 vdd.n3299 19.3944
R19579 vdd.n3299 vdd.n3298 19.3944
R19580 vdd.n3294 vdd.n3293 19.3944
R19581 vdd.n3290 vdd.n3289 19.3944
R19582 vdd.n1761 vdd.n1696 19.0066
R19583 vdd.n2317 vdd.n1218 19.0066
R19584 vdd.n550 vdd.n547 19.0066
R19585 vdd.n3331 vdd.n722 19.0066
R19586 vdd.n1829 vdd.n1599 18.5924
R19587 vdd.n2275 vdd.n1112 18.5924
R19588 vdd.n3417 vdd.n658 18.5924
R19589 vdd.n3526 vdd.n3525 18.5924
R19590 vdd.n1287 vdd.n1286 16.0975
R19591 vdd.n982 vdd.n981 16.0975
R19592 vdd.n1604 vdd.n1603 16.0975
R19593 vdd.n1760 vdd.n1759 16.0975
R19594 vdd.n1796 vdd.n1795 16.0975
R19595 vdd.n2280 vdd.n2279 16.0975
R19596 vdd.n1220 vdd.n1219 16.0975
R19597 vdd.n1180 vdd.n1179 16.0975
R19598 vdd.n1291 vdd.n1290 16.0975
R19599 vdd.n973 vdd.n972 16.0975
R19600 vdd.n2741 vdd.n2740 16.0975
R19601 vdd.n406 vdd.n405 16.0975
R19602 vdd.n420 vdd.n419 16.0975
R19603 vdd.n432 vdd.n431 16.0975
R19604 vdd.n724 vdd.n723 16.0975
R19605 vdd.n687 vdd.n686 16.0975
R19606 vdd.n805 vdd.n804 16.0975
R19607 vdd.n2738 vdd.n2737 16.0975
R19608 vdd.n3286 vdd.n3285 16.0975
R19609 vdd.n769 vdd.n768 16.0975
R19610 vdd.t30 vdd.n2701 15.4182
R19611 vdd.n3005 vdd.t17 15.4182
R19612 vdd.n28 vdd.n27 14.7341
R19613 vdd.n316 vdd.n281 13.1884
R19614 vdd.n261 vdd.n226 13.1884
R19615 vdd.n218 vdd.n183 13.1884
R19616 vdd.n163 vdd.n128 13.1884
R19617 vdd.n121 vdd.n86 13.1884
R19618 vdd.n66 vdd.n31 13.1884
R19619 vdd.n2140 vdd.n2105 13.1884
R19620 vdd.n2195 vdd.n2160 13.1884
R19621 vdd.n2042 vdd.n2007 13.1884
R19622 vdd.n2097 vdd.n2062 13.1884
R19623 vdd.n1945 vdd.n1910 13.1884
R19624 vdd.n2000 vdd.n1965 13.1884
R19625 vdd.n2423 vdd.n1105 13.1509
R19626 vdd.n3248 vdd.n756 13.1509
R19627 vdd.n1797 vdd.n1792 12.9944
R19628 vdd.n1797 vdd.n1663 12.9944
R19629 vdd.n2356 vdd.n1178 12.9944
R19630 vdd.n2357 vdd.n2356 12.9944
R19631 vdd.n496 vdd.n433 12.9944
R19632 vdd.n490 vdd.n433 12.9944
R19633 vdd.n3372 vdd.n688 12.9944
R19634 vdd.n3378 vdd.n688 12.9944
R19635 vdd.n317 vdd.n279 12.8005
R19636 vdd.n312 vdd.n283 12.8005
R19637 vdd.n262 vdd.n224 12.8005
R19638 vdd.n257 vdd.n228 12.8005
R19639 vdd.n219 vdd.n181 12.8005
R19640 vdd.n214 vdd.n185 12.8005
R19641 vdd.n164 vdd.n126 12.8005
R19642 vdd.n159 vdd.n130 12.8005
R19643 vdd.n122 vdd.n84 12.8005
R19644 vdd.n117 vdd.n88 12.8005
R19645 vdd.n67 vdd.n29 12.8005
R19646 vdd.n62 vdd.n33 12.8005
R19647 vdd.n2141 vdd.n2103 12.8005
R19648 vdd.n2136 vdd.n2107 12.8005
R19649 vdd.n2196 vdd.n2158 12.8005
R19650 vdd.n2191 vdd.n2162 12.8005
R19651 vdd.n2043 vdd.n2005 12.8005
R19652 vdd.n2038 vdd.n2009 12.8005
R19653 vdd.n2098 vdd.n2060 12.8005
R19654 vdd.n2093 vdd.n2064 12.8005
R19655 vdd.n1946 vdd.n1908 12.8005
R19656 vdd.n1941 vdd.n1912 12.8005
R19657 vdd.n2001 vdd.n1963 12.8005
R19658 vdd.n1996 vdd.n1967 12.8005
R19659 vdd.n311 vdd.n284 12.0247
R19660 vdd.n256 vdd.n229 12.0247
R19661 vdd.n213 vdd.n186 12.0247
R19662 vdd.n158 vdd.n131 12.0247
R19663 vdd.n116 vdd.n89 12.0247
R19664 vdd.n61 vdd.n34 12.0247
R19665 vdd.n2135 vdd.n2108 12.0247
R19666 vdd.n2190 vdd.n2163 12.0247
R19667 vdd.n2037 vdd.n2010 12.0247
R19668 vdd.n2092 vdd.n2065 12.0247
R19669 vdd.n1940 vdd.n1913 12.0247
R19670 vdd.n1995 vdd.n1968 12.0247
R19671 vdd.n1837 vdd.n1599 11.337
R19672 vdd.n1845 vdd.n1593 11.337
R19673 vdd.n1845 vdd.n1587 11.337
R19674 vdd.n1854 vdd.n1587 11.337
R19675 vdd.n1862 vdd.n1581 11.337
R19676 vdd.n1871 vdd.n1870 11.337
R19677 vdd.n1887 vdd.n1565 11.337
R19678 vdd.n1895 vdd.n1558 11.337
R19679 vdd.n1904 vdd.n1903 11.337
R19680 vdd.n2207 vdd.n1547 11.337
R19681 vdd.n2223 vdd.n1536 11.337
R19682 vdd.n2232 vdd.n1530 11.337
R19683 vdd.n2240 vdd.n1524 11.337
R19684 vdd.n2249 vdd.n2248 11.337
R19685 vdd.n2257 vdd.n1507 11.337
R19686 vdd.n2267 vdd.n1507 11.337
R19687 vdd.n2275 vdd.n1500 11.337
R19688 vdd.n3417 vdd.n659 11.337
R19689 vdd.n3425 vdd.n648 11.337
R19690 vdd.n3433 vdd.n648 11.337
R19691 vdd.n3441 vdd.n642 11.337
R19692 vdd.n3449 vdd.n635 11.337
R19693 vdd.n3458 vdd.n3457 11.337
R19694 vdd.n3466 vdd.n624 11.337
R19695 vdd.n3485 vdd.n613 11.337
R19696 vdd.n3559 vdd.n328 11.337
R19697 vdd.n3557 vdd.n332 11.337
R19698 vdd.n3551 vdd.n3550 11.337
R19699 vdd.n3543 vdd.n349 11.337
R19700 vdd.n3542 vdd.n3541 11.337
R19701 vdd.n3535 vdd.n3534 11.337
R19702 vdd.n3534 vdd.n3533 11.337
R19703 vdd.n3533 vdd.n363 11.337
R19704 vdd.n3527 vdd.n3526 11.337
R19705 vdd.n308 vdd.n307 11.249
R19706 vdd.n253 vdd.n252 11.249
R19707 vdd.n210 vdd.n209 11.249
R19708 vdd.n155 vdd.n154 11.249
R19709 vdd.n113 vdd.n112 11.249
R19710 vdd.n58 vdd.n57 11.249
R19711 vdd.n2132 vdd.n2131 11.249
R19712 vdd.n2187 vdd.n2186 11.249
R19713 vdd.n2034 vdd.n2033 11.249
R19714 vdd.n2089 vdd.n2088 11.249
R19715 vdd.n1937 vdd.n1936 11.249
R19716 vdd.n1992 vdd.n1991 11.249
R19717 vdd.n2257 vdd.t68 10.7702
R19718 vdd.n3433 vdd.t129 10.7702
R19719 vdd.n293 vdd.n292 10.7238
R19720 vdd.n238 vdd.n237 10.7238
R19721 vdd.n195 vdd.n194 10.7238
R19722 vdd.n140 vdd.n139 10.7238
R19723 vdd.n98 vdd.n97 10.7238
R19724 vdd.n43 vdd.n42 10.7238
R19725 vdd.n2117 vdd.n2116 10.7238
R19726 vdd.n2172 vdd.n2171 10.7238
R19727 vdd.n2019 vdd.n2018 10.7238
R19728 vdd.n2074 vdd.n2073 10.7238
R19729 vdd.n1922 vdd.n1921 10.7238
R19730 vdd.n1977 vdd.n1976 10.7238
R19731 vdd.n2428 vdd.n2427 10.6151
R19732 vdd.n2428 vdd.n1098 10.6151
R19733 vdd.n2438 vdd.n1098 10.6151
R19734 vdd.n2439 vdd.n2438 10.6151
R19735 vdd.n2440 vdd.n2439 10.6151
R19736 vdd.n2440 vdd.n1085 10.6151
R19737 vdd.n2450 vdd.n1085 10.6151
R19738 vdd.n2451 vdd.n2450 10.6151
R19739 vdd.n2452 vdd.n2451 10.6151
R19740 vdd.n2452 vdd.n1073 10.6151
R19741 vdd.n2462 vdd.n1073 10.6151
R19742 vdd.n2463 vdd.n2462 10.6151
R19743 vdd.n2464 vdd.n2463 10.6151
R19744 vdd.n2464 vdd.n1062 10.6151
R19745 vdd.n2474 vdd.n1062 10.6151
R19746 vdd.n2475 vdd.n2474 10.6151
R19747 vdd.n2476 vdd.n2475 10.6151
R19748 vdd.n2476 vdd.n1049 10.6151
R19749 vdd.n2486 vdd.n1049 10.6151
R19750 vdd.n2487 vdd.n2486 10.6151
R19751 vdd.n2488 vdd.n2487 10.6151
R19752 vdd.n2488 vdd.n1037 10.6151
R19753 vdd.n2499 vdd.n1037 10.6151
R19754 vdd.n2500 vdd.n2499 10.6151
R19755 vdd.n2501 vdd.n2500 10.6151
R19756 vdd.n2501 vdd.n1025 10.6151
R19757 vdd.n2511 vdd.n1025 10.6151
R19758 vdd.n2512 vdd.n2511 10.6151
R19759 vdd.n2513 vdd.n2512 10.6151
R19760 vdd.n2513 vdd.n1013 10.6151
R19761 vdd.n2523 vdd.n1013 10.6151
R19762 vdd.n2524 vdd.n2523 10.6151
R19763 vdd.n2525 vdd.n2524 10.6151
R19764 vdd.n2525 vdd.n1003 10.6151
R19765 vdd.n2535 vdd.n1003 10.6151
R19766 vdd.n2536 vdd.n2535 10.6151
R19767 vdd.n2537 vdd.n2536 10.6151
R19768 vdd.n2537 vdd.n990 10.6151
R19769 vdd.n2549 vdd.n990 10.6151
R19770 vdd.n2550 vdd.n2549 10.6151
R19771 vdd.n2552 vdd.n2550 10.6151
R19772 vdd.n2552 vdd.n2551 10.6151
R19773 vdd.n2551 vdd.n971 10.6151
R19774 vdd.n2699 vdd.n2698 10.6151
R19775 vdd.n2698 vdd.n2697 10.6151
R19776 vdd.n2697 vdd.n2694 10.6151
R19777 vdd.n2694 vdd.n2693 10.6151
R19778 vdd.n2693 vdd.n2690 10.6151
R19779 vdd.n2690 vdd.n2689 10.6151
R19780 vdd.n2689 vdd.n2686 10.6151
R19781 vdd.n2686 vdd.n2685 10.6151
R19782 vdd.n2685 vdd.n2682 10.6151
R19783 vdd.n2682 vdd.n2681 10.6151
R19784 vdd.n2681 vdd.n2678 10.6151
R19785 vdd.n2678 vdd.n2677 10.6151
R19786 vdd.n2677 vdd.n2674 10.6151
R19787 vdd.n2674 vdd.n2673 10.6151
R19788 vdd.n2673 vdd.n2670 10.6151
R19789 vdd.n2670 vdd.n2669 10.6151
R19790 vdd.n2669 vdd.n2666 10.6151
R19791 vdd.n2666 vdd.n2665 10.6151
R19792 vdd.n2665 vdd.n2662 10.6151
R19793 vdd.n2662 vdd.n2661 10.6151
R19794 vdd.n2661 vdd.n2658 10.6151
R19795 vdd.n2658 vdd.n2657 10.6151
R19796 vdd.n2657 vdd.n2654 10.6151
R19797 vdd.n2654 vdd.n2653 10.6151
R19798 vdd.n2653 vdd.n2650 10.6151
R19799 vdd.n2650 vdd.n2649 10.6151
R19800 vdd.n2649 vdd.n2646 10.6151
R19801 vdd.n2646 vdd.n2645 10.6151
R19802 vdd.n2645 vdd.n2642 10.6151
R19803 vdd.n2642 vdd.n2641 10.6151
R19804 vdd.n2641 vdd.n2638 10.6151
R19805 vdd.n2636 vdd.n2633 10.6151
R19806 vdd.n2633 vdd.n2632 10.6151
R19807 vdd.n1328 vdd.n1327 10.6151
R19808 vdd.n1330 vdd.n1328 10.6151
R19809 vdd.n1331 vdd.n1330 10.6151
R19810 vdd.n1333 vdd.n1331 10.6151
R19811 vdd.n1334 vdd.n1333 10.6151
R19812 vdd.n1336 vdd.n1334 10.6151
R19813 vdd.n1337 vdd.n1336 10.6151
R19814 vdd.n1339 vdd.n1337 10.6151
R19815 vdd.n1340 vdd.n1339 10.6151
R19816 vdd.n1342 vdd.n1340 10.6151
R19817 vdd.n1343 vdd.n1342 10.6151
R19818 vdd.n1345 vdd.n1343 10.6151
R19819 vdd.n1346 vdd.n1345 10.6151
R19820 vdd.n1348 vdd.n1346 10.6151
R19821 vdd.n1349 vdd.n1348 10.6151
R19822 vdd.n1351 vdd.n1349 10.6151
R19823 vdd.n1352 vdd.n1351 10.6151
R19824 vdd.n1354 vdd.n1352 10.6151
R19825 vdd.n1355 vdd.n1354 10.6151
R19826 vdd.n1357 vdd.n1355 10.6151
R19827 vdd.n1358 vdd.n1357 10.6151
R19828 vdd.n1360 vdd.n1358 10.6151
R19829 vdd.n1361 vdd.n1360 10.6151
R19830 vdd.n1363 vdd.n1361 10.6151
R19831 vdd.n1364 vdd.n1363 10.6151
R19832 vdd.n1366 vdd.n1364 10.6151
R19833 vdd.n1367 vdd.n1366 10.6151
R19834 vdd.n1406 vdd.n1367 10.6151
R19835 vdd.n1406 vdd.n1405 10.6151
R19836 vdd.n1405 vdd.n1404 10.6151
R19837 vdd.n1404 vdd.n1402 10.6151
R19838 vdd.n1402 vdd.n1401 10.6151
R19839 vdd.n1401 vdd.n1399 10.6151
R19840 vdd.n1399 vdd.n1398 10.6151
R19841 vdd.n1398 vdd.n1379 10.6151
R19842 vdd.n1379 vdd.n1378 10.6151
R19843 vdd.n1378 vdd.n1376 10.6151
R19844 vdd.n1376 vdd.n1375 10.6151
R19845 vdd.n1375 vdd.n1373 10.6151
R19846 vdd.n1373 vdd.n1372 10.6151
R19847 vdd.n1372 vdd.n1369 10.6151
R19848 vdd.n1369 vdd.n1368 10.6151
R19849 vdd.n1368 vdd.n974 10.6151
R19850 vdd.n2426 vdd.n1110 10.6151
R19851 vdd.n2421 vdd.n1110 10.6151
R19852 vdd.n2421 vdd.n2420 10.6151
R19853 vdd.n2420 vdd.n2419 10.6151
R19854 vdd.n2419 vdd.n2416 10.6151
R19855 vdd.n2416 vdd.n2415 10.6151
R19856 vdd.n2415 vdd.n2412 10.6151
R19857 vdd.n2412 vdd.n2411 10.6151
R19858 vdd.n2411 vdd.n2408 10.6151
R19859 vdd.n2408 vdd.n2407 10.6151
R19860 vdd.n2407 vdd.n2404 10.6151
R19861 vdd.n2404 vdd.n2403 10.6151
R19862 vdd.n2403 vdd.n2400 10.6151
R19863 vdd.n2400 vdd.n2399 10.6151
R19864 vdd.n2399 vdd.n2396 10.6151
R19865 vdd.n2396 vdd.n2395 10.6151
R19866 vdd.n2395 vdd.n2392 10.6151
R19867 vdd.n2392 vdd.n1148 10.6151
R19868 vdd.n1294 vdd.n1148 10.6151
R19869 vdd.n1295 vdd.n1294 10.6151
R19870 vdd.n1298 vdd.n1295 10.6151
R19871 vdd.n1299 vdd.n1298 10.6151
R19872 vdd.n1302 vdd.n1299 10.6151
R19873 vdd.n1303 vdd.n1302 10.6151
R19874 vdd.n1306 vdd.n1303 10.6151
R19875 vdd.n1307 vdd.n1306 10.6151
R19876 vdd.n1310 vdd.n1307 10.6151
R19877 vdd.n1311 vdd.n1310 10.6151
R19878 vdd.n1314 vdd.n1311 10.6151
R19879 vdd.n1315 vdd.n1314 10.6151
R19880 vdd.n1318 vdd.n1315 10.6151
R19881 vdd.n1323 vdd.n1320 10.6151
R19882 vdd.n1324 vdd.n1323 10.6151
R19883 vdd.n2937 vdd.n2936 10.6151
R19884 vdd.n2936 vdd.n2935 10.6151
R19885 vdd.n2935 vdd.n2739 10.6151
R19886 vdd.n2817 vdd.n2739 10.6151
R19887 vdd.n2818 vdd.n2817 10.6151
R19888 vdd.n2820 vdd.n2818 10.6151
R19889 vdd.n2821 vdd.n2820 10.6151
R19890 vdd.n2919 vdd.n2821 10.6151
R19891 vdd.n2919 vdd.n2918 10.6151
R19892 vdd.n2918 vdd.n2917 10.6151
R19893 vdd.n2917 vdd.n2865 10.6151
R19894 vdd.n2865 vdd.n2864 10.6151
R19895 vdd.n2864 vdd.n2862 10.6151
R19896 vdd.n2862 vdd.n2861 10.6151
R19897 vdd.n2861 vdd.n2859 10.6151
R19898 vdd.n2859 vdd.n2858 10.6151
R19899 vdd.n2858 vdd.n2856 10.6151
R19900 vdd.n2856 vdd.n2855 10.6151
R19901 vdd.n2855 vdd.n2853 10.6151
R19902 vdd.n2853 vdd.n2852 10.6151
R19903 vdd.n2852 vdd.n2850 10.6151
R19904 vdd.n2850 vdd.n2849 10.6151
R19905 vdd.n2849 vdd.n2847 10.6151
R19906 vdd.n2847 vdd.n2846 10.6151
R19907 vdd.n2846 vdd.n2844 10.6151
R19908 vdd.n2844 vdd.n2843 10.6151
R19909 vdd.n2843 vdd.n2841 10.6151
R19910 vdd.n2841 vdd.n2840 10.6151
R19911 vdd.n2840 vdd.n2838 10.6151
R19912 vdd.n2838 vdd.n2837 10.6151
R19913 vdd.n2837 vdd.n2835 10.6151
R19914 vdd.n2835 vdd.n2834 10.6151
R19915 vdd.n2834 vdd.n2832 10.6151
R19916 vdd.n2832 vdd.n2831 10.6151
R19917 vdd.n2831 vdd.n2829 10.6151
R19918 vdd.n2829 vdd.n2828 10.6151
R19919 vdd.n2828 vdd.n2826 10.6151
R19920 vdd.n2826 vdd.n2825 10.6151
R19921 vdd.n2825 vdd.n2823 10.6151
R19922 vdd.n2823 vdd.n2822 10.6151
R19923 vdd.n2822 vdd.n807 10.6151
R19924 vdd.n3181 vdd.n807 10.6151
R19925 vdd.n3182 vdd.n3181 10.6151
R19926 vdd.n3008 vdd.n932 10.6151
R19927 vdd.n3003 vdd.n932 10.6151
R19928 vdd.n3003 vdd.n3002 10.6151
R19929 vdd.n3002 vdd.n3001 10.6151
R19930 vdd.n3001 vdd.n2998 10.6151
R19931 vdd.n2998 vdd.n2997 10.6151
R19932 vdd.n2997 vdd.n2994 10.6151
R19933 vdd.n2994 vdd.n2993 10.6151
R19934 vdd.n2993 vdd.n2990 10.6151
R19935 vdd.n2990 vdd.n2989 10.6151
R19936 vdd.n2989 vdd.n2986 10.6151
R19937 vdd.n2986 vdd.n2985 10.6151
R19938 vdd.n2985 vdd.n2982 10.6151
R19939 vdd.n2982 vdd.n2981 10.6151
R19940 vdd.n2981 vdd.n2978 10.6151
R19941 vdd.n2978 vdd.n2977 10.6151
R19942 vdd.n2977 vdd.n2974 10.6151
R19943 vdd.n2974 vdd.n2973 10.6151
R19944 vdd.n2973 vdd.n2970 10.6151
R19945 vdd.n2970 vdd.n2969 10.6151
R19946 vdd.n2969 vdd.n2966 10.6151
R19947 vdd.n2966 vdd.n2965 10.6151
R19948 vdd.n2965 vdd.n2962 10.6151
R19949 vdd.n2962 vdd.n2961 10.6151
R19950 vdd.n2961 vdd.n2958 10.6151
R19951 vdd.n2958 vdd.n2957 10.6151
R19952 vdd.n2957 vdd.n2954 10.6151
R19953 vdd.n2954 vdd.n2953 10.6151
R19954 vdd.n2953 vdd.n2950 10.6151
R19955 vdd.n2950 vdd.n2949 10.6151
R19956 vdd.n2949 vdd.n2946 10.6151
R19957 vdd.n2944 vdd.n2941 10.6151
R19958 vdd.n2941 vdd.n2940 10.6151
R19959 vdd.n3010 vdd.n3009 10.6151
R19960 vdd.n3010 vdd.n921 10.6151
R19961 vdd.n3020 vdd.n921 10.6151
R19962 vdd.n3021 vdd.n3020 10.6151
R19963 vdd.n3022 vdd.n3021 10.6151
R19964 vdd.n3022 vdd.n909 10.6151
R19965 vdd.n3032 vdd.n909 10.6151
R19966 vdd.n3033 vdd.n3032 10.6151
R19967 vdd.n3034 vdd.n3033 10.6151
R19968 vdd.n3034 vdd.n898 10.6151
R19969 vdd.n3044 vdd.n898 10.6151
R19970 vdd.n3045 vdd.n3044 10.6151
R19971 vdd.n3046 vdd.n3045 10.6151
R19972 vdd.n3046 vdd.n887 10.6151
R19973 vdd.n3056 vdd.n887 10.6151
R19974 vdd.n3057 vdd.n3056 10.6151
R19975 vdd.n3058 vdd.n3057 10.6151
R19976 vdd.n3058 vdd.n874 10.6151
R19977 vdd.n3069 vdd.n874 10.6151
R19978 vdd.n3070 vdd.n3069 10.6151
R19979 vdd.n3071 vdd.n3070 10.6151
R19980 vdd.n3071 vdd.n862 10.6151
R19981 vdd.n3081 vdd.n862 10.6151
R19982 vdd.n3082 vdd.n3081 10.6151
R19983 vdd.n3083 vdd.n3082 10.6151
R19984 vdd.n3083 vdd.n850 10.6151
R19985 vdd.n3093 vdd.n850 10.6151
R19986 vdd.n3094 vdd.n3093 10.6151
R19987 vdd.n3095 vdd.n3094 10.6151
R19988 vdd.n3095 vdd.n837 10.6151
R19989 vdd.n3105 vdd.n837 10.6151
R19990 vdd.n3106 vdd.n3105 10.6151
R19991 vdd.n3107 vdd.n3106 10.6151
R19992 vdd.n3107 vdd.n826 10.6151
R19993 vdd.n3117 vdd.n826 10.6151
R19994 vdd.n3118 vdd.n3117 10.6151
R19995 vdd.n3119 vdd.n3118 10.6151
R19996 vdd.n3119 vdd.n812 10.6151
R19997 vdd.n3174 vdd.n812 10.6151
R19998 vdd.n3175 vdd.n3174 10.6151
R19999 vdd.n3176 vdd.n3175 10.6151
R20000 vdd.n3176 vdd.n779 10.6151
R20001 vdd.n3246 vdd.n779 10.6151
R20002 vdd.n3245 vdd.n3244 10.6151
R20003 vdd.n3244 vdd.n780 10.6151
R20004 vdd.n781 vdd.n780 10.6151
R20005 vdd.n3237 vdd.n781 10.6151
R20006 vdd.n3237 vdd.n3236 10.6151
R20007 vdd.n3236 vdd.n3235 10.6151
R20008 vdd.n3235 vdd.n783 10.6151
R20009 vdd.n3230 vdd.n783 10.6151
R20010 vdd.n3230 vdd.n3229 10.6151
R20011 vdd.n3229 vdd.n3228 10.6151
R20012 vdd.n3228 vdd.n786 10.6151
R20013 vdd.n3223 vdd.n786 10.6151
R20014 vdd.n3223 vdd.n3222 10.6151
R20015 vdd.n3222 vdd.n3221 10.6151
R20016 vdd.n3221 vdd.n789 10.6151
R20017 vdd.n3216 vdd.n789 10.6151
R20018 vdd.n3216 vdd.n3215 10.6151
R20019 vdd.n3215 vdd.n3213 10.6151
R20020 vdd.n3213 vdd.n792 10.6151
R20021 vdd.n3208 vdd.n792 10.6151
R20022 vdd.n3208 vdd.n3207 10.6151
R20023 vdd.n3207 vdd.n3206 10.6151
R20024 vdd.n3206 vdd.n795 10.6151
R20025 vdd.n3201 vdd.n795 10.6151
R20026 vdd.n3201 vdd.n3200 10.6151
R20027 vdd.n3200 vdd.n3199 10.6151
R20028 vdd.n3199 vdd.n798 10.6151
R20029 vdd.n3194 vdd.n798 10.6151
R20030 vdd.n3194 vdd.n3193 10.6151
R20031 vdd.n3193 vdd.n3192 10.6151
R20032 vdd.n3192 vdd.n801 10.6151
R20033 vdd.n3187 vdd.n3186 10.6151
R20034 vdd.n3186 vdd.n3185 10.6151
R20035 vdd.n3164 vdd.n3125 10.6151
R20036 vdd.n3159 vdd.n3125 10.6151
R20037 vdd.n3159 vdd.n3158 10.6151
R20038 vdd.n3158 vdd.n3157 10.6151
R20039 vdd.n3157 vdd.n3127 10.6151
R20040 vdd.n3152 vdd.n3127 10.6151
R20041 vdd.n3152 vdd.n3151 10.6151
R20042 vdd.n3151 vdd.n3150 10.6151
R20043 vdd.n3150 vdd.n3130 10.6151
R20044 vdd.n3145 vdd.n3130 10.6151
R20045 vdd.n3145 vdd.n3144 10.6151
R20046 vdd.n3144 vdd.n3143 10.6151
R20047 vdd.n3143 vdd.n3133 10.6151
R20048 vdd.n3138 vdd.n3133 10.6151
R20049 vdd.n3138 vdd.n3137 10.6151
R20050 vdd.n3137 vdd.n753 10.6151
R20051 vdd.n3281 vdd.n753 10.6151
R20052 vdd.n3281 vdd.n754 10.6151
R20053 vdd.n757 vdd.n754 10.6151
R20054 vdd.n3274 vdd.n757 10.6151
R20055 vdd.n3274 vdd.n3273 10.6151
R20056 vdd.n3273 vdd.n3272 10.6151
R20057 vdd.n3272 vdd.n759 10.6151
R20058 vdd.n3267 vdd.n759 10.6151
R20059 vdd.n3267 vdd.n3266 10.6151
R20060 vdd.n3266 vdd.n3265 10.6151
R20061 vdd.n3265 vdd.n762 10.6151
R20062 vdd.n3260 vdd.n762 10.6151
R20063 vdd.n3260 vdd.n3259 10.6151
R20064 vdd.n3259 vdd.n3258 10.6151
R20065 vdd.n3258 vdd.n765 10.6151
R20066 vdd.n3253 vdd.n3252 10.6151
R20067 vdd.n3252 vdd.n3251 10.6151
R20068 vdd.n2814 vdd.n2813 10.6151
R20069 vdd.n2931 vdd.n2814 10.6151
R20070 vdd.n2931 vdd.n2930 10.6151
R20071 vdd.n2930 vdd.n2929 10.6151
R20072 vdd.n2929 vdd.n2927 10.6151
R20073 vdd.n2927 vdd.n2926 10.6151
R20074 vdd.n2926 vdd.n2924 10.6151
R20075 vdd.n2924 vdd.n2923 10.6151
R20076 vdd.n2923 vdd.n2815 10.6151
R20077 vdd.n2913 vdd.n2815 10.6151
R20078 vdd.n2913 vdd.n2912 10.6151
R20079 vdd.n2912 vdd.n2911 10.6151
R20080 vdd.n2911 vdd.n2909 10.6151
R20081 vdd.n2909 vdd.n2908 10.6151
R20082 vdd.n2908 vdd.n2906 10.6151
R20083 vdd.n2906 vdd.n2905 10.6151
R20084 vdd.n2905 vdd.n2903 10.6151
R20085 vdd.n2903 vdd.n2902 10.6151
R20086 vdd.n2902 vdd.n2900 10.6151
R20087 vdd.n2900 vdd.n2899 10.6151
R20088 vdd.n2899 vdd.n2897 10.6151
R20089 vdd.n2897 vdd.n2896 10.6151
R20090 vdd.n2896 vdd.n2894 10.6151
R20091 vdd.n2894 vdd.n2893 10.6151
R20092 vdd.n2893 vdd.n2891 10.6151
R20093 vdd.n2891 vdd.n2890 10.6151
R20094 vdd.n2890 vdd.n2888 10.6151
R20095 vdd.n2888 vdd.n2887 10.6151
R20096 vdd.n2887 vdd.n2885 10.6151
R20097 vdd.n2885 vdd.n2884 10.6151
R20098 vdd.n2884 vdd.n2882 10.6151
R20099 vdd.n2882 vdd.n2881 10.6151
R20100 vdd.n2881 vdd.n2879 10.6151
R20101 vdd.n2879 vdd.n2878 10.6151
R20102 vdd.n2878 vdd.n2876 10.6151
R20103 vdd.n2876 vdd.n2875 10.6151
R20104 vdd.n2875 vdd.n2873 10.6151
R20105 vdd.n2873 vdd.n2872 10.6151
R20106 vdd.n2872 vdd.n2870 10.6151
R20107 vdd.n2870 vdd.n2869 10.6151
R20108 vdd.n2869 vdd.n2867 10.6151
R20109 vdd.n2867 vdd.n2866 10.6151
R20110 vdd.n2866 vdd.n771 10.6151
R20111 vdd.n2745 vdd.n2744 10.6151
R20112 vdd.n2748 vdd.n2745 10.6151
R20113 vdd.n2749 vdd.n2748 10.6151
R20114 vdd.n2752 vdd.n2749 10.6151
R20115 vdd.n2753 vdd.n2752 10.6151
R20116 vdd.n2756 vdd.n2753 10.6151
R20117 vdd.n2757 vdd.n2756 10.6151
R20118 vdd.n2760 vdd.n2757 10.6151
R20119 vdd.n2761 vdd.n2760 10.6151
R20120 vdd.n2764 vdd.n2761 10.6151
R20121 vdd.n2765 vdd.n2764 10.6151
R20122 vdd.n2768 vdd.n2765 10.6151
R20123 vdd.n2769 vdd.n2768 10.6151
R20124 vdd.n2772 vdd.n2769 10.6151
R20125 vdd.n2773 vdd.n2772 10.6151
R20126 vdd.n2776 vdd.n2773 10.6151
R20127 vdd.n2777 vdd.n2776 10.6151
R20128 vdd.n2780 vdd.n2777 10.6151
R20129 vdd.n2781 vdd.n2780 10.6151
R20130 vdd.n2784 vdd.n2781 10.6151
R20131 vdd.n2785 vdd.n2784 10.6151
R20132 vdd.n2788 vdd.n2785 10.6151
R20133 vdd.n2789 vdd.n2788 10.6151
R20134 vdd.n2792 vdd.n2789 10.6151
R20135 vdd.n2793 vdd.n2792 10.6151
R20136 vdd.n2796 vdd.n2793 10.6151
R20137 vdd.n2797 vdd.n2796 10.6151
R20138 vdd.n2800 vdd.n2797 10.6151
R20139 vdd.n2801 vdd.n2800 10.6151
R20140 vdd.n2804 vdd.n2801 10.6151
R20141 vdd.n2805 vdd.n2804 10.6151
R20142 vdd.n2810 vdd.n2808 10.6151
R20143 vdd.n2811 vdd.n2810 10.6151
R20144 vdd.n3014 vdd.n926 10.6151
R20145 vdd.n3015 vdd.n3014 10.6151
R20146 vdd.n3016 vdd.n3015 10.6151
R20147 vdd.n3016 vdd.n915 10.6151
R20148 vdd.n3026 vdd.n915 10.6151
R20149 vdd.n3027 vdd.n3026 10.6151
R20150 vdd.n3028 vdd.n3027 10.6151
R20151 vdd.n3028 vdd.n904 10.6151
R20152 vdd.n3038 vdd.n904 10.6151
R20153 vdd.n3039 vdd.n3038 10.6151
R20154 vdd.n3040 vdd.n3039 10.6151
R20155 vdd.n3040 vdd.n892 10.6151
R20156 vdd.n3050 vdd.n892 10.6151
R20157 vdd.n3051 vdd.n3050 10.6151
R20158 vdd.n3052 vdd.n3051 10.6151
R20159 vdd.n3052 vdd.n881 10.6151
R20160 vdd.n3062 vdd.n881 10.6151
R20161 vdd.n3063 vdd.n3062 10.6151
R20162 vdd.n3065 vdd.n3063 10.6151
R20163 vdd.n3065 vdd.n3064 10.6151
R20164 vdd.n3076 vdd.n3075 10.6151
R20165 vdd.n3077 vdd.n3076 10.6151
R20166 vdd.n3077 vdd.n856 10.6151
R20167 vdd.n3087 vdd.n856 10.6151
R20168 vdd.n3088 vdd.n3087 10.6151
R20169 vdd.n3089 vdd.n3088 10.6151
R20170 vdd.n3089 vdd.n843 10.6151
R20171 vdd.n3099 vdd.n843 10.6151
R20172 vdd.n3100 vdd.n3099 10.6151
R20173 vdd.n3101 vdd.n3100 10.6151
R20174 vdd.n3101 vdd.n831 10.6151
R20175 vdd.n3111 vdd.n831 10.6151
R20176 vdd.n3112 vdd.n3111 10.6151
R20177 vdd.n3113 vdd.n3112 10.6151
R20178 vdd.n3113 vdd.n820 10.6151
R20179 vdd.n3123 vdd.n820 10.6151
R20180 vdd.n3124 vdd.n3123 10.6151
R20181 vdd.n3170 vdd.n3124 10.6151
R20182 vdd.n3170 vdd.n3169 10.6151
R20183 vdd.n3169 vdd.n3168 10.6151
R20184 vdd.n3168 vdd.n3167 10.6151
R20185 vdd.n3167 vdd.n3165 10.6151
R20186 vdd.n2432 vdd.n1103 10.6151
R20187 vdd.n2433 vdd.n2432 10.6151
R20188 vdd.n2434 vdd.n2433 10.6151
R20189 vdd.n2434 vdd.n1092 10.6151
R20190 vdd.n2444 vdd.n1092 10.6151
R20191 vdd.n2445 vdd.n2444 10.6151
R20192 vdd.n2446 vdd.n2445 10.6151
R20193 vdd.n2446 vdd.n1079 10.6151
R20194 vdd.n2456 vdd.n1079 10.6151
R20195 vdd.n2457 vdd.n2456 10.6151
R20196 vdd.n2458 vdd.n2457 10.6151
R20197 vdd.n2458 vdd.n1068 10.6151
R20198 vdd.n2468 vdd.n1068 10.6151
R20199 vdd.n2469 vdd.n2468 10.6151
R20200 vdd.n2470 vdd.n2469 10.6151
R20201 vdd.n2470 vdd.n1056 10.6151
R20202 vdd.n2480 vdd.n1056 10.6151
R20203 vdd.n2481 vdd.n2480 10.6151
R20204 vdd.n2482 vdd.n2481 10.6151
R20205 vdd.n2482 vdd.n1043 10.6151
R20206 vdd.n2492 vdd.n1043 10.6151
R20207 vdd.n2493 vdd.n2492 10.6151
R20208 vdd.n2495 vdd.n1031 10.6151
R20209 vdd.n2505 vdd.n1031 10.6151
R20210 vdd.n2506 vdd.n2505 10.6151
R20211 vdd.n2507 vdd.n2506 10.6151
R20212 vdd.n2507 vdd.n1019 10.6151
R20213 vdd.n2517 vdd.n1019 10.6151
R20214 vdd.n2518 vdd.n2517 10.6151
R20215 vdd.n2519 vdd.n2518 10.6151
R20216 vdd.n2519 vdd.n1008 10.6151
R20217 vdd.n2529 vdd.n1008 10.6151
R20218 vdd.n2530 vdd.n2529 10.6151
R20219 vdd.n2531 vdd.n2530 10.6151
R20220 vdd.n2531 vdd.n997 10.6151
R20221 vdd.n2541 vdd.n997 10.6151
R20222 vdd.n2542 vdd.n2541 10.6151
R20223 vdd.n2545 vdd.n2542 10.6151
R20224 vdd.n2545 vdd.n2544 10.6151
R20225 vdd.n2544 vdd.n2543 10.6151
R20226 vdd.n2543 vdd.n980 10.6151
R20227 vdd.n2627 vdd.n980 10.6151
R20228 vdd.n2626 vdd.n2625 10.6151
R20229 vdd.n2625 vdd.n2622 10.6151
R20230 vdd.n2622 vdd.n2621 10.6151
R20231 vdd.n2621 vdd.n2618 10.6151
R20232 vdd.n2618 vdd.n2617 10.6151
R20233 vdd.n2617 vdd.n2614 10.6151
R20234 vdd.n2614 vdd.n2613 10.6151
R20235 vdd.n2613 vdd.n2610 10.6151
R20236 vdd.n2610 vdd.n2609 10.6151
R20237 vdd.n2609 vdd.n2606 10.6151
R20238 vdd.n2606 vdd.n2605 10.6151
R20239 vdd.n2605 vdd.n2602 10.6151
R20240 vdd.n2602 vdd.n2601 10.6151
R20241 vdd.n2601 vdd.n2598 10.6151
R20242 vdd.n2598 vdd.n2597 10.6151
R20243 vdd.n2597 vdd.n2594 10.6151
R20244 vdd.n2594 vdd.n2593 10.6151
R20245 vdd.n2593 vdd.n2590 10.6151
R20246 vdd.n2590 vdd.n2589 10.6151
R20247 vdd.n2589 vdd.n2586 10.6151
R20248 vdd.n2586 vdd.n2585 10.6151
R20249 vdd.n2585 vdd.n2582 10.6151
R20250 vdd.n2582 vdd.n2581 10.6151
R20251 vdd.n2581 vdd.n2578 10.6151
R20252 vdd.n2578 vdd.n2577 10.6151
R20253 vdd.n2577 vdd.n2574 10.6151
R20254 vdd.n2574 vdd.n2573 10.6151
R20255 vdd.n2573 vdd.n2570 10.6151
R20256 vdd.n2570 vdd.n2569 10.6151
R20257 vdd.n2569 vdd.n2566 10.6151
R20258 vdd.n2566 vdd.n2565 10.6151
R20259 vdd.n2562 vdd.n2561 10.6151
R20260 vdd.n2561 vdd.n2559 10.6151
R20261 vdd.n1452 vdd.n1450 10.6151
R20262 vdd.n1450 vdd.n1449 10.6151
R20263 vdd.n1449 vdd.n1447 10.6151
R20264 vdd.n1447 vdd.n1446 10.6151
R20265 vdd.n1446 vdd.n1444 10.6151
R20266 vdd.n1444 vdd.n1443 10.6151
R20267 vdd.n1443 vdd.n1441 10.6151
R20268 vdd.n1441 vdd.n1440 10.6151
R20269 vdd.n1440 vdd.n1438 10.6151
R20270 vdd.n1438 vdd.n1437 10.6151
R20271 vdd.n1437 vdd.n1435 10.6151
R20272 vdd.n1435 vdd.n1434 10.6151
R20273 vdd.n1434 vdd.n1432 10.6151
R20274 vdd.n1432 vdd.n1431 10.6151
R20275 vdd.n1431 vdd.n1429 10.6151
R20276 vdd.n1429 vdd.n1428 10.6151
R20277 vdd.n1428 vdd.n1426 10.6151
R20278 vdd.n1426 vdd.n1425 10.6151
R20279 vdd.n1425 vdd.n1423 10.6151
R20280 vdd.n1423 vdd.n1422 10.6151
R20281 vdd.n1422 vdd.n1420 10.6151
R20282 vdd.n1420 vdd.n1419 10.6151
R20283 vdd.n1419 vdd.n1417 10.6151
R20284 vdd.n1417 vdd.n1416 10.6151
R20285 vdd.n1416 vdd.n1414 10.6151
R20286 vdd.n1414 vdd.n1413 10.6151
R20287 vdd.n1413 vdd.n1411 10.6151
R20288 vdd.n1411 vdd.n1410 10.6151
R20289 vdd.n1410 vdd.n1289 10.6151
R20290 vdd.n1381 vdd.n1289 10.6151
R20291 vdd.n1382 vdd.n1381 10.6151
R20292 vdd.n1384 vdd.n1382 10.6151
R20293 vdd.n1385 vdd.n1384 10.6151
R20294 vdd.n1394 vdd.n1385 10.6151
R20295 vdd.n1394 vdd.n1393 10.6151
R20296 vdd.n1393 vdd.n1392 10.6151
R20297 vdd.n1392 vdd.n1390 10.6151
R20298 vdd.n1390 vdd.n1389 10.6151
R20299 vdd.n1389 vdd.n1387 10.6151
R20300 vdd.n1387 vdd.n1386 10.6151
R20301 vdd.n1386 vdd.n984 10.6151
R20302 vdd.n2557 vdd.n984 10.6151
R20303 vdd.n2558 vdd.n2557 10.6151
R20304 vdd.n1253 vdd.n1252 10.6151
R20305 vdd.n1256 vdd.n1253 10.6151
R20306 vdd.n1257 vdd.n1256 10.6151
R20307 vdd.n1260 vdd.n1257 10.6151
R20308 vdd.n1261 vdd.n1260 10.6151
R20309 vdd.n1264 vdd.n1261 10.6151
R20310 vdd.n1265 vdd.n1264 10.6151
R20311 vdd.n1268 vdd.n1265 10.6151
R20312 vdd.n1269 vdd.n1268 10.6151
R20313 vdd.n1272 vdd.n1269 10.6151
R20314 vdd.n1273 vdd.n1272 10.6151
R20315 vdd.n1276 vdd.n1273 10.6151
R20316 vdd.n1277 vdd.n1276 10.6151
R20317 vdd.n1280 vdd.n1277 10.6151
R20318 vdd.n1281 vdd.n1280 10.6151
R20319 vdd.n1284 vdd.n1281 10.6151
R20320 vdd.n1486 vdd.n1284 10.6151
R20321 vdd.n1486 vdd.n1485 10.6151
R20322 vdd.n1485 vdd.n1483 10.6151
R20323 vdd.n1483 vdd.n1480 10.6151
R20324 vdd.n1480 vdd.n1479 10.6151
R20325 vdd.n1479 vdd.n1476 10.6151
R20326 vdd.n1476 vdd.n1475 10.6151
R20327 vdd.n1475 vdd.n1472 10.6151
R20328 vdd.n1472 vdd.n1471 10.6151
R20329 vdd.n1471 vdd.n1468 10.6151
R20330 vdd.n1468 vdd.n1467 10.6151
R20331 vdd.n1467 vdd.n1464 10.6151
R20332 vdd.n1464 vdd.n1463 10.6151
R20333 vdd.n1463 vdd.n1460 10.6151
R20334 vdd.n1460 vdd.n1459 10.6151
R20335 vdd.n1456 vdd.n1455 10.6151
R20336 vdd.n1455 vdd.n1453 10.6151
R20337 vdd.t78 vdd.n2231 10.5435
R20338 vdd.n636 vdd.t87 10.5435
R20339 vdd.n304 vdd.n286 10.4732
R20340 vdd.n249 vdd.n231 10.4732
R20341 vdd.n206 vdd.n188 10.4732
R20342 vdd.n151 vdd.n133 10.4732
R20343 vdd.n109 vdd.n91 10.4732
R20344 vdd.n54 vdd.n36 10.4732
R20345 vdd.n2128 vdd.n2110 10.4732
R20346 vdd.n2183 vdd.n2165 10.4732
R20347 vdd.n2030 vdd.n2012 10.4732
R20348 vdd.n2085 vdd.n2067 10.4732
R20349 vdd.n1933 vdd.n1915 10.4732
R20350 vdd.n1988 vdd.n1970 10.4732
R20351 vdd.n2215 vdd.t66 10.3167
R20352 vdd.n3477 vdd.t127 10.3167
R20353 vdd.t134 vdd.n1559 10.09
R20354 vdd.n2267 vdd.t202 10.09
R20355 vdd.n3425 vdd.t216 10.09
R20356 vdd.n3558 vdd.t112 10.09
R20357 vdd.n2392 vdd.n2391 9.98956
R20358 vdd.n3215 vdd.n3214 9.98956
R20359 vdd.n3282 vdd.n3281 9.98956
R20360 vdd.n2284 vdd.n1486 9.98956
R20361 vdd.n1879 vdd.t152 9.86327
R20362 vdd.n3549 vdd.t104 9.86327
R20363 vdd.n2629 vdd.t50 9.7499
R20364 vdd.t35 vdd.n928 9.7499
R20365 vdd.n303 vdd.n288 9.69747
R20366 vdd.n248 vdd.n233 9.69747
R20367 vdd.n205 vdd.n190 9.69747
R20368 vdd.n150 vdd.n135 9.69747
R20369 vdd.n108 vdd.n93 9.69747
R20370 vdd.n53 vdd.n38 9.69747
R20371 vdd.n2127 vdd.n2112 9.69747
R20372 vdd.n2182 vdd.n2167 9.69747
R20373 vdd.n2029 vdd.n2014 9.69747
R20374 vdd.n2084 vdd.n2069 9.69747
R20375 vdd.n1932 vdd.n1917 9.69747
R20376 vdd.n1987 vdd.n1972 9.69747
R20377 vdd.t138 vdd.n1853 9.63654
R20378 vdd.n3508 vdd.t80 9.63654
R20379 vdd.n319 vdd.n318 9.45567
R20380 vdd.n264 vdd.n263 9.45567
R20381 vdd.n221 vdd.n220 9.45567
R20382 vdd.n166 vdd.n165 9.45567
R20383 vdd.n124 vdd.n123 9.45567
R20384 vdd.n69 vdd.n68 9.45567
R20385 vdd.n2143 vdd.n2142 9.45567
R20386 vdd.n2198 vdd.n2197 9.45567
R20387 vdd.n2045 vdd.n2044 9.45567
R20388 vdd.n2100 vdd.n2099 9.45567
R20389 vdd.n1948 vdd.n1947 9.45567
R20390 vdd.n2003 vdd.n2002 9.45567
R20391 vdd.n2354 vdd.n1178 9.3005
R20392 vdd.n2353 vdd.n2352 9.3005
R20393 vdd.n1184 vdd.n1183 9.3005
R20394 vdd.n2347 vdd.n1188 9.3005
R20395 vdd.n2346 vdd.n1189 9.3005
R20396 vdd.n2345 vdd.n1190 9.3005
R20397 vdd.n1194 vdd.n1191 9.3005
R20398 vdd.n2340 vdd.n1195 9.3005
R20399 vdd.n2339 vdd.n1196 9.3005
R20400 vdd.n2338 vdd.n1197 9.3005
R20401 vdd.n1201 vdd.n1198 9.3005
R20402 vdd.n2333 vdd.n1202 9.3005
R20403 vdd.n2332 vdd.n1203 9.3005
R20404 vdd.n2331 vdd.n1204 9.3005
R20405 vdd.n1208 vdd.n1205 9.3005
R20406 vdd.n2326 vdd.n1209 9.3005
R20407 vdd.n2325 vdd.n1210 9.3005
R20408 vdd.n2324 vdd.n1211 9.3005
R20409 vdd.n1215 vdd.n1212 9.3005
R20410 vdd.n2319 vdd.n1216 9.3005
R20411 vdd.n2318 vdd.n1217 9.3005
R20412 vdd.n2317 vdd.n2316 9.3005
R20413 vdd.n2315 vdd.n1218 9.3005
R20414 vdd.n2314 vdd.n2313 9.3005
R20415 vdd.n1224 vdd.n1223 9.3005
R20416 vdd.n2308 vdd.n1228 9.3005
R20417 vdd.n2307 vdd.n1229 9.3005
R20418 vdd.n2306 vdd.n1230 9.3005
R20419 vdd.n1234 vdd.n1231 9.3005
R20420 vdd.n2301 vdd.n1235 9.3005
R20421 vdd.n2300 vdd.n1236 9.3005
R20422 vdd.n2299 vdd.n1237 9.3005
R20423 vdd.n1241 vdd.n1238 9.3005
R20424 vdd.n2294 vdd.n1242 9.3005
R20425 vdd.n2293 vdd.n1243 9.3005
R20426 vdd.n2292 vdd.n1244 9.3005
R20427 vdd.n1248 vdd.n1245 9.3005
R20428 vdd.n2287 vdd.n1249 9.3005
R20429 vdd.n2356 vdd.n2355 9.3005
R20430 vdd.n2378 vdd.n1149 9.3005
R20431 vdd.n2377 vdd.n1157 9.3005
R20432 vdd.n1161 vdd.n1158 9.3005
R20433 vdd.n2372 vdd.n1162 9.3005
R20434 vdd.n2371 vdd.n1163 9.3005
R20435 vdd.n2370 vdd.n1164 9.3005
R20436 vdd.n1168 vdd.n1165 9.3005
R20437 vdd.n2365 vdd.n1169 9.3005
R20438 vdd.n2364 vdd.n1170 9.3005
R20439 vdd.n2363 vdd.n1171 9.3005
R20440 vdd.n1175 vdd.n1172 9.3005
R20441 vdd.n2358 vdd.n1176 9.3005
R20442 vdd.n2357 vdd.n1177 9.3005
R20443 vdd.n2390 vdd.n2389 9.3005
R20444 vdd.n1153 vdd.n1152 9.3005
R20445 vdd.n2203 vdd.n1549 9.3005
R20446 vdd.n2205 vdd.n2204 9.3005
R20447 vdd.n1540 vdd.n1539 9.3005
R20448 vdd.n2218 vdd.n2217 9.3005
R20449 vdd.n2219 vdd.n1538 9.3005
R20450 vdd.n2221 vdd.n2220 9.3005
R20451 vdd.n1528 vdd.n1527 9.3005
R20452 vdd.n2235 vdd.n2234 9.3005
R20453 vdd.n2236 vdd.n1526 9.3005
R20454 vdd.n2238 vdd.n2237 9.3005
R20455 vdd.n1517 vdd.n1516 9.3005
R20456 vdd.n2252 vdd.n2251 9.3005
R20457 vdd.n2253 vdd.n1515 9.3005
R20458 vdd.n2255 vdd.n2254 9.3005
R20459 vdd.n1505 vdd.n1504 9.3005
R20460 vdd.n2270 vdd.n2269 9.3005
R20461 vdd.n2271 vdd.n1503 9.3005
R20462 vdd.n2273 vdd.n2272 9.3005
R20463 vdd.n295 vdd.n294 9.3005
R20464 vdd.n290 vdd.n289 9.3005
R20465 vdd.n301 vdd.n300 9.3005
R20466 vdd.n303 vdd.n302 9.3005
R20467 vdd.n286 vdd.n285 9.3005
R20468 vdd.n309 vdd.n308 9.3005
R20469 vdd.n311 vdd.n310 9.3005
R20470 vdd.n283 vdd.n280 9.3005
R20471 vdd.n318 vdd.n317 9.3005
R20472 vdd.n240 vdd.n239 9.3005
R20473 vdd.n235 vdd.n234 9.3005
R20474 vdd.n246 vdd.n245 9.3005
R20475 vdd.n248 vdd.n247 9.3005
R20476 vdd.n231 vdd.n230 9.3005
R20477 vdd.n254 vdd.n253 9.3005
R20478 vdd.n256 vdd.n255 9.3005
R20479 vdd.n228 vdd.n225 9.3005
R20480 vdd.n263 vdd.n262 9.3005
R20481 vdd.n197 vdd.n196 9.3005
R20482 vdd.n192 vdd.n191 9.3005
R20483 vdd.n203 vdd.n202 9.3005
R20484 vdd.n205 vdd.n204 9.3005
R20485 vdd.n188 vdd.n187 9.3005
R20486 vdd.n211 vdd.n210 9.3005
R20487 vdd.n213 vdd.n212 9.3005
R20488 vdd.n185 vdd.n182 9.3005
R20489 vdd.n220 vdd.n219 9.3005
R20490 vdd.n142 vdd.n141 9.3005
R20491 vdd.n137 vdd.n136 9.3005
R20492 vdd.n148 vdd.n147 9.3005
R20493 vdd.n150 vdd.n149 9.3005
R20494 vdd.n133 vdd.n132 9.3005
R20495 vdd.n156 vdd.n155 9.3005
R20496 vdd.n158 vdd.n157 9.3005
R20497 vdd.n130 vdd.n127 9.3005
R20498 vdd.n165 vdd.n164 9.3005
R20499 vdd.n100 vdd.n99 9.3005
R20500 vdd.n95 vdd.n94 9.3005
R20501 vdd.n106 vdd.n105 9.3005
R20502 vdd.n108 vdd.n107 9.3005
R20503 vdd.n91 vdd.n90 9.3005
R20504 vdd.n114 vdd.n113 9.3005
R20505 vdd.n116 vdd.n115 9.3005
R20506 vdd.n88 vdd.n85 9.3005
R20507 vdd.n123 vdd.n122 9.3005
R20508 vdd.n45 vdd.n44 9.3005
R20509 vdd.n40 vdd.n39 9.3005
R20510 vdd.n51 vdd.n50 9.3005
R20511 vdd.n53 vdd.n52 9.3005
R20512 vdd.n36 vdd.n35 9.3005
R20513 vdd.n59 vdd.n58 9.3005
R20514 vdd.n61 vdd.n60 9.3005
R20515 vdd.n33 vdd.n30 9.3005
R20516 vdd.n68 vdd.n67 9.3005
R20517 vdd.n3331 vdd.n3330 9.3005
R20518 vdd.n3332 vdd.n721 9.3005
R20519 vdd.n720 vdd.n718 9.3005
R20520 vdd.n3338 vdd.n717 9.3005
R20521 vdd.n3339 vdd.n716 9.3005
R20522 vdd.n3340 vdd.n715 9.3005
R20523 vdd.n714 vdd.n712 9.3005
R20524 vdd.n3346 vdd.n711 9.3005
R20525 vdd.n3347 vdd.n710 9.3005
R20526 vdd.n3348 vdd.n709 9.3005
R20527 vdd.n708 vdd.n706 9.3005
R20528 vdd.n3354 vdd.n705 9.3005
R20529 vdd.n3355 vdd.n704 9.3005
R20530 vdd.n3356 vdd.n703 9.3005
R20531 vdd.n702 vdd.n700 9.3005
R20532 vdd.n3362 vdd.n699 9.3005
R20533 vdd.n3363 vdd.n698 9.3005
R20534 vdd.n3364 vdd.n697 9.3005
R20535 vdd.n696 vdd.n694 9.3005
R20536 vdd.n3370 vdd.n693 9.3005
R20537 vdd.n3371 vdd.n692 9.3005
R20538 vdd.n3372 vdd.n691 9.3005
R20539 vdd.n690 vdd.n688 9.3005
R20540 vdd.n3378 vdd.n685 9.3005
R20541 vdd.n3379 vdd.n684 9.3005
R20542 vdd.n3380 vdd.n683 9.3005
R20543 vdd.n682 vdd.n680 9.3005
R20544 vdd.n3386 vdd.n679 9.3005
R20545 vdd.n3387 vdd.n678 9.3005
R20546 vdd.n3388 vdd.n677 9.3005
R20547 vdd.n676 vdd.n674 9.3005
R20548 vdd.n3394 vdd.n673 9.3005
R20549 vdd.n3395 vdd.n672 9.3005
R20550 vdd.n3396 vdd.n671 9.3005
R20551 vdd.n670 vdd.n668 9.3005
R20552 vdd.n3401 vdd.n667 9.3005
R20553 vdd.n3411 vdd.n661 9.3005
R20554 vdd.n3413 vdd.n3412 9.3005
R20555 vdd.n652 vdd.n651 9.3005
R20556 vdd.n3428 vdd.n3427 9.3005
R20557 vdd.n3429 vdd.n650 9.3005
R20558 vdd.n3431 vdd.n3430 9.3005
R20559 vdd.n640 vdd.n639 9.3005
R20560 vdd.n3444 vdd.n3443 9.3005
R20561 vdd.n3445 vdd.n638 9.3005
R20562 vdd.n3447 vdd.n3446 9.3005
R20563 vdd.n628 vdd.n627 9.3005
R20564 vdd.n3461 vdd.n3460 9.3005
R20565 vdd.n3462 vdd.n626 9.3005
R20566 vdd.n3464 vdd.n3463 9.3005
R20567 vdd.n617 vdd.n616 9.3005
R20568 vdd.n3480 vdd.n3479 9.3005
R20569 vdd.n3481 vdd.n615 9.3005
R20570 vdd.n3483 vdd.n3482 9.3005
R20571 vdd.n324 vdd.n322 9.3005
R20572 vdd.n3415 vdd.n3414 9.3005
R20573 vdd.n3562 vdd.n3561 9.3005
R20574 vdd.n325 vdd.n323 9.3005
R20575 vdd.n3555 vdd.n334 9.3005
R20576 vdd.n3554 vdd.n335 9.3005
R20577 vdd.n3553 vdd.n336 9.3005
R20578 vdd.n343 vdd.n337 9.3005
R20579 vdd.n3547 vdd.n344 9.3005
R20580 vdd.n3546 vdd.n345 9.3005
R20581 vdd.n3545 vdd.n346 9.3005
R20582 vdd.n354 vdd.n347 9.3005
R20583 vdd.n3539 vdd.n355 9.3005
R20584 vdd.n3538 vdd.n356 9.3005
R20585 vdd.n3537 vdd.n357 9.3005
R20586 vdd.n365 vdd.n358 9.3005
R20587 vdd.n3531 vdd.n366 9.3005
R20588 vdd.n3530 vdd.n367 9.3005
R20589 vdd.n3529 vdd.n368 9.3005
R20590 vdd.n443 vdd.n369 9.3005
R20591 vdd.n447 vdd.n442 9.3005
R20592 vdd.n451 vdd.n450 9.3005
R20593 vdd.n452 vdd.n441 9.3005
R20594 vdd.n456 vdd.n453 9.3005
R20595 vdd.n457 vdd.n440 9.3005
R20596 vdd.n461 vdd.n460 9.3005
R20597 vdd.n462 vdd.n439 9.3005
R20598 vdd.n466 vdd.n463 9.3005
R20599 vdd.n467 vdd.n438 9.3005
R20600 vdd.n471 vdd.n470 9.3005
R20601 vdd.n472 vdd.n437 9.3005
R20602 vdd.n476 vdd.n473 9.3005
R20603 vdd.n477 vdd.n436 9.3005
R20604 vdd.n481 vdd.n480 9.3005
R20605 vdd.n482 vdd.n435 9.3005
R20606 vdd.n486 vdd.n483 9.3005
R20607 vdd.n487 vdd.n434 9.3005
R20608 vdd.n491 vdd.n490 9.3005
R20609 vdd.n492 vdd.n433 9.3005
R20610 vdd.n496 vdd.n493 9.3005
R20611 vdd.n497 vdd.n430 9.3005
R20612 vdd.n501 vdd.n500 9.3005
R20613 vdd.n502 vdd.n429 9.3005
R20614 vdd.n506 vdd.n503 9.3005
R20615 vdd.n507 vdd.n428 9.3005
R20616 vdd.n511 vdd.n510 9.3005
R20617 vdd.n512 vdd.n427 9.3005
R20618 vdd.n516 vdd.n513 9.3005
R20619 vdd.n517 vdd.n426 9.3005
R20620 vdd.n521 vdd.n520 9.3005
R20621 vdd.n522 vdd.n425 9.3005
R20622 vdd.n526 vdd.n523 9.3005
R20623 vdd.n527 vdd.n424 9.3005
R20624 vdd.n531 vdd.n530 9.3005
R20625 vdd.n532 vdd.n423 9.3005
R20626 vdd.n536 vdd.n533 9.3005
R20627 vdd.n537 vdd.n422 9.3005
R20628 vdd.n541 vdd.n540 9.3005
R20629 vdd.n542 vdd.n421 9.3005
R20630 vdd.n546 vdd.n543 9.3005
R20631 vdd.n547 vdd.n418 9.3005
R20632 vdd.n551 vdd.n550 9.3005
R20633 vdd.n552 vdd.n417 9.3005
R20634 vdd.n556 vdd.n553 9.3005
R20635 vdd.n557 vdd.n416 9.3005
R20636 vdd.n561 vdd.n560 9.3005
R20637 vdd.n562 vdd.n415 9.3005
R20638 vdd.n566 vdd.n563 9.3005
R20639 vdd.n567 vdd.n414 9.3005
R20640 vdd.n571 vdd.n570 9.3005
R20641 vdd.n572 vdd.n413 9.3005
R20642 vdd.n576 vdd.n573 9.3005
R20643 vdd.n577 vdd.n412 9.3005
R20644 vdd.n581 vdd.n580 9.3005
R20645 vdd.n582 vdd.n411 9.3005
R20646 vdd.n586 vdd.n583 9.3005
R20647 vdd.n587 vdd.n410 9.3005
R20648 vdd.n591 vdd.n590 9.3005
R20649 vdd.n592 vdd.n409 9.3005
R20650 vdd.n596 vdd.n593 9.3005
R20651 vdd.n598 vdd.n408 9.3005
R20652 vdd.n600 vdd.n599 9.3005
R20653 vdd.n3522 vdd.n3521 9.3005
R20654 vdd.n446 vdd.n444 9.3005
R20655 vdd.n3421 vdd.n655 9.3005
R20656 vdd.n3423 vdd.n3422 9.3005
R20657 vdd.n646 vdd.n645 9.3005
R20658 vdd.n3436 vdd.n3435 9.3005
R20659 vdd.n3437 vdd.n644 9.3005
R20660 vdd.n3439 vdd.n3438 9.3005
R20661 vdd.n633 vdd.n632 9.3005
R20662 vdd.n3452 vdd.n3451 9.3005
R20663 vdd.n3453 vdd.n631 9.3005
R20664 vdd.n3455 vdd.n3454 9.3005
R20665 vdd.n622 vdd.n621 9.3005
R20666 vdd.n3469 vdd.n3468 9.3005
R20667 vdd.n3470 vdd.n620 9.3005
R20668 vdd.n3475 vdd.n3471 9.3005
R20669 vdd.n3474 vdd.n3473 9.3005
R20670 vdd.n3472 vdd.n610 9.3005
R20671 vdd.n3488 vdd.n611 9.3005
R20672 vdd.n3489 vdd.n609 9.3005
R20673 vdd.n3491 vdd.n3490 9.3005
R20674 vdd.n3492 vdd.n608 9.3005
R20675 vdd.n3495 vdd.n3493 9.3005
R20676 vdd.n3496 vdd.n607 9.3005
R20677 vdd.n3498 vdd.n3497 9.3005
R20678 vdd.n3499 vdd.n606 9.3005
R20679 vdd.n3502 vdd.n3500 9.3005
R20680 vdd.n3503 vdd.n605 9.3005
R20681 vdd.n3505 vdd.n3504 9.3005
R20682 vdd.n3506 vdd.n604 9.3005
R20683 vdd.n3510 vdd.n3507 9.3005
R20684 vdd.n3511 vdd.n603 9.3005
R20685 vdd.n3513 vdd.n3512 9.3005
R20686 vdd.n3514 vdd.n602 9.3005
R20687 vdd.n3517 vdd.n3515 9.3005
R20688 vdd.n3518 vdd.n601 9.3005
R20689 vdd.n3520 vdd.n3519 9.3005
R20690 vdd.n3420 vdd.n3419 9.3005
R20691 vdd.n3284 vdd.n656 9.3005
R20692 vdd.n3289 vdd.n3283 9.3005
R20693 vdd.n3299 vdd.n748 9.3005
R20694 vdd.n3300 vdd.n747 9.3005
R20695 vdd.n746 vdd.n744 9.3005
R20696 vdd.n3306 vdd.n743 9.3005
R20697 vdd.n3307 vdd.n742 9.3005
R20698 vdd.n3308 vdd.n741 9.3005
R20699 vdd.n740 vdd.n738 9.3005
R20700 vdd.n3314 vdd.n737 9.3005
R20701 vdd.n3315 vdd.n736 9.3005
R20702 vdd.n3316 vdd.n735 9.3005
R20703 vdd.n734 vdd.n732 9.3005
R20704 vdd.n3321 vdd.n731 9.3005
R20705 vdd.n3322 vdd.n730 9.3005
R20706 vdd.n726 vdd.n725 9.3005
R20707 vdd.n3328 vdd.n3327 9.3005
R20708 vdd.n3329 vdd.n722 9.3005
R20709 vdd.n2283 vdd.n2282 9.3005
R20710 vdd.n2278 vdd.n1488 9.3005
R20711 vdd.n1835 vdd.n1834 9.3005
R20712 vdd.n1591 vdd.n1590 9.3005
R20713 vdd.n1848 vdd.n1847 9.3005
R20714 vdd.n1849 vdd.n1589 9.3005
R20715 vdd.n1851 vdd.n1850 9.3005
R20716 vdd.n1579 vdd.n1578 9.3005
R20717 vdd.n1865 vdd.n1864 9.3005
R20718 vdd.n1866 vdd.n1577 9.3005
R20719 vdd.n1868 vdd.n1867 9.3005
R20720 vdd.n1569 vdd.n1568 9.3005
R20721 vdd.n1882 vdd.n1881 9.3005
R20722 vdd.n1883 vdd.n1567 9.3005
R20723 vdd.n1885 vdd.n1884 9.3005
R20724 vdd.n1556 vdd.n1555 9.3005
R20725 vdd.n1898 vdd.n1897 9.3005
R20726 vdd.n1899 vdd.n1554 9.3005
R20727 vdd.n1901 vdd.n1900 9.3005
R20728 vdd.n1545 vdd.n1544 9.3005
R20729 vdd.n2210 vdd.n2209 9.3005
R20730 vdd.n2211 vdd.n1543 9.3005
R20731 vdd.n2213 vdd.n2212 9.3005
R20732 vdd.n1534 vdd.n1533 9.3005
R20733 vdd.n2226 vdd.n2225 9.3005
R20734 vdd.n2227 vdd.n1532 9.3005
R20735 vdd.n2229 vdd.n2228 9.3005
R20736 vdd.n1522 vdd.n1521 9.3005
R20737 vdd.n2243 vdd.n2242 9.3005
R20738 vdd.n2244 vdd.n1520 9.3005
R20739 vdd.n2246 vdd.n2245 9.3005
R20740 vdd.n1512 vdd.n1511 9.3005
R20741 vdd.n2260 vdd.n2259 9.3005
R20742 vdd.n2261 vdd.n1509 9.3005
R20743 vdd.n2265 vdd.n2264 9.3005
R20744 vdd.n2263 vdd.n1510 9.3005
R20745 vdd.n2262 vdd.n1499 9.3005
R20746 vdd.n1833 vdd.n1601 9.3005
R20747 vdd.n1726 vdd.n1602 9.3005
R20748 vdd.n1728 vdd.n1727 9.3005
R20749 vdd.n1729 vdd.n1721 9.3005
R20750 vdd.n1731 vdd.n1730 9.3005
R20751 vdd.n1732 vdd.n1720 9.3005
R20752 vdd.n1734 vdd.n1733 9.3005
R20753 vdd.n1735 vdd.n1715 9.3005
R20754 vdd.n1737 vdd.n1736 9.3005
R20755 vdd.n1738 vdd.n1714 9.3005
R20756 vdd.n1740 vdd.n1739 9.3005
R20757 vdd.n1741 vdd.n1709 9.3005
R20758 vdd.n1743 vdd.n1742 9.3005
R20759 vdd.n1744 vdd.n1708 9.3005
R20760 vdd.n1746 vdd.n1745 9.3005
R20761 vdd.n1747 vdd.n1703 9.3005
R20762 vdd.n1749 vdd.n1748 9.3005
R20763 vdd.n1750 vdd.n1702 9.3005
R20764 vdd.n1752 vdd.n1751 9.3005
R20765 vdd.n1753 vdd.n1697 9.3005
R20766 vdd.n1755 vdd.n1754 9.3005
R20767 vdd.n1756 vdd.n1696 9.3005
R20768 vdd.n1761 vdd.n1757 9.3005
R20769 vdd.n1762 vdd.n1692 9.3005
R20770 vdd.n1764 vdd.n1763 9.3005
R20771 vdd.n1765 vdd.n1691 9.3005
R20772 vdd.n1767 vdd.n1766 9.3005
R20773 vdd.n1768 vdd.n1686 9.3005
R20774 vdd.n1770 vdd.n1769 9.3005
R20775 vdd.n1771 vdd.n1685 9.3005
R20776 vdd.n1773 vdd.n1772 9.3005
R20777 vdd.n1774 vdd.n1680 9.3005
R20778 vdd.n1776 vdd.n1775 9.3005
R20779 vdd.n1777 vdd.n1679 9.3005
R20780 vdd.n1779 vdd.n1778 9.3005
R20781 vdd.n1780 vdd.n1674 9.3005
R20782 vdd.n1782 vdd.n1781 9.3005
R20783 vdd.n1783 vdd.n1673 9.3005
R20784 vdd.n1785 vdd.n1784 9.3005
R20785 vdd.n1786 vdd.n1668 9.3005
R20786 vdd.n1788 vdd.n1787 9.3005
R20787 vdd.n1789 vdd.n1667 9.3005
R20788 vdd.n1791 vdd.n1790 9.3005
R20789 vdd.n1792 vdd.n1664 9.3005
R20790 vdd.n1798 vdd.n1797 9.3005
R20791 vdd.n1799 vdd.n1663 9.3005
R20792 vdd.n1801 vdd.n1800 9.3005
R20793 vdd.n1802 vdd.n1658 9.3005
R20794 vdd.n1804 vdd.n1803 9.3005
R20795 vdd.n1805 vdd.n1657 9.3005
R20796 vdd.n1807 vdd.n1806 9.3005
R20797 vdd.n1808 vdd.n1652 9.3005
R20798 vdd.n1810 vdd.n1809 9.3005
R20799 vdd.n1811 vdd.n1651 9.3005
R20800 vdd.n1813 vdd.n1812 9.3005
R20801 vdd.n1814 vdd.n1646 9.3005
R20802 vdd.n1816 vdd.n1815 9.3005
R20803 vdd.n1817 vdd.n1645 9.3005
R20804 vdd.n1819 vdd.n1818 9.3005
R20805 vdd.n1820 vdd.n1641 9.3005
R20806 vdd.n1822 vdd.n1821 9.3005
R20807 vdd.n1823 vdd.n1640 9.3005
R20808 vdd.n1825 vdd.n1824 9.3005
R20809 vdd.n1826 vdd.n1639 9.3005
R20810 vdd.n1832 vdd.n1831 9.3005
R20811 vdd.n1840 vdd.n1839 9.3005
R20812 vdd.n1841 vdd.n1595 9.3005
R20813 vdd.n1843 vdd.n1842 9.3005
R20814 vdd.n1585 vdd.n1584 9.3005
R20815 vdd.n1857 vdd.n1856 9.3005
R20816 vdd.n1858 vdd.n1583 9.3005
R20817 vdd.n1860 vdd.n1859 9.3005
R20818 vdd.n1574 vdd.n1573 9.3005
R20819 vdd.n1874 vdd.n1873 9.3005
R20820 vdd.n1875 vdd.n1572 9.3005
R20821 vdd.n1877 vdd.n1876 9.3005
R20822 vdd.n1563 vdd.n1562 9.3005
R20823 vdd.n1890 vdd.n1889 9.3005
R20824 vdd.n1891 vdd.n1561 9.3005
R20825 vdd.n1893 vdd.n1892 9.3005
R20826 vdd.n1551 vdd.n1550 9.3005
R20827 vdd.n1907 vdd.n1906 9.3005
R20828 vdd.n1597 vdd.n1596 9.3005
R20829 vdd.n2119 vdd.n2118 9.3005
R20830 vdd.n2114 vdd.n2113 9.3005
R20831 vdd.n2125 vdd.n2124 9.3005
R20832 vdd.n2127 vdd.n2126 9.3005
R20833 vdd.n2110 vdd.n2109 9.3005
R20834 vdd.n2133 vdd.n2132 9.3005
R20835 vdd.n2135 vdd.n2134 9.3005
R20836 vdd.n2107 vdd.n2104 9.3005
R20837 vdd.n2142 vdd.n2141 9.3005
R20838 vdd.n2174 vdd.n2173 9.3005
R20839 vdd.n2169 vdd.n2168 9.3005
R20840 vdd.n2180 vdd.n2179 9.3005
R20841 vdd.n2182 vdd.n2181 9.3005
R20842 vdd.n2165 vdd.n2164 9.3005
R20843 vdd.n2188 vdd.n2187 9.3005
R20844 vdd.n2190 vdd.n2189 9.3005
R20845 vdd.n2162 vdd.n2159 9.3005
R20846 vdd.n2197 vdd.n2196 9.3005
R20847 vdd.n2021 vdd.n2020 9.3005
R20848 vdd.n2016 vdd.n2015 9.3005
R20849 vdd.n2027 vdd.n2026 9.3005
R20850 vdd.n2029 vdd.n2028 9.3005
R20851 vdd.n2012 vdd.n2011 9.3005
R20852 vdd.n2035 vdd.n2034 9.3005
R20853 vdd.n2037 vdd.n2036 9.3005
R20854 vdd.n2009 vdd.n2006 9.3005
R20855 vdd.n2044 vdd.n2043 9.3005
R20856 vdd.n2076 vdd.n2075 9.3005
R20857 vdd.n2071 vdd.n2070 9.3005
R20858 vdd.n2082 vdd.n2081 9.3005
R20859 vdd.n2084 vdd.n2083 9.3005
R20860 vdd.n2067 vdd.n2066 9.3005
R20861 vdd.n2090 vdd.n2089 9.3005
R20862 vdd.n2092 vdd.n2091 9.3005
R20863 vdd.n2064 vdd.n2061 9.3005
R20864 vdd.n2099 vdd.n2098 9.3005
R20865 vdd.n1924 vdd.n1923 9.3005
R20866 vdd.n1919 vdd.n1918 9.3005
R20867 vdd.n1930 vdd.n1929 9.3005
R20868 vdd.n1932 vdd.n1931 9.3005
R20869 vdd.n1915 vdd.n1914 9.3005
R20870 vdd.n1938 vdd.n1937 9.3005
R20871 vdd.n1940 vdd.n1939 9.3005
R20872 vdd.n1912 vdd.n1909 9.3005
R20873 vdd.n1947 vdd.n1946 9.3005
R20874 vdd.n1979 vdd.n1978 9.3005
R20875 vdd.n1974 vdd.n1973 9.3005
R20876 vdd.n1985 vdd.n1984 9.3005
R20877 vdd.n1987 vdd.n1986 9.3005
R20878 vdd.n1970 vdd.n1969 9.3005
R20879 vdd.n1993 vdd.n1992 9.3005
R20880 vdd.n1995 vdd.n1994 9.3005
R20881 vdd.n1967 vdd.n1964 9.3005
R20882 vdd.n2002 vdd.n2001 9.3005
R20883 vdd.n1853 vdd.t101 9.18308
R20884 vdd.n3508 vdd.t176 9.18308
R20885 vdd.n1879 vdd.t72 8.95635
R20886 vdd.t82 vdd.n3549 8.95635
R20887 vdd.n300 vdd.n299 8.92171
R20888 vdd.n245 vdd.n244 8.92171
R20889 vdd.n202 vdd.n201 8.92171
R20890 vdd.n147 vdd.n146 8.92171
R20891 vdd.n105 vdd.n104 8.92171
R20892 vdd.n50 vdd.n49 8.92171
R20893 vdd.n2124 vdd.n2123 8.92171
R20894 vdd.n2179 vdd.n2178 8.92171
R20895 vdd.n2026 vdd.n2025 8.92171
R20896 vdd.n2081 vdd.n2080 8.92171
R20897 vdd.n1929 vdd.n1928 8.92171
R20898 vdd.n1984 vdd.n1983 8.92171
R20899 vdd.n223 vdd.n125 8.81535
R20900 vdd.n2102 vdd.n2004 8.81535
R20901 vdd.n1559 vdd.t109 8.72962
R20902 vdd.t76 vdd.n3558 8.72962
R20903 vdd.n2215 vdd.t97 8.50289
R20904 vdd.n3477 vdd.t70 8.50289
R20905 vdd.n28 vdd.n14 8.42249
R20906 vdd.n2231 vdd.t140 8.27616
R20907 vdd.t84 vdd.n636 8.27616
R20908 vdd.n3564 vdd.n3563 8.16225
R20909 vdd.n2202 vdd.n2201 8.16225
R20910 vdd.n296 vdd.n290 8.14595
R20911 vdd.n241 vdd.n235 8.14595
R20912 vdd.n198 vdd.n192 8.14595
R20913 vdd.n143 vdd.n137 8.14595
R20914 vdd.n101 vdd.n95 8.14595
R20915 vdd.n46 vdd.n40 8.14595
R20916 vdd.n2120 vdd.n2114 8.14595
R20917 vdd.n2175 vdd.n2169 8.14595
R20918 vdd.n2022 vdd.n2016 8.14595
R20919 vdd.n2077 vdd.n2071 8.14595
R20920 vdd.n1925 vdd.n1919 8.14595
R20921 vdd.n1980 vdd.n1974 8.14595
R20922 vdd.t239 vdd.n1593 7.8227
R20923 vdd.t212 vdd.n363 7.8227
R20924 vdd.n2430 vdd.n1105 7.70933
R20925 vdd.n2430 vdd.n1108 7.70933
R20926 vdd.n2436 vdd.n1094 7.70933
R20927 vdd.n2442 vdd.n1094 7.70933
R20928 vdd.n2442 vdd.n1087 7.70933
R20929 vdd.n2448 vdd.n1087 7.70933
R20930 vdd.n2448 vdd.n1090 7.70933
R20931 vdd.n2454 vdd.n1083 7.70933
R20932 vdd.n2460 vdd.n1077 7.70933
R20933 vdd.n2466 vdd.n1064 7.70933
R20934 vdd.n2472 vdd.n1064 7.70933
R20935 vdd.n2478 vdd.n1058 7.70933
R20936 vdd.n2484 vdd.n1051 7.70933
R20937 vdd.n2484 vdd.n1054 7.70933
R20938 vdd.n2490 vdd.n1047 7.70933
R20939 vdd.n2497 vdd.n1033 7.70933
R20940 vdd.n2503 vdd.n1033 7.70933
R20941 vdd.n2509 vdd.n1027 7.70933
R20942 vdd.n2515 vdd.n1023 7.70933
R20943 vdd.n2521 vdd.n1017 7.70933
R20944 vdd.n2539 vdd.n999 7.70933
R20945 vdd.n2539 vdd.n992 7.70933
R20946 vdd.n2547 vdd.n992 7.70933
R20947 vdd.n2629 vdd.n976 7.70933
R20948 vdd.n3012 vdd.n928 7.70933
R20949 vdd.n3024 vdd.n917 7.70933
R20950 vdd.n3024 vdd.n911 7.70933
R20951 vdd.n3030 vdd.n911 7.70933
R20952 vdd.n3042 vdd.n902 7.70933
R20953 vdd.n3048 vdd.n896 7.70933
R20954 vdd.n3060 vdd.n883 7.70933
R20955 vdd.n3067 vdd.n876 7.70933
R20956 vdd.n3067 vdd.n879 7.70933
R20957 vdd.n3073 vdd.n872 7.70933
R20958 vdd.n3079 vdd.n858 7.70933
R20959 vdd.n3085 vdd.n858 7.70933
R20960 vdd.n3091 vdd.n852 7.70933
R20961 vdd.n3097 vdd.n845 7.70933
R20962 vdd.n3097 vdd.n848 7.70933
R20963 vdd.n3103 vdd.n841 7.70933
R20964 vdd.n3109 vdd.n835 7.70933
R20965 vdd.n3115 vdd.n822 7.70933
R20966 vdd.n3121 vdd.n822 7.70933
R20967 vdd.n3121 vdd.n814 7.70933
R20968 vdd.n3172 vdd.n814 7.70933
R20969 vdd.n3172 vdd.n817 7.70933
R20970 vdd.n3178 vdd.n774 7.70933
R20971 vdd.n3248 vdd.n774 7.70933
R20972 vdd.n295 vdd.n292 7.3702
R20973 vdd.n240 vdd.n237 7.3702
R20974 vdd.n197 vdd.n194 7.3702
R20975 vdd.n142 vdd.n139 7.3702
R20976 vdd.n100 vdd.n97 7.3702
R20977 vdd.n45 vdd.n42 7.3702
R20978 vdd.n2119 vdd.n2116 7.3702
R20979 vdd.n2174 vdd.n2171 7.3702
R20980 vdd.n2021 vdd.n2018 7.3702
R20981 vdd.n2076 vdd.n2073 7.3702
R20982 vdd.n1924 vdd.n1921 7.3702
R20983 vdd.n1979 vdd.n1976 7.3702
R20984 vdd.n1077 vdd.t55 7.36923
R20985 vdd.n3103 vdd.t32 7.36923
R20986 vdd.n2454 vdd.t7 7.1425
R20987 vdd.n1396 vdd.t3 7.1425
R20988 vdd.n3036 vdd.t6 7.1425
R20989 vdd.n835 vdd.t16 7.1425
R20990 vdd.n1762 vdd.n1761 6.98232
R20991 vdd.n2318 vdd.n2317 6.98232
R20992 vdd.n547 vdd.n546 6.98232
R20993 vdd.n3332 vdd.n3331 6.98232
R20994 vdd.n2249 vdd.t136 6.91577
R20995 vdd.n3441 vdd.t106 6.91577
R20996 vdd.n1396 vdd.t4 6.80241
R20997 vdd.n3036 vdd.t48 6.80241
R20998 vdd.t94 vdd.n1530 6.68904
R20999 vdd.n3457 vdd.t154 6.68904
R21000 vdd.n2207 vdd.t74 6.46231
R21001 vdd.n2478 vdd.t14 6.46231
R21002 vdd.t19 vdd.n1027 6.46231
R21003 vdd.n3060 vdd.t24 6.46231
R21004 vdd.t40 vdd.n852 6.46231
R21005 vdd.n3485 vdd.t116 6.46231
R21006 vdd.n2554 vdd.t52 6.34895
R21007 vdd.n2933 vdd.t37 6.34895
R21008 vdd.n3564 vdd.n321 6.32949
R21009 vdd.n2201 vdd.n2200 6.32949
R21010 vdd.n3075 vdd.n868 6.2444
R21011 vdd.n2494 vdd.n2493 6.2444
R21012 vdd.t64 vdd.n1558 6.23558
R21013 vdd.t158 vdd.n332 6.23558
R21014 vdd.n1871 vdd.t124 6.00885
R21015 vdd.n3543 vdd.t122 6.00885
R21016 vdd.n2515 vdd.t45 5.89549
R21017 vdd.n896 vdd.t20 5.89549
R21018 vdd.n296 vdd.n295 5.81868
R21019 vdd.n241 vdd.n240 5.81868
R21020 vdd.n198 vdd.n197 5.81868
R21021 vdd.n143 vdd.n142 5.81868
R21022 vdd.n101 vdd.n100 5.81868
R21023 vdd.n46 vdd.n45 5.81868
R21024 vdd.n2120 vdd.n2119 5.81868
R21025 vdd.n2175 vdd.n2174 5.81868
R21026 vdd.n2022 vdd.n2021 5.81868
R21027 vdd.n2077 vdd.n2076 5.81868
R21028 vdd.n1925 vdd.n1924 5.81868
R21029 vdd.n1980 vdd.n1979 5.81868
R21030 vdd.n2637 vdd.n2636 5.77611
R21031 vdd.n1320 vdd.n1319 5.77611
R21032 vdd.n2945 vdd.n2944 5.77611
R21033 vdd.n3187 vdd.n806 5.77611
R21034 vdd.n3253 vdd.n770 5.77611
R21035 vdd.n2808 vdd.n2742 5.77611
R21036 vdd.n2562 vdd.n983 5.77611
R21037 vdd.n1456 vdd.n1288 5.77611
R21038 vdd.n1831 vdd.n1605 5.62474
R21039 vdd.n2281 vdd.n2278 5.62474
R21040 vdd.n3522 vdd.n407 5.62474
R21041 vdd.n3287 vdd.n3284 5.62474
R21042 vdd.n2490 vdd.t34 5.55539
R21043 vdd.n872 vdd.t10 5.55539
R21044 vdd.n1581 vdd.t124 5.32866
R21045 vdd.t122 vdd.n3542 5.32866
R21046 vdd.n1887 vdd.t64 5.10193
R21047 vdd.n3551 vdd.t158 5.10193
R21048 vdd.n299 vdd.n290 5.04292
R21049 vdd.n244 vdd.n235 5.04292
R21050 vdd.n201 vdd.n192 5.04292
R21051 vdd.n146 vdd.n137 5.04292
R21052 vdd.n104 vdd.n95 5.04292
R21053 vdd.n49 vdd.n40 5.04292
R21054 vdd.n2123 vdd.n2114 5.04292
R21055 vdd.n2178 vdd.n2169 5.04292
R21056 vdd.n2025 vdd.n2016 5.04292
R21057 vdd.n2080 vdd.n2071 5.04292
R21058 vdd.n1928 vdd.n1919 5.04292
R21059 vdd.n1983 vdd.n1974 5.04292
R21060 vdd.n1903 vdd.t74 4.8752
R21061 vdd.t13 vdd.t25 4.8752
R21062 vdd.t56 vdd.t2 4.8752
R21063 vdd.t116 vdd.n328 4.8752
R21064 vdd.n2638 vdd.n2637 4.83952
R21065 vdd.n1319 vdd.n1318 4.83952
R21066 vdd.n2946 vdd.n2945 4.83952
R21067 vdd.n806 vdd.n801 4.83952
R21068 vdd.n770 vdd.n765 4.83952
R21069 vdd.n2805 vdd.n2742 4.83952
R21070 vdd.n2565 vdd.n983 4.83952
R21071 vdd.n1459 vdd.n1288 4.83952
R21072 vdd.n1370 vdd.t22 4.76184
R21073 vdd.n3018 vdd.t8 4.76184
R21074 vdd.n2286 vdd.n2285 4.74817
R21075 vdd.n1492 vdd.n1487 4.74817
R21076 vdd.n1154 vdd.n1151 4.74817
R21077 vdd.n2379 vdd.n1150 4.74817
R21078 vdd.n2384 vdd.n1151 4.74817
R21079 vdd.n2383 vdd.n1150 4.74817
R21080 vdd.n664 vdd.n662 4.74817
R21081 vdd.n3402 vdd.n665 4.74817
R21082 vdd.n3405 vdd.n665 4.74817
R21083 vdd.n3406 vdd.n664 4.74817
R21084 vdd.n3294 vdd.n749 4.74817
R21085 vdd.n3290 vdd.n751 4.74817
R21086 vdd.n3293 vdd.n751 4.74817
R21087 vdd.n3298 vdd.n749 4.74817
R21088 vdd.n2285 vdd.n1250 4.74817
R21089 vdd.n1489 vdd.n1487 4.74817
R21090 vdd.n321 vdd.n320 4.7074
R21091 vdd.n223 vdd.n222 4.7074
R21092 vdd.n2200 vdd.n2199 4.7074
R21093 vdd.n2102 vdd.n2101 4.7074
R21094 vdd.n2223 vdd.t94 4.64847
R21095 vdd.t15 vdd.n1058 4.64847
R21096 vdd.n2509 vdd.t54 4.64847
R21097 vdd.t43 vdd.n883 4.64847
R21098 vdd.n3091 vdd.t39 4.64847
R21099 vdd.n3466 vdd.t154 4.64847
R21100 vdd.n1047 vdd.t257 4.53511
R21101 vdd.n3073 vdd.t220 4.53511
R21102 vdd.n1524 vdd.t136 4.42174
R21103 vdd.n2436 vdd.t198 4.42174
R21104 vdd.n1370 vdd.t243 4.42174
R21105 vdd.n3018 vdd.t250 4.42174
R21106 vdd.n817 vdd.t194 4.42174
R21107 vdd.t106 vdd.n635 4.42174
R21108 vdd.n3064 vdd.n868 4.37123
R21109 vdd.n2495 vdd.n2494 4.37123
R21110 vdd.n2533 vdd.t41 4.30838
R21111 vdd.n2921 vdd.t28 4.30838
R21112 vdd.n300 vdd.n288 4.26717
R21113 vdd.n245 vdd.n233 4.26717
R21114 vdd.n202 vdd.n190 4.26717
R21115 vdd.n147 vdd.n135 4.26717
R21116 vdd.n105 vdd.n93 4.26717
R21117 vdd.n50 vdd.n38 4.26717
R21118 vdd.n2124 vdd.n2112 4.26717
R21119 vdd.n2179 vdd.n2167 4.26717
R21120 vdd.n2026 vdd.n2014 4.26717
R21121 vdd.n2081 vdd.n2069 4.26717
R21122 vdd.n1929 vdd.n1917 4.26717
R21123 vdd.n1984 vdd.n1972 4.26717
R21124 vdd.n321 vdd.n223 4.10845
R21125 vdd.n2200 vdd.n2102 4.10845
R21126 vdd.n277 vdd.t151 4.06363
R21127 vdd.n277 vdd.t184 4.06363
R21128 vdd.n275 vdd.t83 4.06363
R21129 vdd.n275 vdd.t119 4.06363
R21130 vdd.n273 vdd.t121 4.06363
R21131 vdd.n273 vdd.t166 4.06363
R21132 vdd.n271 vdd.t168 4.06363
R21133 vdd.n271 vdd.t77 4.06363
R21134 vdd.n269 vdd.t96 4.06363
R21135 vdd.n269 vdd.t146 4.06363
R21136 vdd.n267 vdd.t169 4.06363
R21137 vdd.n267 vdd.t182 4.06363
R21138 vdd.n265 vdd.t186 4.06363
R21139 vdd.n265 vdd.t103 4.06363
R21140 vdd.n179 vdd.t144 4.06363
R21141 vdd.n179 vdd.t177 4.06363
R21142 vdd.n177 vdd.t190 4.06363
R21143 vdd.n177 vdd.t105 4.06363
R21144 vdd.n175 vdd.t113 4.06363
R21145 vdd.n175 vdd.t159 4.06363
R21146 vdd.n173 vdd.t160 4.06363
R21147 vdd.n173 vdd.t183 4.06363
R21148 vdd.n171 vdd.t71 4.06363
R21149 vdd.n171 vdd.t128 4.06363
R21150 vdd.n169 vdd.t163 4.06363
R21151 vdd.n169 vdd.t170 4.06363
R21152 vdd.n167 vdd.t178 4.06363
R21153 vdd.n167 vdd.t85 4.06363
R21154 vdd.n82 vdd.t123 4.06363
R21155 vdd.n82 vdd.t187 4.06363
R21156 vdd.n80 vdd.t108 4.06363
R21157 vdd.n80 vdd.t173 4.06363
R21158 vdd.n78 vdd.t133 4.06363
R21159 vdd.n78 vdd.t161 4.06363
R21160 vdd.n76 vdd.t117 4.06363
R21161 vdd.n76 vdd.t180 4.06363
R21162 vdd.n74 vdd.t93 4.06363
R21163 vdd.n74 vdd.t167 4.06363
R21164 vdd.n72 vdd.t88 4.06363
R21165 vdd.n72 vdd.t155 4.06363
R21166 vdd.n70 vdd.t107 4.06363
R21167 vdd.n70 vdd.t171 4.06363
R21168 vdd.n2144 vdd.t150 4.06363
R21169 vdd.n2144 vdd.t149 4.06363
R21170 vdd.n2146 vdd.t114 4.06363
R21171 vdd.n2146 vdd.t92 4.06363
R21172 vdd.n2148 vdd.t90 4.06363
R21173 vdd.n2148 vdd.t143 4.06363
R21174 vdd.n2150 vdd.t126 4.06363
R21175 vdd.n2150 vdd.t91 4.06363
R21176 vdd.n2152 vdd.t86 4.06363
R21177 vdd.n2152 vdd.t165 4.06363
R21178 vdd.n2154 vdd.t164 4.06363
R21179 vdd.n2154 vdd.t120 4.06363
R21180 vdd.n2156 vdd.t115 4.06363
R21181 vdd.n2156 vdd.t189 4.06363
R21182 vdd.n2046 vdd.t141 4.06363
R21183 vdd.n2046 vdd.t137 4.06363
R21184 vdd.n2048 vdd.t95 4.06363
R21185 vdd.n2048 vdd.t79 4.06363
R21186 vdd.n2050 vdd.t67 4.06363
R21187 vdd.n2050 vdd.t132 4.06363
R21188 vdd.n2052 vdd.t110 4.06363
R21189 vdd.n2052 vdd.t75 4.06363
R21190 vdd.n2054 vdd.t65 4.06363
R21191 vdd.n2054 vdd.t157 4.06363
R21192 vdd.n2056 vdd.t153 4.06363
R21193 vdd.n2056 vdd.t111 4.06363
R21194 vdd.n2058 vdd.t102 4.06363
R21195 vdd.n2058 vdd.t179 4.06363
R21196 vdd.n1949 vdd.t172 4.06363
R21197 vdd.n1949 vdd.t191 4.06363
R21198 vdd.n1951 vdd.t156 4.06363
R21199 vdd.n1951 vdd.t89 4.06363
R21200 vdd.n1953 vdd.t142 4.06363
R21201 vdd.n1953 vdd.t98 4.06363
R21202 vdd.n1955 vdd.t181 4.06363
R21203 vdd.n1955 vdd.t118 4.06363
R21204 vdd.n1957 vdd.t162 4.06363
R21205 vdd.n1957 vdd.t135 4.06363
R21206 vdd.n1959 vdd.t174 4.06363
R21207 vdd.n1959 vdd.t73 4.06363
R21208 vdd.n1961 vdd.t188 4.06363
R21209 vdd.n1961 vdd.t125 4.06363
R21210 vdd.n1083 vdd.t47 3.96828
R21211 vdd.n2527 vdd.t27 3.96828
R21212 vdd.n2915 vdd.t44 3.96828
R21213 vdd.n3109 vdd.t33 3.96828
R21214 vdd.n26 vdd.t275 3.9605
R21215 vdd.n26 vdd.t192 3.9605
R21216 vdd.n23 vdd.t61 3.9605
R21217 vdd.n23 vdd.t274 3.9605
R21218 vdd.n21 vdd.t273 3.9605
R21219 vdd.n21 vdd.t59 3.9605
R21220 vdd.n20 vdd.t63 3.9605
R21221 vdd.n20 vdd.t270 3.9605
R21222 vdd.n15 vdd.t271 3.9605
R21223 vdd.n15 vdd.t272 3.9605
R21224 vdd.n16 vdd.t62 3.9605
R21225 vdd.n16 vdd.t269 3.9605
R21226 vdd.n18 vdd.t0 3.9605
R21227 vdd.n18 vdd.t60 3.9605
R21228 vdd.n25 vdd.t1 3.9605
R21229 vdd.n25 vdd.t58 3.9605
R21230 vdd.n2460 vdd.t47 3.74155
R21231 vdd.n1017 vdd.t27 3.74155
R21232 vdd.n3042 vdd.t44 3.74155
R21233 vdd.n841 vdd.t33 3.74155
R21234 vdd.n7 vdd.t57 3.61217
R21235 vdd.n7 vdd.t21 3.61217
R21236 vdd.n8 vdd.t29 3.61217
R21237 vdd.n8 vdd.t49 3.61217
R21238 vdd.n10 vdd.t38 3.61217
R21239 vdd.n10 vdd.t9 3.61217
R21240 vdd.n12 vdd.t18 3.61217
R21241 vdd.n12 vdd.t36 3.61217
R21242 vdd.n5 vdd.t51 3.61217
R21243 vdd.n5 vdd.t31 3.61217
R21244 vdd.n3 vdd.t23 3.61217
R21245 vdd.n3 vdd.t53 3.61217
R21246 vdd.n1 vdd.t5 3.61217
R21247 vdd.n1 vdd.t42 3.61217
R21248 vdd.n0 vdd.t46 3.61217
R21249 vdd.n0 vdd.t26 3.61217
R21250 vdd.n1837 vdd.t239 3.51482
R21251 vdd.n3527 vdd.t212 3.51482
R21252 vdd.n304 vdd.n303 3.49141
R21253 vdd.n249 vdd.n248 3.49141
R21254 vdd.n206 vdd.n205 3.49141
R21255 vdd.n151 vdd.n150 3.49141
R21256 vdd.n109 vdd.n108 3.49141
R21257 vdd.n54 vdd.n53 3.49141
R21258 vdd.n2128 vdd.n2127 3.49141
R21259 vdd.n2183 vdd.n2182 3.49141
R21260 vdd.n2030 vdd.n2029 3.49141
R21261 vdd.n2085 vdd.n2084 3.49141
R21262 vdd.n1933 vdd.n1932 3.49141
R21263 vdd.n1988 vdd.n1987 3.49141
R21264 vdd.t41 vdd.n999 3.40145
R21265 vdd.n2701 vdd.t50 3.40145
R21266 vdd.n3005 vdd.t35 3.40145
R21267 vdd.n3030 vdd.t28 3.40145
R21268 vdd.n1108 vdd.t198 3.28809
R21269 vdd.n2554 vdd.t243 3.28809
R21270 vdd.n2933 vdd.t250 3.28809
R21271 vdd.n3178 vdd.t194 3.28809
R21272 vdd.n2240 vdd.t140 3.06136
R21273 vdd.n2472 vdd.t15 3.06136
R21274 vdd.n1408 vdd.t54 3.06136
R21275 vdd.n3054 vdd.t43 3.06136
R21276 vdd.t39 vdd.n845 3.06136
R21277 vdd.n3449 vdd.t84 3.06136
R21278 vdd.n2547 vdd.t22 2.94799
R21279 vdd.t8 vdd.n917 2.94799
R21280 vdd.t97 vdd.n1536 2.83463
R21281 vdd.n624 vdd.t70 2.83463
R21282 vdd.n307 vdd.n286 2.71565
R21283 vdd.n252 vdd.n231 2.71565
R21284 vdd.n209 vdd.n188 2.71565
R21285 vdd.n154 vdd.n133 2.71565
R21286 vdd.n112 vdd.n91 2.71565
R21287 vdd.n57 vdd.n36 2.71565
R21288 vdd.n2131 vdd.n2110 2.71565
R21289 vdd.n2186 vdd.n2165 2.71565
R21290 vdd.n2033 vdd.n2012 2.71565
R21291 vdd.n2088 vdd.n2067 2.71565
R21292 vdd.n1936 vdd.n1915 2.71565
R21293 vdd.n1991 vdd.n1970 2.71565
R21294 vdd.n1904 vdd.t109 2.6079
R21295 vdd.n3559 vdd.t76 2.6079
R21296 vdd.n2521 vdd.t25 2.49453
R21297 vdd.n902 vdd.t56 2.49453
R21298 vdd.n294 vdd.n293 2.4129
R21299 vdd.n239 vdd.n238 2.4129
R21300 vdd.n196 vdd.n195 2.4129
R21301 vdd.n141 vdd.n140 2.4129
R21302 vdd.n99 vdd.n98 2.4129
R21303 vdd.n44 vdd.n43 2.4129
R21304 vdd.n2118 vdd.n2117 2.4129
R21305 vdd.n2173 vdd.n2172 2.4129
R21306 vdd.n2020 vdd.n2019 2.4129
R21307 vdd.n2075 vdd.n2074 2.4129
R21308 vdd.n1923 vdd.n1922 2.4129
R21309 vdd.n1978 vdd.n1977 2.4129
R21310 vdd.t72 vdd.n1565 2.38117
R21311 vdd.n3550 vdd.t82 2.38117
R21312 vdd.n2391 vdd.n1151 2.27742
R21313 vdd.n2391 vdd.n1150 2.27742
R21314 vdd.n3214 vdd.n665 2.27742
R21315 vdd.n3214 vdd.n664 2.27742
R21316 vdd.n3282 vdd.n751 2.27742
R21317 vdd.n3282 vdd.n749 2.27742
R21318 vdd.n2285 vdd.n2284 2.27742
R21319 vdd.n2284 vdd.n1487 2.27742
R21320 vdd.n1862 vdd.t101 2.15444
R21321 vdd.n1054 vdd.t34 2.15444
R21322 vdd.n2497 vdd.t12 2.15444
R21323 vdd.n879 vdd.t11 2.15444
R21324 vdd.n3079 vdd.t10 2.15444
R21325 vdd.n3541 vdd.t176 2.15444
R21326 vdd.n308 vdd.n284 1.93989
R21327 vdd.n253 vdd.n229 1.93989
R21328 vdd.n210 vdd.n186 1.93989
R21329 vdd.n155 vdd.n131 1.93989
R21330 vdd.n113 vdd.n89 1.93989
R21331 vdd.n58 vdd.n34 1.93989
R21332 vdd.n2132 vdd.n2108 1.93989
R21333 vdd.n2187 vdd.n2163 1.93989
R21334 vdd.n2034 vdd.n2010 1.93989
R21335 vdd.n2089 vdd.n2065 1.93989
R21336 vdd.n1937 vdd.n1913 1.93989
R21337 vdd.n1992 vdd.n1968 1.93989
R21338 vdd.n1408 vdd.t45 1.81434
R21339 vdd.n3054 vdd.t20 1.81434
R21340 vdd.n1854 vdd.t138 1.70098
R21341 vdd.n3535 vdd.t80 1.70098
R21342 vdd.n1870 vdd.t152 1.47425
R21343 vdd.n349 vdd.t104 1.47425
R21344 vdd.t52 vdd.n976 1.36088
R21345 vdd.n3012 vdd.t37 1.36088
R21346 vdd.n1895 vdd.t134 1.24752
R21347 vdd.t202 vdd.n1500 1.24752
R21348 vdd.t14 vdd.n1051 1.24752
R21349 vdd.n2503 vdd.t19 1.24752
R21350 vdd.t24 vdd.n876 1.24752
R21351 vdd.n3085 vdd.t40 1.24752
R21352 vdd.n659 vdd.t216 1.24752
R21353 vdd.t112 vdd.n3557 1.24752
R21354 vdd.n2201 vdd.n28 1.16438
R21355 vdd.n319 vdd.n279 1.16414
R21356 vdd.n312 vdd.n311 1.16414
R21357 vdd.n264 vdd.n224 1.16414
R21358 vdd.n257 vdd.n256 1.16414
R21359 vdd.n221 vdd.n181 1.16414
R21360 vdd.n214 vdd.n213 1.16414
R21361 vdd.n166 vdd.n126 1.16414
R21362 vdd.n159 vdd.n158 1.16414
R21363 vdd.n124 vdd.n84 1.16414
R21364 vdd.n117 vdd.n116 1.16414
R21365 vdd.n69 vdd.n29 1.16414
R21366 vdd.n62 vdd.n61 1.16414
R21367 vdd.n2143 vdd.n2103 1.16414
R21368 vdd.n2136 vdd.n2135 1.16414
R21369 vdd.n2198 vdd.n2158 1.16414
R21370 vdd.n2191 vdd.n2190 1.16414
R21371 vdd.n2045 vdd.n2005 1.16414
R21372 vdd.n2038 vdd.n2037 1.16414
R21373 vdd.n2100 vdd.n2060 1.16414
R21374 vdd.n2093 vdd.n2092 1.16414
R21375 vdd.n1948 vdd.n1908 1.16414
R21376 vdd.n1941 vdd.n1940 1.16414
R21377 vdd.n2003 vdd.n1963 1.16414
R21378 vdd.n1996 vdd.n1995 1.16414
R21379 vdd vdd.n3564 1.15654
R21380 vdd.n1547 vdd.t66 1.02079
R21381 vdd.t257 vdd.t12 1.02079
R21382 vdd.t11 vdd.t220 1.02079
R21383 vdd.t127 vdd.n613 1.02079
R21384 vdd.n1726 vdd.n1605 0.970197
R21385 vdd.n2282 vdd.n2281 0.970197
R21386 vdd.n599 vdd.n407 0.970197
R21387 vdd.n3289 vdd.n3287 0.970197
R21388 vdd.n2527 vdd.t4 0.907421
R21389 vdd.n2915 vdd.t48 0.907421
R21390 vdd.n2232 vdd.t78 0.794056
R21391 vdd.n3458 vdd.t87 0.794056
R21392 vdd.n2248 vdd.t68 0.567326
R21393 vdd.n1090 vdd.t7 0.567326
R21394 vdd.n2533 vdd.t3 0.567326
R21395 vdd.n2921 vdd.t6 0.567326
R21396 vdd.n3115 vdd.t16 0.567326
R21397 vdd.t129 vdd.n642 0.567326
R21398 vdd.n2272 vdd.n1152 0.482207
R21399 vdd.n3414 vdd.n3413 0.482207
R21400 vdd.n444 vdd.n443 0.482207
R21401 vdd.n3521 vdd.n3520 0.482207
R21402 vdd.n3420 vdd.n656 0.482207
R21403 vdd.n2262 vdd.n1488 0.482207
R21404 vdd.n1833 vdd.n1832 0.482207
R21405 vdd.n1639 vdd.n1596 0.482207
R21406 vdd.n4 vdd.n2 0.459552
R21407 vdd.n11 vdd.n9 0.459552
R21408 vdd.n317 vdd.n316 0.388379
R21409 vdd.n283 vdd.n281 0.388379
R21410 vdd.n262 vdd.n261 0.388379
R21411 vdd.n228 vdd.n226 0.388379
R21412 vdd.n219 vdd.n218 0.388379
R21413 vdd.n185 vdd.n183 0.388379
R21414 vdd.n164 vdd.n163 0.388379
R21415 vdd.n130 vdd.n128 0.388379
R21416 vdd.n122 vdd.n121 0.388379
R21417 vdd.n88 vdd.n86 0.388379
R21418 vdd.n67 vdd.n66 0.388379
R21419 vdd.n33 vdd.n31 0.388379
R21420 vdd.n2141 vdd.n2140 0.388379
R21421 vdd.n2107 vdd.n2105 0.388379
R21422 vdd.n2196 vdd.n2195 0.388379
R21423 vdd.n2162 vdd.n2160 0.388379
R21424 vdd.n2043 vdd.n2042 0.388379
R21425 vdd.n2009 vdd.n2007 0.388379
R21426 vdd.n2098 vdd.n2097 0.388379
R21427 vdd.n2064 vdd.n2062 0.388379
R21428 vdd.n1946 vdd.n1945 0.388379
R21429 vdd.n1912 vdd.n1910 0.388379
R21430 vdd.n2001 vdd.n2000 0.388379
R21431 vdd.n1967 vdd.n1965 0.388379
R21432 vdd.n19 vdd.n17 0.387128
R21433 vdd.n24 vdd.n22 0.387128
R21434 vdd.n6 vdd.n4 0.358259
R21435 vdd.n13 vdd.n11 0.358259
R21436 vdd.n268 vdd.n266 0.358259
R21437 vdd.n270 vdd.n268 0.358259
R21438 vdd.n272 vdd.n270 0.358259
R21439 vdd.n274 vdd.n272 0.358259
R21440 vdd.n276 vdd.n274 0.358259
R21441 vdd.n278 vdd.n276 0.358259
R21442 vdd.n320 vdd.n278 0.358259
R21443 vdd.n170 vdd.n168 0.358259
R21444 vdd.n172 vdd.n170 0.358259
R21445 vdd.n174 vdd.n172 0.358259
R21446 vdd.n176 vdd.n174 0.358259
R21447 vdd.n178 vdd.n176 0.358259
R21448 vdd.n180 vdd.n178 0.358259
R21449 vdd.n222 vdd.n180 0.358259
R21450 vdd.n73 vdd.n71 0.358259
R21451 vdd.n75 vdd.n73 0.358259
R21452 vdd.n77 vdd.n75 0.358259
R21453 vdd.n79 vdd.n77 0.358259
R21454 vdd.n81 vdd.n79 0.358259
R21455 vdd.n83 vdd.n81 0.358259
R21456 vdd.n125 vdd.n83 0.358259
R21457 vdd.n2199 vdd.n2157 0.358259
R21458 vdd.n2157 vdd.n2155 0.358259
R21459 vdd.n2155 vdd.n2153 0.358259
R21460 vdd.n2153 vdd.n2151 0.358259
R21461 vdd.n2151 vdd.n2149 0.358259
R21462 vdd.n2149 vdd.n2147 0.358259
R21463 vdd.n2147 vdd.n2145 0.358259
R21464 vdd.n2101 vdd.n2059 0.358259
R21465 vdd.n2059 vdd.n2057 0.358259
R21466 vdd.n2057 vdd.n2055 0.358259
R21467 vdd.n2055 vdd.n2053 0.358259
R21468 vdd.n2053 vdd.n2051 0.358259
R21469 vdd.n2051 vdd.n2049 0.358259
R21470 vdd.n2049 vdd.n2047 0.358259
R21471 vdd.n2004 vdd.n1962 0.358259
R21472 vdd.n1962 vdd.n1960 0.358259
R21473 vdd.n1960 vdd.n1958 0.358259
R21474 vdd.n1958 vdd.n1956 0.358259
R21475 vdd.n1956 vdd.n1954 0.358259
R21476 vdd.n1954 vdd.n1952 0.358259
R21477 vdd.n1952 vdd.n1950 0.358259
R21478 vdd.n2466 vdd.t55 0.340595
R21479 vdd.n1023 vdd.t13 0.340595
R21480 vdd.n3048 vdd.t2 0.340595
R21481 vdd.n848 vdd.t32 0.340595
R21482 vdd.n14 vdd.n6 0.334552
R21483 vdd.n14 vdd.n13 0.334552
R21484 vdd.n27 vdd.n19 0.21707
R21485 vdd.n27 vdd.n24 0.21707
R21486 vdd.n318 vdd.n280 0.155672
R21487 vdd.n310 vdd.n280 0.155672
R21488 vdd.n310 vdd.n309 0.155672
R21489 vdd.n309 vdd.n285 0.155672
R21490 vdd.n302 vdd.n285 0.155672
R21491 vdd.n302 vdd.n301 0.155672
R21492 vdd.n301 vdd.n289 0.155672
R21493 vdd.n294 vdd.n289 0.155672
R21494 vdd.n263 vdd.n225 0.155672
R21495 vdd.n255 vdd.n225 0.155672
R21496 vdd.n255 vdd.n254 0.155672
R21497 vdd.n254 vdd.n230 0.155672
R21498 vdd.n247 vdd.n230 0.155672
R21499 vdd.n247 vdd.n246 0.155672
R21500 vdd.n246 vdd.n234 0.155672
R21501 vdd.n239 vdd.n234 0.155672
R21502 vdd.n220 vdd.n182 0.155672
R21503 vdd.n212 vdd.n182 0.155672
R21504 vdd.n212 vdd.n211 0.155672
R21505 vdd.n211 vdd.n187 0.155672
R21506 vdd.n204 vdd.n187 0.155672
R21507 vdd.n204 vdd.n203 0.155672
R21508 vdd.n203 vdd.n191 0.155672
R21509 vdd.n196 vdd.n191 0.155672
R21510 vdd.n165 vdd.n127 0.155672
R21511 vdd.n157 vdd.n127 0.155672
R21512 vdd.n157 vdd.n156 0.155672
R21513 vdd.n156 vdd.n132 0.155672
R21514 vdd.n149 vdd.n132 0.155672
R21515 vdd.n149 vdd.n148 0.155672
R21516 vdd.n148 vdd.n136 0.155672
R21517 vdd.n141 vdd.n136 0.155672
R21518 vdd.n123 vdd.n85 0.155672
R21519 vdd.n115 vdd.n85 0.155672
R21520 vdd.n115 vdd.n114 0.155672
R21521 vdd.n114 vdd.n90 0.155672
R21522 vdd.n107 vdd.n90 0.155672
R21523 vdd.n107 vdd.n106 0.155672
R21524 vdd.n106 vdd.n94 0.155672
R21525 vdd.n99 vdd.n94 0.155672
R21526 vdd.n68 vdd.n30 0.155672
R21527 vdd.n60 vdd.n30 0.155672
R21528 vdd.n60 vdd.n59 0.155672
R21529 vdd.n59 vdd.n35 0.155672
R21530 vdd.n52 vdd.n35 0.155672
R21531 vdd.n52 vdd.n51 0.155672
R21532 vdd.n51 vdd.n39 0.155672
R21533 vdd.n44 vdd.n39 0.155672
R21534 vdd.n2142 vdd.n2104 0.155672
R21535 vdd.n2134 vdd.n2104 0.155672
R21536 vdd.n2134 vdd.n2133 0.155672
R21537 vdd.n2133 vdd.n2109 0.155672
R21538 vdd.n2126 vdd.n2109 0.155672
R21539 vdd.n2126 vdd.n2125 0.155672
R21540 vdd.n2125 vdd.n2113 0.155672
R21541 vdd.n2118 vdd.n2113 0.155672
R21542 vdd.n2197 vdd.n2159 0.155672
R21543 vdd.n2189 vdd.n2159 0.155672
R21544 vdd.n2189 vdd.n2188 0.155672
R21545 vdd.n2188 vdd.n2164 0.155672
R21546 vdd.n2181 vdd.n2164 0.155672
R21547 vdd.n2181 vdd.n2180 0.155672
R21548 vdd.n2180 vdd.n2168 0.155672
R21549 vdd.n2173 vdd.n2168 0.155672
R21550 vdd.n2044 vdd.n2006 0.155672
R21551 vdd.n2036 vdd.n2006 0.155672
R21552 vdd.n2036 vdd.n2035 0.155672
R21553 vdd.n2035 vdd.n2011 0.155672
R21554 vdd.n2028 vdd.n2011 0.155672
R21555 vdd.n2028 vdd.n2027 0.155672
R21556 vdd.n2027 vdd.n2015 0.155672
R21557 vdd.n2020 vdd.n2015 0.155672
R21558 vdd.n2099 vdd.n2061 0.155672
R21559 vdd.n2091 vdd.n2061 0.155672
R21560 vdd.n2091 vdd.n2090 0.155672
R21561 vdd.n2090 vdd.n2066 0.155672
R21562 vdd.n2083 vdd.n2066 0.155672
R21563 vdd.n2083 vdd.n2082 0.155672
R21564 vdd.n2082 vdd.n2070 0.155672
R21565 vdd.n2075 vdd.n2070 0.155672
R21566 vdd.n1947 vdd.n1909 0.155672
R21567 vdd.n1939 vdd.n1909 0.155672
R21568 vdd.n1939 vdd.n1938 0.155672
R21569 vdd.n1938 vdd.n1914 0.155672
R21570 vdd.n1931 vdd.n1914 0.155672
R21571 vdd.n1931 vdd.n1930 0.155672
R21572 vdd.n1930 vdd.n1918 0.155672
R21573 vdd.n1923 vdd.n1918 0.155672
R21574 vdd.n2002 vdd.n1964 0.155672
R21575 vdd.n1994 vdd.n1964 0.155672
R21576 vdd.n1994 vdd.n1993 0.155672
R21577 vdd.n1993 vdd.n1969 0.155672
R21578 vdd.n1986 vdd.n1969 0.155672
R21579 vdd.n1986 vdd.n1985 0.155672
R21580 vdd.n1985 vdd.n1973 0.155672
R21581 vdd.n1978 vdd.n1973 0.155672
R21582 vdd.n1157 vdd.n1149 0.152939
R21583 vdd.n1161 vdd.n1157 0.152939
R21584 vdd.n1162 vdd.n1161 0.152939
R21585 vdd.n1163 vdd.n1162 0.152939
R21586 vdd.n1164 vdd.n1163 0.152939
R21587 vdd.n1168 vdd.n1164 0.152939
R21588 vdd.n1169 vdd.n1168 0.152939
R21589 vdd.n1170 vdd.n1169 0.152939
R21590 vdd.n1171 vdd.n1170 0.152939
R21591 vdd.n1175 vdd.n1171 0.152939
R21592 vdd.n1176 vdd.n1175 0.152939
R21593 vdd.n1177 vdd.n1176 0.152939
R21594 vdd.n2355 vdd.n1177 0.152939
R21595 vdd.n2355 vdd.n2354 0.152939
R21596 vdd.n2354 vdd.n2353 0.152939
R21597 vdd.n2353 vdd.n1183 0.152939
R21598 vdd.n1188 vdd.n1183 0.152939
R21599 vdd.n1189 vdd.n1188 0.152939
R21600 vdd.n1190 vdd.n1189 0.152939
R21601 vdd.n1194 vdd.n1190 0.152939
R21602 vdd.n1195 vdd.n1194 0.152939
R21603 vdd.n1196 vdd.n1195 0.152939
R21604 vdd.n1197 vdd.n1196 0.152939
R21605 vdd.n1201 vdd.n1197 0.152939
R21606 vdd.n1202 vdd.n1201 0.152939
R21607 vdd.n1203 vdd.n1202 0.152939
R21608 vdd.n1204 vdd.n1203 0.152939
R21609 vdd.n1208 vdd.n1204 0.152939
R21610 vdd.n1209 vdd.n1208 0.152939
R21611 vdd.n1210 vdd.n1209 0.152939
R21612 vdd.n1211 vdd.n1210 0.152939
R21613 vdd.n1215 vdd.n1211 0.152939
R21614 vdd.n1216 vdd.n1215 0.152939
R21615 vdd.n1217 vdd.n1216 0.152939
R21616 vdd.n2316 vdd.n1217 0.152939
R21617 vdd.n2316 vdd.n2315 0.152939
R21618 vdd.n2315 vdd.n2314 0.152939
R21619 vdd.n2314 vdd.n1223 0.152939
R21620 vdd.n1228 vdd.n1223 0.152939
R21621 vdd.n1229 vdd.n1228 0.152939
R21622 vdd.n1230 vdd.n1229 0.152939
R21623 vdd.n1234 vdd.n1230 0.152939
R21624 vdd.n1235 vdd.n1234 0.152939
R21625 vdd.n1236 vdd.n1235 0.152939
R21626 vdd.n1237 vdd.n1236 0.152939
R21627 vdd.n1241 vdd.n1237 0.152939
R21628 vdd.n1242 vdd.n1241 0.152939
R21629 vdd.n1243 vdd.n1242 0.152939
R21630 vdd.n1244 vdd.n1243 0.152939
R21631 vdd.n1248 vdd.n1244 0.152939
R21632 vdd.n1249 vdd.n1248 0.152939
R21633 vdd.n2390 vdd.n1152 0.152939
R21634 vdd.n2204 vdd.n2203 0.152939
R21635 vdd.n2204 vdd.n1539 0.152939
R21636 vdd.n2218 vdd.n1539 0.152939
R21637 vdd.n2219 vdd.n2218 0.152939
R21638 vdd.n2220 vdd.n2219 0.152939
R21639 vdd.n2220 vdd.n1527 0.152939
R21640 vdd.n2235 vdd.n1527 0.152939
R21641 vdd.n2236 vdd.n2235 0.152939
R21642 vdd.n2237 vdd.n2236 0.152939
R21643 vdd.n2237 vdd.n1516 0.152939
R21644 vdd.n2252 vdd.n1516 0.152939
R21645 vdd.n2253 vdd.n2252 0.152939
R21646 vdd.n2254 vdd.n2253 0.152939
R21647 vdd.n2254 vdd.n1504 0.152939
R21648 vdd.n2270 vdd.n1504 0.152939
R21649 vdd.n2271 vdd.n2270 0.152939
R21650 vdd.n2272 vdd.n2271 0.152939
R21651 vdd.n670 vdd.n667 0.152939
R21652 vdd.n671 vdd.n670 0.152939
R21653 vdd.n672 vdd.n671 0.152939
R21654 vdd.n673 vdd.n672 0.152939
R21655 vdd.n676 vdd.n673 0.152939
R21656 vdd.n677 vdd.n676 0.152939
R21657 vdd.n678 vdd.n677 0.152939
R21658 vdd.n679 vdd.n678 0.152939
R21659 vdd.n682 vdd.n679 0.152939
R21660 vdd.n683 vdd.n682 0.152939
R21661 vdd.n684 vdd.n683 0.152939
R21662 vdd.n685 vdd.n684 0.152939
R21663 vdd.n690 vdd.n685 0.152939
R21664 vdd.n691 vdd.n690 0.152939
R21665 vdd.n692 vdd.n691 0.152939
R21666 vdd.n693 vdd.n692 0.152939
R21667 vdd.n696 vdd.n693 0.152939
R21668 vdd.n697 vdd.n696 0.152939
R21669 vdd.n698 vdd.n697 0.152939
R21670 vdd.n699 vdd.n698 0.152939
R21671 vdd.n702 vdd.n699 0.152939
R21672 vdd.n703 vdd.n702 0.152939
R21673 vdd.n704 vdd.n703 0.152939
R21674 vdd.n705 vdd.n704 0.152939
R21675 vdd.n708 vdd.n705 0.152939
R21676 vdd.n709 vdd.n708 0.152939
R21677 vdd.n710 vdd.n709 0.152939
R21678 vdd.n711 vdd.n710 0.152939
R21679 vdd.n714 vdd.n711 0.152939
R21680 vdd.n715 vdd.n714 0.152939
R21681 vdd.n716 vdd.n715 0.152939
R21682 vdd.n717 vdd.n716 0.152939
R21683 vdd.n720 vdd.n717 0.152939
R21684 vdd.n721 vdd.n720 0.152939
R21685 vdd.n3330 vdd.n721 0.152939
R21686 vdd.n3330 vdd.n3329 0.152939
R21687 vdd.n3329 vdd.n3328 0.152939
R21688 vdd.n3328 vdd.n725 0.152939
R21689 vdd.n730 vdd.n725 0.152939
R21690 vdd.n731 vdd.n730 0.152939
R21691 vdd.n734 vdd.n731 0.152939
R21692 vdd.n735 vdd.n734 0.152939
R21693 vdd.n736 vdd.n735 0.152939
R21694 vdd.n737 vdd.n736 0.152939
R21695 vdd.n740 vdd.n737 0.152939
R21696 vdd.n741 vdd.n740 0.152939
R21697 vdd.n742 vdd.n741 0.152939
R21698 vdd.n743 vdd.n742 0.152939
R21699 vdd.n746 vdd.n743 0.152939
R21700 vdd.n747 vdd.n746 0.152939
R21701 vdd.n748 vdd.n747 0.152939
R21702 vdd.n3413 vdd.n661 0.152939
R21703 vdd.n3414 vdd.n651 0.152939
R21704 vdd.n3428 vdd.n651 0.152939
R21705 vdd.n3429 vdd.n3428 0.152939
R21706 vdd.n3430 vdd.n3429 0.152939
R21707 vdd.n3430 vdd.n639 0.152939
R21708 vdd.n3444 vdd.n639 0.152939
R21709 vdd.n3445 vdd.n3444 0.152939
R21710 vdd.n3446 vdd.n3445 0.152939
R21711 vdd.n3446 vdd.n627 0.152939
R21712 vdd.n3461 vdd.n627 0.152939
R21713 vdd.n3462 vdd.n3461 0.152939
R21714 vdd.n3463 vdd.n3462 0.152939
R21715 vdd.n3463 vdd.n616 0.152939
R21716 vdd.n3480 vdd.n616 0.152939
R21717 vdd.n3481 vdd.n3480 0.152939
R21718 vdd.n3482 vdd.n3481 0.152939
R21719 vdd.n3482 vdd.n322 0.152939
R21720 vdd.n3562 vdd.n323 0.152939
R21721 vdd.n334 vdd.n323 0.152939
R21722 vdd.n335 vdd.n334 0.152939
R21723 vdd.n336 vdd.n335 0.152939
R21724 vdd.n343 vdd.n336 0.152939
R21725 vdd.n344 vdd.n343 0.152939
R21726 vdd.n345 vdd.n344 0.152939
R21727 vdd.n346 vdd.n345 0.152939
R21728 vdd.n354 vdd.n346 0.152939
R21729 vdd.n355 vdd.n354 0.152939
R21730 vdd.n356 vdd.n355 0.152939
R21731 vdd.n357 vdd.n356 0.152939
R21732 vdd.n365 vdd.n357 0.152939
R21733 vdd.n366 vdd.n365 0.152939
R21734 vdd.n367 vdd.n366 0.152939
R21735 vdd.n368 vdd.n367 0.152939
R21736 vdd.n443 vdd.n368 0.152939
R21737 vdd.n444 vdd.n442 0.152939
R21738 vdd.n451 vdd.n442 0.152939
R21739 vdd.n452 vdd.n451 0.152939
R21740 vdd.n453 vdd.n452 0.152939
R21741 vdd.n453 vdd.n440 0.152939
R21742 vdd.n461 vdd.n440 0.152939
R21743 vdd.n462 vdd.n461 0.152939
R21744 vdd.n463 vdd.n462 0.152939
R21745 vdd.n463 vdd.n438 0.152939
R21746 vdd.n471 vdd.n438 0.152939
R21747 vdd.n472 vdd.n471 0.152939
R21748 vdd.n473 vdd.n472 0.152939
R21749 vdd.n473 vdd.n436 0.152939
R21750 vdd.n481 vdd.n436 0.152939
R21751 vdd.n482 vdd.n481 0.152939
R21752 vdd.n483 vdd.n482 0.152939
R21753 vdd.n483 vdd.n434 0.152939
R21754 vdd.n491 vdd.n434 0.152939
R21755 vdd.n492 vdd.n491 0.152939
R21756 vdd.n493 vdd.n492 0.152939
R21757 vdd.n493 vdd.n430 0.152939
R21758 vdd.n501 vdd.n430 0.152939
R21759 vdd.n502 vdd.n501 0.152939
R21760 vdd.n503 vdd.n502 0.152939
R21761 vdd.n503 vdd.n428 0.152939
R21762 vdd.n511 vdd.n428 0.152939
R21763 vdd.n512 vdd.n511 0.152939
R21764 vdd.n513 vdd.n512 0.152939
R21765 vdd.n513 vdd.n426 0.152939
R21766 vdd.n521 vdd.n426 0.152939
R21767 vdd.n522 vdd.n521 0.152939
R21768 vdd.n523 vdd.n522 0.152939
R21769 vdd.n523 vdd.n424 0.152939
R21770 vdd.n531 vdd.n424 0.152939
R21771 vdd.n532 vdd.n531 0.152939
R21772 vdd.n533 vdd.n532 0.152939
R21773 vdd.n533 vdd.n422 0.152939
R21774 vdd.n541 vdd.n422 0.152939
R21775 vdd.n542 vdd.n541 0.152939
R21776 vdd.n543 vdd.n542 0.152939
R21777 vdd.n543 vdd.n418 0.152939
R21778 vdd.n551 vdd.n418 0.152939
R21779 vdd.n552 vdd.n551 0.152939
R21780 vdd.n553 vdd.n552 0.152939
R21781 vdd.n553 vdd.n416 0.152939
R21782 vdd.n561 vdd.n416 0.152939
R21783 vdd.n562 vdd.n561 0.152939
R21784 vdd.n563 vdd.n562 0.152939
R21785 vdd.n563 vdd.n414 0.152939
R21786 vdd.n571 vdd.n414 0.152939
R21787 vdd.n572 vdd.n571 0.152939
R21788 vdd.n573 vdd.n572 0.152939
R21789 vdd.n573 vdd.n412 0.152939
R21790 vdd.n581 vdd.n412 0.152939
R21791 vdd.n582 vdd.n581 0.152939
R21792 vdd.n583 vdd.n582 0.152939
R21793 vdd.n583 vdd.n410 0.152939
R21794 vdd.n591 vdd.n410 0.152939
R21795 vdd.n592 vdd.n591 0.152939
R21796 vdd.n593 vdd.n592 0.152939
R21797 vdd.n593 vdd.n408 0.152939
R21798 vdd.n600 vdd.n408 0.152939
R21799 vdd.n3521 vdd.n600 0.152939
R21800 vdd.n3421 vdd.n3420 0.152939
R21801 vdd.n3422 vdd.n3421 0.152939
R21802 vdd.n3422 vdd.n645 0.152939
R21803 vdd.n3436 vdd.n645 0.152939
R21804 vdd.n3437 vdd.n3436 0.152939
R21805 vdd.n3438 vdd.n3437 0.152939
R21806 vdd.n3438 vdd.n632 0.152939
R21807 vdd.n3452 vdd.n632 0.152939
R21808 vdd.n3453 vdd.n3452 0.152939
R21809 vdd.n3454 vdd.n3453 0.152939
R21810 vdd.n3454 vdd.n621 0.152939
R21811 vdd.n3469 vdd.n621 0.152939
R21812 vdd.n3470 vdd.n3469 0.152939
R21813 vdd.n3471 vdd.n3470 0.152939
R21814 vdd.n3473 vdd.n3471 0.152939
R21815 vdd.n3473 vdd.n3472 0.152939
R21816 vdd.n3472 vdd.n611 0.152939
R21817 vdd.n611 vdd.n609 0.152939
R21818 vdd.n3491 vdd.n609 0.152939
R21819 vdd.n3492 vdd.n3491 0.152939
R21820 vdd.n3493 vdd.n3492 0.152939
R21821 vdd.n3493 vdd.n607 0.152939
R21822 vdd.n3498 vdd.n607 0.152939
R21823 vdd.n3499 vdd.n3498 0.152939
R21824 vdd.n3500 vdd.n3499 0.152939
R21825 vdd.n3500 vdd.n605 0.152939
R21826 vdd.n3505 vdd.n605 0.152939
R21827 vdd.n3506 vdd.n3505 0.152939
R21828 vdd.n3507 vdd.n3506 0.152939
R21829 vdd.n3507 vdd.n603 0.152939
R21830 vdd.n3513 vdd.n603 0.152939
R21831 vdd.n3514 vdd.n3513 0.152939
R21832 vdd.n3515 vdd.n3514 0.152939
R21833 vdd.n3515 vdd.n601 0.152939
R21834 vdd.n3520 vdd.n601 0.152939
R21835 vdd.n3283 vdd.n656 0.152939
R21836 vdd.n2283 vdd.n1488 0.152939
R21837 vdd.n1834 vdd.n1833 0.152939
R21838 vdd.n1834 vdd.n1590 0.152939
R21839 vdd.n1848 vdd.n1590 0.152939
R21840 vdd.n1849 vdd.n1848 0.152939
R21841 vdd.n1850 vdd.n1849 0.152939
R21842 vdd.n1850 vdd.n1578 0.152939
R21843 vdd.n1865 vdd.n1578 0.152939
R21844 vdd.n1866 vdd.n1865 0.152939
R21845 vdd.n1867 vdd.n1866 0.152939
R21846 vdd.n1867 vdd.n1568 0.152939
R21847 vdd.n1882 vdd.n1568 0.152939
R21848 vdd.n1883 vdd.n1882 0.152939
R21849 vdd.n1884 vdd.n1883 0.152939
R21850 vdd.n1884 vdd.n1555 0.152939
R21851 vdd.n1898 vdd.n1555 0.152939
R21852 vdd.n1899 vdd.n1898 0.152939
R21853 vdd.n1900 vdd.n1899 0.152939
R21854 vdd.n1900 vdd.n1544 0.152939
R21855 vdd.n2210 vdd.n1544 0.152939
R21856 vdd.n2211 vdd.n2210 0.152939
R21857 vdd.n2212 vdd.n2211 0.152939
R21858 vdd.n2212 vdd.n1533 0.152939
R21859 vdd.n2226 vdd.n1533 0.152939
R21860 vdd.n2227 vdd.n2226 0.152939
R21861 vdd.n2228 vdd.n2227 0.152939
R21862 vdd.n2228 vdd.n1521 0.152939
R21863 vdd.n2243 vdd.n1521 0.152939
R21864 vdd.n2244 vdd.n2243 0.152939
R21865 vdd.n2245 vdd.n2244 0.152939
R21866 vdd.n2245 vdd.n1511 0.152939
R21867 vdd.n2260 vdd.n1511 0.152939
R21868 vdd.n2261 vdd.n2260 0.152939
R21869 vdd.n2264 vdd.n2261 0.152939
R21870 vdd.n2264 vdd.n2263 0.152939
R21871 vdd.n2263 vdd.n2262 0.152939
R21872 vdd.n1824 vdd.n1639 0.152939
R21873 vdd.n1824 vdd.n1823 0.152939
R21874 vdd.n1823 vdd.n1822 0.152939
R21875 vdd.n1822 vdd.n1641 0.152939
R21876 vdd.n1818 vdd.n1641 0.152939
R21877 vdd.n1818 vdd.n1817 0.152939
R21878 vdd.n1817 vdd.n1816 0.152939
R21879 vdd.n1816 vdd.n1646 0.152939
R21880 vdd.n1812 vdd.n1646 0.152939
R21881 vdd.n1812 vdd.n1811 0.152939
R21882 vdd.n1811 vdd.n1810 0.152939
R21883 vdd.n1810 vdd.n1652 0.152939
R21884 vdd.n1806 vdd.n1652 0.152939
R21885 vdd.n1806 vdd.n1805 0.152939
R21886 vdd.n1805 vdd.n1804 0.152939
R21887 vdd.n1804 vdd.n1658 0.152939
R21888 vdd.n1800 vdd.n1658 0.152939
R21889 vdd.n1800 vdd.n1799 0.152939
R21890 vdd.n1799 vdd.n1798 0.152939
R21891 vdd.n1798 vdd.n1664 0.152939
R21892 vdd.n1790 vdd.n1664 0.152939
R21893 vdd.n1790 vdd.n1789 0.152939
R21894 vdd.n1789 vdd.n1788 0.152939
R21895 vdd.n1788 vdd.n1668 0.152939
R21896 vdd.n1784 vdd.n1668 0.152939
R21897 vdd.n1784 vdd.n1783 0.152939
R21898 vdd.n1783 vdd.n1782 0.152939
R21899 vdd.n1782 vdd.n1674 0.152939
R21900 vdd.n1778 vdd.n1674 0.152939
R21901 vdd.n1778 vdd.n1777 0.152939
R21902 vdd.n1777 vdd.n1776 0.152939
R21903 vdd.n1776 vdd.n1680 0.152939
R21904 vdd.n1772 vdd.n1680 0.152939
R21905 vdd.n1772 vdd.n1771 0.152939
R21906 vdd.n1771 vdd.n1770 0.152939
R21907 vdd.n1770 vdd.n1686 0.152939
R21908 vdd.n1766 vdd.n1686 0.152939
R21909 vdd.n1766 vdd.n1765 0.152939
R21910 vdd.n1765 vdd.n1764 0.152939
R21911 vdd.n1764 vdd.n1692 0.152939
R21912 vdd.n1757 vdd.n1692 0.152939
R21913 vdd.n1757 vdd.n1756 0.152939
R21914 vdd.n1756 vdd.n1755 0.152939
R21915 vdd.n1755 vdd.n1697 0.152939
R21916 vdd.n1751 vdd.n1697 0.152939
R21917 vdd.n1751 vdd.n1750 0.152939
R21918 vdd.n1750 vdd.n1749 0.152939
R21919 vdd.n1749 vdd.n1703 0.152939
R21920 vdd.n1745 vdd.n1703 0.152939
R21921 vdd.n1745 vdd.n1744 0.152939
R21922 vdd.n1744 vdd.n1743 0.152939
R21923 vdd.n1743 vdd.n1709 0.152939
R21924 vdd.n1739 vdd.n1709 0.152939
R21925 vdd.n1739 vdd.n1738 0.152939
R21926 vdd.n1738 vdd.n1737 0.152939
R21927 vdd.n1737 vdd.n1715 0.152939
R21928 vdd.n1733 vdd.n1715 0.152939
R21929 vdd.n1733 vdd.n1732 0.152939
R21930 vdd.n1732 vdd.n1731 0.152939
R21931 vdd.n1731 vdd.n1721 0.152939
R21932 vdd.n1727 vdd.n1721 0.152939
R21933 vdd.n1727 vdd.n1602 0.152939
R21934 vdd.n1832 vdd.n1602 0.152939
R21935 vdd.n1840 vdd.n1596 0.152939
R21936 vdd.n1841 vdd.n1840 0.152939
R21937 vdd.n1842 vdd.n1841 0.152939
R21938 vdd.n1842 vdd.n1584 0.152939
R21939 vdd.n1857 vdd.n1584 0.152939
R21940 vdd.n1858 vdd.n1857 0.152939
R21941 vdd.n1859 vdd.n1858 0.152939
R21942 vdd.n1859 vdd.n1573 0.152939
R21943 vdd.n1874 vdd.n1573 0.152939
R21944 vdd.n1875 vdd.n1874 0.152939
R21945 vdd.n1876 vdd.n1875 0.152939
R21946 vdd.n1876 vdd.n1562 0.152939
R21947 vdd.n1890 vdd.n1562 0.152939
R21948 vdd.n1891 vdd.n1890 0.152939
R21949 vdd.n1892 vdd.n1891 0.152939
R21950 vdd.n1892 vdd.n1550 0.152939
R21951 vdd.n1907 vdd.n1550 0.152939
R21952 vdd.n2391 vdd.n2390 0.110256
R21953 vdd.n3214 vdd.n661 0.110256
R21954 vdd.n3283 vdd.n3282 0.110256
R21955 vdd.n2284 vdd.n2283 0.110256
R21956 vdd.n2203 vdd.n2202 0.0695946
R21957 vdd.n3563 vdd.n322 0.0695946
R21958 vdd.n3563 vdd.n3562 0.0695946
R21959 vdd.n2202 vdd.n1907 0.0695946
R21960 vdd.n2391 vdd.n1149 0.0431829
R21961 vdd.n2284 vdd.n1249 0.0431829
R21962 vdd.n3214 vdd.n667 0.0431829
R21963 vdd.n3282 vdd.n748 0.0431829
R21964 vdd vdd.n28 0.00833333
R21965 commonsourceibias.n397 commonsourceibias.t184 222.032
R21966 commonsourceibias.n281 commonsourceibias.t134 222.032
R21967 commonsourceibias.n44 commonsourceibias.t26 222.032
R21968 commonsourceibias.n166 commonsourceibias.t140 222.032
R21969 commonsourceibias.n875 commonsourceibias.t191 222.032
R21970 commonsourceibias.n759 commonsourceibias.t98 222.032
R21971 commonsourceibias.n529 commonsourceibias.t68 222.032
R21972 commonsourceibias.n645 commonsourceibias.t177 222.032
R21973 commonsourceibias.n480 commonsourceibias.t183 207.983
R21974 commonsourceibias.n364 commonsourceibias.t88 207.983
R21975 commonsourceibias.n127 commonsourceibias.t16 207.983
R21976 commonsourceibias.n249 commonsourceibias.t151 207.983
R21977 commonsourceibias.n963 commonsourceibias.t101 207.983
R21978 commonsourceibias.n847 commonsourceibias.t189 207.983
R21979 commonsourceibias.n617 commonsourceibias.t40 207.983
R21980 commonsourceibias.n732 commonsourceibias.t112 207.983
R21981 commonsourceibias.n396 commonsourceibias.t150 168.701
R21982 commonsourceibias.n402 commonsourceibias.t155 168.701
R21983 commonsourceibias.n408 commonsourceibias.t199 168.701
R21984 commonsourceibias.n392 commonsourceibias.t175 168.701
R21985 commonsourceibias.n416 commonsourceibias.t165 168.701
R21986 commonsourceibias.n422 commonsourceibias.t96 168.701
R21987 commonsourceibias.n387 commonsourceibias.t187 168.701
R21988 commonsourceibias.n430 commonsourceibias.t168 168.701
R21989 commonsourceibias.n436 commonsourceibias.t172 168.701
R21990 commonsourceibias.n382 commonsourceibias.t80 168.701
R21991 commonsourceibias.n444 commonsourceibias.t173 168.701
R21992 commonsourceibias.n450 commonsourceibias.t182 168.701
R21993 commonsourceibias.n377 commonsourceibias.t149 168.701
R21994 commonsourceibias.n458 commonsourceibias.t110 168.701
R21995 commonsourceibias.n464 commonsourceibias.t194 168.701
R21996 commonsourceibias.n372 commonsourceibias.t157 168.701
R21997 commonsourceibias.n472 commonsourceibias.t163 168.701
R21998 commonsourceibias.n478 commonsourceibias.t92 168.701
R21999 commonsourceibias.n362 commonsourceibias.t198 168.701
R22000 commonsourceibias.n356 commonsourceibias.t186 168.701
R22001 commonsourceibias.n256 commonsourceibias.t95 168.701
R22002 commonsourceibias.n348 commonsourceibias.t196 168.701
R22003 commonsourceibias.n342 commonsourceibias.t105 168.701
R22004 commonsourceibias.n261 commonsourceibias.t94 168.701
R22005 commonsourceibias.n334 commonsourceibias.t197 168.701
R22006 commonsourceibias.n328 commonsourceibias.t115 168.701
R22007 commonsourceibias.n266 commonsourceibias.t141 168.701
R22008 commonsourceibias.n320 commonsourceibias.t195 168.701
R22009 commonsourceibias.n314 commonsourceibias.t113 168.701
R22010 commonsourceibias.n271 commonsourceibias.t138 168.701
R22011 commonsourceibias.n306 commonsourceibias.t130 168.701
R22012 commonsourceibias.n300 commonsourceibias.t114 168.701
R22013 commonsourceibias.n276 commonsourceibias.t139 168.701
R22014 commonsourceibias.n292 commonsourceibias.t129 168.701
R22015 commonsourceibias.n286 commonsourceibias.t125 168.701
R22016 commonsourceibias.n280 commonsourceibias.t147 168.701
R22017 commonsourceibias.n125 commonsourceibias.t60 168.701
R22018 commonsourceibias.n119 commonsourceibias.t4 168.701
R22019 commonsourceibias.n19 commonsourceibias.t14 168.701
R22020 commonsourceibias.n111 commonsourceibias.t74 168.701
R22021 commonsourceibias.n105 commonsourceibias.t20 168.701
R22022 commonsourceibias.n24 commonsourceibias.t34 168.701
R22023 commonsourceibias.n97 commonsourceibias.t10 168.701
R22024 commonsourceibias.n91 commonsourceibias.t18 168.701
R22025 commonsourceibias.n29 commonsourceibias.t54 168.701
R22026 commonsourceibias.n83 commonsourceibias.t30 168.701
R22027 commonsourceibias.n77 commonsourceibias.t36 168.701
R22028 commonsourceibias.n34 commonsourceibias.t70 168.701
R22029 commonsourceibias.n69 commonsourceibias.t22 168.701
R22030 commonsourceibias.n63 commonsourceibias.t62 168.701
R22031 commonsourceibias.n39 commonsourceibias.t0 168.701
R22032 commonsourceibias.n55 commonsourceibias.t42 168.701
R22033 commonsourceibias.n49 commonsourceibias.t52 168.701
R22034 commonsourceibias.n43 commonsourceibias.t58 168.701
R22035 commonsourceibias.n247 commonsourceibias.t83 168.701
R22036 commonsourceibias.n241 commonsourceibias.t161 168.701
R22037 commonsourceibias.n5 commonsourceibias.t152 168.701
R22038 commonsourceibias.n233 commonsourceibias.t171 168.701
R22039 commonsourceibias.n227 commonsourceibias.t145 168.701
R22040 commonsourceibias.n10 commonsourceibias.t124 168.701
R22041 commonsourceibias.n219 commonsourceibias.t158 168.701
R22042 commonsourceibias.n213 commonsourceibias.t148 168.701
R22043 commonsourceibias.n150 commonsourceibias.t93 168.701
R22044 commonsourceibias.n151 commonsourceibias.t131 168.701
R22045 commonsourceibias.n153 commonsourceibias.t117 168.701
R22046 commonsourceibias.n155 commonsourceibias.t176 168.701
R22047 commonsourceibias.n191 commonsourceibias.t144 168.701
R22048 commonsourceibias.n185 commonsourceibias.t190 168.701
R22049 commonsourceibias.n161 commonsourceibias.t164 168.701
R22050 commonsourceibias.n177 commonsourceibias.t111 168.701
R22051 commonsourceibias.n171 commonsourceibias.t100 168.701
R22052 commonsourceibias.n165 commonsourceibias.t84 168.701
R22053 commonsourceibias.n874 commonsourceibias.t156 168.701
R22054 commonsourceibias.n880 commonsourceibias.t146 168.701
R22055 commonsourceibias.n886 commonsourceibias.t126 168.701
R22056 commonsourceibias.n888 commonsourceibias.t91 168.701
R22057 commonsourceibias.n895 commonsourceibias.t181 168.701
R22058 commonsourceibias.n901 commonsourceibias.t136 168.701
R22059 commonsourceibias.n903 commonsourceibias.t107 168.701
R22060 commonsourceibias.n910 commonsourceibias.t192 168.701
R22061 commonsourceibias.n916 commonsourceibias.t167 168.701
R22062 commonsourceibias.n918 commonsourceibias.t127 168.701
R22063 commonsourceibias.n925 commonsourceibias.t87 168.701
R22064 commonsourceibias.n931 commonsourceibias.t99 168.701
R22065 commonsourceibias.n933 commonsourceibias.t137 168.701
R22066 commonsourceibias.n940 commonsourceibias.t143 168.701
R22067 commonsourceibias.n946 commonsourceibias.t122 168.701
R22068 commonsourceibias.n948 commonsourceibias.t170 168.701
R22069 commonsourceibias.n955 commonsourceibias.t153 168.701
R22070 commonsourceibias.n961 commonsourceibias.t133 168.701
R22071 commonsourceibias.n758 commonsourceibias.t123 168.701
R22072 commonsourceibias.n764 commonsourceibias.t132 168.701
R22073 commonsourceibias.n770 commonsourceibias.t104 168.701
R22074 commonsourceibias.n772 commonsourceibias.t118 168.701
R22075 commonsourceibias.n779 commonsourceibias.t85 168.701
R22076 commonsourceibias.n785 commonsourceibias.t106 168.701
R22077 commonsourceibias.n787 commonsourceibias.t119 168.701
R22078 commonsourceibias.n794 commonsourceibias.t86 168.701
R22079 commonsourceibias.n800 commonsourceibias.t97 168.701
R22080 commonsourceibias.n802 commonsourceibias.t120 168.701
R22081 commonsourceibias.n809 commonsourceibias.t89 168.701
R22082 commonsourceibias.n815 commonsourceibias.t178 168.701
R22083 commonsourceibias.n817 commonsourceibias.t121 168.701
R22084 commonsourceibias.n824 commonsourceibias.t81 168.701
R22085 commonsourceibias.n830 commonsourceibias.t179 168.701
R22086 commonsourceibias.n832 commonsourceibias.t193 168.701
R22087 commonsourceibias.n839 commonsourceibias.t82 168.701
R22088 commonsourceibias.n845 commonsourceibias.t180 168.701
R22089 commonsourceibias.n528 commonsourceibias.t8 168.701
R22090 commonsourceibias.n534 commonsourceibias.t6 168.701
R22091 commonsourceibias.n540 commonsourceibias.t66 168.701
R22092 commonsourceibias.n542 commonsourceibias.t28 168.701
R22093 commonsourceibias.n549 commonsourceibias.t78 168.701
R22094 commonsourceibias.n555 commonsourceibias.t48 168.701
R22095 commonsourceibias.n557 commonsourceibias.t2 168.701
R22096 commonsourceibias.n564 commonsourceibias.t64 168.701
R22097 commonsourceibias.n570 commonsourceibias.t50 168.701
R22098 commonsourceibias.n572 commonsourceibias.t72 168.701
R22099 commonsourceibias.n579 commonsourceibias.t44 168.701
R22100 commonsourceibias.n585 commonsourceibias.t32 168.701
R22101 commonsourceibias.n587 commonsourceibias.t56 168.701
R22102 commonsourceibias.n594 commonsourceibias.t46 168.701
R22103 commonsourceibias.n600 commonsourceibias.t12 168.701
R22104 commonsourceibias.n602 commonsourceibias.t38 168.701
R22105 commonsourceibias.n609 commonsourceibias.t24 168.701
R22106 commonsourceibias.n615 commonsourceibias.t76 168.701
R22107 commonsourceibias.n730 commonsourceibias.t169 168.701
R22108 commonsourceibias.n724 commonsourceibias.t142 168.701
R22109 commonsourceibias.n717 commonsourceibias.t116 168.701
R22110 commonsourceibias.n715 commonsourceibias.t154 168.701
R22111 commonsourceibias.n709 commonsourceibias.t108 168.701
R22112 commonsourceibias.n702 commonsourceibias.t90 168.701
R22113 commonsourceibias.n700 commonsourceibias.t128 168.701
R22114 commonsourceibias.n694 commonsourceibias.t109 168.701
R22115 commonsourceibias.n687 commonsourceibias.t174 168.701
R22116 commonsourceibias.n644 commonsourceibias.t159 168.701
R22117 commonsourceibias.n650 commonsourceibias.t160 168.701
R22118 commonsourceibias.n656 commonsourceibias.t185 168.701
R22119 commonsourceibias.n658 commonsourceibias.t135 168.701
R22120 commonsourceibias.n665 commonsourceibias.t166 168.701
R22121 commonsourceibias.n671 commonsourceibias.t103 168.701
R22122 commonsourceibias.n635 commonsourceibias.t162 168.701
R22123 commonsourceibias.n633 commonsourceibias.t188 168.701
R22124 commonsourceibias.n631 commonsourceibias.t102 168.701
R22125 commonsourceibias.n479 commonsourceibias.n367 161.3
R22126 commonsourceibias.n477 commonsourceibias.n476 161.3
R22127 commonsourceibias.n475 commonsourceibias.n368 161.3
R22128 commonsourceibias.n474 commonsourceibias.n473 161.3
R22129 commonsourceibias.n471 commonsourceibias.n369 161.3
R22130 commonsourceibias.n470 commonsourceibias.n469 161.3
R22131 commonsourceibias.n468 commonsourceibias.n370 161.3
R22132 commonsourceibias.n467 commonsourceibias.n466 161.3
R22133 commonsourceibias.n465 commonsourceibias.n371 161.3
R22134 commonsourceibias.n463 commonsourceibias.n462 161.3
R22135 commonsourceibias.n461 commonsourceibias.n373 161.3
R22136 commonsourceibias.n460 commonsourceibias.n459 161.3
R22137 commonsourceibias.n457 commonsourceibias.n374 161.3
R22138 commonsourceibias.n456 commonsourceibias.n455 161.3
R22139 commonsourceibias.n454 commonsourceibias.n375 161.3
R22140 commonsourceibias.n453 commonsourceibias.n452 161.3
R22141 commonsourceibias.n451 commonsourceibias.n376 161.3
R22142 commonsourceibias.n449 commonsourceibias.n448 161.3
R22143 commonsourceibias.n447 commonsourceibias.n378 161.3
R22144 commonsourceibias.n446 commonsourceibias.n445 161.3
R22145 commonsourceibias.n443 commonsourceibias.n379 161.3
R22146 commonsourceibias.n442 commonsourceibias.n441 161.3
R22147 commonsourceibias.n440 commonsourceibias.n380 161.3
R22148 commonsourceibias.n439 commonsourceibias.n438 161.3
R22149 commonsourceibias.n437 commonsourceibias.n381 161.3
R22150 commonsourceibias.n435 commonsourceibias.n434 161.3
R22151 commonsourceibias.n433 commonsourceibias.n383 161.3
R22152 commonsourceibias.n432 commonsourceibias.n431 161.3
R22153 commonsourceibias.n429 commonsourceibias.n384 161.3
R22154 commonsourceibias.n428 commonsourceibias.n427 161.3
R22155 commonsourceibias.n426 commonsourceibias.n385 161.3
R22156 commonsourceibias.n425 commonsourceibias.n424 161.3
R22157 commonsourceibias.n423 commonsourceibias.n386 161.3
R22158 commonsourceibias.n421 commonsourceibias.n420 161.3
R22159 commonsourceibias.n419 commonsourceibias.n388 161.3
R22160 commonsourceibias.n418 commonsourceibias.n417 161.3
R22161 commonsourceibias.n415 commonsourceibias.n389 161.3
R22162 commonsourceibias.n414 commonsourceibias.n413 161.3
R22163 commonsourceibias.n412 commonsourceibias.n390 161.3
R22164 commonsourceibias.n411 commonsourceibias.n410 161.3
R22165 commonsourceibias.n409 commonsourceibias.n391 161.3
R22166 commonsourceibias.n407 commonsourceibias.n406 161.3
R22167 commonsourceibias.n405 commonsourceibias.n393 161.3
R22168 commonsourceibias.n404 commonsourceibias.n403 161.3
R22169 commonsourceibias.n401 commonsourceibias.n394 161.3
R22170 commonsourceibias.n400 commonsourceibias.n399 161.3
R22171 commonsourceibias.n398 commonsourceibias.n395 161.3
R22172 commonsourceibias.n282 commonsourceibias.n279 161.3
R22173 commonsourceibias.n284 commonsourceibias.n283 161.3
R22174 commonsourceibias.n285 commonsourceibias.n278 161.3
R22175 commonsourceibias.n288 commonsourceibias.n287 161.3
R22176 commonsourceibias.n289 commonsourceibias.n277 161.3
R22177 commonsourceibias.n291 commonsourceibias.n290 161.3
R22178 commonsourceibias.n293 commonsourceibias.n275 161.3
R22179 commonsourceibias.n295 commonsourceibias.n294 161.3
R22180 commonsourceibias.n296 commonsourceibias.n274 161.3
R22181 commonsourceibias.n298 commonsourceibias.n297 161.3
R22182 commonsourceibias.n299 commonsourceibias.n273 161.3
R22183 commonsourceibias.n302 commonsourceibias.n301 161.3
R22184 commonsourceibias.n303 commonsourceibias.n272 161.3
R22185 commonsourceibias.n305 commonsourceibias.n304 161.3
R22186 commonsourceibias.n307 commonsourceibias.n270 161.3
R22187 commonsourceibias.n309 commonsourceibias.n308 161.3
R22188 commonsourceibias.n310 commonsourceibias.n269 161.3
R22189 commonsourceibias.n312 commonsourceibias.n311 161.3
R22190 commonsourceibias.n313 commonsourceibias.n268 161.3
R22191 commonsourceibias.n316 commonsourceibias.n315 161.3
R22192 commonsourceibias.n317 commonsourceibias.n267 161.3
R22193 commonsourceibias.n319 commonsourceibias.n318 161.3
R22194 commonsourceibias.n321 commonsourceibias.n265 161.3
R22195 commonsourceibias.n323 commonsourceibias.n322 161.3
R22196 commonsourceibias.n324 commonsourceibias.n264 161.3
R22197 commonsourceibias.n326 commonsourceibias.n325 161.3
R22198 commonsourceibias.n327 commonsourceibias.n263 161.3
R22199 commonsourceibias.n330 commonsourceibias.n329 161.3
R22200 commonsourceibias.n331 commonsourceibias.n262 161.3
R22201 commonsourceibias.n333 commonsourceibias.n332 161.3
R22202 commonsourceibias.n335 commonsourceibias.n260 161.3
R22203 commonsourceibias.n337 commonsourceibias.n336 161.3
R22204 commonsourceibias.n338 commonsourceibias.n259 161.3
R22205 commonsourceibias.n340 commonsourceibias.n339 161.3
R22206 commonsourceibias.n341 commonsourceibias.n258 161.3
R22207 commonsourceibias.n344 commonsourceibias.n343 161.3
R22208 commonsourceibias.n345 commonsourceibias.n257 161.3
R22209 commonsourceibias.n347 commonsourceibias.n346 161.3
R22210 commonsourceibias.n349 commonsourceibias.n255 161.3
R22211 commonsourceibias.n351 commonsourceibias.n350 161.3
R22212 commonsourceibias.n352 commonsourceibias.n254 161.3
R22213 commonsourceibias.n354 commonsourceibias.n353 161.3
R22214 commonsourceibias.n355 commonsourceibias.n253 161.3
R22215 commonsourceibias.n358 commonsourceibias.n357 161.3
R22216 commonsourceibias.n359 commonsourceibias.n252 161.3
R22217 commonsourceibias.n361 commonsourceibias.n360 161.3
R22218 commonsourceibias.n363 commonsourceibias.n251 161.3
R22219 commonsourceibias.n45 commonsourceibias.n42 161.3
R22220 commonsourceibias.n47 commonsourceibias.n46 161.3
R22221 commonsourceibias.n48 commonsourceibias.n41 161.3
R22222 commonsourceibias.n51 commonsourceibias.n50 161.3
R22223 commonsourceibias.n52 commonsourceibias.n40 161.3
R22224 commonsourceibias.n54 commonsourceibias.n53 161.3
R22225 commonsourceibias.n56 commonsourceibias.n38 161.3
R22226 commonsourceibias.n58 commonsourceibias.n57 161.3
R22227 commonsourceibias.n59 commonsourceibias.n37 161.3
R22228 commonsourceibias.n61 commonsourceibias.n60 161.3
R22229 commonsourceibias.n62 commonsourceibias.n36 161.3
R22230 commonsourceibias.n65 commonsourceibias.n64 161.3
R22231 commonsourceibias.n66 commonsourceibias.n35 161.3
R22232 commonsourceibias.n68 commonsourceibias.n67 161.3
R22233 commonsourceibias.n70 commonsourceibias.n33 161.3
R22234 commonsourceibias.n72 commonsourceibias.n71 161.3
R22235 commonsourceibias.n73 commonsourceibias.n32 161.3
R22236 commonsourceibias.n75 commonsourceibias.n74 161.3
R22237 commonsourceibias.n76 commonsourceibias.n31 161.3
R22238 commonsourceibias.n79 commonsourceibias.n78 161.3
R22239 commonsourceibias.n80 commonsourceibias.n30 161.3
R22240 commonsourceibias.n82 commonsourceibias.n81 161.3
R22241 commonsourceibias.n84 commonsourceibias.n28 161.3
R22242 commonsourceibias.n86 commonsourceibias.n85 161.3
R22243 commonsourceibias.n87 commonsourceibias.n27 161.3
R22244 commonsourceibias.n89 commonsourceibias.n88 161.3
R22245 commonsourceibias.n90 commonsourceibias.n26 161.3
R22246 commonsourceibias.n93 commonsourceibias.n92 161.3
R22247 commonsourceibias.n94 commonsourceibias.n25 161.3
R22248 commonsourceibias.n96 commonsourceibias.n95 161.3
R22249 commonsourceibias.n98 commonsourceibias.n23 161.3
R22250 commonsourceibias.n100 commonsourceibias.n99 161.3
R22251 commonsourceibias.n101 commonsourceibias.n22 161.3
R22252 commonsourceibias.n103 commonsourceibias.n102 161.3
R22253 commonsourceibias.n104 commonsourceibias.n21 161.3
R22254 commonsourceibias.n107 commonsourceibias.n106 161.3
R22255 commonsourceibias.n108 commonsourceibias.n20 161.3
R22256 commonsourceibias.n110 commonsourceibias.n109 161.3
R22257 commonsourceibias.n112 commonsourceibias.n18 161.3
R22258 commonsourceibias.n114 commonsourceibias.n113 161.3
R22259 commonsourceibias.n115 commonsourceibias.n17 161.3
R22260 commonsourceibias.n117 commonsourceibias.n116 161.3
R22261 commonsourceibias.n118 commonsourceibias.n16 161.3
R22262 commonsourceibias.n121 commonsourceibias.n120 161.3
R22263 commonsourceibias.n122 commonsourceibias.n15 161.3
R22264 commonsourceibias.n124 commonsourceibias.n123 161.3
R22265 commonsourceibias.n126 commonsourceibias.n14 161.3
R22266 commonsourceibias.n167 commonsourceibias.n164 161.3
R22267 commonsourceibias.n169 commonsourceibias.n168 161.3
R22268 commonsourceibias.n170 commonsourceibias.n163 161.3
R22269 commonsourceibias.n173 commonsourceibias.n172 161.3
R22270 commonsourceibias.n174 commonsourceibias.n162 161.3
R22271 commonsourceibias.n176 commonsourceibias.n175 161.3
R22272 commonsourceibias.n178 commonsourceibias.n160 161.3
R22273 commonsourceibias.n180 commonsourceibias.n179 161.3
R22274 commonsourceibias.n181 commonsourceibias.n159 161.3
R22275 commonsourceibias.n183 commonsourceibias.n182 161.3
R22276 commonsourceibias.n184 commonsourceibias.n158 161.3
R22277 commonsourceibias.n187 commonsourceibias.n186 161.3
R22278 commonsourceibias.n188 commonsourceibias.n157 161.3
R22279 commonsourceibias.n190 commonsourceibias.n189 161.3
R22280 commonsourceibias.n192 commonsourceibias.n156 161.3
R22281 commonsourceibias.n194 commonsourceibias.n193 161.3
R22282 commonsourceibias.n196 commonsourceibias.n195 161.3
R22283 commonsourceibias.n197 commonsourceibias.n154 161.3
R22284 commonsourceibias.n199 commonsourceibias.n198 161.3
R22285 commonsourceibias.n201 commonsourceibias.n200 161.3
R22286 commonsourceibias.n202 commonsourceibias.n152 161.3
R22287 commonsourceibias.n204 commonsourceibias.n203 161.3
R22288 commonsourceibias.n206 commonsourceibias.n205 161.3
R22289 commonsourceibias.n208 commonsourceibias.n207 161.3
R22290 commonsourceibias.n209 commonsourceibias.n13 161.3
R22291 commonsourceibias.n211 commonsourceibias.n210 161.3
R22292 commonsourceibias.n212 commonsourceibias.n12 161.3
R22293 commonsourceibias.n215 commonsourceibias.n214 161.3
R22294 commonsourceibias.n216 commonsourceibias.n11 161.3
R22295 commonsourceibias.n218 commonsourceibias.n217 161.3
R22296 commonsourceibias.n220 commonsourceibias.n9 161.3
R22297 commonsourceibias.n222 commonsourceibias.n221 161.3
R22298 commonsourceibias.n223 commonsourceibias.n8 161.3
R22299 commonsourceibias.n225 commonsourceibias.n224 161.3
R22300 commonsourceibias.n226 commonsourceibias.n7 161.3
R22301 commonsourceibias.n229 commonsourceibias.n228 161.3
R22302 commonsourceibias.n230 commonsourceibias.n6 161.3
R22303 commonsourceibias.n232 commonsourceibias.n231 161.3
R22304 commonsourceibias.n234 commonsourceibias.n4 161.3
R22305 commonsourceibias.n236 commonsourceibias.n235 161.3
R22306 commonsourceibias.n237 commonsourceibias.n3 161.3
R22307 commonsourceibias.n239 commonsourceibias.n238 161.3
R22308 commonsourceibias.n240 commonsourceibias.n2 161.3
R22309 commonsourceibias.n243 commonsourceibias.n242 161.3
R22310 commonsourceibias.n244 commonsourceibias.n1 161.3
R22311 commonsourceibias.n246 commonsourceibias.n245 161.3
R22312 commonsourceibias.n248 commonsourceibias.n0 161.3
R22313 commonsourceibias.n962 commonsourceibias.n850 161.3
R22314 commonsourceibias.n960 commonsourceibias.n959 161.3
R22315 commonsourceibias.n958 commonsourceibias.n851 161.3
R22316 commonsourceibias.n957 commonsourceibias.n956 161.3
R22317 commonsourceibias.n954 commonsourceibias.n852 161.3
R22318 commonsourceibias.n953 commonsourceibias.n952 161.3
R22319 commonsourceibias.n951 commonsourceibias.n853 161.3
R22320 commonsourceibias.n950 commonsourceibias.n949 161.3
R22321 commonsourceibias.n947 commonsourceibias.n854 161.3
R22322 commonsourceibias.n945 commonsourceibias.n944 161.3
R22323 commonsourceibias.n943 commonsourceibias.n855 161.3
R22324 commonsourceibias.n942 commonsourceibias.n941 161.3
R22325 commonsourceibias.n939 commonsourceibias.n856 161.3
R22326 commonsourceibias.n938 commonsourceibias.n937 161.3
R22327 commonsourceibias.n936 commonsourceibias.n857 161.3
R22328 commonsourceibias.n935 commonsourceibias.n934 161.3
R22329 commonsourceibias.n932 commonsourceibias.n858 161.3
R22330 commonsourceibias.n930 commonsourceibias.n929 161.3
R22331 commonsourceibias.n928 commonsourceibias.n859 161.3
R22332 commonsourceibias.n927 commonsourceibias.n926 161.3
R22333 commonsourceibias.n924 commonsourceibias.n860 161.3
R22334 commonsourceibias.n923 commonsourceibias.n922 161.3
R22335 commonsourceibias.n921 commonsourceibias.n861 161.3
R22336 commonsourceibias.n920 commonsourceibias.n919 161.3
R22337 commonsourceibias.n917 commonsourceibias.n862 161.3
R22338 commonsourceibias.n915 commonsourceibias.n914 161.3
R22339 commonsourceibias.n913 commonsourceibias.n863 161.3
R22340 commonsourceibias.n912 commonsourceibias.n911 161.3
R22341 commonsourceibias.n909 commonsourceibias.n864 161.3
R22342 commonsourceibias.n908 commonsourceibias.n907 161.3
R22343 commonsourceibias.n906 commonsourceibias.n865 161.3
R22344 commonsourceibias.n905 commonsourceibias.n904 161.3
R22345 commonsourceibias.n902 commonsourceibias.n866 161.3
R22346 commonsourceibias.n900 commonsourceibias.n899 161.3
R22347 commonsourceibias.n898 commonsourceibias.n867 161.3
R22348 commonsourceibias.n897 commonsourceibias.n896 161.3
R22349 commonsourceibias.n894 commonsourceibias.n868 161.3
R22350 commonsourceibias.n893 commonsourceibias.n892 161.3
R22351 commonsourceibias.n891 commonsourceibias.n869 161.3
R22352 commonsourceibias.n890 commonsourceibias.n889 161.3
R22353 commonsourceibias.n887 commonsourceibias.n870 161.3
R22354 commonsourceibias.n885 commonsourceibias.n884 161.3
R22355 commonsourceibias.n883 commonsourceibias.n871 161.3
R22356 commonsourceibias.n882 commonsourceibias.n881 161.3
R22357 commonsourceibias.n879 commonsourceibias.n872 161.3
R22358 commonsourceibias.n878 commonsourceibias.n877 161.3
R22359 commonsourceibias.n876 commonsourceibias.n873 161.3
R22360 commonsourceibias.n846 commonsourceibias.n734 161.3
R22361 commonsourceibias.n844 commonsourceibias.n843 161.3
R22362 commonsourceibias.n842 commonsourceibias.n735 161.3
R22363 commonsourceibias.n841 commonsourceibias.n840 161.3
R22364 commonsourceibias.n838 commonsourceibias.n736 161.3
R22365 commonsourceibias.n837 commonsourceibias.n836 161.3
R22366 commonsourceibias.n835 commonsourceibias.n737 161.3
R22367 commonsourceibias.n834 commonsourceibias.n833 161.3
R22368 commonsourceibias.n831 commonsourceibias.n738 161.3
R22369 commonsourceibias.n829 commonsourceibias.n828 161.3
R22370 commonsourceibias.n827 commonsourceibias.n739 161.3
R22371 commonsourceibias.n826 commonsourceibias.n825 161.3
R22372 commonsourceibias.n823 commonsourceibias.n740 161.3
R22373 commonsourceibias.n822 commonsourceibias.n821 161.3
R22374 commonsourceibias.n820 commonsourceibias.n741 161.3
R22375 commonsourceibias.n819 commonsourceibias.n818 161.3
R22376 commonsourceibias.n816 commonsourceibias.n742 161.3
R22377 commonsourceibias.n814 commonsourceibias.n813 161.3
R22378 commonsourceibias.n812 commonsourceibias.n743 161.3
R22379 commonsourceibias.n811 commonsourceibias.n810 161.3
R22380 commonsourceibias.n808 commonsourceibias.n744 161.3
R22381 commonsourceibias.n807 commonsourceibias.n806 161.3
R22382 commonsourceibias.n805 commonsourceibias.n745 161.3
R22383 commonsourceibias.n804 commonsourceibias.n803 161.3
R22384 commonsourceibias.n801 commonsourceibias.n746 161.3
R22385 commonsourceibias.n799 commonsourceibias.n798 161.3
R22386 commonsourceibias.n797 commonsourceibias.n747 161.3
R22387 commonsourceibias.n796 commonsourceibias.n795 161.3
R22388 commonsourceibias.n793 commonsourceibias.n748 161.3
R22389 commonsourceibias.n792 commonsourceibias.n791 161.3
R22390 commonsourceibias.n790 commonsourceibias.n749 161.3
R22391 commonsourceibias.n789 commonsourceibias.n788 161.3
R22392 commonsourceibias.n786 commonsourceibias.n750 161.3
R22393 commonsourceibias.n784 commonsourceibias.n783 161.3
R22394 commonsourceibias.n782 commonsourceibias.n751 161.3
R22395 commonsourceibias.n781 commonsourceibias.n780 161.3
R22396 commonsourceibias.n778 commonsourceibias.n752 161.3
R22397 commonsourceibias.n777 commonsourceibias.n776 161.3
R22398 commonsourceibias.n775 commonsourceibias.n753 161.3
R22399 commonsourceibias.n774 commonsourceibias.n773 161.3
R22400 commonsourceibias.n771 commonsourceibias.n754 161.3
R22401 commonsourceibias.n769 commonsourceibias.n768 161.3
R22402 commonsourceibias.n767 commonsourceibias.n755 161.3
R22403 commonsourceibias.n766 commonsourceibias.n765 161.3
R22404 commonsourceibias.n763 commonsourceibias.n756 161.3
R22405 commonsourceibias.n762 commonsourceibias.n761 161.3
R22406 commonsourceibias.n760 commonsourceibias.n757 161.3
R22407 commonsourceibias.n616 commonsourceibias.n504 161.3
R22408 commonsourceibias.n614 commonsourceibias.n613 161.3
R22409 commonsourceibias.n612 commonsourceibias.n505 161.3
R22410 commonsourceibias.n611 commonsourceibias.n610 161.3
R22411 commonsourceibias.n608 commonsourceibias.n506 161.3
R22412 commonsourceibias.n607 commonsourceibias.n606 161.3
R22413 commonsourceibias.n605 commonsourceibias.n507 161.3
R22414 commonsourceibias.n604 commonsourceibias.n603 161.3
R22415 commonsourceibias.n601 commonsourceibias.n508 161.3
R22416 commonsourceibias.n599 commonsourceibias.n598 161.3
R22417 commonsourceibias.n597 commonsourceibias.n509 161.3
R22418 commonsourceibias.n596 commonsourceibias.n595 161.3
R22419 commonsourceibias.n593 commonsourceibias.n510 161.3
R22420 commonsourceibias.n592 commonsourceibias.n591 161.3
R22421 commonsourceibias.n590 commonsourceibias.n511 161.3
R22422 commonsourceibias.n589 commonsourceibias.n588 161.3
R22423 commonsourceibias.n586 commonsourceibias.n512 161.3
R22424 commonsourceibias.n584 commonsourceibias.n583 161.3
R22425 commonsourceibias.n582 commonsourceibias.n513 161.3
R22426 commonsourceibias.n581 commonsourceibias.n580 161.3
R22427 commonsourceibias.n578 commonsourceibias.n514 161.3
R22428 commonsourceibias.n577 commonsourceibias.n576 161.3
R22429 commonsourceibias.n575 commonsourceibias.n515 161.3
R22430 commonsourceibias.n574 commonsourceibias.n573 161.3
R22431 commonsourceibias.n571 commonsourceibias.n516 161.3
R22432 commonsourceibias.n569 commonsourceibias.n568 161.3
R22433 commonsourceibias.n567 commonsourceibias.n517 161.3
R22434 commonsourceibias.n566 commonsourceibias.n565 161.3
R22435 commonsourceibias.n563 commonsourceibias.n518 161.3
R22436 commonsourceibias.n562 commonsourceibias.n561 161.3
R22437 commonsourceibias.n560 commonsourceibias.n519 161.3
R22438 commonsourceibias.n559 commonsourceibias.n558 161.3
R22439 commonsourceibias.n556 commonsourceibias.n520 161.3
R22440 commonsourceibias.n554 commonsourceibias.n553 161.3
R22441 commonsourceibias.n552 commonsourceibias.n521 161.3
R22442 commonsourceibias.n551 commonsourceibias.n550 161.3
R22443 commonsourceibias.n548 commonsourceibias.n522 161.3
R22444 commonsourceibias.n547 commonsourceibias.n546 161.3
R22445 commonsourceibias.n545 commonsourceibias.n523 161.3
R22446 commonsourceibias.n544 commonsourceibias.n543 161.3
R22447 commonsourceibias.n541 commonsourceibias.n524 161.3
R22448 commonsourceibias.n539 commonsourceibias.n538 161.3
R22449 commonsourceibias.n537 commonsourceibias.n525 161.3
R22450 commonsourceibias.n536 commonsourceibias.n535 161.3
R22451 commonsourceibias.n533 commonsourceibias.n526 161.3
R22452 commonsourceibias.n532 commonsourceibias.n531 161.3
R22453 commonsourceibias.n530 commonsourceibias.n527 161.3
R22454 commonsourceibias.n686 commonsourceibias.n685 161.3
R22455 commonsourceibias.n684 commonsourceibias.n683 161.3
R22456 commonsourceibias.n682 commonsourceibias.n632 161.3
R22457 commonsourceibias.n681 commonsourceibias.n680 161.3
R22458 commonsourceibias.n679 commonsourceibias.n678 161.3
R22459 commonsourceibias.n677 commonsourceibias.n634 161.3
R22460 commonsourceibias.n676 commonsourceibias.n675 161.3
R22461 commonsourceibias.n674 commonsourceibias.n673 161.3
R22462 commonsourceibias.n672 commonsourceibias.n636 161.3
R22463 commonsourceibias.n670 commonsourceibias.n669 161.3
R22464 commonsourceibias.n668 commonsourceibias.n637 161.3
R22465 commonsourceibias.n667 commonsourceibias.n666 161.3
R22466 commonsourceibias.n664 commonsourceibias.n638 161.3
R22467 commonsourceibias.n663 commonsourceibias.n662 161.3
R22468 commonsourceibias.n661 commonsourceibias.n639 161.3
R22469 commonsourceibias.n660 commonsourceibias.n659 161.3
R22470 commonsourceibias.n657 commonsourceibias.n640 161.3
R22471 commonsourceibias.n655 commonsourceibias.n654 161.3
R22472 commonsourceibias.n653 commonsourceibias.n641 161.3
R22473 commonsourceibias.n652 commonsourceibias.n651 161.3
R22474 commonsourceibias.n649 commonsourceibias.n642 161.3
R22475 commonsourceibias.n648 commonsourceibias.n647 161.3
R22476 commonsourceibias.n646 commonsourceibias.n643 161.3
R22477 commonsourceibias.n731 commonsourceibias.n483 161.3
R22478 commonsourceibias.n729 commonsourceibias.n728 161.3
R22479 commonsourceibias.n727 commonsourceibias.n484 161.3
R22480 commonsourceibias.n726 commonsourceibias.n725 161.3
R22481 commonsourceibias.n723 commonsourceibias.n485 161.3
R22482 commonsourceibias.n722 commonsourceibias.n721 161.3
R22483 commonsourceibias.n720 commonsourceibias.n486 161.3
R22484 commonsourceibias.n719 commonsourceibias.n718 161.3
R22485 commonsourceibias.n716 commonsourceibias.n487 161.3
R22486 commonsourceibias.n714 commonsourceibias.n713 161.3
R22487 commonsourceibias.n712 commonsourceibias.n488 161.3
R22488 commonsourceibias.n711 commonsourceibias.n710 161.3
R22489 commonsourceibias.n708 commonsourceibias.n489 161.3
R22490 commonsourceibias.n707 commonsourceibias.n706 161.3
R22491 commonsourceibias.n705 commonsourceibias.n490 161.3
R22492 commonsourceibias.n704 commonsourceibias.n703 161.3
R22493 commonsourceibias.n701 commonsourceibias.n491 161.3
R22494 commonsourceibias.n699 commonsourceibias.n698 161.3
R22495 commonsourceibias.n697 commonsourceibias.n492 161.3
R22496 commonsourceibias.n696 commonsourceibias.n695 161.3
R22497 commonsourceibias.n693 commonsourceibias.n493 161.3
R22498 commonsourceibias.n692 commonsourceibias.n691 161.3
R22499 commonsourceibias.n690 commonsourceibias.n494 161.3
R22500 commonsourceibias.n689 commonsourceibias.n688 161.3
R22501 commonsourceibias.n141 commonsourceibias.n139 81.5057
R22502 commonsourceibias.n497 commonsourceibias.n495 81.5057
R22503 commonsourceibias.n141 commonsourceibias.n140 80.9324
R22504 commonsourceibias.n143 commonsourceibias.n142 80.9324
R22505 commonsourceibias.n145 commonsourceibias.n144 80.9324
R22506 commonsourceibias.n147 commonsourceibias.n146 80.9324
R22507 commonsourceibias.n138 commonsourceibias.n137 80.9324
R22508 commonsourceibias.n136 commonsourceibias.n135 80.9324
R22509 commonsourceibias.n134 commonsourceibias.n133 80.9324
R22510 commonsourceibias.n132 commonsourceibias.n131 80.9324
R22511 commonsourceibias.n130 commonsourceibias.n129 80.9324
R22512 commonsourceibias.n620 commonsourceibias.n619 80.9324
R22513 commonsourceibias.n622 commonsourceibias.n621 80.9324
R22514 commonsourceibias.n624 commonsourceibias.n623 80.9324
R22515 commonsourceibias.n626 commonsourceibias.n625 80.9324
R22516 commonsourceibias.n628 commonsourceibias.n627 80.9324
R22517 commonsourceibias.n503 commonsourceibias.n502 80.9324
R22518 commonsourceibias.n501 commonsourceibias.n500 80.9324
R22519 commonsourceibias.n499 commonsourceibias.n498 80.9324
R22520 commonsourceibias.n497 commonsourceibias.n496 80.9324
R22521 commonsourceibias.n481 commonsourceibias.n480 80.6037
R22522 commonsourceibias.n365 commonsourceibias.n364 80.6037
R22523 commonsourceibias.n128 commonsourceibias.n127 80.6037
R22524 commonsourceibias.n250 commonsourceibias.n249 80.6037
R22525 commonsourceibias.n964 commonsourceibias.n963 80.6037
R22526 commonsourceibias.n848 commonsourceibias.n847 80.6037
R22527 commonsourceibias.n618 commonsourceibias.n617 80.6037
R22528 commonsourceibias.n733 commonsourceibias.n732 80.6037
R22529 commonsourceibias.n438 commonsourceibias.n437 56.5617
R22530 commonsourceibias.n452 commonsourceibias.n451 56.5617
R22531 commonsourceibias.n322 commonsourceibias.n321 56.5617
R22532 commonsourceibias.n308 commonsourceibias.n307 56.5617
R22533 commonsourceibias.n85 commonsourceibias.n84 56.5617
R22534 commonsourceibias.n71 commonsourceibias.n70 56.5617
R22535 commonsourceibias.n207 commonsourceibias.n206 56.5617
R22536 commonsourceibias.n193 commonsourceibias.n192 56.5617
R22537 commonsourceibias.n919 commonsourceibias.n917 56.5617
R22538 commonsourceibias.n934 commonsourceibias.n932 56.5617
R22539 commonsourceibias.n803 commonsourceibias.n801 56.5617
R22540 commonsourceibias.n818 commonsourceibias.n816 56.5617
R22541 commonsourceibias.n573 commonsourceibias.n571 56.5617
R22542 commonsourceibias.n588 commonsourceibias.n586 56.5617
R22543 commonsourceibias.n688 commonsourceibias.n686 56.5617
R22544 commonsourceibias.n410 commonsourceibias.n409 56.5617
R22545 commonsourceibias.n424 commonsourceibias.n423 56.5617
R22546 commonsourceibias.n466 commonsourceibias.n465 56.5617
R22547 commonsourceibias.n350 commonsourceibias.n349 56.5617
R22548 commonsourceibias.n336 commonsourceibias.n335 56.5617
R22549 commonsourceibias.n294 commonsourceibias.n293 56.5617
R22550 commonsourceibias.n113 commonsourceibias.n112 56.5617
R22551 commonsourceibias.n99 commonsourceibias.n98 56.5617
R22552 commonsourceibias.n57 commonsourceibias.n56 56.5617
R22553 commonsourceibias.n235 commonsourceibias.n234 56.5617
R22554 commonsourceibias.n221 commonsourceibias.n220 56.5617
R22555 commonsourceibias.n179 commonsourceibias.n178 56.5617
R22556 commonsourceibias.n889 commonsourceibias.n887 56.5617
R22557 commonsourceibias.n904 commonsourceibias.n902 56.5617
R22558 commonsourceibias.n949 commonsourceibias.n947 56.5617
R22559 commonsourceibias.n773 commonsourceibias.n771 56.5617
R22560 commonsourceibias.n788 commonsourceibias.n786 56.5617
R22561 commonsourceibias.n833 commonsourceibias.n831 56.5617
R22562 commonsourceibias.n543 commonsourceibias.n541 56.5617
R22563 commonsourceibias.n558 commonsourceibias.n556 56.5617
R22564 commonsourceibias.n603 commonsourceibias.n601 56.5617
R22565 commonsourceibias.n718 commonsourceibias.n716 56.5617
R22566 commonsourceibias.n703 commonsourceibias.n701 56.5617
R22567 commonsourceibias.n659 commonsourceibias.n657 56.5617
R22568 commonsourceibias.n673 commonsourceibias.n672 56.5617
R22569 commonsourceibias.n401 commonsourceibias.n400 51.2335
R22570 commonsourceibias.n473 commonsourceibias.n368 51.2335
R22571 commonsourceibias.n357 commonsourceibias.n252 51.2335
R22572 commonsourceibias.n285 commonsourceibias.n284 51.2335
R22573 commonsourceibias.n120 commonsourceibias.n15 51.2335
R22574 commonsourceibias.n48 commonsourceibias.n47 51.2335
R22575 commonsourceibias.n242 commonsourceibias.n1 51.2335
R22576 commonsourceibias.n170 commonsourceibias.n169 51.2335
R22577 commonsourceibias.n879 commonsourceibias.n878 51.2335
R22578 commonsourceibias.n956 commonsourceibias.n851 51.2335
R22579 commonsourceibias.n763 commonsourceibias.n762 51.2335
R22580 commonsourceibias.n840 commonsourceibias.n735 51.2335
R22581 commonsourceibias.n533 commonsourceibias.n532 51.2335
R22582 commonsourceibias.n610 commonsourceibias.n505 51.2335
R22583 commonsourceibias.n725 commonsourceibias.n484 51.2335
R22584 commonsourceibias.n649 commonsourceibias.n648 51.2335
R22585 commonsourceibias.n480 commonsourceibias.n479 50.9056
R22586 commonsourceibias.n364 commonsourceibias.n363 50.9056
R22587 commonsourceibias.n127 commonsourceibias.n126 50.9056
R22588 commonsourceibias.n249 commonsourceibias.n248 50.9056
R22589 commonsourceibias.n963 commonsourceibias.n962 50.9056
R22590 commonsourceibias.n847 commonsourceibias.n846 50.9056
R22591 commonsourceibias.n617 commonsourceibias.n616 50.9056
R22592 commonsourceibias.n732 commonsourceibias.n731 50.9056
R22593 commonsourceibias.n415 commonsourceibias.n414 50.2647
R22594 commonsourceibias.n459 commonsourceibias.n373 50.2647
R22595 commonsourceibias.n343 commonsourceibias.n257 50.2647
R22596 commonsourceibias.n299 commonsourceibias.n298 50.2647
R22597 commonsourceibias.n106 commonsourceibias.n20 50.2647
R22598 commonsourceibias.n62 commonsourceibias.n61 50.2647
R22599 commonsourceibias.n228 commonsourceibias.n6 50.2647
R22600 commonsourceibias.n184 commonsourceibias.n183 50.2647
R22601 commonsourceibias.n894 commonsourceibias.n893 50.2647
R22602 commonsourceibias.n941 commonsourceibias.n855 50.2647
R22603 commonsourceibias.n778 commonsourceibias.n777 50.2647
R22604 commonsourceibias.n825 commonsourceibias.n739 50.2647
R22605 commonsourceibias.n548 commonsourceibias.n547 50.2647
R22606 commonsourceibias.n595 commonsourceibias.n509 50.2647
R22607 commonsourceibias.n710 commonsourceibias.n488 50.2647
R22608 commonsourceibias.n664 commonsourceibias.n663 50.2647
R22609 commonsourceibias.n397 commonsourceibias.n396 49.9027
R22610 commonsourceibias.n281 commonsourceibias.n280 49.9027
R22611 commonsourceibias.n44 commonsourceibias.n43 49.9027
R22612 commonsourceibias.n166 commonsourceibias.n165 49.9027
R22613 commonsourceibias.n875 commonsourceibias.n874 49.9027
R22614 commonsourceibias.n759 commonsourceibias.n758 49.9027
R22615 commonsourceibias.n529 commonsourceibias.n528 49.9027
R22616 commonsourceibias.n645 commonsourceibias.n644 49.9027
R22617 commonsourceibias.n429 commonsourceibias.n428 49.296
R22618 commonsourceibias.n445 commonsourceibias.n378 49.296
R22619 commonsourceibias.n329 commonsourceibias.n262 49.296
R22620 commonsourceibias.n313 commonsourceibias.n312 49.296
R22621 commonsourceibias.n92 commonsourceibias.n25 49.296
R22622 commonsourceibias.n76 commonsourceibias.n75 49.296
R22623 commonsourceibias.n214 commonsourceibias.n11 49.296
R22624 commonsourceibias.n198 commonsourceibias.n197 49.296
R22625 commonsourceibias.n909 commonsourceibias.n908 49.296
R22626 commonsourceibias.n926 commonsourceibias.n859 49.296
R22627 commonsourceibias.n793 commonsourceibias.n792 49.296
R22628 commonsourceibias.n810 commonsourceibias.n743 49.296
R22629 commonsourceibias.n563 commonsourceibias.n562 49.296
R22630 commonsourceibias.n580 commonsourceibias.n513 49.296
R22631 commonsourceibias.n695 commonsourceibias.n492 49.296
R22632 commonsourceibias.n678 commonsourceibias.n677 49.296
R22633 commonsourceibias.n431 commonsourceibias.n383 48.3272
R22634 commonsourceibias.n443 commonsourceibias.n442 48.3272
R22635 commonsourceibias.n327 commonsourceibias.n326 48.3272
R22636 commonsourceibias.n315 commonsourceibias.n267 48.3272
R22637 commonsourceibias.n90 commonsourceibias.n89 48.3272
R22638 commonsourceibias.n78 commonsourceibias.n30 48.3272
R22639 commonsourceibias.n212 commonsourceibias.n211 48.3272
R22640 commonsourceibias.n202 commonsourceibias.n201 48.3272
R22641 commonsourceibias.n911 commonsourceibias.n863 48.3272
R22642 commonsourceibias.n924 commonsourceibias.n923 48.3272
R22643 commonsourceibias.n795 commonsourceibias.n747 48.3272
R22644 commonsourceibias.n808 commonsourceibias.n807 48.3272
R22645 commonsourceibias.n565 commonsourceibias.n517 48.3272
R22646 commonsourceibias.n578 commonsourceibias.n577 48.3272
R22647 commonsourceibias.n693 commonsourceibias.n692 48.3272
R22648 commonsourceibias.n682 commonsourceibias.n681 48.3272
R22649 commonsourceibias.n417 commonsourceibias.n388 47.3584
R22650 commonsourceibias.n457 commonsourceibias.n456 47.3584
R22651 commonsourceibias.n341 commonsourceibias.n340 47.3584
R22652 commonsourceibias.n301 commonsourceibias.n272 47.3584
R22653 commonsourceibias.n104 commonsourceibias.n103 47.3584
R22654 commonsourceibias.n64 commonsourceibias.n35 47.3584
R22655 commonsourceibias.n226 commonsourceibias.n225 47.3584
R22656 commonsourceibias.n186 commonsourceibias.n157 47.3584
R22657 commonsourceibias.n896 commonsourceibias.n867 47.3584
R22658 commonsourceibias.n939 commonsourceibias.n938 47.3584
R22659 commonsourceibias.n780 commonsourceibias.n751 47.3584
R22660 commonsourceibias.n823 commonsourceibias.n822 47.3584
R22661 commonsourceibias.n550 commonsourceibias.n521 47.3584
R22662 commonsourceibias.n593 commonsourceibias.n592 47.3584
R22663 commonsourceibias.n708 commonsourceibias.n707 47.3584
R22664 commonsourceibias.n666 commonsourceibias.n637 47.3584
R22665 commonsourceibias.n403 commonsourceibias.n393 46.3896
R22666 commonsourceibias.n471 commonsourceibias.n470 46.3896
R22667 commonsourceibias.n355 commonsourceibias.n354 46.3896
R22668 commonsourceibias.n287 commonsourceibias.n277 46.3896
R22669 commonsourceibias.n118 commonsourceibias.n117 46.3896
R22670 commonsourceibias.n50 commonsourceibias.n40 46.3896
R22671 commonsourceibias.n240 commonsourceibias.n239 46.3896
R22672 commonsourceibias.n172 commonsourceibias.n162 46.3896
R22673 commonsourceibias.n881 commonsourceibias.n871 46.3896
R22674 commonsourceibias.n954 commonsourceibias.n953 46.3896
R22675 commonsourceibias.n765 commonsourceibias.n755 46.3896
R22676 commonsourceibias.n838 commonsourceibias.n837 46.3896
R22677 commonsourceibias.n535 commonsourceibias.n525 46.3896
R22678 commonsourceibias.n608 commonsourceibias.n607 46.3896
R22679 commonsourceibias.n723 commonsourceibias.n722 46.3896
R22680 commonsourceibias.n651 commonsourceibias.n641 46.3896
R22681 commonsourceibias.n398 commonsourceibias.n397 44.7059
R22682 commonsourceibias.n876 commonsourceibias.n875 44.7059
R22683 commonsourceibias.n760 commonsourceibias.n759 44.7059
R22684 commonsourceibias.n530 commonsourceibias.n529 44.7059
R22685 commonsourceibias.n646 commonsourceibias.n645 44.7059
R22686 commonsourceibias.n282 commonsourceibias.n281 44.7059
R22687 commonsourceibias.n45 commonsourceibias.n44 44.7059
R22688 commonsourceibias.n167 commonsourceibias.n166 44.7059
R22689 commonsourceibias.n407 commonsourceibias.n393 34.7644
R22690 commonsourceibias.n470 commonsourceibias.n370 34.7644
R22691 commonsourceibias.n354 commonsourceibias.n254 34.7644
R22692 commonsourceibias.n291 commonsourceibias.n277 34.7644
R22693 commonsourceibias.n117 commonsourceibias.n17 34.7644
R22694 commonsourceibias.n54 commonsourceibias.n40 34.7644
R22695 commonsourceibias.n239 commonsourceibias.n3 34.7644
R22696 commonsourceibias.n176 commonsourceibias.n162 34.7644
R22697 commonsourceibias.n885 commonsourceibias.n871 34.7644
R22698 commonsourceibias.n953 commonsourceibias.n853 34.7644
R22699 commonsourceibias.n769 commonsourceibias.n755 34.7644
R22700 commonsourceibias.n837 commonsourceibias.n737 34.7644
R22701 commonsourceibias.n539 commonsourceibias.n525 34.7644
R22702 commonsourceibias.n607 commonsourceibias.n507 34.7644
R22703 commonsourceibias.n722 commonsourceibias.n486 34.7644
R22704 commonsourceibias.n655 commonsourceibias.n641 34.7644
R22705 commonsourceibias.n421 commonsourceibias.n388 33.7956
R22706 commonsourceibias.n456 commonsourceibias.n375 33.7956
R22707 commonsourceibias.n340 commonsourceibias.n259 33.7956
R22708 commonsourceibias.n305 commonsourceibias.n272 33.7956
R22709 commonsourceibias.n103 commonsourceibias.n22 33.7956
R22710 commonsourceibias.n68 commonsourceibias.n35 33.7956
R22711 commonsourceibias.n225 commonsourceibias.n8 33.7956
R22712 commonsourceibias.n190 commonsourceibias.n157 33.7956
R22713 commonsourceibias.n900 commonsourceibias.n867 33.7956
R22714 commonsourceibias.n938 commonsourceibias.n857 33.7956
R22715 commonsourceibias.n784 commonsourceibias.n751 33.7956
R22716 commonsourceibias.n822 commonsourceibias.n741 33.7956
R22717 commonsourceibias.n554 commonsourceibias.n521 33.7956
R22718 commonsourceibias.n592 commonsourceibias.n511 33.7956
R22719 commonsourceibias.n707 commonsourceibias.n490 33.7956
R22720 commonsourceibias.n670 commonsourceibias.n637 33.7956
R22721 commonsourceibias.n435 commonsourceibias.n383 32.8269
R22722 commonsourceibias.n442 commonsourceibias.n380 32.8269
R22723 commonsourceibias.n326 commonsourceibias.n264 32.8269
R22724 commonsourceibias.n319 commonsourceibias.n267 32.8269
R22725 commonsourceibias.n89 commonsourceibias.n27 32.8269
R22726 commonsourceibias.n82 commonsourceibias.n30 32.8269
R22727 commonsourceibias.n211 commonsourceibias.n13 32.8269
R22728 commonsourceibias.n203 commonsourceibias.n202 32.8269
R22729 commonsourceibias.n915 commonsourceibias.n863 32.8269
R22730 commonsourceibias.n923 commonsourceibias.n861 32.8269
R22731 commonsourceibias.n799 commonsourceibias.n747 32.8269
R22732 commonsourceibias.n807 commonsourceibias.n745 32.8269
R22733 commonsourceibias.n569 commonsourceibias.n517 32.8269
R22734 commonsourceibias.n577 commonsourceibias.n515 32.8269
R22735 commonsourceibias.n692 commonsourceibias.n494 32.8269
R22736 commonsourceibias.n683 commonsourceibias.n682 32.8269
R22737 commonsourceibias.n428 commonsourceibias.n385 31.8581
R22738 commonsourceibias.n449 commonsourceibias.n378 31.8581
R22739 commonsourceibias.n333 commonsourceibias.n262 31.8581
R22740 commonsourceibias.n312 commonsourceibias.n269 31.8581
R22741 commonsourceibias.n96 commonsourceibias.n25 31.8581
R22742 commonsourceibias.n75 commonsourceibias.n32 31.8581
R22743 commonsourceibias.n218 commonsourceibias.n11 31.8581
R22744 commonsourceibias.n197 commonsourceibias.n196 31.8581
R22745 commonsourceibias.n908 commonsourceibias.n865 31.8581
R22746 commonsourceibias.n930 commonsourceibias.n859 31.8581
R22747 commonsourceibias.n792 commonsourceibias.n749 31.8581
R22748 commonsourceibias.n814 commonsourceibias.n743 31.8581
R22749 commonsourceibias.n562 commonsourceibias.n519 31.8581
R22750 commonsourceibias.n584 commonsourceibias.n513 31.8581
R22751 commonsourceibias.n699 commonsourceibias.n492 31.8581
R22752 commonsourceibias.n677 commonsourceibias.n676 31.8581
R22753 commonsourceibias.n414 commonsourceibias.n390 30.8893
R22754 commonsourceibias.n463 commonsourceibias.n373 30.8893
R22755 commonsourceibias.n347 commonsourceibias.n257 30.8893
R22756 commonsourceibias.n298 commonsourceibias.n274 30.8893
R22757 commonsourceibias.n110 commonsourceibias.n20 30.8893
R22758 commonsourceibias.n61 commonsourceibias.n37 30.8893
R22759 commonsourceibias.n232 commonsourceibias.n6 30.8893
R22760 commonsourceibias.n183 commonsourceibias.n159 30.8893
R22761 commonsourceibias.n893 commonsourceibias.n869 30.8893
R22762 commonsourceibias.n945 commonsourceibias.n855 30.8893
R22763 commonsourceibias.n777 commonsourceibias.n753 30.8893
R22764 commonsourceibias.n829 commonsourceibias.n739 30.8893
R22765 commonsourceibias.n547 commonsourceibias.n523 30.8893
R22766 commonsourceibias.n599 commonsourceibias.n509 30.8893
R22767 commonsourceibias.n714 commonsourceibias.n488 30.8893
R22768 commonsourceibias.n663 commonsourceibias.n639 30.8893
R22769 commonsourceibias.n400 commonsourceibias.n395 29.9206
R22770 commonsourceibias.n477 commonsourceibias.n368 29.9206
R22771 commonsourceibias.n361 commonsourceibias.n252 29.9206
R22772 commonsourceibias.n284 commonsourceibias.n279 29.9206
R22773 commonsourceibias.n124 commonsourceibias.n15 29.9206
R22774 commonsourceibias.n47 commonsourceibias.n42 29.9206
R22775 commonsourceibias.n246 commonsourceibias.n1 29.9206
R22776 commonsourceibias.n169 commonsourceibias.n164 29.9206
R22777 commonsourceibias.n878 commonsourceibias.n873 29.9206
R22778 commonsourceibias.n960 commonsourceibias.n851 29.9206
R22779 commonsourceibias.n762 commonsourceibias.n757 29.9206
R22780 commonsourceibias.n844 commonsourceibias.n735 29.9206
R22781 commonsourceibias.n532 commonsourceibias.n527 29.9206
R22782 commonsourceibias.n614 commonsourceibias.n505 29.9206
R22783 commonsourceibias.n729 commonsourceibias.n484 29.9206
R22784 commonsourceibias.n648 commonsourceibias.n643 29.9206
R22785 commonsourceibias.n479 commonsourceibias.n478 21.8872
R22786 commonsourceibias.n363 commonsourceibias.n362 21.8872
R22787 commonsourceibias.n126 commonsourceibias.n125 21.8872
R22788 commonsourceibias.n248 commonsourceibias.n247 21.8872
R22789 commonsourceibias.n962 commonsourceibias.n961 21.8872
R22790 commonsourceibias.n846 commonsourceibias.n845 21.8872
R22791 commonsourceibias.n616 commonsourceibias.n615 21.8872
R22792 commonsourceibias.n731 commonsourceibias.n730 21.8872
R22793 commonsourceibias.n410 commonsourceibias.n392 21.3954
R22794 commonsourceibias.n465 commonsourceibias.n464 21.3954
R22795 commonsourceibias.n349 commonsourceibias.n348 21.3954
R22796 commonsourceibias.n294 commonsourceibias.n276 21.3954
R22797 commonsourceibias.n112 commonsourceibias.n111 21.3954
R22798 commonsourceibias.n57 commonsourceibias.n39 21.3954
R22799 commonsourceibias.n234 commonsourceibias.n233 21.3954
R22800 commonsourceibias.n179 commonsourceibias.n161 21.3954
R22801 commonsourceibias.n889 commonsourceibias.n888 21.3954
R22802 commonsourceibias.n947 commonsourceibias.n946 21.3954
R22803 commonsourceibias.n773 commonsourceibias.n772 21.3954
R22804 commonsourceibias.n831 commonsourceibias.n830 21.3954
R22805 commonsourceibias.n543 commonsourceibias.n542 21.3954
R22806 commonsourceibias.n601 commonsourceibias.n600 21.3954
R22807 commonsourceibias.n716 commonsourceibias.n715 21.3954
R22808 commonsourceibias.n659 commonsourceibias.n658 21.3954
R22809 commonsourceibias.n424 commonsourceibias.n387 20.9036
R22810 commonsourceibias.n451 commonsourceibias.n450 20.9036
R22811 commonsourceibias.n335 commonsourceibias.n334 20.9036
R22812 commonsourceibias.n308 commonsourceibias.n271 20.9036
R22813 commonsourceibias.n98 commonsourceibias.n97 20.9036
R22814 commonsourceibias.n71 commonsourceibias.n34 20.9036
R22815 commonsourceibias.n220 commonsourceibias.n219 20.9036
R22816 commonsourceibias.n193 commonsourceibias.n155 20.9036
R22817 commonsourceibias.n904 commonsourceibias.n903 20.9036
R22818 commonsourceibias.n932 commonsourceibias.n931 20.9036
R22819 commonsourceibias.n788 commonsourceibias.n787 20.9036
R22820 commonsourceibias.n816 commonsourceibias.n815 20.9036
R22821 commonsourceibias.n558 commonsourceibias.n557 20.9036
R22822 commonsourceibias.n586 commonsourceibias.n585 20.9036
R22823 commonsourceibias.n701 commonsourceibias.n700 20.9036
R22824 commonsourceibias.n673 commonsourceibias.n635 20.9036
R22825 commonsourceibias.n437 commonsourceibias.n436 20.4117
R22826 commonsourceibias.n438 commonsourceibias.n382 20.4117
R22827 commonsourceibias.n322 commonsourceibias.n266 20.4117
R22828 commonsourceibias.n321 commonsourceibias.n320 20.4117
R22829 commonsourceibias.n85 commonsourceibias.n29 20.4117
R22830 commonsourceibias.n84 commonsourceibias.n83 20.4117
R22831 commonsourceibias.n207 commonsourceibias.n150 20.4117
R22832 commonsourceibias.n206 commonsourceibias.n151 20.4117
R22833 commonsourceibias.n917 commonsourceibias.n916 20.4117
R22834 commonsourceibias.n919 commonsourceibias.n918 20.4117
R22835 commonsourceibias.n801 commonsourceibias.n800 20.4117
R22836 commonsourceibias.n803 commonsourceibias.n802 20.4117
R22837 commonsourceibias.n571 commonsourceibias.n570 20.4117
R22838 commonsourceibias.n573 commonsourceibias.n572 20.4117
R22839 commonsourceibias.n688 commonsourceibias.n687 20.4117
R22840 commonsourceibias.n686 commonsourceibias.n631 20.4117
R22841 commonsourceibias.n423 commonsourceibias.n422 19.9199
R22842 commonsourceibias.n452 commonsourceibias.n377 19.9199
R22843 commonsourceibias.n336 commonsourceibias.n261 19.9199
R22844 commonsourceibias.n307 commonsourceibias.n306 19.9199
R22845 commonsourceibias.n99 commonsourceibias.n24 19.9199
R22846 commonsourceibias.n70 commonsourceibias.n69 19.9199
R22847 commonsourceibias.n221 commonsourceibias.n10 19.9199
R22848 commonsourceibias.n192 commonsourceibias.n191 19.9199
R22849 commonsourceibias.n902 commonsourceibias.n901 19.9199
R22850 commonsourceibias.n934 commonsourceibias.n933 19.9199
R22851 commonsourceibias.n786 commonsourceibias.n785 19.9199
R22852 commonsourceibias.n818 commonsourceibias.n817 19.9199
R22853 commonsourceibias.n556 commonsourceibias.n555 19.9199
R22854 commonsourceibias.n588 commonsourceibias.n587 19.9199
R22855 commonsourceibias.n703 commonsourceibias.n702 19.9199
R22856 commonsourceibias.n672 commonsourceibias.n671 19.9199
R22857 commonsourceibias.n409 commonsourceibias.n408 19.4281
R22858 commonsourceibias.n466 commonsourceibias.n372 19.4281
R22859 commonsourceibias.n350 commonsourceibias.n256 19.4281
R22860 commonsourceibias.n293 commonsourceibias.n292 19.4281
R22861 commonsourceibias.n113 commonsourceibias.n19 19.4281
R22862 commonsourceibias.n56 commonsourceibias.n55 19.4281
R22863 commonsourceibias.n235 commonsourceibias.n5 19.4281
R22864 commonsourceibias.n178 commonsourceibias.n177 19.4281
R22865 commonsourceibias.n887 commonsourceibias.n886 19.4281
R22866 commonsourceibias.n949 commonsourceibias.n948 19.4281
R22867 commonsourceibias.n771 commonsourceibias.n770 19.4281
R22868 commonsourceibias.n833 commonsourceibias.n832 19.4281
R22869 commonsourceibias.n541 commonsourceibias.n540 19.4281
R22870 commonsourceibias.n603 commonsourceibias.n602 19.4281
R22871 commonsourceibias.n718 commonsourceibias.n717 19.4281
R22872 commonsourceibias.n657 commonsourceibias.n656 19.4281
R22873 commonsourceibias.n402 commonsourceibias.n401 13.526
R22874 commonsourceibias.n473 commonsourceibias.n472 13.526
R22875 commonsourceibias.n357 commonsourceibias.n356 13.526
R22876 commonsourceibias.n286 commonsourceibias.n285 13.526
R22877 commonsourceibias.n120 commonsourceibias.n119 13.526
R22878 commonsourceibias.n49 commonsourceibias.n48 13.526
R22879 commonsourceibias.n242 commonsourceibias.n241 13.526
R22880 commonsourceibias.n171 commonsourceibias.n170 13.526
R22881 commonsourceibias.n880 commonsourceibias.n879 13.526
R22882 commonsourceibias.n956 commonsourceibias.n955 13.526
R22883 commonsourceibias.n764 commonsourceibias.n763 13.526
R22884 commonsourceibias.n840 commonsourceibias.n839 13.526
R22885 commonsourceibias.n534 commonsourceibias.n533 13.526
R22886 commonsourceibias.n610 commonsourceibias.n609 13.526
R22887 commonsourceibias.n725 commonsourceibias.n724 13.526
R22888 commonsourceibias.n650 commonsourceibias.n649 13.526
R22889 commonsourceibias.n130 commonsourceibias.n128 13.2322
R22890 commonsourceibias.n620 commonsourceibias.n618 13.2322
R22891 commonsourceibias.n416 commonsourceibias.n415 13.0342
R22892 commonsourceibias.n459 commonsourceibias.n458 13.0342
R22893 commonsourceibias.n343 commonsourceibias.n342 13.0342
R22894 commonsourceibias.n300 commonsourceibias.n299 13.0342
R22895 commonsourceibias.n106 commonsourceibias.n105 13.0342
R22896 commonsourceibias.n63 commonsourceibias.n62 13.0342
R22897 commonsourceibias.n228 commonsourceibias.n227 13.0342
R22898 commonsourceibias.n185 commonsourceibias.n184 13.0342
R22899 commonsourceibias.n895 commonsourceibias.n894 13.0342
R22900 commonsourceibias.n941 commonsourceibias.n940 13.0342
R22901 commonsourceibias.n779 commonsourceibias.n778 13.0342
R22902 commonsourceibias.n825 commonsourceibias.n824 13.0342
R22903 commonsourceibias.n549 commonsourceibias.n548 13.0342
R22904 commonsourceibias.n595 commonsourceibias.n594 13.0342
R22905 commonsourceibias.n710 commonsourceibias.n709 13.0342
R22906 commonsourceibias.n665 commonsourceibias.n664 13.0342
R22907 commonsourceibias.n430 commonsourceibias.n429 12.5423
R22908 commonsourceibias.n445 commonsourceibias.n444 12.5423
R22909 commonsourceibias.n329 commonsourceibias.n328 12.5423
R22910 commonsourceibias.n314 commonsourceibias.n313 12.5423
R22911 commonsourceibias.n92 commonsourceibias.n91 12.5423
R22912 commonsourceibias.n77 commonsourceibias.n76 12.5423
R22913 commonsourceibias.n214 commonsourceibias.n213 12.5423
R22914 commonsourceibias.n198 commonsourceibias.n153 12.5423
R22915 commonsourceibias.n910 commonsourceibias.n909 12.5423
R22916 commonsourceibias.n926 commonsourceibias.n925 12.5423
R22917 commonsourceibias.n794 commonsourceibias.n793 12.5423
R22918 commonsourceibias.n810 commonsourceibias.n809 12.5423
R22919 commonsourceibias.n564 commonsourceibias.n563 12.5423
R22920 commonsourceibias.n580 commonsourceibias.n579 12.5423
R22921 commonsourceibias.n695 commonsourceibias.n694 12.5423
R22922 commonsourceibias.n678 commonsourceibias.n633 12.5423
R22923 commonsourceibias.n431 commonsourceibias.n430 12.0505
R22924 commonsourceibias.n444 commonsourceibias.n443 12.0505
R22925 commonsourceibias.n328 commonsourceibias.n327 12.0505
R22926 commonsourceibias.n315 commonsourceibias.n314 12.0505
R22927 commonsourceibias.n91 commonsourceibias.n90 12.0505
R22928 commonsourceibias.n78 commonsourceibias.n77 12.0505
R22929 commonsourceibias.n213 commonsourceibias.n212 12.0505
R22930 commonsourceibias.n201 commonsourceibias.n153 12.0505
R22931 commonsourceibias.n911 commonsourceibias.n910 12.0505
R22932 commonsourceibias.n925 commonsourceibias.n924 12.0505
R22933 commonsourceibias.n795 commonsourceibias.n794 12.0505
R22934 commonsourceibias.n809 commonsourceibias.n808 12.0505
R22935 commonsourceibias.n565 commonsourceibias.n564 12.0505
R22936 commonsourceibias.n579 commonsourceibias.n578 12.0505
R22937 commonsourceibias.n694 commonsourceibias.n693 12.0505
R22938 commonsourceibias.n681 commonsourceibias.n633 12.0505
R22939 commonsourceibias.n417 commonsourceibias.n416 11.5587
R22940 commonsourceibias.n458 commonsourceibias.n457 11.5587
R22941 commonsourceibias.n342 commonsourceibias.n341 11.5587
R22942 commonsourceibias.n301 commonsourceibias.n300 11.5587
R22943 commonsourceibias.n105 commonsourceibias.n104 11.5587
R22944 commonsourceibias.n64 commonsourceibias.n63 11.5587
R22945 commonsourceibias.n227 commonsourceibias.n226 11.5587
R22946 commonsourceibias.n186 commonsourceibias.n185 11.5587
R22947 commonsourceibias.n896 commonsourceibias.n895 11.5587
R22948 commonsourceibias.n940 commonsourceibias.n939 11.5587
R22949 commonsourceibias.n780 commonsourceibias.n779 11.5587
R22950 commonsourceibias.n824 commonsourceibias.n823 11.5587
R22951 commonsourceibias.n550 commonsourceibias.n549 11.5587
R22952 commonsourceibias.n594 commonsourceibias.n593 11.5587
R22953 commonsourceibias.n709 commonsourceibias.n708 11.5587
R22954 commonsourceibias.n666 commonsourceibias.n665 11.5587
R22955 commonsourceibias.n403 commonsourceibias.n402 11.0668
R22956 commonsourceibias.n472 commonsourceibias.n471 11.0668
R22957 commonsourceibias.n356 commonsourceibias.n355 11.0668
R22958 commonsourceibias.n287 commonsourceibias.n286 11.0668
R22959 commonsourceibias.n119 commonsourceibias.n118 11.0668
R22960 commonsourceibias.n50 commonsourceibias.n49 11.0668
R22961 commonsourceibias.n241 commonsourceibias.n240 11.0668
R22962 commonsourceibias.n172 commonsourceibias.n171 11.0668
R22963 commonsourceibias.n881 commonsourceibias.n880 11.0668
R22964 commonsourceibias.n955 commonsourceibias.n954 11.0668
R22965 commonsourceibias.n765 commonsourceibias.n764 11.0668
R22966 commonsourceibias.n839 commonsourceibias.n838 11.0668
R22967 commonsourceibias.n535 commonsourceibias.n534 11.0668
R22968 commonsourceibias.n609 commonsourceibias.n608 11.0668
R22969 commonsourceibias.n724 commonsourceibias.n723 11.0668
R22970 commonsourceibias.n651 commonsourceibias.n650 11.0668
R22971 commonsourceibias.n966 commonsourceibias.n482 10.122
R22972 commonsourceibias.n149 commonsourceibias.n148 9.50363
R22973 commonsourceibias.n630 commonsourceibias.n629 9.50363
R22974 commonsourceibias.n366 commonsourceibias.n250 8.76042
R22975 commonsourceibias.n849 commonsourceibias.n733 8.76042
R22976 commonsourceibias.n966 commonsourceibias.n965 8.46921
R22977 commonsourceibias.n408 commonsourceibias.n407 5.16479
R22978 commonsourceibias.n372 commonsourceibias.n370 5.16479
R22979 commonsourceibias.n256 commonsourceibias.n254 5.16479
R22980 commonsourceibias.n292 commonsourceibias.n291 5.16479
R22981 commonsourceibias.n19 commonsourceibias.n17 5.16479
R22982 commonsourceibias.n55 commonsourceibias.n54 5.16479
R22983 commonsourceibias.n5 commonsourceibias.n3 5.16479
R22984 commonsourceibias.n177 commonsourceibias.n176 5.16479
R22985 commonsourceibias.n886 commonsourceibias.n885 5.16479
R22986 commonsourceibias.n948 commonsourceibias.n853 5.16479
R22987 commonsourceibias.n770 commonsourceibias.n769 5.16479
R22988 commonsourceibias.n832 commonsourceibias.n737 5.16479
R22989 commonsourceibias.n540 commonsourceibias.n539 5.16479
R22990 commonsourceibias.n602 commonsourceibias.n507 5.16479
R22991 commonsourceibias.n717 commonsourceibias.n486 5.16479
R22992 commonsourceibias.n656 commonsourceibias.n655 5.16479
R22993 commonsourceibias.n482 commonsourceibias.n481 5.03125
R22994 commonsourceibias.n366 commonsourceibias.n365 5.03125
R22995 commonsourceibias.n965 commonsourceibias.n964 5.03125
R22996 commonsourceibias.n849 commonsourceibias.n848 5.03125
R22997 commonsourceibias.n422 commonsourceibias.n421 4.67295
R22998 commonsourceibias.n377 commonsourceibias.n375 4.67295
R22999 commonsourceibias.n261 commonsourceibias.n259 4.67295
R23000 commonsourceibias.n306 commonsourceibias.n305 4.67295
R23001 commonsourceibias.n24 commonsourceibias.n22 4.67295
R23002 commonsourceibias.n69 commonsourceibias.n68 4.67295
R23003 commonsourceibias.n10 commonsourceibias.n8 4.67295
R23004 commonsourceibias.n191 commonsourceibias.n190 4.67295
R23005 commonsourceibias.n901 commonsourceibias.n900 4.67295
R23006 commonsourceibias.n933 commonsourceibias.n857 4.67295
R23007 commonsourceibias.n785 commonsourceibias.n784 4.67295
R23008 commonsourceibias.n817 commonsourceibias.n741 4.67295
R23009 commonsourceibias.n555 commonsourceibias.n554 4.67295
R23010 commonsourceibias.n587 commonsourceibias.n511 4.67295
R23011 commonsourceibias.n702 commonsourceibias.n490 4.67295
R23012 commonsourceibias.n671 commonsourceibias.n670 4.67295
R23013 commonsourceibias commonsourceibias.n966 4.20978
R23014 commonsourceibias.n436 commonsourceibias.n435 4.18111
R23015 commonsourceibias.n382 commonsourceibias.n380 4.18111
R23016 commonsourceibias.n266 commonsourceibias.n264 4.18111
R23017 commonsourceibias.n320 commonsourceibias.n319 4.18111
R23018 commonsourceibias.n29 commonsourceibias.n27 4.18111
R23019 commonsourceibias.n83 commonsourceibias.n82 4.18111
R23020 commonsourceibias.n150 commonsourceibias.n13 4.18111
R23021 commonsourceibias.n203 commonsourceibias.n151 4.18111
R23022 commonsourceibias.n916 commonsourceibias.n915 4.18111
R23023 commonsourceibias.n918 commonsourceibias.n861 4.18111
R23024 commonsourceibias.n800 commonsourceibias.n799 4.18111
R23025 commonsourceibias.n802 commonsourceibias.n745 4.18111
R23026 commonsourceibias.n570 commonsourceibias.n569 4.18111
R23027 commonsourceibias.n572 commonsourceibias.n515 4.18111
R23028 commonsourceibias.n687 commonsourceibias.n494 4.18111
R23029 commonsourceibias.n683 commonsourceibias.n631 4.18111
R23030 commonsourceibias.n482 commonsourceibias.n366 3.72967
R23031 commonsourceibias.n965 commonsourceibias.n849 3.72967
R23032 commonsourceibias.n387 commonsourceibias.n385 3.68928
R23033 commonsourceibias.n450 commonsourceibias.n449 3.68928
R23034 commonsourceibias.n334 commonsourceibias.n333 3.68928
R23035 commonsourceibias.n271 commonsourceibias.n269 3.68928
R23036 commonsourceibias.n97 commonsourceibias.n96 3.68928
R23037 commonsourceibias.n34 commonsourceibias.n32 3.68928
R23038 commonsourceibias.n219 commonsourceibias.n218 3.68928
R23039 commonsourceibias.n196 commonsourceibias.n155 3.68928
R23040 commonsourceibias.n903 commonsourceibias.n865 3.68928
R23041 commonsourceibias.n931 commonsourceibias.n930 3.68928
R23042 commonsourceibias.n787 commonsourceibias.n749 3.68928
R23043 commonsourceibias.n815 commonsourceibias.n814 3.68928
R23044 commonsourceibias.n557 commonsourceibias.n519 3.68928
R23045 commonsourceibias.n585 commonsourceibias.n584 3.68928
R23046 commonsourceibias.n700 commonsourceibias.n699 3.68928
R23047 commonsourceibias.n676 commonsourceibias.n635 3.68928
R23048 commonsourceibias.n392 commonsourceibias.n390 3.19744
R23049 commonsourceibias.n464 commonsourceibias.n463 3.19744
R23050 commonsourceibias.n348 commonsourceibias.n347 3.19744
R23051 commonsourceibias.n276 commonsourceibias.n274 3.19744
R23052 commonsourceibias.n111 commonsourceibias.n110 3.19744
R23053 commonsourceibias.n39 commonsourceibias.n37 3.19744
R23054 commonsourceibias.n233 commonsourceibias.n232 3.19744
R23055 commonsourceibias.n161 commonsourceibias.n159 3.19744
R23056 commonsourceibias.n888 commonsourceibias.n869 3.19744
R23057 commonsourceibias.n946 commonsourceibias.n945 3.19744
R23058 commonsourceibias.n772 commonsourceibias.n753 3.19744
R23059 commonsourceibias.n830 commonsourceibias.n829 3.19744
R23060 commonsourceibias.n542 commonsourceibias.n523 3.19744
R23061 commonsourceibias.n600 commonsourceibias.n599 3.19744
R23062 commonsourceibias.n715 commonsourceibias.n714 3.19744
R23063 commonsourceibias.n658 commonsourceibias.n639 3.19744
R23064 commonsourceibias.n139 commonsourceibias.t59 2.82907
R23065 commonsourceibias.n139 commonsourceibias.t27 2.82907
R23066 commonsourceibias.n140 commonsourceibias.t43 2.82907
R23067 commonsourceibias.n140 commonsourceibias.t53 2.82907
R23068 commonsourceibias.n142 commonsourceibias.t63 2.82907
R23069 commonsourceibias.n142 commonsourceibias.t1 2.82907
R23070 commonsourceibias.n144 commonsourceibias.t71 2.82907
R23071 commonsourceibias.n144 commonsourceibias.t23 2.82907
R23072 commonsourceibias.n146 commonsourceibias.t31 2.82907
R23073 commonsourceibias.n146 commonsourceibias.t37 2.82907
R23074 commonsourceibias.n137 commonsourceibias.t19 2.82907
R23075 commonsourceibias.n137 commonsourceibias.t55 2.82907
R23076 commonsourceibias.n135 commonsourceibias.t35 2.82907
R23077 commonsourceibias.n135 commonsourceibias.t11 2.82907
R23078 commonsourceibias.n133 commonsourceibias.t75 2.82907
R23079 commonsourceibias.n133 commonsourceibias.t21 2.82907
R23080 commonsourceibias.n131 commonsourceibias.t5 2.82907
R23081 commonsourceibias.n131 commonsourceibias.t15 2.82907
R23082 commonsourceibias.n129 commonsourceibias.t17 2.82907
R23083 commonsourceibias.n129 commonsourceibias.t61 2.82907
R23084 commonsourceibias.n619 commonsourceibias.t77 2.82907
R23085 commonsourceibias.n619 commonsourceibias.t41 2.82907
R23086 commonsourceibias.n621 commonsourceibias.t39 2.82907
R23087 commonsourceibias.n621 commonsourceibias.t25 2.82907
R23088 commonsourceibias.n623 commonsourceibias.t47 2.82907
R23089 commonsourceibias.n623 commonsourceibias.t13 2.82907
R23090 commonsourceibias.n625 commonsourceibias.t33 2.82907
R23091 commonsourceibias.n625 commonsourceibias.t57 2.82907
R23092 commonsourceibias.n627 commonsourceibias.t73 2.82907
R23093 commonsourceibias.n627 commonsourceibias.t45 2.82907
R23094 commonsourceibias.n502 commonsourceibias.t65 2.82907
R23095 commonsourceibias.n502 commonsourceibias.t51 2.82907
R23096 commonsourceibias.n500 commonsourceibias.t49 2.82907
R23097 commonsourceibias.n500 commonsourceibias.t3 2.82907
R23098 commonsourceibias.n498 commonsourceibias.t29 2.82907
R23099 commonsourceibias.n498 commonsourceibias.t79 2.82907
R23100 commonsourceibias.n496 commonsourceibias.t7 2.82907
R23101 commonsourceibias.n496 commonsourceibias.t67 2.82907
R23102 commonsourceibias.n495 commonsourceibias.t69 2.82907
R23103 commonsourceibias.n495 commonsourceibias.t9 2.82907
R23104 commonsourceibias.n396 commonsourceibias.n395 2.7056
R23105 commonsourceibias.n478 commonsourceibias.n477 2.7056
R23106 commonsourceibias.n362 commonsourceibias.n361 2.7056
R23107 commonsourceibias.n280 commonsourceibias.n279 2.7056
R23108 commonsourceibias.n125 commonsourceibias.n124 2.7056
R23109 commonsourceibias.n43 commonsourceibias.n42 2.7056
R23110 commonsourceibias.n247 commonsourceibias.n246 2.7056
R23111 commonsourceibias.n165 commonsourceibias.n164 2.7056
R23112 commonsourceibias.n874 commonsourceibias.n873 2.7056
R23113 commonsourceibias.n961 commonsourceibias.n960 2.7056
R23114 commonsourceibias.n758 commonsourceibias.n757 2.7056
R23115 commonsourceibias.n845 commonsourceibias.n844 2.7056
R23116 commonsourceibias.n528 commonsourceibias.n527 2.7056
R23117 commonsourceibias.n615 commonsourceibias.n614 2.7056
R23118 commonsourceibias.n730 commonsourceibias.n729 2.7056
R23119 commonsourceibias.n644 commonsourceibias.n643 2.7056
R23120 commonsourceibias.n132 commonsourceibias.n130 0.573776
R23121 commonsourceibias.n134 commonsourceibias.n132 0.573776
R23122 commonsourceibias.n136 commonsourceibias.n134 0.573776
R23123 commonsourceibias.n138 commonsourceibias.n136 0.573776
R23124 commonsourceibias.n147 commonsourceibias.n145 0.573776
R23125 commonsourceibias.n145 commonsourceibias.n143 0.573776
R23126 commonsourceibias.n143 commonsourceibias.n141 0.573776
R23127 commonsourceibias.n499 commonsourceibias.n497 0.573776
R23128 commonsourceibias.n501 commonsourceibias.n499 0.573776
R23129 commonsourceibias.n503 commonsourceibias.n501 0.573776
R23130 commonsourceibias.n628 commonsourceibias.n626 0.573776
R23131 commonsourceibias.n626 commonsourceibias.n624 0.573776
R23132 commonsourceibias.n624 commonsourceibias.n622 0.573776
R23133 commonsourceibias.n622 commonsourceibias.n620 0.573776
R23134 commonsourceibias.n148 commonsourceibias.n138 0.287138
R23135 commonsourceibias.n148 commonsourceibias.n147 0.287138
R23136 commonsourceibias.n629 commonsourceibias.n503 0.287138
R23137 commonsourceibias.n629 commonsourceibias.n628 0.287138
R23138 commonsourceibias.n481 commonsourceibias.n367 0.285035
R23139 commonsourceibias.n365 commonsourceibias.n251 0.285035
R23140 commonsourceibias.n128 commonsourceibias.n14 0.285035
R23141 commonsourceibias.n250 commonsourceibias.n0 0.285035
R23142 commonsourceibias.n964 commonsourceibias.n850 0.285035
R23143 commonsourceibias.n848 commonsourceibias.n734 0.285035
R23144 commonsourceibias.n618 commonsourceibias.n504 0.285035
R23145 commonsourceibias.n733 commonsourceibias.n483 0.285035
R23146 commonsourceibias.n476 commonsourceibias.n367 0.189894
R23147 commonsourceibias.n476 commonsourceibias.n475 0.189894
R23148 commonsourceibias.n475 commonsourceibias.n474 0.189894
R23149 commonsourceibias.n474 commonsourceibias.n369 0.189894
R23150 commonsourceibias.n469 commonsourceibias.n369 0.189894
R23151 commonsourceibias.n469 commonsourceibias.n468 0.189894
R23152 commonsourceibias.n468 commonsourceibias.n467 0.189894
R23153 commonsourceibias.n467 commonsourceibias.n371 0.189894
R23154 commonsourceibias.n462 commonsourceibias.n371 0.189894
R23155 commonsourceibias.n462 commonsourceibias.n461 0.189894
R23156 commonsourceibias.n461 commonsourceibias.n460 0.189894
R23157 commonsourceibias.n460 commonsourceibias.n374 0.189894
R23158 commonsourceibias.n455 commonsourceibias.n374 0.189894
R23159 commonsourceibias.n455 commonsourceibias.n454 0.189894
R23160 commonsourceibias.n454 commonsourceibias.n453 0.189894
R23161 commonsourceibias.n453 commonsourceibias.n376 0.189894
R23162 commonsourceibias.n448 commonsourceibias.n376 0.189894
R23163 commonsourceibias.n448 commonsourceibias.n447 0.189894
R23164 commonsourceibias.n447 commonsourceibias.n446 0.189894
R23165 commonsourceibias.n446 commonsourceibias.n379 0.189894
R23166 commonsourceibias.n441 commonsourceibias.n379 0.189894
R23167 commonsourceibias.n441 commonsourceibias.n440 0.189894
R23168 commonsourceibias.n440 commonsourceibias.n439 0.189894
R23169 commonsourceibias.n439 commonsourceibias.n381 0.189894
R23170 commonsourceibias.n434 commonsourceibias.n381 0.189894
R23171 commonsourceibias.n434 commonsourceibias.n433 0.189894
R23172 commonsourceibias.n433 commonsourceibias.n432 0.189894
R23173 commonsourceibias.n432 commonsourceibias.n384 0.189894
R23174 commonsourceibias.n427 commonsourceibias.n384 0.189894
R23175 commonsourceibias.n427 commonsourceibias.n426 0.189894
R23176 commonsourceibias.n426 commonsourceibias.n425 0.189894
R23177 commonsourceibias.n425 commonsourceibias.n386 0.189894
R23178 commonsourceibias.n420 commonsourceibias.n386 0.189894
R23179 commonsourceibias.n420 commonsourceibias.n419 0.189894
R23180 commonsourceibias.n419 commonsourceibias.n418 0.189894
R23181 commonsourceibias.n418 commonsourceibias.n389 0.189894
R23182 commonsourceibias.n413 commonsourceibias.n389 0.189894
R23183 commonsourceibias.n413 commonsourceibias.n412 0.189894
R23184 commonsourceibias.n412 commonsourceibias.n411 0.189894
R23185 commonsourceibias.n411 commonsourceibias.n391 0.189894
R23186 commonsourceibias.n406 commonsourceibias.n391 0.189894
R23187 commonsourceibias.n406 commonsourceibias.n405 0.189894
R23188 commonsourceibias.n405 commonsourceibias.n404 0.189894
R23189 commonsourceibias.n404 commonsourceibias.n394 0.189894
R23190 commonsourceibias.n399 commonsourceibias.n394 0.189894
R23191 commonsourceibias.n399 commonsourceibias.n398 0.189894
R23192 commonsourceibias.n360 commonsourceibias.n251 0.189894
R23193 commonsourceibias.n360 commonsourceibias.n359 0.189894
R23194 commonsourceibias.n359 commonsourceibias.n358 0.189894
R23195 commonsourceibias.n358 commonsourceibias.n253 0.189894
R23196 commonsourceibias.n353 commonsourceibias.n253 0.189894
R23197 commonsourceibias.n353 commonsourceibias.n352 0.189894
R23198 commonsourceibias.n352 commonsourceibias.n351 0.189894
R23199 commonsourceibias.n351 commonsourceibias.n255 0.189894
R23200 commonsourceibias.n346 commonsourceibias.n255 0.189894
R23201 commonsourceibias.n346 commonsourceibias.n345 0.189894
R23202 commonsourceibias.n345 commonsourceibias.n344 0.189894
R23203 commonsourceibias.n344 commonsourceibias.n258 0.189894
R23204 commonsourceibias.n339 commonsourceibias.n258 0.189894
R23205 commonsourceibias.n339 commonsourceibias.n338 0.189894
R23206 commonsourceibias.n338 commonsourceibias.n337 0.189894
R23207 commonsourceibias.n337 commonsourceibias.n260 0.189894
R23208 commonsourceibias.n332 commonsourceibias.n260 0.189894
R23209 commonsourceibias.n332 commonsourceibias.n331 0.189894
R23210 commonsourceibias.n331 commonsourceibias.n330 0.189894
R23211 commonsourceibias.n330 commonsourceibias.n263 0.189894
R23212 commonsourceibias.n325 commonsourceibias.n263 0.189894
R23213 commonsourceibias.n325 commonsourceibias.n324 0.189894
R23214 commonsourceibias.n324 commonsourceibias.n323 0.189894
R23215 commonsourceibias.n323 commonsourceibias.n265 0.189894
R23216 commonsourceibias.n318 commonsourceibias.n265 0.189894
R23217 commonsourceibias.n318 commonsourceibias.n317 0.189894
R23218 commonsourceibias.n317 commonsourceibias.n316 0.189894
R23219 commonsourceibias.n316 commonsourceibias.n268 0.189894
R23220 commonsourceibias.n311 commonsourceibias.n268 0.189894
R23221 commonsourceibias.n311 commonsourceibias.n310 0.189894
R23222 commonsourceibias.n310 commonsourceibias.n309 0.189894
R23223 commonsourceibias.n309 commonsourceibias.n270 0.189894
R23224 commonsourceibias.n304 commonsourceibias.n270 0.189894
R23225 commonsourceibias.n304 commonsourceibias.n303 0.189894
R23226 commonsourceibias.n303 commonsourceibias.n302 0.189894
R23227 commonsourceibias.n302 commonsourceibias.n273 0.189894
R23228 commonsourceibias.n297 commonsourceibias.n273 0.189894
R23229 commonsourceibias.n297 commonsourceibias.n296 0.189894
R23230 commonsourceibias.n296 commonsourceibias.n295 0.189894
R23231 commonsourceibias.n295 commonsourceibias.n275 0.189894
R23232 commonsourceibias.n290 commonsourceibias.n275 0.189894
R23233 commonsourceibias.n290 commonsourceibias.n289 0.189894
R23234 commonsourceibias.n289 commonsourceibias.n288 0.189894
R23235 commonsourceibias.n288 commonsourceibias.n278 0.189894
R23236 commonsourceibias.n283 commonsourceibias.n278 0.189894
R23237 commonsourceibias.n283 commonsourceibias.n282 0.189894
R23238 commonsourceibias.n123 commonsourceibias.n14 0.189894
R23239 commonsourceibias.n123 commonsourceibias.n122 0.189894
R23240 commonsourceibias.n122 commonsourceibias.n121 0.189894
R23241 commonsourceibias.n121 commonsourceibias.n16 0.189894
R23242 commonsourceibias.n116 commonsourceibias.n16 0.189894
R23243 commonsourceibias.n116 commonsourceibias.n115 0.189894
R23244 commonsourceibias.n115 commonsourceibias.n114 0.189894
R23245 commonsourceibias.n114 commonsourceibias.n18 0.189894
R23246 commonsourceibias.n109 commonsourceibias.n18 0.189894
R23247 commonsourceibias.n109 commonsourceibias.n108 0.189894
R23248 commonsourceibias.n108 commonsourceibias.n107 0.189894
R23249 commonsourceibias.n107 commonsourceibias.n21 0.189894
R23250 commonsourceibias.n102 commonsourceibias.n21 0.189894
R23251 commonsourceibias.n102 commonsourceibias.n101 0.189894
R23252 commonsourceibias.n101 commonsourceibias.n100 0.189894
R23253 commonsourceibias.n100 commonsourceibias.n23 0.189894
R23254 commonsourceibias.n95 commonsourceibias.n23 0.189894
R23255 commonsourceibias.n95 commonsourceibias.n94 0.189894
R23256 commonsourceibias.n94 commonsourceibias.n93 0.189894
R23257 commonsourceibias.n93 commonsourceibias.n26 0.189894
R23258 commonsourceibias.n88 commonsourceibias.n26 0.189894
R23259 commonsourceibias.n88 commonsourceibias.n87 0.189894
R23260 commonsourceibias.n87 commonsourceibias.n86 0.189894
R23261 commonsourceibias.n86 commonsourceibias.n28 0.189894
R23262 commonsourceibias.n81 commonsourceibias.n28 0.189894
R23263 commonsourceibias.n81 commonsourceibias.n80 0.189894
R23264 commonsourceibias.n80 commonsourceibias.n79 0.189894
R23265 commonsourceibias.n79 commonsourceibias.n31 0.189894
R23266 commonsourceibias.n74 commonsourceibias.n31 0.189894
R23267 commonsourceibias.n74 commonsourceibias.n73 0.189894
R23268 commonsourceibias.n73 commonsourceibias.n72 0.189894
R23269 commonsourceibias.n72 commonsourceibias.n33 0.189894
R23270 commonsourceibias.n67 commonsourceibias.n33 0.189894
R23271 commonsourceibias.n67 commonsourceibias.n66 0.189894
R23272 commonsourceibias.n66 commonsourceibias.n65 0.189894
R23273 commonsourceibias.n65 commonsourceibias.n36 0.189894
R23274 commonsourceibias.n60 commonsourceibias.n36 0.189894
R23275 commonsourceibias.n60 commonsourceibias.n59 0.189894
R23276 commonsourceibias.n59 commonsourceibias.n58 0.189894
R23277 commonsourceibias.n58 commonsourceibias.n38 0.189894
R23278 commonsourceibias.n53 commonsourceibias.n38 0.189894
R23279 commonsourceibias.n53 commonsourceibias.n52 0.189894
R23280 commonsourceibias.n52 commonsourceibias.n51 0.189894
R23281 commonsourceibias.n51 commonsourceibias.n41 0.189894
R23282 commonsourceibias.n46 commonsourceibias.n41 0.189894
R23283 commonsourceibias.n46 commonsourceibias.n45 0.189894
R23284 commonsourceibias.n205 commonsourceibias.n204 0.189894
R23285 commonsourceibias.n204 commonsourceibias.n152 0.189894
R23286 commonsourceibias.n200 commonsourceibias.n152 0.189894
R23287 commonsourceibias.n200 commonsourceibias.n199 0.189894
R23288 commonsourceibias.n199 commonsourceibias.n154 0.189894
R23289 commonsourceibias.n195 commonsourceibias.n154 0.189894
R23290 commonsourceibias.n195 commonsourceibias.n194 0.189894
R23291 commonsourceibias.n194 commonsourceibias.n156 0.189894
R23292 commonsourceibias.n189 commonsourceibias.n156 0.189894
R23293 commonsourceibias.n189 commonsourceibias.n188 0.189894
R23294 commonsourceibias.n188 commonsourceibias.n187 0.189894
R23295 commonsourceibias.n187 commonsourceibias.n158 0.189894
R23296 commonsourceibias.n182 commonsourceibias.n158 0.189894
R23297 commonsourceibias.n182 commonsourceibias.n181 0.189894
R23298 commonsourceibias.n181 commonsourceibias.n180 0.189894
R23299 commonsourceibias.n180 commonsourceibias.n160 0.189894
R23300 commonsourceibias.n175 commonsourceibias.n160 0.189894
R23301 commonsourceibias.n175 commonsourceibias.n174 0.189894
R23302 commonsourceibias.n174 commonsourceibias.n173 0.189894
R23303 commonsourceibias.n173 commonsourceibias.n163 0.189894
R23304 commonsourceibias.n168 commonsourceibias.n163 0.189894
R23305 commonsourceibias.n168 commonsourceibias.n167 0.189894
R23306 commonsourceibias.n245 commonsourceibias.n0 0.189894
R23307 commonsourceibias.n245 commonsourceibias.n244 0.189894
R23308 commonsourceibias.n244 commonsourceibias.n243 0.189894
R23309 commonsourceibias.n243 commonsourceibias.n2 0.189894
R23310 commonsourceibias.n238 commonsourceibias.n2 0.189894
R23311 commonsourceibias.n238 commonsourceibias.n237 0.189894
R23312 commonsourceibias.n237 commonsourceibias.n236 0.189894
R23313 commonsourceibias.n236 commonsourceibias.n4 0.189894
R23314 commonsourceibias.n231 commonsourceibias.n4 0.189894
R23315 commonsourceibias.n231 commonsourceibias.n230 0.189894
R23316 commonsourceibias.n230 commonsourceibias.n229 0.189894
R23317 commonsourceibias.n229 commonsourceibias.n7 0.189894
R23318 commonsourceibias.n224 commonsourceibias.n7 0.189894
R23319 commonsourceibias.n224 commonsourceibias.n223 0.189894
R23320 commonsourceibias.n223 commonsourceibias.n222 0.189894
R23321 commonsourceibias.n222 commonsourceibias.n9 0.189894
R23322 commonsourceibias.n217 commonsourceibias.n9 0.189894
R23323 commonsourceibias.n217 commonsourceibias.n216 0.189894
R23324 commonsourceibias.n216 commonsourceibias.n215 0.189894
R23325 commonsourceibias.n215 commonsourceibias.n12 0.189894
R23326 commonsourceibias.n210 commonsourceibias.n12 0.189894
R23327 commonsourceibias.n210 commonsourceibias.n209 0.189894
R23328 commonsourceibias.n209 commonsourceibias.n208 0.189894
R23329 commonsourceibias.n877 commonsourceibias.n876 0.189894
R23330 commonsourceibias.n877 commonsourceibias.n872 0.189894
R23331 commonsourceibias.n882 commonsourceibias.n872 0.189894
R23332 commonsourceibias.n883 commonsourceibias.n882 0.189894
R23333 commonsourceibias.n884 commonsourceibias.n883 0.189894
R23334 commonsourceibias.n884 commonsourceibias.n870 0.189894
R23335 commonsourceibias.n890 commonsourceibias.n870 0.189894
R23336 commonsourceibias.n891 commonsourceibias.n890 0.189894
R23337 commonsourceibias.n892 commonsourceibias.n891 0.189894
R23338 commonsourceibias.n892 commonsourceibias.n868 0.189894
R23339 commonsourceibias.n897 commonsourceibias.n868 0.189894
R23340 commonsourceibias.n898 commonsourceibias.n897 0.189894
R23341 commonsourceibias.n899 commonsourceibias.n898 0.189894
R23342 commonsourceibias.n899 commonsourceibias.n866 0.189894
R23343 commonsourceibias.n905 commonsourceibias.n866 0.189894
R23344 commonsourceibias.n906 commonsourceibias.n905 0.189894
R23345 commonsourceibias.n907 commonsourceibias.n906 0.189894
R23346 commonsourceibias.n907 commonsourceibias.n864 0.189894
R23347 commonsourceibias.n912 commonsourceibias.n864 0.189894
R23348 commonsourceibias.n913 commonsourceibias.n912 0.189894
R23349 commonsourceibias.n914 commonsourceibias.n913 0.189894
R23350 commonsourceibias.n914 commonsourceibias.n862 0.189894
R23351 commonsourceibias.n920 commonsourceibias.n862 0.189894
R23352 commonsourceibias.n921 commonsourceibias.n920 0.189894
R23353 commonsourceibias.n922 commonsourceibias.n921 0.189894
R23354 commonsourceibias.n922 commonsourceibias.n860 0.189894
R23355 commonsourceibias.n927 commonsourceibias.n860 0.189894
R23356 commonsourceibias.n928 commonsourceibias.n927 0.189894
R23357 commonsourceibias.n929 commonsourceibias.n928 0.189894
R23358 commonsourceibias.n929 commonsourceibias.n858 0.189894
R23359 commonsourceibias.n935 commonsourceibias.n858 0.189894
R23360 commonsourceibias.n936 commonsourceibias.n935 0.189894
R23361 commonsourceibias.n937 commonsourceibias.n936 0.189894
R23362 commonsourceibias.n937 commonsourceibias.n856 0.189894
R23363 commonsourceibias.n942 commonsourceibias.n856 0.189894
R23364 commonsourceibias.n943 commonsourceibias.n942 0.189894
R23365 commonsourceibias.n944 commonsourceibias.n943 0.189894
R23366 commonsourceibias.n944 commonsourceibias.n854 0.189894
R23367 commonsourceibias.n950 commonsourceibias.n854 0.189894
R23368 commonsourceibias.n951 commonsourceibias.n950 0.189894
R23369 commonsourceibias.n952 commonsourceibias.n951 0.189894
R23370 commonsourceibias.n952 commonsourceibias.n852 0.189894
R23371 commonsourceibias.n957 commonsourceibias.n852 0.189894
R23372 commonsourceibias.n958 commonsourceibias.n957 0.189894
R23373 commonsourceibias.n959 commonsourceibias.n958 0.189894
R23374 commonsourceibias.n959 commonsourceibias.n850 0.189894
R23375 commonsourceibias.n761 commonsourceibias.n760 0.189894
R23376 commonsourceibias.n761 commonsourceibias.n756 0.189894
R23377 commonsourceibias.n766 commonsourceibias.n756 0.189894
R23378 commonsourceibias.n767 commonsourceibias.n766 0.189894
R23379 commonsourceibias.n768 commonsourceibias.n767 0.189894
R23380 commonsourceibias.n768 commonsourceibias.n754 0.189894
R23381 commonsourceibias.n774 commonsourceibias.n754 0.189894
R23382 commonsourceibias.n775 commonsourceibias.n774 0.189894
R23383 commonsourceibias.n776 commonsourceibias.n775 0.189894
R23384 commonsourceibias.n776 commonsourceibias.n752 0.189894
R23385 commonsourceibias.n781 commonsourceibias.n752 0.189894
R23386 commonsourceibias.n782 commonsourceibias.n781 0.189894
R23387 commonsourceibias.n783 commonsourceibias.n782 0.189894
R23388 commonsourceibias.n783 commonsourceibias.n750 0.189894
R23389 commonsourceibias.n789 commonsourceibias.n750 0.189894
R23390 commonsourceibias.n790 commonsourceibias.n789 0.189894
R23391 commonsourceibias.n791 commonsourceibias.n790 0.189894
R23392 commonsourceibias.n791 commonsourceibias.n748 0.189894
R23393 commonsourceibias.n796 commonsourceibias.n748 0.189894
R23394 commonsourceibias.n797 commonsourceibias.n796 0.189894
R23395 commonsourceibias.n798 commonsourceibias.n797 0.189894
R23396 commonsourceibias.n798 commonsourceibias.n746 0.189894
R23397 commonsourceibias.n804 commonsourceibias.n746 0.189894
R23398 commonsourceibias.n805 commonsourceibias.n804 0.189894
R23399 commonsourceibias.n806 commonsourceibias.n805 0.189894
R23400 commonsourceibias.n806 commonsourceibias.n744 0.189894
R23401 commonsourceibias.n811 commonsourceibias.n744 0.189894
R23402 commonsourceibias.n812 commonsourceibias.n811 0.189894
R23403 commonsourceibias.n813 commonsourceibias.n812 0.189894
R23404 commonsourceibias.n813 commonsourceibias.n742 0.189894
R23405 commonsourceibias.n819 commonsourceibias.n742 0.189894
R23406 commonsourceibias.n820 commonsourceibias.n819 0.189894
R23407 commonsourceibias.n821 commonsourceibias.n820 0.189894
R23408 commonsourceibias.n821 commonsourceibias.n740 0.189894
R23409 commonsourceibias.n826 commonsourceibias.n740 0.189894
R23410 commonsourceibias.n827 commonsourceibias.n826 0.189894
R23411 commonsourceibias.n828 commonsourceibias.n827 0.189894
R23412 commonsourceibias.n828 commonsourceibias.n738 0.189894
R23413 commonsourceibias.n834 commonsourceibias.n738 0.189894
R23414 commonsourceibias.n835 commonsourceibias.n834 0.189894
R23415 commonsourceibias.n836 commonsourceibias.n835 0.189894
R23416 commonsourceibias.n836 commonsourceibias.n736 0.189894
R23417 commonsourceibias.n841 commonsourceibias.n736 0.189894
R23418 commonsourceibias.n842 commonsourceibias.n841 0.189894
R23419 commonsourceibias.n843 commonsourceibias.n842 0.189894
R23420 commonsourceibias.n843 commonsourceibias.n734 0.189894
R23421 commonsourceibias.n531 commonsourceibias.n530 0.189894
R23422 commonsourceibias.n531 commonsourceibias.n526 0.189894
R23423 commonsourceibias.n536 commonsourceibias.n526 0.189894
R23424 commonsourceibias.n537 commonsourceibias.n536 0.189894
R23425 commonsourceibias.n538 commonsourceibias.n537 0.189894
R23426 commonsourceibias.n538 commonsourceibias.n524 0.189894
R23427 commonsourceibias.n544 commonsourceibias.n524 0.189894
R23428 commonsourceibias.n545 commonsourceibias.n544 0.189894
R23429 commonsourceibias.n546 commonsourceibias.n545 0.189894
R23430 commonsourceibias.n546 commonsourceibias.n522 0.189894
R23431 commonsourceibias.n551 commonsourceibias.n522 0.189894
R23432 commonsourceibias.n552 commonsourceibias.n551 0.189894
R23433 commonsourceibias.n553 commonsourceibias.n552 0.189894
R23434 commonsourceibias.n553 commonsourceibias.n520 0.189894
R23435 commonsourceibias.n559 commonsourceibias.n520 0.189894
R23436 commonsourceibias.n560 commonsourceibias.n559 0.189894
R23437 commonsourceibias.n561 commonsourceibias.n560 0.189894
R23438 commonsourceibias.n561 commonsourceibias.n518 0.189894
R23439 commonsourceibias.n566 commonsourceibias.n518 0.189894
R23440 commonsourceibias.n567 commonsourceibias.n566 0.189894
R23441 commonsourceibias.n568 commonsourceibias.n567 0.189894
R23442 commonsourceibias.n568 commonsourceibias.n516 0.189894
R23443 commonsourceibias.n574 commonsourceibias.n516 0.189894
R23444 commonsourceibias.n575 commonsourceibias.n574 0.189894
R23445 commonsourceibias.n576 commonsourceibias.n575 0.189894
R23446 commonsourceibias.n576 commonsourceibias.n514 0.189894
R23447 commonsourceibias.n581 commonsourceibias.n514 0.189894
R23448 commonsourceibias.n582 commonsourceibias.n581 0.189894
R23449 commonsourceibias.n583 commonsourceibias.n582 0.189894
R23450 commonsourceibias.n583 commonsourceibias.n512 0.189894
R23451 commonsourceibias.n589 commonsourceibias.n512 0.189894
R23452 commonsourceibias.n590 commonsourceibias.n589 0.189894
R23453 commonsourceibias.n591 commonsourceibias.n590 0.189894
R23454 commonsourceibias.n591 commonsourceibias.n510 0.189894
R23455 commonsourceibias.n596 commonsourceibias.n510 0.189894
R23456 commonsourceibias.n597 commonsourceibias.n596 0.189894
R23457 commonsourceibias.n598 commonsourceibias.n597 0.189894
R23458 commonsourceibias.n598 commonsourceibias.n508 0.189894
R23459 commonsourceibias.n604 commonsourceibias.n508 0.189894
R23460 commonsourceibias.n605 commonsourceibias.n604 0.189894
R23461 commonsourceibias.n606 commonsourceibias.n605 0.189894
R23462 commonsourceibias.n606 commonsourceibias.n506 0.189894
R23463 commonsourceibias.n611 commonsourceibias.n506 0.189894
R23464 commonsourceibias.n612 commonsourceibias.n611 0.189894
R23465 commonsourceibias.n613 commonsourceibias.n612 0.189894
R23466 commonsourceibias.n613 commonsourceibias.n504 0.189894
R23467 commonsourceibias.n647 commonsourceibias.n646 0.189894
R23468 commonsourceibias.n647 commonsourceibias.n642 0.189894
R23469 commonsourceibias.n652 commonsourceibias.n642 0.189894
R23470 commonsourceibias.n653 commonsourceibias.n652 0.189894
R23471 commonsourceibias.n654 commonsourceibias.n653 0.189894
R23472 commonsourceibias.n654 commonsourceibias.n640 0.189894
R23473 commonsourceibias.n660 commonsourceibias.n640 0.189894
R23474 commonsourceibias.n661 commonsourceibias.n660 0.189894
R23475 commonsourceibias.n662 commonsourceibias.n661 0.189894
R23476 commonsourceibias.n662 commonsourceibias.n638 0.189894
R23477 commonsourceibias.n667 commonsourceibias.n638 0.189894
R23478 commonsourceibias.n668 commonsourceibias.n667 0.189894
R23479 commonsourceibias.n669 commonsourceibias.n668 0.189894
R23480 commonsourceibias.n669 commonsourceibias.n636 0.189894
R23481 commonsourceibias.n674 commonsourceibias.n636 0.189894
R23482 commonsourceibias.n675 commonsourceibias.n674 0.189894
R23483 commonsourceibias.n675 commonsourceibias.n634 0.189894
R23484 commonsourceibias.n679 commonsourceibias.n634 0.189894
R23485 commonsourceibias.n680 commonsourceibias.n679 0.189894
R23486 commonsourceibias.n680 commonsourceibias.n632 0.189894
R23487 commonsourceibias.n684 commonsourceibias.n632 0.189894
R23488 commonsourceibias.n685 commonsourceibias.n684 0.189894
R23489 commonsourceibias.n690 commonsourceibias.n689 0.189894
R23490 commonsourceibias.n691 commonsourceibias.n690 0.189894
R23491 commonsourceibias.n691 commonsourceibias.n493 0.189894
R23492 commonsourceibias.n696 commonsourceibias.n493 0.189894
R23493 commonsourceibias.n697 commonsourceibias.n696 0.189894
R23494 commonsourceibias.n698 commonsourceibias.n697 0.189894
R23495 commonsourceibias.n698 commonsourceibias.n491 0.189894
R23496 commonsourceibias.n704 commonsourceibias.n491 0.189894
R23497 commonsourceibias.n705 commonsourceibias.n704 0.189894
R23498 commonsourceibias.n706 commonsourceibias.n705 0.189894
R23499 commonsourceibias.n706 commonsourceibias.n489 0.189894
R23500 commonsourceibias.n711 commonsourceibias.n489 0.189894
R23501 commonsourceibias.n712 commonsourceibias.n711 0.189894
R23502 commonsourceibias.n713 commonsourceibias.n712 0.189894
R23503 commonsourceibias.n713 commonsourceibias.n487 0.189894
R23504 commonsourceibias.n719 commonsourceibias.n487 0.189894
R23505 commonsourceibias.n720 commonsourceibias.n719 0.189894
R23506 commonsourceibias.n721 commonsourceibias.n720 0.189894
R23507 commonsourceibias.n721 commonsourceibias.n485 0.189894
R23508 commonsourceibias.n726 commonsourceibias.n485 0.189894
R23509 commonsourceibias.n727 commonsourceibias.n726 0.189894
R23510 commonsourceibias.n728 commonsourceibias.n727 0.189894
R23511 commonsourceibias.n728 commonsourceibias.n483 0.189894
R23512 commonsourceibias.n205 commonsourceibias.n149 0.0762576
R23513 commonsourceibias.n208 commonsourceibias.n149 0.0762576
R23514 commonsourceibias.n685 commonsourceibias.n630 0.0762576
R23515 commonsourceibias.n689 commonsourceibias.n630 0.0762576
R23516 CSoutput.n19 CSoutput.t235 184.661
R23517 CSoutput.n78 CSoutput.n77 165.8
R23518 CSoutput.n76 CSoutput.n0 165.8
R23519 CSoutput.n75 CSoutput.n74 165.8
R23520 CSoutput.n73 CSoutput.n72 165.8
R23521 CSoutput.n71 CSoutput.n2 165.8
R23522 CSoutput.n69 CSoutput.n68 165.8
R23523 CSoutput.n67 CSoutput.n3 165.8
R23524 CSoutput.n66 CSoutput.n65 165.8
R23525 CSoutput.n63 CSoutput.n4 165.8
R23526 CSoutput.n61 CSoutput.n60 165.8
R23527 CSoutput.n59 CSoutput.n5 165.8
R23528 CSoutput.n58 CSoutput.n57 165.8
R23529 CSoutput.n55 CSoutput.n6 165.8
R23530 CSoutput.n54 CSoutput.n53 165.8
R23531 CSoutput.n52 CSoutput.n51 165.8
R23532 CSoutput.n50 CSoutput.n8 165.8
R23533 CSoutput.n48 CSoutput.n47 165.8
R23534 CSoutput.n46 CSoutput.n9 165.8
R23535 CSoutput.n45 CSoutput.n44 165.8
R23536 CSoutput.n42 CSoutput.n10 165.8
R23537 CSoutput.n41 CSoutput.n40 165.8
R23538 CSoutput.n39 CSoutput.n38 165.8
R23539 CSoutput.n37 CSoutput.n12 165.8
R23540 CSoutput.n35 CSoutput.n34 165.8
R23541 CSoutput.n33 CSoutput.n13 165.8
R23542 CSoutput.n32 CSoutput.n31 165.8
R23543 CSoutput.n29 CSoutput.n14 165.8
R23544 CSoutput.n28 CSoutput.n27 165.8
R23545 CSoutput.n26 CSoutput.n25 165.8
R23546 CSoutput.n24 CSoutput.n16 165.8
R23547 CSoutput.n22 CSoutput.n21 165.8
R23548 CSoutput.n20 CSoutput.n17 165.8
R23549 CSoutput.n77 CSoutput.t236 162.194
R23550 CSoutput.n18 CSoutput.t225 120.501
R23551 CSoutput.n23 CSoutput.t227 120.501
R23552 CSoutput.n15 CSoutput.t220 120.501
R23553 CSoutput.n30 CSoutput.t233 120.501
R23554 CSoutput.n36 CSoutput.t228 120.501
R23555 CSoutput.n11 CSoutput.t223 120.501
R23556 CSoutput.n43 CSoutput.t218 120.501
R23557 CSoutput.n49 CSoutput.t229 120.501
R23558 CSoutput.n7 CSoutput.t231 120.501
R23559 CSoutput.n56 CSoutput.t221 120.501
R23560 CSoutput.n62 CSoutput.t217 120.501
R23561 CSoutput.n64 CSoutput.t234 120.501
R23562 CSoutput.n70 CSoutput.t224 120.501
R23563 CSoutput.n1 CSoutput.t226 120.501
R23564 CSoutput.n310 CSoutput.n308 103.469
R23565 CSoutput.n294 CSoutput.n292 103.469
R23566 CSoutput.n279 CSoutput.n277 103.469
R23567 CSoutput.n112 CSoutput.n110 103.469
R23568 CSoutput.n96 CSoutput.n94 103.469
R23569 CSoutput.n81 CSoutput.n79 103.469
R23570 CSoutput.n320 CSoutput.n319 103.111
R23571 CSoutput.n318 CSoutput.n317 103.111
R23572 CSoutput.n316 CSoutput.n315 103.111
R23573 CSoutput.n314 CSoutput.n313 103.111
R23574 CSoutput.n312 CSoutput.n311 103.111
R23575 CSoutput.n310 CSoutput.n309 103.111
R23576 CSoutput.n306 CSoutput.n305 103.111
R23577 CSoutput.n304 CSoutput.n303 103.111
R23578 CSoutput.n302 CSoutput.n301 103.111
R23579 CSoutput.n300 CSoutput.n299 103.111
R23580 CSoutput.n298 CSoutput.n297 103.111
R23581 CSoutput.n296 CSoutput.n295 103.111
R23582 CSoutput.n294 CSoutput.n293 103.111
R23583 CSoutput.n291 CSoutput.n290 103.111
R23584 CSoutput.n289 CSoutput.n288 103.111
R23585 CSoutput.n287 CSoutput.n286 103.111
R23586 CSoutput.n285 CSoutput.n284 103.111
R23587 CSoutput.n283 CSoutput.n282 103.111
R23588 CSoutput.n281 CSoutput.n280 103.111
R23589 CSoutput.n279 CSoutput.n278 103.111
R23590 CSoutput.n112 CSoutput.n111 103.111
R23591 CSoutput.n114 CSoutput.n113 103.111
R23592 CSoutput.n116 CSoutput.n115 103.111
R23593 CSoutput.n118 CSoutput.n117 103.111
R23594 CSoutput.n120 CSoutput.n119 103.111
R23595 CSoutput.n122 CSoutput.n121 103.111
R23596 CSoutput.n124 CSoutput.n123 103.111
R23597 CSoutput.n96 CSoutput.n95 103.111
R23598 CSoutput.n98 CSoutput.n97 103.111
R23599 CSoutput.n100 CSoutput.n99 103.111
R23600 CSoutput.n102 CSoutput.n101 103.111
R23601 CSoutput.n104 CSoutput.n103 103.111
R23602 CSoutput.n106 CSoutput.n105 103.111
R23603 CSoutput.n108 CSoutput.n107 103.111
R23604 CSoutput.n81 CSoutput.n80 103.111
R23605 CSoutput.n83 CSoutput.n82 103.111
R23606 CSoutput.n85 CSoutput.n84 103.111
R23607 CSoutput.n87 CSoutput.n86 103.111
R23608 CSoutput.n89 CSoutput.n88 103.111
R23609 CSoutput.n91 CSoutput.n90 103.111
R23610 CSoutput.n93 CSoutput.n92 103.111
R23611 CSoutput.n322 CSoutput.n321 103.111
R23612 CSoutput.n366 CSoutput.n364 81.5057
R23613 CSoutput.n346 CSoutput.n344 81.5057
R23614 CSoutput.n327 CSoutput.n325 81.5057
R23615 CSoutput.n426 CSoutput.n424 81.5057
R23616 CSoutput.n406 CSoutput.n404 81.5057
R23617 CSoutput.n387 CSoutput.n385 81.5057
R23618 CSoutput.n382 CSoutput.n381 80.9324
R23619 CSoutput.n380 CSoutput.n379 80.9324
R23620 CSoutput.n378 CSoutput.n377 80.9324
R23621 CSoutput.n376 CSoutput.n375 80.9324
R23622 CSoutput.n374 CSoutput.n373 80.9324
R23623 CSoutput.n372 CSoutput.n371 80.9324
R23624 CSoutput.n370 CSoutput.n369 80.9324
R23625 CSoutput.n368 CSoutput.n367 80.9324
R23626 CSoutput.n366 CSoutput.n365 80.9324
R23627 CSoutput.n362 CSoutput.n361 80.9324
R23628 CSoutput.n360 CSoutput.n359 80.9324
R23629 CSoutput.n358 CSoutput.n357 80.9324
R23630 CSoutput.n356 CSoutput.n355 80.9324
R23631 CSoutput.n354 CSoutput.n353 80.9324
R23632 CSoutput.n352 CSoutput.n351 80.9324
R23633 CSoutput.n350 CSoutput.n349 80.9324
R23634 CSoutput.n348 CSoutput.n347 80.9324
R23635 CSoutput.n346 CSoutput.n345 80.9324
R23636 CSoutput.n343 CSoutput.n342 80.9324
R23637 CSoutput.n341 CSoutput.n340 80.9324
R23638 CSoutput.n339 CSoutput.n338 80.9324
R23639 CSoutput.n337 CSoutput.n336 80.9324
R23640 CSoutput.n335 CSoutput.n334 80.9324
R23641 CSoutput.n333 CSoutput.n332 80.9324
R23642 CSoutput.n331 CSoutput.n330 80.9324
R23643 CSoutput.n329 CSoutput.n328 80.9324
R23644 CSoutput.n327 CSoutput.n326 80.9324
R23645 CSoutput.n426 CSoutput.n425 80.9324
R23646 CSoutput.n428 CSoutput.n427 80.9324
R23647 CSoutput.n430 CSoutput.n429 80.9324
R23648 CSoutput.n432 CSoutput.n431 80.9324
R23649 CSoutput.n434 CSoutput.n433 80.9324
R23650 CSoutput.n436 CSoutput.n435 80.9324
R23651 CSoutput.n438 CSoutput.n437 80.9324
R23652 CSoutput.n440 CSoutput.n439 80.9324
R23653 CSoutput.n442 CSoutput.n441 80.9324
R23654 CSoutput.n406 CSoutput.n405 80.9324
R23655 CSoutput.n408 CSoutput.n407 80.9324
R23656 CSoutput.n410 CSoutput.n409 80.9324
R23657 CSoutput.n412 CSoutput.n411 80.9324
R23658 CSoutput.n414 CSoutput.n413 80.9324
R23659 CSoutput.n416 CSoutput.n415 80.9324
R23660 CSoutput.n418 CSoutput.n417 80.9324
R23661 CSoutput.n420 CSoutput.n419 80.9324
R23662 CSoutput.n422 CSoutput.n421 80.9324
R23663 CSoutput.n387 CSoutput.n386 80.9324
R23664 CSoutput.n389 CSoutput.n388 80.9324
R23665 CSoutput.n391 CSoutput.n390 80.9324
R23666 CSoutput.n393 CSoutput.n392 80.9324
R23667 CSoutput.n395 CSoutput.n394 80.9324
R23668 CSoutput.n397 CSoutput.n396 80.9324
R23669 CSoutput.n399 CSoutput.n398 80.9324
R23670 CSoutput.n401 CSoutput.n400 80.9324
R23671 CSoutput.n403 CSoutput.n402 80.9324
R23672 CSoutput.n25 CSoutput.n24 48.1486
R23673 CSoutput.n69 CSoutput.n3 48.1486
R23674 CSoutput.n38 CSoutput.n37 48.1486
R23675 CSoutput.n42 CSoutput.n41 48.1486
R23676 CSoutput.n51 CSoutput.n50 48.1486
R23677 CSoutput.n55 CSoutput.n54 48.1486
R23678 CSoutput.n22 CSoutput.n17 46.462
R23679 CSoutput.n72 CSoutput.n71 46.462
R23680 CSoutput.n20 CSoutput.n19 44.9055
R23681 CSoutput.n29 CSoutput.n28 43.7635
R23682 CSoutput.n65 CSoutput.n63 43.7635
R23683 CSoutput.n35 CSoutput.n13 41.7396
R23684 CSoutput.n57 CSoutput.n5 41.7396
R23685 CSoutput.n44 CSoutput.n9 37.0171
R23686 CSoutput.n48 CSoutput.n9 37.0171
R23687 CSoutput.n76 CSoutput.n75 34.9932
R23688 CSoutput.n31 CSoutput.n13 32.2947
R23689 CSoutput.n61 CSoutput.n5 32.2947
R23690 CSoutput.n30 CSoutput.n29 29.6014
R23691 CSoutput.n63 CSoutput.n62 29.6014
R23692 CSoutput.n19 CSoutput.n18 28.4085
R23693 CSoutput.n18 CSoutput.n17 25.1176
R23694 CSoutput.n72 CSoutput.n1 25.1176
R23695 CSoutput.n43 CSoutput.n42 22.0922
R23696 CSoutput.n50 CSoutput.n49 22.0922
R23697 CSoutput.n77 CSoutput.n76 21.8586
R23698 CSoutput.n37 CSoutput.n36 18.9681
R23699 CSoutput.n56 CSoutput.n55 18.9681
R23700 CSoutput.n25 CSoutput.n15 17.6292
R23701 CSoutput.n64 CSoutput.n3 17.6292
R23702 CSoutput.n24 CSoutput.n23 15.844
R23703 CSoutput.n70 CSoutput.n69 15.844
R23704 CSoutput.n38 CSoutput.n11 14.5051
R23705 CSoutput.n54 CSoutput.n7 14.5051
R23706 CSoutput.n445 CSoutput.n78 11.4982
R23707 CSoutput.n41 CSoutput.n11 11.3811
R23708 CSoutput.n51 CSoutput.n7 11.3811
R23709 CSoutput.n23 CSoutput.n22 10.0422
R23710 CSoutput.n71 CSoutput.n70 10.0422
R23711 CSoutput.n307 CSoutput.n291 9.25285
R23712 CSoutput.n109 CSoutput.n93 9.25285
R23713 CSoutput.n363 CSoutput.n343 8.98182
R23714 CSoutput.n423 CSoutput.n403 8.98182
R23715 CSoutput.n384 CSoutput.n324 8.74155
R23716 CSoutput.n28 CSoutput.n15 8.25698
R23717 CSoutput.n65 CSoutput.n64 8.25698
R23718 CSoutput.n324 CSoutput.n323 7.12641
R23719 CSoutput.n126 CSoutput.n125 7.12641
R23720 CSoutput.n36 CSoutput.n35 6.91809
R23721 CSoutput.n57 CSoutput.n56 6.91809
R23722 CSoutput.n384 CSoutput.n383 6.02792
R23723 CSoutput.n444 CSoutput.n443 6.02792
R23724 CSoutput.n383 CSoutput.n382 5.25266
R23725 CSoutput.n363 CSoutput.n362 5.25266
R23726 CSoutput.n443 CSoutput.n442 5.25266
R23727 CSoutput.n423 CSoutput.n422 5.25266
R23728 CSoutput.n445 CSoutput.n126 5.14911
R23729 CSoutput.n323 CSoutput.n322 5.1449
R23730 CSoutput.n307 CSoutput.n306 5.1449
R23731 CSoutput.n125 CSoutput.n124 5.1449
R23732 CSoutput.n109 CSoutput.n108 5.1449
R23733 CSoutput.n217 CSoutput.n170 4.5005
R23734 CSoutput.n186 CSoutput.n170 4.5005
R23735 CSoutput.n181 CSoutput.n165 4.5005
R23736 CSoutput.n181 CSoutput.n167 4.5005
R23737 CSoutput.n181 CSoutput.n164 4.5005
R23738 CSoutput.n181 CSoutput.n168 4.5005
R23739 CSoutput.n181 CSoutput.n163 4.5005
R23740 CSoutput.n181 CSoutput.t237 4.5005
R23741 CSoutput.n181 CSoutput.n162 4.5005
R23742 CSoutput.n181 CSoutput.n169 4.5005
R23743 CSoutput.n181 CSoutput.n170 4.5005
R23744 CSoutput.n179 CSoutput.n165 4.5005
R23745 CSoutput.n179 CSoutput.n167 4.5005
R23746 CSoutput.n179 CSoutput.n164 4.5005
R23747 CSoutput.n179 CSoutput.n168 4.5005
R23748 CSoutput.n179 CSoutput.n163 4.5005
R23749 CSoutput.n179 CSoutput.t237 4.5005
R23750 CSoutput.n179 CSoutput.n162 4.5005
R23751 CSoutput.n179 CSoutput.n169 4.5005
R23752 CSoutput.n179 CSoutput.n170 4.5005
R23753 CSoutput.n178 CSoutput.n165 4.5005
R23754 CSoutput.n178 CSoutput.n167 4.5005
R23755 CSoutput.n178 CSoutput.n164 4.5005
R23756 CSoutput.n178 CSoutput.n168 4.5005
R23757 CSoutput.n178 CSoutput.n163 4.5005
R23758 CSoutput.n178 CSoutput.t237 4.5005
R23759 CSoutput.n178 CSoutput.n162 4.5005
R23760 CSoutput.n178 CSoutput.n169 4.5005
R23761 CSoutput.n178 CSoutput.n170 4.5005
R23762 CSoutput.n263 CSoutput.n165 4.5005
R23763 CSoutput.n263 CSoutput.n167 4.5005
R23764 CSoutput.n263 CSoutput.n164 4.5005
R23765 CSoutput.n263 CSoutput.n168 4.5005
R23766 CSoutput.n263 CSoutput.n163 4.5005
R23767 CSoutput.n263 CSoutput.t237 4.5005
R23768 CSoutput.n263 CSoutput.n162 4.5005
R23769 CSoutput.n263 CSoutput.n169 4.5005
R23770 CSoutput.n263 CSoutput.n170 4.5005
R23771 CSoutput.n261 CSoutput.n165 4.5005
R23772 CSoutput.n261 CSoutput.n167 4.5005
R23773 CSoutput.n261 CSoutput.n164 4.5005
R23774 CSoutput.n261 CSoutput.n168 4.5005
R23775 CSoutput.n261 CSoutput.n163 4.5005
R23776 CSoutput.n261 CSoutput.t237 4.5005
R23777 CSoutput.n261 CSoutput.n162 4.5005
R23778 CSoutput.n261 CSoutput.n169 4.5005
R23779 CSoutput.n259 CSoutput.n165 4.5005
R23780 CSoutput.n259 CSoutput.n167 4.5005
R23781 CSoutput.n259 CSoutput.n164 4.5005
R23782 CSoutput.n259 CSoutput.n168 4.5005
R23783 CSoutput.n259 CSoutput.n163 4.5005
R23784 CSoutput.n259 CSoutput.t237 4.5005
R23785 CSoutput.n259 CSoutput.n162 4.5005
R23786 CSoutput.n259 CSoutput.n169 4.5005
R23787 CSoutput.n189 CSoutput.n165 4.5005
R23788 CSoutput.n189 CSoutput.n167 4.5005
R23789 CSoutput.n189 CSoutput.n164 4.5005
R23790 CSoutput.n189 CSoutput.n168 4.5005
R23791 CSoutput.n189 CSoutput.n163 4.5005
R23792 CSoutput.n189 CSoutput.t237 4.5005
R23793 CSoutput.n189 CSoutput.n162 4.5005
R23794 CSoutput.n189 CSoutput.n169 4.5005
R23795 CSoutput.n189 CSoutput.n170 4.5005
R23796 CSoutput.n188 CSoutput.n165 4.5005
R23797 CSoutput.n188 CSoutput.n167 4.5005
R23798 CSoutput.n188 CSoutput.n164 4.5005
R23799 CSoutput.n188 CSoutput.n168 4.5005
R23800 CSoutput.n188 CSoutput.n163 4.5005
R23801 CSoutput.n188 CSoutput.t237 4.5005
R23802 CSoutput.n188 CSoutput.n162 4.5005
R23803 CSoutput.n188 CSoutput.n169 4.5005
R23804 CSoutput.n188 CSoutput.n170 4.5005
R23805 CSoutput.n192 CSoutput.n165 4.5005
R23806 CSoutput.n192 CSoutput.n167 4.5005
R23807 CSoutput.n192 CSoutput.n164 4.5005
R23808 CSoutput.n192 CSoutput.n168 4.5005
R23809 CSoutput.n192 CSoutput.n163 4.5005
R23810 CSoutput.n192 CSoutput.t237 4.5005
R23811 CSoutput.n192 CSoutput.n162 4.5005
R23812 CSoutput.n192 CSoutput.n169 4.5005
R23813 CSoutput.n192 CSoutput.n170 4.5005
R23814 CSoutput.n191 CSoutput.n165 4.5005
R23815 CSoutput.n191 CSoutput.n167 4.5005
R23816 CSoutput.n191 CSoutput.n164 4.5005
R23817 CSoutput.n191 CSoutput.n168 4.5005
R23818 CSoutput.n191 CSoutput.n163 4.5005
R23819 CSoutput.n191 CSoutput.t237 4.5005
R23820 CSoutput.n191 CSoutput.n162 4.5005
R23821 CSoutput.n191 CSoutput.n169 4.5005
R23822 CSoutput.n191 CSoutput.n170 4.5005
R23823 CSoutput.n174 CSoutput.n165 4.5005
R23824 CSoutput.n174 CSoutput.n167 4.5005
R23825 CSoutput.n174 CSoutput.n164 4.5005
R23826 CSoutput.n174 CSoutput.n168 4.5005
R23827 CSoutput.n174 CSoutput.n163 4.5005
R23828 CSoutput.n174 CSoutput.t237 4.5005
R23829 CSoutput.n174 CSoutput.n162 4.5005
R23830 CSoutput.n174 CSoutput.n169 4.5005
R23831 CSoutput.n174 CSoutput.n170 4.5005
R23832 CSoutput.n266 CSoutput.n165 4.5005
R23833 CSoutput.n266 CSoutput.n167 4.5005
R23834 CSoutput.n266 CSoutput.n164 4.5005
R23835 CSoutput.n266 CSoutput.n168 4.5005
R23836 CSoutput.n266 CSoutput.n163 4.5005
R23837 CSoutput.n266 CSoutput.t237 4.5005
R23838 CSoutput.n266 CSoutput.n162 4.5005
R23839 CSoutput.n266 CSoutput.n169 4.5005
R23840 CSoutput.n266 CSoutput.n170 4.5005
R23841 CSoutput.n253 CSoutput.n224 4.5005
R23842 CSoutput.n253 CSoutput.n230 4.5005
R23843 CSoutput.n211 CSoutput.n200 4.5005
R23844 CSoutput.n211 CSoutput.n202 4.5005
R23845 CSoutput.n211 CSoutput.n199 4.5005
R23846 CSoutput.n211 CSoutput.n203 4.5005
R23847 CSoutput.n211 CSoutput.n198 4.5005
R23848 CSoutput.n211 CSoutput.t232 4.5005
R23849 CSoutput.n211 CSoutput.n197 4.5005
R23850 CSoutput.n211 CSoutput.n204 4.5005
R23851 CSoutput.n253 CSoutput.n211 4.5005
R23852 CSoutput.n232 CSoutput.n200 4.5005
R23853 CSoutput.n232 CSoutput.n202 4.5005
R23854 CSoutput.n232 CSoutput.n199 4.5005
R23855 CSoutput.n232 CSoutput.n203 4.5005
R23856 CSoutput.n232 CSoutput.n198 4.5005
R23857 CSoutput.n232 CSoutput.t232 4.5005
R23858 CSoutput.n232 CSoutput.n197 4.5005
R23859 CSoutput.n232 CSoutput.n204 4.5005
R23860 CSoutput.n253 CSoutput.n232 4.5005
R23861 CSoutput.n210 CSoutput.n200 4.5005
R23862 CSoutput.n210 CSoutput.n202 4.5005
R23863 CSoutput.n210 CSoutput.n199 4.5005
R23864 CSoutput.n210 CSoutput.n203 4.5005
R23865 CSoutput.n210 CSoutput.n198 4.5005
R23866 CSoutput.n210 CSoutput.t232 4.5005
R23867 CSoutput.n210 CSoutput.n197 4.5005
R23868 CSoutput.n210 CSoutput.n204 4.5005
R23869 CSoutput.n253 CSoutput.n210 4.5005
R23870 CSoutput.n234 CSoutput.n200 4.5005
R23871 CSoutput.n234 CSoutput.n202 4.5005
R23872 CSoutput.n234 CSoutput.n199 4.5005
R23873 CSoutput.n234 CSoutput.n203 4.5005
R23874 CSoutput.n234 CSoutput.n198 4.5005
R23875 CSoutput.n234 CSoutput.t232 4.5005
R23876 CSoutput.n234 CSoutput.n197 4.5005
R23877 CSoutput.n234 CSoutput.n204 4.5005
R23878 CSoutput.n253 CSoutput.n234 4.5005
R23879 CSoutput.n200 CSoutput.n195 4.5005
R23880 CSoutput.n202 CSoutput.n195 4.5005
R23881 CSoutput.n199 CSoutput.n195 4.5005
R23882 CSoutput.n203 CSoutput.n195 4.5005
R23883 CSoutput.n198 CSoutput.n195 4.5005
R23884 CSoutput.t232 CSoutput.n195 4.5005
R23885 CSoutput.n197 CSoutput.n195 4.5005
R23886 CSoutput.n204 CSoutput.n195 4.5005
R23887 CSoutput.n256 CSoutput.n200 4.5005
R23888 CSoutput.n256 CSoutput.n202 4.5005
R23889 CSoutput.n256 CSoutput.n199 4.5005
R23890 CSoutput.n256 CSoutput.n203 4.5005
R23891 CSoutput.n256 CSoutput.n198 4.5005
R23892 CSoutput.n256 CSoutput.t232 4.5005
R23893 CSoutput.n256 CSoutput.n197 4.5005
R23894 CSoutput.n256 CSoutput.n204 4.5005
R23895 CSoutput.n254 CSoutput.n200 4.5005
R23896 CSoutput.n254 CSoutput.n202 4.5005
R23897 CSoutput.n254 CSoutput.n199 4.5005
R23898 CSoutput.n254 CSoutput.n203 4.5005
R23899 CSoutput.n254 CSoutput.n198 4.5005
R23900 CSoutput.n254 CSoutput.t232 4.5005
R23901 CSoutput.n254 CSoutput.n197 4.5005
R23902 CSoutput.n254 CSoutput.n204 4.5005
R23903 CSoutput.n254 CSoutput.n253 4.5005
R23904 CSoutput.n236 CSoutput.n200 4.5005
R23905 CSoutput.n236 CSoutput.n202 4.5005
R23906 CSoutput.n236 CSoutput.n199 4.5005
R23907 CSoutput.n236 CSoutput.n203 4.5005
R23908 CSoutput.n236 CSoutput.n198 4.5005
R23909 CSoutput.n236 CSoutput.t232 4.5005
R23910 CSoutput.n236 CSoutput.n197 4.5005
R23911 CSoutput.n236 CSoutput.n204 4.5005
R23912 CSoutput.n253 CSoutput.n236 4.5005
R23913 CSoutput.n208 CSoutput.n200 4.5005
R23914 CSoutput.n208 CSoutput.n202 4.5005
R23915 CSoutput.n208 CSoutput.n199 4.5005
R23916 CSoutput.n208 CSoutput.n203 4.5005
R23917 CSoutput.n208 CSoutput.n198 4.5005
R23918 CSoutput.n208 CSoutput.t232 4.5005
R23919 CSoutput.n208 CSoutput.n197 4.5005
R23920 CSoutput.n208 CSoutput.n204 4.5005
R23921 CSoutput.n253 CSoutput.n208 4.5005
R23922 CSoutput.n238 CSoutput.n200 4.5005
R23923 CSoutput.n238 CSoutput.n202 4.5005
R23924 CSoutput.n238 CSoutput.n199 4.5005
R23925 CSoutput.n238 CSoutput.n203 4.5005
R23926 CSoutput.n238 CSoutput.n198 4.5005
R23927 CSoutput.n238 CSoutput.t232 4.5005
R23928 CSoutput.n238 CSoutput.n197 4.5005
R23929 CSoutput.n238 CSoutput.n204 4.5005
R23930 CSoutput.n253 CSoutput.n238 4.5005
R23931 CSoutput.n207 CSoutput.n200 4.5005
R23932 CSoutput.n207 CSoutput.n202 4.5005
R23933 CSoutput.n207 CSoutput.n199 4.5005
R23934 CSoutput.n207 CSoutput.n203 4.5005
R23935 CSoutput.n207 CSoutput.n198 4.5005
R23936 CSoutput.n207 CSoutput.t232 4.5005
R23937 CSoutput.n207 CSoutput.n197 4.5005
R23938 CSoutput.n207 CSoutput.n204 4.5005
R23939 CSoutput.n253 CSoutput.n207 4.5005
R23940 CSoutput.n252 CSoutput.n200 4.5005
R23941 CSoutput.n252 CSoutput.n202 4.5005
R23942 CSoutput.n252 CSoutput.n199 4.5005
R23943 CSoutput.n252 CSoutput.n203 4.5005
R23944 CSoutput.n252 CSoutput.n198 4.5005
R23945 CSoutput.n252 CSoutput.t232 4.5005
R23946 CSoutput.n252 CSoutput.n197 4.5005
R23947 CSoutput.n252 CSoutput.n204 4.5005
R23948 CSoutput.n253 CSoutput.n252 4.5005
R23949 CSoutput.n251 CSoutput.n136 4.5005
R23950 CSoutput.n152 CSoutput.n136 4.5005
R23951 CSoutput.n147 CSoutput.n131 4.5005
R23952 CSoutput.n147 CSoutput.n133 4.5005
R23953 CSoutput.n147 CSoutput.n130 4.5005
R23954 CSoutput.n147 CSoutput.n134 4.5005
R23955 CSoutput.n147 CSoutput.n129 4.5005
R23956 CSoutput.n147 CSoutput.t230 4.5005
R23957 CSoutput.n147 CSoutput.n128 4.5005
R23958 CSoutput.n147 CSoutput.n135 4.5005
R23959 CSoutput.n147 CSoutput.n136 4.5005
R23960 CSoutput.n145 CSoutput.n131 4.5005
R23961 CSoutput.n145 CSoutput.n133 4.5005
R23962 CSoutput.n145 CSoutput.n130 4.5005
R23963 CSoutput.n145 CSoutput.n134 4.5005
R23964 CSoutput.n145 CSoutput.n129 4.5005
R23965 CSoutput.n145 CSoutput.t230 4.5005
R23966 CSoutput.n145 CSoutput.n128 4.5005
R23967 CSoutput.n145 CSoutput.n135 4.5005
R23968 CSoutput.n145 CSoutput.n136 4.5005
R23969 CSoutput.n144 CSoutput.n131 4.5005
R23970 CSoutput.n144 CSoutput.n133 4.5005
R23971 CSoutput.n144 CSoutput.n130 4.5005
R23972 CSoutput.n144 CSoutput.n134 4.5005
R23973 CSoutput.n144 CSoutput.n129 4.5005
R23974 CSoutput.n144 CSoutput.t230 4.5005
R23975 CSoutput.n144 CSoutput.n128 4.5005
R23976 CSoutput.n144 CSoutput.n135 4.5005
R23977 CSoutput.n144 CSoutput.n136 4.5005
R23978 CSoutput.n273 CSoutput.n131 4.5005
R23979 CSoutput.n273 CSoutput.n133 4.5005
R23980 CSoutput.n273 CSoutput.n130 4.5005
R23981 CSoutput.n273 CSoutput.n134 4.5005
R23982 CSoutput.n273 CSoutput.n129 4.5005
R23983 CSoutput.n273 CSoutput.t230 4.5005
R23984 CSoutput.n273 CSoutput.n128 4.5005
R23985 CSoutput.n273 CSoutput.n135 4.5005
R23986 CSoutput.n273 CSoutput.n136 4.5005
R23987 CSoutput.n271 CSoutput.n131 4.5005
R23988 CSoutput.n271 CSoutput.n133 4.5005
R23989 CSoutput.n271 CSoutput.n130 4.5005
R23990 CSoutput.n271 CSoutput.n134 4.5005
R23991 CSoutput.n271 CSoutput.n129 4.5005
R23992 CSoutput.n271 CSoutput.t230 4.5005
R23993 CSoutput.n271 CSoutput.n128 4.5005
R23994 CSoutput.n271 CSoutput.n135 4.5005
R23995 CSoutput.n269 CSoutput.n131 4.5005
R23996 CSoutput.n269 CSoutput.n133 4.5005
R23997 CSoutput.n269 CSoutput.n130 4.5005
R23998 CSoutput.n269 CSoutput.n134 4.5005
R23999 CSoutput.n269 CSoutput.n129 4.5005
R24000 CSoutput.n269 CSoutput.t230 4.5005
R24001 CSoutput.n269 CSoutput.n128 4.5005
R24002 CSoutput.n269 CSoutput.n135 4.5005
R24003 CSoutput.n155 CSoutput.n131 4.5005
R24004 CSoutput.n155 CSoutput.n133 4.5005
R24005 CSoutput.n155 CSoutput.n130 4.5005
R24006 CSoutput.n155 CSoutput.n134 4.5005
R24007 CSoutput.n155 CSoutput.n129 4.5005
R24008 CSoutput.n155 CSoutput.t230 4.5005
R24009 CSoutput.n155 CSoutput.n128 4.5005
R24010 CSoutput.n155 CSoutput.n135 4.5005
R24011 CSoutput.n155 CSoutput.n136 4.5005
R24012 CSoutput.n154 CSoutput.n131 4.5005
R24013 CSoutput.n154 CSoutput.n133 4.5005
R24014 CSoutput.n154 CSoutput.n130 4.5005
R24015 CSoutput.n154 CSoutput.n134 4.5005
R24016 CSoutput.n154 CSoutput.n129 4.5005
R24017 CSoutput.n154 CSoutput.t230 4.5005
R24018 CSoutput.n154 CSoutput.n128 4.5005
R24019 CSoutput.n154 CSoutput.n135 4.5005
R24020 CSoutput.n154 CSoutput.n136 4.5005
R24021 CSoutput.n158 CSoutput.n131 4.5005
R24022 CSoutput.n158 CSoutput.n133 4.5005
R24023 CSoutput.n158 CSoutput.n130 4.5005
R24024 CSoutput.n158 CSoutput.n134 4.5005
R24025 CSoutput.n158 CSoutput.n129 4.5005
R24026 CSoutput.n158 CSoutput.t230 4.5005
R24027 CSoutput.n158 CSoutput.n128 4.5005
R24028 CSoutput.n158 CSoutput.n135 4.5005
R24029 CSoutput.n158 CSoutput.n136 4.5005
R24030 CSoutput.n157 CSoutput.n131 4.5005
R24031 CSoutput.n157 CSoutput.n133 4.5005
R24032 CSoutput.n157 CSoutput.n130 4.5005
R24033 CSoutput.n157 CSoutput.n134 4.5005
R24034 CSoutput.n157 CSoutput.n129 4.5005
R24035 CSoutput.n157 CSoutput.t230 4.5005
R24036 CSoutput.n157 CSoutput.n128 4.5005
R24037 CSoutput.n157 CSoutput.n135 4.5005
R24038 CSoutput.n157 CSoutput.n136 4.5005
R24039 CSoutput.n140 CSoutput.n131 4.5005
R24040 CSoutput.n140 CSoutput.n133 4.5005
R24041 CSoutput.n140 CSoutput.n130 4.5005
R24042 CSoutput.n140 CSoutput.n134 4.5005
R24043 CSoutput.n140 CSoutput.n129 4.5005
R24044 CSoutput.n140 CSoutput.t230 4.5005
R24045 CSoutput.n140 CSoutput.n128 4.5005
R24046 CSoutput.n140 CSoutput.n135 4.5005
R24047 CSoutput.n140 CSoutput.n136 4.5005
R24048 CSoutput.n276 CSoutput.n131 4.5005
R24049 CSoutput.n276 CSoutput.n133 4.5005
R24050 CSoutput.n276 CSoutput.n130 4.5005
R24051 CSoutput.n276 CSoutput.n134 4.5005
R24052 CSoutput.n276 CSoutput.n129 4.5005
R24053 CSoutput.n276 CSoutput.t230 4.5005
R24054 CSoutput.n276 CSoutput.n128 4.5005
R24055 CSoutput.n276 CSoutput.n135 4.5005
R24056 CSoutput.n276 CSoutput.n136 4.5005
R24057 CSoutput.n323 CSoutput.n307 4.10845
R24058 CSoutput.n125 CSoutput.n109 4.10845
R24059 CSoutput.n321 CSoutput.t89 4.06363
R24060 CSoutput.n321 CSoutput.t19 4.06363
R24061 CSoutput.n319 CSoutput.t35 4.06363
R24062 CSoutput.n319 CSoutput.t59 4.06363
R24063 CSoutput.n317 CSoutput.t71 4.06363
R24064 CSoutput.n317 CSoutput.t6 4.06363
R24065 CSoutput.n315 CSoutput.t2 4.06363
R24066 CSoutput.n315 CSoutput.t37 4.06363
R24067 CSoutput.n313 CSoutput.t53 4.06363
R24068 CSoutput.n313 CSoutput.t73 4.06363
R24069 CSoutput.n311 CSoutput.t86 4.06363
R24070 CSoutput.n311 CSoutput.t16 4.06363
R24071 CSoutput.n309 CSoutput.t22 4.06363
R24072 CSoutput.n309 CSoutput.t74 4.06363
R24073 CSoutput.n308 CSoutput.t88 4.06363
R24074 CSoutput.n308 CSoutput.t90 4.06363
R24075 CSoutput.n305 CSoutput.t81 4.06363
R24076 CSoutput.n305 CSoutput.t7 4.06363
R24077 CSoutput.n303 CSoutput.t23 4.06363
R24078 CSoutput.n303 CSoutput.t51 4.06363
R24079 CSoutput.n301 CSoutput.t64 4.06363
R24080 CSoutput.n301 CSoutput.t94 4.06363
R24081 CSoutput.n299 CSoutput.t87 4.06363
R24082 CSoutput.n299 CSoutput.t28 4.06363
R24083 CSoutput.n297 CSoutput.t41 4.06363
R24084 CSoutput.n297 CSoutput.t65 4.06363
R24085 CSoutput.n295 CSoutput.t75 4.06363
R24086 CSoutput.n295 CSoutput.t5 4.06363
R24087 CSoutput.n293 CSoutput.t8 4.06363
R24088 CSoutput.n293 CSoutput.t68 4.06363
R24089 CSoutput.n292 CSoutput.t80 4.06363
R24090 CSoutput.n292 CSoutput.t82 4.06363
R24091 CSoutput.n290 CSoutput.t91 4.06363
R24092 CSoutput.n290 CSoutput.t52 4.06363
R24093 CSoutput.n288 CSoutput.t78 4.06363
R24094 CSoutput.n288 CSoutput.t38 4.06363
R24095 CSoutput.n286 CSoutput.t66 4.06363
R24096 CSoutput.n286 CSoutput.t26 4.06363
R24097 CSoutput.n284 CSoutput.t84 4.06363
R24098 CSoutput.n284 CSoutput.t45 4.06363
R24099 CSoutput.n282 CSoutput.t72 4.06363
R24100 CSoutput.n282 CSoutput.t33 4.06363
R24101 CSoutput.n280 CSoutput.t61 4.06363
R24102 CSoutput.n280 CSoutput.t15 4.06363
R24103 CSoutput.n278 CSoutput.t76 4.06363
R24104 CSoutput.n278 CSoutput.t10 4.06363
R24105 CSoutput.n277 CSoutput.t42 4.06363
R24106 CSoutput.n277 CSoutput.t24 4.06363
R24107 CSoutput.n110 CSoutput.t57 4.06363
R24108 CSoutput.n110 CSoutput.t32 4.06363
R24109 CSoutput.n111 CSoutput.t14 4.06363
R24110 CSoutput.n111 CSoutput.t58 4.06363
R24111 CSoutput.n113 CSoutput.t55 4.06363
R24112 CSoutput.n113 CSoutput.t29 4.06363
R24113 CSoutput.n115 CSoutput.t13 4.06363
R24114 CSoutput.n115 CSoutput.t12 4.06363
R24115 CSoutput.n117 CSoutput.t70 4.06363
R24116 CSoutput.n117 CSoutput.t40 4.06363
R24117 CSoutput.n119 CSoutput.t36 4.06363
R24118 CSoutput.n119 CSoutput.t9 4.06363
R24119 CSoutput.n121 CSoutput.t93 4.06363
R24120 CSoutput.n121 CSoutput.t69 4.06363
R24121 CSoutput.n123 CSoutput.t56 4.06363
R24122 CSoutput.n123 CSoutput.t31 4.06363
R24123 CSoutput.n94 CSoutput.t47 4.06363
R24124 CSoutput.n94 CSoutput.t20 4.06363
R24125 CSoutput.n95 CSoutput.t4 4.06363
R24126 CSoutput.n95 CSoutput.t49 4.06363
R24127 CSoutput.n97 CSoutput.t44 4.06363
R24128 CSoutput.n97 CSoutput.t17 4.06363
R24129 CSoutput.n99 CSoutput.t3 4.06363
R24130 CSoutput.n99 CSoutput.t1 4.06363
R24131 CSoutput.n101 CSoutput.t63 4.06363
R24132 CSoutput.n101 CSoutput.t30 4.06363
R24133 CSoutput.n103 CSoutput.t27 4.06363
R24134 CSoutput.n103 CSoutput.t0 4.06363
R24135 CSoutput.n105 CSoutput.t83 4.06363
R24136 CSoutput.n105 CSoutput.t60 4.06363
R24137 CSoutput.n107 CSoutput.t48 4.06363
R24138 CSoutput.n107 CSoutput.t21 4.06363
R24139 CSoutput.n79 CSoutput.t95 4.06363
R24140 CSoutput.n79 CSoutput.t43 4.06363
R24141 CSoutput.n80 CSoutput.t11 4.06363
R24142 CSoutput.n80 CSoutput.t77 4.06363
R24143 CSoutput.n82 CSoutput.t18 4.06363
R24144 CSoutput.n82 CSoutput.t62 4.06363
R24145 CSoutput.n84 CSoutput.t34 4.06363
R24146 CSoutput.n84 CSoutput.t50 4.06363
R24147 CSoutput.n86 CSoutput.t46 4.06363
R24148 CSoutput.n86 CSoutput.t85 4.06363
R24149 CSoutput.n88 CSoutput.t25 4.06363
R24150 CSoutput.n88 CSoutput.t67 4.06363
R24151 CSoutput.n90 CSoutput.t39 4.06363
R24152 CSoutput.n90 CSoutput.t79 4.06363
R24153 CSoutput.n92 CSoutput.t54 4.06363
R24154 CSoutput.n92 CSoutput.t92 4.06363
R24155 CSoutput.n44 CSoutput.n43 3.79402
R24156 CSoutput.n49 CSoutput.n48 3.79402
R24157 CSoutput.n383 CSoutput.n363 3.72967
R24158 CSoutput.n443 CSoutput.n423 3.72967
R24159 CSoutput.n445 CSoutput.n444 3.57343
R24160 CSoutput.n444 CSoutput.n384 3.42304
R24161 CSoutput.n324 CSoutput.n126 2.99158
R24162 CSoutput.n381 CSoutput.t145 2.82907
R24163 CSoutput.n381 CSoutput.t111 2.82907
R24164 CSoutput.n379 CSoutput.t96 2.82907
R24165 CSoutput.n379 CSoutput.t140 2.82907
R24166 CSoutput.n377 CSoutput.t130 2.82907
R24167 CSoutput.n377 CSoutput.t120 2.82907
R24168 CSoutput.n375 CSoutput.t108 2.82907
R24169 CSoutput.n375 CSoutput.t199 2.82907
R24170 CSoutput.n373 CSoutput.t123 2.82907
R24171 CSoutput.n373 CSoutput.t127 2.82907
R24172 CSoutput.n371 CSoutput.t122 2.82907
R24173 CSoutput.n371 CSoutput.t215 2.82907
R24174 CSoutput.n369 CSoutput.t146 2.82907
R24175 CSoutput.n369 CSoutput.t113 2.82907
R24176 CSoutput.n367 CSoutput.t101 2.82907
R24177 CSoutput.n367 CSoutput.t185 2.82907
R24178 CSoutput.n365 CSoutput.t132 2.82907
R24179 CSoutput.n365 CSoutput.t138 2.82907
R24180 CSoutput.n364 CSoutput.t112 2.82907
R24181 CSoutput.n364 CSoutput.t203 2.82907
R24182 CSoutput.n361 CSoutput.t148 2.82907
R24183 CSoutput.n361 CSoutput.t161 2.82907
R24184 CSoutput.n359 CSoutput.t166 2.82907
R24185 CSoutput.n359 CSoutput.t170 2.82907
R24186 CSoutput.n357 CSoutput.t181 2.82907
R24187 CSoutput.n357 CSoutput.t156 2.82907
R24188 CSoutput.n355 CSoutput.t157 2.82907
R24189 CSoutput.n355 CSoutput.t165 2.82907
R24190 CSoutput.n353 CSoutput.t100 2.82907
R24191 CSoutput.n353 CSoutput.t182 2.82907
R24192 CSoutput.n351 CSoutput.t180 2.82907
R24193 CSoutput.n351 CSoutput.t154 2.82907
R24194 CSoutput.n349 CSoutput.t201 2.82907
R24195 CSoutput.n349 CSoutput.t98 2.82907
R24196 CSoutput.n347 CSoutput.t99 2.82907
R24197 CSoutput.n347 CSoutput.t190 2.82907
R24198 CSoutput.n345 CSoutput.t109 2.82907
R24199 CSoutput.n345 CSoutput.t200 2.82907
R24200 CSoutput.n344 CSoutput.t207 2.82907
R24201 CSoutput.n344 CSoutput.t97 2.82907
R24202 CSoutput.n342 CSoutput.t211 2.82907
R24203 CSoutput.n342 CSoutput.t155 2.82907
R24204 CSoutput.n340 CSoutput.t184 2.82907
R24205 CSoutput.n340 CSoutput.t195 2.82907
R24206 CSoutput.n338 CSoutput.t105 2.82907
R24207 CSoutput.n338 CSoutput.t131 2.82907
R24208 CSoutput.n336 CSoutput.t119 2.82907
R24209 CSoutput.n336 CSoutput.t151 2.82907
R24210 CSoutput.n334 CSoutput.t164 2.82907
R24211 CSoutput.n334 CSoutput.t178 2.82907
R24212 CSoutput.n332 CSoutput.t147 2.82907
R24213 CSoutput.n332 CSoutput.t202 2.82907
R24214 CSoutput.n330 CSoutput.t171 2.82907
R24215 CSoutput.n330 CSoutput.t137 2.82907
R24216 CSoutput.n328 CSoutput.t124 2.82907
R24217 CSoutput.n328 CSoutput.t150 2.82907
R24218 CSoutput.n326 CSoutput.t134 2.82907
R24219 CSoutput.n326 CSoutput.t143 2.82907
R24220 CSoutput.n325 CSoutput.t144 2.82907
R24221 CSoutput.n325 CSoutput.t212 2.82907
R24222 CSoutput.n424 CSoutput.t162 2.82907
R24223 CSoutput.n424 CSoutput.t194 2.82907
R24224 CSoutput.n425 CSoutput.t125 2.82907
R24225 CSoutput.n425 CSoutput.t142 2.82907
R24226 CSoutput.n427 CSoutput.t152 2.82907
R24227 CSoutput.n427 CSoutput.t173 2.82907
R24228 CSoutput.n429 CSoutput.t196 2.82907
R24229 CSoutput.n429 CSoutput.t158 2.82907
R24230 CSoutput.n431 CSoutput.t168 2.82907
R24231 CSoutput.n431 CSoutput.t208 2.82907
R24232 CSoutput.n433 CSoutput.t103 2.82907
R24233 CSoutput.n433 CSoutput.t128 2.82907
R24234 CSoutput.n435 CSoutput.t159 2.82907
R24235 CSoutput.n435 CSoutput.t188 2.82907
R24236 CSoutput.n437 CSoutput.t204 2.82907
R24237 CSoutput.n437 CSoutput.t114 2.82907
R24238 CSoutput.n439 CSoutput.t149 2.82907
R24239 CSoutput.n439 CSoutput.t169 2.82907
R24240 CSoutput.n441 CSoutput.t104 2.82907
R24241 CSoutput.n441 CSoutput.t139 2.82907
R24242 CSoutput.n404 CSoutput.t115 2.82907
R24243 CSoutput.n404 CSoutput.t106 2.82907
R24244 CSoutput.n405 CSoutput.t102 2.82907
R24245 CSoutput.n405 CSoutput.t213 2.82907
R24246 CSoutput.n407 CSoutput.t214 2.82907
R24247 CSoutput.n407 CSoutput.t116 2.82907
R24248 CSoutput.n409 CSoutput.t117 2.82907
R24249 CSoutput.n409 CSoutput.t174 2.82907
R24250 CSoutput.n411 CSoutput.t175 2.82907
R24251 CSoutput.n411 CSoutput.t206 2.82907
R24252 CSoutput.n413 CSoutput.t209 2.82907
R24253 CSoutput.n413 CSoutput.t198 2.82907
R24254 CSoutput.n415 CSoutput.t189 2.82907
R24255 CSoutput.n415 CSoutput.t176 2.82907
R24256 CSoutput.n417 CSoutput.t177 2.82907
R24257 CSoutput.n417 CSoutput.t210 2.82907
R24258 CSoutput.n419 CSoutput.t163 2.82907
R24259 CSoutput.n419 CSoutput.t191 2.82907
R24260 CSoutput.n421 CSoutput.t197 2.82907
R24261 CSoutput.n421 CSoutput.t172 2.82907
R24262 CSoutput.n385 CSoutput.t126 2.82907
R24263 CSoutput.n385 CSoutput.t183 2.82907
R24264 CSoutput.n386 CSoutput.t179 2.82907
R24265 CSoutput.n386 CSoutput.t153 2.82907
R24266 CSoutput.n388 CSoutput.t187 2.82907
R24267 CSoutput.n388 CSoutput.t141 2.82907
R24268 CSoutput.n390 CSoutput.t167 2.82907
R24269 CSoutput.n390 CSoutput.t205 2.82907
R24270 CSoutput.n392 CSoutput.t121 2.82907
R24271 CSoutput.n392 CSoutput.t186 2.82907
R24272 CSoutput.n394 CSoutput.t107 2.82907
R24273 CSoutput.n394 CSoutput.t193 2.82907
R24274 CSoutput.n396 CSoutput.t192 2.82907
R24275 CSoutput.n396 CSoutput.t133 2.82907
R24276 CSoutput.n398 CSoutput.t160 2.82907
R24277 CSoutput.n398 CSoutput.t129 2.82907
R24278 CSoutput.n400 CSoutput.t135 2.82907
R24279 CSoutput.n400 CSoutput.t110 2.82907
R24280 CSoutput.n402 CSoutput.t118 2.82907
R24281 CSoutput.n402 CSoutput.t136 2.82907
R24282 CSoutput.n75 CSoutput.n1 2.45513
R24283 CSoutput.n217 CSoutput.n215 2.251
R24284 CSoutput.n217 CSoutput.n214 2.251
R24285 CSoutput.n217 CSoutput.n213 2.251
R24286 CSoutput.n217 CSoutput.n212 2.251
R24287 CSoutput.n186 CSoutput.n185 2.251
R24288 CSoutput.n186 CSoutput.n184 2.251
R24289 CSoutput.n186 CSoutput.n183 2.251
R24290 CSoutput.n186 CSoutput.n182 2.251
R24291 CSoutput.n259 CSoutput.n258 2.251
R24292 CSoutput.n224 CSoutput.n222 2.251
R24293 CSoutput.n224 CSoutput.n221 2.251
R24294 CSoutput.n224 CSoutput.n220 2.251
R24295 CSoutput.n242 CSoutput.n224 2.251
R24296 CSoutput.n230 CSoutput.n229 2.251
R24297 CSoutput.n230 CSoutput.n228 2.251
R24298 CSoutput.n230 CSoutput.n227 2.251
R24299 CSoutput.n230 CSoutput.n226 2.251
R24300 CSoutput.n256 CSoutput.n196 2.251
R24301 CSoutput.n251 CSoutput.n249 2.251
R24302 CSoutput.n251 CSoutput.n248 2.251
R24303 CSoutput.n251 CSoutput.n247 2.251
R24304 CSoutput.n251 CSoutput.n246 2.251
R24305 CSoutput.n152 CSoutput.n151 2.251
R24306 CSoutput.n152 CSoutput.n150 2.251
R24307 CSoutput.n152 CSoutput.n149 2.251
R24308 CSoutput.n152 CSoutput.n148 2.251
R24309 CSoutput.n269 CSoutput.n268 2.251
R24310 CSoutput.n186 CSoutput.n166 2.2505
R24311 CSoutput.n181 CSoutput.n166 2.2505
R24312 CSoutput.n179 CSoutput.n166 2.2505
R24313 CSoutput.n178 CSoutput.n166 2.2505
R24314 CSoutput.n263 CSoutput.n166 2.2505
R24315 CSoutput.n261 CSoutput.n166 2.2505
R24316 CSoutput.n259 CSoutput.n166 2.2505
R24317 CSoutput.n189 CSoutput.n166 2.2505
R24318 CSoutput.n188 CSoutput.n166 2.2505
R24319 CSoutput.n192 CSoutput.n166 2.2505
R24320 CSoutput.n191 CSoutput.n166 2.2505
R24321 CSoutput.n174 CSoutput.n166 2.2505
R24322 CSoutput.n266 CSoutput.n166 2.2505
R24323 CSoutput.n266 CSoutput.n265 2.2505
R24324 CSoutput.n230 CSoutput.n201 2.2505
R24325 CSoutput.n211 CSoutput.n201 2.2505
R24326 CSoutput.n232 CSoutput.n201 2.2505
R24327 CSoutput.n210 CSoutput.n201 2.2505
R24328 CSoutput.n234 CSoutput.n201 2.2505
R24329 CSoutput.n201 CSoutput.n195 2.2505
R24330 CSoutput.n256 CSoutput.n201 2.2505
R24331 CSoutput.n254 CSoutput.n201 2.2505
R24332 CSoutput.n236 CSoutput.n201 2.2505
R24333 CSoutput.n208 CSoutput.n201 2.2505
R24334 CSoutput.n238 CSoutput.n201 2.2505
R24335 CSoutput.n207 CSoutput.n201 2.2505
R24336 CSoutput.n252 CSoutput.n201 2.2505
R24337 CSoutput.n252 CSoutput.n205 2.2505
R24338 CSoutput.n152 CSoutput.n132 2.2505
R24339 CSoutput.n147 CSoutput.n132 2.2505
R24340 CSoutput.n145 CSoutput.n132 2.2505
R24341 CSoutput.n144 CSoutput.n132 2.2505
R24342 CSoutput.n273 CSoutput.n132 2.2505
R24343 CSoutput.n271 CSoutput.n132 2.2505
R24344 CSoutput.n269 CSoutput.n132 2.2505
R24345 CSoutput.n155 CSoutput.n132 2.2505
R24346 CSoutput.n154 CSoutput.n132 2.2505
R24347 CSoutput.n158 CSoutput.n132 2.2505
R24348 CSoutput.n157 CSoutput.n132 2.2505
R24349 CSoutput.n140 CSoutput.n132 2.2505
R24350 CSoutput.n276 CSoutput.n132 2.2505
R24351 CSoutput.n276 CSoutput.n275 2.2505
R24352 CSoutput.n194 CSoutput.n187 2.25024
R24353 CSoutput.n194 CSoutput.n180 2.25024
R24354 CSoutput.n262 CSoutput.n194 2.25024
R24355 CSoutput.n194 CSoutput.n190 2.25024
R24356 CSoutput.n194 CSoutput.n193 2.25024
R24357 CSoutput.n194 CSoutput.n161 2.25024
R24358 CSoutput.n244 CSoutput.n241 2.25024
R24359 CSoutput.n244 CSoutput.n240 2.25024
R24360 CSoutput.n244 CSoutput.n239 2.25024
R24361 CSoutput.n244 CSoutput.n206 2.25024
R24362 CSoutput.n244 CSoutput.n243 2.25024
R24363 CSoutput.n245 CSoutput.n244 2.25024
R24364 CSoutput.n160 CSoutput.n153 2.25024
R24365 CSoutput.n160 CSoutput.n146 2.25024
R24366 CSoutput.n272 CSoutput.n160 2.25024
R24367 CSoutput.n160 CSoutput.n156 2.25024
R24368 CSoutput.n160 CSoutput.n159 2.25024
R24369 CSoutput.n160 CSoutput.n127 2.25024
R24370 CSoutput.n261 CSoutput.n171 1.50111
R24371 CSoutput.n209 CSoutput.n195 1.50111
R24372 CSoutput.n271 CSoutput.n137 1.50111
R24373 CSoutput.n217 CSoutput.n216 1.501
R24374 CSoutput.n224 CSoutput.n223 1.501
R24375 CSoutput.n251 CSoutput.n250 1.501
R24376 CSoutput.n265 CSoutput.n176 1.12536
R24377 CSoutput.n265 CSoutput.n177 1.12536
R24378 CSoutput.n265 CSoutput.n264 1.12536
R24379 CSoutput.n225 CSoutput.n205 1.12536
R24380 CSoutput.n231 CSoutput.n205 1.12536
R24381 CSoutput.n233 CSoutput.n205 1.12536
R24382 CSoutput.n275 CSoutput.n142 1.12536
R24383 CSoutput.n275 CSoutput.n143 1.12536
R24384 CSoutput.n275 CSoutput.n274 1.12536
R24385 CSoutput.n265 CSoutput.n172 1.12536
R24386 CSoutput.n265 CSoutput.n173 1.12536
R24387 CSoutput.n265 CSoutput.n175 1.12536
R24388 CSoutput.n255 CSoutput.n205 1.12536
R24389 CSoutput.n235 CSoutput.n205 1.12536
R24390 CSoutput.n237 CSoutput.n205 1.12536
R24391 CSoutput.n275 CSoutput.n138 1.12536
R24392 CSoutput.n275 CSoutput.n139 1.12536
R24393 CSoutput.n275 CSoutput.n141 1.12536
R24394 CSoutput.n31 CSoutput.n30 0.669944
R24395 CSoutput.n62 CSoutput.n61 0.669944
R24396 CSoutput.n368 CSoutput.n366 0.573776
R24397 CSoutput.n370 CSoutput.n368 0.573776
R24398 CSoutput.n372 CSoutput.n370 0.573776
R24399 CSoutput.n374 CSoutput.n372 0.573776
R24400 CSoutput.n376 CSoutput.n374 0.573776
R24401 CSoutput.n378 CSoutput.n376 0.573776
R24402 CSoutput.n380 CSoutput.n378 0.573776
R24403 CSoutput.n382 CSoutput.n380 0.573776
R24404 CSoutput.n348 CSoutput.n346 0.573776
R24405 CSoutput.n350 CSoutput.n348 0.573776
R24406 CSoutput.n352 CSoutput.n350 0.573776
R24407 CSoutput.n354 CSoutput.n352 0.573776
R24408 CSoutput.n356 CSoutput.n354 0.573776
R24409 CSoutput.n358 CSoutput.n356 0.573776
R24410 CSoutput.n360 CSoutput.n358 0.573776
R24411 CSoutput.n362 CSoutput.n360 0.573776
R24412 CSoutput.n329 CSoutput.n327 0.573776
R24413 CSoutput.n331 CSoutput.n329 0.573776
R24414 CSoutput.n333 CSoutput.n331 0.573776
R24415 CSoutput.n335 CSoutput.n333 0.573776
R24416 CSoutput.n337 CSoutput.n335 0.573776
R24417 CSoutput.n339 CSoutput.n337 0.573776
R24418 CSoutput.n341 CSoutput.n339 0.573776
R24419 CSoutput.n343 CSoutput.n341 0.573776
R24420 CSoutput.n442 CSoutput.n440 0.573776
R24421 CSoutput.n440 CSoutput.n438 0.573776
R24422 CSoutput.n438 CSoutput.n436 0.573776
R24423 CSoutput.n436 CSoutput.n434 0.573776
R24424 CSoutput.n434 CSoutput.n432 0.573776
R24425 CSoutput.n432 CSoutput.n430 0.573776
R24426 CSoutput.n430 CSoutput.n428 0.573776
R24427 CSoutput.n428 CSoutput.n426 0.573776
R24428 CSoutput.n422 CSoutput.n420 0.573776
R24429 CSoutput.n420 CSoutput.n418 0.573776
R24430 CSoutput.n418 CSoutput.n416 0.573776
R24431 CSoutput.n416 CSoutput.n414 0.573776
R24432 CSoutput.n414 CSoutput.n412 0.573776
R24433 CSoutput.n412 CSoutput.n410 0.573776
R24434 CSoutput.n410 CSoutput.n408 0.573776
R24435 CSoutput.n408 CSoutput.n406 0.573776
R24436 CSoutput.n403 CSoutput.n401 0.573776
R24437 CSoutput.n401 CSoutput.n399 0.573776
R24438 CSoutput.n399 CSoutput.n397 0.573776
R24439 CSoutput.n397 CSoutput.n395 0.573776
R24440 CSoutput.n395 CSoutput.n393 0.573776
R24441 CSoutput.n393 CSoutput.n391 0.573776
R24442 CSoutput.n391 CSoutput.n389 0.573776
R24443 CSoutput.n389 CSoutput.n387 0.573776
R24444 CSoutput.n445 CSoutput.n276 0.53442
R24445 CSoutput.n312 CSoutput.n310 0.358259
R24446 CSoutput.n314 CSoutput.n312 0.358259
R24447 CSoutput.n316 CSoutput.n314 0.358259
R24448 CSoutput.n318 CSoutput.n316 0.358259
R24449 CSoutput.n320 CSoutput.n318 0.358259
R24450 CSoutput.n322 CSoutput.n320 0.358259
R24451 CSoutput.n296 CSoutput.n294 0.358259
R24452 CSoutput.n298 CSoutput.n296 0.358259
R24453 CSoutput.n300 CSoutput.n298 0.358259
R24454 CSoutput.n302 CSoutput.n300 0.358259
R24455 CSoutput.n304 CSoutput.n302 0.358259
R24456 CSoutput.n306 CSoutput.n304 0.358259
R24457 CSoutput.n281 CSoutput.n279 0.358259
R24458 CSoutput.n283 CSoutput.n281 0.358259
R24459 CSoutput.n285 CSoutput.n283 0.358259
R24460 CSoutput.n287 CSoutput.n285 0.358259
R24461 CSoutput.n289 CSoutput.n287 0.358259
R24462 CSoutput.n291 CSoutput.n289 0.358259
R24463 CSoutput.n124 CSoutput.n122 0.358259
R24464 CSoutput.n122 CSoutput.n120 0.358259
R24465 CSoutput.n120 CSoutput.n118 0.358259
R24466 CSoutput.n118 CSoutput.n116 0.358259
R24467 CSoutput.n116 CSoutput.n114 0.358259
R24468 CSoutput.n114 CSoutput.n112 0.358259
R24469 CSoutput.n108 CSoutput.n106 0.358259
R24470 CSoutput.n106 CSoutput.n104 0.358259
R24471 CSoutput.n104 CSoutput.n102 0.358259
R24472 CSoutput.n102 CSoutput.n100 0.358259
R24473 CSoutput.n100 CSoutput.n98 0.358259
R24474 CSoutput.n98 CSoutput.n96 0.358259
R24475 CSoutput.n93 CSoutput.n91 0.358259
R24476 CSoutput.n91 CSoutput.n89 0.358259
R24477 CSoutput.n89 CSoutput.n87 0.358259
R24478 CSoutput.n87 CSoutput.n85 0.358259
R24479 CSoutput.n85 CSoutput.n83 0.358259
R24480 CSoutput.n83 CSoutput.n81 0.358259
R24481 CSoutput.n21 CSoutput.n20 0.169105
R24482 CSoutput.n21 CSoutput.n16 0.169105
R24483 CSoutput.n26 CSoutput.n16 0.169105
R24484 CSoutput.n27 CSoutput.n26 0.169105
R24485 CSoutput.n27 CSoutput.n14 0.169105
R24486 CSoutput.n32 CSoutput.n14 0.169105
R24487 CSoutput.n33 CSoutput.n32 0.169105
R24488 CSoutput.n34 CSoutput.n33 0.169105
R24489 CSoutput.n34 CSoutput.n12 0.169105
R24490 CSoutput.n39 CSoutput.n12 0.169105
R24491 CSoutput.n40 CSoutput.n39 0.169105
R24492 CSoutput.n40 CSoutput.n10 0.169105
R24493 CSoutput.n45 CSoutput.n10 0.169105
R24494 CSoutput.n46 CSoutput.n45 0.169105
R24495 CSoutput.n47 CSoutput.n46 0.169105
R24496 CSoutput.n47 CSoutput.n8 0.169105
R24497 CSoutput.n52 CSoutput.n8 0.169105
R24498 CSoutput.n53 CSoutput.n52 0.169105
R24499 CSoutput.n53 CSoutput.n6 0.169105
R24500 CSoutput.n58 CSoutput.n6 0.169105
R24501 CSoutput.n59 CSoutput.n58 0.169105
R24502 CSoutput.n60 CSoutput.n59 0.169105
R24503 CSoutput.n60 CSoutput.n4 0.169105
R24504 CSoutput.n66 CSoutput.n4 0.169105
R24505 CSoutput.n67 CSoutput.n66 0.169105
R24506 CSoutput.n68 CSoutput.n67 0.169105
R24507 CSoutput.n68 CSoutput.n2 0.169105
R24508 CSoutput.n73 CSoutput.n2 0.169105
R24509 CSoutput.n74 CSoutput.n73 0.169105
R24510 CSoutput.n74 CSoutput.n0 0.169105
R24511 CSoutput.n78 CSoutput.n0 0.169105
R24512 CSoutput.n219 CSoutput.n218 0.0910737
R24513 CSoutput.n270 CSoutput.n267 0.0723685
R24514 CSoutput.n224 CSoutput.n219 0.0522944
R24515 CSoutput.n267 CSoutput.n266 0.0499135
R24516 CSoutput.n218 CSoutput.n217 0.0499135
R24517 CSoutput.n252 CSoutput.n251 0.0464294
R24518 CSoutput.n260 CSoutput.n257 0.0391444
R24519 CSoutput.n219 CSoutput.t216 0.023435
R24520 CSoutput.n267 CSoutput.t219 0.02262
R24521 CSoutput.n218 CSoutput.t222 0.02262
R24522 CSoutput CSoutput.n445 0.0052
R24523 CSoutput.n189 CSoutput.n172 0.00365111
R24524 CSoutput.n192 CSoutput.n173 0.00365111
R24525 CSoutput.n175 CSoutput.n174 0.00365111
R24526 CSoutput.n217 CSoutput.n176 0.00365111
R24527 CSoutput.n181 CSoutput.n177 0.00365111
R24528 CSoutput.n264 CSoutput.n178 0.00365111
R24529 CSoutput.n255 CSoutput.n254 0.00365111
R24530 CSoutput.n235 CSoutput.n208 0.00365111
R24531 CSoutput.n237 CSoutput.n207 0.00365111
R24532 CSoutput.n225 CSoutput.n224 0.00365111
R24533 CSoutput.n231 CSoutput.n211 0.00365111
R24534 CSoutput.n233 CSoutput.n210 0.00365111
R24535 CSoutput.n155 CSoutput.n138 0.00365111
R24536 CSoutput.n158 CSoutput.n139 0.00365111
R24537 CSoutput.n141 CSoutput.n140 0.00365111
R24538 CSoutput.n251 CSoutput.n142 0.00365111
R24539 CSoutput.n147 CSoutput.n143 0.00365111
R24540 CSoutput.n274 CSoutput.n144 0.00365111
R24541 CSoutput.n186 CSoutput.n176 0.00340054
R24542 CSoutput.n179 CSoutput.n177 0.00340054
R24543 CSoutput.n264 CSoutput.n263 0.00340054
R24544 CSoutput.n259 CSoutput.n172 0.00340054
R24545 CSoutput.n188 CSoutput.n173 0.00340054
R24546 CSoutput.n191 CSoutput.n175 0.00340054
R24547 CSoutput.n230 CSoutput.n225 0.00340054
R24548 CSoutput.n232 CSoutput.n231 0.00340054
R24549 CSoutput.n234 CSoutput.n233 0.00340054
R24550 CSoutput.n256 CSoutput.n255 0.00340054
R24551 CSoutput.n236 CSoutput.n235 0.00340054
R24552 CSoutput.n238 CSoutput.n237 0.00340054
R24553 CSoutput.n152 CSoutput.n142 0.00340054
R24554 CSoutput.n145 CSoutput.n143 0.00340054
R24555 CSoutput.n274 CSoutput.n273 0.00340054
R24556 CSoutput.n269 CSoutput.n138 0.00340054
R24557 CSoutput.n154 CSoutput.n139 0.00340054
R24558 CSoutput.n157 CSoutput.n141 0.00340054
R24559 CSoutput.n187 CSoutput.n181 0.00252698
R24560 CSoutput.n180 CSoutput.n178 0.00252698
R24561 CSoutput.n262 CSoutput.n261 0.00252698
R24562 CSoutput.n190 CSoutput.n188 0.00252698
R24563 CSoutput.n193 CSoutput.n191 0.00252698
R24564 CSoutput.n266 CSoutput.n161 0.00252698
R24565 CSoutput.n187 CSoutput.n186 0.00252698
R24566 CSoutput.n180 CSoutput.n179 0.00252698
R24567 CSoutput.n263 CSoutput.n262 0.00252698
R24568 CSoutput.n190 CSoutput.n189 0.00252698
R24569 CSoutput.n193 CSoutput.n192 0.00252698
R24570 CSoutput.n174 CSoutput.n161 0.00252698
R24571 CSoutput.n241 CSoutput.n211 0.00252698
R24572 CSoutput.n240 CSoutput.n210 0.00252698
R24573 CSoutput.n239 CSoutput.n195 0.00252698
R24574 CSoutput.n236 CSoutput.n206 0.00252698
R24575 CSoutput.n243 CSoutput.n238 0.00252698
R24576 CSoutput.n252 CSoutput.n245 0.00252698
R24577 CSoutput.n241 CSoutput.n230 0.00252698
R24578 CSoutput.n240 CSoutput.n232 0.00252698
R24579 CSoutput.n239 CSoutput.n234 0.00252698
R24580 CSoutput.n254 CSoutput.n206 0.00252698
R24581 CSoutput.n243 CSoutput.n208 0.00252698
R24582 CSoutput.n245 CSoutput.n207 0.00252698
R24583 CSoutput.n153 CSoutput.n147 0.00252698
R24584 CSoutput.n146 CSoutput.n144 0.00252698
R24585 CSoutput.n272 CSoutput.n271 0.00252698
R24586 CSoutput.n156 CSoutput.n154 0.00252698
R24587 CSoutput.n159 CSoutput.n157 0.00252698
R24588 CSoutput.n276 CSoutput.n127 0.00252698
R24589 CSoutput.n153 CSoutput.n152 0.00252698
R24590 CSoutput.n146 CSoutput.n145 0.00252698
R24591 CSoutput.n273 CSoutput.n272 0.00252698
R24592 CSoutput.n156 CSoutput.n155 0.00252698
R24593 CSoutput.n159 CSoutput.n158 0.00252698
R24594 CSoutput.n140 CSoutput.n127 0.00252698
R24595 CSoutput.n261 CSoutput.n260 0.0020275
R24596 CSoutput.n260 CSoutput.n259 0.0020275
R24597 CSoutput.n257 CSoutput.n195 0.0020275
R24598 CSoutput.n257 CSoutput.n256 0.0020275
R24599 CSoutput.n271 CSoutput.n270 0.0020275
R24600 CSoutput.n270 CSoutput.n269 0.0020275
R24601 CSoutput.n171 CSoutput.n170 0.00166668
R24602 CSoutput.n253 CSoutput.n209 0.00166668
R24603 CSoutput.n137 CSoutput.n136 0.00166668
R24604 CSoutput.n275 CSoutput.n137 0.00133328
R24605 CSoutput.n209 CSoutput.n205 0.00133328
R24606 CSoutput.n265 CSoutput.n171 0.00133328
R24607 CSoutput.n268 CSoutput.n160 0.001
R24608 CSoutput.n246 CSoutput.n160 0.001
R24609 CSoutput.n148 CSoutput.n128 0.001
R24610 CSoutput.n247 CSoutput.n128 0.001
R24611 CSoutput.n149 CSoutput.n129 0.001
R24612 CSoutput.n248 CSoutput.n129 0.001
R24613 CSoutput.n150 CSoutput.n130 0.001
R24614 CSoutput.n249 CSoutput.n130 0.001
R24615 CSoutput.n151 CSoutput.n131 0.001
R24616 CSoutput.n250 CSoutput.n131 0.001
R24617 CSoutput.n244 CSoutput.n196 0.001
R24618 CSoutput.n244 CSoutput.n242 0.001
R24619 CSoutput.n226 CSoutput.n197 0.001
R24620 CSoutput.n220 CSoutput.n197 0.001
R24621 CSoutput.n227 CSoutput.n198 0.001
R24622 CSoutput.n221 CSoutput.n198 0.001
R24623 CSoutput.n228 CSoutput.n199 0.001
R24624 CSoutput.n222 CSoutput.n199 0.001
R24625 CSoutput.n229 CSoutput.n200 0.001
R24626 CSoutput.n223 CSoutput.n200 0.001
R24627 CSoutput.n258 CSoutput.n194 0.001
R24628 CSoutput.n212 CSoutput.n194 0.001
R24629 CSoutput.n182 CSoutput.n162 0.001
R24630 CSoutput.n213 CSoutput.n162 0.001
R24631 CSoutput.n183 CSoutput.n163 0.001
R24632 CSoutput.n214 CSoutput.n163 0.001
R24633 CSoutput.n184 CSoutput.n164 0.001
R24634 CSoutput.n215 CSoutput.n164 0.001
R24635 CSoutput.n185 CSoutput.n165 0.001
R24636 CSoutput.n216 CSoutput.n165 0.001
R24637 CSoutput.n216 CSoutput.n166 0.001
R24638 CSoutput.n215 CSoutput.n167 0.001
R24639 CSoutput.n214 CSoutput.n168 0.001
R24640 CSoutput.n213 CSoutput.t237 0.001
R24641 CSoutput.n212 CSoutput.n169 0.001
R24642 CSoutput.n185 CSoutput.n167 0.001
R24643 CSoutput.n184 CSoutput.n168 0.001
R24644 CSoutput.n183 CSoutput.t237 0.001
R24645 CSoutput.n182 CSoutput.n169 0.001
R24646 CSoutput.n258 CSoutput.n170 0.001
R24647 CSoutput.n223 CSoutput.n201 0.001
R24648 CSoutput.n222 CSoutput.n202 0.001
R24649 CSoutput.n221 CSoutput.n203 0.001
R24650 CSoutput.n220 CSoutput.t232 0.001
R24651 CSoutput.n242 CSoutput.n204 0.001
R24652 CSoutput.n229 CSoutput.n202 0.001
R24653 CSoutput.n228 CSoutput.n203 0.001
R24654 CSoutput.n227 CSoutput.t232 0.001
R24655 CSoutput.n226 CSoutput.n204 0.001
R24656 CSoutput.n253 CSoutput.n196 0.001
R24657 CSoutput.n250 CSoutput.n132 0.001
R24658 CSoutput.n249 CSoutput.n133 0.001
R24659 CSoutput.n248 CSoutput.n134 0.001
R24660 CSoutput.n247 CSoutput.t230 0.001
R24661 CSoutput.n246 CSoutput.n135 0.001
R24662 CSoutput.n151 CSoutput.n133 0.001
R24663 CSoutput.n150 CSoutput.n134 0.001
R24664 CSoutput.n149 CSoutput.t230 0.001
R24665 CSoutput.n148 CSoutput.n135 0.001
R24666 CSoutput.n268 CSoutput.n136 0.001
R24667 a_n2982_8322.n12 a_n2982_8322.t27 74.6477
R24668 a_n2982_8322.n1 a_n2982_8322.t6 74.6477
R24669 a_n2982_8322.n28 a_n2982_8322.t21 74.6474
R24670 a_n2982_8322.n20 a_n2982_8322.t1 74.2899
R24671 a_n2982_8322.n13 a_n2982_8322.t25 74.2899
R24672 a_n2982_8322.n14 a_n2982_8322.t28 74.2899
R24673 a_n2982_8322.n17 a_n2982_8322.t29 74.2899
R24674 a_n2982_8322.n10 a_n2982_8322.t0 74.2899
R24675 a_n2982_8322.n28 a_n2982_8322.n27 70.6783
R24676 a_n2982_8322.n26 a_n2982_8322.n25 70.6783
R24677 a_n2982_8322.n24 a_n2982_8322.n23 70.6783
R24678 a_n2982_8322.n22 a_n2982_8322.n21 70.6783
R24679 a_n2982_8322.n12 a_n2982_8322.n11 70.6783
R24680 a_n2982_8322.n16 a_n2982_8322.n15 70.6783
R24681 a_n2982_8322.n1 a_n2982_8322.n0 70.6783
R24682 a_n2982_8322.n3 a_n2982_8322.n2 70.6783
R24683 a_n2982_8322.n5 a_n2982_8322.n4 70.6783
R24684 a_n2982_8322.n7 a_n2982_8322.n6 70.6783
R24685 a_n2982_8322.n9 a_n2982_8322.n8 70.6783
R24686 a_n2982_8322.n30 a_n2982_8322.n29 70.6782
R24687 a_n2982_8322.n18 a_n2982_8322.n10 24.9022
R24688 a_n2982_8322.n19 a_n2982_8322.t37 9.81851
R24689 a_n2982_8322.n18 a_n2982_8322.n17 8.38735
R24690 a_n2982_8322.n20 a_n2982_8322.n19 6.90998
R24691 a_n2982_8322.n19 a_n2982_8322.n18 5.3452
R24692 a_n2982_8322.n27 a_n2982_8322.t14 3.61217
R24693 a_n2982_8322.n27 a_n2982_8322.t10 3.61217
R24694 a_n2982_8322.n25 a_n2982_8322.t20 3.61217
R24695 a_n2982_8322.n25 a_n2982_8322.t8 3.61217
R24696 a_n2982_8322.n23 a_n2982_8322.t5 3.61217
R24697 a_n2982_8322.n23 a_n2982_8322.t4 3.61217
R24698 a_n2982_8322.n21 a_n2982_8322.t18 3.61217
R24699 a_n2982_8322.n21 a_n2982_8322.t17 3.61217
R24700 a_n2982_8322.n11 a_n2982_8322.t31 3.61217
R24701 a_n2982_8322.n11 a_n2982_8322.t30 3.61217
R24702 a_n2982_8322.n15 a_n2982_8322.t26 3.61217
R24703 a_n2982_8322.n15 a_n2982_8322.t24 3.61217
R24704 a_n2982_8322.n0 a_n2982_8322.t19 3.61217
R24705 a_n2982_8322.n0 a_n2982_8322.t15 3.61217
R24706 a_n2982_8322.n2 a_n2982_8322.t22 3.61217
R24707 a_n2982_8322.n2 a_n2982_8322.t12 3.61217
R24708 a_n2982_8322.n4 a_n2982_8322.t3 3.61217
R24709 a_n2982_8322.n4 a_n2982_8322.t2 3.61217
R24710 a_n2982_8322.n6 a_n2982_8322.t16 3.61217
R24711 a_n2982_8322.n6 a_n2982_8322.t9 3.61217
R24712 a_n2982_8322.n8 a_n2982_8322.t13 3.61217
R24713 a_n2982_8322.n8 a_n2982_8322.t11 3.61217
R24714 a_n2982_8322.n30 a_n2982_8322.t7 3.61217
R24715 a_n2982_8322.t23 a_n2982_8322.n30 3.61217
R24716 a_n2982_8322.n17 a_n2982_8322.n16 0.358259
R24717 a_n2982_8322.n16 a_n2982_8322.n14 0.358259
R24718 a_n2982_8322.n13 a_n2982_8322.n12 0.358259
R24719 a_n2982_8322.n10 a_n2982_8322.n9 0.358259
R24720 a_n2982_8322.n9 a_n2982_8322.n7 0.358259
R24721 a_n2982_8322.n7 a_n2982_8322.n5 0.358259
R24722 a_n2982_8322.n5 a_n2982_8322.n3 0.358259
R24723 a_n2982_8322.n3 a_n2982_8322.n1 0.358259
R24724 a_n2982_8322.n22 a_n2982_8322.n20 0.358259
R24725 a_n2982_8322.n24 a_n2982_8322.n22 0.358259
R24726 a_n2982_8322.n26 a_n2982_8322.n24 0.358259
R24727 a_n2982_8322.n29 a_n2982_8322.n26 0.358259
R24728 a_n2982_8322.n29 a_n2982_8322.n28 0.358259
R24729 a_n2982_8322.n14 a_n2982_8322.n13 0.101793
R24730 a_n2982_8322.t36 a_n2982_8322.t34 0.0788333
R24731 a_n2982_8322.t32 a_n2982_8322.t33 0.0788333
R24732 a_n2982_8322.t37 a_n2982_8322.t35 0.0788333
R24733 a_n2982_8322.t32 a_n2982_8322.t36 0.0318333
R24734 a_n2982_8322.t37 a_n2982_8322.t33 0.0318333
R24735 a_n2982_8322.t34 a_n2982_8322.t33 0.0318333
R24736 a_n2982_8322.t35 a_n2982_8322.t32 0.0318333
R24737 output.n41 output.n15 289.615
R24738 output.n72 output.n46 289.615
R24739 output.n104 output.n78 289.615
R24740 output.n136 output.n110 289.615
R24741 output.n77 output.n45 197.26
R24742 output.n77 output.n76 196.298
R24743 output.n109 output.n108 196.298
R24744 output.n141 output.n140 196.298
R24745 output.n42 output.n41 185
R24746 output.n40 output.n39 185
R24747 output.n19 output.n18 185
R24748 output.n34 output.n33 185
R24749 output.n32 output.n31 185
R24750 output.n23 output.n22 185
R24751 output.n26 output.n25 185
R24752 output.n73 output.n72 185
R24753 output.n71 output.n70 185
R24754 output.n50 output.n49 185
R24755 output.n65 output.n64 185
R24756 output.n63 output.n62 185
R24757 output.n54 output.n53 185
R24758 output.n57 output.n56 185
R24759 output.n105 output.n104 185
R24760 output.n103 output.n102 185
R24761 output.n82 output.n81 185
R24762 output.n97 output.n96 185
R24763 output.n95 output.n94 185
R24764 output.n86 output.n85 185
R24765 output.n89 output.n88 185
R24766 output.n137 output.n136 185
R24767 output.n135 output.n134 185
R24768 output.n114 output.n113 185
R24769 output.n129 output.n128 185
R24770 output.n127 output.n126 185
R24771 output.n118 output.n117 185
R24772 output.n121 output.n120 185
R24773 output.t1 output.n24 147.661
R24774 output.t19 output.n55 147.661
R24775 output.t0 output.n87 147.661
R24776 output.t2 output.n119 147.661
R24777 output.n41 output.n40 104.615
R24778 output.n40 output.n18 104.615
R24779 output.n33 output.n18 104.615
R24780 output.n33 output.n32 104.615
R24781 output.n32 output.n22 104.615
R24782 output.n25 output.n22 104.615
R24783 output.n72 output.n71 104.615
R24784 output.n71 output.n49 104.615
R24785 output.n64 output.n49 104.615
R24786 output.n64 output.n63 104.615
R24787 output.n63 output.n53 104.615
R24788 output.n56 output.n53 104.615
R24789 output.n104 output.n103 104.615
R24790 output.n103 output.n81 104.615
R24791 output.n96 output.n81 104.615
R24792 output.n96 output.n95 104.615
R24793 output.n95 output.n85 104.615
R24794 output.n88 output.n85 104.615
R24795 output.n136 output.n135 104.615
R24796 output.n135 output.n113 104.615
R24797 output.n128 output.n113 104.615
R24798 output.n128 output.n127 104.615
R24799 output.n127 output.n117 104.615
R24800 output.n120 output.n117 104.615
R24801 output.n1 output.t3 77.056
R24802 output.n14 output.t4 76.6694
R24803 output.n1 output.n0 72.7095
R24804 output.n3 output.n2 72.7095
R24805 output.n5 output.n4 72.7095
R24806 output.n7 output.n6 72.7095
R24807 output.n9 output.n8 72.7095
R24808 output.n11 output.n10 72.7095
R24809 output.n13 output.n12 72.7095
R24810 output.n25 output.t1 52.3082
R24811 output.n56 output.t19 52.3082
R24812 output.n88 output.t0 52.3082
R24813 output.n120 output.t2 52.3082
R24814 output.n26 output.n24 15.6674
R24815 output.n57 output.n55 15.6674
R24816 output.n89 output.n87 15.6674
R24817 output.n121 output.n119 15.6674
R24818 output.n27 output.n23 12.8005
R24819 output.n58 output.n54 12.8005
R24820 output.n90 output.n86 12.8005
R24821 output.n122 output.n118 12.8005
R24822 output.n31 output.n30 12.0247
R24823 output.n62 output.n61 12.0247
R24824 output.n94 output.n93 12.0247
R24825 output.n126 output.n125 12.0247
R24826 output.n34 output.n21 11.249
R24827 output.n65 output.n52 11.249
R24828 output.n97 output.n84 11.249
R24829 output.n129 output.n116 11.249
R24830 output.n35 output.n19 10.4732
R24831 output.n66 output.n50 10.4732
R24832 output.n98 output.n82 10.4732
R24833 output.n130 output.n114 10.4732
R24834 output.n39 output.n38 9.69747
R24835 output.n70 output.n69 9.69747
R24836 output.n102 output.n101 9.69747
R24837 output.n134 output.n133 9.69747
R24838 output.n45 output.n44 9.45567
R24839 output.n76 output.n75 9.45567
R24840 output.n108 output.n107 9.45567
R24841 output.n140 output.n139 9.45567
R24842 output.n44 output.n43 9.3005
R24843 output.n17 output.n16 9.3005
R24844 output.n38 output.n37 9.3005
R24845 output.n36 output.n35 9.3005
R24846 output.n21 output.n20 9.3005
R24847 output.n30 output.n29 9.3005
R24848 output.n28 output.n27 9.3005
R24849 output.n75 output.n74 9.3005
R24850 output.n48 output.n47 9.3005
R24851 output.n69 output.n68 9.3005
R24852 output.n67 output.n66 9.3005
R24853 output.n52 output.n51 9.3005
R24854 output.n61 output.n60 9.3005
R24855 output.n59 output.n58 9.3005
R24856 output.n107 output.n106 9.3005
R24857 output.n80 output.n79 9.3005
R24858 output.n101 output.n100 9.3005
R24859 output.n99 output.n98 9.3005
R24860 output.n84 output.n83 9.3005
R24861 output.n93 output.n92 9.3005
R24862 output.n91 output.n90 9.3005
R24863 output.n139 output.n138 9.3005
R24864 output.n112 output.n111 9.3005
R24865 output.n133 output.n132 9.3005
R24866 output.n131 output.n130 9.3005
R24867 output.n116 output.n115 9.3005
R24868 output.n125 output.n124 9.3005
R24869 output.n123 output.n122 9.3005
R24870 output.n42 output.n17 8.92171
R24871 output.n73 output.n48 8.92171
R24872 output.n105 output.n80 8.92171
R24873 output.n137 output.n112 8.92171
R24874 output output.n141 8.15037
R24875 output.n43 output.n15 8.14595
R24876 output.n74 output.n46 8.14595
R24877 output.n106 output.n78 8.14595
R24878 output.n138 output.n110 8.14595
R24879 output.n45 output.n15 5.81868
R24880 output.n76 output.n46 5.81868
R24881 output.n108 output.n78 5.81868
R24882 output.n140 output.n110 5.81868
R24883 output.n43 output.n42 5.04292
R24884 output.n74 output.n73 5.04292
R24885 output.n106 output.n105 5.04292
R24886 output.n138 output.n137 5.04292
R24887 output.n28 output.n24 4.38594
R24888 output.n59 output.n55 4.38594
R24889 output.n91 output.n87 4.38594
R24890 output.n123 output.n119 4.38594
R24891 output.n39 output.n17 4.26717
R24892 output.n70 output.n48 4.26717
R24893 output.n102 output.n80 4.26717
R24894 output.n134 output.n112 4.26717
R24895 output.n0 output.t13 3.9605
R24896 output.n0 output.t11 3.9605
R24897 output.n2 output.t18 3.9605
R24898 output.n2 output.t5 3.9605
R24899 output.n4 output.t7 3.9605
R24900 output.n4 output.t15 3.9605
R24901 output.n6 output.t17 3.9605
R24902 output.n6 output.t8 3.9605
R24903 output.n8 output.t9 3.9605
R24904 output.n8 output.t14 3.9605
R24905 output.n10 output.t16 3.9605
R24906 output.n10 output.t6 3.9605
R24907 output.n12 output.t12 3.9605
R24908 output.n12 output.t10 3.9605
R24909 output.n38 output.n19 3.49141
R24910 output.n69 output.n50 3.49141
R24911 output.n101 output.n82 3.49141
R24912 output.n133 output.n114 3.49141
R24913 output.n35 output.n34 2.71565
R24914 output.n66 output.n65 2.71565
R24915 output.n98 output.n97 2.71565
R24916 output.n130 output.n129 2.71565
R24917 output.n31 output.n21 1.93989
R24918 output.n62 output.n52 1.93989
R24919 output.n94 output.n84 1.93989
R24920 output.n126 output.n116 1.93989
R24921 output.n30 output.n23 1.16414
R24922 output.n61 output.n54 1.16414
R24923 output.n93 output.n86 1.16414
R24924 output.n125 output.n118 1.16414
R24925 output.n141 output.n109 0.962709
R24926 output.n109 output.n77 0.962709
R24927 output.n27 output.n26 0.388379
R24928 output.n58 output.n57 0.388379
R24929 output.n90 output.n89 0.388379
R24930 output.n122 output.n121 0.388379
R24931 output.n14 output.n13 0.387128
R24932 output.n13 output.n11 0.387128
R24933 output.n11 output.n9 0.387128
R24934 output.n9 output.n7 0.387128
R24935 output.n7 output.n5 0.387128
R24936 output.n5 output.n3 0.387128
R24937 output.n3 output.n1 0.387128
R24938 output.n44 output.n16 0.155672
R24939 output.n37 output.n16 0.155672
R24940 output.n37 output.n36 0.155672
R24941 output.n36 output.n20 0.155672
R24942 output.n29 output.n20 0.155672
R24943 output.n29 output.n28 0.155672
R24944 output.n75 output.n47 0.155672
R24945 output.n68 output.n47 0.155672
R24946 output.n68 output.n67 0.155672
R24947 output.n67 output.n51 0.155672
R24948 output.n60 output.n51 0.155672
R24949 output.n60 output.n59 0.155672
R24950 output.n107 output.n79 0.155672
R24951 output.n100 output.n79 0.155672
R24952 output.n100 output.n99 0.155672
R24953 output.n99 output.n83 0.155672
R24954 output.n92 output.n83 0.155672
R24955 output.n92 output.n91 0.155672
R24956 output.n139 output.n111 0.155672
R24957 output.n132 output.n111 0.155672
R24958 output.n132 output.n131 0.155672
R24959 output.n131 output.n115 0.155672
R24960 output.n124 output.n115 0.155672
R24961 output.n124 output.n123 0.155672
R24962 output output.n14 0.126227
R24963 minus.n33 minus.t20 321.495
R24964 minus.n7 minus.t6 321.495
R24965 minus.n50 minus.t18 297.12
R24966 minus.n48 minus.t15 297.12
R24967 minus.n28 minus.t16 297.12
R24968 minus.n42 minus.t11 297.12
R24969 minus.n30 minus.t12 297.12
R24970 minus.n36 minus.t7 297.12
R24971 minus.n32 minus.t19 297.12
R24972 minus.n6 minus.t5 297.12
R24973 minus.n10 minus.t9 297.12
R24974 minus.n12 minus.t8 297.12
R24975 minus.n16 minus.t10 297.12
R24976 minus.n18 minus.t14 297.12
R24977 minus.n22 minus.t13 297.12
R24978 minus.n24 minus.t17 297.12
R24979 minus.n56 minus.t4 243.255
R24980 minus.n55 minus.n53 224.169
R24981 minus.n55 minus.n54 223.454
R24982 minus.n35 minus.n34 161.3
R24983 minus.n36 minus.n31 161.3
R24984 minus.n38 minus.n37 161.3
R24985 minus.n39 minus.n30 161.3
R24986 minus.n41 minus.n40 161.3
R24987 minus.n42 minus.n29 161.3
R24988 minus.n44 minus.n43 161.3
R24989 minus.n45 minus.n28 161.3
R24990 minus.n47 minus.n46 161.3
R24991 minus.n48 minus.n27 161.3
R24992 minus.n49 minus.n26 161.3
R24993 minus.n51 minus.n50 161.3
R24994 minus.n25 minus.n24 161.3
R24995 minus.n23 minus.n0 161.3
R24996 minus.n22 minus.n21 161.3
R24997 minus.n20 minus.n1 161.3
R24998 minus.n19 minus.n18 161.3
R24999 minus.n17 minus.n2 161.3
R25000 minus.n16 minus.n15 161.3
R25001 minus.n14 minus.n3 161.3
R25002 minus.n13 minus.n12 161.3
R25003 minus.n11 minus.n4 161.3
R25004 minus.n10 minus.n9 161.3
R25005 minus.n8 minus.n5 161.3
R25006 minus.n8 minus.n7 44.9377
R25007 minus.n34 minus.n33 44.9377
R25008 minus.n50 minus.n49 37.246
R25009 minus.n24 minus.n23 37.246
R25010 minus.n48 minus.n47 32.8641
R25011 minus.n35 minus.n32 32.8641
R25012 minus.n6 minus.n5 32.8641
R25013 minus.n22 minus.n1 32.8641
R25014 minus.n52 minus.n51 30.2486
R25015 minus.n43 minus.n28 28.4823
R25016 minus.n37 minus.n36 28.4823
R25017 minus.n11 minus.n10 28.4823
R25018 minus.n18 minus.n17 28.4823
R25019 minus.n42 minus.n41 24.1005
R25020 minus.n41 minus.n30 24.1005
R25021 minus.n12 minus.n3 24.1005
R25022 minus.n16 minus.n3 24.1005
R25023 minus.n54 minus.t3 19.8005
R25024 minus.n54 minus.t2 19.8005
R25025 minus.n53 minus.t1 19.8005
R25026 minus.n53 minus.t0 19.8005
R25027 minus.n43 minus.n42 19.7187
R25028 minus.n37 minus.n30 19.7187
R25029 minus.n12 minus.n11 19.7187
R25030 minus.n17 minus.n16 19.7187
R25031 minus.n33 minus.n32 17.0522
R25032 minus.n7 minus.n6 17.0522
R25033 minus.n47 minus.n28 15.3369
R25034 minus.n36 minus.n35 15.3369
R25035 minus.n10 minus.n5 15.3369
R25036 minus.n18 minus.n1 15.3369
R25037 minus.n52 minus.n25 12.0706
R25038 minus minus.n57 12.0012
R25039 minus.n49 minus.n48 10.955
R25040 minus.n23 minus.n22 10.955
R25041 minus.n57 minus.n56 4.80222
R25042 minus.n57 minus.n52 0.972091
R25043 minus.n56 minus.n55 0.716017
R25044 minus.n51 minus.n26 0.189894
R25045 minus.n27 minus.n26 0.189894
R25046 minus.n46 minus.n27 0.189894
R25047 minus.n46 minus.n45 0.189894
R25048 minus.n45 minus.n44 0.189894
R25049 minus.n44 minus.n29 0.189894
R25050 minus.n40 minus.n29 0.189894
R25051 minus.n40 minus.n39 0.189894
R25052 minus.n39 minus.n38 0.189894
R25053 minus.n38 minus.n31 0.189894
R25054 minus.n34 minus.n31 0.189894
R25055 minus.n9 minus.n8 0.189894
R25056 minus.n9 minus.n4 0.189894
R25057 minus.n13 minus.n4 0.189894
R25058 minus.n14 minus.n13 0.189894
R25059 minus.n15 minus.n14 0.189894
R25060 minus.n15 minus.n2 0.189894
R25061 minus.n19 minus.n2 0.189894
R25062 minus.n20 minus.n19 0.189894
R25063 minus.n21 minus.n20 0.189894
R25064 minus.n21 minus.n0 0.189894
R25065 minus.n25 minus.n0 0.189894
R25066 diffpairibias.n0 diffpairibias.t18 436.822
R25067 diffpairibias.n21 diffpairibias.t19 435.479
R25068 diffpairibias.n20 diffpairibias.t16 435.479
R25069 diffpairibias.n19 diffpairibias.t17 435.479
R25070 diffpairibias.n18 diffpairibias.t21 435.479
R25071 diffpairibias.n0 diffpairibias.t22 435.479
R25072 diffpairibias.n1 diffpairibias.t20 435.479
R25073 diffpairibias.n2 diffpairibias.t23 435.479
R25074 diffpairibias.n10 diffpairibias.t0 377.536
R25075 diffpairibias.n10 diffpairibias.t8 376.193
R25076 diffpairibias.n11 diffpairibias.t10 376.193
R25077 diffpairibias.n12 diffpairibias.t6 376.193
R25078 diffpairibias.n13 diffpairibias.t2 376.193
R25079 diffpairibias.n14 diffpairibias.t12 376.193
R25080 diffpairibias.n15 diffpairibias.t4 376.193
R25081 diffpairibias.n16 diffpairibias.t14 376.193
R25082 diffpairibias.n3 diffpairibias.t1 113.368
R25083 diffpairibias.n3 diffpairibias.t9 112.698
R25084 diffpairibias.n4 diffpairibias.t11 112.698
R25085 diffpairibias.n5 diffpairibias.t7 112.698
R25086 diffpairibias.n6 diffpairibias.t3 112.698
R25087 diffpairibias.n7 diffpairibias.t13 112.698
R25088 diffpairibias.n8 diffpairibias.t5 112.698
R25089 diffpairibias.n9 diffpairibias.t15 112.698
R25090 diffpairibias.n17 diffpairibias.n16 4.77242
R25091 diffpairibias.n17 diffpairibias.n9 4.30807
R25092 diffpairibias.n18 diffpairibias.n17 4.13945
R25093 diffpairibias.n16 diffpairibias.n15 1.34352
R25094 diffpairibias.n15 diffpairibias.n14 1.34352
R25095 diffpairibias.n14 diffpairibias.n13 1.34352
R25096 diffpairibias.n13 diffpairibias.n12 1.34352
R25097 diffpairibias.n12 diffpairibias.n11 1.34352
R25098 diffpairibias.n11 diffpairibias.n10 1.34352
R25099 diffpairibias.n2 diffpairibias.n1 1.34352
R25100 diffpairibias.n1 diffpairibias.n0 1.34352
R25101 diffpairibias.n19 diffpairibias.n18 1.34352
R25102 diffpairibias.n20 diffpairibias.n19 1.34352
R25103 diffpairibias.n21 diffpairibias.n20 1.34352
R25104 diffpairibias.n22 diffpairibias.n21 0.862419
R25105 diffpairibias diffpairibias.n22 0.684875
R25106 diffpairibias.n9 diffpairibias.n8 0.672012
R25107 diffpairibias.n8 diffpairibias.n7 0.672012
R25108 diffpairibias.n7 diffpairibias.n6 0.672012
R25109 diffpairibias.n6 diffpairibias.n5 0.672012
R25110 diffpairibias.n5 diffpairibias.n4 0.672012
R25111 diffpairibias.n4 diffpairibias.n3 0.672012
R25112 diffpairibias.n22 diffpairibias.n2 0.190907
R25113 outputibias.n27 outputibias.n1 289.615
R25114 outputibias.n58 outputibias.n32 289.615
R25115 outputibias.n90 outputibias.n64 289.615
R25116 outputibias.n122 outputibias.n96 289.615
R25117 outputibias.n28 outputibias.n27 185
R25118 outputibias.n26 outputibias.n25 185
R25119 outputibias.n5 outputibias.n4 185
R25120 outputibias.n20 outputibias.n19 185
R25121 outputibias.n18 outputibias.n17 185
R25122 outputibias.n9 outputibias.n8 185
R25123 outputibias.n12 outputibias.n11 185
R25124 outputibias.n59 outputibias.n58 185
R25125 outputibias.n57 outputibias.n56 185
R25126 outputibias.n36 outputibias.n35 185
R25127 outputibias.n51 outputibias.n50 185
R25128 outputibias.n49 outputibias.n48 185
R25129 outputibias.n40 outputibias.n39 185
R25130 outputibias.n43 outputibias.n42 185
R25131 outputibias.n91 outputibias.n90 185
R25132 outputibias.n89 outputibias.n88 185
R25133 outputibias.n68 outputibias.n67 185
R25134 outputibias.n83 outputibias.n82 185
R25135 outputibias.n81 outputibias.n80 185
R25136 outputibias.n72 outputibias.n71 185
R25137 outputibias.n75 outputibias.n74 185
R25138 outputibias.n123 outputibias.n122 185
R25139 outputibias.n121 outputibias.n120 185
R25140 outputibias.n100 outputibias.n99 185
R25141 outputibias.n115 outputibias.n114 185
R25142 outputibias.n113 outputibias.n112 185
R25143 outputibias.n104 outputibias.n103 185
R25144 outputibias.n107 outputibias.n106 185
R25145 outputibias.n0 outputibias.t8 178.945
R25146 outputibias.n133 outputibias.t11 177.018
R25147 outputibias.n132 outputibias.t9 177.018
R25148 outputibias.n0 outputibias.t10 177.018
R25149 outputibias.t7 outputibias.n10 147.661
R25150 outputibias.t1 outputibias.n41 147.661
R25151 outputibias.t3 outputibias.n73 147.661
R25152 outputibias.t5 outputibias.n105 147.661
R25153 outputibias.n128 outputibias.t6 132.363
R25154 outputibias.n128 outputibias.t0 130.436
R25155 outputibias.n129 outputibias.t2 130.436
R25156 outputibias.n130 outputibias.t4 130.436
R25157 outputibias.n27 outputibias.n26 104.615
R25158 outputibias.n26 outputibias.n4 104.615
R25159 outputibias.n19 outputibias.n4 104.615
R25160 outputibias.n19 outputibias.n18 104.615
R25161 outputibias.n18 outputibias.n8 104.615
R25162 outputibias.n11 outputibias.n8 104.615
R25163 outputibias.n58 outputibias.n57 104.615
R25164 outputibias.n57 outputibias.n35 104.615
R25165 outputibias.n50 outputibias.n35 104.615
R25166 outputibias.n50 outputibias.n49 104.615
R25167 outputibias.n49 outputibias.n39 104.615
R25168 outputibias.n42 outputibias.n39 104.615
R25169 outputibias.n90 outputibias.n89 104.615
R25170 outputibias.n89 outputibias.n67 104.615
R25171 outputibias.n82 outputibias.n67 104.615
R25172 outputibias.n82 outputibias.n81 104.615
R25173 outputibias.n81 outputibias.n71 104.615
R25174 outputibias.n74 outputibias.n71 104.615
R25175 outputibias.n122 outputibias.n121 104.615
R25176 outputibias.n121 outputibias.n99 104.615
R25177 outputibias.n114 outputibias.n99 104.615
R25178 outputibias.n114 outputibias.n113 104.615
R25179 outputibias.n113 outputibias.n103 104.615
R25180 outputibias.n106 outputibias.n103 104.615
R25181 outputibias.n63 outputibias.n31 95.6354
R25182 outputibias.n63 outputibias.n62 94.6732
R25183 outputibias.n95 outputibias.n94 94.6732
R25184 outputibias.n127 outputibias.n126 94.6732
R25185 outputibias.n11 outputibias.t7 52.3082
R25186 outputibias.n42 outputibias.t1 52.3082
R25187 outputibias.n74 outputibias.t3 52.3082
R25188 outputibias.n106 outputibias.t5 52.3082
R25189 outputibias.n12 outputibias.n10 15.6674
R25190 outputibias.n43 outputibias.n41 15.6674
R25191 outputibias.n75 outputibias.n73 15.6674
R25192 outputibias.n107 outputibias.n105 15.6674
R25193 outputibias.n13 outputibias.n9 12.8005
R25194 outputibias.n44 outputibias.n40 12.8005
R25195 outputibias.n76 outputibias.n72 12.8005
R25196 outputibias.n108 outputibias.n104 12.8005
R25197 outputibias.n17 outputibias.n16 12.0247
R25198 outputibias.n48 outputibias.n47 12.0247
R25199 outputibias.n80 outputibias.n79 12.0247
R25200 outputibias.n112 outputibias.n111 12.0247
R25201 outputibias.n20 outputibias.n7 11.249
R25202 outputibias.n51 outputibias.n38 11.249
R25203 outputibias.n83 outputibias.n70 11.249
R25204 outputibias.n115 outputibias.n102 11.249
R25205 outputibias.n21 outputibias.n5 10.4732
R25206 outputibias.n52 outputibias.n36 10.4732
R25207 outputibias.n84 outputibias.n68 10.4732
R25208 outputibias.n116 outputibias.n100 10.4732
R25209 outputibias.n25 outputibias.n24 9.69747
R25210 outputibias.n56 outputibias.n55 9.69747
R25211 outputibias.n88 outputibias.n87 9.69747
R25212 outputibias.n120 outputibias.n119 9.69747
R25213 outputibias.n31 outputibias.n30 9.45567
R25214 outputibias.n62 outputibias.n61 9.45567
R25215 outputibias.n94 outputibias.n93 9.45567
R25216 outputibias.n126 outputibias.n125 9.45567
R25217 outputibias.n30 outputibias.n29 9.3005
R25218 outputibias.n3 outputibias.n2 9.3005
R25219 outputibias.n24 outputibias.n23 9.3005
R25220 outputibias.n22 outputibias.n21 9.3005
R25221 outputibias.n7 outputibias.n6 9.3005
R25222 outputibias.n16 outputibias.n15 9.3005
R25223 outputibias.n14 outputibias.n13 9.3005
R25224 outputibias.n61 outputibias.n60 9.3005
R25225 outputibias.n34 outputibias.n33 9.3005
R25226 outputibias.n55 outputibias.n54 9.3005
R25227 outputibias.n53 outputibias.n52 9.3005
R25228 outputibias.n38 outputibias.n37 9.3005
R25229 outputibias.n47 outputibias.n46 9.3005
R25230 outputibias.n45 outputibias.n44 9.3005
R25231 outputibias.n93 outputibias.n92 9.3005
R25232 outputibias.n66 outputibias.n65 9.3005
R25233 outputibias.n87 outputibias.n86 9.3005
R25234 outputibias.n85 outputibias.n84 9.3005
R25235 outputibias.n70 outputibias.n69 9.3005
R25236 outputibias.n79 outputibias.n78 9.3005
R25237 outputibias.n77 outputibias.n76 9.3005
R25238 outputibias.n125 outputibias.n124 9.3005
R25239 outputibias.n98 outputibias.n97 9.3005
R25240 outputibias.n119 outputibias.n118 9.3005
R25241 outputibias.n117 outputibias.n116 9.3005
R25242 outputibias.n102 outputibias.n101 9.3005
R25243 outputibias.n111 outputibias.n110 9.3005
R25244 outputibias.n109 outputibias.n108 9.3005
R25245 outputibias.n28 outputibias.n3 8.92171
R25246 outputibias.n59 outputibias.n34 8.92171
R25247 outputibias.n91 outputibias.n66 8.92171
R25248 outputibias.n123 outputibias.n98 8.92171
R25249 outputibias.n29 outputibias.n1 8.14595
R25250 outputibias.n60 outputibias.n32 8.14595
R25251 outputibias.n92 outputibias.n64 8.14595
R25252 outputibias.n124 outputibias.n96 8.14595
R25253 outputibias.n31 outputibias.n1 5.81868
R25254 outputibias.n62 outputibias.n32 5.81868
R25255 outputibias.n94 outputibias.n64 5.81868
R25256 outputibias.n126 outputibias.n96 5.81868
R25257 outputibias.n131 outputibias.n130 5.20947
R25258 outputibias.n29 outputibias.n28 5.04292
R25259 outputibias.n60 outputibias.n59 5.04292
R25260 outputibias.n92 outputibias.n91 5.04292
R25261 outputibias.n124 outputibias.n123 5.04292
R25262 outputibias.n131 outputibias.n127 4.42209
R25263 outputibias.n14 outputibias.n10 4.38594
R25264 outputibias.n45 outputibias.n41 4.38594
R25265 outputibias.n77 outputibias.n73 4.38594
R25266 outputibias.n109 outputibias.n105 4.38594
R25267 outputibias.n132 outputibias.n131 4.28454
R25268 outputibias.n25 outputibias.n3 4.26717
R25269 outputibias.n56 outputibias.n34 4.26717
R25270 outputibias.n88 outputibias.n66 4.26717
R25271 outputibias.n120 outputibias.n98 4.26717
R25272 outputibias.n24 outputibias.n5 3.49141
R25273 outputibias.n55 outputibias.n36 3.49141
R25274 outputibias.n87 outputibias.n68 3.49141
R25275 outputibias.n119 outputibias.n100 3.49141
R25276 outputibias.n21 outputibias.n20 2.71565
R25277 outputibias.n52 outputibias.n51 2.71565
R25278 outputibias.n84 outputibias.n83 2.71565
R25279 outputibias.n116 outputibias.n115 2.71565
R25280 outputibias.n17 outputibias.n7 1.93989
R25281 outputibias.n48 outputibias.n38 1.93989
R25282 outputibias.n80 outputibias.n70 1.93989
R25283 outputibias.n112 outputibias.n102 1.93989
R25284 outputibias.n130 outputibias.n129 1.9266
R25285 outputibias.n129 outputibias.n128 1.9266
R25286 outputibias.n133 outputibias.n132 1.92658
R25287 outputibias.n134 outputibias.n133 1.29913
R25288 outputibias.n16 outputibias.n9 1.16414
R25289 outputibias.n47 outputibias.n40 1.16414
R25290 outputibias.n79 outputibias.n72 1.16414
R25291 outputibias.n111 outputibias.n104 1.16414
R25292 outputibias.n127 outputibias.n95 0.962709
R25293 outputibias.n95 outputibias.n63 0.962709
R25294 outputibias.n13 outputibias.n12 0.388379
R25295 outputibias.n44 outputibias.n43 0.388379
R25296 outputibias.n76 outputibias.n75 0.388379
R25297 outputibias.n108 outputibias.n107 0.388379
R25298 outputibias.n134 outputibias.n0 0.337251
R25299 outputibias outputibias.n134 0.302375
R25300 outputibias.n30 outputibias.n2 0.155672
R25301 outputibias.n23 outputibias.n2 0.155672
R25302 outputibias.n23 outputibias.n22 0.155672
R25303 outputibias.n22 outputibias.n6 0.155672
R25304 outputibias.n15 outputibias.n6 0.155672
R25305 outputibias.n15 outputibias.n14 0.155672
R25306 outputibias.n61 outputibias.n33 0.155672
R25307 outputibias.n54 outputibias.n33 0.155672
R25308 outputibias.n54 outputibias.n53 0.155672
R25309 outputibias.n53 outputibias.n37 0.155672
R25310 outputibias.n46 outputibias.n37 0.155672
R25311 outputibias.n46 outputibias.n45 0.155672
R25312 outputibias.n93 outputibias.n65 0.155672
R25313 outputibias.n86 outputibias.n65 0.155672
R25314 outputibias.n86 outputibias.n85 0.155672
R25315 outputibias.n85 outputibias.n69 0.155672
R25316 outputibias.n78 outputibias.n69 0.155672
R25317 outputibias.n78 outputibias.n77 0.155672
R25318 outputibias.n125 outputibias.n97 0.155672
R25319 outputibias.n118 outputibias.n97 0.155672
R25320 outputibias.n118 outputibias.n117 0.155672
R25321 outputibias.n117 outputibias.n101 0.155672
R25322 outputibias.n110 outputibias.n101 0.155672
R25323 outputibias.n110 outputibias.n109 0.155672
C0 plus commonsourceibias 0.273048f
C1 output outputibias 2.34152f
C2 vdd output 7.23429f
C3 CSoutput output 6.13881f
C4 CSoutput outputibias 0.032386f
C5 vdd CSoutput 0.117233p
C6 minus diffpairibias 3.1e-19
C7 commonsourceibias output 0.006808f
C8 CSoutput minus 3.13952f
C9 vdd plus 0.090904f
C10 commonsourceibias outputibias 0.003832f
C11 plus diffpairibias 3.12e-19
C12 vdd commonsourceibias 0.004218f
C13 CSoutput plus 0.862911f
C14 commonsourceibias diffpairibias 0.06482f
C15 CSoutput commonsourceibias 66.33679f
C16 minus plus 9.237121f
C17 minus commonsourceibias 0.318966f
C18 diffpairibias gnd 48.980038f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.222615p
C22 plus gnd 31.7302f
C23 minus gnd 27.363628f
C24 CSoutput gnd 0.143035p
C25 vdd gnd 0.511372p
C26 outputibias.t10 gnd 0.11477f
C27 outputibias.t8 gnd 0.115567f
C28 outputibias.n0 gnd 0.130108f
C29 outputibias.n1 gnd 0.001372f
C30 outputibias.n2 gnd 9.76e-19
C31 outputibias.n3 gnd 5.24e-19
C32 outputibias.n4 gnd 0.001239f
C33 outputibias.n5 gnd 5.55e-19
C34 outputibias.n6 gnd 9.76e-19
C35 outputibias.n7 gnd 5.24e-19
C36 outputibias.n8 gnd 0.001239f
C37 outputibias.n9 gnd 5.55e-19
C38 outputibias.n10 gnd 0.004176f
C39 outputibias.t7 gnd 0.00202f
C40 outputibias.n11 gnd 9.3e-19
C41 outputibias.n12 gnd 7.32e-19
C42 outputibias.n13 gnd 5.24e-19
C43 outputibias.n14 gnd 0.02322f
C44 outputibias.n15 gnd 9.76e-19
C45 outputibias.n16 gnd 5.24e-19
C46 outputibias.n17 gnd 5.55e-19
C47 outputibias.n18 gnd 0.001239f
C48 outputibias.n19 gnd 0.001239f
C49 outputibias.n20 gnd 5.55e-19
C50 outputibias.n21 gnd 5.24e-19
C51 outputibias.n22 gnd 9.76e-19
C52 outputibias.n23 gnd 9.76e-19
C53 outputibias.n24 gnd 5.24e-19
C54 outputibias.n25 gnd 5.55e-19
C55 outputibias.n26 gnd 0.001239f
C56 outputibias.n27 gnd 0.002683f
C57 outputibias.n28 gnd 5.55e-19
C58 outputibias.n29 gnd 5.24e-19
C59 outputibias.n30 gnd 0.002256f
C60 outputibias.n31 gnd 0.005781f
C61 outputibias.n32 gnd 0.001372f
C62 outputibias.n33 gnd 9.76e-19
C63 outputibias.n34 gnd 5.24e-19
C64 outputibias.n35 gnd 0.001239f
C65 outputibias.n36 gnd 5.55e-19
C66 outputibias.n37 gnd 9.76e-19
C67 outputibias.n38 gnd 5.24e-19
C68 outputibias.n39 gnd 0.001239f
C69 outputibias.n40 gnd 5.55e-19
C70 outputibias.n41 gnd 0.004176f
C71 outputibias.t1 gnd 0.00202f
C72 outputibias.n42 gnd 9.3e-19
C73 outputibias.n43 gnd 7.32e-19
C74 outputibias.n44 gnd 5.24e-19
C75 outputibias.n45 gnd 0.02322f
C76 outputibias.n46 gnd 9.76e-19
C77 outputibias.n47 gnd 5.24e-19
C78 outputibias.n48 gnd 5.55e-19
C79 outputibias.n49 gnd 0.001239f
C80 outputibias.n50 gnd 0.001239f
C81 outputibias.n51 gnd 5.55e-19
C82 outputibias.n52 gnd 5.24e-19
C83 outputibias.n53 gnd 9.76e-19
C84 outputibias.n54 gnd 9.76e-19
C85 outputibias.n55 gnd 5.24e-19
C86 outputibias.n56 gnd 5.55e-19
C87 outputibias.n57 gnd 0.001239f
C88 outputibias.n58 gnd 0.002683f
C89 outputibias.n59 gnd 5.55e-19
C90 outputibias.n60 gnd 5.24e-19
C91 outputibias.n61 gnd 0.002256f
C92 outputibias.n62 gnd 0.005197f
C93 outputibias.n63 gnd 0.121892f
C94 outputibias.n64 gnd 0.001372f
C95 outputibias.n65 gnd 9.76e-19
C96 outputibias.n66 gnd 5.24e-19
C97 outputibias.n67 gnd 0.001239f
C98 outputibias.n68 gnd 5.55e-19
C99 outputibias.n69 gnd 9.76e-19
C100 outputibias.n70 gnd 5.24e-19
C101 outputibias.n71 gnd 0.001239f
C102 outputibias.n72 gnd 5.55e-19
C103 outputibias.n73 gnd 0.004176f
C104 outputibias.t3 gnd 0.00202f
C105 outputibias.n74 gnd 9.3e-19
C106 outputibias.n75 gnd 7.32e-19
C107 outputibias.n76 gnd 5.24e-19
C108 outputibias.n77 gnd 0.02322f
C109 outputibias.n78 gnd 9.76e-19
C110 outputibias.n79 gnd 5.24e-19
C111 outputibias.n80 gnd 5.55e-19
C112 outputibias.n81 gnd 0.001239f
C113 outputibias.n82 gnd 0.001239f
C114 outputibias.n83 gnd 5.55e-19
C115 outputibias.n84 gnd 5.24e-19
C116 outputibias.n85 gnd 9.76e-19
C117 outputibias.n86 gnd 9.76e-19
C118 outputibias.n87 gnd 5.24e-19
C119 outputibias.n88 gnd 5.55e-19
C120 outputibias.n89 gnd 0.001239f
C121 outputibias.n90 gnd 0.002683f
C122 outputibias.n91 gnd 5.55e-19
C123 outputibias.n92 gnd 5.24e-19
C124 outputibias.n93 gnd 0.002256f
C125 outputibias.n94 gnd 0.005197f
C126 outputibias.n95 gnd 0.064513f
C127 outputibias.n96 gnd 0.001372f
C128 outputibias.n97 gnd 9.76e-19
C129 outputibias.n98 gnd 5.24e-19
C130 outputibias.n99 gnd 0.001239f
C131 outputibias.n100 gnd 5.55e-19
C132 outputibias.n101 gnd 9.76e-19
C133 outputibias.n102 gnd 5.24e-19
C134 outputibias.n103 gnd 0.001239f
C135 outputibias.n104 gnd 5.55e-19
C136 outputibias.n105 gnd 0.004176f
C137 outputibias.t5 gnd 0.00202f
C138 outputibias.n106 gnd 9.3e-19
C139 outputibias.n107 gnd 7.32e-19
C140 outputibias.n108 gnd 5.24e-19
C141 outputibias.n109 gnd 0.02322f
C142 outputibias.n110 gnd 9.76e-19
C143 outputibias.n111 gnd 5.24e-19
C144 outputibias.n112 gnd 5.55e-19
C145 outputibias.n113 gnd 0.001239f
C146 outputibias.n114 gnd 0.001239f
C147 outputibias.n115 gnd 5.55e-19
C148 outputibias.n116 gnd 5.24e-19
C149 outputibias.n117 gnd 9.76e-19
C150 outputibias.n118 gnd 9.76e-19
C151 outputibias.n119 gnd 5.24e-19
C152 outputibias.n120 gnd 5.55e-19
C153 outputibias.n121 gnd 0.001239f
C154 outputibias.n122 gnd 0.002683f
C155 outputibias.n123 gnd 5.55e-19
C156 outputibias.n124 gnd 5.24e-19
C157 outputibias.n125 gnd 0.002256f
C158 outputibias.n126 gnd 0.005197f
C159 outputibias.n127 gnd 0.084814f
C160 outputibias.t4 gnd 0.108319f
C161 outputibias.t2 gnd 0.108319f
C162 outputibias.t0 gnd 0.108319f
C163 outputibias.t6 gnd 0.109238f
C164 outputibias.n128 gnd 0.134674f
C165 outputibias.n129 gnd 0.07244f
C166 outputibias.n130 gnd 0.079818f
C167 outputibias.n131 gnd 0.164901f
C168 outputibias.t9 gnd 0.11477f
C169 outputibias.n132 gnd 0.067481f
C170 outputibias.t11 gnd 0.11477f
C171 outputibias.n133 gnd 0.065115f
C172 outputibias.n134 gnd 0.029159f
C173 diffpairibias.t18 gnd 0.087401f
C174 diffpairibias.t22 gnd 0.087239f
C175 diffpairibias.n0 gnd 0.102784f
C176 diffpairibias.t20 gnd 0.087239f
C177 diffpairibias.n1 gnd 0.050171f
C178 diffpairibias.t23 gnd 0.087239f
C179 diffpairibias.n2 gnd 0.039841f
C180 diffpairibias.t1 gnd 0.083757f
C181 diffpairibias.t9 gnd 0.083392f
C182 diffpairibias.n3 gnd 0.131682f
C183 diffpairibias.t11 gnd 0.083392f
C184 diffpairibias.n4 gnd 0.07027f
C185 diffpairibias.t7 gnd 0.083392f
C186 diffpairibias.n5 gnd 0.07027f
C187 diffpairibias.t3 gnd 0.083392f
C188 diffpairibias.n6 gnd 0.07027f
C189 diffpairibias.t13 gnd 0.083392f
C190 diffpairibias.n7 gnd 0.07027f
C191 diffpairibias.t5 gnd 0.083392f
C192 diffpairibias.n8 gnd 0.07027f
C193 diffpairibias.t15 gnd 0.083392f
C194 diffpairibias.n9 gnd 0.099771f
C195 diffpairibias.t0 gnd 0.08427f
C196 diffpairibias.t8 gnd 0.084123f
C197 diffpairibias.n10 gnd 0.091784f
C198 diffpairibias.t10 gnd 0.084123f
C199 diffpairibias.n11 gnd 0.050681f
C200 diffpairibias.t6 gnd 0.084123f
C201 diffpairibias.n12 gnd 0.050681f
C202 diffpairibias.t2 gnd 0.084123f
C203 diffpairibias.n13 gnd 0.050681f
C204 diffpairibias.t12 gnd 0.084123f
C205 diffpairibias.n14 gnd 0.050681f
C206 diffpairibias.t4 gnd 0.084123f
C207 diffpairibias.n15 gnd 0.050681f
C208 diffpairibias.t14 gnd 0.084123f
C209 diffpairibias.n16 gnd 0.059977f
C210 diffpairibias.n17 gnd 0.226448f
C211 diffpairibias.t21 gnd 0.087239f
C212 diffpairibias.n18 gnd 0.050181f
C213 diffpairibias.t17 gnd 0.087239f
C214 diffpairibias.n19 gnd 0.050171f
C215 diffpairibias.t16 gnd 0.087239f
C216 diffpairibias.n20 gnd 0.050171f
C217 diffpairibias.t19 gnd 0.087239f
C218 diffpairibias.n21 gnd 0.045859f
C219 diffpairibias.n22 gnd 0.046268f
C220 minus.n0 gnd 0.030081f
C221 minus.n1 gnd 0.006826f
C222 minus.n2 gnd 0.030081f
C223 minus.n3 gnd 0.006826f
C224 minus.n4 gnd 0.030081f
C225 minus.n5 gnd 0.006826f
C226 minus.t6 gnd 0.439814f
C227 minus.t5 gnd 0.425475f
C228 minus.n6 gnd 0.19313f
C229 minus.n7 gnd 0.177173f
C230 minus.n8 gnd 0.127298f
C231 minus.n9 gnd 0.030081f
C232 minus.t9 gnd 0.425475f
C233 minus.n10 gnd 0.189009f
C234 minus.n11 gnd 0.006826f
C235 minus.t8 gnd 0.425475f
C236 minus.n12 gnd 0.189009f
C237 minus.n13 gnd 0.030081f
C238 minus.n14 gnd 0.030081f
C239 minus.n15 gnd 0.030081f
C240 minus.t10 gnd 0.425475f
C241 minus.n16 gnd 0.189009f
C242 minus.n17 gnd 0.006826f
C243 minus.t14 gnd 0.425475f
C244 minus.n18 gnd 0.189009f
C245 minus.n19 gnd 0.030081f
C246 minus.n20 gnd 0.030081f
C247 minus.n21 gnd 0.030081f
C248 minus.t13 gnd 0.425475f
C249 minus.n22 gnd 0.189009f
C250 minus.n23 gnd 0.006826f
C251 minus.t17 gnd 0.425475f
C252 minus.n24 gnd 0.188175f
C253 minus.n25 gnd 0.346762f
C254 minus.n26 gnd 0.030081f
C255 minus.t18 gnd 0.425475f
C256 minus.t15 gnd 0.425475f
C257 minus.n27 gnd 0.030081f
C258 minus.t16 gnd 0.425475f
C259 minus.n28 gnd 0.189009f
C260 minus.n29 gnd 0.030081f
C261 minus.t11 gnd 0.425475f
C262 minus.t12 gnd 0.425475f
C263 minus.n30 gnd 0.189009f
C264 minus.n31 gnd 0.030081f
C265 minus.t7 gnd 0.425475f
C266 minus.t19 gnd 0.425475f
C267 minus.n32 gnd 0.19313f
C268 minus.t20 gnd 0.439814f
C269 minus.n33 gnd 0.177173f
C270 minus.n34 gnd 0.127298f
C271 minus.n35 gnd 0.006826f
C272 minus.n36 gnd 0.189009f
C273 minus.n37 gnd 0.006826f
C274 minus.n38 gnd 0.030081f
C275 minus.n39 gnd 0.030081f
C276 minus.n40 gnd 0.030081f
C277 minus.n41 gnd 0.006826f
C278 minus.n42 gnd 0.189009f
C279 minus.n43 gnd 0.006826f
C280 minus.n44 gnd 0.030081f
C281 minus.n45 gnd 0.030081f
C282 minus.n46 gnd 0.030081f
C283 minus.n47 gnd 0.006826f
C284 minus.n48 gnd 0.189009f
C285 minus.n49 gnd 0.006826f
C286 minus.n50 gnd 0.188175f
C287 minus.n51 gnd 0.873119f
C288 minus.n52 gnd 1.3277f
C289 minus.t1 gnd 0.009273f
C290 minus.t0 gnd 0.009273f
C291 minus.n53 gnd 0.030493f
C292 minus.t3 gnd 0.009273f
C293 minus.t2 gnd 0.009273f
C294 minus.n54 gnd 0.030075f
C295 minus.n55 gnd 0.256674f
C296 minus.t4 gnd 0.051614f
C297 minus.n56 gnd 0.140065f
C298 minus.n57 gnd 2.20692f
C299 output.t3 gnd 0.464308f
C300 output.t13 gnd 0.044422f
C301 output.t11 gnd 0.044422f
C302 output.n0 gnd 0.364624f
C303 output.n1 gnd 0.614102f
C304 output.t18 gnd 0.044422f
C305 output.t5 gnd 0.044422f
C306 output.n2 gnd 0.364624f
C307 output.n3 gnd 0.350265f
C308 output.t7 gnd 0.044422f
C309 output.t15 gnd 0.044422f
C310 output.n4 gnd 0.364624f
C311 output.n5 gnd 0.350265f
C312 output.t17 gnd 0.044422f
C313 output.t8 gnd 0.044422f
C314 output.n6 gnd 0.364624f
C315 output.n7 gnd 0.350265f
C316 output.t9 gnd 0.044422f
C317 output.t14 gnd 0.044422f
C318 output.n8 gnd 0.364624f
C319 output.n9 gnd 0.350265f
C320 output.t16 gnd 0.044422f
C321 output.t6 gnd 0.044422f
C322 output.n10 gnd 0.364624f
C323 output.n11 gnd 0.350265f
C324 output.t12 gnd 0.044422f
C325 output.t10 gnd 0.044422f
C326 output.n12 gnd 0.364624f
C327 output.n13 gnd 0.350265f
C328 output.t4 gnd 0.462979f
C329 output.n14 gnd 0.28994f
C330 output.n15 gnd 0.015803f
C331 output.n16 gnd 0.011243f
C332 output.n17 gnd 0.006041f
C333 output.n18 gnd 0.01428f
C334 output.n19 gnd 0.006397f
C335 output.n20 gnd 0.011243f
C336 output.n21 gnd 0.006041f
C337 output.n22 gnd 0.01428f
C338 output.n23 gnd 0.006397f
C339 output.n24 gnd 0.048111f
C340 output.t1 gnd 0.023274f
C341 output.n25 gnd 0.01071f
C342 output.n26 gnd 0.008435f
C343 output.n27 gnd 0.006041f
C344 output.n28 gnd 0.267512f
C345 output.n29 gnd 0.011243f
C346 output.n30 gnd 0.006041f
C347 output.n31 gnd 0.006397f
C348 output.n32 gnd 0.01428f
C349 output.n33 gnd 0.01428f
C350 output.n34 gnd 0.006397f
C351 output.n35 gnd 0.006041f
C352 output.n36 gnd 0.011243f
C353 output.n37 gnd 0.011243f
C354 output.n38 gnd 0.006041f
C355 output.n39 gnd 0.006397f
C356 output.n40 gnd 0.01428f
C357 output.n41 gnd 0.030913f
C358 output.n42 gnd 0.006397f
C359 output.n43 gnd 0.006041f
C360 output.n44 gnd 0.025987f
C361 output.n45 gnd 0.097665f
C362 output.n46 gnd 0.015803f
C363 output.n47 gnd 0.011243f
C364 output.n48 gnd 0.006041f
C365 output.n49 gnd 0.01428f
C366 output.n50 gnd 0.006397f
C367 output.n51 gnd 0.011243f
C368 output.n52 gnd 0.006041f
C369 output.n53 gnd 0.01428f
C370 output.n54 gnd 0.006397f
C371 output.n55 gnd 0.048111f
C372 output.t19 gnd 0.023274f
C373 output.n56 gnd 0.01071f
C374 output.n57 gnd 0.008435f
C375 output.n58 gnd 0.006041f
C376 output.n59 gnd 0.267512f
C377 output.n60 gnd 0.011243f
C378 output.n61 gnd 0.006041f
C379 output.n62 gnd 0.006397f
C380 output.n63 gnd 0.01428f
C381 output.n64 gnd 0.01428f
C382 output.n65 gnd 0.006397f
C383 output.n66 gnd 0.006041f
C384 output.n67 gnd 0.011243f
C385 output.n68 gnd 0.011243f
C386 output.n69 gnd 0.006041f
C387 output.n70 gnd 0.006397f
C388 output.n71 gnd 0.01428f
C389 output.n72 gnd 0.030913f
C390 output.n73 gnd 0.006397f
C391 output.n74 gnd 0.006041f
C392 output.n75 gnd 0.025987f
C393 output.n76 gnd 0.09306f
C394 output.n77 gnd 1.65264f
C395 output.n78 gnd 0.015803f
C396 output.n79 gnd 0.011243f
C397 output.n80 gnd 0.006041f
C398 output.n81 gnd 0.01428f
C399 output.n82 gnd 0.006397f
C400 output.n83 gnd 0.011243f
C401 output.n84 gnd 0.006041f
C402 output.n85 gnd 0.01428f
C403 output.n86 gnd 0.006397f
C404 output.n87 gnd 0.048111f
C405 output.t0 gnd 0.023274f
C406 output.n88 gnd 0.01071f
C407 output.n89 gnd 0.008435f
C408 output.n90 gnd 0.006041f
C409 output.n91 gnd 0.267512f
C410 output.n92 gnd 0.011243f
C411 output.n93 gnd 0.006041f
C412 output.n94 gnd 0.006397f
C413 output.n95 gnd 0.01428f
C414 output.n96 gnd 0.01428f
C415 output.n97 gnd 0.006397f
C416 output.n98 gnd 0.006041f
C417 output.n99 gnd 0.011243f
C418 output.n100 gnd 0.011243f
C419 output.n101 gnd 0.006041f
C420 output.n102 gnd 0.006397f
C421 output.n103 gnd 0.01428f
C422 output.n104 gnd 0.030913f
C423 output.n105 gnd 0.006397f
C424 output.n106 gnd 0.006041f
C425 output.n107 gnd 0.025987f
C426 output.n108 gnd 0.09306f
C427 output.n109 gnd 0.713089f
C428 output.n110 gnd 0.015803f
C429 output.n111 gnd 0.011243f
C430 output.n112 gnd 0.006041f
C431 output.n113 gnd 0.01428f
C432 output.n114 gnd 0.006397f
C433 output.n115 gnd 0.011243f
C434 output.n116 gnd 0.006041f
C435 output.n117 gnd 0.01428f
C436 output.n118 gnd 0.006397f
C437 output.n119 gnd 0.048111f
C438 output.t2 gnd 0.023274f
C439 output.n120 gnd 0.01071f
C440 output.n121 gnd 0.008435f
C441 output.n122 gnd 0.006041f
C442 output.n123 gnd 0.267512f
C443 output.n124 gnd 0.011243f
C444 output.n125 gnd 0.006041f
C445 output.n126 gnd 0.006397f
C446 output.n127 gnd 0.01428f
C447 output.n128 gnd 0.01428f
C448 output.n129 gnd 0.006397f
C449 output.n130 gnd 0.006041f
C450 output.n131 gnd 0.011243f
C451 output.n132 gnd 0.011243f
C452 output.n133 gnd 0.006041f
C453 output.n134 gnd 0.006397f
C454 output.n135 gnd 0.01428f
C455 output.n136 gnd 0.030913f
C456 output.n137 gnd 0.006397f
C457 output.n138 gnd 0.006041f
C458 output.n139 gnd 0.025987f
C459 output.n140 gnd 0.09306f
C460 output.n141 gnd 1.67353f
C461 a_n2982_8322.t7 gnd 0.100149f
C462 a_n2982_8322.t33 gnd 20.7769f
C463 a_n2982_8322.t34 gnd 20.631199f
C464 a_n2982_8322.t36 gnd 20.631199f
C465 a_n2982_8322.t32 gnd 20.7769f
C466 a_n2982_8322.t35 gnd 20.631199f
C467 a_n2982_8322.t37 gnd 29.5576f
C468 a_n2982_8322.t6 gnd 0.937748f
C469 a_n2982_8322.t19 gnd 0.100149f
C470 a_n2982_8322.t15 gnd 0.100149f
C471 a_n2982_8322.n0 gnd 0.705452f
C472 a_n2982_8322.n1 gnd 0.788239f
C473 a_n2982_8322.t22 gnd 0.100149f
C474 a_n2982_8322.t12 gnd 0.100149f
C475 a_n2982_8322.n2 gnd 0.705452f
C476 a_n2982_8322.n3 gnd 0.400494f
C477 a_n2982_8322.t3 gnd 0.100149f
C478 a_n2982_8322.t2 gnd 0.100149f
C479 a_n2982_8322.n4 gnd 0.705452f
C480 a_n2982_8322.n5 gnd 0.400494f
C481 a_n2982_8322.t16 gnd 0.100149f
C482 a_n2982_8322.t9 gnd 0.100149f
C483 a_n2982_8322.n6 gnd 0.705452f
C484 a_n2982_8322.n7 gnd 0.400494f
C485 a_n2982_8322.t13 gnd 0.100149f
C486 a_n2982_8322.t11 gnd 0.100149f
C487 a_n2982_8322.n8 gnd 0.705452f
C488 a_n2982_8322.n9 gnd 0.400494f
C489 a_n2982_8322.t0 gnd 0.935881f
C490 a_n2982_8322.n10 gnd 1.8712f
C491 a_n2982_8322.t27 gnd 0.937748f
C492 a_n2982_8322.t31 gnd 0.100149f
C493 a_n2982_8322.t30 gnd 0.100149f
C494 a_n2982_8322.n11 gnd 0.705452f
C495 a_n2982_8322.n12 gnd 0.788239f
C496 a_n2982_8322.t25 gnd 0.935881f
C497 a_n2982_8322.n13 gnd 0.396653f
C498 a_n2982_8322.t28 gnd 0.935881f
C499 a_n2982_8322.n14 gnd 0.396653f
C500 a_n2982_8322.t26 gnd 0.100149f
C501 a_n2982_8322.t24 gnd 0.100149f
C502 a_n2982_8322.n15 gnd 0.705452f
C503 a_n2982_8322.n16 gnd 0.400494f
C504 a_n2982_8322.t29 gnd 0.935881f
C505 a_n2982_8322.n17 gnd 1.47125f
C506 a_n2982_8322.n18 gnd 2.3511f
C507 a_n2982_8322.n19 gnd 3.56583f
C508 a_n2982_8322.t1 gnd 0.935881f
C509 a_n2982_8322.n20 gnd 1.11135f
C510 a_n2982_8322.t18 gnd 0.100149f
C511 a_n2982_8322.t17 gnd 0.100149f
C512 a_n2982_8322.n21 gnd 0.705452f
C513 a_n2982_8322.n22 gnd 0.400494f
C514 a_n2982_8322.t5 gnd 0.100149f
C515 a_n2982_8322.t4 gnd 0.100149f
C516 a_n2982_8322.n23 gnd 0.705452f
C517 a_n2982_8322.n24 gnd 0.400494f
C518 a_n2982_8322.t20 gnd 0.100149f
C519 a_n2982_8322.t8 gnd 0.100149f
C520 a_n2982_8322.n25 gnd 0.705452f
C521 a_n2982_8322.n26 gnd 0.400494f
C522 a_n2982_8322.t21 gnd 0.937745f
C523 a_n2982_8322.t14 gnd 0.100149f
C524 a_n2982_8322.t10 gnd 0.100149f
C525 a_n2982_8322.n27 gnd 0.705452f
C526 a_n2982_8322.n28 gnd 0.788241f
C527 a_n2982_8322.n29 gnd 0.400492f
C528 a_n2982_8322.n30 gnd 0.705454f
C529 a_n2982_8322.t23 gnd 0.100149f
C530 CSoutput.n0 gnd 0.045881f
C531 CSoutput.t226 gnd 0.303495f
C532 CSoutput.n1 gnd 0.137043f
C533 CSoutput.n2 gnd 0.045881f
C534 CSoutput.t224 gnd 0.303495f
C535 CSoutput.n3 gnd 0.036365f
C536 CSoutput.n4 gnd 0.045881f
C537 CSoutput.t217 gnd 0.303495f
C538 CSoutput.n5 gnd 0.031358f
C539 CSoutput.n6 gnd 0.045881f
C540 CSoutput.t221 gnd 0.303495f
C541 CSoutput.t231 gnd 0.303495f
C542 CSoutput.n7 gnd 0.135549f
C543 CSoutput.n8 gnd 0.045881f
C544 CSoutput.t229 gnd 0.303495f
C545 CSoutput.n9 gnd 0.029898f
C546 CSoutput.n10 gnd 0.045881f
C547 CSoutput.t218 gnd 0.303495f
C548 CSoutput.t223 gnd 0.303495f
C549 CSoutput.n11 gnd 0.135549f
C550 CSoutput.n12 gnd 0.045881f
C551 CSoutput.t228 gnd 0.303495f
C552 CSoutput.n13 gnd 0.031358f
C553 CSoutput.n14 gnd 0.045881f
C554 CSoutput.t233 gnd 0.303495f
C555 CSoutput.t220 gnd 0.303495f
C556 CSoutput.n15 gnd 0.135549f
C557 CSoutput.n16 gnd 0.045881f
C558 CSoutput.t227 gnd 0.303495f
C559 CSoutput.n17 gnd 0.033491f
C560 CSoutput.t235 gnd 0.362684f
C561 CSoutput.t225 gnd 0.303495f
C562 CSoutput.n18 gnd 0.173044f
C563 CSoutput.n19 gnd 0.167912f
C564 CSoutput.n20 gnd 0.194798f
C565 CSoutput.n21 gnd 0.045881f
C566 CSoutput.n22 gnd 0.038293f
C567 CSoutput.n23 gnd 0.135549f
C568 CSoutput.n24 gnd 0.036913f
C569 CSoutput.n25 gnd 0.036365f
C570 CSoutput.n26 gnd 0.045881f
C571 CSoutput.n27 gnd 0.045881f
C572 CSoutput.n28 gnd 0.037999f
C573 CSoutput.n29 gnd 0.032262f
C574 CSoutput.n30 gnd 0.138567f
C575 CSoutput.n31 gnd 0.032706f
C576 CSoutput.n32 gnd 0.045881f
C577 CSoutput.n33 gnd 0.045881f
C578 CSoutput.n34 gnd 0.045881f
C579 CSoutput.n35 gnd 0.037594f
C580 CSoutput.n36 gnd 0.135549f
C581 CSoutput.n37 gnd 0.035953f
C582 CSoutput.n38 gnd 0.037325f
C583 CSoutput.n39 gnd 0.045881f
C584 CSoutput.n40 gnd 0.045881f
C585 CSoutput.n41 gnd 0.038285f
C586 CSoutput.n42 gnd 0.034993f
C587 CSoutput.n43 gnd 0.135549f
C588 CSoutput.n44 gnd 0.03588f
C589 CSoutput.n45 gnd 0.045881f
C590 CSoutput.n46 gnd 0.045881f
C591 CSoutput.n47 gnd 0.045881f
C592 CSoutput.n48 gnd 0.03588f
C593 CSoutput.n49 gnd 0.135549f
C594 CSoutput.n50 gnd 0.034993f
C595 CSoutput.n51 gnd 0.038285f
C596 CSoutput.n52 gnd 0.045881f
C597 CSoutput.n53 gnd 0.045881f
C598 CSoutput.n54 gnd 0.037325f
C599 CSoutput.n55 gnd 0.035953f
C600 CSoutput.n56 gnd 0.135549f
C601 CSoutput.n57 gnd 0.037594f
C602 CSoutput.n58 gnd 0.045881f
C603 CSoutput.n59 gnd 0.045881f
C604 CSoutput.n60 gnd 0.045881f
C605 CSoutput.n61 gnd 0.032706f
C606 CSoutput.n62 gnd 0.138567f
C607 CSoutput.n63 gnd 0.032262f
C608 CSoutput.t234 gnd 0.303495f
C609 CSoutput.n64 gnd 0.135549f
C610 CSoutput.n65 gnd 0.037999f
C611 CSoutput.n66 gnd 0.045881f
C612 CSoutput.n67 gnd 0.045881f
C613 CSoutput.n68 gnd 0.045881f
C614 CSoutput.n69 gnd 0.036913f
C615 CSoutput.n70 gnd 0.135549f
C616 CSoutput.n71 gnd 0.038293f
C617 CSoutput.n72 gnd 0.033491f
C618 CSoutput.n73 gnd 0.045881f
C619 CSoutput.n74 gnd 0.045881f
C620 CSoutput.n75 gnd 0.034733f
C621 CSoutput.n76 gnd 0.020628f
C622 CSoutput.t236 gnd 0.340998f
C623 CSoutput.n77 gnd 0.169394f
C624 CSoutput.n78 gnd 0.692982f
C625 CSoutput.t95 gnd 0.05723f
C626 CSoutput.t43 gnd 0.05723f
C627 CSoutput.n79 gnd 0.443097f
C628 CSoutput.t11 gnd 0.05723f
C629 CSoutput.t77 gnd 0.05723f
C630 CSoutput.n80 gnd 0.442307f
C631 CSoutput.n81 gnd 0.448941f
C632 CSoutput.t18 gnd 0.05723f
C633 CSoutput.t62 gnd 0.05723f
C634 CSoutput.n82 gnd 0.442307f
C635 CSoutput.n83 gnd 0.221219f
C636 CSoutput.t34 gnd 0.05723f
C637 CSoutput.t50 gnd 0.05723f
C638 CSoutput.n84 gnd 0.442307f
C639 CSoutput.n85 gnd 0.221219f
C640 CSoutput.t46 gnd 0.05723f
C641 CSoutput.t85 gnd 0.05723f
C642 CSoutput.n86 gnd 0.442307f
C643 CSoutput.n87 gnd 0.221219f
C644 CSoutput.t25 gnd 0.05723f
C645 CSoutput.t67 gnd 0.05723f
C646 CSoutput.n88 gnd 0.442307f
C647 CSoutput.n89 gnd 0.221219f
C648 CSoutput.t39 gnd 0.05723f
C649 CSoutput.t79 gnd 0.05723f
C650 CSoutput.n90 gnd 0.442307f
C651 CSoutput.n91 gnd 0.221219f
C652 CSoutput.t54 gnd 0.05723f
C653 CSoutput.t92 gnd 0.05723f
C654 CSoutput.n92 gnd 0.442307f
C655 CSoutput.n93 gnd 0.405665f
C656 CSoutput.t47 gnd 0.05723f
C657 CSoutput.t20 gnd 0.05723f
C658 CSoutput.n94 gnd 0.443097f
C659 CSoutput.t4 gnd 0.05723f
C660 CSoutput.t49 gnd 0.05723f
C661 CSoutput.n95 gnd 0.442307f
C662 CSoutput.n96 gnd 0.448941f
C663 CSoutput.t44 gnd 0.05723f
C664 CSoutput.t17 gnd 0.05723f
C665 CSoutput.n97 gnd 0.442307f
C666 CSoutput.n98 gnd 0.221219f
C667 CSoutput.t3 gnd 0.05723f
C668 CSoutput.t1 gnd 0.05723f
C669 CSoutput.n99 gnd 0.442307f
C670 CSoutput.n100 gnd 0.221219f
C671 CSoutput.t63 gnd 0.05723f
C672 CSoutput.t30 gnd 0.05723f
C673 CSoutput.n101 gnd 0.442307f
C674 CSoutput.n102 gnd 0.221219f
C675 CSoutput.t27 gnd 0.05723f
C676 CSoutput.t0 gnd 0.05723f
C677 CSoutput.n103 gnd 0.442307f
C678 CSoutput.n104 gnd 0.221219f
C679 CSoutput.t83 gnd 0.05723f
C680 CSoutput.t60 gnd 0.05723f
C681 CSoutput.n105 gnd 0.442307f
C682 CSoutput.n106 gnd 0.221219f
C683 CSoutput.t48 gnd 0.05723f
C684 CSoutput.t21 gnd 0.05723f
C685 CSoutput.n107 gnd 0.442307f
C686 CSoutput.n108 gnd 0.329893f
C687 CSoutput.n109 gnd 0.415993f
C688 CSoutput.t57 gnd 0.05723f
C689 CSoutput.t32 gnd 0.05723f
C690 CSoutput.n110 gnd 0.443097f
C691 CSoutput.t14 gnd 0.05723f
C692 CSoutput.t58 gnd 0.05723f
C693 CSoutput.n111 gnd 0.442307f
C694 CSoutput.n112 gnd 0.448941f
C695 CSoutput.t55 gnd 0.05723f
C696 CSoutput.t29 gnd 0.05723f
C697 CSoutput.n113 gnd 0.442307f
C698 CSoutput.n114 gnd 0.221219f
C699 CSoutput.t13 gnd 0.05723f
C700 CSoutput.t12 gnd 0.05723f
C701 CSoutput.n115 gnd 0.442307f
C702 CSoutput.n116 gnd 0.221219f
C703 CSoutput.t70 gnd 0.05723f
C704 CSoutput.t40 gnd 0.05723f
C705 CSoutput.n117 gnd 0.442307f
C706 CSoutput.n118 gnd 0.221219f
C707 CSoutput.t36 gnd 0.05723f
C708 CSoutput.t9 gnd 0.05723f
C709 CSoutput.n119 gnd 0.442307f
C710 CSoutput.n120 gnd 0.221219f
C711 CSoutput.t93 gnd 0.05723f
C712 CSoutput.t69 gnd 0.05723f
C713 CSoutput.n121 gnd 0.442307f
C714 CSoutput.n122 gnd 0.221219f
C715 CSoutput.t56 gnd 0.05723f
C716 CSoutput.t31 gnd 0.05723f
C717 CSoutput.n123 gnd 0.442307f
C718 CSoutput.n124 gnd 0.329893f
C719 CSoutput.n125 gnd 0.464974f
C720 CSoutput.n126 gnd 9.317969f
C721 CSoutput.n128 gnd 0.811631f
C722 CSoutput.n129 gnd 0.608723f
C723 CSoutput.n130 gnd 0.811631f
C724 CSoutput.n131 gnd 0.811631f
C725 CSoutput.n132 gnd 2.18516f
C726 CSoutput.n133 gnd 0.811631f
C727 CSoutput.n134 gnd 0.811631f
C728 CSoutput.t230 gnd 1.01454f
C729 CSoutput.n135 gnd 0.811631f
C730 CSoutput.n136 gnd 0.811631f
C731 CSoutput.n140 gnd 0.811631f
C732 CSoutput.n144 gnd 0.811631f
C733 CSoutput.n145 gnd 0.811631f
C734 CSoutput.n147 gnd 0.811631f
C735 CSoutput.n152 gnd 0.811631f
C736 CSoutput.n154 gnd 0.811631f
C737 CSoutput.n155 gnd 0.811631f
C738 CSoutput.n157 gnd 0.811631f
C739 CSoutput.n158 gnd 0.811631f
C740 CSoutput.n160 gnd 0.811631f
C741 CSoutput.t219 gnd 13.562301f
C742 CSoutput.n162 gnd 0.811631f
C743 CSoutput.n163 gnd 0.608723f
C744 CSoutput.n164 gnd 0.811631f
C745 CSoutput.n165 gnd 0.811631f
C746 CSoutput.n166 gnd 2.18516f
C747 CSoutput.n167 gnd 0.811631f
C748 CSoutput.n168 gnd 0.811631f
C749 CSoutput.t237 gnd 1.01454f
C750 CSoutput.n169 gnd 0.811631f
C751 CSoutput.n170 gnd 0.811631f
C752 CSoutput.n174 gnd 0.811631f
C753 CSoutput.n178 gnd 0.811631f
C754 CSoutput.n179 gnd 0.811631f
C755 CSoutput.n181 gnd 0.811631f
C756 CSoutput.n186 gnd 0.811631f
C757 CSoutput.n188 gnd 0.811631f
C758 CSoutput.n189 gnd 0.811631f
C759 CSoutput.n191 gnd 0.811631f
C760 CSoutput.n192 gnd 0.811631f
C761 CSoutput.n194 gnd 0.811631f
C762 CSoutput.n195 gnd 0.608723f
C763 CSoutput.n197 gnd 0.811631f
C764 CSoutput.n198 gnd 0.608723f
C765 CSoutput.n199 gnd 0.811631f
C766 CSoutput.n200 gnd 0.811631f
C767 CSoutput.n201 gnd 2.18516f
C768 CSoutput.n202 gnd 0.811631f
C769 CSoutput.n203 gnd 0.811631f
C770 CSoutput.t232 gnd 1.01454f
C771 CSoutput.n204 gnd 0.811631f
C772 CSoutput.n205 gnd 2.18516f
C773 CSoutput.n207 gnd 0.811631f
C774 CSoutput.n208 gnd 0.811631f
C775 CSoutput.n210 gnd 0.811631f
C776 CSoutput.n211 gnd 0.811631f
C777 CSoutput.t216 gnd 13.3412f
C778 CSoutput.t222 gnd 13.562301f
C779 CSoutput.n217 gnd 2.54621f
C780 CSoutput.n218 gnd 10.372299f
C781 CSoutput.n219 gnd 10.8063f
C782 CSoutput.n224 gnd 2.75823f
C783 CSoutput.n230 gnd 0.811631f
C784 CSoutput.n232 gnd 0.811631f
C785 CSoutput.n234 gnd 0.811631f
C786 CSoutput.n236 gnd 0.811631f
C787 CSoutput.n238 gnd 0.811631f
C788 CSoutput.n244 gnd 0.811631f
C789 CSoutput.n251 gnd 1.48903f
C790 CSoutput.n252 gnd 1.48903f
C791 CSoutput.n253 gnd 0.811631f
C792 CSoutput.n254 gnd 0.811631f
C793 CSoutput.n256 gnd 0.608723f
C794 CSoutput.n257 gnd 0.521317f
C795 CSoutput.n259 gnd 0.608723f
C796 CSoutput.n260 gnd 0.521317f
C797 CSoutput.n261 gnd 0.608723f
C798 CSoutput.n263 gnd 0.811631f
C799 CSoutput.n265 gnd 2.18516f
C800 CSoutput.n266 gnd 2.54621f
C801 CSoutput.n267 gnd 9.53986f
C802 CSoutput.n269 gnd 0.608723f
C803 CSoutput.n270 gnd 1.56628f
C804 CSoutput.n271 gnd 0.608723f
C805 CSoutput.n273 gnd 0.811631f
C806 CSoutput.n275 gnd 2.18516f
C807 CSoutput.n276 gnd 4.75963f
C808 CSoutput.t42 gnd 0.05723f
C809 CSoutput.t24 gnd 0.05723f
C810 CSoutput.n277 gnd 0.443097f
C811 CSoutput.t76 gnd 0.05723f
C812 CSoutput.t10 gnd 0.05723f
C813 CSoutput.n278 gnd 0.442307f
C814 CSoutput.n279 gnd 0.448941f
C815 CSoutput.t61 gnd 0.05723f
C816 CSoutput.t15 gnd 0.05723f
C817 CSoutput.n280 gnd 0.442307f
C818 CSoutput.n281 gnd 0.221219f
C819 CSoutput.t72 gnd 0.05723f
C820 CSoutput.t33 gnd 0.05723f
C821 CSoutput.n282 gnd 0.442307f
C822 CSoutput.n283 gnd 0.221219f
C823 CSoutput.t84 gnd 0.05723f
C824 CSoutput.t45 gnd 0.05723f
C825 CSoutput.n284 gnd 0.442307f
C826 CSoutput.n285 gnd 0.221219f
C827 CSoutput.t66 gnd 0.05723f
C828 CSoutput.t26 gnd 0.05723f
C829 CSoutput.n286 gnd 0.442307f
C830 CSoutput.n287 gnd 0.221219f
C831 CSoutput.t78 gnd 0.05723f
C832 CSoutput.t38 gnd 0.05723f
C833 CSoutput.n288 gnd 0.442307f
C834 CSoutput.n289 gnd 0.221219f
C835 CSoutput.t91 gnd 0.05723f
C836 CSoutput.t52 gnd 0.05723f
C837 CSoutput.n290 gnd 0.442307f
C838 CSoutput.n291 gnd 0.405665f
C839 CSoutput.t80 gnd 0.05723f
C840 CSoutput.t82 gnd 0.05723f
C841 CSoutput.n292 gnd 0.443097f
C842 CSoutput.t8 gnd 0.05723f
C843 CSoutput.t68 gnd 0.05723f
C844 CSoutput.n293 gnd 0.442307f
C845 CSoutput.n294 gnd 0.448941f
C846 CSoutput.t75 gnd 0.05723f
C847 CSoutput.t5 gnd 0.05723f
C848 CSoutput.n295 gnd 0.442307f
C849 CSoutput.n296 gnd 0.221219f
C850 CSoutput.t41 gnd 0.05723f
C851 CSoutput.t65 gnd 0.05723f
C852 CSoutput.n297 gnd 0.442307f
C853 CSoutput.n298 gnd 0.221219f
C854 CSoutput.t87 gnd 0.05723f
C855 CSoutput.t28 gnd 0.05723f
C856 CSoutput.n299 gnd 0.442307f
C857 CSoutput.n300 gnd 0.221219f
C858 CSoutput.t64 gnd 0.05723f
C859 CSoutput.t94 gnd 0.05723f
C860 CSoutput.n301 gnd 0.442307f
C861 CSoutput.n302 gnd 0.221219f
C862 CSoutput.t23 gnd 0.05723f
C863 CSoutput.t51 gnd 0.05723f
C864 CSoutput.n303 gnd 0.442307f
C865 CSoutput.n304 gnd 0.221219f
C866 CSoutput.t81 gnd 0.05723f
C867 CSoutput.t7 gnd 0.05723f
C868 CSoutput.n305 gnd 0.442307f
C869 CSoutput.n306 gnd 0.329893f
C870 CSoutput.n307 gnd 0.415993f
C871 CSoutput.t88 gnd 0.05723f
C872 CSoutput.t90 gnd 0.05723f
C873 CSoutput.n308 gnd 0.443097f
C874 CSoutput.t22 gnd 0.05723f
C875 CSoutput.t74 gnd 0.05723f
C876 CSoutput.n309 gnd 0.442307f
C877 CSoutput.n310 gnd 0.448941f
C878 CSoutput.t86 gnd 0.05723f
C879 CSoutput.t16 gnd 0.05723f
C880 CSoutput.n311 gnd 0.442307f
C881 CSoutput.n312 gnd 0.221219f
C882 CSoutput.t53 gnd 0.05723f
C883 CSoutput.t73 gnd 0.05723f
C884 CSoutput.n313 gnd 0.442307f
C885 CSoutput.n314 gnd 0.221219f
C886 CSoutput.t2 gnd 0.05723f
C887 CSoutput.t37 gnd 0.05723f
C888 CSoutput.n315 gnd 0.442307f
C889 CSoutput.n316 gnd 0.221219f
C890 CSoutput.t71 gnd 0.05723f
C891 CSoutput.t6 gnd 0.05723f
C892 CSoutput.n317 gnd 0.442307f
C893 CSoutput.n318 gnd 0.221219f
C894 CSoutput.t35 gnd 0.05723f
C895 CSoutput.t59 gnd 0.05723f
C896 CSoutput.n319 gnd 0.442307f
C897 CSoutput.n320 gnd 0.221219f
C898 CSoutput.t89 gnd 0.05723f
C899 CSoutput.t19 gnd 0.05723f
C900 CSoutput.n321 gnd 0.442305f
C901 CSoutput.n322 gnd 0.329895f
C902 CSoutput.n323 gnd 0.464974f
C903 CSoutput.n324 gnd 13.0127f
C904 CSoutput.t144 gnd 0.050077f
C905 CSoutput.t212 gnd 0.050077f
C906 CSoutput.n325 gnd 0.443975f
C907 CSoutput.t134 gnd 0.050077f
C908 CSoutput.t143 gnd 0.050077f
C909 CSoutput.n326 gnd 0.442494f
C910 CSoutput.n327 gnd 0.412322f
C911 CSoutput.t124 gnd 0.050077f
C912 CSoutput.t150 gnd 0.050077f
C913 CSoutput.n328 gnd 0.442494f
C914 CSoutput.n329 gnd 0.203255f
C915 CSoutput.t171 gnd 0.050077f
C916 CSoutput.t137 gnd 0.050077f
C917 CSoutput.n330 gnd 0.442494f
C918 CSoutput.n331 gnd 0.203255f
C919 CSoutput.t147 gnd 0.050077f
C920 CSoutput.t202 gnd 0.050077f
C921 CSoutput.n332 gnd 0.442494f
C922 CSoutput.n333 gnd 0.203255f
C923 CSoutput.t164 gnd 0.050077f
C924 CSoutput.t178 gnd 0.050077f
C925 CSoutput.n334 gnd 0.442494f
C926 CSoutput.n335 gnd 0.203255f
C927 CSoutput.t119 gnd 0.050077f
C928 CSoutput.t151 gnd 0.050077f
C929 CSoutput.n336 gnd 0.442494f
C930 CSoutput.n337 gnd 0.203255f
C931 CSoutput.t105 gnd 0.050077f
C932 CSoutput.t131 gnd 0.050077f
C933 CSoutput.n338 gnd 0.442494f
C934 CSoutput.n339 gnd 0.203255f
C935 CSoutput.t184 gnd 0.050077f
C936 CSoutput.t195 gnd 0.050077f
C937 CSoutput.n340 gnd 0.442494f
C938 CSoutput.n341 gnd 0.203255f
C939 CSoutput.t211 gnd 0.050077f
C940 CSoutput.t155 gnd 0.050077f
C941 CSoutput.n342 gnd 0.442494f
C942 CSoutput.n343 gnd 0.374893f
C943 CSoutput.t207 gnd 0.050077f
C944 CSoutput.t97 gnd 0.050077f
C945 CSoutput.n344 gnd 0.443975f
C946 CSoutput.t109 gnd 0.050077f
C947 CSoutput.t200 gnd 0.050077f
C948 CSoutput.n345 gnd 0.442494f
C949 CSoutput.n346 gnd 0.412322f
C950 CSoutput.t99 gnd 0.050077f
C951 CSoutput.t190 gnd 0.050077f
C952 CSoutput.n347 gnd 0.442494f
C953 CSoutput.n348 gnd 0.203255f
C954 CSoutput.t201 gnd 0.050077f
C955 CSoutput.t98 gnd 0.050077f
C956 CSoutput.n349 gnd 0.442494f
C957 CSoutput.n350 gnd 0.203255f
C958 CSoutput.t180 gnd 0.050077f
C959 CSoutput.t154 gnd 0.050077f
C960 CSoutput.n351 gnd 0.442494f
C961 CSoutput.n352 gnd 0.203255f
C962 CSoutput.t100 gnd 0.050077f
C963 CSoutput.t182 gnd 0.050077f
C964 CSoutput.n353 gnd 0.442494f
C965 CSoutput.n354 gnd 0.203255f
C966 CSoutput.t157 gnd 0.050077f
C967 CSoutput.t165 gnd 0.050077f
C968 CSoutput.n355 gnd 0.442494f
C969 CSoutput.n356 gnd 0.203255f
C970 CSoutput.t181 gnd 0.050077f
C971 CSoutput.t156 gnd 0.050077f
C972 CSoutput.n357 gnd 0.442494f
C973 CSoutput.n358 gnd 0.203255f
C974 CSoutput.t166 gnd 0.050077f
C975 CSoutput.t170 gnd 0.050077f
C976 CSoutput.n359 gnd 0.442494f
C977 CSoutput.n360 gnd 0.203255f
C978 CSoutput.t148 gnd 0.050077f
C979 CSoutput.t161 gnd 0.050077f
C980 CSoutput.n361 gnd 0.442494f
C981 CSoutput.n362 gnd 0.308585f
C982 CSoutput.n363 gnd 0.389222f
C983 CSoutput.t112 gnd 0.050077f
C984 CSoutput.t203 gnd 0.050077f
C985 CSoutput.n364 gnd 0.443975f
C986 CSoutput.t132 gnd 0.050077f
C987 CSoutput.t138 gnd 0.050077f
C988 CSoutput.n365 gnd 0.442494f
C989 CSoutput.n366 gnd 0.412322f
C990 CSoutput.t101 gnd 0.050077f
C991 CSoutput.t185 gnd 0.050077f
C992 CSoutput.n367 gnd 0.442494f
C993 CSoutput.n368 gnd 0.203255f
C994 CSoutput.t146 gnd 0.050077f
C995 CSoutput.t113 gnd 0.050077f
C996 CSoutput.n369 gnd 0.442494f
C997 CSoutput.n370 gnd 0.203255f
C998 CSoutput.t122 gnd 0.050077f
C999 CSoutput.t215 gnd 0.050077f
C1000 CSoutput.n371 gnd 0.442494f
C1001 CSoutput.n372 gnd 0.203255f
C1002 CSoutput.t123 gnd 0.050077f
C1003 CSoutput.t127 gnd 0.050077f
C1004 CSoutput.n373 gnd 0.442494f
C1005 CSoutput.n374 gnd 0.203255f
C1006 CSoutput.t108 gnd 0.050077f
C1007 CSoutput.t199 gnd 0.050077f
C1008 CSoutput.n375 gnd 0.442494f
C1009 CSoutput.n376 gnd 0.203255f
C1010 CSoutput.t130 gnd 0.050077f
C1011 CSoutput.t120 gnd 0.050077f
C1012 CSoutput.n377 gnd 0.442494f
C1013 CSoutput.n378 gnd 0.203255f
C1014 CSoutput.t96 gnd 0.050077f
C1015 CSoutput.t140 gnd 0.050077f
C1016 CSoutput.n379 gnd 0.442494f
C1017 CSoutput.n380 gnd 0.203255f
C1018 CSoutput.t145 gnd 0.050077f
C1019 CSoutput.t111 gnd 0.050077f
C1020 CSoutput.n381 gnd 0.442494f
C1021 CSoutput.n382 gnd 0.308585f
C1022 CSoutput.n383 gnd 0.417963f
C1023 CSoutput.n384 gnd 13.2788f
C1024 CSoutput.t126 gnd 0.050077f
C1025 CSoutput.t183 gnd 0.050077f
C1026 CSoutput.n385 gnd 0.443975f
C1027 CSoutput.t179 gnd 0.050077f
C1028 CSoutput.t153 gnd 0.050077f
C1029 CSoutput.n386 gnd 0.442494f
C1030 CSoutput.n387 gnd 0.412322f
C1031 CSoutput.t187 gnd 0.050077f
C1032 CSoutput.t141 gnd 0.050077f
C1033 CSoutput.n388 gnd 0.442494f
C1034 CSoutput.n389 gnd 0.203255f
C1035 CSoutput.t167 gnd 0.050077f
C1036 CSoutput.t205 gnd 0.050077f
C1037 CSoutput.n390 gnd 0.442494f
C1038 CSoutput.n391 gnd 0.203255f
C1039 CSoutput.t121 gnd 0.050077f
C1040 CSoutput.t186 gnd 0.050077f
C1041 CSoutput.n392 gnd 0.442494f
C1042 CSoutput.n393 gnd 0.203255f
C1043 CSoutput.t107 gnd 0.050077f
C1044 CSoutput.t193 gnd 0.050077f
C1045 CSoutput.n394 gnd 0.442494f
C1046 CSoutput.n395 gnd 0.203255f
C1047 CSoutput.t192 gnd 0.050077f
C1048 CSoutput.t133 gnd 0.050077f
C1049 CSoutput.n396 gnd 0.442494f
C1050 CSoutput.n397 gnd 0.203255f
C1051 CSoutput.t160 gnd 0.050077f
C1052 CSoutput.t129 gnd 0.050077f
C1053 CSoutput.n398 gnd 0.442494f
C1054 CSoutput.n399 gnd 0.203255f
C1055 CSoutput.t135 gnd 0.050077f
C1056 CSoutput.t110 gnd 0.050077f
C1057 CSoutput.n400 gnd 0.442494f
C1058 CSoutput.n401 gnd 0.203255f
C1059 CSoutput.t118 gnd 0.050077f
C1060 CSoutput.t136 gnd 0.050077f
C1061 CSoutput.n402 gnd 0.442494f
C1062 CSoutput.n403 gnd 0.374893f
C1063 CSoutput.t115 gnd 0.050077f
C1064 CSoutput.t106 gnd 0.050077f
C1065 CSoutput.n404 gnd 0.443975f
C1066 CSoutput.t102 gnd 0.050077f
C1067 CSoutput.t213 gnd 0.050077f
C1068 CSoutput.n405 gnd 0.442494f
C1069 CSoutput.n406 gnd 0.412322f
C1070 CSoutput.t214 gnd 0.050077f
C1071 CSoutput.t116 gnd 0.050077f
C1072 CSoutput.n407 gnd 0.442494f
C1073 CSoutput.n408 gnd 0.203255f
C1074 CSoutput.t117 gnd 0.050077f
C1075 CSoutput.t174 gnd 0.050077f
C1076 CSoutput.n409 gnd 0.442494f
C1077 CSoutput.n410 gnd 0.203255f
C1078 CSoutput.t175 gnd 0.050077f
C1079 CSoutput.t206 gnd 0.050077f
C1080 CSoutput.n411 gnd 0.442494f
C1081 CSoutput.n412 gnd 0.203255f
C1082 CSoutput.t209 gnd 0.050077f
C1083 CSoutput.t198 gnd 0.050077f
C1084 CSoutput.n413 gnd 0.442494f
C1085 CSoutput.n414 gnd 0.203255f
C1086 CSoutput.t189 gnd 0.050077f
C1087 CSoutput.t176 gnd 0.050077f
C1088 CSoutput.n415 gnd 0.442494f
C1089 CSoutput.n416 gnd 0.203255f
C1090 CSoutput.t177 gnd 0.050077f
C1091 CSoutput.t210 gnd 0.050077f
C1092 CSoutput.n417 gnd 0.442494f
C1093 CSoutput.n418 gnd 0.203255f
C1094 CSoutput.t163 gnd 0.050077f
C1095 CSoutput.t191 gnd 0.050077f
C1096 CSoutput.n419 gnd 0.442494f
C1097 CSoutput.n420 gnd 0.203255f
C1098 CSoutput.t197 gnd 0.050077f
C1099 CSoutput.t172 gnd 0.050077f
C1100 CSoutput.n421 gnd 0.442494f
C1101 CSoutput.n422 gnd 0.308585f
C1102 CSoutput.n423 gnd 0.389222f
C1103 CSoutput.t162 gnd 0.050077f
C1104 CSoutput.t194 gnd 0.050077f
C1105 CSoutput.n424 gnd 0.443975f
C1106 CSoutput.t125 gnd 0.050077f
C1107 CSoutput.t142 gnd 0.050077f
C1108 CSoutput.n425 gnd 0.442494f
C1109 CSoutput.n426 gnd 0.412322f
C1110 CSoutput.t152 gnd 0.050077f
C1111 CSoutput.t173 gnd 0.050077f
C1112 CSoutput.n427 gnd 0.442494f
C1113 CSoutput.n428 gnd 0.203255f
C1114 CSoutput.t196 gnd 0.050077f
C1115 CSoutput.t158 gnd 0.050077f
C1116 CSoutput.n429 gnd 0.442494f
C1117 CSoutput.n430 gnd 0.203255f
C1118 CSoutput.t168 gnd 0.050077f
C1119 CSoutput.t208 gnd 0.050077f
C1120 CSoutput.n431 gnd 0.442494f
C1121 CSoutput.n432 gnd 0.203255f
C1122 CSoutput.t103 gnd 0.050077f
C1123 CSoutput.t128 gnd 0.050077f
C1124 CSoutput.n433 gnd 0.442494f
C1125 CSoutput.n434 gnd 0.203255f
C1126 CSoutput.t159 gnd 0.050077f
C1127 CSoutput.t188 gnd 0.050077f
C1128 CSoutput.n435 gnd 0.442494f
C1129 CSoutput.n436 gnd 0.203255f
C1130 CSoutput.t204 gnd 0.050077f
C1131 CSoutput.t114 gnd 0.050077f
C1132 CSoutput.n437 gnd 0.442494f
C1133 CSoutput.n438 gnd 0.203255f
C1134 CSoutput.t149 gnd 0.050077f
C1135 CSoutput.t169 gnd 0.050077f
C1136 CSoutput.n439 gnd 0.442494f
C1137 CSoutput.n440 gnd 0.203255f
C1138 CSoutput.t104 gnd 0.050077f
C1139 CSoutput.t139 gnd 0.050077f
C1140 CSoutput.n441 gnd 0.442494f
C1141 CSoutput.n442 gnd 0.308585f
C1142 CSoutput.n443 gnd 0.417963f
C1143 CSoutput.n444 gnd 7.98289f
C1144 CSoutput.n445 gnd 13.8985f
C1145 commonsourceibias.n0 gnd 0.012817f
C1146 commonsourceibias.t151 gnd 0.194086f
C1147 commonsourceibias.t83 gnd 0.17946f
C1148 commonsourceibias.n1 gnd 0.009349f
C1149 commonsourceibias.n2 gnd 0.009605f
C1150 commonsourceibias.t161 gnd 0.17946f
C1151 commonsourceibias.n3 gnd 0.012358f
C1152 commonsourceibias.n4 gnd 0.009605f
C1153 commonsourceibias.t152 gnd 0.17946f
C1154 commonsourceibias.n5 gnd 0.071604f
C1155 commonsourceibias.t171 gnd 0.17946f
C1156 commonsourceibias.n6 gnd 0.009057f
C1157 commonsourceibias.n7 gnd 0.009605f
C1158 commonsourceibias.t145 gnd 0.17946f
C1159 commonsourceibias.n8 gnd 0.012174f
C1160 commonsourceibias.n9 gnd 0.009605f
C1161 commonsourceibias.t124 gnd 0.17946f
C1162 commonsourceibias.n10 gnd 0.071604f
C1163 commonsourceibias.t158 gnd 0.17946f
C1164 commonsourceibias.n11 gnd 0.008798f
C1165 commonsourceibias.n12 gnd 0.009605f
C1166 commonsourceibias.t148 gnd 0.17946f
C1167 commonsourceibias.n13 gnd 0.01197f
C1168 commonsourceibias.n14 gnd 0.012817f
C1169 commonsourceibias.t16 gnd 0.194086f
C1170 commonsourceibias.t60 gnd 0.17946f
C1171 commonsourceibias.n15 gnd 0.009349f
C1172 commonsourceibias.n16 gnd 0.009605f
C1173 commonsourceibias.t4 gnd 0.17946f
C1174 commonsourceibias.n17 gnd 0.012358f
C1175 commonsourceibias.n18 gnd 0.009605f
C1176 commonsourceibias.t14 gnd 0.17946f
C1177 commonsourceibias.n19 gnd 0.071604f
C1178 commonsourceibias.t74 gnd 0.17946f
C1179 commonsourceibias.n20 gnd 0.009057f
C1180 commonsourceibias.n21 gnd 0.009605f
C1181 commonsourceibias.t20 gnd 0.17946f
C1182 commonsourceibias.n22 gnd 0.012174f
C1183 commonsourceibias.n23 gnd 0.009605f
C1184 commonsourceibias.t34 gnd 0.17946f
C1185 commonsourceibias.n24 gnd 0.071604f
C1186 commonsourceibias.t10 gnd 0.17946f
C1187 commonsourceibias.n25 gnd 0.008798f
C1188 commonsourceibias.n26 gnd 0.009605f
C1189 commonsourceibias.t18 gnd 0.17946f
C1190 commonsourceibias.n27 gnd 0.01197f
C1191 commonsourceibias.n28 gnd 0.009605f
C1192 commonsourceibias.t54 gnd 0.17946f
C1193 commonsourceibias.n29 gnd 0.071604f
C1194 commonsourceibias.t30 gnd 0.17946f
C1195 commonsourceibias.n30 gnd 0.008571f
C1196 commonsourceibias.n31 gnd 0.009605f
C1197 commonsourceibias.t36 gnd 0.17946f
C1198 commonsourceibias.n32 gnd 0.011742f
C1199 commonsourceibias.n33 gnd 0.009605f
C1200 commonsourceibias.t70 gnd 0.17946f
C1201 commonsourceibias.n34 gnd 0.071604f
C1202 commonsourceibias.t22 gnd 0.17946f
C1203 commonsourceibias.n35 gnd 0.008375f
C1204 commonsourceibias.n36 gnd 0.009605f
C1205 commonsourceibias.t62 gnd 0.17946f
C1206 commonsourceibias.n37 gnd 0.011489f
C1207 commonsourceibias.n38 gnd 0.009605f
C1208 commonsourceibias.t0 gnd 0.17946f
C1209 commonsourceibias.n39 gnd 0.071604f
C1210 commonsourceibias.t42 gnd 0.17946f
C1211 commonsourceibias.n40 gnd 0.008208f
C1212 commonsourceibias.n41 gnd 0.009605f
C1213 commonsourceibias.t52 gnd 0.17946f
C1214 commonsourceibias.n42 gnd 0.011208f
C1215 commonsourceibias.t26 gnd 0.199526f
C1216 commonsourceibias.t58 gnd 0.17946f
C1217 commonsourceibias.n43 gnd 0.078221f
C1218 commonsourceibias.n44 gnd 0.085838f
C1219 commonsourceibias.n45 gnd 0.03983f
C1220 commonsourceibias.n46 gnd 0.009605f
C1221 commonsourceibias.n47 gnd 0.009349f
C1222 commonsourceibias.n48 gnd 0.013398f
C1223 commonsourceibias.n49 gnd 0.071604f
C1224 commonsourceibias.n50 gnd 0.013389f
C1225 commonsourceibias.n51 gnd 0.009605f
C1226 commonsourceibias.n52 gnd 0.009605f
C1227 commonsourceibias.n53 gnd 0.009605f
C1228 commonsourceibias.n54 gnd 0.012358f
C1229 commonsourceibias.n55 gnd 0.071604f
C1230 commonsourceibias.n56 gnd 0.012648f
C1231 commonsourceibias.n57 gnd 0.012288f
C1232 commonsourceibias.n58 gnd 0.009605f
C1233 commonsourceibias.n59 gnd 0.009605f
C1234 commonsourceibias.n60 gnd 0.009605f
C1235 commonsourceibias.n61 gnd 0.009057f
C1236 commonsourceibias.n62 gnd 0.01341f
C1237 commonsourceibias.n63 gnd 0.071604f
C1238 commonsourceibias.n64 gnd 0.013406f
C1239 commonsourceibias.n65 gnd 0.009605f
C1240 commonsourceibias.n66 gnd 0.009605f
C1241 commonsourceibias.n67 gnd 0.009605f
C1242 commonsourceibias.n68 gnd 0.012174f
C1243 commonsourceibias.n69 gnd 0.071604f
C1244 commonsourceibias.n70 gnd 0.012558f
C1245 commonsourceibias.n71 gnd 0.012378f
C1246 commonsourceibias.n72 gnd 0.009605f
C1247 commonsourceibias.n73 gnd 0.009605f
C1248 commonsourceibias.n74 gnd 0.009605f
C1249 commonsourceibias.n75 gnd 0.008798f
C1250 commonsourceibias.n76 gnd 0.013415f
C1251 commonsourceibias.n77 gnd 0.071604f
C1252 commonsourceibias.n78 gnd 0.013414f
C1253 commonsourceibias.n79 gnd 0.009605f
C1254 commonsourceibias.n80 gnd 0.009605f
C1255 commonsourceibias.n81 gnd 0.009605f
C1256 commonsourceibias.n82 gnd 0.01197f
C1257 commonsourceibias.n83 gnd 0.071604f
C1258 commonsourceibias.n84 gnd 0.012468f
C1259 commonsourceibias.n85 gnd 0.012468f
C1260 commonsourceibias.n86 gnd 0.009605f
C1261 commonsourceibias.n87 gnd 0.009605f
C1262 commonsourceibias.n88 gnd 0.009605f
C1263 commonsourceibias.n89 gnd 0.008571f
C1264 commonsourceibias.n90 gnd 0.013414f
C1265 commonsourceibias.n91 gnd 0.071604f
C1266 commonsourceibias.n92 gnd 0.013415f
C1267 commonsourceibias.n93 gnd 0.009605f
C1268 commonsourceibias.n94 gnd 0.009605f
C1269 commonsourceibias.n95 gnd 0.009605f
C1270 commonsourceibias.n96 gnd 0.011742f
C1271 commonsourceibias.n97 gnd 0.071604f
C1272 commonsourceibias.n98 gnd 0.012378f
C1273 commonsourceibias.n99 gnd 0.012558f
C1274 commonsourceibias.n100 gnd 0.009605f
C1275 commonsourceibias.n101 gnd 0.009605f
C1276 commonsourceibias.n102 gnd 0.009605f
C1277 commonsourceibias.n103 gnd 0.008375f
C1278 commonsourceibias.n104 gnd 0.013406f
C1279 commonsourceibias.n105 gnd 0.071604f
C1280 commonsourceibias.n106 gnd 0.01341f
C1281 commonsourceibias.n107 gnd 0.009605f
C1282 commonsourceibias.n108 gnd 0.009605f
C1283 commonsourceibias.n109 gnd 0.009605f
C1284 commonsourceibias.n110 gnd 0.011489f
C1285 commonsourceibias.n111 gnd 0.071604f
C1286 commonsourceibias.n112 gnd 0.012288f
C1287 commonsourceibias.n113 gnd 0.012648f
C1288 commonsourceibias.n114 gnd 0.009605f
C1289 commonsourceibias.n115 gnd 0.009605f
C1290 commonsourceibias.n116 gnd 0.009605f
C1291 commonsourceibias.n117 gnd 0.008208f
C1292 commonsourceibias.n118 gnd 0.013389f
C1293 commonsourceibias.n119 gnd 0.071604f
C1294 commonsourceibias.n120 gnd 0.013398f
C1295 commonsourceibias.n121 gnd 0.009605f
C1296 commonsourceibias.n122 gnd 0.009605f
C1297 commonsourceibias.n123 gnd 0.009605f
C1298 commonsourceibias.n124 gnd 0.011208f
C1299 commonsourceibias.n125 gnd 0.071604f
C1300 commonsourceibias.n126 gnd 0.011785f
C1301 commonsourceibias.n127 gnd 0.085919f
C1302 commonsourceibias.n128 gnd 0.095702f
C1303 commonsourceibias.t17 gnd 0.020728f
C1304 commonsourceibias.t61 gnd 0.020728f
C1305 commonsourceibias.n129 gnd 0.183157f
C1306 commonsourceibias.n130 gnd 0.158432f
C1307 commonsourceibias.t5 gnd 0.020728f
C1308 commonsourceibias.t15 gnd 0.020728f
C1309 commonsourceibias.n131 gnd 0.183157f
C1310 commonsourceibias.n132 gnd 0.084131f
C1311 commonsourceibias.t75 gnd 0.020728f
C1312 commonsourceibias.t21 gnd 0.020728f
C1313 commonsourceibias.n133 gnd 0.183157f
C1314 commonsourceibias.n134 gnd 0.084131f
C1315 commonsourceibias.t35 gnd 0.020728f
C1316 commonsourceibias.t11 gnd 0.020728f
C1317 commonsourceibias.n135 gnd 0.183157f
C1318 commonsourceibias.n136 gnd 0.084131f
C1319 commonsourceibias.t19 gnd 0.020728f
C1320 commonsourceibias.t55 gnd 0.020728f
C1321 commonsourceibias.n137 gnd 0.183157f
C1322 commonsourceibias.n138 gnd 0.070287f
C1323 commonsourceibias.t59 gnd 0.020728f
C1324 commonsourceibias.t27 gnd 0.020728f
C1325 commonsourceibias.n139 gnd 0.18377f
C1326 commonsourceibias.t43 gnd 0.020728f
C1327 commonsourceibias.t53 gnd 0.020728f
C1328 commonsourceibias.n140 gnd 0.183157f
C1329 commonsourceibias.n141 gnd 0.170668f
C1330 commonsourceibias.t63 gnd 0.020728f
C1331 commonsourceibias.t1 gnd 0.020728f
C1332 commonsourceibias.n142 gnd 0.183157f
C1333 commonsourceibias.n143 gnd 0.084131f
C1334 commonsourceibias.t71 gnd 0.020728f
C1335 commonsourceibias.t23 gnd 0.020728f
C1336 commonsourceibias.n144 gnd 0.183157f
C1337 commonsourceibias.n145 gnd 0.084131f
C1338 commonsourceibias.t31 gnd 0.020728f
C1339 commonsourceibias.t37 gnd 0.020728f
C1340 commonsourceibias.n146 gnd 0.183157f
C1341 commonsourceibias.n147 gnd 0.070287f
C1342 commonsourceibias.n148 gnd 0.085111f
C1343 commonsourceibias.n149 gnd 0.062167f
C1344 commonsourceibias.t93 gnd 0.17946f
C1345 commonsourceibias.n150 gnd 0.071604f
C1346 commonsourceibias.t131 gnd 0.17946f
C1347 commonsourceibias.n151 gnd 0.071604f
C1348 commonsourceibias.n152 gnd 0.009605f
C1349 commonsourceibias.t117 gnd 0.17946f
C1350 commonsourceibias.n153 gnd 0.071604f
C1351 commonsourceibias.n154 gnd 0.009605f
C1352 commonsourceibias.t176 gnd 0.17946f
C1353 commonsourceibias.n155 gnd 0.071604f
C1354 commonsourceibias.n156 gnd 0.009605f
C1355 commonsourceibias.t144 gnd 0.17946f
C1356 commonsourceibias.n157 gnd 0.008375f
C1357 commonsourceibias.n158 gnd 0.009605f
C1358 commonsourceibias.t190 gnd 0.17946f
C1359 commonsourceibias.n159 gnd 0.011489f
C1360 commonsourceibias.n160 gnd 0.009605f
C1361 commonsourceibias.t164 gnd 0.17946f
C1362 commonsourceibias.n161 gnd 0.071604f
C1363 commonsourceibias.t111 gnd 0.17946f
C1364 commonsourceibias.n162 gnd 0.008208f
C1365 commonsourceibias.n163 gnd 0.009605f
C1366 commonsourceibias.t100 gnd 0.17946f
C1367 commonsourceibias.n164 gnd 0.011208f
C1368 commonsourceibias.t140 gnd 0.199526f
C1369 commonsourceibias.t84 gnd 0.17946f
C1370 commonsourceibias.n165 gnd 0.078221f
C1371 commonsourceibias.n166 gnd 0.085838f
C1372 commonsourceibias.n167 gnd 0.03983f
C1373 commonsourceibias.n168 gnd 0.009605f
C1374 commonsourceibias.n169 gnd 0.009349f
C1375 commonsourceibias.n170 gnd 0.013398f
C1376 commonsourceibias.n171 gnd 0.071604f
C1377 commonsourceibias.n172 gnd 0.013389f
C1378 commonsourceibias.n173 gnd 0.009605f
C1379 commonsourceibias.n174 gnd 0.009605f
C1380 commonsourceibias.n175 gnd 0.009605f
C1381 commonsourceibias.n176 gnd 0.012358f
C1382 commonsourceibias.n177 gnd 0.071604f
C1383 commonsourceibias.n178 gnd 0.012648f
C1384 commonsourceibias.n179 gnd 0.012288f
C1385 commonsourceibias.n180 gnd 0.009605f
C1386 commonsourceibias.n181 gnd 0.009605f
C1387 commonsourceibias.n182 gnd 0.009605f
C1388 commonsourceibias.n183 gnd 0.009057f
C1389 commonsourceibias.n184 gnd 0.01341f
C1390 commonsourceibias.n185 gnd 0.071604f
C1391 commonsourceibias.n186 gnd 0.013406f
C1392 commonsourceibias.n187 gnd 0.009605f
C1393 commonsourceibias.n188 gnd 0.009605f
C1394 commonsourceibias.n189 gnd 0.009605f
C1395 commonsourceibias.n190 gnd 0.012174f
C1396 commonsourceibias.n191 gnd 0.071604f
C1397 commonsourceibias.n192 gnd 0.012558f
C1398 commonsourceibias.n193 gnd 0.012378f
C1399 commonsourceibias.n194 gnd 0.009605f
C1400 commonsourceibias.n195 gnd 0.009605f
C1401 commonsourceibias.n196 gnd 0.011742f
C1402 commonsourceibias.n197 gnd 0.008798f
C1403 commonsourceibias.n198 gnd 0.013415f
C1404 commonsourceibias.n199 gnd 0.009605f
C1405 commonsourceibias.n200 gnd 0.009605f
C1406 commonsourceibias.n201 gnd 0.013414f
C1407 commonsourceibias.n202 gnd 0.008571f
C1408 commonsourceibias.n203 gnd 0.01197f
C1409 commonsourceibias.n204 gnd 0.009605f
C1410 commonsourceibias.n205 gnd 0.008391f
C1411 commonsourceibias.n206 gnd 0.012468f
C1412 commonsourceibias.n207 gnd 0.012468f
C1413 commonsourceibias.n208 gnd 0.008391f
C1414 commonsourceibias.n209 gnd 0.009605f
C1415 commonsourceibias.n210 gnd 0.009605f
C1416 commonsourceibias.n211 gnd 0.008571f
C1417 commonsourceibias.n212 gnd 0.013414f
C1418 commonsourceibias.n213 gnd 0.071604f
C1419 commonsourceibias.n214 gnd 0.013415f
C1420 commonsourceibias.n215 gnd 0.009605f
C1421 commonsourceibias.n216 gnd 0.009605f
C1422 commonsourceibias.n217 gnd 0.009605f
C1423 commonsourceibias.n218 gnd 0.011742f
C1424 commonsourceibias.n219 gnd 0.071604f
C1425 commonsourceibias.n220 gnd 0.012378f
C1426 commonsourceibias.n221 gnd 0.012558f
C1427 commonsourceibias.n222 gnd 0.009605f
C1428 commonsourceibias.n223 gnd 0.009605f
C1429 commonsourceibias.n224 gnd 0.009605f
C1430 commonsourceibias.n225 gnd 0.008375f
C1431 commonsourceibias.n226 gnd 0.013406f
C1432 commonsourceibias.n227 gnd 0.071604f
C1433 commonsourceibias.n228 gnd 0.01341f
C1434 commonsourceibias.n229 gnd 0.009605f
C1435 commonsourceibias.n230 gnd 0.009605f
C1436 commonsourceibias.n231 gnd 0.009605f
C1437 commonsourceibias.n232 gnd 0.011489f
C1438 commonsourceibias.n233 gnd 0.071604f
C1439 commonsourceibias.n234 gnd 0.012288f
C1440 commonsourceibias.n235 gnd 0.012648f
C1441 commonsourceibias.n236 gnd 0.009605f
C1442 commonsourceibias.n237 gnd 0.009605f
C1443 commonsourceibias.n238 gnd 0.009605f
C1444 commonsourceibias.n239 gnd 0.008208f
C1445 commonsourceibias.n240 gnd 0.013389f
C1446 commonsourceibias.n241 gnd 0.071604f
C1447 commonsourceibias.n242 gnd 0.013398f
C1448 commonsourceibias.n243 gnd 0.009605f
C1449 commonsourceibias.n244 gnd 0.009605f
C1450 commonsourceibias.n245 gnd 0.009605f
C1451 commonsourceibias.n246 gnd 0.011208f
C1452 commonsourceibias.n247 gnd 0.071604f
C1453 commonsourceibias.n248 gnd 0.011785f
C1454 commonsourceibias.n249 gnd 0.085919f
C1455 commonsourceibias.n250 gnd 0.056156f
C1456 commonsourceibias.n251 gnd 0.012817f
C1457 commonsourceibias.t88 gnd 0.194086f
C1458 commonsourceibias.t198 gnd 0.17946f
C1459 commonsourceibias.n252 gnd 0.009349f
C1460 commonsourceibias.n253 gnd 0.009605f
C1461 commonsourceibias.t186 gnd 0.17946f
C1462 commonsourceibias.n254 gnd 0.012358f
C1463 commonsourceibias.n255 gnd 0.009605f
C1464 commonsourceibias.t95 gnd 0.17946f
C1465 commonsourceibias.n256 gnd 0.071604f
C1466 commonsourceibias.t196 gnd 0.17946f
C1467 commonsourceibias.n257 gnd 0.009057f
C1468 commonsourceibias.n258 gnd 0.009605f
C1469 commonsourceibias.t105 gnd 0.17946f
C1470 commonsourceibias.n259 gnd 0.012174f
C1471 commonsourceibias.n260 gnd 0.009605f
C1472 commonsourceibias.t94 gnd 0.17946f
C1473 commonsourceibias.n261 gnd 0.071604f
C1474 commonsourceibias.t197 gnd 0.17946f
C1475 commonsourceibias.n262 gnd 0.008798f
C1476 commonsourceibias.n263 gnd 0.009605f
C1477 commonsourceibias.t115 gnd 0.17946f
C1478 commonsourceibias.n264 gnd 0.01197f
C1479 commonsourceibias.n265 gnd 0.009605f
C1480 commonsourceibias.t141 gnd 0.17946f
C1481 commonsourceibias.n266 gnd 0.071604f
C1482 commonsourceibias.t195 gnd 0.17946f
C1483 commonsourceibias.n267 gnd 0.008571f
C1484 commonsourceibias.n268 gnd 0.009605f
C1485 commonsourceibias.t113 gnd 0.17946f
C1486 commonsourceibias.n269 gnd 0.011742f
C1487 commonsourceibias.n270 gnd 0.009605f
C1488 commonsourceibias.t138 gnd 0.17946f
C1489 commonsourceibias.n271 gnd 0.071604f
C1490 commonsourceibias.t130 gnd 0.17946f
C1491 commonsourceibias.n272 gnd 0.008375f
C1492 commonsourceibias.n273 gnd 0.009605f
C1493 commonsourceibias.t114 gnd 0.17946f
C1494 commonsourceibias.n274 gnd 0.011489f
C1495 commonsourceibias.n275 gnd 0.009605f
C1496 commonsourceibias.t139 gnd 0.17946f
C1497 commonsourceibias.n276 gnd 0.071604f
C1498 commonsourceibias.t129 gnd 0.17946f
C1499 commonsourceibias.n277 gnd 0.008208f
C1500 commonsourceibias.n278 gnd 0.009605f
C1501 commonsourceibias.t125 gnd 0.17946f
C1502 commonsourceibias.n279 gnd 0.011208f
C1503 commonsourceibias.t134 gnd 0.199526f
C1504 commonsourceibias.t147 gnd 0.17946f
C1505 commonsourceibias.n280 gnd 0.078221f
C1506 commonsourceibias.n281 gnd 0.085838f
C1507 commonsourceibias.n282 gnd 0.03983f
C1508 commonsourceibias.n283 gnd 0.009605f
C1509 commonsourceibias.n284 gnd 0.009349f
C1510 commonsourceibias.n285 gnd 0.013398f
C1511 commonsourceibias.n286 gnd 0.071604f
C1512 commonsourceibias.n287 gnd 0.013389f
C1513 commonsourceibias.n288 gnd 0.009605f
C1514 commonsourceibias.n289 gnd 0.009605f
C1515 commonsourceibias.n290 gnd 0.009605f
C1516 commonsourceibias.n291 gnd 0.012358f
C1517 commonsourceibias.n292 gnd 0.071604f
C1518 commonsourceibias.n293 gnd 0.012648f
C1519 commonsourceibias.n294 gnd 0.012288f
C1520 commonsourceibias.n295 gnd 0.009605f
C1521 commonsourceibias.n296 gnd 0.009605f
C1522 commonsourceibias.n297 gnd 0.009605f
C1523 commonsourceibias.n298 gnd 0.009057f
C1524 commonsourceibias.n299 gnd 0.01341f
C1525 commonsourceibias.n300 gnd 0.071604f
C1526 commonsourceibias.n301 gnd 0.013406f
C1527 commonsourceibias.n302 gnd 0.009605f
C1528 commonsourceibias.n303 gnd 0.009605f
C1529 commonsourceibias.n304 gnd 0.009605f
C1530 commonsourceibias.n305 gnd 0.012174f
C1531 commonsourceibias.n306 gnd 0.071604f
C1532 commonsourceibias.n307 gnd 0.012558f
C1533 commonsourceibias.n308 gnd 0.012378f
C1534 commonsourceibias.n309 gnd 0.009605f
C1535 commonsourceibias.n310 gnd 0.009605f
C1536 commonsourceibias.n311 gnd 0.009605f
C1537 commonsourceibias.n312 gnd 0.008798f
C1538 commonsourceibias.n313 gnd 0.013415f
C1539 commonsourceibias.n314 gnd 0.071604f
C1540 commonsourceibias.n315 gnd 0.013414f
C1541 commonsourceibias.n316 gnd 0.009605f
C1542 commonsourceibias.n317 gnd 0.009605f
C1543 commonsourceibias.n318 gnd 0.009605f
C1544 commonsourceibias.n319 gnd 0.01197f
C1545 commonsourceibias.n320 gnd 0.071604f
C1546 commonsourceibias.n321 gnd 0.012468f
C1547 commonsourceibias.n322 gnd 0.012468f
C1548 commonsourceibias.n323 gnd 0.009605f
C1549 commonsourceibias.n324 gnd 0.009605f
C1550 commonsourceibias.n325 gnd 0.009605f
C1551 commonsourceibias.n326 gnd 0.008571f
C1552 commonsourceibias.n327 gnd 0.013414f
C1553 commonsourceibias.n328 gnd 0.071604f
C1554 commonsourceibias.n329 gnd 0.013415f
C1555 commonsourceibias.n330 gnd 0.009605f
C1556 commonsourceibias.n331 gnd 0.009605f
C1557 commonsourceibias.n332 gnd 0.009605f
C1558 commonsourceibias.n333 gnd 0.011742f
C1559 commonsourceibias.n334 gnd 0.071604f
C1560 commonsourceibias.n335 gnd 0.012378f
C1561 commonsourceibias.n336 gnd 0.012558f
C1562 commonsourceibias.n337 gnd 0.009605f
C1563 commonsourceibias.n338 gnd 0.009605f
C1564 commonsourceibias.n339 gnd 0.009605f
C1565 commonsourceibias.n340 gnd 0.008375f
C1566 commonsourceibias.n341 gnd 0.013406f
C1567 commonsourceibias.n342 gnd 0.071604f
C1568 commonsourceibias.n343 gnd 0.01341f
C1569 commonsourceibias.n344 gnd 0.009605f
C1570 commonsourceibias.n345 gnd 0.009605f
C1571 commonsourceibias.n346 gnd 0.009605f
C1572 commonsourceibias.n347 gnd 0.011489f
C1573 commonsourceibias.n348 gnd 0.071604f
C1574 commonsourceibias.n349 gnd 0.012288f
C1575 commonsourceibias.n350 gnd 0.012648f
C1576 commonsourceibias.n351 gnd 0.009605f
C1577 commonsourceibias.n352 gnd 0.009605f
C1578 commonsourceibias.n353 gnd 0.009605f
C1579 commonsourceibias.n354 gnd 0.008208f
C1580 commonsourceibias.n355 gnd 0.013389f
C1581 commonsourceibias.n356 gnd 0.071604f
C1582 commonsourceibias.n357 gnd 0.013398f
C1583 commonsourceibias.n358 gnd 0.009605f
C1584 commonsourceibias.n359 gnd 0.009605f
C1585 commonsourceibias.n360 gnd 0.009605f
C1586 commonsourceibias.n361 gnd 0.011208f
C1587 commonsourceibias.n362 gnd 0.071604f
C1588 commonsourceibias.n363 gnd 0.011785f
C1589 commonsourceibias.n364 gnd 0.085919f
C1590 commonsourceibias.n365 gnd 0.029883f
C1591 commonsourceibias.n366 gnd 0.153509f
C1592 commonsourceibias.n367 gnd 0.012817f
C1593 commonsourceibias.t92 gnd 0.17946f
C1594 commonsourceibias.n368 gnd 0.009349f
C1595 commonsourceibias.n369 gnd 0.009605f
C1596 commonsourceibias.t163 gnd 0.17946f
C1597 commonsourceibias.n370 gnd 0.012358f
C1598 commonsourceibias.n371 gnd 0.009605f
C1599 commonsourceibias.t157 gnd 0.17946f
C1600 commonsourceibias.n372 gnd 0.071604f
C1601 commonsourceibias.t194 gnd 0.17946f
C1602 commonsourceibias.n373 gnd 0.009057f
C1603 commonsourceibias.n374 gnd 0.009605f
C1604 commonsourceibias.t110 gnd 0.17946f
C1605 commonsourceibias.n375 gnd 0.012174f
C1606 commonsourceibias.n376 gnd 0.009605f
C1607 commonsourceibias.t149 gnd 0.17946f
C1608 commonsourceibias.n377 gnd 0.071604f
C1609 commonsourceibias.t182 gnd 0.17946f
C1610 commonsourceibias.n378 gnd 0.008798f
C1611 commonsourceibias.n379 gnd 0.009605f
C1612 commonsourceibias.t173 gnd 0.17946f
C1613 commonsourceibias.n380 gnd 0.01197f
C1614 commonsourceibias.n381 gnd 0.009605f
C1615 commonsourceibias.t80 gnd 0.17946f
C1616 commonsourceibias.n382 gnd 0.071604f
C1617 commonsourceibias.t172 gnd 0.17946f
C1618 commonsourceibias.n383 gnd 0.008571f
C1619 commonsourceibias.n384 gnd 0.009605f
C1620 commonsourceibias.t168 gnd 0.17946f
C1621 commonsourceibias.n385 gnd 0.011742f
C1622 commonsourceibias.n386 gnd 0.009605f
C1623 commonsourceibias.t187 gnd 0.17946f
C1624 commonsourceibias.n387 gnd 0.071604f
C1625 commonsourceibias.t96 gnd 0.17946f
C1626 commonsourceibias.n388 gnd 0.008375f
C1627 commonsourceibias.n389 gnd 0.009605f
C1628 commonsourceibias.t165 gnd 0.17946f
C1629 commonsourceibias.n390 gnd 0.011489f
C1630 commonsourceibias.n391 gnd 0.009605f
C1631 commonsourceibias.t175 gnd 0.17946f
C1632 commonsourceibias.n392 gnd 0.071604f
C1633 commonsourceibias.t199 gnd 0.17946f
C1634 commonsourceibias.n393 gnd 0.008208f
C1635 commonsourceibias.n394 gnd 0.009605f
C1636 commonsourceibias.t155 gnd 0.17946f
C1637 commonsourceibias.n395 gnd 0.011208f
C1638 commonsourceibias.t184 gnd 0.199526f
C1639 commonsourceibias.t150 gnd 0.17946f
C1640 commonsourceibias.n396 gnd 0.078221f
C1641 commonsourceibias.n397 gnd 0.085838f
C1642 commonsourceibias.n398 gnd 0.03983f
C1643 commonsourceibias.n399 gnd 0.009605f
C1644 commonsourceibias.n400 gnd 0.009349f
C1645 commonsourceibias.n401 gnd 0.013398f
C1646 commonsourceibias.n402 gnd 0.071604f
C1647 commonsourceibias.n403 gnd 0.013389f
C1648 commonsourceibias.n404 gnd 0.009605f
C1649 commonsourceibias.n405 gnd 0.009605f
C1650 commonsourceibias.n406 gnd 0.009605f
C1651 commonsourceibias.n407 gnd 0.012358f
C1652 commonsourceibias.n408 gnd 0.071604f
C1653 commonsourceibias.n409 gnd 0.012648f
C1654 commonsourceibias.n410 gnd 0.012288f
C1655 commonsourceibias.n411 gnd 0.009605f
C1656 commonsourceibias.n412 gnd 0.009605f
C1657 commonsourceibias.n413 gnd 0.009605f
C1658 commonsourceibias.n414 gnd 0.009057f
C1659 commonsourceibias.n415 gnd 0.01341f
C1660 commonsourceibias.n416 gnd 0.071604f
C1661 commonsourceibias.n417 gnd 0.013406f
C1662 commonsourceibias.n418 gnd 0.009605f
C1663 commonsourceibias.n419 gnd 0.009605f
C1664 commonsourceibias.n420 gnd 0.009605f
C1665 commonsourceibias.n421 gnd 0.012174f
C1666 commonsourceibias.n422 gnd 0.071604f
C1667 commonsourceibias.n423 gnd 0.012558f
C1668 commonsourceibias.n424 gnd 0.012378f
C1669 commonsourceibias.n425 gnd 0.009605f
C1670 commonsourceibias.n426 gnd 0.009605f
C1671 commonsourceibias.n427 gnd 0.009605f
C1672 commonsourceibias.n428 gnd 0.008798f
C1673 commonsourceibias.n429 gnd 0.013415f
C1674 commonsourceibias.n430 gnd 0.071604f
C1675 commonsourceibias.n431 gnd 0.013414f
C1676 commonsourceibias.n432 gnd 0.009605f
C1677 commonsourceibias.n433 gnd 0.009605f
C1678 commonsourceibias.n434 gnd 0.009605f
C1679 commonsourceibias.n435 gnd 0.01197f
C1680 commonsourceibias.n436 gnd 0.071604f
C1681 commonsourceibias.n437 gnd 0.012468f
C1682 commonsourceibias.n438 gnd 0.012468f
C1683 commonsourceibias.n439 gnd 0.009605f
C1684 commonsourceibias.n440 gnd 0.009605f
C1685 commonsourceibias.n441 gnd 0.009605f
C1686 commonsourceibias.n442 gnd 0.008571f
C1687 commonsourceibias.n443 gnd 0.013414f
C1688 commonsourceibias.n444 gnd 0.071604f
C1689 commonsourceibias.n445 gnd 0.013415f
C1690 commonsourceibias.n446 gnd 0.009605f
C1691 commonsourceibias.n447 gnd 0.009605f
C1692 commonsourceibias.n448 gnd 0.009605f
C1693 commonsourceibias.n449 gnd 0.011742f
C1694 commonsourceibias.n450 gnd 0.071604f
C1695 commonsourceibias.n451 gnd 0.012378f
C1696 commonsourceibias.n452 gnd 0.012558f
C1697 commonsourceibias.n453 gnd 0.009605f
C1698 commonsourceibias.n454 gnd 0.009605f
C1699 commonsourceibias.n455 gnd 0.009605f
C1700 commonsourceibias.n456 gnd 0.008375f
C1701 commonsourceibias.n457 gnd 0.013406f
C1702 commonsourceibias.n458 gnd 0.071604f
C1703 commonsourceibias.n459 gnd 0.01341f
C1704 commonsourceibias.n460 gnd 0.009605f
C1705 commonsourceibias.n461 gnd 0.009605f
C1706 commonsourceibias.n462 gnd 0.009605f
C1707 commonsourceibias.n463 gnd 0.011489f
C1708 commonsourceibias.n464 gnd 0.071604f
C1709 commonsourceibias.n465 gnd 0.012288f
C1710 commonsourceibias.n466 gnd 0.012648f
C1711 commonsourceibias.n467 gnd 0.009605f
C1712 commonsourceibias.n468 gnd 0.009605f
C1713 commonsourceibias.n469 gnd 0.009605f
C1714 commonsourceibias.n470 gnd 0.008208f
C1715 commonsourceibias.n471 gnd 0.013389f
C1716 commonsourceibias.n472 gnd 0.071604f
C1717 commonsourceibias.n473 gnd 0.013398f
C1718 commonsourceibias.n474 gnd 0.009605f
C1719 commonsourceibias.n475 gnd 0.009605f
C1720 commonsourceibias.n476 gnd 0.009605f
C1721 commonsourceibias.n477 gnd 0.011208f
C1722 commonsourceibias.n478 gnd 0.071604f
C1723 commonsourceibias.n479 gnd 0.011785f
C1724 commonsourceibias.t183 gnd 0.194086f
C1725 commonsourceibias.n480 gnd 0.085919f
C1726 commonsourceibias.n481 gnd 0.029883f
C1727 commonsourceibias.n482 gnd 0.456424f
C1728 commonsourceibias.n483 gnd 0.012817f
C1729 commonsourceibias.t112 gnd 0.194086f
C1730 commonsourceibias.t169 gnd 0.17946f
C1731 commonsourceibias.n484 gnd 0.009349f
C1732 commonsourceibias.n485 gnd 0.009605f
C1733 commonsourceibias.t142 gnd 0.17946f
C1734 commonsourceibias.n486 gnd 0.012358f
C1735 commonsourceibias.n487 gnd 0.009605f
C1736 commonsourceibias.t154 gnd 0.17946f
C1737 commonsourceibias.n488 gnd 0.009057f
C1738 commonsourceibias.n489 gnd 0.009605f
C1739 commonsourceibias.t108 gnd 0.17946f
C1740 commonsourceibias.n490 gnd 0.012174f
C1741 commonsourceibias.n491 gnd 0.009605f
C1742 commonsourceibias.t128 gnd 0.17946f
C1743 commonsourceibias.n492 gnd 0.008798f
C1744 commonsourceibias.n493 gnd 0.009605f
C1745 commonsourceibias.t109 gnd 0.17946f
C1746 commonsourceibias.n494 gnd 0.01197f
C1747 commonsourceibias.t69 gnd 0.020728f
C1748 commonsourceibias.t9 gnd 0.020728f
C1749 commonsourceibias.n495 gnd 0.18377f
C1750 commonsourceibias.t7 gnd 0.020728f
C1751 commonsourceibias.t67 gnd 0.020728f
C1752 commonsourceibias.n496 gnd 0.183157f
C1753 commonsourceibias.n497 gnd 0.170668f
C1754 commonsourceibias.t29 gnd 0.020728f
C1755 commonsourceibias.t79 gnd 0.020728f
C1756 commonsourceibias.n498 gnd 0.183157f
C1757 commonsourceibias.n499 gnd 0.084131f
C1758 commonsourceibias.t49 gnd 0.020728f
C1759 commonsourceibias.t3 gnd 0.020728f
C1760 commonsourceibias.n500 gnd 0.183157f
C1761 commonsourceibias.n501 gnd 0.084131f
C1762 commonsourceibias.t65 gnd 0.020728f
C1763 commonsourceibias.t51 gnd 0.020728f
C1764 commonsourceibias.n502 gnd 0.183157f
C1765 commonsourceibias.n503 gnd 0.070287f
C1766 commonsourceibias.n504 gnd 0.012817f
C1767 commonsourceibias.t76 gnd 0.17946f
C1768 commonsourceibias.n505 gnd 0.009349f
C1769 commonsourceibias.n506 gnd 0.009605f
C1770 commonsourceibias.t24 gnd 0.17946f
C1771 commonsourceibias.n507 gnd 0.012358f
C1772 commonsourceibias.n508 gnd 0.009605f
C1773 commonsourceibias.t12 gnd 0.17946f
C1774 commonsourceibias.n509 gnd 0.009057f
C1775 commonsourceibias.n510 gnd 0.009605f
C1776 commonsourceibias.t46 gnd 0.17946f
C1777 commonsourceibias.n511 gnd 0.012174f
C1778 commonsourceibias.n512 gnd 0.009605f
C1779 commonsourceibias.t32 gnd 0.17946f
C1780 commonsourceibias.n513 gnd 0.008798f
C1781 commonsourceibias.n514 gnd 0.009605f
C1782 commonsourceibias.t44 gnd 0.17946f
C1783 commonsourceibias.n515 gnd 0.01197f
C1784 commonsourceibias.n516 gnd 0.009605f
C1785 commonsourceibias.t50 gnd 0.17946f
C1786 commonsourceibias.n517 gnd 0.008571f
C1787 commonsourceibias.n518 gnd 0.009605f
C1788 commonsourceibias.t64 gnd 0.17946f
C1789 commonsourceibias.n519 gnd 0.011742f
C1790 commonsourceibias.n520 gnd 0.009605f
C1791 commonsourceibias.t48 gnd 0.17946f
C1792 commonsourceibias.n521 gnd 0.008375f
C1793 commonsourceibias.n522 gnd 0.009605f
C1794 commonsourceibias.t78 gnd 0.17946f
C1795 commonsourceibias.n523 gnd 0.011489f
C1796 commonsourceibias.n524 gnd 0.009605f
C1797 commonsourceibias.t66 gnd 0.17946f
C1798 commonsourceibias.n525 gnd 0.008208f
C1799 commonsourceibias.n526 gnd 0.009605f
C1800 commonsourceibias.t6 gnd 0.17946f
C1801 commonsourceibias.n527 gnd 0.011208f
C1802 commonsourceibias.t68 gnd 0.199526f
C1803 commonsourceibias.t8 gnd 0.17946f
C1804 commonsourceibias.n528 gnd 0.078221f
C1805 commonsourceibias.n529 gnd 0.085838f
C1806 commonsourceibias.n530 gnd 0.03983f
C1807 commonsourceibias.n531 gnd 0.009605f
C1808 commonsourceibias.n532 gnd 0.009349f
C1809 commonsourceibias.n533 gnd 0.013398f
C1810 commonsourceibias.n534 gnd 0.071604f
C1811 commonsourceibias.n535 gnd 0.013389f
C1812 commonsourceibias.n536 gnd 0.009605f
C1813 commonsourceibias.n537 gnd 0.009605f
C1814 commonsourceibias.n538 gnd 0.009605f
C1815 commonsourceibias.n539 gnd 0.012358f
C1816 commonsourceibias.n540 gnd 0.071604f
C1817 commonsourceibias.n541 gnd 0.012648f
C1818 commonsourceibias.t28 gnd 0.17946f
C1819 commonsourceibias.n542 gnd 0.071604f
C1820 commonsourceibias.n543 gnd 0.012288f
C1821 commonsourceibias.n544 gnd 0.009605f
C1822 commonsourceibias.n545 gnd 0.009605f
C1823 commonsourceibias.n546 gnd 0.009605f
C1824 commonsourceibias.n547 gnd 0.009057f
C1825 commonsourceibias.n548 gnd 0.01341f
C1826 commonsourceibias.n549 gnd 0.071604f
C1827 commonsourceibias.n550 gnd 0.013406f
C1828 commonsourceibias.n551 gnd 0.009605f
C1829 commonsourceibias.n552 gnd 0.009605f
C1830 commonsourceibias.n553 gnd 0.009605f
C1831 commonsourceibias.n554 gnd 0.012174f
C1832 commonsourceibias.n555 gnd 0.071604f
C1833 commonsourceibias.n556 gnd 0.012558f
C1834 commonsourceibias.t2 gnd 0.17946f
C1835 commonsourceibias.n557 gnd 0.071604f
C1836 commonsourceibias.n558 gnd 0.012378f
C1837 commonsourceibias.n559 gnd 0.009605f
C1838 commonsourceibias.n560 gnd 0.009605f
C1839 commonsourceibias.n561 gnd 0.009605f
C1840 commonsourceibias.n562 gnd 0.008798f
C1841 commonsourceibias.n563 gnd 0.013415f
C1842 commonsourceibias.n564 gnd 0.071604f
C1843 commonsourceibias.n565 gnd 0.013414f
C1844 commonsourceibias.n566 gnd 0.009605f
C1845 commonsourceibias.n567 gnd 0.009605f
C1846 commonsourceibias.n568 gnd 0.009605f
C1847 commonsourceibias.n569 gnd 0.01197f
C1848 commonsourceibias.n570 gnd 0.071604f
C1849 commonsourceibias.n571 gnd 0.012468f
C1850 commonsourceibias.t72 gnd 0.17946f
C1851 commonsourceibias.n572 gnd 0.071604f
C1852 commonsourceibias.n573 gnd 0.012468f
C1853 commonsourceibias.n574 gnd 0.009605f
C1854 commonsourceibias.n575 gnd 0.009605f
C1855 commonsourceibias.n576 gnd 0.009605f
C1856 commonsourceibias.n577 gnd 0.008571f
C1857 commonsourceibias.n578 gnd 0.013414f
C1858 commonsourceibias.n579 gnd 0.071604f
C1859 commonsourceibias.n580 gnd 0.013415f
C1860 commonsourceibias.n581 gnd 0.009605f
C1861 commonsourceibias.n582 gnd 0.009605f
C1862 commonsourceibias.n583 gnd 0.009605f
C1863 commonsourceibias.n584 gnd 0.011742f
C1864 commonsourceibias.n585 gnd 0.071604f
C1865 commonsourceibias.n586 gnd 0.012378f
C1866 commonsourceibias.t56 gnd 0.17946f
C1867 commonsourceibias.n587 gnd 0.071604f
C1868 commonsourceibias.n588 gnd 0.012558f
C1869 commonsourceibias.n589 gnd 0.009605f
C1870 commonsourceibias.n590 gnd 0.009605f
C1871 commonsourceibias.n591 gnd 0.009605f
C1872 commonsourceibias.n592 gnd 0.008375f
C1873 commonsourceibias.n593 gnd 0.013406f
C1874 commonsourceibias.n594 gnd 0.071604f
C1875 commonsourceibias.n595 gnd 0.01341f
C1876 commonsourceibias.n596 gnd 0.009605f
C1877 commonsourceibias.n597 gnd 0.009605f
C1878 commonsourceibias.n598 gnd 0.009605f
C1879 commonsourceibias.n599 gnd 0.011489f
C1880 commonsourceibias.n600 gnd 0.071604f
C1881 commonsourceibias.n601 gnd 0.012288f
C1882 commonsourceibias.t38 gnd 0.17946f
C1883 commonsourceibias.n602 gnd 0.071604f
C1884 commonsourceibias.n603 gnd 0.012648f
C1885 commonsourceibias.n604 gnd 0.009605f
C1886 commonsourceibias.n605 gnd 0.009605f
C1887 commonsourceibias.n606 gnd 0.009605f
C1888 commonsourceibias.n607 gnd 0.008208f
C1889 commonsourceibias.n608 gnd 0.013389f
C1890 commonsourceibias.n609 gnd 0.071604f
C1891 commonsourceibias.n610 gnd 0.013398f
C1892 commonsourceibias.n611 gnd 0.009605f
C1893 commonsourceibias.n612 gnd 0.009605f
C1894 commonsourceibias.n613 gnd 0.009605f
C1895 commonsourceibias.n614 gnd 0.011208f
C1896 commonsourceibias.n615 gnd 0.071604f
C1897 commonsourceibias.n616 gnd 0.011785f
C1898 commonsourceibias.t40 gnd 0.194086f
C1899 commonsourceibias.n617 gnd 0.085919f
C1900 commonsourceibias.n618 gnd 0.095702f
C1901 commonsourceibias.t77 gnd 0.020728f
C1902 commonsourceibias.t41 gnd 0.020728f
C1903 commonsourceibias.n619 gnd 0.183157f
C1904 commonsourceibias.n620 gnd 0.158432f
C1905 commonsourceibias.t39 gnd 0.020728f
C1906 commonsourceibias.t25 gnd 0.020728f
C1907 commonsourceibias.n621 gnd 0.183157f
C1908 commonsourceibias.n622 gnd 0.084131f
C1909 commonsourceibias.t47 gnd 0.020728f
C1910 commonsourceibias.t13 gnd 0.020728f
C1911 commonsourceibias.n623 gnd 0.183157f
C1912 commonsourceibias.n624 gnd 0.084131f
C1913 commonsourceibias.t33 gnd 0.020728f
C1914 commonsourceibias.t57 gnd 0.020728f
C1915 commonsourceibias.n625 gnd 0.183157f
C1916 commonsourceibias.n626 gnd 0.084131f
C1917 commonsourceibias.t73 gnd 0.020728f
C1918 commonsourceibias.t45 gnd 0.020728f
C1919 commonsourceibias.n627 gnd 0.183157f
C1920 commonsourceibias.n628 gnd 0.070287f
C1921 commonsourceibias.n629 gnd 0.085111f
C1922 commonsourceibias.n630 gnd 0.062167f
C1923 commonsourceibias.t102 gnd 0.17946f
C1924 commonsourceibias.n631 gnd 0.071604f
C1925 commonsourceibias.n632 gnd 0.009605f
C1926 commonsourceibias.t188 gnd 0.17946f
C1927 commonsourceibias.n633 gnd 0.071604f
C1928 commonsourceibias.n634 gnd 0.009605f
C1929 commonsourceibias.t162 gnd 0.17946f
C1930 commonsourceibias.n635 gnd 0.071604f
C1931 commonsourceibias.n636 gnd 0.009605f
C1932 commonsourceibias.t103 gnd 0.17946f
C1933 commonsourceibias.n637 gnd 0.008375f
C1934 commonsourceibias.n638 gnd 0.009605f
C1935 commonsourceibias.t166 gnd 0.17946f
C1936 commonsourceibias.n639 gnd 0.011489f
C1937 commonsourceibias.n640 gnd 0.009605f
C1938 commonsourceibias.t185 gnd 0.17946f
C1939 commonsourceibias.n641 gnd 0.008208f
C1940 commonsourceibias.n642 gnd 0.009605f
C1941 commonsourceibias.t160 gnd 0.17946f
C1942 commonsourceibias.n643 gnd 0.011208f
C1943 commonsourceibias.t177 gnd 0.199526f
C1944 commonsourceibias.t159 gnd 0.17946f
C1945 commonsourceibias.n644 gnd 0.078221f
C1946 commonsourceibias.n645 gnd 0.085838f
C1947 commonsourceibias.n646 gnd 0.03983f
C1948 commonsourceibias.n647 gnd 0.009605f
C1949 commonsourceibias.n648 gnd 0.009349f
C1950 commonsourceibias.n649 gnd 0.013398f
C1951 commonsourceibias.n650 gnd 0.071604f
C1952 commonsourceibias.n651 gnd 0.013389f
C1953 commonsourceibias.n652 gnd 0.009605f
C1954 commonsourceibias.n653 gnd 0.009605f
C1955 commonsourceibias.n654 gnd 0.009605f
C1956 commonsourceibias.n655 gnd 0.012358f
C1957 commonsourceibias.n656 gnd 0.071604f
C1958 commonsourceibias.n657 gnd 0.012648f
C1959 commonsourceibias.t135 gnd 0.17946f
C1960 commonsourceibias.n658 gnd 0.071604f
C1961 commonsourceibias.n659 gnd 0.012288f
C1962 commonsourceibias.n660 gnd 0.009605f
C1963 commonsourceibias.n661 gnd 0.009605f
C1964 commonsourceibias.n662 gnd 0.009605f
C1965 commonsourceibias.n663 gnd 0.009057f
C1966 commonsourceibias.n664 gnd 0.01341f
C1967 commonsourceibias.n665 gnd 0.071604f
C1968 commonsourceibias.n666 gnd 0.013406f
C1969 commonsourceibias.n667 gnd 0.009605f
C1970 commonsourceibias.n668 gnd 0.009605f
C1971 commonsourceibias.n669 gnd 0.009605f
C1972 commonsourceibias.n670 gnd 0.012174f
C1973 commonsourceibias.n671 gnd 0.071604f
C1974 commonsourceibias.n672 gnd 0.012558f
C1975 commonsourceibias.n673 gnd 0.012378f
C1976 commonsourceibias.n674 gnd 0.009605f
C1977 commonsourceibias.n675 gnd 0.009605f
C1978 commonsourceibias.n676 gnd 0.011742f
C1979 commonsourceibias.n677 gnd 0.008798f
C1980 commonsourceibias.n678 gnd 0.013415f
C1981 commonsourceibias.n679 gnd 0.009605f
C1982 commonsourceibias.n680 gnd 0.009605f
C1983 commonsourceibias.n681 gnd 0.013414f
C1984 commonsourceibias.n682 gnd 0.008571f
C1985 commonsourceibias.n683 gnd 0.01197f
C1986 commonsourceibias.n684 gnd 0.009605f
C1987 commonsourceibias.n685 gnd 0.008391f
C1988 commonsourceibias.n686 gnd 0.012468f
C1989 commonsourceibias.t174 gnd 0.17946f
C1990 commonsourceibias.n687 gnd 0.071604f
C1991 commonsourceibias.n688 gnd 0.012468f
C1992 commonsourceibias.n689 gnd 0.008391f
C1993 commonsourceibias.n690 gnd 0.009605f
C1994 commonsourceibias.n691 gnd 0.009605f
C1995 commonsourceibias.n692 gnd 0.008571f
C1996 commonsourceibias.n693 gnd 0.013414f
C1997 commonsourceibias.n694 gnd 0.071604f
C1998 commonsourceibias.n695 gnd 0.013415f
C1999 commonsourceibias.n696 gnd 0.009605f
C2000 commonsourceibias.n697 gnd 0.009605f
C2001 commonsourceibias.n698 gnd 0.009605f
C2002 commonsourceibias.n699 gnd 0.011742f
C2003 commonsourceibias.n700 gnd 0.071604f
C2004 commonsourceibias.n701 gnd 0.012378f
C2005 commonsourceibias.t90 gnd 0.17946f
C2006 commonsourceibias.n702 gnd 0.071604f
C2007 commonsourceibias.n703 gnd 0.012558f
C2008 commonsourceibias.n704 gnd 0.009605f
C2009 commonsourceibias.n705 gnd 0.009605f
C2010 commonsourceibias.n706 gnd 0.009605f
C2011 commonsourceibias.n707 gnd 0.008375f
C2012 commonsourceibias.n708 gnd 0.013406f
C2013 commonsourceibias.n709 gnd 0.071604f
C2014 commonsourceibias.n710 gnd 0.01341f
C2015 commonsourceibias.n711 gnd 0.009605f
C2016 commonsourceibias.n712 gnd 0.009605f
C2017 commonsourceibias.n713 gnd 0.009605f
C2018 commonsourceibias.n714 gnd 0.011489f
C2019 commonsourceibias.n715 gnd 0.071604f
C2020 commonsourceibias.n716 gnd 0.012288f
C2021 commonsourceibias.t116 gnd 0.17946f
C2022 commonsourceibias.n717 gnd 0.071604f
C2023 commonsourceibias.n718 gnd 0.012648f
C2024 commonsourceibias.n719 gnd 0.009605f
C2025 commonsourceibias.n720 gnd 0.009605f
C2026 commonsourceibias.n721 gnd 0.009605f
C2027 commonsourceibias.n722 gnd 0.008208f
C2028 commonsourceibias.n723 gnd 0.013389f
C2029 commonsourceibias.n724 gnd 0.071604f
C2030 commonsourceibias.n725 gnd 0.013398f
C2031 commonsourceibias.n726 gnd 0.009605f
C2032 commonsourceibias.n727 gnd 0.009605f
C2033 commonsourceibias.n728 gnd 0.009605f
C2034 commonsourceibias.n729 gnd 0.011208f
C2035 commonsourceibias.n730 gnd 0.071604f
C2036 commonsourceibias.n731 gnd 0.011785f
C2037 commonsourceibias.n732 gnd 0.085919f
C2038 commonsourceibias.n733 gnd 0.056156f
C2039 commonsourceibias.n734 gnd 0.012817f
C2040 commonsourceibias.t180 gnd 0.17946f
C2041 commonsourceibias.n735 gnd 0.009349f
C2042 commonsourceibias.n736 gnd 0.009605f
C2043 commonsourceibias.t82 gnd 0.17946f
C2044 commonsourceibias.n737 gnd 0.012358f
C2045 commonsourceibias.n738 gnd 0.009605f
C2046 commonsourceibias.t179 gnd 0.17946f
C2047 commonsourceibias.n739 gnd 0.009057f
C2048 commonsourceibias.n740 gnd 0.009605f
C2049 commonsourceibias.t81 gnd 0.17946f
C2050 commonsourceibias.n741 gnd 0.012174f
C2051 commonsourceibias.n742 gnd 0.009605f
C2052 commonsourceibias.t178 gnd 0.17946f
C2053 commonsourceibias.n743 gnd 0.008798f
C2054 commonsourceibias.n744 gnd 0.009605f
C2055 commonsourceibias.t89 gnd 0.17946f
C2056 commonsourceibias.n745 gnd 0.01197f
C2057 commonsourceibias.n746 gnd 0.009605f
C2058 commonsourceibias.t97 gnd 0.17946f
C2059 commonsourceibias.n747 gnd 0.008571f
C2060 commonsourceibias.n748 gnd 0.009605f
C2061 commonsourceibias.t86 gnd 0.17946f
C2062 commonsourceibias.n749 gnd 0.011742f
C2063 commonsourceibias.n750 gnd 0.009605f
C2064 commonsourceibias.t106 gnd 0.17946f
C2065 commonsourceibias.n751 gnd 0.008375f
C2066 commonsourceibias.n752 gnd 0.009605f
C2067 commonsourceibias.t85 gnd 0.17946f
C2068 commonsourceibias.n753 gnd 0.011489f
C2069 commonsourceibias.n754 gnd 0.009605f
C2070 commonsourceibias.t104 gnd 0.17946f
C2071 commonsourceibias.n755 gnd 0.008208f
C2072 commonsourceibias.n756 gnd 0.009605f
C2073 commonsourceibias.t132 gnd 0.17946f
C2074 commonsourceibias.n757 gnd 0.011208f
C2075 commonsourceibias.t98 gnd 0.199526f
C2076 commonsourceibias.t123 gnd 0.17946f
C2077 commonsourceibias.n758 gnd 0.078221f
C2078 commonsourceibias.n759 gnd 0.085838f
C2079 commonsourceibias.n760 gnd 0.03983f
C2080 commonsourceibias.n761 gnd 0.009605f
C2081 commonsourceibias.n762 gnd 0.009349f
C2082 commonsourceibias.n763 gnd 0.013398f
C2083 commonsourceibias.n764 gnd 0.071604f
C2084 commonsourceibias.n765 gnd 0.013389f
C2085 commonsourceibias.n766 gnd 0.009605f
C2086 commonsourceibias.n767 gnd 0.009605f
C2087 commonsourceibias.n768 gnd 0.009605f
C2088 commonsourceibias.n769 gnd 0.012358f
C2089 commonsourceibias.n770 gnd 0.071604f
C2090 commonsourceibias.n771 gnd 0.012648f
C2091 commonsourceibias.t118 gnd 0.17946f
C2092 commonsourceibias.n772 gnd 0.071604f
C2093 commonsourceibias.n773 gnd 0.012288f
C2094 commonsourceibias.n774 gnd 0.009605f
C2095 commonsourceibias.n775 gnd 0.009605f
C2096 commonsourceibias.n776 gnd 0.009605f
C2097 commonsourceibias.n777 gnd 0.009057f
C2098 commonsourceibias.n778 gnd 0.01341f
C2099 commonsourceibias.n779 gnd 0.071604f
C2100 commonsourceibias.n780 gnd 0.013406f
C2101 commonsourceibias.n781 gnd 0.009605f
C2102 commonsourceibias.n782 gnd 0.009605f
C2103 commonsourceibias.n783 gnd 0.009605f
C2104 commonsourceibias.n784 gnd 0.012174f
C2105 commonsourceibias.n785 gnd 0.071604f
C2106 commonsourceibias.n786 gnd 0.012558f
C2107 commonsourceibias.t119 gnd 0.17946f
C2108 commonsourceibias.n787 gnd 0.071604f
C2109 commonsourceibias.n788 gnd 0.012378f
C2110 commonsourceibias.n789 gnd 0.009605f
C2111 commonsourceibias.n790 gnd 0.009605f
C2112 commonsourceibias.n791 gnd 0.009605f
C2113 commonsourceibias.n792 gnd 0.008798f
C2114 commonsourceibias.n793 gnd 0.013415f
C2115 commonsourceibias.n794 gnd 0.071604f
C2116 commonsourceibias.n795 gnd 0.013414f
C2117 commonsourceibias.n796 gnd 0.009605f
C2118 commonsourceibias.n797 gnd 0.009605f
C2119 commonsourceibias.n798 gnd 0.009605f
C2120 commonsourceibias.n799 gnd 0.01197f
C2121 commonsourceibias.n800 gnd 0.071604f
C2122 commonsourceibias.n801 gnd 0.012468f
C2123 commonsourceibias.t120 gnd 0.17946f
C2124 commonsourceibias.n802 gnd 0.071604f
C2125 commonsourceibias.n803 gnd 0.012468f
C2126 commonsourceibias.n804 gnd 0.009605f
C2127 commonsourceibias.n805 gnd 0.009605f
C2128 commonsourceibias.n806 gnd 0.009605f
C2129 commonsourceibias.n807 gnd 0.008571f
C2130 commonsourceibias.n808 gnd 0.013414f
C2131 commonsourceibias.n809 gnd 0.071604f
C2132 commonsourceibias.n810 gnd 0.013415f
C2133 commonsourceibias.n811 gnd 0.009605f
C2134 commonsourceibias.n812 gnd 0.009605f
C2135 commonsourceibias.n813 gnd 0.009605f
C2136 commonsourceibias.n814 gnd 0.011742f
C2137 commonsourceibias.n815 gnd 0.071604f
C2138 commonsourceibias.n816 gnd 0.012378f
C2139 commonsourceibias.t121 gnd 0.17946f
C2140 commonsourceibias.n817 gnd 0.071604f
C2141 commonsourceibias.n818 gnd 0.012558f
C2142 commonsourceibias.n819 gnd 0.009605f
C2143 commonsourceibias.n820 gnd 0.009605f
C2144 commonsourceibias.n821 gnd 0.009605f
C2145 commonsourceibias.n822 gnd 0.008375f
C2146 commonsourceibias.n823 gnd 0.013406f
C2147 commonsourceibias.n824 gnd 0.071604f
C2148 commonsourceibias.n825 gnd 0.01341f
C2149 commonsourceibias.n826 gnd 0.009605f
C2150 commonsourceibias.n827 gnd 0.009605f
C2151 commonsourceibias.n828 gnd 0.009605f
C2152 commonsourceibias.n829 gnd 0.011489f
C2153 commonsourceibias.n830 gnd 0.071604f
C2154 commonsourceibias.n831 gnd 0.012288f
C2155 commonsourceibias.t193 gnd 0.17946f
C2156 commonsourceibias.n832 gnd 0.071604f
C2157 commonsourceibias.n833 gnd 0.012648f
C2158 commonsourceibias.n834 gnd 0.009605f
C2159 commonsourceibias.n835 gnd 0.009605f
C2160 commonsourceibias.n836 gnd 0.009605f
C2161 commonsourceibias.n837 gnd 0.008208f
C2162 commonsourceibias.n838 gnd 0.013389f
C2163 commonsourceibias.n839 gnd 0.071604f
C2164 commonsourceibias.n840 gnd 0.013398f
C2165 commonsourceibias.n841 gnd 0.009605f
C2166 commonsourceibias.n842 gnd 0.009605f
C2167 commonsourceibias.n843 gnd 0.009605f
C2168 commonsourceibias.n844 gnd 0.011208f
C2169 commonsourceibias.n845 gnd 0.071604f
C2170 commonsourceibias.n846 gnd 0.011785f
C2171 commonsourceibias.t189 gnd 0.194086f
C2172 commonsourceibias.n847 gnd 0.085919f
C2173 commonsourceibias.n848 gnd 0.029883f
C2174 commonsourceibias.n849 gnd 0.153509f
C2175 commonsourceibias.n850 gnd 0.012817f
C2176 commonsourceibias.t133 gnd 0.17946f
C2177 commonsourceibias.n851 gnd 0.009349f
C2178 commonsourceibias.n852 gnd 0.009605f
C2179 commonsourceibias.t153 gnd 0.17946f
C2180 commonsourceibias.n853 gnd 0.012358f
C2181 commonsourceibias.n854 gnd 0.009605f
C2182 commonsourceibias.t122 gnd 0.17946f
C2183 commonsourceibias.n855 gnd 0.009057f
C2184 commonsourceibias.n856 gnd 0.009605f
C2185 commonsourceibias.t143 gnd 0.17946f
C2186 commonsourceibias.n857 gnd 0.012174f
C2187 commonsourceibias.n858 gnd 0.009605f
C2188 commonsourceibias.t99 gnd 0.17946f
C2189 commonsourceibias.n859 gnd 0.008798f
C2190 commonsourceibias.n860 gnd 0.009605f
C2191 commonsourceibias.t87 gnd 0.17946f
C2192 commonsourceibias.n861 gnd 0.01197f
C2193 commonsourceibias.n862 gnd 0.009605f
C2194 commonsourceibias.t167 gnd 0.17946f
C2195 commonsourceibias.n863 gnd 0.008571f
C2196 commonsourceibias.n864 gnd 0.009605f
C2197 commonsourceibias.t192 gnd 0.17946f
C2198 commonsourceibias.n865 gnd 0.011742f
C2199 commonsourceibias.n866 gnd 0.009605f
C2200 commonsourceibias.t136 gnd 0.17946f
C2201 commonsourceibias.n867 gnd 0.008375f
C2202 commonsourceibias.n868 gnd 0.009605f
C2203 commonsourceibias.t181 gnd 0.17946f
C2204 commonsourceibias.n869 gnd 0.011489f
C2205 commonsourceibias.n870 gnd 0.009605f
C2206 commonsourceibias.t126 gnd 0.17946f
C2207 commonsourceibias.n871 gnd 0.008208f
C2208 commonsourceibias.n872 gnd 0.009605f
C2209 commonsourceibias.t146 gnd 0.17946f
C2210 commonsourceibias.n873 gnd 0.011208f
C2211 commonsourceibias.t191 gnd 0.199526f
C2212 commonsourceibias.t156 gnd 0.17946f
C2213 commonsourceibias.n874 gnd 0.078221f
C2214 commonsourceibias.n875 gnd 0.085838f
C2215 commonsourceibias.n876 gnd 0.03983f
C2216 commonsourceibias.n877 gnd 0.009605f
C2217 commonsourceibias.n878 gnd 0.009349f
C2218 commonsourceibias.n879 gnd 0.013398f
C2219 commonsourceibias.n880 gnd 0.071604f
C2220 commonsourceibias.n881 gnd 0.013389f
C2221 commonsourceibias.n882 gnd 0.009605f
C2222 commonsourceibias.n883 gnd 0.009605f
C2223 commonsourceibias.n884 gnd 0.009605f
C2224 commonsourceibias.n885 gnd 0.012358f
C2225 commonsourceibias.n886 gnd 0.071604f
C2226 commonsourceibias.n887 gnd 0.012648f
C2227 commonsourceibias.t91 gnd 0.17946f
C2228 commonsourceibias.n888 gnd 0.071604f
C2229 commonsourceibias.n889 gnd 0.012288f
C2230 commonsourceibias.n890 gnd 0.009605f
C2231 commonsourceibias.n891 gnd 0.009605f
C2232 commonsourceibias.n892 gnd 0.009605f
C2233 commonsourceibias.n893 gnd 0.009057f
C2234 commonsourceibias.n894 gnd 0.01341f
C2235 commonsourceibias.n895 gnd 0.071604f
C2236 commonsourceibias.n896 gnd 0.013406f
C2237 commonsourceibias.n897 gnd 0.009605f
C2238 commonsourceibias.n898 gnd 0.009605f
C2239 commonsourceibias.n899 gnd 0.009605f
C2240 commonsourceibias.n900 gnd 0.012174f
C2241 commonsourceibias.n901 gnd 0.071604f
C2242 commonsourceibias.n902 gnd 0.012558f
C2243 commonsourceibias.t107 gnd 0.17946f
C2244 commonsourceibias.n903 gnd 0.071604f
C2245 commonsourceibias.n904 gnd 0.012378f
C2246 commonsourceibias.n905 gnd 0.009605f
C2247 commonsourceibias.n906 gnd 0.009605f
C2248 commonsourceibias.n907 gnd 0.009605f
C2249 commonsourceibias.n908 gnd 0.008798f
C2250 commonsourceibias.n909 gnd 0.013415f
C2251 commonsourceibias.n910 gnd 0.071604f
C2252 commonsourceibias.n911 gnd 0.013414f
C2253 commonsourceibias.n912 gnd 0.009605f
C2254 commonsourceibias.n913 gnd 0.009605f
C2255 commonsourceibias.n914 gnd 0.009605f
C2256 commonsourceibias.n915 gnd 0.01197f
C2257 commonsourceibias.n916 gnd 0.071604f
C2258 commonsourceibias.n917 gnd 0.012468f
C2259 commonsourceibias.t127 gnd 0.17946f
C2260 commonsourceibias.n918 gnd 0.071604f
C2261 commonsourceibias.n919 gnd 0.012468f
C2262 commonsourceibias.n920 gnd 0.009605f
C2263 commonsourceibias.n921 gnd 0.009605f
C2264 commonsourceibias.n922 gnd 0.009605f
C2265 commonsourceibias.n923 gnd 0.008571f
C2266 commonsourceibias.n924 gnd 0.013414f
C2267 commonsourceibias.n925 gnd 0.071604f
C2268 commonsourceibias.n926 gnd 0.013415f
C2269 commonsourceibias.n927 gnd 0.009605f
C2270 commonsourceibias.n928 gnd 0.009605f
C2271 commonsourceibias.n929 gnd 0.009605f
C2272 commonsourceibias.n930 gnd 0.011742f
C2273 commonsourceibias.n931 gnd 0.071604f
C2274 commonsourceibias.n932 gnd 0.012378f
C2275 commonsourceibias.t137 gnd 0.17946f
C2276 commonsourceibias.n933 gnd 0.071604f
C2277 commonsourceibias.n934 gnd 0.012558f
C2278 commonsourceibias.n935 gnd 0.009605f
C2279 commonsourceibias.n936 gnd 0.009605f
C2280 commonsourceibias.n937 gnd 0.009605f
C2281 commonsourceibias.n938 gnd 0.008375f
C2282 commonsourceibias.n939 gnd 0.013406f
C2283 commonsourceibias.n940 gnd 0.071604f
C2284 commonsourceibias.n941 gnd 0.01341f
C2285 commonsourceibias.n942 gnd 0.009605f
C2286 commonsourceibias.n943 gnd 0.009605f
C2287 commonsourceibias.n944 gnd 0.009605f
C2288 commonsourceibias.n945 gnd 0.011489f
C2289 commonsourceibias.n946 gnd 0.071604f
C2290 commonsourceibias.n947 gnd 0.012288f
C2291 commonsourceibias.t170 gnd 0.17946f
C2292 commonsourceibias.n948 gnd 0.071604f
C2293 commonsourceibias.n949 gnd 0.012648f
C2294 commonsourceibias.n950 gnd 0.009605f
C2295 commonsourceibias.n951 gnd 0.009605f
C2296 commonsourceibias.n952 gnd 0.009605f
C2297 commonsourceibias.n953 gnd 0.008208f
C2298 commonsourceibias.n954 gnd 0.013389f
C2299 commonsourceibias.n955 gnd 0.071604f
C2300 commonsourceibias.n956 gnd 0.013398f
C2301 commonsourceibias.n957 gnd 0.009605f
C2302 commonsourceibias.n958 gnd 0.009605f
C2303 commonsourceibias.n959 gnd 0.009605f
C2304 commonsourceibias.n960 gnd 0.011208f
C2305 commonsourceibias.n961 gnd 0.071604f
C2306 commonsourceibias.n962 gnd 0.011785f
C2307 commonsourceibias.t101 gnd 0.194086f
C2308 commonsourceibias.n963 gnd 0.085919f
C2309 commonsourceibias.n964 gnd 0.029883f
C2310 commonsourceibias.n965 gnd 0.202572f
C2311 commonsourceibias.n966 gnd 5.28148f
C2312 vdd.t46 gnd 0.034846f
C2313 vdd.t26 gnd 0.034846f
C2314 vdd.n0 gnd 0.274839f
C2315 vdd.t5 gnd 0.034846f
C2316 vdd.t42 gnd 0.034846f
C2317 vdd.n1 gnd 0.274385f
C2318 vdd.n2 gnd 0.253035f
C2319 vdd.t23 gnd 0.034846f
C2320 vdd.t53 gnd 0.034846f
C2321 vdd.n3 gnd 0.274385f
C2322 vdd.n4 gnd 0.127969f
C2323 vdd.t51 gnd 0.034846f
C2324 vdd.t31 gnd 0.034846f
C2325 vdd.n5 gnd 0.274385f
C2326 vdd.n6 gnd 0.120076f
C2327 vdd.t57 gnd 0.034846f
C2328 vdd.t21 gnd 0.034846f
C2329 vdd.n7 gnd 0.274839f
C2330 vdd.t29 gnd 0.034846f
C2331 vdd.t49 gnd 0.034846f
C2332 vdd.n8 gnd 0.274385f
C2333 vdd.n9 gnd 0.253035f
C2334 vdd.t38 gnd 0.034846f
C2335 vdd.t9 gnd 0.034846f
C2336 vdd.n10 gnd 0.274385f
C2337 vdd.n11 gnd 0.127969f
C2338 vdd.t18 gnd 0.034846f
C2339 vdd.t36 gnd 0.034846f
C2340 vdd.n12 gnd 0.274385f
C2341 vdd.n13 gnd 0.120076f
C2342 vdd.n14 gnd 0.084891f
C2343 vdd.t271 gnd 0.019359f
C2344 vdd.t272 gnd 0.019359f
C2345 vdd.n15 gnd 0.178192f
C2346 vdd.t62 gnd 0.019359f
C2347 vdd.t269 gnd 0.019359f
C2348 vdd.n16 gnd 0.177671f
C2349 vdd.n17 gnd 0.309202f
C2350 vdd.t0 gnd 0.019359f
C2351 vdd.t60 gnd 0.019359f
C2352 vdd.n18 gnd 0.177671f
C2353 vdd.n19 gnd 0.127921f
C2354 vdd.t63 gnd 0.019359f
C2355 vdd.t270 gnd 0.019359f
C2356 vdd.n20 gnd 0.178192f
C2357 vdd.t273 gnd 0.019359f
C2358 vdd.t59 gnd 0.019359f
C2359 vdd.n21 gnd 0.177671f
C2360 vdd.n22 gnd 0.309202f
C2361 vdd.t61 gnd 0.019359f
C2362 vdd.t274 gnd 0.019359f
C2363 vdd.n23 gnd 0.177671f
C2364 vdd.n24 gnd 0.127921f
C2365 vdd.t1 gnd 0.019359f
C2366 vdd.t58 gnd 0.019359f
C2367 vdd.n25 gnd 0.177671f
C2368 vdd.t275 gnd 0.019359f
C2369 vdd.t192 gnd 0.019359f
C2370 vdd.n26 gnd 0.177671f
C2371 vdd.n27 gnd 19.6921f
C2372 vdd.n28 gnd 7.906759f
C2373 vdd.n29 gnd 0.00528f
C2374 vdd.n30 gnd 0.0049f
C2375 vdd.n31 gnd 0.00271f
C2376 vdd.n32 gnd 0.006223f
C2377 vdd.n33 gnd 0.002633f
C2378 vdd.n34 gnd 0.002788f
C2379 vdd.n35 gnd 0.0049f
C2380 vdd.n36 gnd 0.002633f
C2381 vdd.n37 gnd 0.006223f
C2382 vdd.n38 gnd 0.002788f
C2383 vdd.n39 gnd 0.0049f
C2384 vdd.n40 gnd 0.002633f
C2385 vdd.n41 gnd 0.004667f
C2386 vdd.n42 gnd 0.004681f
C2387 vdd.t130 gnd 0.01337f
C2388 vdd.n43 gnd 0.029747f
C2389 vdd.n44 gnd 0.154813f
C2390 vdd.n45 gnd 0.002633f
C2391 vdd.n46 gnd 0.002788f
C2392 vdd.n47 gnd 0.006223f
C2393 vdd.n48 gnd 0.006223f
C2394 vdd.n49 gnd 0.002788f
C2395 vdd.n50 gnd 0.002633f
C2396 vdd.n51 gnd 0.0049f
C2397 vdd.n52 gnd 0.0049f
C2398 vdd.n53 gnd 0.002633f
C2399 vdd.n54 gnd 0.002788f
C2400 vdd.n55 gnd 0.006223f
C2401 vdd.n56 gnd 0.006223f
C2402 vdd.n57 gnd 0.002788f
C2403 vdd.n58 gnd 0.002633f
C2404 vdd.n59 gnd 0.0049f
C2405 vdd.n60 gnd 0.0049f
C2406 vdd.n61 gnd 0.002633f
C2407 vdd.n62 gnd 0.002788f
C2408 vdd.n63 gnd 0.006223f
C2409 vdd.n64 gnd 0.006223f
C2410 vdd.n65 gnd 0.014713f
C2411 vdd.n66 gnd 0.00271f
C2412 vdd.n67 gnd 0.002633f
C2413 vdd.n68 gnd 0.012664f
C2414 vdd.n69 gnd 0.008841f
C2415 vdd.t107 gnd 0.030974f
C2416 vdd.t171 gnd 0.030974f
C2417 vdd.n70 gnd 0.212878f
C2418 vdd.n71 gnd 0.167396f
C2419 vdd.t88 gnd 0.030974f
C2420 vdd.t155 gnd 0.030974f
C2421 vdd.n72 gnd 0.212878f
C2422 vdd.n73 gnd 0.135088f
C2423 vdd.t93 gnd 0.030974f
C2424 vdd.t167 gnd 0.030974f
C2425 vdd.n74 gnd 0.212878f
C2426 vdd.n75 gnd 0.135088f
C2427 vdd.t117 gnd 0.030974f
C2428 vdd.t180 gnd 0.030974f
C2429 vdd.n76 gnd 0.212878f
C2430 vdd.n77 gnd 0.135088f
C2431 vdd.t133 gnd 0.030974f
C2432 vdd.t161 gnd 0.030974f
C2433 vdd.n78 gnd 0.212878f
C2434 vdd.n79 gnd 0.135088f
C2435 vdd.t108 gnd 0.030974f
C2436 vdd.t173 gnd 0.030974f
C2437 vdd.n80 gnd 0.212878f
C2438 vdd.n81 gnd 0.135088f
C2439 vdd.t123 gnd 0.030974f
C2440 vdd.t187 gnd 0.030974f
C2441 vdd.n82 gnd 0.212878f
C2442 vdd.n83 gnd 0.135088f
C2443 vdd.n84 gnd 0.00528f
C2444 vdd.n85 gnd 0.0049f
C2445 vdd.n86 gnd 0.00271f
C2446 vdd.n87 gnd 0.006223f
C2447 vdd.n88 gnd 0.002633f
C2448 vdd.n89 gnd 0.002788f
C2449 vdd.n90 gnd 0.0049f
C2450 vdd.n91 gnd 0.002633f
C2451 vdd.n92 gnd 0.006223f
C2452 vdd.n93 gnd 0.002788f
C2453 vdd.n94 gnd 0.0049f
C2454 vdd.n95 gnd 0.002633f
C2455 vdd.n96 gnd 0.004667f
C2456 vdd.n97 gnd 0.004681f
C2457 vdd.t145 gnd 0.01337f
C2458 vdd.n98 gnd 0.029747f
C2459 vdd.n99 gnd 0.154813f
C2460 vdd.n100 gnd 0.002633f
C2461 vdd.n101 gnd 0.002788f
C2462 vdd.n102 gnd 0.006223f
C2463 vdd.n103 gnd 0.006223f
C2464 vdd.n104 gnd 0.002788f
C2465 vdd.n105 gnd 0.002633f
C2466 vdd.n106 gnd 0.0049f
C2467 vdd.n107 gnd 0.0049f
C2468 vdd.n108 gnd 0.002633f
C2469 vdd.n109 gnd 0.002788f
C2470 vdd.n110 gnd 0.006223f
C2471 vdd.n111 gnd 0.006223f
C2472 vdd.n112 gnd 0.002788f
C2473 vdd.n113 gnd 0.002633f
C2474 vdd.n114 gnd 0.0049f
C2475 vdd.n115 gnd 0.0049f
C2476 vdd.n116 gnd 0.002633f
C2477 vdd.n117 gnd 0.002788f
C2478 vdd.n118 gnd 0.006223f
C2479 vdd.n119 gnd 0.006223f
C2480 vdd.n120 gnd 0.014713f
C2481 vdd.n121 gnd 0.00271f
C2482 vdd.n122 gnd 0.002633f
C2483 vdd.n123 gnd 0.012664f
C2484 vdd.n124 gnd 0.008564f
C2485 vdd.n125 gnd 0.100506f
C2486 vdd.n126 gnd 0.00528f
C2487 vdd.n127 gnd 0.0049f
C2488 vdd.n128 gnd 0.00271f
C2489 vdd.n129 gnd 0.006223f
C2490 vdd.n130 gnd 0.002633f
C2491 vdd.n131 gnd 0.002788f
C2492 vdd.n132 gnd 0.0049f
C2493 vdd.n133 gnd 0.002633f
C2494 vdd.n134 gnd 0.006223f
C2495 vdd.n135 gnd 0.002788f
C2496 vdd.n136 gnd 0.0049f
C2497 vdd.n137 gnd 0.002633f
C2498 vdd.n138 gnd 0.004667f
C2499 vdd.n139 gnd 0.004681f
C2500 vdd.t175 gnd 0.01337f
C2501 vdd.n140 gnd 0.029747f
C2502 vdd.n141 gnd 0.154813f
C2503 vdd.n142 gnd 0.002633f
C2504 vdd.n143 gnd 0.002788f
C2505 vdd.n144 gnd 0.006223f
C2506 vdd.n145 gnd 0.006223f
C2507 vdd.n146 gnd 0.002788f
C2508 vdd.n147 gnd 0.002633f
C2509 vdd.n148 gnd 0.0049f
C2510 vdd.n149 gnd 0.0049f
C2511 vdd.n150 gnd 0.002633f
C2512 vdd.n151 gnd 0.002788f
C2513 vdd.n152 gnd 0.006223f
C2514 vdd.n153 gnd 0.006223f
C2515 vdd.n154 gnd 0.002788f
C2516 vdd.n155 gnd 0.002633f
C2517 vdd.n156 gnd 0.0049f
C2518 vdd.n157 gnd 0.0049f
C2519 vdd.n158 gnd 0.002633f
C2520 vdd.n159 gnd 0.002788f
C2521 vdd.n160 gnd 0.006223f
C2522 vdd.n161 gnd 0.006223f
C2523 vdd.n162 gnd 0.014713f
C2524 vdd.n163 gnd 0.00271f
C2525 vdd.n164 gnd 0.002633f
C2526 vdd.n165 gnd 0.012664f
C2527 vdd.n166 gnd 0.008841f
C2528 vdd.t178 gnd 0.030974f
C2529 vdd.t85 gnd 0.030974f
C2530 vdd.n167 gnd 0.212878f
C2531 vdd.n168 gnd 0.167396f
C2532 vdd.t163 gnd 0.030974f
C2533 vdd.t170 gnd 0.030974f
C2534 vdd.n169 gnd 0.212878f
C2535 vdd.n170 gnd 0.135088f
C2536 vdd.t71 gnd 0.030974f
C2537 vdd.t128 gnd 0.030974f
C2538 vdd.n171 gnd 0.212878f
C2539 vdd.n172 gnd 0.135088f
C2540 vdd.t160 gnd 0.030974f
C2541 vdd.t183 gnd 0.030974f
C2542 vdd.n173 gnd 0.212878f
C2543 vdd.n174 gnd 0.135088f
C2544 vdd.t113 gnd 0.030974f
C2545 vdd.t159 gnd 0.030974f
C2546 vdd.n175 gnd 0.212878f
C2547 vdd.n176 gnd 0.135088f
C2548 vdd.t190 gnd 0.030974f
C2549 vdd.t105 gnd 0.030974f
C2550 vdd.n177 gnd 0.212878f
C2551 vdd.n178 gnd 0.135088f
C2552 vdd.t144 gnd 0.030974f
C2553 vdd.t177 gnd 0.030974f
C2554 vdd.n179 gnd 0.212878f
C2555 vdd.n180 gnd 0.135088f
C2556 vdd.n181 gnd 0.00528f
C2557 vdd.n182 gnd 0.0049f
C2558 vdd.n183 gnd 0.00271f
C2559 vdd.n184 gnd 0.006223f
C2560 vdd.n185 gnd 0.002633f
C2561 vdd.n186 gnd 0.002788f
C2562 vdd.n187 gnd 0.0049f
C2563 vdd.n188 gnd 0.002633f
C2564 vdd.n189 gnd 0.006223f
C2565 vdd.n190 gnd 0.002788f
C2566 vdd.n191 gnd 0.0049f
C2567 vdd.n192 gnd 0.002633f
C2568 vdd.n193 gnd 0.004667f
C2569 vdd.n194 gnd 0.004681f
C2570 vdd.t81 gnd 0.01337f
C2571 vdd.n195 gnd 0.029747f
C2572 vdd.n196 gnd 0.154813f
C2573 vdd.n197 gnd 0.002633f
C2574 vdd.n198 gnd 0.002788f
C2575 vdd.n199 gnd 0.006223f
C2576 vdd.n200 gnd 0.006223f
C2577 vdd.n201 gnd 0.002788f
C2578 vdd.n202 gnd 0.002633f
C2579 vdd.n203 gnd 0.0049f
C2580 vdd.n204 gnd 0.0049f
C2581 vdd.n205 gnd 0.002633f
C2582 vdd.n206 gnd 0.002788f
C2583 vdd.n207 gnd 0.006223f
C2584 vdd.n208 gnd 0.006223f
C2585 vdd.n209 gnd 0.002788f
C2586 vdd.n210 gnd 0.002633f
C2587 vdd.n211 gnd 0.0049f
C2588 vdd.n212 gnd 0.0049f
C2589 vdd.n213 gnd 0.002633f
C2590 vdd.n214 gnd 0.002788f
C2591 vdd.n215 gnd 0.006223f
C2592 vdd.n216 gnd 0.006223f
C2593 vdd.n217 gnd 0.014713f
C2594 vdd.n218 gnd 0.00271f
C2595 vdd.n219 gnd 0.002633f
C2596 vdd.n220 gnd 0.012664f
C2597 vdd.n221 gnd 0.008564f
C2598 vdd.n222 gnd 0.059791f
C2599 vdd.n223 gnd 0.215442f
C2600 vdd.n224 gnd 0.00528f
C2601 vdd.n225 gnd 0.0049f
C2602 vdd.n226 gnd 0.00271f
C2603 vdd.n227 gnd 0.006223f
C2604 vdd.n228 gnd 0.002633f
C2605 vdd.n229 gnd 0.002788f
C2606 vdd.n230 gnd 0.0049f
C2607 vdd.n231 gnd 0.002633f
C2608 vdd.n232 gnd 0.006223f
C2609 vdd.n233 gnd 0.002788f
C2610 vdd.n234 gnd 0.0049f
C2611 vdd.n235 gnd 0.002633f
C2612 vdd.n236 gnd 0.004667f
C2613 vdd.n237 gnd 0.004681f
C2614 vdd.t185 gnd 0.01337f
C2615 vdd.n238 gnd 0.029747f
C2616 vdd.n239 gnd 0.154813f
C2617 vdd.n240 gnd 0.002633f
C2618 vdd.n241 gnd 0.002788f
C2619 vdd.n242 gnd 0.006223f
C2620 vdd.n243 gnd 0.006223f
C2621 vdd.n244 gnd 0.002788f
C2622 vdd.n245 gnd 0.002633f
C2623 vdd.n246 gnd 0.0049f
C2624 vdd.n247 gnd 0.0049f
C2625 vdd.n248 gnd 0.002633f
C2626 vdd.n249 gnd 0.002788f
C2627 vdd.n250 gnd 0.006223f
C2628 vdd.n251 gnd 0.006223f
C2629 vdd.n252 gnd 0.002788f
C2630 vdd.n253 gnd 0.002633f
C2631 vdd.n254 gnd 0.0049f
C2632 vdd.n255 gnd 0.0049f
C2633 vdd.n256 gnd 0.002633f
C2634 vdd.n257 gnd 0.002788f
C2635 vdd.n258 gnd 0.006223f
C2636 vdd.n259 gnd 0.006223f
C2637 vdd.n260 gnd 0.014713f
C2638 vdd.n261 gnd 0.00271f
C2639 vdd.n262 gnd 0.002633f
C2640 vdd.n263 gnd 0.012664f
C2641 vdd.n264 gnd 0.008841f
C2642 vdd.t186 gnd 0.030974f
C2643 vdd.t103 gnd 0.030974f
C2644 vdd.n265 gnd 0.212878f
C2645 vdd.n266 gnd 0.167396f
C2646 vdd.t169 gnd 0.030974f
C2647 vdd.t182 gnd 0.030974f
C2648 vdd.n267 gnd 0.212878f
C2649 vdd.n268 gnd 0.135088f
C2650 vdd.t96 gnd 0.030974f
C2651 vdd.t146 gnd 0.030974f
C2652 vdd.n269 gnd 0.212878f
C2653 vdd.n270 gnd 0.135088f
C2654 vdd.t168 gnd 0.030974f
C2655 vdd.t77 gnd 0.030974f
C2656 vdd.n271 gnd 0.212878f
C2657 vdd.n272 gnd 0.135088f
C2658 vdd.t121 gnd 0.030974f
C2659 vdd.t166 gnd 0.030974f
C2660 vdd.n273 gnd 0.212878f
C2661 vdd.n274 gnd 0.135088f
C2662 vdd.t83 gnd 0.030974f
C2663 vdd.t119 gnd 0.030974f
C2664 vdd.n275 gnd 0.212878f
C2665 vdd.n276 gnd 0.135088f
C2666 vdd.t151 gnd 0.030974f
C2667 vdd.t184 gnd 0.030974f
C2668 vdd.n277 gnd 0.212878f
C2669 vdd.n278 gnd 0.135088f
C2670 vdd.n279 gnd 0.00528f
C2671 vdd.n280 gnd 0.0049f
C2672 vdd.n281 gnd 0.00271f
C2673 vdd.n282 gnd 0.006223f
C2674 vdd.n283 gnd 0.002633f
C2675 vdd.n284 gnd 0.002788f
C2676 vdd.n285 gnd 0.0049f
C2677 vdd.n286 gnd 0.002633f
C2678 vdd.n287 gnd 0.006223f
C2679 vdd.n288 gnd 0.002788f
C2680 vdd.n289 gnd 0.0049f
C2681 vdd.n290 gnd 0.002633f
C2682 vdd.n291 gnd 0.004667f
C2683 vdd.n292 gnd 0.004681f
C2684 vdd.t99 gnd 0.01337f
C2685 vdd.n293 gnd 0.029747f
C2686 vdd.n294 gnd 0.154813f
C2687 vdd.n295 gnd 0.002633f
C2688 vdd.n296 gnd 0.002788f
C2689 vdd.n297 gnd 0.006223f
C2690 vdd.n298 gnd 0.006223f
C2691 vdd.n299 gnd 0.002788f
C2692 vdd.n300 gnd 0.002633f
C2693 vdd.n301 gnd 0.0049f
C2694 vdd.n302 gnd 0.0049f
C2695 vdd.n303 gnd 0.002633f
C2696 vdd.n304 gnd 0.002788f
C2697 vdd.n305 gnd 0.006223f
C2698 vdd.n306 gnd 0.006223f
C2699 vdd.n307 gnd 0.002788f
C2700 vdd.n308 gnd 0.002633f
C2701 vdd.n309 gnd 0.0049f
C2702 vdd.n310 gnd 0.0049f
C2703 vdd.n311 gnd 0.002633f
C2704 vdd.n312 gnd 0.002788f
C2705 vdd.n313 gnd 0.006223f
C2706 vdd.n314 gnd 0.006223f
C2707 vdd.n315 gnd 0.014713f
C2708 vdd.n316 gnd 0.00271f
C2709 vdd.n317 gnd 0.002633f
C2710 vdd.n318 gnd 0.012664f
C2711 vdd.n319 gnd 0.008564f
C2712 vdd.n320 gnd 0.059791f
C2713 vdd.n321 gnd 0.241267f
C2714 vdd.n322 gnd 0.007394f
C2715 vdd.n323 gnd 0.009621f
C2716 vdd.n324 gnd 0.007744f
C2717 vdd.n325 gnd 0.007744f
C2718 vdd.n326 gnd 0.009621f
C2719 vdd.n327 gnd 0.009621f
C2720 vdd.n328 gnd 0.702993f
C2721 vdd.n329 gnd 0.009621f
C2722 vdd.n330 gnd 0.009621f
C2723 vdd.n331 gnd 0.009621f
C2724 vdd.n332 gnd 0.761985f
C2725 vdd.n333 gnd 0.009621f
C2726 vdd.n334 gnd 0.009621f
C2727 vdd.n335 gnd 0.009621f
C2728 vdd.n336 gnd 0.009621f
C2729 vdd.n337 gnd 0.007744f
C2730 vdd.n338 gnd 0.009621f
C2731 vdd.t158 gnd 0.491603f
C2732 vdd.n339 gnd 0.009621f
C2733 vdd.n340 gnd 0.009621f
C2734 vdd.n341 gnd 0.009621f
C2735 vdd.t104 gnd 0.491603f
C2736 vdd.n342 gnd 0.009621f
C2737 vdd.n343 gnd 0.009621f
C2738 vdd.n344 gnd 0.009621f
C2739 vdd.n345 gnd 0.009621f
C2740 vdd.n346 gnd 0.009621f
C2741 vdd.n347 gnd 0.007744f
C2742 vdd.n348 gnd 0.009621f
C2743 vdd.n349 gnd 0.555512f
C2744 vdd.n350 gnd 0.009621f
C2745 vdd.n351 gnd 0.009621f
C2746 vdd.n352 gnd 0.009621f
C2747 vdd.t176 gnd 0.491603f
C2748 vdd.n353 gnd 0.009621f
C2749 vdd.n354 gnd 0.009621f
C2750 vdd.n355 gnd 0.009621f
C2751 vdd.n356 gnd 0.009621f
C2752 vdd.n357 gnd 0.009621f
C2753 vdd.n358 gnd 0.007744f
C2754 vdd.n359 gnd 0.009621f
C2755 vdd.t80 gnd 0.491603f
C2756 vdd.n360 gnd 0.009621f
C2757 vdd.n361 gnd 0.009621f
C2758 vdd.n362 gnd 0.009621f
C2759 vdd.n363 gnd 0.830809f
C2760 vdd.n364 gnd 0.009621f
C2761 vdd.n365 gnd 0.009621f
C2762 vdd.n366 gnd 0.009621f
C2763 vdd.n367 gnd 0.009621f
C2764 vdd.n368 gnd 0.009621f
C2765 vdd.n369 gnd 0.006427f
C2766 vdd.n370 gnd 0.021909f
C2767 vdd.t212 gnd 0.491603f
C2768 vdd.n371 gnd 0.009621f
C2769 vdd.n372 gnd 0.021909f
C2770 vdd.n404 gnd 0.009621f
C2771 vdd.t237 gnd 0.118362f
C2772 vdd.t236 gnd 0.126496f
C2773 vdd.t235 gnd 0.154579f
C2774 vdd.n405 gnd 0.198149f
C2775 vdd.n406 gnd 0.167255f
C2776 vdd.n407 gnd 0.0127f
C2777 vdd.n408 gnd 0.009621f
C2778 vdd.n409 gnd 0.007744f
C2779 vdd.n410 gnd 0.009621f
C2780 vdd.n411 gnd 0.007744f
C2781 vdd.n412 gnd 0.009621f
C2782 vdd.n413 gnd 0.007744f
C2783 vdd.n414 gnd 0.009621f
C2784 vdd.n415 gnd 0.007744f
C2785 vdd.n416 gnd 0.009621f
C2786 vdd.n417 gnd 0.007744f
C2787 vdd.n418 gnd 0.009621f
C2788 vdd.t214 gnd 0.118362f
C2789 vdd.t213 gnd 0.126496f
C2790 vdd.t211 gnd 0.154579f
C2791 vdd.n419 gnd 0.198149f
C2792 vdd.n420 gnd 0.167255f
C2793 vdd.n421 gnd 0.007744f
C2794 vdd.n422 gnd 0.009621f
C2795 vdd.n423 gnd 0.007744f
C2796 vdd.n424 gnd 0.009621f
C2797 vdd.n425 gnd 0.007744f
C2798 vdd.n426 gnd 0.009621f
C2799 vdd.n427 gnd 0.007744f
C2800 vdd.n428 gnd 0.009621f
C2801 vdd.n429 gnd 0.007744f
C2802 vdd.n430 gnd 0.009621f
C2803 vdd.t228 gnd 0.118362f
C2804 vdd.t227 gnd 0.126496f
C2805 vdd.t226 gnd 0.154579f
C2806 vdd.n431 gnd 0.198149f
C2807 vdd.n432 gnd 0.167255f
C2808 vdd.n433 gnd 0.016571f
C2809 vdd.n434 gnd 0.009621f
C2810 vdd.n435 gnd 0.007744f
C2811 vdd.n436 gnd 0.009621f
C2812 vdd.n437 gnd 0.007744f
C2813 vdd.n438 gnd 0.009621f
C2814 vdd.n439 gnd 0.007744f
C2815 vdd.n440 gnd 0.009621f
C2816 vdd.n441 gnd 0.007744f
C2817 vdd.n442 gnd 0.009621f
C2818 vdd.n443 gnd 0.021909f
C2819 vdd.n444 gnd 0.022059f
C2820 vdd.n445 gnd 0.022059f
C2821 vdd.n446 gnd 0.006427f
C2822 vdd.n447 gnd 0.007744f
C2823 vdd.n448 gnd 0.009621f
C2824 vdd.n449 gnd 0.009621f
C2825 vdd.n450 gnd 0.007744f
C2826 vdd.n451 gnd 0.009621f
C2827 vdd.n452 gnd 0.009621f
C2828 vdd.n453 gnd 0.009621f
C2829 vdd.n454 gnd 0.009621f
C2830 vdd.n455 gnd 0.009621f
C2831 vdd.n456 gnd 0.007744f
C2832 vdd.n457 gnd 0.007744f
C2833 vdd.n458 gnd 0.009621f
C2834 vdd.n459 gnd 0.009621f
C2835 vdd.n460 gnd 0.007744f
C2836 vdd.n461 gnd 0.009621f
C2837 vdd.n462 gnd 0.009621f
C2838 vdd.n463 gnd 0.009621f
C2839 vdd.n464 gnd 0.009621f
C2840 vdd.n465 gnd 0.009621f
C2841 vdd.n466 gnd 0.007744f
C2842 vdd.n467 gnd 0.007744f
C2843 vdd.n468 gnd 0.009621f
C2844 vdd.n469 gnd 0.009621f
C2845 vdd.n470 gnd 0.007744f
C2846 vdd.n471 gnd 0.009621f
C2847 vdd.n472 gnd 0.009621f
C2848 vdd.n473 gnd 0.009621f
C2849 vdd.n474 gnd 0.009621f
C2850 vdd.n475 gnd 0.009621f
C2851 vdd.n476 gnd 0.007744f
C2852 vdd.n477 gnd 0.007744f
C2853 vdd.n478 gnd 0.009621f
C2854 vdd.n479 gnd 0.009621f
C2855 vdd.n480 gnd 0.007744f
C2856 vdd.n481 gnd 0.009621f
C2857 vdd.n482 gnd 0.009621f
C2858 vdd.n483 gnd 0.009621f
C2859 vdd.n484 gnd 0.009621f
C2860 vdd.n485 gnd 0.009621f
C2861 vdd.n486 gnd 0.007744f
C2862 vdd.n487 gnd 0.007744f
C2863 vdd.n488 gnd 0.009621f
C2864 vdd.n489 gnd 0.009621f
C2865 vdd.n490 gnd 0.006466f
C2866 vdd.n491 gnd 0.009621f
C2867 vdd.n492 gnd 0.009621f
C2868 vdd.n493 gnd 0.009621f
C2869 vdd.n494 gnd 0.009621f
C2870 vdd.n495 gnd 0.009621f
C2871 vdd.n496 gnd 0.006466f
C2872 vdd.n497 gnd 0.007744f
C2873 vdd.n498 gnd 0.009621f
C2874 vdd.n499 gnd 0.009621f
C2875 vdd.n500 gnd 0.007744f
C2876 vdd.n501 gnd 0.009621f
C2877 vdd.n502 gnd 0.009621f
C2878 vdd.n503 gnd 0.009621f
C2879 vdd.n504 gnd 0.009621f
C2880 vdd.n505 gnd 0.009621f
C2881 vdd.n506 gnd 0.007744f
C2882 vdd.n507 gnd 0.007744f
C2883 vdd.n508 gnd 0.009621f
C2884 vdd.n509 gnd 0.009621f
C2885 vdd.n510 gnd 0.007744f
C2886 vdd.n511 gnd 0.009621f
C2887 vdd.n512 gnd 0.009621f
C2888 vdd.n513 gnd 0.009621f
C2889 vdd.n514 gnd 0.009621f
C2890 vdd.n515 gnd 0.009621f
C2891 vdd.n516 gnd 0.007744f
C2892 vdd.n517 gnd 0.007744f
C2893 vdd.n518 gnd 0.009621f
C2894 vdd.n519 gnd 0.009621f
C2895 vdd.n520 gnd 0.007744f
C2896 vdd.n521 gnd 0.009621f
C2897 vdd.n522 gnd 0.009621f
C2898 vdd.n523 gnd 0.009621f
C2899 vdd.n524 gnd 0.009621f
C2900 vdd.n525 gnd 0.009621f
C2901 vdd.n526 gnd 0.007744f
C2902 vdd.n527 gnd 0.007744f
C2903 vdd.n528 gnd 0.009621f
C2904 vdd.n529 gnd 0.009621f
C2905 vdd.n530 gnd 0.007744f
C2906 vdd.n531 gnd 0.009621f
C2907 vdd.n532 gnd 0.009621f
C2908 vdd.n533 gnd 0.009621f
C2909 vdd.n534 gnd 0.009621f
C2910 vdd.n535 gnd 0.009621f
C2911 vdd.n536 gnd 0.007744f
C2912 vdd.n537 gnd 0.007744f
C2913 vdd.n538 gnd 0.009621f
C2914 vdd.n539 gnd 0.009621f
C2915 vdd.n540 gnd 0.007744f
C2916 vdd.n541 gnd 0.009621f
C2917 vdd.n542 gnd 0.009621f
C2918 vdd.n543 gnd 0.009621f
C2919 vdd.n544 gnd 0.009621f
C2920 vdd.n545 gnd 0.009621f
C2921 vdd.n546 gnd 0.005266f
C2922 vdd.n547 gnd 0.016571f
C2923 vdd.n548 gnd 0.009621f
C2924 vdd.n549 gnd 0.009621f
C2925 vdd.n550 gnd 0.007666f
C2926 vdd.n551 gnd 0.009621f
C2927 vdd.n552 gnd 0.009621f
C2928 vdd.n553 gnd 0.009621f
C2929 vdd.n554 gnd 0.009621f
C2930 vdd.n555 gnd 0.009621f
C2931 vdd.n556 gnd 0.007744f
C2932 vdd.n557 gnd 0.007744f
C2933 vdd.n558 gnd 0.009621f
C2934 vdd.n559 gnd 0.009621f
C2935 vdd.n560 gnd 0.007744f
C2936 vdd.n561 gnd 0.009621f
C2937 vdd.n562 gnd 0.009621f
C2938 vdd.n563 gnd 0.009621f
C2939 vdd.n564 gnd 0.009621f
C2940 vdd.n565 gnd 0.009621f
C2941 vdd.n566 gnd 0.007744f
C2942 vdd.n567 gnd 0.007744f
C2943 vdd.n568 gnd 0.009621f
C2944 vdd.n569 gnd 0.009621f
C2945 vdd.n570 gnd 0.007744f
C2946 vdd.n571 gnd 0.009621f
C2947 vdd.n572 gnd 0.009621f
C2948 vdd.n573 gnd 0.009621f
C2949 vdd.n574 gnd 0.009621f
C2950 vdd.n575 gnd 0.009621f
C2951 vdd.n576 gnd 0.007744f
C2952 vdd.n577 gnd 0.007744f
C2953 vdd.n578 gnd 0.009621f
C2954 vdd.n579 gnd 0.009621f
C2955 vdd.n580 gnd 0.007744f
C2956 vdd.n581 gnd 0.009621f
C2957 vdd.n582 gnd 0.009621f
C2958 vdd.n583 gnd 0.009621f
C2959 vdd.n584 gnd 0.009621f
C2960 vdd.n585 gnd 0.009621f
C2961 vdd.n586 gnd 0.007744f
C2962 vdd.n587 gnd 0.007744f
C2963 vdd.n588 gnd 0.009621f
C2964 vdd.n589 gnd 0.009621f
C2965 vdd.n590 gnd 0.007744f
C2966 vdd.n591 gnd 0.009621f
C2967 vdd.n592 gnd 0.009621f
C2968 vdd.n593 gnd 0.009621f
C2969 vdd.n594 gnd 0.009621f
C2970 vdd.n595 gnd 0.009621f
C2971 vdd.n596 gnd 0.007744f
C2972 vdd.n597 gnd 0.009621f
C2973 vdd.n598 gnd 0.007744f
C2974 vdd.n599 gnd 0.004065f
C2975 vdd.n600 gnd 0.009621f
C2976 vdd.n601 gnd 0.009621f
C2977 vdd.n602 gnd 0.007744f
C2978 vdd.n603 gnd 0.009621f
C2979 vdd.n604 gnd 0.007744f
C2980 vdd.n605 gnd 0.009621f
C2981 vdd.n606 gnd 0.007744f
C2982 vdd.n607 gnd 0.009621f
C2983 vdd.n608 gnd 0.007744f
C2984 vdd.n609 gnd 0.009621f
C2985 vdd.n610 gnd 0.007744f
C2986 vdd.n611 gnd 0.009621f
C2987 vdd.n612 gnd 0.009621f
C2988 vdd.n613 gnd 0.535848f
C2989 vdd.t116 gnd 0.491603f
C2990 vdd.n614 gnd 0.009621f
C2991 vdd.n615 gnd 0.007744f
C2992 vdd.n616 gnd 0.009621f
C2993 vdd.n617 gnd 0.007744f
C2994 vdd.n618 gnd 0.009621f
C2995 vdd.t70 gnd 0.491603f
C2996 vdd.n619 gnd 0.009621f
C2997 vdd.n620 gnd 0.007744f
C2998 vdd.n621 gnd 0.009621f
C2999 vdd.n622 gnd 0.007744f
C3000 vdd.n623 gnd 0.009621f
C3001 vdd.t154 gnd 0.491603f
C3002 vdd.n624 gnd 0.614504f
C3003 vdd.n625 gnd 0.009621f
C3004 vdd.n626 gnd 0.007744f
C3005 vdd.n627 gnd 0.009621f
C3006 vdd.n628 gnd 0.007744f
C3007 vdd.n629 gnd 0.009621f
C3008 vdd.t87 gnd 0.491603f
C3009 vdd.n630 gnd 0.009621f
C3010 vdd.n631 gnd 0.007744f
C3011 vdd.n632 gnd 0.009621f
C3012 vdd.n633 gnd 0.007744f
C3013 vdd.n634 gnd 0.009621f
C3014 vdd.n635 gnd 0.683328f
C3015 vdd.n636 gnd 0.816061f
C3016 vdd.t84 gnd 0.491603f
C3017 vdd.n637 gnd 0.009621f
C3018 vdd.n638 gnd 0.007744f
C3019 vdd.n639 gnd 0.009621f
C3020 vdd.n640 gnd 0.007744f
C3021 vdd.n641 gnd 0.009621f
C3022 vdd.n642 gnd 0.516183f
C3023 vdd.n643 gnd 0.009621f
C3024 vdd.n644 gnd 0.007744f
C3025 vdd.n645 gnd 0.009621f
C3026 vdd.n646 gnd 0.007744f
C3027 vdd.n647 gnd 0.009621f
C3028 vdd.n648 gnd 0.983206f
C3029 vdd.t129 gnd 0.491603f
C3030 vdd.n649 gnd 0.009621f
C3031 vdd.n650 gnd 0.007744f
C3032 vdd.n651 gnd 0.009621f
C3033 vdd.n652 gnd 0.007744f
C3034 vdd.n653 gnd 0.009621f
C3035 vdd.t216 gnd 0.491603f
C3036 vdd.n654 gnd 0.009621f
C3037 vdd.n655 gnd 0.007744f
C3038 vdd.n656 gnd 0.022059f
C3039 vdd.n657 gnd 0.022059f
C3040 vdd.n658 gnd 11.8476f
C3041 vdd.n659 gnd 0.54568f
C3042 vdd.n660 gnd 0.022059f
C3043 vdd.n661 gnd 0.008274f
C3044 vdd.n662 gnd 0.007744f
C3045 vdd.n667 gnd 0.006157f
C3046 vdd.n668 gnd 0.007744f
C3047 vdd.n669 gnd 0.009621f
C3048 vdd.n670 gnd 0.009621f
C3049 vdd.n671 gnd 0.009621f
C3050 vdd.n672 gnd 0.009621f
C3051 vdd.n673 gnd 0.009621f
C3052 vdd.n674 gnd 0.007744f
C3053 vdd.n675 gnd 0.009621f
C3054 vdd.n676 gnd 0.009621f
C3055 vdd.n677 gnd 0.009621f
C3056 vdd.n678 gnd 0.009621f
C3057 vdd.n679 gnd 0.009621f
C3058 vdd.n680 gnd 0.007744f
C3059 vdd.n681 gnd 0.009621f
C3060 vdd.n682 gnd 0.009621f
C3061 vdd.n683 gnd 0.009621f
C3062 vdd.n684 gnd 0.009621f
C3063 vdd.n685 gnd 0.009621f
C3064 vdd.t247 gnd 0.118362f
C3065 vdd.t248 gnd 0.126496f
C3066 vdd.t246 gnd 0.154579f
C3067 vdd.n686 gnd 0.198149f
C3068 vdd.n687 gnd 0.166481f
C3069 vdd.n688 gnd 0.015797f
C3070 vdd.n689 gnd 0.009621f
C3071 vdd.n690 gnd 0.009621f
C3072 vdd.n691 gnd 0.009621f
C3073 vdd.n692 gnd 0.009621f
C3074 vdd.n693 gnd 0.009621f
C3075 vdd.n694 gnd 0.007744f
C3076 vdd.n695 gnd 0.009621f
C3077 vdd.n696 gnd 0.009621f
C3078 vdd.n697 gnd 0.009621f
C3079 vdd.n698 gnd 0.009621f
C3080 vdd.n699 gnd 0.009621f
C3081 vdd.n700 gnd 0.007744f
C3082 vdd.n701 gnd 0.009621f
C3083 vdd.n702 gnd 0.009621f
C3084 vdd.n703 gnd 0.009621f
C3085 vdd.n704 gnd 0.009621f
C3086 vdd.n705 gnd 0.009621f
C3087 vdd.n706 gnd 0.007744f
C3088 vdd.n707 gnd 0.009621f
C3089 vdd.n708 gnd 0.009621f
C3090 vdd.n709 gnd 0.009621f
C3091 vdd.n710 gnd 0.009621f
C3092 vdd.n711 gnd 0.009621f
C3093 vdd.n712 gnd 0.007744f
C3094 vdd.n713 gnd 0.009621f
C3095 vdd.n714 gnd 0.009621f
C3096 vdd.n715 gnd 0.009621f
C3097 vdd.n716 gnd 0.009621f
C3098 vdd.n717 gnd 0.009621f
C3099 vdd.n718 gnd 0.007744f
C3100 vdd.n719 gnd 0.009621f
C3101 vdd.n720 gnd 0.009621f
C3102 vdd.n721 gnd 0.009621f
C3103 vdd.n722 gnd 0.007666f
C3104 vdd.t230 gnd 0.118362f
C3105 vdd.t231 gnd 0.126496f
C3106 vdd.t229 gnd 0.154579f
C3107 vdd.n723 gnd 0.198149f
C3108 vdd.n724 gnd 0.166481f
C3109 vdd.n725 gnd 0.009621f
C3110 vdd.n726 gnd 0.007744f
C3111 vdd.n728 gnd 0.009621f
C3112 vdd.n730 gnd 0.009621f
C3113 vdd.n731 gnd 0.009621f
C3114 vdd.n732 gnd 0.007744f
C3115 vdd.n733 gnd 0.009621f
C3116 vdd.n734 gnd 0.009621f
C3117 vdd.n735 gnd 0.009621f
C3118 vdd.n736 gnd 0.009621f
C3119 vdd.n737 gnd 0.009621f
C3120 vdd.n738 gnd 0.007744f
C3121 vdd.n739 gnd 0.009621f
C3122 vdd.n740 gnd 0.009621f
C3123 vdd.n741 gnd 0.009621f
C3124 vdd.n742 gnd 0.009621f
C3125 vdd.n743 gnd 0.009621f
C3126 vdd.n744 gnd 0.007744f
C3127 vdd.n745 gnd 0.009621f
C3128 vdd.n746 gnd 0.009621f
C3129 vdd.n747 gnd 0.009621f
C3130 vdd.n748 gnd 0.006157f
C3131 vdd.n753 gnd 0.006542f
C3132 vdd.n754 gnd 0.006542f
C3133 vdd.n755 gnd 0.006542f
C3134 vdd.n756 gnd 11.6117f
C3135 vdd.n757 gnd 0.006542f
C3136 vdd.n758 gnd 0.006542f
C3137 vdd.n759 gnd 0.006542f
C3138 vdd.n761 gnd 0.006542f
C3139 vdd.n762 gnd 0.006542f
C3140 vdd.n764 gnd 0.006542f
C3141 vdd.n765 gnd 0.004762f
C3142 vdd.n767 gnd 0.006542f
C3143 vdd.t196 gnd 0.264369f
C3144 vdd.t195 gnd 0.270614f
C3145 vdd.t193 gnd 0.17259f
C3146 vdd.n768 gnd 0.093276f
C3147 vdd.n769 gnd 0.052909f
C3148 vdd.n770 gnd 0.00935f
C3149 vdd.n771 gnd 0.014855f
C3150 vdd.n773 gnd 0.006542f
C3151 vdd.n774 gnd 0.66858f
C3152 vdd.n775 gnd 0.014008f
C3153 vdd.n776 gnd 0.014008f
C3154 vdd.n777 gnd 0.006542f
C3155 vdd.n778 gnd 0.014855f
C3156 vdd.n779 gnd 0.006542f
C3157 vdd.n780 gnd 0.006542f
C3158 vdd.n781 gnd 0.006542f
C3159 vdd.n782 gnd 0.006542f
C3160 vdd.n783 gnd 0.006542f
C3161 vdd.n785 gnd 0.006542f
C3162 vdd.n786 gnd 0.006542f
C3163 vdd.n788 gnd 0.006542f
C3164 vdd.n789 gnd 0.006542f
C3165 vdd.n791 gnd 0.006542f
C3166 vdd.n792 gnd 0.006542f
C3167 vdd.n794 gnd 0.006542f
C3168 vdd.n795 gnd 0.006542f
C3169 vdd.n797 gnd 0.006542f
C3170 vdd.n798 gnd 0.006542f
C3171 vdd.n800 gnd 0.006542f
C3172 vdd.n801 gnd 0.004762f
C3173 vdd.n803 gnd 0.006542f
C3174 vdd.t210 gnd 0.264369f
C3175 vdd.t209 gnd 0.270614f
C3176 vdd.t208 gnd 0.17259f
C3177 vdd.n804 gnd 0.093276f
C3178 vdd.n805 gnd 0.052909f
C3179 vdd.n806 gnd 0.00935f
C3180 vdd.n807 gnd 0.006542f
C3181 vdd.n808 gnd 0.006542f
C3182 vdd.t194 gnd 0.33429f
C3183 vdd.n809 gnd 0.006542f
C3184 vdd.n810 gnd 0.006542f
C3185 vdd.n811 gnd 0.006542f
C3186 vdd.n812 gnd 0.006542f
C3187 vdd.n813 gnd 0.006542f
C3188 vdd.n814 gnd 0.66858f
C3189 vdd.n815 gnd 0.006542f
C3190 vdd.n816 gnd 0.006542f
C3191 vdd.n817 gnd 0.526015f
C3192 vdd.n818 gnd 0.006542f
C3193 vdd.n819 gnd 0.006542f
C3194 vdd.n820 gnd 0.006542f
C3195 vdd.n821 gnd 0.006542f
C3196 vdd.n822 gnd 0.66858f
C3197 vdd.n823 gnd 0.006542f
C3198 vdd.n824 gnd 0.006542f
C3199 vdd.n825 gnd 0.006542f
C3200 vdd.n826 gnd 0.006542f
C3201 vdd.n827 gnd 0.006542f
C3202 vdd.t16 gnd 0.33429f
C3203 vdd.n828 gnd 0.006542f
C3204 vdd.n829 gnd 0.006542f
C3205 vdd.n830 gnd 0.006542f
C3206 vdd.n831 gnd 0.006542f
C3207 vdd.n832 gnd 0.006542f
C3208 vdd.t33 gnd 0.33429f
C3209 vdd.n833 gnd 0.006542f
C3210 vdd.n834 gnd 0.006542f
C3211 vdd.n835 gnd 0.644f
C3212 vdd.n836 gnd 0.006542f
C3213 vdd.n837 gnd 0.006542f
C3214 vdd.n838 gnd 0.006542f
C3215 vdd.t32 gnd 0.33429f
C3216 vdd.n839 gnd 0.006542f
C3217 vdd.n840 gnd 0.006542f
C3218 vdd.n841 gnd 0.496519f
C3219 vdd.n842 gnd 0.006542f
C3220 vdd.n843 gnd 0.006542f
C3221 vdd.n844 gnd 0.006542f
C3222 vdd.n845 gnd 0.467023f
C3223 vdd.n846 gnd 0.006542f
C3224 vdd.n847 gnd 0.006542f
C3225 vdd.n848 gnd 0.349038f
C3226 vdd.n849 gnd 0.006542f
C3227 vdd.n850 gnd 0.006542f
C3228 vdd.n851 gnd 0.006542f
C3229 vdd.n852 gnd 0.614504f
C3230 vdd.n853 gnd 0.006542f
C3231 vdd.n854 gnd 0.006542f
C3232 vdd.t39 gnd 0.33429f
C3233 vdd.n855 gnd 0.006542f
C3234 vdd.n856 gnd 0.006542f
C3235 vdd.n857 gnd 0.006542f
C3236 vdd.n858 gnd 0.66858f
C3237 vdd.n859 gnd 0.006542f
C3238 vdd.n860 gnd 0.006542f
C3239 vdd.t40 gnd 0.33429f
C3240 vdd.n861 gnd 0.006542f
C3241 vdd.n862 gnd 0.006542f
C3242 vdd.n863 gnd 0.006542f
C3243 vdd.t10 gnd 0.33429f
C3244 vdd.n864 gnd 0.006542f
C3245 vdd.n865 gnd 0.006542f
C3246 vdd.n866 gnd 0.006542f
C3247 vdd.t221 gnd 0.270614f
C3248 vdd.t219 gnd 0.17259f
C3249 vdd.t222 gnd 0.270614f
C3250 vdd.n867 gnd 0.152096f
C3251 vdd.n868 gnd 0.018952f
C3252 vdd.n869 gnd 0.006542f
C3253 vdd.t220 gnd 0.240886f
C3254 vdd.n870 gnd 0.006542f
C3255 vdd.n871 gnd 0.006542f
C3256 vdd.n872 gnd 0.575176f
C3257 vdd.n873 gnd 0.006542f
C3258 vdd.n874 gnd 0.006542f
C3259 vdd.n875 gnd 0.006542f
C3260 vdd.n876 gnd 0.388367f
C3261 vdd.n877 gnd 0.006542f
C3262 vdd.n878 gnd 0.006542f
C3263 vdd.t11 gnd 0.137649f
C3264 vdd.n879 gnd 0.427695f
C3265 vdd.n880 gnd 0.006542f
C3266 vdd.n881 gnd 0.006542f
C3267 vdd.n882 gnd 0.006542f
C3268 vdd.n883 gnd 0.535848f
C3269 vdd.n884 gnd 0.006542f
C3270 vdd.n885 gnd 0.006542f
C3271 vdd.t24 gnd 0.33429f
C3272 vdd.n886 gnd 0.006542f
C3273 vdd.n887 gnd 0.006542f
C3274 vdd.n888 gnd 0.006542f
C3275 vdd.t20 gnd 0.33429f
C3276 vdd.n889 gnd 0.006542f
C3277 vdd.n890 gnd 0.006542f
C3278 vdd.t43 gnd 0.33429f
C3279 vdd.n891 gnd 0.006542f
C3280 vdd.n892 gnd 0.006542f
C3281 vdd.n893 gnd 0.006542f
C3282 vdd.t2 gnd 0.226137f
C3283 vdd.n894 gnd 0.006542f
C3284 vdd.n895 gnd 0.006542f
C3285 vdd.n896 gnd 0.589924f
C3286 vdd.n897 gnd 0.006542f
C3287 vdd.n898 gnd 0.006542f
C3288 vdd.n899 gnd 0.006542f
C3289 vdd.t44 gnd 0.33429f
C3290 vdd.n900 gnd 0.006542f
C3291 vdd.n901 gnd 0.006542f
C3292 vdd.t56 gnd 0.319542f
C3293 vdd.n902 gnd 0.442443f
C3294 vdd.n903 gnd 0.006542f
C3295 vdd.n904 gnd 0.006542f
C3296 vdd.n905 gnd 0.006542f
C3297 vdd.t6 gnd 0.33429f
C3298 vdd.n906 gnd 0.006542f
C3299 vdd.n907 gnd 0.006542f
C3300 vdd.t48 gnd 0.33429f
C3301 vdd.n908 gnd 0.006542f
C3302 vdd.n909 gnd 0.006542f
C3303 vdd.n910 gnd 0.006542f
C3304 vdd.n911 gnd 0.66858f
C3305 vdd.n912 gnd 0.006542f
C3306 vdd.n913 gnd 0.006542f
C3307 vdd.t28 gnd 0.33429f
C3308 vdd.n914 gnd 0.006542f
C3309 vdd.n915 gnd 0.006542f
C3310 vdd.n916 gnd 0.006542f
C3311 vdd.n917 gnd 0.462107f
C3312 vdd.n918 gnd 0.006542f
C3313 vdd.n919 gnd 0.006542f
C3314 vdd.n920 gnd 0.006542f
C3315 vdd.n921 gnd 0.006542f
C3316 vdd.n922 gnd 0.006542f
C3317 vdd.t250 gnd 0.33429f
C3318 vdd.n923 gnd 0.006542f
C3319 vdd.n924 gnd 0.006542f
C3320 vdd.t8 gnd 0.33429f
C3321 vdd.n925 gnd 0.006542f
C3322 vdd.n926 gnd 0.014008f
C3323 vdd.n927 gnd 0.014008f
C3324 vdd.n928 gnd 0.757069f
C3325 vdd.n929 gnd 0.006542f
C3326 vdd.n930 gnd 0.006542f
C3327 vdd.t37 gnd 0.33429f
C3328 vdd.n931 gnd 0.014008f
C3329 vdd.n932 gnd 0.006542f
C3330 vdd.n933 gnd 0.006542f
C3331 vdd.t50 gnd 0.57026f
C3332 vdd.n951 gnd 0.014855f
C3333 vdd.n969 gnd 0.014008f
C3334 vdd.n970 gnd 0.006542f
C3335 vdd.n971 gnd 0.014008f
C3336 vdd.t268 gnd 0.264369f
C3337 vdd.t267 gnd 0.270614f
C3338 vdd.t266 gnd 0.17259f
C3339 vdd.n972 gnd 0.093276f
C3340 vdd.n973 gnd 0.052909f
C3341 vdd.n974 gnd 0.014855f
C3342 vdd.n975 gnd 0.006542f
C3343 vdd.n976 gnd 0.393283f
C3344 vdd.n977 gnd 0.014008f
C3345 vdd.n978 gnd 0.006542f
C3346 vdd.n979 gnd 0.014855f
C3347 vdd.n980 gnd 0.006542f
C3348 vdd.t245 gnd 0.264369f
C3349 vdd.t244 gnd 0.270614f
C3350 vdd.t242 gnd 0.17259f
C3351 vdd.n981 gnd 0.093276f
C3352 vdd.n982 gnd 0.052909f
C3353 vdd.n983 gnd 0.00935f
C3354 vdd.n984 gnd 0.006542f
C3355 vdd.n985 gnd 0.006542f
C3356 vdd.t243 gnd 0.33429f
C3357 vdd.n986 gnd 0.006542f
C3358 vdd.t52 gnd 0.33429f
C3359 vdd.n987 gnd 0.006542f
C3360 vdd.n988 gnd 0.006542f
C3361 vdd.n989 gnd 0.006542f
C3362 vdd.n990 gnd 0.006542f
C3363 vdd.n991 gnd 0.006542f
C3364 vdd.n992 gnd 0.66858f
C3365 vdd.n993 gnd 0.006542f
C3366 vdd.n994 gnd 0.006542f
C3367 vdd.t22 gnd 0.33429f
C3368 vdd.n995 gnd 0.006542f
C3369 vdd.n996 gnd 0.006542f
C3370 vdd.n997 gnd 0.006542f
C3371 vdd.n998 gnd 0.006542f
C3372 vdd.n999 gnd 0.481771f
C3373 vdd.n1000 gnd 0.006542f
C3374 vdd.n1001 gnd 0.006542f
C3375 vdd.n1002 gnd 0.006542f
C3376 vdd.n1003 gnd 0.006542f
C3377 vdd.n1004 gnd 0.006542f
C3378 vdd.t3 gnd 0.33429f
C3379 vdd.n1005 gnd 0.006542f
C3380 vdd.n1006 gnd 0.006542f
C3381 vdd.t41 gnd 0.33429f
C3382 vdd.n1007 gnd 0.006542f
C3383 vdd.n1008 gnd 0.006542f
C3384 vdd.n1009 gnd 0.006542f
C3385 vdd.t27 gnd 0.33429f
C3386 vdd.n1010 gnd 0.006542f
C3387 vdd.n1011 gnd 0.006542f
C3388 vdd.t4 gnd 0.33429f
C3389 vdd.n1012 gnd 0.006542f
C3390 vdd.n1013 gnd 0.006542f
C3391 vdd.n1014 gnd 0.006542f
C3392 vdd.t25 gnd 0.319542f
C3393 vdd.n1015 gnd 0.006542f
C3394 vdd.n1016 gnd 0.006542f
C3395 vdd.n1017 gnd 0.496519f
C3396 vdd.n1018 gnd 0.006542f
C3397 vdd.n1019 gnd 0.006542f
C3398 vdd.n1020 gnd 0.006542f
C3399 vdd.t45 gnd 0.33429f
C3400 vdd.n1021 gnd 0.006542f
C3401 vdd.n1022 gnd 0.006542f
C3402 vdd.t13 gnd 0.226137f
C3403 vdd.n1023 gnd 0.349038f
C3404 vdd.n1024 gnd 0.006542f
C3405 vdd.n1025 gnd 0.006542f
C3406 vdd.n1026 gnd 0.006542f
C3407 vdd.n1027 gnd 0.614504f
C3408 vdd.n1028 gnd 0.006542f
C3409 vdd.n1029 gnd 0.006542f
C3410 vdd.t54 gnd 0.33429f
C3411 vdd.n1030 gnd 0.006542f
C3412 vdd.n1031 gnd 0.006542f
C3413 vdd.n1032 gnd 0.006542f
C3414 vdd.n1033 gnd 0.66858f
C3415 vdd.n1034 gnd 0.006542f
C3416 vdd.n1035 gnd 0.006542f
C3417 vdd.t19 gnd 0.33429f
C3418 vdd.n1036 gnd 0.006542f
C3419 vdd.n1037 gnd 0.006542f
C3420 vdd.n1038 gnd 0.006542f
C3421 vdd.t12 gnd 0.137649f
C3422 vdd.n1039 gnd 0.006542f
C3423 vdd.n1040 gnd 0.006542f
C3424 vdd.n1041 gnd 0.006542f
C3425 vdd.t258 gnd 0.270614f
C3426 vdd.t256 gnd 0.17259f
C3427 vdd.t259 gnd 0.270614f
C3428 vdd.n1042 gnd 0.152096f
C3429 vdd.n1043 gnd 0.006542f
C3430 vdd.n1044 gnd 0.006542f
C3431 vdd.t34 gnd 0.33429f
C3432 vdd.n1045 gnd 0.006542f
C3433 vdd.n1046 gnd 0.006542f
C3434 vdd.t257 gnd 0.240886f
C3435 vdd.n1047 gnd 0.530931f
C3436 vdd.n1048 gnd 0.006542f
C3437 vdd.n1049 gnd 0.006542f
C3438 vdd.n1050 gnd 0.006542f
C3439 vdd.n1051 gnd 0.388367f
C3440 vdd.n1052 gnd 0.006542f
C3441 vdd.n1053 gnd 0.006542f
C3442 vdd.n1054 gnd 0.427695f
C3443 vdd.n1055 gnd 0.006542f
C3444 vdd.n1056 gnd 0.006542f
C3445 vdd.n1057 gnd 0.006542f
C3446 vdd.n1058 gnd 0.535848f
C3447 vdd.n1059 gnd 0.006542f
C3448 vdd.n1060 gnd 0.006542f
C3449 vdd.t14 gnd 0.33429f
C3450 vdd.n1061 gnd 0.006542f
C3451 vdd.n1062 gnd 0.006542f
C3452 vdd.n1063 gnd 0.006542f
C3453 vdd.n1064 gnd 0.66858f
C3454 vdd.n1065 gnd 0.006542f
C3455 vdd.n1066 gnd 0.006542f
C3456 vdd.t15 gnd 0.33429f
C3457 vdd.n1067 gnd 0.006542f
C3458 vdd.n1068 gnd 0.006542f
C3459 vdd.n1069 gnd 0.006542f
C3460 vdd.t55 gnd 0.33429f
C3461 vdd.n1070 gnd 0.006542f
C3462 vdd.n1071 gnd 0.006542f
C3463 vdd.n1072 gnd 0.006542f
C3464 vdd.n1073 gnd 0.006542f
C3465 vdd.n1074 gnd 0.006542f
C3466 vdd.t47 gnd 0.33429f
C3467 vdd.n1075 gnd 0.006542f
C3468 vdd.n1076 gnd 0.006542f
C3469 vdd.n1077 gnd 0.653832f
C3470 vdd.n1078 gnd 0.006542f
C3471 vdd.n1079 gnd 0.006542f
C3472 vdd.n1080 gnd 0.006542f
C3473 vdd.t7 gnd 0.33429f
C3474 vdd.n1081 gnd 0.006542f
C3475 vdd.n1082 gnd 0.006542f
C3476 vdd.n1083 gnd 0.506351f
C3477 vdd.n1084 gnd 0.006542f
C3478 vdd.n1085 gnd 0.006542f
C3479 vdd.n1086 gnd 0.006542f
C3480 vdd.n1087 gnd 0.66858f
C3481 vdd.n1088 gnd 0.006542f
C3482 vdd.n1089 gnd 0.006542f
C3483 vdd.n1090 gnd 0.35887f
C3484 vdd.n1091 gnd 0.006542f
C3485 vdd.n1092 gnd 0.006542f
C3486 vdd.n1093 gnd 0.006542f
C3487 vdd.n1094 gnd 0.66858f
C3488 vdd.n1095 gnd 0.006542f
C3489 vdd.n1096 gnd 0.006542f
C3490 vdd.n1097 gnd 0.006542f
C3491 vdd.n1098 gnd 0.006542f
C3492 vdd.n1099 gnd 0.006542f
C3493 vdd.t198 gnd 0.33429f
C3494 vdd.n1100 gnd 0.006542f
C3495 vdd.n1101 gnd 0.006542f
C3496 vdd.n1102 gnd 0.006542f
C3497 vdd.n1103 gnd 0.014008f
C3498 vdd.n1104 gnd 0.014008f
C3499 vdd.n1105 gnd 0.90455f
C3500 vdd.n1106 gnd 0.006542f
C3501 vdd.n1107 gnd 0.006542f
C3502 vdd.n1108 gnd 0.476855f
C3503 vdd.n1109 gnd 0.014008f
C3504 vdd.n1110 gnd 0.006542f
C3505 vdd.n1111 gnd 0.006542f
C3506 vdd.n1112 gnd 11.8476f
C3507 vdd.n1146 gnd 0.014855f
C3508 vdd.n1147 gnd 0.006542f
C3509 vdd.n1148 gnd 0.006542f
C3510 vdd.n1149 gnd 0.006157f
C3511 vdd.n1152 gnd 0.022059f
C3512 vdd.n1153 gnd 0.006427f
C3513 vdd.n1154 gnd 0.007744f
C3514 vdd.n1156 gnd 0.009621f
C3515 vdd.n1157 gnd 0.009621f
C3516 vdd.n1158 gnd 0.007744f
C3517 vdd.n1160 gnd 0.009621f
C3518 vdd.n1161 gnd 0.009621f
C3519 vdd.n1162 gnd 0.009621f
C3520 vdd.n1163 gnd 0.009621f
C3521 vdd.n1164 gnd 0.009621f
C3522 vdd.n1165 gnd 0.007744f
C3523 vdd.n1167 gnd 0.009621f
C3524 vdd.n1168 gnd 0.009621f
C3525 vdd.n1169 gnd 0.009621f
C3526 vdd.n1170 gnd 0.009621f
C3527 vdd.n1171 gnd 0.009621f
C3528 vdd.n1172 gnd 0.007744f
C3529 vdd.n1174 gnd 0.009621f
C3530 vdd.n1175 gnd 0.009621f
C3531 vdd.n1176 gnd 0.009621f
C3532 vdd.n1177 gnd 0.009621f
C3533 vdd.n1178 gnd 0.006466f
C3534 vdd.t207 gnd 0.118362f
C3535 vdd.t206 gnd 0.126496f
C3536 vdd.t205 gnd 0.154579f
C3537 vdd.n1179 gnd 0.198149f
C3538 vdd.n1180 gnd 0.166481f
C3539 vdd.n1182 gnd 0.009621f
C3540 vdd.n1183 gnd 0.009621f
C3541 vdd.n1184 gnd 0.007744f
C3542 vdd.n1185 gnd 0.009621f
C3543 vdd.n1187 gnd 0.009621f
C3544 vdd.n1188 gnd 0.009621f
C3545 vdd.n1189 gnd 0.009621f
C3546 vdd.n1190 gnd 0.009621f
C3547 vdd.n1191 gnd 0.007744f
C3548 vdd.n1193 gnd 0.009621f
C3549 vdd.n1194 gnd 0.009621f
C3550 vdd.n1195 gnd 0.009621f
C3551 vdd.n1196 gnd 0.009621f
C3552 vdd.n1197 gnd 0.009621f
C3553 vdd.n1198 gnd 0.007744f
C3554 vdd.n1200 gnd 0.009621f
C3555 vdd.n1201 gnd 0.009621f
C3556 vdd.n1202 gnd 0.009621f
C3557 vdd.n1203 gnd 0.009621f
C3558 vdd.n1204 gnd 0.009621f
C3559 vdd.n1205 gnd 0.007744f
C3560 vdd.n1207 gnd 0.009621f
C3561 vdd.n1208 gnd 0.009621f
C3562 vdd.n1209 gnd 0.009621f
C3563 vdd.n1210 gnd 0.009621f
C3564 vdd.n1211 gnd 0.009621f
C3565 vdd.n1212 gnd 0.007744f
C3566 vdd.n1214 gnd 0.009621f
C3567 vdd.n1215 gnd 0.009621f
C3568 vdd.n1216 gnd 0.009621f
C3569 vdd.n1217 gnd 0.009621f
C3570 vdd.n1218 gnd 0.007666f
C3571 vdd.t204 gnd 0.118362f
C3572 vdd.t203 gnd 0.126496f
C3573 vdd.t201 gnd 0.154579f
C3574 vdd.n1219 gnd 0.198149f
C3575 vdd.n1220 gnd 0.166481f
C3576 vdd.n1222 gnd 0.009621f
C3577 vdd.n1223 gnd 0.009621f
C3578 vdd.n1224 gnd 0.007744f
C3579 vdd.n1225 gnd 0.009621f
C3580 vdd.n1227 gnd 0.009621f
C3581 vdd.n1228 gnd 0.009621f
C3582 vdd.n1229 gnd 0.009621f
C3583 vdd.n1230 gnd 0.009621f
C3584 vdd.n1231 gnd 0.007744f
C3585 vdd.n1233 gnd 0.009621f
C3586 vdd.n1234 gnd 0.009621f
C3587 vdd.n1235 gnd 0.009621f
C3588 vdd.n1236 gnd 0.009621f
C3589 vdd.n1237 gnd 0.009621f
C3590 vdd.n1238 gnd 0.007744f
C3591 vdd.n1240 gnd 0.009621f
C3592 vdd.n1241 gnd 0.009621f
C3593 vdd.n1242 gnd 0.009621f
C3594 vdd.n1243 gnd 0.009621f
C3595 vdd.n1244 gnd 0.009621f
C3596 vdd.n1245 gnd 0.007744f
C3597 vdd.n1247 gnd 0.009621f
C3598 vdd.n1248 gnd 0.009621f
C3599 vdd.n1249 gnd 0.006157f
C3600 vdd.n1250 gnd 0.007744f
C3601 vdd.n1251 gnd 0.014855f
C3602 vdd.n1252 gnd 0.014855f
C3603 vdd.n1253 gnd 0.006542f
C3604 vdd.n1254 gnd 0.006542f
C3605 vdd.n1255 gnd 0.006542f
C3606 vdd.n1256 gnd 0.006542f
C3607 vdd.n1257 gnd 0.006542f
C3608 vdd.n1258 gnd 0.006542f
C3609 vdd.n1259 gnd 0.006542f
C3610 vdd.n1260 gnd 0.006542f
C3611 vdd.n1261 gnd 0.006542f
C3612 vdd.n1262 gnd 0.006542f
C3613 vdd.n1263 gnd 0.006542f
C3614 vdd.n1264 gnd 0.006542f
C3615 vdd.n1265 gnd 0.006542f
C3616 vdd.n1266 gnd 0.006542f
C3617 vdd.n1267 gnd 0.006542f
C3618 vdd.n1268 gnd 0.006542f
C3619 vdd.n1269 gnd 0.006542f
C3620 vdd.n1270 gnd 0.006542f
C3621 vdd.n1271 gnd 0.006542f
C3622 vdd.n1272 gnd 0.006542f
C3623 vdd.n1273 gnd 0.006542f
C3624 vdd.n1274 gnd 0.006542f
C3625 vdd.n1275 gnd 0.006542f
C3626 vdd.n1276 gnd 0.006542f
C3627 vdd.n1277 gnd 0.006542f
C3628 vdd.n1278 gnd 0.006542f
C3629 vdd.n1279 gnd 0.006542f
C3630 vdd.n1280 gnd 0.006542f
C3631 vdd.n1281 gnd 0.006542f
C3632 vdd.n1282 gnd 0.006542f
C3633 vdd.n1283 gnd 0.006542f
C3634 vdd.n1284 gnd 0.006542f
C3635 vdd.n1285 gnd 0.006542f
C3636 vdd.t199 gnd 0.264369f
C3637 vdd.t200 gnd 0.270614f
C3638 vdd.t197 gnd 0.17259f
C3639 vdd.n1286 gnd 0.093276f
C3640 vdd.n1287 gnd 0.052909f
C3641 vdd.n1288 gnd 0.00935f
C3642 vdd.n1289 gnd 0.006542f
C3643 vdd.t233 gnd 0.264369f
C3644 vdd.t234 gnd 0.270614f
C3645 vdd.t232 gnd 0.17259f
C3646 vdd.n1290 gnd 0.093276f
C3647 vdd.n1291 gnd 0.052909f
C3648 vdd.n1292 gnd 0.006542f
C3649 vdd.n1293 gnd 0.006542f
C3650 vdd.n1294 gnd 0.006542f
C3651 vdd.n1295 gnd 0.006542f
C3652 vdd.n1296 gnd 0.006542f
C3653 vdd.n1297 gnd 0.006542f
C3654 vdd.n1298 gnd 0.006542f
C3655 vdd.n1299 gnd 0.006542f
C3656 vdd.n1300 gnd 0.006542f
C3657 vdd.n1301 gnd 0.006542f
C3658 vdd.n1302 gnd 0.006542f
C3659 vdd.n1303 gnd 0.006542f
C3660 vdd.n1304 gnd 0.006542f
C3661 vdd.n1305 gnd 0.006542f
C3662 vdd.n1306 gnd 0.006542f
C3663 vdd.n1307 gnd 0.006542f
C3664 vdd.n1308 gnd 0.006542f
C3665 vdd.n1309 gnd 0.006542f
C3666 vdd.n1310 gnd 0.006542f
C3667 vdd.n1311 gnd 0.006542f
C3668 vdd.n1312 gnd 0.006542f
C3669 vdd.n1313 gnd 0.006542f
C3670 vdd.n1314 gnd 0.006542f
C3671 vdd.n1315 gnd 0.006542f
C3672 vdd.n1316 gnd 0.006542f
C3673 vdd.n1317 gnd 0.006542f
C3674 vdd.n1318 gnd 0.004762f
C3675 vdd.n1319 gnd 0.00935f
C3676 vdd.n1320 gnd 0.005051f
C3677 vdd.n1321 gnd 0.006542f
C3678 vdd.n1322 gnd 0.006542f
C3679 vdd.n1323 gnd 0.006542f
C3680 vdd.n1324 gnd 0.014855f
C3681 vdd.n1325 gnd 0.014855f
C3682 vdd.n1326 gnd 0.014008f
C3683 vdd.n1327 gnd 0.014008f
C3684 vdd.n1328 gnd 0.006542f
C3685 vdd.n1329 gnd 0.006542f
C3686 vdd.n1330 gnd 0.006542f
C3687 vdd.n1331 gnd 0.006542f
C3688 vdd.n1332 gnd 0.006542f
C3689 vdd.n1333 gnd 0.006542f
C3690 vdd.n1334 gnd 0.006542f
C3691 vdd.n1335 gnd 0.006542f
C3692 vdd.n1336 gnd 0.006542f
C3693 vdd.n1337 gnd 0.006542f
C3694 vdd.n1338 gnd 0.006542f
C3695 vdd.n1339 gnd 0.006542f
C3696 vdd.n1340 gnd 0.006542f
C3697 vdd.n1341 gnd 0.006542f
C3698 vdd.n1342 gnd 0.006542f
C3699 vdd.n1343 gnd 0.006542f
C3700 vdd.n1344 gnd 0.006542f
C3701 vdd.n1345 gnd 0.006542f
C3702 vdd.n1346 gnd 0.006542f
C3703 vdd.n1347 gnd 0.006542f
C3704 vdd.n1348 gnd 0.006542f
C3705 vdd.n1349 gnd 0.006542f
C3706 vdd.n1350 gnd 0.006542f
C3707 vdd.n1351 gnd 0.006542f
C3708 vdd.n1352 gnd 0.006542f
C3709 vdd.n1353 gnd 0.006542f
C3710 vdd.n1354 gnd 0.006542f
C3711 vdd.n1355 gnd 0.006542f
C3712 vdd.n1356 gnd 0.006542f
C3713 vdd.n1357 gnd 0.006542f
C3714 vdd.n1358 gnd 0.006542f
C3715 vdd.n1359 gnd 0.006542f
C3716 vdd.n1360 gnd 0.006542f
C3717 vdd.n1361 gnd 0.006542f
C3718 vdd.n1362 gnd 0.006542f
C3719 vdd.n1363 gnd 0.006542f
C3720 vdd.n1364 gnd 0.006542f
C3721 vdd.n1365 gnd 0.006542f
C3722 vdd.n1366 gnd 0.006542f
C3723 vdd.n1367 gnd 0.006542f
C3724 vdd.n1368 gnd 0.006542f
C3725 vdd.n1369 gnd 0.006542f
C3726 vdd.n1370 gnd 0.398199f
C3727 vdd.n1371 gnd 0.006542f
C3728 vdd.n1372 gnd 0.006542f
C3729 vdd.n1373 gnd 0.006542f
C3730 vdd.n1374 gnd 0.006542f
C3731 vdd.n1375 gnd 0.006542f
C3732 vdd.n1376 gnd 0.006542f
C3733 vdd.n1377 gnd 0.006542f
C3734 vdd.n1378 gnd 0.006542f
C3735 vdd.n1379 gnd 0.006542f
C3736 vdd.n1380 gnd 0.006542f
C3737 vdd.n1381 gnd 0.006542f
C3738 vdd.n1382 gnd 0.006542f
C3739 vdd.n1383 gnd 0.006542f
C3740 vdd.n1384 gnd 0.006542f
C3741 vdd.n1385 gnd 0.006542f
C3742 vdd.n1386 gnd 0.006542f
C3743 vdd.n1387 gnd 0.006542f
C3744 vdd.n1388 gnd 0.006542f
C3745 vdd.n1389 gnd 0.006542f
C3746 vdd.n1390 gnd 0.006542f
C3747 vdd.n1391 gnd 0.006542f
C3748 vdd.n1392 gnd 0.006542f
C3749 vdd.n1393 gnd 0.006542f
C3750 vdd.n1394 gnd 0.006542f
C3751 vdd.n1395 gnd 0.006542f
C3752 vdd.n1396 gnd 0.604672f
C3753 vdd.n1397 gnd 0.006542f
C3754 vdd.n1398 gnd 0.006542f
C3755 vdd.n1399 gnd 0.006542f
C3756 vdd.n1400 gnd 0.006542f
C3757 vdd.n1401 gnd 0.006542f
C3758 vdd.n1402 gnd 0.006542f
C3759 vdd.n1403 gnd 0.006542f
C3760 vdd.n1404 gnd 0.006542f
C3761 vdd.n1405 gnd 0.006542f
C3762 vdd.n1406 gnd 0.006542f
C3763 vdd.n1407 gnd 0.006542f
C3764 vdd.n1408 gnd 0.211389f
C3765 vdd.n1409 gnd 0.006542f
C3766 vdd.n1410 gnd 0.006542f
C3767 vdd.n1411 gnd 0.006542f
C3768 vdd.n1412 gnd 0.006542f
C3769 vdd.n1413 gnd 0.006542f
C3770 vdd.n1414 gnd 0.006542f
C3771 vdd.n1415 gnd 0.006542f
C3772 vdd.n1416 gnd 0.006542f
C3773 vdd.n1417 gnd 0.006542f
C3774 vdd.n1418 gnd 0.006542f
C3775 vdd.n1419 gnd 0.006542f
C3776 vdd.n1420 gnd 0.006542f
C3777 vdd.n1421 gnd 0.006542f
C3778 vdd.n1422 gnd 0.006542f
C3779 vdd.n1423 gnd 0.006542f
C3780 vdd.n1424 gnd 0.006542f
C3781 vdd.n1425 gnd 0.006542f
C3782 vdd.n1426 gnd 0.006542f
C3783 vdd.n1427 gnd 0.006542f
C3784 vdd.n1428 gnd 0.006542f
C3785 vdd.n1429 gnd 0.006542f
C3786 vdd.n1430 gnd 0.006542f
C3787 vdd.n1431 gnd 0.006542f
C3788 vdd.n1432 gnd 0.006542f
C3789 vdd.n1433 gnd 0.006542f
C3790 vdd.n1434 gnd 0.006542f
C3791 vdd.n1435 gnd 0.006542f
C3792 vdd.n1436 gnd 0.006542f
C3793 vdd.n1437 gnd 0.006542f
C3794 vdd.n1438 gnd 0.006542f
C3795 vdd.n1439 gnd 0.006542f
C3796 vdd.n1440 gnd 0.006542f
C3797 vdd.n1441 gnd 0.006542f
C3798 vdd.n1442 gnd 0.006542f
C3799 vdd.n1443 gnd 0.006542f
C3800 vdd.n1444 gnd 0.006542f
C3801 vdd.n1445 gnd 0.006542f
C3802 vdd.n1446 gnd 0.006542f
C3803 vdd.n1447 gnd 0.006542f
C3804 vdd.n1448 gnd 0.006542f
C3805 vdd.n1449 gnd 0.006542f
C3806 vdd.n1450 gnd 0.006542f
C3807 vdd.n1451 gnd 0.014008f
C3808 vdd.n1452 gnd 0.014008f
C3809 vdd.n1453 gnd 0.014855f
C3810 vdd.n1454 gnd 0.006542f
C3811 vdd.n1455 gnd 0.006542f
C3812 vdd.n1456 gnd 0.005051f
C3813 vdd.n1457 gnd 0.006542f
C3814 vdd.n1458 gnd 0.006542f
C3815 vdd.n1459 gnd 0.004762f
C3816 vdd.n1460 gnd 0.006542f
C3817 vdd.n1461 gnd 0.006542f
C3818 vdd.n1462 gnd 0.006542f
C3819 vdd.n1463 gnd 0.006542f
C3820 vdd.n1464 gnd 0.006542f
C3821 vdd.n1465 gnd 0.006542f
C3822 vdd.n1466 gnd 0.006542f
C3823 vdd.n1467 gnd 0.006542f
C3824 vdd.n1468 gnd 0.006542f
C3825 vdd.n1469 gnd 0.006542f
C3826 vdd.n1470 gnd 0.006542f
C3827 vdd.n1471 gnd 0.006542f
C3828 vdd.n1472 gnd 0.006542f
C3829 vdd.n1473 gnd 0.006542f
C3830 vdd.n1474 gnd 0.006542f
C3831 vdd.n1475 gnd 0.006542f
C3832 vdd.n1476 gnd 0.006542f
C3833 vdd.n1477 gnd 0.006542f
C3834 vdd.n1478 gnd 0.006542f
C3835 vdd.n1479 gnd 0.006542f
C3836 vdd.n1480 gnd 0.006542f
C3837 vdd.n1481 gnd 0.006542f
C3838 vdd.n1482 gnd 0.006542f
C3839 vdd.n1483 gnd 0.006542f
C3840 vdd.n1484 gnd 0.006542f
C3841 vdd.n1485 gnd 0.006542f
C3842 vdd.n1486 gnd 0.044072f
C3843 vdd.n1488 gnd 0.022059f
C3844 vdd.n1489 gnd 0.007744f
C3845 vdd.n1491 gnd 0.009621f
C3846 vdd.n1492 gnd 0.007744f
C3847 vdd.n1493 gnd 0.009621f
C3848 vdd.n1495 gnd 0.009621f
C3849 vdd.n1496 gnd 0.009621f
C3850 vdd.n1498 gnd 0.009621f
C3851 vdd.n1499 gnd 0.006427f
C3852 vdd.n1500 gnd 0.54568f
C3853 vdd.n1501 gnd 0.009621f
C3854 vdd.n1502 gnd 0.022059f
C3855 vdd.n1503 gnd 0.007744f
C3856 vdd.n1504 gnd 0.009621f
C3857 vdd.n1505 gnd 0.007744f
C3858 vdd.n1506 gnd 0.009621f
C3859 vdd.n1507 gnd 0.983206f
C3860 vdd.n1508 gnd 0.009621f
C3861 vdd.n1509 gnd 0.007744f
C3862 vdd.n1510 gnd 0.007744f
C3863 vdd.n1511 gnd 0.009621f
C3864 vdd.n1512 gnd 0.007744f
C3865 vdd.n1513 gnd 0.009621f
C3866 vdd.t68 gnd 0.491603f
C3867 vdd.n1514 gnd 0.009621f
C3868 vdd.n1515 gnd 0.007744f
C3869 vdd.n1516 gnd 0.009621f
C3870 vdd.n1517 gnd 0.007744f
C3871 vdd.n1518 gnd 0.009621f
C3872 vdd.t136 gnd 0.491603f
C3873 vdd.n1519 gnd 0.009621f
C3874 vdd.n1520 gnd 0.007744f
C3875 vdd.n1521 gnd 0.009621f
C3876 vdd.n1522 gnd 0.007744f
C3877 vdd.n1523 gnd 0.009621f
C3878 vdd.t140 gnd 0.491603f
C3879 vdd.n1524 gnd 0.683328f
C3880 vdd.n1525 gnd 0.009621f
C3881 vdd.n1526 gnd 0.007744f
C3882 vdd.n1527 gnd 0.009621f
C3883 vdd.n1528 gnd 0.007744f
C3884 vdd.n1529 gnd 0.009621f
C3885 vdd.n1530 gnd 0.781649f
C3886 vdd.n1531 gnd 0.009621f
C3887 vdd.n1532 gnd 0.007744f
C3888 vdd.n1533 gnd 0.009621f
C3889 vdd.n1534 gnd 0.007744f
C3890 vdd.n1535 gnd 0.009621f
C3891 vdd.n1536 gnd 0.614504f
C3892 vdd.t94 gnd 0.491603f
C3893 vdd.n1537 gnd 0.009621f
C3894 vdd.n1538 gnd 0.007744f
C3895 vdd.n1539 gnd 0.009621f
C3896 vdd.n1540 gnd 0.007744f
C3897 vdd.n1541 gnd 0.009621f
C3898 vdd.t66 gnd 0.491603f
C3899 vdd.n1542 gnd 0.009621f
C3900 vdd.n1543 gnd 0.007744f
C3901 vdd.n1544 gnd 0.009621f
C3902 vdd.n1545 gnd 0.007744f
C3903 vdd.n1546 gnd 0.009621f
C3904 vdd.t74 gnd 0.491603f
C3905 vdd.n1547 gnd 0.535848f
C3906 vdd.n1548 gnd 0.009621f
C3907 vdd.n1549 gnd 0.007744f
C3908 vdd.n1550 gnd 0.009621f
C3909 vdd.n1551 gnd 0.007744f
C3910 vdd.n1552 gnd 0.009621f
C3911 vdd.t109 gnd 0.491603f
C3912 vdd.n1553 gnd 0.009621f
C3913 vdd.n1554 gnd 0.007744f
C3914 vdd.n1555 gnd 0.009621f
C3915 vdd.n1556 gnd 0.007744f
C3916 vdd.n1557 gnd 0.009621f
C3917 vdd.n1558 gnd 0.761985f
C3918 vdd.n1559 gnd 0.816061f
C3919 vdd.t134 gnd 0.491603f
C3920 vdd.n1560 gnd 0.009621f
C3921 vdd.n1561 gnd 0.007744f
C3922 vdd.n1562 gnd 0.009621f
C3923 vdd.n1563 gnd 0.007744f
C3924 vdd.n1564 gnd 0.009621f
C3925 vdd.n1565 gnd 0.59484f
C3926 vdd.n1566 gnd 0.009621f
C3927 vdd.n1567 gnd 0.007744f
C3928 vdd.n1568 gnd 0.009621f
C3929 vdd.n1569 gnd 0.007744f
C3930 vdd.n1570 gnd 0.009621f
C3931 vdd.t152 gnd 0.491603f
C3932 vdd.t72 gnd 0.491603f
C3933 vdd.n1571 gnd 0.009621f
C3934 vdd.n1572 gnd 0.007744f
C3935 vdd.n1573 gnd 0.009621f
C3936 vdd.n1574 gnd 0.007744f
C3937 vdd.n1575 gnd 0.009621f
C3938 vdd.t124 gnd 0.491603f
C3939 vdd.n1576 gnd 0.009621f
C3940 vdd.n1577 gnd 0.007744f
C3941 vdd.n1578 gnd 0.009621f
C3942 vdd.n1579 gnd 0.007744f
C3943 vdd.n1580 gnd 0.009621f
C3944 vdd.t101 gnd 0.491603f
C3945 vdd.n1581 gnd 0.722657f
C3946 vdd.n1582 gnd 0.009621f
C3947 vdd.n1583 gnd 0.007744f
C3948 vdd.n1584 gnd 0.009621f
C3949 vdd.n1585 gnd 0.007744f
C3950 vdd.n1586 gnd 0.009621f
C3951 vdd.n1587 gnd 0.983206f
C3952 vdd.n1588 gnd 0.009621f
C3953 vdd.n1589 gnd 0.007744f
C3954 vdd.n1590 gnd 0.009621f
C3955 vdd.n1591 gnd 0.007744f
C3956 vdd.n1592 gnd 0.009621f
C3957 vdd.n1593 gnd 0.830809f
C3958 vdd.n1594 gnd 0.009621f
C3959 vdd.n1595 gnd 0.007744f
C3960 vdd.n1596 gnd 0.021909f
C3961 vdd.n1597 gnd 0.006427f
C3962 vdd.n1598 gnd 0.021909f
C3963 vdd.n1599 gnd 1.29783f
C3964 vdd.n1600 gnd 0.021909f
C3965 vdd.n1601 gnd 0.006427f
C3966 vdd.n1602 gnd 0.009621f
C3967 vdd.t240 gnd 0.118362f
C3968 vdd.t241 gnd 0.126496f
C3969 vdd.t238 gnd 0.154579f
C3970 vdd.n1603 gnd 0.198149f
C3971 vdd.n1604 gnd 0.167255f
C3972 vdd.n1605 gnd 0.0127f
C3973 vdd.n1606 gnd 0.009621f
C3974 vdd.n1637 gnd 0.009621f
C3975 vdd.n1638 gnd 0.009621f
C3976 vdd.n1639 gnd 0.022059f
C3977 vdd.n1640 gnd 0.007744f
C3978 vdd.n1641 gnd 0.009621f
C3979 vdd.n1642 gnd 0.009621f
C3980 vdd.n1643 gnd 0.009621f
C3981 vdd.n1644 gnd 0.009621f
C3982 vdd.n1645 gnd 0.007744f
C3983 vdd.n1646 gnd 0.009621f
C3984 vdd.n1647 gnd 0.009621f
C3985 vdd.n1648 gnd 0.009621f
C3986 vdd.n1649 gnd 0.009621f
C3987 vdd.n1650 gnd 0.009621f
C3988 vdd.n1651 gnd 0.007744f
C3989 vdd.n1652 gnd 0.009621f
C3990 vdd.n1653 gnd 0.009621f
C3991 vdd.n1654 gnd 0.009621f
C3992 vdd.n1655 gnd 0.009621f
C3993 vdd.n1656 gnd 0.009621f
C3994 vdd.n1657 gnd 0.007744f
C3995 vdd.n1658 gnd 0.009621f
C3996 vdd.n1659 gnd 0.009621f
C3997 vdd.n1660 gnd 0.009621f
C3998 vdd.n1661 gnd 0.009621f
C3999 vdd.n1662 gnd 0.009621f
C4000 vdd.n1663 gnd 0.006466f
C4001 vdd.n1664 gnd 0.009621f
C4002 vdd.n1665 gnd 0.009621f
C4003 vdd.n1666 gnd 0.009621f
C4004 vdd.n1667 gnd 0.007744f
C4005 vdd.n1668 gnd 0.009621f
C4006 vdd.n1669 gnd 0.009621f
C4007 vdd.n1670 gnd 0.009621f
C4008 vdd.n1671 gnd 0.009621f
C4009 vdd.n1672 gnd 0.009621f
C4010 vdd.n1673 gnd 0.007744f
C4011 vdd.n1674 gnd 0.009621f
C4012 vdd.n1675 gnd 0.009621f
C4013 vdd.n1676 gnd 0.009621f
C4014 vdd.n1677 gnd 0.009621f
C4015 vdd.n1678 gnd 0.009621f
C4016 vdd.n1679 gnd 0.007744f
C4017 vdd.n1680 gnd 0.009621f
C4018 vdd.n1681 gnd 0.009621f
C4019 vdd.n1682 gnd 0.009621f
C4020 vdd.n1683 gnd 0.009621f
C4021 vdd.n1684 gnd 0.009621f
C4022 vdd.n1685 gnd 0.007744f
C4023 vdd.n1686 gnd 0.009621f
C4024 vdd.n1687 gnd 0.009621f
C4025 vdd.n1688 gnd 0.009621f
C4026 vdd.n1689 gnd 0.009621f
C4027 vdd.n1690 gnd 0.009621f
C4028 vdd.n1691 gnd 0.007744f
C4029 vdd.n1692 gnd 0.009621f
C4030 vdd.n1693 gnd 0.009621f
C4031 vdd.n1694 gnd 0.009621f
C4032 vdd.n1695 gnd 0.009621f
C4033 vdd.n1696 gnd 0.007666f
C4034 vdd.n1697 gnd 0.009621f
C4035 vdd.n1698 gnd 0.009621f
C4036 vdd.n1699 gnd 0.009621f
C4037 vdd.n1700 gnd 0.009621f
C4038 vdd.n1701 gnd 0.009621f
C4039 vdd.n1702 gnd 0.007744f
C4040 vdd.n1703 gnd 0.009621f
C4041 vdd.n1704 gnd 0.009621f
C4042 vdd.n1705 gnd 0.009621f
C4043 vdd.n1706 gnd 0.009621f
C4044 vdd.n1707 gnd 0.009621f
C4045 vdd.n1708 gnd 0.007744f
C4046 vdd.n1709 gnd 0.009621f
C4047 vdd.n1710 gnd 0.009621f
C4048 vdd.n1711 gnd 0.009621f
C4049 vdd.n1712 gnd 0.009621f
C4050 vdd.n1713 gnd 0.009621f
C4051 vdd.n1714 gnd 0.007744f
C4052 vdd.n1715 gnd 0.009621f
C4053 vdd.n1716 gnd 0.009621f
C4054 vdd.n1717 gnd 0.009621f
C4055 vdd.n1718 gnd 0.009621f
C4056 vdd.n1719 gnd 0.009621f
C4057 vdd.n1720 gnd 0.007744f
C4058 vdd.n1721 gnd 0.009621f
C4059 vdd.n1722 gnd 0.009621f
C4060 vdd.n1723 gnd 0.009621f
C4061 vdd.n1724 gnd 0.009621f
C4062 vdd.n1725 gnd 0.009621f
C4063 vdd.n1726 gnd 0.004065f
C4064 vdd.n1727 gnd 0.009621f
C4065 vdd.n1728 gnd 0.007744f
C4066 vdd.n1729 gnd 0.007744f
C4067 vdd.n1730 gnd 0.007744f
C4068 vdd.n1731 gnd 0.009621f
C4069 vdd.n1732 gnd 0.009621f
C4070 vdd.n1733 gnd 0.009621f
C4071 vdd.n1734 gnd 0.007744f
C4072 vdd.n1735 gnd 0.007744f
C4073 vdd.n1736 gnd 0.007744f
C4074 vdd.n1737 gnd 0.009621f
C4075 vdd.n1738 gnd 0.009621f
C4076 vdd.n1739 gnd 0.009621f
C4077 vdd.n1740 gnd 0.007744f
C4078 vdd.n1741 gnd 0.007744f
C4079 vdd.n1742 gnd 0.007744f
C4080 vdd.n1743 gnd 0.009621f
C4081 vdd.n1744 gnd 0.009621f
C4082 vdd.n1745 gnd 0.009621f
C4083 vdd.n1746 gnd 0.007744f
C4084 vdd.n1747 gnd 0.007744f
C4085 vdd.n1748 gnd 0.007744f
C4086 vdd.n1749 gnd 0.009621f
C4087 vdd.n1750 gnd 0.009621f
C4088 vdd.n1751 gnd 0.009621f
C4089 vdd.n1752 gnd 0.007744f
C4090 vdd.n1753 gnd 0.007744f
C4091 vdd.n1754 gnd 0.007744f
C4092 vdd.n1755 gnd 0.009621f
C4093 vdd.n1756 gnd 0.009621f
C4094 vdd.n1757 gnd 0.009621f
C4095 vdd.n1758 gnd 0.009621f
C4096 vdd.t254 gnd 0.118362f
C4097 vdd.t255 gnd 0.126496f
C4098 vdd.t253 gnd 0.154579f
C4099 vdd.n1759 gnd 0.198149f
C4100 vdd.n1760 gnd 0.167255f
C4101 vdd.n1761 gnd 0.016571f
C4102 vdd.n1762 gnd 0.005266f
C4103 vdd.n1763 gnd 0.007744f
C4104 vdd.n1764 gnd 0.009621f
C4105 vdd.n1765 gnd 0.009621f
C4106 vdd.n1766 gnd 0.009621f
C4107 vdd.n1767 gnd 0.007744f
C4108 vdd.n1768 gnd 0.007744f
C4109 vdd.n1769 gnd 0.007744f
C4110 vdd.n1770 gnd 0.009621f
C4111 vdd.n1771 gnd 0.009621f
C4112 vdd.n1772 gnd 0.009621f
C4113 vdd.n1773 gnd 0.007744f
C4114 vdd.n1774 gnd 0.007744f
C4115 vdd.n1775 gnd 0.007744f
C4116 vdd.n1776 gnd 0.009621f
C4117 vdd.n1777 gnd 0.009621f
C4118 vdd.n1778 gnd 0.009621f
C4119 vdd.n1779 gnd 0.007744f
C4120 vdd.n1780 gnd 0.007744f
C4121 vdd.n1781 gnd 0.007744f
C4122 vdd.n1782 gnd 0.009621f
C4123 vdd.n1783 gnd 0.009621f
C4124 vdd.n1784 gnd 0.009621f
C4125 vdd.n1785 gnd 0.007744f
C4126 vdd.n1786 gnd 0.007744f
C4127 vdd.n1787 gnd 0.007744f
C4128 vdd.n1788 gnd 0.009621f
C4129 vdd.n1789 gnd 0.009621f
C4130 vdd.n1790 gnd 0.009621f
C4131 vdd.n1791 gnd 0.007744f
C4132 vdd.n1792 gnd 0.006466f
C4133 vdd.n1793 gnd 0.009621f
C4134 vdd.n1794 gnd 0.009621f
C4135 vdd.t264 gnd 0.118362f
C4136 vdd.t265 gnd 0.126496f
C4137 vdd.t263 gnd 0.154579f
C4138 vdd.n1795 gnd 0.198149f
C4139 vdd.n1796 gnd 0.167255f
C4140 vdd.n1797 gnd 0.016571f
C4141 vdd.n1798 gnd 0.009621f
C4142 vdd.n1799 gnd 0.009621f
C4143 vdd.n1800 gnd 0.009621f
C4144 vdd.n1801 gnd 0.007744f
C4145 vdd.n1802 gnd 0.007744f
C4146 vdd.n1803 gnd 0.007744f
C4147 vdd.n1804 gnd 0.009621f
C4148 vdd.n1805 gnd 0.009621f
C4149 vdd.n1806 gnd 0.009621f
C4150 vdd.n1807 gnd 0.007744f
C4151 vdd.n1808 gnd 0.007744f
C4152 vdd.n1809 gnd 0.007744f
C4153 vdd.n1810 gnd 0.009621f
C4154 vdd.n1811 gnd 0.009621f
C4155 vdd.n1812 gnd 0.009621f
C4156 vdd.n1813 gnd 0.007744f
C4157 vdd.n1814 gnd 0.007744f
C4158 vdd.n1815 gnd 0.007744f
C4159 vdd.n1816 gnd 0.009621f
C4160 vdd.n1817 gnd 0.009621f
C4161 vdd.n1818 gnd 0.009621f
C4162 vdd.n1819 gnd 0.007744f
C4163 vdd.n1820 gnd 0.007744f
C4164 vdd.n1821 gnd 0.007744f
C4165 vdd.n1822 gnd 0.009621f
C4166 vdd.n1823 gnd 0.009621f
C4167 vdd.n1824 gnd 0.009621f
C4168 vdd.n1825 gnd 0.007744f
C4169 vdd.n1826 gnd 0.006427f
C4170 vdd.n1827 gnd 0.022059f
C4171 vdd.n1829 gnd 2.17289f
C4172 vdd.n1830 gnd 0.022059f
C4173 vdd.n1831 gnd 0.003678f
C4174 vdd.n1832 gnd 0.022059f
C4175 vdd.n1833 gnd 0.021909f
C4176 vdd.n1834 gnd 0.009621f
C4177 vdd.n1835 gnd 0.007744f
C4178 vdd.n1836 gnd 0.009621f
C4179 vdd.t239 gnd 0.491603f
C4180 vdd.n1837 gnd 0.644f
C4181 vdd.n1838 gnd 0.009621f
C4182 vdd.n1839 gnd 0.007744f
C4183 vdd.n1840 gnd 0.009621f
C4184 vdd.n1841 gnd 0.009621f
C4185 vdd.n1842 gnd 0.009621f
C4186 vdd.n1843 gnd 0.007744f
C4187 vdd.n1844 gnd 0.009621f
C4188 vdd.n1845 gnd 0.983206f
C4189 vdd.n1846 gnd 0.009621f
C4190 vdd.n1847 gnd 0.007744f
C4191 vdd.n1848 gnd 0.009621f
C4192 vdd.n1849 gnd 0.009621f
C4193 vdd.n1850 gnd 0.009621f
C4194 vdd.n1851 gnd 0.007744f
C4195 vdd.n1852 gnd 0.009621f
C4196 vdd.n1853 gnd 0.816061f
C4197 vdd.t138 gnd 0.491603f
C4198 vdd.n1854 gnd 0.565344f
C4199 vdd.n1855 gnd 0.009621f
C4200 vdd.n1856 gnd 0.007744f
C4201 vdd.n1857 gnd 0.009621f
C4202 vdd.n1858 gnd 0.009621f
C4203 vdd.n1859 gnd 0.009621f
C4204 vdd.n1860 gnd 0.007744f
C4205 vdd.n1861 gnd 0.009621f
C4206 vdd.n1862 gnd 0.585008f
C4207 vdd.n1863 gnd 0.009621f
C4208 vdd.n1864 gnd 0.007744f
C4209 vdd.n1865 gnd 0.009621f
C4210 vdd.n1866 gnd 0.009621f
C4211 vdd.n1867 gnd 0.009621f
C4212 vdd.n1868 gnd 0.007744f
C4213 vdd.n1869 gnd 0.009621f
C4214 vdd.n1870 gnd 0.555512f
C4215 vdd.n1871 gnd 0.752153f
C4216 vdd.n1872 gnd 0.009621f
C4217 vdd.n1873 gnd 0.007744f
C4218 vdd.n1874 gnd 0.009621f
C4219 vdd.n1875 gnd 0.009621f
C4220 vdd.n1876 gnd 0.009621f
C4221 vdd.n1877 gnd 0.007744f
C4222 vdd.n1878 gnd 0.009621f
C4223 vdd.n1879 gnd 0.816061f
C4224 vdd.n1880 gnd 0.009621f
C4225 vdd.n1881 gnd 0.007744f
C4226 vdd.n1882 gnd 0.009621f
C4227 vdd.n1883 gnd 0.009621f
C4228 vdd.n1884 gnd 0.009621f
C4229 vdd.n1885 gnd 0.007744f
C4230 vdd.n1886 gnd 0.009621f
C4231 vdd.t64 gnd 0.491603f
C4232 vdd.n1887 gnd 0.712825f
C4233 vdd.n1888 gnd 0.009621f
C4234 vdd.n1889 gnd 0.007744f
C4235 vdd.n1890 gnd 0.009621f
C4236 vdd.n1891 gnd 0.009621f
C4237 vdd.n1892 gnd 0.009621f
C4238 vdd.n1893 gnd 0.007744f
C4239 vdd.n1894 gnd 0.009621f
C4240 vdd.n1895 gnd 0.54568f
C4241 vdd.n1896 gnd 0.009621f
C4242 vdd.n1897 gnd 0.007744f
C4243 vdd.n1898 gnd 0.009621f
C4244 vdd.n1899 gnd 0.009621f
C4245 vdd.n1900 gnd 0.009621f
C4246 vdd.n1901 gnd 0.007744f
C4247 vdd.n1902 gnd 0.009621f
C4248 vdd.n1903 gnd 0.702993f
C4249 vdd.n1904 gnd 0.604672f
C4250 vdd.n1905 gnd 0.009621f
C4251 vdd.n1906 gnd 0.007744f
C4252 vdd.n1907 gnd 0.007394f
C4253 vdd.n1908 gnd 0.00528f
C4254 vdd.n1909 gnd 0.0049f
C4255 vdd.n1910 gnd 0.00271f
C4256 vdd.n1911 gnd 0.006223f
C4257 vdd.n1912 gnd 0.002633f
C4258 vdd.n1913 gnd 0.002788f
C4259 vdd.n1914 gnd 0.0049f
C4260 vdd.n1915 gnd 0.002633f
C4261 vdd.n1916 gnd 0.006223f
C4262 vdd.n1917 gnd 0.002788f
C4263 vdd.n1918 gnd 0.0049f
C4264 vdd.n1919 gnd 0.002633f
C4265 vdd.n1920 gnd 0.004667f
C4266 vdd.n1921 gnd 0.004681f
C4267 vdd.t131 gnd 0.01337f
C4268 vdd.n1922 gnd 0.029747f
C4269 vdd.n1923 gnd 0.154813f
C4270 vdd.n1924 gnd 0.002633f
C4271 vdd.n1925 gnd 0.002788f
C4272 vdd.n1926 gnd 0.006223f
C4273 vdd.n1927 gnd 0.006223f
C4274 vdd.n1928 gnd 0.002788f
C4275 vdd.n1929 gnd 0.002633f
C4276 vdd.n1930 gnd 0.0049f
C4277 vdd.n1931 gnd 0.0049f
C4278 vdd.n1932 gnd 0.002633f
C4279 vdd.n1933 gnd 0.002788f
C4280 vdd.n1934 gnd 0.006223f
C4281 vdd.n1935 gnd 0.006223f
C4282 vdd.n1936 gnd 0.002788f
C4283 vdd.n1937 gnd 0.002633f
C4284 vdd.n1938 gnd 0.0049f
C4285 vdd.n1939 gnd 0.0049f
C4286 vdd.n1940 gnd 0.002633f
C4287 vdd.n1941 gnd 0.002788f
C4288 vdd.n1942 gnd 0.006223f
C4289 vdd.n1943 gnd 0.006223f
C4290 vdd.n1944 gnd 0.014713f
C4291 vdd.n1945 gnd 0.00271f
C4292 vdd.n1946 gnd 0.002633f
C4293 vdd.n1947 gnd 0.012664f
C4294 vdd.n1948 gnd 0.008841f
C4295 vdd.t172 gnd 0.030974f
C4296 vdd.t191 gnd 0.030974f
C4297 vdd.n1949 gnd 0.212878f
C4298 vdd.n1950 gnd 0.167396f
C4299 vdd.t156 gnd 0.030974f
C4300 vdd.t89 gnd 0.030974f
C4301 vdd.n1951 gnd 0.212878f
C4302 vdd.n1952 gnd 0.135088f
C4303 vdd.t142 gnd 0.030974f
C4304 vdd.t98 gnd 0.030974f
C4305 vdd.n1953 gnd 0.212878f
C4306 vdd.n1954 gnd 0.135088f
C4307 vdd.t181 gnd 0.030974f
C4308 vdd.t118 gnd 0.030974f
C4309 vdd.n1955 gnd 0.212878f
C4310 vdd.n1956 gnd 0.135088f
C4311 vdd.t162 gnd 0.030974f
C4312 vdd.t135 gnd 0.030974f
C4313 vdd.n1957 gnd 0.212878f
C4314 vdd.n1958 gnd 0.135088f
C4315 vdd.t174 gnd 0.030974f
C4316 vdd.t73 gnd 0.030974f
C4317 vdd.n1959 gnd 0.212878f
C4318 vdd.n1960 gnd 0.135088f
C4319 vdd.t188 gnd 0.030974f
C4320 vdd.t125 gnd 0.030974f
C4321 vdd.n1961 gnd 0.212878f
C4322 vdd.n1962 gnd 0.135088f
C4323 vdd.n1963 gnd 0.00528f
C4324 vdd.n1964 gnd 0.0049f
C4325 vdd.n1965 gnd 0.00271f
C4326 vdd.n1966 gnd 0.006223f
C4327 vdd.n1967 gnd 0.002633f
C4328 vdd.n1968 gnd 0.002788f
C4329 vdd.n1969 gnd 0.0049f
C4330 vdd.n1970 gnd 0.002633f
C4331 vdd.n1971 gnd 0.006223f
C4332 vdd.n1972 gnd 0.002788f
C4333 vdd.n1973 gnd 0.0049f
C4334 vdd.n1974 gnd 0.002633f
C4335 vdd.n1975 gnd 0.004667f
C4336 vdd.n1976 gnd 0.004681f
C4337 vdd.t147 gnd 0.01337f
C4338 vdd.n1977 gnd 0.029747f
C4339 vdd.n1978 gnd 0.154813f
C4340 vdd.n1979 gnd 0.002633f
C4341 vdd.n1980 gnd 0.002788f
C4342 vdd.n1981 gnd 0.006223f
C4343 vdd.n1982 gnd 0.006223f
C4344 vdd.n1983 gnd 0.002788f
C4345 vdd.n1984 gnd 0.002633f
C4346 vdd.n1985 gnd 0.0049f
C4347 vdd.n1986 gnd 0.0049f
C4348 vdd.n1987 gnd 0.002633f
C4349 vdd.n1988 gnd 0.002788f
C4350 vdd.n1989 gnd 0.006223f
C4351 vdd.n1990 gnd 0.006223f
C4352 vdd.n1991 gnd 0.002788f
C4353 vdd.n1992 gnd 0.002633f
C4354 vdd.n1993 gnd 0.0049f
C4355 vdd.n1994 gnd 0.0049f
C4356 vdd.n1995 gnd 0.002633f
C4357 vdd.n1996 gnd 0.002788f
C4358 vdd.n1997 gnd 0.006223f
C4359 vdd.n1998 gnd 0.006223f
C4360 vdd.n1999 gnd 0.014713f
C4361 vdd.n2000 gnd 0.00271f
C4362 vdd.n2001 gnd 0.002633f
C4363 vdd.n2002 gnd 0.012664f
C4364 vdd.n2003 gnd 0.008564f
C4365 vdd.n2004 gnd 0.100506f
C4366 vdd.n2005 gnd 0.00528f
C4367 vdd.n2006 gnd 0.0049f
C4368 vdd.n2007 gnd 0.00271f
C4369 vdd.n2008 gnd 0.006223f
C4370 vdd.n2009 gnd 0.002633f
C4371 vdd.n2010 gnd 0.002788f
C4372 vdd.n2011 gnd 0.0049f
C4373 vdd.n2012 gnd 0.002633f
C4374 vdd.n2013 gnd 0.006223f
C4375 vdd.n2014 gnd 0.002788f
C4376 vdd.n2015 gnd 0.0049f
C4377 vdd.n2016 gnd 0.002633f
C4378 vdd.n2017 gnd 0.004667f
C4379 vdd.n2018 gnd 0.004681f
C4380 vdd.t100 gnd 0.01337f
C4381 vdd.n2019 gnd 0.029747f
C4382 vdd.n2020 gnd 0.154813f
C4383 vdd.n2021 gnd 0.002633f
C4384 vdd.n2022 gnd 0.002788f
C4385 vdd.n2023 gnd 0.006223f
C4386 vdd.n2024 gnd 0.006223f
C4387 vdd.n2025 gnd 0.002788f
C4388 vdd.n2026 gnd 0.002633f
C4389 vdd.n2027 gnd 0.0049f
C4390 vdd.n2028 gnd 0.0049f
C4391 vdd.n2029 gnd 0.002633f
C4392 vdd.n2030 gnd 0.002788f
C4393 vdd.n2031 gnd 0.006223f
C4394 vdd.n2032 gnd 0.006223f
C4395 vdd.n2033 gnd 0.002788f
C4396 vdd.n2034 gnd 0.002633f
C4397 vdd.n2035 gnd 0.0049f
C4398 vdd.n2036 gnd 0.0049f
C4399 vdd.n2037 gnd 0.002633f
C4400 vdd.n2038 gnd 0.002788f
C4401 vdd.n2039 gnd 0.006223f
C4402 vdd.n2040 gnd 0.006223f
C4403 vdd.n2041 gnd 0.014713f
C4404 vdd.n2042 gnd 0.00271f
C4405 vdd.n2043 gnd 0.002633f
C4406 vdd.n2044 gnd 0.012664f
C4407 vdd.n2045 gnd 0.008841f
C4408 vdd.t141 gnd 0.030974f
C4409 vdd.t137 gnd 0.030974f
C4410 vdd.n2046 gnd 0.212878f
C4411 vdd.n2047 gnd 0.167396f
C4412 vdd.t95 gnd 0.030974f
C4413 vdd.t79 gnd 0.030974f
C4414 vdd.n2048 gnd 0.212878f
C4415 vdd.n2049 gnd 0.135088f
C4416 vdd.t67 gnd 0.030974f
C4417 vdd.t132 gnd 0.030974f
C4418 vdd.n2050 gnd 0.212878f
C4419 vdd.n2051 gnd 0.135088f
C4420 vdd.t110 gnd 0.030974f
C4421 vdd.t75 gnd 0.030974f
C4422 vdd.n2052 gnd 0.212878f
C4423 vdd.n2053 gnd 0.135088f
C4424 vdd.t65 gnd 0.030974f
C4425 vdd.t157 gnd 0.030974f
C4426 vdd.n2054 gnd 0.212878f
C4427 vdd.n2055 gnd 0.135088f
C4428 vdd.t153 gnd 0.030974f
C4429 vdd.t111 gnd 0.030974f
C4430 vdd.n2056 gnd 0.212878f
C4431 vdd.n2057 gnd 0.135088f
C4432 vdd.t102 gnd 0.030974f
C4433 vdd.t179 gnd 0.030974f
C4434 vdd.n2058 gnd 0.212878f
C4435 vdd.n2059 gnd 0.135088f
C4436 vdd.n2060 gnd 0.00528f
C4437 vdd.n2061 gnd 0.0049f
C4438 vdd.n2062 gnd 0.00271f
C4439 vdd.n2063 gnd 0.006223f
C4440 vdd.n2064 gnd 0.002633f
C4441 vdd.n2065 gnd 0.002788f
C4442 vdd.n2066 gnd 0.0049f
C4443 vdd.n2067 gnd 0.002633f
C4444 vdd.n2068 gnd 0.006223f
C4445 vdd.n2069 gnd 0.002788f
C4446 vdd.n2070 gnd 0.0049f
C4447 vdd.n2071 gnd 0.002633f
C4448 vdd.n2072 gnd 0.004667f
C4449 vdd.n2073 gnd 0.004681f
C4450 vdd.t139 gnd 0.01337f
C4451 vdd.n2074 gnd 0.029747f
C4452 vdd.n2075 gnd 0.154813f
C4453 vdd.n2076 gnd 0.002633f
C4454 vdd.n2077 gnd 0.002788f
C4455 vdd.n2078 gnd 0.006223f
C4456 vdd.n2079 gnd 0.006223f
C4457 vdd.n2080 gnd 0.002788f
C4458 vdd.n2081 gnd 0.002633f
C4459 vdd.n2082 gnd 0.0049f
C4460 vdd.n2083 gnd 0.0049f
C4461 vdd.n2084 gnd 0.002633f
C4462 vdd.n2085 gnd 0.002788f
C4463 vdd.n2086 gnd 0.006223f
C4464 vdd.n2087 gnd 0.006223f
C4465 vdd.n2088 gnd 0.002788f
C4466 vdd.n2089 gnd 0.002633f
C4467 vdd.n2090 gnd 0.0049f
C4468 vdd.n2091 gnd 0.0049f
C4469 vdd.n2092 gnd 0.002633f
C4470 vdd.n2093 gnd 0.002788f
C4471 vdd.n2094 gnd 0.006223f
C4472 vdd.n2095 gnd 0.006223f
C4473 vdd.n2096 gnd 0.014713f
C4474 vdd.n2097 gnd 0.00271f
C4475 vdd.n2098 gnd 0.002633f
C4476 vdd.n2099 gnd 0.012664f
C4477 vdd.n2100 gnd 0.008564f
C4478 vdd.n2101 gnd 0.059791f
C4479 vdd.n2102 gnd 0.215442f
C4480 vdd.n2103 gnd 0.00528f
C4481 vdd.n2104 gnd 0.0049f
C4482 vdd.n2105 gnd 0.00271f
C4483 vdd.n2106 gnd 0.006223f
C4484 vdd.n2107 gnd 0.002633f
C4485 vdd.n2108 gnd 0.002788f
C4486 vdd.n2109 gnd 0.0049f
C4487 vdd.n2110 gnd 0.002633f
C4488 vdd.n2111 gnd 0.006223f
C4489 vdd.n2112 gnd 0.002788f
C4490 vdd.n2113 gnd 0.0049f
C4491 vdd.n2114 gnd 0.002633f
C4492 vdd.n2115 gnd 0.004667f
C4493 vdd.n2116 gnd 0.004681f
C4494 vdd.t69 gnd 0.01337f
C4495 vdd.n2117 gnd 0.029747f
C4496 vdd.n2118 gnd 0.154813f
C4497 vdd.n2119 gnd 0.002633f
C4498 vdd.n2120 gnd 0.002788f
C4499 vdd.n2121 gnd 0.006223f
C4500 vdd.n2122 gnd 0.006223f
C4501 vdd.n2123 gnd 0.002788f
C4502 vdd.n2124 gnd 0.002633f
C4503 vdd.n2125 gnd 0.0049f
C4504 vdd.n2126 gnd 0.0049f
C4505 vdd.n2127 gnd 0.002633f
C4506 vdd.n2128 gnd 0.002788f
C4507 vdd.n2129 gnd 0.006223f
C4508 vdd.n2130 gnd 0.006223f
C4509 vdd.n2131 gnd 0.002788f
C4510 vdd.n2132 gnd 0.002633f
C4511 vdd.n2133 gnd 0.0049f
C4512 vdd.n2134 gnd 0.0049f
C4513 vdd.n2135 gnd 0.002633f
C4514 vdd.n2136 gnd 0.002788f
C4515 vdd.n2137 gnd 0.006223f
C4516 vdd.n2138 gnd 0.006223f
C4517 vdd.n2139 gnd 0.014713f
C4518 vdd.n2140 gnd 0.00271f
C4519 vdd.n2141 gnd 0.002633f
C4520 vdd.n2142 gnd 0.012664f
C4521 vdd.n2143 gnd 0.008841f
C4522 vdd.t150 gnd 0.030974f
C4523 vdd.t149 gnd 0.030974f
C4524 vdd.n2144 gnd 0.212878f
C4525 vdd.n2145 gnd 0.167396f
C4526 vdd.t114 gnd 0.030974f
C4527 vdd.t92 gnd 0.030974f
C4528 vdd.n2146 gnd 0.212878f
C4529 vdd.n2147 gnd 0.135088f
C4530 vdd.t90 gnd 0.030974f
C4531 vdd.t143 gnd 0.030974f
C4532 vdd.n2148 gnd 0.212878f
C4533 vdd.n2149 gnd 0.135088f
C4534 vdd.t126 gnd 0.030974f
C4535 vdd.t91 gnd 0.030974f
C4536 vdd.n2150 gnd 0.212878f
C4537 vdd.n2151 gnd 0.135088f
C4538 vdd.t86 gnd 0.030974f
C4539 vdd.t165 gnd 0.030974f
C4540 vdd.n2152 gnd 0.212878f
C4541 vdd.n2153 gnd 0.135088f
C4542 vdd.t164 gnd 0.030974f
C4543 vdd.t120 gnd 0.030974f
C4544 vdd.n2154 gnd 0.212878f
C4545 vdd.n2155 gnd 0.135088f
C4546 vdd.t115 gnd 0.030974f
C4547 vdd.t189 gnd 0.030974f
C4548 vdd.n2156 gnd 0.212878f
C4549 vdd.n2157 gnd 0.135088f
C4550 vdd.n2158 gnd 0.00528f
C4551 vdd.n2159 gnd 0.0049f
C4552 vdd.n2160 gnd 0.00271f
C4553 vdd.n2161 gnd 0.006223f
C4554 vdd.n2162 gnd 0.002633f
C4555 vdd.n2163 gnd 0.002788f
C4556 vdd.n2164 gnd 0.0049f
C4557 vdd.n2165 gnd 0.002633f
C4558 vdd.n2166 gnd 0.006223f
C4559 vdd.n2167 gnd 0.002788f
C4560 vdd.n2168 gnd 0.0049f
C4561 vdd.n2169 gnd 0.002633f
C4562 vdd.n2170 gnd 0.004667f
C4563 vdd.n2171 gnd 0.004681f
C4564 vdd.t148 gnd 0.01337f
C4565 vdd.n2172 gnd 0.029747f
C4566 vdd.n2173 gnd 0.154813f
C4567 vdd.n2174 gnd 0.002633f
C4568 vdd.n2175 gnd 0.002788f
C4569 vdd.n2176 gnd 0.006223f
C4570 vdd.n2177 gnd 0.006223f
C4571 vdd.n2178 gnd 0.002788f
C4572 vdd.n2179 gnd 0.002633f
C4573 vdd.n2180 gnd 0.0049f
C4574 vdd.n2181 gnd 0.0049f
C4575 vdd.n2182 gnd 0.002633f
C4576 vdd.n2183 gnd 0.002788f
C4577 vdd.n2184 gnd 0.006223f
C4578 vdd.n2185 gnd 0.006223f
C4579 vdd.n2186 gnd 0.002788f
C4580 vdd.n2187 gnd 0.002633f
C4581 vdd.n2188 gnd 0.0049f
C4582 vdd.n2189 gnd 0.0049f
C4583 vdd.n2190 gnd 0.002633f
C4584 vdd.n2191 gnd 0.002788f
C4585 vdd.n2192 gnd 0.006223f
C4586 vdd.n2193 gnd 0.006223f
C4587 vdd.n2194 gnd 0.014713f
C4588 vdd.n2195 gnd 0.00271f
C4589 vdd.n2196 gnd 0.002633f
C4590 vdd.n2197 gnd 0.012664f
C4591 vdd.n2198 gnd 0.008564f
C4592 vdd.n2199 gnd 0.059791f
C4593 vdd.n2200 gnd 0.241267f
C4594 vdd.n2201 gnd 2.6504f
C4595 vdd.n2202 gnd 0.567475f
C4596 vdd.n2203 gnd 0.007394f
C4597 vdd.n2204 gnd 0.009621f
C4598 vdd.n2205 gnd 0.007744f
C4599 vdd.n2206 gnd 0.009621f
C4600 vdd.n2207 gnd 0.771817f
C4601 vdd.n2208 gnd 0.009621f
C4602 vdd.n2209 gnd 0.007744f
C4603 vdd.n2210 gnd 0.009621f
C4604 vdd.n2211 gnd 0.009621f
C4605 vdd.n2212 gnd 0.009621f
C4606 vdd.n2213 gnd 0.007744f
C4607 vdd.n2214 gnd 0.009621f
C4608 vdd.t97 gnd 0.491603f
C4609 vdd.n2215 gnd 0.816061f
C4610 vdd.n2216 gnd 0.009621f
C4611 vdd.n2217 gnd 0.007744f
C4612 vdd.n2218 gnd 0.009621f
C4613 vdd.n2219 gnd 0.009621f
C4614 vdd.n2220 gnd 0.009621f
C4615 vdd.n2221 gnd 0.007744f
C4616 vdd.n2222 gnd 0.009621f
C4617 vdd.n2223 gnd 0.693161f
C4618 vdd.n2224 gnd 0.009621f
C4619 vdd.n2225 gnd 0.007744f
C4620 vdd.n2226 gnd 0.009621f
C4621 vdd.n2227 gnd 0.009621f
C4622 vdd.n2228 gnd 0.009621f
C4623 vdd.n2229 gnd 0.007744f
C4624 vdd.n2230 gnd 0.009621f
C4625 vdd.n2231 gnd 0.816061f
C4626 vdd.t78 gnd 0.491603f
C4627 vdd.n2232 gnd 0.526015f
C4628 vdd.n2233 gnd 0.009621f
C4629 vdd.n2234 gnd 0.007744f
C4630 vdd.n2235 gnd 0.009621f
C4631 vdd.n2236 gnd 0.009621f
C4632 vdd.n2237 gnd 0.009621f
C4633 vdd.n2238 gnd 0.007744f
C4634 vdd.n2239 gnd 0.009621f
C4635 vdd.n2240 gnd 0.624336f
C4636 vdd.n2241 gnd 0.009621f
C4637 vdd.n2242 gnd 0.007744f
C4638 vdd.n2243 gnd 0.009621f
C4639 vdd.n2244 gnd 0.009621f
C4640 vdd.n2245 gnd 0.009621f
C4641 vdd.n2246 gnd 0.007744f
C4642 vdd.n2247 gnd 0.009621f
C4643 vdd.n2248 gnd 0.516183f
C4644 vdd.n2249 gnd 0.791481f
C4645 vdd.n2250 gnd 0.009621f
C4646 vdd.n2251 gnd 0.007744f
C4647 vdd.n2252 gnd 0.009621f
C4648 vdd.n2253 gnd 0.009621f
C4649 vdd.n2254 gnd 0.009621f
C4650 vdd.n2255 gnd 0.007744f
C4651 vdd.n2256 gnd 0.009621f
C4652 vdd.n2257 gnd 0.958626f
C4653 vdd.n2258 gnd 0.009621f
C4654 vdd.n2259 gnd 0.007744f
C4655 vdd.n2260 gnd 0.009621f
C4656 vdd.n2261 gnd 0.009621f
C4657 vdd.n2262 gnd 0.021909f
C4658 vdd.n2263 gnd 0.009621f
C4659 vdd.n2264 gnd 0.009621f
C4660 vdd.n2265 gnd 0.007744f
C4661 vdd.n2266 gnd 0.009621f
C4662 vdd.t202 gnd 0.491603f
C4663 vdd.n2267 gnd 0.92913f
C4664 vdd.n2268 gnd 0.009621f
C4665 vdd.n2269 gnd 0.007744f
C4666 vdd.n2270 gnd 0.009621f
C4667 vdd.n2271 gnd 0.009621f
C4668 vdd.n2272 gnd 0.021909f
C4669 vdd.n2273 gnd 0.006427f
C4670 vdd.n2274 gnd 0.021909f
C4671 vdd.n2275 gnd 1.29783f
C4672 vdd.n2276 gnd 0.021909f
C4673 vdd.n2277 gnd 0.022059f
C4674 vdd.n2278 gnd 0.003678f
C4675 vdd.t225 gnd 0.118362f
C4676 vdd.t224 gnd 0.126496f
C4677 vdd.t223 gnd 0.154579f
C4678 vdd.n2279 gnd 0.198149f
C4679 vdd.n2280 gnd 0.166481f
C4680 vdd.n2281 gnd 0.011925f
C4681 vdd.n2282 gnd 0.004065f
C4682 vdd.n2283 gnd 0.008274f
C4683 vdd.n2284 gnd 1.02135f
C4684 vdd.n2286 gnd 0.007744f
C4685 vdd.n2287 gnd 0.007744f
C4686 vdd.n2288 gnd 0.009621f
C4687 vdd.n2290 gnd 0.009621f
C4688 vdd.n2291 gnd 0.009621f
C4689 vdd.n2292 gnd 0.007744f
C4690 vdd.n2293 gnd 0.007744f
C4691 vdd.n2294 gnd 0.007744f
C4692 vdd.n2295 gnd 0.009621f
C4693 vdd.n2297 gnd 0.009621f
C4694 vdd.n2298 gnd 0.009621f
C4695 vdd.n2299 gnd 0.007744f
C4696 vdd.n2300 gnd 0.007744f
C4697 vdd.n2301 gnd 0.007744f
C4698 vdd.n2302 gnd 0.009621f
C4699 vdd.n2304 gnd 0.009621f
C4700 vdd.n2305 gnd 0.009621f
C4701 vdd.n2306 gnd 0.007744f
C4702 vdd.n2307 gnd 0.007744f
C4703 vdd.n2308 gnd 0.007744f
C4704 vdd.n2309 gnd 0.009621f
C4705 vdd.n2311 gnd 0.009621f
C4706 vdd.n2312 gnd 0.009621f
C4707 vdd.n2313 gnd 0.007744f
C4708 vdd.n2314 gnd 0.009621f
C4709 vdd.n2315 gnd 0.009621f
C4710 vdd.n2316 gnd 0.009621f
C4711 vdd.n2317 gnd 0.015797f
C4712 vdd.n2318 gnd 0.005266f
C4713 vdd.n2319 gnd 0.007744f
C4714 vdd.n2320 gnd 0.009621f
C4715 vdd.n2322 gnd 0.009621f
C4716 vdd.n2323 gnd 0.009621f
C4717 vdd.n2324 gnd 0.007744f
C4718 vdd.n2325 gnd 0.007744f
C4719 vdd.n2326 gnd 0.007744f
C4720 vdd.n2327 gnd 0.009621f
C4721 vdd.n2329 gnd 0.009621f
C4722 vdd.n2330 gnd 0.009621f
C4723 vdd.n2331 gnd 0.007744f
C4724 vdd.n2332 gnd 0.007744f
C4725 vdd.n2333 gnd 0.007744f
C4726 vdd.n2334 gnd 0.009621f
C4727 vdd.n2336 gnd 0.009621f
C4728 vdd.n2337 gnd 0.009621f
C4729 vdd.n2338 gnd 0.007744f
C4730 vdd.n2339 gnd 0.007744f
C4731 vdd.n2340 gnd 0.007744f
C4732 vdd.n2341 gnd 0.009621f
C4733 vdd.n2343 gnd 0.009621f
C4734 vdd.n2344 gnd 0.009621f
C4735 vdd.n2345 gnd 0.007744f
C4736 vdd.n2346 gnd 0.007744f
C4737 vdd.n2347 gnd 0.007744f
C4738 vdd.n2348 gnd 0.009621f
C4739 vdd.n2350 gnd 0.009621f
C4740 vdd.n2351 gnd 0.009621f
C4741 vdd.n2352 gnd 0.007744f
C4742 vdd.n2353 gnd 0.009621f
C4743 vdd.n2354 gnd 0.009621f
C4744 vdd.n2355 gnd 0.009621f
C4745 vdd.n2356 gnd 0.015797f
C4746 vdd.n2357 gnd 0.006466f
C4747 vdd.n2358 gnd 0.007744f
C4748 vdd.n2359 gnd 0.009621f
C4749 vdd.n2361 gnd 0.009621f
C4750 vdd.n2362 gnd 0.009621f
C4751 vdd.n2363 gnd 0.007744f
C4752 vdd.n2364 gnd 0.007744f
C4753 vdd.n2365 gnd 0.007744f
C4754 vdd.n2366 gnd 0.009621f
C4755 vdd.n2368 gnd 0.009621f
C4756 vdd.n2369 gnd 0.009621f
C4757 vdd.n2370 gnd 0.007744f
C4758 vdd.n2371 gnd 0.007744f
C4759 vdd.n2372 gnd 0.007744f
C4760 vdd.n2373 gnd 0.009621f
C4761 vdd.n2375 gnd 0.009621f
C4762 vdd.n2376 gnd 0.009621f
C4763 vdd.n2377 gnd 0.007744f
C4764 vdd.n2378 gnd 0.007744f
C4765 vdd.n2379 gnd 0.007744f
C4766 vdd.n2380 gnd 0.009621f
C4767 vdd.n2382 gnd 0.009621f
C4768 vdd.n2383 gnd 0.007744f
C4769 vdd.n2384 gnd 0.007744f
C4770 vdd.n2385 gnd 0.009621f
C4771 vdd.n2387 gnd 0.009621f
C4772 vdd.n2388 gnd 0.009621f
C4773 vdd.n2389 gnd 0.007744f
C4774 vdd.n2390 gnd 0.008274f
C4775 vdd.n2391 gnd 1.02135f
C4776 vdd.n2392 gnd 0.044072f
C4777 vdd.n2393 gnd 0.006542f
C4778 vdd.n2394 gnd 0.006542f
C4779 vdd.n2395 gnd 0.006542f
C4780 vdd.n2396 gnd 0.006542f
C4781 vdd.n2397 gnd 0.006542f
C4782 vdd.n2398 gnd 0.006542f
C4783 vdd.n2399 gnd 0.006542f
C4784 vdd.n2400 gnd 0.006542f
C4785 vdd.n2401 gnd 0.006542f
C4786 vdd.n2402 gnd 0.006542f
C4787 vdd.n2403 gnd 0.006542f
C4788 vdd.n2404 gnd 0.006542f
C4789 vdd.n2405 gnd 0.006542f
C4790 vdd.n2406 gnd 0.006542f
C4791 vdd.n2407 gnd 0.006542f
C4792 vdd.n2408 gnd 0.006542f
C4793 vdd.n2409 gnd 0.006542f
C4794 vdd.n2410 gnd 0.006542f
C4795 vdd.n2411 gnd 0.006542f
C4796 vdd.n2412 gnd 0.006542f
C4797 vdd.n2413 gnd 0.006542f
C4798 vdd.n2414 gnd 0.006542f
C4799 vdd.n2415 gnd 0.006542f
C4800 vdd.n2416 gnd 0.006542f
C4801 vdd.n2417 gnd 0.006542f
C4802 vdd.n2418 gnd 0.006542f
C4803 vdd.n2419 gnd 0.006542f
C4804 vdd.n2420 gnd 0.006542f
C4805 vdd.n2421 gnd 0.006542f
C4806 vdd.n2422 gnd 0.006542f
C4807 vdd.n2423 gnd 11.6117f
C4808 vdd.n2425 gnd 0.014855f
C4809 vdd.n2426 gnd 0.014855f
C4810 vdd.n2427 gnd 0.014008f
C4811 vdd.n2428 gnd 0.006542f
C4812 vdd.n2429 gnd 0.006542f
C4813 vdd.n2430 gnd 0.66858f
C4814 vdd.n2431 gnd 0.006542f
C4815 vdd.n2432 gnd 0.006542f
C4816 vdd.n2433 gnd 0.006542f
C4817 vdd.n2434 gnd 0.006542f
C4818 vdd.n2435 gnd 0.006542f
C4819 vdd.n2436 gnd 0.526015f
C4820 vdd.n2437 gnd 0.006542f
C4821 vdd.n2438 gnd 0.006542f
C4822 vdd.n2439 gnd 0.006542f
C4823 vdd.n2440 gnd 0.006542f
C4824 vdd.n2441 gnd 0.006542f
C4825 vdd.n2442 gnd 0.66858f
C4826 vdd.n2443 gnd 0.006542f
C4827 vdd.n2444 gnd 0.006542f
C4828 vdd.n2445 gnd 0.006542f
C4829 vdd.n2446 gnd 0.006542f
C4830 vdd.n2447 gnd 0.006542f
C4831 vdd.n2448 gnd 0.66858f
C4832 vdd.n2449 gnd 0.006542f
C4833 vdd.n2450 gnd 0.006542f
C4834 vdd.n2451 gnd 0.006542f
C4835 vdd.n2452 gnd 0.006542f
C4836 vdd.n2453 gnd 0.006542f
C4837 vdd.n2454 gnd 0.644f
C4838 vdd.n2455 gnd 0.006542f
C4839 vdd.n2456 gnd 0.006542f
C4840 vdd.n2457 gnd 0.006542f
C4841 vdd.n2458 gnd 0.006542f
C4842 vdd.n2459 gnd 0.006542f
C4843 vdd.n2460 gnd 0.496519f
C4844 vdd.n2461 gnd 0.006542f
C4845 vdd.n2462 gnd 0.006542f
C4846 vdd.n2463 gnd 0.006542f
C4847 vdd.n2464 gnd 0.006542f
C4848 vdd.n2465 gnd 0.006542f
C4849 vdd.n2466 gnd 0.349038f
C4850 vdd.n2467 gnd 0.006542f
C4851 vdd.n2468 gnd 0.006542f
C4852 vdd.n2469 gnd 0.006542f
C4853 vdd.n2470 gnd 0.006542f
C4854 vdd.n2471 gnd 0.006542f
C4855 vdd.n2472 gnd 0.467023f
C4856 vdd.n2473 gnd 0.006542f
C4857 vdd.n2474 gnd 0.006542f
C4858 vdd.n2475 gnd 0.006542f
C4859 vdd.n2476 gnd 0.006542f
C4860 vdd.n2477 gnd 0.006542f
C4861 vdd.n2478 gnd 0.614504f
C4862 vdd.n2479 gnd 0.006542f
C4863 vdd.n2480 gnd 0.006542f
C4864 vdd.n2481 gnd 0.006542f
C4865 vdd.n2482 gnd 0.006542f
C4866 vdd.n2483 gnd 0.006542f
C4867 vdd.n2484 gnd 0.66858f
C4868 vdd.n2485 gnd 0.006542f
C4869 vdd.n2486 gnd 0.006542f
C4870 vdd.n2487 gnd 0.006542f
C4871 vdd.n2488 gnd 0.006542f
C4872 vdd.n2489 gnd 0.006542f
C4873 vdd.n2490 gnd 0.575176f
C4874 vdd.n2491 gnd 0.006542f
C4875 vdd.n2492 gnd 0.006542f
C4876 vdd.n2493 gnd 0.005195f
C4877 vdd.n2494 gnd 0.018952f
C4878 vdd.n2495 gnd 0.004618f
C4879 vdd.n2496 gnd 0.006542f
C4880 vdd.n2497 gnd 0.427695f
C4881 vdd.n2498 gnd 0.006542f
C4882 vdd.n2499 gnd 0.006542f
C4883 vdd.n2500 gnd 0.006542f
C4884 vdd.n2501 gnd 0.006542f
C4885 vdd.n2502 gnd 0.006542f
C4886 vdd.n2503 gnd 0.388367f
C4887 vdd.n2504 gnd 0.006542f
C4888 vdd.n2505 gnd 0.006542f
C4889 vdd.n2506 gnd 0.006542f
C4890 vdd.n2507 gnd 0.006542f
C4891 vdd.n2508 gnd 0.006542f
C4892 vdd.n2509 gnd 0.535848f
C4893 vdd.n2510 gnd 0.006542f
C4894 vdd.n2511 gnd 0.006542f
C4895 vdd.n2512 gnd 0.006542f
C4896 vdd.n2513 gnd 0.006542f
C4897 vdd.n2514 gnd 0.006542f
C4898 vdd.n2515 gnd 0.589924f
C4899 vdd.n2516 gnd 0.006542f
C4900 vdd.n2517 gnd 0.006542f
C4901 vdd.n2518 gnd 0.006542f
C4902 vdd.n2519 gnd 0.006542f
C4903 vdd.n2520 gnd 0.006542f
C4904 vdd.n2521 gnd 0.442443f
C4905 vdd.n2522 gnd 0.006542f
C4906 vdd.n2523 gnd 0.006542f
C4907 vdd.n2524 gnd 0.006542f
C4908 vdd.n2525 gnd 0.006542f
C4909 vdd.n2526 gnd 0.006542f
C4910 vdd.n2527 gnd 0.211389f
C4911 vdd.n2528 gnd 0.006542f
C4912 vdd.n2529 gnd 0.006542f
C4913 vdd.n2530 gnd 0.006542f
C4914 vdd.n2531 gnd 0.006542f
C4915 vdd.n2532 gnd 0.006542f
C4916 vdd.n2533 gnd 0.211389f
C4917 vdd.n2534 gnd 0.006542f
C4918 vdd.n2535 gnd 0.006542f
C4919 vdd.n2536 gnd 0.006542f
C4920 vdd.n2537 gnd 0.006542f
C4921 vdd.n2538 gnd 0.006542f
C4922 vdd.n2539 gnd 0.66858f
C4923 vdd.n2540 gnd 0.006542f
C4924 vdd.n2541 gnd 0.006542f
C4925 vdd.n2542 gnd 0.006542f
C4926 vdd.n2543 gnd 0.006542f
C4927 vdd.n2544 gnd 0.006542f
C4928 vdd.n2545 gnd 0.006542f
C4929 vdd.n2546 gnd 0.006542f
C4930 vdd.n2547 gnd 0.462107f
C4931 vdd.n2548 gnd 0.006542f
C4932 vdd.n2549 gnd 0.006542f
C4933 vdd.n2550 gnd 0.006542f
C4934 vdd.n2551 gnd 0.006542f
C4935 vdd.n2552 gnd 0.006542f
C4936 vdd.n2553 gnd 0.006542f
C4937 vdd.n2554 gnd 0.417863f
C4938 vdd.n2555 gnd 0.006542f
C4939 vdd.n2556 gnd 0.006542f
C4940 vdd.n2557 gnd 0.006542f
C4941 vdd.n2558 gnd 0.014855f
C4942 vdd.n2559 gnd 0.014008f
C4943 vdd.n2560 gnd 0.006542f
C4944 vdd.n2561 gnd 0.006542f
C4945 vdd.n2562 gnd 0.005051f
C4946 vdd.n2563 gnd 0.006542f
C4947 vdd.n2564 gnd 0.006542f
C4948 vdd.n2565 gnd 0.004762f
C4949 vdd.n2566 gnd 0.006542f
C4950 vdd.n2567 gnd 0.006542f
C4951 vdd.n2568 gnd 0.006542f
C4952 vdd.n2569 gnd 0.006542f
C4953 vdd.n2570 gnd 0.006542f
C4954 vdd.n2571 gnd 0.006542f
C4955 vdd.n2572 gnd 0.006542f
C4956 vdd.n2573 gnd 0.006542f
C4957 vdd.n2574 gnd 0.006542f
C4958 vdd.n2575 gnd 0.006542f
C4959 vdd.n2576 gnd 0.006542f
C4960 vdd.n2577 gnd 0.006542f
C4961 vdd.n2578 gnd 0.006542f
C4962 vdd.n2579 gnd 0.006542f
C4963 vdd.n2580 gnd 0.006542f
C4964 vdd.n2581 gnd 0.006542f
C4965 vdd.n2582 gnd 0.006542f
C4966 vdd.n2583 gnd 0.006542f
C4967 vdd.n2584 gnd 0.006542f
C4968 vdd.n2585 gnd 0.006542f
C4969 vdd.n2586 gnd 0.006542f
C4970 vdd.n2587 gnd 0.006542f
C4971 vdd.n2588 gnd 0.006542f
C4972 vdd.n2589 gnd 0.006542f
C4973 vdd.n2590 gnd 0.006542f
C4974 vdd.n2591 gnd 0.006542f
C4975 vdd.n2592 gnd 0.006542f
C4976 vdd.n2593 gnd 0.006542f
C4977 vdd.n2594 gnd 0.006542f
C4978 vdd.n2595 gnd 0.006542f
C4979 vdd.n2596 gnd 0.006542f
C4980 vdd.n2597 gnd 0.006542f
C4981 vdd.n2598 gnd 0.006542f
C4982 vdd.n2599 gnd 0.006542f
C4983 vdd.n2600 gnd 0.006542f
C4984 vdd.n2601 gnd 0.006542f
C4985 vdd.n2602 gnd 0.006542f
C4986 vdd.n2603 gnd 0.006542f
C4987 vdd.n2604 gnd 0.006542f
C4988 vdd.n2605 gnd 0.006542f
C4989 vdd.n2606 gnd 0.006542f
C4990 vdd.n2607 gnd 0.006542f
C4991 vdd.n2608 gnd 0.006542f
C4992 vdd.n2609 gnd 0.006542f
C4993 vdd.n2610 gnd 0.006542f
C4994 vdd.n2611 gnd 0.006542f
C4995 vdd.n2612 gnd 0.006542f
C4996 vdd.n2613 gnd 0.006542f
C4997 vdd.n2614 gnd 0.006542f
C4998 vdd.n2615 gnd 0.006542f
C4999 vdd.n2616 gnd 0.006542f
C5000 vdd.n2617 gnd 0.006542f
C5001 vdd.n2618 gnd 0.006542f
C5002 vdd.n2619 gnd 0.006542f
C5003 vdd.n2620 gnd 0.006542f
C5004 vdd.n2621 gnd 0.006542f
C5005 vdd.n2622 gnd 0.006542f
C5006 vdd.n2623 gnd 0.006542f
C5007 vdd.n2624 gnd 0.006542f
C5008 vdd.n2625 gnd 0.006542f
C5009 vdd.n2626 gnd 0.014855f
C5010 vdd.n2627 gnd 0.014008f
C5011 vdd.n2628 gnd 0.014008f
C5012 vdd.n2629 gnd 0.757069f
C5013 vdd.n2630 gnd 0.014008f
C5014 vdd.n2631 gnd 0.014855f
C5015 vdd.n2632 gnd 0.014008f
C5016 vdd.n2633 gnd 0.006542f
C5017 vdd.n2634 gnd 0.006542f
C5018 vdd.n2635 gnd 0.006542f
C5019 vdd.n2636 gnd 0.005051f
C5020 vdd.n2637 gnd 0.00935f
C5021 vdd.n2638 gnd 0.004762f
C5022 vdd.n2639 gnd 0.006542f
C5023 vdd.n2640 gnd 0.006542f
C5024 vdd.n2641 gnd 0.006542f
C5025 vdd.n2642 gnd 0.006542f
C5026 vdd.n2643 gnd 0.006542f
C5027 vdd.n2644 gnd 0.006542f
C5028 vdd.n2645 gnd 0.006542f
C5029 vdd.n2646 gnd 0.006542f
C5030 vdd.n2647 gnd 0.006542f
C5031 vdd.n2648 gnd 0.006542f
C5032 vdd.n2649 gnd 0.006542f
C5033 vdd.n2650 gnd 0.006542f
C5034 vdd.n2651 gnd 0.006542f
C5035 vdd.n2652 gnd 0.006542f
C5036 vdd.n2653 gnd 0.006542f
C5037 vdd.n2654 gnd 0.006542f
C5038 vdd.n2655 gnd 0.006542f
C5039 vdd.n2656 gnd 0.006542f
C5040 vdd.n2657 gnd 0.006542f
C5041 vdd.n2658 gnd 0.006542f
C5042 vdd.n2659 gnd 0.006542f
C5043 vdd.n2660 gnd 0.006542f
C5044 vdd.n2661 gnd 0.006542f
C5045 vdd.n2662 gnd 0.006542f
C5046 vdd.n2663 gnd 0.006542f
C5047 vdd.n2664 gnd 0.006542f
C5048 vdd.n2665 gnd 0.006542f
C5049 vdd.n2666 gnd 0.006542f
C5050 vdd.n2667 gnd 0.006542f
C5051 vdd.n2668 gnd 0.006542f
C5052 vdd.n2669 gnd 0.006542f
C5053 vdd.n2670 gnd 0.006542f
C5054 vdd.n2671 gnd 0.006542f
C5055 vdd.n2672 gnd 0.006542f
C5056 vdd.n2673 gnd 0.006542f
C5057 vdd.n2674 gnd 0.006542f
C5058 vdd.n2675 gnd 0.006542f
C5059 vdd.n2676 gnd 0.006542f
C5060 vdd.n2677 gnd 0.006542f
C5061 vdd.n2678 gnd 0.006542f
C5062 vdd.n2679 gnd 0.006542f
C5063 vdd.n2680 gnd 0.006542f
C5064 vdd.n2681 gnd 0.006542f
C5065 vdd.n2682 gnd 0.006542f
C5066 vdd.n2683 gnd 0.006542f
C5067 vdd.n2684 gnd 0.006542f
C5068 vdd.n2685 gnd 0.006542f
C5069 vdd.n2686 gnd 0.006542f
C5070 vdd.n2687 gnd 0.006542f
C5071 vdd.n2688 gnd 0.006542f
C5072 vdd.n2689 gnd 0.006542f
C5073 vdd.n2690 gnd 0.006542f
C5074 vdd.n2691 gnd 0.006542f
C5075 vdd.n2692 gnd 0.006542f
C5076 vdd.n2693 gnd 0.006542f
C5077 vdd.n2694 gnd 0.006542f
C5078 vdd.n2695 gnd 0.006542f
C5079 vdd.n2696 gnd 0.006542f
C5080 vdd.n2697 gnd 0.006542f
C5081 vdd.n2698 gnd 0.006542f
C5082 vdd.n2699 gnd 0.014855f
C5083 vdd.n2700 gnd 0.014855f
C5084 vdd.n2701 gnd 0.816061f
C5085 vdd.t30 gnd 2.90046f
C5086 vdd.t17 gnd 2.90046f
C5087 vdd.n2735 gnd 0.014855f
C5088 vdd.t35 gnd 0.57026f
C5089 vdd.n2736 gnd 0.006542f
C5090 vdd.t251 gnd 0.264369f
C5091 vdd.t252 gnd 0.270614f
C5092 vdd.t249 gnd 0.17259f
C5093 vdd.n2737 gnd 0.093276f
C5094 vdd.n2738 gnd 0.052909f
C5095 vdd.n2739 gnd 0.006542f
C5096 vdd.t261 gnd 0.264369f
C5097 vdd.t262 gnd 0.270614f
C5098 vdd.t260 gnd 0.17259f
C5099 vdd.n2740 gnd 0.093276f
C5100 vdd.n2741 gnd 0.052909f
C5101 vdd.n2742 gnd 0.00935f
C5102 vdd.n2743 gnd 0.014855f
C5103 vdd.n2744 gnd 0.014855f
C5104 vdd.n2745 gnd 0.006542f
C5105 vdd.n2746 gnd 0.006542f
C5106 vdd.n2747 gnd 0.006542f
C5107 vdd.n2748 gnd 0.006542f
C5108 vdd.n2749 gnd 0.006542f
C5109 vdd.n2750 gnd 0.006542f
C5110 vdd.n2751 gnd 0.006542f
C5111 vdd.n2752 gnd 0.006542f
C5112 vdd.n2753 gnd 0.006542f
C5113 vdd.n2754 gnd 0.006542f
C5114 vdd.n2755 gnd 0.006542f
C5115 vdd.n2756 gnd 0.006542f
C5116 vdd.n2757 gnd 0.006542f
C5117 vdd.n2758 gnd 0.006542f
C5118 vdd.n2759 gnd 0.006542f
C5119 vdd.n2760 gnd 0.006542f
C5120 vdd.n2761 gnd 0.006542f
C5121 vdd.n2762 gnd 0.006542f
C5122 vdd.n2763 gnd 0.006542f
C5123 vdd.n2764 gnd 0.006542f
C5124 vdd.n2765 gnd 0.006542f
C5125 vdd.n2766 gnd 0.006542f
C5126 vdd.n2767 gnd 0.006542f
C5127 vdd.n2768 gnd 0.006542f
C5128 vdd.n2769 gnd 0.006542f
C5129 vdd.n2770 gnd 0.006542f
C5130 vdd.n2771 gnd 0.006542f
C5131 vdd.n2772 gnd 0.006542f
C5132 vdd.n2773 gnd 0.006542f
C5133 vdd.n2774 gnd 0.006542f
C5134 vdd.n2775 gnd 0.006542f
C5135 vdd.n2776 gnd 0.006542f
C5136 vdd.n2777 gnd 0.006542f
C5137 vdd.n2778 gnd 0.006542f
C5138 vdd.n2779 gnd 0.006542f
C5139 vdd.n2780 gnd 0.006542f
C5140 vdd.n2781 gnd 0.006542f
C5141 vdd.n2782 gnd 0.006542f
C5142 vdd.n2783 gnd 0.006542f
C5143 vdd.n2784 gnd 0.006542f
C5144 vdd.n2785 gnd 0.006542f
C5145 vdd.n2786 gnd 0.006542f
C5146 vdd.n2787 gnd 0.006542f
C5147 vdd.n2788 gnd 0.006542f
C5148 vdd.n2789 gnd 0.006542f
C5149 vdd.n2790 gnd 0.006542f
C5150 vdd.n2791 gnd 0.006542f
C5151 vdd.n2792 gnd 0.006542f
C5152 vdd.n2793 gnd 0.006542f
C5153 vdd.n2794 gnd 0.006542f
C5154 vdd.n2795 gnd 0.006542f
C5155 vdd.n2796 gnd 0.006542f
C5156 vdd.n2797 gnd 0.006542f
C5157 vdd.n2798 gnd 0.006542f
C5158 vdd.n2799 gnd 0.006542f
C5159 vdd.n2800 gnd 0.006542f
C5160 vdd.n2801 gnd 0.006542f
C5161 vdd.n2802 gnd 0.006542f
C5162 vdd.n2803 gnd 0.006542f
C5163 vdd.n2804 gnd 0.006542f
C5164 vdd.n2805 gnd 0.004762f
C5165 vdd.n2806 gnd 0.006542f
C5166 vdd.n2807 gnd 0.006542f
C5167 vdd.n2808 gnd 0.005051f
C5168 vdd.n2809 gnd 0.006542f
C5169 vdd.n2810 gnd 0.006542f
C5170 vdd.n2811 gnd 0.014855f
C5171 vdd.n2812 gnd 0.014008f
C5172 vdd.n2813 gnd 0.014008f
C5173 vdd.n2814 gnd 0.006542f
C5174 vdd.n2815 gnd 0.006542f
C5175 vdd.n2816 gnd 0.006542f
C5176 vdd.n2817 gnd 0.006542f
C5177 vdd.n2818 gnd 0.006542f
C5178 vdd.n2819 gnd 0.006542f
C5179 vdd.n2820 gnd 0.006542f
C5180 vdd.n2821 gnd 0.006542f
C5181 vdd.n2822 gnd 0.006542f
C5182 vdd.n2823 gnd 0.006542f
C5183 vdd.n2824 gnd 0.006542f
C5184 vdd.n2825 gnd 0.006542f
C5185 vdd.n2826 gnd 0.006542f
C5186 vdd.n2827 gnd 0.006542f
C5187 vdd.n2828 gnd 0.006542f
C5188 vdd.n2829 gnd 0.006542f
C5189 vdd.n2830 gnd 0.006542f
C5190 vdd.n2831 gnd 0.006542f
C5191 vdd.n2832 gnd 0.006542f
C5192 vdd.n2833 gnd 0.006542f
C5193 vdd.n2834 gnd 0.006542f
C5194 vdd.n2835 gnd 0.006542f
C5195 vdd.n2836 gnd 0.006542f
C5196 vdd.n2837 gnd 0.006542f
C5197 vdd.n2838 gnd 0.006542f
C5198 vdd.n2839 gnd 0.006542f
C5199 vdd.n2840 gnd 0.006542f
C5200 vdd.n2841 gnd 0.006542f
C5201 vdd.n2842 gnd 0.006542f
C5202 vdd.n2843 gnd 0.006542f
C5203 vdd.n2844 gnd 0.006542f
C5204 vdd.n2845 gnd 0.006542f
C5205 vdd.n2846 gnd 0.006542f
C5206 vdd.n2847 gnd 0.006542f
C5207 vdd.n2848 gnd 0.006542f
C5208 vdd.n2849 gnd 0.006542f
C5209 vdd.n2850 gnd 0.006542f
C5210 vdd.n2851 gnd 0.006542f
C5211 vdd.n2852 gnd 0.006542f
C5212 vdd.n2853 gnd 0.006542f
C5213 vdd.n2854 gnd 0.006542f
C5214 vdd.n2855 gnd 0.006542f
C5215 vdd.n2856 gnd 0.006542f
C5216 vdd.n2857 gnd 0.006542f
C5217 vdd.n2858 gnd 0.006542f
C5218 vdd.n2859 gnd 0.006542f
C5219 vdd.n2860 gnd 0.006542f
C5220 vdd.n2861 gnd 0.006542f
C5221 vdd.n2862 gnd 0.006542f
C5222 vdd.n2863 gnd 0.006542f
C5223 vdd.n2864 gnd 0.006542f
C5224 vdd.n2865 gnd 0.006542f
C5225 vdd.n2866 gnd 0.006542f
C5226 vdd.n2867 gnd 0.006542f
C5227 vdd.n2868 gnd 0.006542f
C5228 vdd.n2869 gnd 0.006542f
C5229 vdd.n2870 gnd 0.006542f
C5230 vdd.n2871 gnd 0.006542f
C5231 vdd.n2872 gnd 0.006542f
C5232 vdd.n2873 gnd 0.006542f
C5233 vdd.n2874 gnd 0.006542f
C5234 vdd.n2875 gnd 0.006542f
C5235 vdd.n2876 gnd 0.006542f
C5236 vdd.n2877 gnd 0.006542f
C5237 vdd.n2878 gnd 0.006542f
C5238 vdd.n2879 gnd 0.006542f
C5239 vdd.n2880 gnd 0.006542f
C5240 vdd.n2881 gnd 0.006542f
C5241 vdd.n2882 gnd 0.006542f
C5242 vdd.n2883 gnd 0.006542f
C5243 vdd.n2884 gnd 0.006542f
C5244 vdd.n2885 gnd 0.006542f
C5245 vdd.n2886 gnd 0.006542f
C5246 vdd.n2887 gnd 0.006542f
C5247 vdd.n2888 gnd 0.006542f
C5248 vdd.n2889 gnd 0.006542f
C5249 vdd.n2890 gnd 0.006542f
C5250 vdd.n2891 gnd 0.006542f
C5251 vdd.n2892 gnd 0.006542f
C5252 vdd.n2893 gnd 0.006542f
C5253 vdd.n2894 gnd 0.006542f
C5254 vdd.n2895 gnd 0.006542f
C5255 vdd.n2896 gnd 0.006542f
C5256 vdd.n2897 gnd 0.006542f
C5257 vdd.n2898 gnd 0.006542f
C5258 vdd.n2899 gnd 0.006542f
C5259 vdd.n2900 gnd 0.006542f
C5260 vdd.n2901 gnd 0.006542f
C5261 vdd.n2902 gnd 0.006542f
C5262 vdd.n2903 gnd 0.006542f
C5263 vdd.n2904 gnd 0.006542f
C5264 vdd.n2905 gnd 0.006542f
C5265 vdd.n2906 gnd 0.006542f
C5266 vdd.n2907 gnd 0.006542f
C5267 vdd.n2908 gnd 0.006542f
C5268 vdd.n2909 gnd 0.006542f
C5269 vdd.n2910 gnd 0.006542f
C5270 vdd.n2911 gnd 0.006542f
C5271 vdd.n2912 gnd 0.006542f
C5272 vdd.n2913 gnd 0.006542f
C5273 vdd.n2914 gnd 0.006542f
C5274 vdd.n2915 gnd 0.211389f
C5275 vdd.n2916 gnd 0.006542f
C5276 vdd.n2917 gnd 0.006542f
C5277 vdd.n2918 gnd 0.006542f
C5278 vdd.n2919 gnd 0.006542f
C5279 vdd.n2920 gnd 0.006542f
C5280 vdd.n2921 gnd 0.211389f
C5281 vdd.n2922 gnd 0.006542f
C5282 vdd.n2923 gnd 0.006542f
C5283 vdd.n2924 gnd 0.006542f
C5284 vdd.n2925 gnd 0.006542f
C5285 vdd.n2926 gnd 0.006542f
C5286 vdd.n2927 gnd 0.006542f
C5287 vdd.n2928 gnd 0.006542f
C5288 vdd.n2929 gnd 0.006542f
C5289 vdd.n2930 gnd 0.006542f
C5290 vdd.n2931 gnd 0.006542f
C5291 vdd.n2932 gnd 0.006542f
C5292 vdd.n2933 gnd 0.417863f
C5293 vdd.n2934 gnd 0.006542f
C5294 vdd.n2935 gnd 0.006542f
C5295 vdd.n2936 gnd 0.006542f
C5296 vdd.n2937 gnd 0.014008f
C5297 vdd.n2938 gnd 0.014008f
C5298 vdd.n2939 gnd 0.014855f
C5299 vdd.n2940 gnd 0.014855f
C5300 vdd.n2941 gnd 0.006542f
C5301 vdd.n2942 gnd 0.006542f
C5302 vdd.n2943 gnd 0.006542f
C5303 vdd.n2944 gnd 0.005051f
C5304 vdd.n2945 gnd 0.00935f
C5305 vdd.n2946 gnd 0.004762f
C5306 vdd.n2947 gnd 0.006542f
C5307 vdd.n2948 gnd 0.006542f
C5308 vdd.n2949 gnd 0.006542f
C5309 vdd.n2950 gnd 0.006542f
C5310 vdd.n2951 gnd 0.006542f
C5311 vdd.n2952 gnd 0.006542f
C5312 vdd.n2953 gnd 0.006542f
C5313 vdd.n2954 gnd 0.006542f
C5314 vdd.n2955 gnd 0.006542f
C5315 vdd.n2956 gnd 0.006542f
C5316 vdd.n2957 gnd 0.006542f
C5317 vdd.n2958 gnd 0.006542f
C5318 vdd.n2959 gnd 0.006542f
C5319 vdd.n2960 gnd 0.006542f
C5320 vdd.n2961 gnd 0.006542f
C5321 vdd.n2962 gnd 0.006542f
C5322 vdd.n2963 gnd 0.006542f
C5323 vdd.n2964 gnd 0.006542f
C5324 vdd.n2965 gnd 0.006542f
C5325 vdd.n2966 gnd 0.006542f
C5326 vdd.n2967 gnd 0.006542f
C5327 vdd.n2968 gnd 0.006542f
C5328 vdd.n2969 gnd 0.006542f
C5329 vdd.n2970 gnd 0.006542f
C5330 vdd.n2971 gnd 0.006542f
C5331 vdd.n2972 gnd 0.006542f
C5332 vdd.n2973 gnd 0.006542f
C5333 vdd.n2974 gnd 0.006542f
C5334 vdd.n2975 gnd 0.006542f
C5335 vdd.n2976 gnd 0.006542f
C5336 vdd.n2977 gnd 0.006542f
C5337 vdd.n2978 gnd 0.006542f
C5338 vdd.n2979 gnd 0.006542f
C5339 vdd.n2980 gnd 0.006542f
C5340 vdd.n2981 gnd 0.006542f
C5341 vdd.n2982 gnd 0.006542f
C5342 vdd.n2983 gnd 0.006542f
C5343 vdd.n2984 gnd 0.006542f
C5344 vdd.n2985 gnd 0.006542f
C5345 vdd.n2986 gnd 0.006542f
C5346 vdd.n2987 gnd 0.006542f
C5347 vdd.n2988 gnd 0.006542f
C5348 vdd.n2989 gnd 0.006542f
C5349 vdd.n2990 gnd 0.006542f
C5350 vdd.n2991 gnd 0.006542f
C5351 vdd.n2992 gnd 0.006542f
C5352 vdd.n2993 gnd 0.006542f
C5353 vdd.n2994 gnd 0.006542f
C5354 vdd.n2995 gnd 0.006542f
C5355 vdd.n2996 gnd 0.006542f
C5356 vdd.n2997 gnd 0.006542f
C5357 vdd.n2998 gnd 0.006542f
C5358 vdd.n2999 gnd 0.006542f
C5359 vdd.n3000 gnd 0.006542f
C5360 vdd.n3001 gnd 0.006542f
C5361 vdd.n3002 gnd 0.006542f
C5362 vdd.n3003 gnd 0.006542f
C5363 vdd.n3004 gnd 0.006542f
C5364 vdd.n3005 gnd 0.816061f
C5365 vdd.n3007 gnd 0.014855f
C5366 vdd.n3008 gnd 0.014855f
C5367 vdd.n3009 gnd 0.014008f
C5368 vdd.n3010 gnd 0.006542f
C5369 vdd.n3011 gnd 0.006542f
C5370 vdd.n3012 gnd 0.393283f
C5371 vdd.n3013 gnd 0.006542f
C5372 vdd.n3014 gnd 0.006542f
C5373 vdd.n3015 gnd 0.006542f
C5374 vdd.n3016 gnd 0.006542f
C5375 vdd.n3017 gnd 0.006542f
C5376 vdd.n3018 gnd 0.398199f
C5377 vdd.n3019 gnd 0.006542f
C5378 vdd.n3020 gnd 0.006542f
C5379 vdd.n3021 gnd 0.006542f
C5380 vdd.n3022 gnd 0.006542f
C5381 vdd.n3023 gnd 0.006542f
C5382 vdd.n3024 gnd 0.66858f
C5383 vdd.n3025 gnd 0.006542f
C5384 vdd.n3026 gnd 0.006542f
C5385 vdd.n3027 gnd 0.006542f
C5386 vdd.n3028 gnd 0.006542f
C5387 vdd.n3029 gnd 0.006542f
C5388 vdd.n3030 gnd 0.481771f
C5389 vdd.n3031 gnd 0.006542f
C5390 vdd.n3032 gnd 0.006542f
C5391 vdd.n3033 gnd 0.006542f
C5392 vdd.n3034 gnd 0.006542f
C5393 vdd.n3035 gnd 0.006542f
C5394 vdd.n3036 gnd 0.604672f
C5395 vdd.n3037 gnd 0.006542f
C5396 vdd.n3038 gnd 0.006542f
C5397 vdd.n3039 gnd 0.006542f
C5398 vdd.n3040 gnd 0.006542f
C5399 vdd.n3041 gnd 0.006542f
C5400 vdd.n3042 gnd 0.496519f
C5401 vdd.n3043 gnd 0.006542f
C5402 vdd.n3044 gnd 0.006542f
C5403 vdd.n3045 gnd 0.006542f
C5404 vdd.n3046 gnd 0.006542f
C5405 vdd.n3047 gnd 0.006542f
C5406 vdd.n3048 gnd 0.349038f
C5407 vdd.n3049 gnd 0.006542f
C5408 vdd.n3050 gnd 0.006542f
C5409 vdd.n3051 gnd 0.006542f
C5410 vdd.n3052 gnd 0.006542f
C5411 vdd.n3053 gnd 0.006542f
C5412 vdd.n3054 gnd 0.211389f
C5413 vdd.n3055 gnd 0.006542f
C5414 vdd.n3056 gnd 0.006542f
C5415 vdd.n3057 gnd 0.006542f
C5416 vdd.n3058 gnd 0.006542f
C5417 vdd.n3059 gnd 0.006542f
C5418 vdd.n3060 gnd 0.614504f
C5419 vdd.n3061 gnd 0.006542f
C5420 vdd.n3062 gnd 0.006542f
C5421 vdd.n3063 gnd 0.006542f
C5422 vdd.n3064 gnd 0.004618f
C5423 vdd.n3065 gnd 0.006542f
C5424 vdd.n3066 gnd 0.006542f
C5425 vdd.n3067 gnd 0.66858f
C5426 vdd.n3068 gnd 0.006542f
C5427 vdd.n3069 gnd 0.006542f
C5428 vdd.n3070 gnd 0.006542f
C5429 vdd.n3071 gnd 0.006542f
C5430 vdd.n3072 gnd 0.006542f
C5431 vdd.n3073 gnd 0.530931f
C5432 vdd.n3074 gnd 0.006542f
C5433 vdd.n3075 gnd 0.005195f
C5434 vdd.n3076 gnd 0.006542f
C5435 vdd.n3077 gnd 0.006542f
C5436 vdd.n3078 gnd 0.006542f
C5437 vdd.n3079 gnd 0.427695f
C5438 vdd.n3080 gnd 0.006542f
C5439 vdd.n3081 gnd 0.006542f
C5440 vdd.n3082 gnd 0.006542f
C5441 vdd.n3083 gnd 0.006542f
C5442 vdd.n3084 gnd 0.006542f
C5443 vdd.n3085 gnd 0.388367f
C5444 vdd.n3086 gnd 0.006542f
C5445 vdd.n3087 gnd 0.006542f
C5446 vdd.n3088 gnd 0.006542f
C5447 vdd.n3089 gnd 0.006542f
C5448 vdd.n3090 gnd 0.006542f
C5449 vdd.n3091 gnd 0.535848f
C5450 vdd.n3092 gnd 0.006542f
C5451 vdd.n3093 gnd 0.006542f
C5452 vdd.n3094 gnd 0.006542f
C5453 vdd.n3095 gnd 0.006542f
C5454 vdd.n3096 gnd 0.006542f
C5455 vdd.n3097 gnd 0.66858f
C5456 vdd.n3098 gnd 0.006542f
C5457 vdd.n3099 gnd 0.006542f
C5458 vdd.n3100 gnd 0.006542f
C5459 vdd.n3101 gnd 0.006542f
C5460 vdd.n3102 gnd 0.006542f
C5461 vdd.n3103 gnd 0.653832f
C5462 vdd.n3104 gnd 0.006542f
C5463 vdd.n3105 gnd 0.006542f
C5464 vdd.n3106 gnd 0.006542f
C5465 vdd.n3107 gnd 0.006542f
C5466 vdd.n3108 gnd 0.006542f
C5467 vdd.n3109 gnd 0.506351f
C5468 vdd.n3110 gnd 0.006542f
C5469 vdd.n3111 gnd 0.006542f
C5470 vdd.n3112 gnd 0.006542f
C5471 vdd.n3113 gnd 0.006542f
C5472 vdd.n3114 gnd 0.006542f
C5473 vdd.n3115 gnd 0.35887f
C5474 vdd.n3116 gnd 0.006542f
C5475 vdd.n3117 gnd 0.006542f
C5476 vdd.n3118 gnd 0.006542f
C5477 vdd.n3119 gnd 0.006542f
C5478 vdd.n3120 gnd 0.006542f
C5479 vdd.n3121 gnd 0.66858f
C5480 vdd.n3122 gnd 0.006542f
C5481 vdd.n3123 gnd 0.006542f
C5482 vdd.n3124 gnd 0.006542f
C5483 vdd.n3125 gnd 0.006542f
C5484 vdd.n3126 gnd 0.006542f
C5485 vdd.n3127 gnd 0.006542f
C5486 vdd.n3129 gnd 0.006542f
C5487 vdd.n3130 gnd 0.006542f
C5488 vdd.n3132 gnd 0.006542f
C5489 vdd.n3133 gnd 0.006542f
C5490 vdd.n3136 gnd 0.006542f
C5491 vdd.n3137 gnd 0.006542f
C5492 vdd.n3138 gnd 0.006542f
C5493 vdd.n3139 gnd 0.006542f
C5494 vdd.n3141 gnd 0.006542f
C5495 vdd.n3142 gnd 0.006542f
C5496 vdd.n3143 gnd 0.006542f
C5497 vdd.n3144 gnd 0.006542f
C5498 vdd.n3145 gnd 0.006542f
C5499 vdd.n3146 gnd 0.006542f
C5500 vdd.n3148 gnd 0.006542f
C5501 vdd.n3149 gnd 0.006542f
C5502 vdd.n3150 gnd 0.006542f
C5503 vdd.n3151 gnd 0.006542f
C5504 vdd.n3152 gnd 0.006542f
C5505 vdd.n3153 gnd 0.006542f
C5506 vdd.n3155 gnd 0.006542f
C5507 vdd.n3156 gnd 0.006542f
C5508 vdd.n3157 gnd 0.006542f
C5509 vdd.n3158 gnd 0.006542f
C5510 vdd.n3159 gnd 0.006542f
C5511 vdd.n3160 gnd 0.006542f
C5512 vdd.n3162 gnd 0.006542f
C5513 vdd.n3163 gnd 0.014855f
C5514 vdd.n3164 gnd 0.014855f
C5515 vdd.n3165 gnd 0.014008f
C5516 vdd.n3166 gnd 0.006542f
C5517 vdd.n3167 gnd 0.006542f
C5518 vdd.n3168 gnd 0.006542f
C5519 vdd.n3169 gnd 0.006542f
C5520 vdd.n3170 gnd 0.006542f
C5521 vdd.n3171 gnd 0.006542f
C5522 vdd.n3172 gnd 0.66858f
C5523 vdd.n3173 gnd 0.006542f
C5524 vdd.n3174 gnd 0.006542f
C5525 vdd.n3175 gnd 0.006542f
C5526 vdd.n3176 gnd 0.006542f
C5527 vdd.n3177 gnd 0.006542f
C5528 vdd.n3178 gnd 0.476855f
C5529 vdd.n3179 gnd 0.006542f
C5530 vdd.n3180 gnd 0.006542f
C5531 vdd.n3181 gnd 0.006542f
C5532 vdd.n3182 gnd 0.014855f
C5533 vdd.n3184 gnd 0.014855f
C5534 vdd.n3185 gnd 0.014008f
C5535 vdd.n3186 gnd 0.006542f
C5536 vdd.n3187 gnd 0.005051f
C5537 vdd.n3188 gnd 0.006542f
C5538 vdd.n3190 gnd 0.006542f
C5539 vdd.n3191 gnd 0.006542f
C5540 vdd.n3192 gnd 0.006542f
C5541 vdd.n3193 gnd 0.006542f
C5542 vdd.n3194 gnd 0.006542f
C5543 vdd.n3195 gnd 0.006542f
C5544 vdd.n3197 gnd 0.006542f
C5545 vdd.n3198 gnd 0.006542f
C5546 vdd.n3199 gnd 0.006542f
C5547 vdd.n3200 gnd 0.006542f
C5548 vdd.n3201 gnd 0.006542f
C5549 vdd.n3202 gnd 0.006542f
C5550 vdd.n3204 gnd 0.006542f
C5551 vdd.n3205 gnd 0.006542f
C5552 vdd.n3206 gnd 0.006542f
C5553 vdd.n3207 gnd 0.006542f
C5554 vdd.n3208 gnd 0.006542f
C5555 vdd.n3209 gnd 0.006542f
C5556 vdd.n3211 gnd 0.006542f
C5557 vdd.n3212 gnd 0.006542f
C5558 vdd.n3213 gnd 0.006542f
C5559 vdd.n3214 gnd 1.02503f
C5560 vdd.n3215 gnd 0.040397f
C5561 vdd.n3216 gnd 0.006542f
C5562 vdd.n3217 gnd 0.006542f
C5563 vdd.n3219 gnd 0.006542f
C5564 vdd.n3220 gnd 0.006542f
C5565 vdd.n3221 gnd 0.006542f
C5566 vdd.n3222 gnd 0.006542f
C5567 vdd.n3223 gnd 0.006542f
C5568 vdd.n3224 gnd 0.006542f
C5569 vdd.n3226 gnd 0.006542f
C5570 vdd.n3227 gnd 0.006542f
C5571 vdd.n3228 gnd 0.006542f
C5572 vdd.n3229 gnd 0.006542f
C5573 vdd.n3230 gnd 0.006542f
C5574 vdd.n3231 gnd 0.006542f
C5575 vdd.n3233 gnd 0.006542f
C5576 vdd.n3234 gnd 0.006542f
C5577 vdd.n3235 gnd 0.006542f
C5578 vdd.n3236 gnd 0.006542f
C5579 vdd.n3237 gnd 0.006542f
C5580 vdd.n3238 gnd 0.006542f
C5581 vdd.n3240 gnd 0.006542f
C5582 vdd.n3241 gnd 0.006542f
C5583 vdd.n3243 gnd 0.006542f
C5584 vdd.n3244 gnd 0.006542f
C5585 vdd.n3245 gnd 0.014855f
C5586 vdd.n3246 gnd 0.014008f
C5587 vdd.n3247 gnd 0.014008f
C5588 vdd.n3248 gnd 0.90455f
C5589 vdd.n3249 gnd 0.014008f
C5590 vdd.n3250 gnd 0.014855f
C5591 vdd.n3251 gnd 0.014008f
C5592 vdd.n3252 gnd 0.006542f
C5593 vdd.n3253 gnd 0.005051f
C5594 vdd.n3254 gnd 0.006542f
C5595 vdd.n3256 gnd 0.006542f
C5596 vdd.n3257 gnd 0.006542f
C5597 vdd.n3258 gnd 0.006542f
C5598 vdd.n3259 gnd 0.006542f
C5599 vdd.n3260 gnd 0.006542f
C5600 vdd.n3261 gnd 0.006542f
C5601 vdd.n3263 gnd 0.006542f
C5602 vdd.n3264 gnd 0.006542f
C5603 vdd.n3265 gnd 0.006542f
C5604 vdd.n3266 gnd 0.006542f
C5605 vdd.n3267 gnd 0.006542f
C5606 vdd.n3268 gnd 0.006542f
C5607 vdd.n3270 gnd 0.006542f
C5608 vdd.n3271 gnd 0.006542f
C5609 vdd.n3272 gnd 0.006542f
C5610 vdd.n3273 gnd 0.006542f
C5611 vdd.n3274 gnd 0.006542f
C5612 vdd.n3275 gnd 0.006542f
C5613 vdd.n3277 gnd 0.006542f
C5614 vdd.n3278 gnd 0.006542f
C5615 vdd.n3280 gnd 0.006542f
C5616 vdd.n3281 gnd 0.040397f
C5617 vdd.n3282 gnd 1.02503f
C5618 vdd.n3283 gnd 0.008274f
C5619 vdd.n3284 gnd 0.003678f
C5620 vdd.t217 gnd 0.118362f
C5621 vdd.t218 gnd 0.126496f
C5622 vdd.t215 gnd 0.154579f
C5623 vdd.n3285 gnd 0.198149f
C5624 vdd.n3286 gnd 0.166481f
C5625 vdd.n3287 gnd 0.011925f
C5626 vdd.n3288 gnd 0.009621f
C5627 vdd.n3289 gnd 0.004065f
C5628 vdd.n3290 gnd 0.007744f
C5629 vdd.n3291 gnd 0.009621f
C5630 vdd.n3292 gnd 0.009621f
C5631 vdd.n3293 gnd 0.007744f
C5632 vdd.n3294 gnd 0.007744f
C5633 vdd.n3295 gnd 0.009621f
C5634 vdd.n3297 gnd 0.009621f
C5635 vdd.n3298 gnd 0.007744f
C5636 vdd.n3299 gnd 0.007744f
C5637 vdd.n3300 gnd 0.007744f
C5638 vdd.n3301 gnd 0.009621f
C5639 vdd.n3303 gnd 0.009621f
C5640 vdd.n3305 gnd 0.009621f
C5641 vdd.n3306 gnd 0.007744f
C5642 vdd.n3307 gnd 0.007744f
C5643 vdd.n3308 gnd 0.007744f
C5644 vdd.n3309 gnd 0.009621f
C5645 vdd.n3311 gnd 0.009621f
C5646 vdd.n3313 gnd 0.009621f
C5647 vdd.n3314 gnd 0.007744f
C5648 vdd.n3315 gnd 0.007744f
C5649 vdd.n3316 gnd 0.007744f
C5650 vdd.n3317 gnd 0.009621f
C5651 vdd.n3319 gnd 0.009621f
C5652 vdd.n3320 gnd 0.009621f
C5653 vdd.n3321 gnd 0.007744f
C5654 vdd.n3322 gnd 0.007744f
C5655 vdd.n3323 gnd 0.009621f
C5656 vdd.n3324 gnd 0.009621f
C5657 vdd.n3326 gnd 0.009621f
C5658 vdd.n3327 gnd 0.007744f
C5659 vdd.n3328 gnd 0.009621f
C5660 vdd.n3329 gnd 0.009621f
C5661 vdd.n3330 gnd 0.009621f
C5662 vdd.n3331 gnd 0.015797f
C5663 vdd.n3332 gnd 0.005266f
C5664 vdd.n3333 gnd 0.009621f
C5665 vdd.n3335 gnd 0.009621f
C5666 vdd.n3337 gnd 0.009621f
C5667 vdd.n3338 gnd 0.007744f
C5668 vdd.n3339 gnd 0.007744f
C5669 vdd.n3340 gnd 0.007744f
C5670 vdd.n3341 gnd 0.009621f
C5671 vdd.n3343 gnd 0.009621f
C5672 vdd.n3345 gnd 0.009621f
C5673 vdd.n3346 gnd 0.007744f
C5674 vdd.n3347 gnd 0.007744f
C5675 vdd.n3348 gnd 0.007744f
C5676 vdd.n3349 gnd 0.009621f
C5677 vdd.n3351 gnd 0.009621f
C5678 vdd.n3353 gnd 0.009621f
C5679 vdd.n3354 gnd 0.007744f
C5680 vdd.n3355 gnd 0.007744f
C5681 vdd.n3356 gnd 0.007744f
C5682 vdd.n3357 gnd 0.009621f
C5683 vdd.n3359 gnd 0.009621f
C5684 vdd.n3361 gnd 0.009621f
C5685 vdd.n3362 gnd 0.007744f
C5686 vdd.n3363 gnd 0.007744f
C5687 vdd.n3364 gnd 0.007744f
C5688 vdd.n3365 gnd 0.009621f
C5689 vdd.n3367 gnd 0.009621f
C5690 vdd.n3369 gnd 0.009621f
C5691 vdd.n3370 gnd 0.007744f
C5692 vdd.n3371 gnd 0.007744f
C5693 vdd.n3372 gnd 0.006466f
C5694 vdd.n3373 gnd 0.009621f
C5695 vdd.n3375 gnd 0.009621f
C5696 vdd.n3377 gnd 0.009621f
C5697 vdd.n3378 gnd 0.006466f
C5698 vdd.n3379 gnd 0.007744f
C5699 vdd.n3380 gnd 0.007744f
C5700 vdd.n3381 gnd 0.009621f
C5701 vdd.n3383 gnd 0.009621f
C5702 vdd.n3385 gnd 0.009621f
C5703 vdd.n3386 gnd 0.007744f
C5704 vdd.n3387 gnd 0.007744f
C5705 vdd.n3388 gnd 0.007744f
C5706 vdd.n3389 gnd 0.009621f
C5707 vdd.n3391 gnd 0.009621f
C5708 vdd.n3393 gnd 0.009621f
C5709 vdd.n3394 gnd 0.007744f
C5710 vdd.n3395 gnd 0.007744f
C5711 vdd.n3396 gnd 0.007744f
C5712 vdd.n3397 gnd 0.009621f
C5713 vdd.n3399 gnd 0.009621f
C5714 vdd.n3400 gnd 0.009621f
C5715 vdd.n3401 gnd 0.007744f
C5716 vdd.n3402 gnd 0.007744f
C5717 vdd.n3403 gnd 0.009621f
C5718 vdd.n3404 gnd 0.009621f
C5719 vdd.n3405 gnd 0.007744f
C5720 vdd.n3406 gnd 0.007744f
C5721 vdd.n3407 gnd 0.009621f
C5722 vdd.n3408 gnd 0.009621f
C5723 vdd.n3410 gnd 0.009621f
C5724 vdd.n3411 gnd 0.007744f
C5725 vdd.n3412 gnd 0.006427f
C5726 vdd.n3413 gnd 0.022059f
C5727 vdd.n3414 gnd 0.021909f
C5728 vdd.n3415 gnd 0.006427f
C5729 vdd.n3416 gnd 0.021909f
C5730 vdd.n3417 gnd 1.29783f
C5731 vdd.n3418 gnd 0.021909f
C5732 vdd.n3419 gnd 0.006427f
C5733 vdd.n3420 gnd 0.021909f
C5734 vdd.n3421 gnd 0.009621f
C5735 vdd.n3422 gnd 0.009621f
C5736 vdd.n3423 gnd 0.007744f
C5737 vdd.n3424 gnd 0.009621f
C5738 vdd.n3425 gnd 0.92913f
C5739 vdd.n3426 gnd 0.009621f
C5740 vdd.n3427 gnd 0.007744f
C5741 vdd.n3428 gnd 0.009621f
C5742 vdd.n3429 gnd 0.009621f
C5743 vdd.n3430 gnd 0.009621f
C5744 vdd.n3431 gnd 0.007744f
C5745 vdd.n3432 gnd 0.009621f
C5746 vdd.n3433 gnd 0.958626f
C5747 vdd.n3434 gnd 0.009621f
C5748 vdd.n3435 gnd 0.007744f
C5749 vdd.n3436 gnd 0.009621f
C5750 vdd.n3437 gnd 0.009621f
C5751 vdd.n3438 gnd 0.009621f
C5752 vdd.n3439 gnd 0.007744f
C5753 vdd.n3440 gnd 0.009621f
C5754 vdd.t106 gnd 0.491603f
C5755 vdd.n3441 gnd 0.791481f
C5756 vdd.n3442 gnd 0.009621f
C5757 vdd.n3443 gnd 0.007744f
C5758 vdd.n3444 gnd 0.009621f
C5759 vdd.n3445 gnd 0.009621f
C5760 vdd.n3446 gnd 0.009621f
C5761 vdd.n3447 gnd 0.007744f
C5762 vdd.n3448 gnd 0.009621f
C5763 vdd.n3449 gnd 0.624336f
C5764 vdd.n3450 gnd 0.009621f
C5765 vdd.n3451 gnd 0.007744f
C5766 vdd.n3452 gnd 0.009621f
C5767 vdd.n3453 gnd 0.009621f
C5768 vdd.n3454 gnd 0.009621f
C5769 vdd.n3455 gnd 0.007744f
C5770 vdd.n3456 gnd 0.009621f
C5771 vdd.n3457 gnd 0.781649f
C5772 vdd.n3458 gnd 0.526015f
C5773 vdd.n3459 gnd 0.009621f
C5774 vdd.n3460 gnd 0.007744f
C5775 vdd.n3461 gnd 0.009621f
C5776 vdd.n3462 gnd 0.009621f
C5777 vdd.n3463 gnd 0.009621f
C5778 vdd.n3464 gnd 0.007744f
C5779 vdd.n3465 gnd 0.009621f
C5780 vdd.n3466 gnd 0.693161f
C5781 vdd.n3467 gnd 0.009621f
C5782 vdd.n3468 gnd 0.007744f
C5783 vdd.n3469 gnd 0.009621f
C5784 vdd.n3470 gnd 0.009621f
C5785 vdd.n3471 gnd 0.009621f
C5786 vdd.n3472 gnd 0.009621f
C5787 vdd.n3473 gnd 0.009621f
C5788 vdd.n3474 gnd 0.007744f
C5789 vdd.n3475 gnd 0.007744f
C5790 vdd.n3476 gnd 0.009621f
C5791 vdd.t127 gnd 0.491603f
C5792 vdd.n3477 gnd 0.816061f
C5793 vdd.n3478 gnd 0.009621f
C5794 vdd.n3479 gnd 0.007744f
C5795 vdd.n3480 gnd 0.009621f
C5796 vdd.n3481 gnd 0.009621f
C5797 vdd.n3482 gnd 0.009621f
C5798 vdd.n3483 gnd 0.007744f
C5799 vdd.n3484 gnd 0.009621f
C5800 vdd.n3485 gnd 0.771817f
C5801 vdd.n3486 gnd 0.009621f
C5802 vdd.n3487 gnd 0.009621f
C5803 vdd.n3488 gnd 0.007744f
C5804 vdd.n3489 gnd 0.007744f
C5805 vdd.n3490 gnd 0.007744f
C5806 vdd.n3491 gnd 0.009621f
C5807 vdd.n3492 gnd 0.009621f
C5808 vdd.n3493 gnd 0.009621f
C5809 vdd.n3494 gnd 0.009621f
C5810 vdd.n3495 gnd 0.007744f
C5811 vdd.n3496 gnd 0.007744f
C5812 vdd.n3497 gnd 0.007744f
C5813 vdd.n3498 gnd 0.009621f
C5814 vdd.n3499 gnd 0.009621f
C5815 vdd.n3500 gnd 0.009621f
C5816 vdd.n3501 gnd 0.009621f
C5817 vdd.n3502 gnd 0.007744f
C5818 vdd.n3503 gnd 0.007744f
C5819 vdd.n3504 gnd 0.007744f
C5820 vdd.n3505 gnd 0.009621f
C5821 vdd.n3506 gnd 0.009621f
C5822 vdd.n3507 gnd 0.009621f
C5823 vdd.n3508 gnd 0.816061f
C5824 vdd.n3509 gnd 0.009621f
C5825 vdd.n3510 gnd 0.007744f
C5826 vdd.n3511 gnd 0.007744f
C5827 vdd.n3512 gnd 0.007744f
C5828 vdd.n3513 gnd 0.009621f
C5829 vdd.n3514 gnd 0.009621f
C5830 vdd.n3515 gnd 0.009621f
C5831 vdd.n3516 gnd 0.009621f
C5832 vdd.n3517 gnd 0.007744f
C5833 vdd.n3518 gnd 0.007744f
C5834 vdd.n3519 gnd 0.006427f
C5835 vdd.n3520 gnd 0.021909f
C5836 vdd.n3521 gnd 0.022059f
C5837 vdd.n3522 gnd 0.003678f
C5838 vdd.n3523 gnd 0.022059f
C5839 vdd.n3525 gnd 2.17289f
C5840 vdd.n3526 gnd 1.29783f
C5841 vdd.n3527 gnd 0.644f
C5842 vdd.n3528 gnd 0.009621f
C5843 vdd.n3529 gnd 0.007744f
C5844 vdd.n3530 gnd 0.007744f
C5845 vdd.n3531 gnd 0.007744f
C5846 vdd.n3532 gnd 0.009621f
C5847 vdd.n3533 gnd 0.983206f
C5848 vdd.n3534 gnd 0.983206f
C5849 vdd.n3535 gnd 0.565344f
C5850 vdd.n3536 gnd 0.009621f
C5851 vdd.n3537 gnd 0.007744f
C5852 vdd.n3538 gnd 0.007744f
C5853 vdd.n3539 gnd 0.007744f
C5854 vdd.n3540 gnd 0.009621f
C5855 vdd.n3541 gnd 0.585008f
C5856 vdd.n3542 gnd 0.722657f
C5857 vdd.t122 gnd 0.491603f
C5858 vdd.n3543 gnd 0.752153f
C5859 vdd.n3544 gnd 0.009621f
C5860 vdd.n3545 gnd 0.007744f
C5861 vdd.n3546 gnd 0.007744f
C5862 vdd.n3547 gnd 0.007744f
C5863 vdd.n3548 gnd 0.009621f
C5864 vdd.n3549 gnd 0.816061f
C5865 vdd.t82 gnd 0.491603f
C5866 vdd.n3550 gnd 0.59484f
C5867 vdd.n3551 gnd 0.712825f
C5868 vdd.n3552 gnd 0.009621f
C5869 vdd.n3553 gnd 0.007744f
C5870 vdd.n3554 gnd 0.007744f
C5871 vdd.n3555 gnd 0.007744f
C5872 vdd.n3556 gnd 0.009621f
C5873 vdd.n3557 gnd 0.54568f
C5874 vdd.t112 gnd 0.491603f
C5875 vdd.n3558 gnd 0.816061f
C5876 vdd.t76 gnd 0.491603f
C5877 vdd.n3559 gnd 0.604672f
C5878 vdd.n3560 gnd 0.009621f
C5879 vdd.n3561 gnd 0.007744f
C5880 vdd.n3562 gnd 0.007394f
C5881 vdd.n3563 gnd 0.567475f
C5882 vdd.n3564 gnd 2.64002f
C5883 a_n2804_13878.t19 gnd 0.194556f
C5884 a_n2804_13878.t6 gnd 0.194556f
C5885 a_n2804_13878.t16 gnd 0.194556f
C5886 a_n2804_13878.n0 gnd 1.53358f
C5887 a_n2804_13878.t21 gnd 0.194556f
C5888 a_n2804_13878.t11 gnd 0.194556f
C5889 a_n2804_13878.n1 gnd 1.53196f
C5890 a_n2804_13878.n2 gnd 2.14061f
C5891 a_n2804_13878.t17 gnd 0.194556f
C5892 a_n2804_13878.t10 gnd 0.194556f
C5893 a_n2804_13878.n3 gnd 1.53196f
C5894 a_n2804_13878.n4 gnd 1.04414f
C5895 a_n2804_13878.t4 gnd 0.194556f
C5896 a_n2804_13878.t7 gnd 0.194556f
C5897 a_n2804_13878.n5 gnd 1.53196f
C5898 a_n2804_13878.n6 gnd 1.04414f
C5899 a_n2804_13878.t20 gnd 0.194556f
C5900 a_n2804_13878.t5 gnd 0.194556f
C5901 a_n2804_13878.n7 gnd 1.53196f
C5902 a_n2804_13878.n8 gnd 1.04414f
C5903 a_n2804_13878.t15 gnd 0.194556f
C5904 a_n2804_13878.t3 gnd 0.194556f
C5905 a_n2804_13878.n9 gnd 1.53196f
C5906 a_n2804_13878.n10 gnd 4.90178f
C5907 a_n2804_13878.t27 gnd 1.82172f
C5908 a_n2804_13878.t28 gnd 0.194556f
C5909 a_n2804_13878.t31 gnd 0.194556f
C5910 a_n2804_13878.n11 gnd 1.37045f
C5911 a_n2804_13878.n12 gnd 1.53128f
C5912 a_n2804_13878.t1 gnd 1.81809f
C5913 a_n2804_13878.n13 gnd 0.770559f
C5914 a_n2804_13878.t0 gnd 1.81809f
C5915 a_n2804_13878.n14 gnd 0.770559f
C5916 a_n2804_13878.t29 gnd 0.194556f
C5917 a_n2804_13878.t30 gnd 0.194556f
C5918 a_n2804_13878.n15 gnd 1.37045f
C5919 a_n2804_13878.n16 gnd 0.778022f
C5920 a_n2804_13878.t26 gnd 1.81809f
C5921 a_n2804_13878.n17 gnd 2.85814f
C5922 a_n2804_13878.n18 gnd 3.74876f
C5923 a_n2804_13878.t9 gnd 0.194556f
C5924 a_n2804_13878.t18 gnd 0.194556f
C5925 a_n2804_13878.n19 gnd 1.53195f
C5926 a_n2804_13878.n20 gnd 2.50239f
C5927 a_n2804_13878.t22 gnd 0.194556f
C5928 a_n2804_13878.t8 gnd 0.194556f
C5929 a_n2804_13878.n21 gnd 1.53196f
C5930 a_n2804_13878.n22 gnd 0.678771f
C5931 a_n2804_13878.t12 gnd 0.194556f
C5932 a_n2804_13878.t13 gnd 0.194556f
C5933 a_n2804_13878.n23 gnd 1.53196f
C5934 a_n2804_13878.n24 gnd 0.678771f
C5935 a_n2804_13878.t23 gnd 0.194556f
C5936 a_n2804_13878.t24 gnd 0.194556f
C5937 a_n2804_13878.n25 gnd 1.53196f
C5938 a_n2804_13878.n26 gnd 0.678771f
C5939 a_n2804_13878.t2 gnd 0.194556f
C5940 a_n2804_13878.t14 gnd 0.194556f
C5941 a_n2804_13878.n27 gnd 1.53196f
C5942 a_n2804_13878.n28 gnd 1.37704f
C5943 a_n2804_13878.n29 gnd 1.5345f
C5944 a_n2804_13878.t25 gnd 0.194556f
C5945 a_n2982_13878.n0 gnd 2.53375f
C5946 a_n2982_13878.n1 gnd 3.78544f
C5947 a_n2982_13878.n2 gnd 3.42813f
C5948 a_n2982_13878.n3 gnd 0.20945f
C5949 a_n2982_13878.n4 gnd 0.20945f
C5950 a_n2982_13878.n5 gnd 0.791576f
C5951 a_n2982_13878.n6 gnd 0.20945f
C5952 a_n2982_13878.n7 gnd 0.971817f
C5953 a_n2982_13878.n8 gnd 0.20945f
C5954 a_n2982_13878.n9 gnd 0.20945f
C5955 a_n2982_13878.n10 gnd 0.458033f
C5956 a_n2982_13878.n11 gnd 0.20945f
C5957 a_n2982_13878.n12 gnd 0.27462f
C5958 a_n2982_13878.n13 gnd 0.90404f
C5959 a_n2982_13878.n14 gnd 0.198733f
C5960 a_n2982_13878.n15 gnd 0.146371f
C5961 a_n2982_13878.n16 gnd 0.230048f
C5962 a_n2982_13878.n17 gnd 0.177686f
C5963 a_n2982_13878.n18 gnd 0.198733f
C5964 a_n2982_13878.n19 gnd 1.32386f
C5965 a_n2982_13878.n20 gnd 0.146371f
C5966 a_n2982_13878.n21 gnd 0.956403f
C5967 a_n2982_13878.n22 gnd 0.20945f
C5968 a_n2982_13878.n23 gnd 0.73719f
C5969 a_n2982_13878.n24 gnd 0.20945f
C5970 a_n2982_13878.n25 gnd 0.20945f
C5971 a_n2982_13878.n26 gnd 0.477018f
C5972 a_n2982_13878.n27 gnd 0.27462f
C5973 a_n2982_13878.n28 gnd 0.20945f
C5974 a_n2982_13878.n29 gnd 0.529381f
C5975 a_n2982_13878.n30 gnd 0.20945f
C5976 a_n2982_13878.n31 gnd 0.20945f
C5977 a_n2982_13878.n32 gnd 0.931898f
C5978 a_n2982_13878.n33 gnd 0.27462f
C5979 a_n2982_13878.n34 gnd 3.08362f
C5980 a_n2982_13878.n35 gnd 0.27462f
C5981 a_n2982_13878.n36 gnd 1.72437f
C5982 a_n2982_13878.n37 gnd 1.16191f
C5983 a_n2982_13878.n38 gnd 2.32061f
C5984 a_n2982_13878.n39 gnd 2.12168f
C5985 a_n2982_13878.n40 gnd 1.72437f
C5986 a_n2982_13878.n41 gnd 1.16191f
C5987 a_n2982_13878.n42 gnd 0.008404f
C5988 a_n2982_13878.n43 gnd 4.05e-19
C5989 a_n2982_13878.n45 gnd 0.008109f
C5990 a_n2982_13878.n46 gnd 0.011792f
C5991 a_n2982_13878.n47 gnd 0.007801f
C5992 a_n2982_13878.n49 gnd 0.277816f
C5993 a_n2982_13878.n50 gnd 0.008404f
C5994 a_n2982_13878.n51 gnd 4.05e-19
C5995 a_n2982_13878.n53 gnd 0.008109f
C5996 a_n2982_13878.n54 gnd 0.011792f
C5997 a_n2982_13878.n55 gnd 0.007801f
C5998 a_n2982_13878.n57 gnd 0.277816f
C5999 a_n2982_13878.n58 gnd 0.008109f
C6000 a_n2982_13878.n59 gnd 0.276683f
C6001 a_n2982_13878.n60 gnd 0.008109f
C6002 a_n2982_13878.n61 gnd 0.276683f
C6003 a_n2982_13878.n62 gnd 0.008109f
C6004 a_n2982_13878.n63 gnd 0.276683f
C6005 a_n2982_13878.n64 gnd 0.008109f
C6006 a_n2982_13878.n65 gnd 0.276683f
C6007 a_n2982_13878.n66 gnd 0.008404f
C6008 a_n2982_13878.n67 gnd 4.05e-19
C6009 a_n2982_13878.n69 gnd 0.008109f
C6010 a_n2982_13878.n70 gnd 0.011792f
C6011 a_n2982_13878.n71 gnd 0.007801f
C6012 a_n2982_13878.n73 gnd 0.277816f
C6013 a_n2982_13878.n74 gnd 0.277816f
C6014 a_n2982_13878.n76 gnd 0.007801f
C6015 a_n2982_13878.n77 gnd 0.011792f
C6016 a_n2982_13878.n78 gnd 0.008109f
C6017 a_n2982_13878.n80 gnd 4.05e-19
C6018 a_n2982_13878.n81 gnd 0.008404f
C6019 a_n2982_13878.n82 gnd 0.104725f
C6020 a_n2982_13878.t51 gnd 0.145277f
C6021 a_n2982_13878.t12 gnd 0.686627f
C6022 a_n2982_13878.t10 gnd 0.675756f
C6023 a_n2982_13878.t30 gnd 0.675756f
C6024 a_n2982_13878.t26 gnd 0.675756f
C6025 a_n2982_13878.n83 gnd 0.293584f
C6026 a_n2982_13878.t48 gnd 0.675756f
C6027 a_n2982_13878.t6 gnd 0.675756f
C6028 a_n2982_13878.t50 gnd 0.675756f
C6029 a_n2982_13878.n84 gnd 0.297105f
C6030 a_n2982_13878.t34 gnd 0.675756f
C6031 a_n2982_13878.t22 gnd 0.675756f
C6032 a_n2982_13878.t38 gnd 0.675756f
C6033 a_n2982_13878.n85 gnd 0.293009f
C6034 a_n2982_13878.t42 gnd 0.675756f
C6035 a_n2982_13878.t40 gnd 0.689824f
C6036 a_n2982_13878.t102 gnd 0.689824f
C6037 a_n2982_13878.t79 gnd 0.675756f
C6038 a_n2982_13878.t84 gnd 0.675756f
C6039 a_n2982_13878.t72 gnd 0.675756f
C6040 a_n2982_13878.n86 gnd 0.296971f
C6041 a_n2982_13878.t89 gnd 0.675756f
C6042 a_n2982_13878.t98 gnd 0.675756f
C6043 a_n2982_13878.t99 gnd 0.675756f
C6044 a_n2982_13878.n87 gnd 0.293332f
C6045 a_n2982_13878.t66 gnd 0.675756f
C6046 a_n2982_13878.t81 gnd 0.675756f
C6047 a_n2982_13878.t69 gnd 0.675756f
C6048 a_n2982_13878.n88 gnd 0.29709f
C6049 a_n2982_13878.t76 gnd 0.675756f
C6050 a_n2982_13878.t95 gnd 0.686627f
C6051 a_n2982_13878.t9 gnd 1.3603f
C6052 a_n2982_13878.t45 gnd 0.145277f
C6053 a_n2982_13878.t53 gnd 0.145277f
C6054 a_n2982_13878.n89 gnd 1.02333f
C6055 a_n2982_13878.t47 gnd 0.145277f
C6056 a_n2982_13878.t21 gnd 0.145277f
C6057 a_n2982_13878.n90 gnd 1.02333f
C6058 a_n2982_13878.t33 gnd 0.145277f
C6059 a_n2982_13878.t15 gnd 0.145277f
C6060 a_n2982_13878.n91 gnd 1.02333f
C6061 a_n2982_13878.t37 gnd 0.145277f
C6062 a_n2982_13878.t17 gnd 0.145277f
C6063 a_n2982_13878.n92 gnd 1.02333f
C6064 a_n2982_13878.t25 gnd 0.145277f
C6065 a_n2982_13878.t29 gnd 0.145277f
C6066 a_n2982_13878.n93 gnd 1.02333f
C6067 a_n2982_13878.t19 gnd 1.35758f
C6068 a_n2982_13878.t24 gnd 0.675756f
C6069 a_n2982_13878.n94 gnd 0.29709f
C6070 a_n2982_13878.t28 gnd 0.675756f
C6071 a_n2982_13878.t36 gnd 0.675756f
C6072 a_n2982_13878.n95 gnd 0.288167f
C6073 a_n2982_13878.t20 gnd 0.675756f
C6074 a_n2982_13878.n96 gnd 0.299644f
C6075 a_n2982_13878.t32 gnd 0.675756f
C6076 a_n2982_13878.t52 gnd 0.675756f
C6077 a_n2982_13878.n97 gnd 0.293009f
C6078 a_n2982_13878.t8 gnd 0.689824f
C6079 a_n2982_13878.t78 gnd 0.675756f
C6080 a_n2982_13878.n98 gnd 0.29709f
C6081 a_n2982_13878.t87 gnd 0.675756f
C6082 a_n2982_13878.t93 gnd 0.675756f
C6083 a_n2982_13878.n99 gnd 0.288167f
C6084 a_n2982_13878.t97 gnd 0.675756f
C6085 a_n2982_13878.n100 gnd 0.299644f
C6086 a_n2982_13878.t68 gnd 0.675756f
C6087 a_n2982_13878.t71 gnd 0.675756f
C6088 a_n2982_13878.n101 gnd 0.293009f
C6089 a_n2982_13878.t101 gnd 0.689824f
C6090 a_n2982_13878.t70 gnd 0.675756f
C6091 a_n2982_13878.n102 gnd 0.299205f
C6092 a_n2982_13878.t96 gnd 0.675756f
C6093 a_n2982_13878.n103 gnd 0.296971f
C6094 a_n2982_13878.n104 gnd 0.297105f
C6095 a_n2982_13878.t92 gnd 0.675756f
C6096 a_n2982_13878.n105 gnd 0.293332f
C6097 a_n2982_13878.t65 gnd 0.675756f
C6098 a_n2982_13878.n106 gnd 0.293584f
C6099 a_n2982_13878.n107 gnd 0.299206f
C6100 a_n2982_13878.t67 gnd 0.686627f
C6101 a_n2982_13878.t44 gnd 0.675756f
C6102 a_n2982_13878.n108 gnd 0.299205f
C6103 a_n2982_13878.t46 gnd 0.675756f
C6104 a_n2982_13878.n109 gnd 0.296971f
C6105 a_n2982_13878.n110 gnd 0.297105f
C6106 a_n2982_13878.t14 gnd 0.675756f
C6107 a_n2982_13878.n111 gnd 0.293332f
C6108 a_n2982_13878.t16 gnd 0.675756f
C6109 a_n2982_13878.n112 gnd 0.293584f
C6110 a_n2982_13878.n113 gnd 0.299206f
C6111 a_n2982_13878.t18 gnd 0.686627f
C6112 a_n2982_13878.n114 gnd 1.30834f
C6113 a_n2982_13878.t75 gnd 0.675756f
C6114 a_n2982_13878.n115 gnd 0.293332f
C6115 a_n2982_13878.t83 gnd 0.675756f
C6116 a_n2982_13878.n116 gnd 0.293332f
C6117 a_n2982_13878.t73 gnd 0.675756f
C6118 a_n2982_13878.n117 gnd 0.293332f
C6119 a_n2982_13878.t88 gnd 0.675756f
C6120 a_n2982_13878.n118 gnd 0.293332f
C6121 a_n2982_13878.t77 gnd 0.675756f
C6122 a_n2982_13878.n119 gnd 0.288005f
C6123 a_n2982_13878.t103 gnd 0.675756f
C6124 a_n2982_13878.n120 gnd 0.297105f
C6125 a_n2982_13878.t80 gnd 0.687079f
C6126 a_n2982_13878.t90 gnd 0.675756f
C6127 a_n2982_13878.n121 gnd 0.288005f
C6128 a_n2982_13878.t74 gnd 0.675756f
C6129 a_n2982_13878.n122 gnd 0.297105f
C6130 a_n2982_13878.t85 gnd 0.687079f
C6131 a_n2982_13878.t94 gnd 0.675756f
C6132 a_n2982_13878.n123 gnd 0.288005f
C6133 a_n2982_13878.t82 gnd 0.675756f
C6134 a_n2982_13878.n124 gnd 0.297105f
C6135 a_n2982_13878.t100 gnd 0.687079f
C6136 a_n2982_13878.t86 gnd 0.675756f
C6137 a_n2982_13878.n125 gnd 0.288005f
C6138 a_n2982_13878.t64 gnd 0.675756f
C6139 a_n2982_13878.n126 gnd 0.297105f
C6140 a_n2982_13878.t91 gnd 0.687079f
C6141 a_n2982_13878.n127 gnd 1.64574f
C6142 a_n2982_13878.n128 gnd 0.299206f
C6143 a_n2982_13878.n129 gnd 0.293584f
C6144 a_n2982_13878.n130 gnd 0.288167f
C6145 a_n2982_13878.n131 gnd 0.297105f
C6146 a_n2982_13878.n132 gnd 0.299644f
C6147 a_n2982_13878.n133 gnd 0.293009f
C6148 a_n2982_13878.n134 gnd 0.299205f
C6149 a_n2982_13878.t5 gnd 0.112993f
C6150 a_n2982_13878.t63 gnd 0.112993f
C6151 a_n2982_13878.n135 gnd 1.00066f
C6152 a_n2982_13878.t4 gnd 0.112993f
C6153 a_n2982_13878.t58 gnd 0.112993f
C6154 a_n2982_13878.n136 gnd 0.998444f
C6155 a_n2982_13878.t54 gnd 0.112993f
C6156 a_n2982_13878.t56 gnd 0.112993f
C6157 a_n2982_13878.n137 gnd 1.00066f
C6158 a_n2982_13878.t61 gnd 0.112993f
C6159 a_n2982_13878.t60 gnd 0.112993f
C6160 a_n2982_13878.n138 gnd 0.998444f
C6161 a_n2982_13878.t59 gnd 0.112993f
C6162 a_n2982_13878.t55 gnd 0.112993f
C6163 a_n2982_13878.n139 gnd 0.998444f
C6164 a_n2982_13878.t62 gnd 0.112993f
C6165 a_n2982_13878.t57 gnd 0.112993f
C6166 a_n2982_13878.n140 gnd 0.998444f
C6167 a_n2982_13878.t1 gnd 0.112993f
C6168 a_n2982_13878.t2 gnd 0.112993f
C6169 a_n2982_13878.n141 gnd 1.00066f
C6170 a_n2982_13878.t3 gnd 0.112993f
C6171 a_n2982_13878.t0 gnd 0.112993f
C6172 a_n2982_13878.n142 gnd 0.998444f
C6173 a_n2982_13878.n143 gnd 0.299205f
C6174 a_n2982_13878.n144 gnd 0.296971f
C6175 a_n2982_13878.n145 gnd 0.299644f
C6176 a_n2982_13878.n146 gnd 0.293332f
C6177 a_n2982_13878.n147 gnd 0.288167f
C6178 a_n2982_13878.n148 gnd 0.29709f
C6179 a_n2982_13878.n149 gnd 0.299206f
C6180 a_n2982_13878.n150 gnd 0.994805f
C6181 a_n2982_13878.t13 gnd 1.35759f
C6182 a_n2982_13878.t11 gnd 0.145277f
C6183 a_n2982_13878.t31 gnd 0.145277f
C6184 a_n2982_13878.n151 gnd 1.02333f
C6185 a_n2982_13878.t27 gnd 0.145277f
C6186 a_n2982_13878.t49 gnd 0.145277f
C6187 a_n2982_13878.n152 gnd 1.02333f
C6188 a_n2982_13878.t41 gnd 1.3603f
C6189 a_n2982_13878.t39 gnd 0.145277f
C6190 a_n2982_13878.t43 gnd 0.145277f
C6191 a_n2982_13878.n153 gnd 1.02333f
C6192 a_n2982_13878.t35 gnd 0.145277f
C6193 a_n2982_13878.t23 gnd 0.145277f
C6194 a_n2982_13878.n154 gnd 1.02333f
C6195 a_n2982_13878.n155 gnd 1.02333f
C6196 a_n2982_13878.t7 gnd 0.145277f
C6197 a_n8964_8799.t33 gnd 0.112902f
C6198 a_n8964_8799.t17 gnd 0.145159f
C6199 a_n8964_8799.t19 gnd 0.145159f
C6200 a_n8964_8799.n0 gnd 1.14489f
C6201 a_n8964_8799.t0 gnd 0.145159f
C6202 a_n8964_8799.t15 gnd 0.145159f
C6203 a_n8964_8799.n1 gnd 1.143f
C6204 a_n8964_8799.n2 gnd 1.02742f
C6205 a_n8964_8799.t7 gnd 0.145159f
C6206 a_n8964_8799.t2 gnd 0.145159f
C6207 a_n8964_8799.n3 gnd 1.143f
C6208 a_n8964_8799.n4 gnd 0.506435f
C6209 a_n8964_8799.t21 gnd 0.145159f
C6210 a_n8964_8799.t9 gnd 0.145159f
C6211 a_n8964_8799.n5 gnd 1.143f
C6212 a_n8964_8799.n6 gnd 0.506435f
C6213 a_n8964_8799.t14 gnd 0.145159f
C6214 a_n8964_8799.t20 gnd 0.145159f
C6215 a_n8964_8799.n7 gnd 1.143f
C6216 a_n8964_8799.n8 gnd 0.506435f
C6217 a_n8964_8799.t10 gnd 0.145159f
C6218 a_n8964_8799.t16 gnd 0.145159f
C6219 a_n8964_8799.n9 gnd 1.143f
C6220 a_n8964_8799.n10 gnd 3.67991f
C6221 a_n8964_8799.t8 gnd 0.145159f
C6222 a_n8964_8799.t38 gnd 0.145159f
C6223 a_n8964_8799.n11 gnd 1.14489f
C6224 a_n8964_8799.t6 gnd 0.145159f
C6225 a_n8964_8799.t39 gnd 0.145159f
C6226 a_n8964_8799.n12 gnd 1.143f
C6227 a_n8964_8799.n13 gnd 1.02742f
C6228 a_n8964_8799.t4 gnd 0.145159f
C6229 a_n8964_8799.t11 gnd 0.145159f
C6230 a_n8964_8799.n14 gnd 1.143f
C6231 a_n8964_8799.n15 gnd 0.506435f
C6232 a_n8964_8799.t3 gnd 0.145159f
C6233 a_n8964_8799.t18 gnd 0.145159f
C6234 a_n8964_8799.n16 gnd 1.143f
C6235 a_n8964_8799.n17 gnd 0.506435f
C6236 a_n8964_8799.t5 gnd 0.145159f
C6237 a_n8964_8799.t1 gnd 0.145159f
C6238 a_n8964_8799.n18 gnd 1.143f
C6239 a_n8964_8799.n19 gnd 0.506435f
C6240 a_n8964_8799.t12 gnd 0.145159f
C6241 a_n8964_8799.t13 gnd 0.145159f
C6242 a_n8964_8799.n20 gnd 1.143f
C6243 a_n8964_8799.n21 gnd 2.55489f
C6244 a_n8964_8799.n22 gnd 7.68275f
C6245 a_n8964_8799.n23 gnd 0.05232f
C6246 a_n8964_8799.t77 gnd 0.601897f
C6247 a_n8964_8799.n24 gnd 0.268819f
C6248 a_n8964_8799.n25 gnd 0.05232f
C6249 a_n8964_8799.n26 gnd 0.011873f
C6250 a_n8964_8799.t106 gnd 0.601897f
C6251 a_n8964_8799.n27 gnd 0.05232f
C6252 a_n8964_8799.t122 gnd 0.601897f
C6253 a_n8964_8799.n28 gnd 0.268658f
C6254 a_n8964_8799.t123 gnd 0.601897f
C6255 a_n8964_8799.n29 gnd 0.05232f
C6256 a_n8964_8799.n30 gnd 0.011873f
C6257 a_n8964_8799.t65 gnd 0.601897f
C6258 a_n8964_8799.n31 gnd 0.05232f
C6259 a_n8964_8799.t66 gnd 0.601897f
C6260 a_n8964_8799.n32 gnd 0.263819f
C6261 a_n8964_8799.t99 gnd 0.601897f
C6262 a_n8964_8799.n33 gnd 0.05232f
C6263 a_n8964_8799.t104 gnd 0.601897f
C6264 a_n8964_8799.n34 gnd 0.268012f
C6265 a_n8964_8799.t79 gnd 0.613289f
C6266 a_n8964_8799.n35 gnd 0.252342f
C6267 a_n8964_8799.n36 gnd 0.171077f
C6268 a_n8964_8799.n37 gnd 0.011873f
C6269 a_n8964_8799.t42 gnd 0.601897f
C6270 a_n8964_8799.n38 gnd 0.268819f
C6271 a_n8964_8799.n39 gnd 0.011873f
C6272 a_n8964_8799.n40 gnd 0.05232f
C6273 a_n8964_8799.n41 gnd 0.05232f
C6274 a_n8964_8799.n42 gnd 0.05232f
C6275 a_n8964_8799.n43 gnd 0.268335f
C6276 a_n8964_8799.n44 gnd 0.011873f
C6277 a_n8964_8799.t126 gnd 0.601897f
C6278 a_n8964_8799.n45 gnd 0.268819f
C6279 a_n8964_8799.n46 gnd 0.05232f
C6280 a_n8964_8799.n47 gnd 0.05232f
C6281 a_n8964_8799.n48 gnd 0.05232f
C6282 a_n8964_8799.n49 gnd 0.263496f
C6283 a_n8964_8799.t95 gnd 0.601897f
C6284 a_n8964_8799.n50 gnd 0.268658f
C6285 a_n8964_8799.n51 gnd 0.011873f
C6286 a_n8964_8799.n52 gnd 0.05232f
C6287 a_n8964_8799.n53 gnd 0.05232f
C6288 a_n8964_8799.n54 gnd 0.05232f
C6289 a_n8964_8799.n55 gnd 0.263496f
C6290 a_n8964_8799.n56 gnd 0.011873f
C6291 a_n8964_8799.t80 gnd 0.601897f
C6292 a_n8964_8799.n57 gnd 0.268819f
C6293 a_n8964_8799.n58 gnd 0.05232f
C6294 a_n8964_8799.n59 gnd 0.05232f
C6295 a_n8964_8799.n60 gnd 0.05232f
C6296 a_n8964_8799.n61 gnd 0.268335f
C6297 a_n8964_8799.t121 gnd 0.601897f
C6298 a_n8964_8799.n62 gnd 0.263819f
C6299 a_n8964_8799.n63 gnd 0.011873f
C6300 a_n8964_8799.n64 gnd 0.05232f
C6301 a_n8964_8799.n65 gnd 0.05232f
C6302 a_n8964_8799.n66 gnd 0.05232f
C6303 a_n8964_8799.n67 gnd 0.011873f
C6304 a_n8964_8799.t78 gnd 0.601897f
C6305 a_n8964_8799.n68 gnd 0.268012f
C6306 a_n8964_8799.t103 gnd 0.601897f
C6307 a_n8964_8799.n69 gnd 0.263335f
C6308 a_n8964_8799.n70 gnd 0.301459f
C6309 a_n8964_8799.n71 gnd 0.05232f
C6310 a_n8964_8799.t86 gnd 0.601897f
C6311 a_n8964_8799.n72 gnd 0.268819f
C6312 a_n8964_8799.n73 gnd 0.05232f
C6313 a_n8964_8799.n74 gnd 0.011873f
C6314 a_n8964_8799.t118 gnd 0.601897f
C6315 a_n8964_8799.n75 gnd 0.05232f
C6316 a_n8964_8799.t132 gnd 0.601897f
C6317 a_n8964_8799.n76 gnd 0.268658f
C6318 a_n8964_8799.t134 gnd 0.601897f
C6319 a_n8964_8799.n77 gnd 0.05232f
C6320 a_n8964_8799.n78 gnd 0.011873f
C6321 a_n8964_8799.t72 gnd 0.601897f
C6322 a_n8964_8799.n79 gnd 0.05232f
C6323 a_n8964_8799.t75 gnd 0.601897f
C6324 a_n8964_8799.n80 gnd 0.263819f
C6325 a_n8964_8799.t108 gnd 0.601897f
C6326 a_n8964_8799.n81 gnd 0.05232f
C6327 a_n8964_8799.t114 gnd 0.601897f
C6328 a_n8964_8799.n82 gnd 0.268012f
C6329 a_n8964_8799.t87 gnd 0.613289f
C6330 a_n8964_8799.n83 gnd 0.252342f
C6331 a_n8964_8799.n84 gnd 0.171077f
C6332 a_n8964_8799.n85 gnd 0.011873f
C6333 a_n8964_8799.t52 gnd 0.601897f
C6334 a_n8964_8799.n86 gnd 0.268819f
C6335 a_n8964_8799.n87 gnd 0.011873f
C6336 a_n8964_8799.n88 gnd 0.05232f
C6337 a_n8964_8799.n89 gnd 0.05232f
C6338 a_n8964_8799.n90 gnd 0.05232f
C6339 a_n8964_8799.n91 gnd 0.268335f
C6340 a_n8964_8799.n92 gnd 0.011873f
C6341 a_n8964_8799.t135 gnd 0.601897f
C6342 a_n8964_8799.n93 gnd 0.268819f
C6343 a_n8964_8799.n94 gnd 0.05232f
C6344 a_n8964_8799.n95 gnd 0.05232f
C6345 a_n8964_8799.n96 gnd 0.05232f
C6346 a_n8964_8799.n97 gnd 0.263496f
C6347 a_n8964_8799.t105 gnd 0.601897f
C6348 a_n8964_8799.n98 gnd 0.268658f
C6349 a_n8964_8799.n99 gnd 0.011873f
C6350 a_n8964_8799.n100 gnd 0.05232f
C6351 a_n8964_8799.n101 gnd 0.05232f
C6352 a_n8964_8799.n102 gnd 0.05232f
C6353 a_n8964_8799.n103 gnd 0.263496f
C6354 a_n8964_8799.n104 gnd 0.011873f
C6355 a_n8964_8799.t91 gnd 0.601897f
C6356 a_n8964_8799.n105 gnd 0.268819f
C6357 a_n8964_8799.n106 gnd 0.05232f
C6358 a_n8964_8799.n107 gnd 0.05232f
C6359 a_n8964_8799.n108 gnd 0.05232f
C6360 a_n8964_8799.n109 gnd 0.268335f
C6361 a_n8964_8799.t131 gnd 0.601897f
C6362 a_n8964_8799.n110 gnd 0.263819f
C6363 a_n8964_8799.n111 gnd 0.011873f
C6364 a_n8964_8799.n112 gnd 0.05232f
C6365 a_n8964_8799.n113 gnd 0.05232f
C6366 a_n8964_8799.n114 gnd 0.05232f
C6367 a_n8964_8799.n115 gnd 0.011873f
C6368 a_n8964_8799.t88 gnd 0.601897f
C6369 a_n8964_8799.n116 gnd 0.268012f
C6370 a_n8964_8799.t115 gnd 0.601897f
C6371 a_n8964_8799.n117 gnd 0.263335f
C6372 a_n8964_8799.n118 gnd 0.135549f
C6373 a_n8964_8799.n119 gnd 0.906524f
C6374 a_n8964_8799.n120 gnd 0.05232f
C6375 a_n8964_8799.t58 gnd 0.601897f
C6376 a_n8964_8799.n121 gnd 0.268819f
C6377 a_n8964_8799.n122 gnd 0.05232f
C6378 a_n8964_8799.n123 gnd 0.011873f
C6379 a_n8964_8799.t73 gnd 0.601897f
C6380 a_n8964_8799.n124 gnd 0.05232f
C6381 a_n8964_8799.t101 gnd 0.601897f
C6382 a_n8964_8799.n125 gnd 0.268658f
C6383 a_n8964_8799.t85 gnd 0.601897f
C6384 a_n8964_8799.n126 gnd 0.05232f
C6385 a_n8964_8799.n127 gnd 0.011873f
C6386 a_n8964_8799.t89 gnd 0.601897f
C6387 a_n8964_8799.n128 gnd 0.05232f
C6388 a_n8964_8799.t56 gnd 0.601897f
C6389 a_n8964_8799.n129 gnd 0.263819f
C6390 a_n8964_8799.t110 gnd 0.601897f
C6391 a_n8964_8799.n130 gnd 0.05232f
C6392 a_n8964_8799.t43 gnd 0.601897f
C6393 a_n8964_8799.n131 gnd 0.268012f
C6394 a_n8964_8799.t81 gnd 0.613289f
C6395 a_n8964_8799.n132 gnd 0.252342f
C6396 a_n8964_8799.n133 gnd 0.171077f
C6397 a_n8964_8799.n134 gnd 0.011873f
C6398 a_n8964_8799.t96 gnd 0.601897f
C6399 a_n8964_8799.n135 gnd 0.268819f
C6400 a_n8964_8799.n136 gnd 0.011873f
C6401 a_n8964_8799.n137 gnd 0.05232f
C6402 a_n8964_8799.n138 gnd 0.05232f
C6403 a_n8964_8799.n139 gnd 0.05232f
C6404 a_n8964_8799.n140 gnd 0.268335f
C6405 a_n8964_8799.n141 gnd 0.011873f
C6406 a_n8964_8799.t68 gnd 0.601897f
C6407 a_n8964_8799.n142 gnd 0.268819f
C6408 a_n8964_8799.n143 gnd 0.05232f
C6409 a_n8964_8799.n144 gnd 0.05232f
C6410 a_n8964_8799.n145 gnd 0.05232f
C6411 a_n8964_8799.n146 gnd 0.263496f
C6412 a_n8964_8799.t50 gnd 0.601897f
C6413 a_n8964_8799.n147 gnd 0.268658f
C6414 a_n8964_8799.n148 gnd 0.011873f
C6415 a_n8964_8799.n149 gnd 0.05232f
C6416 a_n8964_8799.n150 gnd 0.05232f
C6417 a_n8964_8799.n151 gnd 0.05232f
C6418 a_n8964_8799.n152 gnd 0.263496f
C6419 a_n8964_8799.n153 gnd 0.011873f
C6420 a_n8964_8799.t117 gnd 0.601897f
C6421 a_n8964_8799.n154 gnd 0.268819f
C6422 a_n8964_8799.n155 gnd 0.05232f
C6423 a_n8964_8799.n156 gnd 0.05232f
C6424 a_n8964_8799.n157 gnd 0.05232f
C6425 a_n8964_8799.n158 gnd 0.268335f
C6426 a_n8964_8799.t124 gnd 0.601897f
C6427 a_n8964_8799.n159 gnd 0.263819f
C6428 a_n8964_8799.n160 gnd 0.011873f
C6429 a_n8964_8799.n161 gnd 0.05232f
C6430 a_n8964_8799.n162 gnd 0.05232f
C6431 a_n8964_8799.n163 gnd 0.05232f
C6432 a_n8964_8799.n164 gnd 0.011873f
C6433 a_n8964_8799.t40 gnd 0.601897f
C6434 a_n8964_8799.n165 gnd 0.268012f
C6435 a_n8964_8799.t92 gnd 0.601897f
C6436 a_n8964_8799.n166 gnd 0.263335f
C6437 a_n8964_8799.n167 gnd 0.135549f
C6438 a_n8964_8799.n168 gnd 1.82134f
C6439 a_n8964_8799.n169 gnd 0.05232f
C6440 a_n8964_8799.t47 gnd 0.601897f
C6441 a_n8964_8799.t45 gnd 0.601897f
C6442 a_n8964_8799.t113 gnd 0.601897f
C6443 a_n8964_8799.n170 gnd 0.268819f
C6444 a_n8964_8799.n171 gnd 0.05232f
C6445 a_n8964_8799.t61 gnd 0.601897f
C6446 a_n8964_8799.t49 gnd 0.601897f
C6447 a_n8964_8799.n172 gnd 0.05232f
C6448 a_n8964_8799.t119 gnd 0.601897f
C6449 a_n8964_8799.n173 gnd 0.268819f
C6450 a_n8964_8799.n174 gnd 0.05232f
C6451 a_n8964_8799.t82 gnd 0.601897f
C6452 a_n8964_8799.t62 gnd 0.601897f
C6453 a_n8964_8799.n175 gnd 0.05232f
C6454 a_n8964_8799.t133 gnd 0.601897f
C6455 a_n8964_8799.n176 gnd 0.268658f
C6456 a_n8964_8799.n177 gnd 0.05232f
C6457 a_n8964_8799.t98 gnd 0.601897f
C6458 a_n8964_8799.t64 gnd 0.601897f
C6459 a_n8964_8799.n178 gnd 0.05232f
C6460 a_n8964_8799.t129 gnd 0.601897f
C6461 a_n8964_8799.n179 gnd 0.268335f
C6462 a_n8964_8799.n180 gnd 0.05232f
C6463 a_n8964_8799.t100 gnd 0.601897f
C6464 a_n8964_8799.t76 gnd 0.601897f
C6465 a_n8964_8799.n181 gnd 0.05232f
C6466 a_n8964_8799.t46 gnd 0.601897f
C6467 a_n8964_8799.n182 gnd 0.268012f
C6468 a_n8964_8799.t116 gnd 0.613289f
C6469 a_n8964_8799.n183 gnd 0.252342f
C6470 a_n8964_8799.n184 gnd 0.171077f
C6471 a_n8964_8799.n185 gnd 0.011873f
C6472 a_n8964_8799.n186 gnd 0.268819f
C6473 a_n8964_8799.n187 gnd 0.011873f
C6474 a_n8964_8799.n188 gnd 0.263819f
C6475 a_n8964_8799.n189 gnd 0.05232f
C6476 a_n8964_8799.n190 gnd 0.05232f
C6477 a_n8964_8799.n191 gnd 0.05232f
C6478 a_n8964_8799.n192 gnd 0.011873f
C6479 a_n8964_8799.n193 gnd 0.268819f
C6480 a_n8964_8799.n194 gnd 0.011873f
C6481 a_n8964_8799.n195 gnd 0.263496f
C6482 a_n8964_8799.n196 gnd 0.05232f
C6483 a_n8964_8799.n197 gnd 0.05232f
C6484 a_n8964_8799.n198 gnd 0.05232f
C6485 a_n8964_8799.n199 gnd 0.011873f
C6486 a_n8964_8799.n200 gnd 0.268658f
C6487 a_n8964_8799.n201 gnd 0.263496f
C6488 a_n8964_8799.n202 gnd 0.011873f
C6489 a_n8964_8799.n203 gnd 0.05232f
C6490 a_n8964_8799.n204 gnd 0.05232f
C6491 a_n8964_8799.n205 gnd 0.05232f
C6492 a_n8964_8799.n206 gnd 0.011873f
C6493 a_n8964_8799.n207 gnd 0.268335f
C6494 a_n8964_8799.n208 gnd 0.263819f
C6495 a_n8964_8799.n209 gnd 0.011873f
C6496 a_n8964_8799.n210 gnd 0.05232f
C6497 a_n8964_8799.n211 gnd 0.05232f
C6498 a_n8964_8799.n212 gnd 0.05232f
C6499 a_n8964_8799.n213 gnd 0.011873f
C6500 a_n8964_8799.n214 gnd 0.268012f
C6501 a_n8964_8799.n215 gnd 0.263335f
C6502 a_n8964_8799.n216 gnd 0.301459f
C6503 a_n8964_8799.n217 gnd 0.05232f
C6504 a_n8964_8799.t55 gnd 0.601897f
C6505 a_n8964_8799.t53 gnd 0.601897f
C6506 a_n8964_8799.t127 gnd 0.601897f
C6507 a_n8964_8799.n218 gnd 0.268819f
C6508 a_n8964_8799.n219 gnd 0.05232f
C6509 a_n8964_8799.t67 gnd 0.601897f
C6510 a_n8964_8799.t60 gnd 0.601897f
C6511 a_n8964_8799.n220 gnd 0.05232f
C6512 a_n8964_8799.t130 gnd 0.601897f
C6513 a_n8964_8799.n221 gnd 0.268819f
C6514 a_n8964_8799.n222 gnd 0.05232f
C6515 a_n8964_8799.t94 gnd 0.601897f
C6516 a_n8964_8799.t70 gnd 0.601897f
C6517 a_n8964_8799.n223 gnd 0.05232f
C6518 a_n8964_8799.t48 gnd 0.601897f
C6519 a_n8964_8799.n224 gnd 0.268658f
C6520 a_n8964_8799.n225 gnd 0.05232f
C6521 a_n8964_8799.t107 gnd 0.601897f
C6522 a_n8964_8799.t71 gnd 0.601897f
C6523 a_n8964_8799.n226 gnd 0.05232f
C6524 a_n8964_8799.t41 gnd 0.601897f
C6525 a_n8964_8799.n227 gnd 0.268335f
C6526 a_n8964_8799.n228 gnd 0.05232f
C6527 a_n8964_8799.t112 gnd 0.601897f
C6528 a_n8964_8799.t84 gnd 0.601897f
C6529 a_n8964_8799.n229 gnd 0.05232f
C6530 a_n8964_8799.t54 gnd 0.601897f
C6531 a_n8964_8799.n230 gnd 0.268012f
C6532 a_n8964_8799.t128 gnd 0.613289f
C6533 a_n8964_8799.n231 gnd 0.252342f
C6534 a_n8964_8799.n232 gnd 0.171077f
C6535 a_n8964_8799.n233 gnd 0.011873f
C6536 a_n8964_8799.n234 gnd 0.268819f
C6537 a_n8964_8799.n235 gnd 0.011873f
C6538 a_n8964_8799.n236 gnd 0.263819f
C6539 a_n8964_8799.n237 gnd 0.05232f
C6540 a_n8964_8799.n238 gnd 0.05232f
C6541 a_n8964_8799.n239 gnd 0.05232f
C6542 a_n8964_8799.n240 gnd 0.011873f
C6543 a_n8964_8799.n241 gnd 0.268819f
C6544 a_n8964_8799.n242 gnd 0.011873f
C6545 a_n8964_8799.n243 gnd 0.263496f
C6546 a_n8964_8799.n244 gnd 0.05232f
C6547 a_n8964_8799.n245 gnd 0.05232f
C6548 a_n8964_8799.n246 gnd 0.05232f
C6549 a_n8964_8799.n247 gnd 0.011873f
C6550 a_n8964_8799.n248 gnd 0.268658f
C6551 a_n8964_8799.n249 gnd 0.263496f
C6552 a_n8964_8799.n250 gnd 0.011873f
C6553 a_n8964_8799.n251 gnd 0.05232f
C6554 a_n8964_8799.n252 gnd 0.05232f
C6555 a_n8964_8799.n253 gnd 0.05232f
C6556 a_n8964_8799.n254 gnd 0.011873f
C6557 a_n8964_8799.n255 gnd 0.268335f
C6558 a_n8964_8799.n256 gnd 0.263819f
C6559 a_n8964_8799.n257 gnd 0.011873f
C6560 a_n8964_8799.n258 gnd 0.05232f
C6561 a_n8964_8799.n259 gnd 0.05232f
C6562 a_n8964_8799.n260 gnd 0.05232f
C6563 a_n8964_8799.n261 gnd 0.011873f
C6564 a_n8964_8799.n262 gnd 0.268012f
C6565 a_n8964_8799.n263 gnd 0.263335f
C6566 a_n8964_8799.n264 gnd 0.135549f
C6567 a_n8964_8799.n265 gnd 0.906524f
C6568 a_n8964_8799.n266 gnd 0.05232f
C6569 a_n8964_8799.t93 gnd 0.601897f
C6570 a_n8964_8799.t111 gnd 0.601897f
C6571 a_n8964_8799.t59 gnd 0.601897f
C6572 a_n8964_8799.n267 gnd 0.268819f
C6573 a_n8964_8799.n268 gnd 0.05232f
C6574 a_n8964_8799.t125 gnd 0.601897f
C6575 a_n8964_8799.t74 gnd 0.601897f
C6576 a_n8964_8799.n269 gnd 0.05232f
C6577 a_n8964_8799.t120 gnd 0.601897f
C6578 a_n8964_8799.n270 gnd 0.268819f
C6579 a_n8964_8799.n271 gnd 0.05232f
C6580 a_n8964_8799.t63 gnd 0.601897f
C6581 a_n8964_8799.t102 gnd 0.601897f
C6582 a_n8964_8799.n272 gnd 0.05232f
C6583 a_n8964_8799.t51 gnd 0.601897f
C6584 a_n8964_8799.n273 gnd 0.268658f
C6585 a_n8964_8799.n274 gnd 0.05232f
C6586 a_n8964_8799.t90 gnd 0.601897f
C6587 a_n8964_8799.t69 gnd 0.601897f
C6588 a_n8964_8799.n275 gnd 0.05232f
C6589 a_n8964_8799.t109 gnd 0.601897f
C6590 a_n8964_8799.n276 gnd 0.268335f
C6591 a_n8964_8799.n277 gnd 0.05232f
C6592 a_n8964_8799.t57 gnd 0.601897f
C6593 a_n8964_8799.t97 gnd 0.601897f
C6594 a_n8964_8799.n278 gnd 0.05232f
C6595 a_n8964_8799.t44 gnd 0.601897f
C6596 a_n8964_8799.n279 gnd 0.268012f
C6597 a_n8964_8799.t83 gnd 0.613289f
C6598 a_n8964_8799.n280 gnd 0.252342f
C6599 a_n8964_8799.n281 gnd 0.171077f
C6600 a_n8964_8799.n282 gnd 0.011873f
C6601 a_n8964_8799.n283 gnd 0.268819f
C6602 a_n8964_8799.n284 gnd 0.011873f
C6603 a_n8964_8799.n285 gnd 0.263819f
C6604 a_n8964_8799.n286 gnd 0.05232f
C6605 a_n8964_8799.n287 gnd 0.05232f
C6606 a_n8964_8799.n288 gnd 0.05232f
C6607 a_n8964_8799.n289 gnd 0.011873f
C6608 a_n8964_8799.n290 gnd 0.268819f
C6609 a_n8964_8799.n291 gnd 0.011873f
C6610 a_n8964_8799.n292 gnd 0.263496f
C6611 a_n8964_8799.n293 gnd 0.05232f
C6612 a_n8964_8799.n294 gnd 0.05232f
C6613 a_n8964_8799.n295 gnd 0.05232f
C6614 a_n8964_8799.n296 gnd 0.011873f
C6615 a_n8964_8799.n297 gnd 0.268658f
C6616 a_n8964_8799.n298 gnd 0.263496f
C6617 a_n8964_8799.n299 gnd 0.011873f
C6618 a_n8964_8799.n300 gnd 0.05232f
C6619 a_n8964_8799.n301 gnd 0.05232f
C6620 a_n8964_8799.n302 gnd 0.05232f
C6621 a_n8964_8799.n303 gnd 0.011873f
C6622 a_n8964_8799.n304 gnd 0.268335f
C6623 a_n8964_8799.n305 gnd 0.263819f
C6624 a_n8964_8799.n306 gnd 0.011873f
C6625 a_n8964_8799.n307 gnd 0.05232f
C6626 a_n8964_8799.n308 gnd 0.05232f
C6627 a_n8964_8799.n309 gnd 0.05232f
C6628 a_n8964_8799.n310 gnd 0.011873f
C6629 a_n8964_8799.n311 gnd 0.268012f
C6630 a_n8964_8799.n312 gnd 0.263335f
C6631 a_n8964_8799.n313 gnd 0.135549f
C6632 a_n8964_8799.n314 gnd 1.45602f
C6633 a_n8964_8799.n315 gnd 17.5023f
C6634 a_n8964_8799.n316 gnd 4.40501f
C6635 a_n8964_8799.t27 gnd 0.112902f
C6636 a_n8964_8799.t28 gnd 0.112902f
C6637 a_n8964_8799.n317 gnd 0.999856f
C6638 a_n8964_8799.t23 gnd 0.112902f
C6639 a_n8964_8799.t24 gnd 0.112902f
C6640 a_n8964_8799.n318 gnd 0.997638f
C6641 a_n8964_8799.n319 gnd 0.736268f
C6642 a_n8964_8799.n320 gnd 0.473739f
C6643 a_n8964_8799.t22 gnd 0.112902f
C6644 a_n8964_8799.t34 gnd 0.112902f
C6645 a_n8964_8799.n321 gnd 0.997638f
C6646 a_n8964_8799.n322 gnd 0.331824f
C6647 a_n8964_8799.t35 gnd 0.112902f
C6648 a_n8964_8799.t31 gnd 0.112902f
C6649 a_n8964_8799.n323 gnd 0.997638f
C6650 a_n8964_8799.n324 gnd 2.587f
C6651 a_n8964_8799.t32 gnd 0.112902f
C6652 a_n8964_8799.t30 gnd 0.112902f
C6653 a_n8964_8799.n325 gnd 0.999855f
C6654 a_n8964_8799.t25 gnd 0.112902f
C6655 a_n8964_8799.t29 gnd 0.112902f
C6656 a_n8964_8799.n326 gnd 0.997637f
C6657 a_n8964_8799.n327 gnd 0.73627f
C6658 a_n8964_8799.n328 gnd 2.00302f
C6659 a_n8964_8799.t36 gnd 0.112902f
C6660 a_n8964_8799.t26 gnd 0.112902f
C6661 a_n8964_8799.n329 gnd 0.997637f
C6662 a_n8964_8799.n330 gnd 0.736272f
C6663 a_n8964_8799.n331 gnd 0.999853f
C6664 a_n8964_8799.t37 gnd 0.112902f
C6665 a_n2903_n3924.n0 gnd 1.85226f
C6666 a_n2903_n3924.n1 gnd 1.55666f
C6667 a_n2903_n3924.n2 gnd 1.22094f
C6668 a_n2903_n3924.n3 gnd 1.34544f
C6669 a_n2903_n3924.n4 gnd 1.97724f
C6670 a_n2903_n3924.n5 gnd 1.64424f
C6671 a_n2903_n3924.n6 gnd 0.82212f
C6672 a_n2903_n3924.n7 gnd 2.30935f
C6673 a_n2903_n3924.n8 gnd 1.00973f
C6674 a_n2903_n3924.n9 gnd 1.18081f
C6675 a_n2903_n3924.t1 gnd 0.090392f
C6676 a_n2903_n3924.t13 gnd 0.090392f
C6677 a_n2903_n3924.t3 gnd 0.090392f
C6678 a_n2903_n3924.n10 gnd 0.738247f
C6679 a_n2903_n3924.t18 gnd 1.16889f
C6680 a_n2903_n3924.t10 gnd 0.090392f
C6681 a_n2903_n3924.t38 gnd 0.090392f
C6682 a_n2903_n3924.n11 gnd 0.738247f
C6683 a_n2903_n3924.t16 gnd 0.939461f
C6684 a_n2903_n3924.t14 gnd 1.16892f
C6685 a_n2903_n3924.t9 gnd 1.16726f
C6686 a_n2903_n3924.t11 gnd 1.16726f
C6687 a_n2903_n3924.t20 gnd 1.16726f
C6688 a_n2903_n3924.t6 gnd 1.16726f
C6689 a_n2903_n3924.t4 gnd 1.16726f
C6690 a_n2903_n3924.t21 gnd 1.16726f
C6691 a_n2903_n3924.n12 gnd 0.847907f
C6692 a_n2903_n3924.t24 gnd 0.939457f
C6693 a_n2903_n3924.t35 gnd 0.090392f
C6694 a_n2903_n3924.t31 gnd 0.090392f
C6695 a_n2903_n3924.n13 gnd 0.738246f
C6696 a_n2903_n3924.t32 gnd 0.090392f
C6697 a_n2903_n3924.t29 gnd 0.090392f
C6698 a_n2903_n3924.n14 gnd 0.738246f
C6699 a_n2903_n3924.t23 gnd 0.090392f
C6700 a_n2903_n3924.t37 gnd 0.090392f
C6701 a_n2903_n3924.n15 gnd 0.738246f
C6702 a_n2903_n3924.t36 gnd 0.939457f
C6703 a_n2903_n3924.t7 gnd 0.939457f
C6704 a_n2903_n3924.t39 gnd 0.090392f
C6705 a_n2903_n3924.t5 gnd 0.090392f
C6706 a_n2903_n3924.n16 gnd 0.738246f
C6707 a_n2903_n3924.t15 gnd 0.090392f
C6708 a_n2903_n3924.t19 gnd 0.090392f
C6709 a_n2903_n3924.n17 gnd 0.738246f
C6710 a_n2903_n3924.t17 gnd 0.090392f
C6711 a_n2903_n3924.t8 gnd 0.090392f
C6712 a_n2903_n3924.n18 gnd 0.738246f
C6713 a_n2903_n3924.t12 gnd 0.939457f
C6714 a_n2903_n3924.n19 gnd 0.847907f
C6715 a_n2903_n3924.t22 gnd 0.939457f
C6716 a_n2903_n3924.t27 gnd 0.090392f
C6717 a_n2903_n3924.t26 gnd 0.090392f
C6718 a_n2903_n3924.n20 gnd 0.738247f
C6719 a_n2903_n3924.t25 gnd 0.090392f
C6720 a_n2903_n3924.t33 gnd 0.090392f
C6721 a_n2903_n3924.n21 gnd 0.738247f
C6722 a_n2903_n3924.t30 gnd 0.090392f
C6723 a_n2903_n3924.t34 gnd 0.090392f
C6724 a_n2903_n3924.n22 gnd 0.738247f
C6725 a_n2903_n3924.t28 gnd 0.939461f
C6726 a_n2903_n3924.t2 gnd 0.939461f
C6727 a_n2903_n3924.n23 gnd 0.738248f
C6728 a_n2903_n3924.t0 gnd 0.090392f
C6729 plus.n0 gnd 0.021868f
C6730 plus.t9 gnd 0.309306f
C6731 plus.n1 gnd 0.021868f
C6732 plus.t5 gnd 0.309306f
C6733 plus.t6 gnd 0.309306f
C6734 plus.n2 gnd 0.137403f
C6735 plus.n3 gnd 0.021868f
C6736 plus.t16 gnd 0.309306f
C6737 plus.t17 gnd 0.309306f
C6738 plus.n4 gnd 0.137403f
C6739 plus.n5 gnd 0.021868f
C6740 plus.t13 gnd 0.309306f
C6741 plus.t10 gnd 0.309306f
C6742 plus.n6 gnd 0.140399f
C6743 plus.t12 gnd 0.31973f
C6744 plus.n7 gnd 0.128799f
C6745 plus.n8 gnd 0.092541f
C6746 plus.n9 gnd 0.004962f
C6747 plus.n10 gnd 0.137403f
C6748 plus.n11 gnd 0.004962f
C6749 plus.n12 gnd 0.021868f
C6750 plus.n13 gnd 0.021868f
C6751 plus.n14 gnd 0.021868f
C6752 plus.n15 gnd 0.004962f
C6753 plus.n16 gnd 0.137403f
C6754 plus.n17 gnd 0.004962f
C6755 plus.n18 gnd 0.021868f
C6756 plus.n19 gnd 0.021868f
C6757 plus.n20 gnd 0.021868f
C6758 plus.n21 gnd 0.004962f
C6759 plus.n22 gnd 0.137403f
C6760 plus.n23 gnd 0.004962f
C6761 plus.n24 gnd 0.136797f
C6762 plus.n25 gnd 0.24645f
C6763 plus.n26 gnd 0.021868f
C6764 plus.n27 gnd 0.004962f
C6765 plus.t7 gnd 0.309306f
C6766 plus.n28 gnd 0.021868f
C6767 plus.n29 gnd 0.004962f
C6768 plus.t20 gnd 0.309306f
C6769 plus.n30 gnd 0.021868f
C6770 plus.n31 gnd 0.004962f
C6771 plus.t19 gnd 0.309306f
C6772 plus.t15 gnd 0.31973f
C6773 plus.t14 gnd 0.309306f
C6774 plus.n32 gnd 0.140399f
C6775 plus.n33 gnd 0.128799f
C6776 plus.n34 gnd 0.092541f
C6777 plus.n35 gnd 0.021868f
C6778 plus.n36 gnd 0.137403f
C6779 plus.n37 gnd 0.004962f
C6780 plus.t18 gnd 0.309306f
C6781 plus.n38 gnd 0.137403f
C6782 plus.n39 gnd 0.021868f
C6783 plus.n40 gnd 0.021868f
C6784 plus.n41 gnd 0.021868f
C6785 plus.n42 gnd 0.137403f
C6786 plus.n43 gnd 0.004962f
C6787 plus.t8 gnd 0.309306f
C6788 plus.n44 gnd 0.137403f
C6789 plus.n45 gnd 0.021868f
C6790 plus.n46 gnd 0.021868f
C6791 plus.n47 gnd 0.021868f
C6792 plus.n48 gnd 0.137403f
C6793 plus.n49 gnd 0.004962f
C6794 plus.t11 gnd 0.309306f
C6795 plus.n50 gnd 0.136797f
C6796 plus.n51 gnd 0.625951f
C6797 plus.n52 gnd 0.956547f
C6798 plus.t4 gnd 0.037751f
C6799 plus.t2 gnd 0.006741f
C6800 plus.t3 gnd 0.006741f
C6801 plus.n53 gnd 0.021863f
C6802 plus.n54 gnd 0.169727f
C6803 plus.t1 gnd 0.006741f
C6804 plus.t0 gnd 0.006741f
C6805 plus.n55 gnd 0.021863f
C6806 plus.n56 gnd 0.127401f
C6807 plus.n57 gnd 2.6083f
.ends

